/*

c5315:
	jxor: 109
	jspl: 308
	jspl3: 385
	jnot: 226
	jdff: 4692
	jand: 605
	jor: 419

Summary:
	jxor: 109
	jspl: 308
	jspl3: 385
	jnot: 226
	jdff: 4692
	jand: 605
	jor: 419
*/

module c5315(gclk, G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37, G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79, G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106, G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G140, G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170, G173, G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206, G209, G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248, G251, G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292, G293, G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335, G338, G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386, G389, G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514, G523, G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691, G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717, G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115, G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843, G882, G767, G807, G658, G690);
	input gclk;
	input G1;
	input G4;
	input G11;
	input G14;
	input G17;
	input G20;
	input G23;
	input G24;
	input G25;
	input G26;
	input G27;
	input G31;
	input G34;
	input G37;
	input G40;
	input G43;
	input G46;
	input G49;
	input G52;
	input G53;
	input G54;
	input G61;
	input G64;
	input G67;
	input G70;
	input G73;
	input G76;
	input G79;
	input G80;
	input G81;
	input G82;
	input G83;
	input G86;
	input G87;
	input G88;
	input G91;
	input G94;
	input G97;
	input G100;
	input G103;
	input G106;
	input G109;
	input G112;
	input G113;
	input G114;
	input G115;
	input G116;
	input G117;
	input G118;
	input G119;
	input G120;
	input G121;
	input G122;
	input G123;
	input G126;
	input G127;
	input G128;
	input G129;
	input G130;
	input G131;
	input G132;
	input G135;
	input G136;
	input G137;
	input G140;
	input G141;
	input G145;
	input G146;
	input G149;
	input G152;
	input G155;
	input G158;
	input G161;
	input G164;
	input G167;
	input G170;
	input G173;
	input G176;
	input G179;
	input G182;
	input G185;
	input G188;
	input G191;
	input G194;
	input G197;
	input G200;
	input G203;
	input G206;
	input G209;
	input G210;
	input G217;
	input G218;
	input G225;
	input G226;
	input G233;
	input G234;
	input G241;
	input G242;
	input G245;
	input G248;
	input G251;
	input G254;
	input G257;
	input G264;
	input G265;
	input G272;
	input G273;
	input G280;
	input G281;
	input G288;
	input G289;
	input G292;
	input G293;
	input G299;
	input G302;
	input G307;
	input G308;
	input G315;
	input G316;
	input G323;
	input G324;
	input G331;
	input G332;
	input G335;
	input G338;
	input G341;
	input G348;
	input G351;
	input G358;
	input G361;
	input G366;
	input G369;
	input G372;
	input G373;
	input G374;
	input G386;
	input G389;
	input G400;
	input G411;
	input G422;
	input G435;
	input G446;
	input G457;
	input G468;
	input G479;
	input G490;
	input G503;
	input G514;
	input G523;
	input G534;
	input G545;
	input G549;
	input G552;
	input G556;
	input G559;
	input G562;
	input G1497;
	input G1689;
	input G1690;
	input G1691;
	input G1694;
	input G2174;
	input G2358;
	input G2824;
	input G3173;
	input G3546;
	input G3548;
	input G3550;
	input G3552;
	input G3717;
	input G3724;
	input G4087;
	input G4088;
	input G4089;
	input G4090;
	input G4091;
	input G4092;
	input G4115;
	output G144;
	output G298;
	output G973;
	output G594;
	output G599;
	output G600;
	output G601;
	output G602;
	output G603;
	output G604;
	output G611;
	output G612;
	output G810;
	output G848;
	output G849;
	output G850;
	output G851;
	output G634;
	output G815;
	output G845;
	output G847;
	output G926;
	output G923;
	output G921;
	output G892;
	output G887;
	output G606;
	output G656;
	output G809;
	output G993;
	output G978;
	output G949;
	output G939;
	output G889;
	output G593;
	output G636;
	output G704;
	output G717;
	output G820;
	output G639;
	output G673;
	output G707;
	output G715;
	output G598;
	output G610;
	output G588;
	output G615;
	output G626;
	output G632;
	output G1002;
	output G1004;
	output G591;
	output G618;
	output G621;
	output G629;
	output G822;
	output G838;
	output G861;
	output G623;
	output G722;
	output G832;
	output G834;
	output G836;
	output G859;
	output G871;
	output G873;
	output G875;
	output G877;
	output G998;
	output G1000;
	output G575;
	output G585;
	output G661;
	output G693;
	output G747;
	output G752;
	output G757;
	output G762;
	output G787;
	output G792;
	output G797;
	output G802;
	output G642;
	output G664;
	output G667;
	output G670;
	output G676;
	output G696;
	output G699;
	output G702;
	output G818;
	output G813;
	output G824;
	output G826;
	output G828;
	output G830;
	output G854;
	output G863;
	output G865;
	output G867;
	output G869;
	output G712;
	output G727;
	output G732;
	output G737;
	output G742;
	output G772;
	output G777;
	output G782;
	output G645;
	output G648;
	output G651;
	output G654;
	output G679;
	output G682;
	output G685;
	output G688;
	output G843;
	output G882;
	output G767;
	output G807;
	output G658;
	output G690;
	wire n314;
	wire n316;
	wire n318;
	wire n320;
	wire n321;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n338;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1157;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire[2:0] w_G1_0;
	wire[2:0] w_G1_1;
	wire[1:0] w_G1_2;
	wire[2:0] w_G4_0;
	wire[1:0] w_G4_1;
	wire[1:0] w_G11_0;
	wire[1:0] w_G14_0;
	wire[1:0] w_G17_0;
	wire[1:0] w_G20_0;
	wire[1:0] w_G37_0;
	wire[1:0] w_G40_0;
	wire[1:0] w_G43_0;
	wire[1:0] w_G46_0;
	wire[1:0] w_G49_0;
	wire[1:0] w_G54_0;
	wire[1:0] w_G61_0;
	wire[1:0] w_G64_0;
	wire[1:0] w_G67_0;
	wire[1:0] w_G70_0;
	wire[1:0] w_G73_0;
	wire[1:0] w_G76_0;
	wire[1:0] w_G91_0;
	wire[1:0] w_G100_0;
	wire[1:0] w_G103_0;
	wire[1:0] w_G106_0;
	wire[1:0] w_G109_0;
	wire[1:0] w_G123_0;
	wire[1:0] w_G132_0;
	wire[2:0] w_G137_0;
	wire[2:0] w_G137_1;
	wire[2:0] w_G137_2;
	wire[2:0] w_G137_3;
	wire[2:0] w_G137_4;
	wire[2:0] w_G137_5;
	wire[2:0] w_G137_6;
	wire[2:0] w_G137_7;
	wire[2:0] w_G137_8;
	wire[1:0] w_G137_9;
	wire[2:0] w_G141_0;
	wire[2:0] w_G141_1;
	wire[2:0] w_G141_2;
	wire[1:0] w_G146_0;
	wire[1:0] w_G149_0;
	wire[1:0] w_G152_0;
	wire[1:0] w_G155_0;
	wire[1:0] w_G158_0;
	wire[1:0] w_G161_0;
	wire[1:0] w_G164_0;
	wire[1:0] w_G167_0;
	wire[1:0] w_G170_0;
	wire[1:0] w_G173_0;
	wire[1:0] w_G182_0;
	wire[1:0] w_G185_0;
	wire[1:0] w_G188_0;
	wire[1:0] w_G191_0;
	wire[1:0] w_G194_0;
	wire[1:0] w_G197_0;
	wire[1:0] w_G200_0;
	wire[1:0] w_G203_0;
	wire[2:0] w_G206_0;
	wire[2:0] w_G210_0;
	wire[2:0] w_G210_1;
	wire[2:0] w_G210_2;
	wire[2:0] w_G218_0;
	wire[2:0] w_G218_1;
	wire[2:0] w_G218_2;
	wire[2:0] w_G226_0;
	wire[2:0] w_G226_1;
	wire[2:0] w_G226_2;
	wire[2:0] w_G234_0;
	wire[2:0] w_G234_1;
	wire[1:0] w_G234_2;
	wire[2:0] w_G242_0;
	wire[2:0] w_G242_1;
	wire[1:0] w_G245_0;
	wire[2:0] w_G248_0;
	wire[2:0] w_G248_1;
	wire[2:0] w_G248_2;
	wire[2:0] w_G248_3;
	wire[2:0] w_G248_4;
	wire[1:0] w_G248_5;
	wire[2:0] w_G251_0;
	wire[2:0] w_G251_1;
	wire[2:0] w_G251_2;
	wire[2:0] w_G251_3;
	wire[2:0] w_G251_4;
	wire[2:0] w_G254_0;
	wire[2:0] w_G254_1;
	wire[2:0] w_G257_0;
	wire[2:0] w_G257_1;
	wire[2:0] w_G257_2;
	wire[2:0] w_G265_0;
	wire[2:0] w_G265_1;
	wire[1:0] w_G265_2;
	wire[2:0] w_G273_0;
	wire[2:0] w_G273_1;
	wire[2:0] w_G273_2;
	wire[1:0] w_G280_0;
	wire[2:0] w_G281_0;
	wire[2:0] w_G281_1;
	wire[1:0] w_G281_2;
	wire[1:0] w_G289_0;
	wire[2:0] w_G293_0;
	wire[2:0] w_G299_0;
	wire[2:0] w_G302_0;
	wire[2:0] w_G308_0;
	wire[2:0] w_G308_1;
	wire[2:0] w_G316_0;
	wire[2:0] w_G316_1;
	wire[2:0] w_G324_0;
	wire[2:0] w_G324_1;
	wire[1:0] w_G331_0;
	wire[2:0] w_G332_0;
	wire[2:0] w_G332_1;
	wire[2:0] w_G332_2;
	wire[2:0] w_G332_3;
	wire[2:0] w_G332_4;
	wire[2:0] w_G335_0;
	wire[2:0] w_G335_1;
	wire[2:0] w_G335_2;
	wire[2:0] w_G335_3;
	wire[1:0] w_G335_4;
	wire[2:0] w_G341_0;
	wire[2:0] w_G341_1;
	wire[2:0] w_G341_2;
	wire[1:0] w_G348_0;
	wire[2:0] w_G351_0;
	wire[2:0] w_G351_1;
	wire[2:0] w_G351_2;
	wire[1:0] w_G358_0;
	wire[2:0] w_G361_0;
	wire[1:0] w_G369_0;
	wire[2:0] w_G374_0;
	wire[2:0] w_G389_0;
	wire[2:0] w_G400_0;
	wire[1:0] w_G400_1;
	wire[2:0] w_G411_0;
	wire[2:0] w_G422_0;
	wire[2:0] w_G422_1;
	wire[1:0] w_G422_2;
	wire[2:0] w_G435_0;
	wire[2:0] w_G435_1;
	wire[2:0] w_G446_0;
	wire[2:0] w_G446_1;
	wire[2:0] w_G457_0;
	wire[2:0] w_G457_1;
	wire[1:0] w_G457_2;
	wire[2:0] w_G468_0;
	wire[2:0] w_G468_1;
	wire[2:0] w_G479_0;
	wire[1:0] w_G479_1;
	wire[2:0] w_G490_0;
	wire[2:0] w_G490_1;
	wire[2:0] w_G503_0;
	wire[2:0] w_G503_1;
	wire[2:0] w_G514_0;
	wire[1:0] w_G514_1;
	wire[2:0] w_G523_0;
	wire[1:0] w_G523_1;
	wire[2:0] w_G534_0;
	wire[2:0] w_G534_1;
	wire[2:0] w_G545_0;
	wire[2:0] w_G549_0;
	wire[1:0] w_G552_0;
	wire[1:0] w_G559_0;
	wire[1:0] w_G562_0;
	wire[2:0] w_G1497_0;
	wire[2:0] w_G1689_0;
	wire[2:0] w_G1690_0;
	wire[2:0] w_G1691_0;
	wire[2:0] w_G1694_0;
	wire[2:0] w_G2174_0;
	wire[2:0] w_G2358_0;
	wire[2:0] w_G2358_1;
	wire[2:0] w_G2358_2;
	wire[1:0] w_G3173_0;
	wire[2:0] w_G3546_0;
	wire[2:0] w_G3546_1;
	wire[2:0] w_G3546_2;
	wire[2:0] w_G3546_3;
	wire[2:0] w_G3546_4;
	wire[1:0] w_G3546_5;
	wire[2:0] w_G3548_0;
	wire[2:0] w_G3548_1;
	wire[2:0] w_G3548_2;
	wire[2:0] w_G3548_3;
	wire[2:0] w_G3548_4;
	wire[1:0] w_G3552_0;
	wire[1:0] w_G3717_0;
	wire[2:0] w_G3724_0;
	wire[2:0] w_G4087_0;
	wire[2:0] w_G4088_0;
	wire[2:0] w_G4089_0;
	wire[2:0] w_G4090_0;
	wire[2:0] w_G4091_0;
	wire[2:0] w_G4091_1;
	wire[2:0] w_G4091_2;
	wire[2:0] w_G4092_0;
	wire[2:0] w_G4092_1;
	wire w_G599_0;
	wire G599_fa_;
	wire w_G600_0;
	wire G600_fa_;
	wire w_G601_0;
	wire G601_fa_;
	wire w_G611_0;
	wire G611_fa_;
	wire w_G612_0;
	wire G612_fa_;
	wire[2:0] w_G809_0;
	wire[2:0] w_G809_1;
	wire[2:0] w_G809_2;
	wire[1:0] w_G809_3;
	wire G809_fa_;
	wire w_G593_0;
	wire G593_fa_;
	wire w_G822_0;
	wire G822_fa_;
	wire w_G838_0;
	wire G838_fa_;
	wire w_G861_0;
	wire G861_fa_;
	wire w_G832_0;
	wire G832_fa_;
	wire w_G834_0;
	wire G834_fa_;
	wire w_G836_0;
	wire G836_fa_;
	wire w_G871_0;
	wire G871_fa_;
	wire w_G873_0;
	wire G873_fa_;
	wire w_G875_0;
	wire G875_fa_;
	wire w_G877_0;
	wire G877_fa_;
	wire w_G1000_0;
	wire G1000_fa_;
	wire w_G826_0;
	wire G826_fa_;
	wire w_G828_0;
	wire G828_fa_;
	wire w_G830_0;
	wire G830_fa_;
	wire w_G867_0;
	wire G867_fa_;
	wire w_G869_0;
	wire G869_fa_;
	wire[1:0] w_n316_0;
	wire[1:0] w_n318_0;
	wire[2:0] w_n326_0;
	wire[2:0] w_n326_1;
	wire[1:0] w_n326_2;
	wire[1:0] w_n333_0;
	wire[1:0] w_n336_0;
	wire[1:0] w_n360_0;
	wire[1:0] w_n362_0;
	wire[2:0] w_n366_0;
	wire[2:0] w_n366_1;
	wire[2:0] w_n366_2;
	wire[2:0] w_n366_3;
	wire[2:0] w_n366_4;
	wire[2:0] w_n368_0;
	wire[2:0] w_n368_1;
	wire[2:0] w_n368_2;
	wire[2:0] w_n368_3;
	wire[2:0] w_n368_4;
	wire[1:0] w_n368_5;
	wire[2:0] w_n372_0;
	wire[1:0] w_n373_0;
	wire[2:0] w_n383_0;
	wire[2:0] w_n385_0;
	wire[2:0] w_n385_1;
	wire[2:0] w_n386_0;
	wire[2:0] w_n386_1;
	wire[2:0] w_n386_2;
	wire[2:0] w_n386_3;
	wire[2:0] w_n386_4;
	wire[2:0] w_n388_0;
	wire[2:0] w_n388_1;
	wire[2:0] w_n389_0;
	wire[2:0] w_n389_1;
	wire[2:0] w_n389_2;
	wire[2:0] w_n389_3;
	wire[2:0] w_n389_4;
	wire[1:0] w_n397_0;
	wire[2:0] w_n398_0;
	wire[2:0] w_n401_0;
	wire[2:0] w_n402_0;
	wire[2:0] w_n402_1;
	wire[1:0] w_n402_2;
	wire[1:0] w_n403_0;
	wire[2:0] w_n405_0;
	wire[2:0] w_n405_1;
	wire[1:0] w_n405_2;
	wire[1:0] w_n407_0;
	wire[1:0] w_n408_0;
	wire[2:0] w_n410_0;
	wire[1:0] w_n410_1;
	wire[1:0] w_n414_0;
	wire[1:0] w_n416_0;
	wire[2:0] w_n419_0;
	wire[2:0] w_n424_0;
	wire[2:0] w_n424_1;
	wire[1:0] w_n424_2;
	wire[1:0] w_n426_0;
	wire[1:0] w_n434_0;
	wire[2:0] w_n435_0;
	wire[2:0] w_n435_1;
	wire[2:0] w_n437_0;
	wire[2:0] w_n437_1;
	wire[1:0] w_n445_0;
	wire[2:0] w_n449_0;
	wire[2:0] w_n449_1;
	wire[2:0] w_n451_0;
	wire[1:0] w_n451_1;
	wire[1:0] w_n459_0;
	wire[2:0] w_n460_0;
	wire[2:0] w_n460_1;
	wire[2:0] w_n462_0;
	wire[1:0] w_n470_0;
	wire[2:0] w_n471_0;
	wire[1:0] w_n471_1;
	wire[2:0] w_n473_0;
	wire[2:0] w_n473_1;
	wire[1:0] w_n481_0;
	wire[2:0] w_n484_0;
	wire[1:0] w_n484_1;
	wire[2:0] w_n486_0;
	wire[1:0] w_n486_1;
	wire[1:0] w_n494_0;
	wire[2:0] w_n495_0;
	wire[2:0] w_n495_1;
	wire[2:0] w_n497_0;
	wire[1:0] w_n497_1;
	wire[1:0] w_n505_0;
	wire[2:0] w_n507_0;
	wire[1:0] w_n507_1;
	wire[1:0] w_n509_0;
	wire[1:0] w_n517_0;
	wire[2:0] w_n518_0;
	wire[1:0] w_n518_1;
	wire[2:0] w_n528_0;
	wire[2:0] w_n530_0;
	wire[1:0] w_n530_1;
	wire[1:0] w_n532_0;
	wire[1:0] w_n540_0;
	wire[2:0] w_n541_0;
	wire[1:0] w_n541_1;
	wire[1:0] w_n543_0;
	wire[1:0] w_n551_0;
	wire[2:0] w_n556_0;
	wire[2:0] w_n556_1;
	wire[2:0] w_n556_2;
	wire[2:0] w_n556_3;
	wire[2:0] w_n556_4;
	wire[1:0] w_n556_5;
	wire[2:0] w_n560_0;
	wire[1:0] w_n560_1;
	wire[2:0] w_n561_0;
	wire[1:0] w_n562_0;
	wire[2:0] w_n566_0;
	wire[2:0] w_n567_0;
	wire[1:0] w_n567_1;
	wire[1:0] w_n569_0;
	wire[1:0] w_n570_0;
	wire[2:0] w_n571_0;
	wire[1:0] w_n571_1;
	wire[2:0] w_n572_0;
	wire[2:0] w_n574_0;
	wire[2:0] w_n577_0;
	wire[2:0] w_n578_0;
	wire[2:0] w_n582_0;
	wire[1:0] w_n582_1;
	wire[2:0] w_n583_0;
	wire[1:0] w_n583_1;
	wire[1:0] w_n585_0;
	wire[2:0] w_n587_0;
	wire[1:0] w_n587_1;
	wire[2:0] w_n590_0;
	wire[1:0] w_n590_1;
	wire[1:0] w_n591_0;
	wire[2:0] w_n595_0;
	wire[1:0] w_n595_1;
	wire[2:0] w_n596_0;
	wire[2:0] w_n600_0;
	wire[1:0] w_n600_1;
	wire[1:0] w_n601_0;
	wire[2:0] w_n604_0;
	wire[2:0] w_n605_0;
	wire[2:0] w_n605_1;
	wire[2:0] w_n605_2;
	wire[2:0] w_n607_0;
	wire[2:0] w_n609_0;
	wire[2:0] w_n609_1;
	wire[2:0] w_n609_2;
	wire[2:0] w_n609_3;
	wire[2:0] w_n609_4;
	wire[2:0] w_n609_5;
	wire[2:0] w_n613_0;
	wire[2:0] w_n614_0;
	wire[2:0] w_n614_1;
	wire[1:0] w_n614_2;
	wire[2:0] w_n617_0;
	wire[1:0] w_n617_1;
	wire[2:0] w_n618_0;
	wire[1:0] w_n618_1;
	wire[2:0] w_n621_0;
	wire[2:0] w_n621_1;
	wire[1:0] w_n621_2;
	wire[2:0] w_n622_0;
	wire[1:0] w_n622_1;
	wire[1:0] w_n623_0;
	wire[2:0] w_n624_0;
	wire[2:0] w_n624_1;
	wire[2:0] w_n625_0;
	wire[2:0] w_n628_0;
	wire[2:0] w_n629_0;
	wire[1:0] w_n631_0;
	wire[2:0] w_n633_0;
	wire[1:0] w_n633_1;
	wire[2:0] w_n636_0;
	wire[1:0] w_n636_1;
	wire[2:0] w_n640_0;
	wire[2:0] w_n640_1;
	wire[1:0] w_n641_0;
	wire[1:0] w_n642_0;
	wire[2:0] w_n645_0;
	wire[2:0] w_n646_0;
	wire[2:0] w_n649_0;
	wire[1:0] w_n649_1;
	wire[1:0] w_n650_0;
	wire[2:0] w_n651_0;
	wire[1:0] w_n651_1;
	wire[1:0] w_n652_0;
	wire[1:0] w_n661_0;
	wire[1:0] w_n671_0;
	wire[1:0] w_n677_0;
	wire[1:0] w_n678_0;
	wire[1:0] w_n679_0;
	wire[1:0] w_n680_0;
	wire[2:0] w_n681_0;
	wire[2:0] w_n681_1;
	wire[1:0] w_n681_2;
	wire[1:0] w_n682_0;
	wire[2:0] w_n687_0;
	wire[1:0] w_n689_0;
	wire[2:0] w_n691_0;
	wire[2:0] w_n693_0;
	wire[2:0] w_n696_0;
	wire[1:0] w_n697_0;
	wire[1:0] w_n700_0;
	wire[1:0] w_n702_0;
	wire[2:0] w_n703_0;
	wire[1:0] w_n705_0;
	wire[1:0] w_n706_0;
	wire[2:0] w_n707_0;
	wire[1:0] w_n709_0;
	wire[1:0] w_n716_0;
	wire[2:0] w_n717_0;
	wire[1:0] w_n720_0;
	wire[2:0] w_n721_0;
	wire[1:0] w_n723_0;
	wire[1:0] w_n726_0;
	wire[2:0] w_n727_0;
	wire[2:0] w_n729_0;
	wire[1:0] w_n729_1;
	wire[2:0] w_n732_0;
	wire[1:0] w_n733_0;
	wire[1:0] w_n735_0;
	wire[1:0] w_n736_0;
	wire[2:0] w_n739_0;
	wire[1:0] w_n739_1;
	wire[1:0] w_n740_0;
	wire[1:0] w_n741_0;
	wire[1:0] w_n742_0;
	wire[2:0] w_n744_0;
	wire[2:0] w_n744_1;
	wire[2:0] w_n746_0;
	wire[2:0] w_n746_1;
	wire[2:0] w_n747_0;
	wire[2:0] w_n747_1;
	wire[2:0] w_n747_2;
	wire[2:0] w_n747_3;
	wire[2:0] w_n748_0;
	wire[2:0] w_n748_1;
	wire[2:0] w_n748_2;
	wire[2:0] w_n748_3;
	wire[1:0] w_n748_4;
	wire[2:0] w_n750_0;
	wire[1:0] w_n750_1;
	wire[2:0] w_n751_0;
	wire[2:0] w_n751_1;
	wire[1:0] w_n751_2;
	wire[2:0] w_n753_0;
	wire[2:0] w_n753_1;
	wire[2:0] w_n753_2;
	wire[2:0] w_n753_3;
	wire[2:0] w_n753_4;
	wire[2:0] w_n753_5;
	wire[2:0] w_n753_6;
	wire[2:0] w_n753_7;
	wire[1:0] w_n753_8;
	wire[1:0] w_n759_0;
	wire[1:0] w_n760_0;
	wire[1:0] w_n761_0;
	wire[2:0] w_n765_0;
	wire[2:0] w_n765_1;
	wire[2:0] w_n765_2;
	wire[2:0] w_n765_3;
	wire[2:0] w_n765_4;
	wire[2:0] w_n765_5;
	wire[1:0] w_n771_0;
	wire[1:0] w_n779_0;
	wire[2:0] w_n781_0;
	wire[2:0] w_n783_0;
	wire[1:0] w_n783_1;
	wire[1:0] w_n786_0;
	wire[1:0] w_n787_0;
	wire[2:0] w_n789_0;
	wire[2:0] w_n791_0;
	wire[1:0] w_n791_1;
	wire[1:0] w_n792_0;
	wire[2:0] w_n793_0;
	wire[2:0] w_n793_1;
	wire[2:0] w_n793_2;
	wire[2:0] w_n793_3;
	wire[1:0] w_n793_4;
	wire[2:0] w_n795_0;
	wire[1:0] w_n795_1;
	wire[1:0] w_n796_0;
	wire[2:0] w_n797_0;
	wire[2:0] w_n797_1;
	wire[2:0] w_n797_2;
	wire[2:0] w_n797_3;
	wire[1:0] w_n797_4;
	wire[2:0] w_n799_0;
	wire[2:0] w_n799_1;
	wire[2:0] w_n799_2;
	wire[2:0] w_n799_3;
	wire[1:0] w_n799_4;
	wire[2:0] w_n801_0;
	wire[2:0] w_n801_1;
	wire[2:0] w_n801_2;
	wire[2:0] w_n801_3;
	wire[1:0] w_n801_4;
	wire[2:0] w_n806_0;
	wire[1:0] w_n809_0;
	wire[1:0] w_n819_0;
	wire[1:0] w_n821_0;
	wire[2:0] w_n828_0;
	wire[1:0] w_n829_0;
	wire[1:0] w_n832_0;
	wire[1:0] w_n839_0;
	wire[2:0] w_n840_0;
	wire[2:0] w_n840_1;
	wire[2:0] w_n840_2;
	wire[2:0] w_n840_3;
	wire[1:0] w_n840_4;
	wire[1:0] w_n842_0;
	wire[2:0] w_n843_0;
	wire[2:0] w_n843_1;
	wire[2:0] w_n843_2;
	wire[2:0] w_n843_3;
	wire[1:0] w_n843_4;
	wire[2:0] w_n845_0;
	wire[2:0] w_n845_1;
	wire[2:0] w_n845_2;
	wire[2:0] w_n845_3;
	wire[1:0] w_n845_4;
	wire[2:0] w_n847_0;
	wire[2:0] w_n847_1;
	wire[2:0] w_n847_2;
	wire[2:0] w_n847_3;
	wire[1:0] w_n847_4;
	wire[1:0] w_n853_0;
	wire[1:0] w_n855_0;
	wire[1:0] w_n856_0;
	wire[1:0] w_n857_0;
	wire[1:0] w_n859_0;
	wire[1:0] w_n862_0;
	wire[1:0] w_n869_0;
	wire[1:0] w_n877_0;
	wire[1:0] w_n879_0;
	wire[1:0] w_n881_0;
	wire[1:0] w_n892_0;
	wire[1:0] w_n914_0;
	wire[1:0] w_n928_0;
	wire[2:0] w_n930_0;
	wire[1:0] w_n932_0;
	wire[2:0] w_n936_0;
	wire[1:0] w_n938_0;
	wire[1:0] w_n941_0;
	wire[1:0] w_n943_0;
	wire[1:0] w_n944_0;
	wire[1:0] w_n946_0;
	wire[2:0] w_n948_0;
	wire[1:0] w_n953_0;
	wire[1:0] w_n954_0;
	wire[1:0] w_n968_0;
	wire[1:0] w_n971_0;
	wire[1:0] w_n972_0;
	wire[1:0] w_n973_0;
	wire[1:0] w_n984_0;
	wire[2:0] w_n985_0;
	wire[2:0] w_n985_1;
	wire[2:0] w_n985_2;
	wire[2:0] w_n985_3;
	wire[1:0] w_n985_4;
	wire[1:0] w_n987_0;
	wire[2:0] w_n988_0;
	wire[2:0] w_n988_1;
	wire[2:0] w_n988_2;
	wire[2:0] w_n988_3;
	wire[1:0] w_n988_4;
	wire[2:0] w_n990_0;
	wire[2:0] w_n990_1;
	wire[2:0] w_n990_2;
	wire[2:0] w_n990_3;
	wire[1:0] w_n990_4;
	wire[2:0] w_n992_0;
	wire[2:0] w_n992_1;
	wire[2:0] w_n992_2;
	wire[2:0] w_n992_3;
	wire[1:0] w_n992_4;
	wire[1:0] w_n998_0;
	wire[2:0] w_n999_0;
	wire[2:0] w_n999_1;
	wire[2:0] w_n999_2;
	wire[2:0] w_n999_3;
	wire[1:0] w_n999_4;
	wire[1:0] w_n1001_0;
	wire[2:0] w_n1002_0;
	wire[2:0] w_n1002_1;
	wire[2:0] w_n1002_2;
	wire[2:0] w_n1002_3;
	wire[1:0] w_n1002_4;
	wire[2:0] w_n1004_0;
	wire[2:0] w_n1004_1;
	wire[2:0] w_n1004_2;
	wire[2:0] w_n1004_3;
	wire[1:0] w_n1004_4;
	wire[2:0] w_n1006_0;
	wire[2:0] w_n1006_1;
	wire[2:0] w_n1006_2;
	wire[2:0] w_n1006_3;
	wire[1:0] w_n1006_4;
	wire[2:0] w_n1012_0;
	wire[1:0] w_n1012_1;
	wire[2:0] w_n1014_0;
	wire[1:0] w_n1014_1;
	wire[2:0] w_n1021_0;
	wire[1:0] w_n1021_1;
	wire[2:0] w_n1023_0;
	wire[1:0] w_n1023_1;
	wire[2:0] w_n1030_0;
	wire[1:0] w_n1030_1;
	wire[2:0] w_n1032_0;
	wire[1:0] w_n1032_1;
	wire[2:0] w_n1039_0;
	wire[1:0] w_n1039_1;
	wire[2:0] w_n1041_0;
	wire[1:0] w_n1041_1;
	wire[1:0] w_n1142_0;
	wire[1:0] w_n1151_0;
	wire[2:0] w_n1163_0;
	wire[2:0] w_n1163_1;
	wire[2:0] w_n1197_0;
	wire[2:0] w_n1197_1;
	wire[2:0] w_n1205_0;
	wire[2:0] w_n1205_1;
	wire[2:0] w_n1235_0;
	wire[1:0] w_n1235_1;
	wire[2:0] w_n1242_0;
	wire[1:0] w_n1242_1;
	wire[2:0] w_n1244_0;
	wire[1:0] w_n1244_1;
	wire[2:0] w_n1251_0;
	wire[1:0] w_n1251_1;
	wire[2:0] w_n1253_0;
	wire[1:0] w_n1253_1;
	wire[1:0] w_n1358_0;
	wire[1:0] w_n1383_0;
	wire[1:0] w_n1391_0;
	wire[1:0] w_n1394_0;
	wire[1:0] w_n1398_0;
	wire[1:0] w_n1399_0;
	wire[1:0] w_n1409_0;
	wire[1:0] w_n1410_0;
	wire[1:0] w_n1411_0;
	wire[1:0] w_n1421_0;
	wire[1:0] w_n1425_0;
	wire[1:0] w_n1434_0;
	wire[1:0] w_n1438_0;
	wire[1:0] w_n1445_0;
	wire[1:0] w_n1446_0;
	wire[1:0] w_n1447_0;
	wire[1:0] w_n1452_0;
	wire[1:0] w_n1494_0;
	wire[1:0] w_n1533_0;
	wire[1:0] w_n1543_0;
	wire[1:0] w_n1545_0;
	wire[1:0] w_n1553_0;
	wire[1:0] w_n1555_0;
	wire[1:0] w_n1560_0;
	wire[1:0] w_n1568_0;
	wire[1:0] w_n1591_0;
	wire[1:0] w_n1597_0;
	wire[2:0] w_n1601_0;
	wire[1:0] w_n1602_0;
	wire[1:0] w_n1609_0;
	wire[1:0] w_n1610_0;
	wire[1:0] w_n1624_0;
	wire[1:0] w_n1629_0;
	wire[1:0] w_n1631_0;
	wire[1:0] w_n1634_0;
	wire w_dff_B_jHQBTdJq4_1;
	wire w_dff_B_Anr4sdjm6_0;
	wire w_dff_B_IMmybuoF8_1;
	wire w_dff_B_NU61lJJ87_1;
	wire w_dff_B_UXVU0Ypt4_2;
	wire w_dff_B_gm4p0GP46_1;
	wire w_dff_B_623LmuQ12_1;
	wire w_dff_B_wR4gaxUk6_0;
	wire w_dff_B_vHWIvW9o5_1;
	wire w_dff_B_pHBgUaoW0_1;
	wire w_dff_B_IxahGZvQ1_0;
	wire w_dff_B_vtIH2h1n6_1;
	wire w_dff_A_ttLXDYX95_0;
	wire w_dff_A_biDTaEoA3_0;
	wire w_dff_A_YeISUY517_0;
	wire w_dff_A_IMIxIDym3_0;
	wire w_dff_A_f89PYxzO7_1;
	wire w_dff_A_hYDteRYp4_1;
	wire w_dff_A_nBSVcUOf5_1;
	wire w_dff_A_Uix9emZd8_1;
	wire w_dff_B_aqsw1dbN5_1;
	wire w_dff_B_DHaR4A7J8_0;
	wire w_dff_B_gnNJIjpj5_1;
	wire w_dff_B_KqiineDQ9_1;
	wire w_dff_B_PDQFZ4RW9_0;
	wire w_dff_B_4YYVXK1V0_1;
	wire w_dff_A_5EOTA0Rs8_0;
	wire w_dff_A_BkHOyTil1_1;
	wire w_dff_A_yzdqWlka0_1;
	wire w_dff_A_kX2rJmue8_1;
	wire w_dff_A_ys9Qfu3j7_1;
	wire w_dff_A_FVxwN3J96_1;
	wire w_dff_A_CxbGlPds6_2;
	wire w_dff_A_rAKqKSGo9_2;
	wire w_dff_A_A6FfpvXM3_2;
	wire w_dff_A_JcqojU074_2;
	wire w_dff_B_ltj41sKF6_1;
	wire w_dff_B_f3ch99Z31_1;
	wire w_dff_B_eAqgYHn04_0;
	wire w_dff_B_5mlsIGkR7_1;
	wire w_dff_B_uVRcF1Sl0_1;
	wire w_dff_B_7iy6Kj3D8_2;
	wire w_dff_B_pPvj2W9G7_2;
	wire w_dff_B_UJrFruSB3_2;
	wire w_dff_B_aRARWFLQ8_2;
	wire w_dff_B_3yN88npG8_1;
	wire w_dff_B_pEkfxiGf8_1;
	wire w_dff_B_SmeA8bAj8_1;
	wire w_dff_B_pRP80RRX9_1;
	wire w_dff_B_1amRu1IJ8_1;
	wire w_dff_B_Zpe9KJPW8_1;
	wire w_dff_B_NZ2J9zDL7_1;
	wire w_dff_A_Xin0Blvm9_1;
	wire w_dff_A_I5VwRkAh7_1;
	wire w_dff_B_ZINqSSK07_3;
	wire w_dff_B_7Esi7QlS2_3;
	wire w_dff_B_t1QjbpLO5_3;
	wire w_dff_B_hGOH1ICO8_0;
	wire w_dff_B_8Hj9RYZR3_2;
	wire w_dff_B_B8YsHfHS2_2;
	wire w_dff_B_UDI6drwr2_2;
	wire w_dff_B_ZUBpmoAa7_2;
	wire w_dff_B_jfeEQVgx4_2;
	wire w_dff_A_iJp98zHA5_0;
	wire w_dff_A_LAQ99uND5_0;
	wire w_dff_A_b9W3XuLC8_0;
	wire w_dff_A_RNM0zKFw2_0;
	wire w_dff_A_0kVWVmWh9_0;
	wire w_dff_A_IG1CENs25_0;
	wire w_dff_B_vG7gIifi5_0;
	wire w_dff_B_oEWPo6Ko6_0;
	wire w_dff_B_rwu1TT7A8_0;
	wire w_dff_B_nP2d2A7c6_0;
	wire w_dff_B_jUkZISbW0_0;
	wire w_dff_B_zMkpzVqJ5_0;
	wire w_dff_B_z7dgp7jw4_0;
	wire w_dff_B_MZks48Sf6_0;
	wire w_dff_B_gg7adqYB2_0;
	wire w_dff_B_roUtmP064_0;
	wire w_dff_B_hYePd4Ob5_0;
	wire w_dff_B_Mt1TyOcg4_0;
	wire w_dff_B_nWHyNTeU4_2;
	wire w_dff_B_CGOjwWy20_2;
	wire w_dff_B_LLUKbs4O8_2;
	wire w_dff_B_HAwExXEz6_0;
	wire w_dff_B_UP050EU05_0;
	wire w_dff_B_TVnOlHoq5_0;
	wire w_dff_B_YZtlb9hF8_1;
	wire w_dff_B_w7DtqsC31_1;
	wire w_dff_B_7g3InhJ04_1;
	wire w_dff_B_qfGQmnHK9_1;
	wire w_dff_B_4Nihpq5s8_0;
	wire w_dff_B_IJUhH4ns3_0;
	wire w_dff_B_HrMMq4VJ6_0;
	wire w_dff_B_KMqjl7ai9_0;
	wire w_dff_B_XrSWrNTy2_0;
	wire w_dff_B_CGVCrTK19_0;
	wire w_dff_B_UEhCmxNW0_0;
	wire w_dff_B_uATN87N69_0;
	wire w_dff_B_ByQQJMxZ3_0;
	wire w_dff_B_mZX2pVJF1_0;
	wire w_dff_B_X5Rb88TQ7_0;
	wire w_dff_B_ryjvrocQ2_0;
	wire w_dff_B_cj0VNEgI1_0;
	wire w_dff_B_aspS6po80_0;
	wire w_dff_B_PpZaZXXs6_0;
	wire w_dff_B_RRch3qeI3_0;
	wire w_dff_B_4EEW3udA8_0;
	wire w_dff_B_EbjnnGtL5_0;
	wire w_dff_B_EftrGcDC3_2;
	wire w_dff_B_a96C1oTs3_2;
	wire w_dff_B_qds7jQhf3_2;
	wire w_dff_B_oJLhhSj89_1;
	wire w_dff_B_PFf9ptfD2_0;
	wire w_dff_B_31XDNprI8_1;
	wire w_dff_B_BOB3AgmJ6_1;
	wire w_dff_B_QO11U0RQ4_0;
	wire w_dff_B_QnR3iPsJ1_0;
	wire w_dff_B_RJNpD09T1_1;
	wire w_dff_B_pIbDnPuQ1_1;
	wire w_dff_B_OCIN2bTo6_0;
	wire w_dff_B_jwquK25w5_1;
	wire w_dff_B_ce2DHmUC9_0;
	wire w_dff_B_lHQ5ViY04_0;
	wire w_dff_B_CfaUw6c81_0;
	wire w_dff_B_lpwUEjfF0_0;
	wire w_dff_B_Jt3xcbBB6_0;
	wire w_dff_B_1knAGKCk6_0;
	wire w_dff_B_XrFOhDIu0_0;
	wire w_dff_B_3AsR27S58_0;
	wire w_dff_B_orBbCIVg6_0;
	wire w_dff_B_6LIagr1I1_0;
	wire w_dff_B_ZjDAteSM8_0;
	wire w_dff_B_DOJq9JIz6_0;
	wire w_dff_B_ITRFDaAA8_0;
	wire w_dff_B_Q0VfgMkX4_0;
	wire w_dff_A_0rf7psYY1_0;
	wire w_dff_A_AW4savrb3_0;
	wire w_dff_A_gkNdMhPI6_0;
	wire w_dff_A_vj2YgRVs5_0;
	wire w_dff_A_RN1eUI9Y0_0;
	wire w_dff_A_ACvQgDkR0_0;
	wire w_dff_A_yGyRJSXA9_0;
	wire w_dff_A_trJ3JV1b3_0;
	wire w_dff_A_TaAECb3k8_0;
	wire w_dff_A_JmnIQOFK1_0;
	wire w_dff_A_Ypf1M73J5_0;
	wire w_dff_A_cLKTDLD97_0;
	wire w_dff_A_vq5XQZJv8_0;
	wire w_dff_A_bCGTqDzo5_0;
	wire w_dff_A_zKo6lCdE9_0;
	wire w_dff_B_plgG2qC08_0;
	wire w_dff_B_m3Rr661J6_0;
	wire w_dff_B_9Z7rjXjx7_0;
	wire w_dff_B_6IdFPoG57_0;
	wire w_dff_B_OYphEQiZ5_0;
	wire w_dff_B_3zQhCRk18_0;
	wire w_dff_B_hMqcxCjY6_0;
	wire w_dff_B_X4zi9jxB5_0;
	wire w_dff_B_RhiIaZXb6_0;
	wire w_dff_B_K9Mfqw101_0;
	wire w_dff_B_SBR2JHGD2_0;
	wire w_dff_B_yJdSPpJm7_0;
	wire w_dff_B_vUQkrHzj0_0;
	wire w_dff_B_LN2JCHDe2_0;
	wire w_dff_B_u22uWexP5_0;
	wire w_dff_B_nHTc1oyJ6_0;
	wire w_dff_B_rS1GjpzH9_0;
	wire w_dff_B_ZBJWExEA4_0;
	wire w_dff_B_zX6Zn8ZF2_0;
	wire w_dff_B_lWqwbSZy1_0;
	wire w_dff_B_yH1IjA8i5_0;
	wire w_dff_B_b1Bo3pNX3_0;
	wire w_dff_B_FTDf6ngq6_0;
	wire w_dff_B_mNjZmzVF3_0;
	wire w_dff_B_0jpKrJJW7_0;
	wire w_dff_B_yvilTlyr0_0;
	wire w_dff_B_sIGWFB6b0_0;
	wire w_dff_B_3ksMGvfV8_0;
	wire w_dff_B_xJJ6kDRm3_0;
	wire w_dff_B_PDhjoWO68_0;
	wire w_dff_B_vnKuuCMV3_0;
	wire w_dff_B_vpAFIKRV2_0;
	wire w_dff_B_d4K1Bo386_0;
	wire w_dff_A_7JrfLBXL2_1;
	wire w_dff_A_RzFTeu7T9_1;
	wire w_dff_A_85wekFvO6_2;
	wire w_dff_A_qLmNRbxh1_2;
	wire w_dff_A_76Z9Oaut4_2;
	wire w_dff_A_ryKJwIR74_2;
	wire w_dff_A_cyhATo4q5_1;
	wire w_dff_A_wxcAGRZI2_2;
	wire w_dff_A_Z3YaYsW56_2;
	wire w_dff_B_x28AR9oc9_0;
	wire w_dff_B_LaWn1N7U4_0;
	wire w_dff_B_ZrmOjU6m7_0;
	wire w_dff_B_loOHNNpY6_0;
	wire w_dff_B_ROeYGZA83_0;
	wire w_dff_B_HqruB29x5_0;
	wire w_dff_B_f3GWPNL62_0;
	wire w_dff_B_p4vcI9nz8_0;
	wire w_dff_B_H8zwpshB5_0;
	wire w_dff_B_tzFAyP2l8_0;
	wire w_dff_B_sGlEKDiE9_0;
	wire w_dff_B_aUQ55GmA8_0;
	wire w_dff_B_1rrl11Yh9_0;
	wire w_dff_B_9M5xc7r91_0;
	wire w_dff_B_IvRLvBDD0_2;
	wire w_dff_B_7tPDAO0p0_2;
	wire w_dff_B_aMcOYz5D7_2;
	wire w_dff_A_nRNZJ5p44_0;
	wire w_dff_A_ExQoIyrZ9_0;
	wire w_dff_A_INilhmeI0_0;
	wire w_dff_A_AbgE24Bn4_0;
	wire w_dff_A_Vpfju6Nd8_0;
	wire w_dff_A_1Eq9JByu5_0;
	wire w_dff_A_xlSSDrBy9_0;
	wire w_dff_A_hfEVaF540_0;
	wire w_dff_A_iNpUN3Wl3_0;
	wire w_dff_A_ESEnQAr29_0;
	wire w_dff_A_ePefduiP3_0;
	wire w_dff_A_6aeXJ5yw8_0;
	wire w_dff_A_fdUw5kI28_0;
	wire w_dff_A_NWVKWA597_0;
	wire w_dff_A_QcC28Cyj4_0;
	wire w_dff_B_mytJ3CSB9_0;
	wire w_dff_B_STI7cpBA1_0;
	wire w_dff_B_craCbSdK1_0;
	wire w_dff_B_C4JaHRpC0_0;
	wire w_dff_B_6QMXdnGr6_0;
	wire w_dff_B_2HZQdbdX4_0;
	wire w_dff_B_PU0Xr1cP7_0;
	wire w_dff_B_TSbbCI2R9_0;
	wire w_dff_B_QZ7gkqiz8_0;
	wire w_dff_B_OBjHl8bY0_0;
	wire w_dff_B_cfNDjJPe0_0;
	wire w_dff_B_4YYQYK7A9_0;
	wire w_dff_B_u64XRs6s1_2;
	wire w_dff_B_fRvmqErS7_2;
	wire w_dff_B_XzoOlpDi0_2;
	wire w_dff_B_iROGU24a0_0;
	wire w_dff_B_GrUuGhbS2_0;
	wire w_dff_B_RN01pbPJ3_0;
	wire w_dff_B_VgKMD2p48_0;
	wire w_dff_B_wSU9UURo8_0;
	wire w_dff_B_eeh6DvYa5_0;
	wire w_dff_B_TBZmTWlY8_0;
	wire w_dff_B_EWjObTSD2_0;
	wire w_dff_B_5wCpzg9F2_0;
	wire w_dff_B_v63e2pER8_0;
	wire w_dff_B_pwMPdJHW0_0;
	wire w_dff_B_e6C6fCKi5_2;
	wire w_dff_B_gF9J4mhZ7_2;
	wire w_dff_B_cUq7hYYo7_2;
	wire w_dff_B_U01SPKza4_0;
	wire w_dff_B_HNulD6EV5_0;
	wire w_dff_B_pIpn7ApU6_0;
	wire w_dff_B_HBzwF5yD2_0;
	wire w_dff_B_hGLN6FZ34_0;
	wire w_dff_B_GC3UT7hB7_0;
	wire w_dff_B_TiArMLyD8_0;
	wire w_dff_B_Kz42r3AX1_0;
	wire w_dff_B_YZqsccn93_0;
	wire w_dff_B_4tTd2lKx5_0;
	wire w_dff_B_9xJiJbm46_2;
	wire w_dff_B_d0nNtj9g6_2;
	wire w_dff_B_PKSteptA6_2;
	wire w_dff_A_32xajYbh3_1;
	wire w_dff_A_J7Dd7AbO5_1;
	wire w_dff_A_eoTcwGK65_2;
	wire w_dff_A_gYXcvBaG9_2;
	wire w_dff_A_vflnmgKr7_2;
	wire w_dff_A_8OsilrIV3_2;
	wire w_dff_A_dRZ0fmRA0_1;
	wire w_dff_A_Ye90dm7A3_2;
	wire w_dff_A_oajukjWu6_2;
	wire w_dff_B_i4lPnUWI4_0;
	wire w_dff_B_eYCPyy3l6_0;
	wire w_dff_B_NQvq1k092_0;
	wire w_dff_B_JvAyIygj0_0;
	wire w_dff_B_sAN1nCmR0_0;
	wire w_dff_B_3cwXepcK3_0;
	wire w_dff_B_J6ocffbi6_0;
	wire w_dff_B_R98uW9kW2_0;
	wire w_dff_B_LsWCv4p96_0;
	wire w_dff_B_qfU9wApL3_0;
	wire w_dff_B_b48h3PoD0_0;
	wire w_dff_B_kCdUc63p2_0;
	wire w_dff_B_NZAe3sJK5_0;
	wire w_dff_B_Rge1IOJ90_0;
	wire w_dff_A_EjGxEXaG5_0;
	wire w_dff_A_Nkrkw3fs8_0;
	wire w_dff_A_t2RnZ8zQ1_0;
	wire w_dff_A_75LsJQEN2_0;
	wire w_dff_A_cYHaD0Dj2_0;
	wire w_dff_A_gQgyRyRP6_0;
	wire w_dff_A_EpbnYmIi7_0;
	wire w_dff_A_jIUiAxKc8_0;
	wire w_dff_A_GVHxFxes7_0;
	wire w_dff_A_Z2SXCxO75_0;
	wire w_dff_A_G6LaeZFv6_0;
	wire w_dff_A_4slQe8Pt6_0;
	wire w_dff_A_DdZU23Bq4_0;
	wire w_dff_A_ew1ezB1N1_0;
	wire w_dff_A_uIUJ1IzD8_0;
	wire w_dff_B_2Pb3NNG52_0;
	wire w_dff_B_FMadaEYd7_0;
	wire w_dff_B_1H19wOa74_0;
	wire w_dff_B_hYM7vp0g1_0;
	wire w_dff_B_7KwvDgKt5_0;
	wire w_dff_B_l66hWUEN6_0;
	wire w_dff_B_3cejkBvY1_0;
	wire w_dff_B_0G81fxKi8_0;
	wire w_dff_B_jFd1qzXD8_0;
	wire w_dff_B_KuXXw29b6_0;
	wire w_dff_B_4ZNA6fgK6_0;
	wire w_dff_B_aVoZ8Ga37_0;
	wire w_dff_B_pF19CPtU6_0;
	wire w_dff_B_ViHDmc1t2_0;
	wire w_dff_B_hMZc7jZp0_0;
	wire w_dff_B_uVxzigAs6_0;
	wire w_dff_B_QR9s0JAM1_0;
	wire w_dff_B_0PBDAjt86_0;
	wire w_dff_B_59nsSvop7_0;
	wire w_dff_B_j2lnXHmC3_0;
	wire w_dff_B_JL4tlOpu9_0;
	wire w_dff_A_tpjrM7qL1_0;
	wire w_dff_A_AOW9vASK1_2;
	wire w_dff_A_7nfAVQrl2_2;
	wire w_dff_A_y0Z6Nrwr3_2;
	wire w_dff_A_73R8StKX9_2;
	wire w_dff_B_9CDm9T0x5_0;
	wire w_dff_B_vlVnsMvO5_0;
	wire w_dff_B_BLw0u94p0_0;
	wire w_dff_B_1FajR0dB6_0;
	wire w_dff_B_YSqoDrPk3_0;
	wire w_dff_B_tVkZpNZL2_0;
	wire w_dff_B_m89Tvkcf8_0;
	wire w_dff_B_7ydwjWxg0_0;
	wire w_dff_B_lg9jCVoM4_0;
	wire w_dff_B_t7Nkqp0I4_0;
	wire w_dff_B_6HOKj66b5_0;
	wire w_dff_B_ZRYI2TIt9_0;
	wire w_dff_A_DHoUckhx8_0;
	wire w_dff_A_TqZ9U7wu1_0;
	wire w_dff_A_sO5VoXT98_0;
	wire w_dff_A_xOGvZE8S0_0;
	wire w_dff_A_Ufuh4jZt8_1;
	wire w_dff_A_60Bj9an54_1;
	wire w_dff_A_uWTwpn385_0;
	wire w_dff_A_9ez9Zel48_0;
	wire w_dff_A_nznAk0ZQ3_1;
	wire w_dff_B_l1zv4hd97_0;
	wire w_dff_B_O7nBV4Ua1_0;
	wire w_dff_B_vLLMvwMo3_0;
	wire w_dff_B_bKARqemA7_0;
	wire w_dff_B_Smt4RTLZ0_0;
	wire w_dff_B_zXRJjpeM1_0;
	wire w_dff_B_DtqhJbsK6_0;
	wire w_dff_B_gX4stcmz0_0;
	wire w_dff_B_sbCtviuo5_0;
	wire w_dff_B_gnfciyQk9_0;
	wire w_dff_B_eCOwXywu2_0;
	wire w_dff_B_taxkirQY8_0;
	wire w_dff_B_SbyRTDjy5_0;
	wire w_dff_B_Gg9m0Kkv7_0;
	wire w_dff_B_K0FZ46m73_2;
	wire w_dff_B_nGol4eN09_2;
	wire w_dff_B_twHeLHGu2_2;
	wire w_dff_A_pP48pqUT3_0;
	wire w_dff_A_iWfVGpi39_0;
	wire w_dff_A_SqWgLEWl4_0;
	wire w_dff_A_uQP2s3dW3_0;
	wire w_dff_A_3rDjW8yQ0_0;
	wire w_dff_A_vjN9xg9H3_0;
	wire w_dff_A_JvDkBFwb9_0;
	wire w_dff_B_TmoIExVY3_0;
	wire w_dff_B_E9SCZhH61_0;
	wire w_dff_B_5QvAAI5y1_0;
	wire w_dff_B_F3FTmgG70_0;
	wire w_dff_B_bZPZhxkA1_0;
	wire w_dff_B_XsD4gAUV9_0;
	wire w_dff_B_rOEIVskU0_0;
	wire w_dff_B_IgbdpG980_0;
	wire w_dff_B_gbIj66MZ7_1;
	wire w_dff_B_SuVya2Y11_1;
	wire w_dff_B_9zStGqWt6_0;
	wire w_dff_B_axKllIrL3_1;
	wire w_dff_A_xlue22Q54_0;
	wire w_dff_A_KdOGbMLL6_0;
	wire w_dff_A_80YT3jAo2_0;
	wire w_dff_A_zU6SIoox2_0;
	wire w_dff_A_M8aBhL1B2_0;
	wire w_dff_A_1pmCv7j60_0;
	wire w_dff_A_6GGIEMOB6_0;
	wire w_dff_A_HWZNkgDO3_0;
	wire w_dff_B_DZkZdZUp1_0;
	wire w_dff_B_mhqjkvYJ0_0;
	wire w_dff_B_UtB3UMPE8_0;
	wire w_dff_B_EEa1HfNm6_0;
	wire w_dff_B_iUyJeIbm4_0;
	wire w_dff_B_kSsGghPM6_0;
	wire w_dff_B_uvfMouT79_0;
	wire w_dff_B_tCVmtduJ1_0;
	wire w_dff_B_7CGqfLAq3_0;
	wire w_dff_B_fidH2dRX4_0;
	wire w_dff_B_ZC1X76HY8_1;
	wire w_dff_B_5w8VRhtv0_1;
	wire w_dff_B_0p97Hk5s7_0;
	wire w_dff_B_xgN6JT9C7_1;
	wire w_dff_B_attAywGa0_1;
	wire w_dff_B_uJk4IlmZ2_1;
	wire w_dff_B_jX659Nua3_1;
	wire w_dff_B_zOSiBFZS0_1;
	wire w_dff_B_YmxJ9Gyc1_1;
	wire w_dff_B_6IfT1C051_1;
	wire w_dff_B_pzdm031y7_0;
	wire w_dff_B_VmOlFNzb2_0;
	wire w_dff_B_i29EUwTc3_0;
	wire w_dff_B_nOiZL7CW0_0;
	wire w_dff_B_4T0K47LW5_0;
	wire w_dff_B_znoCPcj97_0;
	wire w_dff_B_CgxpWkET1_0;
	wire w_dff_B_GosTMdDX1_0;
	wire w_dff_B_FCy4cNJc8_0;
	wire w_dff_B_dLAyJeXu7_0;
	wire w_dff_B_Xx8Rvxsi8_2;
	wire w_dff_B_OpNkcJd51_2;
	wire w_dff_B_AmPL2t1L6_2;
	wire w_dff_B_p2GlV8Jy7_0;
	wire w_dff_B_I3ZfaRf29_0;
	wire w_dff_B_XtwerSJ70_1;
	wire w_dff_B_4HXG8lg23_1;
	wire w_dff_A_63OKJmVU5_1;
	wire w_dff_B_xSRV8uDk0_0;
	wire w_dff_B_VYhf0rRg0_1;
	wire w_dff_A_iUVppLLC3_0;
	wire w_dff_B_Kyt5Sm5b4_0;
	wire w_dff_B_mk7f2KNx4_0;
	wire w_dff_B_4ecwqkZP1_0;
	wire w_dff_B_vNdBs2kk8_0;
	wire w_dff_B_Tk4bzhyF1_0;
	wire w_dff_B_RCstnGuM4_0;
	wire w_dff_B_StH4f6bM9_1;
	wire w_dff_B_HudtHNcR4_1;
	wire w_dff_B_jgVxFdhx8_0;
	wire w_dff_B_aqDUyMwi0_1;
	wire w_dff_B_L93O4wiF6_0;
	wire w_dff_A_mnovzVWq8_1;
	wire w_dff_A_TgrU2gMY9_1;
	wire w_dff_A_83YjOvyh2_1;
	wire w_dff_A_JJMcdgTq7_1;
	wire w_dff_A_Bo1joco45_2;
	wire w_dff_A_3Z2ePtAG1_2;
	wire w_dff_A_JQQuOTlV8_0;
	wire w_dff_A_dE52QEdm5_0;
	wire w_dff_A_dgFbPYSa1_0;
	wire w_dff_A_lp1paIgS1_0;
	wire w_dff_A_gbgVv3vG8_1;
	wire w_dff_A_M96opvhU6_1;
	wire w_dff_A_y4CvdwjM4_1;
	wire w_dff_A_HWQavakt8_1;
	wire w_dff_B_8NqKbRgT0_0;
	wire w_dff_B_db45aS7f7_0;
	wire w_dff_B_b2Kv6wiO3_0;
	wire w_dff_B_4K5w1RAJ4_0;
	wire w_dff_B_8WeFoxZH2_0;
	wire w_dff_B_IZ8sqVnY6_0;
	wire w_dff_B_1lDDg48k9_0;
	wire w_dff_B_kQPD1IDn1_0;
	wire w_dff_B_KRHTHDfL9_0;
	wire w_dff_B_DgGrCXuz6_0;
	wire w_dff_B_iywwfrfp0_0;
	wire w_dff_B_nJEeufId6_2;
	wire w_dff_B_cPKK66sL5_2;
	wire w_dff_B_Hr5Ef1GE8_2;
	wire w_dff_B_eTOjnUJH1_0;
	wire w_dff_B_Y9Tox2yI6_0;
	wire w_dff_B_d2tuIZ0h6_0;
	wire w_dff_B_0cnio3gY3_0;
	wire w_dff_B_soVvpI2f9_1;
	wire w_dff_B_6P5kMzZz0_1;
	wire w_dff_B_Ub8q9oaB2_0;
	wire w_dff_B_8S4t6fQz2_1;
	wire w_dff_A_ifTUOtl82_0;
	wire w_dff_A_zmsw4He95_0;
	wire w_dff_A_v2FYbrdu1_0;
	wire w_dff_A_uCaByIzH4_0;
	wire w_dff_A_f9tb60g82_0;
	wire w_dff_A_4v02IntC4_0;
	wire w_dff_B_zk4Cjs9z8_0;
	wire w_dff_B_qGCxqqTx3_0;
	wire w_dff_B_DTINZc7i8_0;
	wire w_dff_B_A4XoTYjY2_0;
	wire w_dff_B_fCDC6jCd4_0;
	wire w_dff_B_7f9Yqb9p3_0;
	wire w_dff_B_SUKWI2E52_0;
	wire w_dff_B_O8ilfwh16_1;
	wire w_dff_B_JkvKrsif8_1;
	wire w_dff_A_9vwwXxKD4_1;
	wire w_dff_B_aqqTLBTb6_0;
	wire w_dff_B_YQcTVDeX3_1;
	wire w_dff_B_wvmvDo3N4_0;
	wire w_dff_B_fIZA17lP3_0;
	wire w_dff_B_DvjY02gE6_0;
	wire w_dff_B_XYgIO2Lu7_0;
	wire w_dff_B_679AlWQc6_0;
	wire w_dff_B_V8jDugkm8_0;
	wire w_dff_B_Y3TkIGnK5_0;
	wire w_dff_B_onUrTJDO2_0;
	wire w_dff_B_2iN4p2J15_0;
	wire w_dff_B_rERWmI323_0;
	wire w_dff_B_WWmRkjpa6_0;
	wire w_dff_B_V1GNE4et7_0;
	wire w_dff_B_p5VKIVOZ9_2;
	wire w_dff_B_ykPNCXRN2_2;
	wire w_dff_B_VdpNh2Zg3_2;
	wire w_dff_A_zULHyfoe2_0;
	wire w_dff_A_XenlyZdW2_0;
	wire w_dff_A_bwyYPt6z6_0;
	wire w_dff_A_kfhIpUYa8_0;
	wire w_dff_A_GiaJWmrs0_1;
	wire w_dff_A_lDdfJqoX7_1;
	wire w_dff_B_9TjBKOBe6_0;
	wire w_dff_B_YpB0HddL0_0;
	wire w_dff_B_lorW02c28_0;
	wire w_dff_B_8lKEEDpE1_0;
	wire w_dff_B_Ny5gWR5V1_0;
	wire w_dff_B_SfDirKpW0_0;
	wire w_dff_B_QzOQW9zY4_1;
	wire w_dff_B_MZ5fi9cp2_1;
	wire w_dff_B_lTcAT0Ce7_0;
	wire w_dff_B_VORGvKop1_1;
	wire w_dff_B_Sk8udyQC8_1;
	wire w_dff_B_h6bF9BiN0_1;
	wire w_dff_B_SbwYihbX8_1;
	wire w_dff_B_exRqFS4L6_1;
	wire w_dff_A_PPOdDa8V8_2;
	wire w_dff_A_ICgvkPBk2_2;
	wire w_dff_A_eYXBz0vJ8_2;
	wire w_dff_A_AhU7oceG6_2;
	wire w_dff_B_n7jQxknP7_3;
	wire w_dff_B_IRVa1Pmb5_3;
	wire w_dff_A_2uWg91iH6_1;
	wire w_dff_A_8g0vU4iT8_1;
	wire w_dff_A_zbzUghjV0_2;
	wire w_dff_A_EJ0STCnJ7_2;
	wire w_dff_A_lzzscTAx1_2;
	wire w_dff_A_4NeCTvRO6_2;
	wire w_dff_A_lRHEjDTu5_0;
	wire w_dff_A_33UYVb7Q4_0;
	wire w_dff_A_1nYUCOUx3_1;
	wire w_dff_B_HxKjyXgw0_0;
	wire w_dff_B_xC1SjRwX8_0;
	wire w_dff_B_OyxPJ0tF4_0;
	wire w_dff_B_mIpnp5UF0_0;
	wire w_dff_B_HQ3sJb4f2_0;
	wire w_dff_B_DggdxiwR2_0;
	wire w_dff_B_N2QLohcD1_0;
	wire w_dff_B_xHXuatwA1_0;
	wire w_dff_B_sBsDkjNf9_1;
	wire w_dff_B_RdiaBO6R4_1;
	wire w_dff_B_SzZAg0xl2_0;
	wire w_dff_B_Owewop3E6_1;
	wire w_dff_B_5todjbo18_0;
	wire w_dff_A_hmZACMxk8_0;
	wire w_dff_A_R9unRN3k7_0;
	wire w_dff_A_YeufBsyB9_0;
	wire w_dff_A_Xsi80K702_0;
	wire w_dff_B_OQo50X6U1_0;
	wire w_dff_B_Ilzeax6d3_0;
	wire w_dff_B_bOa9Utrz7_0;
	wire w_dff_B_uHTSgQkm2_0;
	wire w_dff_B_MsNhVbX91_0;
	wire w_dff_B_AHIgh2vR2_0;
	wire w_dff_B_iziWwFyk4_0;
	wire w_dff_B_kPhERWyU0_0;
	wire w_dff_B_KBIWN7di2_0;
	wire w_dff_B_DxHOchE57_0;
	wire w_dff_B_adloSAdU0_0;
	wire w_dff_B_j74uReLR5_0;
	wire w_dff_B_yblj741h6_1;
	wire w_dff_B_9VscNHJl5_1;
	wire w_dff_B_gqoiLU3g3_1;
	wire w_dff_B_gQw9j5Cc2_1;
	wire w_dff_B_eI2359Qg3_1;
	wire w_dff_B_HixqNAtj8_1;
	wire w_dff_B_I1nJ34tq1_0;
	wire w_dff_B_zK58RImn5_0;
	wire w_dff_B_ILi98yKd8_0;
	wire w_dff_B_S2mQ5caC3_0;
	wire w_dff_B_iZqf4yul8_0;
	wire w_dff_B_UHrS96262_0;
	wire w_dff_B_Zuaqtahp2_0;
	wire w_dff_B_7JSgG3i04_0;
	wire w_dff_B_ebQFglhz0_0;
	wire w_dff_B_hHIZ0iXp5_0;
	wire w_dff_B_VDvsx6FZ6_0;
	wire w_dff_B_5UYAlVGf3_0;
	wire w_dff_B_cGTaa0N48_0;
	wire w_dff_B_4YmmOZDP2_0;
	wire w_dff_B_JaxA3jff9_0;
	wire w_dff_B_i7iBOFlZ4_0;
	wire w_dff_B_ugPAGpWl0_1;
	wire w_dff_A_4XsvK0hY4_0;
	wire w_dff_A_VELsOET54_0;
	wire w_dff_A_QgDlqxAf5_0;
	wire w_dff_A_NuwZW70N1_0;
	wire w_dff_A_93rcbJ8W5_0;
	wire w_dff_A_LFMcXJ298_0;
	wire w_dff_A_OA0AK7At2_0;
	wire w_dff_A_iA5EtpUZ7_0;
	wire w_dff_A_HcqOZvGd0_0;
	wire w_dff_A_IHhhvd3w7_0;
	wire w_dff_A_aZL3SwJX9_0;
	wire w_dff_A_f94wbbgQ4_0;
	wire w_dff_A_88dYPDEu9_2;
	wire w_dff_A_yIsJvCgR8_2;
	wire w_dff_A_i2oHWcU87_2;
	wire w_dff_A_00MZFfXb4_2;
	wire w_dff_A_LJ05JdEi1_2;
	wire w_dff_A_nEs3OTwA1_2;
	wire w_dff_A_sefpTJnz7_2;
	wire w_dff_A_rSzX3Gc14_2;
	wire w_dff_A_3xtNxIFQ1_2;
	wire w_dff_A_9Nfi2wJt9_2;
	wire w_dff_A_fIgYN3Ul8_2;
	wire w_dff_A_urRTYDO26_2;
	wire w_dff_A_xf66lUCa1_2;
	wire w_dff_A_OxNUh6XI1_2;
	wire w_dff_A_O0lssmRo2_2;
	wire w_dff_A_Z9sIK7Ul3_2;
	wire w_dff_A_L7UmcHcD4_2;
	wire w_dff_A_QtV3GtD43_2;
	wire w_dff_A_MIOownFJ9_0;
	wire w_dff_A_1MSLH93I7_0;
	wire w_dff_A_CauE5RpT8_0;
	wire w_dff_A_yMnJDmyu7_0;
	wire w_dff_A_nL85My2h9_0;
	wire w_dff_A_BgO5cR615_0;
	wire w_dff_A_DYNBgs530_0;
	wire w_dff_A_rLHIpSQp7_0;
	wire w_dff_A_rSC5yAMZ6_0;
	wire w_dff_A_m5ONKO6z3_0;
	wire w_dff_A_TTPrAq6q7_0;
	wire w_dff_A_nOXqYiFV2_0;
	wire w_dff_A_1gwjD4y12_0;
	wire w_dff_B_Dv6mIgGh6_2;
	wire w_dff_B_SdFwrvQ83_2;
	wire w_dff_B_EIYVk1i47_2;
	wire w_dff_B_GjqMQ1wZ2_1;
	wire w_dff_B_9It1tp8z4_0;
	wire w_dff_B_6yWgKtOw7_0;
	wire w_dff_B_7qWwFGV17_0;
	wire w_dff_A_24pca0HV7_0;
	wire w_dff_B_9v0UvJns1_1;
	wire w_dff_A_tO90tMmr9_0;
	wire w_dff_B_zK5lCcxZ2_1;
	wire w_dff_B_bZ2YK1Iu4_1;
	wire w_dff_B_IrMKE7qT9_1;
	wire w_dff_B_fsiWhS0U1_1;
	wire w_dff_B_u60iEu935_0;
	wire w_dff_B_ZpFDWVFP4_1;
	wire w_dff_B_XwVNHKM36_0;
	wire w_dff_A_5m1sBFBP3_0;
	wire w_dff_A_2gEbBQhW3_0;
	wire w_dff_A_5sB5Qmdb9_0;
	wire w_dff_A_1raUQNaH4_0;
	wire w_dff_B_WwIkTV058_0;
	wire w_dff_A_X2w1lQ6U1_0;
	wire w_dff_B_5gaPbxNb7_0;
	wire w_dff_B_LZUjBD4E1_0;
	wire w_dff_B_iHCHDIPS1_0;
	wire w_dff_B_f6Ui00f27_0;
	wire w_dff_B_jAc165sS2_0;
	wire w_dff_B_smLObfyz5_0;
	wire w_dff_B_Werem8sL7_0;
	wire w_dff_B_49EIEMAo1_0;
	wire w_dff_B_0mHTzpry5_0;
	wire w_dff_B_NqxXKWV73_0;
	wire w_dff_B_WBZdrwGk0_0;
	wire w_dff_B_J9pkYxVq4_0;
	wire w_dff_B_CWM73GqH0_0;
	wire w_dff_B_VYpWjlrd2_0;
	wire w_dff_B_nwXDeyvS8_0;
	wire w_dff_B_dTt7e69l8_0;
	wire w_dff_B_foFSaU8A0_0;
	wire w_dff_B_WQeYJm0f2_0;
	wire w_dff_B_neDWcCt91_0;
	wire w_dff_B_9PRc625b3_0;
	wire w_dff_B_fBhAPvB28_0;
	wire w_dff_B_LSRApeyK8_0;
	wire w_dff_B_p8y7SmDH3_0;
	wire w_dff_B_IIjg4NL32_0;
	wire w_dff_B_pgMHeisA8_0;
	wire w_dff_B_tc7Bs2wn5_0;
	wire w_dff_B_IauBRnPd9_0;
	wire w_dff_B_YsrTa2460_0;
	wire w_dff_B_vojdUPDY4_0;
	wire w_dff_B_g0jx4bv50_0;
	wire w_dff_B_Zt4fGQ628_0;
	wire w_dff_B_IJ7dlnse4_0;
	wire w_dff_B_tFx1AYRP1_0;
	wire w_dff_B_Bb1YNwW11_0;
	wire w_dff_B_ZNrBUawd7_0;
	wire w_dff_B_8rv1HNPK0_0;
	wire w_dff_B_VJUTrNHT7_2;
	wire w_dff_B_BL3JyIJS4_2;
	wire w_dff_B_LlnZ7Dqk4_2;
	wire w_dff_B_2jIm1a6Y6_0;
	wire w_dff_B_4eHGq9aF2_0;
	wire w_dff_B_Obs0PbIK9_0;
	wire w_dff_B_HU9STO0D6_0;
	wire w_dff_B_BOUBNzSk6_0;
	wire w_dff_B_GawIDrEg5_0;
	wire w_dff_B_bK1DZHkL5_0;
	wire w_dff_B_gdrQ4hA06_0;
	wire w_dff_B_C46Yp5rT9_0;
	wire w_dff_B_RsQmhCZC4_0;
	wire w_dff_B_WRs12aCC1_0;
	wire w_dff_B_2FPcrCAD0_0;
	wire w_dff_B_iLdb7h6h5_0;
	wire w_dff_B_JS5YIbSr7_0;
	wire w_dff_B_Alg2lQr27_0;
	wire w_dff_B_bexrAVvW0_0;
	wire w_dff_B_Wf1pMfSH9_0;
	wire w_dff_B_3GoT8bjo8_0;
	wire w_dff_B_3oHSvQGF6_0;
	wire w_dff_B_2dd9hNeQ1_0;
	wire w_dff_B_FdpjtFuW3_0;
	wire w_dff_B_w3V5Omow0_0;
	wire w_dff_B_bINVdSBt0_0;
	wire w_dff_B_aunuScad6_0;
	wire w_dff_B_y5HChuQV8_0;
	wire w_dff_B_EuoWpmdw5_0;
	wire w_dff_B_lOIOp8TB2_0;
	wire w_dff_B_QTrQBzim1_0;
	wire w_dff_B_51ll5nqO0_0;
	wire w_dff_B_rtGJoXJ30_0;
	wire w_dff_B_ShkG2wNF7_0;
	wire w_dff_B_4lzrQbwA2_0;
	wire w_dff_B_gAKDul2C1_0;
	wire w_dff_B_leJxw7Py9_0;
	wire w_dff_A_sFWHDYan7_2;
	wire w_dff_A_pjgPQuD18_2;
	wire w_dff_B_20x9tGxk2_0;
	wire w_dff_B_y6yL2sl84_0;
	wire w_dff_B_8QSHNWlh4_0;
	wire w_dff_B_K9XhQCve7_0;
	wire w_dff_B_JVr4qkUt1_0;
	wire w_dff_B_4iGO9YDx5_0;
	wire w_dff_B_ADhVyGKw3_0;
	wire w_dff_B_4U7IAqCH5_0;
	wire w_dff_B_GcBshYe89_0;
	wire w_dff_B_QuHuM2o98_0;
	wire w_dff_B_jvQLPQR05_0;
	wire w_dff_B_DBQzuKY78_0;
	wire w_dff_B_KUzCtUsv5_0;
	wire w_dff_B_HAZEoKtx6_0;
	wire w_dff_B_kbBNPsoE5_0;
	wire w_dff_B_8wzj2M7N8_0;
	wire w_dff_B_Sw2dCsV19_0;
	wire w_dff_B_UO6PmPVD3_0;
	wire w_dff_B_yhbITnzf3_0;
	wire w_dff_B_aZePPmIH4_0;
	wire w_dff_B_jrpvn6094_0;
	wire w_dff_B_GsUGTxeN9_0;
	wire w_dff_B_o94m2jSD3_0;
	wire w_dff_B_fk177KwR8_0;
	wire w_dff_B_kcVxM77C7_0;
	wire w_dff_B_kW3zZLNS6_0;
	wire w_dff_B_XGvfQ2Gc5_0;
	wire w_dff_B_R4JQJ6dt9_0;
	wire w_dff_B_WXwKa3HZ3_0;
	wire w_dff_B_L102BejT7_0;
	wire w_dff_B_zS322e1s8_0;
	wire w_dff_B_OeaKwgd32_0;
	wire w_dff_B_EykvKAbE6_0;
	wire w_dff_B_VMkJNZAT8_2;
	wire w_dff_B_id5mtwnl2_2;
	wire w_dff_B_CWb2MDZp4_2;
	wire w_dff_B_gl2MfgDg6_0;
	wire w_dff_B_By8RYdoW4_0;
	wire w_dff_B_kHZhQ3vZ7_0;
	wire w_dff_B_LywzKnL92_0;
	wire w_dff_B_BfgtXapc5_0;
	wire w_dff_B_TpSRZBrM4_0;
	wire w_dff_B_3zPE5ibu4_0;
	wire w_dff_B_RxqksCYE5_0;
	wire w_dff_B_PeCSNeRq8_0;
	wire w_dff_B_Wx5yXMqj3_0;
	wire w_dff_B_clMW8Zes3_0;
	wire w_dff_B_1cntyA2A5_0;
	wire w_dff_B_kF3Pzrva1_0;
	wire w_dff_B_Ijqvewyn4_0;
	wire w_dff_B_PCNzElJv1_0;
	wire w_dff_B_gqepe3so4_0;
	wire w_dff_B_TUIbUdjG8_0;
	wire w_dff_B_XnPH5e6I5_2;
	wire w_dff_B_U5rumXto4_2;
	wire w_dff_B_dCjbwhYg7_2;
	wire w_dff_A_SmbNmyt81_2;
	wire w_dff_A_Hz1qLP2O7_2;
	wire w_dff_B_p2Cx5lnN1_0;
	wire w_dff_B_cxMWjz5X1_0;
	wire w_dff_B_ASmHS2gG4_0;
	wire w_dff_B_Gr4XG9np8_0;
	wire w_dff_B_oTwodoID6_0;
	wire w_dff_B_Zmo8yTop6_0;
	wire w_dff_B_Vift5rqO8_0;
	wire w_dff_B_aMnyNwJM8_0;
	wire w_dff_B_EjvB9dRC0_0;
	wire w_dff_B_3XYKE3Vl7_0;
	wire w_dff_B_SxJqGZvK2_0;
	wire w_dff_B_DZXUIWvj3_0;
	wire w_dff_B_I3htXaNh3_0;
	wire w_dff_B_j5zEbwX24_0;
	wire w_dff_B_k1BaaJBX6_0;
	wire w_dff_B_O0tS13sh8_0;
	wire w_dff_B_Mo8eHblO3_2;
	wire w_dff_B_gjtDFMWi6_2;
	wire w_dff_B_el6Qlaq36_2;
	wire w_dff_B_YlXyAUM25_0;
	wire w_dff_B_aVj4Kkp72_0;
	wire w_dff_B_yq5DeBgq9_0;
	wire w_dff_B_sEJqdaGv0_0;
	wire w_dff_B_GLVIhucX2_0;
	wire w_dff_B_o72YPEzF5_0;
	wire w_dff_B_jw7iBpqr7_0;
	wire w_dff_B_NzQpgOY98_0;
	wire w_dff_B_De4INmgk8_0;
	wire w_dff_B_gXtEZGjE4_0;
	wire w_dff_B_eXUOmbkv6_0;
	wire w_dff_B_pc9SxJp39_0;
	wire w_dff_B_HVwaOk6v1_0;
	wire w_dff_B_FAtq4dTe0_0;
	wire w_dff_B_qH4ghL7g7_0;
	wire w_dff_B_ATcF3x672_0;
	wire w_dff_A_P1d707Og2_0;
	wire w_dff_A_i0nhRt9V4_0;
	wire w_dff_A_5z3ezwth3_0;
	wire w_dff_A_zyfe1BjJ8_0;
	wire w_dff_A_hwg82l3u4_0;
	wire w_dff_A_6cW6CQ4E5_1;
	wire w_dff_B_YNCVFuse0_0;
	wire w_dff_B_xN5Dk6JH0_0;
	wire w_dff_B_QgUyiywD0_0;
	wire w_dff_B_F0e6Rtjo2_0;
	wire w_dff_B_o1fgI3in6_0;
	wire w_dff_B_BEmcUTEZ6_0;
	wire w_dff_B_Ujy3i7h34_0;
	wire w_dff_B_VmXc9wwG0_0;
	wire w_dff_B_mY58C45M5_0;
	wire w_dff_B_ZOYtNVIT5_0;
	wire w_dff_B_op6k6ob95_0;
	wire w_dff_B_VD1RIM4u9_0;
	wire w_dff_B_K6oArLI90_0;
	wire w_dff_B_cxOX2idm5_0;
	wire w_dff_B_lSPkGAlU4_0;
	wire w_dff_B_M3NHt4gJ0_0;
	wire w_dff_B_QiyBP5GP1_0;
	wire w_dff_B_4msxmbml3_0;
	wire w_dff_B_zT7HkHPO6_0;
	wire w_dff_B_IRW2hMpD2_0;
	wire w_dff_B_LkrIOcYJ0_0;
	wire w_dff_B_aIZyJHXx4_0;
	wire w_dff_B_UhoOIOAq9_0;
	wire w_dff_B_ng5hXrky7_0;
	wire w_dff_B_TAghHFYQ5_0;
	wire w_dff_B_5ha3oELz4_0;
	wire w_dff_B_PlyUo6wp5_0;
	wire w_dff_B_yIo92Wkk0_0;
	wire w_dff_B_P2y9kksI0_0;
	wire w_dff_B_bOuWH4Eb6_0;
	wire w_dff_B_OdQbqyHw6_0;
	wire w_dff_B_t6jvK84v4_0;
	wire w_dff_B_3harrfKT3_0;
	wire w_dff_B_utLN8AQu0_0;
	wire w_dff_A_kniqA7ph3_0;
	wire w_dff_A_9abkvoqm3_1;
	wire w_dff_A_tC8auo9X0_0;
	wire w_dff_A_JLEfot5E1_1;
	wire w_dff_B_k8f7HUkw4_0;
	wire w_dff_B_XXqDlLwL6_0;
	wire w_dff_B_InhiICYY6_0;
	wire w_dff_B_reJt5BAK4_0;
	wire w_dff_B_2RNbhanw1_0;
	wire w_dff_B_5HpS8KsX8_0;
	wire w_dff_B_udvZJu4k1_0;
	wire w_dff_B_p9dWWpY59_0;
	wire w_dff_B_GJIH3AXz6_0;
	wire w_dff_B_HOEg0NhJ5_0;
	wire w_dff_B_pIsb6NzU4_0;
	wire w_dff_B_5VbBwoJ82_0;
	wire w_dff_B_lugxgPWM9_0;
	wire w_dff_B_U8AA5nKf2_0;
	wire w_dff_B_fAEC05d99_0;
	wire w_dff_B_AfURZYz12_0;
	wire w_dff_B_5tYYOmDO1_0;
	wire w_dff_B_GkzyK1x01_0;
	wire w_dff_A_a3Hw78NH0_0;
	wire w_dff_B_12U1LPE12_0;
	wire w_dff_B_KboSwyh90_0;
	wire w_dff_B_lkw6DABr2_0;
	wire w_dff_B_Ujyp9KRj3_0;
	wire w_dff_B_XYuEFKGi6_0;
	wire w_dff_B_2mBpvFFB1_0;
	wire w_dff_B_kiAnCau14_0;
	wire w_dff_B_gLUmyhuQ8_0;
	wire w_dff_B_vuir9hZV3_0;
	wire w_dff_B_iSZ1uR1d2_0;
	wire w_dff_B_Qdk5EYEE6_0;
	wire w_dff_B_Bzp7SjmF5_0;
	wire w_dff_B_iC0h8nva9_0;
	wire w_dff_B_bRY6WnYk0_0;
	wire w_dff_B_cvumRequ5_0;
	wire w_dff_B_MjGKjvwP7_0;
	wire w_dff_B_SurJZRrC4_2;
	wire w_dff_B_p7Wfqv4N3_2;
	wire w_dff_B_hcqlBw8G8_2;
	wire w_dff_B_w7B4ucgx9_0;
	wire w_dff_B_7VQL5rZ74_0;
	wire w_dff_B_S9c7Ccw26_0;
	wire w_dff_B_QNNNQo5B6_0;
	wire w_dff_B_GkqvVYFW1_0;
	wire w_dff_B_7gm4x91E5_0;
	wire w_dff_B_H2oYONkY2_0;
	wire w_dff_B_Ssvhphfd4_0;
	wire w_dff_B_Z8qSrzYS1_0;
	wire w_dff_B_q2OBw3WY3_0;
	wire w_dff_B_rFDNt3jY9_0;
	wire w_dff_B_bdJBNayM5_1;
	wire w_dff_B_ITDwAj4G9_1;
	wire w_dff_B_E8g3QzHa4_0;
	wire w_dff_B_lqrPEihh4_0;
	wire w_dff_B_jmxu1wD30_0;
	wire w_dff_B_TkLFjQNn8_0;
	wire w_dff_B_fc0m9S6j5_0;
	wire w_dff_B_Zki4KhR49_0;
	wire w_dff_B_HYYn7Udg2_0;
	wire w_dff_B_J2lMJmb59_0;
	wire w_dff_B_ixx83PVO8_0;
	wire w_dff_B_CoRr7QPr6_0;
	wire w_dff_B_WqfnwOen3_0;
	wire w_dff_B_D0xwtLV79_0;
	wire w_dff_B_LEUCKzil8_1;
	wire w_dff_B_cJA6FlcG8_1;
	wire w_dff_B_4nckjkxE7_0;
	wire w_dff_B_uOxuyozF6_1;
	wire w_dff_B_I4KrkMhc7_0;
	wire w_dff_B_HS4BqWTz7_0;
	wire w_dff_B_5akhSlJ55_0;
	wire w_dff_B_HMaARgkk1_0;
	wire w_dff_B_fT54kYaw2_0;
	wire w_dff_B_Tb9HEADJ3_0;
	wire w_dff_B_iCdtjdEr4_0;
	wire w_dff_B_aIP1Qrtr9_0;
	wire w_dff_B_xyU3yWxr2_0;
	wire w_dff_B_Bg74AEqj0_0;
	wire w_dff_B_PQ5jmQuJ6_0;
	wire w_dff_B_5r3plSjt2_0;
	wire w_dff_B_YHPm9qSs4_0;
	wire w_dff_B_ajDbJ6IJ9_0;
	wire w_dff_B_nOP5mOmz5_0;
	wire w_dff_B_7xflPzTx9_0;
	wire w_dff_B_Nh4RGfHi0_0;
	wire w_dff_B_HwkqESHD8_2;
	wire w_dff_B_I8wy6ybV9_2;
	wire w_dff_B_xpzfz9bn8_2;
	wire w_dff_B_pGEWszLa2_0;
	wire w_dff_B_70mbkrCG6_0;
	wire w_dff_B_82aZFgDR1_0;
	wire w_dff_B_l3VHYHKN3_0;
	wire w_dff_B_SqEKtrOP0_0;
	wire w_dff_B_vnhBaksL6_0;
	wire w_dff_B_I5EIZfyO6_0;
	wire w_dff_B_rjIdWvdH7_0;
	wire w_dff_B_YxpToVNN0_0;
	wire w_dff_B_brMOSBEK6_0;
	wire w_dff_B_lqayjOb33_0;
	wire w_dff_B_UWtMXrMa8_0;
	wire w_dff_B_EgurrhzS3_1;
	wire w_dff_B_qH7SRKVN3_1;
	wire w_dff_A_DNotvZS61_1;
	wire w_dff_B_0uH6sVWG8_1;
	wire w_dff_B_UuRwrD601_1;
	wire w_dff_B_zznk1NDg9_1;
	wire w_dff_B_6PAokJul5_1;
	wire w_dff_B_carxNRFb2_1;
	wire w_dff_B_Znrzi2Jp6_1;
	wire w_dff_B_TQCUVPUU7_1;
	wire w_dff_B_sAY3s7jv2_1;
	wire w_dff_B_OOTinskz4_1;
	wire w_dff_B_DrJsBLWi0_1;
	wire w_dff_B_knbxOmLs0_0;
	wire w_dff_B_VFdQSXig9_0;
	wire w_dff_B_u7GkHHnL4_0;
	wire w_dff_B_cjLvs0lE2_0;
	wire w_dff_B_wh4YQLXe2_0;
	wire w_dff_B_XIHeVgmt9_0;
	wire w_dff_B_gGeo0y4J5_0;
	wire w_dff_B_QCmH1uUZ1_0;
	wire w_dff_B_UbmoN6sJ0_0;
	wire w_dff_B_YMzSjBaa5_0;
	wire w_dff_B_N1JcnImR0_0;
	wire w_dff_B_4sIPjaQH0_0;
	wire w_dff_B_cTovec442_0;
	wire w_dff_B_h4nnryEP7_1;
	wire w_dff_B_pPteiRlH7_1;
	wire w_dff_B_5azsRgP08_0;
	wire w_dff_B_8ngaOgZp0_1;
	wire w_dff_B_ghmy57IS4_1;
	wire w_dff_B_ulSZtaFu8_1;
	wire w_dff_B_6IZ25oof1_1;
	wire w_dff_B_rqgEC4XS4_1;
	wire w_dff_B_qrbp3l5i8_1;
	wire w_dff_B_Z5TGiR6n4_1;
	wire w_dff_B_X8We1c0a4_1;
	wire w_dff_B_x7A8Np4n0_1;
	wire w_dff_B_UDifye6W0_1;
	wire w_dff_B_VGJ83NmS9_1;
	wire w_dff_B_nsf7sUfc3_1;
	wire w_dff_B_Ui9iQyjd0_1;
	wire w_dff_B_2jmTBkcx4_1;
	wire w_dff_B_Q7f9PXUA6_1;
	wire w_dff_B_ZQO9pmoP6_1;
	wire w_dff_B_5Ot26uPJ7_1;
	wire w_dff_B_6ZwNLYnp6_1;
	wire w_dff_B_7J51VwjJ9_1;
	wire w_dff_B_JasYwprn6_1;
	wire w_dff_A_eTIhmptp4_1;
	wire w_dff_A_0ABgA4ZH5_1;
	wire w_dff_A_nWwNMmAl9_1;
	wire w_dff_A_e5sfyIm04_1;
	wire w_dff_A_WmOrV3Fc7_1;
	wire w_dff_A_TxbQkaMK3_1;
	wire w_dff_A_pUdYOU2L4_1;
	wire w_dff_A_fT9ePtr77_1;
	wire w_dff_A_uLpVJ25x2_1;
	wire w_dff_A_fGyFZUvc5_1;
	wire w_dff_A_59LsnX7Q3_1;
	wire w_dff_A_018LXOWc5_1;
	wire w_dff_A_pVTYFNtE9_1;
	wire w_dff_A_eTYBwnWT9_2;
	wire w_dff_A_Nsw36ZaJ8_2;
	wire w_dff_A_srXh94j66_2;
	wire w_dff_A_iOykxtBa3_2;
	wire w_dff_A_r0gtHvQl2_2;
	wire w_dff_A_5Oo6AbkR6_2;
	wire w_dff_A_1HpV4mEj0_2;
	wire w_dff_A_mJ6drfkE6_2;
	wire w_dff_A_dkLkqm3k4_2;
	wire w_dff_A_xnxpTREI0_2;
	wire w_dff_A_1Go8PI2h1_2;
	wire w_dff_A_38LaT17l8_2;
	wire w_dff_B_AZprxqzJ0_0;
	wire w_dff_B_mJ1j1gTD0_0;
	wire w_dff_B_7HZIShAY0_0;
	wire w_dff_B_n1wrDYVY5_0;
	wire w_dff_B_1RR1CZsP4_0;
	wire w_dff_B_tfpD0Udf2_0;
	wire w_dff_B_vSj85tUk1_0;
	wire w_dff_B_pVt6E6em8_0;
	wire w_dff_B_7zjMzTiS5_0;
	wire w_dff_B_oScitRmT1_0;
	wire w_dff_B_yFm1JmTH9_0;
	wire w_dff_B_2dJWhgjF7_0;
	wire w_dff_B_qLHmevy57_0;
	wire w_dff_B_TuGE8FT87_0;
	wire w_dff_B_tKJwDoLf8_0;
	wire w_dff_B_r8jmrCwB8_0;
	wire w_dff_B_b4LZq0Iw7_0;
	wire w_dff_B_8Rzw76ML0_2;
	wire w_dff_B_UxgFEG5G5_2;
	wire w_dff_B_kg6O6kvQ3_2;
	wire w_dff_B_BzXtCudD3_0;
	wire w_dff_B_64ZAyU2B5_0;
	wire w_dff_B_1yU9SCky0_0;
	wire w_dff_B_eeKeqSw40_0;
	wire w_dff_B_g1Qpje6Z1_0;
	wire w_dff_B_tzWsAc6R7_0;
	wire w_dff_B_ytQDl9nC8_0;
	wire w_dff_B_Myw9mLdh9_0;
	wire w_dff_B_8XhrK0Hx5_0;
	wire w_dff_B_cJFTjYXl4_0;
	wire w_dff_B_5EJPR0oB7_0;
	wire w_dff_B_e3bAn2re2_0;
	wire w_dff_B_CUFbrsfo3_1;
	wire w_dff_B_qIHigijf7_1;
	wire w_dff_A_zHdw3oJE0_0;
	wire w_dff_A_AFXfzUH98_0;
	wire w_dff_A_Uhkbv8Pc0_0;
	wire w_dff_A_xIckdFqs7_0;
	wire w_dff_A_oaUSor5k9_2;
	wire w_dff_A_6f8Kk6ui9_2;
	wire w_dff_A_hm8qYiz91_1;
	wire w_dff_A_w7FT3ZHn7_1;
	wire w_dff_A_vZuh13DQ2_1;
	wire w_dff_A_GSd6Hx7u4_1;
	wire w_dff_A_tA1UrYIt4_1;
	wire w_dff_A_bHU8Cxld7_1;
	wire w_dff_A_MDJfGGFF6_1;
	wire w_dff_A_UfZ86a0w8_1;
	wire w_dff_A_iUdpGVFf1_2;
	wire w_dff_A_SRHHe0ma6_2;
	wire w_dff_A_DGzWvVuZ2_2;
	wire w_dff_A_N4ptuOW26_2;
	wire w_dff_B_ihQVpXUD7_3;
	wire w_dff_A_RVWRKP4u1_0;
	wire w_dff_A_UsOp91Lb7_0;
	wire w_dff_A_J08NF0FU0_0;
	wire w_dff_A_2BCbV1iz5_0;
	wire w_dff_A_Iy73Tv2g0_0;
	wire w_dff_A_MOpsaM2X7_0;
	wire w_dff_A_v7q9nTJl1_0;
	wire w_dff_A_COGThtqU9_0;
	wire w_dff_A_pFbXiNEm7_1;
	wire w_dff_A_eKidrWQg0_1;
	wire w_dff_A_mE9sZeDh0_1;
	wire w_dff_A_rcHSEw7v8_0;
	wire w_dff_A_BDAlbrwS2_1;
	wire w_dff_B_CQd7OXAe5_0;
	wire w_dff_B_5QXWSjRb3_0;
	wire w_dff_B_R7dNp7hJ7_0;
	wire w_dff_B_n3xBIV976_0;
	wire w_dff_B_LIfP6j794_0;
	wire w_dff_B_BpP2UyFK0_0;
	wire w_dff_B_nKDMICHL9_0;
	wire w_dff_B_dT3YUtLv0_0;
	wire w_dff_B_xDE9Jiw79_0;
	wire w_dff_B_9aBtAWWI9_0;
	wire w_dff_B_pRA1cafs6_0;
	wire w_dff_B_ZvN6PyDk5_0;
	wire w_dff_B_8vNbqRXJ6_0;
	wire w_dff_B_eHQunb1k9_1;
	wire w_dff_B_evsv9m3f0_1;
	wire w_dff_B_AlfhYG632_3;
	wire w_dff_B_zVEI9lAu4_3;
	wire w_dff_A_wIJmSegh5_1;
	wire w_dff_B_Lm8hocjk6_0;
	wire w_dff_B_r7DXClUe9_3;
	wire w_dff_B_3iQ4hjCX7_1;
	wire w_dff_A_CohO1dF46_0;
	wire w_dff_A_pvudMBQF0_1;
	wire w_dff_A_eo9C9SN44_0;
	wire w_dff_A_nd61yT9j0_1;
	wire w_dff_A_el7JVLJ86_0;
	wire w_dff_A_OSLWcwJ35_0;
	wire w_dff_A_Cs21iRWK2_0;
	wire w_dff_A_GF7DKR0k2_0;
	wire w_dff_A_bi3X8rNv0_0;
	wire w_dff_A_46Zjjtm19_1;
	wire w_dff_A_2wQNXJ733_1;
	wire w_dff_A_ll5qnhqY0_1;
	wire w_dff_A_thSmdNK93_1;
	wire w_dff_A_cblSsHYI7_1;
	wire w_dff_A_ooNgcASa8_1;
	wire w_dff_B_almq03eI8_0;
	wire w_dff_B_IRLgO7kt4_0;
	wire w_dff_B_Blybwakb8_0;
	wire w_dff_B_0RFEi9ci0_0;
	wire w_dff_B_MeIY2g1J9_0;
	wire w_dff_B_wirLnp5Y7_0;
	wire w_dff_B_sZFEaVQg0_0;
	wire w_dff_B_NMbhQSno3_0;
	wire w_dff_B_f1WBGkjH6_0;
	wire w_dff_B_r142rHGR1_0;
	wire w_dff_B_QXlYfsDA3_0;
	wire w_dff_B_qINY983G6_0;
	wire w_dff_B_ITqUOcel1_0;
	wire w_dff_B_wjxWFONT5_0;
	wire w_dff_B_t7Yetd7S2_0;
	wire w_dff_B_Rly3K5lm9_0;
	wire w_dff_B_Cz04OjIr1_0;
	wire w_dff_B_vnyIMFO61_0;
	wire w_dff_B_FiyemRXA2_2;
	wire w_dff_B_px3atMtj6_2;
	wire w_dff_B_PNYWUf4z8_2;
	wire w_dff_B_IT0FyqTn8_0;
	wire w_dff_B_aYFo1R831_0;
	wire w_dff_B_9oEZ1EmU6_0;
	wire w_dff_B_oGgbRWhq1_0;
	wire w_dff_B_5vOD4vSr4_0;
	wire w_dff_B_RuDVHECz3_0;
	wire w_dff_B_J1fDPc8v1_0;
	wire w_dff_B_DnvMvUNs7_0;
	wire w_dff_B_8QCisCFT2_0;
	wire w_dff_B_ntq2q3TZ1_0;
	wire w_dff_B_YsrSnTeg1_0;
	wire w_dff_B_QLeuCNyl6_0;
	wire w_dff_B_dJTTVpsB3_0;
	wire w_dff_B_cF4ZbbJB2_1;
	wire w_dff_B_WSVXGEBq2_1;
	wire w_dff_A_3ZPaxM2o1_1;
	wire w_dff_A_knKS0aNM9_0;
	wire w_dff_B_YztjzzMN1_2;
	wire w_dff_B_gcIRcr813_0;
	wire w_dff_B_GVlAryBp3_0;
	wire w_dff_B_GUlMS4gv6_0;
	wire w_dff_B_3RXYZWmb0_0;
	wire w_dff_A_ux3c2iUQ5_0;
	wire w_dff_A_xHdeIjsH5_0;
	wire w_dff_A_Ptqp5SJG7_0;
	wire w_dff_A_NWYkjshc5_0;
	wire w_dff_A_SjLtKWoS8_0;
	wire w_dff_A_7xOfXmXs0_0;
	wire w_dff_A_25C853gH3_0;
	wire w_dff_A_arY8dTIP6_0;
	wire w_dff_A_dMhfcUjY7_0;
	wire w_dff_A_PvX7XXFv4_0;
	wire w_dff_A_DiOMKzrL1_0;
	wire w_dff_A_OuHO2q7r5_0;
	wire w_dff_A_K7AyFFeR1_0;
	wire w_dff_A_dwYZuPoa4_0;
	wire w_dff_A_S50wsJSu9_0;
	wire w_dff_A_7ZMgPdB88_0;
	wire w_dff_A_uFZ7ilqp2_0;
	wire w_dff_A_xoQKAynq0_0;
	wire w_dff_A_WZJHD5gS9_0;
	wire w_dff_A_NrSQtPIH1_0;
	wire w_dff_A_B3mCpQCe6_1;
	wire w_dff_A_oBdeOxA45_1;
	wire w_dff_A_zkzI0MoW7_1;
	wire w_dff_A_jSgBYgoR4_1;
	wire w_dff_A_FBWiu6sb3_1;
	wire w_dff_A_LYNo2ASk7_1;
	wire w_dff_A_ACD1nKsc4_1;
	wire w_dff_A_GAKN05Nq0_1;
	wire w_dff_A_46KeFG3T5_1;
	wire w_dff_B_mqZHnNjT7_0;
	wire w_dff_B_zVHJlvIO3_0;
	wire w_dff_B_xUFYXKgH2_0;
	wire w_dff_B_XUtwgCBg4_0;
	wire w_dff_B_l6lm0sY73_0;
	wire w_dff_B_iuwMfApg1_0;
	wire w_dff_B_huMTkWf36_0;
	wire w_dff_B_jhuFUAdV5_0;
	wire w_dff_B_KOlIZRFo4_0;
	wire w_dff_B_D592iDCk4_0;
	wire w_dff_B_zqJOUQM15_0;
	wire w_dff_B_2XMIVhUw3_0;
	wire w_dff_B_kfM8BBMH2_0;
	wire w_dff_B_rRV3MrUo5_0;
	wire w_dff_B_xtfFS7ya0_0;
	wire w_dff_B_KwgV3T4n3_0;
	wire w_dff_B_RQTw2CmT4_1;
	wire w_dff_B_CjpD4YzR1_1;
	wire w_dff_A_b3F2XRIP3_0;
	wire w_dff_A_i2MhnlsV3_2;
	wire w_dff_A_SswdMDB54_2;
	wire w_dff_A_wqPfTT917_2;
	wire w_dff_A_uIcXy7Ld2_2;
	wire w_dff_B_KmBIXJZD9_1;
	wire w_dff_B_vABTjAim3_1;
	wire w_dff_B_lE0fHd272_1;
	wire w_dff_B_mG22AAd94_1;
	wire w_dff_B_sHr3FexY7_1;
	wire w_dff_B_ZC0Suado3_1;
	wire w_dff_B_1MX1hrpz6_1;
	wire w_dff_B_n8WOJk9M0_1;
	wire w_dff_B_gcQBnGqx9_1;
	wire w_dff_B_5BahILlN4_1;
	wire w_dff_B_0DZi2YVH6_1;
	wire w_dff_B_eG2B8B5I5_1;
	wire w_dff_B_X582oZyd9_1;
	wire w_dff_B_P2Tlkxjg6_1;
	wire w_dff_B_tXbYhoQQ6_1;
	wire w_dff_B_VezKcuRz7_1;
	wire w_dff_B_VH3KISCb2_1;
	wire w_dff_B_Apat5Bi87_1;
	wire w_dff_B_NtUiBiVq2_0;
	wire w_dff_A_2Sfp7Nqg3_1;
	wire w_dff_A_5jwWtI1F4_1;
	wire w_dff_A_yDS8hk1Y9_1;
	wire w_dff_A_W9Ozmo8a0_1;
	wire w_dff_A_lYjkwI1V6_1;
	wire w_dff_A_9Gi1pbWn9_1;
	wire w_dff_B_g3IckT5T9_3;
	wire w_dff_B_4eX0Co9w0_3;
	wire w_dff_B_2CffgmCk6_3;
	wire w_dff_B_K8ORnOKd0_3;
	wire w_dff_B_DAKqQrDa0_2;
	wire w_dff_B_LuVljHUT6_2;
	wire w_dff_B_Ppqaer007_2;
	wire w_dff_B_gNUNXADe4_2;
	wire w_dff_B_ricpX7Rv7_2;
	wire w_dff_B_ugLXr8VB4_2;
	wire w_dff_B_gknoEShI4_2;
	wire w_dff_B_RFcK7kxy9_2;
	wire w_dff_B_yjprOUEj0_2;
	wire w_dff_A_SgNHVH5Z3_1;
	wire w_dff_A_iFVfDNt66_1;
	wire w_dff_A_vsXEra7e3_1;
	wire w_dff_A_W2DtHLXz9_2;
	wire w_dff_A_pvl3mcel0_2;
	wire w_dff_A_03Umby7w5_2;
	wire w_dff_A_iT9fQLBz5_2;
	wire w_dff_A_v34TugCi6_0;
	wire w_dff_A_mBnxGzrR9_0;
	wire w_dff_A_CSeudXrA7_0;
	wire w_dff_A_thU9StEt9_0;
	wire w_dff_A_gIZTJ2SD4_0;
	wire w_dff_A_4GamQ0Jp2_0;
	wire w_dff_A_hvvYB3n21_0;
	wire w_dff_A_TWQEc8XZ8_0;
	wire w_dff_A_pczc4ae96_0;
	wire w_dff_A_BmndQNu78_0;
	wire w_dff_A_vPbLhE3F2_0;
	wire w_dff_A_75gcu1mL0_0;
	wire w_dff_A_4H65fA2y3_0;
	wire w_dff_A_sJR2gL3C3_1;
	wire w_dff_A_CgSBUOBR4_1;
	wire w_dff_A_YtMPeKmw1_1;
	wire w_dff_A_PNQ1jMf32_1;
	wire w_dff_A_lWU3J0Ge3_1;
	wire w_dff_A_evCurInq7_1;
	wire w_dff_A_gZRPnmG56_1;
	wire w_dff_B_5RGa8LMP9_1;
	wire w_dff_B_HxLhjqH88_1;
	wire w_dff_B_74sPFeaY7_1;
	wire w_dff_B_27JaNkQl8_1;
	wire w_dff_B_8oTVzDsz9_1;
	wire w_dff_B_YGBlsYku1_1;
	wire w_dff_B_uxi4rQSK1_1;
	wire w_dff_B_TBbHLIV76_1;
	wire w_dff_B_Uvt2fEHQ9_1;
	wire w_dff_B_Hmj92KV31_1;
	wire w_dff_B_ax4oRnWb1_1;
	wire w_dff_B_gGG5PQ2J1_1;
	wire w_dff_B_q2KJSj7E7_1;
	wire w_dff_B_NCck7nZb0_1;
	wire w_dff_B_rW0Q9rgF2_1;
	wire w_dff_B_aHHJLOyA5_1;
	wire w_dff_B_uazdRGXM7_1;
	wire w_dff_B_zOwdtIAm3_1;
	wire w_dff_B_jxny4ArA6_1;
	wire w_dff_B_qGfkV9Ns6_1;
	wire w_dff_B_eGcvvx9E1_1;
	wire w_dff_B_4f5py8GE0_1;
	wire w_dff_B_S69VBAbw0_1;
	wire w_dff_B_2qZ4r7xt4_1;
	wire w_dff_B_wHqDGhkw3_1;
	wire w_dff_B_gdxU8hfz6_1;
	wire w_dff_B_t2cExOin3_1;
	wire w_dff_B_gMbUnIvW5_1;
	wire w_dff_B_7BMQW0dG5_1;
	wire w_dff_B_5tJKBy3B1_1;
	wire w_dff_B_Hwg6UBlW5_1;
	wire w_dff_B_8dbasd5t4_1;
	wire w_dff_B_FStOYtq33_1;
	wire w_dff_B_vYN0ROCC7_1;
	wire w_dff_B_UR5UkB7Z1_1;
	wire w_dff_B_crLcOZlU7_1;
	wire w_dff_B_OU4yaq7L3_1;
	wire w_dff_B_nIpOyoey8_1;
	wire w_dff_B_fRM4cHqM2_0;
	wire w_dff_B_kitt4geg0_0;
	wire w_dff_B_liwupeu76_0;
	wire w_dff_B_bvWzRpva7_0;
	wire w_dff_B_kbArhJW13_0;
	wire w_dff_B_liTFATlW4_0;
	wire w_dff_B_Kj340Lus6_0;
	wire w_dff_B_1fzNq9SA6_0;
	wire w_dff_B_GbUkwzVG5_0;
	wire w_dff_B_IIaOuqWc4_0;
	wire w_dff_B_MC0H8Sk78_0;
	wire w_dff_B_UqiGo2xb0_0;
	wire w_dff_B_h8W123E12_0;
	wire w_dff_B_vpAbq5Po0_0;
	wire w_dff_B_dK9GxTrQ6_0;
	wire w_dff_B_P8zjaeIw7_0;
	wire w_dff_B_lZI4WODN9_0;
	wire w_dff_B_I5IH0MMJ2_0;
	wire w_dff_B_4rHYBAdE5_0;
	wire w_dff_B_h1ssQCLb9_0;
	wire w_dff_A_62QowrCK3_1;
	wire w_dff_A_44HAr5Qh2_1;
	wire w_dff_A_4j65zlAi8_1;
	wire w_dff_A_e1fNy4Ma2_1;
	wire w_dff_A_kBPdLRwq7_1;
	wire w_dff_A_dwd6FNwR2_1;
	wire w_dff_A_4ZMbzVX56_1;
	wire w_dff_A_cKUj5x8V8_1;
	wire w_dff_A_LzInWdmJ3_1;
	wire w_dff_A_s6I1a9Su3_1;
	wire w_dff_A_sOa87aUo4_1;
	wire w_dff_A_oNDKrWIW1_1;
	wire w_dff_A_3gVy0WKl4_1;
	wire w_dff_A_1PVE3DRf5_1;
	wire w_dff_A_ZBIsONhY0_2;
	wire w_dff_A_LSJWrf1e7_2;
	wire w_dff_A_P1hkd3J18_2;
	wire w_dff_A_Vrm60Fkm3_2;
	wire w_dff_A_64DEMkZ58_2;
	wire w_dff_A_1bZSorDu6_2;
	wire w_dff_A_JUoG50SJ8_2;
	wire w_dff_A_7praynRV6_2;
	wire w_dff_A_7CIQBXyA2_2;
	wire w_dff_A_hL4526bv5_2;
	wire w_dff_A_qAJnDHiJ4_1;
	wire w_dff_A_K9DS2KSS3_1;
	wire w_dff_A_qlCUkixp0_1;
	wire w_dff_A_VFR3Wbyt5_1;
	wire w_dff_A_mroUqqRB1_1;
	wire w_dff_A_KglxCDra0_1;
	wire w_dff_A_O26fNIRH7_1;
	wire w_dff_A_IPQ2NA3F8_1;
	wire w_dff_A_4JxQ5gnA4_1;
	wire w_dff_A_r2w5kEW48_1;
	wire w_dff_A_vufs09fJ5_1;
	wire w_dff_A_V3S91piA1_2;
	wire w_dff_B_zVz0njuI9_3;
	wire w_dff_B_853ihHdN7_3;
	wire w_dff_B_l2KaA5Gl2_3;
	wire w_dff_B_9YBJuyUI5_3;
	wire w_dff_B_JRRagGoi5_3;
	wire w_dff_B_p44IFa8m3_3;
	wire w_dff_A_kio7HzqD0_1;
	wire w_dff_A_89JhneNF5_1;
	wire w_dff_A_oxxJBvXz8_1;
	wire w_dff_A_V93YUqWD9_1;
	wire w_dff_A_Cgt4QIfM0_1;
	wire w_dff_A_9AN431Ud5_1;
	wire w_dff_A_IMcBrGU46_1;
	wire w_dff_A_waABEiXy6_1;
	wire w_dff_A_23tbKixm2_1;
	wire w_dff_A_vIgoic5m5_1;
	wire w_dff_A_sazGto2U8_1;
	wire w_dff_A_shYT65ez1_1;
	wire w_dff_A_RKl2ve8Q2_1;
	wire w_dff_A_wYf4CRIS1_1;
	wire w_dff_A_UVlzuZWb8_2;
	wire w_dff_A_QzRlgLRO8_2;
	wire w_dff_A_yzc1uo0F6_2;
	wire w_dff_A_eEqAMYCR9_2;
	wire w_dff_A_XYjok7qO5_2;
	wire w_dff_A_y9yAjSAU3_2;
	wire w_dff_A_PGi66FSw6_2;
	wire w_dff_A_isx0Vjju4_2;
	wire w_dff_A_SVYFXeQF0_2;
	wire w_dff_A_0Wy3drpl8_2;
	wire w_dff_A_jkVu3gCc7_1;
	wire w_dff_A_M74dmBav1_1;
	wire w_dff_A_KelRrALB2_1;
	wire w_dff_A_PwFCSI5r0_1;
	wire w_dff_A_V2Y6lBwb6_1;
	wire w_dff_A_8JskB42r8_1;
	wire w_dff_A_kTF9EuCu8_1;
	wire w_dff_A_SYAEVGV86_1;
	wire w_dff_A_KbIqXLc50_1;
	wire w_dff_A_J17m2agI0_1;
	wire w_dff_A_dYGaO07l1_1;
	wire w_dff_A_j69jbkpN2_2;
	wire w_dff_A_HyK6inpt4_2;
	wire w_dff_A_5PWCTDXZ9_2;
	wire w_dff_A_AeEiZwLg7_2;
	wire w_dff_B_Vz2IWRYo0_3;
	wire w_dff_B_lKYooOn52_3;
	wire w_dff_B_7Y5UojCy3_3;
	wire w_dff_B_Ki2i9Lgb6_3;
	wire w_dff_B_LsMfgfUp1_3;
	wire w_dff_B_QcBZguBB0_3;
	wire w_dff_B_yK95vB9c5_3;
	wire w_dff_A_tXtXJkyC4_2;
	wire w_dff_A_bHB1uaTW0_1;
	wire w_dff_B_R330pzjb9_0;
	wire w_dff_B_416ZNeiT5_0;
	wire w_dff_B_qHzkM02Y0_0;
	wire w_dff_B_UK0QYkxR1_0;
	wire w_dff_B_oMITCUFG6_0;
	wire w_dff_B_a5esy9Ro8_0;
	wire w_dff_B_dldAmf1U9_0;
	wire w_dff_B_HU89f4DN3_0;
	wire w_dff_B_w8mBglBD0_0;
	wire w_dff_B_vZIkUZa78_0;
	wire w_dff_B_C30ova2w0_0;
	wire w_dff_B_lpjfJTRG5_0;
	wire w_dff_B_eNMxXgBn3_0;
	wire w_dff_B_XCIH7Gjk7_0;
	wire w_dff_B_5GKH6wMV0_0;
	wire w_dff_B_E4TLQkV22_0;
	wire w_dff_B_8PIr0QJx3_0;
	wire w_dff_B_2UCQuvcd7_0;
	wire w_dff_B_8D5LGT767_0;
	wire w_dff_B_RTVcvQFq5_0;
	wire w_dff_B_J9TBYGZH4_2;
	wire w_dff_B_nFTGIpDI1_2;
	wire w_dff_B_CaICsnEX1_2;
	wire w_dff_A_PGw1EWcz1_1;
	wire w_dff_A_cq3UHFCW8_1;
	wire w_dff_A_PVEWL3WN6_1;
	wire w_dff_A_eiIao9IU9_1;
	wire w_dff_A_TU0tkgSz0_1;
	wire w_dff_A_uOmx0oVi4_1;
	wire w_dff_A_KKUldiPv3_1;
	wire w_dff_A_vqAPTctO8_1;
	wire w_dff_A_07gJrxt32_1;
	wire w_dff_A_7lNkLDfZ5_1;
	wire w_dff_A_qjUNg49A8_1;
	wire w_dff_A_PAhiSHvw1_1;
	wire w_dff_A_tflyMCkZ3_1;
	wire w_dff_A_cLm3788F5_1;
	wire w_dff_A_XA3SDY189_2;
	wire w_dff_A_d5uhTrnv5_2;
	wire w_dff_A_PdeTCBKx7_2;
	wire w_dff_A_n41sYB646_2;
	wire w_dff_A_9Paqwd7y9_2;
	wire w_dff_A_YCzmOSG41_2;
	wire w_dff_A_GExw5Bi55_2;
	wire w_dff_A_IGyNVtjA3_2;
	wire w_dff_A_KVtIpd1a3_2;
	wire w_dff_A_e0Ih2LcX7_2;
	wire w_dff_A_zKvsHlYu4_1;
	wire w_dff_A_odlVhcBS1_1;
	wire w_dff_A_0sGSeRAR2_1;
	wire w_dff_A_VlmWAUTu7_1;
	wire w_dff_A_wTZE1LMp4_1;
	wire w_dff_A_jMtItFaU1_1;
	wire w_dff_A_7r37JUvU9_1;
	wire w_dff_A_PKjuOhSd0_1;
	wire w_dff_A_IaLfFmXh7_1;
	wire w_dff_A_47JVa2709_1;
	wire w_dff_A_EW7Rn3p67_1;
	wire w_dff_A_bYMz636x6_2;
	wire w_dff_B_wp8dM40r5_3;
	wire w_dff_B_tuhr30Vj1_3;
	wire w_dff_B_J8rV2HTe9_3;
	wire w_dff_B_rVkRGztn0_3;
	wire w_dff_B_i0e3EPfR9_3;
	wire w_dff_B_Yt0cDv956_3;
	wire w_dff_A_6al98zBo1_1;
	wire w_dff_A_KznqRwtA5_1;
	wire w_dff_A_iSVqMZcw6_1;
	wire w_dff_A_G4snWQlh7_1;
	wire w_dff_A_Hd6fwTqp3_1;
	wire w_dff_A_d5fkMHs96_1;
	wire w_dff_A_UvbRpELu2_1;
	wire w_dff_A_woVgbpwc3_1;
	wire w_dff_A_yuZPb1Ar7_1;
	wire w_dff_A_jJNAynl08_1;
	wire w_dff_A_j9d07eNU4_1;
	wire w_dff_A_M0bkpkk80_1;
	wire w_dff_A_1AGjTaxK9_1;
	wire w_dff_A_XrgxLxLA5_1;
	wire w_dff_A_YJYuMKOa9_2;
	wire w_dff_A_USTdVEhM2_2;
	wire w_dff_A_NZQwyrq54_2;
	wire w_dff_A_t7TaXIc05_2;
	wire w_dff_A_MGSQUssF7_2;
	wire w_dff_A_uYJht2rJ8_2;
	wire w_dff_A_qPHr3S106_2;
	wire w_dff_A_ej6mg8YW9_2;
	wire w_dff_A_HxmgycGO8_2;
	wire w_dff_A_CkR3Lkis6_2;
	wire w_dff_A_CY8HBJaz8_1;
	wire w_dff_A_gqvYkV7F0_1;
	wire w_dff_A_vhFkP5jC4_1;
	wire w_dff_A_ACkO4bKS0_1;
	wire w_dff_A_0Be0J8de3_1;
	wire w_dff_A_gGllZOSn2_1;
	wire w_dff_A_yqQWdsBy9_1;
	wire w_dff_A_iPOZRX7i5_1;
	wire w_dff_A_fdth1E2X9_1;
	wire w_dff_A_QyQBBsOP3_1;
	wire w_dff_A_UvlIyvVv4_1;
	wire w_dff_A_pdKeiF792_2;
	wire w_dff_A_yd5hhSny7_2;
	wire w_dff_A_7W3Zxmuo6_2;
	wire w_dff_A_r4VlKp9Y2_2;
	wire w_dff_B_EUSU9yvi1_3;
	wire w_dff_B_7oV083Ax8_3;
	wire w_dff_B_fEauzMyq9_3;
	wire w_dff_B_ZTw2ET2C5_3;
	wire w_dff_B_dyjCc6uR2_3;
	wire w_dff_B_x1X5DVsv4_3;
	wire w_dff_B_o0TO8GKR4_3;
	wire w_dff_A_cq0xHiKF9_1;
	wire w_dff_A_KdvOQBlZ5_2;
	wire w_dff_B_NR8kUKjf6_1;
	wire w_dff_B_WhQnq5sJ4_0;
	wire w_dff_B_KZ5ZqctT0_0;
	wire w_dff_B_SFZ16NJx3_0;
	wire w_dff_B_gtxJtZeV9_0;
	wire w_dff_B_O3ZZ2U2y0_0;
	wire w_dff_B_luJSb5d74_0;
	wire w_dff_B_pX3fj7mK9_0;
	wire w_dff_B_O1SrJoJK7_0;
	wire w_dff_B_slhLsD888_0;
	wire w_dff_B_HD260L7R7_0;
	wire w_dff_B_lMkKxrOG9_0;
	wire w_dff_B_S8Ko5jJ31_0;
	wire w_dff_B_JB0jJLuj6_0;
	wire w_dff_B_AwwbHqDV9_0;
	wire w_dff_B_Iv89Bw3L1_0;
	wire w_dff_B_qCy93SKL0_0;
	wire w_dff_B_Q8YlNiuX2_0;
	wire w_dff_B_N3bhsw929_0;
	wire w_dff_B_Y2zKwqgq8_1;
	wire w_dff_B_OaTQ7bdM2_1;
	wire w_dff_B_gTnF0hhZ1_1;
	wire w_dff_B_XmbERwBF2_1;
	wire w_dff_B_Yn4fCEHl0_1;
	wire w_dff_B_x24QcgoJ7_1;
	wire w_dff_B_om6QDEp21_1;
	wire w_dff_B_8CjxlMrm4_1;
	wire w_dff_B_GJRJsd8C2_1;
	wire w_dff_B_MQ5E8njR0_1;
	wire w_dff_B_cMWd1y872_1;
	wire w_dff_B_UChMHbeZ7_1;
	wire w_dff_B_e3dfbYO75_1;
	wire w_dff_B_7eugVS2t5_1;
	wire w_dff_B_arJRmmGp6_1;
	wire w_dff_B_KpvqEHQ73_1;
	wire w_dff_B_cPfKSmq26_1;
	wire w_dff_B_h1YwIRpF1_1;
	wire w_dff_B_ser3Szfs2_1;
	wire w_dff_B_6DkHFI564_1;
	wire w_dff_A_b2HyIx4X7_0;
	wire w_dff_A_l1KzmhGt6_0;
	wire w_dff_A_bfPMpFec3_0;
	wire w_dff_A_7wTMAY2a4_0;
	wire w_dff_A_5zgI1F9C6_0;
	wire w_dff_A_9hkTMXuv6_0;
	wire w_dff_A_6nWnQ8WQ2_2;
	wire w_dff_A_JIqhdBQF0_2;
	wire w_dff_A_aOpzuHuB4_2;
	wire w_dff_A_hP5MfCMH7_2;
	wire w_dff_A_iPooV75A1_2;
	wire w_dff_A_CBESp0Zv8_2;
	wire w_dff_A_lRH3KiF76_2;
	wire w_dff_A_4orQVfpH8_2;
	wire w_dff_A_FuUeHiEx8_2;
	wire w_dff_A_79McScpt7_2;
	wire w_dff_A_XBJgKqPn5_2;
	wire w_dff_A_zowD7kYJ3_2;
	wire w_dff_A_hlS3TIUR2_2;
	wire w_dff_A_y1aAJKTm9_2;
	wire w_dff_A_DUCTwtbJ8_2;
	wire w_dff_A_WSAtZebq9_2;
	wire w_dff_A_VE9dbpK31_2;
	wire w_dff_A_05E4x0Ju7_2;
	wire w_dff_A_BDhw5niW5_1;
	wire w_dff_A_4EjTNEXI4_1;
	wire w_dff_A_nVPydCPI0_1;
	wire w_dff_A_b7mgi8hu3_1;
	wire w_dff_A_Su36576Z0_1;
	wire w_dff_A_7z0UyjIh7_1;
	wire w_dff_A_BVgrDzBA1_1;
	wire w_dff_A_xQGBG9ho0_1;
	wire w_dff_A_Dv96yhB60_1;
	wire w_dff_A_2n6c2x286_1;
	wire w_dff_A_801GmJsc4_1;
	wire w_dff_A_DxVimEqQ5_1;
	wire w_dff_A_Vzv5zBV12_1;
	wire w_dff_A_UeDiK38c1_1;
	wire w_dff_A_uA8EBtVp2_1;
	wire w_dff_A_E0FEgWNI2_1;
	wire w_dff_A_MOLNIlYw8_2;
	wire w_dff_A_tZT1IM5d1_2;
	wire w_dff_A_32gvR2nv3_2;
	wire w_dff_A_hMyA9hSm9_2;
	wire w_dff_A_HQlyKJhr0_2;
	wire w_dff_A_g576yzHV3_2;
	wire w_dff_A_TM4UFaXR3_2;
	wire w_dff_B_uX6fm1yp9_1;
	wire w_dff_B_l55ac3zf1_1;
	wire w_dff_B_k85U420F9_1;
	wire w_dff_B_dOQvKVCU2_1;
	wire w_dff_B_Z5MpaPjb9_1;
	wire w_dff_B_eL2i8GMT5_1;
	wire w_dff_B_BKYNshWs5_1;
	wire w_dff_B_LdmblYQH9_1;
	wire w_dff_B_gqxdiTH57_1;
	wire w_dff_B_hF5jwuWr3_1;
	wire w_dff_B_S2gX7Guz7_1;
	wire w_dff_B_OJRHRCdZ1_1;
	wire w_dff_B_3YWEuYjq6_1;
	wire w_dff_B_JdvvhKqA7_1;
	wire w_dff_B_JDlRFUv94_1;
	wire w_dff_B_8dg9T0ZE7_1;
	wire w_dff_B_bjbOQTVL5_1;
	wire w_dff_B_swLcmRVK0_1;
	wire w_dff_B_yj6s74DZ0_1;
	wire w_dff_A_3aoepQuQ6_0;
	wire w_dff_A_MaiT6gHE5_0;
	wire w_dff_A_eHoJOWCv1_0;
	wire w_dff_A_vT4XYbAy8_0;
	wire w_dff_A_rN21rD7D0_0;
	wire w_dff_A_BvsbVYay0_0;
	wire w_dff_A_mIXe8xdZ8_0;
	wire w_dff_A_2gLfNMss4_2;
	wire w_dff_A_qxkoWRMr5_2;
	wire w_dff_A_kF9n7W9F8_2;
	wire w_dff_A_XGsl4uvd2_2;
	wire w_dff_A_C94puwKL4_2;
	wire w_dff_A_WGqOagTa3_2;
	wire w_dff_A_92Z6vrxQ4_2;
	wire w_dff_A_h28ilWMj8_2;
	wire w_dff_A_gXW1EJ6i6_2;
	wire w_dff_A_Zled6e9F0_2;
	wire w_dff_A_mm6LFWM94_2;
	wire w_dff_A_E9NYpw2J6_2;
	wire w_dff_A_HWRYfVeP3_2;
	wire w_dff_A_2AYdM0B88_2;
	wire w_dff_A_9ces2Q0F2_2;
	wire w_dff_A_8gVRgFJw9_2;
	wire w_dff_A_saL2bOkE4_2;
	wire w_dff_A_IqvSwh3X0_2;
	wire w_dff_A_KvJpBKkq7_2;
	wire w_dff_A_pQDVWf7y9_1;
	wire w_dff_A_yII1lfT33_1;
	wire w_dff_A_niGQDmtC9_1;
	wire w_dff_A_bAhZVycI6_1;
	wire w_dff_A_bCsgbZr89_1;
	wire w_dff_A_9VZLBhhS3_1;
	wire w_dff_A_t7GbPZJz4_1;
	wire w_dff_A_r84M9yzz2_1;
	wire w_dff_A_HKHY9Xyz9_1;
	wire w_dff_A_2eIHalnS0_1;
	wire w_dff_A_GKxW2dKs6_1;
	wire w_dff_A_mlGq3BEF8_1;
	wire w_dff_A_e6EBoZ4o1_1;
	wire w_dff_A_Qyllv4ZZ3_1;
	wire w_dff_A_UTIaLtJJ8_1;
	wire w_dff_A_OtcaZTIm7_1;
	wire w_dff_A_b0r6wlAP8_1;
	wire w_dff_A_xQFUmvbJ1_2;
	wire w_dff_A_waD4hJNb6_2;
	wire w_dff_A_OI4vDBoZ9_2;
	wire w_dff_A_XWwaykSg4_2;
	wire w_dff_A_gN2WVd530_2;
	wire w_dff_A_zj42el4G8_2;
	wire w_dff_A_vAAavfTv4_2;
	wire w_dff_A_DSuEjwyl4_2;
	wire w_dff_A_kZwk6EeY7_2;
	wire w_dff_A_YLufA5ov7_2;
	wire w_dff_A_8kV4NODC1_2;
	wire w_dff_A_hAuu7uOo4_1;
	wire w_dff_A_4K5utaxy6_2;
	wire w_dff_B_bUIEw9Ht9_1;
	wire w_dff_B_MFqRftBj7_0;
	wire w_dff_B_wwN2ZWMl5_0;
	wire w_dff_B_5HLcBw6a1_0;
	wire w_dff_B_0vi24xSR5_0;
	wire w_dff_B_WtlxMSEY0_0;
	wire w_dff_B_HA87sxbP3_0;
	wire w_dff_B_6QZC9LO09_0;
	wire w_dff_B_R1knWCXl8_0;
	wire w_dff_B_FGfREHID0_0;
	wire w_dff_B_XkOSzIVb3_0;
	wire w_dff_B_7lFzwO0I2_0;
	wire w_dff_B_NTH83tE10_0;
	wire w_dff_B_ZFAznCmj2_0;
	wire w_dff_B_4BVnWiFU5_0;
	wire w_dff_B_wet4wW6b3_0;
	wire w_dff_B_fxuBubNH2_0;
	wire w_dff_B_OiZopLEY6_0;
	wire w_dff_B_oAXzuI4Y3_0;
	wire w_dff_B_rptlmaIn4_1;
	wire w_dff_B_PEdQ3EmT9_2;
	wire w_dff_B_Ae5xATey6_2;
	wire w_dff_B_tg4sOAdy4_2;
	wire w_dff_B_wFafgjDp1_1;
	wire w_dff_B_vJYesSgQ2_1;
	wire w_dff_B_1hL04zqt9_1;
	wire w_dff_B_1XAG4UB94_1;
	wire w_dff_B_XIBLpbuT5_1;
	wire w_dff_B_7xXww1s13_1;
	wire w_dff_B_20GffJfk8_1;
	wire w_dff_B_kOF44eMj7_1;
	wire w_dff_B_FcE3S7Hb0_1;
	wire w_dff_B_ohPMvGva8_1;
	wire w_dff_B_kt67avJ57_1;
	wire w_dff_B_v4LIvFRX2_1;
	wire w_dff_B_IAUSHcP70_1;
	wire w_dff_B_rCJXoSVM0_1;
	wire w_dff_B_fI3iXvtQ8_1;
	wire w_dff_B_DRCfWsLp8_1;
	wire w_dff_B_0eWZonhG5_1;
	wire w_dff_B_SlYcJ2tf3_1;
	wire w_dff_B_cRFX9r2w7_1;
	wire w_dff_B_mPT6U0vQ3_0;
	wire w_dff_B_PxBszWCK7_0;
	wire w_dff_B_GCtCjRgK1_0;
	wire w_dff_B_A9LejHtE9_0;
	wire w_dff_B_qgpV7zM45_0;
	wire w_dff_B_zcSyOTBC1_0;
	wire w_dff_B_RRbwzLUp8_0;
	wire w_dff_B_pV9SSINE3_0;
	wire w_dff_B_H4xIpi0f4_0;
	wire w_dff_B_n41wXQkQ7_0;
	wire w_dff_B_qB89Bdb28_0;
	wire w_dff_B_sRa9pirE5_0;
	wire w_dff_B_cZ5Z913j9_0;
	wire w_dff_B_5adj63mH4_0;
	wire w_dff_B_raffp4Gz1_0;
	wire w_dff_B_DStWDLom9_0;
	wire w_dff_B_nOi1Eb6f7_0;
	wire w_dff_B_LiCEL3ez6_0;
	wire w_dff_B_ndLxsYM54_0;
	wire w_dff_A_vIxuH3bn2_1;
	wire w_dff_A_ySeyDz0k8_1;
	wire w_dff_A_sYySZKhM7_1;
	wire w_dff_A_iAeNujxT2_1;
	wire w_dff_A_GuEfVYmM7_1;
	wire w_dff_A_nngtRCkn2_1;
	wire w_dff_A_28AHSCOU8_1;
	wire w_dff_A_ljhqv3wv9_1;
	wire w_dff_A_of8p1i5s4_1;
	wire w_dff_A_V7FRgrat5_1;
	wire w_dff_A_G7nwF14k6_1;
	wire w_dff_A_h5shk5OM9_1;
	wire w_dff_A_kssqCnv77_1;
	wire w_dff_A_Qq1Quq655_1;
	wire w_dff_A_aEH3TtKE1_1;
	wire w_dff_A_zUepeZO53_1;
	wire w_dff_A_Pfw3SXlD2_1;
	wire w_dff_A_3XaApVro6_1;
	wire w_dff_A_1waapGIX9_1;
	wire w_dff_A_iMMMSng30_1;
	wire w_dff_B_BHeKXnXZ2_1;
	wire w_dff_B_KVlBrTpP5_1;
	wire w_dff_B_WefEbtTG6_1;
	wire w_dff_B_jam0XCMa2_1;
	wire w_dff_B_5n2VQ88Z8_1;
	wire w_dff_B_jqjgnu9Y6_1;
	wire w_dff_A_0WWrV3Qm4_1;
	wire w_dff_B_0IsRCJ7J0_1;
	wire w_dff_B_ToTGSQCL8_1;
	wire w_dff_B_B9H9mwxN9_1;
	wire w_dff_B_5T2WGnII4_1;
	wire w_dff_B_8GDfDaZf7_1;
	wire w_dff_B_9VPRZAvV0_1;
	wire w_dff_B_jqkJz3wv9_1;
	wire w_dff_B_Ot29YlhJ6_1;
	wire w_dff_B_Ot9mHkHa8_1;
	wire w_dff_B_tMFsKl7A6_1;
	wire w_dff_B_eVVXfIIu3_0;
	wire w_dff_B_kNcJBDK78_0;
	wire w_dff_A_QDCpwcuD4_1;
	wire w_dff_A_WZ674L7l1_1;
	wire w_dff_A_oUO70yLF7_1;
	wire w_dff_B_E8ELHlzE2_0;
	wire w_dff_B_hmBEblHa7_1;
	wire w_dff_B_IYst7Amn4_1;
	wire w_dff_B_8uPzYekn1_1;
	wire w_dff_B_g9ldojdN6_1;
	wire w_dff_B_aC24Z1dY1_1;
	wire w_dff_B_BZbrv8zs5_1;
	wire w_dff_B_Tn6q7SvF2_1;
	wire w_dff_B_42Ps8CYr7_1;
	wire w_dff_B_WbCOkQ0C7_1;
	wire w_dff_B_CnHwM22T6_1;
	wire w_dff_B_41ZhxqkA9_1;
	wire w_dff_B_nf95VBKY2_1;
	wire w_dff_B_3XZyGNpK2_1;
	wire w_dff_B_UFy47rG22_1;
	wire w_dff_B_fiyu5Gxj7_1;
	wire w_dff_B_y49ND7CU4_1;
	wire w_dff_B_OTErftW91_1;
	wire w_dff_B_1KhJuAEY4_0;
	wire w_dff_A_4fcUXYff2_0;
	wire w_dff_A_brSy7YNQ1_0;
	wire w_dff_A_XpGcU9sY8_0;
	wire w_dff_B_76ZUcUfQ7_1;
	wire w_dff_A_FkPSMB6o6_1;
	wire w_dff_A_zZCI2VO65_0;
	wire w_dff_A_xMc5mXMI1_0;
	wire w_dff_A_QI8vLCMf4_0;
	wire w_dff_A_FdhXM2JR2_0;
	wire w_dff_A_VCistAtS2_0;
	wire w_dff_A_09s7L97M0_2;
	wire w_dff_A_FTyIHLeY4_2;
	wire w_dff_A_qYfta7xC9_2;
	wire w_dff_A_hH9bAMMd6_2;
	wire w_dff_A_oyGDJ2Jt1_2;
	wire w_dff_A_p8xOZy5d0_2;
	wire w_dff_A_BCiL83yU1_1;
	wire w_dff_A_6d1ddAg80_1;
	wire w_dff_A_C3xtNIXA3_1;
	wire w_dff_A_iRhT1CDt2_1;
	wire w_dff_A_7FCyCoJM5_1;
	wire w_dff_A_7jdad2lW2_1;
	wire w_dff_A_T5NMb1MX1_2;
	wire w_dff_A_OJIT8lba9_2;
	wire w_dff_B_Mh3JndIn2_2;
	wire w_dff_B_MZQNFqqM5_2;
	wire w_dff_B_rNOq08aD8_2;
	wire w_dff_B_Yd3RaHDl1_2;
	wire w_dff_B_TVIXFEki8_2;
	wire w_dff_B_phM7qrV39_2;
	wire w_dff_B_GgWPJpw72_2;
	wire w_dff_B_ROTYPJsD2_2;
	wire w_dff_B_FSISOWg23_2;
	wire w_dff_A_rcpRD7dV0_1;
	wire w_dff_A_nLpx2NTb8_1;
	wire w_dff_A_yCOEN5au0_1;
	wire w_dff_A_Ml2bBaEz1_1;
	wire w_dff_A_67u18kr91_1;
	wire w_dff_A_c7oDginB8_1;
	wire w_dff_A_wClsaO2M6_1;
	wire w_dff_A_iWVUUbPu3_1;
	wire w_dff_A_cYWoVSJP6_1;
	wire w_dff_A_ddv5fYwH6_1;
	wire w_dff_A_k26LsMPL1_1;
	wire w_dff_A_MaU7TXpH9_1;
	wire w_dff_A_ZP4UbCEf5_1;
	wire w_dff_A_l10nIiRm6_1;
	wire w_dff_A_6BEI3sAR2_2;
	wire w_dff_A_4B1mheP25_0;
	wire w_dff_A_Gqh8Jh6F4_0;
	wire w_dff_A_fLXyLqX78_0;
	wire w_dff_A_Of2vPbt25_0;
	wire w_dff_A_z6De8r066_0;
	wire w_dff_A_hVQnnvja8_0;
	wire w_dff_A_59eggMik5_0;
	wire w_dff_A_rsD7FIMN5_0;
	wire w_dff_A_RcUXlHWv0_0;
	wire w_dff_A_WaAZAjwT5_0;
	wire w_dff_A_7HpJId9l8_0;
	wire w_dff_A_nLPM3D7D0_0;
	wire w_dff_B_uCKs5HVf6_1;
	wire w_dff_B_wtl9Oema5_0;
	wire w_dff_B_Flsaga4c0_0;
	wire w_dff_B_nXVhM1Rx0_0;
	wire w_dff_B_qscW8IVx3_0;
	wire w_dff_A_iLfKEUtW7_1;
	wire w_dff_A_PXyvd2ks5_1;
	wire w_dff_A_9O5UXZ154_1;
	wire w_dff_A_qFTtFlRi2_1;
	wire w_dff_A_RjAXddZ37_1;
	wire w_dff_B_kt9B0qJD9_2;
	wire w_dff_B_MOfdpE6P9_2;
	wire w_dff_B_Nj8WUajz9_2;
	wire w_dff_B_SLMTPtCs1_2;
	wire w_dff_B_BywBpOYm8_2;
	wire w_dff_B_rZr6ZrTy5_0;
	wire w_dff_B_3RbFhSx97_0;
	wire w_dff_B_c2AMwgBo0_1;
	wire w_dff_B_0prXEDw41_1;
	wire w_dff_B_ztEuUki02_1;
	wire w_dff_A_Cka2V7856_1;
	wire w_dff_A_3wpdnrIV2_1;
	wire w_dff_A_tPlTKaWH6_1;
	wire w_dff_A_dhReTvlB7_2;
	wire w_dff_A_ePq601SJ4_2;
	wire w_dff_A_GxFhgmSn1_2;
	wire w_dff_A_CsVBg2om0_2;
	wire w_dff_A_fREJw3An9_2;
	wire w_dff_A_U6OwVIsN2_2;
	wire w_dff_A_HqFGmp4m9_2;
	wire w_dff_B_HqYOc0uM0_3;
	wire w_dff_A_y7xTsVOc6_0;
	wire w_dff_A_kun5VUET6_0;
	wire w_dff_A_tBp2Hsn68_0;
	wire w_dff_A_jYxV5az43_0;
	wire w_dff_A_ssGrBkRW2_0;
	wire w_dff_A_axq4HGjQ0_0;
	wire w_dff_A_Ussb0dT78_0;
	wire w_dff_A_L14DxMQa2_0;
	wire w_dff_A_Td0FQIsI3_0;
	wire w_dff_B_4M2MQAlr4_1;
	wire w_dff_A_NgjfhL585_1;
	wire w_dff_A_9b00a6Wm0_0;
	wire w_dff_A_WM9O4aQN3_0;
	wire w_dff_A_PziGP8hv4_0;
	wire w_dff_A_R3Yk2wKz5_0;
	wire w_dff_A_ZSZNXX9l0_0;
	wire w_dff_A_VEFizTQq6_0;
	wire w_dff_A_D3LNxEph9_0;
	wire w_dff_A_7OoVbUce7_0;
	wire w_dff_A_0Yj7e50W7_0;
	wire w_dff_A_rcOAliD40_2;
	wire w_dff_A_vuGKH9bt2_2;
	wire w_dff_A_3fHr742m8_2;
	wire w_dff_A_rjE4E3PC6_2;
	wire w_dff_A_ZiHBGFqw1_2;
	wire w_dff_A_h601iIzf1_2;
	wire w_dff_B_ajomxJhW9_0;
	wire w_dff_B_OVby5Z5C3_1;
	wire w_dff_A_9Z8YzaJR0_0;
	wire w_dff_A_hoLr25wI1_0;
	wire w_dff_A_333dDAbD8_0;
	wire w_dff_A_1Cp6KO1i0_0;
	wire w_dff_A_HHnB3VB34_0;
	wire w_dff_A_neDUdMgU6_0;
	wire w_dff_A_VNnF3vLh9_0;
	wire w_dff_A_Ucl5ZpZa5_0;
	wire w_dff_A_78w0CKoW7_0;
	wire w_dff_A_Ln1P0pbx4_0;
	wire w_dff_A_D7AxmQ9P6_0;
	wire w_dff_A_4ZtY3t7X9_0;
	wire w_dff_A_6BIevfPr4_0;
	wire w_dff_B_UOnL0LPK6_0;
	wire w_dff_B_5Qogf0L47_1;
	wire w_dff_A_1SvuEk1l6_1;
	wire w_dff_A_T34XIiGr7_2;
	wire w_dff_A_Un4by8Su6_2;
	wire w_dff_A_TBuxjPfM6_2;
	wire w_dff_A_PZ46vJmd6_2;
	wire w_dff_A_b6iIEez91_2;
	wire w_dff_A_tE1zBRHh8_2;
	wire w_dff_A_gpHzgrZb4_2;
	wire w_dff_A_Nj4cffsC8_2;
	wire w_dff_A_zDCSsXC69_2;
	wire w_dff_A_FCeaU0Lj3_2;
	wire w_dff_A_LO8JhS1b5_2;
	wire w_dff_B_wQ37Nmac5_1;
	wire w_dff_B_Cqd1kKUi5_1;
	wire w_dff_B_ueR6QxYH8_0;
	wire w_dff_B_0n2iSvza1_0;
	wire w_dff_B_sTEgEJtc9_0;
	wire w_dff_A_tVf5I4i34_0;
	wire w_dff_A_TGiwqkbc7_0;
	wire w_dff_A_BHyEiyWj8_0;
	wire w_dff_A_gRJu8dra0_1;
	wire w_dff_A_PaftL0gZ0_1;
	wire w_dff_A_t9pJYt2t9_1;
	wire w_dff_A_OuIvP6MH8_1;
	wire w_dff_B_sy6KjLuo3_0;
	wire w_dff_A_6FBPsbun8_0;
	wire w_dff_A_zIdAlXXi9_2;
	wire w_dff_A_VdAWrNPu1_0;
	wire w_dff_B_rRKEK39E6_0;
	wire w_dff_A_3lcgRqEX1_0;
	wire w_dff_A_Pf5VAkFP8_0;
	wire w_dff_A_sXQc0UB34_0;
	wire w_dff_A_bGQnNttp7_0;
	wire w_dff_A_NTRfhQdx2_0;
	wire w_dff_A_hgT2m9R40_0;
	wire w_dff_A_x0rP3c8Z5_0;
	wire w_dff_A_FRltRma56_0;
	wire w_dff_A_Px5ZGXrK0_0;
	wire w_dff_A_uaJnVHqy2_0;
	wire w_dff_A_Z08EWguM7_0;
	wire w_dff_A_l5bz6pxi6_2;
	wire w_dff_A_16V4Hxzh5_2;
	wire w_dff_A_fixQuJMB8_2;
	wire w_dff_A_hoAfj9jr7_2;
	wire w_dff_A_4GDP5TXL1_2;
	wire w_dff_A_1wQP34qU5_2;
	wire w_dff_A_LwJ5T8GU8_2;
	wire w_dff_A_5KgIyjV38_2;
	wire w_dff_B_nwTId6tV3_1;
	wire w_dff_B_TNNtcrsm6_1;
	wire w_dff_B_BWdDp12D4_1;
	wire w_dff_B_pZXcCq6v4_1;
	wire w_dff_B_j3t6z3pP4_1;
	wire w_dff_B_37SCrA0S9_1;
	wire w_dff_B_3iwYDHDS5_1;
	wire w_dff_B_36KGz4ig5_1;
	wire w_dff_B_N3s96bPx9_1;
	wire w_dff_B_wvi7Aap69_1;
	wire w_dff_B_s7NA25D62_1;
	wire w_dff_B_geJVyNwW7_1;
	wire w_dff_B_32HAyE5l5_1;
	wire w_dff_B_RUmbkIb40_1;
	wire w_dff_B_zFRFbdqH0_1;
	wire w_dff_A_2osJTg5r6_0;
	wire w_dff_A_64zhRRF94_0;
	wire w_dff_A_lKBBG9nc4_1;
	wire w_dff_A_iIioO9lY3_1;
	wire w_dff_A_TpbrnZoO6_1;
	wire w_dff_A_0gVNNokL9_1;
	wire w_dff_A_1Lie9nTu7_1;
	wire w_dff_A_RRSfynhV3_1;
	wire w_dff_A_EcPFPxEC7_0;
	wire w_dff_A_HIVMkKha8_0;
	wire w_dff_A_sYehwKfj0_1;
	wire w_dff_A_6ITWIBCe7_1;
	wire w_dff_A_41tmBw654_1;
	wire w_dff_A_b8mN4CkN8_1;
	wire w_dff_A_tphtfBPB4_2;
	wire w_dff_A_VhxFh8dI9_2;
	wire w_dff_A_F1MW2BrB7_0;
	wire w_dff_A_SjAokIeW6_0;
	wire w_dff_A_wnFGLyFC2_0;
	wire w_dff_A_W8kNSJ959_1;
	wire w_dff_A_CrsoojyL3_0;
	wire w_dff_A_iDRi8Z7q6_2;
	wire w_dff_A_RHDn8gJ77_0;
	wire w_dff_A_NGjVTmbe1_0;
	wire w_dff_A_Vfr0JD8t2_0;
	wire w_dff_A_sPNwFVsy2_0;
	wire w_dff_A_qTO4q7QN5_1;
	wire w_dff_A_5lRKS5Go0_1;
	wire w_dff_A_vZh9OXyE6_2;
	wire w_dff_A_DThUBnis6_2;
	wire w_dff_A_OnmdS1oM1_2;
	wire w_dff_A_0LLucqvu0_2;
	wire w_dff_B_Tse1RMZe5_1;
	wire w_dff_A_EeOoDiHL9_0;
	wire w_dff_A_XlcVMFwu1_2;
	wire w_dff_A_AvITlxYr9_1;
	wire w_dff_A_8snwYWZG3_0;
	wire w_dff_A_j84CDqMi4_0;
	wire w_dff_A_sF3fyNOK1_0;
	wire w_dff_A_6suxaqd71_0;
	wire w_dff_A_1771ZTwu0_0;
	wire w_dff_A_miAybj3Y3_0;
	wire w_dff_A_EZ2RwlKo8_0;
	wire w_dff_B_CbKVzz7k2_1;
	wire w_dff_B_r7EWpylQ1_1;
	wire w_dff_A_yTm2tt4S6_1;
	wire w_dff_A_3oiJsFeB4_1;
	wire w_dff_A_yupCMjfw9_1;
	wire w_dff_A_CUzQPcYa0_1;
	wire w_dff_A_82YZAv663_1;
	wire w_dff_A_GKwyiBR81_1;
	wire w_dff_A_nIvZjjzB4_1;
	wire w_dff_A_2aYNoF4G8_1;
	wire w_dff_A_FUbKw7eB0_1;
	wire w_dff_A_UBRmLcbE0_1;
	wire w_dff_A_oXLwo3uF8_1;
	wire w_dff_A_y5ZDPO9D8_1;
	wire w_dff_A_3fzlM4684_1;
	wire w_dff_A_WZaGHca36_1;
	wire w_dff_A_FVXWl3FD7_1;
	wire w_dff_A_kjImmVOb9_1;
	wire w_dff_A_6SFRLNe67_1;
	wire w_dff_A_hl1WHQlu0_1;
	wire w_dff_A_D3C8o9HN8_2;
	wire w_dff_A_fYMbMDMp3_2;
	wire w_dff_A_BgaD9RHb7_2;
	wire w_dff_A_2p0oSSNB8_2;
	wire w_dff_A_0e6U2DBd6_2;
	wire w_dff_A_Xuznx5uz1_2;
	wire w_dff_A_rTU8kwPP7_2;
	wire w_dff_A_d4unRuEc8_2;
	wire w_dff_A_Nia2hEuS7_2;
	wire w_dff_A_Dcor2tS24_2;
	wire w_dff_A_om3N0AQY7_0;
	wire w_dff_A_sN4mtC7W7_0;
	wire w_dff_B_PByhN64L5_1;
	wire w_dff_B_sPMlff716_1;
	wire w_dff_B_nHvIWuat9_1;
	wire w_dff_B_MPpmLCTT3_1;
	wire w_dff_A_t9VyOwxo3_1;
	wire w_dff_A_KI74boHH4_0;
	wire w_dff_A_JLWgZOeG5_0;
	wire w_dff_A_Xge3qlDa3_0;
	wire w_dff_A_FFQSG4AZ9_0;
	wire w_dff_A_R2qompgH1_1;
	wire w_dff_A_5HmmIuF97_1;
	wire w_dff_A_84OCqbd11_1;
	wire w_dff_A_vrlvvKg91_2;
	wire w_dff_A_5zYvxq7W2_2;
	wire w_dff_A_LGtPvX8K8_2;
	wire w_dff_A_HyLyg6kX7_2;
	wire w_dff_A_f2Bes9Bs9_1;
	wire w_dff_A_X2o6mQP26_1;
	wire w_dff_B_pk6zXsK44_1;
	wire w_dff_B_QKm8l0wr0_1;
	wire w_dff_A_a3hhoJix0_2;
	wire w_dff_B_yHrQBdqF8_3;
	wire w_dff_A_xzOc3OnQ6_0;
	wire w_dff_A_Bv3pi35O0_0;
	wire w_dff_A_FFhWWLlg1_0;
	wire w_dff_A_DX0O2Syd8_1;
	wire w_dff_B_LBOSmfTe1_1;
	wire w_dff_A_HY2aFV2P3_1;
	wire w_dff_A_ELM8S4fv3_1;
	wire w_dff_A_vd4oStN78_1;
	wire w_dff_A_JjHqfE2P8_2;
	wire w_dff_A_4gOKqh2V3_2;
	wire w_dff_A_ogSajMlJ4_2;
	wire w_dff_A_hXqnvGe07_0;
	wire w_dff_A_tVLIpjof3_2;
	wire w_dff_A_tg6NZPpn6_1;
	wire w_dff_A_HajIFmL30_2;
	wire w_dff_A_Z4IRXIZx4_2;
	wire w_dff_A_2gyqCwep7_1;
	wire w_dff_B_Q9sxPbQ39_1;
	wire w_dff_B_Xn8RU2f01_1;
	wire w_dff_B_hVArdk7n8_1;
	wire w_dff_B_mR1RJ9Tk9_1;
	wire w_dff_B_MzvEPU5s9_1;
	wire w_dff_A_A5X5yhsF9_0;
	wire w_dff_A_v7GQKGqV5_0;
	wire w_dff_A_XRPK02d44_0;
	wire w_dff_A_p6vRd7Fz8_1;
	wire w_dff_A_nzThzmNM3_1;
	wire w_dff_A_VpsuK4DU7_1;
	wire w_dff_A_KPhwFbOo5_1;
	wire w_dff_A_wQ07uUHs9_1;
	wire w_dff_A_5b5e9Wvx1_2;
	wire w_dff_A_x4tZzhZR6_2;
	wire w_dff_A_OJtfwC613_2;
	wire w_dff_A_WRca75ot1_0;
	wire w_dff_B_65tFn0Ix8_1;
	wire w_dff_B_eBibGzSN8_1;
	wire w_dff_A_AO0pwfjq9_0;
	wire w_dff_A_lWn202HJ2_0;
	wire w_dff_A_E50FNLHQ9_0;
	wire w_dff_A_5vLUvMLA7_0;
	wire w_dff_A_38xu0fvJ7_0;
	wire w_dff_A_srWn93J30_1;
	wire w_dff_A_LUrWZIuz1_1;
	wire w_dff_A_wvmDIRuM7_1;
	wire w_dff_A_QPWzXnZF4_2;
	wire w_dff_A_3IDIkQpR3_2;
	wire w_dff_A_YYBiyCFM4_2;
	wire w_dff_A_Z06Ba6Xd8_0;
	wire w_dff_A_FTOzRZ710_0;
	wire w_dff_A_5EZWNJ094_1;
	wire w_dff_A_tYEALtjI1_0;
	wire w_dff_A_55YIOMal5_2;
	wire w_dff_A_ClLpTeIE1_1;
	wire w_dff_B_ZC3lkNWB4_1;
	wire w_dff_B_G3JSTTyC0_1;
	wire w_dff_A_ugTUNeBj5_0;
	wire w_dff_A_hiWDEWT99_2;
	wire w_dff_A_UKFq0IAf2_2;
	wire w_dff_A_7maiGc5N3_0;
	wire w_dff_A_sDHb6b4O3_1;
	wire w_dff_A_R93ISZ5k6_1;
	wire w_dff_A_Jk1aUJmI7_1;
	wire w_dff_A_6jMeSYC38_2;
	wire w_dff_A_7dGOx6od9_2;
	wire w_dff_A_YGYkLDhj5_1;
	wire w_dff_A_YiyeAhCF0_2;
	wire w_dff_A_9Oadu2nu0_2;
	wire w_dff_A_9AB4Gv7c2_2;
	wire w_dff_A_H74xHTCF5_2;
	wire w_dff_A_5GfGXW058_2;
	wire w_dff_A_mqFVnjb22_2;
	wire w_dff_A_dfRVq1zI3_2;
	wire w_dff_A_ej7CPOa77_2;
	wire w_dff_A_zipsQr5v1_2;
	wire w_dff_A_YM6urWMD0_2;
	wire w_dff_A_BDSPxLJq6_2;
	wire w_dff_A_mTgfSlbB7_2;
	wire w_dff_A_7ggp5Ux39_0;
	wire w_dff_A_nnZXttfa8_0;
	wire w_dff_A_0tyBVRu23_0;
	wire w_dff_A_CSjwxdJN3_0;
	wire w_dff_A_D1dy12dg0_0;
	wire w_dff_A_966KkFoe3_0;
	wire w_dff_A_KW6NuIfj9_2;
	wire w_dff_A_nCKZH5oX1_2;
	wire w_dff_A_lT6JCe9K1_2;
	wire w_dff_A_QGWsjoSk8_2;
	wire w_dff_A_Q1kJlyPq1_2;
	wire w_dff_A_O5b5TPBz6_2;
	wire w_dff_A_zVpT7JMg6_2;
	wire w_dff_A_hvbSankV7_2;
	wire w_dff_A_ZMoQtbfK2_2;
	wire w_dff_A_cjfNjDfN8_2;
	wire w_dff_A_5M8zWWMe8_2;
	wire w_dff_A_rANZesdT1_2;
	wire w_dff_A_hYVvEH8k1_2;
	wire w_dff_A_DRiJzPKp3_2;
	wire w_dff_A_MzHK8kA45_2;
	wire w_dff_A_ovlJJ6Mc1_2;
	wire w_dff_A_Dfx2R6WO6_2;
	wire w_dff_A_q93wqV3h6_2;
	wire w_dff_A_voDyk4lD2_1;
	wire w_dff_A_cIlpqCWR9_1;
	wire w_dff_A_RUOoy5O83_1;
	wire w_dff_A_WdZ9Phl33_1;
	wire w_dff_A_MIbnbtuL8_1;
	wire w_dff_A_AF624G4h9_1;
	wire w_dff_A_XrkqKJF24_1;
	wire w_dff_A_yt3tsEhN3_1;
	wire w_dff_A_xHk4giye6_1;
	wire w_dff_A_qSiXrfL87_1;
	wire w_dff_A_tlpMJSzr4_1;
	wire w_dff_A_RQnR9Z2z7_1;
	wire w_dff_A_8NeluTTn1_1;
	wire w_dff_A_Bz2T7az03_1;
	wire w_dff_A_tPdzturL8_1;
	wire w_dff_A_IJvihPOl2_1;
	wire w_dff_A_RVqfX0ie3_2;
	wire w_dff_A_FRwjEamb9_2;
	wire w_dff_A_MMUzKkQ14_2;
	wire w_dff_A_xSw0jKL40_2;
	wire w_dff_A_aC7ZYpJE6_2;
	wire w_dff_A_ZpM9mmJf0_2;
	wire w_dff_A_Qs8lUsEQ2_2;
	wire w_dff_B_liGyRj4Q1_1;
	wire w_dff_B_OJ5HfNRL9_1;
	wire w_dff_B_0TEmTxzM6_1;
	wire w_dff_B_0aP2VCWM6_1;
	wire w_dff_B_08P3VPFK4_1;
	wire w_dff_B_omhSyZ459_1;
	wire w_dff_B_jckNwaR91_1;
	wire w_dff_B_MLQIsMuH8_1;
	wire w_dff_B_7jWKwy5r6_1;
	wire w_dff_B_UE95Re2t4_1;
	wire w_dff_B_ddPsgluX1_1;
	wire w_dff_B_M7gHhWNt2_1;
	wire w_dff_B_1JIu4NRL5_1;
	wire w_dff_B_bkC1scp71_1;
	wire w_dff_B_lw3J3g0N6_1;
	wire w_dff_B_Vss8iiPJ5_1;
	wire w_dff_B_65m2zDPh4_1;
	wire w_dff_B_FcdK7Hcj1_1;
	wire w_dff_B_pR7GSL0Y7_1;
	wire w_dff_B_e0zrZFup3_0;
	wire w_dff_B_6O7fnQNo2_0;
	wire w_dff_B_zWB4DmA52_0;
	wire w_dff_B_XBWlxRN51_0;
	wire w_dff_B_dl97fqRg4_0;
	wire w_dff_B_lSCZGfZS8_0;
	wire w_dff_B_FolDlFxt7_0;
	wire w_dff_B_ovF0zvai4_0;
	wire w_dff_B_FUwn0LRS8_0;
	wire w_dff_B_7f94zMcT0_0;
	wire w_dff_B_o3gIcTf50_0;
	wire w_dff_B_ipHBBiCP9_0;
	wire w_dff_B_JYjRxzTa0_0;
	wire w_dff_B_2f0bdyTH6_0;
	wire w_dff_B_5qGAiS8O8_0;
	wire w_dff_B_K8rmROJK2_0;
	wire w_dff_B_2huLCqb88_0;
	wire w_dff_B_NPy4TpUC3_0;
	wire w_dff_B_Yrygy9EL4_0;
	wire w_dff_B_yCq0ZVJN9_1;
	wire w_dff_B_JbFcHKGO0_1;
	wire w_dff_B_zuUBF6Gq3_1;
	wire w_dff_B_WhspaehD7_1;
	wire w_dff_B_B2x6Xiyd7_1;
	wire w_dff_B_lEtp34gp1_1;
	wire w_dff_B_tYi7udAD2_1;
	wire w_dff_B_QcHQcyID4_1;
	wire w_dff_B_s4uYJj257_0;
	wire w_dff_B_iCRNtnLO0_0;
	wire w_dff_B_EtojTeXx9_1;
	wire w_dff_B_ohrudmbV7_0;
	wire w_dff_B_XxUMWEiy2_0;
	wire w_dff_B_aWwzQuXm1_0;
	wire w_dff_B_OZLQFGTU9_0;
	wire w_dff_B_1ugzbJt42_1;
	wire w_dff_B_yhPL1mvI4_1;
	wire w_dff_B_fiXlRQhm6_1;
	wire w_dff_B_U7FZVWcd5_1;
	wire w_dff_B_bxgfQRrM6_1;
	wire w_dff_B_SUWRyUAo3_1;
	wire w_dff_B_5PhlypIg2_1;
	wire w_dff_B_rYGBZQAS1_1;
	wire w_dff_B_9ndrnDAh8_1;
	wire w_dff_B_nnE2UKrf0_1;
	wire w_dff_B_xgf0Q80y2_1;
	wire w_dff_B_cMf6aa0h5_1;
	wire w_dff_B_KYhvU6y66_1;
	wire w_dff_B_dTFJsWoQ6_1;
	wire w_dff_B_8wmzcDz37_1;
	wire w_dff_B_BY6gYS6B7_1;
	wire w_dff_B_s14nKBMl3_1;
	wire w_dff_B_Gq9c9ON17_1;
	wire w_dff_B_ilc10LQn9_1;
	wire w_dff_B_PpbW6kti0_1;
	wire w_dff_B_ECree2Cn4_1;
	wire w_dff_B_gi6eUhAL8_1;
	wire w_dff_B_KctnXjBN9_1;
	wire w_dff_A_XXL0aiQW4_0;
	wire w_dff_A_an92ggBv9_1;
	wire w_dff_B_swnD9oMO4_2;
	wire w_dff_B_WUOsOuwl1_2;
	wire w_dff_B_t5ysg7OS6_2;
	wire w_dff_B_P1SYit4Z8_2;
	wire w_dff_A_UFU9iMn87_0;
	wire w_dff_A_VBWCWI629_0;
	wire w_dff_A_3QGKgOPX4_0;
	wire w_dff_A_5ZnwEata7_0;
	wire w_dff_A_IznMhbn49_1;
	wire w_dff_A_QBOcDrZP2_1;
	wire w_dff_B_yPRmIuMF4_1;
	wire w_dff_B_bPw4S0de1_0;
	wire w_dff_B_tJK6alD19_1;
	wire w_dff_A_TQPcLq8Y1_0;
	wire w_dff_A_qVskqiBq8_0;
	wire w_dff_B_5mIHG5uh0_2;
	wire w_dff_B_dTE99gFY9_2;
	wire w_dff_B_M0lIgbye8_2;
	wire w_dff_B_g7CoFDCG5_2;
	wire w_dff_B_i2ziskj46_2;
	wire w_dff_B_g7uquTPI9_2;
	wire w_dff_B_szxuXp6g0_0;
	wire w_dff_B_Bv05TyMV1_0;
	wire w_dff_B_znBonFDJ3_0;
	wire w_dff_B_2MSOpb3o0_0;
	wire w_dff_B_JzQBGI5E3_0;
	wire w_dff_B_M7YL1Mkh1_0;
	wire w_dff_B_2CZqcMtj8_0;
	wire w_dff_B_rbzmz5CZ9_0;
	wire w_dff_A_6UUSTrVX6_2;
	wire w_dff_A_3etelolD8_2;
	wire w_dff_A_3caDZTan3_2;
	wire w_dff_A_X1Meqaci4_2;
	wire w_dff_A_KQupukqT0_2;
	wire w_dff_A_uIv2YcRA2_2;
	wire w_dff_A_yybsGvv85_2;
	wire w_dff_A_xsWpch2G5_2;
	wire w_dff_A_XWtA6UuR0_2;
	wire w_dff_A_sfWyFTcT3_2;
	wire w_dff_A_JVPgjwDp8_2;
	wire w_dff_A_Aw2TO8zp6_2;
	wire w_dff_A_eEZ6ClbX2_1;
	wire w_dff_A_vPpa6Jj87_1;
	wire w_dff_A_ZpyLbyDc0_1;
	wire w_dff_A_8kukiMfi7_1;
	wire w_dff_A_A497m73K3_1;
	wire w_dff_A_SbvhoUPS6_1;
	wire w_dff_A_ZFnKkMIO5_1;
	wire w_dff_A_Wf9am40F1_1;
	wire w_dff_A_QwGW2V7L3_1;
	wire w_dff_A_wYlswrCS8_2;
	wire w_dff_A_51KeTvav3_2;
	wire w_dff_A_Wp43asRs1_2;
	wire w_dff_A_23vj8eKw1_2;
	wire w_dff_A_1i58seqN6_2;
	wire w_dff_A_HkAEoIV02_2;
	wire w_dff_A_tVodmN4C5_2;
	wire w_dff_A_iimUTs6z2_2;
	wire w_dff_A_knsfbCJo1_2;
	wire w_dff_B_JYxjRNqs6_3;
	wire w_dff_B_3ijbnRXv9_3;
	wire w_dff_A_Hy1lOvfA7_1;
	wire w_dff_A_AAFa1FuD2_1;
	wire w_dff_A_PPHdl43q8_1;
	wire w_dff_A_Lg42zLWs3_0;
	wire w_dff_B_jWVFJh3J6_1;
	wire w_dff_B_fJkWUVKm7_1;
	wire w_dff_B_k5g8YeC02_0;
	wire w_dff_B_XgANFRu84_1;
	wire w_dff_B_rsIdIZLY8_2;
	wire w_dff_A_qxb4VXKh9_0;
	wire w_dff_B_rlpoLhJZ6_0;
	wire w_dff_B_Od3WhJOn7_1;
	wire w_dff_A_3Xzr9Mok0_1;
	wire w_dff_A_COxX6Hug9_1;
	wire w_dff_A_H5f7fWQY6_1;
	wire w_dff_A_Eq4TaIX45_1;
	wire w_dff_A_V3yLGFNH1_1;
	wire w_dff_A_ZkPL7UUL6_1;
	wire w_dff_A_459UX8bo9_1;
	wire w_dff_A_xUmdKPGb9_1;
	wire w_dff_A_G8ZG0IOT3_1;
	wire w_dff_B_od7BNBhR9_2;
	wire w_dff_B_dPTIeqpS1_2;
	wire w_dff_B_r59SndGa8_2;
	wire w_dff_A_vyfh7V7W4_0;
	wire w_dff_A_eBUFyfDL9_0;
	wire w_dff_A_7wscXeRN4_0;
	wire w_dff_A_AutBRX7P6_0;
	wire w_dff_A_Hgu7Ljw35_0;
	wire w_dff_B_sQt5zr0P4_1;
	wire w_dff_B_VZOWUMFk6_1;
	wire w_dff_B_j6uxmmWU0_0;
	wire w_dff_A_oyEdJAoc4_0;
	wire w_dff_B_MrI0xqPx9_0;
	wire w_dff_B_CLDgGND10_0;
	wire w_dff_A_srezomRw5_0;
	wire w_dff_A_LnIAdAHM9_0;
	wire w_dff_A_mTq4iD9w4_0;
	wire w_dff_A_B2mDDxTW7_0;
	wire w_dff_A_claZv6Kr0_0;
	wire w_dff_A_kAGnBtDr9_0;
	wire w_dff_A_vOM2tzt18_0;
	wire w_dff_A_T1e90f7s3_1;
	wire w_dff_A_r9gdVtro5_1;
	wire w_dff_A_Uk9XHvCw3_1;
	wire w_dff_A_aqXlXeOX2_1;
	wire w_dff_A_Post4hJQ0_0;
	wire w_dff_A_67razSdm1_0;
	wire w_dff_A_ZUyMMdJq0_0;
	wire w_dff_A_pnldaA2v3_0;
	wire w_dff_A_hfuoI0jo8_0;
	wire w_dff_A_uQZAZQvC3_0;
	wire w_dff_B_ussOJq4x6_2;
	wire w_dff_B_Al0hJv4B7_2;
	wire w_dff_A_im8jegML9_0;
	wire w_dff_A_CyFevzjJ5_1;
	wire w_dff_A_BZcAxFcO4_1;
	wire w_dff_A_zoXmK7Iz9_1;
	wire w_dff_A_nvPNabXU6_0;
	wire w_dff_A_sGYejoD97_0;
	wire w_dff_A_A30FOO4l2_0;
	wire w_dff_A_mryewm2Q4_0;
	wire w_dff_A_8pyzMGoY5_0;
	wire w_dff_A_NgA305G65_0;
	wire w_dff_A_DB7W0JUv0_0;
	wire w_dff_A_gPrNeSA64_0;
	wire w_dff_A_nLKpNx1b7_0;
	wire w_dff_A_atBJ4bHd9_0;
	wire w_dff_A_OTWRGP8Y7_0;
	wire w_dff_A_YEIBHXyR5_0;
	wire w_dff_A_XXcrqkgg2_2;
	wire w_dff_A_AHaBidWx0_2;
	wire w_dff_A_m2xroV9f9_2;
	wire w_dff_A_NdBLsNQB4_2;
	wire w_dff_A_YJvAUXfQ2_2;
	wire w_dff_A_MG58C1ah5_2;
	wire w_dff_A_Jaq0R8y90_2;
	wire w_dff_A_fqtU4tWr0_2;
	wire w_dff_A_JYsk3MQM5_2;
	wire w_dff_A_dHQDRExs4_2;
	wire w_dff_B_VYjxetyZ9_1;
	wire w_dff_B_l5JERaAC2_1;
	wire w_dff_B_DPpmcpte9_1;
	wire w_dff_B_DeBgD0QU3_1;
	wire w_dff_B_6tPrnNlL0_1;
	wire w_dff_B_GAskT40k0_1;
	wire w_dff_B_Mr5vgPFN9_1;
	wire w_dff_B_lJf389oy3_1;
	wire w_dff_B_Db1QQsdW2_1;
	wire w_dff_A_8wQEgTCA2_1;
	wire w_dff_A_UIiibPO25_0;
	wire w_dff_A_geAXsMnP2_0;
	wire w_dff_A_JJrjz0nd1_1;
	wire w_dff_A_YuoYuwoU9_1;
	wire w_dff_A_8a6PCgz73_1;
	wire w_dff_A_DcXsmqnS8_1;
	wire w_dff_A_C6bAeuK52_2;
	wire w_dff_A_omfJLI8Y4_2;
	wire w_dff_A_xmhvvj0Z8_2;
	wire w_dff_A_MsUDDw1v4_1;
	wire w_dff_A_o9qhUCMZ1_1;
	wire w_dff_A_Iw5jiIn26_0;
	wire w_dff_A_zfHbfcdg1_0;
	wire w_dff_A_7EVxPVdw9_0;
	wire w_dff_A_gIyESD6S9_1;
	wire w_dff_B_JaGxgQWT2_2;
	wire w_dff_A_yGT0P50w9_0;
	wire w_dff_A_EgTalk5v9_1;
	wire w_dff_A_4qE7KPEQ0_1;
	wire w_dff_A_iH4CnHb29_1;
	wire w_dff_A_o6BsNIX50_1;
	wire w_dff_A_8N7eNG3U7_1;
	wire w_dff_B_KJPtpKsx2_1;
	wire w_dff_B_KBAynGeM1_1;
	wire w_dff_B_HPOgCEnt4_2;
	wire w_dff_B_JXXNJSkA4_2;
	wire w_dff_B_KzH9yKB38_2;
	wire w_dff_B_j90GPViM9_2;
	wire w_dff_B_W5NYCNTJ1_2;
	wire w_dff_B_xf1oSZ5z0_2;
	wire w_dff_B_pNYRD1394_2;
	wire w_dff_B_oqpHiaKM8_2;
	wire w_dff_B_12Zklbrq1_2;
	wire w_dff_B_ev8wgKxz4_2;
	wire w_dff_A_Ts12P0AV9_2;
	wire w_dff_A_0qwZDuaV1_2;
	wire w_dff_A_2dhCT1Wk4_2;
	wire w_dff_A_5TKP5dxK2_2;
	wire w_dff_A_crk6p3iG6_2;
	wire w_dff_A_kd1v6NbK6_1;
	wire w_dff_A_y0pz9t1g3_1;
	wire w_dff_A_8cro9meK8_1;
	wire w_dff_A_Rura2hEo7_1;
	wire w_dff_A_2VGnmVt25_1;
	wire w_dff_A_JOdOdnOj3_1;
	wire w_dff_A_FaJwG62n8_1;
	wire w_dff_B_tbhq58vP9_0;
	wire w_dff_A_D4JVfPTQ7_0;
	wire w_dff_B_LFNFrl5q5_1;
	wire w_dff_A_Nf3spo5L7_0;
	wire w_dff_A_M1zNiXjj5_0;
	wire w_dff_A_5qs9epFC4_1;
	wire w_dff_A_9nVRPNt67_1;
	wire w_dff_A_pdR9RIH36_1;
	wire w_dff_A_by5yijvO9_1;
	wire w_dff_A_bU9h8p941_1;
	wire w_dff_A_kbQ3KtJP4_1;
	wire w_dff_A_et7Eq4Wx6_1;
	wire w_dff_A_IreSGpQ86_1;
	wire w_dff_A_PmNSlo4L5_1;
	wire w_dff_A_waBRAppj0_1;
	wire w_dff_A_J9WXGZ522_1;
	wire w_dff_A_dt1Fa41b3_1;
	wire w_dff_A_WZBf4SCa2_1;
	wire w_dff_A_lDjO1o2S5_1;
	wire w_dff_A_f8CAGVsM8_1;
	wire w_dff_A_FWYweYQo4_1;
	wire w_dff_B_uFZfeLal0_0;
	wire w_dff_B_hfdQdMaW8_1;
	wire w_dff_A_dINxCVap4_0;
	wire w_dff_A_z285s69A9_2;
	wire w_dff_A_I24ibmv85_1;
	wire w_dff_A_yEZO1IIM9_1;
	wire w_dff_A_DGq2Bw4E3_1;
	wire w_dff_A_p0aJPN2Z1_1;
	wire w_dff_A_36lCpSwf6_1;
	wire w_dff_A_4yC9fNkP6_1;
	wire w_dff_A_hPcV7d4t9_1;
	wire w_dff_A_GpGtVjMW1_1;
	wire w_dff_A_WXAGokCV2_1;
	wire w_dff_A_nPYokcY65_1;
	wire w_dff_A_zZjDeUYC9_1;
	wire w_dff_A_PSuEwDMR0_1;
	wire w_dff_A_4pP9wztx5_1;
	wire w_dff_A_qDVqyDDb1_1;
	wire w_dff_A_jTz3AAI64_1;
	wire w_dff_A_7x98A8be8_1;
	wire w_dff_A_PqAu7HDC8_1;
	wire w_dff_A_pJHP8ukH6_2;
	wire w_dff_A_cElaUkoG5_2;
	wire w_dff_A_9KbYkFrg0_2;
	wire w_dff_A_W9O4aZ8K8_2;
	wire w_dff_A_vqtsjzzj7_2;
	wire w_dff_A_dAwaBqhc0_2;
	wire w_dff_A_MGXlMyfQ4_2;
	wire w_dff_A_7VL5Q9WW4_2;
	wire w_dff_A_AAaitIOj4_2;
	wire w_dff_A_Yc6PNerJ2_2;
	wire w_dff_A_4nFkwIba8_2;
	wire w_dff_A_4C3HrD6y1_2;
	wire w_dff_A_Z7fQ9pbj9_2;
	wire w_dff_A_ijIv27JT2_2;
	wire w_dff_A_kksTxhOK8_2;
	wire w_dff_A_2SGXp0oM2_2;
	wire w_dff_A_4HolBZtJ9_2;
	wire w_dff_A_edmQBWUx8_2;
	wire w_dff_A_QhwQfpfa2_2;
	wire w_dff_A_677S7Hut9_2;
	wire w_dff_A_6cJ6o5721_2;
	wire w_dff_A_273yAYLc6_2;
	wire w_dff_A_DUGoD5AN0_2;
	wire w_dff_A_xPdKTMWM8_2;
	wire w_dff_A_pqofm7Rs6_2;
	wire w_dff_A_5s3u3bZC2_2;
	wire w_dff_A_p7lWIDlr6_2;
	wire w_dff_B_8CK6fxJ17_2;
	wire w_dff_B_ICVIfdOc7_1;
	wire w_dff_B_wUIvTA2e6_1;
	wire w_dff_A_MVXiMlLm6_0;
	wire w_dff_A_2vz3W4HZ9_2;
	wire w_dff_A_B8oHIgWy0_2;
	wire w_dff_A_THdHVtNs4_0;
	wire w_dff_A_lp8KMlFN7_0;
	wire w_dff_A_jOqVUj9t0_1;
	wire w_dff_A_CgprWX050_1;
	wire w_dff_A_NUBUx68D1_2;
	wire w_dff_B_er0lYqO62_1;
	wire w_dff_B_OicV9Q9v5_1;
	wire w_dff_A_EGI21scW8_2;
	wire w_dff_A_4959dTQj2_2;
	wire w_dff_B_cNjfOzIY2_3;
	wire w_dff_B_10meFRAC4_1;
	wire w_dff_A_xKkvtONz0_1;
	wire w_dff_A_VTAY7AXp1_0;
	wire w_dff_A_deWhamyq0_0;
	wire w_dff_A_bdsLIN204_1;
	wire w_dff_A_bANAr1uV7_0;
	wire w_dff_B_cCsAviXl1_1;
	wire w_dff_B_NJxDURGC2_1;
	wire w_dff_A_gVE6PJP04_0;
	wire w_dff_A_cyAvUDdr7_2;
	wire w_dff_A_E1z9zFPw6_2;
	wire w_dff_A_MVwIv0GP9_0;
	wire w_dff_A_UwK3clxq8_1;
	wire w_dff_A_9GNBrGGm0_1;
	wire w_dff_A_MBcWebB95_2;
	wire w_dff_A_DefNt8va7_2;
	wire w_dff_A_cF42Pl3q4_2;
	wire w_dff_A_a10Qzhlk4_0;
	wire w_dff_A_CWikI4PP6_2;
	wire w_dff_B_GixM5bZd1_1;
	wire w_dff_B_SAipD6aa6_1;
	wire w_dff_A_t8GskBuY4_0;
	wire w_dff_A_n8hXXRMk4_2;
	wire w_dff_A_BgIz9GOx3_2;
	wire w_dff_A_0MVFq6Xk6_0;
	wire w_dff_A_EA789TRI2_0;
	wire w_dff_A_iAcg0cnm8_1;
	wire w_dff_A_AAuUKy352_0;
	wire w_dff_A_3ZfCYEqE6_2;
	wire w_dff_B_DBmktnb60_1;
	wire w_dff_B_TxKrL9ni2_1;
	wire w_dff_B_xxXRhAoH8_1;
	wire w_dff_B_0aMwDOAT0_1;
	wire w_dff_A_IV5zb80V7_1;
	wire w_dff_A_SCGFeEfB8_1;
	wire w_dff_A_73sXI6kO5_0;
	wire w_dff_A_AePJaZQz2_0;
	wire w_dff_A_Xc6ft2vN3_0;
	wire w_dff_A_Jut5NXeM6_0;
	wire w_dff_A_fejT3bwL7_2;
	wire w_dff_A_xZYFZW7P3_2;
	wire w_dff_A_0Pys0NPO7_1;
	wire w_dff_A_BgefP6GH8_2;
	wire w_dff_B_yoonln1B9_1;
	wire w_dff_B_kkKjk15J7_1;
	wire w_dff_B_Jr6O50Gx2_2;
	wire w_dff_A_y3avN7Kb8_0;
	wire w_dff_A_6yDkhFjs5_0;
	wire w_dff_A_3uU7QwdY8_0;
	wire w_dff_A_UkQVmX7O7_1;
	wire w_dff_B_QPKBkYa50_1;
	wire w_dff_A_dhGTwRnI9_1;
	wire w_dff_A_vPjgPKnP4_1;
	wire w_dff_A_2Rm7Aary5_1;
	wire w_dff_A_IyTfIq1V5_2;
	wire w_dff_A_pIPAGnXt1_2;
	wire w_dff_A_YXV3NzWV7_2;
	wire w_dff_A_nXUQGQHM8_0;
	wire w_dff_B_gjMBR40Q7_1;
	wire w_dff_B_A8uZyRAU6_1;
	wire w_dff_B_3kpYIH2t1_2;
	wire w_dff_A_yRJKABJA7_0;
	wire w_dff_B_Tu4nLu7q1_1;
	wire w_dff_A_kG5zjPzZ4_1;
	wire w_dff_A_NhkLcVSS1_0;
	wire w_dff_A_kFFPNKen1_0;
	wire w_dff_A_J4a6OJl35_0;
	wire w_dff_A_fI3DVBQl6_2;
	wire w_dff_A_LuvEiM885_2;
	wire w_dff_A_OUwJ3ss06_1;
	wire w_dff_A_JLvkYXd86_2;
	wire w_dff_A_FE7aTk4H4_1;
	wire w_dff_A_5yJTXELi2_2;
	wire w_dff_A_OpqiR3Vc2_0;
	wire w_dff_B_DM8NHtC44_1;
	wire w_dff_B_ERk43COR3_1;
	wire w_dff_A_csDIYLrv1_0;
	wire w_dff_A_V4NBYffl6_0;
	wire w_dff_A_uwAD3Z5m5_0;
	wire w_dff_A_bbab6R4y3_0;
	wire w_dff_A_Zv5HTxQ87_1;
	wire w_dff_A_hEVKOsBS8_1;
	wire w_dff_A_CI9viVWJ3_1;
	wire w_dff_A_jGnHbOL21_1;
	wire w_dff_A_l4IzvBjI0_1;
	wire w_dff_A_89vNui0Q7_1;
	wire w_dff_A_W4AvdWoO1_2;
	wire w_dff_A_TE3jcuxM9_2;
	wire w_dff_A_Ys9Fg2av1_2;
	wire w_dff_A_I0myafGa7_2;
	wire w_dff_A_eMdGojBb4_0;
	wire w_dff_B_ts6ctaUK2_1;
	wire w_dff_B_XmZ1eiIF8_1;
	wire w_dff_A_1cbmMLvm9_0;
	wire w_dff_A_iYvooa9B2_1;
	wire w_dff_A_NOh48NUa9_1;
	wire w_dff_A_o2DKDKw12_2;
	wire w_dff_A_i7B6QyWf9_2;
	wire w_dff_A_zw1S1KHt6_1;
	wire w_dff_A_3ks3UEbD4_1;
	wire w_dff_A_qpkDTumY8_1;
	wire w_dff_A_wrTCqjNx6_1;
	wire w_dff_A_Kn1bkS712_2;
	wire w_dff_A_iq7LmbY75_0;
	wire w_dff_A_s8E2cyjG5_0;
	wire w_dff_A_jouJrXEr8_0;
	wire w_dff_A_veECLmaf3_0;
	wire w_dff_A_SBOE7Fke9_1;
	wire w_dff_A_3V0Vm0B15_1;
	wire w_dff_A_8bvJuRvx0_1;
	wire w_dff_A_LHiAelBe1_2;
	wire w_dff_A_sD1utwgA9_2;
	wire w_dff_A_w2R1iwmP6_2;
	wire w_dff_A_tGhJKCd82_2;
	wire w_dff_A_qJLIzwhg0_1;
	wire w_dff_A_w4RxTup30_2;
	wire w_dff_A_s2t4eMkx3_0;
	wire w_dff_A_q9w38W3Z5_2;
	wire w_dff_A_SssbdDsk4_0;
	wire w_dff_A_UtUx6igc9_0;
	wire w_dff_A_RudJcVFx6_0;
	wire w_dff_A_mH82zFvq4_0;
	wire w_dff_A_MT1G3OY36_0;
	wire w_dff_A_GQbrbEcQ3_0;
	wire w_dff_A_Vil1QuFM0_0;
	wire w_dff_A_Bx9SpO2Z4_0;
	wire w_dff_A_fGb21stF5_0;
	wire w_dff_A_UFHV60qe1_0;
	wire w_dff_A_HioiWyno7_0;
	wire w_dff_A_tiqr3PDH6_1;
	wire w_dff_A_aCo5Gh4Y6_0;
	wire w_dff_A_MsqheXaF3_0;
	wire w_dff_A_hXX5za0E7_0;
	wire w_dff_A_VJssQblt5_0;
	wire w_dff_A_ARmYp1xD2_0;
	wire w_dff_A_kqWYIkrs0_0;
	wire w_dff_A_i8oAcA1P3_0;
	wire w_dff_A_nW5w3hZ52_2;
	wire w_dff_A_Hry0ZRis6_2;
	wire w_dff_A_yTLYQhWh3_2;
	wire w_dff_A_sfrbuVF69_2;
	wire w_dff_A_dGpCHngu8_2;
	wire w_dff_A_P2nNnnMx7_2;
	wire w_dff_A_3ySoJ11v1_2;
	wire w_dff_A_fRvdGumS9_2;
	wire w_dff_A_mRQKqnyj6_2;
	wire w_dff_A_wVpZ0ypX9_2;
	wire w_dff_A_yG9WEfH69_2;
	wire w_dff_A_WeqxlSju4_2;
	wire w_dff_A_v5LyskgL4_2;
	wire w_dff_A_JA6O6dTh1_2;
	wire w_dff_A_sTG3Glzy5_2;
	wire w_dff_A_GjC3orH78_2;
	wire w_dff_A_vnnaMtET6_2;
	wire w_dff_A_0C7rssIX6_2;
	wire w_dff_A_x1eHhxId0_2;
	wire w_dff_A_ZtLGQnYV7_1;
	wire w_dff_A_ZvDFzrbu4_1;
	wire w_dff_A_wiZYGcvl5_1;
	wire w_dff_A_QU304iMb2_1;
	wire w_dff_A_BQyx0Emi5_1;
	wire w_dff_A_UoNcJO6G7_1;
	wire w_dff_A_Cybi2LeB9_1;
	wire w_dff_A_RoEvyOu82_1;
	wire w_dff_A_5k0j8sKn3_1;
	wire w_dff_A_gUTMHAdq3_1;
	wire w_dff_A_yoOkNbya8_1;
	wire w_dff_A_9fe40RVz0_1;
	wire w_dff_A_zanh6Atf6_1;
	wire w_dff_A_c0KHvXL23_1;
	wire w_dff_A_L2YAXgQa0_1;
	wire w_dff_A_rLVuhbm90_1;
	wire w_dff_A_3K6GrN4X4_1;
	wire w_dff_A_iI4S3sc08_2;
	wire w_dff_A_1cobA0TI7_2;
	wire w_dff_A_Vlr5r1QO1_2;
	wire w_dff_A_XsHFxLCG5_2;
	wire w_dff_A_TfcDO0ZB1_2;
	wire w_dff_A_aA9mping5_2;
	wire w_dff_A_dMpSaAdQ9_2;
	wire w_dff_A_y2qxMShh2_2;
	wire w_dff_A_yrOUtYlm7_2;
	wire w_dff_A_3t3whZ2Y3_2;
	wire w_dff_A_dahGnmyB9_2;
	wire w_dff_A_IaEcCyU10_1;
	wire w_dff_A_zWSyWcJh3_2;
	wire w_dff_B_PaArHjYw6_2;
	wire w_dff_B_zdbVsq0K2_2;
	wire w_dff_B_VKhCWsLv7_2;
	wire w_dff_B_MeLGRvv19_2;
	wire w_dff_B_DeWhxuHb4_2;
	wire w_dff_B_hyVuRBW98_2;
	wire w_dff_B_a8R01oOk4_2;
	wire w_dff_B_ZgqPkHwa6_2;
	wire w_dff_B_0fV5U8zh0_2;
	wire w_dff_B_IH5kUP9c2_2;
	wire w_dff_B_np9OwCyc2_2;
	wire w_dff_B_lcY3qdge8_2;
	wire w_dff_B_j0zQEHMk1_2;
	wire w_dff_B_Z66bq53k5_2;
	wire w_dff_B_czvFAzS05_2;
	wire w_dff_B_4T5ih9X59_2;
	wire w_dff_B_0gAnX0VS6_2;
	wire w_dff_B_uAU7InlV9_2;
	wire w_dff_B_hDQiykh92_2;
	wire w_dff_B_leXMfk1o1_2;
	wire w_dff_B_4nDZVYd27_2;
	wire w_dff_B_z5pUiMO61_2;
	wire w_dff_B_FIxQMkhB5_2;
	wire w_dff_B_HJ0gmp534_2;
	wire w_dff_A_hWHP13Na3_2;
	wire w_dff_A_yWb9TyGp6_2;
	wire w_dff_A_3Jn64Rcv4_2;
	wire w_dff_A_fNDQtBoU9_2;
	wire w_dff_A_1oiwm1U34_2;
	wire w_dff_A_wmJ7KXU28_2;
	wire w_dff_A_g2NadnpD6_2;
	wire w_dff_A_8N7lv18q8_2;
	wire w_dff_A_QfF5VCWS8_2;
	wire w_dff_A_QB9sNRC20_2;
	wire w_dff_A_rgcB032A9_2;
	wire w_dff_A_2kXcv5EP4_2;
	wire w_dff_A_ELTcECpr2_2;
	wire w_dff_A_8lGAZe4P5_2;
	wire w_dff_A_am4IBHpH9_2;
	wire w_dff_A_Sp41L3gm8_2;
	wire w_dff_A_qNgS8F394_2;
	wire w_dff_A_iqdgmdfO7_2;
	wire w_dff_A_RXfGAZfL9_2;
	wire w_dff_A_hCrS64lY0_2;
	wire w_dff_A_NICqD9a91_2;
	wire w_dff_A_KJlkTg9i7_2;
	wire w_dff_A_QGAAvwDb4_2;
	wire w_dff_A_tU1ov6fD1_0;
	wire w_dff_A_dJhWGqua3_0;
	wire w_dff_A_bISyXt4b5_0;
	wire w_dff_A_F6sRyIu06_0;
	wire w_dff_A_nKozoKNF7_0;
	wire w_dff_A_4g0sPfdQ3_0;
	wire w_dff_A_hMi0SqkB0_0;
	wire w_dff_A_uom8rbJg7_0;
	wire w_dff_A_i8ENp6xF8_0;
	wire w_dff_A_ntJvPZ7t5_0;
	wire w_dff_A_7w2cHXdd8_0;
	wire w_dff_A_nTlvFufY7_0;
	wire w_dff_A_7SJP1IDB0_0;
	wire w_dff_A_IcvyyfZm0_0;
	wire w_dff_A_nAywAc2n6_0;
	wire w_dff_A_y8EKslp71_0;
	wire w_dff_A_7M70bVjP4_1;
	wire w_dff_A_6zeM2juR0_1;
	wire w_dff_A_W0s8m6Dw6_1;
	wire w_dff_A_J80eq6C52_1;
	wire w_dff_A_M0S4rPp63_1;
	wire w_dff_A_tD29lgOE2_1;
	wire w_dff_A_1ZsIH3Tu9_1;
	wire w_dff_A_N89QNPHs4_1;
	wire w_dff_A_BweG7lt36_1;
	wire w_dff_A_55ArJU9c9_1;
	wire w_dff_A_7BUQRPrB0_1;
	wire w_dff_A_okV472fm6_1;
	wire w_dff_A_ogv3lNCr0_0;
	wire w_dff_A_oV1uorzV5_0;
	wire w_dff_A_6ezAHKGO0_0;
	wire w_dff_A_mfQVpu4y6_0;
	wire w_dff_A_5XrMRjGZ9_0;
	wire w_dff_A_QSIOIiXg8_0;
	wire w_dff_A_IIrlkdnD9_0;
	wire w_dff_A_kJYYLnkk0_0;
	wire w_dff_A_2KhvLaZT1_0;
	wire w_dff_A_zknnBtXH6_0;
	wire w_dff_A_163sYPsF4_0;
	wire w_dff_A_3llhc7En7_0;
	wire w_dff_A_KXjDxkDD7_0;
	wire w_dff_A_XiqObUWP7_0;
	wire w_dff_A_StNbPVKd8_0;
	wire w_dff_A_p2lsyuUi2_0;
	wire w_dff_A_qM7m0ZwE3_0;
	wire w_dff_A_asfHprWw6_0;
	wire w_dff_A_rA6LTo662_0;
	wire w_dff_A_LTWHRYH73_0;
	wire w_dff_A_hpVaIVDg6_0;
	wire w_dff_A_eJ703AlT6_0;
	wire w_dff_A_glrjwNps1_0;
	wire w_dff_A_HkFzjxmf8_0;
	wire w_dff_A_Vfdcr69x0_0;
	wire w_dff_A_NZDPOgPm2_1;
	wire w_dff_A_ZyfyjtQ58_0;
	wire w_dff_A_xUsn0j0M1_0;
	wire w_dff_A_ZemeG7VO1_0;
	wire w_dff_A_8hP8GLcc6_0;
	wire w_dff_A_7IS9ToZb2_0;
	wire w_dff_A_kZamQdsq8_0;
	wire w_dff_A_8wx8sm6s8_0;
	wire w_dff_A_gJV0myzi1_0;
	wire w_dff_A_a6epFmHE2_0;
	wire w_dff_A_zZxeVQxT1_0;
	wire w_dff_A_uocuKcTo0_0;
	wire w_dff_A_ZVEl00kN4_0;
	wire w_dff_A_LHnIaVZn7_0;
	wire w_dff_A_I6zfqJfT1_0;
	wire w_dff_A_C9SvRgiR4_0;
	wire w_dff_A_krBIP1DP1_0;
	wire w_dff_A_6WtM4WiY7_0;
	wire w_dff_A_NnYtvDvs9_0;
	wire w_dff_A_n6teTyJa8_0;
	wire w_dff_A_yztdqtqJ6_0;
	wire w_dff_A_IrafUO6r5_0;
	wire w_dff_A_wExJG9WZ4_0;
	wire w_dff_A_YYGfBxpA6_0;
	wire w_dff_A_SMhb38CL7_0;
	wire w_dff_A_BZ2jFIPl8_0;
	wire w_dff_A_8SfPKRXf1_1;
	wire w_dff_A_LlC6qNoO9_0;
	wire w_dff_A_HqNFrRRt4_0;
	wire w_dff_A_yvZDnkZh2_0;
	wire w_dff_A_9t4xMM6Z8_0;
	wire w_dff_A_Kt8rJOXo9_0;
	wire w_dff_A_Jm1bYKHC5_0;
	wire w_dff_A_mqLiPzgE7_0;
	wire w_dff_A_14G34L1o0_0;
	wire w_dff_A_GZudCT3D3_0;
	wire w_dff_A_c7FLgvys3_0;
	wire w_dff_A_uUgr2uCA1_0;
	wire w_dff_A_eScK2o8I6_0;
	wire w_dff_A_XRUibDmM2_0;
	wire w_dff_A_j7RkDJ4j3_0;
	wire w_dff_A_K3BJWmvQ8_0;
	wire w_dff_A_xK8qpfUj2_0;
	wire w_dff_A_6rP5M31f8_0;
	wire w_dff_A_K2sNMlaT7_0;
	wire w_dff_A_E2qBVsr26_0;
	wire w_dff_A_jXxYKFhQ5_0;
	wire w_dff_A_QFhRrDUe9_0;
	wire w_dff_A_8tPwtVAx0_0;
	wire w_dff_A_0R8davIi8_0;
	wire w_dff_A_6WpTeIW55_0;
	wire w_dff_A_mZUjYeH90_0;
	wire w_dff_A_V5AYLoBR3_1;
	wire w_dff_A_cK7bFte06_0;
	wire w_dff_A_bEIyv3CV0_0;
	wire w_dff_A_SvnUPLiK5_0;
	wire w_dff_A_dIn0g7Gl1_0;
	wire w_dff_A_y6CqniDP2_0;
	wire w_dff_A_HP5Z9x121_0;
	wire w_dff_A_o2wPvOQr5_0;
	wire w_dff_A_vjXx6cGV7_0;
	wire w_dff_A_WC6WBIOd7_0;
	wire w_dff_A_O6BdxDHu8_0;
	wire w_dff_A_MLAbcBpK0_0;
	wire w_dff_A_JTrxyZqm5_0;
	wire w_dff_A_DMMdjmFM7_0;
	wire w_dff_A_8L68Y3DV7_0;
	wire w_dff_A_dYTMK3Rp9_0;
	wire w_dff_A_MmXwx7mn3_0;
	wire w_dff_A_yf4b1s9v4_0;
	wire w_dff_A_VHClbzyf3_0;
	wire w_dff_A_MMnRv6694_0;
	wire w_dff_A_pH0bz1jt6_0;
	wire w_dff_A_JXJiJwas5_0;
	wire w_dff_A_6Z1n3bKR4_0;
	wire w_dff_A_4bxgWxj34_0;
	wire w_dff_A_hRtNzZgp9_0;
	wire w_dff_A_3L9jc5wg9_1;
	wire w_dff_A_vEKKRsGd7_0;
	wire w_dff_A_Wkh1cTgd0_0;
	wire w_dff_A_V4AD3w623_0;
	wire w_dff_A_sEdITJI15_0;
	wire w_dff_A_KZojZsK95_0;
	wire w_dff_A_ME6bXSDU7_0;
	wire w_dff_A_372uKjDW6_0;
	wire w_dff_A_4ATw8BM06_0;
	wire w_dff_A_LFNjDd318_0;
	wire w_dff_A_dTxQpufI2_0;
	wire w_dff_A_chJmIE7D0_0;
	wire w_dff_A_8BImmkCY5_0;
	wire w_dff_A_ORCTvjGy5_0;
	wire w_dff_A_onIyKMjz1_0;
	wire w_dff_A_o5ccFe7B0_0;
	wire w_dff_A_IrbJFcy67_0;
	wire w_dff_A_Foi1f5FH9_0;
	wire w_dff_A_7hkYaTDD6_0;
	wire w_dff_A_cfovHEdE4_0;
	wire w_dff_A_t7dss5vg3_0;
	wire w_dff_A_Q2ijlehy2_0;
	wire w_dff_A_rkNQ3HYH3_0;
	wire w_dff_A_IBfoackQ7_0;
	wire w_dff_A_jEwMu9cN4_0;
	wire w_dff_A_p2Avj4Ok5_1;
	wire w_dff_A_PvkSDAGn4_0;
	wire w_dff_A_jGTmYm5E9_0;
	wire w_dff_A_B0ncpjQE1_0;
	wire w_dff_A_nqm7mEeW9_0;
	wire w_dff_A_17ehKx0R9_0;
	wire w_dff_A_Z4ZJUrZ52_0;
	wire w_dff_A_yUxjOSnH4_0;
	wire w_dff_A_56DkgF726_0;
	wire w_dff_A_LbyzknDR6_0;
	wire w_dff_A_hR7vLwDL6_0;
	wire w_dff_A_xRInDINj1_0;
	wire w_dff_A_5A3jwpn55_0;
	wire w_dff_A_LOftf9yg5_0;
	wire w_dff_A_s7wkQ6Hz1_0;
	wire w_dff_A_T6XvvGTH9_0;
	wire w_dff_A_eoPN4I3c5_0;
	wire w_dff_A_TBM72KVF3_0;
	wire w_dff_A_nBhgTgC88_0;
	wire w_dff_A_r6YHjFLu7_0;
	wire w_dff_A_wpx4jmy09_0;
	wire w_dff_A_HyFR7HTm2_0;
	wire w_dff_A_3tnw3Zr51_0;
	wire w_dff_A_O6WhPV7G1_0;
	wire w_dff_A_WLQln4x22_0;
	wire w_dff_A_dz8Ft8Lm5_1;
	wire w_dff_A_JSDsn5kA7_0;
	wire w_dff_A_YLSG9GNz5_0;
	wire w_dff_A_7F0UaqCH5_0;
	wire w_dff_A_zatp2yiT1_0;
	wire w_dff_A_9B6YAoJi9_0;
	wire w_dff_A_czAkkZYJ4_0;
	wire w_dff_A_aVAMlb7C0_0;
	wire w_dff_A_1g9QgtAa1_0;
	wire w_dff_A_mvp3yt8P4_0;
	wire w_dff_A_5P0tR7P50_0;
	wire w_dff_A_4IeFLxLt1_0;
	wire w_dff_A_71tAsMEu9_0;
	wire w_dff_A_CU8oE03d1_0;
	wire w_dff_A_U0PMj6Bc6_0;
	wire w_dff_A_fOQcQTle7_0;
	wire w_dff_A_6aSEVCcj7_0;
	wire w_dff_A_1PUlN2gS0_0;
	wire w_dff_A_2oKprsdt4_0;
	wire w_dff_A_Ob9qltBQ5_0;
	wire w_dff_A_bQC6ySv07_0;
	wire w_dff_A_QkI0g3Hq5_0;
	wire w_dff_A_sIJyTJWJ8_0;
	wire w_dff_A_UTG4Somq5_0;
	wire w_dff_A_6VZBjnF37_0;
	wire w_dff_A_s2RVKcId6_1;
	wire w_dff_A_tATd9YJz8_0;
	wire w_dff_A_6NubUDHE1_0;
	wire w_dff_A_rUf7Mbw61_0;
	wire w_dff_A_uXM7UcU86_0;
	wire w_dff_A_MrQoWlc55_0;
	wire w_dff_A_UudJEs7V8_0;
	wire w_dff_A_hNPCBG3p9_0;
	wire w_dff_A_VqGfESAb5_0;
	wire w_dff_A_ngFzu4ba5_0;
	wire w_dff_A_DmAxYJDc0_0;
	wire w_dff_A_f2DKxFer1_0;
	wire w_dff_A_5oPoE5Ht3_0;
	wire w_dff_A_EaksyIGh6_0;
	wire w_dff_A_h5j7dwQU7_0;
	wire w_dff_A_h1g6MR6z3_0;
	wire w_dff_A_UbL2vsxL3_0;
	wire w_dff_A_BIH5wCk30_0;
	wire w_dff_A_GXcw6zQD2_0;
	wire w_dff_A_uSOO17m51_0;
	wire w_dff_A_XpFWsEE17_0;
	wire w_dff_A_DPFy6FRM4_0;
	wire w_dff_A_tbLsQrJW9_0;
	wire w_dff_A_DAXSPrcr1_0;
	wire w_dff_A_Y1x8Pt0Y4_0;
	wire w_dff_A_kcOoDOTs8_1;
	wire w_dff_A_2DVT02543_0;
	wire w_dff_A_ZQqX4Lkn5_0;
	wire w_dff_A_Jq4xC4fU9_0;
	wire w_dff_A_b6NtChoc4_0;
	wire w_dff_A_XHXmZc7H3_0;
	wire w_dff_A_zPnjCGk42_0;
	wire w_dff_A_7zeZws047_0;
	wire w_dff_A_fsXqtNpA0_0;
	wire w_dff_A_gAnHUW3u7_0;
	wire w_dff_A_DmeUCcow5_0;
	wire w_dff_A_2Mu281sQ3_0;
	wire w_dff_A_DbcBmpOW3_0;
	wire w_dff_A_OjVjaU0Q9_0;
	wire w_dff_A_jecQuqw36_0;
	wire w_dff_A_HqIFvB276_0;
	wire w_dff_A_tE3NpQdt1_0;
	wire w_dff_A_PwQp3b3Q5_0;
	wire w_dff_A_k9yQ1RNl7_0;
	wire w_dff_A_Wm0gzxWe2_0;
	wire w_dff_A_t2Gusbyd9_0;
	wire w_dff_A_fwRGXway1_0;
	wire w_dff_A_ZH1r2eSj6_0;
	wire w_dff_A_50evll2s5_0;
	wire w_dff_A_4LggUN8F5_0;
	wire w_dff_A_hDMD60wB6_1;
	wire w_dff_A_BCtwA5XO2_0;
	wire w_dff_A_L27Jgo6W3_0;
	wire w_dff_A_lKDAFeTZ4_0;
	wire w_dff_A_B36YSzB13_0;
	wire w_dff_A_lOCQ4mXJ2_0;
	wire w_dff_A_zSFbqrLS6_0;
	wire w_dff_A_dqrBGxKs8_0;
	wire w_dff_A_Yqw9PheB4_0;
	wire w_dff_A_Azg8u7so6_0;
	wire w_dff_A_dDD3VMX70_0;
	wire w_dff_A_PzNrCIkj1_0;
	wire w_dff_A_oAPoFMC03_0;
	wire w_dff_A_UVrokZLl8_0;
	wire w_dff_A_HJ6gta4a1_0;
	wire w_dff_A_Mn9BlPf28_0;
	wire w_dff_A_0jTRirf47_0;
	wire w_dff_A_PWTnVoTw6_0;
	wire w_dff_A_o3iDkmJj6_0;
	wire w_dff_A_pvYdX6aT8_0;
	wire w_dff_A_DwpUNVel8_0;
	wire w_dff_A_leUowjKv2_0;
	wire w_dff_A_7XJp0Tgc2_0;
	wire w_dff_A_9AvTUtQC3_0;
	wire w_dff_A_QAO211s71_0;
	wire w_dff_A_u0F4vmwG6_1;
	wire w_dff_A_9iV7etma1_0;
	wire w_dff_A_xR1CDCiH4_0;
	wire w_dff_A_9mkTrHY12_0;
	wire w_dff_A_gWCQvCZl6_0;
	wire w_dff_A_GyU4E6NA8_0;
	wire w_dff_A_w4vdD8iZ6_0;
	wire w_dff_A_6vkkNFpX1_0;
	wire w_dff_A_aZqO8c5F7_0;
	wire w_dff_A_XLjHdiyH6_0;
	wire w_dff_A_jGsUjMvm1_0;
	wire w_dff_A_J2f4JC6P8_0;
	wire w_dff_A_HI9stvvD5_0;
	wire w_dff_A_eUrec72X5_0;
	wire w_dff_A_g1yjhV022_0;
	wire w_dff_A_IcadDF6t1_0;
	wire w_dff_A_Q2HGDxci3_0;
	wire w_dff_A_TzHKWsDc2_0;
	wire w_dff_A_XeaXkH5p3_0;
	wire w_dff_A_1KQqB91M8_0;
	wire w_dff_A_m0ZEIDAx1_0;
	wire w_dff_A_nhN7O2Om4_0;
	wire w_dff_A_CBXEhqr40_0;
	wire w_dff_A_NlbAecwD3_0;
	wire w_dff_A_y4uxC6nd1_0;
	wire w_dff_A_vV76YNP35_1;
	wire w_dff_A_lziMPqTj0_0;
	wire w_dff_A_5F9DPMfw0_0;
	wire w_dff_A_EBWMsjJe0_0;
	wire w_dff_A_VT7EMWLc4_0;
	wire w_dff_A_O5E1qDJi2_0;
	wire w_dff_A_8qnEGAZC1_0;
	wire w_dff_A_MQsAG5lq6_0;
	wire w_dff_A_c6Vsn3OW2_0;
	wire w_dff_A_YL86j1d33_0;
	wire w_dff_A_0jrsovDC6_0;
	wire w_dff_A_L6iIM8QM3_0;
	wire w_dff_A_tKlmUtQS7_0;
	wire w_dff_A_BpTMQnj98_0;
	wire w_dff_A_KHT5ooBw7_0;
	wire w_dff_A_sx1oMZqH1_0;
	wire w_dff_A_fci6eniY4_0;
	wire w_dff_A_YU9eLELf6_0;
	wire w_dff_A_T0WxmrKV1_0;
	wire w_dff_A_XgHagHai4_0;
	wire w_dff_A_vuCuXbVo5_0;
	wire w_dff_A_Cs3hiT9K0_0;
	wire w_dff_A_1nJyn9qk6_0;
	wire w_dff_A_uD2KJBVk3_0;
	wire w_dff_A_UOomnUKF3_0;
	wire w_dff_A_GlKmi3Mx5_2;
	wire w_dff_A_FoF28rke4_0;
	wire w_dff_A_kc5WQBGy2_0;
	wire w_dff_A_LmKqX8Mj9_0;
	wire w_dff_A_pGUnQGn94_0;
	wire w_dff_A_EZegEoFd7_0;
	wire w_dff_A_GfQslj0o0_0;
	wire w_dff_A_XIFE8IBm9_0;
	wire w_dff_A_tIPzgF7l9_0;
	wire w_dff_A_wJC5mJQg8_0;
	wire w_dff_A_b5NydUYV6_0;
	wire w_dff_A_wIskXDYU2_0;
	wire w_dff_A_AjpMm4TS2_0;
	wire w_dff_A_l9i4VvN49_0;
	wire w_dff_A_85K5QOOH6_0;
	wire w_dff_A_fF3m1NiH2_0;
	wire w_dff_A_Z7MDiG8V9_0;
	wire w_dff_A_nR1ZUh5U2_0;
	wire w_dff_A_baKoa0Ig6_0;
	wire w_dff_A_Yzmkfj7N6_0;
	wire w_dff_A_mQCLBEtB0_0;
	wire w_dff_A_Z5MYojyL4_0;
	wire w_dff_A_qHp9fiAq2_0;
	wire w_dff_A_ASFLD3OY1_0;
	wire w_dff_A_b2dglj631_0;
	wire w_dff_A_xyLwOATF7_1;
	wire w_dff_A_eNvCPr9i4_0;
	wire w_dff_A_8oRD8j3h4_0;
	wire w_dff_A_ibAyT6ij0_0;
	wire w_dff_A_vxof0kK68_0;
	wire w_dff_A_x7g8EHZc3_0;
	wire w_dff_A_pKxM4MRV2_0;
	wire w_dff_A_nkl7Wo2H5_0;
	wire w_dff_A_hpLOQV0C5_0;
	wire w_dff_A_Nyq8fd0V1_0;
	wire w_dff_A_WsWtyNfe4_0;
	wire w_dff_A_10sVEysO1_0;
	wire w_dff_A_MKWPLyAp1_0;
	wire w_dff_A_WkFiKJKM7_0;
	wire w_dff_A_JhzUAlvL1_0;
	wire w_dff_A_mGg9XuzS9_0;
	wire w_dff_A_6sR7H9hy4_0;
	wire w_dff_A_CrtDy2rj8_0;
	wire w_dff_A_Ng0nP9Pz8_0;
	wire w_dff_A_m95qoQ9p1_0;
	wire w_dff_A_dh9HbEoW8_0;
	wire w_dff_A_hCYOeZJR5_0;
	wire w_dff_A_tJcdIU2f8_0;
	wire w_dff_A_RW53ZOK86_0;
	wire w_dff_A_ZsI0AaUQ5_0;
	wire w_dff_A_H8rH6ICZ3_1;
	wire w_dff_A_nOtMmBbK9_0;
	wire w_dff_A_OtbwNwYB6_0;
	wire w_dff_A_2khSAweJ4_0;
	wire w_dff_A_dyVsIhlv3_0;
	wire w_dff_A_oDPWNfAa3_0;
	wire w_dff_A_gQMW51AI1_0;
	wire w_dff_A_HPcxssCH8_0;
	wire w_dff_A_bMNuzee73_0;
	wire w_dff_A_musNaZm99_0;
	wire w_dff_A_I9eo0zv08_0;
	wire w_dff_A_Y9g00JQ24_0;
	wire w_dff_A_z0mWXjxE3_0;
	wire w_dff_A_CImKJKok4_0;
	wire w_dff_A_VaSZNCj75_0;
	wire w_dff_A_WHcI2w6f8_0;
	wire w_dff_A_GqwwfeYl1_0;
	wire w_dff_A_TRjxx3Lq9_0;
	wire w_dff_A_cZa8AnBW9_0;
	wire w_dff_A_pqDlsAvc7_0;
	wire w_dff_A_kzcHeqM82_0;
	wire w_dff_A_goHCHCuz3_0;
	wire w_dff_A_CdK5SyKL2_0;
	wire w_dff_A_akEnMZTu2_0;
	wire w_dff_A_bRKOe4wl6_0;
	wire w_dff_A_Xusarkiy7_1;
	wire w_dff_A_hrBPrJ3k4_0;
	wire w_dff_A_aaPWOIIu8_0;
	wire w_dff_A_werb8YnI4_0;
	wire w_dff_A_mYezHKSE6_0;
	wire w_dff_A_vvgoF3Lp1_0;
	wire w_dff_A_S60DZFUn0_0;
	wire w_dff_A_IoM7ebW96_0;
	wire w_dff_A_hNOh6rtH1_0;
	wire w_dff_A_YuxYtkDv0_0;
	wire w_dff_A_JmG6gYIf4_0;
	wire w_dff_A_MRP53ePZ5_0;
	wire w_dff_A_BzvS1uvv3_0;
	wire w_dff_A_icKZ0k6n3_0;
	wire w_dff_A_LNQpHKrV1_0;
	wire w_dff_A_GZAhTFVz3_0;
	wire w_dff_A_uNsXvIKA0_0;
	wire w_dff_A_8IQsyxm79_0;
	wire w_dff_A_3qu5WyOD6_0;
	wire w_dff_A_JcX9TJoS0_0;
	wire w_dff_A_i4BeRQuP4_0;
	wire w_dff_A_JRIPggxw5_0;
	wire w_dff_A_4QOfRiWB4_0;
	wire w_dff_A_X1jHTkfH9_0;
	wire w_dff_A_MxEkLznI2_0;
	wire w_dff_A_pmLPKsfd4_1;
	wire w_dff_A_suFphxG97_0;
	wire w_dff_A_lOTGBhQ59_0;
	wire w_dff_A_lgW7zxz77_0;
	wire w_dff_A_1wEnSzqF5_0;
	wire w_dff_A_CeNpf4TS3_0;
	wire w_dff_A_J1Bvu7ZZ0_0;
	wire w_dff_A_g5njZi7L8_0;
	wire w_dff_A_ik80OX237_0;
	wire w_dff_A_PLfaf77S1_0;
	wire w_dff_A_9GR8uVrz7_0;
	wire w_dff_A_1KyUeUtZ2_0;
	wire w_dff_A_euXqnPdk9_0;
	wire w_dff_A_RQvKvLTV1_0;
	wire w_dff_A_zEYokS6w1_0;
	wire w_dff_A_iyIxatti8_0;
	wire w_dff_A_gTrcipWg2_0;
	wire w_dff_A_ixKCXnwZ3_0;
	wire w_dff_A_MVwL5dF71_0;
	wire w_dff_A_BjiThJyY8_0;
	wire w_dff_A_GyPH7zPK1_0;
	wire w_dff_A_0nUYBNEz8_0;
	wire w_dff_A_D8IQuX735_0;
	wire w_dff_A_BnMfACOa4_0;
	wire w_dff_A_pAd7P8mQ8_0;
	wire w_dff_A_RYNJc9DE7_2;
	wire w_dff_A_K0Gp274N1_0;
	wire w_dff_A_MPy72eiW4_0;
	wire w_dff_A_LvSJJ4uN7_0;
	wire w_dff_A_PicTrorG4_0;
	wire w_dff_A_bJmFwyF66_0;
	wire w_dff_A_kK0Iytzo9_0;
	wire w_dff_A_7HUGsfuw3_0;
	wire w_dff_A_zoTMS6al2_0;
	wire w_dff_A_5Tikg5i43_0;
	wire w_dff_A_eYqwXIcD6_0;
	wire w_dff_A_Am5Z8qri4_0;
	wire w_dff_A_k5QkWKsX2_0;
	wire w_dff_A_nQB22ICq8_0;
	wire w_dff_A_ErQaohi93_0;
	wire w_dff_A_DF8xFxXn1_0;
	wire w_dff_A_PBoDfIGd6_0;
	wire w_dff_A_BuOOO1na7_0;
	wire w_dff_A_V9mPnqth7_0;
	wire w_dff_A_44bQQigm3_0;
	wire w_dff_A_gdzRynCj5_0;
	wire w_dff_A_1EuwGAOE6_0;
	wire w_dff_A_V2pChiko1_0;
	wire w_dff_A_xMavVPiU9_0;
	wire w_dff_A_usp0TRLn9_0;
	wire w_dff_A_yXw8OWlh0_2;
	wire w_dff_A_6jWmU8vg1_0;
	wire w_dff_A_bF6tchFU2_0;
	wire w_dff_A_9iJdGgTj6_0;
	wire w_dff_A_8LdQTxzS7_0;
	wire w_dff_A_0eLUeaiW9_0;
	wire w_dff_A_Ceyaryv07_0;
	wire w_dff_A_Ubbj64qM5_0;
	wire w_dff_A_79uyTPsg2_0;
	wire w_dff_A_GZgr1Pdm2_0;
	wire w_dff_A_MYrR1AiH1_0;
	wire w_dff_A_LYcd1Qc95_0;
	wire w_dff_A_sUhUoX0H5_0;
	wire w_dff_A_ad0N5twf0_0;
	wire w_dff_A_sVhWGoNO2_0;
	wire w_dff_A_QY3ozO4E2_0;
	wire w_dff_A_V66hZaVM6_0;
	wire w_dff_A_r2go5Xi55_0;
	wire w_dff_A_2gr0sy7n1_0;
	wire w_dff_A_xLR3sFmw6_0;
	wire w_dff_A_BwEWsH041_0;
	wire w_dff_A_H1QIBT7v8_0;
	wire w_dff_A_mJNNPMaw0_0;
	wire w_dff_A_ve09drHw3_0;
	wire w_dff_A_QrS0w1hc9_2;
	wire w_dff_A_v0R7cT3A2_0;
	wire w_dff_A_qnf4sQky6_0;
	wire w_dff_A_Kb0UWdzr6_0;
	wire w_dff_A_fmGQrk6p4_0;
	wire w_dff_A_v0Xaxmzn5_0;
	wire w_dff_A_DeGVkzQk2_0;
	wire w_dff_A_JVSjm7gC7_0;
	wire w_dff_A_wV771ojw7_0;
	wire w_dff_A_cauunzu24_0;
	wire w_dff_A_eFetDvas1_0;
	wire w_dff_A_Vf76mOl43_0;
	wire w_dff_A_WsAz6DbW6_0;
	wire w_dff_A_7XNVSPDS9_0;
	wire w_dff_A_DFSGgDvy2_0;
	wire w_dff_A_BLedsIhK0_0;
	wire w_dff_A_inFCm5b98_0;
	wire w_dff_A_L10plpC43_0;
	wire w_dff_A_Xx8EgXT19_0;
	wire w_dff_A_STM1ZcFU2_0;
	wire w_dff_A_jc5rUWe24_0;
	wire w_dff_A_NiTD0wdi5_0;
	wire w_dff_A_dDlBSleA7_0;
	wire w_dff_A_khFgEntc2_0;
	wire w_dff_A_LSvafEGP1_1;
	wire w_dff_A_YQv15aTr9_0;
	wire w_dff_A_8OrmuQq63_0;
	wire w_dff_A_hSOEr44i2_0;
	wire w_dff_A_yIVB93VL1_0;
	wire w_dff_A_SKCuxarp6_0;
	wire w_dff_A_1wO0lHia8_0;
	wire w_dff_A_BLaFsW7q7_0;
	wire w_dff_A_TeVbRD8X4_0;
	wire w_dff_A_IUuOibde7_0;
	wire w_dff_A_mR1x8Z0y0_0;
	wire w_dff_A_Au8xFoSx1_0;
	wire w_dff_A_LnQZhrv18_0;
	wire w_dff_A_5VicGoJH0_0;
	wire w_dff_A_tkRk2qtZ4_0;
	wire w_dff_A_Sk04FQP71_0;
	wire w_dff_A_30QA9Yde5_0;
	wire w_dff_A_1XokZoC53_0;
	wire w_dff_A_WT4Cl0NM0_0;
	wire w_dff_A_CcE17NJy0_0;
	wire w_dff_A_OsiQXJQo9_0;
	wire w_dff_A_zXP9mh6c1_0;
	wire w_dff_A_qCE6IiTW5_0;
	wire w_dff_A_ekCsCMJB8_0;
	wire w_dff_A_01NRIr0n5_1;
	wire w_dff_A_T0KCI0Br3_0;
	wire w_dff_A_JIqo6lAF5_0;
	wire w_dff_A_HAOSnCqu0_0;
	wire w_dff_A_lJbLgato8_0;
	wire w_dff_A_QgPb02XW2_0;
	wire w_dff_A_bPrzDpx25_0;
	wire w_dff_A_HZEVDcEq9_0;
	wire w_dff_A_tKnN1aix3_0;
	wire w_dff_A_oJlQzsHm4_0;
	wire w_dff_A_quIB8Cb39_0;
	wire w_dff_A_pazK6p7m6_0;
	wire w_dff_A_zXBOdUVV8_0;
	wire w_dff_A_y4fXJ6dx2_0;
	wire w_dff_A_C3vpuTLt0_0;
	wire w_dff_A_l9MOsyXH0_0;
	wire w_dff_A_mnOm5jxk3_0;
	wire w_dff_A_vDZEMzXW4_0;
	wire w_dff_A_2EtgvZrm1_0;
	wire w_dff_A_GjBOM3mV0_0;
	wire w_dff_A_2jLytp936_0;
	wire w_dff_A_Vz8iP4Hr0_0;
	wire w_dff_A_o86rQLXx9_0;
	wire w_dff_A_UB2FYZMP8_0;
	wire w_dff_A_YnJ1tJzk2_0;
	wire w_dff_A_pRwshihh7_0;
	wire w_dff_A_BnnZ8yRL2_1;
	wire w_dff_A_1EQsAT453_0;
	wire w_dff_A_QCNTUIu25_0;
	wire w_dff_A_oWBKiZVp8_0;
	wire w_dff_A_BYFycvHY6_0;
	wire w_dff_A_V0026irJ5_0;
	wire w_dff_A_jdCPur5z9_0;
	wire w_dff_A_XhD97bkX3_0;
	wire w_dff_A_piGLnmpn8_0;
	wire w_dff_A_Kgi0SGy95_0;
	wire w_dff_A_SJYGjweE5_0;
	wire w_dff_A_VYbr9uzs3_0;
	wire w_dff_A_PKCIma1I4_0;
	wire w_dff_A_lqCx9CMD5_0;
	wire w_dff_A_bjgza2BL2_0;
	wire w_dff_A_IEAjRMro8_0;
	wire w_dff_A_Ba2UnCps9_0;
	wire w_dff_A_YElEShL60_0;
	wire w_dff_A_dFSTVjYn2_0;
	wire w_dff_A_AYz8fusT0_0;
	wire w_dff_A_TY7K932o2_0;
	wire w_dff_A_CPD6Efrp8_0;
	wire w_dff_A_hpefC9ae1_0;
	wire w_dff_A_0zIeliN32_0;
	wire w_dff_A_ZDS7IzTM6_0;
	wire w_dff_A_DaHO4N7T2_0;
	wire w_dff_A_Lh3AxbIW3_1;
	wire w_dff_A_ImlrT97C3_0;
	wire w_dff_A_SCYZ5BkE7_0;
	wire w_dff_A_qSgrRCIc4_0;
	wire w_dff_A_a5YIGvpc7_0;
	wire w_dff_A_NxQ5Bbpb9_0;
	wire w_dff_A_MmIiKObK2_0;
	wire w_dff_A_avlQfnii2_0;
	wire w_dff_A_iAhmQvPT1_0;
	wire w_dff_A_Tq5F952u4_0;
	wire w_dff_A_mSSI74u32_0;
	wire w_dff_A_qF0E5Cdl7_0;
	wire w_dff_A_W6LOQr1W9_0;
	wire w_dff_A_b3VcpK2n0_0;
	wire w_dff_A_b3CdZCJ50_0;
	wire w_dff_A_mroB81Cj5_0;
	wire w_dff_A_nhVwgCod1_0;
	wire w_dff_A_UNby12XJ2_0;
	wire w_dff_A_VFkGOxeG0_0;
	wire w_dff_A_f71d8YOX5_0;
	wire w_dff_A_d4u2VCCL9_0;
	wire w_dff_A_ks86YvjL4_0;
	wire w_dff_A_6ASGuWde8_0;
	wire w_dff_A_wugflzAV7_0;
	wire w_dff_A_QZ6xIBF59_0;
	wire w_dff_A_MPSd35nE2_0;
	wire w_dff_A_J5XkOm3N6_1;
	wire w_dff_A_myOflQGG3_0;
	wire w_dff_A_FOQwnEDt2_0;
	wire w_dff_A_xs7nUafR2_0;
	wire w_dff_A_88eakqhA7_0;
	wire w_dff_A_lpmANb3k2_0;
	wire w_dff_A_so9lmTyb8_0;
	wire w_dff_A_Z5jBZ53w8_0;
	wire w_dff_A_uT4eruv50_0;
	wire w_dff_A_1EBmzuvu6_0;
	wire w_dff_A_Pjrjv0Rx3_0;
	wire w_dff_A_gDSMpamd6_0;
	wire w_dff_A_YGtJp68q5_0;
	wire w_dff_A_fTe3itQ76_0;
	wire w_dff_A_BTTZFMKc3_0;
	wire w_dff_A_BXhTVqsY9_0;
	wire w_dff_A_mMNki7lP1_0;
	wire w_dff_A_MvxY6Iah0_0;
	wire w_dff_A_FRRRTgtz2_0;
	wire w_dff_A_wxG9MtEi6_0;
	wire w_dff_A_y74yrhsH9_0;
	wire w_dff_A_lwAAOZ8e9_0;
	wire w_dff_A_HuiI7CWG0_0;
	wire w_dff_A_2mFCOca89_0;
	wire w_dff_A_ta3JEm181_0;
	wire w_dff_A_yKxRKaqF8_0;
	wire w_dff_A_DyvXlmRo5_1;
	wire w_dff_A_tLXdturw1_0;
	wire w_dff_A_3hodUwyi5_0;
	wire w_dff_A_ZwlNl2494_0;
	wire w_dff_A_sn0h8oOY2_0;
	wire w_dff_A_QnKjVoYS2_0;
	wire w_dff_A_ORld5hr40_0;
	wire w_dff_A_wffqNnzy9_0;
	wire w_dff_A_knN7M2ZI9_0;
	wire w_dff_A_h2AQVlxP7_0;
	wire w_dff_A_3EPTT3hI8_0;
	wire w_dff_A_V0VRm04v5_0;
	wire w_dff_A_WyWQ5rCf3_0;
	wire w_dff_A_xFHIHZRf1_0;
	wire w_dff_A_09qoeox29_0;
	wire w_dff_A_6EqdFl8v8_0;
	wire w_dff_A_qW2PdEIs8_0;
	wire w_dff_A_1b82hlNA8_0;
	wire w_dff_A_tO5O59357_0;
	wire w_dff_A_ZHPBeITe7_0;
	wire w_dff_A_h04npl922_0;
	wire w_dff_A_jfQCWTci0_0;
	wire w_dff_A_Rgsvvq4d7_0;
	wire w_dff_A_fMpYah1y6_0;
	wire w_dff_A_9vSzsBJX8_0;
	wire w_dff_A_bEhDIrq66_0;
	wire w_dff_A_nvgG7fE58_1;
	wire w_dff_A_N3hu5bC12_0;
	wire w_dff_A_KPOicwMq5_0;
	wire w_dff_A_OCKymEXB1_0;
	wire w_dff_A_ucdGveD86_0;
	wire w_dff_A_bXE7E3GN4_0;
	wire w_dff_A_Txy0aA5D9_0;
	wire w_dff_A_2U2VnnSb3_0;
	wire w_dff_A_zFLFNVP43_0;
	wire w_dff_A_452iNvR68_0;
	wire w_dff_A_Qm3VKH1a3_0;
	wire w_dff_A_MRj4ygRT9_0;
	wire w_dff_A_fiZrchch4_0;
	wire w_dff_A_3kIM8ibh6_0;
	wire w_dff_A_AVLyIPyA1_0;
	wire w_dff_A_S0LhnmTs7_0;
	wire w_dff_A_3dkV0ct89_0;
	wire w_dff_A_JWLLaUqB4_0;
	wire w_dff_A_4JLrEYuS9_0;
	wire w_dff_A_Lrjjx16v3_0;
	wire w_dff_A_IeJ6ryVi6_0;
	wire w_dff_A_ZJFFcWwp6_0;
	wire w_dff_A_SZ3yWRj41_0;
	wire w_dff_A_J6zAg7lC5_0;
	wire w_dff_A_cNWvPRCi8_0;
	wire w_dff_A_dtpCUlzB5_2;
	wire w_dff_A_5Eh2GO9F2_0;
	wire w_dff_A_3suHmsej5_0;
	wire w_dff_A_ksBNEb8g7_0;
	wire w_dff_A_tJNslEAo5_0;
	wire w_dff_A_niiULae75_0;
	wire w_dff_A_ZexcCbco4_0;
	wire w_dff_A_c8l4WoxB8_0;
	wire w_dff_A_QXxPXL2C1_0;
	wire w_dff_A_1LWx9mDd8_0;
	wire w_dff_A_DfgroJEz6_0;
	wire w_dff_A_OXozIfOx0_0;
	wire w_dff_A_DQsS3MaV7_0;
	wire w_dff_A_3C9QpG8a6_0;
	wire w_dff_A_J4ZLPBDi8_0;
	wire w_dff_A_EjPBXT596_0;
	wire w_dff_A_LnaG41ak7_0;
	wire w_dff_A_Q1XUl7WF2_0;
	wire w_dff_A_kvcSJhn63_0;
	wire w_dff_A_3YyCJeWj3_0;
	wire w_dff_A_tpObOz4f2_0;
	wire w_dff_A_CGMV944R3_0;
	wire w_dff_A_akhxLudq6_0;
	wire w_dff_A_Wkcf8uO35_2;
	wire w_dff_A_nVQkj7KY2_0;
	wire w_dff_A_XrIZB1W39_0;
	wire w_dff_A_2RAvaipf5_0;
	wire w_dff_A_L5qTC1Tz5_0;
	wire w_dff_A_tkrlteuN8_0;
	wire w_dff_A_PjIRoYcv5_0;
	wire w_dff_A_PXAjyjue2_0;
	wire w_dff_A_bQtcwnco8_0;
	wire w_dff_A_1xfS7pJG0_0;
	wire w_dff_A_iC1qYZAI9_0;
	wire w_dff_A_RvJEUfeB5_0;
	wire w_dff_A_4ECh9uD13_0;
	wire w_dff_A_i0x8pCV67_0;
	wire w_dff_A_azu69xyF1_0;
	wire w_dff_A_ge2p8Y7j5_0;
	wire w_dff_A_WtbNT1NZ1_0;
	wire w_dff_A_uRqDqbqv6_0;
	wire w_dff_A_AmbNLimM7_0;
	wire w_dff_A_7Jy3zYRO0_0;
	wire w_dff_A_H2s2XOom2_0;
	wire w_dff_A_61abACHB9_0;
	wire w_dff_A_BJ2ZWDW55_0;
	wire w_dff_A_4AybJTNt1_0;
	wire w_dff_A_cVuHOXky3_1;
	wire w_dff_A_oNXFHuPE6_0;
	wire w_dff_A_MkyAEXfM5_0;
	wire w_dff_A_wbm6SpU57_0;
	wire w_dff_A_GEQHmbgQ0_0;
	wire w_dff_A_oaA25qda8_0;
	wire w_dff_A_DaZs9uKh2_0;
	wire w_dff_A_U9NpTuD58_0;
	wire w_dff_A_zK3GZtg69_0;
	wire w_dff_A_4WNNsVql6_0;
	wire w_dff_A_m5YsQizm3_0;
	wire w_dff_A_l7ISEKSu8_0;
	wire w_dff_A_OtdfU1Pj1_0;
	wire w_dff_A_mue8HkJW4_0;
	wire w_dff_A_yqGfCi8F5_0;
	wire w_dff_A_uoUYJGq24_0;
	wire w_dff_A_acO3YlaP4_0;
	wire w_dff_A_ctM2dYWb6_0;
	wire w_dff_A_GRk5yzkq3_0;
	wire w_dff_A_pYljRpJX2_0;
	wire w_dff_A_o3rCca0V4_0;
	wire w_dff_A_FSbSJtL34_0;
	wire w_dff_A_3xBXSfal7_0;
	wire w_dff_A_gUEw0R6k7_0;
	wire w_dff_A_nFWSTKc02_0;
	wire w_dff_A_MpCT5jKU2_0;
	wire w_dff_A_iX0YGi3V0_1;
	wire w_dff_A_uPMFkgiK0_0;
	wire w_dff_A_Rwek7Y8j2_0;
	wire w_dff_A_5ZD3t5XU0_0;
	wire w_dff_A_ZcMaCXiN7_0;
	wire w_dff_A_nack7WKD7_0;
	wire w_dff_A_rF0C75SO9_0;
	wire w_dff_A_CdkQSd1x3_0;
	wire w_dff_A_4OuDYHoh8_0;
	wire w_dff_A_zSZ3q2jN6_0;
	wire w_dff_A_nhVGhS5G2_0;
	wire w_dff_A_jFQXGY4W0_0;
	wire w_dff_A_OxYy07Nz4_0;
	wire w_dff_A_TuZ54p393_0;
	wire w_dff_A_Q3b3frXR6_0;
	wire w_dff_A_73WZmY8t9_0;
	wire w_dff_A_XTVnZnC67_0;
	wire w_dff_A_jmRj4X3v9_0;
	wire w_dff_A_9OS8w7ag8_0;
	wire w_dff_A_vGK8cV1X4_0;
	wire w_dff_A_io1MLuGf8_0;
	wire w_dff_A_ZT50cMaF1_0;
	wire w_dff_A_KnGPUazE0_0;
	wire w_dff_A_fsCTBilZ2_0;
	wire w_dff_A_LRw983rV2_0;
	wire w_dff_A_JNJ830t24_0;
	wire w_dff_A_FzCJlgsD0_1;
	wire w_dff_A_dmqgJdYK4_0;
	wire w_dff_A_2QQJPzUD8_0;
	wire w_dff_A_uE8It0L95_0;
	wire w_dff_A_s7llUBAs4_0;
	wire w_dff_A_AEfoKEYj8_0;
	wire w_dff_A_Pr9QXGPp1_0;
	wire w_dff_A_kRCdJWnq7_0;
	wire w_dff_A_ajdiTEoj5_0;
	wire w_dff_A_GB3TSgUR4_0;
	wire w_dff_A_swdJ8koh8_0;
	wire w_dff_A_ilnXyLGe7_0;
	wire w_dff_A_gIZtQk7r6_0;
	wire w_dff_A_lWwMjQo36_0;
	wire w_dff_A_O7eCQBbb2_0;
	wire w_dff_A_xTEGNqlA5_0;
	wire w_dff_A_uUZh42M83_0;
	wire w_dff_A_AerjJxn55_0;
	wire w_dff_A_YktjNGhO8_0;
	wire w_dff_A_68Z6taLk3_0;
	wire w_dff_A_A1Uvqxpg2_0;
	wire w_dff_A_fmycmVYt0_0;
	wire w_dff_A_rz93mtqB6_0;
	wire w_dff_A_U97nWb8Q7_0;
	wire w_dff_A_DZWc4IE48_0;
	wire w_dff_A_Gub68ra10_0;
	wire w_dff_A_PtVtnSx29_1;
	wire w_dff_A_fkZ5MK9m3_0;
	wire w_dff_A_B0Cr4v9X6_0;
	wire w_dff_A_1N53pl6k6_0;
	wire w_dff_A_Gr0SZmbl3_0;
	wire w_dff_A_408Dljpk0_0;
	wire w_dff_A_SPm3Y7r77_0;
	wire w_dff_A_1CJ1iw1z4_0;
	wire w_dff_A_jFjpe5yW0_0;
	wire w_dff_A_9S70EFcj0_0;
	wire w_dff_A_1qU3BK194_0;
	wire w_dff_A_uLbWhK2j7_0;
	wire w_dff_A_ZCHuBAbr1_0;
	wire w_dff_A_JJOFqeDL5_0;
	wire w_dff_A_fWbAKXRj8_0;
	wire w_dff_A_7JKVIISd5_0;
	wire w_dff_A_QF20WGQF1_0;
	wire w_dff_A_jZt2ctxf9_0;
	wire w_dff_A_BNRjKA9u5_0;
	wire w_dff_A_xUHN77XW6_0;
	wire w_dff_A_NheApzMZ7_0;
	wire w_dff_A_5lhFs6f03_0;
	wire w_dff_A_A1jHp2lW7_0;
	wire w_dff_A_UOzIG68G1_0;
	wire w_dff_A_YBjhP92M7_0;
	wire w_dff_A_M83qPGpc7_0;
	wire w_dff_A_bcmCouej6_1;
	wire w_dff_A_0jyR4lP04_0;
	wire w_dff_A_gmKLIKev7_0;
	wire w_dff_A_YTLtTUxd2_0;
	wire w_dff_A_Ap2Le9Ou7_0;
	wire w_dff_A_h6xfBR1K8_0;
	wire w_dff_A_Wb3ghfmV5_0;
	wire w_dff_A_iQxqBBte5_0;
	wire w_dff_A_I7gTCGFI3_0;
	wire w_dff_A_B294Nn5X4_0;
	wire w_dff_A_ZZyr5BFy2_0;
	wire w_dff_A_DbAQnLHE3_0;
	wire w_dff_A_1wRDI2Yz8_0;
	wire w_dff_A_Y8fz1tEs0_0;
	wire w_dff_A_3rMu2ikH3_0;
	wire w_dff_A_a1lF7Oo46_0;
	wire w_dff_A_hVQg70iO8_0;
	wire w_dff_A_XMlaIjP11_0;
	wire w_dff_A_mU4Kjgeb7_0;
	wire w_dff_A_A92cHQJO4_0;
	wire w_dff_A_4PJwjazR5_0;
	wire w_dff_A_VcHY7LOQ3_0;
	wire w_dff_A_jYKzQ7hn3_0;
	wire w_dff_A_HA24eAHg9_0;
	wire w_dff_A_ndTmpEou3_0;
	wire w_dff_A_dFui7bHY3_0;
	wire w_dff_A_iy5NfA8p1_1;
	wire w_dff_A_WnizSuDl5_0;
	wire w_dff_A_jqAJpjmk0_0;
	wire w_dff_A_5ShCLTLz2_0;
	wire w_dff_A_edl3g0y16_0;
	wire w_dff_A_F23wutM29_0;
	wire w_dff_A_fCjuVgCk7_0;
	wire w_dff_A_Wd3bmiyF4_0;
	wire w_dff_A_NlFev7FY6_0;
	wire w_dff_A_r32K8gd08_0;
	wire w_dff_A_2fj1LZui6_0;
	wire w_dff_A_eMI39XM03_0;
	wire w_dff_A_J7yENLvS0_0;
	wire w_dff_A_njOTFXhz2_0;
	wire w_dff_A_JmBlk7qa4_0;
	wire w_dff_A_xbHFW4oG3_0;
	wire w_dff_A_cXk9f2aw7_0;
	wire w_dff_A_XF12hza79_0;
	wire w_dff_A_Pc8IWniA8_0;
	wire w_dff_A_HvLlkRkW3_0;
	wire w_dff_A_kTiCZk2C8_0;
	wire w_dff_A_WOCNomxj0_0;
	wire w_dff_A_xQE2EbN35_0;
	wire w_dff_A_HB62ZxmB8_0;
	wire w_dff_A_QnMQBUgv3_0;
	wire w_dff_A_DH3gqMbd6_2;
	wire w_dff_A_CmMV3JTc6_0;
	wire w_dff_A_4sAg2tf42_0;
	wire w_dff_A_6TuJaMJU3_0;
	wire w_dff_A_SJq7rbG52_0;
	wire w_dff_A_zR1ClXM12_0;
	wire w_dff_A_7QSNtk6c3_0;
	wire w_dff_A_0RIaDIDr2_0;
	wire w_dff_A_3ye0t4pd9_0;
	wire w_dff_A_pjsRGaGO3_0;
	wire w_dff_A_0GUbYCaN5_0;
	wire w_dff_A_g5no8Ieu0_0;
	wire w_dff_A_ovphpXRL6_0;
	wire w_dff_A_w0Ofdea05_0;
	wire w_dff_A_7O0dIBuK8_0;
	wire w_dff_A_hoZIqJxi2_0;
	wire w_dff_A_BWLc6lkr4_0;
	wire w_dff_A_n32w4r7Q7_0;
	wire w_dff_A_QqrZRL7u9_0;
	wire w_dff_A_VovFy6QC9_0;
	wire w_dff_A_KDKlOLjc6_0;
	wire w_dff_A_eCjy2DTL6_0;
	wire w_dff_A_4mIO0Omj6_2;
	wire w_dff_A_42libba56_0;
	wire w_dff_A_ICpZIEjr2_0;
	wire w_dff_A_myNgd3T04_0;
	wire w_dff_A_LECBlswP2_0;
	wire w_dff_A_i4mh0IRK1_0;
	wire w_dff_A_8dB4UqgM0_0;
	wire w_dff_A_SaT244wW4_0;
	wire w_dff_A_d5BNXPMn3_0;
	wire w_dff_A_7ifcpMUb6_0;
	wire w_dff_A_7yauADEk4_0;
	wire w_dff_A_hFthHK0W8_0;
	wire w_dff_A_ZqPdSjTr7_0;
	wire w_dff_A_vnJaF1wA2_0;
	wire w_dff_A_OTwb2gWc9_0;
	wire w_dff_A_ByzumVJf7_0;
	wire w_dff_A_3sFOxuGv5_0;
	wire w_dff_A_eDC7b2zl8_0;
	wire w_dff_A_7mLwgt455_0;
	wire w_dff_A_x2eiRihv3_0;
	wire w_dff_A_mYNzs6kq8_0;
	wire w_dff_A_vw4iXDjF4_0;
	wire w_dff_A_2Em61F4H5_2;
	wire w_dff_A_xiUguW3E1_0;
	wire w_dff_A_40YbK28V7_0;
	wire w_dff_A_x7HYhBMb5_0;
	wire w_dff_A_pgxDGr2p1_0;
	wire w_dff_A_6sFEABCs6_0;
	wire w_dff_A_O85zz5Yw9_0;
	wire w_dff_A_aNcka0Tf5_0;
	wire w_dff_A_FyvA1L460_0;
	wire w_dff_A_btOH0xby6_0;
	wire w_dff_A_tgUyvSwV0_0;
	wire w_dff_A_V6IfQMwu5_0;
	wire w_dff_A_DrrzWTJH3_0;
	wire w_dff_A_1Ds676rs7_0;
	wire w_dff_A_8NHAdBE15_0;
	wire w_dff_A_9ngVJhHv1_0;
	wire w_dff_A_ggvqsBZ73_0;
	wire w_dff_A_f1588PC83_0;
	wire w_dff_A_sHuAMXua5_0;
	wire w_dff_A_iG8A7Kc61_0;
	wire w_dff_A_sYQDF5Ft9_0;
	wire w_dff_A_4jhY0ozW6_0;
	wire w_dff_A_A5LKfscm0_2;
	wire w_dff_A_8UVu3P1o4_0;
	wire w_dff_A_IgtMrHSH0_0;
	wire w_dff_A_eQ7ytHvT5_0;
	wire w_dff_A_BvcAjru20_0;
	wire w_dff_A_Tqws9Go98_0;
	wire w_dff_A_dO9ENwZc2_0;
	wire w_dff_A_BsssJlFj5_0;
	wire w_dff_A_WvTHqim74_0;
	wire w_dff_A_nvkX9kGY8_0;
	wire w_dff_A_Obspi6Qb8_0;
	wire w_dff_A_Nar49g3h6_0;
	wire w_dff_A_zvRhIdJR3_0;
	wire w_dff_A_SFGJmORD5_0;
	wire w_dff_A_cJtRRpLy3_0;
	wire w_dff_A_DGuOGsEF6_0;
	wire w_dff_A_zT3UutYA1_0;
	wire w_dff_A_YIwsOfxn3_0;
	wire w_dff_A_0ZjIJTIx7_0;
	wire w_dff_A_wGrbOC296_0;
	wire w_dff_A_xp30hxAN5_0;
	wire w_dff_A_lIQFrxW29_0;
	wire w_dff_A_NbbBuFK88_0;
	wire w_dff_A_Dmxui67i6_2;
	wire w_dff_A_x9gktYI57_0;
	wire w_dff_A_mVo6lrbu5_0;
	wire w_dff_A_JkoDpI2e9_0;
	wire w_dff_A_mxCGr4qK7_0;
	wire w_dff_A_Z5KuMd7A3_0;
	wire w_dff_A_jqUCwjqE2_0;
	wire w_dff_A_KdDENeJl7_0;
	wire w_dff_A_GrJflWi90_0;
	wire w_dff_A_w5EN2PPQ6_0;
	wire w_dff_A_fzftObhP6_0;
	wire w_dff_A_2dgtgsxt5_0;
	wire w_dff_A_8hesfdpX0_0;
	wire w_dff_A_FCsUu0T63_0;
	wire w_dff_A_BbL73qQO2_0;
	wire w_dff_A_6xhh7bEr9_0;
	wire w_dff_A_o5NfWBeA1_0;
	wire w_dff_A_FZ1sBM308_0;
	wire w_dff_A_rcd1sCUV5_0;
	wire w_dff_A_rDNfw0bc1_0;
	wire w_dff_A_fKR6z7ZD4_0;
	wire w_dff_A_HfINcbMs5_2;
	wire w_dff_A_NjjlIWWp7_0;
	wire w_dff_A_wLhg0KgC0_0;
	wire w_dff_A_M5ihDUVK3_0;
	wire w_dff_A_uyJTWQvZ5_0;
	wire w_dff_A_Q6myFDG04_0;
	wire w_dff_A_J1IczByK7_0;
	wire w_dff_A_JDQLBS9Q9_0;
	wire w_dff_A_IFH4fHVJ4_0;
	wire w_dff_A_XdVlqxEw6_0;
	wire w_dff_A_yPvTAhhl9_0;
	wire w_dff_A_yFrkmDoC2_0;
	wire w_dff_A_Gpofob8w1_0;
	wire w_dff_A_8IqI5o9d3_0;
	wire w_dff_A_JY65UEty4_0;
	wire w_dff_A_mWIv4CyH7_0;
	wire w_dff_A_JL5VW8MT2_0;
	wire w_dff_A_MajAAWAF6_0;
	wire w_dff_A_zvTHwCxX2_0;
	wire w_dff_A_bf9cG4Uh4_0;
	wire w_dff_A_XBBAZAtX5_0;
	wire w_dff_A_tqTmAX2J9_2;
	wire w_dff_A_FbKda17C0_0;
	wire w_dff_A_vy1dXzfE3_0;
	wire w_dff_A_GwgnK8Ip5_0;
	wire w_dff_A_KBcoGBz02_0;
	wire w_dff_A_4tPiuj820_0;
	wire w_dff_A_c38XK2fk1_0;
	wire w_dff_A_nGzWbQt52_0;
	wire w_dff_A_oJAor8DH0_0;
	wire w_dff_A_cmJn8vqh7_0;
	wire w_dff_A_dOlrK4WA8_0;
	wire w_dff_A_E9yatNKt3_0;
	wire w_dff_A_3gHNAW3k5_0;
	wire w_dff_A_dTjKujKg0_0;
	wire w_dff_A_ZnhYaYrQ4_0;
	wire w_dff_A_vAwl76YB2_0;
	wire w_dff_A_V9f7g9746_0;
	wire w_dff_A_XlSktFXb4_0;
	wire w_dff_A_qIno74EG6_0;
	wire w_dff_A_sPYnRjJ17_0;
	wire w_dff_A_1mtzjYA46_0;
	wire w_dff_A_q4HuDZnG7_2;
	wire w_dff_A_TWZc9Xtm3_0;
	wire w_dff_A_Rx6lPAWf1_0;
	wire w_dff_A_VIBZPs6z8_0;
	wire w_dff_A_MKzonvyp8_0;
	wire w_dff_A_5MHi83Gz0_0;
	wire w_dff_A_53XiVxZg0_0;
	wire w_dff_A_Kmxau93S9_0;
	wire w_dff_A_nGzfsclY7_0;
	wire w_dff_A_T1cJwZ1b2_0;
	wire w_dff_A_iJIqBvhn6_0;
	wire w_dff_A_HgjWojgE0_0;
	wire w_dff_A_XwsWGQLh1_0;
	wire w_dff_A_avTfQtX47_0;
	wire w_dff_A_CdzOsXks1_0;
	wire w_dff_A_0pycos278_0;
	wire w_dff_A_yWTR9anx7_0;
	wire w_dff_A_REVqGbwf5_0;
	wire w_dff_A_tmagXIk38_0;
	wire w_dff_A_LmZjFiPI6_0;
	wire w_dff_A_U8gfVIhp5_0;
	wire w_dff_A_heVA6OvF9_2;
	wire w_dff_A_t8mItqJ92_0;
	wire w_dff_A_vosmfmve7_0;
	wire w_dff_A_mdYMnQ570_0;
	wire w_dff_A_F6s3PHqc5_0;
	wire w_dff_A_xceauyHw8_0;
	wire w_dff_A_3VmWHgRi8_0;
	wire w_dff_A_N5nTT7Wf7_0;
	wire w_dff_A_EAuFS8nH9_0;
	wire w_dff_A_PfbEqwEC2_0;
	wire w_dff_A_yMf15lEb7_0;
	wire w_dff_A_0czaHG583_0;
	wire w_dff_A_NOk9F1RR3_0;
	wire w_dff_A_4hbYQgSX9_0;
	wire w_dff_A_74pB983h9_0;
	wire w_dff_A_jUnLpZRw1_0;
	wire w_dff_A_JdlXYvSK0_0;
	wire w_dff_A_98gOsWEt3_2;
	wire w_dff_A_B0OFEQIp4_0;
	wire w_dff_A_pZowCQg91_0;
	wire w_dff_A_JxmTd9VK4_0;
	wire w_dff_A_KDWIDx9X5_0;
	wire w_dff_A_NO8x4lF96_0;
	wire w_dff_A_LHnw3tqh2_0;
	wire w_dff_A_dFRJKTIY3_0;
	wire w_dff_A_jjWsjl0j0_0;
	wire w_dff_A_JSZIaNST4_0;
	wire w_dff_A_JGkX3g258_0;
	wire w_dff_A_p3EM4PfW2_0;
	wire w_dff_A_lk1kbily6_0;
	wire w_dff_A_fFQcJEqi8_0;
	wire w_dff_A_3aJOuQ8I3_0;
	wire w_dff_A_fnbxQkNv3_0;
	wire w_dff_A_W5jSJ4eO7_0;
	wire w_dff_A_a8FPstR07_2;
	wire w_dff_A_Y76EPjOu1_0;
	wire w_dff_A_4sK39zaX6_0;
	wire w_dff_A_SmKTwjui8_0;
	wire w_dff_A_QCPup3ZN5_0;
	wire w_dff_A_lsmNFQ1N9_0;
	wire w_dff_A_Tf6AjAa66_0;
	wire w_dff_A_cnKgS36D6_0;
	wire w_dff_A_4qn29nex5_0;
	wire w_dff_A_hkN3Y5US3_0;
	wire w_dff_A_YUuRk3Tf1_0;
	wire w_dff_A_54INVPiv3_0;
	wire w_dff_A_J4ZslZdO7_0;
	wire w_dff_A_TptopMkg5_0;
	wire w_dff_A_oXwBPp741_0;
	wire w_dff_A_iLCWaaL96_2;
	wire w_dff_A_0RjeCt8U2_0;
	wire w_dff_A_6FaBFqCk0_0;
	wire w_dff_A_usc74RgE8_0;
	wire w_dff_A_4ihPoDKK8_0;
	wire w_dff_A_14ba03835_0;
	wire w_dff_A_KYCdHPsg0_0;
	wire w_dff_A_UBujfgeH7_0;
	wire w_dff_A_pYNG3d568_0;
	wire w_dff_A_Cv7jV60I6_0;
	wire w_dff_A_b6iYVehc4_0;
	wire w_dff_A_N1ZFTzWl2_0;
	wire w_dff_A_IHL1tGRu8_0;
	wire w_dff_A_0twmngdc0_0;
	wire w_dff_A_5zaUQwQ88_0;
	wire w_dff_A_9IYrsimw1_0;
	wire w_dff_A_AAXedV3U9_0;
	wire w_dff_A_Y2JNsu3g3_2;
	wire w_dff_A_vUBCUwcC5_0;
	wire w_dff_A_QYMabMA04_0;
	wire w_dff_A_Fp0HoExl9_0;
	wire w_dff_A_jw9xzuQn0_0;
	wire w_dff_A_V9msACep6_0;
	wire w_dff_A_s5Ti432w4_0;
	wire w_dff_A_HSgIQdQZ1_0;
	wire w_dff_A_pyUPLJAW7_0;
	wire w_dff_A_upNVlbE39_0;
	wire w_dff_A_dwo7mkOJ1_0;
	wire w_dff_A_WpLPLNHG7_0;
	wire w_dff_A_rd5YAnOU5_0;
	wire w_dff_A_xV3QuAoi6_0;
	wire w_dff_A_tZrQMKIb6_0;
	wire w_dff_A_omVFdhgg0_0;
	wire w_dff_A_LW7XAMXs6_0;
	wire w_dff_A_ILZVgwZy8_2;
	wire w_dff_A_PQlf6GMd2_0;
	wire w_dff_A_Mwot3wa29_0;
	wire w_dff_A_JRabvF5G4_0;
	wire w_dff_A_vW0Eyizj4_0;
	wire w_dff_A_6d9O58BP4_0;
	wire w_dff_A_50drFKUZ0_0;
	wire w_dff_A_mszFQdJs6_0;
	wire w_dff_A_Ew9C0ilo8_0;
	wire w_dff_A_tkIG6ZIX9_0;
	wire w_dff_A_DhgW0GUa4_0;
	wire w_dff_A_SRsdwpud5_0;
	wire w_dff_A_jQSc5UrE5_0;
	wire w_dff_A_2YFZ3K0t2_0;
	wire w_dff_A_OLiViglB7_0;
	wire w_dff_A_1v2VW66l6_1;
	wire w_dff_A_Ira4mwGl4_0;
	wire w_dff_A_KjHPCE8R2_0;
	wire w_dff_A_b0b7x1cQ1_0;
	wire w_dff_A_5thJ7mpQ6_0;
	wire w_dff_A_nzSsYxOa7_0;
	wire w_dff_A_wnSh4jIM9_0;
	wire w_dff_A_oIUb7XkB7_0;
	wire w_dff_A_Iy5RohBW1_0;
	wire w_dff_A_fagOtbE00_0;
	wire w_dff_A_gPSsUOWk0_0;
	wire w_dff_A_REk4iN1w1_0;
	wire w_dff_A_Xgayo0G98_0;
	wire w_dff_A_isge7Zwi0_0;
	wire w_dff_A_GXS5mcUB4_0;
	wire w_dff_A_SGceFbLn2_0;
	wire w_dff_A_dEhmY3mf2_0;
	wire w_dff_A_AXx7NQnL9_0;
	wire w_dff_A_lkZKFyOo3_0;
	wire w_dff_A_QUueERQi5_0;
	wire w_dff_A_aZNTGliG6_0;
	wire w_dff_A_nMfNfIJ88_1;
	wire w_dff_A_aia6tAyR1_0;
	wire w_dff_A_3ZJMfTKa0_0;
	wire w_dff_A_BqJGGqG23_0;
	wire w_dff_A_QQOReGzZ6_0;
	wire w_dff_A_vTtqk7PU2_0;
	wire w_dff_A_xHaQ98584_0;
	wire w_dff_A_tax63zYn0_0;
	wire w_dff_A_OuQBdFaA4_0;
	wire w_dff_A_vAKZcCet1_0;
	wire w_dff_A_iMuTPVJI2_0;
	wire w_dff_A_KboyahDh7_0;
	wire w_dff_A_rtJ5pmdO1_0;
	wire w_dff_A_gcRAxrbN8_0;
	wire w_dff_A_g4C1Kh1p8_0;
	wire w_dff_A_KEATrYLB3_0;
	wire w_dff_A_U7D0JHqV1_0;
	wire w_dff_A_PTdGLIUt1_0;
	wire w_dff_A_dLTj28wV3_0;
	wire w_dff_A_RuScc4Lg1_0;
	wire w_dff_A_oLmbBiYt2_0;
	wire w_dff_A_oGRN7NsA0_2;
	wire w_dff_A_HCSwzBOJ5_0;
	wire w_dff_A_fN03UcI28_0;
	wire w_dff_A_htbl4Arh5_0;
	wire w_dff_A_qikab3oX8_0;
	wire w_dff_A_WWLLOsE74_0;
	wire w_dff_A_k5QyiATD7_0;
	wire w_dff_A_T3WfK5JS4_0;
	wire w_dff_A_HgUm4Wfm5_0;
	wire w_dff_A_PIB0gAmo8_0;
	wire w_dff_A_iUmsnd2u0_0;
	wire w_dff_A_LgYyAyff6_0;
	wire w_dff_A_M3kaUjHO8_2;
	wire w_dff_A_od9CFQac1_0;
	wire w_dff_A_nX9SPcRE3_0;
	wire w_dff_A_2n5ueYHb8_0;
	wire w_dff_A_JBAlqqQD3_0;
	wire w_dff_A_K7Le8zQa2_0;
	wire w_dff_A_QDFoqplF2_0;
	wire w_dff_A_LgqFVPYY7_0;
	wire w_dff_A_xfAN4HbR0_0;
	wire w_dff_A_Pwbwltpl3_0;
	wire w_dff_A_3Lxeulcw4_0;
	wire w_dff_A_ikhfFZ2b7_0;
	wire w_dff_A_k90aNcvw2_2;
	wire w_dff_A_kcddZhXl0_0;
	wire w_dff_A_oMly865h2_0;
	wire w_dff_A_RBF4SVrQ4_0;
	wire w_dff_A_6lx0kjh80_0;
	wire w_dff_A_u5xUUkRd4_0;
	wire w_dff_A_K4xHwNqM3_0;
	wire w_dff_A_OAC6sqxy9_0;
	wire w_dff_A_XUAquFlY9_0;
	wire w_dff_A_9mtx4GaW5_0;
	wire w_dff_A_zkJmKRXE4_0;
	wire w_dff_A_WfnNI6MR0_0;
	wire w_dff_A_zku3LX0f7_2;
	wire w_dff_A_JkRydBe31_0;
	wire w_dff_A_NvZPpkuv9_0;
	wire w_dff_A_icD3YL3o2_0;
	wire w_dff_A_sEqoTvZ97_0;
	wire w_dff_A_k3vzIK5t7_0;
	wire w_dff_A_UWZkjq8E7_0;
	wire w_dff_A_9oCgsZoT0_0;
	wire w_dff_A_ibtOhAEi6_0;
	wire w_dff_A_daXPEoIA9_0;
	wire w_dff_A_cPbU9v4P8_0;
	wire w_dff_A_EXRv7mO53_0;
	wire w_dff_A_q1tFT8lp8_1;
	wire w_dff_A_P44sLowh2_0;
	wire w_dff_A_eOPioVdF8_0;
	wire w_dff_A_Jlrw9ktA1_0;
	wire w_dff_A_8F5vlDrx5_0;
	wire w_dff_A_h3laRYog9_0;
	wire w_dff_A_MdCieRsr0_0;
	wire w_dff_A_r547ROxf8_0;
	wire w_dff_A_P4DjLPsY8_0;
	wire w_dff_A_aO3i0XEV3_0;
	wire w_dff_A_95qOkN0M0_0;
	wire w_dff_A_N84C3P9f2_0;
	wire w_dff_A_QkcwueYH6_0;
	wire w_dff_A_WrAYzFoG5_0;
	wire w_dff_A_8mFoipho1_0;
	wire w_dff_A_wHXTGEO89_0;
	wire w_dff_A_2zND4OGL2_0;
	wire w_dff_A_9PbdJEEm1_0;
	wire w_dff_A_2wxje0ys9_0;
	wire w_dff_A_AYO72yhU1_1;
	wire w_dff_A_XywcEaJ49_0;
	wire w_dff_A_s3udFBJ43_0;
	wire w_dff_A_dLPwlqWd0_0;
	wire w_dff_A_jWz8xjl01_0;
	wire w_dff_A_C6ioL0HG9_0;
	wire w_dff_A_hCN6uBsO0_0;
	wire w_dff_A_Uggwwmxa7_0;
	wire w_dff_A_zkIZLCHX2_0;
	wire w_dff_A_W9cNDRiU2_0;
	wire w_dff_A_yFpiiRYf5_0;
	wire w_dff_A_TxhCSyiI7_0;
	wire w_dff_A_FAHrZ0hJ6_0;
	wire w_dff_A_FPqdRuPV2_0;
	wire w_dff_A_o2HfYUVo3_0;
	wire w_dff_A_W5WvkQ2T0_0;
	wire w_dff_A_2L03ORBx3_0;
	wire w_dff_A_zh0iCaZF6_0;
	wire w_dff_A_KfJFor9N7_1;
	wire w_dff_A_NN2k55lL9_0;
	wire w_dff_A_86GzOnGp2_0;
	wire w_dff_A_DZ79gRgf2_0;
	wire w_dff_A_3bLamFKY7_0;
	wire w_dff_A_5tuFy5kO6_0;
	wire w_dff_A_PHA3kwzM4_0;
	wire w_dff_A_wGvFnnkW3_0;
	wire w_dff_A_Tj2n1Jc63_0;
	wire w_dff_A_r2RlglYq9_0;
	wire w_dff_A_4CCKekpJ0_0;
	wire w_dff_A_FZGNVepn3_0;
	wire w_dff_A_JOfdidDz0_0;
	wire w_dff_A_UschAx5w8_0;
	wire w_dff_A_HOSW48Mq9_0;
	wire w_dff_A_wBkrJtwD1_0;
	wire w_dff_A_iAVYVYPd1_0;
	wire w_dff_A_Mhtqgaee2_0;
	wire w_dff_A_i69PVv1d1_1;
	wire w_dff_A_wOAaABEf7_0;
	wire w_dff_A_AktMmHI74_0;
	wire w_dff_A_HO4H0c6d9_0;
	wire w_dff_A_vaiEItOd4_0;
	wire w_dff_A_EIDCrBcL4_0;
	wire w_dff_A_G45eVPtF1_0;
	wire w_dff_A_sV8pytjm1_2;
	wire w_dff_A_GTZ7yswP5_0;
	wire w_dff_A_smA2jgin7_0;
	wire w_dff_A_hEttIOEH2_0;
	wire w_dff_A_NoHJkvAX1_0;
	wire w_dff_A_VRsR3txa9_0;
	wire w_dff_A_JD23QiaJ4_0;
	wire w_dff_A_gDWVLIAC8_0;
	wire w_dff_A_O4Px5IhQ0_0;
	wire w_dff_A_Gfh6MIS83_0;
	wire w_dff_A_yiJOh81W8_0;
	wire w_dff_A_rxWA0Uww8_0;
	wire w_dff_A_KXxs2KMA3_0;
	wire w_dff_A_NlauAOvK1_0;
	wire w_dff_A_2PY7AmP71_0;
	wire w_dff_A_0wXNdgG84_1;
	wire w_dff_A_Fv9CePF61_0;
	wire w_dff_A_9RJTjqSd6_0;
	wire w_dff_A_8mtJ3sJX8_0;
	wire w_dff_A_23Sc72Pf9_0;
	wire w_dff_A_nKORoGTi4_0;
	wire w_dff_A_Z1vwV1fg9_0;
	wire w_dff_A_6JVam7T38_0;
	wire w_dff_A_kqO1J8L91_0;
	wire w_dff_A_aC3wlJzx9_0;
	wire w_dff_A_SdBkTOWy7_0;
	wire w_dff_A_1RqMgdJa1_0;
	wire w_dff_A_wKLlrNjI5_1;
	wire w_dff_A_MFK3SxBP6_0;
	wire w_dff_A_s4jXqwk55_0;
	wire w_dff_A_n5q1i7FY9_0;
	wire w_dff_A_ep3x9ehP5_0;
	wire w_dff_A_018dXP870_0;
	wire w_dff_A_7Ldy8DOA4_0;
	wire w_dff_A_4OqwkNU43_0;
	wire w_dff_A_OQiNf4Hy1_0;
	wire w_dff_A_KXP7UABL8_0;
	wire w_dff_A_Gqcwnt1r2_0;
	wire w_dff_A_GJf4cJnl9_0;
	wire w_dff_A_uhzzR6FF1_0;
	wire w_dff_A_Bv7ww4kQ5_0;
	wire w_dff_A_ScVFdJA46_1;
	wire w_dff_A_8lyBC1yo0_0;
	wire w_dff_A_3rpw4Cls2_0;
	wire w_dff_A_IwlMcOzk0_0;
	wire w_dff_A_DQZ2UmjT7_0;
	wire w_dff_A_a4mf9Bax4_0;
	wire w_dff_A_gB1E08NY5_0;
	wire w_dff_A_0PM042256_0;
	wire w_dff_A_LQ7uBeoz3_0;
	wire w_dff_A_dkVtVOUx5_0;
	wire w_dff_A_HJzGzpIc0_0;
	wire w_dff_A_S4dd3pon7_0;
	wire w_dff_A_6vceczxd9_0;
	wire w_dff_A_uUkxmizt2_0;
	wire w_dff_A_JD0ybVW66_0;
	wire w_dff_A_zo8Acg4y6_0;
	wire w_dff_A_V0Jxk4lg2_2;
	wire w_dff_A_3fAq5jVR5_0;
	wire w_dff_A_JreTsS6M8_0;
	wire w_dff_A_F36WOgGT9_0;
	wire w_dff_A_6RaYDjH62_0;
	wire w_dff_A_0JSxN4jW6_0;
	wire w_dff_A_NGaX2Gbd8_0;
	wire w_dff_A_icfMg0JI1_0;
	wire w_dff_A_8rfjwdNr7_0;
	wire w_dff_A_cwR4FYFA7_0;
	wire w_dff_A_VD44ma169_0;
	wire w_dff_A_tcCrlzQ04_0;
	wire w_dff_A_rvBYlond9_0;
	wire w_dff_A_kqInnoN63_0;
	wire w_dff_A_2jvwvDog9_0;
	wire w_dff_A_xqc4ukvK3_1;
	wire w_dff_A_lN3QgUuj6_0;
	wire w_dff_A_qlI3RfQY3_0;
	wire w_dff_A_OVUrvpWZ7_0;
	wire w_dff_A_DPxXXKgb9_0;
	wire w_dff_A_PRENhfcU9_0;
	wire w_dff_A_c6EHn7EM2_0;
	wire w_dff_A_9YirO3EP8_0;
	wire w_dff_A_e3LLgrUR6_0;
	wire w_dff_A_YdeDvYTh5_0;
	wire w_dff_A_R11IaAAo2_1;
	wire w_dff_A_34wxYVgv2_0;
	wire w_dff_A_aMsFzV8k2_0;
	wire w_dff_A_f2iSOEjN8_0;
	wire w_dff_A_4jZyDO4a2_0;
	wire w_dff_A_6KvbrMhZ3_0;
	wire w_dff_A_yn9p9jYD3_0;
	wire w_dff_A_BI9Q3Wlq4_0;
	wire w_dff_A_iFNhOtGr8_0;
	wire w_dff_A_PumRsgop7_0;
	wire w_dff_A_pPGSV0VE7_0;
	wire w_dff_A_VrTxVwbE1_0;
	wire w_dff_A_UWtWUJzu5_1;
	wire w_dff_A_39IcbON36_0;
	wire w_dff_A_FYxACZtd5_0;
	wire w_dff_A_ayPqb62j7_0;
	wire w_dff_A_nkWawfgl9_0;
	wire w_dff_A_35pPbuLW8_0;
	wire w_dff_A_PV0eDmLD2_0;
	wire w_dff_A_Q5O5yeK04_0;
	wire w_dff_A_dPif8dpM3_0;
	wire w_dff_A_lSAPL9oN3_0;
	wire w_dff_A_Aptn8CNa9_0;
	wire w_dff_A_JaIYGaxb7_0;
	wire w_dff_A_NhEquGyl5_0;
	wire w_dff_A_cO0UkzHS2_1;
	wire w_dff_A_ip7BzEE51_0;
	wire w_dff_A_BAXNnSZN6_0;
	wire w_dff_A_uvL9Ps9j7_0;
	wire w_dff_A_Niz0Sftl6_0;
	wire w_dff_A_AbRH6wS81_0;
	wire w_dff_A_52SqaebH2_0;
	wire w_dff_A_0z11elp72_0;
	wire w_dff_A_wbxJ4dX05_0;
	wire w_dff_A_PhSOUEfc0_0;
	wire w_dff_A_bEapAac94_0;
	wire w_dff_A_H8DrywDq1_0;
	wire w_dff_A_gGj9Yd925_0;
	wire w_dff_A_OiVSYWaj6_0;
	wire w_dff_A_XkoNU5Q13_1;
	wire w_dff_A_RKrC5ZHB3_0;
	wire w_dff_A_Czml2uA94_0;
	wire w_dff_A_B0VxtW2z7_0;
	wire w_dff_A_5gFIGXCd4_0;
	wire w_dff_A_g1LOYUUf7_0;
	wire w_dff_A_zQTHNMeU9_0;
	wire w_dff_A_irAHEeFG0_0;
	wire w_dff_A_n8FKUin47_0;
	wire w_dff_A_MWSLrTf99_0;
	wire w_dff_A_9qqlxDDT8_0;
	wire w_dff_A_LCOpbfAy6_0;
	wire w_dff_A_izv6SuXY7_0;
	wire w_dff_A_7KmsnVih6_0;
	wire w_dff_A_bvKln7vL9_0;
	wire w_dff_A_RphIj3Cg1_0;
	wire w_dff_A_gsdpr9LF7_0;
	wire w_dff_A_yoQ7gBu71_1;
	wire w_dff_A_iSYEqmS21_0;
	wire w_dff_A_uNS3x3oT3_0;
	wire w_dff_A_Lx3rdpWJ6_0;
	wire w_dff_A_vZ4IEJ8v7_0;
	wire w_dff_A_hEIGV5SA4_0;
	wire w_dff_A_weId0Al02_0;
	wire w_dff_A_D9x0JpWX4_0;
	wire w_dff_A_S0O6gJBc6_0;
	wire w_dff_A_YAUmi3wI3_0;
	wire w_dff_A_HEe99Rb48_0;
	wire w_dff_A_7YMUW1C25_0;
	wire w_dff_A_xZWHCZ1w7_0;
	wire w_dff_A_S2M7FuCm3_0;
	wire w_dff_A_zfigGTY95_0;
	wire w_dff_A_xE6rwWB77_0;
	wire w_dff_A_DyG2AYCJ2_0;
	wire w_dff_A_KYIcgXZK9_0;
	wire w_dff_A_DE0qVNGK7_0;
	wire w_dff_A_BkWFxhEB2_2;
	wire w_dff_A_LIHDGeJw9_0;
	wire w_dff_A_Q2z2mpl82_0;
	wire w_dff_A_FK5KjLBy5_0;
	wire w_dff_A_nus5Dde81_0;
	wire w_dff_A_XLGJ52ZR5_2;
	wire w_dff_A_yO4CAvnu2_0;
	wire w_dff_A_pxA9yVPv5_0;
	wire w_dff_A_dLK0pC1x3_0;
	wire w_dff_A_o0Jw7GZ85_0;
	wire w_dff_A_IGgCN6zc6_0;
	wire w_dff_A_tYqxSV9P9_0;
	wire w_dff_A_Gm6tIDHY6_0;
	wire w_dff_A_e2padhDy3_2;
	wire w_dff_A_uBXnkbt63_0;
	wire w_dff_A_eEPrYxCc7_0;
	wire w_dff_A_FD3nYQMz1_0;
	wire w_dff_A_KoTCeSlk2_0;
	wire w_dff_A_QonrsW5u4_0;
	wire w_dff_A_5T2T07X71_0;
	wire w_dff_A_I7e5AaJw5_0;
	wire w_dff_A_qZnUxT0U4_0;
	wire w_dff_A_FpbqjnAy5_0;
	wire w_dff_A_feb7IkaZ7_0;
	wire w_dff_A_OxP4DydG3_0;
	wire w_dff_A_F5nQuhG97_0;
	wire w_dff_A_cJoOyBTr8_0;
	wire w_dff_A_G2chA7m48_2;
	wire w_dff_A_wVK0n5eK1_0;
	wire w_dff_A_W2JuKv913_0;
	wire w_dff_A_xoMZBcXG3_0;
	wire w_dff_A_JwSLsdri0_0;
	wire w_dff_A_nSVnXpew0_0;
	wire w_dff_A_W6ZacWyL9_0;
	wire w_dff_A_rYbRjz7Y4_0;
	wire w_dff_A_Pf22BUOx2_0;
	wire w_dff_A_aScrGtdP7_0;
	wire w_dff_A_DjvQs8ro6_0;
	wire w_dff_A_YNj8iHuq2_0;
	wire w_dff_A_IeYx8ogJ0_0;
	wire w_dff_A_P0pqoz6w3_0;
	wire w_dff_A_KfeUhVrq5_2;
	wire w_dff_A_sw9TurKs6_0;
	wire w_dff_A_gdKEuIgu0_0;
	wire w_dff_A_6TAhwbi33_0;
	wire w_dff_A_f8wdPuSn7_0;
	wire w_dff_A_PPEJbsS00_0;
	wire w_dff_A_VcBBHN7L5_0;
	wire w_dff_A_PcgqmF0C8_2;
	wire w_dff_A_LlYxkoFK2_0;
	wire w_dff_A_PrxaREaY1_0;
	wire w_dff_A_WrM61pGw6_0;
	wire w_dff_A_6Agh3nae8_0;
	wire w_dff_A_ZDzdhXwH2_0;
	wire w_dff_A_ubzKpfvl7_0;
	wire w_dff_A_IoZq34576_0;
	wire w_dff_A_zt1aQIae0_0;
	wire w_dff_A_m0ajpebn0_2;
	wire w_dff_A_H21ayT7A1_0;
	wire w_dff_A_9qftIk2h8_0;
	wire w_dff_A_CEZNUDmR0_0;
	wire w_dff_A_LF3C5FvE0_0;
	wire w_dff_A_O2C8IRlZ2_0;
	wire w_dff_A_MtlKiWrl1_0;
	wire w_dff_A_Rnp7sFGs3_0;
	wire w_dff_A_hv5YRrBr0_0;
	wire w_dff_A_79skVkXk9_0;
	wire w_dff_A_XI6uvqqZ6_2;
	wire w_dff_A_3m7y0daf0_0;
	wire w_dff_A_cfPFmr3Q8_0;
	wire w_dff_A_AT7wuAsi5_0;
	wire w_dff_A_d0gbtnvA0_0;
	wire w_dff_A_o4BH9woU7_0;
	wire w_dff_A_IyjwKG330_0;
	wire w_dff_A_4rkMP9574_0;
	wire w_dff_A_CGycL2bp0_0;
	wire w_dff_A_Ekrj35rS5_0;
	wire w_dff_A_YdVTRq8h2_0;
	wire w_dff_A_DLFcmILU9_2;
	wire w_dff_A_7DsRj9d82_0;
	wire w_dff_A_IZWbhzad0_0;
	wire w_dff_A_07IHCwMa5_0;
	wire w_dff_A_j941N7RO1_0;
	wire w_dff_A_CQJAyi6Z7_0;
	wire w_dff_A_TuKixy3M7_0;
	wire w_dff_A_YktHXzVq0_2;
	wire w_dff_A_re5PmL8l6_0;
	wire w_dff_A_AmdGjX9a3_0;
	wire w_dff_A_L8VBNfcp8_0;
	wire w_dff_A_R4aHEPUq6_0;
	wire w_dff_A_7uUWhyxP3_0;
	wire w_dff_A_IfoUIBxR7_0;
	wire w_dff_A_CmysDfHQ4_0;
	wire w_dff_A_QLxuj4PK5_0;
	wire w_dff_A_cyMtHO7V5_2;
	wire w_dff_A_sUutweHT1_0;
	wire w_dff_A_fBhiAi4m1_0;
	wire w_dff_A_yovYQJGz1_0;
	wire w_dff_A_nw5VLl9K3_0;
	wire w_dff_A_Nj7wgGHs1_0;
	wire w_dff_A_JdRDKO1R0_0;
	wire w_dff_A_N7F4nlJd9_0;
	wire w_dff_A_gforHNgk5_0;
	wire w_dff_A_TqNE87JS0_0;
	wire w_dff_A_UsxZO5xA4_2;
	wire w_dff_A_G4UTTrst8_0;
	wire w_dff_A_1npkqYoq4_0;
	wire w_dff_A_ycIUmILo3_0;
	wire w_dff_A_RmDXIECh4_0;
	wire w_dff_A_z1RsAgon6_0;
	wire w_dff_A_10lPO5b46_0;
	wire w_dff_A_2WgqWnaS6_0;
	wire w_dff_A_E6rFXZc67_0;
	wire w_dff_A_SCaJMEFS6_0;
	wire w_dff_A_R4zKaMHj4_0;
	wire w_dff_A_6jd38nub0_2;
	wire w_dff_A_HUUyLBEI8_0;
	wire w_dff_A_NJWHBOQZ2_0;
	wire w_dff_A_8bF9mKUP4_0;
	wire w_dff_A_IkevpuYe7_0;
	wire w_dff_A_33ApNxvO6_0;
	wire w_dff_A_OpM8B9au0_2;
	wire w_dff_A_aI0b3nHX3_0;
	wire w_dff_A_eOUS4aCB5_0;
	wire w_dff_A_Movwvcct3_0;
	wire w_dff_A_WU3jNiUi5_0;
	wire w_dff_A_QBGXEpzD3_0;
	wire w_dff_A_g0GIViA89_0;
	wire w_dff_A_amorDON28_0;
	wire w_dff_A_TezhaO5U8_0;
	wire w_dff_A_bMCyt9rB7_0;
	wire w_dff_A_udMizoxK1_2;
	wire w_dff_A_yBkPGO3U5_0;
	wire w_dff_A_wEysfK7J6_0;
	wire w_dff_A_zETBLhsg2_0;
	wire w_dff_A_3V4LSvAs7_0;
	wire w_dff_A_xMKSsKJY5_0;
	wire w_dff_A_vzrUmWJS2_0;
	wire w_dff_A_92m1C4v31_0;
	wire w_dff_A_fy4KqLWz1_0;
	wire w_dff_A_TCP58EKm3_2;
	wire w_dff_A_iqqhNhl31_0;
	wire w_dff_A_9P5V4bFX5_0;
	wire w_dff_A_DRJfTUuy4_0;
	wire w_dff_A_LQhoXsez3_0;
	wire w_dff_A_27r3yQnt9_0;
	wire w_dff_A_jm2Pknel3_0;
	wire w_dff_A_aNCUmeGx3_0;
	wire w_dff_A_QvBFmF6Z6_2;
	wire w_dff_A_0fdGEpoZ3_0;
	wire w_dff_A_O3kUIhD13_0;
	wire w_dff_A_YqtBKm4R3_0;
	wire w_dff_A_nowEBGt29_0;
	wire w_dff_A_paLQIGTv9_0;
	wire w_dff_A_njPQMHMP1_2;
	wire w_dff_A_8caSmFim4_0;
	wire w_dff_A_ZIDX8myp7_0;
	wire w_dff_A_yt2ugcf46_0;
	wire w_dff_A_1hHPdofn0_0;
	wire w_dff_A_ABEYC4pv5_0;
	wire w_dff_A_HfBsieBw1_0;
	wire w_dff_A_MeHZ2idK8_0;
	wire w_dff_A_BucchbI89_0;
	wire w_dff_A_Mrg8eEnt9_0;
	wire w_dff_A_ZS1XpX9r3_2;
	wire w_dff_A_zdlHojwO9_0;
	wire w_dff_A_rXAFWKTq6_0;
	wire w_dff_A_NaHH3ghF9_0;
	wire w_dff_A_HGPSY1TS8_0;
	wire w_dff_A_sZZ8GS4z4_0;
	wire w_dff_A_0TPxsssF6_0;
	wire w_dff_A_yox6R9RO2_0;
	wire w_dff_A_DSeg5Ow66_0;
	wire w_dff_A_zWSShnYZ7_2;
	wire w_dff_A_wKc1AnBc5_0;
	wire w_dff_A_psyDHTXp7_0;
	wire w_dff_A_NBLqhgg33_0;
	wire w_dff_A_go4tHWlx0_0;
	wire w_dff_A_c9CRuBSl9_0;
	wire w_dff_A_Gjjnfko22_0;
	wire w_dff_A_86oNSgpI9_0;
	wire w_dff_A_l4yz9gMX7_2;
	wire w_dff_A_zkYGFyXL7_0;
	wire w_dff_A_VRRIksgD8_0;
	wire w_dff_A_r3tqBjKz0_0;
	wire w_dff_A_OY81yL1H5_0;
	wire w_dff_A_L9zsaGmQ8_2;
	wire w_dff_A_LYpe9dVu2_0;
	wire w_dff_A_fuy1ln707_0;
	wire w_dff_A_qIv0wFGT5_0;
	wire w_dff_A_THk1K6z39_0;
	wire w_dff_A_9YHmGWnu8_0;
	wire w_dff_A_k3ttNZWg1_0;
	wire w_dff_A_USZW6DS72_0;
	wire w_dff_A_JzIb8vCp1_0;
	wire w_dff_A_9EZjqA4L7_1;
	wire w_dff_A_bQrR0xJV0_0;
	wire w_dff_A_pCvGfdx16_0;
	wire w_dff_A_YYRBnywg7_0;
	wire w_dff_A_wj5tLXI33_0;
	wire w_dff_A_dwolBJTY9_1;
	wire w_dff_A_BKpGG5iG4_0;
	wire w_dff_A_Hpep7J3y2_0;
	wire w_dff_A_JRdwbNRh2_0;
	wire w_dff_A_vjXltcIc1_0;
	wire w_dff_A_AlalE32A0_0;
	wire w_dff_A_m8FZdKM60_0;
	wire w_dff_A_p1awfmKN1_0;
	wire w_dff_A_3wJHFv7k4_1;
	wire w_dff_A_VkfNnmTx6_0;
	wire w_dff_A_3XnJbGon3_0;
	wire w_dff_A_VIfu4nsG8_0;
	wire w_dff_A_92RiWWjv9_0;
	wire w_dff_A_IGMm0hw32_0;
	wire w_dff_A_M8CvIGpZ2_0;
	wire w_dff_A_6fxtla8y5_0;
	wire w_dff_A_MBb3kScK9_1;
	wire w_dff_A_UGF4B9OL7_0;
	wire w_dff_A_5cW82O3G2_0;
	wire w_dff_A_2DXE5XMF0_0;
	wire w_dff_A_zGdrRZ2t6_0;
	wire w_dff_A_7kQy0GeY2_0;
	wire w_dff_A_i08W0axm3_0;
	wire w_dff_A_EsSEP6TS5_0;
	wire w_dff_A_fmwDIW7V4_0;
	wire w_dff_A_nqVLCUVr3_2;
	wire w_dff_A_0VfPSdb12_0;
	wire w_dff_A_Iagi2dte9_0;
	wire w_dff_A_FlMEXxlu2_0;
	wire w_dff_A_sBiLunp72_0;
	wire w_dff_A_A0adeJyV5_0;
	wire w_dff_A_Od26WcvR8_0;
	wire w_dff_A_na0vV0mC1_0;
	wire w_dff_A_cfghQrmU8_0;
	wire w_dff_A_lU2XKDt26_0;
	wire w_dff_A_p1ahxHWL0_0;
	wire w_dff_A_xDQ8vvcq9_0;
	wire w_dff_A_38UsTg3g7_0;
	wire w_dff_A_PV3dgX6G1_0;
	wire w_dff_A_QFuOL9ih1_0;
	wire w_dff_A_aoOEAbmr5_0;
	wire w_dff_A_O5MACyFk6_1;
	wire w_dff_A_NZNHPMkf8_0;
	wire w_dff_A_nrSWo5Hn7_0;
	wire w_dff_A_5l5XOZcE6_0;
	wire w_dff_A_qeZz187w9_1;
	wire w_dff_A_SsNyH2IT6_0;
	wire w_dff_A_aRHYR99A4_0;
	wire w_dff_A_5X9sX5nS6_0;
	wire w_dff_A_v0mXYtEf6_0;
	wire w_dff_A_JgOw3Pju8_1;
	wire w_dff_A_sJ5zsEQo0_0;
	wire w_dff_A_FV1ZoX9j0_0;
	wire w_dff_A_u57xHKBL7_0;
	wire w_dff_A_Vsy9ohhV8_0;
	wire w_dff_A_yVWuYFiZ9_0;
	wire w_dff_A_1POWETG96_0;
	wire w_dff_A_4kASBhIa2_1;
	wire w_dff_A_ALiaipha0_0;
	wire w_dff_A_ULjYCfey9_0;
	wire w_dff_A_YwmtFct39_0;
	wire w_dff_A_Ax9852qS7_0;
	wire w_dff_A_Lv5BfZpU2_0;
	wire w_dff_A_PVNJ4laq9_0;
	wire w_dff_A_JnOKkwIw7_0;
	wire w_dff_A_EPXAZVpy7_2;
	wire w_dff_A_U2KV2y4S7_0;
	wire w_dff_A_8rFUIk6B2_0;
	wire w_dff_A_A0bT2Z0q4_2;
	wire w_dff_A_a1LOtgJo5_0;
	wire w_dff_A_AonfvHhS2_0;
	wire w_dff_A_aSx5mPAn3_2;
	wire w_dff_A_98miXHfY4_0;
	wire w_dff_A_N8kAfbe75_0;
	wire w_dff_A_B9YxbKYa1_0;
	wire w_dff_A_EvzIhjy47_2;
	wire w_dff_A_lE73QFUH6_0;
	wire w_dff_A_brAqeK2M2_0;
	wire w_dff_A_gmj7bXCZ4_0;
	wire w_dff_A_5IAg5QGE8_2;
	wire w_dff_A_cczKyqNy3_0;
	wire w_dff_A_6fF4pLax1_0;
	wire w_dff_A_IUweG6cp8_0;
	wire w_dff_A_YPI6aWDE5_0;
	wire w_dff_A_KRUM41us5_2;
	wire w_dff_A_Z4Js1zJe9_0;
	wire w_dff_A_XS2z2DUo2_0;
	wire w_dff_A_uO8HpWfq1_0;
	wire w_dff_A_RrTJUjUs0_2;
	wire w_dff_A_uaTZb3Xr7_0;
	wire w_dff_A_Yb1mhufn6_0;
	wire w_dff_A_FRtqdOhg9_0;
	wire w_dff_A_sdnfD5209_2;
	wire w_dff_A_MxF9yI1R1_0;
	wire w_dff_A_oHh2Qmiy7_0;
	wire w_dff_A_MnACyr4n1_0;
	wire w_dff_A_RgW3IAYd3_0;
	wire w_dff_A_Gwj90k1Q2_2;
	wire w_dff_A_9ysUNOTD0_0;
	wire w_dff_A_QHls6gRw0_0;
	wire w_dff_A_0GymOqF51_0;
	wire w_dff_A_G2E6wyy35_2;
	wire w_dff_A_LNUwRMhl1_0;
	wire w_dff_A_7VnH1jEX5_0;
	wire w_dff_A_sGgb8Vsx5_2;
	wire w_dff_A_Ln59w4Pj7_0;
	wire w_dff_A_OapA63Vb1_0;
	wire w_dff_A_7PhnTXaZ8_2;
	wire w_dff_A_U3jvNd3r3_0;
	wire w_dff_A_RjIELs5s6_2;
	wire w_dff_A_lDl6L8a50_0;
	wire w_dff_A_G4lu5pDk8_0;
	wire w_dff_A_JLHAKdxX1_0;
	wire w_dff_A_nq2iXq3a8_2;
	wire w_dff_A_AaUtWyPQ7_0;
	wire w_dff_A_sqk5T6Ib0_0;
	wire w_dff_A_LZXvWiyX4_2;
	wire w_dff_A_W7owOvbo8_0;
	wire w_dff_A_rCUTpasy5_0;
	wire w_dff_A_wCM0Ubje4_2;
	wire w_dff_A_G8P3GmPF3_0;
	wire w_dff_A_NFX8Ro7t6_2;
	wire w_dff_A_PLc1xrpK6_0;
	wire w_dff_A_C7vfaVHx9_0;
	wire w_dff_A_CTAO9IKv4_0;
	wire w_dff_A_bDIpSuPb9_2;
	wire w_dff_A_lrlwHHYA8_0;
	wire w_dff_A_mKw851y78_0;
	wire w_dff_A_VCgMwWwu9_0;
	wire w_dff_A_5NIX1Iv46_2;
	wire w_dff_A_X47nM5mB6_2;
	jnot g0000(.din(w_G545_0[2]),.dout(w_dff_A_V5AYLoBR3_1),.clk(gclk));
	jnot g0001(.din(w_G348_0[1]),.dout(G599_fa_),.clk(gclk));
	jnot g0002(.din(G366),.dout(G600_fa_),.clk(gclk));
	jand g0003(.dina(w_G562_0[1]),.dinb(w_G552_0[1]),.dout(G601_fa_),.clk(gclk));
	jnot g0004(.din(w_G549_0[2]),.dout(w_dff_A_s2RVKcId6_1),.clk(gclk));
	jnot g0005(.din(G338),.dout(G611_fa_),.clk(gclk));
	jnot g0006(.din(w_G358_0[1]),.dout(G612_fa_),.clk(gclk));
	jand g0007(.dina(G145),.dinb(w_G141_2[2]),.dout(w_dff_A_GlKmi3Mx5_2),.clk(gclk));
	jnot g0008(.din(w_G245_0[1]),.dout(w_dff_A_xyLwOATF7_1),.clk(gclk));
	jnot g0009(.din(w_G552_0[0]),.dout(w_dff_A_H8rH6ICZ3_1),.clk(gclk));
	jnot g0010(.din(w_G562_0[0]),.dout(w_dff_A_Xusarkiy7_1),.clk(gclk));
	jnot g0011(.din(w_G559_0[1]),.dout(w_dff_A_pmLPKsfd4_1),.clk(gclk));
	jand g0012(.dina(G373),.dinb(w_G1_2[1]),.dout(w_dff_A_RYNJc9DE7_2),.clk(gclk));
	jnot g0013(.din(w_G3173_0[1]),.dout(n314),.clk(gclk));
	jand g0014(.dina(n314),.dinb(w_dff_B_jHQBTdJq4_1),.dout(w_dff_A_yXw8OWlh0_2),.clk(gclk));
	jnot g0015(.din(G27),.dout(n316),.clk(gclk));
	jor g0016(.dina(w_dff_B_Anr4sdjm6_0),.dinb(w_n316_0[1]),.dout(w_dff_A_QrS0w1hc9_2),.clk(gclk));
	jand g0017(.dina(G556),.dinb(G386),.dout(n318),.clk(gclk));
	jnot g0018(.din(w_n318_0[1]),.dout(w_dff_A_LSvafEGP1_1),.clk(gclk));
	jnot g0019(.din(G140),.dout(n320),.clk(gclk));
	jnot g0020(.din(G31),.dout(n321),.clk(gclk));
	jor g0021(.dina(n321),.dinb(w_n316_0[0]),.dout(G809_fa_),.clk(gclk));
	jor g0022(.dina(w_G809_3[1]),.dinb(w_dff_B_IMmybuoF8_1),.dout(w_dff_A_dtpCUlzB5_2),.clk(gclk));
	jnot g0023(.din(w_G299_0[2]),.dout(G593_fa_),.clk(gclk));
	jnot g0024(.din(G86),.dout(n325),.clk(gclk));
	jnot g0025(.din(w_G2358_2[2]),.dout(n326),.clk(gclk));
	jand g0026(.dina(w_n326_2[1]),.dinb(n325),.dout(n327),.clk(gclk));
	jnot g0027(.din(G87),.dout(n328),.clk(gclk));
	jand g0028(.dina(w_G2358_2[1]),.dinb(n328),.dout(n329),.clk(gclk));
	jor g0029(.dina(n329),.dinb(w_G809_3[0]),.dout(n330),.clk(gclk));
	jor g0030(.dina(n330),.dinb(w_dff_B_NU61lJJ87_1),.dout(w_dff_A_DH3gqMbd6_2),.clk(gclk));
	jnot g0031(.din(G88),.dout(n332),.clk(gclk));
	jand g0032(.dina(w_n326_2[0]),.dinb(n332),.dout(n333),.clk(gclk));
	jnot g0033(.din(G34),.dout(n334),.clk(gclk));
	jand g0034(.dina(w_G2358_2[0]),.dinb(n334),.dout(n335),.clk(gclk));
	jor g0035(.dina(n335),.dinb(w_G809_2[2]),.dout(n336),.clk(gclk));
	jor g0036(.dina(w_n336_0[1]),.dinb(w_n333_0[1]),.dout(w_dff_A_4mIO0Omj6_2),.clk(gclk));
	jnot g0037(.din(G83),.dout(n338),.clk(gclk));
	jor g0038(.dina(w_G809_2[1]),.dinb(w_dff_B_gm4p0GP46_1),.dout(w_dff_A_A5LKfscm0_2),.clk(gclk));
	jand g0039(.dina(w_n326_1[2]),.dinb(w_dff_B_vHWIvW9o5_1),.dout(n340),.clk(gclk));
	jand g0040(.dina(w_G2358_1[2]),.dinb(G25),.dout(n341),.clk(gclk));
	jor g0041(.dina(w_dff_B_wR4gaxUk6_0),.dinb(w_G809_2[0]),.dout(n342),.clk(gclk));
	jor g0042(.dina(n342),.dinb(w_dff_B_623LmuQ12_1),.dout(n343),.clk(gclk));
	jand g0043(.dina(n343),.dinb(w_G141_2[1]),.dout(w_dff_A_Dmxui67i6_2),.clk(gclk));
	jand g0044(.dina(w_n326_1[1]),.dinb(w_dff_B_vtIH2h1n6_1),.dout(n345),.clk(gclk));
	jand g0045(.dina(w_G2358_1[1]),.dinb(G81),.dout(n346),.clk(gclk));
	jor g0046(.dina(w_dff_B_IxahGZvQ1_0),.dinb(w_G809_1[2]),.dout(n347),.clk(gclk));
	jor g0047(.dina(n347),.dinb(w_dff_B_pHBgUaoW0_1),.dout(n348),.clk(gclk));
	jand g0048(.dina(n348),.dinb(w_G141_2[0]),.dout(w_dff_A_HfINcbMs5_2),.clk(gclk));
	jand g0049(.dina(w_n326_1[0]),.dinb(w_dff_B_gnNJIjpj5_1),.dout(n350),.clk(gclk));
	jand g0050(.dina(w_G2358_1[0]),.dinb(G23),.dout(n351),.clk(gclk));
	jor g0051(.dina(w_dff_B_DHaR4A7J8_0),.dinb(w_G809_1[1]),.dout(n352),.clk(gclk));
	jor g0052(.dina(n352),.dinb(w_dff_B_aqsw1dbN5_1),.dout(n353),.clk(gclk));
	jand g0053(.dina(n353),.dinb(w_G141_1[2]),.dout(w_dff_A_tqTmAX2J9_2),.clk(gclk));
	jand g0054(.dina(w_n326_0[2]),.dinb(w_dff_B_4YYVXK1V0_1),.dout(n355),.clk(gclk));
	jand g0055(.dina(w_G2358_0[2]),.dinb(G80),.dout(n356),.clk(gclk));
	jor g0056(.dina(w_dff_B_PDQFZ4RW9_0),.dinb(w_G809_1[0]),.dout(n357),.clk(gclk));
	jor g0057(.dina(n357),.dinb(w_dff_B_KqiineDQ9_1),.dout(n358),.clk(gclk));
	jand g0058(.dina(n358),.dinb(w_G141_1[1]),.dout(w_dff_A_q4HuDZnG7_2),.clk(gclk));
	jnot g0059(.din(w_G308_1[2]),.dout(n360),.clk(gclk));
	jand g0060(.dina(w_n360_0[1]),.dinb(w_G251_4[2]),.dout(n361),.clk(gclk));
	jnot g0061(.din(w_G479_1[1]),.dout(n362),.clk(gclk));
	jand g0062(.dina(w_G308_1[1]),.dinb(w_G248_5[1]),.dout(n363),.clk(gclk));
	jor g0063(.dina(n363),.dinb(w_n362_0[1]),.dout(n364),.clk(gclk));
	jor g0064(.dina(n364),.dinb(n361),.dout(n365),.clk(gclk));
	jnot g0065(.din(w_G254_1[2]),.dout(n366),.clk(gclk));
	jand g0066(.dina(w_n360_0[0]),.dinb(w_n366_4[2]),.dout(n367),.clk(gclk));
	jnot g0067(.din(w_G242_1[2]),.dout(n368),.clk(gclk));
	jand g0068(.dina(w_G308_1[0]),.dinb(w_n368_5[1]),.dout(n369),.clk(gclk));
	jor g0069(.dina(n369),.dinb(w_G479_1[0]),.dout(n370),.clk(gclk));
	jor g0070(.dina(n370),.dinb(w_dff_B_eBibGzSN8_1),.dout(n371),.clk(gclk));
	jand g0071(.dina(n371),.dinb(w_dff_B_65tFn0Ix8_1),.dout(n372),.clk(gclk));
	jnot g0072(.din(w_G316_1[2]),.dout(n373),.clk(gclk));
	jand g0073(.dina(w_n373_0[1]),.dinb(w_G251_4[1]),.dout(n374),.clk(gclk));
	jnot g0074(.din(w_G490_1[2]),.dout(n375),.clk(gclk));
	jand g0075(.dina(w_G316_1[1]),.dinb(w_G248_5[0]),.dout(n376),.clk(gclk));
	jor g0076(.dina(n376),.dinb(n375),.dout(n377),.clk(gclk));
	jor g0077(.dina(n377),.dinb(n374),.dout(n378),.clk(gclk));
	jand g0078(.dina(w_n373_0[0]),.dinb(w_n366_4[1]),.dout(n379),.clk(gclk));
	jand g0079(.dina(w_G316_1[0]),.dinb(w_n368_5[0]),.dout(n380),.clk(gclk));
	jor g0080(.dina(n380),.dinb(w_G490_1[1]),.dout(n381),.clk(gclk));
	jor g0081(.dina(n381),.dinb(w_dff_B_MzvEPU5s9_1),.dout(n382),.clk(gclk));
	jand g0082(.dina(n382),.dinb(w_dff_B_mR1RJ9Tk9_1),.dout(n383),.clk(gclk));
	jand g0083(.dina(w_n383_0[2]),.dinb(w_n372_0[2]),.dout(n384),.clk(gclk));
	jnot g0084(.din(w_G351_2[2]),.dout(n385),.clk(gclk));
	jnot g0085(.din(G3550),.dout(n386),.clk(gclk));
	jand g0086(.dina(w_n386_4[2]),.dinb(w_n385_1[2]),.dout(n387),.clk(gclk));
	jnot g0087(.din(w_G534_1[2]),.dout(n388),.clk(gclk));
	jnot g0088(.din(w_G3552_0[1]),.dout(n389),.clk(gclk));
	jand g0089(.dina(w_n389_4[2]),.dinb(w_G351_2[1]),.dout(n390),.clk(gclk));
	jor g0090(.dina(n390),.dinb(w_n388_1[2]),.dout(n391),.clk(gclk));
	jor g0091(.dina(n391),.dinb(w_dff_B_VYhf0rRg0_1),.dout(n392),.clk(gclk));
	jand g0092(.dina(w_G3548_4[2]),.dinb(w_n385_1[1]),.dout(n393),.clk(gclk));
	jand g0093(.dina(w_G3546_5[1]),.dinb(w_G351_2[0]),.dout(n394),.clk(gclk));
	jor g0094(.dina(n394),.dinb(w_G534_1[1]),.dout(n395),.clk(gclk));
	jor g0095(.dina(n395),.dinb(n393),.dout(n396),.clk(gclk));
	jand g0096(.dina(w_dff_B_xSRV8uDk0_0),.dinb(n392),.dout(n397),.clk(gclk));
	jnot g0097(.din(w_G293_0[2]),.dout(n398),.clk(gclk));
	jand g0098(.dina(w_n398_0[2]),.dinb(w_n366_4[0]),.dout(n399),.clk(gclk));
	jand g0099(.dina(w_G293_0[1]),.dinb(w_n368_4[2]),.dout(n400),.clk(gclk));
	jor g0100(.dina(n400),.dinb(n399),.dout(n401),.clk(gclk));
	jnot g0101(.din(w_G251_4[0]),.dout(n402),.clk(gclk));
	jnot g0102(.din(w_G302_0[2]),.dout(n403),.clk(gclk));
	jand g0103(.dina(w_n403_0[1]),.dinb(w_n402_2[1]),.dout(n404),.clk(gclk));
	jnot g0104(.din(w_G248_4[2]),.dout(n405),.clk(gclk));
	jand g0105(.dina(w_G302_0[1]),.dinb(w_n405_2[1]),.dout(n406),.clk(gclk));
	jor g0106(.dina(n406),.dinb(n404),.dout(n407),.clk(gclk));
	jnot g0107(.din(w_n407_0[1]),.dout(n408),.clk(gclk));
	jand g0108(.dina(w_n408_0[1]),.dinb(w_n401_0[2]),.dout(n409),.clk(gclk));
	jnot g0109(.din(w_G514_1[1]),.dout(n410),.clk(gclk));
	jnot g0110(.din(w_G3546_5[0]),.dout(n411),.clk(gclk));
	jand g0111(.dina(n411),.dinb(w_n410_1[1]),.dout(n412),.clk(gclk));
	jand g0112(.dina(w_G3552_0[0]),.dinb(w_G514_1[0]),.dout(n413),.clk(gclk));
	jor g0113(.dina(w_dff_B_lTcAT0Ce7_0),.dinb(n412),.dout(n414),.clk(gclk));
	jnot g0114(.din(w_n414_0[1]),.dout(n415),.clk(gclk));
	jnot g0115(.din(w_G361_0[2]),.dout(n416),.clk(gclk));
	jand g0116(.dina(w_n416_0[1]),.dinb(w_n402_2[0]),.dout(n417),.clk(gclk));
	jand g0117(.dina(w_G361_0[1]),.dinb(w_n405_2[0]),.dout(n418),.clk(gclk));
	jor g0118(.dina(n418),.dinb(n417),.dout(n419),.clk(gclk));
	jnot g0119(.din(w_n419_0[2]),.dout(n420),.clk(gclk));
	jand g0120(.dina(n420),.dinb(n415),.dout(n421),.clk(gclk));
	jand g0121(.dina(n421),.dinb(n409),.dout(n422),.clk(gclk));
	jand g0122(.dina(n422),.dinb(w_n397_0[1]),.dout(n423),.clk(gclk));
	jnot g0123(.din(w_G324_1[2]),.dout(n424),.clk(gclk));
	jand g0124(.dina(w_n386_4[1]),.dinb(w_n424_2[1]),.dout(n425),.clk(gclk));
	jnot g0125(.din(w_G503_1[2]),.dout(n426),.clk(gclk));
	jand g0126(.dina(w_n389_4[1]),.dinb(w_G324_1[1]),.dout(n427),.clk(gclk));
	jor g0127(.dina(n427),.dinb(w_n426_0[1]),.dout(n428),.clk(gclk));
	jor g0128(.dina(n428),.dinb(w_dff_B_axKllIrL3_1),.dout(n429),.clk(gclk));
	jand g0129(.dina(w_G3548_4[1]),.dinb(w_n424_2[0]),.dout(n430),.clk(gclk));
	jand g0130(.dina(w_G3546_4[2]),.dinb(w_G324_1[0]),.dout(n431),.clk(gclk));
	jor g0131(.dina(n431),.dinb(w_G503_1[1]),.dout(n432),.clk(gclk));
	jor g0132(.dina(n432),.dinb(n430),.dout(n433),.clk(gclk));
	jand g0133(.dina(w_dff_B_9zStGqWt6_0),.dinb(n429),.dout(n434),.clk(gclk));
	jnot g0134(.din(w_G341_2[2]),.dout(n435),.clk(gclk));
	jand g0135(.dina(w_n386_4[0]),.dinb(w_n435_1[2]),.dout(n436),.clk(gclk));
	jnot g0136(.din(w_G523_1[1]),.dout(n437),.clk(gclk));
	jand g0137(.dina(w_n389_4[0]),.dinb(w_G341_2[1]),.dout(n438),.clk(gclk));
	jor g0138(.dina(n438),.dinb(w_n437_1[2]),.dout(n439),.clk(gclk));
	jor g0139(.dina(n439),.dinb(w_dff_B_8S4t6fQz2_1),.dout(n440),.clk(gclk));
	jand g0140(.dina(w_G3548_4[0]),.dinb(w_n435_1[1]),.dout(n441),.clk(gclk));
	jand g0141(.dina(w_G3546_4[1]),.dinb(w_G341_2[0]),.dout(n442),.clk(gclk));
	jor g0142(.dina(n442),.dinb(w_G523_1[0]),.dout(n443),.clk(gclk));
	jor g0143(.dina(n443),.dinb(n441),.dout(n444),.clk(gclk));
	jand g0144(.dina(w_dff_B_Ub8q9oaB2_0),.dinb(n440),.dout(n445),.clk(gclk));
	jand g0145(.dina(w_n445_0[1]),.dinb(w_n434_0[1]),.dout(n446),.clk(gclk));
	jand g0146(.dina(w_dff_B_eAqgYHn04_0),.dinb(n423),.dout(n447),.clk(gclk));
	jand g0147(.dina(n447),.dinb(w_dff_B_f3ch99Z31_1),.dout(w_dff_A_heVA6OvF9_2),.clk(gclk));
	jnot g0148(.din(w_G265_2[1]),.dout(n449),.clk(gclk));
	jand g0149(.dina(w_n386_3[2]),.dinb(w_n449_1[2]),.dout(n450),.clk(gclk));
	jnot g0150(.din(w_G400_1[1]),.dout(n451),.clk(gclk));
	jand g0151(.dina(w_n389_3[2]),.dinb(w_G265_2[0]),.dout(n452),.clk(gclk));
	jor g0152(.dina(n452),.dinb(w_n451_1[1]),.dout(n453),.clk(gclk));
	jor g0153(.dina(n453),.dinb(w_dff_B_YQcTVDeX3_1),.dout(n454),.clk(gclk));
	jand g0154(.dina(w_G3548_3[2]),.dinb(w_n449_1[1]),.dout(n455),.clk(gclk));
	jand g0155(.dina(w_G3546_4[0]),.dinb(w_G265_1[2]),.dout(n456),.clk(gclk));
	jor g0156(.dina(n456),.dinb(w_G400_1[0]),.dout(n457),.clk(gclk));
	jor g0157(.dina(n457),.dinb(n455),.dout(n458),.clk(gclk));
	jand g0158(.dina(w_dff_B_aqqTLBTb6_0),.dinb(n454),.dout(n459),.clk(gclk));
	jnot g0159(.din(w_G234_2[1]),.dout(n460),.clk(gclk));
	jand g0160(.dina(w_n386_3[1]),.dinb(w_n460_1[2]),.dout(n461),.clk(gclk));
	jnot g0161(.din(w_G435_1[2]),.dout(n462),.clk(gclk));
	jand g0162(.dina(w_n389_3[1]),.dinb(w_G234_2[0]),.dout(n463),.clk(gclk));
	jor g0163(.dina(n463),.dinb(w_n462_0[2]),.dout(n464),.clk(gclk));
	jor g0164(.dina(n464),.dinb(w_dff_B_xgN6JT9C7_1),.dout(n465),.clk(gclk));
	jand g0165(.dina(w_G3548_3[1]),.dinb(w_n460_1[1]),.dout(n466),.clk(gclk));
	jand g0166(.dina(w_G3546_3[2]),.dinb(w_G234_1[2]),.dout(n467),.clk(gclk));
	jor g0167(.dina(n467),.dinb(w_G435_1[1]),.dout(n468),.clk(gclk));
	jor g0168(.dina(n468),.dinb(n466),.dout(n469),.clk(gclk));
	jand g0169(.dina(w_dff_B_0p97Hk5s7_0),.dinb(n465),.dout(n470),.clk(gclk));
	jnot g0170(.din(w_G257_2[2]),.dout(n471),.clk(gclk));
	jand g0171(.dina(w_n386_3[0]),.dinb(w_n471_1[1]),.dout(n472),.clk(gclk));
	jnot g0172(.din(w_G389_0[2]),.dout(n473),.clk(gclk));
	jand g0173(.dina(w_n389_3[0]),.dinb(w_G257_2[1]),.dout(n474),.clk(gclk));
	jor g0174(.dina(n474),.dinb(w_n473_1[2]),.dout(n475),.clk(gclk));
	jor g0175(.dina(n475),.dinb(w_dff_B_Owewop3E6_1),.dout(n476),.clk(gclk));
	jand g0176(.dina(w_G3548_3[0]),.dinb(w_n471_1[0]),.dout(n477),.clk(gclk));
	jand g0177(.dina(w_G3546_3[1]),.dinb(w_G257_2[0]),.dout(n478),.clk(gclk));
	jor g0178(.dina(n478),.dinb(w_G389_0[1]),.dout(n479),.clk(gclk));
	jor g0179(.dina(n479),.dinb(n477),.dout(n480),.clk(gclk));
	jand g0180(.dina(w_dff_B_SzZAg0xl2_0),.dinb(n476),.dout(n481),.clk(gclk));
	jand g0181(.dina(w_n481_0[1]),.dinb(w_n470_0[1]),.dout(n482),.clk(gclk));
	jand g0182(.dina(n482),.dinb(w_n459_0[1]),.dout(n483),.clk(gclk));
	jnot g0183(.din(w_G273_2[2]),.dout(n484),.clk(gclk));
	jand g0184(.dina(w_n386_2[2]),.dinb(w_n484_1[1]),.dout(n485),.clk(gclk));
	jnot g0185(.din(w_G411_0[2]),.dout(n486),.clk(gclk));
	jand g0186(.dina(w_n389_2[2]),.dinb(w_G273_2[1]),.dout(n487),.clk(gclk));
	jor g0187(.dina(n487),.dinb(w_n486_1[1]),.dout(n488),.clk(gclk));
	jor g0188(.dina(n488),.dinb(w_dff_B_aqDUyMwi0_1),.dout(n489),.clk(gclk));
	jand g0189(.dina(w_G3548_2[2]),.dinb(w_n484_1[0]),.dout(n490),.clk(gclk));
	jand g0190(.dina(w_G3546_3[0]),.dinb(w_G273_2[0]),.dout(n491),.clk(gclk));
	jor g0191(.dina(n491),.dinb(w_G411_0[1]),.dout(n492),.clk(gclk));
	jor g0192(.dina(n492),.dinb(n490),.dout(n493),.clk(gclk));
	jand g0193(.dina(w_dff_B_jgVxFdhx8_0),.dinb(n489),.dout(n494),.clk(gclk));
	jnot g0194(.din(w_G281_2[1]),.dout(n495),.clk(gclk));
	jand g0195(.dina(w_n386_2[1]),.dinb(w_n495_1[2]),.dout(n496),.clk(gclk));
	jnot g0196(.din(w_G374_0[2]),.dout(n497),.clk(gclk));
	jand g0197(.dina(w_n389_2[1]),.dinb(w_G281_2[0]),.dout(n498),.clk(gclk));
	jor g0198(.dina(n498),.dinb(w_n497_1[1]),.dout(n499),.clk(gclk));
	jor g0199(.dina(n499),.dinb(w_dff_B_jwquK25w5_1),.dout(n500),.clk(gclk));
	jand g0200(.dina(w_G3548_2[1]),.dinb(w_n495_1[1]),.dout(n501),.clk(gclk));
	jand g0201(.dina(w_G3546_2[2]),.dinb(w_G281_1[2]),.dout(n502),.clk(gclk));
	jor g0202(.dina(n502),.dinb(w_G374_0[1]),.dout(n503),.clk(gclk));
	jor g0203(.dina(n503),.dinb(n501),.dout(n504),.clk(gclk));
	jand g0204(.dina(w_dff_B_OCIN2bTo6_0),.dinb(n500),.dout(n505),.clk(gclk));
	jand g0205(.dina(w_n505_0[1]),.dinb(w_n494_0[1]),.dout(n506),.clk(gclk));
	jnot g0206(.din(w_G218_2[2]),.dout(n507),.clk(gclk));
	jand g0207(.dina(w_n386_2[0]),.dinb(w_n507_1[1]),.dout(n508),.clk(gclk));
	jnot g0208(.din(w_G468_1[2]),.dout(n509),.clk(gclk));
	jand g0209(.dina(w_n389_2[0]),.dinb(w_G218_2[1]),.dout(n510),.clk(gclk));
	jor g0210(.dina(n510),.dinb(w_n509_0[1]),.dout(n511),.clk(gclk));
	jor g0211(.dina(n511),.dinb(w_dff_B_8ngaOgZp0_1),.dout(n512),.clk(gclk));
	jand g0212(.dina(w_G3548_2[0]),.dinb(w_n507_1[0]),.dout(n513),.clk(gclk));
	jand g0213(.dina(w_G3546_2[1]),.dinb(w_G218_2[0]),.dout(n514),.clk(gclk));
	jor g0214(.dina(n514),.dinb(w_G468_1[1]),.dout(n515),.clk(gclk));
	jor g0215(.dina(n515),.dinb(n513),.dout(n516),.clk(gclk));
	jand g0216(.dina(w_dff_B_5azsRgP08_0),.dinb(n512),.dout(n517),.clk(gclk));
	jnot g0217(.din(w_G206_0[2]),.dout(n518),.clk(gclk));
	jand g0218(.dina(w_G251_3[2]),.dinb(w_n518_1[1]),.dout(n519),.clk(gclk));
	jnot g0219(.din(w_G446_1[2]),.dout(n520),.clk(gclk));
	jand g0220(.dina(w_G248_4[1]),.dinb(w_G206_0[1]),.dout(n521),.clk(gclk));
	jor g0221(.dina(n521),.dinb(n520),.dout(n522),.clk(gclk));
	jor g0222(.dina(n522),.dinb(n519),.dout(n523),.clk(gclk));
	jand g0223(.dina(w_n366_3[2]),.dinb(w_n518_1[0]),.dout(n524),.clk(gclk));
	jand g0224(.dina(w_n368_4[1]),.dinb(w_G206_0[0]),.dout(n525),.clk(gclk));
	jor g0225(.dina(n525),.dinb(w_G446_1[1]),.dout(n526),.clk(gclk));
	jor g0226(.dina(n526),.dinb(w_dff_B_ERk43COR3_1),.dout(n527),.clk(gclk));
	jand g0227(.dina(n527),.dinb(w_dff_B_DM8NHtC44_1),.dout(n528),.clk(gclk));
	jand g0228(.dina(w_n528_0[2]),.dinb(w_n517_0[1]),.dout(n529),.clk(gclk));
	jnot g0229(.din(w_G226_2[2]),.dout(n530),.clk(gclk));
	jand g0230(.dina(w_n386_1[2]),.dinb(w_n530_1[1]),.dout(n531),.clk(gclk));
	jnot g0231(.din(w_G422_2[1]),.dout(n532),.clk(gclk));
	jand g0232(.dina(w_n389_1[2]),.dinb(w_G226_2[1]),.dout(n533),.clk(gclk));
	jor g0233(.dina(n533),.dinb(w_n532_0[1]),.dout(n534),.clk(gclk));
	jor g0234(.dina(n534),.dinb(w_dff_B_uOxuyozF6_1),.dout(n535),.clk(gclk));
	jand g0235(.dina(w_G3548_1[2]),.dinb(w_n530_1[0]),.dout(n536),.clk(gclk));
	jand g0236(.dina(w_G3546_2[0]),.dinb(w_G226_2[0]),.dout(n537),.clk(gclk));
	jor g0237(.dina(n537),.dinb(w_G422_2[0]),.dout(n538),.clk(gclk));
	jor g0238(.dina(n538),.dinb(n536),.dout(n539),.clk(gclk));
	jand g0239(.dina(w_dff_B_4nckjkxE7_0),.dinb(n535),.dout(n540),.clk(gclk));
	jnot g0240(.din(w_G210_2[2]),.dout(n541),.clk(gclk));
	jand g0241(.dina(w_n386_1[1]),.dinb(w_n541_1[1]),.dout(n542),.clk(gclk));
	jnot g0242(.din(w_G457_2[1]),.dout(n543),.clk(gclk));
	jand g0243(.dina(w_n389_1[1]),.dinb(w_G210_2[1]),.dout(n544),.clk(gclk));
	jor g0244(.dina(n544),.dinb(w_n543_0[1]),.dout(n545),.clk(gclk));
	jor g0245(.dina(n545),.dinb(w_dff_B_3iQ4hjCX7_1),.dout(n546),.clk(gclk));
	jand g0246(.dina(w_G3548_1[1]),.dinb(w_n541_1[0]),.dout(n547),.clk(gclk));
	jand g0247(.dina(w_G3546_1[2]),.dinb(w_G210_2[0]),.dout(n548),.clk(gclk));
	jor g0248(.dina(n548),.dinb(w_G457_2[0]),.dout(n549),.clk(gclk));
	jor g0249(.dina(n549),.dinb(n547),.dout(n550),.clk(gclk));
	jand g0250(.dina(w_dff_B_Lm8hocjk6_0),.dinb(n546),.dout(n551),.clk(gclk));
	jand g0251(.dina(w_n551_0[1]),.dinb(w_n540_0[1]),.dout(n552),.clk(gclk));
	jand g0252(.dina(n552),.dinb(n529),.dout(n553),.clk(gclk));
	jand g0253(.dina(n553),.dinb(w_dff_B_uVRcF1Sl0_1),.dout(n554),.clk(gclk));
	jand g0254(.dina(n554),.dinb(w_dff_B_5mlsIGkR7_1),.dout(w_dff_A_98gOsWEt3_2),.clk(gclk));
	jnot g0255(.din(w_G335_4[1]),.dout(n556),.clk(gclk));
	jor g0256(.dina(w_n556_5[1]),.dinb(w_dff_B_KBAynGeM1_1),.dout(n557),.clk(gclk));
	jand g0257(.dina(w_n556_5[0]),.dinb(w_n460_1[0]),.dout(n558),.clk(gclk));
	jnot g0258(.din(n558),.dout(n559),.clk(gclk));
	jand g0259(.dina(n559),.dinb(w_dff_B_KJPtpKsx2_1),.dout(n560),.clk(gclk));
	jxor g0260(.dina(w_n560_1[1]),.dinb(w_G435_1[0]),.dout(n561),.clk(gclk));
	jnot g0261(.din(w_n561_0[2]),.dout(n562),.clk(gclk));
	jnot g0262(.din(G288),.dout(n563),.clk(gclk));
	jand g0263(.dina(w_G335_4[0]),.dinb(n563),.dout(n564),.clk(gclk));
	jand g0264(.dina(w_n556_4[2]),.dinb(w_n495_1[0]),.dout(n565),.clk(gclk));
	jor g0265(.dina(n565),.dinb(n564),.dout(n566),.clk(gclk));
	jxor g0266(.dina(w_n566_0[2]),.dinb(w_n497_1[0]),.dout(n567),.clk(gclk));
	jor g0267(.dina(w_n556_4[1]),.dinb(w_G280_0[1]),.dout(n568),.clk(gclk));
	jor g0268(.dina(w_G335_3[2]),.dinb(w_G273_1[2]),.dout(n569),.clk(gclk));
	jand g0269(.dina(w_n569_0[1]),.dinb(n568),.dout(n570),.clk(gclk));
	jxor g0270(.dina(w_n570_0[1]),.dinb(w_n486_1[0]),.dout(n571),.clk(gclk));
	jnot g0271(.din(w_n571_1[1]),.dout(n572),.clk(gclk));
	jand g0272(.dina(w_n572_0[2]),.dinb(w_n567_1[1]),.dout(n573),.clk(gclk));
	jnot g0273(.din(n573),.dout(n574),.clk(gclk));
	jor g0274(.dina(w_n556_4[0]),.dinb(w_dff_B_LFNFrl5q5_1),.dout(n575),.clk(gclk));
	jor g0275(.dina(w_G335_3[1]),.dinb(w_G257_1[2]),.dout(n576),.clk(gclk));
	jand g0276(.dina(w_dff_B_tbhq58vP9_0),.dinb(n575),.dout(n577),.clk(gclk));
	jxor g0277(.dina(w_n577_0[2]),.dinb(w_n473_1[1]),.dout(n578),.clk(gclk));
	jnot g0278(.din(G272),.dout(n579),.clk(gclk));
	jand g0279(.dina(w_G335_3[0]),.dinb(n579),.dout(n580),.clk(gclk));
	jand g0280(.dina(w_n556_3[2]),.dinb(w_n449_1[0]),.dout(n581),.clk(gclk));
	jor g0281(.dina(n581),.dinb(n580),.dout(n582),.clk(gclk));
	jxor g0282(.dina(w_n582_1[1]),.dinb(w_G400_0[2]),.dout(n583),.clk(gclk));
	jor g0283(.dina(w_n583_1[1]),.dinb(w_n578_0[2]),.dout(n584),.clk(gclk));
	jor g0284(.dina(w_dff_B_CLDgGND10_0),.dinb(w_n574_0[2]),.dout(n585),.clk(gclk));
	jor g0285(.dina(w_n585_0[1]),.dinb(w_n562_0[1]),.dout(n586),.clk(gclk));
	jnot g0286(.din(n586),.dout(n587),.clk(gclk));
	jor g0287(.dina(w_n556_3[1]),.dinb(w_dff_B_hfdQdMaW8_1),.dout(n588),.clk(gclk));
	jor g0288(.dina(w_G335_2[2]),.dinb(w_G210_1[2]),.dout(n589),.clk(gclk));
	jand g0289(.dina(w_dff_B_uFZfeLal0_0),.dinb(n588),.dout(n590),.clk(gclk));
	jxor g0290(.dina(w_n590_1[1]),.dinb(w_G457_1[2]),.dout(n591),.clk(gclk));
	jor g0291(.dina(w_n556_3[0]),.dinb(w_dff_B_VZOWUMFk6_1),.dout(n592),.clk(gclk));
	jand g0292(.dina(w_n556_2[2]),.dinb(w_n518_0[2]),.dout(n593),.clk(gclk));
	jnot g0293(.din(n593),.dout(n594),.clk(gclk));
	jand g0294(.dina(n594),.dinb(w_dff_B_sQt5zr0P4_1),.dout(n595),.clk(gclk));
	jxor g0295(.dina(w_n595_1[1]),.dinb(w_G446_1[0]),.dout(n596),.clk(gclk));
	jand g0296(.dina(w_n596_0[2]),.dinb(w_n591_0[1]),.dout(n597),.clk(gclk));
	jor g0297(.dina(w_n556_2[1]),.dinb(w_dff_B_XgANFRu84_1),.dout(n598),.clk(gclk));
	jor g0298(.dina(w_G335_2[1]),.dinb(w_G226_1[2]),.dout(n599),.clk(gclk));
	jand g0299(.dina(w_dff_B_k5g8YeC02_0),.dinb(n598),.dout(n600),.clk(gclk));
	jxor g0300(.dina(w_n600_1[1]),.dinb(w_G422_1[2]),.dout(n601),.clk(gclk));
	jor g0301(.dina(w_n556_2[0]),.dinb(w_dff_B_Od3WhJOn7_1),.dout(n602),.clk(gclk));
	jor g0302(.dina(w_G335_2[0]),.dinb(w_G218_1[2]),.dout(n603),.clk(gclk));
	jand g0303(.dina(w_dff_B_rlpoLhJZ6_0),.dinb(n602),.dout(n604),.clk(gclk));
	jxor g0304(.dina(w_n604_0[2]),.dinb(w_G468_1[0]),.dout(n605),.clk(gclk));
	jand g0305(.dina(w_n605_2[2]),.dinb(w_n601_0[1]),.dout(n606),.clk(gclk));
	jand g0306(.dina(w_dff_B_hGOH1ICO8_0),.dinb(n597),.dout(n607),.clk(gclk));
	jand g0307(.dina(w_n607_0[2]),.dinb(w_n587_1[1]),.dout(w_dff_A_a8FPstR07_2),.clk(gclk));
	jnot g0308(.din(w_G332_4[2]),.dout(n609),.clk(gclk));
	jor g0309(.dina(w_n609_5[2]),.dinb(w_G331_0[1]),.dout(n610),.clk(gclk));
	jand g0310(.dina(w_n609_5[1]),.dinb(w_n424_1[2]),.dout(n611),.clk(gclk));
	jnot g0311(.din(n611),.dout(n612),.clk(gclk));
	jand g0312(.dina(n612),.dinb(w_dff_B_Tse1RMZe5_1),.dout(n613),.clk(gclk));
	jxor g0313(.dina(w_n613_0[2]),.dinb(w_G503_1[0]),.dout(n614),.clk(gclk));
	jor g0314(.dina(w_G358_0[0]),.dinb(w_n609_5[0]),.dout(n615),.clk(gclk));
	jor g0315(.dina(w_G351_1[2]),.dinb(w_G332_4[1]),.dout(n616),.clk(gclk));
	jand g0316(.dina(w_dff_B_rRKEK39E6_0),.dinb(n615),.dout(n617),.clk(gclk));
	jxor g0317(.dina(w_n617_1[1]),.dinb(w_n388_1[1]),.dout(n618),.clk(gclk));
	jand g0318(.dina(w_G600_0),.dinb(w_G332_4[0]),.dout(n619),.clk(gclk));
	jand g0319(.dina(w_n416_0[0]),.dinb(w_n609_4[2]),.dout(n620),.clk(gclk));
	jor g0320(.dina(n620),.dinb(n619),.dout(n621),.clk(gclk));
	jnot g0321(.din(w_n621_2[1]),.dout(n622),.clk(gclk));
	jor g0322(.dina(w_n622_1[1]),.dinb(w_n618_1[1]),.dout(n623),.clk(gclk));
	jand g0323(.dina(w_G611_0),.dinb(w_G332_3[2]),.dout(n624),.clk(gclk));
	jxor g0324(.dina(w_n624_1[2]),.dinb(w_G514_0[2]),.dout(n625),.clk(gclk));
	jor g0325(.dina(w_G348_0[0]),.dinb(w_n609_4[1]),.dout(n626),.clk(gclk));
	jor g0326(.dina(w_G341_1[2]),.dinb(w_G332_3[1]),.dout(n627),.clk(gclk));
	jand g0327(.dina(w_dff_B_sy6KjLuo3_0),.dinb(n626),.dout(n628),.clk(gclk));
	jxor g0328(.dina(w_n628_0[2]),.dinb(w_n437_1[1]),.dout(n629),.clk(gclk));
	jor g0329(.dina(w_n629_0[2]),.dinb(w_n625_0[2]),.dout(n630),.clk(gclk));
	jor g0330(.dina(n630),.dinb(w_n623_0[1]),.dout(n631),.clk(gclk));
	jnot g0331(.din(w_n631_0[1]),.dout(n632),.clk(gclk));
	jand g0332(.dina(n632),.dinb(w_n614_2[1]),.dout(n633),.clk(gclk));
	jand g0333(.dina(w_G332_3[0]),.dinb(w_G593_0),.dout(n634),.clk(gclk));
	jand g0334(.dina(w_n609_4[0]),.dinb(w_n398_0[1]),.dout(n635),.clk(gclk));
	jor g0335(.dina(n635),.dinb(n634),.dout(n636),.clk(gclk));
	jor g0336(.dina(w_n609_3[2]),.dinb(w_dff_B_Cqd1kKUi5_1),.dout(n637),.clk(gclk));
	jand g0337(.dina(w_n609_3[1]),.dinb(w_n403_0[0]),.dout(n638),.clk(gclk));
	jnot g0338(.din(n638),.dout(n639),.clk(gclk));
	jand g0339(.dina(n639),.dinb(w_dff_B_wQ37Nmac5_1),.dout(n640),.clk(gclk));
	jnot g0340(.din(w_n640_1[2]),.dout(n641),.clk(gclk));
	jand g0341(.dina(w_n641_0[1]),.dinb(w_n636_1[1]),.dout(n642),.clk(gclk));
	jor g0342(.dina(w_n609_3[0]),.dinb(w_dff_B_5Qogf0L47_1),.dout(n643),.clk(gclk));
	jor g0343(.dina(w_G332_2[2]),.dinb(w_G308_0[2]),.dout(n644),.clk(gclk));
	jand g0344(.dina(w_dff_B_UOnL0LPK6_0),.dinb(n643),.dout(n645),.clk(gclk));
	jxor g0345(.dina(w_n645_0[2]),.dinb(w_G479_0[2]),.dout(n646),.clk(gclk));
	jor g0346(.dina(w_n609_2[2]),.dinb(w_dff_B_OVby5Z5C3_1),.dout(n647),.clk(gclk));
	jor g0347(.dina(w_G332_2[1]),.dinb(w_G316_0[2]),.dout(n648),.clk(gclk));
	jand g0348(.dina(w_dff_B_ajomxJhW9_0),.dinb(n647),.dout(n649),.clk(gclk));
	jxor g0349(.dina(w_n649_1[1]),.dinb(w_G490_1[0]),.dout(n650),.clk(gclk));
	jand g0350(.dina(w_n650_0[1]),.dinb(w_n646_0[2]),.dout(n651),.clk(gclk));
	jand g0351(.dina(w_n651_1[1]),.dinb(w_n642_0[1]),.dout(n652),.clk(gclk));
	jand g0352(.dina(w_n652_0[1]),.dinb(w_n633_1[1]),.dout(w_dff_A_iLCWaaL96_2),.clk(gclk));
	jxor g0353(.dina(w_G316_0[1]),.dinb(w_G308_0[1]),.dout(n654),.clk(gclk));
	jxor g0354(.dina(w_G351_1[1]),.dinb(w_G341_1[1]),.dout(n655),.clk(gclk));
	jxor g0355(.dina(n655),.dinb(n654),.dout(n656),.clk(gclk));
	jxor g0356(.dina(w_G369_0[1]),.dinb(w_G361_0[0]),.dout(n657),.clk(gclk));
	jxor g0357(.dina(n657),.dinb(w_n424_1[1]),.dout(n658),.clk(gclk));
	jxor g0358(.dina(w_G302_0[0]),.dinb(w_n398_0[0]),.dout(n659),.clk(gclk));
	jxor g0359(.dina(n659),.dinb(n658),.dout(n660),.clk(gclk));
	jxor g0360(.dina(n660),.dinb(w_dff_B_9v0UvJns1_1),.dout(n661),.clk(gclk));
	jnot g0361(.din(w_n661_0[1]),.dout(w_dff_A_1v2VW66l6_1),.clk(gclk));
	jxor g0362(.dina(w_G226_1[1]),.dinb(w_G218_1[1]),.dout(n663),.clk(gclk));
	jxor g0363(.dina(w_G273_1[1]),.dinb(w_G265_1[1]),.dout(n664),.clk(gclk));
	jxor g0364(.dina(n664),.dinb(n663),.dout(n665),.clk(gclk));
	jxor g0365(.dina(w_G289_0[1]),.dinb(w_G281_1[1]),.dout(n666),.clk(gclk));
	jxor g0366(.dina(w_G257_1[1]),.dinb(w_G234_1[1]),.dout(n667),.clk(gclk));
	jxor g0367(.dina(n667),.dinb(n666),.dout(n668),.clk(gclk));
	jxor g0368(.dina(w_G210_1[1]),.dinb(w_n518_0[1]),.dout(n669),.clk(gclk));
	jxor g0369(.dina(n669),.dinb(n668),.dout(n670),.clk(gclk));
	jxor g0370(.dina(n670),.dinb(w_dff_B_zK5lCcxZ2_1),.dout(n671),.clk(gclk));
	jnot g0371(.din(w_n671_0[1]),.dout(w_dff_A_nMfNfIJ88_1),.clk(gclk));
	jnot g0372(.din(w_n560_1[0]),.dout(n673),.clk(gclk));
	jand g0373(.dina(n673),.dinb(w_n462_0[1]),.dout(n674),.clk(gclk));
	jnot g0374(.din(n674),.dout(n675),.clk(gclk));
	jand g0375(.dina(w_n560_0[2]),.dinb(w_G435_0[2]),.dout(n676),.clk(gclk));
	jnot g0376(.din(w_n577_0[1]),.dout(n677),.clk(gclk));
	jand g0377(.dina(w_n677_0[1]),.dinb(w_n473_1[0]),.dout(n678),.clk(gclk));
	jor g0378(.dina(w_n677_0[0]),.dinb(w_n473_0[2]),.dout(n679),.clk(gclk));
	jand g0379(.dina(w_n582_1[0]),.dinb(w_n451_1[0]),.dout(n680),.clk(gclk));
	jor g0380(.dina(w_n566_0[1]),.dinb(w_n497_0[2]),.dout(n681),.clk(gclk));
	jor g0381(.dina(w_n571_1[0]),.dinb(w_n681_2[1]),.dout(n682),.clk(gclk));
	jnot g0382(.din(w_G280_0[0]),.dout(n683),.clk(gclk));
	jand g0383(.dina(w_G335_1[2]),.dinb(n683),.dout(n684),.clk(gclk));
	jnot g0384(.din(w_n569_0[0]),.dout(n685),.clk(gclk));
	jor g0385(.dina(n685),.dinb(n684),.dout(n686),.clk(gclk));
	jor g0386(.dina(n686),.dinb(w_n486_0[2]),.dout(n687),.clk(gclk));
	jor g0387(.dina(w_n582_0[2]),.dinb(w_n451_0[2]),.dout(n688),.clk(gclk));
	jand g0388(.dina(n688),.dinb(w_n687_0[2]),.dout(n689),.clk(gclk));
	jand g0389(.dina(w_n689_0[1]),.dinb(w_n682_0[1]),.dout(n690),.clk(gclk));
	jor g0390(.dina(n690),.dinb(w_n680_0[1]),.dout(n691),.clk(gclk));
	jand g0391(.dina(w_n691_0[2]),.dinb(w_n679_0[1]),.dout(n692),.clk(gclk));
	jor g0392(.dina(n692),.dinb(w_n678_0[1]),.dout(n693),.clk(gclk));
	jnot g0393(.din(w_n693_0[2]),.dout(n694),.clk(gclk));
	jor g0394(.dina(n694),.dinb(w_dff_B_Db1QQsdW2_1),.dout(n695),.clk(gclk));
	jand g0395(.dina(n695),.dinb(w_dff_B_DeBgD0QU3_1),.dout(n696),.clk(gclk));
	jand g0396(.dina(w_n696_0[2]),.dinb(w_n607_0[1]),.dout(n697),.clk(gclk));
	jand g0397(.dina(w_n595_1[0]),.dinb(w_G446_0[2]),.dout(n698),.clk(gclk));
	jor g0398(.dina(w_n595_0[2]),.dinb(w_G446_0[1]),.dout(n699),.clk(gclk));
	jor g0399(.dina(w_n590_1[0]),.dinb(w_G457_1[1]),.dout(n700),.clk(gclk));
	jand g0400(.dina(w_n590_0[2]),.dinb(w_G457_1[0]),.dout(n701),.clk(gclk));
	jand g0401(.dina(w_n604_0[1]),.dinb(w_G468_0[2]),.dout(n702),.clk(gclk));
	jand g0402(.dina(w_n600_1[0]),.dinb(w_G422_1[1]),.dout(n703),.clk(gclk));
	jand g0403(.dina(w_n605_2[1]),.dinb(w_n703_0[2]),.dout(n704),.clk(gclk));
	jor g0404(.dina(n704),.dinb(w_n702_0[1]),.dout(n705),.clk(gclk));
	jor g0405(.dina(w_n705_0[1]),.dinb(w_dff_B_fJkWUVKm7_1),.dout(n706),.clk(gclk));
	jand g0406(.dina(w_n706_0[1]),.dinb(w_n700_0[1]),.dout(n707),.clk(gclk));
	jand g0407(.dina(w_n707_0[2]),.dinb(w_dff_B_NZ2J9zDL7_1),.dout(n708),.clk(gclk));
	jor g0408(.dina(n708),.dinb(w_dff_B_pRP80RRX9_1),.dout(n709),.clk(gclk));
	jor g0409(.dina(w_n709_0[1]),.dinb(w_n697_0[1]),.dout(w_dff_A_oGRN7NsA0_2),.clk(gclk));
	jand g0410(.dina(w_n613_0[1]),.dinb(w_G503_0[2]),.dout(n711),.clk(gclk));
	jor g0411(.dina(w_n624_1[1]),.dinb(w_n410_1[0]),.dout(n712),.clk(gclk));
	jand g0412(.dina(w_n624_1[0]),.dinb(w_n410_0[2]),.dout(n713),.clk(gclk));
	jand g0413(.dina(w_G599_0),.dinb(w_G332_2[0]),.dout(n714),.clk(gclk));
	jand g0414(.dina(w_n435_1[0]),.dinb(w_n609_2[1]),.dout(n715),.clk(gclk));
	jor g0415(.dina(n715),.dinb(n714),.dout(n716),.clk(gclk));
	jand g0416(.dina(w_n716_0[1]),.dinb(w_n437_1[0]),.dout(n717),.clk(gclk));
	jand g0417(.dina(w_G612_0),.dinb(w_G332_1[2]),.dout(n718),.clk(gclk));
	jand g0418(.dina(w_n385_1[0]),.dinb(w_n609_2[0]),.dout(n719),.clk(gclk));
	jor g0419(.dina(n719),.dinb(n718),.dout(n720),.clk(gclk));
	jand g0420(.dina(w_n720_0[1]),.dinb(w_n388_1[0]),.dout(n721),.clk(gclk));
	jor g0421(.dina(w_n621_2[0]),.dinb(w_n721_0[2]),.dout(n722),.clk(gclk));
	jor g0422(.dina(w_n720_0[0]),.dinb(w_n388_0[2]),.dout(n723),.clk(gclk));
	jor g0423(.dina(w_n716_0[0]),.dinb(w_n437_0[2]),.dout(n724),.clk(gclk));
	jand g0424(.dina(n724),.dinb(w_n723_0[1]),.dout(n725),.clk(gclk));
	jand g0425(.dina(n725),.dinb(n722),.dout(n726),.clk(gclk));
	jor g0426(.dina(w_n726_0[1]),.dinb(w_n717_0[2]),.dout(n727),.clk(gclk));
	jor g0427(.dina(w_n727_0[2]),.dinb(w_dff_B_zFRFbdqH0_1),.dout(n728),.clk(gclk));
	jand g0428(.dina(n728),.dinb(w_dff_B_s7NA25D62_1),.dout(n729),.clk(gclk));
	jnot g0429(.din(w_n729_1[1]),.dout(n730),.clk(gclk));
	jand g0430(.dina(n730),.dinb(w_n614_2[0]),.dout(n731),.clk(gclk));
	jor g0431(.dina(n731),.dinb(w_dff_B_37SCrA0S9_1),.dout(n732),.clk(gclk));
	jand g0432(.dina(w_n732_0[2]),.dinb(w_n651_1[0]),.dout(n733),.clk(gclk));
	jnot g0433(.din(w_n642_0[0]),.dout(n734),.clk(gclk));
	jnot g0434(.din(w_n645_0[1]),.dout(n735),.clk(gclk));
	jand g0435(.dina(w_n735_0[1]),.dinb(w_n362_0[0]),.dout(n736),.clk(gclk));
	jnot g0436(.din(w_n736_0[1]),.dout(n737),.clk(gclk));
	jand g0437(.dina(w_n645_0[0]),.dinb(w_G479_0[1]),.dout(n738),.clk(gclk));
	jand g0438(.dina(w_n649_1[0]),.dinb(w_G490_0[2]),.dout(n739),.clk(gclk));
	jor g0439(.dina(w_n739_1[1]),.dinb(n738),.dout(n740),.clk(gclk));
	jand g0440(.dina(w_n740_0[1]),.dinb(n737),.dout(n741),.clk(gclk));
	jor g0441(.dina(w_n741_0[1]),.dinb(n734),.dout(n742),.clk(gclk));
	jor g0442(.dina(w_n742_0[1]),.dinb(w_n733_0[1]),.dout(w_dff_A_M3kaUjHO8_2),.clk(gclk));
	jnot g0443(.din(w_G54_0[1]),.dout(n744),.clk(gclk));
	jxor g0444(.dina(w_n621_1[2]),.dinb(w_n744_1[2]),.dout(n745),.clk(gclk));
	jnot g0445(.din(w_G4092_1[2]),.dout(n746),.clk(gclk));
	jand g0446(.dina(w_n746_1[2]),.dinb(w_G4091_2[2]),.dout(n747),.clk(gclk));
	jnot g0447(.din(w_n747_3[2]),.dout(n748),.clk(gclk));
	jor g0448(.dina(w_n748_4[1]),.dinb(n745),.dout(n749),.clk(gclk));
	jnot g0449(.din(w_G4091_2[1]),.dout(n750),.clk(gclk));
	jand g0450(.dina(w_n746_1[1]),.dinb(w_n750_1[1]),.dout(n751),.clk(gclk));
	jand g0451(.dina(w_n751_2[1]),.dinb(w_n419_0[1]),.dout(n752),.clk(gclk));
	jand g0452(.dina(w_G4092_1[1]),.dinb(w_n750_1[0]),.dout(n753),.clk(gclk));
	jand g0453(.dina(w_n753_8[1]),.dinb(w_dff_B_BOB3AgmJ6_1),.dout(n754),.clk(gclk));
	jor g0454(.dina(w_dff_B_PFf9ptfD2_0),.dinb(n752),.dout(n755),.clk(gclk));
	jnot g0455(.din(n755),.dout(n756),.clk(gclk));
	jand g0456(.dina(n756),.dinb(w_dff_B_oJLhhSj89_1),.dout(G822_fa_),.clk(gclk));
	jnot g0457(.din(w_n618_1[0]),.dout(n758),.clk(gclk));
	jand g0458(.dina(w_n621_1[1]),.dinb(w_n744_1[1]),.dout(n759),.clk(gclk));
	jnot g0459(.din(w_n759_0[1]),.dout(n760),.clk(gclk));
	jand g0460(.dina(w_n760_0[1]),.dinb(n758),.dout(n761),.clk(gclk));
	jand g0461(.dina(w_n759_0[0]),.dinb(w_n618_0[2]),.dout(n762),.clk(gclk));
	jor g0462(.dina(n762),.dinb(w_n748_4[0]),.dout(n763),.clk(gclk));
	jor g0463(.dina(n763),.dinb(w_n761_0[1]),.dout(n764),.clk(gclk));
	jnot g0464(.din(w_n751_2[0]),.dout(n765),.clk(gclk));
	jor g0465(.dina(w_n765_5[2]),.dinb(w_n397_0[0]),.dout(n766),.clk(gclk));
	jand g0466(.dina(w_n753_8[0]),.dinb(w_dff_B_4HXG8lg23_1),.dout(n767),.clk(gclk));
	jnot g0467(.din(n767),.dout(n768),.clk(gclk));
	jand g0468(.dina(w_dff_B_I3ZfaRf29_0),.dinb(n766),.dout(n769),.clk(gclk));
	jand g0469(.dina(n769),.dinb(n764),.dout(G838_fa_),.clk(gclk));
	jxor g0470(.dina(w_n567_1[0]),.dinb(w_G4_1[1]),.dout(n771),.clk(gclk));
	jand g0471(.dina(w_n771_0[1]),.dinb(w_n747_3[1]),.dout(n772),.clk(gclk));
	jnot g0472(.din(n772),.dout(n773),.clk(gclk));
	jor g0473(.dina(w_n765_5[1]),.dinb(w_n505_0[0]),.dout(n774),.clk(gclk));
	jand g0474(.dina(w_n753_7[2]),.dinb(w_dff_B_pIbDnPuQ1_1),.dout(n775),.clk(gclk));
	jnot g0475(.din(n775),.dout(n776),.clk(gclk));
	jand g0476(.dina(w_dff_B_QnR3iPsJ1_0),.dinb(n774),.dout(n777),.clk(gclk));
	jand g0477(.dina(n777),.dinb(n773),.dout(G861_fa_),.clk(gclk));
	jnot g0478(.din(w_n636_1[0]),.dout(n779),.clk(gclk));
	jand g0479(.dina(w_n633_1[0]),.dinb(w_G54_0[0]),.dout(n780),.clk(gclk));
	jor g0480(.dina(w_dff_B_3RXYZWmb0_0),.dinb(w_n732_0[1]),.dout(n781),.clk(gclk));
	jand g0481(.dina(w_n781_0[2]),.dinb(w_n651_0[2]),.dout(n782),.clk(gclk));
	jor g0482(.dina(n782),.dinb(w_n741_0[0]),.dout(n783),.clk(gclk));
	jnot g0483(.din(w_n783_1[1]),.dout(n784),.clk(gclk));
	jor g0484(.dina(n784),.dinb(w_n779_0[1]),.dout(n785),.clk(gclk));
	jxor g0485(.dina(w_n640_1[1]),.dinb(w_n779_0[0]),.dout(n786),.clk(gclk));
	jnot g0486(.din(w_n786_0[1]),.dout(n787),.clk(gclk));
	jor g0487(.dina(w_n787_0[1]),.dinb(w_n783_1[0]),.dout(n788),.clk(gclk));
	jand g0488(.dina(w_dff_B_gcIRcr813_0),.dinb(n785),.dout(n789),.clk(gclk));
	jnot g0489(.din(w_n789_0[2]),.dout(w_dff_A_i69PVv1d1_1),.clk(gclk));
	jnot g0490(.din(w_G861_0),.dout(n791),.clk(gclk));
	jnot g0491(.din(w_G4087_0[2]),.dout(n792),.clk(gclk));
	jand g0492(.dina(w_G4088_0[2]),.dinb(w_n792_0[1]),.dout(n793),.clk(gclk));
	jand g0493(.dina(w_n793_4[1]),.dinb(w_n791_1[1]),.dout(n794),.clk(gclk));
	jnot g0494(.din(w_G822_0),.dout(n795),.clk(gclk));
	jnot g0495(.din(w_G4088_0[1]),.dout(n796),.clk(gclk));
	jand g0496(.dina(w_n796_0[1]),.dinb(w_n792_0[0]),.dout(n797),.clk(gclk));
	jand g0497(.dina(w_n797_4[1]),.dinb(w_n795_1[1]),.dout(n798),.clk(gclk));
	jand g0498(.dina(w_n796_0[0]),.dinb(w_G4087_0[1]),.dout(n799),.clk(gclk));
	jand g0499(.dina(w_n799_4[1]),.dinb(w_G11_0[1]),.dout(n800),.clk(gclk));
	jand g0500(.dina(w_G4088_0[0]),.dinb(w_G4087_0[0]),.dout(n801),.clk(gclk));
	jand g0501(.dina(w_n801_4[1]),.dinb(w_G61_0[1]),.dout(n802),.clk(gclk));
	jor g0502(.dina(w_dff_B_zMkpzVqJ5_0),.dinb(n800),.dout(n803),.clk(gclk));
	jor g0503(.dina(w_dff_B_jUkZISbW0_0),.dinb(n798),.dout(n804),.clk(gclk));
	jor g0504(.dina(n804),.dinb(n794),.dout(w_dff_A_sV8pytjm1_2),.clk(gclk));
	jand g0505(.dina(w_n729_1[0]),.dinb(w_n631_0[0]),.dout(n806),.clk(gclk));
	jand g0506(.dina(w_n729_0[2]),.dinb(w_n744_1[0]),.dout(n807),.clk(gclk));
	jor g0507(.dina(n807),.dinb(w_n806_0[2]),.dout(n808),.clk(gclk));
	jxor g0508(.dina(n808),.dinb(w_n614_1[2]),.dout(n809),.clk(gclk));
	jor g0509(.dina(w_n809_0[1]),.dinb(w_n748_3[2]),.dout(n810),.clk(gclk));
	jor g0510(.dina(w_n765_5[0]),.dinb(w_n434_0[0]),.dout(n811),.clk(gclk));
	jand g0511(.dina(w_n753_7[1]),.dinb(w_dff_B_SuVya2Y11_1),.dout(n812),.clk(gclk));
	jnot g0512(.din(n812),.dout(n813),.clk(gclk));
	jand g0513(.dina(w_dff_B_IgbdpG980_0),.dinb(n811),.dout(n814),.clk(gclk));
	jand g0514(.dina(w_dff_B_XsD4gAUV9_0),.dinb(n810),.dout(G832_fa_),.clk(gclk));
	jnot g0515(.din(w_n625_0[1]),.dout(n816),.clk(gclk));
	jand g0516(.dina(w_n727_0[1]),.dinb(w_n744_0[2]),.dout(n817),.clk(gclk));
	jand g0517(.dina(w_n726_0[0]),.dinb(w_n623_0[0]),.dout(n818),.clk(gclk));
	jor g0518(.dina(n818),.dinb(w_n717_0[1]),.dout(n819),.clk(gclk));
	jor g0519(.dina(w_n819_0[1]),.dinb(n817),.dout(n820),.clk(gclk));
	jxor g0520(.dina(n820),.dinb(w_dff_B_exRqFS4L6_1),.dout(n821),.clk(gclk));
	jor g0521(.dina(w_n821_0[1]),.dinb(w_n748_3[1]),.dout(n822),.clk(gclk));
	jand g0522(.dina(w_n751_1[2]),.dinb(w_n414_0[0]),.dout(n823),.clk(gclk));
	jand g0523(.dina(w_n753_7[0]),.dinb(w_dff_B_MZ5fi9cp2_1),.dout(n824),.clk(gclk));
	jor g0524(.dina(w_dff_B_SfDirKpW0_0),.dinb(n823),.dout(n825),.clk(gclk));
	jnot g0525(.din(n825),.dout(n826),.clk(gclk));
	jand g0526(.dina(w_dff_B_Ny5gWR5V1_0),.dinb(n822),.dout(G834_fa_),.clk(gclk));
	jor g0527(.dina(w_n617_1[0]),.dinb(w_G534_1[0]),.dout(n828),.clk(gclk));
	jand g0528(.dina(w_n617_0[2]),.dinb(w_G534_0[2]),.dout(n829),.clk(gclk));
	jor g0529(.dina(w_n760_0[0]),.dinb(w_n829_0[1]),.dout(n830),.clk(gclk));
	jand g0530(.dina(n830),.dinb(w_n828_0[2]),.dout(n831),.clk(gclk));
	jxor g0531(.dina(n831),.dinb(w_n629_0[1]),.dout(n832),.clk(gclk));
	jor g0532(.dina(w_n832_0[1]),.dinb(w_n748_3[0]),.dout(n833),.clk(gclk));
	jor g0533(.dina(w_n765_4[2]),.dinb(w_n445_0[0]),.dout(n834),.clk(gclk));
	jand g0534(.dina(w_n753_6[2]),.dinb(w_dff_B_6P5kMzZz0_1),.dout(n835),.clk(gclk));
	jnot g0535(.din(n835),.dout(n836),.clk(gclk));
	jand g0536(.dina(w_dff_B_0cnio3gY3_0),.dinb(n834),.dout(n837),.clk(gclk));
	jand g0537(.dina(w_dff_B_Y9Tox2yI6_0),.dinb(n833),.dout(G836_fa_),.clk(gclk));
	jnot g0538(.din(w_G4090_0[2]),.dout(n839),.clk(gclk));
	jand g0539(.dina(w_n839_0[1]),.dinb(w_G4089_0[2]),.dout(n840),.clk(gclk));
	jand g0540(.dina(w_n840_4[1]),.dinb(w_n791_1[0]),.dout(n841),.clk(gclk));
	jnot g0541(.din(w_G4089_0[1]),.dout(n842),.clk(gclk));
	jand g0542(.dina(w_n839_0[0]),.dinb(w_n842_0[1]),.dout(n843),.clk(gclk));
	jand g0543(.dina(w_n843_4[1]),.dinb(w_n795_1[0]),.dout(n844),.clk(gclk));
	jand g0544(.dina(w_G4090_0[1]),.dinb(w_n842_0[0]),.dout(n845),.clk(gclk));
	jand g0545(.dina(w_n845_4[1]),.dinb(w_G11_0[0]),.dout(n846),.clk(gclk));
	jand g0546(.dina(w_G4090_0[0]),.dinb(w_G4089_0[0]),.dout(n847),.clk(gclk));
	jand g0547(.dina(w_n847_4[1]),.dinb(w_G61_0[0]),.dout(n848),.clk(gclk));
	jor g0548(.dina(w_dff_B_Mt1TyOcg4_0),.dinb(n846),.dout(n849),.clk(gclk));
	jor g0549(.dina(w_dff_B_hYePd4Ob5_0),.dinb(n844),.dout(n850),.clk(gclk));
	jor g0550(.dina(n850),.dinb(n841),.dout(w_dff_A_V0Jxk4lg2_2),.clk(gclk));
	jnot g0551(.din(w_n678_0[0]),.dout(n852),.clk(gclk));
	jnot g0552(.din(w_n679_0[0]),.dout(n853),.clk(gclk));
	jor g0553(.dina(w_n583_1[0]),.dinb(w_n574_0[1]),.dout(n854),.clk(gclk));
	jand g0554(.dina(n854),.dinb(w_n691_0[1]),.dout(n855),.clk(gclk));
	jnot g0555(.din(w_n855_0[1]),.dout(n856),.clk(gclk));
	jnot g0556(.din(w_n691_0[0]),.dout(n857),.clk(gclk));
	jor g0557(.dina(w_n857_0[1]),.dinb(w_G4_1[0]),.dout(n858),.clk(gclk));
	jand g0558(.dina(w_dff_B_5todjbo18_0),.dinb(w_n856_0[1]),.dout(n859),.clk(gclk));
	jor g0559(.dina(w_n859_0[1]),.dinb(w_n853_0[1]),.dout(n860),.clk(gclk));
	jand g0560(.dina(n860),.dinb(w_dff_B_6IfT1C051_1),.dout(n861),.clk(gclk));
	jxor g0561(.dina(n861),.dinb(w_n562_0[0]),.dout(n862),.clk(gclk));
	jor g0562(.dina(w_n862_0[1]),.dinb(w_n748_2[2]),.dout(n863),.clk(gclk));
	jor g0563(.dina(w_n765_4[1]),.dinb(w_n470_0[0]),.dout(n864),.clk(gclk));
	jand g0564(.dina(w_n753_6[1]),.dinb(w_dff_B_5w8VRhtv0_1),.dout(n865),.clk(gclk));
	jnot g0565(.din(n865),.dout(n866),.clk(gclk));
	jand g0566(.dina(w_dff_B_fidH2dRX4_0),.dinb(n864),.dout(n867),.clk(gclk));
	jand g0567(.dina(w_dff_B_tCVmtduJ1_0),.dinb(n863),.dout(G871_fa_),.clk(gclk));
	jxor g0568(.dina(w_n859_0[0]),.dinb(w_n578_0[1]),.dout(n869),.clk(gclk));
	jor g0569(.dina(w_n869_0[1]),.dinb(w_n748_2[1]),.dout(n870),.clk(gclk));
	jor g0570(.dina(w_n765_4[0]),.dinb(w_n481_0[0]),.dout(n871),.clk(gclk));
	jand g0571(.dina(w_n753_6[0]),.dinb(w_dff_B_RdiaBO6R4_1),.dout(n872),.clk(gclk));
	jnot g0572(.din(n872),.dout(n873),.clk(gclk));
	jand g0573(.dina(w_dff_B_xHXuatwA1_0),.dinb(n871),.dout(n874),.clk(gclk));
	jand g0574(.dina(w_dff_B_DggdxiwR2_0),.dinb(n870),.dout(G873_fa_),.clk(gclk));
	jand g0575(.dina(w_n567_0[2]),.dinb(w_G4_0[2]),.dout(n876),.clk(gclk));
	jnot g0576(.din(n876),.dout(n877),.clk(gclk));
	jand g0577(.dina(w_n877_0[1]),.dinb(w_n681_2[0]),.dout(n878),.clk(gclk));
	jor g0578(.dina(n878),.dinb(w_n571_0[2]),.dout(n879),.clk(gclk));
	jand g0579(.dina(w_n879_0[1]),.dinb(w_n687_0[1]),.dout(n880),.clk(gclk));
	jxor g0580(.dina(n880),.dinb(w_n583_0[2]),.dout(n881),.clk(gclk));
	jand g0581(.dina(w_n881_0[1]),.dinb(w_n747_3[0]),.dout(n882),.clk(gclk));
	jnot g0582(.din(n882),.dout(n883),.clk(gclk));
	jor g0583(.dina(w_n765_3[2]),.dinb(w_n459_0[0]),.dout(n884),.clk(gclk));
	jand g0584(.dina(w_n753_5[2]),.dinb(w_dff_B_JkvKrsif8_1),.dout(n885),.clk(gclk));
	jnot g0585(.din(n885),.dout(n886),.clk(gclk));
	jand g0586(.dina(w_dff_B_SUKWI2E52_0),.dinb(n884),.dout(n887),.clk(gclk));
	jand g0587(.dina(w_dff_B_fCDC6jCd4_0),.dinb(n883),.dout(G875_fa_),.clk(gclk));
	jand g0588(.dina(w_n571_0[1]),.dinb(w_n681_1[2]),.dout(n889),.clk(gclk));
	jand g0589(.dina(w_dff_B_L93O4wiF6_0),.dinb(w_n877_0[0]),.dout(n890),.clk(gclk));
	jnot g0590(.din(n890),.dout(n891),.clk(gclk));
	jand g0591(.dina(n891),.dinb(w_n879_0[0]),.dout(n892),.clk(gclk));
	jand g0592(.dina(w_n892_0[1]),.dinb(w_n747_2[2]),.dout(n893),.clk(gclk));
	jnot g0593(.din(n893),.dout(n894),.clk(gclk));
	jor g0594(.dina(w_n765_3[1]),.dinb(w_n494_0[0]),.dout(n895),.clk(gclk));
	jand g0595(.dina(w_n753_5[1]),.dinb(w_dff_B_HudtHNcR4_1),.dout(n896),.clk(gclk));
	jnot g0596(.din(n896),.dout(n897),.clk(gclk));
	jand g0597(.dina(w_dff_B_RCstnGuM4_0),.dinb(n895),.dout(n898),.clk(gclk));
	jand g0598(.dina(w_dff_B_vNdBs2kk8_0),.dinb(n894),.dout(G877_fa_),.clk(gclk));
	jxor g0599(.dina(w_n649_0[2]),.dinb(w_n735_0[0]),.dout(n900),.clk(gclk));
	jxor g0600(.dina(n900),.dinb(w_n786_0[0]),.dout(n901),.clk(gclk));
	jxor g0601(.dina(n901),.dinb(w_n621_1[0]),.dout(n902),.clk(gclk));
	jand g0602(.dina(w_G369_0[0]),.dinb(w_n609_1[2]),.dout(n903),.clk(gclk));
	jand g0603(.dina(G372),.dinb(w_G332_1[1]),.dout(n904),.clk(gclk));
	jor g0604(.dina(w_dff_B_XwVNHKM36_0),.dinb(n903),.dout(n905),.clk(gclk));
	jxor g0605(.dina(n905),.dinb(w_n617_0[1]),.dout(n906),.clk(gclk));
	jxor g0606(.dina(n906),.dinb(w_n628_0[1]),.dout(n907),.clk(gclk));
	jnot g0607(.din(w_G331_0[0]),.dout(n908),.clk(gclk));
	jand g0608(.dina(w_n624_0[2]),.dinb(w_dff_B_ZpFDWVFP4_1),.dout(n909),.clk(gclk));
	jnot g0609(.din(w_n624_0[1]),.dout(n910),.clk(gclk));
	jand g0610(.dina(w_dff_B_u60iEu935_0),.dinb(w_n613_0[0]),.dout(n911),.clk(gclk));
	jor g0611(.dina(n911),.dinb(w_dff_B_fsiWhS0U1_1),.dout(n912),.clk(gclk));
	jxor g0612(.dina(n912),.dinb(w_dff_B_bZ2YK1Iu4_1),.dout(n913),.clk(gclk));
	jxor g0613(.dina(n913),.dinb(n902),.dout(n914),.clk(gclk));
	jnot g0614(.din(w_n914_0[1]),.dout(w_dff_A_XkoNU5Q13_1),.clk(gclk));
	jxor g0615(.dina(w_n577_0[0]),.dinb(w_n566_0[0]),.dout(n916),.clk(gclk));
	jxor g0616(.dina(w_n582_0[1]),.dinb(w_n570_0[0]),.dout(n917),.clk(gclk));
	jxor g0617(.dina(n917),.dinb(n916),.dout(n918),.clk(gclk));
	jxor g0618(.dina(n918),.dinb(w_n590_0[1]),.dout(n919),.clk(gclk));
	jand g0619(.dina(w_n556_1[2]),.dinb(w_G289_0[0]),.dout(n920),.clk(gclk));
	jand g0620(.dina(w_G335_1[1]),.dinb(G292),.dout(n921),.clk(gclk));
	jor g0621(.dina(w_dff_B_WwIkTV058_0),.dinb(n920),.dout(n922),.clk(gclk));
	jxor g0622(.dina(n922),.dinb(w_n600_0[2]),.dout(n923),.clk(gclk));
	jxor g0623(.dina(n923),.dinb(w_n560_0[1]),.dout(n924),.clk(gclk));
	jxor g0624(.dina(w_n604_0[0]),.dinb(w_n595_0[1]),.dout(n925),.clk(gclk));
	jxor g0625(.dina(n925),.dinb(n924),.dout(n926),.clk(gclk));
	jxor g0626(.dina(n926),.dinb(n919),.dout(G1000_fa_),.clk(gclk));
	jnot g0627(.din(w_n596_0[1]),.dout(n928),.clk(gclk));
	jnot g0628(.din(w_n707_0[1]),.dout(n929),.clk(gclk));
	jnot g0629(.din(w_n700_0[0]),.dout(n930),.clk(gclk));
	jnot g0630(.din(w_n605_2[0]),.dout(n931),.clk(gclk));
	jnot g0631(.din(w_n601_0[0]),.dout(n932),.clk(gclk));
	jnot g0632(.din(w_n696_0[1]),.dout(n933),.clk(gclk));
	jand g0633(.dina(w_n587_1[0]),.dinb(w_G4_0[1]),.dout(n934),.clk(gclk));
	jnot g0634(.din(n934),.dout(n935),.clk(gclk));
	jand g0635(.dina(w_dff_B_NtUiBiVq2_0),.dinb(n933),.dout(n936),.clk(gclk));
	jor g0636(.dina(w_n936_0[2]),.dinb(w_n932_0[1]),.dout(n937),.clk(gclk));
	jor g0637(.dina(n937),.dinb(w_dff_B_Apat5Bi87_1),.dout(n938),.clk(gclk));
	jor g0638(.dina(w_n938_0[1]),.dinb(w_n930_0[2]),.dout(n939),.clk(gclk));
	jand g0639(.dina(n939),.dinb(w_dff_B_n8WOJk9M0_1),.dout(n940),.clk(gclk));
	jxor g0640(.dina(n940),.dinb(w_n928_0[1]),.dout(n941),.clk(gclk));
	jnot g0641(.din(w_n941_0[1]),.dout(n942),.clk(gclk));
	jnot g0642(.din(w_n591_0[0]),.dout(n943),.clk(gclk));
	jnot g0643(.din(w_n705_0[0]),.dout(n944),.clk(gclk));
	jand g0644(.dina(w_n938_0[0]),.dinb(w_n944_0[1]),.dout(n945),.clk(gclk));
	jxor g0645(.dina(n945),.dinb(w_n943_0[1]),.dout(n946),.clk(gclk));
	jnot g0646(.din(w_n946_0[1]),.dout(n947),.clk(gclk));
	jor g0647(.dina(w_n600_0[1]),.dinb(w_G422_1[0]),.dout(n948),.clk(gclk));
	jnot g0648(.din(w_n948_0[2]),.dout(n949),.clk(gclk));
	jnot g0649(.din(w_n703_0[1]),.dout(n950),.clk(gclk));
	jand g0650(.dina(w_n936_0[1]),.dinb(w_dff_B_JasYwprn6_1),.dout(n951),.clk(gclk));
	jor g0651(.dina(n951),.dinb(w_dff_B_VGJ83NmS9_1),.dout(n952),.clk(gclk));
	jxor g0652(.dina(n952),.dinb(w_n605_1[2]),.dout(n953),.clk(gclk));
	jxor g0653(.dina(w_n936_0[0]),.dinb(w_n932_0[0]),.dout(n954),.clk(gclk));
	jnot g0654(.din(w_n954_0[1]),.dout(n955),.clk(gclk));
	jnot g0655(.din(w_n881_0[0]),.dout(n956),.clk(gclk));
	jnot g0656(.din(w_n771_0[0]),.dout(n957),.clk(gclk));
	jnot g0657(.din(w_n892_0[0]),.dout(n958),.clk(gclk));
	jand g0658(.dina(n958),.dinb(w_dff_B_qfGQmnHK9_1),.dout(n959),.clk(gclk));
	jand g0659(.dina(n959),.dinb(n956),.dout(n960),.clk(gclk));
	jand g0660(.dina(n960),.dinb(w_n869_0[0]),.dout(n961),.clk(gclk));
	jand g0661(.dina(w_dff_B_TVnOlHoq5_0),.dinb(w_n862_0[0]),.dout(n962),.clk(gclk));
	jand g0662(.dina(w_dff_B_UP050EU05_0),.dinb(n955),.dout(n963),.clk(gclk));
	jand g0663(.dina(n963),.dinb(w_n953_0[1]),.dout(n964),.clk(gclk));
	jand g0664(.dina(w_dff_B_HAwExXEz6_0),.dinb(n947),.dout(n965),.clk(gclk));
	jand g0665(.dina(n965),.dinb(n942),.dout(w_dff_A_BkWFxhEB2_2),.clk(gclk));
	jnot g0666(.din(w_n646_0[1]),.dout(n967),.clk(gclk));
	jor g0667(.dina(w_n649_0[1]),.dinb(w_G490_0[1]),.dout(n968),.clk(gclk));
	jor g0668(.dina(w_n781_0[1]),.dinb(w_n739_1[0]),.dout(n969),.clk(gclk));
	jand g0669(.dina(n969),.dinb(w_n968_0[1]),.dout(n970),.clk(gclk));
	jxor g0670(.dina(n970),.dinb(w_dff_B_DrJsBLWi0_1),.dout(n971),.clk(gclk));
	jxor g0671(.dina(w_n783_0[2]),.dinb(w_n640_1[0]),.dout(n972),.clk(gclk));
	jxor g0672(.dina(w_n781_0[0]),.dinb(w_n650_0[0]),.dout(n973),.clk(gclk));
	jnot g0673(.din(w_n973_0[1]),.dout(n974),.clk(gclk));
	jor g0674(.dina(w_n621_0[2]),.dinb(w_n744_0[1]),.dout(n975),.clk(gclk));
	jand g0675(.dina(n975),.dinb(w_n636_0[2]),.dout(n976),.clk(gclk));
	jand g0676(.dina(w_dff_B_CGVCrTK19_0),.dinb(w_n761_0[0]),.dout(n977),.clk(gclk));
	jand g0677(.dina(w_dff_B_XrSWrNTy2_0),.dinb(w_n832_0[0]),.dout(n978),.clk(gclk));
	jand g0678(.dina(w_dff_B_KMqjl7ai9_0),.dinb(w_n821_0[0]),.dout(n979),.clk(gclk));
	jand g0679(.dina(w_dff_B_HrMMq4VJ6_0),.dinb(w_n809_0[0]),.dout(n980),.clk(gclk));
	jand g0680(.dina(w_dff_B_IJUhH4ns3_0),.dinb(n974),.dout(n981),.clk(gclk));
	jand g0681(.dina(n981),.dinb(w_n972_0[1]),.dout(n982),.clk(gclk));
	jand g0682(.dina(n982),.dinb(w_n971_0[1]),.dout(w_dff_A_XLGJ52ZR5_2),.clk(gclk));
	jnot g0683(.din(w_G1690_0[2]),.dout(n984),.clk(gclk));
	jand g0684(.dina(w_n984_0[1]),.dinb(w_G1689_0[2]),.dout(n985),.clk(gclk));
	jand g0685(.dina(w_n985_4[1]),.dinb(w_n791_0[2]),.dout(n986),.clk(gclk));
	jnot g0686(.din(w_G1689_0[1]),.dout(n987),.clk(gclk));
	jand g0687(.dina(w_n984_0[0]),.dinb(w_n987_0[1]),.dout(n988),.clk(gclk));
	jand g0688(.dina(w_n988_4[1]),.dinb(w_n795_0[2]),.dout(n989),.clk(gclk));
	jand g0689(.dina(w_G1690_0[1]),.dinb(w_n987_0[0]),.dout(n990),.clk(gclk));
	jand g0690(.dina(w_n990_4[1]),.dinb(w_G182_0[1]),.dout(n991),.clk(gclk));
	jand g0691(.dina(w_G1690_0[0]),.dinb(w_G1689_0[0]),.dout(n992),.clk(gclk));
	jand g0692(.dina(w_n992_4[1]),.dinb(w_G185_0[1]),.dout(n993),.clk(gclk));
	jor g0693(.dina(w_dff_B_ryjvrocQ2_0),.dinb(n991),.dout(n994),.clk(gclk));
	jor g0694(.dina(w_dff_B_X5Rb88TQ7_0),.dinb(n989),.dout(n995),.clk(gclk));
	jor g0695(.dina(n995),.dinb(n986),.dout(n996),.clk(gclk));
	jand g0696(.dina(n996),.dinb(w_G137_9[1]),.dout(w_dff_A_e2padhDy3_2),.clk(gclk));
	jnot g0697(.din(w_G1694_0[2]),.dout(n998),.clk(gclk));
	jand g0698(.dina(w_n998_0[1]),.dinb(w_G1691_0[2]),.dout(n999),.clk(gclk));
	jand g0699(.dina(w_n999_4[1]),.dinb(w_n791_0[1]),.dout(n1000),.clk(gclk));
	jnot g0700(.din(w_G1691_0[1]),.dout(n1001),.clk(gclk));
	jand g0701(.dina(w_n998_0[0]),.dinb(w_n1001_0[1]),.dout(n1002),.clk(gclk));
	jand g0702(.dina(w_n1002_4[1]),.dinb(w_n795_0[1]),.dout(n1003),.clk(gclk));
	jand g0703(.dina(w_G1694_0[1]),.dinb(w_n1001_0[0]),.dout(n1004),.clk(gclk));
	jand g0704(.dina(w_n1004_4[1]),.dinb(w_G182_0[0]),.dout(n1005),.clk(gclk));
	jand g0705(.dina(w_G1694_0[0]),.dinb(w_G1691_0[0]),.dout(n1006),.clk(gclk));
	jand g0706(.dina(w_n1006_4[1]),.dinb(w_G185_0[0]),.dout(n1007),.clk(gclk));
	jor g0707(.dina(w_dff_B_EbjnnGtL5_0),.dinb(n1005),.dout(n1008),.clk(gclk));
	jor g0708(.dina(w_dff_B_4EEW3udA8_0),.dinb(n1003),.dout(n1009),.clk(gclk));
	jor g0709(.dina(n1009),.dinb(n1000),.dout(n1010),.clk(gclk));
	jand g0710(.dina(n1010),.dinb(w_G137_9[0]),.dout(w_dff_A_G2chA7m48_2),.clk(gclk));
	jnot g0711(.din(w_G871_0),.dout(n1012),.clk(gclk));
	jand g0712(.dina(w_n1012_1[1]),.dinb(w_n793_4[0]),.dout(n1013),.clk(gclk));
	jnot g0713(.din(w_G832_0),.dout(n1014),.clk(gclk));
	jand g0714(.dina(w_n1014_1[1]),.dinb(w_n797_4[0]),.dout(n1015),.clk(gclk));
	jand g0715(.dina(w_n799_4[0]),.dinb(w_G43_0[1]),.dout(n1016),.clk(gclk));
	jand g0716(.dina(w_n801_4[0]),.dinb(w_G37_0[1]),.dout(n1017),.clk(gclk));
	jor g0717(.dina(w_dff_B_Q0VfgMkX4_0),.dinb(n1016),.dout(n1018),.clk(gclk));
	jor g0718(.dina(w_dff_B_ITRFDaAA8_0),.dinb(n1015),.dout(n1019),.clk(gclk));
	jor g0719(.dina(w_dff_B_ce2DHmUC9_0),.dinb(n1013),.dout(w_dff_A_KfeUhVrq5_2),.clk(gclk));
	jnot g0720(.din(w_G873_0),.dout(n1021),.clk(gclk));
	jand g0721(.dina(w_n1021_1[1]),.dinb(w_n793_3[2]),.dout(n1022),.clk(gclk));
	jnot g0722(.din(w_G834_0),.dout(n1023),.clk(gclk));
	jand g0723(.dina(w_n1023_1[1]),.dinb(w_n797_3[2]),.dout(n1024),.clk(gclk));
	jand g0724(.dina(w_n799_3[2]),.dinb(w_G76_0[1]),.dout(n1025),.clk(gclk));
	jand g0725(.dina(w_n801_3[2]),.dinb(w_G20_0[1]),.dout(n1026),.clk(gclk));
	jor g0726(.dina(w_dff_B_yJdSPpJm7_0),.dinb(n1025),.dout(n1027),.clk(gclk));
	jor g0727(.dina(w_dff_B_SBR2JHGD2_0),.dinb(n1024),.dout(n1028),.clk(gclk));
	jor g0728(.dina(w_dff_B_plgG2qC08_0),.dinb(n1022),.dout(w_dff_A_PcgqmF0C8_2),.clk(gclk));
	jnot g0729(.din(w_G875_0),.dout(n1030),.clk(gclk));
	jand g0730(.dina(w_n1030_1[1]),.dinb(w_n793_3[1]),.dout(n1031),.clk(gclk));
	jnot g0731(.din(w_G836_0),.dout(n1032),.clk(gclk));
	jand g0732(.dina(w_n1032_1[1]),.dinb(w_n797_3[1]),.dout(n1033),.clk(gclk));
	jand g0733(.dina(w_n799_3[1]),.dinb(w_G73_0[1]),.dout(n1034),.clk(gclk));
	jand g0734(.dina(w_n801_3[1]),.dinb(w_G17_0[1]),.dout(n1035),.clk(gclk));
	jor g0735(.dina(w_dff_B_FTDf6ngq6_0),.dinb(n1034),.dout(n1036),.clk(gclk));
	jor g0736(.dina(w_dff_B_b1Bo3pNX3_0),.dinb(n1033),.dout(n1037),.clk(gclk));
	jor g0737(.dina(w_dff_B_LN2JCHDe2_0),.dinb(n1031),.dout(w_dff_A_m0ajpebn0_2),.clk(gclk));
	jnot g0738(.din(w_G877_0),.dout(n1039),.clk(gclk));
	jand g0739(.dina(w_n1039_1[1]),.dinb(w_n793_3[0]),.dout(n1040),.clk(gclk));
	jnot g0740(.din(w_G838_0),.dout(n1041),.clk(gclk));
	jand g0741(.dina(w_n797_3[0]),.dinb(w_n1041_1[1]),.dout(n1042),.clk(gclk));
	jand g0742(.dina(w_n799_3[0]),.dinb(w_G67_0[1]),.dout(n1043),.clk(gclk));
	jand g0743(.dina(w_n801_3[0]),.dinb(w_G70_0[1]),.dout(n1044),.clk(gclk));
	jor g0744(.dina(w_dff_B_d4K1Bo386_0),.dinb(n1043),.dout(n1045),.clk(gclk));
	jor g0745(.dina(w_dff_B_vpAFIKRV2_0),.dinb(n1042),.dout(n1046),.clk(gclk));
	jor g0746(.dina(w_dff_B_yvilTlyr0_0),.dinb(n1040),.dout(w_dff_A_XI6uvqqZ6_2),.clk(gclk));
	jand g0747(.dina(w_n1012_1[0]),.dinb(w_n840_4[0]),.dout(n1048),.clk(gclk));
	jand g0748(.dina(w_n843_4[0]),.dinb(w_n1014_1[0]),.dout(n1049),.clk(gclk));
	jand g0749(.dina(w_n845_4[0]),.dinb(w_G43_0[0]),.dout(n1050),.clk(gclk));
	jand g0750(.dina(w_n847_4[0]),.dinb(w_G37_0[0]),.dout(n1051),.clk(gclk));
	jor g0751(.dina(w_dff_B_9M5xc7r91_0),.dinb(n1050),.dout(n1052),.clk(gclk));
	jor g0752(.dina(w_dff_B_1rrl11Yh9_0),.dinb(n1049),.dout(n1053),.clk(gclk));
	jor g0753(.dina(w_dff_B_x28AR9oc9_0),.dinb(n1048),.dout(w_dff_A_DLFcmILU9_2),.clk(gclk));
	jand g0754(.dina(w_n1021_1[0]),.dinb(w_n840_3[2]),.dout(n1055),.clk(gclk));
	jand g0755(.dina(w_n843_3[2]),.dinb(w_n1023_1[0]),.dout(n1056),.clk(gclk));
	jand g0756(.dina(w_n845_3[2]),.dinb(w_G76_0[0]),.dout(n1057),.clk(gclk));
	jand g0757(.dina(w_n847_3[2]),.dinb(w_G20_0[0]),.dout(n1058),.clk(gclk));
	jor g0758(.dina(w_dff_B_4YYQYK7A9_0),.dinb(n1057),.dout(n1059),.clk(gclk));
	jor g0759(.dina(w_dff_B_cfNDjJPe0_0),.dinb(n1056),.dout(n1060),.clk(gclk));
	jor g0760(.dina(w_dff_B_mytJ3CSB9_0),.dinb(n1055),.dout(w_dff_A_YktHXzVq0_2),.clk(gclk));
	jand g0761(.dina(w_n1030_1[0]),.dinb(w_n840_3[1]),.dout(n1062),.clk(gclk));
	jand g0762(.dina(w_n843_3[1]),.dinb(w_n1032_1[0]),.dout(n1063),.clk(gclk));
	jand g0763(.dina(w_n845_3[1]),.dinb(w_G73_0[0]),.dout(n1064),.clk(gclk));
	jand g0764(.dina(w_n847_3[1]),.dinb(w_G17_0[0]),.dout(n1065),.clk(gclk));
	jor g0765(.dina(w_dff_B_pwMPdJHW0_0),.dinb(n1064),.dout(n1066),.clk(gclk));
	jor g0766(.dina(w_dff_B_v63e2pER8_0),.dinb(n1063),.dout(n1067),.clk(gclk));
	jor g0767(.dina(w_dff_B_GrUuGhbS2_0),.dinb(n1062),.dout(w_dff_A_cyMtHO7V5_2),.clk(gclk));
	jand g0768(.dina(w_n1039_1[0]),.dinb(w_n840_3[0]),.dout(n1069),.clk(gclk));
	jand g0769(.dina(w_n843_3[0]),.dinb(w_n1041_1[0]),.dout(n1070),.clk(gclk));
	jand g0770(.dina(w_n845_3[0]),.dinb(w_G67_0[0]),.dout(n1071),.clk(gclk));
	jand g0771(.dina(w_n847_3[0]),.dinb(w_G70_0[0]),.dout(n1072),.clk(gclk));
	jor g0772(.dina(w_dff_B_4tTd2lKx5_0),.dinb(n1071),.dout(n1073),.clk(gclk));
	jor g0773(.dina(w_dff_B_YZqsccn93_0),.dinb(n1070),.dout(n1074),.clk(gclk));
	jor g0774(.dina(w_dff_B_pIpn7ApU6_0),.dinb(n1069),.dout(w_dff_A_UsxZO5xA4_2),.clk(gclk));
	jand g0775(.dina(w_n985_4[0]),.dinb(w_n1012_0[2]),.dout(n1076),.clk(gclk));
	jand g0776(.dina(w_n988_4[0]),.dinb(w_n1014_0[2]),.dout(n1077),.clk(gclk));
	jand g0777(.dina(w_n990_4[0]),.dinb(w_G200_0[1]),.dout(n1078),.clk(gclk));
	jand g0778(.dina(w_n992_4[0]),.dinb(w_G170_0[1]),.dout(n1079),.clk(gclk));
	jor g0779(.dina(w_dff_B_Rge1IOJ90_0),.dinb(n1078),.dout(n1080),.clk(gclk));
	jor g0780(.dina(w_dff_B_NZAe3sJK5_0),.dinb(n1077),.dout(n1081),.clk(gclk));
	jor g0781(.dina(w_dff_B_i4lPnUWI4_0),.dinb(n1076),.dout(n1082),.clk(gclk));
	jand g0782(.dina(n1082),.dinb(w_G137_8[2]),.dout(w_dff_A_6jd38nub0_2),.clk(gclk));
	jand g0783(.dina(w_n985_3[2]),.dinb(w_n1039_0[2]),.dout(n1084),.clk(gclk));
	jand g0784(.dina(w_n988_3[2]),.dinb(w_n1041_0[2]),.dout(n1085),.clk(gclk));
	jand g0785(.dina(w_n990_3[2]),.dinb(w_G188_0[1]),.dout(n1086),.clk(gclk));
	jand g0786(.dina(w_n992_3[2]),.dinb(w_G158_0[1]),.dout(n1087),.clk(gclk));
	jor g0787(.dina(w_dff_B_KuXXw29b6_0),.dinb(n1086),.dout(n1088),.clk(gclk));
	jor g0788(.dina(w_dff_B_jFd1qzXD8_0),.dinb(n1085),.dout(n1089),.clk(gclk));
	jor g0789(.dina(w_dff_B_1H19wOa74_0),.dinb(n1084),.dout(n1090),.clk(gclk));
	jand g0790(.dina(n1090),.dinb(w_G137_8[1]),.dout(w_dff_A_OpM8B9au0_2),.clk(gclk));
	jand g0791(.dina(w_n985_3[1]),.dinb(w_n1030_0[2]),.dout(n1092),.clk(gclk));
	jand g0792(.dina(w_n988_3[1]),.dinb(w_n1032_0[2]),.dout(n1093),.clk(gclk));
	jand g0793(.dina(w_n990_3[1]),.dinb(w_G155_0[1]),.dout(n1094),.clk(gclk));
	jand g0794(.dina(w_n992_3[1]),.dinb(w_G152_0[1]),.dout(n1095),.clk(gclk));
	jor g0795(.dina(w_dff_B_JL4tlOpu9_0),.dinb(n1094),.dout(n1096),.clk(gclk));
	jor g0796(.dina(w_dff_B_j2lnXHmC3_0),.dinb(n1093),.dout(n1097),.clk(gclk));
	jor g0797(.dina(w_dff_B_aVoZ8Ga37_0),.dinb(n1092),.dout(n1098),.clk(gclk));
	jand g0798(.dina(n1098),.dinb(w_G137_8[0]),.dout(w_dff_A_udMizoxK1_2),.clk(gclk));
	jand g0799(.dina(w_n985_3[0]),.dinb(w_n1021_0[2]),.dout(n1100),.clk(gclk));
	jand g0800(.dina(w_n988_3[0]),.dinb(w_n1023_0[2]),.dout(n1101),.clk(gclk));
	jand g0801(.dina(w_n990_3[0]),.dinb(w_G149_0[1]),.dout(n1102),.clk(gclk));
	jand g0802(.dina(w_n992_3[0]),.dinb(w_G146_0[1]),.dout(n1103),.clk(gclk));
	jor g0803(.dina(w_dff_B_ZRYI2TIt9_0),.dinb(n1102),.dout(n1104),.clk(gclk));
	jor g0804(.dina(w_dff_B_6HOKj66b5_0),.dinb(n1101),.dout(n1105),.clk(gclk));
	jor g0805(.dina(w_dff_B_9CDm9T0x5_0),.dinb(n1100),.dout(n1106),.clk(gclk));
	jand g0806(.dina(n1106),.dinb(w_G137_7[2]),.dout(w_dff_A_TCP58EKm3_2),.clk(gclk));
	jand g0807(.dina(w_n999_4[0]),.dinb(w_n1012_0[1]),.dout(n1108),.clk(gclk));
	jand g0808(.dina(w_n1002_4[0]),.dinb(w_n1014_0[1]),.dout(n1109),.clk(gclk));
	jand g0809(.dina(w_n1004_4[0]),.dinb(w_G200_0[0]),.dout(n1110),.clk(gclk));
	jand g0810(.dina(w_n1006_4[0]),.dinb(w_G170_0[0]),.dout(n1111),.clk(gclk));
	jor g0811(.dina(w_dff_B_Gg9m0Kkv7_0),.dinb(n1110),.dout(n1112),.clk(gclk));
	jor g0812(.dina(w_dff_B_SbyRTDjy5_0),.dinb(n1109),.dout(n1113),.clk(gclk));
	jor g0813(.dina(w_dff_B_l1zv4hd97_0),.dinb(n1108),.dout(n1114),.clk(gclk));
	jand g0814(.dina(n1114),.dinb(w_G137_7[1]),.dout(w_dff_A_QvBFmF6Z6_2),.clk(gclk));
	jand g0815(.dina(w_n999_3[2]),.dinb(w_n1039_0[1]),.dout(n1116),.clk(gclk));
	jand g0816(.dina(w_n1002_3[2]),.dinb(w_n1041_0[1]),.dout(n1117),.clk(gclk));
	jand g0817(.dina(w_n1004_3[2]),.dinb(w_G188_0[0]),.dout(n1118),.clk(gclk));
	jand g0818(.dina(w_n1006_3[2]),.dinb(w_G158_0[0]),.dout(n1119),.clk(gclk));
	jor g0819(.dina(w_dff_B_dLAyJeXu7_0),.dinb(n1118),.dout(n1120),.clk(gclk));
	jor g0820(.dina(w_dff_B_FCy4cNJc8_0),.dinb(n1117),.dout(n1121),.clk(gclk));
	jor g0821(.dina(w_dff_B_i29EUwTc3_0),.dinb(n1116),.dout(n1122),.clk(gclk));
	jand g0822(.dina(n1122),.dinb(w_G137_7[0]),.dout(w_dff_A_njPQMHMP1_2),.clk(gclk));
	jand g0823(.dina(w_n999_3[1]),.dinb(w_n1030_0[1]),.dout(n1124),.clk(gclk));
	jand g0824(.dina(w_n1002_3[1]),.dinb(w_n1032_0[1]),.dout(n1125),.clk(gclk));
	jand g0825(.dina(w_n1004_3[1]),.dinb(w_G155_0[0]),.dout(n1126),.clk(gclk));
	jand g0826(.dina(w_n1006_3[1]),.dinb(w_G152_0[0]),.dout(n1127),.clk(gclk));
	jor g0827(.dina(w_dff_B_iywwfrfp0_0),.dinb(n1126),.dout(n1128),.clk(gclk));
	jor g0828(.dina(w_dff_B_DgGrCXuz6_0),.dinb(n1125),.dout(n1129),.clk(gclk));
	jor g0829(.dina(w_dff_B_db45aS7f7_0),.dinb(n1124),.dout(n1130),.clk(gclk));
	jand g0830(.dina(n1130),.dinb(w_G137_6[2]),.dout(w_dff_A_ZS1XpX9r3_2),.clk(gclk));
	jand g0831(.dina(w_n999_3[0]),.dinb(w_n1021_0[1]),.dout(n1132),.clk(gclk));
	jand g0832(.dina(w_n1002_3[0]),.dinb(w_n1023_0[1]),.dout(n1133),.clk(gclk));
	jand g0833(.dina(w_n1004_3[0]),.dinb(w_G149_0[0]),.dout(n1134),.clk(gclk));
	jand g0834(.dina(w_n1006_3[0]),.dinb(w_G146_0[0]),.dout(n1135),.clk(gclk));
	jor g0835(.dina(w_dff_B_V1GNE4et7_0),.dinb(n1134),.dout(n1136),.clk(gclk));
	jor g0836(.dina(w_dff_B_WWmRkjpa6_0),.dinb(n1133),.dout(n1137),.clk(gclk));
	jor g0837(.dina(w_dff_B_wvmvDo3N4_0),.dinb(n1132),.dout(n1138),.clk(gclk));
	jand g0838(.dina(n1138),.dinb(w_G137_6[1]),.dout(w_dff_A_zWSShnYZ7_2),.clk(gclk));
	jand g0839(.dina(w_n789_0[1]),.dinb(w_G3724_0[2]),.dout(n1140),.clk(gclk));
	jnot g0840(.din(w_G3717_0[1]),.dout(n1141),.clk(gclk));
	jnot g0841(.din(w_G3724_0[1]),.dout(n1142),.clk(gclk));
	jand g0842(.dina(w_n1142_0[1]),.dinb(w_G123_0[1]),.dout(n1143),.clk(gclk));
	jor g0843(.dina(n1143),.dinb(w_dff_B_ugPAGpWl0_1),.dout(n1144),.clk(gclk));
	jor g0844(.dina(w_dff_B_i7iBOFlZ4_0),.dinb(n1140),.dout(n1145),.clk(gclk));
	jnot g0845(.din(G135),.dout(n1146),.clk(gclk));
	jnot g0846(.din(G4115),.dout(n1147),.clk(gclk));
	jor g0847(.dina(n1147),.dinb(n1146),.dout(n1148),.clk(gclk));
	jxor g0848(.dina(w_n636_0[1]),.dinb(w_G132_0[1]),.dout(n1149),.clk(gclk));
	jand g0849(.dina(n1149),.dinb(w_G3724_0[0]),.dout(n1150),.clk(gclk));
	jnot g0850(.din(w_n401_0[1]),.dout(n1151),.clk(gclk));
	jand g0851(.dina(w_n1151_0[1]),.dinb(w_n1142_0[0]),.dout(n1152),.clk(gclk));
	jor g0852(.dina(n1152),.dinb(w_G3717_0[0]),.dout(n1153),.clk(gclk));
	jor g0853(.dina(n1153),.dinb(w_dff_B_HixqNAtj8_1),.dout(n1154),.clk(gclk));
	jand g0854(.dina(n1154),.dinb(w_dff_B_eI2359Qg3_1),.dout(n1155),.clk(gclk));
	jand g0855(.dina(w_dff_B_j74uReLR5_0),.dinb(n1145),.dout(w_dff_A_l4yz9gMX7_2),.clk(gclk));
	jor g0856(.dina(w_n783_0[1]),.dinb(w_n640_0[2]),.dout(n1157),.clk(gclk));
	jxor g0857(.dina(n1157),.dinb(w_G132_0[0]),.dout(w_dff_A_L9zsaGmQ8_2),.clk(gclk));
	jand g0858(.dina(w_n789_0[0]),.dinb(w_n747_2[1]),.dout(n1159),.clk(gclk));
	jand g0859(.dina(w_n753_5[0]),.dinb(w_G123_0[0]),.dout(n1160),.clk(gclk));
	jand g0860(.dina(w_n751_1[1]),.dinb(w_n1151_0[0]),.dout(n1161),.clk(gclk));
	jor g0861(.dina(n1161),.dinb(w_dff_B_WSVXGEBq2_1),.dout(n1162),.clk(gclk));
	jor g0862(.dina(w_dff_B_dJTTVpsB3_0),.dinb(n1159),.dout(n1163),.clk(gclk));
	jnot g0863(.din(w_n1163_1[2]),.dout(w_dff_A_9EZjqA4L7_1),.clk(gclk));
	jor g0864(.dina(w_n972_0[0]),.dinb(w_n748_2[0]),.dout(n1165),.clk(gclk));
	jand g0865(.dina(w_n751_1[0]),.dinb(w_n407_0[0]),.dout(n1166),.clk(gclk));
	jand g0866(.dina(w_n753_4[2]),.dinb(w_dff_B_qIHigijf7_1),.dout(n1167),.clk(gclk));
	jor g0867(.dina(w_dff_B_e3bAn2re2_0),.dinb(n1166),.dout(n1168),.clk(gclk));
	jnot g0868(.din(n1168),.dout(n1169),.clk(gclk));
	jand g0869(.dina(w_dff_B_5EJPR0oB7_0),.dinb(n1165),.dout(G826_fa_),.clk(gclk));
	jor g0870(.dina(w_n971_0[0]),.dinb(w_n748_1[2]),.dout(n1171),.clk(gclk));
	jor g0871(.dina(w_n765_3[0]),.dinb(w_n372_0[1]),.dout(n1172),.clk(gclk));
	jand g0872(.dina(w_n753_4[1]),.dinb(w_dff_B_qH7SRKVN3_1),.dout(n1173),.clk(gclk));
	jnot g0873(.din(n1173),.dout(n1174),.clk(gclk));
	jand g0874(.dina(w_dff_B_UWtMXrMa8_0),.dinb(n1172),.dout(n1175),.clk(gclk));
	jand g0875(.dina(w_dff_B_brMOSBEK6_0),.dinb(n1171),.dout(G828_fa_),.clk(gclk));
	jand g0876(.dina(w_n973_0[0]),.dinb(w_n747_2[0]),.dout(n1177),.clk(gclk));
	jnot g0877(.din(n1177),.dout(n1178),.clk(gclk));
	jor g0878(.dina(w_n765_2[2]),.dinb(w_n383_0[1]),.dout(n1179),.clk(gclk));
	jand g0879(.dina(w_n753_4[0]),.dinb(w_dff_B_ITDwAj4G9_1),.dout(n1180),.clk(gclk));
	jnot g0880(.din(n1180),.dout(n1181),.clk(gclk));
	jand g0881(.dina(w_dff_B_rFDNt3jY9_0),.dinb(n1179),.dout(n1182),.clk(gclk));
	jand g0882(.dina(w_dff_B_Z8qSrzYS1_0),.dinb(n1178),.dout(G830_fa_),.clk(gclk));
	jnot g0883(.din(w_G1000_0),.dout(n1184),.clk(gclk));
	jand g0884(.dina(w_G559_0[0]),.dinb(w_G245_0[0]),.dout(n1185),.clk(gclk));
	jand g0885(.dina(n1185),.dinb(w_n318_0[0]),.dout(n1186),.clk(gclk));
	jand g0886(.dina(n1186),.dinb(w_G601_0),.dout(n1187),.clk(gclk));
	jand g0887(.dina(w_dff_B_7qWwFGV17_0),.dinb(w_n661_0[0]),.dout(n1188),.clk(gclk));
	jand g0888(.dina(n1188),.dinb(w_n671_0[0]),.dout(n1189),.clk(gclk));
	jand g0889(.dina(w_dff_B_6yWgKtOw7_0),.dinb(w_n914_0[0]),.dout(n1190),.clk(gclk));
	jand g0890(.dina(n1190),.dinb(w_dff_B_GjqMQ1wZ2_1),.dout(w_dff_A_nqVLCUVr3_2),.clk(gclk));
	jand g0891(.dina(w_n941_0[0]),.dinb(w_n747_1[2]),.dout(n1192),.clk(gclk));
	jnot g0892(.din(w_n528_0[1]),.dout(n1193),.clk(gclk));
	jand g0893(.dina(w_n751_0[2]),.dinb(n1193),.dout(n1194),.clk(gclk));
	jand g0894(.dina(w_n753_3[2]),.dinb(w_dff_B_CjpD4YzR1_1),.dout(n1195),.clk(gclk));
	jor g0895(.dina(w_dff_B_KwgV3T4n3_0),.dinb(n1194),.dout(n1196),.clk(gclk));
	jor g0896(.dina(w_dff_B_2XMIVhUw3_0),.dinb(n1192),.dout(n1197),.clk(gclk));
	jnot g0897(.din(w_n1197_1[2]),.dout(w_dff_A_O5MACyFk6_1),.clk(gclk));
	jand g0898(.dina(w_n946_0[0]),.dinb(w_n747_1[1]),.dout(n1199),.clk(gclk));
	jor g0899(.dina(w_n765_2[1]),.dinb(w_n551_0[0]),.dout(n1200),.clk(gclk));
	jand g0900(.dina(w_n753_3[1]),.dinb(w_dff_B_evsv9m3f0_1),.dout(n1201),.clk(gclk));
	jnot g0901(.din(n1201),.dout(n1202),.clk(gclk));
	jand g0902(.dina(w_dff_B_8vNbqRXJ6_0),.dinb(n1200),.dout(n1203),.clk(gclk));
	jnot g0903(.din(n1203),.dout(n1204),.clk(gclk));
	jor g0904(.dina(w_dff_B_pRA1cafs6_0),.dinb(n1199),.dout(n1205),.clk(gclk));
	jnot g0905(.din(w_n1205_1[2]),.dout(w_dff_A_qeZz187w9_1),.clk(gclk));
	jor g0906(.dina(w_n953_0[0]),.dinb(w_n748_1[1]),.dout(n1207),.clk(gclk));
	jor g0907(.dina(w_n765_2[0]),.dinb(w_n517_0[0]),.dout(n1208),.clk(gclk));
	jand g0908(.dina(w_n753_3[0]),.dinb(w_dff_B_pPteiRlH7_1),.dout(n1209),.clk(gclk));
	jnot g0909(.din(n1209),.dout(n1210),.clk(gclk));
	jand g0910(.dina(w_dff_B_cTovec442_0),.dinb(n1208),.dout(n1211),.clk(gclk));
	jand g0911(.dina(w_dff_B_N1JcnImR0_0),.dinb(n1207),.dout(G867_fa_),.clk(gclk));
	jand g0912(.dina(w_n954_0[0]),.dinb(w_n747_1[0]),.dout(n1213),.clk(gclk));
	jnot g0913(.din(n1213),.dout(n1214),.clk(gclk));
	jor g0914(.dina(w_n765_1[2]),.dinb(w_n540_0[0]),.dout(n1215),.clk(gclk));
	jand g0915(.dina(w_n753_2[2]),.dinb(w_dff_B_cJA6FlcG8_1),.dout(n1216),.clk(gclk));
	jnot g0916(.din(n1216),.dout(n1217),.clk(gclk));
	jand g0917(.dina(w_dff_B_D0xwtLV79_0),.dinb(n1215),.dout(n1218),.clk(gclk));
	jand g0918(.dina(w_dff_B_CoRr7QPr6_0),.dinb(n1214),.dout(G869_fa_),.clk(gclk));
	jand g0919(.dina(w_n1197_1[1]),.dinb(w_n840_2[2]),.dout(n1220),.clk(gclk));
	jand g0920(.dina(w_n1163_1[1]),.dinb(w_n843_2[2]),.dout(n1221),.clk(gclk));
	jand g0921(.dina(w_n845_2[2]),.dinb(w_G109_0[1]),.dout(n1222),.clk(gclk));
	jand g0922(.dina(w_n847_2[2]),.dinb(w_G106_0[1]),.dout(n1223),.clk(gclk));
	jor g0923(.dina(w_dff_B_WQeYJm0f2_0),.dinb(n1222),.dout(n1224),.clk(gclk));
	jor g0924(.dina(w_dff_B_foFSaU8A0_0),.dinb(n1221),.dout(n1225),.clk(gclk));
	jor g0925(.dina(n1225),.dinb(n1220),.dout(w_dff_A_EPXAZVpy7_2),.clk(gclk));
	jand g0926(.dina(w_n1197_1[0]),.dinb(w_n793_2[2]),.dout(n1227),.clk(gclk));
	jand g0927(.dina(w_n1163_1[0]),.dinb(w_n797_2[2]),.dout(n1228),.clk(gclk));
	jand g0928(.dina(w_n799_2[2]),.dinb(w_G109_0[0]),.dout(n1229),.clk(gclk));
	jand g0929(.dina(w_n801_2[2]),.dinb(w_G106_0[0]),.dout(n1230),.clk(gclk));
	jor g0930(.dina(w_dff_B_8rv1HNPK0_0),.dinb(n1229),.dout(n1231),.clk(gclk));
	jor g0931(.dina(w_dff_B_ZNrBUawd7_0),.dinb(n1228),.dout(n1232),.clk(gclk));
	jor g0932(.dina(n1232),.dinb(n1227),.dout(w_dff_A_A0bT2Z0q4_2),.clk(gclk));
	jand g0933(.dina(w_n1205_1[1]),.dinb(w_n793_2[1]),.dout(n1234),.clk(gclk));
	jnot g0934(.din(w_G826_0),.dout(n1235),.clk(gclk));
	jand g0935(.dina(w_n1235_1[1]),.dinb(w_n797_2[1]),.dout(n1236),.clk(gclk));
	jand g0936(.dina(w_n799_2[1]),.dinb(w_G46_0[1]),.dout(n1237),.clk(gclk));
	jand g0937(.dina(w_n801_2[1]),.dinb(w_G49_0[1]),.dout(n1238),.clk(gclk));
	jor g0938(.dina(w_dff_B_Wf1pMfSH9_0),.dinb(n1237),.dout(n1239),.clk(gclk));
	jor g0939(.dina(w_dff_B_bexrAVvW0_0),.dinb(n1236),.dout(n1240),.clk(gclk));
	jor g0940(.dina(n1240),.dinb(n1234),.dout(w_dff_A_aSx5mPAn3_2),.clk(gclk));
	jnot g0941(.din(w_G867_0),.dout(n1242),.clk(gclk));
	jand g0942(.dina(w_n1242_1[1]),.dinb(w_n793_2[0]),.dout(n1243),.clk(gclk));
	jnot g0943(.din(w_G828_0),.dout(n1244),.clk(gclk));
	jand g0944(.dina(w_n1244_1[1]),.dinb(w_n797_2[0]),.dout(n1245),.clk(gclk));
	jand g0945(.dina(w_n799_2[0]),.dinb(w_G100_0[1]),.dout(n1246),.clk(gclk));
	jand g0946(.dina(w_n801_2[0]),.dinb(w_G103_0[1]),.dout(n1247),.clk(gclk));
	jor g0947(.dina(w_dff_B_leJxw7Py9_0),.dinb(n1246),.dout(n1248),.clk(gclk));
	jor g0948(.dina(w_dff_B_gAKDul2C1_0),.dinb(n1245),.dout(n1249),.clk(gclk));
	jor g0949(.dina(n1249),.dinb(n1243),.dout(w_dff_A_EvzIhjy47_2),.clk(gclk));
	jnot g0950(.din(w_G869_0),.dout(n1251),.clk(gclk));
	jand g0951(.dina(w_n1251_1[1]),.dinb(w_n793_1[2]),.dout(n1252),.clk(gclk));
	jnot g0952(.din(w_G830_0),.dout(n1253),.clk(gclk));
	jand g0953(.dina(w_n1253_1[1]),.dinb(w_n797_1[2]),.dout(n1254),.clk(gclk));
	jand g0954(.dina(w_n799_1[2]),.dinb(w_G91_0[1]),.dout(n1255),.clk(gclk));
	jand g0955(.dina(w_n801_1[2]),.dinb(w_G40_0[1]),.dout(n1256),.clk(gclk));
	jor g0956(.dina(w_dff_B_8wzj2M7N8_0),.dinb(n1255),.dout(n1257),.clk(gclk));
	jor g0957(.dina(w_dff_B_kbBNPsoE5_0),.dinb(n1254),.dout(n1258),.clk(gclk));
	jor g0958(.dina(n1258),.dinb(n1252),.dout(w_dff_A_5IAg5QGE8_2),.clk(gclk));
	jand g0959(.dina(w_n1205_1[0]),.dinb(w_n840_2[1]),.dout(n1260),.clk(gclk));
	jand g0960(.dina(w_n1235_1[0]),.dinb(w_n843_2[1]),.dout(n1261),.clk(gclk));
	jand g0961(.dina(w_n845_2[1]),.dinb(w_G46_0[0]),.dout(n1262),.clk(gclk));
	jand g0962(.dina(w_n847_2[1]),.dinb(w_G49_0[0]),.dout(n1263),.clk(gclk));
	jor g0963(.dina(w_dff_B_EykvKAbE6_0),.dinb(n1262),.dout(n1264),.clk(gclk));
	jor g0964(.dina(w_dff_B_OeaKwgd32_0),.dinb(n1261),.dout(n1265),.clk(gclk));
	jor g0965(.dina(n1265),.dinb(n1260),.dout(w_dff_A_KRUM41us5_2),.clk(gclk));
	jand g0966(.dina(w_n1242_1[0]),.dinb(w_n840_2[0]),.dout(n1267),.clk(gclk));
	jand g0967(.dina(w_n1244_1[0]),.dinb(w_n843_2[0]),.dout(n1268),.clk(gclk));
	jand g0968(.dina(w_n845_2[0]),.dinb(w_G100_0[0]),.dout(n1269),.clk(gclk));
	jand g0969(.dina(w_n847_2[0]),.dinb(w_G103_0[0]),.dout(n1270),.clk(gclk));
	jor g0970(.dina(w_dff_B_TUIbUdjG8_0),.dinb(n1269),.dout(n1271),.clk(gclk));
	jor g0971(.dina(w_dff_B_gqepe3so4_0),.dinb(n1268),.dout(n1272),.clk(gclk));
	jor g0972(.dina(n1272),.dinb(n1267),.dout(w_dff_A_RrTJUjUs0_2),.clk(gclk));
	jand g0973(.dina(w_n1251_1[0]),.dinb(w_n840_1[2]),.dout(n1274),.clk(gclk));
	jand g0974(.dina(w_n1253_1[0]),.dinb(w_n843_1[2]),.dout(n1275),.clk(gclk));
	jand g0975(.dina(w_n845_1[2]),.dinb(w_G91_0[0]),.dout(n1276),.clk(gclk));
	jand g0976(.dina(w_n847_1[2]),.dinb(w_G40_0[0]),.dout(n1277),.clk(gclk));
	jor g0977(.dina(w_dff_B_O0tS13sh8_0),.dinb(n1276),.dout(n1278),.clk(gclk));
	jor g0978(.dina(w_dff_B_k1BaaJBX6_0),.dinb(n1275),.dout(n1279),.clk(gclk));
	jor g0979(.dina(n1279),.dinb(n1274),.dout(w_dff_A_sdnfD5209_2),.clk(gclk));
	jand g0980(.dina(w_n1251_0[2]),.dinb(w_n985_2[2]),.dout(n1281),.clk(gclk));
	jand g0981(.dina(w_n1253_0[2]),.dinb(w_n988_2[2]),.dout(n1282),.clk(gclk));
	jand g0982(.dina(w_n990_2[2]),.dinb(w_G203_0[1]),.dout(n1283),.clk(gclk));
	jand g0983(.dina(w_n992_2[2]),.dinb(w_G173_0[1]),.dout(n1284),.clk(gclk));
	jor g0984(.dina(w_dff_B_ATcF3x672_0),.dinb(n1283),.dout(n1285),.clk(gclk));
	jor g0985(.dina(w_dff_B_qH4ghL7g7_0),.dinb(n1282),.dout(n1286),.clk(gclk));
	jor g0986(.dina(n1286),.dinb(n1281),.dout(n1287),.clk(gclk));
	jand g0987(.dina(n1287),.dinb(w_G137_6[0]),.dout(w_dff_A_Gwj90k1Q2_2),.clk(gclk));
	jand g0988(.dina(w_n1242_0[2]),.dinb(w_n985_2[1]),.dout(n1289),.clk(gclk));
	jand g0989(.dina(w_n1244_0[2]),.dinb(w_n988_2[1]),.dout(n1290),.clk(gclk));
	jand g0990(.dina(w_n990_2[1]),.dinb(w_G197_0[1]),.dout(n1291),.clk(gclk));
	jand g0991(.dina(w_n992_2[1]),.dinb(w_G167_0[1]),.dout(n1292),.clk(gclk));
	jor g0992(.dina(w_dff_B_QiyBP5GP1_0),.dinb(n1291),.dout(n1293),.clk(gclk));
	jor g0993(.dina(w_dff_B_M3NHt4gJ0_0),.dinb(n1290),.dout(n1294),.clk(gclk));
	jor g0994(.dina(n1294),.dinb(n1289),.dout(n1295),.clk(gclk));
	jand g0995(.dina(n1295),.dinb(w_G137_5[2]),.dout(w_dff_A_G2E6wyy35_2),.clk(gclk));
	jand g0996(.dina(w_n1205_0[2]),.dinb(w_n985_2[0]),.dout(n1297),.clk(gclk));
	jand g0997(.dina(w_n1235_0[2]),.dinb(w_n988_2[0]),.dout(n1298),.clk(gclk));
	jand g0998(.dina(w_n990_2[0]),.dinb(w_G194_0[1]),.dout(n1299),.clk(gclk));
	jand g0999(.dina(w_n992_2[0]),.dinb(w_G164_0[1]),.dout(n1300),.clk(gclk));
	jor g1000(.dina(w_dff_B_utLN8AQu0_0),.dinb(n1299),.dout(n1301),.clk(gclk));
	jor g1001(.dina(w_dff_B_3harrfKT3_0),.dinb(n1298),.dout(n1302),.clk(gclk));
	jor g1002(.dina(n1302),.dinb(n1297),.dout(n1303),.clk(gclk));
	jand g1003(.dina(n1303),.dinb(w_G137_5[1]),.dout(w_dff_A_sGgb8Vsx5_2),.clk(gclk));
	jand g1004(.dina(w_n1197_0[2]),.dinb(w_n985_1[2]),.dout(n1305),.clk(gclk));
	jand g1005(.dina(w_n1163_0[2]),.dinb(w_n988_1[2]),.dout(n1306),.clk(gclk));
	jand g1006(.dina(w_n990_1[2]),.dinb(w_G191_0[1]),.dout(n1307),.clk(gclk));
	jand g1007(.dina(w_n992_1[2]),.dinb(w_G161_0[1]),.dout(n1308),.clk(gclk));
	jor g1008(.dina(w_dff_B_GkzyK1x01_0),.dinb(n1307),.dout(n1309),.clk(gclk));
	jor g1009(.dina(w_dff_B_5tYYOmDO1_0),.dinb(n1306),.dout(n1310),.clk(gclk));
	jor g1010(.dina(n1310),.dinb(n1305),.dout(n1311),.clk(gclk));
	jand g1011(.dina(n1311),.dinb(w_G137_5[0]),.dout(w_dff_A_7PhnTXaZ8_2),.clk(gclk));
	jand g1012(.dina(w_n1251_0[1]),.dinb(w_n999_2[2]),.dout(n1313),.clk(gclk));
	jand g1013(.dina(w_n1253_0[1]),.dinb(w_n1002_2[2]),.dout(n1314),.clk(gclk));
	jand g1014(.dina(w_n1004_2[2]),.dinb(w_G203_0[0]),.dout(n1315),.clk(gclk));
	jand g1015(.dina(w_n1006_2[2]),.dinb(w_G173_0[0]),.dout(n1316),.clk(gclk));
	jor g1016(.dina(w_dff_B_MjGKjvwP7_0),.dinb(n1315),.dout(n1317),.clk(gclk));
	jor g1017(.dina(w_dff_B_cvumRequ5_0),.dinb(n1314),.dout(n1318),.clk(gclk));
	jor g1018(.dina(n1318),.dinb(n1313),.dout(n1319),.clk(gclk));
	jand g1019(.dina(n1319),.dinb(w_G137_4[2]),.dout(w_dff_A_RjIELs5s6_2),.clk(gclk));
	jand g1020(.dina(w_n1242_0[1]),.dinb(w_n999_2[1]),.dout(n1321),.clk(gclk));
	jand g1021(.dina(w_n1244_0[1]),.dinb(w_n1002_2[1]),.dout(n1322),.clk(gclk));
	jand g1022(.dina(w_n1004_2[1]),.dinb(w_G197_0[0]),.dout(n1323),.clk(gclk));
	jand g1023(.dina(w_n1006_2[1]),.dinb(w_G167_0[0]),.dout(n1324),.clk(gclk));
	jor g1024(.dina(w_dff_B_Nh4RGfHi0_0),.dinb(n1323),.dout(n1325),.clk(gclk));
	jor g1025(.dina(w_dff_B_7xflPzTx9_0),.dinb(n1322),.dout(n1326),.clk(gclk));
	jor g1026(.dina(n1326),.dinb(n1321),.dout(n1327),.clk(gclk));
	jand g1027(.dina(n1327),.dinb(w_G137_4[1]),.dout(w_dff_A_nq2iXq3a8_2),.clk(gclk));
	jand g1028(.dina(w_n1205_0[1]),.dinb(w_n999_2[0]),.dout(n1329),.clk(gclk));
	jand g1029(.dina(w_n1235_0[1]),.dinb(w_n1002_2[0]),.dout(n1330),.clk(gclk));
	jand g1030(.dina(w_n1004_2[0]),.dinb(w_G194_0[0]),.dout(n1331),.clk(gclk));
	jand g1031(.dina(w_n1006_2[0]),.dinb(w_G164_0[0]),.dout(n1332),.clk(gclk));
	jor g1032(.dina(w_dff_B_b4LZq0Iw7_0),.dinb(n1331),.dout(n1333),.clk(gclk));
	jor g1033(.dina(w_dff_B_r8jmrCwB8_0),.dinb(n1330),.dout(n1334),.clk(gclk));
	jor g1034(.dina(n1334),.dinb(n1329),.dout(n1335),.clk(gclk));
	jand g1035(.dina(n1335),.dinb(w_G137_4[0]),.dout(w_dff_A_LZXvWiyX4_2),.clk(gclk));
	jand g1036(.dina(w_n1197_0[1]),.dinb(w_n999_1[2]),.dout(n1337),.clk(gclk));
	jand g1037(.dina(w_n1163_0[1]),.dinb(w_n1002_1[2]),.dout(n1338),.clk(gclk));
	jand g1038(.dina(w_n1004_1[2]),.dinb(w_G191_0[0]),.dout(n1339),.clk(gclk));
	jand g1039(.dina(w_n1006_1[2]),.dinb(w_G161_0[0]),.dout(n1340),.clk(gclk));
	jor g1040(.dina(w_dff_B_vnyIMFO61_0),.dinb(n1339),.dout(n1341),.clk(gclk));
	jor g1041(.dina(w_dff_B_Cz04OjIr1_0),.dinb(n1338),.dout(n1342),.clk(gclk));
	jor g1042(.dina(n1342),.dinb(n1337),.dout(n1343),.clk(gclk));
	jand g1043(.dina(n1343),.dinb(w_G137_3[2]),.dout(w_dff_A_wCM0Ubje4_2),.clk(gclk));
	jor g1044(.dina(w_G4091_2[0]),.dinb(G120),.dout(n1345),.clk(gclk));
	jand g1045(.dina(w_n435_0[2]),.dinb(w_G251_3[1]),.dout(n1346),.clk(gclk));
	jand g1046(.dina(w_G341_1[0]),.dinb(w_G248_4[0]),.dout(n1347),.clk(gclk));
	jor g1047(.dina(n1347),.dinb(w_n437_0[1]),.dout(n1348),.clk(gclk));
	jor g1048(.dina(n1348),.dinb(n1346),.dout(n1349),.clk(gclk));
	jand g1049(.dina(w_n435_0[1]),.dinb(w_n366_3[1]),.dout(n1350),.clk(gclk));
	jand g1050(.dina(w_G341_0[2]),.dinb(w_n368_4[0]),.dout(n1351),.clk(gclk));
	jor g1051(.dina(n1351),.dinb(w_G523_0[2]),.dout(n1352),.clk(gclk));
	jor g1052(.dina(n1352),.dinb(w_dff_B_G3JSTTyC0_1),.dout(n1353),.clk(gclk));
	jand g1053(.dina(n1353),.dinb(w_dff_B_ZC3lkNWB4_1),.dout(n1354),.clk(gclk));
	jxor g1054(.dina(w_n408_0[0]),.dinb(w_n401_0[0]),.dout(n1355),.clk(gclk));
	jxor g1055(.dina(w_n383_0[0]),.dinb(w_n372_0[0]),.dout(n1356),.clk(gclk));
	jxor g1056(.dina(n1356),.dinb(w_dff_B_hVArdk7n8_1),.dout(n1357),.clk(gclk));
	jxor g1057(.dina(n1357),.dinb(w_dff_B_Xn8RU2f01_1),.dout(n1358),.clk(gclk));
	jnot g1058(.din(w_n1358_0[1]),.dout(n1359),.clk(gclk));
	jor g1059(.dina(w_n410_0[1]),.dinb(w_G248_3[2]),.dout(n1360),.clk(gclk));
	jor g1060(.dina(w_G514_0[1]),.dinb(w_n368_3[2]),.dout(n1361),.clk(gclk));
	jand g1061(.dina(n1361),.dinb(n1360),.dout(n1362),.clk(gclk));
	jxor g1062(.dina(n1362),.dinb(w_n419_0[0]),.dout(n1363),.clk(gclk));
	jor g1063(.dina(w_G351_1[0]),.dinb(w_n402_1[2]),.dout(n1364),.clk(gclk));
	jor g1064(.dina(w_n385_0[2]),.dinb(w_n405_1[2]),.dout(n1365),.clk(gclk));
	jand g1065(.dina(n1365),.dinb(w_G534_0[1]),.dout(n1366),.clk(gclk));
	jand g1066(.dina(n1366),.dinb(w_dff_B_LBOSmfTe1_1),.dout(n1367),.clk(gclk));
	jor g1067(.dina(w_G351_0[2]),.dinb(w_G254_1[1]),.dout(n1368),.clk(gclk));
	jor g1068(.dina(w_n385_0[1]),.dinb(w_G242_1[1]),.dout(n1369),.clk(gclk));
	jand g1069(.dina(n1369),.dinb(w_n388_0[1]),.dout(n1370),.clk(gclk));
	jand g1070(.dina(n1370),.dinb(w_dff_B_QKm8l0wr0_1),.dout(n1371),.clk(gclk));
	jor g1071(.dina(n1371),.dinb(n1367),.dout(n1372),.clk(gclk));
	jand g1072(.dina(w_n424_1[0]),.dinb(w_G251_3[0]),.dout(n1373),.clk(gclk));
	jand g1073(.dina(w_G324_0[2]),.dinb(w_G248_3[1]),.dout(n1374),.clk(gclk));
	jor g1074(.dina(n1374),.dinb(w_n426_0[0]),.dout(n1375),.clk(gclk));
	jor g1075(.dina(n1375),.dinb(n1373),.dout(n1376),.clk(gclk));
	jand g1076(.dina(w_n424_0[2]),.dinb(w_n366_3[0]),.dout(n1377),.clk(gclk));
	jand g1077(.dina(w_G324_0[1]),.dinb(w_n368_3[1]),.dout(n1378),.clk(gclk));
	jor g1078(.dina(n1378),.dinb(w_G503_0[1]),.dout(n1379),.clk(gclk));
	jor g1079(.dina(n1379),.dinb(w_dff_B_MPpmLCTT3_1),.dout(n1380),.clk(gclk));
	jand g1080(.dina(n1380),.dinb(w_dff_B_nHvIWuat9_1),.dout(n1381),.clk(gclk));
	jxor g1081(.dina(n1381),.dinb(n1372),.dout(n1382),.clk(gclk));
	jxor g1082(.dina(n1382),.dinb(w_dff_B_sPMlff716_1),.dout(n1383),.clk(gclk));
	jnot g1083(.din(w_n1383_0[1]),.dout(n1384),.clk(gclk));
	jand g1084(.dina(w_n1383_0[0]),.dinb(n1359),.dout(n1385),.clk(gclk));
	jor g1085(.dina(n1385),.dinb(w_G4091_1[2]),.dout(n1386),.clk(gclk));
	jor g1086(.dina(n1345),.dinb(w_n746_1[0]),.dout(n1388),.clk(gclk));
	jand g1087(.dina(n1384),.dinb(w_n1358_0[0]),.dout(n1389),.clk(gclk));
	jor g1088(.dina(n1386),.dinb(w_dff_B_r7EWpylQ1_1),.dout(n1390),.clk(gclk));
	jand g1089(.dina(n1390),.dinb(w_n746_0[2]),.dout(n1391),.clk(gclk));
	jnot g1090(.din(w_n1391_0[1]),.dout(n1392),.clk(gclk));
	jand g1091(.dina(w_n633_0[2]),.dinb(w_G2174_0[2]),.dout(n1393),.clk(gclk));
	jor g1092(.dina(w_dff_B_sTEgEJtc9_0),.dinb(w_n732_0[0]),.dout(n1394),.clk(gclk));
	jand g1093(.dina(w_n736_0[0]),.dinb(w_n640_0[1]),.dout(n1395),.clk(gclk));
	jor g1094(.dina(w_n740_0[0]),.dinb(w_n641_0[0]),.dout(n1396),.clk(gclk));
	jand g1095(.dina(n1396),.dinb(w_n646_0[0]),.dout(n1397),.clk(gclk));
	jor g1096(.dina(n1397),.dinb(w_dff_B_4M2MQAlr4_1),.dout(n1398),.clk(gclk));
	jnot g1097(.din(w_n1398_0[1]),.dout(n1399),.clk(gclk));
	jand g1098(.dina(w_n1399_0[1]),.dinb(w_n739_0[2]),.dout(n1400),.clk(gclk));
	jnot g1099(.din(w_n739_0[1]),.dout(n1401),.clk(gclk));
	jand g1100(.dina(w_n1398_0[0]),.dinb(w_dff_B_ztEuUki02_1),.dout(n1402),.clk(gclk));
	jor g1101(.dina(n1402),.dinb(w_n651_0[1]),.dout(n1403),.clk(gclk));
	jor g1102(.dina(n1403),.dinb(n1400),.dout(n1404),.clk(gclk));
	jand g1103(.dina(w_dff_B_3RbFhSx97_0),.dinb(w_n1394_0[1]),.dout(n1405),.clk(gclk));
	jnot g1104(.din(w_n1394_0[0]),.dout(n1406),.clk(gclk));
	jxor g1105(.dina(w_n1399_0[0]),.dinb(w_n968_0[0]),.dout(n1407),.clk(gclk));
	jand g1106(.dina(w_dff_B_qscW8IVx3_0),.dinb(n1406),.dout(n1408),.clk(gclk));
	jor g1107(.dina(n1408),.dinb(w_dff_B_uCKs5HVf6_1),.dout(n1409),.clk(gclk));
	jnot g1108(.din(w_n1409_0[1]),.dout(n1410),.clk(gclk));
	jxor g1109(.dina(w_n629_0[0]),.dinb(w_n625_0[0]),.dout(n1411),.clk(gclk));
	jnot g1110(.din(w_n1411_0[1]),.dout(n1412),.clk(gclk));
	jxor g1111(.dina(w_n806_0[1]),.dinb(w_n828_0[1]),.dout(n1413),.clk(gclk));
	jnot g1112(.din(w_n614_1[1]),.dout(n1414),.clk(gclk));
	jnot g1113(.din(w_n717_0[0]),.dout(n1415),.clk(gclk));
	jand g1114(.dina(w_n622_1[0]),.dinb(w_n828_0[0]),.dout(n1416),.clk(gclk));
	jand g1115(.dina(w_n628_0[0]),.dinb(w_G523_0[1]),.dout(n1417),.clk(gclk));
	jor g1116(.dina(n1417),.dinb(w_n829_0[0]),.dout(n1418),.clk(gclk));
	jor g1117(.dina(n1418),.dinb(n1416),.dout(n1419),.clk(gclk));
	jand g1118(.dina(n1419),.dinb(w_dff_B_76ZUcUfQ7_1),.dout(n1420),.clk(gclk));
	jxor g1119(.dina(w_n622_0[2]),.dinb(w_n618_0[1]),.dout(n1421),.clk(gclk));
	jnot g1120(.din(w_n1421_0[1]),.dout(n1422),.clk(gclk));
	jor g1121(.dina(w_dff_B_1KhJuAEY4_0),.dinb(n1420),.dout(n1423),.clk(gclk));
	jor g1122(.dina(w_n1421_0[0]),.dinb(w_n819_0[0]),.dout(n1424),.clk(gclk));
	jand g1123(.dina(n1424),.dinb(w_dff_B_OTErftW91_1),.dout(n1425),.clk(gclk));
	jxor g1124(.dina(w_n1425_0[1]),.dinb(w_dff_B_y49ND7CU4_1),.dout(n1426),.clk(gclk));
	jand g1125(.dina(n1426),.dinb(n1413),.dout(n1427),.clk(gclk));
	jnot g1126(.din(w_G2174_0[1]),.dout(n1428),.clk(gclk));
	jxor g1127(.dina(w_n806_0[0]),.dinb(w_n721_0[1]),.dout(n1429),.clk(gclk));
	jxor g1128(.dina(w_n1425_0[0]),.dinb(w_n614_1[0]),.dout(n1430),.clk(gclk));
	jand g1129(.dina(n1430),.dinb(n1429),.dout(n1431),.clk(gclk));
	jor g1130(.dina(n1431),.dinb(w_dff_B_nf95VBKY2_1),.dout(n1432),.clk(gclk));
	jor g1131(.dina(n1432),.dinb(w_dff_B_hmBEblHa7_1),.dout(n1433),.clk(gclk));
	jxor g1132(.dina(w_n729_0[1]),.dinb(w_n614_0[2]),.dout(n1434),.clk(gclk));
	jnot g1133(.din(w_n1434_0[1]),.dout(n1435),.clk(gclk));
	jor g1134(.dina(w_n622_0[1]),.dinb(w_n721_0[0]),.dout(n1436),.clk(gclk));
	jand g1135(.dina(n1436),.dinb(w_n723_0[0]),.dout(n1437),.clk(gclk));
	jxor g1136(.dina(w_dff_B_E8ELHlzE2_0),.dinb(w_n727_0[0]),.dout(n1438),.clk(gclk));
	jand g1137(.dina(w_n1438_0[1]),.dinb(n1435),.dout(n1439),.clk(gclk));
	jnot g1138(.din(w_n1438_0[0]),.dout(n1440),.clk(gclk));
	jand g1139(.dina(w_dff_B_kNcJBDK78_0),.dinb(w_n1434_0[0]),.dout(n1441),.clk(gclk));
	jor g1140(.dina(n1441),.dinb(w_G2174_0[0]),.dout(n1442),.clk(gclk));
	jor g1141(.dina(n1442),.dinb(n1439),.dout(n1443),.clk(gclk));
	jand g1142(.dina(w_dff_B_eVVXfIIu3_0),.dinb(n1433),.dout(n1444),.clk(gclk));
	jxor g1143(.dina(n1444),.dinb(w_n787_0[0]),.dout(n1445),.clk(gclk));
	jxor g1144(.dina(w_n1445_0[1]),.dinb(w_dff_B_tMFsKl7A6_1),.dout(n1446),.clk(gclk));
	jor g1145(.dina(w_n1446_0[1]),.dinb(w_n1410_0[1]),.dout(n1447),.clk(gclk));
	jxor g1146(.dina(w_n1445_0[0]),.dinb(w_n1411_0[0]),.dout(n1448),.clk(gclk));
	jor g1147(.dina(n1448),.dinb(w_n1409_0[0]),.dout(n1449),.clk(gclk));
	jand g1148(.dina(n1449),.dinb(w_G4091_1[1]),.dout(n1450),.clk(gclk));
	jand g1149(.dina(n1450),.dinb(w_n1447_0[1]),.dout(n1451),.clk(gclk));
	jor g1150(.dina(n1451),.dinb(w_dff_B_jqjgnu9Y6_1),.dout(n1452),.clk(gclk));
	jand g1151(.dina(w_n1452_0[1]),.dinb(w_dff_B_jxny4ArA6_1),.dout(w_dff_A_NFX8Ro7t6_2),.clk(gclk));
	jor g1152(.dina(w_G4091_1[0]),.dinb(G118),.dout(n1454),.clk(gclk));
	jand g1153(.dina(w_G251_2[2]),.dinb(w_n460_0[2]),.dout(n1455),.clk(gclk));
	jand g1154(.dina(w_G248_3[0]),.dinb(w_G234_1[0]),.dout(n1456),.clk(gclk));
	jor g1155(.dina(n1456),.dinb(w_n462_0[0]),.dout(n1457),.clk(gclk));
	jor g1156(.dina(n1457),.dinb(n1455),.dout(n1458),.clk(gclk));
	jand g1157(.dina(w_n366_2[2]),.dinb(w_n460_0[1]),.dout(n1459),.clk(gclk));
	jand g1158(.dina(w_n368_3[0]),.dinb(w_G234_0[2]),.dout(n1460),.clk(gclk));
	jor g1159(.dina(n1460),.dinb(w_G435_0[1]),.dout(n1461),.clk(gclk));
	jor g1160(.dina(n1461),.dinb(w_dff_B_XmZ1eiIF8_1),.dout(n1462),.clk(gclk));
	jand g1161(.dina(n1462),.dinb(w_dff_B_ts6ctaUK2_1),.dout(n1463),.clk(gclk));
	jor g1162(.dina(w_n402_1[1]),.dinb(w_G226_1[0]),.dout(n1464),.clk(gclk));
	jor g1163(.dina(w_n405_1[1]),.dinb(w_n530_0[2]),.dout(n1465),.clk(gclk));
	jand g1164(.dina(n1465),.dinb(w_G422_0[2]),.dout(n1466),.clk(gclk));
	jand g1165(.dina(n1466),.dinb(w_dff_B_Tu4nLu7q1_1),.dout(n1467),.clk(gclk));
	jor g1166(.dina(w_G254_1[0]),.dinb(w_G226_0[2]),.dout(n1468),.clk(gclk));
	jor g1167(.dina(w_G242_1[0]),.dinb(w_n530_0[1]),.dout(n1469),.clk(gclk));
	jand g1168(.dina(n1469),.dinb(w_n532_0[0]),.dout(n1470),.clk(gclk));
	jand g1169(.dina(n1470),.dinb(w_dff_B_A8uZyRAU6_1),.dout(n1471),.clk(gclk));
	jor g1170(.dina(n1471),.dinb(n1467),.dout(n1472),.clk(gclk));
	jxor g1171(.dina(n1472),.dinb(w_n528_0[0]),.dout(n1473),.clk(gclk));
	jor g1172(.dina(w_n402_1[0]),.dinb(w_G218_1[0]),.dout(n1474),.clk(gclk));
	jor g1173(.dina(w_n405_1[0]),.dinb(w_n507_0[2]),.dout(n1475),.clk(gclk));
	jand g1174(.dina(n1475),.dinb(w_G468_0[1]),.dout(n1476),.clk(gclk));
	jand g1175(.dina(n1476),.dinb(w_dff_B_QPKBkYa50_1),.dout(n1477),.clk(gclk));
	jor g1176(.dina(w_G254_0[2]),.dinb(w_G218_0[2]),.dout(n1478),.clk(gclk));
	jor g1177(.dina(w_G242_0[2]),.dinb(w_n507_0[1]),.dout(n1479),.clk(gclk));
	jand g1178(.dina(n1479),.dinb(w_n509_0[0]),.dout(n1480),.clk(gclk));
	jand g1179(.dina(n1480),.dinb(w_dff_B_kkKjk15J7_1),.dout(n1481),.clk(gclk));
	jor g1180(.dina(n1481),.dinb(n1477),.dout(n1482),.clk(gclk));
	jand g1181(.dina(w_G251_2[1]),.dinb(w_n541_0[2]),.dout(n1483),.clk(gclk));
	jand g1182(.dina(w_G248_2[2]),.dinb(w_G210_1[0]),.dout(n1484),.clk(gclk));
	jor g1183(.dina(n1484),.dinb(w_n543_0[0]),.dout(n1485),.clk(gclk));
	jor g1184(.dina(n1485),.dinb(n1483),.dout(n1486),.clk(gclk));
	jand g1185(.dina(w_n366_2[1]),.dinb(w_n541_0[1]),.dout(n1487),.clk(gclk));
	jand g1186(.dina(w_n368_2[2]),.dinb(w_G210_0[2]),.dout(n1488),.clk(gclk));
	jor g1187(.dina(n1488),.dinb(w_G457_0[2]),.dout(n1489),.clk(gclk));
	jor g1188(.dina(n1489),.dinb(w_dff_B_0aMwDOAT0_1),.dout(n1490),.clk(gclk));
	jand g1189(.dina(n1490),.dinb(w_dff_B_xxXRhAoH8_1),.dout(n1491),.clk(gclk));
	jxor g1190(.dina(n1491),.dinb(n1482),.dout(n1492),.clk(gclk));
	jxor g1191(.dina(n1492),.dinb(n1473),.dout(n1493),.clk(gclk));
	jxor g1192(.dina(n1493),.dinb(w_dff_B_TxKrL9ni2_1),.dout(n1494),.clk(gclk));
	jand g1193(.dina(w_n495_0[2]),.dinb(w_G251_2[0]),.dout(n1495),.clk(gclk));
	jand g1194(.dina(w_G281_1[0]),.dinb(w_G248_2[1]),.dout(n1496),.clk(gclk));
	jor g1195(.dina(n1496),.dinb(w_n497_0[1]),.dout(n1497),.clk(gclk));
	jor g1196(.dina(n1497),.dinb(n1495),.dout(n1498),.clk(gclk));
	jand g1197(.dina(w_n495_0[1]),.dinb(w_n366_2[0]),.dout(n1499),.clk(gclk));
	jand g1198(.dina(w_G281_0[2]),.dinb(w_n368_2[1]),.dout(n1500),.clk(gclk));
	jor g1199(.dina(n1500),.dinb(w_G374_0[0]),.dout(n1501),.clk(gclk));
	jor g1200(.dina(n1501),.dinb(w_dff_B_SAipD6aa6_1),.dout(n1502),.clk(gclk));
	jand g1201(.dina(n1502),.dinb(w_dff_B_GixM5bZd1_1),.dout(n1503),.clk(gclk));
	jand g1202(.dina(w_n449_0[2]),.dinb(w_G251_1[2]),.dout(n1504),.clk(gclk));
	jand g1203(.dina(w_G265_1[0]),.dinb(w_G248_2[0]),.dout(n1505),.clk(gclk));
	jor g1204(.dina(n1505),.dinb(w_n451_0[1]),.dout(n1506),.clk(gclk));
	jor g1205(.dina(n1506),.dinb(n1504),.dout(n1507),.clk(gclk));
	jand g1206(.dina(w_n449_0[1]),.dinb(w_n366_1[2]),.dout(n1508),.clk(gclk));
	jand g1207(.dina(w_G265_0[2]),.dinb(w_n368_2[0]),.dout(n1509),.clk(gclk));
	jor g1208(.dina(n1509),.dinb(w_G400_0[1]),.dout(n1510),.clk(gclk));
	jor g1209(.dina(n1510),.dinb(w_dff_B_NJxDURGC2_1),.dout(n1511),.clk(gclk));
	jand g1210(.dina(n1511),.dinb(w_dff_B_cCsAviXl1_1),.dout(n1512),.clk(gclk));
	jxor g1211(.dina(n1512),.dinb(n1503),.dout(n1513),.clk(gclk));
	jor g1212(.dina(w_G257_1[0]),.dinb(w_n402_0[2]),.dout(n1514),.clk(gclk));
	jor g1213(.dina(w_n471_0[2]),.dinb(w_n405_0[2]),.dout(n1515),.clk(gclk));
	jand g1214(.dina(n1515),.dinb(w_G389_0[0]),.dout(n1516),.clk(gclk));
	jand g1215(.dina(n1516),.dinb(w_dff_B_10meFRAC4_1),.dout(n1517),.clk(gclk));
	jor g1216(.dina(w_G257_0[2]),.dinb(w_G254_0[1]),.dout(n1518),.clk(gclk));
	jor g1217(.dina(w_n471_0[1]),.dinb(w_G242_0[1]),.dout(n1519),.clk(gclk));
	jand g1218(.dina(n1519),.dinb(w_n473_0[1]),.dout(n1520),.clk(gclk));
	jand g1219(.dina(n1520),.dinb(w_dff_B_OicV9Q9v5_1),.dout(n1521),.clk(gclk));
	jor g1220(.dina(n1521),.dinb(n1517),.dout(n1522),.clk(gclk));
	jand g1221(.dina(w_n484_0[2]),.dinb(w_G251_1[1]),.dout(n1523),.clk(gclk));
	jand g1222(.dina(w_G273_1[0]),.dinb(w_G248_1[2]),.dout(n1524),.clk(gclk));
	jor g1223(.dina(n1524),.dinb(w_n486_0[1]),.dout(n1525),.clk(gclk));
	jor g1224(.dina(n1525),.dinb(n1523),.dout(n1526),.clk(gclk));
	jand g1225(.dina(w_n484_0[1]),.dinb(w_n366_1[1]),.dout(n1527),.clk(gclk));
	jand g1226(.dina(w_G273_0[2]),.dinb(w_n368_1[2]),.dout(n1528),.clk(gclk));
	jor g1227(.dina(n1528),.dinb(w_G411_0[0]),.dout(n1529),.clk(gclk));
	jor g1228(.dina(n1529),.dinb(w_dff_B_wUIvTA2e6_1),.dout(n1530),.clk(gclk));
	jand g1229(.dina(n1530),.dinb(w_dff_B_ICVIfdOc7_1),.dout(n1531),.clk(gclk));
	jxor g1230(.dina(n1531),.dinb(n1522),.dout(n1532),.clk(gclk));
	jxor g1231(.dina(n1532),.dinb(n1513),.dout(n1533),.clk(gclk));
	jand g1232(.dina(w_n1533_0[1]),.dinb(w_n1494_0[1]),.dout(n1534),.clk(gclk));
	jnot g1233(.din(n1534),.dout(n1535),.clk(gclk));
	jor g1234(.dina(w_n1533_0[0]),.dinb(w_n1494_0[0]),.dout(n1536),.clk(gclk));
	jand g1235(.dina(n1536),.dinb(w_n750_0[2]),.dout(n1537),.clk(gclk));
	jand g1236(.dina(n1537),.dinb(n1535),.dout(n1538),.clk(gclk));
	jor g1237(.dina(n1454),.dinb(w_n746_0[1]),.dout(n1539),.clk(gclk));
	jor g1238(.dina(n1538),.dinb(w_G4092_1[0]),.dout(n1540),.clk(gclk));
	jxor g1239(.dina(w_n583_0[1]),.dinb(w_n578_0[0]),.dout(n1541),.clk(gclk));
	jxor g1240(.dina(n1541),.dinb(w_n943_0[0]),.dout(n1542),.clk(gclk));
	jnot g1241(.din(n1542),.dout(n1543),.clk(gclk));
	jand g1242(.dina(w_n587_0[2]),.dinb(w_G1497_0[2]),.dout(n1544),.clk(gclk));
	jor g1243(.dina(w_dff_B_j6uxmmWU0_0),.dinb(w_n696_0[0]),.dout(n1545),.clk(gclk));
	jnot g1244(.din(w_n1545_0[1]),.dout(n1546),.clk(gclk));
	jor g1245(.dina(w_n944_0[0]),.dinb(w_n930_0[1]),.dout(n1547),.clk(gclk));
	jand g1246(.dina(n1547),.dinb(w_n706_0[0]),.dout(n1548),.clk(gclk));
	jxor g1247(.dina(n1548),.dinb(w_n928_0[0]),.dout(n1549),.clk(gclk));
	jxor g1248(.dina(w_n605_1[1]),.dinb(w_n948_0[1]),.dout(n1550),.clk(gclk));
	jxor g1249(.dina(w_dff_B_rbzmz5CZ9_0),.dinb(n1549),.dout(n1551),.clk(gclk));
	jand g1250(.dina(w_dff_B_znBonFDJ3_0),.dinb(n1546),.dout(n1552),.clk(gclk));
	jxor g1251(.dina(w_n605_1[0]),.dinb(w_n703_0[0]),.dout(n1553),.clk(gclk));
	jand g1252(.dina(w_n605_0[2]),.dinb(w_n948_0[0]),.dout(n1554),.clk(gclk));
	jor g1253(.dina(n1554),.dinb(w_n702_0[0]),.dout(n1555),.clk(gclk));
	jnot g1254(.din(w_n1555_0[1]),.dout(n1556),.clk(gclk));
	jor g1255(.dina(n1556),.dinb(w_n930_0[0]),.dout(n1557),.clk(gclk));
	jor g1256(.dina(w_n1555_0[0]),.dinb(w_n707_0[0]),.dout(n1558),.clk(gclk));
	jand g1257(.dina(n1558),.dinb(w_dff_B_tJK6alD19_1),.dout(n1559),.clk(gclk));
	jxor g1258(.dina(n1559),.dinb(w_n596_0[0]),.dout(n1560),.clk(gclk));
	jand g1259(.dina(w_n1560_0[1]),.dinb(w_n1553_0[1]),.dout(n1561),.clk(gclk));
	jnot g1260(.din(n1561),.dout(n1562),.clk(gclk));
	jor g1261(.dina(w_n1560_0[0]),.dinb(w_n1553_0[0]),.dout(n1563),.clk(gclk));
	jand g1262(.dina(w_dff_B_bPw4S0de1_0),.dinb(w_n1545_0[0]),.dout(n1564),.clk(gclk));
	jand g1263(.dina(n1564),.dinb(w_dff_B_yPRmIuMF4_1),.dout(n1565),.clk(gclk));
	jor g1264(.dina(n1565),.dinb(n1552),.dout(n1566),.clk(gclk));
	jnot g1265(.din(w_G1497_0[1]),.dout(n1567),.clk(gclk));
	jand g1266(.dina(w_n682_0[0]),.dinb(w_n687_0[0]),.dout(n1568),.clk(gclk));
	jand g1267(.dina(w_n1568_0[1]),.dinb(w_n574_0[0]),.dout(n1569),.clk(gclk));
	jxor g1268(.dina(n1569),.dinb(w_n561_0[1]),.dout(n1570),.clk(gclk));
	jxor g1269(.dina(w_n572_0[1]),.dinb(w_n681_1[1]),.dout(n1571),.clk(gclk));
	jor g1270(.dina(w_n856_0[0]),.dinb(w_n853_0[0]),.dout(n1572),.clk(gclk));
	jand g1271(.dina(w_n693_0[1]),.dinb(w_n585_0[0]),.dout(n1573),.clk(gclk));
	jor g1272(.dina(n1573),.dinb(w_n855_0[0]),.dout(n1574),.clk(gclk));
	jand g1273(.dina(n1574),.dinb(n1572),.dout(n1575),.clk(gclk));
	jxor g1274(.dina(n1575),.dinb(w_dff_B_KctnXjBN9_1),.dout(n1576),.clk(gclk));
	jxor g1275(.dina(n1576),.dinb(w_dff_B_s14nKBMl3_1),.dout(n1577),.clk(gclk));
	jor g1276(.dina(n1577),.dinb(w_dff_B_KYhvU6y66_1),.dout(n1578),.clk(gclk));
	jxor g1277(.dina(w_n693_0[0]),.dinb(w_n572_0[0]),.dout(n1579),.clk(gclk));
	jor g1278(.dina(w_n857_0[0]),.dinb(w_n681_1[0]),.dout(n1580),.clk(gclk));
	jnot g1279(.din(w_n681_0[2]),.dout(n1581),.clk(gclk));
	jor g1280(.dina(w_n680_0[0]),.dinb(n1581),.dout(n1582),.clk(gclk));
	jor g1281(.dina(n1582),.dinb(w_n689_0[0]),.dout(n1583),.clk(gclk));
	jxor g1282(.dina(n1583),.dinb(w_n567_0[1]),.dout(n1584),.clk(gclk));
	jand g1283(.dina(w_dff_B_OZLQFGTU9_0),.dinb(n1580),.dout(n1585),.clk(gclk));
	jxor g1284(.dina(w_n1568_0[0]),.dinb(w_n561_0[0]),.dout(n1586),.clk(gclk));
	jxor g1285(.dina(w_dff_B_aWwzQuXm1_0),.dinb(n1585),.dout(n1587),.clk(gclk));
	jxor g1286(.dina(n1587),.dinb(w_dff_B_EtojTeXx9_1),.dout(n1588),.clk(gclk));
	jor g1287(.dina(n1588),.dinb(w_G1497_0[0]),.dout(n1589),.clk(gclk));
	jand g1288(.dina(w_dff_B_iCRNtnLO0_0),.dinb(n1578),.dout(n1590),.clk(gclk));
	jxor g1289(.dina(n1590),.dinb(n1566),.dout(n1591),.clk(gclk));
	jand g1290(.dina(w_n1591_0[1]),.dinb(w_n1543_0[1]),.dout(n1592),.clk(gclk));
	jnot g1291(.din(n1592),.dout(n1593),.clk(gclk));
	jor g1292(.dina(w_n1591_0[0]),.dinb(w_n1543_0[0]),.dout(n1594),.clk(gclk));
	jand g1293(.dina(n1594),.dinb(w_G4091_0[2]),.dout(n1595),.clk(gclk));
	jand g1294(.dina(n1595),.dinb(n1593),.dout(n1596),.clk(gclk));
	jor g1295(.dina(n1596),.dinb(w_dff_B_QcHQcyID4_1),.dout(n1597),.clk(gclk));
	jand g1296(.dina(w_n1597_0[1]),.dinb(w_dff_B_nIpOyoey8_1),.dout(w_dff_A_bDIpSuPb9_2),.clk(gclk));
	jand g1297(.dina(w_G4092_0[2]),.dinb(G97),.dout(n1599),.clk(gclk));
	jnot g1298(.din(n1599),.dout(n1600),.clk(gclk));
	jand g1299(.dina(w_dff_B_Yrygy9EL4_0),.dinb(w_n1597_0[0]),.dout(n1601),.clk(gclk));
	jnot g1300(.din(w_n1601_0[2]),.dout(n1602),.clk(gclk));
	jand g1301(.dina(w_n1602_0[1]),.dinb(w_n793_1[1]),.dout(n1603),.clk(gclk));
	jnot g1302(.din(w_n1447_0[0]),.dout(n1604),.clk(gclk));
	jand g1303(.dina(w_n1446_0[0]),.dinb(w_n1410_0[0]),.dout(n1605),.clk(gclk));
	jor g1304(.dina(n1605),.dinb(w_n750_0[1]),.dout(n1606),.clk(gclk));
	jor g1305(.dina(n1606),.dinb(n1604),.dout(n1607),.clk(gclk));
	jand g1306(.dina(n1607),.dinb(w_n1391_0[0]),.dout(n1608),.clk(gclk));
	jand g1307(.dina(w_G4092_0[1]),.dinb(G94),.dout(n1609),.clk(gclk));
	jor g1308(.dina(w_n1609_0[1]),.dinb(n1608),.dout(n1610),.clk(gclk));
	jand g1309(.dina(w_n1610_0[1]),.dinb(w_n797_1[1]),.dout(n1611),.clk(gclk));
	jand g1310(.dina(w_n799_1[1]),.dinb(w_G14_0[1]),.dout(n1612),.clk(gclk));
	jand g1311(.dina(w_n801_1[1]),.dinb(w_G64_0[1]),.dout(n1613),.clk(gclk));
	jor g1312(.dina(w_dff_B_h1ssQCLb9_0),.dinb(n1612),.dout(n1614),.clk(gclk));
	jor g1313(.dina(w_dff_B_4rHYBAdE5_0),.dinb(n1611),.dout(n1615),.clk(gclk));
	jor g1314(.dina(n1615),.dinb(n1603),.dout(w_dff_A_5NIX1Iv46_2),.clk(gclk));
	jand g1315(.dina(w_n1602_0[0]),.dinb(w_n840_1[1]),.dout(n1617),.clk(gclk));
	jand g1316(.dina(w_n1610_0[0]),.dinb(w_n843_1[1]),.dout(n1618),.clk(gclk));
	jand g1317(.dina(w_n845_1[1]),.dinb(w_G14_0[0]),.dout(n1619),.clk(gclk));
	jand g1318(.dina(w_n847_1[1]),.dinb(w_G64_0[0]),.dout(n1620),.clk(gclk));
	jor g1319(.dina(w_dff_B_RTVcvQFq5_0),.dinb(n1619),.dout(n1621),.clk(gclk));
	jor g1320(.dina(w_dff_B_8D5LGT767_0),.dinb(n1618),.dout(n1622),.clk(gclk));
	jor g1321(.dina(n1622),.dinb(n1617),.dout(w_dff_A_X47nM5mB6_2),.clk(gclk));
	jnot g1322(.din(w_G137_3[1]),.dout(n1624),.clk(gclk));
	jnot g1323(.din(w_n985_1[1]),.dout(n1625),.clk(gclk));
	jor g1324(.dina(w_n1601_0[1]),.dinb(w_dff_B_yj6s74DZ0_1),.dout(n1626),.clk(gclk));
	jnot g1325(.din(w_n988_1[1]),.dout(n1627),.clk(gclk));
	jnot g1326(.din(w_n1609_0[0]),.dout(n1628),.clk(gclk));
	jand g1327(.dina(w_dff_B_ndLxsYM54_0),.dinb(w_n1452_0[0]),.dout(n1629),.clk(gclk));
	jor g1328(.dina(w_n1629_0[1]),.dinb(w_dff_B_6DkHFI564_1),.dout(n1630),.clk(gclk));
	jnot g1329(.din(G179),.dout(n1631),.clk(gclk));
	jnot g1330(.din(w_n992_1[1]),.dout(n1632),.clk(gclk));
	jor g1331(.dina(n1632),.dinb(w_n1631_0[1]),.dout(n1633),.clk(gclk));
	jnot g1332(.din(G176),.dout(n1634),.clk(gclk));
	jnot g1333(.din(w_n990_1[1]),.dout(n1635),.clk(gclk));
	jor g1334(.dina(n1635),.dinb(w_n1634_0[1]),.dout(n1636),.clk(gclk));
	jand g1335(.dina(n1636),.dinb(w_dff_B_Y2zKwqgq8_1),.dout(n1637),.clk(gclk));
	jand g1336(.dina(w_dff_B_N3bhsw929_0),.dinb(n1630),.dout(n1638),.clk(gclk));
	jand g1337(.dina(n1638),.dinb(w_dff_B_NR8kUKjf6_1),.dout(n1639),.clk(gclk));
	jor g1338(.dina(n1639),.dinb(w_n1624_0[1]),.dout(G658),.clk(gclk));
	jnot g1339(.din(w_n999_1[1]),.dout(n1641),.clk(gclk));
	jor g1340(.dina(w_n1601_0[0]),.dinb(w_dff_B_pR7GSL0Y7_1),.dout(n1642),.clk(gclk));
	jnot g1341(.din(w_n1002_1[1]),.dout(n1643),.clk(gclk));
	jor g1342(.dina(w_n1629_0[0]),.dinb(w_dff_B_cRFX9r2w7_1),.dout(n1644),.clk(gclk));
	jnot g1343(.din(w_n1006_1[1]),.dout(n1645),.clk(gclk));
	jor g1344(.dina(n1645),.dinb(w_n1631_0[0]),.dout(n1646),.clk(gclk));
	jnot g1345(.din(w_n1004_1[1]),.dout(n1647),.clk(gclk));
	jor g1346(.dina(n1647),.dinb(w_n1634_0[0]),.dout(n1648),.clk(gclk));
	jand g1347(.dina(n1648),.dinb(w_dff_B_rptlmaIn4_1),.dout(n1649),.clk(gclk));
	jand g1348(.dina(w_dff_B_oAXzuI4Y3_0),.dinb(n1644),.dout(n1650),.clk(gclk));
	jand g1349(.dina(n1650),.dinb(w_dff_B_bUIEw9Ht9_1),.dout(n1651),.clk(gclk));
	jor g1350(.dina(n1651),.dinb(w_n1624_0[0]),.dout(G690),.clk(gclk));
	buf g1351(.din(w_G141_1[0]),.dout(w_dff_A_okV472fm6_1));
	buf g1352(.din(w_G293_0[0]),.dout(w_dff_A_NZDPOgPm2_1));
	buf g1353(.din(w_G3173_0[0]),.dout(w_dff_A_8SfPKRXf1_1));
	jnot g1354(.din(w_G545_0[1]),.dout(w_dff_A_kcOoDOTs8_1),.clk(gclk));
	jnot g1355(.din(w_G545_0[0]),.dout(w_dff_A_hDMD60wB6_1),.clk(gclk));
	buf g1356(.din(w_G137_3[0]),.dout(w_dff_A_01NRIr0n5_1));
	buf g1357(.din(w_G141_0[2]),.dout(w_dff_A_BnnZ8yRL2_1));
	buf g1358(.din(w_G1_2[0]),.dout(w_dff_A_Lh3AxbIW3_1));
	buf g1359(.din(w_G549_0[1]),.dout(w_dff_A_J5XkOm3N6_1));
	buf g1360(.din(w_G299_0[1]),.dout(w_dff_A_DyvXlmRo5_1));
	jnot g1361(.din(w_G549_0[0]),.dout(w_dff_A_nvgG7fE58_1),.clk(gclk));
	buf g1362(.din(w_G1_1[2]),.dout(w_dff_A_cVuHOXky3_1));
	buf g1363(.din(w_G1_1[1]),.dout(w_dff_A_iX0YGi3V0_1));
	buf g1364(.din(w_G1_1[0]),.dout(w_dff_A_FzCJlgsD0_1));
	buf g1365(.din(w_G1_0[2]),.dout(w_dff_A_PtVtnSx29_1));
	buf g1366(.din(w_G299_0[0]),.dout(w_dff_A_bcmCouej6_1));
	jor g1367(.dina(w_n336_0[0]),.dinb(w_n333_0[0]),.dout(w_dff_A_2Em61F4H5_2),.clk(gclk));
	jand g1368(.dina(w_n652_0[0]),.dinb(w_n633_0[1]),.dout(w_dff_A_Y2JNsu3g3_2),.clk(gclk));
	jand g1369(.dina(w_n607_0[0]),.dinb(w_n587_0[1]),.dout(w_dff_A_ILZVgwZy8_2),.clk(gclk));
	jor g1370(.dina(w_n709_0[0]),.dinb(w_n697_0[0]),.dout(w_dff_A_k90aNcvw2_2),.clk(gclk));
	jor g1371(.dina(w_n742_0[0]),.dinb(w_n733_0[0]),.dout(w_dff_A_zku3LX0f7_2),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_G1_0[0]),.doutb(w_G1_0[1]),.doutc(w_G1_0[2]),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_G1_1[0]),.doutb(w_G1_1[1]),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl jspl_w_G1_2(.douta(w_G1_2[0]),.doutb(w_G1_2[1]),.din(w_G1_0[1]));
	jspl3 jspl3_w_G4_0(.douta(w_G4_0[0]),.doutb(w_dff_A_9Gi1pbWn9_1),.doutc(w_G4_0[2]),.din(w_dff_B_K8ORnOKd0_3));
	jspl jspl_w_G4_1(.douta(w_dff_A_Xsi80K702_0),.doutb(w_G4_1[1]),.din(w_G4_0[0]));
	jspl jspl_w_G11_0(.douta(w_G11_0[0]),.doutb(w_G11_0[1]),.din(w_dff_B_LLUKbs4O8_2));
	jspl jspl_w_G14_0(.douta(w_G14_0[0]),.doutb(w_G14_0[1]),.din(w_dff_B_CaICsnEX1_2));
	jspl jspl_w_G17_0(.douta(w_G17_0[0]),.doutb(w_G17_0[1]),.din(w_dff_B_e6C6fCKi5_2));
	jspl jspl_w_G20_0(.douta(w_G20_0[0]),.doutb(w_G20_0[1]),.din(w_dff_B_u64XRs6s1_2));
	jspl jspl_w_G37_0(.douta(w_G37_0[0]),.doutb(w_G37_0[1]),.din(w_dff_B_IvRLvBDD0_2));
	jspl jspl_w_G40_0(.douta(w_G40_0[0]),.doutb(w_G40_0[1]),.din(w_dff_B_Mo8eHblO3_2));
	jspl jspl_w_G43_0(.douta(w_G43_0[0]),.doutb(w_G43_0[1]),.din(w_dff_B_aMcOYz5D7_2));
	jspl jspl_w_G46_0(.douta(w_G46_0[0]),.doutb(w_G46_0[1]),.din(w_dff_B_CWb2MDZp4_2));
	jspl jspl_w_G49_0(.douta(w_G49_0[0]),.doutb(w_G49_0[1]),.din(w_dff_B_VMkJNZAT8_2));
	jspl jspl_w_G54_0(.douta(w_dff_A_arY8dTIP6_0),.doutb(w_G54_0[1]),.din(G54));
	jspl jspl_w_G61_0(.douta(w_G61_0[0]),.doutb(w_G61_0[1]),.din(w_dff_B_nWHyNTeU4_2));
	jspl jspl_w_G64_0(.douta(w_G64_0[0]),.doutb(w_G64_0[1]),.din(w_dff_B_J9TBYGZH4_2));
	jspl jspl_w_G67_0(.douta(w_G67_0[0]),.doutb(w_G67_0[1]),.din(w_dff_B_PKSteptA6_2));
	jspl jspl_w_G70_0(.douta(w_G70_0[0]),.doutb(w_G70_0[1]),.din(w_dff_B_9xJiJbm46_2));
	jspl jspl_w_G73_0(.douta(w_G73_0[0]),.doutb(w_G73_0[1]),.din(w_dff_B_cUq7hYYo7_2));
	jspl jspl_w_G76_0(.douta(w_G76_0[0]),.doutb(w_G76_0[1]),.din(w_dff_B_XzoOlpDi0_2));
	jspl jspl_w_G91_0(.douta(w_G91_0[0]),.doutb(w_G91_0[1]),.din(w_dff_B_el6Qlaq36_2));
	jspl jspl_w_G100_0(.douta(w_G100_0[0]),.doutb(w_G100_0[1]),.din(w_dff_B_dCjbwhYg7_2));
	jspl jspl_w_G103_0(.douta(w_G103_0[0]),.doutb(w_G103_0[1]),.din(w_dff_B_XnPH5e6I5_2));
	jspl jspl_w_G106_0(.douta(w_G106_0[0]),.doutb(w_G106_0[1]),.din(w_dff_B_VJUTrNHT7_2));
	jspl jspl_w_G109_0(.douta(w_G109_0[0]),.doutb(w_G109_0[1]),.din(w_dff_B_LlnZ7Dqk4_2));
	jspl jspl_w_G123_0(.douta(w_dff_A_knKS0aNM9_0),.doutb(w_G123_0[1]),.din(w_dff_B_YztjzzMN1_2));
	jspl jspl_w_G132_0(.douta(w_dff_A_1gwjD4y12_0),.doutb(w_G132_0[1]),.din(w_dff_B_EIYVk1i47_2));
	jspl3 jspl3_w_G137_0(.douta(w_dff_A_y8EKslp71_0),.doutb(w_dff_A_7BUQRPrB0_1),.doutc(w_G137_0[2]),.din(G137));
	jspl3 jspl3_w_G137_1(.douta(w_dff_A_bi3X8rNv0_0),.doutb(w_dff_A_ooNgcASa8_1),.doutc(w_G137_1[2]),.din(w_G137_0[0]));
	jspl3 jspl3_w_G137_2(.douta(w_dff_A_lp1paIgS1_0),.doutb(w_dff_A_HWQavakt8_1),.doutc(w_G137_2[2]),.din(w_G137_0[1]));
	jspl3 jspl3_w_G137_3(.douta(w_G137_3[0]),.doutb(w_G137_3[1]),.doutc(w_dff_A_QGAAvwDb4_2),.din(w_G137_0[2]));
	jspl3 jspl3_w_G137_4(.douta(w_dff_A_eo9C9SN44_0),.doutb(w_dff_A_nd61yT9j0_1),.doutc(w_G137_4[2]),.din(w_G137_1[0]));
	jspl3 jspl3_w_G137_5(.douta(w_dff_A_a3Hw78NH0_0),.doutb(w_G137_5[1]),.doutc(w_G137_5[2]),.din(w_G137_1[1]));
	jspl3 jspl3_w_G137_6(.douta(w_dff_A_hwg82l3u4_0),.doutb(w_dff_A_6cW6CQ4E5_1),.doutc(w_G137_6[2]),.din(w_G137_1[2]));
	jspl3 jspl3_w_G137_7(.douta(w_G137_7[0]),.doutb(w_dff_A_JJMcdgTq7_1),.doutc(w_dff_A_3Z2ePtAG1_2),.din(w_G137_2[0]));
	jspl3 jspl3_w_G137_8(.douta(w_dff_A_tpjrM7qL1_0),.doutb(w_G137_8[1]),.doutc(w_dff_A_73R8StKX9_2),.din(w_G137_2[1]));
	jspl jspl_w_G137_9(.douta(w_G137_9[0]),.doutb(w_G137_9[1]),.din(w_G137_2[2]));
	jspl3 jspl3_w_G141_0(.douta(w_G141_0[0]),.doutb(w_G141_0[1]),.doutc(w_G141_0[2]),.din(G141));
	jspl3 jspl3_w_G141_1(.douta(w_G141_1[0]),.doutb(w_dff_A_FVxwN3J96_1),.doutc(w_dff_A_JcqojU074_2),.din(w_G141_0[0]));
	jspl3 jspl3_w_G141_2(.douta(w_dff_A_IMIxIDym3_0),.doutb(w_dff_A_Uix9emZd8_1),.doutc(w_G141_2[2]),.din(w_G141_0[1]));
	jspl jspl_w_G146_0(.douta(w_G146_0[0]),.doutb(w_G146_0[1]),.din(w_dff_B_p5VKIVOZ9_2));
	jspl jspl_w_G149_0(.douta(w_G149_0[0]),.doutb(w_G149_0[1]),.din(w_dff_B_VdpNh2Zg3_2));
	jspl jspl_w_G152_0(.douta(w_G152_0[0]),.doutb(w_G152_0[1]),.din(w_dff_B_nJEeufId6_2));
	jspl jspl_w_G155_0(.douta(w_G155_0[0]),.doutb(w_G155_0[1]),.din(w_dff_B_Hr5Ef1GE8_2));
	jspl jspl_w_G158_0(.douta(w_G158_0[0]),.doutb(w_G158_0[1]),.din(w_dff_B_Xx8Rvxsi8_2));
	jspl jspl_w_G161_0(.douta(w_G161_0[0]),.doutb(w_G161_0[1]),.din(w_dff_B_FiyemRXA2_2));
	jspl jspl_w_G164_0(.douta(w_G164_0[0]),.doutb(w_G164_0[1]),.din(w_dff_B_8Rzw76ML0_2));
	jspl jspl_w_G167_0(.douta(w_G167_0[0]),.doutb(w_G167_0[1]),.din(w_dff_B_HwkqESHD8_2));
	jspl jspl_w_G170_0(.douta(w_G170_0[0]),.doutb(w_G170_0[1]),.din(w_dff_B_K0FZ46m73_2));
	jspl jspl_w_G173_0(.douta(w_G173_0[0]),.doutb(w_G173_0[1]),.din(w_dff_B_SurJZRrC4_2));
	jspl jspl_w_G182_0(.douta(w_G182_0[0]),.doutb(w_G182_0[1]),.din(w_dff_B_qds7jQhf3_2));
	jspl jspl_w_G185_0(.douta(w_G185_0[0]),.doutb(w_G185_0[1]),.din(w_dff_B_EftrGcDC3_2));
	jspl jspl_w_G188_0(.douta(w_G188_0[0]),.doutb(w_G188_0[1]),.din(w_dff_B_AmPL2t1L6_2));
	jspl jspl_w_G191_0(.douta(w_G191_0[0]),.doutb(w_G191_0[1]),.din(w_dff_B_PNYWUf4z8_2));
	jspl jspl_w_G194_0(.douta(w_G194_0[0]),.doutb(w_G194_0[1]),.din(w_dff_B_kg6O6kvQ3_2));
	jspl jspl_w_G197_0(.douta(w_G197_0[0]),.doutb(w_G197_0[1]),.din(w_dff_B_xpzfz9bn8_2));
	jspl jspl_w_G200_0(.douta(w_G200_0[0]),.doutb(w_G200_0[1]),.din(w_dff_B_twHeLHGu2_2));
	jspl jspl_w_G203_0(.douta(w_G203_0[0]),.doutb(w_G203_0[1]),.din(w_dff_B_hcqlBw8G8_2));
	jspl3 jspl3_w_G206_0(.douta(w_dff_A_eMdGojBb4_0),.doutb(w_G206_0[1]),.doutc(w_G206_0[2]),.din(G206));
	jspl3 jspl3_w_G210_0(.douta(w_G210_0[0]),.doutb(w_G210_0[1]),.doutc(w_dff_A_BgefP6GH8_2),.din(G210));
	jspl3 jspl3_w_G210_1(.douta(w_G210_1[0]),.doutb(w_dff_A_IV5zb80V7_1),.doutc(w_G210_1[2]),.din(w_G210_0[0]));
	jspl3 jspl3_w_G210_2(.douta(w_G210_2[0]),.doutb(w_dff_A_0Pys0NPO7_1),.doutc(w_G210_2[2]),.din(w_G210_0[1]));
	jspl3 jspl3_w_G218_0(.douta(w_G218_0[0]),.doutb(w_G218_0[1]),.doutc(w_G218_0[2]),.din(G218));
	jspl3 jspl3_w_G218_1(.douta(w_dff_A_nXUQGQHM8_0),.doutb(w_G218_1[1]),.doutc(w_G218_1[2]),.din(w_G218_0[0]));
	jspl3 jspl3_w_G218_2(.douta(w_G218_2[0]),.doutb(w_dff_A_dhGTwRnI9_1),.doutc(w_G218_2[2]),.din(w_G218_0[1]));
	jspl3 jspl3_w_G226_0(.douta(w_G226_0[0]),.doutb(w_G226_0[1]),.doutc(w_G226_0[2]),.din(G226));
	jspl3 jspl3_w_G226_1(.douta(w_dff_A_OpqiR3Vc2_0),.doutb(w_G226_1[1]),.doutc(w_G226_1[2]),.din(w_G226_0[0]));
	jspl3 jspl3_w_G226_2(.douta(w_G226_2[0]),.doutb(w_dff_A_kG5zjPzZ4_1),.doutc(w_G226_2[2]),.din(w_G226_0[1]));
	jspl3 jspl3_w_G234_0(.douta(w_G234_0[0]),.doutb(w_G234_0[1]),.doutc(w_dff_A_q9w38W3Z5_2),.din(G234));
	jspl3 jspl3_w_G234_1(.douta(w_G234_1[0]),.doutb(w_G234_1[1]),.doutc(w_G234_1[2]),.din(w_G234_0[0]));
	jspl jspl_w_G234_2(.douta(w_dff_A_s2t4eMkx3_0),.doutb(w_G234_2[1]),.din(w_G234_0[1]));
	jspl3 jspl3_w_G242_0(.douta(w_G242_0[0]),.doutb(w_dff_A_NOh48NUa9_1),.doutc(w_dff_A_o2DKDKw12_2),.din(G242));
	jspl3 jspl3_w_G242_1(.douta(w_dff_A_1cbmMLvm9_0),.doutb(w_dff_A_iYvooa9B2_1),.doutc(w_G242_1[2]),.din(w_G242_0[0]));
	jspl jspl_w_G245_0(.douta(w_G245_0[0]),.doutb(w_G245_0[1]),.din(G245));
	jspl3 jspl3_w_G248_0(.douta(w_G248_0[0]),.doutb(w_G248_0[1]),.doutc(w_G248_0[2]),.din(G248));
	jspl3 jspl3_w_G248_1(.douta(w_G248_1[0]),.doutb(w_G248_1[1]),.doutc(w_G248_1[2]),.din(w_G248_0[0]));
	jspl3 jspl3_w_G248_2(.douta(w_G248_2[0]),.doutb(w_G248_2[1]),.doutc(w_G248_2[2]),.din(w_G248_0[1]));
	jspl3 jspl3_w_G248_3(.douta(w_G248_3[0]),.doutb(w_G248_3[1]),.doutc(w_dff_A_i7B6QyWf9_2),.din(w_G248_0[2]));
	jspl3 jspl3_w_G248_4(.douta(w_G248_4[0]),.doutb(w_G248_4[1]),.doutc(w_G248_4[2]),.din(w_G248_1[0]));
	jspl jspl_w_G248_5(.douta(w_G248_5[0]),.doutb(w_G248_5[1]),.din(w_G248_1[1]));
	jspl3 jspl3_w_G251_0(.douta(w_G251_0[0]),.doutb(w_dff_A_qJLIzwhg0_1),.doutc(w_dff_A_w4RxTup30_2),.din(G251));
	jspl3 jspl3_w_G251_1(.douta(w_G251_1[0]),.doutb(w_dff_A_FE7aTk4H4_1),.doutc(w_dff_A_5yJTXELi2_2),.din(w_G251_0[0]));
	jspl3 jspl3_w_G251_2(.douta(w_G251_2[0]),.doutb(w_G251_2[1]),.doutc(w_G251_2[2]),.din(w_G251_0[1]));
	jspl3 jspl3_w_G251_3(.douta(w_G251_3[0]),.doutb(w_G251_3[1]),.doutc(w_G251_3[2]),.din(w_G251_0[2]));
	jspl3 jspl3_w_G251_4(.douta(w_G251_4[0]),.doutb(w_dff_A_OUwJ3ss06_1),.doutc(w_dff_A_JLvkYXd86_2),.din(w_G251_1[0]));
	jspl3 jspl3_w_G254_0(.douta(w_G254_0[0]),.doutb(w_G254_0[1]),.doutc(w_G254_0[2]),.din(G254));
	jspl3 jspl3_w_G254_1(.douta(w_G254_1[0]),.doutb(w_G254_1[1]),.doutc(w_G254_1[2]),.din(w_G254_0[0]));
	jspl3 jspl3_w_G257_0(.douta(w_G257_0[0]),.doutb(w_G257_0[1]),.doutc(w_G257_0[2]),.din(G257));
	jspl3 jspl3_w_G257_1(.douta(w_dff_A_bANAr1uV7_0),.doutb(w_G257_1[1]),.doutc(w_G257_1[2]),.din(w_G257_0[0]));
	jspl3 jspl3_w_G257_2(.douta(w_G257_2[0]),.doutb(w_dff_A_xKkvtONz0_1),.doutc(w_G257_2[2]),.din(w_G257_0[1]));
	jspl3 jspl3_w_G265_0(.douta(w_G265_0[0]),.doutb(w_G265_0[1]),.doutc(w_dff_A_CWikI4PP6_2),.din(G265));
	jspl3 jspl3_w_G265_1(.douta(w_G265_1[0]),.doutb(w_G265_1[1]),.doutc(w_G265_1[2]),.din(w_G265_0[0]));
	jspl jspl_w_G265_2(.douta(w_dff_A_a10Qzhlk4_0),.doutb(w_G265_2[1]),.din(w_G265_0[1]));
	jspl3 jspl3_w_G273_0(.douta(w_G273_0[0]),.doutb(w_G273_0[1]),.doutc(w_dff_A_NUBUx68D1_2),.din(G273));
	jspl3 jspl3_w_G273_1(.douta(w_G273_1[0]),.doutb(w_G273_1[1]),.doutc(w_G273_1[2]),.din(w_G273_0[0]));
	jspl3 jspl3_w_G273_2(.douta(w_G273_2[0]),.doutb(w_dff_A_CgprWX050_1),.doutc(w_G273_2[2]),.din(w_G273_0[1]));
	jspl jspl_w_G280_0(.douta(w_G280_0[0]),.doutb(w_dff_A_o9qhUCMZ1_1),.din(G280));
	jspl3 jspl3_w_G281_0(.douta(w_G281_0[0]),.doutb(w_G281_0[1]),.doutc(w_dff_A_3ZfCYEqE6_2),.din(G281));
	jspl3 jspl3_w_G281_1(.douta(w_G281_1[0]),.doutb(w_G281_1[1]),.doutc(w_G281_1[2]),.din(w_G281_0[0]));
	jspl jspl_w_G281_2(.douta(w_dff_A_AAuUKy352_0),.doutb(w_G281_2[1]),.din(w_G281_0[1]));
	jspl jspl_w_G289_0(.douta(w_dff_A_X2w1lQ6U1_0),.doutb(w_G289_0[1]),.din(G289));
	jspl3 jspl3_w_G293_0(.douta(w_G293_0[0]),.doutb(w_dff_A_ClLpTeIE1_1),.doutc(w_G293_0[2]),.din(G293));
	jspl3 jspl3_w_G299_0(.douta(w_G299_0[0]),.doutb(w_G299_0[1]),.doutc(w_G299_0[2]),.din(G299));
	jspl3 jspl3_w_G302_0(.douta(w_dff_A_FTOzRZ710_0),.doutb(w_dff_A_5EZWNJ094_1),.doutc(w_G302_0[2]),.din(G302));
	jspl3 jspl3_w_G308_0(.douta(w_G308_0[0]),.doutb(w_G308_0[1]),.doutc(w_G308_0[2]),.din(G308));
	jspl3 jspl3_w_G308_1(.douta(w_dff_A_Z06Ba6Xd8_0),.doutb(w_G308_1[1]),.doutc(w_G308_1[2]),.din(w_G308_0[0]));
	jspl3 jspl3_w_G316_0(.douta(w_G316_0[0]),.doutb(w_G316_0[1]),.doutc(w_G316_0[2]),.din(G316));
	jspl3 jspl3_w_G316_1(.douta(w_dff_A_WRca75ot1_0),.doutb(w_G316_1[1]),.doutc(w_G316_1[2]),.din(w_G316_0[0]));
	jspl3 jspl3_w_G324_0(.douta(w_G324_0[0]),.doutb(w_dff_A_X2o6mQP26_1),.doutc(w_G324_0[2]),.din(G324));
	jspl3 jspl3_w_G324_1(.douta(w_G324_1[0]),.doutb(w_dff_A_f2Bes9Bs9_1),.doutc(w_G324_1[2]),.din(w_G324_0[0]));
	jspl jspl_w_G331_0(.douta(w_G331_0[0]),.doutb(w_dff_A_AvITlxYr9_1),.din(G331));
	jspl3 jspl3_w_G332_0(.douta(w_G332_0[0]),.doutb(w_G332_0[1]),.doutc(w_G332_0[2]),.din(G332));
	jspl3 jspl3_w_G332_1(.douta(w_G332_1[0]),.doutb(w_G332_1[1]),.doutc(w_dff_A_XlcVMFwu1_2),.din(w_G332_0[0]));
	jspl3 jspl3_w_G332_2(.douta(w_dff_A_SjAokIeW6_0),.doutb(w_G332_2[1]),.doutc(w_G332_2[2]),.din(w_G332_0[1]));
	jspl3 jspl3_w_G332_3(.douta(w_dff_A_CrsoojyL3_0),.doutb(w_G332_3[1]),.doutc(w_dff_A_iDRi8Z7q6_2),.din(w_G332_0[2]));
	jspl3 jspl3_w_G332_4(.douta(w_dff_A_EeOoDiHL9_0),.doutb(w_G332_4[1]),.doutc(w_G332_4[2]),.din(w_G332_1[0]));
	jspl3 jspl3_w_G335_0(.douta(w_G335_0[0]),.doutb(w_G335_0[1]),.doutc(w_G335_0[2]),.din(G335));
	jspl3 jspl3_w_G335_1(.douta(w_G335_1[0]),.doutb(w_G335_1[1]),.doutc(w_dff_A_z285s69A9_2),.din(w_G335_0[0]));
	jspl3 jspl3_w_G335_2(.douta(w_G335_2[0]),.doutb(w_G335_2[1]),.doutc(w_G335_2[2]),.din(w_G335_0[1]));
	jspl3 jspl3_w_G335_3(.douta(w_dff_A_D4JVfPTQ7_0),.doutb(w_G335_3[1]),.doutc(w_G335_3[2]),.din(w_G335_0[2]));
	jspl jspl_w_G335_4(.douta(w_dff_A_dINxCVap4_0),.doutb(w_G335_4[1]),.din(w_G335_1[0]));
	jspl3 jspl3_w_G341_0(.douta(w_G341_0[0]),.doutb(w_G341_0[1]),.doutc(w_dff_A_YiyeAhCF0_2),.din(G341));
	jspl3 jspl3_w_G341_1(.douta(w_G341_1[0]),.doutb(w_G341_1[1]),.doutc(w_G341_1[2]),.din(w_G341_0[0]));
	jspl3 jspl3_w_G341_2(.douta(w_G341_2[0]),.doutb(w_dff_A_YGYkLDhj5_1),.doutc(w_G341_2[2]),.din(w_G341_0[1]));
	jspl jspl_w_G348_0(.douta(w_dff_A_F1MW2BrB7_0),.doutb(w_G348_0[1]),.din(G348));
	jspl3 jspl3_w_G351_0(.douta(w_G351_0[0]),.doutb(w_G351_0[1]),.doutc(w_G351_0[2]),.din(G351));
	jspl3 jspl3_w_G351_1(.douta(w_dff_A_hXqnvGe07_0),.doutb(w_G351_1[1]),.doutc(w_G351_1[2]),.din(w_G351_0[0]));
	jspl3 jspl3_w_G351_2(.douta(w_G351_2[0]),.doutb(w_dff_A_HY2aFV2P3_1),.doutc(w_G351_2[2]),.din(w_G351_0[1]));
	jspl jspl_w_G358_0(.douta(w_dff_A_EcPFPxEC7_0),.doutb(w_G358_0[1]),.din(G358));
	jspl3 jspl3_w_G361_0(.douta(w_G361_0[0]),.doutb(w_dff_A_2gyqCwep7_1),.doutc(w_G361_0[2]),.din(G361));
	jspl jspl_w_G369_0(.douta(w_dff_A_5m1sBFBP3_0),.doutb(w_G369_0[1]),.din(G369));
	jspl3 jspl3_w_G374_0(.douta(w_dff_A_EA789TRI2_0),.doutb(w_dff_A_iAcg0cnm8_1),.doutc(w_G374_0[2]),.din(G374));
	jspl3 jspl3_w_G389_0(.douta(w_dff_A_deWhamyq0_0),.doutb(w_dff_A_bdsLIN204_1),.doutc(w_G389_0[2]),.din(G389));
	jspl3 jspl3_w_G400_0(.douta(w_G400_0[0]),.doutb(w_dff_A_9GNBrGGm0_1),.doutc(w_dff_A_cF42Pl3q4_2),.din(G400));
	jspl jspl_w_G400_1(.douta(w_dff_A_MVwIv0GP9_0),.doutb(w_G400_1[1]),.din(w_G400_0[0]));
	jspl3 jspl3_w_G411_0(.douta(w_dff_A_lp8KMlFN7_0),.doutb(w_dff_A_jOqVUj9t0_1),.doutc(w_G411_0[2]),.din(G411));
	jspl3 jspl3_w_G422_0(.douta(w_dff_A_J4a6OJl35_0),.doutb(w_G422_0[1]),.doutc(w_dff_A_LuvEiM885_2),.din(G422));
	jspl3 jspl3_w_G422_1(.douta(w_G422_1[0]),.doutb(w_G422_1[1]),.doutc(w_G422_1[2]),.din(w_G422_0[0]));
	jspl jspl_w_G422_2(.douta(w_dff_A_yRJKABJA7_0),.doutb(w_G422_2[1]),.din(w_G422_0[1]));
	jspl3 jspl3_w_G435_0(.douta(w_G435_0[0]),.doutb(w_dff_A_8bvJuRvx0_1),.doutc(w_dff_A_tGhJKCd82_2),.din(G435));
	jspl3 jspl3_w_G435_1(.douta(w_dff_A_veECLmaf3_0),.doutb(w_dff_A_SBOE7Fke9_1),.doutc(w_G435_1[2]),.din(w_G435_0[0]));
	jspl3 jspl3_w_G446_0(.douta(w_G446_0[0]),.doutb(w_dff_A_89vNui0Q7_1),.doutc(w_dff_A_I0myafGa7_2),.din(G446));
	jspl3 jspl3_w_G446_1(.douta(w_dff_A_bbab6R4y3_0),.doutb(w_dff_A_hEVKOsBS8_1),.doutc(w_G446_1[2]),.din(w_G446_0[0]));
	jspl3 jspl3_w_G457_0(.douta(w_dff_A_Jut5NXeM6_0),.doutb(w_G457_0[1]),.doutc(w_dff_A_xZYFZW7P3_2),.din(G457));
	jspl3 jspl3_w_G457_1(.douta(w_G457_1[0]),.doutb(w_G457_1[1]),.doutc(w_G457_1[2]),.din(w_G457_0[0]));
	jspl jspl_w_G457_2(.douta(w_dff_A_73sXI6kO5_0),.doutb(w_G457_2[1]),.din(w_G457_0[1]));
	jspl3 jspl3_w_G468_0(.douta(w_G468_0[0]),.doutb(w_dff_A_2Rm7Aary5_1),.doutc(w_dff_A_YXV3NzWV7_2),.din(G468));
	jspl3 jspl3_w_G468_1(.douta(w_dff_A_3uU7QwdY8_0),.doutb(w_dff_A_UkQVmX7O7_1),.doutc(w_G468_1[2]),.din(w_G468_0[0]));
	jspl3 jspl3_w_G479_0(.douta(w_G479_0[0]),.doutb(w_dff_A_wvmDIRuM7_1),.doutc(w_dff_A_YYBiyCFM4_2),.din(G479));
	jspl jspl_w_G479_1(.douta(w_dff_A_38xu0fvJ7_0),.doutb(w_G479_1[1]),.din(w_G479_0[0]));
	jspl3 jspl3_w_G490_0(.douta(w_G490_0[0]),.doutb(w_dff_A_wQ07uUHs9_1),.doutc(w_dff_A_OJtfwC613_2),.din(G490));
	jspl3 jspl3_w_G490_1(.douta(w_dff_A_XRPK02d44_0),.doutb(w_dff_A_nzThzmNM3_1),.doutc(w_G490_1[2]),.din(w_G490_0[0]));
	jspl3 jspl3_w_G503_0(.douta(w_G503_0[0]),.doutb(w_dff_A_84OCqbd11_1),.doutc(w_dff_A_HyLyg6kX7_2),.din(G503));
	jspl3 jspl3_w_G503_1(.douta(w_dff_A_FFQSG4AZ9_0),.doutb(w_dff_A_R2qompgH1_1),.doutc(w_G503_1[2]),.din(w_G503_0[0]));
	jspl3 jspl3_w_G514_0(.douta(w_G514_0[0]),.doutb(w_dff_A_tg6NZPpn6_1),.doutc(w_dff_A_Z4IRXIZx4_2),.din(G514));
	jspl jspl_w_G514_1(.douta(w_G514_1[0]),.doutb(w_G514_1[1]),.din(w_G514_0[0]));
	jspl3 jspl3_w_G523_0(.douta(w_G523_0[0]),.doutb(w_dff_A_Jk1aUJmI7_1),.doutc(w_dff_A_7dGOx6od9_2),.din(G523));
	jspl jspl_w_G523_1(.douta(w_dff_A_7maiGc5N3_0),.doutb(w_G523_1[1]),.din(w_G523_0[0]));
	jspl3 jspl3_w_G534_0(.douta(w_G534_0[0]),.doutb(w_dff_A_vd4oStN78_1),.doutc(w_dff_A_ogSajMlJ4_2),.din(G534));
	jspl3 jspl3_w_G534_1(.douta(w_dff_A_FFhWWLlg1_0),.doutb(w_dff_A_DX0O2Syd8_1),.doutc(w_G534_1[2]),.din(w_G534_0[0]));
	jspl3 jspl3_w_G545_0(.douta(w_G545_0[0]),.doutb(w_G545_0[1]),.doutc(w_G545_0[2]),.din(G545));
	jspl3 jspl3_w_G549_0(.douta(w_G549_0[0]),.doutb(w_G549_0[1]),.doutc(w_G549_0[2]),.din(G549));
	jspl jspl_w_G552_0(.douta(w_G552_0[0]),.doutb(w_G552_0[1]),.din(G552));
	jspl jspl_w_G559_0(.douta(w_G559_0[0]),.doutb(w_G559_0[1]),.din(G559));
	jspl jspl_w_G562_0(.douta(w_G562_0[0]),.doutb(w_G562_0[1]),.din(G562));
	jspl3 jspl3_w_G1497_0(.douta(w_dff_A_YEIBHXyR5_0),.doutb(w_G1497_0[1]),.doutc(w_dff_A_dHQDRExs4_2),.din(G1497));
	jspl3 jspl3_w_G1689_0(.douta(w_G1689_0[0]),.doutb(w_G1689_0[1]),.doutc(w_dff_A_4K5utaxy6_2),.din(G1689));
	jspl3 jspl3_w_G1690_0(.douta(w_G1690_0[0]),.doutb(w_dff_A_hAuu7uOo4_1),.doutc(w_G1690_0[2]),.din(G1690));
	jspl3 jspl3_w_G1691_0(.douta(w_G1691_0[0]),.doutb(w_G1691_0[1]),.doutc(w_dff_A_zWSyWcJh3_2),.din(G1691));
	jspl3 jspl3_w_G1694_0(.douta(w_G1694_0[0]),.doutb(w_dff_A_IaEcCyU10_1),.doutc(w_G1694_0[2]),.din(G1694));
	jspl3 jspl3_w_G2174_0(.douta(w_dff_A_Z08EWguM7_0),.doutb(w_G2174_0[1]),.doutc(w_dff_A_5KgIyjV38_2),.din(G2174));
	jspl3 jspl3_w_G2358_0(.douta(w_G2358_0[0]),.doutb(w_G2358_0[1]),.doutc(w_G2358_0[2]),.din(G2358));
	jspl3 jspl3_w_G2358_1(.douta(w_G2358_1[0]),.doutb(w_G2358_1[1]),.doutc(w_G2358_1[2]),.din(w_G2358_0[0]));
	jspl3 jspl3_w_G2358_2(.douta(w_dff_A_5EOTA0Rs8_0),.doutb(w_dff_A_BkHOyTil1_1),.doutc(w_G2358_2[2]),.din(w_G2358_0[1]));
	jspl jspl_w_G3173_0(.douta(w_G3173_0[0]),.doutb(w_G3173_0[1]),.din(G3173));
	jspl3 jspl3_w_G3546_0(.douta(w_G3546_0[0]),.doutb(w_G3546_0[1]),.doutc(w_G3546_0[2]),.din(G3546));
	jspl3 jspl3_w_G3546_1(.douta(w_G3546_1[0]),.doutb(w_G3546_1[1]),.doutc(w_G3546_1[2]),.din(w_G3546_0[0]));
	jspl3 jspl3_w_G3546_2(.douta(w_G3546_2[0]),.doutb(w_G3546_2[1]),.doutc(w_G3546_2[2]),.din(w_G3546_0[1]));
	jspl3 jspl3_w_G3546_3(.douta(w_G3546_3[0]),.doutb(w_G3546_3[1]),.doutc(w_G3546_3[2]),.din(w_G3546_0[2]));
	jspl3 jspl3_w_G3546_4(.douta(w_G3546_4[0]),.doutb(w_G3546_4[1]),.doutc(w_G3546_4[2]),.din(w_G3546_1[0]));
	jspl jspl_w_G3546_5(.douta(w_G3546_5[0]),.doutb(w_G3546_5[1]),.din(w_G3546_1[1]));
	jspl3 jspl3_w_G3548_0(.douta(w_G3548_0[0]),.doutb(w_G3548_0[1]),.doutc(w_G3548_0[2]),.din(w_dff_B_r7DXClUe9_3));
	jspl3 jspl3_w_G3548_1(.douta(w_G3548_1[0]),.doutb(w_G3548_1[1]),.doutc(w_G3548_1[2]),.din(w_G3548_0[0]));
	jspl3 jspl3_w_G3548_2(.douta(w_G3548_2[0]),.doutb(w_G3548_2[1]),.doutc(w_G3548_2[2]),.din(w_G3548_0[1]));
	jspl3 jspl3_w_G3548_3(.douta(w_G3548_3[0]),.doutb(w_G3548_3[1]),.doutc(w_G3548_3[2]),.din(w_G3548_0[2]));
	jspl3 jspl3_w_G3548_4(.douta(w_G3548_4[0]),.doutb(w_G3548_4[1]),.doutc(w_G3548_4[2]),.din(w_G3548_1[0]));
	jspl jspl_w_G3552_0(.douta(w_G3552_0[0]),.doutb(w_G3552_0[1]),.din(G3552));
	jspl jspl_w_G3717_0(.douta(w_dff_A_iA5EtpUZ7_0),.doutb(w_G3717_0[1]),.din(G3717));
	jspl3 jspl3_w_G3724_0(.douta(w_dff_A_f94wbbgQ4_0),.doutb(w_G3724_0[1]),.doutc(w_dff_A_QtV3GtD43_2),.din(G3724));
	jspl3 jspl3_w_G4087_0(.douta(w_G4087_0[0]),.doutb(w_dff_A_bHB1uaTW0_1),.doutc(w_G4087_0[2]),.din(G4087));
	jspl3 jspl3_w_G4088_0(.douta(w_G4088_0[0]),.doutb(w_G4088_0[1]),.doutc(w_dff_A_tXtXJkyC4_2),.din(G4088));
	jspl3 jspl3_w_G4089_0(.douta(w_G4089_0[0]),.doutb(w_G4089_0[1]),.doutc(w_dff_A_KdvOQBlZ5_2),.din(G4089));
	jspl3 jspl3_w_G4090_0(.douta(w_G4090_0[0]),.doutb(w_dff_A_cq0xHiKF9_1),.doutc(w_G4090_0[2]),.din(G4090));
	jspl3 jspl3_w_G4091_0(.douta(w_G4091_0[0]),.doutb(w_G4091_0[1]),.doutc(w_dff_A_p7lWIDlr6_2),.din(G4091));
	jspl3 jspl3_w_G4091_1(.douta(w_G4091_1[0]),.doutb(w_dff_A_hl1WHQlu0_1),.doutc(w_dff_A_Dcor2tS24_2),.din(w_G4091_0[0]));
	jspl3 jspl3_w_G4091_2(.douta(w_G4091_2[0]),.doutb(w_G4091_2[1]),.doutc(w_dff_A_AAaitIOj4_2),.din(w_G4091_0[1]));
	jspl3 jspl3_w_G4092_0(.douta(w_G4092_0[0]),.doutb(w_G4092_0[1]),.doutc(w_G4092_0[2]),.din(G4092));
	jspl3 jspl3_w_G4092_1(.douta(w_dff_A_HioiWyno7_0),.doutb(w_dff_A_tiqr3PDH6_1),.doutc(w_G4092_1[2]),.din(w_G4092_0[0]));
	jspl jspl_w_G599_0(.douta(w_G599_0),.doutb(w_dff_A_3L9jc5wg9_1),.din(G599_fa_));
	jspl jspl_w_G600_0(.douta(w_G600_0),.doutb(w_dff_A_p2Avj4Ok5_1),.din(G600_fa_));
	jspl jspl_w_G601_0(.douta(w_dff_A_24pca0HV7_0),.doutb(w_dff_A_dz8Ft8Lm5_1),.din(G601_fa_));
	jspl jspl_w_G611_0(.douta(w_G611_0),.doutb(w_dff_A_u0F4vmwG6_1),.din(G611_fa_));
	jspl jspl_w_G612_0(.douta(w_G612_0),.doutb(w_dff_A_vV76YNP35_1),.din(G612_fa_));
	jspl3 jspl3_w_G809_0(.douta(w_G809_0[0]),.doutb(w_G809_0[1]),.doutc(w_G809_0[2]),.din(G809_fa_));
	jspl3 jspl3_w_G809_1(.douta(w_G809_1[0]),.doutb(w_G809_1[1]),.doutc(w_G809_1[2]),.din(w_G809_0[0]));
	jspl3 jspl3_w_G809_2(.douta(w_G809_2[0]),.doutb(w_G809_2[1]),.doutc(w_G809_2[2]),.din(w_G809_0[1]));
	jspl3 jspl3_w_G809_3(.douta(w_G809_3[0]),.doutb(w_G809_3[1]),.doutc(w_dff_A_Wkcf8uO35_2),.din(w_G809_0[2]));
	jspl jspl_w_G593_0(.douta(w_G593_0),.doutb(w_dff_A_iy5NfA8p1_1),.din(G593_fa_));
	jspl jspl_w_G822_0(.douta(w_G822_0),.doutb(w_dff_A_q1tFT8lp8_1),.din(G822_fa_));
	jspl jspl_w_G838_0(.douta(w_G838_0),.doutb(w_dff_A_AYO72yhU1_1),.din(G838_fa_));
	jspl jspl_w_G861_0(.douta(w_G861_0),.doutb(w_dff_A_KfJFor9N7_1),.din(G861_fa_));
	jspl jspl_w_G832_0(.douta(w_G832_0),.doutb(w_dff_A_0wXNdgG84_1),.din(G832_fa_));
	jspl jspl_w_G834_0(.douta(w_G834_0),.doutb(w_dff_A_wKLlrNjI5_1),.din(G834_fa_));
	jspl jspl_w_G836_0(.douta(w_G836_0),.doutb(w_dff_A_ScVFdJA46_1),.din(G836_fa_));
	jspl jspl_w_G871_0(.douta(w_G871_0),.doutb(w_dff_A_xqc4ukvK3_1),.din(G871_fa_));
	jspl jspl_w_G873_0(.douta(w_G873_0),.doutb(w_dff_A_R11IaAAo2_1),.din(G873_fa_));
	jspl jspl_w_G875_0(.douta(w_G875_0),.doutb(w_dff_A_UWtWUJzu5_1),.din(G875_fa_));
	jspl jspl_w_G877_0(.douta(w_G877_0),.doutb(w_dff_A_cO0UkzHS2_1),.din(G877_fa_));
	jspl jspl_w_G1000_0(.douta(w_G1000_0),.doutb(w_dff_A_yoQ7gBu71_1),.din(G1000_fa_));
	jspl jspl_w_G826_0(.douta(w_G826_0),.doutb(w_dff_A_dwolBJTY9_1),.din(G826_fa_));
	jspl jspl_w_G828_0(.douta(w_G828_0),.doutb(w_dff_A_3wJHFv7k4_1),.din(G828_fa_));
	jspl jspl_w_G830_0(.douta(w_G830_0),.doutb(w_dff_A_MBb3kScK9_1),.din(G830_fa_));
	jspl jspl_w_G867_0(.douta(w_G867_0),.doutb(w_dff_A_JgOw3Pju8_1),.din(G867_fa_));
	jspl jspl_w_G869_0(.douta(w_G869_0),.doutb(w_dff_A_4kASBhIa2_1),.din(G869_fa_));
	jspl jspl_w_n316_0(.douta(w_n316_0[0]),.doutb(w_n316_0[1]),.din(n316));
	jspl jspl_w_n318_0(.douta(w_n318_0[0]),.doutb(w_n318_0[1]),.din(n318));
	jspl3 jspl3_w_n326_0(.douta(w_n326_0[0]),.doutb(w_n326_0[1]),.doutc(w_n326_0[2]),.din(n326));
	jspl3 jspl3_w_n326_1(.douta(w_n326_1[0]),.doutb(w_n326_1[1]),.doutc(w_n326_1[2]),.din(w_n326_0[0]));
	jspl jspl_w_n326_2(.douta(w_n326_2[0]),.doutb(w_n326_2[1]),.din(w_n326_0[1]));
	jspl jspl_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.din(w_dff_B_UXVU0Ypt4_2));
	jspl jspl_w_n336_0(.douta(w_n336_0[0]),.doutb(w_n336_0[1]),.din(n336));
	jspl jspl_w_n360_0(.douta(w_n360_0[0]),.doutb(w_n360_0[1]),.din(n360));
	jspl jspl_w_n362_0(.douta(w_dff_A_E50FNLHQ9_0),.doutb(w_n362_0[1]),.din(n362));
	jspl3 jspl3_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.doutc(w_n366_0[2]),.din(n366));
	jspl3 jspl3_w_n366_1(.douta(w_n366_1[0]),.doutb(w_n366_1[1]),.doutc(w_n366_1[2]),.din(w_n366_0[0]));
	jspl3 jspl3_w_n366_2(.douta(w_n366_2[0]),.doutb(w_n366_2[1]),.doutc(w_n366_2[2]),.din(w_n366_0[1]));
	jspl3 jspl3_w_n366_3(.douta(w_n366_3[0]),.doutb(w_n366_3[1]),.doutc(w_n366_3[2]),.din(w_n366_0[2]));
	jspl3 jspl3_w_n366_4(.douta(w_n366_4[0]),.doutb(w_n366_4[1]),.doutc(w_n366_4[2]),.din(w_n366_1[0]));
	jspl3 jspl3_w_n368_0(.douta(w_n368_0[0]),.doutb(w_n368_0[1]),.doutc(w_n368_0[2]),.din(n368));
	jspl3 jspl3_w_n368_1(.douta(w_n368_1[0]),.doutb(w_n368_1[1]),.doutc(w_n368_1[2]),.din(w_n368_0[0]));
	jspl3 jspl3_w_n368_2(.douta(w_n368_2[0]),.doutb(w_n368_2[1]),.doutc(w_n368_2[2]),.din(w_n368_0[1]));
	jspl3 jspl3_w_n368_3(.douta(w_n368_3[0]),.doutb(w_n368_3[1]),.doutc(w_n368_3[2]),.din(w_n368_0[2]));
	jspl3 jspl3_w_n368_4(.douta(w_n368_4[0]),.doutb(w_n368_4[1]),.doutc(w_n368_4[2]),.din(w_n368_1[0]));
	jspl jspl_w_n368_5(.douta(w_n368_5[0]),.doutb(w_n368_5[1]),.din(w_n368_1[1]));
	jspl3 jspl3_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.doutc(w_n372_0[2]),.din(n372));
	jspl jspl_w_n373_0(.douta(w_n373_0[0]),.doutb(w_n373_0[1]),.din(n373));
	jspl3 jspl3_w_n383_0(.douta(w_n383_0[0]),.doutb(w_n383_0[1]),.doutc(w_n383_0[2]),.din(n383));
	jspl3 jspl3_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.doutc(w_n385_0[2]),.din(n385));
	jspl3 jspl3_w_n385_1(.douta(w_n385_1[0]),.doutb(w_n385_1[1]),.doutc(w_n385_1[2]),.din(w_n385_0[0]));
	jspl3 jspl3_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.doutc(w_n386_0[2]),.din(n386));
	jspl3 jspl3_w_n386_1(.douta(w_n386_1[0]),.doutb(w_n386_1[1]),.doutc(w_n386_1[2]),.din(w_n386_0[0]));
	jspl3 jspl3_w_n386_2(.douta(w_n386_2[0]),.doutb(w_n386_2[1]),.doutc(w_n386_2[2]),.din(w_n386_0[1]));
	jspl3 jspl3_w_n386_3(.douta(w_n386_3[0]),.doutb(w_n386_3[1]),.doutc(w_n386_3[2]),.din(w_n386_0[2]));
	jspl3 jspl3_w_n386_4(.douta(w_n386_4[0]),.doutb(w_n386_4[1]),.doutc(w_n386_4[2]),.din(w_n386_1[0]));
	jspl3 jspl3_w_n388_0(.douta(w_n388_0[0]),.doutb(w_n388_0[1]),.doutc(w_dff_A_a3hhoJix0_2),.din(w_dff_B_yHrQBdqF8_3));
	jspl3 jspl3_w_n388_1(.douta(w_dff_A_HIVMkKha8_0),.doutb(w_dff_A_sYehwKfj0_1),.doutc(w_n388_1[2]),.din(w_n388_0[0]));
	jspl3 jspl3_w_n389_0(.douta(w_n389_0[0]),.doutb(w_n389_0[1]),.doutc(w_n389_0[2]),.din(n389));
	jspl3 jspl3_w_n389_1(.douta(w_n389_1[0]),.doutb(w_n389_1[1]),.doutc(w_n389_1[2]),.din(w_n389_0[0]));
	jspl3 jspl3_w_n389_2(.douta(w_n389_2[0]),.doutb(w_n389_2[1]),.doutc(w_n389_2[2]),.din(w_n389_0[1]));
	jspl3 jspl3_w_n389_3(.douta(w_n389_3[0]),.doutb(w_n389_3[1]),.doutc(w_n389_3[2]),.din(w_n389_0[2]));
	jspl3 jspl3_w_n389_4(.douta(w_n389_4[0]),.doutb(w_n389_4[1]),.doutc(w_n389_4[2]),.din(w_n389_1[0]));
	jspl jspl_w_n397_0(.douta(w_n397_0[0]),.doutb(w_dff_A_63OKJmVU5_1),.din(n397));
	jspl3 jspl3_w_n398_0(.douta(w_n398_0[0]),.doutb(w_n398_0[1]),.doutc(w_n398_0[2]),.din(n398));
	jspl3 jspl3_w_n401_0(.douta(w_dff_A_tYEALtjI1_0),.doutb(w_n401_0[1]),.doutc(w_dff_A_55YIOMal5_2),.din(n401));
	jspl3 jspl3_w_n402_0(.douta(w_n402_0[0]),.doutb(w_n402_0[1]),.doutc(w_n402_0[2]),.din(n402));
	jspl3 jspl3_w_n402_1(.douta(w_n402_1[0]),.doutb(w_n402_1[1]),.doutc(w_n402_1[2]),.din(w_n402_0[0]));
	jspl jspl_w_n402_2(.douta(w_n402_2[0]),.doutb(w_n402_2[1]),.din(w_n402_0[1]));
	jspl jspl_w_n403_0(.douta(w_n403_0[0]),.doutb(w_n403_0[1]),.din(n403));
	jspl3 jspl3_w_n405_0(.douta(w_n405_0[0]),.doutb(w_n405_0[1]),.doutc(w_n405_0[2]),.din(n405));
	jspl3 jspl3_w_n405_1(.douta(w_n405_1[0]),.doutb(w_n405_1[1]),.doutc(w_n405_1[2]),.din(w_n405_0[0]));
	jspl jspl_w_n405_2(.douta(w_n405_2[0]),.doutb(w_n405_2[1]),.din(w_n405_0[1]));
	jspl jspl_w_n407_0(.douta(w_n407_0[0]),.doutb(w_n407_0[1]),.din(n407));
	jspl jspl_w_n408_0(.douta(w_n408_0[0]),.doutb(w_n408_0[1]),.din(n408));
	jspl3 jspl3_w_n410_0(.douta(w_n410_0[0]),.doutb(w_n410_0[1]),.doutc(w_dff_A_tVLIpjof3_2),.din(n410));
	jspl jspl_w_n410_1(.douta(w_dff_A_RHDn8gJ77_0),.doutb(w_n410_1[1]),.din(w_n410_0[0]));
	jspl jspl_w_n414_0(.douta(w_n414_0[0]),.doutb(w_n414_0[1]),.din(n414));
	jspl jspl_w_n416_0(.douta(w_n416_0[0]),.doutb(w_n416_0[1]),.din(n416));
	jspl3 jspl3_w_n419_0(.douta(w_n419_0[0]),.doutb(w_n419_0[1]),.doutc(w_n419_0[2]),.din(n419));
	jspl3 jspl3_w_n424_0(.douta(w_n424_0[0]),.doutb(w_n424_0[1]),.doutc(w_n424_0[2]),.din(n424));
	jspl3 jspl3_w_n424_1(.douta(w_n424_1[0]),.doutb(w_n424_1[1]),.doutc(w_n424_1[2]),.din(w_n424_0[0]));
	jspl jspl_w_n424_2(.douta(w_n424_2[0]),.doutb(w_n424_2[1]),.din(w_n424_0[1]));
	jspl jspl_w_n426_0(.douta(w_n426_0[0]),.doutb(w_dff_A_t9VyOwxo3_1),.din(n426));
	jspl jspl_w_n434_0(.douta(w_n434_0[0]),.doutb(w_n434_0[1]),.din(n434));
	jspl3 jspl3_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.doutc(w_n435_0[2]),.din(n435));
	jspl3 jspl3_w_n435_1(.douta(w_n435_1[0]),.doutb(w_n435_1[1]),.doutc(w_n435_1[2]),.din(w_n435_0[0]));
	jspl3 jspl3_w_n437_0(.douta(w_dff_A_ugTUNeBj5_0),.doutb(w_n437_0[1]),.doutc(w_dff_A_UKFq0IAf2_2),.din(n437));
	jspl3 jspl3_w_n437_1(.douta(w_dff_A_wnFGLyFC2_0),.doutb(w_dff_A_W8kNSJ959_1),.doutc(w_n437_1[2]),.din(w_n437_0[0]));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl3 jspl3_w_n449_0(.douta(w_n449_0[0]),.doutb(w_n449_0[1]),.doutc(w_n449_0[2]),.din(n449));
	jspl3 jspl3_w_n449_1(.douta(w_n449_1[0]),.doutb(w_n449_1[1]),.doutc(w_n449_1[2]),.din(w_n449_0[0]));
	jspl3 jspl3_w_n451_0(.douta(w_dff_A_gVE6PJP04_0),.doutb(w_n451_0[1]),.doutc(w_dff_A_E1z9zFPw6_2),.din(n451));
	jspl jspl_w_n451_1(.douta(w_dff_A_yGT0P50w9_0),.doutb(w_n451_1[1]),.din(w_n451_0[0]));
	jspl jspl_w_n459_0(.douta(w_n459_0[0]),.doutb(w_dff_A_9vwwXxKD4_1),.din(n459));
	jspl3 jspl3_w_n460_0(.douta(w_n460_0[0]),.doutb(w_n460_0[1]),.doutc(w_n460_0[2]),.din(n460));
	jspl3 jspl3_w_n460_1(.douta(w_n460_1[0]),.doutb(w_n460_1[1]),.doutc(w_n460_1[2]),.din(w_n460_0[0]));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_dff_A_wrTCqjNx6_1),.doutc(w_dff_A_Kn1bkS712_2),.din(n462));
	jspl jspl_w_n470_0(.douta(w_n470_0[0]),.doutb(w_n470_0[1]),.din(n470));
	jspl3 jspl3_w_n471_0(.douta(w_n471_0[0]),.doutb(w_n471_0[1]),.doutc(w_n471_0[2]),.din(n471));
	jspl jspl_w_n471_1(.douta(w_n471_1[0]),.doutb(w_n471_1[1]),.din(w_n471_0[0]));
	jspl3 jspl3_w_n473_0(.douta(w_n473_0[0]),.doutb(w_n473_0[1]),.doutc(w_dff_A_4959dTQj2_2),.din(w_dff_B_cNjfOzIY2_3));
	jspl3 jspl3_w_n473_1(.douta(w_dff_A_M1zNiXjj5_0),.doutb(w_dff_A_5qs9epFC4_1),.doutc(w_n473_1[2]),.din(w_n473_0[0]));
	jspl jspl_w_n481_0(.douta(w_n481_0[0]),.doutb(w_n481_0[1]),.din(n481));
	jspl3 jspl3_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.doutc(w_n484_0[2]),.din(n484));
	jspl jspl_w_n484_1(.douta(w_n484_1[0]),.doutb(w_n484_1[1]),.din(w_n484_0[0]));
	jspl3 jspl3_w_n486_0(.douta(w_dff_A_MVXiMlLm6_0),.doutb(w_n486_0[1]),.doutc(w_dff_A_B8oHIgWy0_2),.din(n486));
	jspl jspl_w_n486_1(.douta(w_dff_A_Iw5jiIn26_0),.doutb(w_n486_1[1]),.din(w_n486_0[0]));
	jspl jspl_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.din(n494));
	jspl3 jspl3_w_n495_0(.douta(w_n495_0[0]),.doutb(w_n495_0[1]),.doutc(w_n495_0[2]),.din(n495));
	jspl3 jspl3_w_n495_1(.douta(w_n495_1[0]),.doutb(w_n495_1[1]),.doutc(w_n495_1[2]),.din(w_n495_0[0]));
	jspl3 jspl3_w_n497_0(.douta(w_dff_A_t8GskBuY4_0),.doutb(w_n497_0[1]),.doutc(w_dff_A_BgIz9GOx3_2),.din(n497));
	jspl jspl_w_n497_1(.douta(w_dff_A_Post4hJQ0_0),.doutb(w_n497_1[1]),.din(w_n497_0[0]));
	jspl jspl_w_n505_0(.douta(w_n505_0[0]),.doutb(w_n505_0[1]),.din(n505));
	jspl3 jspl3_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.doutc(w_n507_0[2]),.din(n507));
	jspl jspl_w_n507_1(.douta(w_n507_1[0]),.doutb(w_n507_1[1]),.din(w_n507_0[0]));
	jspl jspl_w_n509_0(.douta(w_n509_0[0]),.doutb(w_n509_0[1]),.din(w_dff_B_Jr6O50Gx2_2));
	jspl jspl_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.din(n517));
	jspl3 jspl3_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.doutc(w_n518_0[2]),.din(n518));
	jspl jspl_w_n518_1(.douta(w_n518_1[0]),.doutb(w_n518_1[1]),.din(w_n518_0[0]));
	jspl3 jspl3_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.doutc(w_n528_0[2]),.din(n528));
	jspl3 jspl3_w_n530_0(.douta(w_n530_0[0]),.doutb(w_n530_0[1]),.doutc(w_n530_0[2]),.din(n530));
	jspl jspl_w_n530_1(.douta(w_n530_1[0]),.doutb(w_n530_1[1]),.din(w_n530_0[0]));
	jspl jspl_w_n532_0(.douta(w_n532_0[0]),.doutb(w_n532_0[1]),.din(w_dff_B_3kpYIH2t1_2));
	jspl jspl_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.din(n540));
	jspl3 jspl3_w_n541_0(.douta(w_n541_0[0]),.doutb(w_n541_0[1]),.doutc(w_n541_0[2]),.din(n541));
	jspl jspl_w_n541_1(.douta(w_n541_1[0]),.doutb(w_n541_1[1]),.din(w_n541_0[0]));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_dff_A_SCGFeEfB8_1),.din(n543));
	jspl jspl_w_n551_0(.douta(w_n551_0[0]),.doutb(w_n551_0[1]),.din(n551));
	jspl3 jspl3_w_n556_0(.douta(w_n556_0[0]),.doutb(w_n556_0[1]),.doutc(w_n556_0[2]),.din(n556));
	jspl3 jspl3_w_n556_1(.douta(w_n556_1[0]),.doutb(w_n556_1[1]),.doutc(w_n556_1[2]),.din(w_n556_0[0]));
	jspl3 jspl3_w_n556_2(.douta(w_n556_2[0]),.doutb(w_n556_2[1]),.doutc(w_n556_2[2]),.din(w_n556_0[1]));
	jspl3 jspl3_w_n556_3(.douta(w_n556_3[0]),.doutb(w_n556_3[1]),.doutc(w_n556_3[2]),.din(w_n556_0[2]));
	jspl3 jspl3_w_n556_4(.douta(w_n556_4[0]),.doutb(w_n556_4[1]),.doutc(w_n556_4[2]),.din(w_n556_1[0]));
	jspl jspl_w_n556_5(.douta(w_n556_5[0]),.doutb(w_n556_5[1]),.din(w_n556_1[1]));
	jspl3 jspl3_w_n560_0(.douta(w_n560_0[0]),.doutb(w_n560_0[1]),.doutc(w_n560_0[2]),.din(n560));
	jspl jspl_w_n560_1(.douta(w_n560_1[0]),.doutb(w_n560_1[1]),.din(w_n560_0[0]));
	jspl3 jspl3_w_n561_0(.douta(w_dff_A_im8jegML9_0),.doutb(w_dff_A_zoXmK7Iz9_1),.doutc(w_n561_0[2]),.din(n561));
	jspl jspl_w_n562_0(.douta(w_dff_A_uQZAZQvC3_0),.doutb(w_n562_0[1]),.din(w_dff_B_Al0hJv4B7_2));
	jspl3 jspl3_w_n566_0(.douta(w_n566_0[0]),.doutb(w_n566_0[1]),.doutc(w_n566_0[2]),.din(n566));
	jspl3 jspl3_w_n567_0(.douta(w_n567_0[0]),.doutb(w_dff_A_aqXlXeOX2_1),.doutc(w_n567_0[2]),.din(n567));
	jspl jspl_w_n567_1(.douta(w_n567_1[0]),.doutb(w_dff_A_T1e90f7s3_1),.din(w_n567_0[0]));
	jspl jspl_w_n569_0(.douta(w_n569_0[0]),.doutb(w_dff_A_MsUDDw1v4_1),.din(n569));
	jspl jspl_w_n570_0(.douta(w_n570_0[0]),.doutb(w_n570_0[1]),.din(n570));
	jspl3 jspl3_w_n571_0(.douta(w_n571_0[0]),.doutb(w_n571_0[1]),.doutc(w_dff_A_xmhvvj0Z8_2),.din(n571));
	jspl jspl_w_n571_1(.douta(w_n571_1[0]),.doutb(w_n571_1[1]),.din(w_n571_0[0]));
	jspl3 jspl3_w_n572_0(.douta(w_dff_A_vOM2tzt18_0),.doutb(w_n572_0[1]),.doutc(w_n572_0[2]),.din(n572));
	jspl3 jspl3_w_n574_0(.douta(w_n574_0[0]),.doutb(w_n574_0[1]),.doutc(w_n574_0[2]),.din(n574));
	jspl3 jspl3_w_n577_0(.douta(w_n577_0[0]),.doutb(w_n577_0[1]),.doutc(w_n577_0[2]),.din(n577));
	jspl3 jspl3_w_n578_0(.douta(w_n578_0[0]),.doutb(w_dff_A_FaJwG62n8_1),.doutc(w_n578_0[2]),.din(n578));
	jspl3 jspl3_w_n582_0(.douta(w_n582_0[0]),.doutb(w_n582_0[1]),.doutc(w_n582_0[2]),.din(n582));
	jspl jspl_w_n582_1(.douta(w_n582_1[0]),.doutb(w_n582_1[1]),.din(w_n582_0[0]));
	jspl3 jspl3_w_n583_0(.douta(w_n583_0[0]),.doutb(w_n583_0[1]),.doutc(w_dff_A_crk6p3iG6_2),.din(n583));
	jspl jspl_w_n583_1(.douta(w_dff_A_mTq4iD9w4_0),.doutb(w_n583_1[1]),.din(w_n583_0[0]));
	jspl jspl_w_n585_0(.douta(w_dff_A_oyEdJAoc4_0),.doutb(w_n585_0[1]),.din(n585));
	jspl3 jspl3_w_n587_0(.douta(w_n587_0[0]),.doutb(w_n587_0[1]),.doutc(w_n587_0[2]),.din(n587));
	jspl jspl_w_n587_1(.douta(w_n587_1[0]),.doutb(w_n587_1[1]),.din(w_n587_0[0]));
	jspl3 jspl3_w_n590_0(.douta(w_n590_0[0]),.doutb(w_dff_A_FWYweYQo4_1),.doutc(w_n590_0[2]),.din(n590));
	jspl jspl_w_n590_1(.douta(w_n590_1[0]),.doutb(w_n590_1[1]),.din(w_n590_0[0]));
	jspl jspl_w_n591_0(.douta(w_n591_0[0]),.doutb(w_dff_A_lDjO1o2S5_1),.din(n591));
	jspl3 jspl3_w_n595_0(.douta(w_n595_0[0]),.doutb(w_n595_0[1]),.doutc(w_n595_0[2]),.din(n595));
	jspl jspl_w_n595_1(.douta(w_n595_1[0]),.doutb(w_n595_1[1]),.din(w_n595_0[0]));
	jspl3 jspl3_w_n596_0(.douta(w_dff_A_Hgu7Ljw35_0),.doutb(w_n596_0[1]),.doutc(w_n596_0[2]),.din(n596));
	jspl3 jspl3_w_n600_0(.douta(w_n600_0[0]),.doutb(w_n600_0[1]),.doutc(w_n600_0[2]),.din(n600));
	jspl jspl_w_n600_1(.douta(w_n600_1[0]),.doutb(w_n600_1[1]),.din(w_n600_0[0]));
	jspl jspl_w_n601_0(.douta(w_n601_0[0]),.doutb(w_n601_0[1]),.din(n601));
	jspl3 jspl3_w_n604_0(.douta(w_dff_A_qxb4VXKh9_0),.doutb(w_n604_0[1]),.doutc(w_n604_0[2]),.din(n604));
	jspl3 jspl3_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.doutc(w_n605_0[2]),.din(n605));
	jspl3 jspl3_w_n605_1(.douta(w_n605_1[0]),.doutb(w_n605_1[1]),.doutc(w_dff_A_Aw2TO8zp6_2),.din(w_n605_0[0]));
	jspl3 jspl3_w_n605_2(.douta(w_n605_2[0]),.doutb(w_n605_2[1]),.doutc(w_n605_2[2]),.din(w_n605_0[1]));
	jspl3 jspl3_w_n607_0(.douta(w_n607_0[0]),.doutb(w_dff_A_I5VwRkAh7_1),.doutc(w_n607_0[2]),.din(w_dff_B_t1QjbpLO5_3));
	jspl3 jspl3_w_n609_0(.douta(w_n609_0[0]),.doutb(w_n609_0[1]),.doutc(w_n609_0[2]),.din(n609));
	jspl3 jspl3_w_n609_1(.douta(w_n609_1[0]),.doutb(w_n609_1[1]),.doutc(w_n609_1[2]),.din(w_n609_0[0]));
	jspl3 jspl3_w_n609_2(.douta(w_n609_2[0]),.doutb(w_n609_2[1]),.doutc(w_n609_2[2]),.din(w_n609_0[1]));
	jspl3 jspl3_w_n609_3(.douta(w_n609_3[0]),.doutb(w_n609_3[1]),.doutc(w_n609_3[2]),.din(w_n609_0[2]));
	jspl3 jspl3_w_n609_4(.douta(w_n609_4[0]),.doutb(w_n609_4[1]),.doutc(w_n609_4[2]),.din(w_n609_1[0]));
	jspl3 jspl3_w_n609_5(.douta(w_n609_5[0]),.doutb(w_n609_5[1]),.doutc(w_n609_5[2]),.din(w_n609_1[1]));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.doutc(w_n613_0[2]),.din(n613));
	jspl3 jspl3_w_n614_0(.douta(w_n614_0[0]),.doutb(w_dff_A_5lRKS5Go0_1),.doutc(w_dff_A_0LLucqvu0_2),.din(n614));
	jspl3 jspl3_w_n614_1(.douta(w_dff_A_VCistAtS2_0),.doutb(w_n614_1[1]),.doutc(w_dff_A_p8xOZy5d0_2),.din(w_n614_0[0]));
	jspl jspl_w_n614_2(.douta(w_dff_A_sPNwFVsy2_0),.doutb(w_n614_2[1]),.din(w_n614_0[1]));
	jspl3 jspl3_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.doutc(w_n617_0[2]),.din(n617));
	jspl jspl_w_n617_1(.douta(w_n617_1[0]),.doutb(w_n617_1[1]),.din(w_n617_0[0]));
	jspl3 jspl3_w_n618_0(.douta(w_n618_0[0]),.doutb(w_n618_0[1]),.doutc(w_n618_0[2]),.din(n618));
	jspl jspl_w_n618_1(.douta(w_n618_1[0]),.doutb(w_n618_1[1]),.din(w_n618_0[0]));
	jspl3 jspl3_w_n621_0(.douta(w_n621_0[0]),.doutb(w_n621_0[1]),.doutc(w_n621_0[2]),.din(n621));
	jspl3 jspl3_w_n621_1(.douta(w_dff_A_1raUQNaH4_0),.doutb(w_n621_1[1]),.doutc(w_n621_1[2]),.din(w_n621_0[0]));
	jspl jspl_w_n621_2(.douta(w_dff_A_64zhRRF94_0),.doutb(w_n621_2[1]),.din(w_n621_0[1]));
	jspl3 jspl3_w_n622_0(.douta(w_n622_0[0]),.doutb(w_n622_0[1]),.doutc(w_n622_0[2]),.din(n622));
	jspl jspl_w_n622_1(.douta(w_n622_1[0]),.doutb(w_n622_1[1]),.din(w_n622_0[0]));
	jspl jspl_w_n623_0(.douta(w_dff_A_VdAWrNPu1_0),.doutb(w_n623_0[1]),.din(n623));
	jspl3 jspl3_w_n624_0(.douta(w_n624_0[0]),.doutb(w_n624_0[1]),.doutc(w_n624_0[2]),.din(n624));
	jspl3 jspl3_w_n624_1(.douta(w_n624_1[0]),.doutb(w_n624_1[1]),.doutc(w_n624_1[2]),.din(w_n624_0[0]));
	jspl3 jspl3_w_n625_0(.douta(w_dff_A_6FBPsbun8_0),.doutb(w_n625_0[1]),.doutc(w_dff_A_zIdAlXXi9_2),.din(n625));
	jspl3 jspl3_w_n628_0(.douta(w_n628_0[0]),.doutb(w_dff_A_OuIvP6MH8_1),.doutc(w_n628_0[2]),.din(n628));
	jspl3 jspl3_w_n629_0(.douta(w_n629_0[0]),.doutb(w_dff_A_t9pJYt2t9_1),.doutc(w_n629_0[2]),.din(n629));
	jspl jspl_w_n631_0(.douta(w_dff_A_BHyEiyWj8_0),.doutb(w_n631_0[1]),.din(n631));
	jspl3 jspl3_w_n633_0(.douta(w_n633_0[0]),.doutb(w_n633_0[1]),.doutc(w_n633_0[2]),.din(n633));
	jspl jspl_w_n633_1(.douta(w_n633_1[0]),.doutb(w_n633_1[1]),.din(w_n633_0[0]));
	jspl3 jspl3_w_n636_0(.douta(w_n636_0[0]),.doutb(w_n636_0[1]),.doutc(w_dff_A_6BEI3sAR2_2),.din(n636));
	jspl jspl_w_n636_1(.douta(w_n636_1[0]),.doutb(w_dff_A_l10nIiRm6_1),.din(w_n636_0[0]));
	jspl3 jspl3_w_n640_0(.douta(w_n640_0[0]),.doutb(w_dff_A_1SvuEk1l6_1),.doutc(w_dff_A_LO8JhS1b5_2),.din(n640));
	jspl3 jspl3_w_n640_1(.douta(w_dff_A_D7AxmQ9P6_0),.doutb(w_n640_1[1]),.doutc(w_n640_1[2]),.din(w_n640_0[0]));
	jspl jspl_w_n641_0(.douta(w_n641_0[0]),.doutb(w_n641_0[1]),.din(n641));
	jspl jspl_w_n642_0(.douta(w_n642_0[0]),.doutb(w_n642_0[1]),.din(n642));
	jspl3 jspl3_w_n645_0(.douta(w_n645_0[0]),.doutb(w_n645_0[1]),.doutc(w_n645_0[2]),.din(n645));
	jspl3 jspl3_w_n646_0(.douta(w_dff_A_6BIevfPr4_0),.doutb(w_n646_0[1]),.doutc(w_n646_0[2]),.din(n646));
	jspl3 jspl3_w_n649_0(.douta(w_n649_0[0]),.doutb(w_n649_0[1]),.doutc(w_dff_A_h601iIzf1_2),.din(n649));
	jspl jspl_w_n649_1(.douta(w_n649_1[0]),.doutb(w_n649_1[1]),.din(w_n649_0[0]));
	jspl jspl_w_n650_0(.douta(w_dff_A_Td0FQIsI3_0),.doutb(w_n650_0[1]),.din(n650));
	jspl3 jspl3_w_n651_0(.douta(w_n651_0[0]),.doutb(w_dff_A_tPlTKaWH6_1),.doutc(w_dff_A_HqFGmp4m9_2),.din(w_dff_B_HqYOc0uM0_3));
	jspl jspl_w_n651_1(.douta(w_dff_A_IG1CENs25_0),.doutb(w_n651_1[1]),.din(w_n651_0[0]));
	jspl jspl_w_n652_0(.douta(w_n652_0[0]),.doutb(w_n652_0[1]),.din(w_dff_B_7iy6Kj3D8_2));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_n661_0[1]),.din(n661));
	jspl jspl_w_n671_0(.douta(w_dff_A_tO90tMmr9_0),.doutb(w_n671_0[1]),.din(n671));
	jspl jspl_w_n677_0(.douta(w_n677_0[0]),.doutb(w_n677_0[1]),.din(n677));
	jspl jspl_w_n678_0(.douta(w_n678_0[0]),.doutb(w_dff_A_8N7eNG3U7_1),.din(n678));
	jspl jspl_w_n679_0(.douta(w_n679_0[0]),.doutb(w_dff_A_4qE7KPEQ0_1),.din(n679));
	jspl jspl_w_n680_0(.douta(w_n680_0[0]),.doutb(w_dff_A_gIyESD6S9_1),.din(w_dff_B_JaGxgQWT2_2));
	jspl3 jspl3_w_n681_0(.douta(w_n681_0[0]),.doutb(w_n681_0[1]),.doutc(w_n681_0[2]),.din(n681));
	jspl3 jspl3_w_n681_1(.douta(w_dff_A_5ZnwEata7_0),.doutb(w_dff_A_IznMhbn49_1),.doutc(w_n681_1[2]),.din(w_n681_0[0]));
	jspl jspl_w_n681_2(.douta(w_dff_A_7EVxPVdw9_0),.doutb(w_n681_2[1]),.din(w_n681_0[1]));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.din(n682));
	jspl3 jspl3_w_n687_0(.douta(w_dff_A_geAXsMnP2_0),.doutb(w_dff_A_DcXsmqnS8_1),.doutc(w_n687_0[2]),.din(n687));
	jspl jspl_w_n689_0(.douta(w_dff_A_UIiibPO25_0),.doutb(w_n689_0[1]),.din(n689));
	jspl3 jspl3_w_n691_0(.douta(w_n691_0[0]),.doutb(w_dff_A_8wQEgTCA2_1),.doutc(w_n691_0[2]),.din(n691));
	jspl3 jspl3_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.doutc(w_n693_0[2]),.din(n693));
	jspl3 jspl3_w_n696_0(.douta(w_n696_0[0]),.doutb(w_n696_0[1]),.doutc(w_n696_0[2]),.din(n696));
	jspl jspl_w_n697_0(.douta(w_n697_0[0]),.doutb(w_n697_0[1]),.din(n697));
	jspl jspl_w_n700_0(.douta(w_n700_0[0]),.doutb(w_dff_A_PPHdl43q8_1),.din(n700));
	jspl jspl_w_n702_0(.douta(w_n702_0[0]),.doutb(w_n702_0[1]),.din(w_dff_B_rsIdIZLY8_2));
	jspl3 jspl3_w_n703_0(.douta(w_n703_0[0]),.doutb(w_n703_0[1]),.doutc(w_n703_0[2]),.din(n703));
	jspl jspl_w_n705_0(.douta(w_n705_0[0]),.doutb(w_n705_0[1]),.din(n705));
	jspl jspl_w_n706_0(.douta(w_dff_A_Lg42zLWs3_0),.doutb(w_n706_0[1]),.din(n706));
	jspl3 jspl3_w_n707_0(.douta(w_n707_0[0]),.doutb(w_n707_0[1]),.doutc(w_n707_0[2]),.din(n707));
	jspl jspl_w_n709_0(.douta(w_n709_0[0]),.doutb(w_n709_0[1]),.din(w_dff_B_aRARWFLQ8_2));
	jspl jspl_w_n716_0(.douta(w_n716_0[0]),.doutb(w_n716_0[1]),.din(n716));
	jspl3 jspl3_w_n717_0(.douta(w_n717_0[0]),.doutb(w_dff_A_b8mN4CkN8_1),.doutc(w_dff_A_VhxFh8dI9_2),.din(n717));
	jspl jspl_w_n720_0(.douta(w_n720_0[0]),.doutb(w_n720_0[1]),.din(n720));
	jspl3 jspl3_w_n721_0(.douta(w_n721_0[0]),.doutb(w_dff_A_RRSfynhV3_1),.doutc(w_n721_0[2]),.din(n721));
	jspl jspl_w_n723_0(.douta(w_dff_A_2osJTg5r6_0),.doutb(w_n723_0[1]),.din(n723));
	jspl jspl_w_n726_0(.douta(w_n726_0[0]),.doutb(w_n726_0[1]),.din(n726));
	jspl3 jspl3_w_n727_0(.douta(w_n727_0[0]),.doutb(w_n727_0[1]),.doutc(w_n727_0[2]),.din(n727));
	jspl3 jspl3_w_n729_0(.douta(w_n729_0[0]),.doutb(w_n729_0[1]),.doutc(w_n729_0[2]),.din(n729));
	jspl jspl_w_n729_1(.douta(w_n729_1[0]),.doutb(w_n729_1[1]),.din(w_n729_0[0]));
	jspl3 jspl3_w_n732_0(.douta(w_n732_0[0]),.doutb(w_n732_0[1]),.doutc(w_n732_0[2]),.din(n732));
	jspl jspl_w_n733_0(.douta(w_n733_0[0]),.doutb(w_n733_0[1]),.din(n733));
	jspl jspl_w_n735_0(.douta(w_n735_0[0]),.doutb(w_n735_0[1]),.din(n735));
	jspl jspl_w_n736_0(.douta(w_n736_0[0]),.doutb(w_n736_0[1]),.din(n736));
	jspl3 jspl3_w_n739_0(.douta(w_n739_0[0]),.doutb(w_n739_0[1]),.doutc(w_dff_A_ZiHBGFqw1_2),.din(n739));
	jspl jspl_w_n739_1(.douta(w_dff_A_0Yj7e50W7_0),.doutb(w_n739_1[1]),.din(w_n739_0[0]));
	jspl jspl_w_n740_0(.douta(w_n740_0[0]),.doutb(w_dff_A_NgjfhL585_1),.din(n740));
	jspl jspl_w_n741_0(.douta(w_dff_A_S50wsJSu9_0),.doutb(w_n741_0[1]),.din(n741));
	jspl jspl_w_n742_0(.douta(w_n742_0[0]),.doutb(w_n742_0[1]),.din(w_dff_B_jfeEQVgx4_2));
	jspl3 jspl3_w_n744_0(.douta(w_n744_0[0]),.doutb(w_n744_0[1]),.doutc(w_dff_A_AhU7oceG6_2),.din(w_dff_B_IRVa1Pmb5_3));
	jspl3 jspl3_w_n744_1(.douta(w_dff_A_4v02IntC4_0),.doutb(w_n744_1[1]),.doutc(w_n744_1[2]),.din(w_n744_0[0]));
	jspl3 jspl3_w_n746_0(.douta(w_n746_0[0]),.doutb(w_n746_0[1]),.doutc(w_dff_A_mTgfSlbB7_2),.din(n746));
	jspl3 jspl3_w_n746_1(.douta(w_n746_1[0]),.doutb(w_n746_1[1]),.doutc(w_n746_1[2]),.din(w_n746_0[0]));
	jspl3 jspl3_w_n747_0(.douta(w_dff_A_4H65fA2y3_0),.doutb(w_dff_A_gZRPnmG56_1),.doutc(w_n747_0[2]),.din(n747));
	jspl3 jspl3_w_n747_1(.douta(w_n747_1[0]),.doutb(w_dff_A_vsXEra7e3_1),.doutc(w_dff_A_iT9fQLBz5_2),.din(w_n747_0[0]));
	jspl3 jspl3_w_n747_2(.douta(w_dff_A_NrSQtPIH1_0),.doutb(w_dff_A_46KeFG3T5_1),.doutc(w_n747_2[2]),.din(w_n747_0[1]));
	jspl3 jspl3_w_n747_3(.douta(w_dff_A_COGThtqU9_0),.doutb(w_dff_A_mE9sZeDh0_1),.doutc(w_n747_3[2]),.din(w_n747_0[2]));
	jspl3 jspl3_w_n748_0(.douta(w_n748_0[0]),.doutb(w_dff_A_UfZ86a0w8_1),.doutc(w_dff_A_N4ptuOW26_2),.din(w_dff_B_ihQVpXUD7_3));
	jspl3 jspl3_w_n748_1(.douta(w_n748_1[0]),.doutb(w_dff_A_pVTYFNtE9_1),.doutc(w_dff_A_38LaT17l8_2),.din(w_n748_0[0]));
	jspl3 jspl3_w_n748_2(.douta(w_dff_A_xIckdFqs7_0),.doutb(w_n748_2[1]),.doutc(w_dff_A_6f8Kk6ui9_2),.din(w_n748_0[1]));
	jspl3 jspl3_w_n748_3(.douta(w_n748_3[0]),.doutb(w_dff_A_8g0vU4iT8_1),.doutc(w_dff_A_4NeCTvRO6_2),.din(w_n748_0[2]));
	jspl jspl_w_n748_4(.douta(w_dff_A_iUVppLLC3_0),.doutb(w_n748_4[1]),.din(w_n748_1[0]));
	jspl3 jspl3_w_n750_0(.douta(w_n750_0[0]),.doutb(w_dff_A_PqAu7HDC8_1),.doutc(w_dff_A_7VL5Q9WW4_2),.din(n750));
	jspl jspl_w_n750_1(.douta(w_n750_1[0]),.doutb(w_n750_1[1]),.din(w_n750_0[0]));
	jspl3 jspl3_w_n751_0(.douta(w_dff_A_b3F2XRIP3_0),.doutb(w_n751_0[1]),.doutc(w_dff_A_uIcXy7Ld2_2),.din(n751));
	jspl3 jspl3_w_n751_1(.douta(w_n751_1[0]),.doutb(w_dff_A_3ZPaxM2o1_1),.doutc(w_n751_1[2]),.din(w_n751_0[0]));
	jspl jspl_w_n751_2(.douta(w_n751_2[0]),.doutb(w_dff_A_wIJmSegh5_1),.din(w_n751_0[1]));
	jspl3 jspl3_w_n753_0(.douta(w_n753_0[0]),.doutb(w_n753_0[1]),.doutc(w_n753_0[2]),.din(n753));
	jspl3 jspl3_w_n753_1(.douta(w_n753_1[0]),.doutb(w_n753_1[1]),.doutc(w_n753_1[2]),.din(w_n753_0[0]));
	jspl3 jspl3_w_n753_2(.douta(w_n753_2[0]),.doutb(w_n753_2[1]),.doutc(w_n753_2[2]),.din(w_n753_0[1]));
	jspl3 jspl3_w_n753_3(.douta(w_n753_3[0]),.doutb(w_n753_3[1]),.doutc(w_n753_3[2]),.din(w_n753_0[2]));
	jspl3 jspl3_w_n753_4(.douta(w_n753_4[0]),.doutb(w_n753_4[1]),.doutc(w_n753_4[2]),.din(w_n753_1[0]));
	jspl3 jspl3_w_n753_5(.douta(w_n753_5[0]),.doutb(w_n753_5[1]),.doutc(w_n753_5[2]),.din(w_n753_1[1]));
	jspl3 jspl3_w_n753_6(.douta(w_n753_6[0]),.doutb(w_n753_6[1]),.doutc(w_n753_6[2]),.din(w_n753_1[2]));
	jspl3 jspl3_w_n753_7(.douta(w_n753_7[0]),.doutb(w_n753_7[1]),.doutc(w_n753_7[2]),.din(w_n753_2[0]));
	jspl jspl_w_n753_8(.douta(w_n753_8[0]),.doutb(w_n753_8[1]),.din(w_n753_2[1]));
	jspl jspl_w_n759_0(.douta(w_n759_0[0]),.doutb(w_n759_0[1]),.din(n759));
	jspl jspl_w_n760_0(.douta(w_n760_0[0]),.doutb(w_n760_0[1]),.din(n760));
	jspl jspl_w_n761_0(.douta(w_n761_0[0]),.doutb(w_n761_0[1]),.din(n761));
	jspl3 jspl3_w_n765_0(.douta(w_n765_0[0]),.doutb(w_n765_0[1]),.doutc(w_n765_0[2]),.din(w_dff_B_zVEI9lAu4_3));
	jspl3 jspl3_w_n765_1(.douta(w_n765_1[0]),.doutb(w_n765_1[1]),.doutc(w_n765_1[2]),.din(w_n765_0[0]));
	jspl3 jspl3_w_n765_2(.douta(w_n765_2[0]),.doutb(w_n765_2[1]),.doutc(w_n765_2[2]),.din(w_n765_0[1]));
	jspl3 jspl3_w_n765_3(.douta(w_n765_3[0]),.doutb(w_n765_3[1]),.doutc(w_n765_3[2]),.din(w_n765_0[2]));
	jspl3 jspl3_w_n765_4(.douta(w_n765_4[0]),.doutb(w_n765_4[1]),.doutc(w_n765_4[2]),.din(w_n765_1[0]));
	jspl3 jspl3_w_n765_5(.douta(w_n765_5[0]),.doutb(w_n765_5[1]),.doutc(w_n765_5[2]),.din(w_n765_1[1]));
	jspl jspl_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.din(n771));
	jspl jspl_w_n779_0(.douta(w_n779_0[0]),.doutb(w_dff_A_MaU7TXpH9_1),.din(n779));
	jspl3 jspl3_w_n781_0(.douta(w_n781_0[0]),.doutb(w_n781_0[1]),.doutc(w_n781_0[2]),.din(n781));
	jspl3 jspl3_w_n783_0(.douta(w_n783_0[0]),.doutb(w_n783_0[1]),.doutc(w_n783_0[2]),.din(n783));
	jspl jspl_w_n783_1(.douta(w_n783_1[0]),.doutb(w_n783_1[1]),.din(w_n783_0[0]));
	jspl jspl_w_n786_0(.douta(w_n786_0[0]),.doutb(w_n786_0[1]),.din(n786));
	jspl jspl_w_n787_0(.douta(w_n787_0[0]),.doutb(w_n787_0[1]),.din(w_dff_B_FSISOWg23_2));
	jspl3 jspl3_w_n789_0(.douta(w_n789_0[0]),.doutb(w_n789_0[1]),.doutc(w_n789_0[2]),.din(n789));
	jspl3 jspl3_w_n791_0(.douta(w_n791_0[0]),.doutb(w_n791_0[1]),.doutc(w_n791_0[2]),.din(n791));
	jspl jspl_w_n791_1(.douta(w_n791_1[0]),.doutb(w_n791_1[1]),.din(w_n791_0[0]));
	jspl jspl_w_n792_0(.douta(w_n792_0[0]),.doutb(w_n792_0[1]),.din(n792));
	jspl3 jspl3_w_n793_0(.douta(w_n793_0[0]),.doutb(w_dff_A_dYGaO07l1_1),.doutc(w_dff_A_AeEiZwLg7_2),.din(w_dff_B_yK95vB9c5_3));
	jspl3 jspl3_w_n793_1(.douta(w_n793_1[0]),.doutb(w_dff_A_wYf4CRIS1_1),.doutc(w_dff_A_0Wy3drpl8_2),.din(w_n793_0[0]));
	jspl3 jspl3_w_n793_2(.douta(w_n793_2[0]),.doutb(w_n793_2[1]),.doutc(w_dff_A_pjgPQuD18_2),.din(w_n793_0[1]));
	jspl3 jspl3_w_n793_3(.douta(w_n793_3[0]),.doutb(w_dff_A_cyhATo4q5_1),.doutc(w_dff_A_Z3YaYsW56_2),.din(w_n793_0[2]));
	jspl jspl_w_n793_4(.douta(w_dff_A_zKo6lCdE9_0),.doutb(w_n793_4[1]),.din(w_n793_1[0]));
	jspl3 jspl3_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.doutc(w_n795_0[2]),.din(n795));
	jspl jspl_w_n795_1(.douta(w_n795_1[0]),.doutb(w_n795_1[1]),.din(w_n795_0[0]));
	jspl jspl_w_n796_0(.douta(w_n796_0[0]),.doutb(w_n796_0[1]),.din(n796));
	jspl3 jspl3_w_n797_0(.douta(w_n797_0[0]),.doutb(w_dff_A_vufs09fJ5_1),.doutc(w_dff_A_V3S91piA1_2),.din(w_dff_B_p44IFa8m3_3));
	jspl3 jspl3_w_n797_1(.douta(w_n797_1[0]),.doutb(w_dff_A_1PVE3DRf5_1),.doutc(w_dff_A_hL4526bv5_2),.din(w_n797_0[0]));
	jspl3 jspl3_w_n797_2(.douta(w_n797_2[0]),.doutb(w_n797_2[1]),.doutc(w_dff_A_sFWHDYan7_2),.din(w_n797_0[1]));
	jspl3 jspl3_w_n797_3(.douta(w_n797_3[0]),.doutb(w_dff_A_RzFTeu7T9_1),.doutc(w_dff_A_ryKJwIR74_2),.din(w_n797_0[2]));
	jspl jspl_w_n797_4(.douta(w_dff_A_yGyRJSXA9_0),.doutb(w_n797_4[1]),.din(w_n797_1[0]));
	jspl3 jspl3_w_n799_0(.douta(w_n799_0[0]),.doutb(w_n799_0[1]),.doutc(w_n799_0[2]),.din(n799));
	jspl3 jspl3_w_n799_1(.douta(w_n799_1[0]),.doutb(w_n799_1[1]),.doutc(w_n799_1[2]),.din(w_n799_0[0]));
	jspl3 jspl3_w_n799_2(.douta(w_n799_2[0]),.doutb(w_n799_2[1]),.doutc(w_n799_2[2]),.din(w_n799_0[1]));
	jspl3 jspl3_w_n799_3(.douta(w_n799_3[0]),.doutb(w_n799_3[1]),.doutc(w_n799_3[2]),.din(w_n799_0[2]));
	jspl jspl_w_n799_4(.douta(w_n799_4[0]),.doutb(w_n799_4[1]),.din(w_n799_1[0]));
	jspl3 jspl3_w_n801_0(.douta(w_n801_0[0]),.doutb(w_n801_0[1]),.doutc(w_n801_0[2]),.din(n801));
	jspl3 jspl3_w_n801_1(.douta(w_n801_1[0]),.doutb(w_n801_1[1]),.doutc(w_n801_1[2]),.din(w_n801_0[0]));
	jspl3 jspl3_w_n801_2(.douta(w_n801_2[0]),.doutb(w_n801_2[1]),.doutc(w_n801_2[2]),.din(w_n801_0[1]));
	jspl3 jspl3_w_n801_3(.douta(w_n801_3[0]),.doutb(w_n801_3[1]),.doutc(w_n801_3[2]),.din(w_n801_0[2]));
	jspl jspl_w_n801_4(.douta(w_n801_4[0]),.doutb(w_n801_4[1]),.din(w_n801_1[0]));
	jspl3 jspl3_w_n806_0(.douta(w_n806_0[0]),.doutb(w_n806_0[1]),.doutc(w_n806_0[2]),.din(n806));
	jspl jspl_w_n809_0(.douta(w_n809_0[0]),.doutb(w_n809_0[1]),.din(n809));
	jspl jspl_w_n819_0(.douta(w_n819_0[0]),.doutb(w_n819_0[1]),.din(n819));
	jspl jspl_w_n821_0(.douta(w_n821_0[0]),.doutb(w_n821_0[1]),.din(n821));
	jspl3 jspl3_w_n828_0(.douta(w_n828_0[0]),.doutb(w_dff_A_7jdad2lW2_1),.doutc(w_dff_A_OJIT8lba9_2),.din(n828));
	jspl jspl_w_n829_0(.douta(w_n829_0[0]),.doutb(w_dff_A_FkPSMB6o6_1),.din(n829));
	jspl jspl_w_n832_0(.douta(w_n832_0[0]),.doutb(w_n832_0[1]),.din(n832));
	jspl jspl_w_n839_0(.douta(w_n839_0[0]),.doutb(w_n839_0[1]),.din(n839));
	jspl3 jspl3_w_n840_0(.douta(w_n840_0[0]),.doutb(w_dff_A_UvlIyvVv4_1),.doutc(w_dff_A_r4VlKp9Y2_2),.din(w_dff_B_o0TO8GKR4_3));
	jspl3 jspl3_w_n840_1(.douta(w_n840_1[0]),.doutb(w_dff_A_XrgxLxLA5_1),.doutc(w_dff_A_CkR3Lkis6_2),.din(w_n840_0[0]));
	jspl3 jspl3_w_n840_2(.douta(w_n840_2[0]),.doutb(w_n840_2[1]),.doutc(w_dff_A_Hz1qLP2O7_2),.din(w_n840_0[1]));
	jspl3 jspl3_w_n840_3(.douta(w_n840_3[0]),.doutb(w_dff_A_dRZ0fmRA0_1),.doutc(w_dff_A_oajukjWu6_2),.din(w_n840_0[2]));
	jspl jspl_w_n840_4(.douta(w_dff_A_QcC28Cyj4_0),.doutb(w_n840_4[1]),.din(w_n840_1[0]));
	jspl jspl_w_n842_0(.douta(w_n842_0[0]),.doutb(w_n842_0[1]),.din(n842));
	jspl3 jspl3_w_n843_0(.douta(w_n843_0[0]),.doutb(w_dff_A_EW7Rn3p67_1),.doutc(w_dff_A_bYMz636x6_2),.din(w_dff_B_Yt0cDv956_3));
	jspl3 jspl3_w_n843_1(.douta(w_n843_1[0]),.doutb(w_dff_A_cLm3788F5_1),.doutc(w_dff_A_e0Ih2LcX7_2),.din(w_n843_0[0]));
	jspl3 jspl3_w_n843_2(.douta(w_n843_2[0]),.doutb(w_n843_2[1]),.doutc(w_dff_A_SmbNmyt81_2),.din(w_n843_0[1]));
	jspl3 jspl3_w_n843_3(.douta(w_n843_3[0]),.doutb(w_dff_A_J7Dd7AbO5_1),.doutc(w_dff_A_8OsilrIV3_2),.din(w_n843_0[2]));
	jspl jspl_w_n843_4(.douta(w_dff_A_xlSSDrBy9_0),.doutb(w_n843_4[1]),.din(w_n843_1[0]));
	jspl3 jspl3_w_n845_0(.douta(w_n845_0[0]),.doutb(w_n845_0[1]),.doutc(w_n845_0[2]),.din(n845));
	jspl3 jspl3_w_n845_1(.douta(w_n845_1[0]),.doutb(w_n845_1[1]),.doutc(w_n845_1[2]),.din(w_n845_0[0]));
	jspl3 jspl3_w_n845_2(.douta(w_n845_2[0]),.doutb(w_n845_2[1]),.doutc(w_n845_2[2]),.din(w_n845_0[1]));
	jspl3 jspl3_w_n845_3(.douta(w_n845_3[0]),.doutb(w_n845_3[1]),.doutc(w_n845_3[2]),.din(w_n845_0[2]));
	jspl jspl_w_n845_4(.douta(w_n845_4[0]),.doutb(w_n845_4[1]),.din(w_n845_1[0]));
	jspl3 jspl3_w_n847_0(.douta(w_n847_0[0]),.doutb(w_n847_0[1]),.doutc(w_n847_0[2]),.din(n847));
	jspl3 jspl3_w_n847_1(.douta(w_n847_1[0]),.doutb(w_n847_1[1]),.doutc(w_n847_1[2]),.din(w_n847_0[0]));
	jspl3 jspl3_w_n847_2(.douta(w_n847_2[0]),.doutb(w_n847_2[1]),.doutc(w_n847_2[2]),.din(w_n847_0[1]));
	jspl3 jspl3_w_n847_3(.douta(w_n847_3[0]),.doutb(w_n847_3[1]),.doutc(w_n847_3[2]),.din(w_n847_0[2]));
	jspl jspl_w_n847_4(.douta(w_n847_4[0]),.doutb(w_n847_4[1]),.din(w_n847_1[0]));
	jspl jspl_w_n853_0(.douta(w_n853_0[0]),.doutb(w_dff_A_an92ggBv9_1),.din(w_dff_B_P1SYit4Z8_2));
	jspl jspl_w_n855_0(.douta(w_dff_A_XXL0aiQW4_0),.doutb(w_n855_0[1]),.din(n855));
	jspl jspl_w_n856_0(.douta(w_n856_0[0]),.doutb(w_n856_0[1]),.din(n856));
	jspl jspl_w_n857_0(.douta(w_n857_0[0]),.doutb(w_n857_0[1]),.din(n857));
	jspl jspl_w_n859_0(.douta(w_n859_0[0]),.doutb(w_n859_0[1]),.din(n859));
	jspl jspl_w_n862_0(.douta(w_n862_0[0]),.doutb(w_n862_0[1]),.din(n862));
	jspl jspl_w_n869_0(.douta(w_n869_0[0]),.doutb(w_n869_0[1]),.din(n869));
	jspl jspl_w_n877_0(.douta(w_n877_0[0]),.doutb(w_n877_0[1]),.din(n877));
	jspl jspl_w_n879_0(.douta(w_n879_0[0]),.doutb(w_n879_0[1]),.din(n879));
	jspl jspl_w_n881_0(.douta(w_n881_0[0]),.doutb(w_n881_0[1]),.din(n881));
	jspl jspl_w_n892_0(.douta(w_n892_0[0]),.doutb(w_n892_0[1]),.din(n892));
	jspl jspl_w_n914_0(.douta(w_n914_0[0]),.doutb(w_n914_0[1]),.din(n914));
	jspl jspl_w_n928_0(.douta(w_n928_0[0]),.doutb(w_dff_A_G8ZG0IOT3_1),.din(w_dff_B_r59SndGa8_2));
	jspl3 jspl3_w_n930_0(.douta(w_n930_0[0]),.doutb(w_n930_0[1]),.doutc(w_dff_A_knsfbCJo1_2),.din(w_dff_B_3ijbnRXv9_3));
	jspl jspl_w_n932_0(.douta(w_n932_0[0]),.doutb(w_n932_0[1]),.din(w_dff_B_yjprOUEj0_2));
	jspl3 jspl3_w_n936_0(.douta(w_n936_0[0]),.doutb(w_n936_0[1]),.doutc(w_n936_0[2]),.din(n936));
	jspl jspl_w_n938_0(.douta(w_n938_0[0]),.doutb(w_n938_0[1]),.din(n938));
	jspl jspl_w_n941_0(.douta(w_n941_0[0]),.doutb(w_n941_0[1]),.din(n941));
	jspl jspl_w_n943_0(.douta(w_n943_0[0]),.doutb(w_dff_A_WZBf4SCa2_1),.din(n943));
	jspl jspl_w_n944_0(.douta(w_n944_0[0]),.doutb(w_dff_A_QwGW2V7L3_1),.din(n944));
	jspl jspl_w_n946_0(.douta(w_n946_0[0]),.doutb(w_n946_0[1]),.din(n946));
	jspl3 jspl3_w_n948_0(.douta(w_n948_0[0]),.doutb(w_n948_0[1]),.doutc(w_n948_0[2]),.din(n948));
	jspl jspl_w_n953_0(.douta(w_n953_0[0]),.doutb(w_n953_0[1]),.din(n953));
	jspl jspl_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.din(n954));
	jspl jspl_w_n968_0(.douta(w_n968_0[0]),.doutb(w_dff_A_RjAXddZ37_1),.din(w_dff_B_BywBpOYm8_2));
	jspl jspl_w_n971_0(.douta(w_n971_0[0]),.doutb(w_dff_A_DNotvZS61_1),.din(n971));
	jspl jspl_w_n972_0(.douta(w_n972_0[0]),.doutb(w_n972_0[1]),.din(n972));
	jspl jspl_w_n973_0(.douta(w_n973_0[0]),.doutb(w_n973_0[1]),.din(n973));
	jspl jspl_w_n984_0(.douta(w_n984_0[0]),.doutb(w_n984_0[1]),.din(n984));
	jspl3 jspl3_w_n985_0(.douta(w_n985_0[0]),.doutb(w_dff_A_b0r6wlAP8_1),.doutc(w_dff_A_8kV4NODC1_2),.din(n985));
	jspl3 jspl3_w_n985_1(.douta(w_dff_A_mIXe8xdZ8_0),.doutb(w_n985_1[1]),.doutc(w_dff_A_KvJpBKkq7_2),.din(w_n985_0[0]));
	jspl3 jspl3_w_n985_2(.douta(w_dff_A_tC8auo9X0_0),.doutb(w_dff_A_JLEfot5E1_1),.doutc(w_n985_2[2]),.din(w_n985_0[1]));
	jspl3 jspl3_w_n985_3(.douta(w_dff_A_9ez9Zel48_0),.doutb(w_dff_A_nznAk0ZQ3_1),.doutc(w_n985_3[2]),.din(w_n985_0[2]));
	jspl jspl_w_n985_4(.douta(w_dff_A_uIUJ1IzD8_0),.doutb(w_n985_4[1]),.din(w_n985_1[0]));
	jspl jspl_w_n987_0(.douta(w_n987_0[0]),.doutb(w_n987_0[1]),.din(n987));
	jspl3 jspl3_w_n988_0(.douta(w_n988_0[0]),.doutb(w_dff_A_E0FEgWNI2_1),.doutc(w_dff_A_TM4UFaXR3_2),.din(n988));
	jspl3 jspl3_w_n988_1(.douta(w_dff_A_9hkTMXuv6_0),.doutb(w_n988_1[1]),.doutc(w_dff_A_05E4x0Ju7_2),.din(w_n988_0[0]));
	jspl3 jspl3_w_n988_2(.douta(w_dff_A_kniqA7ph3_0),.doutb(w_dff_A_9abkvoqm3_1),.doutc(w_n988_2[2]),.din(w_n988_0[1]));
	jspl3 jspl3_w_n988_3(.douta(w_dff_A_xOGvZE8S0_0),.doutb(w_dff_A_60Bj9an54_1),.doutc(w_n988_3[2]),.din(w_n988_0[2]));
	jspl jspl_w_n988_4(.douta(w_dff_A_EpbnYmIi7_0),.doutb(w_n988_4[1]),.din(w_n988_1[0]));
	jspl3 jspl3_w_n990_0(.douta(w_n990_0[0]),.doutb(w_n990_0[1]),.doutc(w_n990_0[2]),.din(n990));
	jspl3 jspl3_w_n990_1(.douta(w_n990_1[0]),.doutb(w_n990_1[1]),.doutc(w_n990_1[2]),.din(w_n990_0[0]));
	jspl3 jspl3_w_n990_2(.douta(w_n990_2[0]),.doutb(w_n990_2[1]),.doutc(w_n990_2[2]),.din(w_n990_0[1]));
	jspl3 jspl3_w_n990_3(.douta(w_n990_3[0]),.doutb(w_n990_3[1]),.doutc(w_n990_3[2]),.din(w_n990_0[2]));
	jspl jspl_w_n990_4(.douta(w_n990_4[0]),.doutb(w_n990_4[1]),.din(w_n990_1[0]));
	jspl3 jspl3_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.doutc(w_n992_0[2]),.din(n992));
	jspl3 jspl3_w_n992_1(.douta(w_n992_1[0]),.doutb(w_n992_1[1]),.doutc(w_n992_1[2]),.din(w_n992_0[0]));
	jspl3 jspl3_w_n992_2(.douta(w_n992_2[0]),.doutb(w_n992_2[1]),.doutc(w_n992_2[2]),.din(w_n992_0[1]));
	jspl3 jspl3_w_n992_3(.douta(w_n992_3[0]),.doutb(w_n992_3[1]),.doutc(w_n992_3[2]),.din(w_n992_0[2]));
	jspl jspl_w_n992_4(.douta(w_n992_4[0]),.doutb(w_n992_4[1]),.din(w_n992_1[0]));
	jspl jspl_w_n998_0(.douta(w_n998_0[0]),.doutb(w_n998_0[1]),.din(n998));
	jspl3 jspl3_w_n999_0(.douta(w_n999_0[0]),.doutb(w_dff_A_3K6GrN4X4_1),.doutc(w_dff_A_dahGnmyB9_2),.din(n999));
	jspl3 jspl3_w_n999_1(.douta(w_dff_A_i8oAcA1P3_0),.doutb(w_n999_1[1]),.doutc(w_dff_A_x1eHhxId0_2),.din(w_n999_0[0]));
	jspl3 jspl3_w_n999_2(.douta(w_dff_A_CohO1dF46_0),.doutb(w_dff_A_pvudMBQF0_1),.doutc(w_n999_2[2]),.din(w_n999_0[1]));
	jspl3 jspl3_w_n999_3(.douta(w_dff_A_33UYVb7Q4_0),.doutb(w_dff_A_1nYUCOUx3_1),.doutc(w_n999_3[2]),.din(w_n999_0[2]));
	jspl jspl_w_n999_4(.douta(w_dff_A_HWZNkgDO3_0),.doutb(w_n999_4[1]),.din(w_n999_1[0]));
	jspl jspl_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.din(n1001));
	jspl3 jspl3_w_n1002_0(.douta(w_n1002_0[0]),.doutb(w_dff_A_IJvihPOl2_1),.doutc(w_dff_A_Qs8lUsEQ2_2),.din(n1002));
	jspl3 jspl3_w_n1002_1(.douta(w_dff_A_966KkFoe3_0),.doutb(w_n1002_1[1]),.doutc(w_dff_A_q93wqV3h6_2),.din(w_n1002_0[0]));
	jspl3 jspl3_w_n1002_2(.douta(w_dff_A_rcHSEw7v8_0),.doutb(w_dff_A_BDAlbrwS2_1),.doutc(w_n1002_2[2]),.din(w_n1002_0[1]));
	jspl3 jspl3_w_n1002_3(.douta(w_dff_A_kfhIpUYa8_0),.doutb(w_dff_A_lDdfJqoX7_1),.doutc(w_n1002_3[2]),.din(w_n1002_0[2]));
	jspl jspl_w_n1002_4(.douta(w_dff_A_JvDkBFwb9_0),.doutb(w_n1002_4[1]),.din(w_n1002_1[0]));
	jspl3 jspl3_w_n1004_0(.douta(w_n1004_0[0]),.doutb(w_n1004_0[1]),.doutc(w_n1004_0[2]),.din(n1004));
	jspl3 jspl3_w_n1004_1(.douta(w_n1004_1[0]),.doutb(w_n1004_1[1]),.doutc(w_n1004_1[2]),.din(w_n1004_0[0]));
	jspl3 jspl3_w_n1004_2(.douta(w_n1004_2[0]),.doutb(w_n1004_2[1]),.doutc(w_n1004_2[2]),.din(w_n1004_0[1]));
	jspl3 jspl3_w_n1004_3(.douta(w_n1004_3[0]),.doutb(w_n1004_3[1]),.doutc(w_n1004_3[2]),.din(w_n1004_0[2]));
	jspl jspl_w_n1004_4(.douta(w_n1004_4[0]),.doutb(w_n1004_4[1]),.din(w_n1004_1[0]));
	jspl3 jspl3_w_n1006_0(.douta(w_n1006_0[0]),.doutb(w_n1006_0[1]),.doutc(w_n1006_0[2]),.din(n1006));
	jspl3 jspl3_w_n1006_1(.douta(w_n1006_1[0]),.doutb(w_n1006_1[1]),.doutc(w_n1006_1[2]),.din(w_n1006_0[0]));
	jspl3 jspl3_w_n1006_2(.douta(w_n1006_2[0]),.doutb(w_n1006_2[1]),.doutc(w_n1006_2[2]),.din(w_n1006_0[1]));
	jspl3 jspl3_w_n1006_3(.douta(w_n1006_3[0]),.doutb(w_n1006_3[1]),.doutc(w_n1006_3[2]),.din(w_n1006_0[2]));
	jspl jspl_w_n1006_4(.douta(w_n1006_4[0]),.doutb(w_n1006_4[1]),.din(w_n1006_1[0]));
	jspl3 jspl3_w_n1012_0(.douta(w_n1012_0[0]),.doutb(w_n1012_0[1]),.doutc(w_n1012_0[2]),.din(n1012));
	jspl jspl_w_n1012_1(.douta(w_n1012_1[0]),.doutb(w_n1012_1[1]),.din(w_n1012_0[0]));
	jspl3 jspl3_w_n1014_0(.douta(w_n1014_0[0]),.doutb(w_n1014_0[1]),.doutc(w_n1014_0[2]),.din(n1014));
	jspl jspl_w_n1014_1(.douta(w_n1014_1[0]),.doutb(w_n1014_1[1]),.din(w_n1014_0[0]));
	jspl3 jspl3_w_n1021_0(.douta(w_n1021_0[0]),.doutb(w_n1021_0[1]),.doutc(w_n1021_0[2]),.din(n1021));
	jspl jspl_w_n1021_1(.douta(w_n1021_1[0]),.doutb(w_n1021_1[1]),.din(w_n1021_0[0]));
	jspl3 jspl3_w_n1023_0(.douta(w_n1023_0[0]),.doutb(w_n1023_0[1]),.doutc(w_n1023_0[2]),.din(n1023));
	jspl jspl_w_n1023_1(.douta(w_n1023_1[0]),.doutb(w_n1023_1[1]),.din(w_n1023_0[0]));
	jspl3 jspl3_w_n1030_0(.douta(w_n1030_0[0]),.doutb(w_n1030_0[1]),.doutc(w_n1030_0[2]),.din(n1030));
	jspl jspl_w_n1030_1(.douta(w_n1030_1[0]),.doutb(w_n1030_1[1]),.din(w_n1030_0[0]));
	jspl3 jspl3_w_n1032_0(.douta(w_n1032_0[0]),.doutb(w_n1032_0[1]),.doutc(w_n1032_0[2]),.din(n1032));
	jspl jspl_w_n1032_1(.douta(w_n1032_1[0]),.doutb(w_n1032_1[1]),.din(w_n1032_0[0]));
	jspl3 jspl3_w_n1039_0(.douta(w_n1039_0[0]),.doutb(w_n1039_0[1]),.doutc(w_n1039_0[2]),.din(n1039));
	jspl jspl_w_n1039_1(.douta(w_n1039_1[0]),.doutb(w_n1039_1[1]),.din(w_n1039_0[0]));
	jspl3 jspl3_w_n1041_0(.douta(w_n1041_0[0]),.doutb(w_n1041_0[1]),.doutc(w_n1041_0[2]),.din(n1041));
	jspl jspl_w_n1041_1(.douta(w_n1041_1[0]),.doutb(w_n1041_1[1]),.din(w_n1041_0[0]));
	jspl jspl_w_n1142_0(.douta(w_dff_A_QgDlqxAf5_0),.doutb(w_n1142_0[1]),.din(n1142));
	jspl jspl_w_n1151_0(.douta(w_n1151_0[0]),.doutb(w_n1151_0[1]),.din(n1151));
	jspl3 jspl3_w_n1163_0(.douta(w_n1163_0[0]),.doutb(w_n1163_0[1]),.doutc(w_n1163_0[2]),.din(n1163));
	jspl3 jspl3_w_n1163_1(.douta(w_n1163_1[0]),.doutb(w_n1163_1[1]),.doutc(w_n1163_1[2]),.din(w_n1163_0[0]));
	jspl3 jspl3_w_n1197_0(.douta(w_n1197_0[0]),.doutb(w_n1197_0[1]),.doutc(w_n1197_0[2]),.din(n1197));
	jspl3 jspl3_w_n1197_1(.douta(w_n1197_1[0]),.doutb(w_n1197_1[1]),.doutc(w_n1197_1[2]),.din(w_n1197_0[0]));
	jspl3 jspl3_w_n1205_0(.douta(w_n1205_0[0]),.doutb(w_n1205_0[1]),.doutc(w_n1205_0[2]),.din(n1205));
	jspl3 jspl3_w_n1205_1(.douta(w_n1205_1[0]),.doutb(w_n1205_1[1]),.doutc(w_n1205_1[2]),.din(w_n1205_0[0]));
	jspl3 jspl3_w_n1235_0(.douta(w_n1235_0[0]),.doutb(w_n1235_0[1]),.doutc(w_n1235_0[2]),.din(n1235));
	jspl jspl_w_n1235_1(.douta(w_n1235_1[0]),.doutb(w_n1235_1[1]),.din(w_n1235_0[0]));
	jspl3 jspl3_w_n1242_0(.douta(w_n1242_0[0]),.doutb(w_n1242_0[1]),.doutc(w_n1242_0[2]),.din(n1242));
	jspl jspl_w_n1242_1(.douta(w_n1242_1[0]),.doutb(w_n1242_1[1]),.din(w_n1242_0[0]));
	jspl3 jspl3_w_n1244_0(.douta(w_n1244_0[0]),.doutb(w_n1244_0[1]),.doutc(w_n1244_0[2]),.din(n1244));
	jspl jspl_w_n1244_1(.douta(w_n1244_1[0]),.doutb(w_n1244_1[1]),.din(w_n1244_0[0]));
	jspl3 jspl3_w_n1251_0(.douta(w_n1251_0[0]),.doutb(w_n1251_0[1]),.doutc(w_n1251_0[2]),.din(n1251));
	jspl jspl_w_n1251_1(.douta(w_n1251_1[0]),.doutb(w_n1251_1[1]),.din(w_n1251_0[0]));
	jspl3 jspl3_w_n1253_0(.douta(w_n1253_0[0]),.doutb(w_n1253_0[1]),.doutc(w_n1253_0[2]),.din(n1253));
	jspl jspl_w_n1253_1(.douta(w_n1253_1[0]),.doutb(w_n1253_1[1]),.din(w_n1253_0[0]));
	jspl jspl_w_n1358_0(.douta(w_n1358_0[0]),.doutb(w_n1358_0[1]),.din(n1358));
	jspl jspl_w_n1383_0(.douta(w_dff_A_sN4mtC7W7_0),.doutb(w_n1383_0[1]),.din(n1383));
	jspl jspl_w_n1391_0(.douta(w_dff_A_EZ2RwlKo8_0),.doutb(w_n1391_0[1]),.din(n1391));
	jspl jspl_w_n1394_0(.douta(w_n1394_0[0]),.doutb(w_n1394_0[1]),.din(n1394));
	jspl jspl_w_n1398_0(.douta(w_n1398_0[0]),.doutb(w_n1398_0[1]),.din(n1398));
	jspl jspl_w_n1399_0(.douta(w_n1399_0[0]),.doutb(w_n1399_0[1]),.din(n1399));
	jspl jspl_w_n1409_0(.douta(w_dff_A_nLPM3D7D0_0),.doutb(w_n1409_0[1]),.din(n1409));
	jspl jspl_w_n1410_0(.douta(w_n1410_0[0]),.doutb(w_n1410_0[1]),.din(n1410));
	jspl jspl_w_n1411_0(.douta(w_dff_A_7HpJId9l8_0),.doutb(w_n1411_0[1]),.din(n1411));
	jspl jspl_w_n1421_0(.douta(w_dff_A_XpGcU9sY8_0),.doutb(w_n1421_0[1]),.din(n1421));
	jspl jspl_w_n1425_0(.douta(w_n1425_0[0]),.doutb(w_n1425_0[1]),.din(n1425));
	jspl jspl_w_n1434_0(.douta(w_n1434_0[0]),.doutb(w_n1434_0[1]),.din(n1434));
	jspl jspl_w_n1438_0(.douta(w_n1438_0[0]),.doutb(w_dff_A_oUO70yLF7_1),.din(n1438));
	jspl jspl_w_n1445_0(.douta(w_n1445_0[0]),.doutb(w_n1445_0[1]),.din(n1445));
	jspl jspl_w_n1446_0(.douta(w_n1446_0[0]),.doutb(w_n1446_0[1]),.din(n1446));
	jspl jspl_w_n1447_0(.douta(w_n1447_0[0]),.doutb(w_dff_A_0WWrV3Qm4_1),.din(n1447));
	jspl jspl_w_n1452_0(.douta(w_n1452_0[0]),.doutb(w_n1452_0[1]),.din(n1452));
	jspl jspl_w_n1494_0(.douta(w_n1494_0[0]),.doutb(w_n1494_0[1]),.din(n1494));
	jspl jspl_w_n1533_0(.douta(w_n1533_0[0]),.doutb(w_n1533_0[1]),.din(w_dff_B_8CK6fxJ17_2));
	jspl jspl_w_n1543_0(.douta(w_n1543_0[0]),.doutb(w_n1543_0[1]),.din(w_dff_B_ev8wgKxz4_2));
	jspl jspl_w_n1545_0(.douta(w_n1545_0[0]),.doutb(w_n1545_0[1]),.din(n1545));
	jspl jspl_w_n1553_0(.douta(w_n1553_0[0]),.doutb(w_n1553_0[1]),.din(w_dff_B_g7uquTPI9_2));
	jspl jspl_w_n1555_0(.douta(w_dff_A_qVskqiBq8_0),.doutb(w_n1555_0[1]),.din(n1555));
	jspl jspl_w_n1560_0(.douta(w_n1560_0[0]),.doutb(w_n1560_0[1]),.din(n1560));
	jspl jspl_w_n1568_0(.douta(w_n1568_0[0]),.doutb(w_dff_A_QBOcDrZP2_1),.din(n1568));
	jspl jspl_w_n1591_0(.douta(w_n1591_0[0]),.doutb(w_n1591_0[1]),.din(n1591));
	jspl jspl_w_n1597_0(.douta(w_n1597_0[0]),.doutb(w_n1597_0[1]),.din(n1597));
	jspl3 jspl3_w_n1601_0(.douta(w_n1601_0[0]),.doutb(w_n1601_0[1]),.doutc(w_n1601_0[2]),.din(n1601));
	jspl jspl_w_n1602_0(.douta(w_n1602_0[0]),.doutb(w_n1602_0[1]),.din(n1602));
	jspl jspl_w_n1609_0(.douta(w_n1609_0[0]),.doutb(w_dff_A_iMMMSng30_1),.din(n1609));
	jspl jspl_w_n1610_0(.douta(w_n1610_0[0]),.doutb(w_n1610_0[1]),.din(n1610));
	jspl jspl_w_n1624_0(.douta(w_n1624_0[0]),.doutb(w_n1624_0[1]),.din(w_dff_B_HJ0gmp534_2));
	jspl jspl_w_n1629_0(.douta(w_n1629_0[0]),.doutb(w_n1629_0[1]),.din(n1629));
	jspl jspl_w_n1631_0(.douta(w_n1631_0[0]),.doutb(w_n1631_0[1]),.din(w_dff_B_tg4sOAdy4_2));
	jspl jspl_w_n1634_0(.douta(w_n1634_0[0]),.doutb(w_n1634_0[1]),.din(w_dff_B_Ae5xATey6_2));
	jdff dff_B_jHQBTdJq4_1(.din(G136),.dout(w_dff_B_jHQBTdJq4_1),.clk(gclk));
	jdff dff_B_Anr4sdjm6_0(.din(G2824),.dout(w_dff_B_Anr4sdjm6_0),.clk(gclk));
	jdff dff_B_IMmybuoF8_1(.din(n320),.dout(w_dff_B_IMmybuoF8_1),.clk(gclk));
	jdff dff_B_NU61lJJ87_1(.din(n327),.dout(w_dff_B_NU61lJJ87_1),.clk(gclk));
	jdff dff_B_UXVU0Ypt4_2(.din(n333),.dout(w_dff_B_UXVU0Ypt4_2),.clk(gclk));
	jdff dff_B_gm4p0GP46_1(.din(n338),.dout(w_dff_B_gm4p0GP46_1),.clk(gclk));
	jdff dff_B_623LmuQ12_1(.din(n340),.dout(w_dff_B_623LmuQ12_1),.clk(gclk));
	jdff dff_B_wR4gaxUk6_0(.din(n341),.dout(w_dff_B_wR4gaxUk6_0),.clk(gclk));
	jdff dff_B_vHWIvW9o5_1(.din(G24),.dout(w_dff_B_vHWIvW9o5_1),.clk(gclk));
	jdff dff_B_pHBgUaoW0_1(.din(n345),.dout(w_dff_B_pHBgUaoW0_1),.clk(gclk));
	jdff dff_B_IxahGZvQ1_0(.din(n346),.dout(w_dff_B_IxahGZvQ1_0),.clk(gclk));
	jdff dff_B_vtIH2h1n6_1(.din(G26),.dout(w_dff_B_vtIH2h1n6_1),.clk(gclk));
	jdff dff_A_ttLXDYX95_0(.dout(w_G141_2[0]),.din(w_dff_A_ttLXDYX95_0),.clk(gclk));
	jdff dff_A_biDTaEoA3_0(.dout(w_dff_A_ttLXDYX95_0),.din(w_dff_A_biDTaEoA3_0),.clk(gclk));
	jdff dff_A_YeISUY517_0(.dout(w_dff_A_biDTaEoA3_0),.din(w_dff_A_YeISUY517_0),.clk(gclk));
	jdff dff_A_IMIxIDym3_0(.dout(w_dff_A_YeISUY517_0),.din(w_dff_A_IMIxIDym3_0),.clk(gclk));
	jdff dff_A_f89PYxzO7_1(.dout(w_G141_2[1]),.din(w_dff_A_f89PYxzO7_1),.clk(gclk));
	jdff dff_A_hYDteRYp4_1(.dout(w_dff_A_f89PYxzO7_1),.din(w_dff_A_hYDteRYp4_1),.clk(gclk));
	jdff dff_A_nBSVcUOf5_1(.dout(w_dff_A_hYDteRYp4_1),.din(w_dff_A_nBSVcUOf5_1),.clk(gclk));
	jdff dff_A_Uix9emZd8_1(.dout(w_dff_A_nBSVcUOf5_1),.din(w_dff_A_Uix9emZd8_1),.clk(gclk));
	jdff dff_B_aqsw1dbN5_1(.din(n350),.dout(w_dff_B_aqsw1dbN5_1),.clk(gclk));
	jdff dff_B_DHaR4A7J8_0(.din(n351),.dout(w_dff_B_DHaR4A7J8_0),.clk(gclk));
	jdff dff_B_gnNJIjpj5_1(.din(G79),.dout(w_dff_B_gnNJIjpj5_1),.clk(gclk));
	jdff dff_B_KqiineDQ9_1(.din(n355),.dout(w_dff_B_KqiineDQ9_1),.clk(gclk));
	jdff dff_B_PDQFZ4RW9_0(.din(n356),.dout(w_dff_B_PDQFZ4RW9_0),.clk(gclk));
	jdff dff_B_4YYVXK1V0_1(.din(G82),.dout(w_dff_B_4YYVXK1V0_1),.clk(gclk));
	jdff dff_A_5EOTA0Rs8_0(.dout(w_G2358_2[0]),.din(w_dff_A_5EOTA0Rs8_0),.clk(gclk));
	jdff dff_A_BkHOyTil1_1(.dout(w_G2358_2[1]),.din(w_dff_A_BkHOyTil1_1),.clk(gclk));
	jdff dff_A_yzdqWlka0_1(.dout(w_G141_1[1]),.din(w_dff_A_yzdqWlka0_1),.clk(gclk));
	jdff dff_A_kX2rJmue8_1(.dout(w_dff_A_yzdqWlka0_1),.din(w_dff_A_kX2rJmue8_1),.clk(gclk));
	jdff dff_A_ys9Qfu3j7_1(.dout(w_dff_A_kX2rJmue8_1),.din(w_dff_A_ys9Qfu3j7_1),.clk(gclk));
	jdff dff_A_FVxwN3J96_1(.dout(w_dff_A_ys9Qfu3j7_1),.din(w_dff_A_FVxwN3J96_1),.clk(gclk));
	jdff dff_A_CxbGlPds6_2(.dout(w_G141_1[2]),.din(w_dff_A_CxbGlPds6_2),.clk(gclk));
	jdff dff_A_rAKqKSGo9_2(.dout(w_dff_A_CxbGlPds6_2),.din(w_dff_A_rAKqKSGo9_2),.clk(gclk));
	jdff dff_A_A6FfpvXM3_2(.dout(w_dff_A_rAKqKSGo9_2),.din(w_dff_A_A6FfpvXM3_2),.clk(gclk));
	jdff dff_A_JcqojU074_2(.dout(w_dff_A_A6FfpvXM3_2),.din(w_dff_A_JcqojU074_2),.clk(gclk));
	jdff dff_B_ltj41sKF6_1(.din(n384),.dout(w_dff_B_ltj41sKF6_1),.clk(gclk));
	jdff dff_B_f3ch99Z31_1(.din(w_dff_B_ltj41sKF6_1),.dout(w_dff_B_f3ch99Z31_1),.clk(gclk));
	jdff dff_B_eAqgYHn04_0(.din(n446),.dout(w_dff_B_eAqgYHn04_0),.clk(gclk));
	jdff dff_B_5mlsIGkR7_1(.din(n483),.dout(w_dff_B_5mlsIGkR7_1),.clk(gclk));
	jdff dff_B_uVRcF1Sl0_1(.din(n506),.dout(w_dff_B_uVRcF1Sl0_1),.clk(gclk));
	jdff dff_B_7iy6Kj3D8_2(.din(n652),.dout(w_dff_B_7iy6Kj3D8_2),.clk(gclk));
	jdff dff_B_pPvj2W9G7_2(.din(n709),.dout(w_dff_B_pPvj2W9G7_2),.clk(gclk));
	jdff dff_B_UJrFruSB3_2(.din(w_dff_B_pPvj2W9G7_2),.dout(w_dff_B_UJrFruSB3_2),.clk(gclk));
	jdff dff_B_aRARWFLQ8_2(.din(w_dff_B_UJrFruSB3_2),.dout(w_dff_B_aRARWFLQ8_2),.clk(gclk));
	jdff dff_B_3yN88npG8_1(.din(n698),.dout(w_dff_B_3yN88npG8_1),.clk(gclk));
	jdff dff_B_pEkfxiGf8_1(.din(w_dff_B_3yN88npG8_1),.dout(w_dff_B_pEkfxiGf8_1),.clk(gclk));
	jdff dff_B_SmeA8bAj8_1(.din(w_dff_B_pEkfxiGf8_1),.dout(w_dff_B_SmeA8bAj8_1),.clk(gclk));
	jdff dff_B_pRP80RRX9_1(.din(w_dff_B_SmeA8bAj8_1),.dout(w_dff_B_pRP80RRX9_1),.clk(gclk));
	jdff dff_B_1amRu1IJ8_1(.din(n699),.dout(w_dff_B_1amRu1IJ8_1),.clk(gclk));
	jdff dff_B_Zpe9KJPW8_1(.din(w_dff_B_1amRu1IJ8_1),.dout(w_dff_B_Zpe9KJPW8_1),.clk(gclk));
	jdff dff_B_NZ2J9zDL7_1(.din(w_dff_B_Zpe9KJPW8_1),.dout(w_dff_B_NZ2J9zDL7_1),.clk(gclk));
	jdff dff_A_Xin0Blvm9_1(.dout(w_n607_0[1]),.din(w_dff_A_Xin0Blvm9_1),.clk(gclk));
	jdff dff_A_I5VwRkAh7_1(.dout(w_dff_A_Xin0Blvm9_1),.din(w_dff_A_I5VwRkAh7_1),.clk(gclk));
	jdff dff_B_ZINqSSK07_3(.din(n607),.dout(w_dff_B_ZINqSSK07_3),.clk(gclk));
	jdff dff_B_7Esi7QlS2_3(.din(w_dff_B_ZINqSSK07_3),.dout(w_dff_B_7Esi7QlS2_3),.clk(gclk));
	jdff dff_B_t1QjbpLO5_3(.din(w_dff_B_7Esi7QlS2_3),.dout(w_dff_B_t1QjbpLO5_3),.clk(gclk));
	jdff dff_B_hGOH1ICO8_0(.din(n606),.dout(w_dff_B_hGOH1ICO8_0),.clk(gclk));
	jdff dff_B_8Hj9RYZR3_2(.din(n742),.dout(w_dff_B_8Hj9RYZR3_2),.clk(gclk));
	jdff dff_B_B8YsHfHS2_2(.din(w_dff_B_8Hj9RYZR3_2),.dout(w_dff_B_B8YsHfHS2_2),.clk(gclk));
	jdff dff_B_UDI6drwr2_2(.din(w_dff_B_B8YsHfHS2_2),.dout(w_dff_B_UDI6drwr2_2),.clk(gclk));
	jdff dff_B_ZUBpmoAa7_2(.din(w_dff_B_UDI6drwr2_2),.dout(w_dff_B_ZUBpmoAa7_2),.clk(gclk));
	jdff dff_B_jfeEQVgx4_2(.din(w_dff_B_ZUBpmoAa7_2),.dout(w_dff_B_jfeEQVgx4_2),.clk(gclk));
	jdff dff_A_iJp98zHA5_0(.dout(w_n651_1[0]),.din(w_dff_A_iJp98zHA5_0),.clk(gclk));
	jdff dff_A_LAQ99uND5_0(.dout(w_dff_A_iJp98zHA5_0),.din(w_dff_A_LAQ99uND5_0),.clk(gclk));
	jdff dff_A_b9W3XuLC8_0(.dout(w_dff_A_LAQ99uND5_0),.din(w_dff_A_b9W3XuLC8_0),.clk(gclk));
	jdff dff_A_RNM0zKFw2_0(.dout(w_dff_A_b9W3XuLC8_0),.din(w_dff_A_RNM0zKFw2_0),.clk(gclk));
	jdff dff_A_0kVWVmWh9_0(.dout(w_dff_A_RNM0zKFw2_0),.din(w_dff_A_0kVWVmWh9_0),.clk(gclk));
	jdff dff_A_IG1CENs25_0(.dout(w_dff_A_0kVWVmWh9_0),.din(w_dff_A_IG1CENs25_0),.clk(gclk));
	jdff dff_B_vG7gIifi5_0(.din(n803),.dout(w_dff_B_vG7gIifi5_0),.clk(gclk));
	jdff dff_B_oEWPo6Ko6_0(.din(w_dff_B_vG7gIifi5_0),.dout(w_dff_B_oEWPo6Ko6_0),.clk(gclk));
	jdff dff_B_rwu1TT7A8_0(.din(w_dff_B_oEWPo6Ko6_0),.dout(w_dff_B_rwu1TT7A8_0),.clk(gclk));
	jdff dff_B_nP2d2A7c6_0(.din(w_dff_B_rwu1TT7A8_0),.dout(w_dff_B_nP2d2A7c6_0),.clk(gclk));
	jdff dff_B_jUkZISbW0_0(.din(w_dff_B_nP2d2A7c6_0),.dout(w_dff_B_jUkZISbW0_0),.clk(gclk));
	jdff dff_B_zMkpzVqJ5_0(.din(n802),.dout(w_dff_B_zMkpzVqJ5_0),.clk(gclk));
	jdff dff_B_z7dgp7jw4_0(.din(n849),.dout(w_dff_B_z7dgp7jw4_0),.clk(gclk));
	jdff dff_B_MZks48Sf6_0(.din(w_dff_B_z7dgp7jw4_0),.dout(w_dff_B_MZks48Sf6_0),.clk(gclk));
	jdff dff_B_gg7adqYB2_0(.din(w_dff_B_MZks48Sf6_0),.dout(w_dff_B_gg7adqYB2_0),.clk(gclk));
	jdff dff_B_roUtmP064_0(.din(w_dff_B_gg7adqYB2_0),.dout(w_dff_B_roUtmP064_0),.clk(gclk));
	jdff dff_B_hYePd4Ob5_0(.din(w_dff_B_roUtmP064_0),.dout(w_dff_B_hYePd4Ob5_0),.clk(gclk));
	jdff dff_B_Mt1TyOcg4_0(.din(n848),.dout(w_dff_B_Mt1TyOcg4_0),.clk(gclk));
	jdff dff_B_nWHyNTeU4_2(.din(G61),.dout(w_dff_B_nWHyNTeU4_2),.clk(gclk));
	jdff dff_B_CGOjwWy20_2(.din(G11),.dout(w_dff_B_CGOjwWy20_2),.clk(gclk));
	jdff dff_B_LLUKbs4O8_2(.din(w_dff_B_CGOjwWy20_2),.dout(w_dff_B_LLUKbs4O8_2),.clk(gclk));
	jdff dff_B_HAwExXEz6_0(.din(n964),.dout(w_dff_B_HAwExXEz6_0),.clk(gclk));
	jdff dff_B_UP050EU05_0(.din(n962),.dout(w_dff_B_UP050EU05_0),.clk(gclk));
	jdff dff_B_TVnOlHoq5_0(.din(n961),.dout(w_dff_B_TVnOlHoq5_0),.clk(gclk));
	jdff dff_B_YZtlb9hF8_1(.din(n957),.dout(w_dff_B_YZtlb9hF8_1),.clk(gclk));
	jdff dff_B_w7DtqsC31_1(.din(w_dff_B_YZtlb9hF8_1),.dout(w_dff_B_w7DtqsC31_1),.clk(gclk));
	jdff dff_B_7g3InhJ04_1(.din(w_dff_B_w7DtqsC31_1),.dout(w_dff_B_7g3InhJ04_1),.clk(gclk));
	jdff dff_B_qfGQmnHK9_1(.din(w_dff_B_7g3InhJ04_1),.dout(w_dff_B_qfGQmnHK9_1),.clk(gclk));
	jdff dff_B_4Nihpq5s8_0(.din(n980),.dout(w_dff_B_4Nihpq5s8_0),.clk(gclk));
	jdff dff_B_IJUhH4ns3_0(.din(w_dff_B_4Nihpq5s8_0),.dout(w_dff_B_IJUhH4ns3_0),.clk(gclk));
	jdff dff_B_HrMMq4VJ6_0(.din(n979),.dout(w_dff_B_HrMMq4VJ6_0),.clk(gclk));
	jdff dff_B_KMqjl7ai9_0(.din(n978),.dout(w_dff_B_KMqjl7ai9_0),.clk(gclk));
	jdff dff_B_XrSWrNTy2_0(.din(n977),.dout(w_dff_B_XrSWrNTy2_0),.clk(gclk));
	jdff dff_B_CGVCrTK19_0(.din(n976),.dout(w_dff_B_CGVCrTK19_0),.clk(gclk));
	jdff dff_B_UEhCmxNW0_0(.din(n994),.dout(w_dff_B_UEhCmxNW0_0),.clk(gclk));
	jdff dff_B_uATN87N69_0(.din(w_dff_B_UEhCmxNW0_0),.dout(w_dff_B_uATN87N69_0),.clk(gclk));
	jdff dff_B_ByQQJMxZ3_0(.din(w_dff_B_uATN87N69_0),.dout(w_dff_B_ByQQJMxZ3_0),.clk(gclk));
	jdff dff_B_mZX2pVJF1_0(.din(w_dff_B_ByQQJMxZ3_0),.dout(w_dff_B_mZX2pVJF1_0),.clk(gclk));
	jdff dff_B_X5Rb88TQ7_0(.din(w_dff_B_mZX2pVJF1_0),.dout(w_dff_B_X5Rb88TQ7_0),.clk(gclk));
	jdff dff_B_ryjvrocQ2_0(.din(n993),.dout(w_dff_B_ryjvrocQ2_0),.clk(gclk));
	jdff dff_B_cj0VNEgI1_0(.din(n1008),.dout(w_dff_B_cj0VNEgI1_0),.clk(gclk));
	jdff dff_B_aspS6po80_0(.din(w_dff_B_cj0VNEgI1_0),.dout(w_dff_B_aspS6po80_0),.clk(gclk));
	jdff dff_B_PpZaZXXs6_0(.din(w_dff_B_aspS6po80_0),.dout(w_dff_B_PpZaZXXs6_0),.clk(gclk));
	jdff dff_B_RRch3qeI3_0(.din(w_dff_B_PpZaZXXs6_0),.dout(w_dff_B_RRch3qeI3_0),.clk(gclk));
	jdff dff_B_4EEW3udA8_0(.din(w_dff_B_RRch3qeI3_0),.dout(w_dff_B_4EEW3udA8_0),.clk(gclk));
	jdff dff_B_EbjnnGtL5_0(.din(n1007),.dout(w_dff_B_EbjnnGtL5_0),.clk(gclk));
	jdff dff_B_EftrGcDC3_2(.din(G185),.dout(w_dff_B_EftrGcDC3_2),.clk(gclk));
	jdff dff_B_a96C1oTs3_2(.din(G182),.dout(w_dff_B_a96C1oTs3_2),.clk(gclk));
	jdff dff_B_qds7jQhf3_2(.din(w_dff_B_a96C1oTs3_2),.dout(w_dff_B_qds7jQhf3_2),.clk(gclk));
	jdff dff_B_oJLhhSj89_1(.din(n749),.dout(w_dff_B_oJLhhSj89_1),.clk(gclk));
	jdff dff_B_PFf9ptfD2_0(.din(n754),.dout(w_dff_B_PFf9ptfD2_0),.clk(gclk));
	jdff dff_B_31XDNprI8_1(.din(G131),.dout(w_dff_B_31XDNprI8_1),.clk(gclk));
	jdff dff_B_BOB3AgmJ6_1(.din(w_dff_B_31XDNprI8_1),.dout(w_dff_B_BOB3AgmJ6_1),.clk(gclk));
	jdff dff_B_QO11U0RQ4_0(.din(n776),.dout(w_dff_B_QO11U0RQ4_0),.clk(gclk));
	jdff dff_B_QnR3iPsJ1_0(.din(w_dff_B_QO11U0RQ4_0),.dout(w_dff_B_QnR3iPsJ1_0),.clk(gclk));
	jdff dff_B_RJNpD09T1_1(.din(G117),.dout(w_dff_B_RJNpD09T1_1),.clk(gclk));
	jdff dff_B_pIbDnPuQ1_1(.din(w_dff_B_RJNpD09T1_1),.dout(w_dff_B_pIbDnPuQ1_1),.clk(gclk));
	jdff dff_B_OCIN2bTo6_0(.din(n504),.dout(w_dff_B_OCIN2bTo6_0),.clk(gclk));
	jdff dff_B_jwquK25w5_1(.din(n496),.dout(w_dff_B_jwquK25w5_1),.clk(gclk));
	jdff dff_B_ce2DHmUC9_0(.din(n1019),.dout(w_dff_B_ce2DHmUC9_0),.clk(gclk));
	jdff dff_B_lHQ5ViY04_0(.din(n1018),.dout(w_dff_B_lHQ5ViY04_0),.clk(gclk));
	jdff dff_B_CfaUw6c81_0(.din(w_dff_B_lHQ5ViY04_0),.dout(w_dff_B_CfaUw6c81_0),.clk(gclk));
	jdff dff_B_lpwUEjfF0_0(.din(w_dff_B_CfaUw6c81_0),.dout(w_dff_B_lpwUEjfF0_0),.clk(gclk));
	jdff dff_B_Jt3xcbBB6_0(.din(w_dff_B_lpwUEjfF0_0),.dout(w_dff_B_Jt3xcbBB6_0),.clk(gclk));
	jdff dff_B_1knAGKCk6_0(.din(w_dff_B_Jt3xcbBB6_0),.dout(w_dff_B_1knAGKCk6_0),.clk(gclk));
	jdff dff_B_XrFOhDIu0_0(.din(w_dff_B_1knAGKCk6_0),.dout(w_dff_B_XrFOhDIu0_0),.clk(gclk));
	jdff dff_B_3AsR27S58_0(.din(w_dff_B_XrFOhDIu0_0),.dout(w_dff_B_3AsR27S58_0),.clk(gclk));
	jdff dff_B_orBbCIVg6_0(.din(w_dff_B_3AsR27S58_0),.dout(w_dff_B_orBbCIVg6_0),.clk(gclk));
	jdff dff_B_6LIagr1I1_0(.din(w_dff_B_orBbCIVg6_0),.dout(w_dff_B_6LIagr1I1_0),.clk(gclk));
	jdff dff_B_ZjDAteSM8_0(.din(w_dff_B_6LIagr1I1_0),.dout(w_dff_B_ZjDAteSM8_0),.clk(gclk));
	jdff dff_B_DOJq9JIz6_0(.din(w_dff_B_ZjDAteSM8_0),.dout(w_dff_B_DOJq9JIz6_0),.clk(gclk));
	jdff dff_B_ITRFDaAA8_0(.din(w_dff_B_DOJq9JIz6_0),.dout(w_dff_B_ITRFDaAA8_0),.clk(gclk));
	jdff dff_B_Q0VfgMkX4_0(.din(n1017),.dout(w_dff_B_Q0VfgMkX4_0),.clk(gclk));
	jdff dff_A_0rf7psYY1_0(.dout(w_n797_4[0]),.din(w_dff_A_0rf7psYY1_0),.clk(gclk));
	jdff dff_A_AW4savrb3_0(.dout(w_dff_A_0rf7psYY1_0),.din(w_dff_A_AW4savrb3_0),.clk(gclk));
	jdff dff_A_gkNdMhPI6_0(.dout(w_dff_A_AW4savrb3_0),.din(w_dff_A_gkNdMhPI6_0),.clk(gclk));
	jdff dff_A_vj2YgRVs5_0(.dout(w_dff_A_gkNdMhPI6_0),.din(w_dff_A_vj2YgRVs5_0),.clk(gclk));
	jdff dff_A_RN1eUI9Y0_0(.dout(w_dff_A_vj2YgRVs5_0),.din(w_dff_A_RN1eUI9Y0_0),.clk(gclk));
	jdff dff_A_ACvQgDkR0_0(.dout(w_dff_A_RN1eUI9Y0_0),.din(w_dff_A_ACvQgDkR0_0),.clk(gclk));
	jdff dff_A_yGyRJSXA9_0(.dout(w_dff_A_ACvQgDkR0_0),.din(w_dff_A_yGyRJSXA9_0),.clk(gclk));
	jdff dff_A_trJ3JV1b3_0(.dout(w_n793_4[0]),.din(w_dff_A_trJ3JV1b3_0),.clk(gclk));
	jdff dff_A_TaAECb3k8_0(.dout(w_dff_A_trJ3JV1b3_0),.din(w_dff_A_TaAECb3k8_0),.clk(gclk));
	jdff dff_A_JmnIQOFK1_0(.dout(w_dff_A_TaAECb3k8_0),.din(w_dff_A_JmnIQOFK1_0),.clk(gclk));
	jdff dff_A_Ypf1M73J5_0(.dout(w_dff_A_JmnIQOFK1_0),.din(w_dff_A_Ypf1M73J5_0),.clk(gclk));
	jdff dff_A_cLKTDLD97_0(.dout(w_dff_A_Ypf1M73J5_0),.din(w_dff_A_cLKTDLD97_0),.clk(gclk));
	jdff dff_A_vq5XQZJv8_0(.dout(w_dff_A_cLKTDLD97_0),.din(w_dff_A_vq5XQZJv8_0),.clk(gclk));
	jdff dff_A_bCGTqDzo5_0(.dout(w_dff_A_vq5XQZJv8_0),.din(w_dff_A_bCGTqDzo5_0),.clk(gclk));
	jdff dff_A_zKo6lCdE9_0(.dout(w_dff_A_bCGTqDzo5_0),.din(w_dff_A_zKo6lCdE9_0),.clk(gclk));
	jdff dff_B_plgG2qC08_0(.din(n1028),.dout(w_dff_B_plgG2qC08_0),.clk(gclk));
	jdff dff_B_m3Rr661J6_0(.din(n1027),.dout(w_dff_B_m3Rr661J6_0),.clk(gclk));
	jdff dff_B_9Z7rjXjx7_0(.din(w_dff_B_m3Rr661J6_0),.dout(w_dff_B_9Z7rjXjx7_0),.clk(gclk));
	jdff dff_B_6IdFPoG57_0(.din(w_dff_B_9Z7rjXjx7_0),.dout(w_dff_B_6IdFPoG57_0),.clk(gclk));
	jdff dff_B_OYphEQiZ5_0(.din(w_dff_B_6IdFPoG57_0),.dout(w_dff_B_OYphEQiZ5_0),.clk(gclk));
	jdff dff_B_3zQhCRk18_0(.din(w_dff_B_OYphEQiZ5_0),.dout(w_dff_B_3zQhCRk18_0),.clk(gclk));
	jdff dff_B_hMqcxCjY6_0(.din(w_dff_B_3zQhCRk18_0),.dout(w_dff_B_hMqcxCjY6_0),.clk(gclk));
	jdff dff_B_X4zi9jxB5_0(.din(w_dff_B_hMqcxCjY6_0),.dout(w_dff_B_X4zi9jxB5_0),.clk(gclk));
	jdff dff_B_RhiIaZXb6_0(.din(w_dff_B_X4zi9jxB5_0),.dout(w_dff_B_RhiIaZXb6_0),.clk(gclk));
	jdff dff_B_K9Mfqw101_0(.din(w_dff_B_RhiIaZXb6_0),.dout(w_dff_B_K9Mfqw101_0),.clk(gclk));
	jdff dff_B_SBR2JHGD2_0(.din(w_dff_B_K9Mfqw101_0),.dout(w_dff_B_SBR2JHGD2_0),.clk(gclk));
	jdff dff_B_yJdSPpJm7_0(.din(n1026),.dout(w_dff_B_yJdSPpJm7_0),.clk(gclk));
	jdff dff_B_vUQkrHzj0_0(.din(n1037),.dout(w_dff_B_vUQkrHzj0_0),.clk(gclk));
	jdff dff_B_LN2JCHDe2_0(.din(w_dff_B_vUQkrHzj0_0),.dout(w_dff_B_LN2JCHDe2_0),.clk(gclk));
	jdff dff_B_u22uWexP5_0(.din(n1036),.dout(w_dff_B_u22uWexP5_0),.clk(gclk));
	jdff dff_B_nHTc1oyJ6_0(.din(w_dff_B_u22uWexP5_0),.dout(w_dff_B_nHTc1oyJ6_0),.clk(gclk));
	jdff dff_B_rS1GjpzH9_0(.din(w_dff_B_nHTc1oyJ6_0),.dout(w_dff_B_rS1GjpzH9_0),.clk(gclk));
	jdff dff_B_ZBJWExEA4_0(.din(w_dff_B_rS1GjpzH9_0),.dout(w_dff_B_ZBJWExEA4_0),.clk(gclk));
	jdff dff_B_zX6Zn8ZF2_0(.din(w_dff_B_ZBJWExEA4_0),.dout(w_dff_B_zX6Zn8ZF2_0),.clk(gclk));
	jdff dff_B_lWqwbSZy1_0(.din(w_dff_B_zX6Zn8ZF2_0),.dout(w_dff_B_lWqwbSZy1_0),.clk(gclk));
	jdff dff_B_yH1IjA8i5_0(.din(w_dff_B_lWqwbSZy1_0),.dout(w_dff_B_yH1IjA8i5_0),.clk(gclk));
	jdff dff_B_b1Bo3pNX3_0(.din(w_dff_B_yH1IjA8i5_0),.dout(w_dff_B_b1Bo3pNX3_0),.clk(gclk));
	jdff dff_B_FTDf6ngq6_0(.din(n1035),.dout(w_dff_B_FTDf6ngq6_0),.clk(gclk));
	jdff dff_B_mNjZmzVF3_0(.din(n1046),.dout(w_dff_B_mNjZmzVF3_0),.clk(gclk));
	jdff dff_B_0jpKrJJW7_0(.din(w_dff_B_mNjZmzVF3_0),.dout(w_dff_B_0jpKrJJW7_0),.clk(gclk));
	jdff dff_B_yvilTlyr0_0(.din(w_dff_B_0jpKrJJW7_0),.dout(w_dff_B_yvilTlyr0_0),.clk(gclk));
	jdff dff_B_sIGWFB6b0_0(.din(n1045),.dout(w_dff_B_sIGWFB6b0_0),.clk(gclk));
	jdff dff_B_3ksMGvfV8_0(.din(w_dff_B_sIGWFB6b0_0),.dout(w_dff_B_3ksMGvfV8_0),.clk(gclk));
	jdff dff_B_xJJ6kDRm3_0(.din(w_dff_B_3ksMGvfV8_0),.dout(w_dff_B_xJJ6kDRm3_0),.clk(gclk));
	jdff dff_B_PDhjoWO68_0(.din(w_dff_B_xJJ6kDRm3_0),.dout(w_dff_B_PDhjoWO68_0),.clk(gclk));
	jdff dff_B_vnKuuCMV3_0(.din(w_dff_B_PDhjoWO68_0),.dout(w_dff_B_vnKuuCMV3_0),.clk(gclk));
	jdff dff_B_vpAFIKRV2_0(.din(w_dff_B_vnKuuCMV3_0),.dout(w_dff_B_vpAFIKRV2_0),.clk(gclk));
	jdff dff_B_d4K1Bo386_0(.din(n1044),.dout(w_dff_B_d4K1Bo386_0),.clk(gclk));
	jdff dff_A_7JrfLBXL2_1(.dout(w_n797_3[1]),.din(w_dff_A_7JrfLBXL2_1),.clk(gclk));
	jdff dff_A_RzFTeu7T9_1(.dout(w_dff_A_7JrfLBXL2_1),.din(w_dff_A_RzFTeu7T9_1),.clk(gclk));
	jdff dff_A_85wekFvO6_2(.dout(w_n797_3[2]),.din(w_dff_A_85wekFvO6_2),.clk(gclk));
	jdff dff_A_qLmNRbxh1_2(.dout(w_dff_A_85wekFvO6_2),.din(w_dff_A_qLmNRbxh1_2),.clk(gclk));
	jdff dff_A_76Z9Oaut4_2(.dout(w_dff_A_qLmNRbxh1_2),.din(w_dff_A_76Z9Oaut4_2),.clk(gclk));
	jdff dff_A_ryKJwIR74_2(.dout(w_dff_A_76Z9Oaut4_2),.din(w_dff_A_ryKJwIR74_2),.clk(gclk));
	jdff dff_A_cyhATo4q5_1(.dout(w_n793_3[1]),.din(w_dff_A_cyhATo4q5_1),.clk(gclk));
	jdff dff_A_wxcAGRZI2_2(.dout(w_n793_3[2]),.din(w_dff_A_wxcAGRZI2_2),.clk(gclk));
	jdff dff_A_Z3YaYsW56_2(.dout(w_dff_A_wxcAGRZI2_2),.din(w_dff_A_Z3YaYsW56_2),.clk(gclk));
	jdff dff_B_x28AR9oc9_0(.din(n1053),.dout(w_dff_B_x28AR9oc9_0),.clk(gclk));
	jdff dff_B_LaWn1N7U4_0(.din(n1052),.dout(w_dff_B_LaWn1N7U4_0),.clk(gclk));
	jdff dff_B_ZrmOjU6m7_0(.din(w_dff_B_LaWn1N7U4_0),.dout(w_dff_B_ZrmOjU6m7_0),.clk(gclk));
	jdff dff_B_loOHNNpY6_0(.din(w_dff_B_ZrmOjU6m7_0),.dout(w_dff_B_loOHNNpY6_0),.clk(gclk));
	jdff dff_B_ROeYGZA83_0(.din(w_dff_B_loOHNNpY6_0),.dout(w_dff_B_ROeYGZA83_0),.clk(gclk));
	jdff dff_B_HqruB29x5_0(.din(w_dff_B_ROeYGZA83_0),.dout(w_dff_B_HqruB29x5_0),.clk(gclk));
	jdff dff_B_f3GWPNL62_0(.din(w_dff_B_HqruB29x5_0),.dout(w_dff_B_f3GWPNL62_0),.clk(gclk));
	jdff dff_B_p4vcI9nz8_0(.din(w_dff_B_f3GWPNL62_0),.dout(w_dff_B_p4vcI9nz8_0),.clk(gclk));
	jdff dff_B_H8zwpshB5_0(.din(w_dff_B_p4vcI9nz8_0),.dout(w_dff_B_H8zwpshB5_0),.clk(gclk));
	jdff dff_B_tzFAyP2l8_0(.din(w_dff_B_H8zwpshB5_0),.dout(w_dff_B_tzFAyP2l8_0),.clk(gclk));
	jdff dff_B_sGlEKDiE9_0(.din(w_dff_B_tzFAyP2l8_0),.dout(w_dff_B_sGlEKDiE9_0),.clk(gclk));
	jdff dff_B_aUQ55GmA8_0(.din(w_dff_B_sGlEKDiE9_0),.dout(w_dff_B_aUQ55GmA8_0),.clk(gclk));
	jdff dff_B_1rrl11Yh9_0(.din(w_dff_B_aUQ55GmA8_0),.dout(w_dff_B_1rrl11Yh9_0),.clk(gclk));
	jdff dff_B_9M5xc7r91_0(.din(n1051),.dout(w_dff_B_9M5xc7r91_0),.clk(gclk));
	jdff dff_B_IvRLvBDD0_2(.din(G37),.dout(w_dff_B_IvRLvBDD0_2),.clk(gclk));
	jdff dff_B_7tPDAO0p0_2(.din(G43),.dout(w_dff_B_7tPDAO0p0_2),.clk(gclk));
	jdff dff_B_aMcOYz5D7_2(.din(w_dff_B_7tPDAO0p0_2),.dout(w_dff_B_aMcOYz5D7_2),.clk(gclk));
	jdff dff_A_nRNZJ5p44_0(.dout(w_n843_4[0]),.din(w_dff_A_nRNZJ5p44_0),.clk(gclk));
	jdff dff_A_ExQoIyrZ9_0(.dout(w_dff_A_nRNZJ5p44_0),.din(w_dff_A_ExQoIyrZ9_0),.clk(gclk));
	jdff dff_A_INilhmeI0_0(.dout(w_dff_A_ExQoIyrZ9_0),.din(w_dff_A_INilhmeI0_0),.clk(gclk));
	jdff dff_A_AbgE24Bn4_0(.dout(w_dff_A_INilhmeI0_0),.din(w_dff_A_AbgE24Bn4_0),.clk(gclk));
	jdff dff_A_Vpfju6Nd8_0(.dout(w_dff_A_AbgE24Bn4_0),.din(w_dff_A_Vpfju6Nd8_0),.clk(gclk));
	jdff dff_A_1Eq9JByu5_0(.dout(w_dff_A_Vpfju6Nd8_0),.din(w_dff_A_1Eq9JByu5_0),.clk(gclk));
	jdff dff_A_xlSSDrBy9_0(.dout(w_dff_A_1Eq9JByu5_0),.din(w_dff_A_xlSSDrBy9_0),.clk(gclk));
	jdff dff_A_hfEVaF540_0(.dout(w_n840_4[0]),.din(w_dff_A_hfEVaF540_0),.clk(gclk));
	jdff dff_A_iNpUN3Wl3_0(.dout(w_dff_A_hfEVaF540_0),.din(w_dff_A_iNpUN3Wl3_0),.clk(gclk));
	jdff dff_A_ESEnQAr29_0(.dout(w_dff_A_iNpUN3Wl3_0),.din(w_dff_A_ESEnQAr29_0),.clk(gclk));
	jdff dff_A_ePefduiP3_0(.dout(w_dff_A_ESEnQAr29_0),.din(w_dff_A_ePefduiP3_0),.clk(gclk));
	jdff dff_A_6aeXJ5yw8_0(.dout(w_dff_A_ePefduiP3_0),.din(w_dff_A_6aeXJ5yw8_0),.clk(gclk));
	jdff dff_A_fdUw5kI28_0(.dout(w_dff_A_6aeXJ5yw8_0),.din(w_dff_A_fdUw5kI28_0),.clk(gclk));
	jdff dff_A_NWVKWA597_0(.dout(w_dff_A_fdUw5kI28_0),.din(w_dff_A_NWVKWA597_0),.clk(gclk));
	jdff dff_A_QcC28Cyj4_0(.dout(w_dff_A_NWVKWA597_0),.din(w_dff_A_QcC28Cyj4_0),.clk(gclk));
	jdff dff_B_mytJ3CSB9_0(.din(n1060),.dout(w_dff_B_mytJ3CSB9_0),.clk(gclk));
	jdff dff_B_STI7cpBA1_0(.din(n1059),.dout(w_dff_B_STI7cpBA1_0),.clk(gclk));
	jdff dff_B_craCbSdK1_0(.din(w_dff_B_STI7cpBA1_0),.dout(w_dff_B_craCbSdK1_0),.clk(gclk));
	jdff dff_B_C4JaHRpC0_0(.din(w_dff_B_craCbSdK1_0),.dout(w_dff_B_C4JaHRpC0_0),.clk(gclk));
	jdff dff_B_6QMXdnGr6_0(.din(w_dff_B_C4JaHRpC0_0),.dout(w_dff_B_6QMXdnGr6_0),.clk(gclk));
	jdff dff_B_2HZQdbdX4_0(.din(w_dff_B_6QMXdnGr6_0),.dout(w_dff_B_2HZQdbdX4_0),.clk(gclk));
	jdff dff_B_PU0Xr1cP7_0(.din(w_dff_B_2HZQdbdX4_0),.dout(w_dff_B_PU0Xr1cP7_0),.clk(gclk));
	jdff dff_B_TSbbCI2R9_0(.din(w_dff_B_PU0Xr1cP7_0),.dout(w_dff_B_TSbbCI2R9_0),.clk(gclk));
	jdff dff_B_QZ7gkqiz8_0(.din(w_dff_B_TSbbCI2R9_0),.dout(w_dff_B_QZ7gkqiz8_0),.clk(gclk));
	jdff dff_B_OBjHl8bY0_0(.din(w_dff_B_QZ7gkqiz8_0),.dout(w_dff_B_OBjHl8bY0_0),.clk(gclk));
	jdff dff_B_cfNDjJPe0_0(.din(w_dff_B_OBjHl8bY0_0),.dout(w_dff_B_cfNDjJPe0_0),.clk(gclk));
	jdff dff_B_4YYQYK7A9_0(.din(n1058),.dout(w_dff_B_4YYQYK7A9_0),.clk(gclk));
	jdff dff_B_u64XRs6s1_2(.din(G20),.dout(w_dff_B_u64XRs6s1_2),.clk(gclk));
	jdff dff_B_fRvmqErS7_2(.din(G76),.dout(w_dff_B_fRvmqErS7_2),.clk(gclk));
	jdff dff_B_XzoOlpDi0_2(.din(w_dff_B_fRvmqErS7_2),.dout(w_dff_B_XzoOlpDi0_2),.clk(gclk));
	jdff dff_B_iROGU24a0_0(.din(n1067),.dout(w_dff_B_iROGU24a0_0),.clk(gclk));
	jdff dff_B_GrUuGhbS2_0(.din(w_dff_B_iROGU24a0_0),.dout(w_dff_B_GrUuGhbS2_0),.clk(gclk));
	jdff dff_B_RN01pbPJ3_0(.din(n1066),.dout(w_dff_B_RN01pbPJ3_0),.clk(gclk));
	jdff dff_B_VgKMD2p48_0(.din(w_dff_B_RN01pbPJ3_0),.dout(w_dff_B_VgKMD2p48_0),.clk(gclk));
	jdff dff_B_wSU9UURo8_0(.din(w_dff_B_VgKMD2p48_0),.dout(w_dff_B_wSU9UURo8_0),.clk(gclk));
	jdff dff_B_eeh6DvYa5_0(.din(w_dff_B_wSU9UURo8_0),.dout(w_dff_B_eeh6DvYa5_0),.clk(gclk));
	jdff dff_B_TBZmTWlY8_0(.din(w_dff_B_eeh6DvYa5_0),.dout(w_dff_B_TBZmTWlY8_0),.clk(gclk));
	jdff dff_B_EWjObTSD2_0(.din(w_dff_B_TBZmTWlY8_0),.dout(w_dff_B_EWjObTSD2_0),.clk(gclk));
	jdff dff_B_5wCpzg9F2_0(.din(w_dff_B_EWjObTSD2_0),.dout(w_dff_B_5wCpzg9F2_0),.clk(gclk));
	jdff dff_B_v63e2pER8_0(.din(w_dff_B_5wCpzg9F2_0),.dout(w_dff_B_v63e2pER8_0),.clk(gclk));
	jdff dff_B_pwMPdJHW0_0(.din(n1065),.dout(w_dff_B_pwMPdJHW0_0),.clk(gclk));
	jdff dff_B_e6C6fCKi5_2(.din(G17),.dout(w_dff_B_e6C6fCKi5_2),.clk(gclk));
	jdff dff_B_gF9J4mhZ7_2(.din(G73),.dout(w_dff_B_gF9J4mhZ7_2),.clk(gclk));
	jdff dff_B_cUq7hYYo7_2(.din(w_dff_B_gF9J4mhZ7_2),.dout(w_dff_B_cUq7hYYo7_2),.clk(gclk));
	jdff dff_B_U01SPKza4_0(.din(n1074),.dout(w_dff_B_U01SPKza4_0),.clk(gclk));
	jdff dff_B_HNulD6EV5_0(.din(w_dff_B_U01SPKza4_0),.dout(w_dff_B_HNulD6EV5_0),.clk(gclk));
	jdff dff_B_pIpn7ApU6_0(.din(w_dff_B_HNulD6EV5_0),.dout(w_dff_B_pIpn7ApU6_0),.clk(gclk));
	jdff dff_B_HBzwF5yD2_0(.din(n1073),.dout(w_dff_B_HBzwF5yD2_0),.clk(gclk));
	jdff dff_B_hGLN6FZ34_0(.din(w_dff_B_HBzwF5yD2_0),.dout(w_dff_B_hGLN6FZ34_0),.clk(gclk));
	jdff dff_B_GC3UT7hB7_0(.din(w_dff_B_hGLN6FZ34_0),.dout(w_dff_B_GC3UT7hB7_0),.clk(gclk));
	jdff dff_B_TiArMLyD8_0(.din(w_dff_B_GC3UT7hB7_0),.dout(w_dff_B_TiArMLyD8_0),.clk(gclk));
	jdff dff_B_Kz42r3AX1_0(.din(w_dff_B_TiArMLyD8_0),.dout(w_dff_B_Kz42r3AX1_0),.clk(gclk));
	jdff dff_B_YZqsccn93_0(.din(w_dff_B_Kz42r3AX1_0),.dout(w_dff_B_YZqsccn93_0),.clk(gclk));
	jdff dff_B_4tTd2lKx5_0(.din(n1072),.dout(w_dff_B_4tTd2lKx5_0),.clk(gclk));
	jdff dff_B_9xJiJbm46_2(.din(G70),.dout(w_dff_B_9xJiJbm46_2),.clk(gclk));
	jdff dff_B_d0nNtj9g6_2(.din(G67),.dout(w_dff_B_d0nNtj9g6_2),.clk(gclk));
	jdff dff_B_PKSteptA6_2(.din(w_dff_B_d0nNtj9g6_2),.dout(w_dff_B_PKSteptA6_2),.clk(gclk));
	jdff dff_A_32xajYbh3_1(.dout(w_n843_3[1]),.din(w_dff_A_32xajYbh3_1),.clk(gclk));
	jdff dff_A_J7Dd7AbO5_1(.dout(w_dff_A_32xajYbh3_1),.din(w_dff_A_J7Dd7AbO5_1),.clk(gclk));
	jdff dff_A_eoTcwGK65_2(.dout(w_n843_3[2]),.din(w_dff_A_eoTcwGK65_2),.clk(gclk));
	jdff dff_A_gYXcvBaG9_2(.dout(w_dff_A_eoTcwGK65_2),.din(w_dff_A_gYXcvBaG9_2),.clk(gclk));
	jdff dff_A_vflnmgKr7_2(.dout(w_dff_A_gYXcvBaG9_2),.din(w_dff_A_vflnmgKr7_2),.clk(gclk));
	jdff dff_A_8OsilrIV3_2(.dout(w_dff_A_vflnmgKr7_2),.din(w_dff_A_8OsilrIV3_2),.clk(gclk));
	jdff dff_A_dRZ0fmRA0_1(.dout(w_n840_3[1]),.din(w_dff_A_dRZ0fmRA0_1),.clk(gclk));
	jdff dff_A_Ye90dm7A3_2(.dout(w_n840_3[2]),.din(w_dff_A_Ye90dm7A3_2),.clk(gclk));
	jdff dff_A_oajukjWu6_2(.dout(w_dff_A_Ye90dm7A3_2),.din(w_dff_A_oajukjWu6_2),.clk(gclk));
	jdff dff_B_i4lPnUWI4_0(.din(n1081),.dout(w_dff_B_i4lPnUWI4_0),.clk(gclk));
	jdff dff_B_eYCPyy3l6_0(.din(n1080),.dout(w_dff_B_eYCPyy3l6_0),.clk(gclk));
	jdff dff_B_NQvq1k092_0(.din(w_dff_B_eYCPyy3l6_0),.dout(w_dff_B_NQvq1k092_0),.clk(gclk));
	jdff dff_B_JvAyIygj0_0(.din(w_dff_B_NQvq1k092_0),.dout(w_dff_B_JvAyIygj0_0),.clk(gclk));
	jdff dff_B_sAN1nCmR0_0(.din(w_dff_B_JvAyIygj0_0),.dout(w_dff_B_sAN1nCmR0_0),.clk(gclk));
	jdff dff_B_3cwXepcK3_0(.din(w_dff_B_sAN1nCmR0_0),.dout(w_dff_B_3cwXepcK3_0),.clk(gclk));
	jdff dff_B_J6ocffbi6_0(.din(w_dff_B_3cwXepcK3_0),.dout(w_dff_B_J6ocffbi6_0),.clk(gclk));
	jdff dff_B_R98uW9kW2_0(.din(w_dff_B_J6ocffbi6_0),.dout(w_dff_B_R98uW9kW2_0),.clk(gclk));
	jdff dff_B_LsWCv4p96_0(.din(w_dff_B_R98uW9kW2_0),.dout(w_dff_B_LsWCv4p96_0),.clk(gclk));
	jdff dff_B_qfU9wApL3_0(.din(w_dff_B_LsWCv4p96_0),.dout(w_dff_B_qfU9wApL3_0),.clk(gclk));
	jdff dff_B_b48h3PoD0_0(.din(w_dff_B_qfU9wApL3_0),.dout(w_dff_B_b48h3PoD0_0),.clk(gclk));
	jdff dff_B_kCdUc63p2_0(.din(w_dff_B_b48h3PoD0_0),.dout(w_dff_B_kCdUc63p2_0),.clk(gclk));
	jdff dff_B_NZAe3sJK5_0(.din(w_dff_B_kCdUc63p2_0),.dout(w_dff_B_NZAe3sJK5_0),.clk(gclk));
	jdff dff_B_Rge1IOJ90_0(.din(n1079),.dout(w_dff_B_Rge1IOJ90_0),.clk(gclk));
	jdff dff_A_EjGxEXaG5_0(.dout(w_n988_4[0]),.din(w_dff_A_EjGxEXaG5_0),.clk(gclk));
	jdff dff_A_Nkrkw3fs8_0(.dout(w_dff_A_EjGxEXaG5_0),.din(w_dff_A_Nkrkw3fs8_0),.clk(gclk));
	jdff dff_A_t2RnZ8zQ1_0(.dout(w_dff_A_Nkrkw3fs8_0),.din(w_dff_A_t2RnZ8zQ1_0),.clk(gclk));
	jdff dff_A_75LsJQEN2_0(.dout(w_dff_A_t2RnZ8zQ1_0),.din(w_dff_A_75LsJQEN2_0),.clk(gclk));
	jdff dff_A_cYHaD0Dj2_0(.dout(w_dff_A_75LsJQEN2_0),.din(w_dff_A_cYHaD0Dj2_0),.clk(gclk));
	jdff dff_A_gQgyRyRP6_0(.dout(w_dff_A_cYHaD0Dj2_0),.din(w_dff_A_gQgyRyRP6_0),.clk(gclk));
	jdff dff_A_EpbnYmIi7_0(.dout(w_dff_A_gQgyRyRP6_0),.din(w_dff_A_EpbnYmIi7_0),.clk(gclk));
	jdff dff_A_jIUiAxKc8_0(.dout(w_n985_4[0]),.din(w_dff_A_jIUiAxKc8_0),.clk(gclk));
	jdff dff_A_GVHxFxes7_0(.dout(w_dff_A_jIUiAxKc8_0),.din(w_dff_A_GVHxFxes7_0),.clk(gclk));
	jdff dff_A_Z2SXCxO75_0(.dout(w_dff_A_GVHxFxes7_0),.din(w_dff_A_Z2SXCxO75_0),.clk(gclk));
	jdff dff_A_G6LaeZFv6_0(.dout(w_dff_A_Z2SXCxO75_0),.din(w_dff_A_G6LaeZFv6_0),.clk(gclk));
	jdff dff_A_4slQe8Pt6_0(.dout(w_dff_A_G6LaeZFv6_0),.din(w_dff_A_4slQe8Pt6_0),.clk(gclk));
	jdff dff_A_DdZU23Bq4_0(.dout(w_dff_A_4slQe8Pt6_0),.din(w_dff_A_DdZU23Bq4_0),.clk(gclk));
	jdff dff_A_ew1ezB1N1_0(.dout(w_dff_A_DdZU23Bq4_0),.din(w_dff_A_ew1ezB1N1_0),.clk(gclk));
	jdff dff_A_uIUJ1IzD8_0(.dout(w_dff_A_ew1ezB1N1_0),.din(w_dff_A_uIUJ1IzD8_0),.clk(gclk));
	jdff dff_B_2Pb3NNG52_0(.din(n1089),.dout(w_dff_B_2Pb3NNG52_0),.clk(gclk));
	jdff dff_B_FMadaEYd7_0(.din(w_dff_B_2Pb3NNG52_0),.dout(w_dff_B_FMadaEYd7_0),.clk(gclk));
	jdff dff_B_1H19wOa74_0(.din(w_dff_B_FMadaEYd7_0),.dout(w_dff_B_1H19wOa74_0),.clk(gclk));
	jdff dff_B_hYM7vp0g1_0(.din(n1088),.dout(w_dff_B_hYM7vp0g1_0),.clk(gclk));
	jdff dff_B_7KwvDgKt5_0(.din(w_dff_B_hYM7vp0g1_0),.dout(w_dff_B_7KwvDgKt5_0),.clk(gclk));
	jdff dff_B_l66hWUEN6_0(.din(w_dff_B_7KwvDgKt5_0),.dout(w_dff_B_l66hWUEN6_0),.clk(gclk));
	jdff dff_B_3cejkBvY1_0(.din(w_dff_B_l66hWUEN6_0),.dout(w_dff_B_3cejkBvY1_0),.clk(gclk));
	jdff dff_B_0G81fxKi8_0(.din(w_dff_B_3cejkBvY1_0),.dout(w_dff_B_0G81fxKi8_0),.clk(gclk));
	jdff dff_B_jFd1qzXD8_0(.din(w_dff_B_0G81fxKi8_0),.dout(w_dff_B_jFd1qzXD8_0),.clk(gclk));
	jdff dff_B_KuXXw29b6_0(.din(n1087),.dout(w_dff_B_KuXXw29b6_0),.clk(gclk));
	jdff dff_B_4ZNA6fgK6_0(.din(n1097),.dout(w_dff_B_4ZNA6fgK6_0),.clk(gclk));
	jdff dff_B_aVoZ8Ga37_0(.din(w_dff_B_4ZNA6fgK6_0),.dout(w_dff_B_aVoZ8Ga37_0),.clk(gclk));
	jdff dff_B_pF19CPtU6_0(.din(n1096),.dout(w_dff_B_pF19CPtU6_0),.clk(gclk));
	jdff dff_B_ViHDmc1t2_0(.din(w_dff_B_pF19CPtU6_0),.dout(w_dff_B_ViHDmc1t2_0),.clk(gclk));
	jdff dff_B_hMZc7jZp0_0(.din(w_dff_B_ViHDmc1t2_0),.dout(w_dff_B_hMZc7jZp0_0),.clk(gclk));
	jdff dff_B_uVxzigAs6_0(.din(w_dff_B_hMZc7jZp0_0),.dout(w_dff_B_uVxzigAs6_0),.clk(gclk));
	jdff dff_B_QR9s0JAM1_0(.din(w_dff_B_uVxzigAs6_0),.dout(w_dff_B_QR9s0JAM1_0),.clk(gclk));
	jdff dff_B_0PBDAjt86_0(.din(w_dff_B_QR9s0JAM1_0),.dout(w_dff_B_0PBDAjt86_0),.clk(gclk));
	jdff dff_B_59nsSvop7_0(.din(w_dff_B_0PBDAjt86_0),.dout(w_dff_B_59nsSvop7_0),.clk(gclk));
	jdff dff_B_j2lnXHmC3_0(.din(w_dff_B_59nsSvop7_0),.dout(w_dff_B_j2lnXHmC3_0),.clk(gclk));
	jdff dff_B_JL4tlOpu9_0(.din(n1095),.dout(w_dff_B_JL4tlOpu9_0),.clk(gclk));
	jdff dff_A_tpjrM7qL1_0(.dout(w_G137_8[0]),.din(w_dff_A_tpjrM7qL1_0),.clk(gclk));
	jdff dff_A_AOW9vASK1_2(.dout(w_G137_8[2]),.din(w_dff_A_AOW9vASK1_2),.clk(gclk));
	jdff dff_A_7nfAVQrl2_2(.dout(w_dff_A_AOW9vASK1_2),.din(w_dff_A_7nfAVQrl2_2),.clk(gclk));
	jdff dff_A_y0Z6Nrwr3_2(.dout(w_dff_A_7nfAVQrl2_2),.din(w_dff_A_y0Z6Nrwr3_2),.clk(gclk));
	jdff dff_A_73R8StKX9_2(.dout(w_dff_A_y0Z6Nrwr3_2),.din(w_dff_A_73R8StKX9_2),.clk(gclk));
	jdff dff_B_9CDm9T0x5_0(.din(n1105),.dout(w_dff_B_9CDm9T0x5_0),.clk(gclk));
	jdff dff_B_vlVnsMvO5_0(.din(n1104),.dout(w_dff_B_vlVnsMvO5_0),.clk(gclk));
	jdff dff_B_BLw0u94p0_0(.din(w_dff_B_vlVnsMvO5_0),.dout(w_dff_B_BLw0u94p0_0),.clk(gclk));
	jdff dff_B_1FajR0dB6_0(.din(w_dff_B_BLw0u94p0_0),.dout(w_dff_B_1FajR0dB6_0),.clk(gclk));
	jdff dff_B_YSqoDrPk3_0(.din(w_dff_B_1FajR0dB6_0),.dout(w_dff_B_YSqoDrPk3_0),.clk(gclk));
	jdff dff_B_tVkZpNZL2_0(.din(w_dff_B_YSqoDrPk3_0),.dout(w_dff_B_tVkZpNZL2_0),.clk(gclk));
	jdff dff_B_m89Tvkcf8_0(.din(w_dff_B_tVkZpNZL2_0),.dout(w_dff_B_m89Tvkcf8_0),.clk(gclk));
	jdff dff_B_7ydwjWxg0_0(.din(w_dff_B_m89Tvkcf8_0),.dout(w_dff_B_7ydwjWxg0_0),.clk(gclk));
	jdff dff_B_lg9jCVoM4_0(.din(w_dff_B_7ydwjWxg0_0),.dout(w_dff_B_lg9jCVoM4_0),.clk(gclk));
	jdff dff_B_t7Nkqp0I4_0(.din(w_dff_B_lg9jCVoM4_0),.dout(w_dff_B_t7Nkqp0I4_0),.clk(gclk));
	jdff dff_B_6HOKj66b5_0(.din(w_dff_B_t7Nkqp0I4_0),.dout(w_dff_B_6HOKj66b5_0),.clk(gclk));
	jdff dff_B_ZRYI2TIt9_0(.din(n1103),.dout(w_dff_B_ZRYI2TIt9_0),.clk(gclk));
	jdff dff_A_DHoUckhx8_0(.dout(w_n988_3[0]),.din(w_dff_A_DHoUckhx8_0),.clk(gclk));
	jdff dff_A_TqZ9U7wu1_0(.dout(w_dff_A_DHoUckhx8_0),.din(w_dff_A_TqZ9U7wu1_0),.clk(gclk));
	jdff dff_A_sO5VoXT98_0(.dout(w_dff_A_TqZ9U7wu1_0),.din(w_dff_A_sO5VoXT98_0),.clk(gclk));
	jdff dff_A_xOGvZE8S0_0(.dout(w_dff_A_sO5VoXT98_0),.din(w_dff_A_xOGvZE8S0_0),.clk(gclk));
	jdff dff_A_Ufuh4jZt8_1(.dout(w_n988_3[1]),.din(w_dff_A_Ufuh4jZt8_1),.clk(gclk));
	jdff dff_A_60Bj9an54_1(.dout(w_dff_A_Ufuh4jZt8_1),.din(w_dff_A_60Bj9an54_1),.clk(gclk));
	jdff dff_A_uWTwpn385_0(.dout(w_n985_3[0]),.din(w_dff_A_uWTwpn385_0),.clk(gclk));
	jdff dff_A_9ez9Zel48_0(.dout(w_dff_A_uWTwpn385_0),.din(w_dff_A_9ez9Zel48_0),.clk(gclk));
	jdff dff_A_nznAk0ZQ3_1(.dout(w_n985_3[1]),.din(w_dff_A_nznAk0ZQ3_1),.clk(gclk));
	jdff dff_B_l1zv4hd97_0(.din(n1113),.dout(w_dff_B_l1zv4hd97_0),.clk(gclk));
	jdff dff_B_O7nBV4Ua1_0(.din(n1112),.dout(w_dff_B_O7nBV4Ua1_0),.clk(gclk));
	jdff dff_B_vLLMvwMo3_0(.din(w_dff_B_O7nBV4Ua1_0),.dout(w_dff_B_vLLMvwMo3_0),.clk(gclk));
	jdff dff_B_bKARqemA7_0(.din(w_dff_B_vLLMvwMo3_0),.dout(w_dff_B_bKARqemA7_0),.clk(gclk));
	jdff dff_B_Smt4RTLZ0_0(.din(w_dff_B_bKARqemA7_0),.dout(w_dff_B_Smt4RTLZ0_0),.clk(gclk));
	jdff dff_B_zXRJjpeM1_0(.din(w_dff_B_Smt4RTLZ0_0),.dout(w_dff_B_zXRJjpeM1_0),.clk(gclk));
	jdff dff_B_DtqhJbsK6_0(.din(w_dff_B_zXRJjpeM1_0),.dout(w_dff_B_DtqhJbsK6_0),.clk(gclk));
	jdff dff_B_gX4stcmz0_0(.din(w_dff_B_DtqhJbsK6_0),.dout(w_dff_B_gX4stcmz0_0),.clk(gclk));
	jdff dff_B_sbCtviuo5_0(.din(w_dff_B_gX4stcmz0_0),.dout(w_dff_B_sbCtviuo5_0),.clk(gclk));
	jdff dff_B_gnfciyQk9_0(.din(w_dff_B_sbCtviuo5_0),.dout(w_dff_B_gnfciyQk9_0),.clk(gclk));
	jdff dff_B_eCOwXywu2_0(.din(w_dff_B_gnfciyQk9_0),.dout(w_dff_B_eCOwXywu2_0),.clk(gclk));
	jdff dff_B_taxkirQY8_0(.din(w_dff_B_eCOwXywu2_0),.dout(w_dff_B_taxkirQY8_0),.clk(gclk));
	jdff dff_B_SbyRTDjy5_0(.din(w_dff_B_taxkirQY8_0),.dout(w_dff_B_SbyRTDjy5_0),.clk(gclk));
	jdff dff_B_Gg9m0Kkv7_0(.din(n1111),.dout(w_dff_B_Gg9m0Kkv7_0),.clk(gclk));
	jdff dff_B_K0FZ46m73_2(.din(G170),.dout(w_dff_B_K0FZ46m73_2),.clk(gclk));
	jdff dff_B_nGol4eN09_2(.din(G200),.dout(w_dff_B_nGol4eN09_2),.clk(gclk));
	jdff dff_B_twHeLHGu2_2(.din(w_dff_B_nGol4eN09_2),.dout(w_dff_B_twHeLHGu2_2),.clk(gclk));
	jdff dff_A_pP48pqUT3_0(.dout(w_n1002_4[0]),.din(w_dff_A_pP48pqUT3_0),.clk(gclk));
	jdff dff_A_iWfVGpi39_0(.dout(w_dff_A_pP48pqUT3_0),.din(w_dff_A_iWfVGpi39_0),.clk(gclk));
	jdff dff_A_SqWgLEWl4_0(.dout(w_dff_A_iWfVGpi39_0),.din(w_dff_A_SqWgLEWl4_0),.clk(gclk));
	jdff dff_A_uQP2s3dW3_0(.dout(w_dff_A_SqWgLEWl4_0),.din(w_dff_A_uQP2s3dW3_0),.clk(gclk));
	jdff dff_A_3rDjW8yQ0_0(.dout(w_dff_A_uQP2s3dW3_0),.din(w_dff_A_3rDjW8yQ0_0),.clk(gclk));
	jdff dff_A_vjN9xg9H3_0(.dout(w_dff_A_3rDjW8yQ0_0),.din(w_dff_A_vjN9xg9H3_0),.clk(gclk));
	jdff dff_A_JvDkBFwb9_0(.dout(w_dff_A_vjN9xg9H3_0),.din(w_dff_A_JvDkBFwb9_0),.clk(gclk));
	jdff dff_B_TmoIExVY3_0(.din(n814),.dout(w_dff_B_TmoIExVY3_0),.clk(gclk));
	jdff dff_B_E9SCZhH61_0(.din(w_dff_B_TmoIExVY3_0),.dout(w_dff_B_E9SCZhH61_0),.clk(gclk));
	jdff dff_B_5QvAAI5y1_0(.din(w_dff_B_E9SCZhH61_0),.dout(w_dff_B_5QvAAI5y1_0),.clk(gclk));
	jdff dff_B_F3FTmgG70_0(.din(w_dff_B_5QvAAI5y1_0),.dout(w_dff_B_F3FTmgG70_0),.clk(gclk));
	jdff dff_B_bZPZhxkA1_0(.din(w_dff_B_F3FTmgG70_0),.dout(w_dff_B_bZPZhxkA1_0),.clk(gclk));
	jdff dff_B_XsD4gAUV9_0(.din(w_dff_B_bZPZhxkA1_0),.dout(w_dff_B_XsD4gAUV9_0),.clk(gclk));
	jdff dff_B_rOEIVskU0_0(.din(n813),.dout(w_dff_B_rOEIVskU0_0),.clk(gclk));
	jdff dff_B_IgbdpG980_0(.din(w_dff_B_rOEIVskU0_0),.dout(w_dff_B_IgbdpG980_0),.clk(gclk));
	jdff dff_B_gbIj66MZ7_1(.din(G52),.dout(w_dff_B_gbIj66MZ7_1),.clk(gclk));
	jdff dff_B_SuVya2Y11_1(.din(w_dff_B_gbIj66MZ7_1),.dout(w_dff_B_SuVya2Y11_1),.clk(gclk));
	jdff dff_B_9zStGqWt6_0(.din(n433),.dout(w_dff_B_9zStGqWt6_0),.clk(gclk));
	jdff dff_B_axKllIrL3_1(.din(n425),.dout(w_dff_B_axKllIrL3_1),.clk(gclk));
	jdff dff_A_xlue22Q54_0(.dout(w_n999_4[0]),.din(w_dff_A_xlue22Q54_0),.clk(gclk));
	jdff dff_A_KdOGbMLL6_0(.dout(w_dff_A_xlue22Q54_0),.din(w_dff_A_KdOGbMLL6_0),.clk(gclk));
	jdff dff_A_80YT3jAo2_0(.dout(w_dff_A_KdOGbMLL6_0),.din(w_dff_A_80YT3jAo2_0),.clk(gclk));
	jdff dff_A_zU6SIoox2_0(.dout(w_dff_A_80YT3jAo2_0),.din(w_dff_A_zU6SIoox2_0),.clk(gclk));
	jdff dff_A_M8aBhL1B2_0(.dout(w_dff_A_zU6SIoox2_0),.din(w_dff_A_M8aBhL1B2_0),.clk(gclk));
	jdff dff_A_1pmCv7j60_0(.dout(w_dff_A_M8aBhL1B2_0),.din(w_dff_A_1pmCv7j60_0),.clk(gclk));
	jdff dff_A_6GGIEMOB6_0(.dout(w_dff_A_1pmCv7j60_0),.din(w_dff_A_6GGIEMOB6_0),.clk(gclk));
	jdff dff_A_HWZNkgDO3_0(.dout(w_dff_A_6GGIEMOB6_0),.din(w_dff_A_HWZNkgDO3_0),.clk(gclk));
	jdff dff_B_DZkZdZUp1_0(.din(n867),.dout(w_dff_B_DZkZdZUp1_0),.clk(gclk));
	jdff dff_B_mhqjkvYJ0_0(.din(w_dff_B_DZkZdZUp1_0),.dout(w_dff_B_mhqjkvYJ0_0),.clk(gclk));
	jdff dff_B_UtB3UMPE8_0(.din(w_dff_B_mhqjkvYJ0_0),.dout(w_dff_B_UtB3UMPE8_0),.clk(gclk));
	jdff dff_B_EEa1HfNm6_0(.din(w_dff_B_UtB3UMPE8_0),.dout(w_dff_B_EEa1HfNm6_0),.clk(gclk));
	jdff dff_B_iUyJeIbm4_0(.din(w_dff_B_EEa1HfNm6_0),.dout(w_dff_B_iUyJeIbm4_0),.clk(gclk));
	jdff dff_B_kSsGghPM6_0(.din(w_dff_B_iUyJeIbm4_0),.dout(w_dff_B_kSsGghPM6_0),.clk(gclk));
	jdff dff_B_uvfMouT79_0(.din(w_dff_B_kSsGghPM6_0),.dout(w_dff_B_uvfMouT79_0),.clk(gclk));
	jdff dff_B_tCVmtduJ1_0(.din(w_dff_B_uvfMouT79_0),.dout(w_dff_B_tCVmtduJ1_0),.clk(gclk));
	jdff dff_B_7CGqfLAq3_0(.din(n866),.dout(w_dff_B_7CGqfLAq3_0),.clk(gclk));
	jdff dff_B_fidH2dRX4_0(.din(w_dff_B_7CGqfLAq3_0),.dout(w_dff_B_fidH2dRX4_0),.clk(gclk));
	jdff dff_B_ZC1X76HY8_1(.din(G122),.dout(w_dff_B_ZC1X76HY8_1),.clk(gclk));
	jdff dff_B_5w8VRhtv0_1(.din(w_dff_B_ZC1X76HY8_1),.dout(w_dff_B_5w8VRhtv0_1),.clk(gclk));
	jdff dff_B_0p97Hk5s7_0(.din(n469),.dout(w_dff_B_0p97Hk5s7_0),.clk(gclk));
	jdff dff_B_xgN6JT9C7_1(.din(n461),.dout(w_dff_B_xgN6JT9C7_1),.clk(gclk));
	jdff dff_B_attAywGa0_1(.din(n852),.dout(w_dff_B_attAywGa0_1),.clk(gclk));
	jdff dff_B_uJk4IlmZ2_1(.din(w_dff_B_attAywGa0_1),.dout(w_dff_B_uJk4IlmZ2_1),.clk(gclk));
	jdff dff_B_jX659Nua3_1(.din(w_dff_B_uJk4IlmZ2_1),.dout(w_dff_B_jX659Nua3_1),.clk(gclk));
	jdff dff_B_zOSiBFZS0_1(.din(w_dff_B_jX659Nua3_1),.dout(w_dff_B_zOSiBFZS0_1),.clk(gclk));
	jdff dff_B_YmxJ9Gyc1_1(.din(w_dff_B_zOSiBFZS0_1),.dout(w_dff_B_YmxJ9Gyc1_1),.clk(gclk));
	jdff dff_B_6IfT1C051_1(.din(w_dff_B_YmxJ9Gyc1_1),.dout(w_dff_B_6IfT1C051_1),.clk(gclk));
	jdff dff_B_pzdm031y7_0(.din(n1121),.dout(w_dff_B_pzdm031y7_0),.clk(gclk));
	jdff dff_B_VmOlFNzb2_0(.din(w_dff_B_pzdm031y7_0),.dout(w_dff_B_VmOlFNzb2_0),.clk(gclk));
	jdff dff_B_i29EUwTc3_0(.din(w_dff_B_VmOlFNzb2_0),.dout(w_dff_B_i29EUwTc3_0),.clk(gclk));
	jdff dff_B_nOiZL7CW0_0(.din(n1120),.dout(w_dff_B_nOiZL7CW0_0),.clk(gclk));
	jdff dff_B_4T0K47LW5_0(.din(w_dff_B_nOiZL7CW0_0),.dout(w_dff_B_4T0K47LW5_0),.clk(gclk));
	jdff dff_B_znoCPcj97_0(.din(w_dff_B_4T0K47LW5_0),.dout(w_dff_B_znoCPcj97_0),.clk(gclk));
	jdff dff_B_CgxpWkET1_0(.din(w_dff_B_znoCPcj97_0),.dout(w_dff_B_CgxpWkET1_0),.clk(gclk));
	jdff dff_B_GosTMdDX1_0(.din(w_dff_B_CgxpWkET1_0),.dout(w_dff_B_GosTMdDX1_0),.clk(gclk));
	jdff dff_B_FCy4cNJc8_0(.din(w_dff_B_GosTMdDX1_0),.dout(w_dff_B_FCy4cNJc8_0),.clk(gclk));
	jdff dff_B_dLAyJeXu7_0(.din(n1119),.dout(w_dff_B_dLAyJeXu7_0),.clk(gclk));
	jdff dff_B_Xx8Rvxsi8_2(.din(G158),.dout(w_dff_B_Xx8Rvxsi8_2),.clk(gclk));
	jdff dff_B_OpNkcJd51_2(.din(G188),.dout(w_dff_B_OpNkcJd51_2),.clk(gclk));
	jdff dff_B_AmPL2t1L6_2(.din(w_dff_B_OpNkcJd51_2),.dout(w_dff_B_AmPL2t1L6_2),.clk(gclk));
	jdff dff_B_p2GlV8Jy7_0(.din(n768),.dout(w_dff_B_p2GlV8Jy7_0),.clk(gclk));
	jdff dff_B_I3ZfaRf29_0(.din(w_dff_B_p2GlV8Jy7_0),.dout(w_dff_B_I3ZfaRf29_0),.clk(gclk));
	jdff dff_B_XtwerSJ70_1(.din(G129),.dout(w_dff_B_XtwerSJ70_1),.clk(gclk));
	jdff dff_B_4HXG8lg23_1(.din(w_dff_B_XtwerSJ70_1),.dout(w_dff_B_4HXG8lg23_1),.clk(gclk));
	jdff dff_A_63OKJmVU5_1(.dout(w_n397_0[1]),.din(w_dff_A_63OKJmVU5_1),.clk(gclk));
	jdff dff_B_xSRV8uDk0_0(.din(n396),.dout(w_dff_B_xSRV8uDk0_0),.clk(gclk));
	jdff dff_B_VYhf0rRg0_1(.din(n387),.dout(w_dff_B_VYhf0rRg0_1),.clk(gclk));
	jdff dff_A_iUVppLLC3_0(.dout(w_n748_4[0]),.din(w_dff_A_iUVppLLC3_0),.clk(gclk));
	jdff dff_B_Kyt5Sm5b4_0(.din(n898),.dout(w_dff_B_Kyt5Sm5b4_0),.clk(gclk));
	jdff dff_B_mk7f2KNx4_0(.din(w_dff_B_Kyt5Sm5b4_0),.dout(w_dff_B_mk7f2KNx4_0),.clk(gclk));
	jdff dff_B_4ecwqkZP1_0(.din(w_dff_B_mk7f2KNx4_0),.dout(w_dff_B_4ecwqkZP1_0),.clk(gclk));
	jdff dff_B_vNdBs2kk8_0(.din(w_dff_B_4ecwqkZP1_0),.dout(w_dff_B_vNdBs2kk8_0),.clk(gclk));
	jdff dff_B_Tk4bzhyF1_0(.din(n897),.dout(w_dff_B_Tk4bzhyF1_0),.clk(gclk));
	jdff dff_B_RCstnGuM4_0(.din(w_dff_B_Tk4bzhyF1_0),.dout(w_dff_B_RCstnGuM4_0),.clk(gclk));
	jdff dff_B_StH4f6bM9_1(.din(G126),.dout(w_dff_B_StH4f6bM9_1),.clk(gclk));
	jdff dff_B_HudtHNcR4_1(.din(w_dff_B_StH4f6bM9_1),.dout(w_dff_B_HudtHNcR4_1),.clk(gclk));
	jdff dff_B_jgVxFdhx8_0(.din(n493),.dout(w_dff_B_jgVxFdhx8_0),.clk(gclk));
	jdff dff_B_aqDUyMwi0_1(.din(n485),.dout(w_dff_B_aqDUyMwi0_1),.clk(gclk));
	jdff dff_B_L93O4wiF6_0(.din(n889),.dout(w_dff_B_L93O4wiF6_0),.clk(gclk));
	jdff dff_A_mnovzVWq8_1(.dout(w_G137_7[1]),.din(w_dff_A_mnovzVWq8_1),.clk(gclk));
	jdff dff_A_TgrU2gMY9_1(.dout(w_dff_A_mnovzVWq8_1),.din(w_dff_A_TgrU2gMY9_1),.clk(gclk));
	jdff dff_A_83YjOvyh2_1(.dout(w_dff_A_TgrU2gMY9_1),.din(w_dff_A_83YjOvyh2_1),.clk(gclk));
	jdff dff_A_JJMcdgTq7_1(.dout(w_dff_A_83YjOvyh2_1),.din(w_dff_A_JJMcdgTq7_1),.clk(gclk));
	jdff dff_A_Bo1joco45_2(.dout(w_G137_7[2]),.din(w_dff_A_Bo1joco45_2),.clk(gclk));
	jdff dff_A_3Z2ePtAG1_2(.dout(w_dff_A_Bo1joco45_2),.din(w_dff_A_3Z2ePtAG1_2),.clk(gclk));
	jdff dff_A_JQQuOTlV8_0(.dout(w_G137_2[0]),.din(w_dff_A_JQQuOTlV8_0),.clk(gclk));
	jdff dff_A_dE52QEdm5_0(.dout(w_dff_A_JQQuOTlV8_0),.din(w_dff_A_dE52QEdm5_0),.clk(gclk));
	jdff dff_A_dgFbPYSa1_0(.dout(w_dff_A_dE52QEdm5_0),.din(w_dff_A_dgFbPYSa1_0),.clk(gclk));
	jdff dff_A_lp1paIgS1_0(.dout(w_dff_A_dgFbPYSa1_0),.din(w_dff_A_lp1paIgS1_0),.clk(gclk));
	jdff dff_A_gbgVv3vG8_1(.dout(w_G137_2[1]),.din(w_dff_A_gbgVv3vG8_1),.clk(gclk));
	jdff dff_A_M96opvhU6_1(.dout(w_dff_A_gbgVv3vG8_1),.din(w_dff_A_M96opvhU6_1),.clk(gclk));
	jdff dff_A_y4CvdwjM4_1(.dout(w_dff_A_M96opvhU6_1),.din(w_dff_A_y4CvdwjM4_1),.clk(gclk));
	jdff dff_A_HWQavakt8_1(.dout(w_dff_A_y4CvdwjM4_1),.din(w_dff_A_HWQavakt8_1),.clk(gclk));
	jdff dff_B_8NqKbRgT0_0(.din(n1129),.dout(w_dff_B_8NqKbRgT0_0),.clk(gclk));
	jdff dff_B_db45aS7f7_0(.din(w_dff_B_8NqKbRgT0_0),.dout(w_dff_B_db45aS7f7_0),.clk(gclk));
	jdff dff_B_b2Kv6wiO3_0(.din(n1128),.dout(w_dff_B_b2Kv6wiO3_0),.clk(gclk));
	jdff dff_B_4K5w1RAJ4_0(.din(w_dff_B_b2Kv6wiO3_0),.dout(w_dff_B_4K5w1RAJ4_0),.clk(gclk));
	jdff dff_B_8WeFoxZH2_0(.din(w_dff_B_4K5w1RAJ4_0),.dout(w_dff_B_8WeFoxZH2_0),.clk(gclk));
	jdff dff_B_IZ8sqVnY6_0(.din(w_dff_B_8WeFoxZH2_0),.dout(w_dff_B_IZ8sqVnY6_0),.clk(gclk));
	jdff dff_B_1lDDg48k9_0(.din(w_dff_B_IZ8sqVnY6_0),.dout(w_dff_B_1lDDg48k9_0),.clk(gclk));
	jdff dff_B_kQPD1IDn1_0(.din(w_dff_B_1lDDg48k9_0),.dout(w_dff_B_kQPD1IDn1_0),.clk(gclk));
	jdff dff_B_KRHTHDfL9_0(.din(w_dff_B_kQPD1IDn1_0),.dout(w_dff_B_KRHTHDfL9_0),.clk(gclk));
	jdff dff_B_DgGrCXuz6_0(.din(w_dff_B_KRHTHDfL9_0),.dout(w_dff_B_DgGrCXuz6_0),.clk(gclk));
	jdff dff_B_iywwfrfp0_0(.din(n1127),.dout(w_dff_B_iywwfrfp0_0),.clk(gclk));
	jdff dff_B_nJEeufId6_2(.din(G152),.dout(w_dff_B_nJEeufId6_2),.clk(gclk));
	jdff dff_B_cPKK66sL5_2(.din(G155),.dout(w_dff_B_cPKK66sL5_2),.clk(gclk));
	jdff dff_B_Hr5Ef1GE8_2(.din(w_dff_B_cPKK66sL5_2),.dout(w_dff_B_Hr5Ef1GE8_2),.clk(gclk));
	jdff dff_B_eTOjnUJH1_0(.din(n837),.dout(w_dff_B_eTOjnUJH1_0),.clk(gclk));
	jdff dff_B_Y9Tox2yI6_0(.din(w_dff_B_eTOjnUJH1_0),.dout(w_dff_B_Y9Tox2yI6_0),.clk(gclk));
	jdff dff_B_d2tuIZ0h6_0(.din(n836),.dout(w_dff_B_d2tuIZ0h6_0),.clk(gclk));
	jdff dff_B_0cnio3gY3_0(.din(w_dff_B_d2tuIZ0h6_0),.dout(w_dff_B_0cnio3gY3_0),.clk(gclk));
	jdff dff_B_soVvpI2f9_1(.din(G119),.dout(w_dff_B_soVvpI2f9_1),.clk(gclk));
	jdff dff_B_6P5kMzZz0_1(.din(w_dff_B_soVvpI2f9_1),.dout(w_dff_B_6P5kMzZz0_1),.clk(gclk));
	jdff dff_B_Ub8q9oaB2_0(.din(n444),.dout(w_dff_B_Ub8q9oaB2_0),.clk(gclk));
	jdff dff_B_8S4t6fQz2_1(.din(n436),.dout(w_dff_B_8S4t6fQz2_1),.clk(gclk));
	jdff dff_A_ifTUOtl82_0(.dout(w_n744_1[0]),.din(w_dff_A_ifTUOtl82_0),.clk(gclk));
	jdff dff_A_zmsw4He95_0(.dout(w_dff_A_ifTUOtl82_0),.din(w_dff_A_zmsw4He95_0),.clk(gclk));
	jdff dff_A_v2FYbrdu1_0(.dout(w_dff_A_zmsw4He95_0),.din(w_dff_A_v2FYbrdu1_0),.clk(gclk));
	jdff dff_A_uCaByIzH4_0(.dout(w_dff_A_v2FYbrdu1_0),.din(w_dff_A_uCaByIzH4_0),.clk(gclk));
	jdff dff_A_f9tb60g82_0(.dout(w_dff_A_uCaByIzH4_0),.din(w_dff_A_f9tb60g82_0),.clk(gclk));
	jdff dff_A_4v02IntC4_0(.dout(w_dff_A_f9tb60g82_0),.din(w_dff_A_4v02IntC4_0),.clk(gclk));
	jdff dff_B_zk4Cjs9z8_0(.din(n887),.dout(w_dff_B_zk4Cjs9z8_0),.clk(gclk));
	jdff dff_B_qGCxqqTx3_0(.din(w_dff_B_zk4Cjs9z8_0),.dout(w_dff_B_qGCxqqTx3_0),.clk(gclk));
	jdff dff_B_DTINZc7i8_0(.din(w_dff_B_qGCxqqTx3_0),.dout(w_dff_B_DTINZc7i8_0),.clk(gclk));
	jdff dff_B_A4XoTYjY2_0(.din(w_dff_B_DTINZc7i8_0),.dout(w_dff_B_A4XoTYjY2_0),.clk(gclk));
	jdff dff_B_fCDC6jCd4_0(.din(w_dff_B_A4XoTYjY2_0),.dout(w_dff_B_fCDC6jCd4_0),.clk(gclk));
	jdff dff_B_7f9Yqb9p3_0(.din(n886),.dout(w_dff_B_7f9Yqb9p3_0),.clk(gclk));
	jdff dff_B_SUKWI2E52_0(.din(w_dff_B_7f9Yqb9p3_0),.dout(w_dff_B_SUKWI2E52_0),.clk(gclk));
	jdff dff_B_O8ilfwh16_1(.din(G127),.dout(w_dff_B_O8ilfwh16_1),.clk(gclk));
	jdff dff_B_JkvKrsif8_1(.din(w_dff_B_O8ilfwh16_1),.dout(w_dff_B_JkvKrsif8_1),.clk(gclk));
	jdff dff_A_9vwwXxKD4_1(.dout(w_n459_0[1]),.din(w_dff_A_9vwwXxKD4_1),.clk(gclk));
	jdff dff_B_aqqTLBTb6_0(.din(n458),.dout(w_dff_B_aqqTLBTb6_0),.clk(gclk));
	jdff dff_B_YQcTVDeX3_1(.din(n450),.dout(w_dff_B_YQcTVDeX3_1),.clk(gclk));
	jdff dff_B_wvmvDo3N4_0(.din(n1137),.dout(w_dff_B_wvmvDo3N4_0),.clk(gclk));
	jdff dff_B_fIZA17lP3_0(.din(n1136),.dout(w_dff_B_fIZA17lP3_0),.clk(gclk));
	jdff dff_B_DvjY02gE6_0(.din(w_dff_B_fIZA17lP3_0),.dout(w_dff_B_DvjY02gE6_0),.clk(gclk));
	jdff dff_B_XYgIO2Lu7_0(.din(w_dff_B_DvjY02gE6_0),.dout(w_dff_B_XYgIO2Lu7_0),.clk(gclk));
	jdff dff_B_679AlWQc6_0(.din(w_dff_B_XYgIO2Lu7_0),.dout(w_dff_B_679AlWQc6_0),.clk(gclk));
	jdff dff_B_V8jDugkm8_0(.din(w_dff_B_679AlWQc6_0),.dout(w_dff_B_V8jDugkm8_0),.clk(gclk));
	jdff dff_B_Y3TkIGnK5_0(.din(w_dff_B_V8jDugkm8_0),.dout(w_dff_B_Y3TkIGnK5_0),.clk(gclk));
	jdff dff_B_onUrTJDO2_0(.din(w_dff_B_Y3TkIGnK5_0),.dout(w_dff_B_onUrTJDO2_0),.clk(gclk));
	jdff dff_B_2iN4p2J15_0(.din(w_dff_B_onUrTJDO2_0),.dout(w_dff_B_2iN4p2J15_0),.clk(gclk));
	jdff dff_B_rERWmI323_0(.din(w_dff_B_2iN4p2J15_0),.dout(w_dff_B_rERWmI323_0),.clk(gclk));
	jdff dff_B_WWmRkjpa6_0(.din(w_dff_B_rERWmI323_0),.dout(w_dff_B_WWmRkjpa6_0),.clk(gclk));
	jdff dff_B_V1GNE4et7_0(.din(n1135),.dout(w_dff_B_V1GNE4et7_0),.clk(gclk));
	jdff dff_B_p5VKIVOZ9_2(.din(G146),.dout(w_dff_B_p5VKIVOZ9_2),.clk(gclk));
	jdff dff_B_ykPNCXRN2_2(.din(G149),.dout(w_dff_B_ykPNCXRN2_2),.clk(gclk));
	jdff dff_B_VdpNh2Zg3_2(.din(w_dff_B_ykPNCXRN2_2),.dout(w_dff_B_VdpNh2Zg3_2),.clk(gclk));
	jdff dff_A_zULHyfoe2_0(.dout(w_n1002_3[0]),.din(w_dff_A_zULHyfoe2_0),.clk(gclk));
	jdff dff_A_XenlyZdW2_0(.dout(w_dff_A_zULHyfoe2_0),.din(w_dff_A_XenlyZdW2_0),.clk(gclk));
	jdff dff_A_bwyYPt6z6_0(.dout(w_dff_A_XenlyZdW2_0),.din(w_dff_A_bwyYPt6z6_0),.clk(gclk));
	jdff dff_A_kfhIpUYa8_0(.dout(w_dff_A_bwyYPt6z6_0),.din(w_dff_A_kfhIpUYa8_0),.clk(gclk));
	jdff dff_A_GiaJWmrs0_1(.dout(w_n1002_3[1]),.din(w_dff_A_GiaJWmrs0_1),.clk(gclk));
	jdff dff_A_lDdfJqoX7_1(.dout(w_dff_A_GiaJWmrs0_1),.din(w_dff_A_lDdfJqoX7_1),.clk(gclk));
	jdff dff_B_9TjBKOBe6_0(.din(n826),.dout(w_dff_B_9TjBKOBe6_0),.clk(gclk));
	jdff dff_B_YpB0HddL0_0(.din(w_dff_B_9TjBKOBe6_0),.dout(w_dff_B_YpB0HddL0_0),.clk(gclk));
	jdff dff_B_lorW02c28_0(.din(w_dff_B_YpB0HddL0_0),.dout(w_dff_B_lorW02c28_0),.clk(gclk));
	jdff dff_B_8lKEEDpE1_0(.din(w_dff_B_lorW02c28_0),.dout(w_dff_B_8lKEEDpE1_0),.clk(gclk));
	jdff dff_B_Ny5gWR5V1_0(.din(w_dff_B_8lKEEDpE1_0),.dout(w_dff_B_Ny5gWR5V1_0),.clk(gclk));
	jdff dff_B_SfDirKpW0_0(.din(n824),.dout(w_dff_B_SfDirKpW0_0),.clk(gclk));
	jdff dff_B_QzOQW9zY4_1(.din(G130),.dout(w_dff_B_QzOQW9zY4_1),.clk(gclk));
	jdff dff_B_MZ5fi9cp2_1(.din(w_dff_B_QzOQW9zY4_1),.dout(w_dff_B_MZ5fi9cp2_1),.clk(gclk));
	jdff dff_B_lTcAT0Ce7_0(.din(n413),.dout(w_dff_B_lTcAT0Ce7_0),.clk(gclk));
	jdff dff_B_VORGvKop1_1(.din(n816),.dout(w_dff_B_VORGvKop1_1),.clk(gclk));
	jdff dff_B_Sk8udyQC8_1(.din(w_dff_B_VORGvKop1_1),.dout(w_dff_B_Sk8udyQC8_1),.clk(gclk));
	jdff dff_B_h6bF9BiN0_1(.din(w_dff_B_Sk8udyQC8_1),.dout(w_dff_B_h6bF9BiN0_1),.clk(gclk));
	jdff dff_B_SbwYihbX8_1(.din(w_dff_B_h6bF9BiN0_1),.dout(w_dff_B_SbwYihbX8_1),.clk(gclk));
	jdff dff_B_exRqFS4L6_1(.din(w_dff_B_SbwYihbX8_1),.dout(w_dff_B_exRqFS4L6_1),.clk(gclk));
	jdff dff_A_PPOdDa8V8_2(.dout(w_n744_0[2]),.din(w_dff_A_PPOdDa8V8_2),.clk(gclk));
	jdff dff_A_ICgvkPBk2_2(.dout(w_dff_A_PPOdDa8V8_2),.din(w_dff_A_ICgvkPBk2_2),.clk(gclk));
	jdff dff_A_eYXBz0vJ8_2(.dout(w_dff_A_ICgvkPBk2_2),.din(w_dff_A_eYXBz0vJ8_2),.clk(gclk));
	jdff dff_A_AhU7oceG6_2(.dout(w_dff_A_eYXBz0vJ8_2),.din(w_dff_A_AhU7oceG6_2),.clk(gclk));
	jdff dff_B_n7jQxknP7_3(.din(n744),.dout(w_dff_B_n7jQxknP7_3),.clk(gclk));
	jdff dff_B_IRVa1Pmb5_3(.din(w_dff_B_n7jQxknP7_3),.dout(w_dff_B_IRVa1Pmb5_3),.clk(gclk));
	jdff dff_A_2uWg91iH6_1(.dout(w_n748_3[1]),.din(w_dff_A_2uWg91iH6_1),.clk(gclk));
	jdff dff_A_8g0vU4iT8_1(.dout(w_dff_A_2uWg91iH6_1),.din(w_dff_A_8g0vU4iT8_1),.clk(gclk));
	jdff dff_A_zbzUghjV0_2(.dout(w_n748_3[2]),.din(w_dff_A_zbzUghjV0_2),.clk(gclk));
	jdff dff_A_EJ0STCnJ7_2(.dout(w_dff_A_zbzUghjV0_2),.din(w_dff_A_EJ0STCnJ7_2),.clk(gclk));
	jdff dff_A_lzzscTAx1_2(.dout(w_dff_A_EJ0STCnJ7_2),.din(w_dff_A_lzzscTAx1_2),.clk(gclk));
	jdff dff_A_4NeCTvRO6_2(.dout(w_dff_A_lzzscTAx1_2),.din(w_dff_A_4NeCTvRO6_2),.clk(gclk));
	jdff dff_A_lRHEjDTu5_0(.dout(w_n999_3[0]),.din(w_dff_A_lRHEjDTu5_0),.clk(gclk));
	jdff dff_A_33UYVb7Q4_0(.dout(w_dff_A_lRHEjDTu5_0),.din(w_dff_A_33UYVb7Q4_0),.clk(gclk));
	jdff dff_A_1nYUCOUx3_1(.dout(w_n999_3[1]),.din(w_dff_A_1nYUCOUx3_1),.clk(gclk));
	jdff dff_B_HxKjyXgw0_0(.din(n874),.dout(w_dff_B_HxKjyXgw0_0),.clk(gclk));
	jdff dff_B_xC1SjRwX8_0(.din(w_dff_B_HxKjyXgw0_0),.dout(w_dff_B_xC1SjRwX8_0),.clk(gclk));
	jdff dff_B_OyxPJ0tF4_0(.din(w_dff_B_xC1SjRwX8_0),.dout(w_dff_B_OyxPJ0tF4_0),.clk(gclk));
	jdff dff_B_mIpnp5UF0_0(.din(w_dff_B_OyxPJ0tF4_0),.dout(w_dff_B_mIpnp5UF0_0),.clk(gclk));
	jdff dff_B_HQ3sJb4f2_0(.din(w_dff_B_mIpnp5UF0_0),.dout(w_dff_B_HQ3sJb4f2_0),.clk(gclk));
	jdff dff_B_DggdxiwR2_0(.din(w_dff_B_HQ3sJb4f2_0),.dout(w_dff_B_DggdxiwR2_0),.clk(gclk));
	jdff dff_B_N2QLohcD1_0(.din(n873),.dout(w_dff_B_N2QLohcD1_0),.clk(gclk));
	jdff dff_B_xHXuatwA1_0(.din(w_dff_B_N2QLohcD1_0),.dout(w_dff_B_xHXuatwA1_0),.clk(gclk));
	jdff dff_B_sBsDkjNf9_1(.din(G128),.dout(w_dff_B_sBsDkjNf9_1),.clk(gclk));
	jdff dff_B_RdiaBO6R4_1(.din(w_dff_B_sBsDkjNf9_1),.dout(w_dff_B_RdiaBO6R4_1),.clk(gclk));
	jdff dff_B_SzZAg0xl2_0(.din(n480),.dout(w_dff_B_SzZAg0xl2_0),.clk(gclk));
	jdff dff_B_Owewop3E6_1(.din(n472),.dout(w_dff_B_Owewop3E6_1),.clk(gclk));
	jdff dff_B_5todjbo18_0(.din(n858),.dout(w_dff_B_5todjbo18_0),.clk(gclk));
	jdff dff_A_hmZACMxk8_0(.dout(w_G4_1[0]),.din(w_dff_A_hmZACMxk8_0),.clk(gclk));
	jdff dff_A_R9unRN3k7_0(.dout(w_dff_A_hmZACMxk8_0),.din(w_dff_A_R9unRN3k7_0),.clk(gclk));
	jdff dff_A_YeufBsyB9_0(.dout(w_dff_A_R9unRN3k7_0),.din(w_dff_A_YeufBsyB9_0),.clk(gclk));
	jdff dff_A_Xsi80K702_0(.dout(w_dff_A_YeufBsyB9_0),.din(w_dff_A_Xsi80K702_0),.clk(gclk));
	jdff dff_B_OQo50X6U1_0(.din(n1155),.dout(w_dff_B_OQo50X6U1_0),.clk(gclk));
	jdff dff_B_Ilzeax6d3_0(.din(w_dff_B_OQo50X6U1_0),.dout(w_dff_B_Ilzeax6d3_0),.clk(gclk));
	jdff dff_B_bOa9Utrz7_0(.din(w_dff_B_Ilzeax6d3_0),.dout(w_dff_B_bOa9Utrz7_0),.clk(gclk));
	jdff dff_B_uHTSgQkm2_0(.din(w_dff_B_bOa9Utrz7_0),.dout(w_dff_B_uHTSgQkm2_0),.clk(gclk));
	jdff dff_B_MsNhVbX91_0(.din(w_dff_B_uHTSgQkm2_0),.dout(w_dff_B_MsNhVbX91_0),.clk(gclk));
	jdff dff_B_AHIgh2vR2_0(.din(w_dff_B_MsNhVbX91_0),.dout(w_dff_B_AHIgh2vR2_0),.clk(gclk));
	jdff dff_B_iziWwFyk4_0(.din(w_dff_B_AHIgh2vR2_0),.dout(w_dff_B_iziWwFyk4_0),.clk(gclk));
	jdff dff_B_kPhERWyU0_0(.din(w_dff_B_iziWwFyk4_0),.dout(w_dff_B_kPhERWyU0_0),.clk(gclk));
	jdff dff_B_KBIWN7di2_0(.din(w_dff_B_kPhERWyU0_0),.dout(w_dff_B_KBIWN7di2_0),.clk(gclk));
	jdff dff_B_DxHOchE57_0(.din(w_dff_B_KBIWN7di2_0),.dout(w_dff_B_DxHOchE57_0),.clk(gclk));
	jdff dff_B_adloSAdU0_0(.din(w_dff_B_DxHOchE57_0),.dout(w_dff_B_adloSAdU0_0),.clk(gclk));
	jdff dff_B_j74uReLR5_0(.din(w_dff_B_adloSAdU0_0),.dout(w_dff_B_j74uReLR5_0),.clk(gclk));
	jdff dff_B_yblj741h6_1(.din(n1148),.dout(w_dff_B_yblj741h6_1),.clk(gclk));
	jdff dff_B_9VscNHJl5_1(.din(w_dff_B_yblj741h6_1),.dout(w_dff_B_9VscNHJl5_1),.clk(gclk));
	jdff dff_B_gqoiLU3g3_1(.din(w_dff_B_9VscNHJl5_1),.dout(w_dff_B_gqoiLU3g3_1),.clk(gclk));
	jdff dff_B_gQw9j5Cc2_1(.din(w_dff_B_gqoiLU3g3_1),.dout(w_dff_B_gQw9j5Cc2_1),.clk(gclk));
	jdff dff_B_eI2359Qg3_1(.din(w_dff_B_gQw9j5Cc2_1),.dout(w_dff_B_eI2359Qg3_1),.clk(gclk));
	jdff dff_B_HixqNAtj8_1(.din(n1150),.dout(w_dff_B_HixqNAtj8_1),.clk(gclk));
	jdff dff_B_I1nJ34tq1_0(.din(n1144),.dout(w_dff_B_I1nJ34tq1_0),.clk(gclk));
	jdff dff_B_zK58RImn5_0(.din(w_dff_B_I1nJ34tq1_0),.dout(w_dff_B_zK58RImn5_0),.clk(gclk));
	jdff dff_B_ILi98yKd8_0(.din(w_dff_B_zK58RImn5_0),.dout(w_dff_B_ILi98yKd8_0),.clk(gclk));
	jdff dff_B_S2mQ5caC3_0(.din(w_dff_B_ILi98yKd8_0),.dout(w_dff_B_S2mQ5caC3_0),.clk(gclk));
	jdff dff_B_iZqf4yul8_0(.din(w_dff_B_S2mQ5caC3_0),.dout(w_dff_B_iZqf4yul8_0),.clk(gclk));
	jdff dff_B_UHrS96262_0(.din(w_dff_B_iZqf4yul8_0),.dout(w_dff_B_UHrS96262_0),.clk(gclk));
	jdff dff_B_Zuaqtahp2_0(.din(w_dff_B_UHrS96262_0),.dout(w_dff_B_Zuaqtahp2_0),.clk(gclk));
	jdff dff_B_7JSgG3i04_0(.din(w_dff_B_Zuaqtahp2_0),.dout(w_dff_B_7JSgG3i04_0),.clk(gclk));
	jdff dff_B_ebQFglhz0_0(.din(w_dff_B_7JSgG3i04_0),.dout(w_dff_B_ebQFglhz0_0),.clk(gclk));
	jdff dff_B_hHIZ0iXp5_0(.din(w_dff_B_ebQFglhz0_0),.dout(w_dff_B_hHIZ0iXp5_0),.clk(gclk));
	jdff dff_B_VDvsx6FZ6_0(.din(w_dff_B_hHIZ0iXp5_0),.dout(w_dff_B_VDvsx6FZ6_0),.clk(gclk));
	jdff dff_B_5UYAlVGf3_0(.din(w_dff_B_VDvsx6FZ6_0),.dout(w_dff_B_5UYAlVGf3_0),.clk(gclk));
	jdff dff_B_cGTaa0N48_0(.din(w_dff_B_5UYAlVGf3_0),.dout(w_dff_B_cGTaa0N48_0),.clk(gclk));
	jdff dff_B_4YmmOZDP2_0(.din(w_dff_B_cGTaa0N48_0),.dout(w_dff_B_4YmmOZDP2_0),.clk(gclk));
	jdff dff_B_JaxA3jff9_0(.din(w_dff_B_4YmmOZDP2_0),.dout(w_dff_B_JaxA3jff9_0),.clk(gclk));
	jdff dff_B_i7iBOFlZ4_0(.din(w_dff_B_JaxA3jff9_0),.dout(w_dff_B_i7iBOFlZ4_0),.clk(gclk));
	jdff dff_B_ugPAGpWl0_1(.din(n1141),.dout(w_dff_B_ugPAGpWl0_1),.clk(gclk));
	jdff dff_A_4XsvK0hY4_0(.dout(w_n1142_0[0]),.din(w_dff_A_4XsvK0hY4_0),.clk(gclk));
	jdff dff_A_VELsOET54_0(.dout(w_dff_A_4XsvK0hY4_0),.din(w_dff_A_VELsOET54_0),.clk(gclk));
	jdff dff_A_QgDlqxAf5_0(.dout(w_dff_A_VELsOET54_0),.din(w_dff_A_QgDlqxAf5_0),.clk(gclk));
	jdff dff_A_NuwZW70N1_0(.dout(w_G3717_0[0]),.din(w_dff_A_NuwZW70N1_0),.clk(gclk));
	jdff dff_A_93rcbJ8W5_0(.dout(w_dff_A_NuwZW70N1_0),.din(w_dff_A_93rcbJ8W5_0),.clk(gclk));
	jdff dff_A_LFMcXJ298_0(.dout(w_dff_A_93rcbJ8W5_0),.din(w_dff_A_LFMcXJ298_0),.clk(gclk));
	jdff dff_A_OA0AK7At2_0(.dout(w_dff_A_LFMcXJ298_0),.din(w_dff_A_OA0AK7At2_0),.clk(gclk));
	jdff dff_A_iA5EtpUZ7_0(.dout(w_dff_A_OA0AK7At2_0),.din(w_dff_A_iA5EtpUZ7_0),.clk(gclk));
	jdff dff_A_HcqOZvGd0_0(.dout(w_G3724_0[0]),.din(w_dff_A_HcqOZvGd0_0),.clk(gclk));
	jdff dff_A_IHhhvd3w7_0(.dout(w_dff_A_HcqOZvGd0_0),.din(w_dff_A_IHhhvd3w7_0),.clk(gclk));
	jdff dff_A_aZL3SwJX9_0(.dout(w_dff_A_IHhhvd3w7_0),.din(w_dff_A_aZL3SwJX9_0),.clk(gclk));
	jdff dff_A_f94wbbgQ4_0(.dout(w_dff_A_aZL3SwJX9_0),.din(w_dff_A_f94wbbgQ4_0),.clk(gclk));
	jdff dff_A_88dYPDEu9_2(.dout(w_G3724_0[2]),.din(w_dff_A_88dYPDEu9_2),.clk(gclk));
	jdff dff_A_yIsJvCgR8_2(.dout(w_dff_A_88dYPDEu9_2),.din(w_dff_A_yIsJvCgR8_2),.clk(gclk));
	jdff dff_A_i2oHWcU87_2(.dout(w_dff_A_yIsJvCgR8_2),.din(w_dff_A_i2oHWcU87_2),.clk(gclk));
	jdff dff_A_00MZFfXb4_2(.dout(w_dff_A_i2oHWcU87_2),.din(w_dff_A_00MZFfXb4_2),.clk(gclk));
	jdff dff_A_LJ05JdEi1_2(.dout(w_dff_A_00MZFfXb4_2),.din(w_dff_A_LJ05JdEi1_2),.clk(gclk));
	jdff dff_A_nEs3OTwA1_2(.dout(w_dff_A_LJ05JdEi1_2),.din(w_dff_A_nEs3OTwA1_2),.clk(gclk));
	jdff dff_A_sefpTJnz7_2(.dout(w_dff_A_nEs3OTwA1_2),.din(w_dff_A_sefpTJnz7_2),.clk(gclk));
	jdff dff_A_rSzX3Gc14_2(.dout(w_dff_A_sefpTJnz7_2),.din(w_dff_A_rSzX3Gc14_2),.clk(gclk));
	jdff dff_A_3xtNxIFQ1_2(.dout(w_dff_A_rSzX3Gc14_2),.din(w_dff_A_3xtNxIFQ1_2),.clk(gclk));
	jdff dff_A_9Nfi2wJt9_2(.dout(w_dff_A_3xtNxIFQ1_2),.din(w_dff_A_9Nfi2wJt9_2),.clk(gclk));
	jdff dff_A_fIgYN3Ul8_2(.dout(w_dff_A_9Nfi2wJt9_2),.din(w_dff_A_fIgYN3Ul8_2),.clk(gclk));
	jdff dff_A_urRTYDO26_2(.dout(w_dff_A_fIgYN3Ul8_2),.din(w_dff_A_urRTYDO26_2),.clk(gclk));
	jdff dff_A_xf66lUCa1_2(.dout(w_dff_A_urRTYDO26_2),.din(w_dff_A_xf66lUCa1_2),.clk(gclk));
	jdff dff_A_OxNUh6XI1_2(.dout(w_dff_A_xf66lUCa1_2),.din(w_dff_A_OxNUh6XI1_2),.clk(gclk));
	jdff dff_A_O0lssmRo2_2(.dout(w_dff_A_OxNUh6XI1_2),.din(w_dff_A_O0lssmRo2_2),.clk(gclk));
	jdff dff_A_Z9sIK7Ul3_2(.dout(w_dff_A_O0lssmRo2_2),.din(w_dff_A_Z9sIK7Ul3_2),.clk(gclk));
	jdff dff_A_L7UmcHcD4_2(.dout(w_dff_A_Z9sIK7Ul3_2),.din(w_dff_A_L7UmcHcD4_2),.clk(gclk));
	jdff dff_A_QtV3GtD43_2(.dout(w_dff_A_L7UmcHcD4_2),.din(w_dff_A_QtV3GtD43_2),.clk(gclk));
	jdff dff_A_MIOownFJ9_0(.dout(w_G132_0[0]),.din(w_dff_A_MIOownFJ9_0),.clk(gclk));
	jdff dff_A_1MSLH93I7_0(.dout(w_dff_A_MIOownFJ9_0),.din(w_dff_A_1MSLH93I7_0),.clk(gclk));
	jdff dff_A_CauE5RpT8_0(.dout(w_dff_A_1MSLH93I7_0),.din(w_dff_A_CauE5RpT8_0),.clk(gclk));
	jdff dff_A_yMnJDmyu7_0(.dout(w_dff_A_CauE5RpT8_0),.din(w_dff_A_yMnJDmyu7_0),.clk(gclk));
	jdff dff_A_nL85My2h9_0(.dout(w_dff_A_yMnJDmyu7_0),.din(w_dff_A_nL85My2h9_0),.clk(gclk));
	jdff dff_A_BgO5cR615_0(.dout(w_dff_A_nL85My2h9_0),.din(w_dff_A_BgO5cR615_0),.clk(gclk));
	jdff dff_A_DYNBgs530_0(.dout(w_dff_A_BgO5cR615_0),.din(w_dff_A_DYNBgs530_0),.clk(gclk));
	jdff dff_A_rLHIpSQp7_0(.dout(w_dff_A_DYNBgs530_0),.din(w_dff_A_rLHIpSQp7_0),.clk(gclk));
	jdff dff_A_rSC5yAMZ6_0(.dout(w_dff_A_rLHIpSQp7_0),.din(w_dff_A_rSC5yAMZ6_0),.clk(gclk));
	jdff dff_A_m5ONKO6z3_0(.dout(w_dff_A_rSC5yAMZ6_0),.din(w_dff_A_m5ONKO6z3_0),.clk(gclk));
	jdff dff_A_TTPrAq6q7_0(.dout(w_dff_A_m5ONKO6z3_0),.din(w_dff_A_TTPrAq6q7_0),.clk(gclk));
	jdff dff_A_nOXqYiFV2_0(.dout(w_dff_A_TTPrAq6q7_0),.din(w_dff_A_nOXqYiFV2_0),.clk(gclk));
	jdff dff_A_1gwjD4y12_0(.dout(w_dff_A_nOXqYiFV2_0),.din(w_dff_A_1gwjD4y12_0),.clk(gclk));
	jdff dff_B_Dv6mIgGh6_2(.din(G132),.dout(w_dff_B_Dv6mIgGh6_2),.clk(gclk));
	jdff dff_B_SdFwrvQ83_2(.din(w_dff_B_Dv6mIgGh6_2),.dout(w_dff_B_SdFwrvQ83_2),.clk(gclk));
	jdff dff_B_EIYVk1i47_2(.din(w_dff_B_SdFwrvQ83_2),.dout(w_dff_B_EIYVk1i47_2),.clk(gclk));
	jdff dff_B_GjqMQ1wZ2_1(.din(n1184),.dout(w_dff_B_GjqMQ1wZ2_1),.clk(gclk));
	jdff dff_B_9It1tp8z4_0(.din(n1189),.dout(w_dff_B_9It1tp8z4_0),.clk(gclk));
	jdff dff_B_6yWgKtOw7_0(.din(w_dff_B_9It1tp8z4_0),.dout(w_dff_B_6yWgKtOw7_0),.clk(gclk));
	jdff dff_B_7qWwFGV17_0(.din(n1187),.dout(w_dff_B_7qWwFGV17_0),.clk(gclk));
	jdff dff_A_24pca0HV7_0(.dout(w_G601_0),.din(w_dff_A_24pca0HV7_0),.clk(gclk));
	jdff dff_B_9v0UvJns1_1(.din(n656),.dout(w_dff_B_9v0UvJns1_1),.clk(gclk));
	jdff dff_A_tO90tMmr9_0(.dout(w_n671_0[0]),.din(w_dff_A_tO90tMmr9_0),.clk(gclk));
	jdff dff_B_zK5lCcxZ2_1(.din(n665),.dout(w_dff_B_zK5lCcxZ2_1),.clk(gclk));
	jdff dff_B_bZ2YK1Iu4_1(.din(n907),.dout(w_dff_B_bZ2YK1Iu4_1),.clk(gclk));
	jdff dff_B_IrMKE7qT9_1(.din(n909),.dout(w_dff_B_IrMKE7qT9_1),.clk(gclk));
	jdff dff_B_fsiWhS0U1_1(.din(w_dff_B_IrMKE7qT9_1),.dout(w_dff_B_fsiWhS0U1_1),.clk(gclk));
	jdff dff_B_u60iEu935_0(.din(n910),.dout(w_dff_B_u60iEu935_0),.clk(gclk));
	jdff dff_B_ZpFDWVFP4_1(.din(n908),.dout(w_dff_B_ZpFDWVFP4_1),.clk(gclk));
	jdff dff_B_XwVNHKM36_0(.din(n904),.dout(w_dff_B_XwVNHKM36_0),.clk(gclk));
	jdff dff_A_5m1sBFBP3_0(.dout(w_G369_0[0]),.din(w_dff_A_5m1sBFBP3_0),.clk(gclk));
	jdff dff_A_2gEbBQhW3_0(.dout(w_n621_1[0]),.din(w_dff_A_2gEbBQhW3_0),.clk(gclk));
	jdff dff_A_5sB5Qmdb9_0(.dout(w_dff_A_2gEbBQhW3_0),.din(w_dff_A_5sB5Qmdb9_0),.clk(gclk));
	jdff dff_A_1raUQNaH4_0(.dout(w_dff_A_5sB5Qmdb9_0),.din(w_dff_A_1raUQNaH4_0),.clk(gclk));
	jdff dff_B_WwIkTV058_0(.din(n921),.dout(w_dff_B_WwIkTV058_0),.clk(gclk));
	jdff dff_A_X2w1lQ6U1_0(.dout(w_G289_0[0]),.din(w_dff_A_X2w1lQ6U1_0),.clk(gclk));
	jdff dff_B_5gaPbxNb7_0(.din(n1224),.dout(w_dff_B_5gaPbxNb7_0),.clk(gclk));
	jdff dff_B_LZUjBD4E1_0(.din(w_dff_B_5gaPbxNb7_0),.dout(w_dff_B_LZUjBD4E1_0),.clk(gclk));
	jdff dff_B_iHCHDIPS1_0(.din(w_dff_B_LZUjBD4E1_0),.dout(w_dff_B_iHCHDIPS1_0),.clk(gclk));
	jdff dff_B_f6Ui00f27_0(.din(w_dff_B_iHCHDIPS1_0),.dout(w_dff_B_f6Ui00f27_0),.clk(gclk));
	jdff dff_B_jAc165sS2_0(.din(w_dff_B_f6Ui00f27_0),.dout(w_dff_B_jAc165sS2_0),.clk(gclk));
	jdff dff_B_smLObfyz5_0(.din(w_dff_B_jAc165sS2_0),.dout(w_dff_B_smLObfyz5_0),.clk(gclk));
	jdff dff_B_Werem8sL7_0(.din(w_dff_B_smLObfyz5_0),.dout(w_dff_B_Werem8sL7_0),.clk(gclk));
	jdff dff_B_49EIEMAo1_0(.din(w_dff_B_Werem8sL7_0),.dout(w_dff_B_49EIEMAo1_0),.clk(gclk));
	jdff dff_B_0mHTzpry5_0(.din(w_dff_B_49EIEMAo1_0),.dout(w_dff_B_0mHTzpry5_0),.clk(gclk));
	jdff dff_B_NqxXKWV73_0(.din(w_dff_B_0mHTzpry5_0),.dout(w_dff_B_NqxXKWV73_0),.clk(gclk));
	jdff dff_B_WBZdrwGk0_0(.din(w_dff_B_NqxXKWV73_0),.dout(w_dff_B_WBZdrwGk0_0),.clk(gclk));
	jdff dff_B_J9pkYxVq4_0(.din(w_dff_B_WBZdrwGk0_0),.dout(w_dff_B_J9pkYxVq4_0),.clk(gclk));
	jdff dff_B_CWM73GqH0_0(.din(w_dff_B_J9pkYxVq4_0),.dout(w_dff_B_CWM73GqH0_0),.clk(gclk));
	jdff dff_B_VYpWjlrd2_0(.din(w_dff_B_CWM73GqH0_0),.dout(w_dff_B_VYpWjlrd2_0),.clk(gclk));
	jdff dff_B_nwXDeyvS8_0(.din(w_dff_B_VYpWjlrd2_0),.dout(w_dff_B_nwXDeyvS8_0),.clk(gclk));
	jdff dff_B_dTt7e69l8_0(.din(w_dff_B_nwXDeyvS8_0),.dout(w_dff_B_dTt7e69l8_0),.clk(gclk));
	jdff dff_B_foFSaU8A0_0(.din(w_dff_B_dTt7e69l8_0),.dout(w_dff_B_foFSaU8A0_0),.clk(gclk));
	jdff dff_B_WQeYJm0f2_0(.din(n1223),.dout(w_dff_B_WQeYJm0f2_0),.clk(gclk));
	jdff dff_B_neDWcCt91_0(.din(n1231),.dout(w_dff_B_neDWcCt91_0),.clk(gclk));
	jdff dff_B_9PRc625b3_0(.din(w_dff_B_neDWcCt91_0),.dout(w_dff_B_9PRc625b3_0),.clk(gclk));
	jdff dff_B_fBhAPvB28_0(.din(w_dff_B_9PRc625b3_0),.dout(w_dff_B_fBhAPvB28_0),.clk(gclk));
	jdff dff_B_LSRApeyK8_0(.din(w_dff_B_fBhAPvB28_0),.dout(w_dff_B_LSRApeyK8_0),.clk(gclk));
	jdff dff_B_p8y7SmDH3_0(.din(w_dff_B_LSRApeyK8_0),.dout(w_dff_B_p8y7SmDH3_0),.clk(gclk));
	jdff dff_B_IIjg4NL32_0(.din(w_dff_B_p8y7SmDH3_0),.dout(w_dff_B_IIjg4NL32_0),.clk(gclk));
	jdff dff_B_pgMHeisA8_0(.din(w_dff_B_IIjg4NL32_0),.dout(w_dff_B_pgMHeisA8_0),.clk(gclk));
	jdff dff_B_tc7Bs2wn5_0(.din(w_dff_B_pgMHeisA8_0),.dout(w_dff_B_tc7Bs2wn5_0),.clk(gclk));
	jdff dff_B_IauBRnPd9_0(.din(w_dff_B_tc7Bs2wn5_0),.dout(w_dff_B_IauBRnPd9_0),.clk(gclk));
	jdff dff_B_YsrTa2460_0(.din(w_dff_B_IauBRnPd9_0),.dout(w_dff_B_YsrTa2460_0),.clk(gclk));
	jdff dff_B_vojdUPDY4_0(.din(w_dff_B_YsrTa2460_0),.dout(w_dff_B_vojdUPDY4_0),.clk(gclk));
	jdff dff_B_g0jx4bv50_0(.din(w_dff_B_vojdUPDY4_0),.dout(w_dff_B_g0jx4bv50_0),.clk(gclk));
	jdff dff_B_Zt4fGQ628_0(.din(w_dff_B_g0jx4bv50_0),.dout(w_dff_B_Zt4fGQ628_0),.clk(gclk));
	jdff dff_B_IJ7dlnse4_0(.din(w_dff_B_Zt4fGQ628_0),.dout(w_dff_B_IJ7dlnse4_0),.clk(gclk));
	jdff dff_B_tFx1AYRP1_0(.din(w_dff_B_IJ7dlnse4_0),.dout(w_dff_B_tFx1AYRP1_0),.clk(gclk));
	jdff dff_B_Bb1YNwW11_0(.din(w_dff_B_tFx1AYRP1_0),.dout(w_dff_B_Bb1YNwW11_0),.clk(gclk));
	jdff dff_B_ZNrBUawd7_0(.din(w_dff_B_Bb1YNwW11_0),.dout(w_dff_B_ZNrBUawd7_0),.clk(gclk));
	jdff dff_B_8rv1HNPK0_0(.din(n1230),.dout(w_dff_B_8rv1HNPK0_0),.clk(gclk));
	jdff dff_B_VJUTrNHT7_2(.din(G106),.dout(w_dff_B_VJUTrNHT7_2),.clk(gclk));
	jdff dff_B_BL3JyIJS4_2(.din(G109),.dout(w_dff_B_BL3JyIJS4_2),.clk(gclk));
	jdff dff_B_LlnZ7Dqk4_2(.din(w_dff_B_BL3JyIJS4_2),.dout(w_dff_B_LlnZ7Dqk4_2),.clk(gclk));
	jdff dff_B_2jIm1a6Y6_0(.din(n1239),.dout(w_dff_B_2jIm1a6Y6_0),.clk(gclk));
	jdff dff_B_4eHGq9aF2_0(.din(w_dff_B_2jIm1a6Y6_0),.dout(w_dff_B_4eHGq9aF2_0),.clk(gclk));
	jdff dff_B_Obs0PbIK9_0(.din(w_dff_B_4eHGq9aF2_0),.dout(w_dff_B_Obs0PbIK9_0),.clk(gclk));
	jdff dff_B_HU9STO0D6_0(.din(w_dff_B_Obs0PbIK9_0),.dout(w_dff_B_HU9STO0D6_0),.clk(gclk));
	jdff dff_B_BOUBNzSk6_0(.din(w_dff_B_HU9STO0D6_0),.dout(w_dff_B_BOUBNzSk6_0),.clk(gclk));
	jdff dff_B_GawIDrEg5_0(.din(w_dff_B_BOUBNzSk6_0),.dout(w_dff_B_GawIDrEg5_0),.clk(gclk));
	jdff dff_B_bK1DZHkL5_0(.din(w_dff_B_GawIDrEg5_0),.dout(w_dff_B_bK1DZHkL5_0),.clk(gclk));
	jdff dff_B_gdrQ4hA06_0(.din(w_dff_B_bK1DZHkL5_0),.dout(w_dff_B_gdrQ4hA06_0),.clk(gclk));
	jdff dff_B_C46Yp5rT9_0(.din(w_dff_B_gdrQ4hA06_0),.dout(w_dff_B_C46Yp5rT9_0),.clk(gclk));
	jdff dff_B_RsQmhCZC4_0(.din(w_dff_B_C46Yp5rT9_0),.dout(w_dff_B_RsQmhCZC4_0),.clk(gclk));
	jdff dff_B_WRs12aCC1_0(.din(w_dff_B_RsQmhCZC4_0),.dout(w_dff_B_WRs12aCC1_0),.clk(gclk));
	jdff dff_B_2FPcrCAD0_0(.din(w_dff_B_WRs12aCC1_0),.dout(w_dff_B_2FPcrCAD0_0),.clk(gclk));
	jdff dff_B_iLdb7h6h5_0(.din(w_dff_B_2FPcrCAD0_0),.dout(w_dff_B_iLdb7h6h5_0),.clk(gclk));
	jdff dff_B_JS5YIbSr7_0(.din(w_dff_B_iLdb7h6h5_0),.dout(w_dff_B_JS5YIbSr7_0),.clk(gclk));
	jdff dff_B_Alg2lQr27_0(.din(w_dff_B_JS5YIbSr7_0),.dout(w_dff_B_Alg2lQr27_0),.clk(gclk));
	jdff dff_B_bexrAVvW0_0(.din(w_dff_B_Alg2lQr27_0),.dout(w_dff_B_bexrAVvW0_0),.clk(gclk));
	jdff dff_B_Wf1pMfSH9_0(.din(n1238),.dout(w_dff_B_Wf1pMfSH9_0),.clk(gclk));
	jdff dff_B_3GoT8bjo8_0(.din(n1248),.dout(w_dff_B_3GoT8bjo8_0),.clk(gclk));
	jdff dff_B_3oHSvQGF6_0(.din(w_dff_B_3GoT8bjo8_0),.dout(w_dff_B_3oHSvQGF6_0),.clk(gclk));
	jdff dff_B_2dd9hNeQ1_0(.din(w_dff_B_3oHSvQGF6_0),.dout(w_dff_B_2dd9hNeQ1_0),.clk(gclk));
	jdff dff_B_FdpjtFuW3_0(.din(w_dff_B_2dd9hNeQ1_0),.dout(w_dff_B_FdpjtFuW3_0),.clk(gclk));
	jdff dff_B_w3V5Omow0_0(.din(w_dff_B_FdpjtFuW3_0),.dout(w_dff_B_w3V5Omow0_0),.clk(gclk));
	jdff dff_B_bINVdSBt0_0(.din(w_dff_B_w3V5Omow0_0),.dout(w_dff_B_bINVdSBt0_0),.clk(gclk));
	jdff dff_B_aunuScad6_0(.din(w_dff_B_bINVdSBt0_0),.dout(w_dff_B_aunuScad6_0),.clk(gclk));
	jdff dff_B_y5HChuQV8_0(.din(w_dff_B_aunuScad6_0),.dout(w_dff_B_y5HChuQV8_0),.clk(gclk));
	jdff dff_B_EuoWpmdw5_0(.din(w_dff_B_y5HChuQV8_0),.dout(w_dff_B_EuoWpmdw5_0),.clk(gclk));
	jdff dff_B_lOIOp8TB2_0(.din(w_dff_B_EuoWpmdw5_0),.dout(w_dff_B_lOIOp8TB2_0),.clk(gclk));
	jdff dff_B_QTrQBzim1_0(.din(w_dff_B_lOIOp8TB2_0),.dout(w_dff_B_QTrQBzim1_0),.clk(gclk));
	jdff dff_B_51ll5nqO0_0(.din(w_dff_B_QTrQBzim1_0),.dout(w_dff_B_51ll5nqO0_0),.clk(gclk));
	jdff dff_B_rtGJoXJ30_0(.din(w_dff_B_51ll5nqO0_0),.dout(w_dff_B_rtGJoXJ30_0),.clk(gclk));
	jdff dff_B_ShkG2wNF7_0(.din(w_dff_B_rtGJoXJ30_0),.dout(w_dff_B_ShkG2wNF7_0),.clk(gclk));
	jdff dff_B_4lzrQbwA2_0(.din(w_dff_B_ShkG2wNF7_0),.dout(w_dff_B_4lzrQbwA2_0),.clk(gclk));
	jdff dff_B_gAKDul2C1_0(.din(w_dff_B_4lzrQbwA2_0),.dout(w_dff_B_gAKDul2C1_0),.clk(gclk));
	jdff dff_B_leJxw7Py9_0(.din(n1247),.dout(w_dff_B_leJxw7Py9_0),.clk(gclk));
	jdff dff_A_sFWHDYan7_2(.dout(w_n797_2[2]),.din(w_dff_A_sFWHDYan7_2),.clk(gclk));
	jdff dff_A_pjgPQuD18_2(.dout(w_n793_2[2]),.din(w_dff_A_pjgPQuD18_2),.clk(gclk));
	jdff dff_B_20x9tGxk2_0(.din(n1257),.dout(w_dff_B_20x9tGxk2_0),.clk(gclk));
	jdff dff_B_y6yL2sl84_0(.din(w_dff_B_20x9tGxk2_0),.dout(w_dff_B_y6yL2sl84_0),.clk(gclk));
	jdff dff_B_8QSHNWlh4_0(.din(w_dff_B_y6yL2sl84_0),.dout(w_dff_B_8QSHNWlh4_0),.clk(gclk));
	jdff dff_B_K9XhQCve7_0(.din(w_dff_B_8QSHNWlh4_0),.dout(w_dff_B_K9XhQCve7_0),.clk(gclk));
	jdff dff_B_JVr4qkUt1_0(.din(w_dff_B_K9XhQCve7_0),.dout(w_dff_B_JVr4qkUt1_0),.clk(gclk));
	jdff dff_B_4iGO9YDx5_0(.din(w_dff_B_JVr4qkUt1_0),.dout(w_dff_B_4iGO9YDx5_0),.clk(gclk));
	jdff dff_B_ADhVyGKw3_0(.din(w_dff_B_4iGO9YDx5_0),.dout(w_dff_B_ADhVyGKw3_0),.clk(gclk));
	jdff dff_B_4U7IAqCH5_0(.din(w_dff_B_ADhVyGKw3_0),.dout(w_dff_B_4U7IAqCH5_0),.clk(gclk));
	jdff dff_B_GcBshYe89_0(.din(w_dff_B_4U7IAqCH5_0),.dout(w_dff_B_GcBshYe89_0),.clk(gclk));
	jdff dff_B_QuHuM2o98_0(.din(w_dff_B_GcBshYe89_0),.dout(w_dff_B_QuHuM2o98_0),.clk(gclk));
	jdff dff_B_jvQLPQR05_0(.din(w_dff_B_QuHuM2o98_0),.dout(w_dff_B_jvQLPQR05_0),.clk(gclk));
	jdff dff_B_DBQzuKY78_0(.din(w_dff_B_jvQLPQR05_0),.dout(w_dff_B_DBQzuKY78_0),.clk(gclk));
	jdff dff_B_KUzCtUsv5_0(.din(w_dff_B_DBQzuKY78_0),.dout(w_dff_B_KUzCtUsv5_0),.clk(gclk));
	jdff dff_B_HAZEoKtx6_0(.din(w_dff_B_KUzCtUsv5_0),.dout(w_dff_B_HAZEoKtx6_0),.clk(gclk));
	jdff dff_B_kbBNPsoE5_0(.din(w_dff_B_HAZEoKtx6_0),.dout(w_dff_B_kbBNPsoE5_0),.clk(gclk));
	jdff dff_B_8wzj2M7N8_0(.din(n1256),.dout(w_dff_B_8wzj2M7N8_0),.clk(gclk));
	jdff dff_B_Sw2dCsV19_0(.din(n1264),.dout(w_dff_B_Sw2dCsV19_0),.clk(gclk));
	jdff dff_B_UO6PmPVD3_0(.din(w_dff_B_Sw2dCsV19_0),.dout(w_dff_B_UO6PmPVD3_0),.clk(gclk));
	jdff dff_B_yhbITnzf3_0(.din(w_dff_B_UO6PmPVD3_0),.dout(w_dff_B_yhbITnzf3_0),.clk(gclk));
	jdff dff_B_aZePPmIH4_0(.din(w_dff_B_yhbITnzf3_0),.dout(w_dff_B_aZePPmIH4_0),.clk(gclk));
	jdff dff_B_jrpvn6094_0(.din(w_dff_B_aZePPmIH4_0),.dout(w_dff_B_jrpvn6094_0),.clk(gclk));
	jdff dff_B_GsUGTxeN9_0(.din(w_dff_B_jrpvn6094_0),.dout(w_dff_B_GsUGTxeN9_0),.clk(gclk));
	jdff dff_B_o94m2jSD3_0(.din(w_dff_B_GsUGTxeN9_0),.dout(w_dff_B_o94m2jSD3_0),.clk(gclk));
	jdff dff_B_fk177KwR8_0(.din(w_dff_B_o94m2jSD3_0),.dout(w_dff_B_fk177KwR8_0),.clk(gclk));
	jdff dff_B_kcVxM77C7_0(.din(w_dff_B_fk177KwR8_0),.dout(w_dff_B_kcVxM77C7_0),.clk(gclk));
	jdff dff_B_kW3zZLNS6_0(.din(w_dff_B_kcVxM77C7_0),.dout(w_dff_B_kW3zZLNS6_0),.clk(gclk));
	jdff dff_B_XGvfQ2Gc5_0(.din(w_dff_B_kW3zZLNS6_0),.dout(w_dff_B_XGvfQ2Gc5_0),.clk(gclk));
	jdff dff_B_R4JQJ6dt9_0(.din(w_dff_B_XGvfQ2Gc5_0),.dout(w_dff_B_R4JQJ6dt9_0),.clk(gclk));
	jdff dff_B_WXwKa3HZ3_0(.din(w_dff_B_R4JQJ6dt9_0),.dout(w_dff_B_WXwKa3HZ3_0),.clk(gclk));
	jdff dff_B_L102BejT7_0(.din(w_dff_B_WXwKa3HZ3_0),.dout(w_dff_B_L102BejT7_0),.clk(gclk));
	jdff dff_B_zS322e1s8_0(.din(w_dff_B_L102BejT7_0),.dout(w_dff_B_zS322e1s8_0),.clk(gclk));
	jdff dff_B_OeaKwgd32_0(.din(w_dff_B_zS322e1s8_0),.dout(w_dff_B_OeaKwgd32_0),.clk(gclk));
	jdff dff_B_EykvKAbE6_0(.din(n1263),.dout(w_dff_B_EykvKAbE6_0),.clk(gclk));
	jdff dff_B_VMkJNZAT8_2(.din(G49),.dout(w_dff_B_VMkJNZAT8_2),.clk(gclk));
	jdff dff_B_id5mtwnl2_2(.din(G46),.dout(w_dff_B_id5mtwnl2_2),.clk(gclk));
	jdff dff_B_CWb2MDZp4_2(.din(w_dff_B_id5mtwnl2_2),.dout(w_dff_B_CWb2MDZp4_2),.clk(gclk));
	jdff dff_B_gl2MfgDg6_0(.din(n1271),.dout(w_dff_B_gl2MfgDg6_0),.clk(gclk));
	jdff dff_B_By8RYdoW4_0(.din(w_dff_B_gl2MfgDg6_0),.dout(w_dff_B_By8RYdoW4_0),.clk(gclk));
	jdff dff_B_kHZhQ3vZ7_0(.din(w_dff_B_By8RYdoW4_0),.dout(w_dff_B_kHZhQ3vZ7_0),.clk(gclk));
	jdff dff_B_LywzKnL92_0(.din(w_dff_B_kHZhQ3vZ7_0),.dout(w_dff_B_LywzKnL92_0),.clk(gclk));
	jdff dff_B_BfgtXapc5_0(.din(w_dff_B_LywzKnL92_0),.dout(w_dff_B_BfgtXapc5_0),.clk(gclk));
	jdff dff_B_TpSRZBrM4_0(.din(w_dff_B_BfgtXapc5_0),.dout(w_dff_B_TpSRZBrM4_0),.clk(gclk));
	jdff dff_B_3zPE5ibu4_0(.din(w_dff_B_TpSRZBrM4_0),.dout(w_dff_B_3zPE5ibu4_0),.clk(gclk));
	jdff dff_B_RxqksCYE5_0(.din(w_dff_B_3zPE5ibu4_0),.dout(w_dff_B_RxqksCYE5_0),.clk(gclk));
	jdff dff_B_PeCSNeRq8_0(.din(w_dff_B_RxqksCYE5_0),.dout(w_dff_B_PeCSNeRq8_0),.clk(gclk));
	jdff dff_B_Wx5yXMqj3_0(.din(w_dff_B_PeCSNeRq8_0),.dout(w_dff_B_Wx5yXMqj3_0),.clk(gclk));
	jdff dff_B_clMW8Zes3_0(.din(w_dff_B_Wx5yXMqj3_0),.dout(w_dff_B_clMW8Zes3_0),.clk(gclk));
	jdff dff_B_1cntyA2A5_0(.din(w_dff_B_clMW8Zes3_0),.dout(w_dff_B_1cntyA2A5_0),.clk(gclk));
	jdff dff_B_kF3Pzrva1_0(.din(w_dff_B_1cntyA2A5_0),.dout(w_dff_B_kF3Pzrva1_0),.clk(gclk));
	jdff dff_B_Ijqvewyn4_0(.din(w_dff_B_kF3Pzrva1_0),.dout(w_dff_B_Ijqvewyn4_0),.clk(gclk));
	jdff dff_B_PCNzElJv1_0(.din(w_dff_B_Ijqvewyn4_0),.dout(w_dff_B_PCNzElJv1_0),.clk(gclk));
	jdff dff_B_gqepe3so4_0(.din(w_dff_B_PCNzElJv1_0),.dout(w_dff_B_gqepe3so4_0),.clk(gclk));
	jdff dff_B_TUIbUdjG8_0(.din(n1270),.dout(w_dff_B_TUIbUdjG8_0),.clk(gclk));
	jdff dff_B_XnPH5e6I5_2(.din(G103),.dout(w_dff_B_XnPH5e6I5_2),.clk(gclk));
	jdff dff_B_U5rumXto4_2(.din(G100),.dout(w_dff_B_U5rumXto4_2),.clk(gclk));
	jdff dff_B_dCjbwhYg7_2(.din(w_dff_B_U5rumXto4_2),.dout(w_dff_B_dCjbwhYg7_2),.clk(gclk));
	jdff dff_A_SmbNmyt81_2(.dout(w_n843_2[2]),.din(w_dff_A_SmbNmyt81_2),.clk(gclk));
	jdff dff_A_Hz1qLP2O7_2(.dout(w_n840_2[2]),.din(w_dff_A_Hz1qLP2O7_2),.clk(gclk));
	jdff dff_B_p2Cx5lnN1_0(.din(n1278),.dout(w_dff_B_p2Cx5lnN1_0),.clk(gclk));
	jdff dff_B_cxMWjz5X1_0(.din(w_dff_B_p2Cx5lnN1_0),.dout(w_dff_B_cxMWjz5X1_0),.clk(gclk));
	jdff dff_B_ASmHS2gG4_0(.din(w_dff_B_cxMWjz5X1_0),.dout(w_dff_B_ASmHS2gG4_0),.clk(gclk));
	jdff dff_B_Gr4XG9np8_0(.din(w_dff_B_ASmHS2gG4_0),.dout(w_dff_B_Gr4XG9np8_0),.clk(gclk));
	jdff dff_B_oTwodoID6_0(.din(w_dff_B_Gr4XG9np8_0),.dout(w_dff_B_oTwodoID6_0),.clk(gclk));
	jdff dff_B_Zmo8yTop6_0(.din(w_dff_B_oTwodoID6_0),.dout(w_dff_B_Zmo8yTop6_0),.clk(gclk));
	jdff dff_B_Vift5rqO8_0(.din(w_dff_B_Zmo8yTop6_0),.dout(w_dff_B_Vift5rqO8_0),.clk(gclk));
	jdff dff_B_aMnyNwJM8_0(.din(w_dff_B_Vift5rqO8_0),.dout(w_dff_B_aMnyNwJM8_0),.clk(gclk));
	jdff dff_B_EjvB9dRC0_0(.din(w_dff_B_aMnyNwJM8_0),.dout(w_dff_B_EjvB9dRC0_0),.clk(gclk));
	jdff dff_B_3XYKE3Vl7_0(.din(w_dff_B_EjvB9dRC0_0),.dout(w_dff_B_3XYKE3Vl7_0),.clk(gclk));
	jdff dff_B_SxJqGZvK2_0(.din(w_dff_B_3XYKE3Vl7_0),.dout(w_dff_B_SxJqGZvK2_0),.clk(gclk));
	jdff dff_B_DZXUIWvj3_0(.din(w_dff_B_SxJqGZvK2_0),.dout(w_dff_B_DZXUIWvj3_0),.clk(gclk));
	jdff dff_B_I3htXaNh3_0(.din(w_dff_B_DZXUIWvj3_0),.dout(w_dff_B_I3htXaNh3_0),.clk(gclk));
	jdff dff_B_j5zEbwX24_0(.din(w_dff_B_I3htXaNh3_0),.dout(w_dff_B_j5zEbwX24_0),.clk(gclk));
	jdff dff_B_k1BaaJBX6_0(.din(w_dff_B_j5zEbwX24_0),.dout(w_dff_B_k1BaaJBX6_0),.clk(gclk));
	jdff dff_B_O0tS13sh8_0(.din(n1277),.dout(w_dff_B_O0tS13sh8_0),.clk(gclk));
	jdff dff_B_Mo8eHblO3_2(.din(G40),.dout(w_dff_B_Mo8eHblO3_2),.clk(gclk));
	jdff dff_B_gjtDFMWi6_2(.din(G91),.dout(w_dff_B_gjtDFMWi6_2),.clk(gclk));
	jdff dff_B_el6Qlaq36_2(.din(w_dff_B_gjtDFMWi6_2),.dout(w_dff_B_el6Qlaq36_2),.clk(gclk));
	jdff dff_B_YlXyAUM25_0(.din(n1285),.dout(w_dff_B_YlXyAUM25_0),.clk(gclk));
	jdff dff_B_aVj4Kkp72_0(.din(w_dff_B_YlXyAUM25_0),.dout(w_dff_B_aVj4Kkp72_0),.clk(gclk));
	jdff dff_B_yq5DeBgq9_0(.din(w_dff_B_aVj4Kkp72_0),.dout(w_dff_B_yq5DeBgq9_0),.clk(gclk));
	jdff dff_B_sEJqdaGv0_0(.din(w_dff_B_yq5DeBgq9_0),.dout(w_dff_B_sEJqdaGv0_0),.clk(gclk));
	jdff dff_B_GLVIhucX2_0(.din(w_dff_B_sEJqdaGv0_0),.dout(w_dff_B_GLVIhucX2_0),.clk(gclk));
	jdff dff_B_o72YPEzF5_0(.din(w_dff_B_GLVIhucX2_0),.dout(w_dff_B_o72YPEzF5_0),.clk(gclk));
	jdff dff_B_jw7iBpqr7_0(.din(w_dff_B_o72YPEzF5_0),.dout(w_dff_B_jw7iBpqr7_0),.clk(gclk));
	jdff dff_B_NzQpgOY98_0(.din(w_dff_B_jw7iBpqr7_0),.dout(w_dff_B_NzQpgOY98_0),.clk(gclk));
	jdff dff_B_De4INmgk8_0(.din(w_dff_B_NzQpgOY98_0),.dout(w_dff_B_De4INmgk8_0),.clk(gclk));
	jdff dff_B_gXtEZGjE4_0(.din(w_dff_B_De4INmgk8_0),.dout(w_dff_B_gXtEZGjE4_0),.clk(gclk));
	jdff dff_B_eXUOmbkv6_0(.din(w_dff_B_gXtEZGjE4_0),.dout(w_dff_B_eXUOmbkv6_0),.clk(gclk));
	jdff dff_B_pc9SxJp39_0(.din(w_dff_B_eXUOmbkv6_0),.dout(w_dff_B_pc9SxJp39_0),.clk(gclk));
	jdff dff_B_HVwaOk6v1_0(.din(w_dff_B_pc9SxJp39_0),.dout(w_dff_B_HVwaOk6v1_0),.clk(gclk));
	jdff dff_B_FAtq4dTe0_0(.din(w_dff_B_HVwaOk6v1_0),.dout(w_dff_B_FAtq4dTe0_0),.clk(gclk));
	jdff dff_B_qH4ghL7g7_0(.din(w_dff_B_FAtq4dTe0_0),.dout(w_dff_B_qH4ghL7g7_0),.clk(gclk));
	jdff dff_B_ATcF3x672_0(.din(n1284),.dout(w_dff_B_ATcF3x672_0),.clk(gclk));
	jdff dff_A_P1d707Og2_0(.dout(w_G137_6[0]),.din(w_dff_A_P1d707Og2_0),.clk(gclk));
	jdff dff_A_i0nhRt9V4_0(.dout(w_dff_A_P1d707Og2_0),.din(w_dff_A_i0nhRt9V4_0),.clk(gclk));
	jdff dff_A_5z3ezwth3_0(.dout(w_dff_A_i0nhRt9V4_0),.din(w_dff_A_5z3ezwth3_0),.clk(gclk));
	jdff dff_A_zyfe1BjJ8_0(.dout(w_dff_A_5z3ezwth3_0),.din(w_dff_A_zyfe1BjJ8_0),.clk(gclk));
	jdff dff_A_hwg82l3u4_0(.dout(w_dff_A_zyfe1BjJ8_0),.din(w_dff_A_hwg82l3u4_0),.clk(gclk));
	jdff dff_A_6cW6CQ4E5_1(.dout(w_G137_6[1]),.din(w_dff_A_6cW6CQ4E5_1),.clk(gclk));
	jdff dff_B_YNCVFuse0_0(.din(n1293),.dout(w_dff_B_YNCVFuse0_0),.clk(gclk));
	jdff dff_B_xN5Dk6JH0_0(.din(w_dff_B_YNCVFuse0_0),.dout(w_dff_B_xN5Dk6JH0_0),.clk(gclk));
	jdff dff_B_QgUyiywD0_0(.din(w_dff_B_xN5Dk6JH0_0),.dout(w_dff_B_QgUyiywD0_0),.clk(gclk));
	jdff dff_B_F0e6Rtjo2_0(.din(w_dff_B_QgUyiywD0_0),.dout(w_dff_B_F0e6Rtjo2_0),.clk(gclk));
	jdff dff_B_o1fgI3in6_0(.din(w_dff_B_F0e6Rtjo2_0),.dout(w_dff_B_o1fgI3in6_0),.clk(gclk));
	jdff dff_B_BEmcUTEZ6_0(.din(w_dff_B_o1fgI3in6_0),.dout(w_dff_B_BEmcUTEZ6_0),.clk(gclk));
	jdff dff_B_Ujy3i7h34_0(.din(w_dff_B_BEmcUTEZ6_0),.dout(w_dff_B_Ujy3i7h34_0),.clk(gclk));
	jdff dff_B_VmXc9wwG0_0(.din(w_dff_B_Ujy3i7h34_0),.dout(w_dff_B_VmXc9wwG0_0),.clk(gclk));
	jdff dff_B_mY58C45M5_0(.din(w_dff_B_VmXc9wwG0_0),.dout(w_dff_B_mY58C45M5_0),.clk(gclk));
	jdff dff_B_ZOYtNVIT5_0(.din(w_dff_B_mY58C45M5_0),.dout(w_dff_B_ZOYtNVIT5_0),.clk(gclk));
	jdff dff_B_op6k6ob95_0(.din(w_dff_B_ZOYtNVIT5_0),.dout(w_dff_B_op6k6ob95_0),.clk(gclk));
	jdff dff_B_VD1RIM4u9_0(.din(w_dff_B_op6k6ob95_0),.dout(w_dff_B_VD1RIM4u9_0),.clk(gclk));
	jdff dff_B_K6oArLI90_0(.din(w_dff_B_VD1RIM4u9_0),.dout(w_dff_B_K6oArLI90_0),.clk(gclk));
	jdff dff_B_cxOX2idm5_0(.din(w_dff_B_K6oArLI90_0),.dout(w_dff_B_cxOX2idm5_0),.clk(gclk));
	jdff dff_B_lSPkGAlU4_0(.din(w_dff_B_cxOX2idm5_0),.dout(w_dff_B_lSPkGAlU4_0),.clk(gclk));
	jdff dff_B_M3NHt4gJ0_0(.din(w_dff_B_lSPkGAlU4_0),.dout(w_dff_B_M3NHt4gJ0_0),.clk(gclk));
	jdff dff_B_QiyBP5GP1_0(.din(n1292),.dout(w_dff_B_QiyBP5GP1_0),.clk(gclk));
	jdff dff_B_4msxmbml3_0(.din(n1301),.dout(w_dff_B_4msxmbml3_0),.clk(gclk));
	jdff dff_B_zT7HkHPO6_0(.din(w_dff_B_4msxmbml3_0),.dout(w_dff_B_zT7HkHPO6_0),.clk(gclk));
	jdff dff_B_IRW2hMpD2_0(.din(w_dff_B_zT7HkHPO6_0),.dout(w_dff_B_IRW2hMpD2_0),.clk(gclk));
	jdff dff_B_LkrIOcYJ0_0(.din(w_dff_B_IRW2hMpD2_0),.dout(w_dff_B_LkrIOcYJ0_0),.clk(gclk));
	jdff dff_B_aIZyJHXx4_0(.din(w_dff_B_LkrIOcYJ0_0),.dout(w_dff_B_aIZyJHXx4_0),.clk(gclk));
	jdff dff_B_UhoOIOAq9_0(.din(w_dff_B_aIZyJHXx4_0),.dout(w_dff_B_UhoOIOAq9_0),.clk(gclk));
	jdff dff_B_ng5hXrky7_0(.din(w_dff_B_UhoOIOAq9_0),.dout(w_dff_B_ng5hXrky7_0),.clk(gclk));
	jdff dff_B_TAghHFYQ5_0(.din(w_dff_B_ng5hXrky7_0),.dout(w_dff_B_TAghHFYQ5_0),.clk(gclk));
	jdff dff_B_5ha3oELz4_0(.din(w_dff_B_TAghHFYQ5_0),.dout(w_dff_B_5ha3oELz4_0),.clk(gclk));
	jdff dff_B_PlyUo6wp5_0(.din(w_dff_B_5ha3oELz4_0),.dout(w_dff_B_PlyUo6wp5_0),.clk(gclk));
	jdff dff_B_yIo92Wkk0_0(.din(w_dff_B_PlyUo6wp5_0),.dout(w_dff_B_yIo92Wkk0_0),.clk(gclk));
	jdff dff_B_P2y9kksI0_0(.din(w_dff_B_yIo92Wkk0_0),.dout(w_dff_B_P2y9kksI0_0),.clk(gclk));
	jdff dff_B_bOuWH4Eb6_0(.din(w_dff_B_P2y9kksI0_0),.dout(w_dff_B_bOuWH4Eb6_0),.clk(gclk));
	jdff dff_B_OdQbqyHw6_0(.din(w_dff_B_bOuWH4Eb6_0),.dout(w_dff_B_OdQbqyHw6_0),.clk(gclk));
	jdff dff_B_t6jvK84v4_0(.din(w_dff_B_OdQbqyHw6_0),.dout(w_dff_B_t6jvK84v4_0),.clk(gclk));
	jdff dff_B_3harrfKT3_0(.din(w_dff_B_t6jvK84v4_0),.dout(w_dff_B_3harrfKT3_0),.clk(gclk));
	jdff dff_B_utLN8AQu0_0(.din(n1300),.dout(w_dff_B_utLN8AQu0_0),.clk(gclk));
	jdff dff_A_kniqA7ph3_0(.dout(w_n988_2[0]),.din(w_dff_A_kniqA7ph3_0),.clk(gclk));
	jdff dff_A_9abkvoqm3_1(.dout(w_n988_2[1]),.din(w_dff_A_9abkvoqm3_1),.clk(gclk));
	jdff dff_A_tC8auo9X0_0(.dout(w_n985_2[0]),.din(w_dff_A_tC8auo9X0_0),.clk(gclk));
	jdff dff_A_JLEfot5E1_1(.dout(w_n985_2[1]),.din(w_dff_A_JLEfot5E1_1),.clk(gclk));
	jdff dff_B_k8f7HUkw4_0(.din(n1309),.dout(w_dff_B_k8f7HUkw4_0),.clk(gclk));
	jdff dff_B_XXqDlLwL6_0(.din(w_dff_B_k8f7HUkw4_0),.dout(w_dff_B_XXqDlLwL6_0),.clk(gclk));
	jdff dff_B_InhiICYY6_0(.din(w_dff_B_XXqDlLwL6_0),.dout(w_dff_B_InhiICYY6_0),.clk(gclk));
	jdff dff_B_reJt5BAK4_0(.din(w_dff_B_InhiICYY6_0),.dout(w_dff_B_reJt5BAK4_0),.clk(gclk));
	jdff dff_B_2RNbhanw1_0(.din(w_dff_B_reJt5BAK4_0),.dout(w_dff_B_2RNbhanw1_0),.clk(gclk));
	jdff dff_B_5HpS8KsX8_0(.din(w_dff_B_2RNbhanw1_0),.dout(w_dff_B_5HpS8KsX8_0),.clk(gclk));
	jdff dff_B_udvZJu4k1_0(.din(w_dff_B_5HpS8KsX8_0),.dout(w_dff_B_udvZJu4k1_0),.clk(gclk));
	jdff dff_B_p9dWWpY59_0(.din(w_dff_B_udvZJu4k1_0),.dout(w_dff_B_p9dWWpY59_0),.clk(gclk));
	jdff dff_B_GJIH3AXz6_0(.din(w_dff_B_p9dWWpY59_0),.dout(w_dff_B_GJIH3AXz6_0),.clk(gclk));
	jdff dff_B_HOEg0NhJ5_0(.din(w_dff_B_GJIH3AXz6_0),.dout(w_dff_B_HOEg0NhJ5_0),.clk(gclk));
	jdff dff_B_pIsb6NzU4_0(.din(w_dff_B_HOEg0NhJ5_0),.dout(w_dff_B_pIsb6NzU4_0),.clk(gclk));
	jdff dff_B_5VbBwoJ82_0(.din(w_dff_B_pIsb6NzU4_0),.dout(w_dff_B_5VbBwoJ82_0),.clk(gclk));
	jdff dff_B_lugxgPWM9_0(.din(w_dff_B_5VbBwoJ82_0),.dout(w_dff_B_lugxgPWM9_0),.clk(gclk));
	jdff dff_B_U8AA5nKf2_0(.din(w_dff_B_lugxgPWM9_0),.dout(w_dff_B_U8AA5nKf2_0),.clk(gclk));
	jdff dff_B_fAEC05d99_0(.din(w_dff_B_U8AA5nKf2_0),.dout(w_dff_B_fAEC05d99_0),.clk(gclk));
	jdff dff_B_AfURZYz12_0(.din(w_dff_B_fAEC05d99_0),.dout(w_dff_B_AfURZYz12_0),.clk(gclk));
	jdff dff_B_5tYYOmDO1_0(.din(w_dff_B_AfURZYz12_0),.dout(w_dff_B_5tYYOmDO1_0),.clk(gclk));
	jdff dff_B_GkzyK1x01_0(.din(n1308),.dout(w_dff_B_GkzyK1x01_0),.clk(gclk));
	jdff dff_A_a3Hw78NH0_0(.dout(w_G137_5[0]),.din(w_dff_A_a3Hw78NH0_0),.clk(gclk));
	jdff dff_B_12U1LPE12_0(.din(n1317),.dout(w_dff_B_12U1LPE12_0),.clk(gclk));
	jdff dff_B_KboSwyh90_0(.din(w_dff_B_12U1LPE12_0),.dout(w_dff_B_KboSwyh90_0),.clk(gclk));
	jdff dff_B_lkw6DABr2_0(.din(w_dff_B_KboSwyh90_0),.dout(w_dff_B_lkw6DABr2_0),.clk(gclk));
	jdff dff_B_Ujyp9KRj3_0(.din(w_dff_B_lkw6DABr2_0),.dout(w_dff_B_Ujyp9KRj3_0),.clk(gclk));
	jdff dff_B_XYuEFKGi6_0(.din(w_dff_B_Ujyp9KRj3_0),.dout(w_dff_B_XYuEFKGi6_0),.clk(gclk));
	jdff dff_B_2mBpvFFB1_0(.din(w_dff_B_XYuEFKGi6_0),.dout(w_dff_B_2mBpvFFB1_0),.clk(gclk));
	jdff dff_B_kiAnCau14_0(.din(w_dff_B_2mBpvFFB1_0),.dout(w_dff_B_kiAnCau14_0),.clk(gclk));
	jdff dff_B_gLUmyhuQ8_0(.din(w_dff_B_kiAnCau14_0),.dout(w_dff_B_gLUmyhuQ8_0),.clk(gclk));
	jdff dff_B_vuir9hZV3_0(.din(w_dff_B_gLUmyhuQ8_0),.dout(w_dff_B_vuir9hZV3_0),.clk(gclk));
	jdff dff_B_iSZ1uR1d2_0(.din(w_dff_B_vuir9hZV3_0),.dout(w_dff_B_iSZ1uR1d2_0),.clk(gclk));
	jdff dff_B_Qdk5EYEE6_0(.din(w_dff_B_iSZ1uR1d2_0),.dout(w_dff_B_Qdk5EYEE6_0),.clk(gclk));
	jdff dff_B_Bzp7SjmF5_0(.din(w_dff_B_Qdk5EYEE6_0),.dout(w_dff_B_Bzp7SjmF5_0),.clk(gclk));
	jdff dff_B_iC0h8nva9_0(.din(w_dff_B_Bzp7SjmF5_0),.dout(w_dff_B_iC0h8nva9_0),.clk(gclk));
	jdff dff_B_bRY6WnYk0_0(.din(w_dff_B_iC0h8nva9_0),.dout(w_dff_B_bRY6WnYk0_0),.clk(gclk));
	jdff dff_B_cvumRequ5_0(.din(w_dff_B_bRY6WnYk0_0),.dout(w_dff_B_cvumRequ5_0),.clk(gclk));
	jdff dff_B_MjGKjvwP7_0(.din(n1316),.dout(w_dff_B_MjGKjvwP7_0),.clk(gclk));
	jdff dff_B_SurJZRrC4_2(.din(G173),.dout(w_dff_B_SurJZRrC4_2),.clk(gclk));
	jdff dff_B_p7Wfqv4N3_2(.din(G203),.dout(w_dff_B_p7Wfqv4N3_2),.clk(gclk));
	jdff dff_B_hcqlBw8G8_2(.din(w_dff_B_p7Wfqv4N3_2),.dout(w_dff_B_hcqlBw8G8_2),.clk(gclk));
	jdff dff_B_w7B4ucgx9_0(.din(n1182),.dout(w_dff_B_w7B4ucgx9_0),.clk(gclk));
	jdff dff_B_7VQL5rZ74_0(.din(w_dff_B_w7B4ucgx9_0),.dout(w_dff_B_7VQL5rZ74_0),.clk(gclk));
	jdff dff_B_S9c7Ccw26_0(.din(w_dff_B_7VQL5rZ74_0),.dout(w_dff_B_S9c7Ccw26_0),.clk(gclk));
	jdff dff_B_QNNNQo5B6_0(.din(w_dff_B_S9c7Ccw26_0),.dout(w_dff_B_QNNNQo5B6_0),.clk(gclk));
	jdff dff_B_GkqvVYFW1_0(.din(w_dff_B_QNNNQo5B6_0),.dout(w_dff_B_GkqvVYFW1_0),.clk(gclk));
	jdff dff_B_7gm4x91E5_0(.din(w_dff_B_GkqvVYFW1_0),.dout(w_dff_B_7gm4x91E5_0),.clk(gclk));
	jdff dff_B_H2oYONkY2_0(.din(w_dff_B_7gm4x91E5_0),.dout(w_dff_B_H2oYONkY2_0),.clk(gclk));
	jdff dff_B_Ssvhphfd4_0(.din(w_dff_B_H2oYONkY2_0),.dout(w_dff_B_Ssvhphfd4_0),.clk(gclk));
	jdff dff_B_Z8qSrzYS1_0(.din(w_dff_B_Ssvhphfd4_0),.dout(w_dff_B_Z8qSrzYS1_0),.clk(gclk));
	jdff dff_B_q2OBw3WY3_0(.din(n1181),.dout(w_dff_B_q2OBw3WY3_0),.clk(gclk));
	jdff dff_B_rFDNt3jY9_0(.din(w_dff_B_q2OBw3WY3_0),.dout(w_dff_B_rFDNt3jY9_0),.clk(gclk));
	jdff dff_B_bdJBNayM5_1(.din(G112),.dout(w_dff_B_bdJBNayM5_1),.clk(gclk));
	jdff dff_B_ITDwAj4G9_1(.din(w_dff_B_bdJBNayM5_1),.dout(w_dff_B_ITDwAj4G9_1),.clk(gclk));
	jdff dff_B_E8g3QzHa4_0(.din(n1218),.dout(w_dff_B_E8g3QzHa4_0),.clk(gclk));
	jdff dff_B_lqrPEihh4_0(.din(w_dff_B_E8g3QzHa4_0),.dout(w_dff_B_lqrPEihh4_0),.clk(gclk));
	jdff dff_B_jmxu1wD30_0(.din(w_dff_B_lqrPEihh4_0),.dout(w_dff_B_jmxu1wD30_0),.clk(gclk));
	jdff dff_B_TkLFjQNn8_0(.din(w_dff_B_jmxu1wD30_0),.dout(w_dff_B_TkLFjQNn8_0),.clk(gclk));
	jdff dff_B_fc0m9S6j5_0(.din(w_dff_B_TkLFjQNn8_0),.dout(w_dff_B_fc0m9S6j5_0),.clk(gclk));
	jdff dff_B_Zki4KhR49_0(.din(w_dff_B_fc0m9S6j5_0),.dout(w_dff_B_Zki4KhR49_0),.clk(gclk));
	jdff dff_B_HYYn7Udg2_0(.din(w_dff_B_Zki4KhR49_0),.dout(w_dff_B_HYYn7Udg2_0),.clk(gclk));
	jdff dff_B_J2lMJmb59_0(.din(w_dff_B_HYYn7Udg2_0),.dout(w_dff_B_J2lMJmb59_0),.clk(gclk));
	jdff dff_B_ixx83PVO8_0(.din(w_dff_B_J2lMJmb59_0),.dout(w_dff_B_ixx83PVO8_0),.clk(gclk));
	jdff dff_B_CoRr7QPr6_0(.din(w_dff_B_ixx83PVO8_0),.dout(w_dff_B_CoRr7QPr6_0),.clk(gclk));
	jdff dff_B_WqfnwOen3_0(.din(n1217),.dout(w_dff_B_WqfnwOen3_0),.clk(gclk));
	jdff dff_B_D0xwtLV79_0(.din(w_dff_B_WqfnwOen3_0),.dout(w_dff_B_D0xwtLV79_0),.clk(gclk));
	jdff dff_B_LEUCKzil8_1(.din(G113),.dout(w_dff_B_LEUCKzil8_1),.clk(gclk));
	jdff dff_B_cJA6FlcG8_1(.din(w_dff_B_LEUCKzil8_1),.dout(w_dff_B_cJA6FlcG8_1),.clk(gclk));
	jdff dff_B_4nckjkxE7_0(.din(n539),.dout(w_dff_B_4nckjkxE7_0),.clk(gclk));
	jdff dff_B_uOxuyozF6_1(.din(n531),.dout(w_dff_B_uOxuyozF6_1),.clk(gclk));
	jdff dff_B_I4KrkMhc7_0(.din(n1325),.dout(w_dff_B_I4KrkMhc7_0),.clk(gclk));
	jdff dff_B_HS4BqWTz7_0(.din(w_dff_B_I4KrkMhc7_0),.dout(w_dff_B_HS4BqWTz7_0),.clk(gclk));
	jdff dff_B_5akhSlJ55_0(.din(w_dff_B_HS4BqWTz7_0),.dout(w_dff_B_5akhSlJ55_0),.clk(gclk));
	jdff dff_B_HMaARgkk1_0(.din(w_dff_B_5akhSlJ55_0),.dout(w_dff_B_HMaARgkk1_0),.clk(gclk));
	jdff dff_B_fT54kYaw2_0(.din(w_dff_B_HMaARgkk1_0),.dout(w_dff_B_fT54kYaw2_0),.clk(gclk));
	jdff dff_B_Tb9HEADJ3_0(.din(w_dff_B_fT54kYaw2_0),.dout(w_dff_B_Tb9HEADJ3_0),.clk(gclk));
	jdff dff_B_iCdtjdEr4_0(.din(w_dff_B_Tb9HEADJ3_0),.dout(w_dff_B_iCdtjdEr4_0),.clk(gclk));
	jdff dff_B_aIP1Qrtr9_0(.din(w_dff_B_iCdtjdEr4_0),.dout(w_dff_B_aIP1Qrtr9_0),.clk(gclk));
	jdff dff_B_xyU3yWxr2_0(.din(w_dff_B_aIP1Qrtr9_0),.dout(w_dff_B_xyU3yWxr2_0),.clk(gclk));
	jdff dff_B_Bg74AEqj0_0(.din(w_dff_B_xyU3yWxr2_0),.dout(w_dff_B_Bg74AEqj0_0),.clk(gclk));
	jdff dff_B_PQ5jmQuJ6_0(.din(w_dff_B_Bg74AEqj0_0),.dout(w_dff_B_PQ5jmQuJ6_0),.clk(gclk));
	jdff dff_B_5r3plSjt2_0(.din(w_dff_B_PQ5jmQuJ6_0),.dout(w_dff_B_5r3plSjt2_0),.clk(gclk));
	jdff dff_B_YHPm9qSs4_0(.din(w_dff_B_5r3plSjt2_0),.dout(w_dff_B_YHPm9qSs4_0),.clk(gclk));
	jdff dff_B_ajDbJ6IJ9_0(.din(w_dff_B_YHPm9qSs4_0),.dout(w_dff_B_ajDbJ6IJ9_0),.clk(gclk));
	jdff dff_B_nOP5mOmz5_0(.din(w_dff_B_ajDbJ6IJ9_0),.dout(w_dff_B_nOP5mOmz5_0),.clk(gclk));
	jdff dff_B_7xflPzTx9_0(.din(w_dff_B_nOP5mOmz5_0),.dout(w_dff_B_7xflPzTx9_0),.clk(gclk));
	jdff dff_B_Nh4RGfHi0_0(.din(n1324),.dout(w_dff_B_Nh4RGfHi0_0),.clk(gclk));
	jdff dff_B_HwkqESHD8_2(.din(G167),.dout(w_dff_B_HwkqESHD8_2),.clk(gclk));
	jdff dff_B_I8wy6ybV9_2(.din(G197),.dout(w_dff_B_I8wy6ybV9_2),.clk(gclk));
	jdff dff_B_xpzfz9bn8_2(.din(w_dff_B_I8wy6ybV9_2),.dout(w_dff_B_xpzfz9bn8_2),.clk(gclk));
	jdff dff_B_pGEWszLa2_0(.din(n1175),.dout(w_dff_B_pGEWszLa2_0),.clk(gclk));
	jdff dff_B_70mbkrCG6_0(.din(w_dff_B_pGEWszLa2_0),.dout(w_dff_B_70mbkrCG6_0),.clk(gclk));
	jdff dff_B_82aZFgDR1_0(.din(w_dff_B_70mbkrCG6_0),.dout(w_dff_B_82aZFgDR1_0),.clk(gclk));
	jdff dff_B_l3VHYHKN3_0(.din(w_dff_B_82aZFgDR1_0),.dout(w_dff_B_l3VHYHKN3_0),.clk(gclk));
	jdff dff_B_SqEKtrOP0_0(.din(w_dff_B_l3VHYHKN3_0),.dout(w_dff_B_SqEKtrOP0_0),.clk(gclk));
	jdff dff_B_vnhBaksL6_0(.din(w_dff_B_SqEKtrOP0_0),.dout(w_dff_B_vnhBaksL6_0),.clk(gclk));
	jdff dff_B_I5EIZfyO6_0(.din(w_dff_B_vnhBaksL6_0),.dout(w_dff_B_I5EIZfyO6_0),.clk(gclk));
	jdff dff_B_rjIdWvdH7_0(.din(w_dff_B_I5EIZfyO6_0),.dout(w_dff_B_rjIdWvdH7_0),.clk(gclk));
	jdff dff_B_YxpToVNN0_0(.din(w_dff_B_rjIdWvdH7_0),.dout(w_dff_B_YxpToVNN0_0),.clk(gclk));
	jdff dff_B_brMOSBEK6_0(.din(w_dff_B_YxpToVNN0_0),.dout(w_dff_B_brMOSBEK6_0),.clk(gclk));
	jdff dff_B_lqayjOb33_0(.din(n1174),.dout(w_dff_B_lqayjOb33_0),.clk(gclk));
	jdff dff_B_UWtMXrMa8_0(.din(w_dff_B_lqayjOb33_0),.dout(w_dff_B_UWtMXrMa8_0),.clk(gclk));
	jdff dff_B_EgurrhzS3_1(.din(G116),.dout(w_dff_B_EgurrhzS3_1),.clk(gclk));
	jdff dff_B_qH7SRKVN3_1(.din(w_dff_B_EgurrhzS3_1),.dout(w_dff_B_qH7SRKVN3_1),.clk(gclk));
	jdff dff_A_DNotvZS61_1(.dout(w_n971_0[1]),.din(w_dff_A_DNotvZS61_1),.clk(gclk));
	jdff dff_B_0uH6sVWG8_1(.din(n967),.dout(w_dff_B_0uH6sVWG8_1),.clk(gclk));
	jdff dff_B_UuRwrD601_1(.din(w_dff_B_0uH6sVWG8_1),.dout(w_dff_B_UuRwrD601_1),.clk(gclk));
	jdff dff_B_zznk1NDg9_1(.din(w_dff_B_UuRwrD601_1),.dout(w_dff_B_zznk1NDg9_1),.clk(gclk));
	jdff dff_B_6PAokJul5_1(.din(w_dff_B_zznk1NDg9_1),.dout(w_dff_B_6PAokJul5_1),.clk(gclk));
	jdff dff_B_carxNRFb2_1(.din(w_dff_B_6PAokJul5_1),.dout(w_dff_B_carxNRFb2_1),.clk(gclk));
	jdff dff_B_Znrzi2Jp6_1(.din(w_dff_B_carxNRFb2_1),.dout(w_dff_B_Znrzi2Jp6_1),.clk(gclk));
	jdff dff_B_TQCUVPUU7_1(.din(w_dff_B_Znrzi2Jp6_1),.dout(w_dff_B_TQCUVPUU7_1),.clk(gclk));
	jdff dff_B_sAY3s7jv2_1(.din(w_dff_B_TQCUVPUU7_1),.dout(w_dff_B_sAY3s7jv2_1),.clk(gclk));
	jdff dff_B_OOTinskz4_1(.din(w_dff_B_sAY3s7jv2_1),.dout(w_dff_B_OOTinskz4_1),.clk(gclk));
	jdff dff_B_DrJsBLWi0_1(.din(w_dff_B_OOTinskz4_1),.dout(w_dff_B_DrJsBLWi0_1),.clk(gclk));
	jdff dff_B_knbxOmLs0_0(.din(n1211),.dout(w_dff_B_knbxOmLs0_0),.clk(gclk));
	jdff dff_B_VFdQSXig9_0(.din(w_dff_B_knbxOmLs0_0),.dout(w_dff_B_VFdQSXig9_0),.clk(gclk));
	jdff dff_B_u7GkHHnL4_0(.din(w_dff_B_VFdQSXig9_0),.dout(w_dff_B_u7GkHHnL4_0),.clk(gclk));
	jdff dff_B_cjLvs0lE2_0(.din(w_dff_B_u7GkHHnL4_0),.dout(w_dff_B_cjLvs0lE2_0),.clk(gclk));
	jdff dff_B_wh4YQLXe2_0(.din(w_dff_B_cjLvs0lE2_0),.dout(w_dff_B_wh4YQLXe2_0),.clk(gclk));
	jdff dff_B_XIHeVgmt9_0(.din(w_dff_B_wh4YQLXe2_0),.dout(w_dff_B_XIHeVgmt9_0),.clk(gclk));
	jdff dff_B_gGeo0y4J5_0(.din(w_dff_B_XIHeVgmt9_0),.dout(w_dff_B_gGeo0y4J5_0),.clk(gclk));
	jdff dff_B_QCmH1uUZ1_0(.din(w_dff_B_gGeo0y4J5_0),.dout(w_dff_B_QCmH1uUZ1_0),.clk(gclk));
	jdff dff_B_UbmoN6sJ0_0(.din(w_dff_B_QCmH1uUZ1_0),.dout(w_dff_B_UbmoN6sJ0_0),.clk(gclk));
	jdff dff_B_YMzSjBaa5_0(.din(w_dff_B_UbmoN6sJ0_0),.dout(w_dff_B_YMzSjBaa5_0),.clk(gclk));
	jdff dff_B_N1JcnImR0_0(.din(w_dff_B_YMzSjBaa5_0),.dout(w_dff_B_N1JcnImR0_0),.clk(gclk));
	jdff dff_B_4sIPjaQH0_0(.din(n1210),.dout(w_dff_B_4sIPjaQH0_0),.clk(gclk));
	jdff dff_B_cTovec442_0(.din(w_dff_B_4sIPjaQH0_0),.dout(w_dff_B_cTovec442_0),.clk(gclk));
	jdff dff_B_h4nnryEP7_1(.din(G53),.dout(w_dff_B_h4nnryEP7_1),.clk(gclk));
	jdff dff_B_pPteiRlH7_1(.din(w_dff_B_h4nnryEP7_1),.dout(w_dff_B_pPteiRlH7_1),.clk(gclk));
	jdff dff_B_5azsRgP08_0(.din(n516),.dout(w_dff_B_5azsRgP08_0),.clk(gclk));
	jdff dff_B_8ngaOgZp0_1(.din(n508),.dout(w_dff_B_8ngaOgZp0_1),.clk(gclk));
	jdff dff_B_ghmy57IS4_1(.din(n949),.dout(w_dff_B_ghmy57IS4_1),.clk(gclk));
	jdff dff_B_ulSZtaFu8_1(.din(w_dff_B_ghmy57IS4_1),.dout(w_dff_B_ulSZtaFu8_1),.clk(gclk));
	jdff dff_B_6IZ25oof1_1(.din(w_dff_B_ulSZtaFu8_1),.dout(w_dff_B_6IZ25oof1_1),.clk(gclk));
	jdff dff_B_rqgEC4XS4_1(.din(w_dff_B_6IZ25oof1_1),.dout(w_dff_B_rqgEC4XS4_1),.clk(gclk));
	jdff dff_B_qrbp3l5i8_1(.din(w_dff_B_rqgEC4XS4_1),.dout(w_dff_B_qrbp3l5i8_1),.clk(gclk));
	jdff dff_B_Z5TGiR6n4_1(.din(w_dff_B_qrbp3l5i8_1),.dout(w_dff_B_Z5TGiR6n4_1),.clk(gclk));
	jdff dff_B_X8We1c0a4_1(.din(w_dff_B_Z5TGiR6n4_1),.dout(w_dff_B_X8We1c0a4_1),.clk(gclk));
	jdff dff_B_x7A8Np4n0_1(.din(w_dff_B_X8We1c0a4_1),.dout(w_dff_B_x7A8Np4n0_1),.clk(gclk));
	jdff dff_B_UDifye6W0_1(.din(w_dff_B_x7A8Np4n0_1),.dout(w_dff_B_UDifye6W0_1),.clk(gclk));
	jdff dff_B_VGJ83NmS9_1(.din(w_dff_B_UDifye6W0_1),.dout(w_dff_B_VGJ83NmS9_1),.clk(gclk));
	jdff dff_B_nsf7sUfc3_1(.din(n950),.dout(w_dff_B_nsf7sUfc3_1),.clk(gclk));
	jdff dff_B_Ui9iQyjd0_1(.din(w_dff_B_nsf7sUfc3_1),.dout(w_dff_B_Ui9iQyjd0_1),.clk(gclk));
	jdff dff_B_2jmTBkcx4_1(.din(w_dff_B_Ui9iQyjd0_1),.dout(w_dff_B_2jmTBkcx4_1),.clk(gclk));
	jdff dff_B_Q7f9PXUA6_1(.din(w_dff_B_2jmTBkcx4_1),.dout(w_dff_B_Q7f9PXUA6_1),.clk(gclk));
	jdff dff_B_ZQO9pmoP6_1(.din(w_dff_B_Q7f9PXUA6_1),.dout(w_dff_B_ZQO9pmoP6_1),.clk(gclk));
	jdff dff_B_5Ot26uPJ7_1(.din(w_dff_B_ZQO9pmoP6_1),.dout(w_dff_B_5Ot26uPJ7_1),.clk(gclk));
	jdff dff_B_6ZwNLYnp6_1(.din(w_dff_B_5Ot26uPJ7_1),.dout(w_dff_B_6ZwNLYnp6_1),.clk(gclk));
	jdff dff_B_7J51VwjJ9_1(.din(w_dff_B_6ZwNLYnp6_1),.dout(w_dff_B_7J51VwjJ9_1),.clk(gclk));
	jdff dff_B_JasYwprn6_1(.din(w_dff_B_7J51VwjJ9_1),.dout(w_dff_B_JasYwprn6_1),.clk(gclk));
	jdff dff_A_eTIhmptp4_1(.dout(w_n748_1[1]),.din(w_dff_A_eTIhmptp4_1),.clk(gclk));
	jdff dff_A_0ABgA4ZH5_1(.dout(w_dff_A_eTIhmptp4_1),.din(w_dff_A_0ABgA4ZH5_1),.clk(gclk));
	jdff dff_A_nWwNMmAl9_1(.dout(w_dff_A_0ABgA4ZH5_1),.din(w_dff_A_nWwNMmAl9_1),.clk(gclk));
	jdff dff_A_e5sfyIm04_1(.dout(w_dff_A_nWwNMmAl9_1),.din(w_dff_A_e5sfyIm04_1),.clk(gclk));
	jdff dff_A_WmOrV3Fc7_1(.dout(w_dff_A_e5sfyIm04_1),.din(w_dff_A_WmOrV3Fc7_1),.clk(gclk));
	jdff dff_A_TxbQkaMK3_1(.dout(w_dff_A_WmOrV3Fc7_1),.din(w_dff_A_TxbQkaMK3_1),.clk(gclk));
	jdff dff_A_pUdYOU2L4_1(.dout(w_dff_A_TxbQkaMK3_1),.din(w_dff_A_pUdYOU2L4_1),.clk(gclk));
	jdff dff_A_fT9ePtr77_1(.dout(w_dff_A_pUdYOU2L4_1),.din(w_dff_A_fT9ePtr77_1),.clk(gclk));
	jdff dff_A_uLpVJ25x2_1(.dout(w_dff_A_fT9ePtr77_1),.din(w_dff_A_uLpVJ25x2_1),.clk(gclk));
	jdff dff_A_fGyFZUvc5_1(.dout(w_dff_A_uLpVJ25x2_1),.din(w_dff_A_fGyFZUvc5_1),.clk(gclk));
	jdff dff_A_59LsnX7Q3_1(.dout(w_dff_A_fGyFZUvc5_1),.din(w_dff_A_59LsnX7Q3_1),.clk(gclk));
	jdff dff_A_018LXOWc5_1(.dout(w_dff_A_59LsnX7Q3_1),.din(w_dff_A_018LXOWc5_1),.clk(gclk));
	jdff dff_A_pVTYFNtE9_1(.dout(w_dff_A_018LXOWc5_1),.din(w_dff_A_pVTYFNtE9_1),.clk(gclk));
	jdff dff_A_eTYBwnWT9_2(.dout(w_n748_1[2]),.din(w_dff_A_eTYBwnWT9_2),.clk(gclk));
	jdff dff_A_Nsw36ZaJ8_2(.dout(w_dff_A_eTYBwnWT9_2),.din(w_dff_A_Nsw36ZaJ8_2),.clk(gclk));
	jdff dff_A_srXh94j66_2(.dout(w_dff_A_Nsw36ZaJ8_2),.din(w_dff_A_srXh94j66_2),.clk(gclk));
	jdff dff_A_iOykxtBa3_2(.dout(w_dff_A_srXh94j66_2),.din(w_dff_A_iOykxtBa3_2),.clk(gclk));
	jdff dff_A_r0gtHvQl2_2(.dout(w_dff_A_iOykxtBa3_2),.din(w_dff_A_r0gtHvQl2_2),.clk(gclk));
	jdff dff_A_5Oo6AbkR6_2(.dout(w_dff_A_r0gtHvQl2_2),.din(w_dff_A_5Oo6AbkR6_2),.clk(gclk));
	jdff dff_A_1HpV4mEj0_2(.dout(w_dff_A_5Oo6AbkR6_2),.din(w_dff_A_1HpV4mEj0_2),.clk(gclk));
	jdff dff_A_mJ6drfkE6_2(.dout(w_dff_A_1HpV4mEj0_2),.din(w_dff_A_mJ6drfkE6_2),.clk(gclk));
	jdff dff_A_dkLkqm3k4_2(.dout(w_dff_A_mJ6drfkE6_2),.din(w_dff_A_dkLkqm3k4_2),.clk(gclk));
	jdff dff_A_xnxpTREI0_2(.dout(w_dff_A_dkLkqm3k4_2),.din(w_dff_A_xnxpTREI0_2),.clk(gclk));
	jdff dff_A_1Go8PI2h1_2(.dout(w_dff_A_xnxpTREI0_2),.din(w_dff_A_1Go8PI2h1_2),.clk(gclk));
	jdff dff_A_38LaT17l8_2(.dout(w_dff_A_1Go8PI2h1_2),.din(w_dff_A_38LaT17l8_2),.clk(gclk));
	jdff dff_B_AZprxqzJ0_0(.din(n1333),.dout(w_dff_B_AZprxqzJ0_0),.clk(gclk));
	jdff dff_B_mJ1j1gTD0_0(.din(w_dff_B_AZprxqzJ0_0),.dout(w_dff_B_mJ1j1gTD0_0),.clk(gclk));
	jdff dff_B_7HZIShAY0_0(.din(w_dff_B_mJ1j1gTD0_0),.dout(w_dff_B_7HZIShAY0_0),.clk(gclk));
	jdff dff_B_n1wrDYVY5_0(.din(w_dff_B_7HZIShAY0_0),.dout(w_dff_B_n1wrDYVY5_0),.clk(gclk));
	jdff dff_B_1RR1CZsP4_0(.din(w_dff_B_n1wrDYVY5_0),.dout(w_dff_B_1RR1CZsP4_0),.clk(gclk));
	jdff dff_B_tfpD0Udf2_0(.din(w_dff_B_1RR1CZsP4_0),.dout(w_dff_B_tfpD0Udf2_0),.clk(gclk));
	jdff dff_B_vSj85tUk1_0(.din(w_dff_B_tfpD0Udf2_0),.dout(w_dff_B_vSj85tUk1_0),.clk(gclk));
	jdff dff_B_pVt6E6em8_0(.din(w_dff_B_vSj85tUk1_0),.dout(w_dff_B_pVt6E6em8_0),.clk(gclk));
	jdff dff_B_7zjMzTiS5_0(.din(w_dff_B_pVt6E6em8_0),.dout(w_dff_B_7zjMzTiS5_0),.clk(gclk));
	jdff dff_B_oScitRmT1_0(.din(w_dff_B_7zjMzTiS5_0),.dout(w_dff_B_oScitRmT1_0),.clk(gclk));
	jdff dff_B_yFm1JmTH9_0(.din(w_dff_B_oScitRmT1_0),.dout(w_dff_B_yFm1JmTH9_0),.clk(gclk));
	jdff dff_B_2dJWhgjF7_0(.din(w_dff_B_yFm1JmTH9_0),.dout(w_dff_B_2dJWhgjF7_0),.clk(gclk));
	jdff dff_B_qLHmevy57_0(.din(w_dff_B_2dJWhgjF7_0),.dout(w_dff_B_qLHmevy57_0),.clk(gclk));
	jdff dff_B_TuGE8FT87_0(.din(w_dff_B_qLHmevy57_0),.dout(w_dff_B_TuGE8FT87_0),.clk(gclk));
	jdff dff_B_tKJwDoLf8_0(.din(w_dff_B_TuGE8FT87_0),.dout(w_dff_B_tKJwDoLf8_0),.clk(gclk));
	jdff dff_B_r8jmrCwB8_0(.din(w_dff_B_tKJwDoLf8_0),.dout(w_dff_B_r8jmrCwB8_0),.clk(gclk));
	jdff dff_B_b4LZq0Iw7_0(.din(n1332),.dout(w_dff_B_b4LZq0Iw7_0),.clk(gclk));
	jdff dff_B_8Rzw76ML0_2(.din(G164),.dout(w_dff_B_8Rzw76ML0_2),.clk(gclk));
	jdff dff_B_UxgFEG5G5_2(.din(G194),.dout(w_dff_B_UxgFEG5G5_2),.clk(gclk));
	jdff dff_B_kg6O6kvQ3_2(.din(w_dff_B_UxgFEG5G5_2),.dout(w_dff_B_kg6O6kvQ3_2),.clk(gclk));
	jdff dff_B_BzXtCudD3_0(.din(n1169),.dout(w_dff_B_BzXtCudD3_0),.clk(gclk));
	jdff dff_B_64ZAyU2B5_0(.din(w_dff_B_BzXtCudD3_0),.dout(w_dff_B_64ZAyU2B5_0),.clk(gclk));
	jdff dff_B_1yU9SCky0_0(.din(w_dff_B_64ZAyU2B5_0),.dout(w_dff_B_1yU9SCky0_0),.clk(gclk));
	jdff dff_B_eeKeqSw40_0(.din(w_dff_B_1yU9SCky0_0),.dout(w_dff_B_eeKeqSw40_0),.clk(gclk));
	jdff dff_B_g1Qpje6Z1_0(.din(w_dff_B_eeKeqSw40_0),.dout(w_dff_B_g1Qpje6Z1_0),.clk(gclk));
	jdff dff_B_tzWsAc6R7_0(.din(w_dff_B_g1Qpje6Z1_0),.dout(w_dff_B_tzWsAc6R7_0),.clk(gclk));
	jdff dff_B_ytQDl9nC8_0(.din(w_dff_B_tzWsAc6R7_0),.dout(w_dff_B_ytQDl9nC8_0),.clk(gclk));
	jdff dff_B_Myw9mLdh9_0(.din(w_dff_B_ytQDl9nC8_0),.dout(w_dff_B_Myw9mLdh9_0),.clk(gclk));
	jdff dff_B_8XhrK0Hx5_0(.din(w_dff_B_Myw9mLdh9_0),.dout(w_dff_B_8XhrK0Hx5_0),.clk(gclk));
	jdff dff_B_cJFTjYXl4_0(.din(w_dff_B_8XhrK0Hx5_0),.dout(w_dff_B_cJFTjYXl4_0),.clk(gclk));
	jdff dff_B_5EJPR0oB7_0(.din(w_dff_B_cJFTjYXl4_0),.dout(w_dff_B_5EJPR0oB7_0),.clk(gclk));
	jdff dff_B_e3bAn2re2_0(.din(n1167),.dout(w_dff_B_e3bAn2re2_0),.clk(gclk));
	jdff dff_B_CUFbrsfo3_1(.din(G121),.dout(w_dff_B_CUFbrsfo3_1),.clk(gclk));
	jdff dff_B_qIHigijf7_1(.din(w_dff_B_CUFbrsfo3_1),.dout(w_dff_B_qIHigijf7_1),.clk(gclk));
	jdff dff_A_zHdw3oJE0_0(.dout(w_n748_2[0]),.din(w_dff_A_zHdw3oJE0_0),.clk(gclk));
	jdff dff_A_AFXfzUH98_0(.dout(w_dff_A_zHdw3oJE0_0),.din(w_dff_A_AFXfzUH98_0),.clk(gclk));
	jdff dff_A_Uhkbv8Pc0_0(.dout(w_dff_A_AFXfzUH98_0),.din(w_dff_A_Uhkbv8Pc0_0),.clk(gclk));
	jdff dff_A_xIckdFqs7_0(.dout(w_dff_A_Uhkbv8Pc0_0),.din(w_dff_A_xIckdFqs7_0),.clk(gclk));
	jdff dff_A_oaUSor5k9_2(.dout(w_n748_2[2]),.din(w_dff_A_oaUSor5k9_2),.clk(gclk));
	jdff dff_A_6f8Kk6ui9_2(.dout(w_dff_A_oaUSor5k9_2),.din(w_dff_A_6f8Kk6ui9_2),.clk(gclk));
	jdff dff_A_hm8qYiz91_1(.dout(w_n748_0[1]),.din(w_dff_A_hm8qYiz91_1),.clk(gclk));
	jdff dff_A_w7FT3ZHn7_1(.dout(w_dff_A_hm8qYiz91_1),.din(w_dff_A_w7FT3ZHn7_1),.clk(gclk));
	jdff dff_A_vZuh13DQ2_1(.dout(w_dff_A_w7FT3ZHn7_1),.din(w_dff_A_vZuh13DQ2_1),.clk(gclk));
	jdff dff_A_GSd6Hx7u4_1(.dout(w_dff_A_vZuh13DQ2_1),.din(w_dff_A_GSd6Hx7u4_1),.clk(gclk));
	jdff dff_A_tA1UrYIt4_1(.dout(w_dff_A_GSd6Hx7u4_1),.din(w_dff_A_tA1UrYIt4_1),.clk(gclk));
	jdff dff_A_bHU8Cxld7_1(.dout(w_dff_A_tA1UrYIt4_1),.din(w_dff_A_bHU8Cxld7_1),.clk(gclk));
	jdff dff_A_MDJfGGFF6_1(.dout(w_dff_A_bHU8Cxld7_1),.din(w_dff_A_MDJfGGFF6_1),.clk(gclk));
	jdff dff_A_UfZ86a0w8_1(.dout(w_dff_A_MDJfGGFF6_1),.din(w_dff_A_UfZ86a0w8_1),.clk(gclk));
	jdff dff_A_iUdpGVFf1_2(.dout(w_n748_0[2]),.din(w_dff_A_iUdpGVFf1_2),.clk(gclk));
	jdff dff_A_SRHHe0ma6_2(.dout(w_dff_A_iUdpGVFf1_2),.din(w_dff_A_SRHHe0ma6_2),.clk(gclk));
	jdff dff_A_DGzWvVuZ2_2(.dout(w_dff_A_SRHHe0ma6_2),.din(w_dff_A_DGzWvVuZ2_2),.clk(gclk));
	jdff dff_A_N4ptuOW26_2(.dout(w_dff_A_DGzWvVuZ2_2),.din(w_dff_A_N4ptuOW26_2),.clk(gclk));
	jdff dff_B_ihQVpXUD7_3(.din(n748),.dout(w_dff_B_ihQVpXUD7_3),.clk(gclk));
	jdff dff_A_RVWRKP4u1_0(.dout(w_n747_3[0]),.din(w_dff_A_RVWRKP4u1_0),.clk(gclk));
	jdff dff_A_UsOp91Lb7_0(.dout(w_dff_A_RVWRKP4u1_0),.din(w_dff_A_UsOp91Lb7_0),.clk(gclk));
	jdff dff_A_J08NF0FU0_0(.dout(w_dff_A_UsOp91Lb7_0),.din(w_dff_A_J08NF0FU0_0),.clk(gclk));
	jdff dff_A_2BCbV1iz5_0(.dout(w_dff_A_J08NF0FU0_0),.din(w_dff_A_2BCbV1iz5_0),.clk(gclk));
	jdff dff_A_Iy73Tv2g0_0(.dout(w_dff_A_2BCbV1iz5_0),.din(w_dff_A_Iy73Tv2g0_0),.clk(gclk));
	jdff dff_A_MOpsaM2X7_0(.dout(w_dff_A_Iy73Tv2g0_0),.din(w_dff_A_MOpsaM2X7_0),.clk(gclk));
	jdff dff_A_v7q9nTJl1_0(.dout(w_dff_A_MOpsaM2X7_0),.din(w_dff_A_v7q9nTJl1_0),.clk(gclk));
	jdff dff_A_COGThtqU9_0(.dout(w_dff_A_v7q9nTJl1_0),.din(w_dff_A_COGThtqU9_0),.clk(gclk));
	jdff dff_A_pFbXiNEm7_1(.dout(w_n747_3[1]),.din(w_dff_A_pFbXiNEm7_1),.clk(gclk));
	jdff dff_A_eKidrWQg0_1(.dout(w_dff_A_pFbXiNEm7_1),.din(w_dff_A_eKidrWQg0_1),.clk(gclk));
	jdff dff_A_mE9sZeDh0_1(.dout(w_dff_A_eKidrWQg0_1),.din(w_dff_A_mE9sZeDh0_1),.clk(gclk));
	jdff dff_A_rcHSEw7v8_0(.dout(w_n1002_2[0]),.din(w_dff_A_rcHSEw7v8_0),.clk(gclk));
	jdff dff_A_BDAlbrwS2_1(.dout(w_n1002_2[1]),.din(w_dff_A_BDAlbrwS2_1),.clk(gclk));
	jdff dff_B_CQd7OXAe5_0(.din(n1204),.dout(w_dff_B_CQd7OXAe5_0),.clk(gclk));
	jdff dff_B_5QXWSjRb3_0(.din(w_dff_B_CQd7OXAe5_0),.dout(w_dff_B_5QXWSjRb3_0),.clk(gclk));
	jdff dff_B_R7dNp7hJ7_0(.din(w_dff_B_5QXWSjRb3_0),.dout(w_dff_B_R7dNp7hJ7_0),.clk(gclk));
	jdff dff_B_n3xBIV976_0(.din(w_dff_B_R7dNp7hJ7_0),.dout(w_dff_B_n3xBIV976_0),.clk(gclk));
	jdff dff_B_LIfP6j794_0(.din(w_dff_B_n3xBIV976_0),.dout(w_dff_B_LIfP6j794_0),.clk(gclk));
	jdff dff_B_BpP2UyFK0_0(.din(w_dff_B_LIfP6j794_0),.dout(w_dff_B_BpP2UyFK0_0),.clk(gclk));
	jdff dff_B_nKDMICHL9_0(.din(w_dff_B_BpP2UyFK0_0),.dout(w_dff_B_nKDMICHL9_0),.clk(gclk));
	jdff dff_B_dT3YUtLv0_0(.din(w_dff_B_nKDMICHL9_0),.dout(w_dff_B_dT3YUtLv0_0),.clk(gclk));
	jdff dff_B_xDE9Jiw79_0(.din(w_dff_B_dT3YUtLv0_0),.dout(w_dff_B_xDE9Jiw79_0),.clk(gclk));
	jdff dff_B_9aBtAWWI9_0(.din(w_dff_B_xDE9Jiw79_0),.dout(w_dff_B_9aBtAWWI9_0),.clk(gclk));
	jdff dff_B_pRA1cafs6_0(.din(w_dff_B_9aBtAWWI9_0),.dout(w_dff_B_pRA1cafs6_0),.clk(gclk));
	jdff dff_B_ZvN6PyDk5_0(.din(n1202),.dout(w_dff_B_ZvN6PyDk5_0),.clk(gclk));
	jdff dff_B_8vNbqRXJ6_0(.din(w_dff_B_ZvN6PyDk5_0),.dout(w_dff_B_8vNbqRXJ6_0),.clk(gclk));
	jdff dff_B_eHQunb1k9_1(.din(G114),.dout(w_dff_B_eHQunb1k9_1),.clk(gclk));
	jdff dff_B_evsv9m3f0_1(.din(w_dff_B_eHQunb1k9_1),.dout(w_dff_B_evsv9m3f0_1),.clk(gclk));
	jdff dff_B_AlfhYG632_3(.din(n765),.dout(w_dff_B_AlfhYG632_3),.clk(gclk));
	jdff dff_B_zVEI9lAu4_3(.din(w_dff_B_AlfhYG632_3),.dout(w_dff_B_zVEI9lAu4_3),.clk(gclk));
	jdff dff_A_wIJmSegh5_1(.dout(w_n751_2[1]),.din(w_dff_A_wIJmSegh5_1),.clk(gclk));
	jdff dff_B_Lm8hocjk6_0(.din(n550),.dout(w_dff_B_Lm8hocjk6_0),.clk(gclk));
	jdff dff_B_r7DXClUe9_3(.din(G3548),.dout(w_dff_B_r7DXClUe9_3),.clk(gclk));
	jdff dff_B_3iQ4hjCX7_1(.din(n542),.dout(w_dff_B_3iQ4hjCX7_1),.clk(gclk));
	jdff dff_A_CohO1dF46_0(.dout(w_n999_2[0]),.din(w_dff_A_CohO1dF46_0),.clk(gclk));
	jdff dff_A_pvudMBQF0_1(.dout(w_n999_2[1]),.din(w_dff_A_pvudMBQF0_1),.clk(gclk));
	jdff dff_A_eo9C9SN44_0(.dout(w_G137_4[0]),.din(w_dff_A_eo9C9SN44_0),.clk(gclk));
	jdff dff_A_nd61yT9j0_1(.dout(w_G137_4[1]),.din(w_dff_A_nd61yT9j0_1),.clk(gclk));
	jdff dff_A_el7JVLJ86_0(.dout(w_G137_1[0]),.din(w_dff_A_el7JVLJ86_0),.clk(gclk));
	jdff dff_A_OSLWcwJ35_0(.dout(w_dff_A_el7JVLJ86_0),.din(w_dff_A_OSLWcwJ35_0),.clk(gclk));
	jdff dff_A_Cs21iRWK2_0(.dout(w_dff_A_OSLWcwJ35_0),.din(w_dff_A_Cs21iRWK2_0),.clk(gclk));
	jdff dff_A_GF7DKR0k2_0(.dout(w_dff_A_Cs21iRWK2_0),.din(w_dff_A_GF7DKR0k2_0),.clk(gclk));
	jdff dff_A_bi3X8rNv0_0(.dout(w_dff_A_GF7DKR0k2_0),.din(w_dff_A_bi3X8rNv0_0),.clk(gclk));
	jdff dff_A_46Zjjtm19_1(.dout(w_G137_1[1]),.din(w_dff_A_46Zjjtm19_1),.clk(gclk));
	jdff dff_A_2wQNXJ733_1(.dout(w_dff_A_46Zjjtm19_1),.din(w_dff_A_2wQNXJ733_1),.clk(gclk));
	jdff dff_A_ll5qnhqY0_1(.dout(w_dff_A_2wQNXJ733_1),.din(w_dff_A_ll5qnhqY0_1),.clk(gclk));
	jdff dff_A_thSmdNK93_1(.dout(w_dff_A_ll5qnhqY0_1),.din(w_dff_A_thSmdNK93_1),.clk(gclk));
	jdff dff_A_cblSsHYI7_1(.dout(w_dff_A_thSmdNK93_1),.din(w_dff_A_cblSsHYI7_1),.clk(gclk));
	jdff dff_A_ooNgcASa8_1(.dout(w_dff_A_cblSsHYI7_1),.din(w_dff_A_ooNgcASa8_1),.clk(gclk));
	jdff dff_B_almq03eI8_0(.din(n1341),.dout(w_dff_B_almq03eI8_0),.clk(gclk));
	jdff dff_B_IRLgO7kt4_0(.din(w_dff_B_almq03eI8_0),.dout(w_dff_B_IRLgO7kt4_0),.clk(gclk));
	jdff dff_B_Blybwakb8_0(.din(w_dff_B_IRLgO7kt4_0),.dout(w_dff_B_Blybwakb8_0),.clk(gclk));
	jdff dff_B_0RFEi9ci0_0(.din(w_dff_B_Blybwakb8_0),.dout(w_dff_B_0RFEi9ci0_0),.clk(gclk));
	jdff dff_B_MeIY2g1J9_0(.din(w_dff_B_0RFEi9ci0_0),.dout(w_dff_B_MeIY2g1J9_0),.clk(gclk));
	jdff dff_B_wirLnp5Y7_0(.din(w_dff_B_MeIY2g1J9_0),.dout(w_dff_B_wirLnp5Y7_0),.clk(gclk));
	jdff dff_B_sZFEaVQg0_0(.din(w_dff_B_wirLnp5Y7_0),.dout(w_dff_B_sZFEaVQg0_0),.clk(gclk));
	jdff dff_B_NMbhQSno3_0(.din(w_dff_B_sZFEaVQg0_0),.dout(w_dff_B_NMbhQSno3_0),.clk(gclk));
	jdff dff_B_f1WBGkjH6_0(.din(w_dff_B_NMbhQSno3_0),.dout(w_dff_B_f1WBGkjH6_0),.clk(gclk));
	jdff dff_B_r142rHGR1_0(.din(w_dff_B_f1WBGkjH6_0),.dout(w_dff_B_r142rHGR1_0),.clk(gclk));
	jdff dff_B_QXlYfsDA3_0(.din(w_dff_B_r142rHGR1_0),.dout(w_dff_B_QXlYfsDA3_0),.clk(gclk));
	jdff dff_B_qINY983G6_0(.din(w_dff_B_QXlYfsDA3_0),.dout(w_dff_B_qINY983G6_0),.clk(gclk));
	jdff dff_B_ITqUOcel1_0(.din(w_dff_B_qINY983G6_0),.dout(w_dff_B_ITqUOcel1_0),.clk(gclk));
	jdff dff_B_wjxWFONT5_0(.din(w_dff_B_ITqUOcel1_0),.dout(w_dff_B_wjxWFONT5_0),.clk(gclk));
	jdff dff_B_t7Yetd7S2_0(.din(w_dff_B_wjxWFONT5_0),.dout(w_dff_B_t7Yetd7S2_0),.clk(gclk));
	jdff dff_B_Rly3K5lm9_0(.din(w_dff_B_t7Yetd7S2_0),.dout(w_dff_B_Rly3K5lm9_0),.clk(gclk));
	jdff dff_B_Cz04OjIr1_0(.din(w_dff_B_Rly3K5lm9_0),.dout(w_dff_B_Cz04OjIr1_0),.clk(gclk));
	jdff dff_B_vnyIMFO61_0(.din(n1340),.dout(w_dff_B_vnyIMFO61_0),.clk(gclk));
	jdff dff_B_FiyemRXA2_2(.din(G161),.dout(w_dff_B_FiyemRXA2_2),.clk(gclk));
	jdff dff_B_px3atMtj6_2(.din(G191),.dout(w_dff_B_px3atMtj6_2),.clk(gclk));
	jdff dff_B_PNYWUf4z8_2(.din(w_dff_B_px3atMtj6_2),.dout(w_dff_B_PNYWUf4z8_2),.clk(gclk));
	jdff dff_B_IT0FyqTn8_0(.din(n1162),.dout(w_dff_B_IT0FyqTn8_0),.clk(gclk));
	jdff dff_B_aYFo1R831_0(.din(w_dff_B_IT0FyqTn8_0),.dout(w_dff_B_aYFo1R831_0),.clk(gclk));
	jdff dff_B_9oEZ1EmU6_0(.din(w_dff_B_aYFo1R831_0),.dout(w_dff_B_9oEZ1EmU6_0),.clk(gclk));
	jdff dff_B_oGgbRWhq1_0(.din(w_dff_B_9oEZ1EmU6_0),.dout(w_dff_B_oGgbRWhq1_0),.clk(gclk));
	jdff dff_B_5vOD4vSr4_0(.din(w_dff_B_oGgbRWhq1_0),.dout(w_dff_B_5vOD4vSr4_0),.clk(gclk));
	jdff dff_B_RuDVHECz3_0(.din(w_dff_B_5vOD4vSr4_0),.dout(w_dff_B_RuDVHECz3_0),.clk(gclk));
	jdff dff_B_J1fDPc8v1_0(.din(w_dff_B_RuDVHECz3_0),.dout(w_dff_B_J1fDPc8v1_0),.clk(gclk));
	jdff dff_B_DnvMvUNs7_0(.din(w_dff_B_J1fDPc8v1_0),.dout(w_dff_B_DnvMvUNs7_0),.clk(gclk));
	jdff dff_B_8QCisCFT2_0(.din(w_dff_B_DnvMvUNs7_0),.dout(w_dff_B_8QCisCFT2_0),.clk(gclk));
	jdff dff_B_ntq2q3TZ1_0(.din(w_dff_B_8QCisCFT2_0),.dout(w_dff_B_ntq2q3TZ1_0),.clk(gclk));
	jdff dff_B_YsrSnTeg1_0(.din(w_dff_B_ntq2q3TZ1_0),.dout(w_dff_B_YsrSnTeg1_0),.clk(gclk));
	jdff dff_B_QLeuCNyl6_0(.din(w_dff_B_YsrSnTeg1_0),.dout(w_dff_B_QLeuCNyl6_0),.clk(gclk));
	jdff dff_B_dJTTVpsB3_0(.din(w_dff_B_QLeuCNyl6_0),.dout(w_dff_B_dJTTVpsB3_0),.clk(gclk));
	jdff dff_B_cF4ZbbJB2_1(.din(n1160),.dout(w_dff_B_cF4ZbbJB2_1),.clk(gclk));
	jdff dff_B_WSVXGEBq2_1(.din(w_dff_B_cF4ZbbJB2_1),.dout(w_dff_B_WSVXGEBq2_1),.clk(gclk));
	jdff dff_A_3ZPaxM2o1_1(.dout(w_n751_1[1]),.din(w_dff_A_3ZPaxM2o1_1),.clk(gclk));
	jdff dff_A_knKS0aNM9_0(.dout(w_G123_0[0]),.din(w_dff_A_knKS0aNM9_0),.clk(gclk));
	jdff dff_B_YztjzzMN1_2(.din(G123),.dout(w_dff_B_YztjzzMN1_2),.clk(gclk));
	jdff dff_B_gcIRcr813_0(.din(n788),.dout(w_dff_B_gcIRcr813_0),.clk(gclk));
	jdff dff_B_GVlAryBp3_0(.din(n780),.dout(w_dff_B_GVlAryBp3_0),.clk(gclk));
	jdff dff_B_GUlMS4gv6_0(.din(w_dff_B_GVlAryBp3_0),.dout(w_dff_B_GUlMS4gv6_0),.clk(gclk));
	jdff dff_B_3RXYZWmb0_0(.din(w_dff_B_GUlMS4gv6_0),.dout(w_dff_B_3RXYZWmb0_0),.clk(gclk));
	jdff dff_A_ux3c2iUQ5_0(.dout(w_G54_0[0]),.din(w_dff_A_ux3c2iUQ5_0),.clk(gclk));
	jdff dff_A_xHdeIjsH5_0(.dout(w_dff_A_ux3c2iUQ5_0),.din(w_dff_A_xHdeIjsH5_0),.clk(gclk));
	jdff dff_A_Ptqp5SJG7_0(.dout(w_dff_A_xHdeIjsH5_0),.din(w_dff_A_Ptqp5SJG7_0),.clk(gclk));
	jdff dff_A_NWYkjshc5_0(.dout(w_dff_A_Ptqp5SJG7_0),.din(w_dff_A_NWYkjshc5_0),.clk(gclk));
	jdff dff_A_SjLtKWoS8_0(.dout(w_dff_A_NWYkjshc5_0),.din(w_dff_A_SjLtKWoS8_0),.clk(gclk));
	jdff dff_A_7xOfXmXs0_0(.dout(w_dff_A_SjLtKWoS8_0),.din(w_dff_A_7xOfXmXs0_0),.clk(gclk));
	jdff dff_A_25C853gH3_0(.dout(w_dff_A_7xOfXmXs0_0),.din(w_dff_A_25C853gH3_0),.clk(gclk));
	jdff dff_A_arY8dTIP6_0(.dout(w_dff_A_25C853gH3_0),.din(w_dff_A_arY8dTIP6_0),.clk(gclk));
	jdff dff_A_dMhfcUjY7_0(.dout(w_n741_0[0]),.din(w_dff_A_dMhfcUjY7_0),.clk(gclk));
	jdff dff_A_PvX7XXFv4_0(.dout(w_dff_A_dMhfcUjY7_0),.din(w_dff_A_PvX7XXFv4_0),.clk(gclk));
	jdff dff_A_DiOMKzrL1_0(.dout(w_dff_A_PvX7XXFv4_0),.din(w_dff_A_DiOMKzrL1_0),.clk(gclk));
	jdff dff_A_OuHO2q7r5_0(.dout(w_dff_A_DiOMKzrL1_0),.din(w_dff_A_OuHO2q7r5_0),.clk(gclk));
	jdff dff_A_K7AyFFeR1_0(.dout(w_dff_A_OuHO2q7r5_0),.din(w_dff_A_K7AyFFeR1_0),.clk(gclk));
	jdff dff_A_dwYZuPoa4_0(.dout(w_dff_A_K7AyFFeR1_0),.din(w_dff_A_dwYZuPoa4_0),.clk(gclk));
	jdff dff_A_S50wsJSu9_0(.dout(w_dff_A_dwYZuPoa4_0),.din(w_dff_A_S50wsJSu9_0),.clk(gclk));
	jdff dff_A_7ZMgPdB88_0(.dout(w_n747_2[0]),.din(w_dff_A_7ZMgPdB88_0),.clk(gclk));
	jdff dff_A_uFZ7ilqp2_0(.dout(w_dff_A_7ZMgPdB88_0),.din(w_dff_A_uFZ7ilqp2_0),.clk(gclk));
	jdff dff_A_xoQKAynq0_0(.dout(w_dff_A_uFZ7ilqp2_0),.din(w_dff_A_xoQKAynq0_0),.clk(gclk));
	jdff dff_A_WZJHD5gS9_0(.dout(w_dff_A_xoQKAynq0_0),.din(w_dff_A_WZJHD5gS9_0),.clk(gclk));
	jdff dff_A_NrSQtPIH1_0(.dout(w_dff_A_WZJHD5gS9_0),.din(w_dff_A_NrSQtPIH1_0),.clk(gclk));
	jdff dff_A_B3mCpQCe6_1(.dout(w_n747_2[1]),.din(w_dff_A_B3mCpQCe6_1),.clk(gclk));
	jdff dff_A_oBdeOxA45_1(.dout(w_dff_A_B3mCpQCe6_1),.din(w_dff_A_oBdeOxA45_1),.clk(gclk));
	jdff dff_A_zkzI0MoW7_1(.dout(w_dff_A_oBdeOxA45_1),.din(w_dff_A_zkzI0MoW7_1),.clk(gclk));
	jdff dff_A_jSgBYgoR4_1(.dout(w_dff_A_zkzI0MoW7_1),.din(w_dff_A_jSgBYgoR4_1),.clk(gclk));
	jdff dff_A_FBWiu6sb3_1(.dout(w_dff_A_jSgBYgoR4_1),.din(w_dff_A_FBWiu6sb3_1),.clk(gclk));
	jdff dff_A_LYNo2ASk7_1(.dout(w_dff_A_FBWiu6sb3_1),.din(w_dff_A_LYNo2ASk7_1),.clk(gclk));
	jdff dff_A_ACD1nKsc4_1(.dout(w_dff_A_LYNo2ASk7_1),.din(w_dff_A_ACD1nKsc4_1),.clk(gclk));
	jdff dff_A_GAKN05Nq0_1(.dout(w_dff_A_ACD1nKsc4_1),.din(w_dff_A_GAKN05Nq0_1),.clk(gclk));
	jdff dff_A_46KeFG3T5_1(.dout(w_dff_A_GAKN05Nq0_1),.din(w_dff_A_46KeFG3T5_1),.clk(gclk));
	jdff dff_B_mqZHnNjT7_0(.din(n1196),.dout(w_dff_B_mqZHnNjT7_0),.clk(gclk));
	jdff dff_B_zVHJlvIO3_0(.din(w_dff_B_mqZHnNjT7_0),.dout(w_dff_B_zVHJlvIO3_0),.clk(gclk));
	jdff dff_B_xUFYXKgH2_0(.din(w_dff_B_zVHJlvIO3_0),.dout(w_dff_B_xUFYXKgH2_0),.clk(gclk));
	jdff dff_B_XUtwgCBg4_0(.din(w_dff_B_xUFYXKgH2_0),.dout(w_dff_B_XUtwgCBg4_0),.clk(gclk));
	jdff dff_B_l6lm0sY73_0(.din(w_dff_B_XUtwgCBg4_0),.dout(w_dff_B_l6lm0sY73_0),.clk(gclk));
	jdff dff_B_iuwMfApg1_0(.din(w_dff_B_l6lm0sY73_0),.dout(w_dff_B_iuwMfApg1_0),.clk(gclk));
	jdff dff_B_huMTkWf36_0(.din(w_dff_B_iuwMfApg1_0),.dout(w_dff_B_huMTkWf36_0),.clk(gclk));
	jdff dff_B_jhuFUAdV5_0(.din(w_dff_B_huMTkWf36_0),.dout(w_dff_B_jhuFUAdV5_0),.clk(gclk));
	jdff dff_B_KOlIZRFo4_0(.din(w_dff_B_jhuFUAdV5_0),.dout(w_dff_B_KOlIZRFo4_0),.clk(gclk));
	jdff dff_B_D592iDCk4_0(.din(w_dff_B_KOlIZRFo4_0),.dout(w_dff_B_D592iDCk4_0),.clk(gclk));
	jdff dff_B_zqJOUQM15_0(.din(w_dff_B_D592iDCk4_0),.dout(w_dff_B_zqJOUQM15_0),.clk(gclk));
	jdff dff_B_2XMIVhUw3_0(.din(w_dff_B_zqJOUQM15_0),.dout(w_dff_B_2XMIVhUw3_0),.clk(gclk));
	jdff dff_B_kfM8BBMH2_0(.din(n1195),.dout(w_dff_B_kfM8BBMH2_0),.clk(gclk));
	jdff dff_B_rRV3MrUo5_0(.din(w_dff_B_kfM8BBMH2_0),.dout(w_dff_B_rRV3MrUo5_0),.clk(gclk));
	jdff dff_B_xtfFS7ya0_0(.din(w_dff_B_rRV3MrUo5_0),.dout(w_dff_B_xtfFS7ya0_0),.clk(gclk));
	jdff dff_B_KwgV3T4n3_0(.din(w_dff_B_xtfFS7ya0_0),.dout(w_dff_B_KwgV3T4n3_0),.clk(gclk));
	jdff dff_B_RQTw2CmT4_1(.din(G115),.dout(w_dff_B_RQTw2CmT4_1),.clk(gclk));
	jdff dff_B_CjpD4YzR1_1(.din(w_dff_B_RQTw2CmT4_1),.dout(w_dff_B_CjpD4YzR1_1),.clk(gclk));
	jdff dff_A_b3F2XRIP3_0(.dout(w_n751_0[0]),.din(w_dff_A_b3F2XRIP3_0),.clk(gclk));
	jdff dff_A_i2MhnlsV3_2(.dout(w_n751_0[2]),.din(w_dff_A_i2MhnlsV3_2),.clk(gclk));
	jdff dff_A_SswdMDB54_2(.dout(w_dff_A_i2MhnlsV3_2),.din(w_dff_A_SswdMDB54_2),.clk(gclk));
	jdff dff_A_wqPfTT917_2(.dout(w_dff_A_SswdMDB54_2),.din(w_dff_A_wqPfTT917_2),.clk(gclk));
	jdff dff_A_uIcXy7Ld2_2(.dout(w_dff_A_wqPfTT917_2),.din(w_dff_A_uIcXy7Ld2_2),.clk(gclk));
	jdff dff_B_KmBIXJZD9_1(.din(n929),.dout(w_dff_B_KmBIXJZD9_1),.clk(gclk));
	jdff dff_B_vABTjAim3_1(.din(w_dff_B_KmBIXJZD9_1),.dout(w_dff_B_vABTjAim3_1),.clk(gclk));
	jdff dff_B_lE0fHd272_1(.din(w_dff_B_vABTjAim3_1),.dout(w_dff_B_lE0fHd272_1),.clk(gclk));
	jdff dff_B_mG22AAd94_1(.din(w_dff_B_lE0fHd272_1),.dout(w_dff_B_mG22AAd94_1),.clk(gclk));
	jdff dff_B_sHr3FexY7_1(.din(w_dff_B_mG22AAd94_1),.dout(w_dff_B_sHr3FexY7_1),.clk(gclk));
	jdff dff_B_ZC0Suado3_1(.din(w_dff_B_sHr3FexY7_1),.dout(w_dff_B_ZC0Suado3_1),.clk(gclk));
	jdff dff_B_1MX1hrpz6_1(.din(w_dff_B_ZC0Suado3_1),.dout(w_dff_B_1MX1hrpz6_1),.clk(gclk));
	jdff dff_B_n8WOJk9M0_1(.din(w_dff_B_1MX1hrpz6_1),.dout(w_dff_B_n8WOJk9M0_1),.clk(gclk));
	jdff dff_B_gcQBnGqx9_1(.din(n931),.dout(w_dff_B_gcQBnGqx9_1),.clk(gclk));
	jdff dff_B_5BahILlN4_1(.din(w_dff_B_gcQBnGqx9_1),.dout(w_dff_B_5BahILlN4_1),.clk(gclk));
	jdff dff_B_0DZi2YVH6_1(.din(w_dff_B_5BahILlN4_1),.dout(w_dff_B_0DZi2YVH6_1),.clk(gclk));
	jdff dff_B_eG2B8B5I5_1(.din(w_dff_B_0DZi2YVH6_1),.dout(w_dff_B_eG2B8B5I5_1),.clk(gclk));
	jdff dff_B_X582oZyd9_1(.din(w_dff_B_eG2B8B5I5_1),.dout(w_dff_B_X582oZyd9_1),.clk(gclk));
	jdff dff_B_P2Tlkxjg6_1(.din(w_dff_B_X582oZyd9_1),.dout(w_dff_B_P2Tlkxjg6_1),.clk(gclk));
	jdff dff_B_tXbYhoQQ6_1(.din(w_dff_B_P2Tlkxjg6_1),.dout(w_dff_B_tXbYhoQQ6_1),.clk(gclk));
	jdff dff_B_VezKcuRz7_1(.din(w_dff_B_tXbYhoQQ6_1),.dout(w_dff_B_VezKcuRz7_1),.clk(gclk));
	jdff dff_B_VH3KISCb2_1(.din(w_dff_B_VezKcuRz7_1),.dout(w_dff_B_VH3KISCb2_1),.clk(gclk));
	jdff dff_B_Apat5Bi87_1(.din(w_dff_B_VH3KISCb2_1),.dout(w_dff_B_Apat5Bi87_1),.clk(gclk));
	jdff dff_B_NtUiBiVq2_0(.din(n935),.dout(w_dff_B_NtUiBiVq2_0),.clk(gclk));
	jdff dff_A_2Sfp7Nqg3_1(.dout(w_G4_0[1]),.din(w_dff_A_2Sfp7Nqg3_1),.clk(gclk));
	jdff dff_A_5jwWtI1F4_1(.dout(w_dff_A_2Sfp7Nqg3_1),.din(w_dff_A_5jwWtI1F4_1),.clk(gclk));
	jdff dff_A_yDS8hk1Y9_1(.dout(w_dff_A_5jwWtI1F4_1),.din(w_dff_A_yDS8hk1Y9_1),.clk(gclk));
	jdff dff_A_W9Ozmo8a0_1(.dout(w_dff_A_yDS8hk1Y9_1),.din(w_dff_A_W9Ozmo8a0_1),.clk(gclk));
	jdff dff_A_lYjkwI1V6_1(.dout(w_dff_A_W9Ozmo8a0_1),.din(w_dff_A_lYjkwI1V6_1),.clk(gclk));
	jdff dff_A_9Gi1pbWn9_1(.dout(w_dff_A_lYjkwI1V6_1),.din(w_dff_A_9Gi1pbWn9_1),.clk(gclk));
	jdff dff_B_g3IckT5T9_3(.din(G4),.dout(w_dff_B_g3IckT5T9_3),.clk(gclk));
	jdff dff_B_4eX0Co9w0_3(.din(w_dff_B_g3IckT5T9_3),.dout(w_dff_B_4eX0Co9w0_3),.clk(gclk));
	jdff dff_B_2CffgmCk6_3(.din(w_dff_B_4eX0Co9w0_3),.dout(w_dff_B_2CffgmCk6_3),.clk(gclk));
	jdff dff_B_K8ORnOKd0_3(.din(w_dff_B_2CffgmCk6_3),.dout(w_dff_B_K8ORnOKd0_3),.clk(gclk));
	jdff dff_B_DAKqQrDa0_2(.din(n932),.dout(w_dff_B_DAKqQrDa0_2),.clk(gclk));
	jdff dff_B_LuVljHUT6_2(.din(w_dff_B_DAKqQrDa0_2),.dout(w_dff_B_LuVljHUT6_2),.clk(gclk));
	jdff dff_B_Ppqaer007_2(.din(w_dff_B_LuVljHUT6_2),.dout(w_dff_B_Ppqaer007_2),.clk(gclk));
	jdff dff_B_gNUNXADe4_2(.din(w_dff_B_Ppqaer007_2),.dout(w_dff_B_gNUNXADe4_2),.clk(gclk));
	jdff dff_B_ricpX7Rv7_2(.din(w_dff_B_gNUNXADe4_2),.dout(w_dff_B_ricpX7Rv7_2),.clk(gclk));
	jdff dff_B_ugLXr8VB4_2(.din(w_dff_B_ricpX7Rv7_2),.dout(w_dff_B_ugLXr8VB4_2),.clk(gclk));
	jdff dff_B_gknoEShI4_2(.din(w_dff_B_ugLXr8VB4_2),.dout(w_dff_B_gknoEShI4_2),.clk(gclk));
	jdff dff_B_RFcK7kxy9_2(.din(w_dff_B_gknoEShI4_2),.dout(w_dff_B_RFcK7kxy9_2),.clk(gclk));
	jdff dff_B_yjprOUEj0_2(.din(w_dff_B_RFcK7kxy9_2),.dout(w_dff_B_yjprOUEj0_2),.clk(gclk));
	jdff dff_A_SgNHVH5Z3_1(.dout(w_n747_1[1]),.din(w_dff_A_SgNHVH5Z3_1),.clk(gclk));
	jdff dff_A_iFVfDNt66_1(.dout(w_dff_A_SgNHVH5Z3_1),.din(w_dff_A_iFVfDNt66_1),.clk(gclk));
	jdff dff_A_vsXEra7e3_1(.dout(w_dff_A_iFVfDNt66_1),.din(w_dff_A_vsXEra7e3_1),.clk(gclk));
	jdff dff_A_W2DtHLXz9_2(.dout(w_n747_1[2]),.din(w_dff_A_W2DtHLXz9_2),.clk(gclk));
	jdff dff_A_pvl3mcel0_2(.dout(w_dff_A_W2DtHLXz9_2),.din(w_dff_A_pvl3mcel0_2),.clk(gclk));
	jdff dff_A_03Umby7w5_2(.dout(w_dff_A_pvl3mcel0_2),.din(w_dff_A_03Umby7w5_2),.clk(gclk));
	jdff dff_A_iT9fQLBz5_2(.dout(w_dff_A_03Umby7w5_2),.din(w_dff_A_iT9fQLBz5_2),.clk(gclk));
	jdff dff_A_v34TugCi6_0(.dout(w_n747_0[0]),.din(w_dff_A_v34TugCi6_0),.clk(gclk));
	jdff dff_A_mBnxGzrR9_0(.dout(w_dff_A_v34TugCi6_0),.din(w_dff_A_mBnxGzrR9_0),.clk(gclk));
	jdff dff_A_CSeudXrA7_0(.dout(w_dff_A_mBnxGzrR9_0),.din(w_dff_A_CSeudXrA7_0),.clk(gclk));
	jdff dff_A_thU9StEt9_0(.dout(w_dff_A_CSeudXrA7_0),.din(w_dff_A_thU9StEt9_0),.clk(gclk));
	jdff dff_A_gIZTJ2SD4_0(.dout(w_dff_A_thU9StEt9_0),.din(w_dff_A_gIZTJ2SD4_0),.clk(gclk));
	jdff dff_A_4GamQ0Jp2_0(.dout(w_dff_A_gIZTJ2SD4_0),.din(w_dff_A_4GamQ0Jp2_0),.clk(gclk));
	jdff dff_A_hvvYB3n21_0(.dout(w_dff_A_4GamQ0Jp2_0),.din(w_dff_A_hvvYB3n21_0),.clk(gclk));
	jdff dff_A_TWQEc8XZ8_0(.dout(w_dff_A_hvvYB3n21_0),.din(w_dff_A_TWQEc8XZ8_0),.clk(gclk));
	jdff dff_A_pczc4ae96_0(.dout(w_dff_A_TWQEc8XZ8_0),.din(w_dff_A_pczc4ae96_0),.clk(gclk));
	jdff dff_A_BmndQNu78_0(.dout(w_dff_A_pczc4ae96_0),.din(w_dff_A_BmndQNu78_0),.clk(gclk));
	jdff dff_A_vPbLhE3F2_0(.dout(w_dff_A_BmndQNu78_0),.din(w_dff_A_vPbLhE3F2_0),.clk(gclk));
	jdff dff_A_75gcu1mL0_0(.dout(w_dff_A_vPbLhE3F2_0),.din(w_dff_A_75gcu1mL0_0),.clk(gclk));
	jdff dff_A_4H65fA2y3_0(.dout(w_dff_A_75gcu1mL0_0),.din(w_dff_A_4H65fA2y3_0),.clk(gclk));
	jdff dff_A_sJR2gL3C3_1(.dout(w_n747_0[1]),.din(w_dff_A_sJR2gL3C3_1),.clk(gclk));
	jdff dff_A_CgSBUOBR4_1(.dout(w_dff_A_sJR2gL3C3_1),.din(w_dff_A_CgSBUOBR4_1),.clk(gclk));
	jdff dff_A_YtMPeKmw1_1(.dout(w_dff_A_CgSBUOBR4_1),.din(w_dff_A_YtMPeKmw1_1),.clk(gclk));
	jdff dff_A_PNQ1jMf32_1(.dout(w_dff_A_YtMPeKmw1_1),.din(w_dff_A_PNQ1jMf32_1),.clk(gclk));
	jdff dff_A_lWU3J0Ge3_1(.dout(w_dff_A_PNQ1jMf32_1),.din(w_dff_A_lWU3J0Ge3_1),.clk(gclk));
	jdff dff_A_evCurInq7_1(.dout(w_dff_A_lWU3J0Ge3_1),.din(w_dff_A_evCurInq7_1),.clk(gclk));
	jdff dff_A_gZRPnmG56_1(.dout(w_dff_A_evCurInq7_1),.din(w_dff_A_gZRPnmG56_1),.clk(gclk));
	jdff dff_B_5RGa8LMP9_1(.din(n1388),.dout(w_dff_B_5RGa8LMP9_1),.clk(gclk));
	jdff dff_B_HxLhjqH88_1(.din(w_dff_B_5RGa8LMP9_1),.dout(w_dff_B_HxLhjqH88_1),.clk(gclk));
	jdff dff_B_74sPFeaY7_1(.din(w_dff_B_HxLhjqH88_1),.dout(w_dff_B_74sPFeaY7_1),.clk(gclk));
	jdff dff_B_27JaNkQl8_1(.din(w_dff_B_74sPFeaY7_1),.dout(w_dff_B_27JaNkQl8_1),.clk(gclk));
	jdff dff_B_8oTVzDsz9_1(.din(w_dff_B_27JaNkQl8_1),.dout(w_dff_B_8oTVzDsz9_1),.clk(gclk));
	jdff dff_B_YGBlsYku1_1(.din(w_dff_B_8oTVzDsz9_1),.dout(w_dff_B_YGBlsYku1_1),.clk(gclk));
	jdff dff_B_uxi4rQSK1_1(.din(w_dff_B_YGBlsYku1_1),.dout(w_dff_B_uxi4rQSK1_1),.clk(gclk));
	jdff dff_B_TBbHLIV76_1(.din(w_dff_B_uxi4rQSK1_1),.dout(w_dff_B_TBbHLIV76_1),.clk(gclk));
	jdff dff_B_Uvt2fEHQ9_1(.din(w_dff_B_TBbHLIV76_1),.dout(w_dff_B_Uvt2fEHQ9_1),.clk(gclk));
	jdff dff_B_Hmj92KV31_1(.din(w_dff_B_Uvt2fEHQ9_1),.dout(w_dff_B_Hmj92KV31_1),.clk(gclk));
	jdff dff_B_ax4oRnWb1_1(.din(w_dff_B_Hmj92KV31_1),.dout(w_dff_B_ax4oRnWb1_1),.clk(gclk));
	jdff dff_B_gGG5PQ2J1_1(.din(w_dff_B_ax4oRnWb1_1),.dout(w_dff_B_gGG5PQ2J1_1),.clk(gclk));
	jdff dff_B_q2KJSj7E7_1(.din(w_dff_B_gGG5PQ2J1_1),.dout(w_dff_B_q2KJSj7E7_1),.clk(gclk));
	jdff dff_B_NCck7nZb0_1(.din(w_dff_B_q2KJSj7E7_1),.dout(w_dff_B_NCck7nZb0_1),.clk(gclk));
	jdff dff_B_rW0Q9rgF2_1(.din(w_dff_B_NCck7nZb0_1),.dout(w_dff_B_rW0Q9rgF2_1),.clk(gclk));
	jdff dff_B_aHHJLOyA5_1(.din(w_dff_B_rW0Q9rgF2_1),.dout(w_dff_B_aHHJLOyA5_1),.clk(gclk));
	jdff dff_B_uazdRGXM7_1(.din(w_dff_B_aHHJLOyA5_1),.dout(w_dff_B_uazdRGXM7_1),.clk(gclk));
	jdff dff_B_zOwdtIAm3_1(.din(w_dff_B_uazdRGXM7_1),.dout(w_dff_B_zOwdtIAm3_1),.clk(gclk));
	jdff dff_B_jxny4ArA6_1(.din(w_dff_B_zOwdtIAm3_1),.dout(w_dff_B_jxny4ArA6_1),.clk(gclk));
	jdff dff_B_qGfkV9Ns6_1(.din(n1539),.dout(w_dff_B_qGfkV9Ns6_1),.clk(gclk));
	jdff dff_B_eGcvvx9E1_1(.din(w_dff_B_qGfkV9Ns6_1),.dout(w_dff_B_eGcvvx9E1_1),.clk(gclk));
	jdff dff_B_4f5py8GE0_1(.din(w_dff_B_eGcvvx9E1_1),.dout(w_dff_B_4f5py8GE0_1),.clk(gclk));
	jdff dff_B_S69VBAbw0_1(.din(w_dff_B_4f5py8GE0_1),.dout(w_dff_B_S69VBAbw0_1),.clk(gclk));
	jdff dff_B_2qZ4r7xt4_1(.din(w_dff_B_S69VBAbw0_1),.dout(w_dff_B_2qZ4r7xt4_1),.clk(gclk));
	jdff dff_B_wHqDGhkw3_1(.din(w_dff_B_2qZ4r7xt4_1),.dout(w_dff_B_wHqDGhkw3_1),.clk(gclk));
	jdff dff_B_gdxU8hfz6_1(.din(w_dff_B_wHqDGhkw3_1),.dout(w_dff_B_gdxU8hfz6_1),.clk(gclk));
	jdff dff_B_t2cExOin3_1(.din(w_dff_B_gdxU8hfz6_1),.dout(w_dff_B_t2cExOin3_1),.clk(gclk));
	jdff dff_B_gMbUnIvW5_1(.din(w_dff_B_t2cExOin3_1),.dout(w_dff_B_gMbUnIvW5_1),.clk(gclk));
	jdff dff_B_7BMQW0dG5_1(.din(w_dff_B_gMbUnIvW5_1),.dout(w_dff_B_7BMQW0dG5_1),.clk(gclk));
	jdff dff_B_5tJKBy3B1_1(.din(w_dff_B_7BMQW0dG5_1),.dout(w_dff_B_5tJKBy3B1_1),.clk(gclk));
	jdff dff_B_Hwg6UBlW5_1(.din(w_dff_B_5tJKBy3B1_1),.dout(w_dff_B_Hwg6UBlW5_1),.clk(gclk));
	jdff dff_B_8dbasd5t4_1(.din(w_dff_B_Hwg6UBlW5_1),.dout(w_dff_B_8dbasd5t4_1),.clk(gclk));
	jdff dff_B_FStOYtq33_1(.din(w_dff_B_8dbasd5t4_1),.dout(w_dff_B_FStOYtq33_1),.clk(gclk));
	jdff dff_B_vYN0ROCC7_1(.din(w_dff_B_FStOYtq33_1),.dout(w_dff_B_vYN0ROCC7_1),.clk(gclk));
	jdff dff_B_UR5UkB7Z1_1(.din(w_dff_B_vYN0ROCC7_1),.dout(w_dff_B_UR5UkB7Z1_1),.clk(gclk));
	jdff dff_B_crLcOZlU7_1(.din(w_dff_B_UR5UkB7Z1_1),.dout(w_dff_B_crLcOZlU7_1),.clk(gclk));
	jdff dff_B_OU4yaq7L3_1(.din(w_dff_B_crLcOZlU7_1),.dout(w_dff_B_OU4yaq7L3_1),.clk(gclk));
	jdff dff_B_nIpOyoey8_1(.din(w_dff_B_OU4yaq7L3_1),.dout(w_dff_B_nIpOyoey8_1),.clk(gclk));
	jdff dff_B_fRM4cHqM2_0(.din(n1614),.dout(w_dff_B_fRM4cHqM2_0),.clk(gclk));
	jdff dff_B_kitt4geg0_0(.din(w_dff_B_fRM4cHqM2_0),.dout(w_dff_B_kitt4geg0_0),.clk(gclk));
	jdff dff_B_liwupeu76_0(.din(w_dff_B_kitt4geg0_0),.dout(w_dff_B_liwupeu76_0),.clk(gclk));
	jdff dff_B_bvWzRpva7_0(.din(w_dff_B_liwupeu76_0),.dout(w_dff_B_bvWzRpva7_0),.clk(gclk));
	jdff dff_B_kbArhJW13_0(.din(w_dff_B_bvWzRpva7_0),.dout(w_dff_B_kbArhJW13_0),.clk(gclk));
	jdff dff_B_liTFATlW4_0(.din(w_dff_B_kbArhJW13_0),.dout(w_dff_B_liTFATlW4_0),.clk(gclk));
	jdff dff_B_Kj340Lus6_0(.din(w_dff_B_liTFATlW4_0),.dout(w_dff_B_Kj340Lus6_0),.clk(gclk));
	jdff dff_B_1fzNq9SA6_0(.din(w_dff_B_Kj340Lus6_0),.dout(w_dff_B_1fzNq9SA6_0),.clk(gclk));
	jdff dff_B_GbUkwzVG5_0(.din(w_dff_B_1fzNq9SA6_0),.dout(w_dff_B_GbUkwzVG5_0),.clk(gclk));
	jdff dff_B_IIaOuqWc4_0(.din(w_dff_B_GbUkwzVG5_0),.dout(w_dff_B_IIaOuqWc4_0),.clk(gclk));
	jdff dff_B_MC0H8Sk78_0(.din(w_dff_B_IIaOuqWc4_0),.dout(w_dff_B_MC0H8Sk78_0),.clk(gclk));
	jdff dff_B_UqiGo2xb0_0(.din(w_dff_B_MC0H8Sk78_0),.dout(w_dff_B_UqiGo2xb0_0),.clk(gclk));
	jdff dff_B_h8W123E12_0(.din(w_dff_B_UqiGo2xb0_0),.dout(w_dff_B_h8W123E12_0),.clk(gclk));
	jdff dff_B_vpAbq5Po0_0(.din(w_dff_B_h8W123E12_0),.dout(w_dff_B_vpAbq5Po0_0),.clk(gclk));
	jdff dff_B_dK9GxTrQ6_0(.din(w_dff_B_vpAbq5Po0_0),.dout(w_dff_B_dK9GxTrQ6_0),.clk(gclk));
	jdff dff_B_P8zjaeIw7_0(.din(w_dff_B_dK9GxTrQ6_0),.dout(w_dff_B_P8zjaeIw7_0),.clk(gclk));
	jdff dff_B_lZI4WODN9_0(.din(w_dff_B_P8zjaeIw7_0),.dout(w_dff_B_lZI4WODN9_0),.clk(gclk));
	jdff dff_B_I5IH0MMJ2_0(.din(w_dff_B_lZI4WODN9_0),.dout(w_dff_B_I5IH0MMJ2_0),.clk(gclk));
	jdff dff_B_4rHYBAdE5_0(.din(w_dff_B_I5IH0MMJ2_0),.dout(w_dff_B_4rHYBAdE5_0),.clk(gclk));
	jdff dff_B_h1ssQCLb9_0(.din(n1613),.dout(w_dff_B_h1ssQCLb9_0),.clk(gclk));
	jdff dff_A_62QowrCK3_1(.dout(w_n797_1[1]),.din(w_dff_A_62QowrCK3_1),.clk(gclk));
	jdff dff_A_44HAr5Qh2_1(.dout(w_dff_A_62QowrCK3_1),.din(w_dff_A_44HAr5Qh2_1),.clk(gclk));
	jdff dff_A_4j65zlAi8_1(.dout(w_dff_A_44HAr5Qh2_1),.din(w_dff_A_4j65zlAi8_1),.clk(gclk));
	jdff dff_A_e1fNy4Ma2_1(.dout(w_dff_A_4j65zlAi8_1),.din(w_dff_A_e1fNy4Ma2_1),.clk(gclk));
	jdff dff_A_kBPdLRwq7_1(.dout(w_dff_A_e1fNy4Ma2_1),.din(w_dff_A_kBPdLRwq7_1),.clk(gclk));
	jdff dff_A_dwd6FNwR2_1(.dout(w_dff_A_kBPdLRwq7_1),.din(w_dff_A_dwd6FNwR2_1),.clk(gclk));
	jdff dff_A_4ZMbzVX56_1(.dout(w_dff_A_dwd6FNwR2_1),.din(w_dff_A_4ZMbzVX56_1),.clk(gclk));
	jdff dff_A_cKUj5x8V8_1(.dout(w_dff_A_4ZMbzVX56_1),.din(w_dff_A_cKUj5x8V8_1),.clk(gclk));
	jdff dff_A_LzInWdmJ3_1(.dout(w_dff_A_cKUj5x8V8_1),.din(w_dff_A_LzInWdmJ3_1),.clk(gclk));
	jdff dff_A_s6I1a9Su3_1(.dout(w_dff_A_LzInWdmJ3_1),.din(w_dff_A_s6I1a9Su3_1),.clk(gclk));
	jdff dff_A_sOa87aUo4_1(.dout(w_dff_A_s6I1a9Su3_1),.din(w_dff_A_sOa87aUo4_1),.clk(gclk));
	jdff dff_A_oNDKrWIW1_1(.dout(w_dff_A_sOa87aUo4_1),.din(w_dff_A_oNDKrWIW1_1),.clk(gclk));
	jdff dff_A_3gVy0WKl4_1(.dout(w_dff_A_oNDKrWIW1_1),.din(w_dff_A_3gVy0WKl4_1),.clk(gclk));
	jdff dff_A_1PVE3DRf5_1(.dout(w_dff_A_3gVy0WKl4_1),.din(w_dff_A_1PVE3DRf5_1),.clk(gclk));
	jdff dff_A_ZBIsONhY0_2(.dout(w_n797_1[2]),.din(w_dff_A_ZBIsONhY0_2),.clk(gclk));
	jdff dff_A_LSJWrf1e7_2(.dout(w_dff_A_ZBIsONhY0_2),.din(w_dff_A_LSJWrf1e7_2),.clk(gclk));
	jdff dff_A_P1hkd3J18_2(.dout(w_dff_A_LSJWrf1e7_2),.din(w_dff_A_P1hkd3J18_2),.clk(gclk));
	jdff dff_A_Vrm60Fkm3_2(.dout(w_dff_A_P1hkd3J18_2),.din(w_dff_A_Vrm60Fkm3_2),.clk(gclk));
	jdff dff_A_64DEMkZ58_2(.dout(w_dff_A_Vrm60Fkm3_2),.din(w_dff_A_64DEMkZ58_2),.clk(gclk));
	jdff dff_A_1bZSorDu6_2(.dout(w_dff_A_64DEMkZ58_2),.din(w_dff_A_1bZSorDu6_2),.clk(gclk));
	jdff dff_A_JUoG50SJ8_2(.dout(w_dff_A_1bZSorDu6_2),.din(w_dff_A_JUoG50SJ8_2),.clk(gclk));
	jdff dff_A_7praynRV6_2(.dout(w_dff_A_JUoG50SJ8_2),.din(w_dff_A_7praynRV6_2),.clk(gclk));
	jdff dff_A_7CIQBXyA2_2(.dout(w_dff_A_7praynRV6_2),.din(w_dff_A_7CIQBXyA2_2),.clk(gclk));
	jdff dff_A_hL4526bv5_2(.dout(w_dff_A_7CIQBXyA2_2),.din(w_dff_A_hL4526bv5_2),.clk(gclk));
	jdff dff_A_qAJnDHiJ4_1(.dout(w_n797_0[1]),.din(w_dff_A_qAJnDHiJ4_1),.clk(gclk));
	jdff dff_A_K9DS2KSS3_1(.dout(w_dff_A_qAJnDHiJ4_1),.din(w_dff_A_K9DS2KSS3_1),.clk(gclk));
	jdff dff_A_qlCUkixp0_1(.dout(w_dff_A_K9DS2KSS3_1),.din(w_dff_A_qlCUkixp0_1),.clk(gclk));
	jdff dff_A_VFR3Wbyt5_1(.dout(w_dff_A_qlCUkixp0_1),.din(w_dff_A_VFR3Wbyt5_1),.clk(gclk));
	jdff dff_A_mroUqqRB1_1(.dout(w_dff_A_VFR3Wbyt5_1),.din(w_dff_A_mroUqqRB1_1),.clk(gclk));
	jdff dff_A_KglxCDra0_1(.dout(w_dff_A_mroUqqRB1_1),.din(w_dff_A_KglxCDra0_1),.clk(gclk));
	jdff dff_A_O26fNIRH7_1(.dout(w_dff_A_KglxCDra0_1),.din(w_dff_A_O26fNIRH7_1),.clk(gclk));
	jdff dff_A_IPQ2NA3F8_1(.dout(w_dff_A_O26fNIRH7_1),.din(w_dff_A_IPQ2NA3F8_1),.clk(gclk));
	jdff dff_A_4JxQ5gnA4_1(.dout(w_dff_A_IPQ2NA3F8_1),.din(w_dff_A_4JxQ5gnA4_1),.clk(gclk));
	jdff dff_A_r2w5kEW48_1(.dout(w_dff_A_4JxQ5gnA4_1),.din(w_dff_A_r2w5kEW48_1),.clk(gclk));
	jdff dff_A_vufs09fJ5_1(.dout(w_dff_A_r2w5kEW48_1),.din(w_dff_A_vufs09fJ5_1),.clk(gclk));
	jdff dff_A_V3S91piA1_2(.dout(w_n797_0[2]),.din(w_dff_A_V3S91piA1_2),.clk(gclk));
	jdff dff_B_zVz0njuI9_3(.din(n797),.dout(w_dff_B_zVz0njuI9_3),.clk(gclk));
	jdff dff_B_853ihHdN7_3(.din(w_dff_B_zVz0njuI9_3),.dout(w_dff_B_853ihHdN7_3),.clk(gclk));
	jdff dff_B_l2KaA5Gl2_3(.din(w_dff_B_853ihHdN7_3),.dout(w_dff_B_l2KaA5Gl2_3),.clk(gclk));
	jdff dff_B_9YBJuyUI5_3(.din(w_dff_B_l2KaA5Gl2_3),.dout(w_dff_B_9YBJuyUI5_3),.clk(gclk));
	jdff dff_B_JRRagGoi5_3(.din(w_dff_B_9YBJuyUI5_3),.dout(w_dff_B_JRRagGoi5_3),.clk(gclk));
	jdff dff_B_p44IFa8m3_3(.din(w_dff_B_JRRagGoi5_3),.dout(w_dff_B_p44IFa8m3_3),.clk(gclk));
	jdff dff_A_kio7HzqD0_1(.dout(w_n793_1[1]),.din(w_dff_A_kio7HzqD0_1),.clk(gclk));
	jdff dff_A_89JhneNF5_1(.dout(w_dff_A_kio7HzqD0_1),.din(w_dff_A_89JhneNF5_1),.clk(gclk));
	jdff dff_A_oxxJBvXz8_1(.dout(w_dff_A_89JhneNF5_1),.din(w_dff_A_oxxJBvXz8_1),.clk(gclk));
	jdff dff_A_V93YUqWD9_1(.dout(w_dff_A_oxxJBvXz8_1),.din(w_dff_A_V93YUqWD9_1),.clk(gclk));
	jdff dff_A_Cgt4QIfM0_1(.dout(w_dff_A_V93YUqWD9_1),.din(w_dff_A_Cgt4QIfM0_1),.clk(gclk));
	jdff dff_A_9AN431Ud5_1(.dout(w_dff_A_Cgt4QIfM0_1),.din(w_dff_A_9AN431Ud5_1),.clk(gclk));
	jdff dff_A_IMcBrGU46_1(.dout(w_dff_A_9AN431Ud5_1),.din(w_dff_A_IMcBrGU46_1),.clk(gclk));
	jdff dff_A_waABEiXy6_1(.dout(w_dff_A_IMcBrGU46_1),.din(w_dff_A_waABEiXy6_1),.clk(gclk));
	jdff dff_A_23tbKixm2_1(.dout(w_dff_A_waABEiXy6_1),.din(w_dff_A_23tbKixm2_1),.clk(gclk));
	jdff dff_A_vIgoic5m5_1(.dout(w_dff_A_23tbKixm2_1),.din(w_dff_A_vIgoic5m5_1),.clk(gclk));
	jdff dff_A_sazGto2U8_1(.dout(w_dff_A_vIgoic5m5_1),.din(w_dff_A_sazGto2U8_1),.clk(gclk));
	jdff dff_A_shYT65ez1_1(.dout(w_dff_A_sazGto2U8_1),.din(w_dff_A_shYT65ez1_1),.clk(gclk));
	jdff dff_A_RKl2ve8Q2_1(.dout(w_dff_A_shYT65ez1_1),.din(w_dff_A_RKl2ve8Q2_1),.clk(gclk));
	jdff dff_A_wYf4CRIS1_1(.dout(w_dff_A_RKl2ve8Q2_1),.din(w_dff_A_wYf4CRIS1_1),.clk(gclk));
	jdff dff_A_UVlzuZWb8_2(.dout(w_n793_1[2]),.din(w_dff_A_UVlzuZWb8_2),.clk(gclk));
	jdff dff_A_QzRlgLRO8_2(.dout(w_dff_A_UVlzuZWb8_2),.din(w_dff_A_QzRlgLRO8_2),.clk(gclk));
	jdff dff_A_yzc1uo0F6_2(.dout(w_dff_A_QzRlgLRO8_2),.din(w_dff_A_yzc1uo0F6_2),.clk(gclk));
	jdff dff_A_eEqAMYCR9_2(.dout(w_dff_A_yzc1uo0F6_2),.din(w_dff_A_eEqAMYCR9_2),.clk(gclk));
	jdff dff_A_XYjok7qO5_2(.dout(w_dff_A_eEqAMYCR9_2),.din(w_dff_A_XYjok7qO5_2),.clk(gclk));
	jdff dff_A_y9yAjSAU3_2(.dout(w_dff_A_XYjok7qO5_2),.din(w_dff_A_y9yAjSAU3_2),.clk(gclk));
	jdff dff_A_PGi66FSw6_2(.dout(w_dff_A_y9yAjSAU3_2),.din(w_dff_A_PGi66FSw6_2),.clk(gclk));
	jdff dff_A_isx0Vjju4_2(.dout(w_dff_A_PGi66FSw6_2),.din(w_dff_A_isx0Vjju4_2),.clk(gclk));
	jdff dff_A_SVYFXeQF0_2(.dout(w_dff_A_isx0Vjju4_2),.din(w_dff_A_SVYFXeQF0_2),.clk(gclk));
	jdff dff_A_0Wy3drpl8_2(.dout(w_dff_A_SVYFXeQF0_2),.din(w_dff_A_0Wy3drpl8_2),.clk(gclk));
	jdff dff_A_jkVu3gCc7_1(.dout(w_n793_0[1]),.din(w_dff_A_jkVu3gCc7_1),.clk(gclk));
	jdff dff_A_M74dmBav1_1(.dout(w_dff_A_jkVu3gCc7_1),.din(w_dff_A_M74dmBav1_1),.clk(gclk));
	jdff dff_A_KelRrALB2_1(.dout(w_dff_A_M74dmBav1_1),.din(w_dff_A_KelRrALB2_1),.clk(gclk));
	jdff dff_A_PwFCSI5r0_1(.dout(w_dff_A_KelRrALB2_1),.din(w_dff_A_PwFCSI5r0_1),.clk(gclk));
	jdff dff_A_V2Y6lBwb6_1(.dout(w_dff_A_PwFCSI5r0_1),.din(w_dff_A_V2Y6lBwb6_1),.clk(gclk));
	jdff dff_A_8JskB42r8_1(.dout(w_dff_A_V2Y6lBwb6_1),.din(w_dff_A_8JskB42r8_1),.clk(gclk));
	jdff dff_A_kTF9EuCu8_1(.dout(w_dff_A_8JskB42r8_1),.din(w_dff_A_kTF9EuCu8_1),.clk(gclk));
	jdff dff_A_SYAEVGV86_1(.dout(w_dff_A_kTF9EuCu8_1),.din(w_dff_A_SYAEVGV86_1),.clk(gclk));
	jdff dff_A_KbIqXLc50_1(.dout(w_dff_A_SYAEVGV86_1),.din(w_dff_A_KbIqXLc50_1),.clk(gclk));
	jdff dff_A_J17m2agI0_1(.dout(w_dff_A_KbIqXLc50_1),.din(w_dff_A_J17m2agI0_1),.clk(gclk));
	jdff dff_A_dYGaO07l1_1(.dout(w_dff_A_J17m2agI0_1),.din(w_dff_A_dYGaO07l1_1),.clk(gclk));
	jdff dff_A_j69jbkpN2_2(.dout(w_n793_0[2]),.din(w_dff_A_j69jbkpN2_2),.clk(gclk));
	jdff dff_A_HyK6inpt4_2(.dout(w_dff_A_j69jbkpN2_2),.din(w_dff_A_HyK6inpt4_2),.clk(gclk));
	jdff dff_A_5PWCTDXZ9_2(.dout(w_dff_A_HyK6inpt4_2),.din(w_dff_A_5PWCTDXZ9_2),.clk(gclk));
	jdff dff_A_AeEiZwLg7_2(.dout(w_dff_A_5PWCTDXZ9_2),.din(w_dff_A_AeEiZwLg7_2),.clk(gclk));
	jdff dff_B_Vz2IWRYo0_3(.din(n793),.dout(w_dff_B_Vz2IWRYo0_3),.clk(gclk));
	jdff dff_B_lKYooOn52_3(.din(w_dff_B_Vz2IWRYo0_3),.dout(w_dff_B_lKYooOn52_3),.clk(gclk));
	jdff dff_B_7Y5UojCy3_3(.din(w_dff_B_lKYooOn52_3),.dout(w_dff_B_7Y5UojCy3_3),.clk(gclk));
	jdff dff_B_Ki2i9Lgb6_3(.din(w_dff_B_7Y5UojCy3_3),.dout(w_dff_B_Ki2i9Lgb6_3),.clk(gclk));
	jdff dff_B_LsMfgfUp1_3(.din(w_dff_B_Ki2i9Lgb6_3),.dout(w_dff_B_LsMfgfUp1_3),.clk(gclk));
	jdff dff_B_QcBZguBB0_3(.din(w_dff_B_LsMfgfUp1_3),.dout(w_dff_B_QcBZguBB0_3),.clk(gclk));
	jdff dff_B_yK95vB9c5_3(.din(w_dff_B_QcBZguBB0_3),.dout(w_dff_B_yK95vB9c5_3),.clk(gclk));
	jdff dff_A_tXtXJkyC4_2(.dout(w_G4088_0[2]),.din(w_dff_A_tXtXJkyC4_2),.clk(gclk));
	jdff dff_A_bHB1uaTW0_1(.dout(w_G4087_0[1]),.din(w_dff_A_bHB1uaTW0_1),.clk(gclk));
	jdff dff_B_R330pzjb9_0(.din(n1621),.dout(w_dff_B_R330pzjb9_0),.clk(gclk));
	jdff dff_B_416ZNeiT5_0(.din(w_dff_B_R330pzjb9_0),.dout(w_dff_B_416ZNeiT5_0),.clk(gclk));
	jdff dff_B_qHzkM02Y0_0(.din(w_dff_B_416ZNeiT5_0),.dout(w_dff_B_qHzkM02Y0_0),.clk(gclk));
	jdff dff_B_UK0QYkxR1_0(.din(w_dff_B_qHzkM02Y0_0),.dout(w_dff_B_UK0QYkxR1_0),.clk(gclk));
	jdff dff_B_oMITCUFG6_0(.din(w_dff_B_UK0QYkxR1_0),.dout(w_dff_B_oMITCUFG6_0),.clk(gclk));
	jdff dff_B_a5esy9Ro8_0(.din(w_dff_B_oMITCUFG6_0),.dout(w_dff_B_a5esy9Ro8_0),.clk(gclk));
	jdff dff_B_dldAmf1U9_0(.din(w_dff_B_a5esy9Ro8_0),.dout(w_dff_B_dldAmf1U9_0),.clk(gclk));
	jdff dff_B_HU89f4DN3_0(.din(w_dff_B_dldAmf1U9_0),.dout(w_dff_B_HU89f4DN3_0),.clk(gclk));
	jdff dff_B_w8mBglBD0_0(.din(w_dff_B_HU89f4DN3_0),.dout(w_dff_B_w8mBglBD0_0),.clk(gclk));
	jdff dff_B_vZIkUZa78_0(.din(w_dff_B_w8mBglBD0_0),.dout(w_dff_B_vZIkUZa78_0),.clk(gclk));
	jdff dff_B_C30ova2w0_0(.din(w_dff_B_vZIkUZa78_0),.dout(w_dff_B_C30ova2w0_0),.clk(gclk));
	jdff dff_B_lpjfJTRG5_0(.din(w_dff_B_C30ova2w0_0),.dout(w_dff_B_lpjfJTRG5_0),.clk(gclk));
	jdff dff_B_eNMxXgBn3_0(.din(w_dff_B_lpjfJTRG5_0),.dout(w_dff_B_eNMxXgBn3_0),.clk(gclk));
	jdff dff_B_XCIH7Gjk7_0(.din(w_dff_B_eNMxXgBn3_0),.dout(w_dff_B_XCIH7Gjk7_0),.clk(gclk));
	jdff dff_B_5GKH6wMV0_0(.din(w_dff_B_XCIH7Gjk7_0),.dout(w_dff_B_5GKH6wMV0_0),.clk(gclk));
	jdff dff_B_E4TLQkV22_0(.din(w_dff_B_5GKH6wMV0_0),.dout(w_dff_B_E4TLQkV22_0),.clk(gclk));
	jdff dff_B_8PIr0QJx3_0(.din(w_dff_B_E4TLQkV22_0),.dout(w_dff_B_8PIr0QJx3_0),.clk(gclk));
	jdff dff_B_2UCQuvcd7_0(.din(w_dff_B_8PIr0QJx3_0),.dout(w_dff_B_2UCQuvcd7_0),.clk(gclk));
	jdff dff_B_8D5LGT767_0(.din(w_dff_B_2UCQuvcd7_0),.dout(w_dff_B_8D5LGT767_0),.clk(gclk));
	jdff dff_B_RTVcvQFq5_0(.din(n1620),.dout(w_dff_B_RTVcvQFq5_0),.clk(gclk));
	jdff dff_B_J9TBYGZH4_2(.din(G64),.dout(w_dff_B_J9TBYGZH4_2),.clk(gclk));
	jdff dff_B_nFTGIpDI1_2(.din(G14),.dout(w_dff_B_nFTGIpDI1_2),.clk(gclk));
	jdff dff_B_CaICsnEX1_2(.din(w_dff_B_nFTGIpDI1_2),.dout(w_dff_B_CaICsnEX1_2),.clk(gclk));
	jdff dff_A_PGw1EWcz1_1(.dout(w_n843_1[1]),.din(w_dff_A_PGw1EWcz1_1),.clk(gclk));
	jdff dff_A_cq3UHFCW8_1(.dout(w_dff_A_PGw1EWcz1_1),.din(w_dff_A_cq3UHFCW8_1),.clk(gclk));
	jdff dff_A_PVEWL3WN6_1(.dout(w_dff_A_cq3UHFCW8_1),.din(w_dff_A_PVEWL3WN6_1),.clk(gclk));
	jdff dff_A_eiIao9IU9_1(.dout(w_dff_A_PVEWL3WN6_1),.din(w_dff_A_eiIao9IU9_1),.clk(gclk));
	jdff dff_A_TU0tkgSz0_1(.dout(w_dff_A_eiIao9IU9_1),.din(w_dff_A_TU0tkgSz0_1),.clk(gclk));
	jdff dff_A_uOmx0oVi4_1(.dout(w_dff_A_TU0tkgSz0_1),.din(w_dff_A_uOmx0oVi4_1),.clk(gclk));
	jdff dff_A_KKUldiPv3_1(.dout(w_dff_A_uOmx0oVi4_1),.din(w_dff_A_KKUldiPv3_1),.clk(gclk));
	jdff dff_A_vqAPTctO8_1(.dout(w_dff_A_KKUldiPv3_1),.din(w_dff_A_vqAPTctO8_1),.clk(gclk));
	jdff dff_A_07gJrxt32_1(.dout(w_dff_A_vqAPTctO8_1),.din(w_dff_A_07gJrxt32_1),.clk(gclk));
	jdff dff_A_7lNkLDfZ5_1(.dout(w_dff_A_07gJrxt32_1),.din(w_dff_A_7lNkLDfZ5_1),.clk(gclk));
	jdff dff_A_qjUNg49A8_1(.dout(w_dff_A_7lNkLDfZ5_1),.din(w_dff_A_qjUNg49A8_1),.clk(gclk));
	jdff dff_A_PAhiSHvw1_1(.dout(w_dff_A_qjUNg49A8_1),.din(w_dff_A_PAhiSHvw1_1),.clk(gclk));
	jdff dff_A_tflyMCkZ3_1(.dout(w_dff_A_PAhiSHvw1_1),.din(w_dff_A_tflyMCkZ3_1),.clk(gclk));
	jdff dff_A_cLm3788F5_1(.dout(w_dff_A_tflyMCkZ3_1),.din(w_dff_A_cLm3788F5_1),.clk(gclk));
	jdff dff_A_XA3SDY189_2(.dout(w_n843_1[2]),.din(w_dff_A_XA3SDY189_2),.clk(gclk));
	jdff dff_A_d5uhTrnv5_2(.dout(w_dff_A_XA3SDY189_2),.din(w_dff_A_d5uhTrnv5_2),.clk(gclk));
	jdff dff_A_PdeTCBKx7_2(.dout(w_dff_A_d5uhTrnv5_2),.din(w_dff_A_PdeTCBKx7_2),.clk(gclk));
	jdff dff_A_n41sYB646_2(.dout(w_dff_A_PdeTCBKx7_2),.din(w_dff_A_n41sYB646_2),.clk(gclk));
	jdff dff_A_9Paqwd7y9_2(.dout(w_dff_A_n41sYB646_2),.din(w_dff_A_9Paqwd7y9_2),.clk(gclk));
	jdff dff_A_YCzmOSG41_2(.dout(w_dff_A_9Paqwd7y9_2),.din(w_dff_A_YCzmOSG41_2),.clk(gclk));
	jdff dff_A_GExw5Bi55_2(.dout(w_dff_A_YCzmOSG41_2),.din(w_dff_A_GExw5Bi55_2),.clk(gclk));
	jdff dff_A_IGyNVtjA3_2(.dout(w_dff_A_GExw5Bi55_2),.din(w_dff_A_IGyNVtjA3_2),.clk(gclk));
	jdff dff_A_KVtIpd1a3_2(.dout(w_dff_A_IGyNVtjA3_2),.din(w_dff_A_KVtIpd1a3_2),.clk(gclk));
	jdff dff_A_e0Ih2LcX7_2(.dout(w_dff_A_KVtIpd1a3_2),.din(w_dff_A_e0Ih2LcX7_2),.clk(gclk));
	jdff dff_A_zKvsHlYu4_1(.dout(w_n843_0[1]),.din(w_dff_A_zKvsHlYu4_1),.clk(gclk));
	jdff dff_A_odlVhcBS1_1(.dout(w_dff_A_zKvsHlYu4_1),.din(w_dff_A_odlVhcBS1_1),.clk(gclk));
	jdff dff_A_0sGSeRAR2_1(.dout(w_dff_A_odlVhcBS1_1),.din(w_dff_A_0sGSeRAR2_1),.clk(gclk));
	jdff dff_A_VlmWAUTu7_1(.dout(w_dff_A_0sGSeRAR2_1),.din(w_dff_A_VlmWAUTu7_1),.clk(gclk));
	jdff dff_A_wTZE1LMp4_1(.dout(w_dff_A_VlmWAUTu7_1),.din(w_dff_A_wTZE1LMp4_1),.clk(gclk));
	jdff dff_A_jMtItFaU1_1(.dout(w_dff_A_wTZE1LMp4_1),.din(w_dff_A_jMtItFaU1_1),.clk(gclk));
	jdff dff_A_7r37JUvU9_1(.dout(w_dff_A_jMtItFaU1_1),.din(w_dff_A_7r37JUvU9_1),.clk(gclk));
	jdff dff_A_PKjuOhSd0_1(.dout(w_dff_A_7r37JUvU9_1),.din(w_dff_A_PKjuOhSd0_1),.clk(gclk));
	jdff dff_A_IaLfFmXh7_1(.dout(w_dff_A_PKjuOhSd0_1),.din(w_dff_A_IaLfFmXh7_1),.clk(gclk));
	jdff dff_A_47JVa2709_1(.dout(w_dff_A_IaLfFmXh7_1),.din(w_dff_A_47JVa2709_1),.clk(gclk));
	jdff dff_A_EW7Rn3p67_1(.dout(w_dff_A_47JVa2709_1),.din(w_dff_A_EW7Rn3p67_1),.clk(gclk));
	jdff dff_A_bYMz636x6_2(.dout(w_n843_0[2]),.din(w_dff_A_bYMz636x6_2),.clk(gclk));
	jdff dff_B_wp8dM40r5_3(.din(n843),.dout(w_dff_B_wp8dM40r5_3),.clk(gclk));
	jdff dff_B_tuhr30Vj1_3(.din(w_dff_B_wp8dM40r5_3),.dout(w_dff_B_tuhr30Vj1_3),.clk(gclk));
	jdff dff_B_J8rV2HTe9_3(.din(w_dff_B_tuhr30Vj1_3),.dout(w_dff_B_J8rV2HTe9_3),.clk(gclk));
	jdff dff_B_rVkRGztn0_3(.din(w_dff_B_J8rV2HTe9_3),.dout(w_dff_B_rVkRGztn0_3),.clk(gclk));
	jdff dff_B_i0e3EPfR9_3(.din(w_dff_B_rVkRGztn0_3),.dout(w_dff_B_i0e3EPfR9_3),.clk(gclk));
	jdff dff_B_Yt0cDv956_3(.din(w_dff_B_i0e3EPfR9_3),.dout(w_dff_B_Yt0cDv956_3),.clk(gclk));
	jdff dff_A_6al98zBo1_1(.dout(w_n840_1[1]),.din(w_dff_A_6al98zBo1_1),.clk(gclk));
	jdff dff_A_KznqRwtA5_1(.dout(w_dff_A_6al98zBo1_1),.din(w_dff_A_KznqRwtA5_1),.clk(gclk));
	jdff dff_A_iSVqMZcw6_1(.dout(w_dff_A_KznqRwtA5_1),.din(w_dff_A_iSVqMZcw6_1),.clk(gclk));
	jdff dff_A_G4snWQlh7_1(.dout(w_dff_A_iSVqMZcw6_1),.din(w_dff_A_G4snWQlh7_1),.clk(gclk));
	jdff dff_A_Hd6fwTqp3_1(.dout(w_dff_A_G4snWQlh7_1),.din(w_dff_A_Hd6fwTqp3_1),.clk(gclk));
	jdff dff_A_d5fkMHs96_1(.dout(w_dff_A_Hd6fwTqp3_1),.din(w_dff_A_d5fkMHs96_1),.clk(gclk));
	jdff dff_A_UvbRpELu2_1(.dout(w_dff_A_d5fkMHs96_1),.din(w_dff_A_UvbRpELu2_1),.clk(gclk));
	jdff dff_A_woVgbpwc3_1(.dout(w_dff_A_UvbRpELu2_1),.din(w_dff_A_woVgbpwc3_1),.clk(gclk));
	jdff dff_A_yuZPb1Ar7_1(.dout(w_dff_A_woVgbpwc3_1),.din(w_dff_A_yuZPb1Ar7_1),.clk(gclk));
	jdff dff_A_jJNAynl08_1(.dout(w_dff_A_yuZPb1Ar7_1),.din(w_dff_A_jJNAynl08_1),.clk(gclk));
	jdff dff_A_j9d07eNU4_1(.dout(w_dff_A_jJNAynl08_1),.din(w_dff_A_j9d07eNU4_1),.clk(gclk));
	jdff dff_A_M0bkpkk80_1(.dout(w_dff_A_j9d07eNU4_1),.din(w_dff_A_M0bkpkk80_1),.clk(gclk));
	jdff dff_A_1AGjTaxK9_1(.dout(w_dff_A_M0bkpkk80_1),.din(w_dff_A_1AGjTaxK9_1),.clk(gclk));
	jdff dff_A_XrgxLxLA5_1(.dout(w_dff_A_1AGjTaxK9_1),.din(w_dff_A_XrgxLxLA5_1),.clk(gclk));
	jdff dff_A_YJYuMKOa9_2(.dout(w_n840_1[2]),.din(w_dff_A_YJYuMKOa9_2),.clk(gclk));
	jdff dff_A_USTdVEhM2_2(.dout(w_dff_A_YJYuMKOa9_2),.din(w_dff_A_USTdVEhM2_2),.clk(gclk));
	jdff dff_A_NZQwyrq54_2(.dout(w_dff_A_USTdVEhM2_2),.din(w_dff_A_NZQwyrq54_2),.clk(gclk));
	jdff dff_A_t7TaXIc05_2(.dout(w_dff_A_NZQwyrq54_2),.din(w_dff_A_t7TaXIc05_2),.clk(gclk));
	jdff dff_A_MGSQUssF7_2(.dout(w_dff_A_t7TaXIc05_2),.din(w_dff_A_MGSQUssF7_2),.clk(gclk));
	jdff dff_A_uYJht2rJ8_2(.dout(w_dff_A_MGSQUssF7_2),.din(w_dff_A_uYJht2rJ8_2),.clk(gclk));
	jdff dff_A_qPHr3S106_2(.dout(w_dff_A_uYJht2rJ8_2),.din(w_dff_A_qPHr3S106_2),.clk(gclk));
	jdff dff_A_ej6mg8YW9_2(.dout(w_dff_A_qPHr3S106_2),.din(w_dff_A_ej6mg8YW9_2),.clk(gclk));
	jdff dff_A_HxmgycGO8_2(.dout(w_dff_A_ej6mg8YW9_2),.din(w_dff_A_HxmgycGO8_2),.clk(gclk));
	jdff dff_A_CkR3Lkis6_2(.dout(w_dff_A_HxmgycGO8_2),.din(w_dff_A_CkR3Lkis6_2),.clk(gclk));
	jdff dff_A_CY8HBJaz8_1(.dout(w_n840_0[1]),.din(w_dff_A_CY8HBJaz8_1),.clk(gclk));
	jdff dff_A_gqvYkV7F0_1(.dout(w_dff_A_CY8HBJaz8_1),.din(w_dff_A_gqvYkV7F0_1),.clk(gclk));
	jdff dff_A_vhFkP5jC4_1(.dout(w_dff_A_gqvYkV7F0_1),.din(w_dff_A_vhFkP5jC4_1),.clk(gclk));
	jdff dff_A_ACkO4bKS0_1(.dout(w_dff_A_vhFkP5jC4_1),.din(w_dff_A_ACkO4bKS0_1),.clk(gclk));
	jdff dff_A_0Be0J8de3_1(.dout(w_dff_A_ACkO4bKS0_1),.din(w_dff_A_0Be0J8de3_1),.clk(gclk));
	jdff dff_A_gGllZOSn2_1(.dout(w_dff_A_0Be0J8de3_1),.din(w_dff_A_gGllZOSn2_1),.clk(gclk));
	jdff dff_A_yqQWdsBy9_1(.dout(w_dff_A_gGllZOSn2_1),.din(w_dff_A_yqQWdsBy9_1),.clk(gclk));
	jdff dff_A_iPOZRX7i5_1(.dout(w_dff_A_yqQWdsBy9_1),.din(w_dff_A_iPOZRX7i5_1),.clk(gclk));
	jdff dff_A_fdth1E2X9_1(.dout(w_dff_A_iPOZRX7i5_1),.din(w_dff_A_fdth1E2X9_1),.clk(gclk));
	jdff dff_A_QyQBBsOP3_1(.dout(w_dff_A_fdth1E2X9_1),.din(w_dff_A_QyQBBsOP3_1),.clk(gclk));
	jdff dff_A_UvlIyvVv4_1(.dout(w_dff_A_QyQBBsOP3_1),.din(w_dff_A_UvlIyvVv4_1),.clk(gclk));
	jdff dff_A_pdKeiF792_2(.dout(w_n840_0[2]),.din(w_dff_A_pdKeiF792_2),.clk(gclk));
	jdff dff_A_yd5hhSny7_2(.dout(w_dff_A_pdKeiF792_2),.din(w_dff_A_yd5hhSny7_2),.clk(gclk));
	jdff dff_A_7W3Zxmuo6_2(.dout(w_dff_A_yd5hhSny7_2),.din(w_dff_A_7W3Zxmuo6_2),.clk(gclk));
	jdff dff_A_r4VlKp9Y2_2(.dout(w_dff_A_7W3Zxmuo6_2),.din(w_dff_A_r4VlKp9Y2_2),.clk(gclk));
	jdff dff_B_EUSU9yvi1_3(.din(n840),.dout(w_dff_B_EUSU9yvi1_3),.clk(gclk));
	jdff dff_B_7oV083Ax8_3(.din(w_dff_B_EUSU9yvi1_3),.dout(w_dff_B_7oV083Ax8_3),.clk(gclk));
	jdff dff_B_fEauzMyq9_3(.din(w_dff_B_7oV083Ax8_3),.dout(w_dff_B_fEauzMyq9_3),.clk(gclk));
	jdff dff_B_ZTw2ET2C5_3(.din(w_dff_B_fEauzMyq9_3),.dout(w_dff_B_ZTw2ET2C5_3),.clk(gclk));
	jdff dff_B_dyjCc6uR2_3(.din(w_dff_B_ZTw2ET2C5_3),.dout(w_dff_B_dyjCc6uR2_3),.clk(gclk));
	jdff dff_B_x1X5DVsv4_3(.din(w_dff_B_dyjCc6uR2_3),.dout(w_dff_B_x1X5DVsv4_3),.clk(gclk));
	jdff dff_B_o0TO8GKR4_3(.din(w_dff_B_x1X5DVsv4_3),.dout(w_dff_B_o0TO8GKR4_3),.clk(gclk));
	jdff dff_A_cq0xHiKF9_1(.dout(w_G4090_0[1]),.din(w_dff_A_cq0xHiKF9_1),.clk(gclk));
	jdff dff_A_KdvOQBlZ5_2(.dout(w_G4089_0[2]),.din(w_dff_A_KdvOQBlZ5_2),.clk(gclk));
	jdff dff_B_NR8kUKjf6_1(.din(n1626),.dout(w_dff_B_NR8kUKjf6_1),.clk(gclk));
	jdff dff_B_WhQnq5sJ4_0(.din(n1637),.dout(w_dff_B_WhQnq5sJ4_0),.clk(gclk));
	jdff dff_B_KZ5ZqctT0_0(.din(w_dff_B_WhQnq5sJ4_0),.dout(w_dff_B_KZ5ZqctT0_0),.clk(gclk));
	jdff dff_B_SFZ16NJx3_0(.din(w_dff_B_KZ5ZqctT0_0),.dout(w_dff_B_SFZ16NJx3_0),.clk(gclk));
	jdff dff_B_gtxJtZeV9_0(.din(w_dff_B_SFZ16NJx3_0),.dout(w_dff_B_gtxJtZeV9_0),.clk(gclk));
	jdff dff_B_O3ZZ2U2y0_0(.din(w_dff_B_gtxJtZeV9_0),.dout(w_dff_B_O3ZZ2U2y0_0),.clk(gclk));
	jdff dff_B_luJSb5d74_0(.din(w_dff_B_O3ZZ2U2y0_0),.dout(w_dff_B_luJSb5d74_0),.clk(gclk));
	jdff dff_B_pX3fj7mK9_0(.din(w_dff_B_luJSb5d74_0),.dout(w_dff_B_pX3fj7mK9_0),.clk(gclk));
	jdff dff_B_O1SrJoJK7_0(.din(w_dff_B_pX3fj7mK9_0),.dout(w_dff_B_O1SrJoJK7_0),.clk(gclk));
	jdff dff_B_slhLsD888_0(.din(w_dff_B_O1SrJoJK7_0),.dout(w_dff_B_slhLsD888_0),.clk(gclk));
	jdff dff_B_HD260L7R7_0(.din(w_dff_B_slhLsD888_0),.dout(w_dff_B_HD260L7R7_0),.clk(gclk));
	jdff dff_B_lMkKxrOG9_0(.din(w_dff_B_HD260L7R7_0),.dout(w_dff_B_lMkKxrOG9_0),.clk(gclk));
	jdff dff_B_S8Ko5jJ31_0(.din(w_dff_B_lMkKxrOG9_0),.dout(w_dff_B_S8Ko5jJ31_0),.clk(gclk));
	jdff dff_B_JB0jJLuj6_0(.din(w_dff_B_S8Ko5jJ31_0),.dout(w_dff_B_JB0jJLuj6_0),.clk(gclk));
	jdff dff_B_AwwbHqDV9_0(.din(w_dff_B_JB0jJLuj6_0),.dout(w_dff_B_AwwbHqDV9_0),.clk(gclk));
	jdff dff_B_Iv89Bw3L1_0(.din(w_dff_B_AwwbHqDV9_0),.dout(w_dff_B_Iv89Bw3L1_0),.clk(gclk));
	jdff dff_B_qCy93SKL0_0(.din(w_dff_B_Iv89Bw3L1_0),.dout(w_dff_B_qCy93SKL0_0),.clk(gclk));
	jdff dff_B_Q8YlNiuX2_0(.din(w_dff_B_qCy93SKL0_0),.dout(w_dff_B_Q8YlNiuX2_0),.clk(gclk));
	jdff dff_B_N3bhsw929_0(.din(w_dff_B_Q8YlNiuX2_0),.dout(w_dff_B_N3bhsw929_0),.clk(gclk));
	jdff dff_B_Y2zKwqgq8_1(.din(n1633),.dout(w_dff_B_Y2zKwqgq8_1),.clk(gclk));
	jdff dff_B_OaTQ7bdM2_1(.din(n1627),.dout(w_dff_B_OaTQ7bdM2_1),.clk(gclk));
	jdff dff_B_gTnF0hhZ1_1(.din(w_dff_B_OaTQ7bdM2_1),.dout(w_dff_B_gTnF0hhZ1_1),.clk(gclk));
	jdff dff_B_XmbERwBF2_1(.din(w_dff_B_gTnF0hhZ1_1),.dout(w_dff_B_XmbERwBF2_1),.clk(gclk));
	jdff dff_B_Yn4fCEHl0_1(.din(w_dff_B_XmbERwBF2_1),.dout(w_dff_B_Yn4fCEHl0_1),.clk(gclk));
	jdff dff_B_x24QcgoJ7_1(.din(w_dff_B_Yn4fCEHl0_1),.dout(w_dff_B_x24QcgoJ7_1),.clk(gclk));
	jdff dff_B_om6QDEp21_1(.din(w_dff_B_x24QcgoJ7_1),.dout(w_dff_B_om6QDEp21_1),.clk(gclk));
	jdff dff_B_8CjxlMrm4_1(.din(w_dff_B_om6QDEp21_1),.dout(w_dff_B_8CjxlMrm4_1),.clk(gclk));
	jdff dff_B_GJRJsd8C2_1(.din(w_dff_B_8CjxlMrm4_1),.dout(w_dff_B_GJRJsd8C2_1),.clk(gclk));
	jdff dff_B_MQ5E8njR0_1(.din(w_dff_B_GJRJsd8C2_1),.dout(w_dff_B_MQ5E8njR0_1),.clk(gclk));
	jdff dff_B_cMWd1y872_1(.din(w_dff_B_MQ5E8njR0_1),.dout(w_dff_B_cMWd1y872_1),.clk(gclk));
	jdff dff_B_UChMHbeZ7_1(.din(w_dff_B_cMWd1y872_1),.dout(w_dff_B_UChMHbeZ7_1),.clk(gclk));
	jdff dff_B_e3dfbYO75_1(.din(w_dff_B_UChMHbeZ7_1),.dout(w_dff_B_e3dfbYO75_1),.clk(gclk));
	jdff dff_B_7eugVS2t5_1(.din(w_dff_B_e3dfbYO75_1),.dout(w_dff_B_7eugVS2t5_1),.clk(gclk));
	jdff dff_B_arJRmmGp6_1(.din(w_dff_B_7eugVS2t5_1),.dout(w_dff_B_arJRmmGp6_1),.clk(gclk));
	jdff dff_B_KpvqEHQ73_1(.din(w_dff_B_arJRmmGp6_1),.dout(w_dff_B_KpvqEHQ73_1),.clk(gclk));
	jdff dff_B_cPfKSmq26_1(.din(w_dff_B_KpvqEHQ73_1),.dout(w_dff_B_cPfKSmq26_1),.clk(gclk));
	jdff dff_B_h1YwIRpF1_1(.din(w_dff_B_cPfKSmq26_1),.dout(w_dff_B_h1YwIRpF1_1),.clk(gclk));
	jdff dff_B_ser3Szfs2_1(.din(w_dff_B_h1YwIRpF1_1),.dout(w_dff_B_ser3Szfs2_1),.clk(gclk));
	jdff dff_B_6DkHFI564_1(.din(w_dff_B_ser3Szfs2_1),.dout(w_dff_B_6DkHFI564_1),.clk(gclk));
	jdff dff_A_b2HyIx4X7_0(.dout(w_n988_1[0]),.din(w_dff_A_b2HyIx4X7_0),.clk(gclk));
	jdff dff_A_l1KzmhGt6_0(.dout(w_dff_A_b2HyIx4X7_0),.din(w_dff_A_l1KzmhGt6_0),.clk(gclk));
	jdff dff_A_bfPMpFec3_0(.dout(w_dff_A_l1KzmhGt6_0),.din(w_dff_A_bfPMpFec3_0),.clk(gclk));
	jdff dff_A_7wTMAY2a4_0(.dout(w_dff_A_bfPMpFec3_0),.din(w_dff_A_7wTMAY2a4_0),.clk(gclk));
	jdff dff_A_5zgI1F9C6_0(.dout(w_dff_A_7wTMAY2a4_0),.din(w_dff_A_5zgI1F9C6_0),.clk(gclk));
	jdff dff_A_9hkTMXuv6_0(.dout(w_dff_A_5zgI1F9C6_0),.din(w_dff_A_9hkTMXuv6_0),.clk(gclk));
	jdff dff_A_6nWnQ8WQ2_2(.dout(w_n988_1[2]),.din(w_dff_A_6nWnQ8WQ2_2),.clk(gclk));
	jdff dff_A_JIqhdBQF0_2(.dout(w_dff_A_6nWnQ8WQ2_2),.din(w_dff_A_JIqhdBQF0_2),.clk(gclk));
	jdff dff_A_aOpzuHuB4_2(.dout(w_dff_A_JIqhdBQF0_2),.din(w_dff_A_aOpzuHuB4_2),.clk(gclk));
	jdff dff_A_hP5MfCMH7_2(.dout(w_dff_A_aOpzuHuB4_2),.din(w_dff_A_hP5MfCMH7_2),.clk(gclk));
	jdff dff_A_iPooV75A1_2(.dout(w_dff_A_hP5MfCMH7_2),.din(w_dff_A_iPooV75A1_2),.clk(gclk));
	jdff dff_A_CBESp0Zv8_2(.dout(w_dff_A_iPooV75A1_2),.din(w_dff_A_CBESp0Zv8_2),.clk(gclk));
	jdff dff_A_lRH3KiF76_2(.dout(w_dff_A_CBESp0Zv8_2),.din(w_dff_A_lRH3KiF76_2),.clk(gclk));
	jdff dff_A_4orQVfpH8_2(.dout(w_dff_A_lRH3KiF76_2),.din(w_dff_A_4orQVfpH8_2),.clk(gclk));
	jdff dff_A_FuUeHiEx8_2(.dout(w_dff_A_4orQVfpH8_2),.din(w_dff_A_FuUeHiEx8_2),.clk(gclk));
	jdff dff_A_79McScpt7_2(.dout(w_dff_A_FuUeHiEx8_2),.din(w_dff_A_79McScpt7_2),.clk(gclk));
	jdff dff_A_XBJgKqPn5_2(.dout(w_dff_A_79McScpt7_2),.din(w_dff_A_XBJgKqPn5_2),.clk(gclk));
	jdff dff_A_zowD7kYJ3_2(.dout(w_dff_A_XBJgKqPn5_2),.din(w_dff_A_zowD7kYJ3_2),.clk(gclk));
	jdff dff_A_hlS3TIUR2_2(.dout(w_dff_A_zowD7kYJ3_2),.din(w_dff_A_hlS3TIUR2_2),.clk(gclk));
	jdff dff_A_y1aAJKTm9_2(.dout(w_dff_A_hlS3TIUR2_2),.din(w_dff_A_y1aAJKTm9_2),.clk(gclk));
	jdff dff_A_DUCTwtbJ8_2(.dout(w_dff_A_y1aAJKTm9_2),.din(w_dff_A_DUCTwtbJ8_2),.clk(gclk));
	jdff dff_A_WSAtZebq9_2(.dout(w_dff_A_DUCTwtbJ8_2),.din(w_dff_A_WSAtZebq9_2),.clk(gclk));
	jdff dff_A_VE9dbpK31_2(.dout(w_dff_A_WSAtZebq9_2),.din(w_dff_A_VE9dbpK31_2),.clk(gclk));
	jdff dff_A_05E4x0Ju7_2(.dout(w_dff_A_VE9dbpK31_2),.din(w_dff_A_05E4x0Ju7_2),.clk(gclk));
	jdff dff_A_BDhw5niW5_1(.dout(w_n988_0[1]),.din(w_dff_A_BDhw5niW5_1),.clk(gclk));
	jdff dff_A_4EjTNEXI4_1(.dout(w_dff_A_BDhw5niW5_1),.din(w_dff_A_4EjTNEXI4_1),.clk(gclk));
	jdff dff_A_nVPydCPI0_1(.dout(w_dff_A_4EjTNEXI4_1),.din(w_dff_A_nVPydCPI0_1),.clk(gclk));
	jdff dff_A_b7mgi8hu3_1(.dout(w_dff_A_nVPydCPI0_1),.din(w_dff_A_b7mgi8hu3_1),.clk(gclk));
	jdff dff_A_Su36576Z0_1(.dout(w_dff_A_b7mgi8hu3_1),.din(w_dff_A_Su36576Z0_1),.clk(gclk));
	jdff dff_A_7z0UyjIh7_1(.dout(w_dff_A_Su36576Z0_1),.din(w_dff_A_7z0UyjIh7_1),.clk(gclk));
	jdff dff_A_BVgrDzBA1_1(.dout(w_dff_A_7z0UyjIh7_1),.din(w_dff_A_BVgrDzBA1_1),.clk(gclk));
	jdff dff_A_xQGBG9ho0_1(.dout(w_dff_A_BVgrDzBA1_1),.din(w_dff_A_xQGBG9ho0_1),.clk(gclk));
	jdff dff_A_Dv96yhB60_1(.dout(w_dff_A_xQGBG9ho0_1),.din(w_dff_A_Dv96yhB60_1),.clk(gclk));
	jdff dff_A_2n6c2x286_1(.dout(w_dff_A_Dv96yhB60_1),.din(w_dff_A_2n6c2x286_1),.clk(gclk));
	jdff dff_A_801GmJsc4_1(.dout(w_dff_A_2n6c2x286_1),.din(w_dff_A_801GmJsc4_1),.clk(gclk));
	jdff dff_A_DxVimEqQ5_1(.dout(w_dff_A_801GmJsc4_1),.din(w_dff_A_DxVimEqQ5_1),.clk(gclk));
	jdff dff_A_Vzv5zBV12_1(.dout(w_dff_A_DxVimEqQ5_1),.din(w_dff_A_Vzv5zBV12_1),.clk(gclk));
	jdff dff_A_UeDiK38c1_1(.dout(w_dff_A_Vzv5zBV12_1),.din(w_dff_A_UeDiK38c1_1),.clk(gclk));
	jdff dff_A_uA8EBtVp2_1(.dout(w_dff_A_UeDiK38c1_1),.din(w_dff_A_uA8EBtVp2_1),.clk(gclk));
	jdff dff_A_E0FEgWNI2_1(.dout(w_dff_A_uA8EBtVp2_1),.din(w_dff_A_E0FEgWNI2_1),.clk(gclk));
	jdff dff_A_MOLNIlYw8_2(.dout(w_n988_0[2]),.din(w_dff_A_MOLNIlYw8_2),.clk(gclk));
	jdff dff_A_tZT1IM5d1_2(.dout(w_dff_A_MOLNIlYw8_2),.din(w_dff_A_tZT1IM5d1_2),.clk(gclk));
	jdff dff_A_32gvR2nv3_2(.dout(w_dff_A_tZT1IM5d1_2),.din(w_dff_A_32gvR2nv3_2),.clk(gclk));
	jdff dff_A_hMyA9hSm9_2(.dout(w_dff_A_32gvR2nv3_2),.din(w_dff_A_hMyA9hSm9_2),.clk(gclk));
	jdff dff_A_HQlyKJhr0_2(.dout(w_dff_A_hMyA9hSm9_2),.din(w_dff_A_HQlyKJhr0_2),.clk(gclk));
	jdff dff_A_g576yzHV3_2(.dout(w_dff_A_HQlyKJhr0_2),.din(w_dff_A_g576yzHV3_2),.clk(gclk));
	jdff dff_A_TM4UFaXR3_2(.dout(w_dff_A_g576yzHV3_2),.din(w_dff_A_TM4UFaXR3_2),.clk(gclk));
	jdff dff_B_uX6fm1yp9_1(.din(n1625),.dout(w_dff_B_uX6fm1yp9_1),.clk(gclk));
	jdff dff_B_l55ac3zf1_1(.din(w_dff_B_uX6fm1yp9_1),.dout(w_dff_B_l55ac3zf1_1),.clk(gclk));
	jdff dff_B_k85U420F9_1(.din(w_dff_B_l55ac3zf1_1),.dout(w_dff_B_k85U420F9_1),.clk(gclk));
	jdff dff_B_dOQvKVCU2_1(.din(w_dff_B_k85U420F9_1),.dout(w_dff_B_dOQvKVCU2_1),.clk(gclk));
	jdff dff_B_Z5MpaPjb9_1(.din(w_dff_B_dOQvKVCU2_1),.dout(w_dff_B_Z5MpaPjb9_1),.clk(gclk));
	jdff dff_B_eL2i8GMT5_1(.din(w_dff_B_Z5MpaPjb9_1),.dout(w_dff_B_eL2i8GMT5_1),.clk(gclk));
	jdff dff_B_BKYNshWs5_1(.din(w_dff_B_eL2i8GMT5_1),.dout(w_dff_B_BKYNshWs5_1),.clk(gclk));
	jdff dff_B_LdmblYQH9_1(.din(w_dff_B_BKYNshWs5_1),.dout(w_dff_B_LdmblYQH9_1),.clk(gclk));
	jdff dff_B_gqxdiTH57_1(.din(w_dff_B_LdmblYQH9_1),.dout(w_dff_B_gqxdiTH57_1),.clk(gclk));
	jdff dff_B_hF5jwuWr3_1(.din(w_dff_B_gqxdiTH57_1),.dout(w_dff_B_hF5jwuWr3_1),.clk(gclk));
	jdff dff_B_S2gX7Guz7_1(.din(w_dff_B_hF5jwuWr3_1),.dout(w_dff_B_S2gX7Guz7_1),.clk(gclk));
	jdff dff_B_OJRHRCdZ1_1(.din(w_dff_B_S2gX7Guz7_1),.dout(w_dff_B_OJRHRCdZ1_1),.clk(gclk));
	jdff dff_B_3YWEuYjq6_1(.din(w_dff_B_OJRHRCdZ1_1),.dout(w_dff_B_3YWEuYjq6_1),.clk(gclk));
	jdff dff_B_JdvvhKqA7_1(.din(w_dff_B_3YWEuYjq6_1),.dout(w_dff_B_JdvvhKqA7_1),.clk(gclk));
	jdff dff_B_JDlRFUv94_1(.din(w_dff_B_JdvvhKqA7_1),.dout(w_dff_B_JDlRFUv94_1),.clk(gclk));
	jdff dff_B_8dg9T0ZE7_1(.din(w_dff_B_JDlRFUv94_1),.dout(w_dff_B_8dg9T0ZE7_1),.clk(gclk));
	jdff dff_B_bjbOQTVL5_1(.din(w_dff_B_8dg9T0ZE7_1),.dout(w_dff_B_bjbOQTVL5_1),.clk(gclk));
	jdff dff_B_swLcmRVK0_1(.din(w_dff_B_bjbOQTVL5_1),.dout(w_dff_B_swLcmRVK0_1),.clk(gclk));
	jdff dff_B_yj6s74DZ0_1(.din(w_dff_B_swLcmRVK0_1),.dout(w_dff_B_yj6s74DZ0_1),.clk(gclk));
	jdff dff_A_3aoepQuQ6_0(.dout(w_n985_1[0]),.din(w_dff_A_3aoepQuQ6_0),.clk(gclk));
	jdff dff_A_MaiT6gHE5_0(.dout(w_dff_A_3aoepQuQ6_0),.din(w_dff_A_MaiT6gHE5_0),.clk(gclk));
	jdff dff_A_eHoJOWCv1_0(.dout(w_dff_A_MaiT6gHE5_0),.din(w_dff_A_eHoJOWCv1_0),.clk(gclk));
	jdff dff_A_vT4XYbAy8_0(.dout(w_dff_A_eHoJOWCv1_0),.din(w_dff_A_vT4XYbAy8_0),.clk(gclk));
	jdff dff_A_rN21rD7D0_0(.dout(w_dff_A_vT4XYbAy8_0),.din(w_dff_A_rN21rD7D0_0),.clk(gclk));
	jdff dff_A_BvsbVYay0_0(.dout(w_dff_A_rN21rD7D0_0),.din(w_dff_A_BvsbVYay0_0),.clk(gclk));
	jdff dff_A_mIXe8xdZ8_0(.dout(w_dff_A_BvsbVYay0_0),.din(w_dff_A_mIXe8xdZ8_0),.clk(gclk));
	jdff dff_A_2gLfNMss4_2(.dout(w_n985_1[2]),.din(w_dff_A_2gLfNMss4_2),.clk(gclk));
	jdff dff_A_qxkoWRMr5_2(.dout(w_dff_A_2gLfNMss4_2),.din(w_dff_A_qxkoWRMr5_2),.clk(gclk));
	jdff dff_A_kF9n7W9F8_2(.dout(w_dff_A_qxkoWRMr5_2),.din(w_dff_A_kF9n7W9F8_2),.clk(gclk));
	jdff dff_A_XGsl4uvd2_2(.dout(w_dff_A_kF9n7W9F8_2),.din(w_dff_A_XGsl4uvd2_2),.clk(gclk));
	jdff dff_A_C94puwKL4_2(.dout(w_dff_A_XGsl4uvd2_2),.din(w_dff_A_C94puwKL4_2),.clk(gclk));
	jdff dff_A_WGqOagTa3_2(.dout(w_dff_A_C94puwKL4_2),.din(w_dff_A_WGqOagTa3_2),.clk(gclk));
	jdff dff_A_92Z6vrxQ4_2(.dout(w_dff_A_WGqOagTa3_2),.din(w_dff_A_92Z6vrxQ4_2),.clk(gclk));
	jdff dff_A_h28ilWMj8_2(.dout(w_dff_A_92Z6vrxQ4_2),.din(w_dff_A_h28ilWMj8_2),.clk(gclk));
	jdff dff_A_gXW1EJ6i6_2(.dout(w_dff_A_h28ilWMj8_2),.din(w_dff_A_gXW1EJ6i6_2),.clk(gclk));
	jdff dff_A_Zled6e9F0_2(.dout(w_dff_A_gXW1EJ6i6_2),.din(w_dff_A_Zled6e9F0_2),.clk(gclk));
	jdff dff_A_mm6LFWM94_2(.dout(w_dff_A_Zled6e9F0_2),.din(w_dff_A_mm6LFWM94_2),.clk(gclk));
	jdff dff_A_E9NYpw2J6_2(.dout(w_dff_A_mm6LFWM94_2),.din(w_dff_A_E9NYpw2J6_2),.clk(gclk));
	jdff dff_A_HWRYfVeP3_2(.dout(w_dff_A_E9NYpw2J6_2),.din(w_dff_A_HWRYfVeP3_2),.clk(gclk));
	jdff dff_A_2AYdM0B88_2(.dout(w_dff_A_HWRYfVeP3_2),.din(w_dff_A_2AYdM0B88_2),.clk(gclk));
	jdff dff_A_9ces2Q0F2_2(.dout(w_dff_A_2AYdM0B88_2),.din(w_dff_A_9ces2Q0F2_2),.clk(gclk));
	jdff dff_A_8gVRgFJw9_2(.dout(w_dff_A_9ces2Q0F2_2),.din(w_dff_A_8gVRgFJw9_2),.clk(gclk));
	jdff dff_A_saL2bOkE4_2(.dout(w_dff_A_8gVRgFJw9_2),.din(w_dff_A_saL2bOkE4_2),.clk(gclk));
	jdff dff_A_IqvSwh3X0_2(.dout(w_dff_A_saL2bOkE4_2),.din(w_dff_A_IqvSwh3X0_2),.clk(gclk));
	jdff dff_A_KvJpBKkq7_2(.dout(w_dff_A_IqvSwh3X0_2),.din(w_dff_A_KvJpBKkq7_2),.clk(gclk));
	jdff dff_A_pQDVWf7y9_1(.dout(w_n985_0[1]),.din(w_dff_A_pQDVWf7y9_1),.clk(gclk));
	jdff dff_A_yII1lfT33_1(.dout(w_dff_A_pQDVWf7y9_1),.din(w_dff_A_yII1lfT33_1),.clk(gclk));
	jdff dff_A_niGQDmtC9_1(.dout(w_dff_A_yII1lfT33_1),.din(w_dff_A_niGQDmtC9_1),.clk(gclk));
	jdff dff_A_bAhZVycI6_1(.dout(w_dff_A_niGQDmtC9_1),.din(w_dff_A_bAhZVycI6_1),.clk(gclk));
	jdff dff_A_bCsgbZr89_1(.dout(w_dff_A_bAhZVycI6_1),.din(w_dff_A_bCsgbZr89_1),.clk(gclk));
	jdff dff_A_9VZLBhhS3_1(.dout(w_dff_A_bCsgbZr89_1),.din(w_dff_A_9VZLBhhS3_1),.clk(gclk));
	jdff dff_A_t7GbPZJz4_1(.dout(w_dff_A_9VZLBhhS3_1),.din(w_dff_A_t7GbPZJz4_1),.clk(gclk));
	jdff dff_A_r84M9yzz2_1(.dout(w_dff_A_t7GbPZJz4_1),.din(w_dff_A_r84M9yzz2_1),.clk(gclk));
	jdff dff_A_HKHY9Xyz9_1(.dout(w_dff_A_r84M9yzz2_1),.din(w_dff_A_HKHY9Xyz9_1),.clk(gclk));
	jdff dff_A_2eIHalnS0_1(.dout(w_dff_A_HKHY9Xyz9_1),.din(w_dff_A_2eIHalnS0_1),.clk(gclk));
	jdff dff_A_GKxW2dKs6_1(.dout(w_dff_A_2eIHalnS0_1),.din(w_dff_A_GKxW2dKs6_1),.clk(gclk));
	jdff dff_A_mlGq3BEF8_1(.dout(w_dff_A_GKxW2dKs6_1),.din(w_dff_A_mlGq3BEF8_1),.clk(gclk));
	jdff dff_A_e6EBoZ4o1_1(.dout(w_dff_A_mlGq3BEF8_1),.din(w_dff_A_e6EBoZ4o1_1),.clk(gclk));
	jdff dff_A_Qyllv4ZZ3_1(.dout(w_dff_A_e6EBoZ4o1_1),.din(w_dff_A_Qyllv4ZZ3_1),.clk(gclk));
	jdff dff_A_UTIaLtJJ8_1(.dout(w_dff_A_Qyllv4ZZ3_1),.din(w_dff_A_UTIaLtJJ8_1),.clk(gclk));
	jdff dff_A_OtcaZTIm7_1(.dout(w_dff_A_UTIaLtJJ8_1),.din(w_dff_A_OtcaZTIm7_1),.clk(gclk));
	jdff dff_A_b0r6wlAP8_1(.dout(w_dff_A_OtcaZTIm7_1),.din(w_dff_A_b0r6wlAP8_1),.clk(gclk));
	jdff dff_A_xQFUmvbJ1_2(.dout(w_n985_0[2]),.din(w_dff_A_xQFUmvbJ1_2),.clk(gclk));
	jdff dff_A_waD4hJNb6_2(.dout(w_dff_A_xQFUmvbJ1_2),.din(w_dff_A_waD4hJNb6_2),.clk(gclk));
	jdff dff_A_OI4vDBoZ9_2(.dout(w_dff_A_waD4hJNb6_2),.din(w_dff_A_OI4vDBoZ9_2),.clk(gclk));
	jdff dff_A_XWwaykSg4_2(.dout(w_dff_A_OI4vDBoZ9_2),.din(w_dff_A_XWwaykSg4_2),.clk(gclk));
	jdff dff_A_gN2WVd530_2(.dout(w_dff_A_XWwaykSg4_2),.din(w_dff_A_gN2WVd530_2),.clk(gclk));
	jdff dff_A_zj42el4G8_2(.dout(w_dff_A_gN2WVd530_2),.din(w_dff_A_zj42el4G8_2),.clk(gclk));
	jdff dff_A_vAAavfTv4_2(.dout(w_dff_A_zj42el4G8_2),.din(w_dff_A_vAAavfTv4_2),.clk(gclk));
	jdff dff_A_DSuEjwyl4_2(.dout(w_dff_A_vAAavfTv4_2),.din(w_dff_A_DSuEjwyl4_2),.clk(gclk));
	jdff dff_A_kZwk6EeY7_2(.dout(w_dff_A_DSuEjwyl4_2),.din(w_dff_A_kZwk6EeY7_2),.clk(gclk));
	jdff dff_A_YLufA5ov7_2(.dout(w_dff_A_kZwk6EeY7_2),.din(w_dff_A_YLufA5ov7_2),.clk(gclk));
	jdff dff_A_8kV4NODC1_2(.dout(w_dff_A_YLufA5ov7_2),.din(w_dff_A_8kV4NODC1_2),.clk(gclk));
	jdff dff_A_hAuu7uOo4_1(.dout(w_G1690_0[1]),.din(w_dff_A_hAuu7uOo4_1),.clk(gclk));
	jdff dff_A_4K5utaxy6_2(.dout(w_G1689_0[2]),.din(w_dff_A_4K5utaxy6_2),.clk(gclk));
	jdff dff_B_bUIEw9Ht9_1(.din(n1642),.dout(w_dff_B_bUIEw9Ht9_1),.clk(gclk));
	jdff dff_B_MFqRftBj7_0(.din(n1649),.dout(w_dff_B_MFqRftBj7_0),.clk(gclk));
	jdff dff_B_wwN2ZWMl5_0(.din(w_dff_B_MFqRftBj7_0),.dout(w_dff_B_wwN2ZWMl5_0),.clk(gclk));
	jdff dff_B_5HLcBw6a1_0(.din(w_dff_B_wwN2ZWMl5_0),.dout(w_dff_B_5HLcBw6a1_0),.clk(gclk));
	jdff dff_B_0vi24xSR5_0(.din(w_dff_B_5HLcBw6a1_0),.dout(w_dff_B_0vi24xSR5_0),.clk(gclk));
	jdff dff_B_WtlxMSEY0_0(.din(w_dff_B_0vi24xSR5_0),.dout(w_dff_B_WtlxMSEY0_0),.clk(gclk));
	jdff dff_B_HA87sxbP3_0(.din(w_dff_B_WtlxMSEY0_0),.dout(w_dff_B_HA87sxbP3_0),.clk(gclk));
	jdff dff_B_6QZC9LO09_0(.din(w_dff_B_HA87sxbP3_0),.dout(w_dff_B_6QZC9LO09_0),.clk(gclk));
	jdff dff_B_R1knWCXl8_0(.din(w_dff_B_6QZC9LO09_0),.dout(w_dff_B_R1knWCXl8_0),.clk(gclk));
	jdff dff_B_FGfREHID0_0(.din(w_dff_B_R1knWCXl8_0),.dout(w_dff_B_FGfREHID0_0),.clk(gclk));
	jdff dff_B_XkOSzIVb3_0(.din(w_dff_B_FGfREHID0_0),.dout(w_dff_B_XkOSzIVb3_0),.clk(gclk));
	jdff dff_B_7lFzwO0I2_0(.din(w_dff_B_XkOSzIVb3_0),.dout(w_dff_B_7lFzwO0I2_0),.clk(gclk));
	jdff dff_B_NTH83tE10_0(.din(w_dff_B_7lFzwO0I2_0),.dout(w_dff_B_NTH83tE10_0),.clk(gclk));
	jdff dff_B_ZFAznCmj2_0(.din(w_dff_B_NTH83tE10_0),.dout(w_dff_B_ZFAznCmj2_0),.clk(gclk));
	jdff dff_B_4BVnWiFU5_0(.din(w_dff_B_ZFAznCmj2_0),.dout(w_dff_B_4BVnWiFU5_0),.clk(gclk));
	jdff dff_B_wet4wW6b3_0(.din(w_dff_B_4BVnWiFU5_0),.dout(w_dff_B_wet4wW6b3_0),.clk(gclk));
	jdff dff_B_fxuBubNH2_0(.din(w_dff_B_wet4wW6b3_0),.dout(w_dff_B_fxuBubNH2_0),.clk(gclk));
	jdff dff_B_OiZopLEY6_0(.din(w_dff_B_fxuBubNH2_0),.dout(w_dff_B_OiZopLEY6_0),.clk(gclk));
	jdff dff_B_oAXzuI4Y3_0(.din(w_dff_B_OiZopLEY6_0),.dout(w_dff_B_oAXzuI4Y3_0),.clk(gclk));
	jdff dff_B_rptlmaIn4_1(.din(n1646),.dout(w_dff_B_rptlmaIn4_1),.clk(gclk));
	jdff dff_B_PEdQ3EmT9_2(.din(n1634),.dout(w_dff_B_PEdQ3EmT9_2),.clk(gclk));
	jdff dff_B_Ae5xATey6_2(.din(w_dff_B_PEdQ3EmT9_2),.dout(w_dff_B_Ae5xATey6_2),.clk(gclk));
	jdff dff_B_tg4sOAdy4_2(.din(n1631),.dout(w_dff_B_tg4sOAdy4_2),.clk(gclk));
	jdff dff_B_wFafgjDp1_1(.din(n1643),.dout(w_dff_B_wFafgjDp1_1),.clk(gclk));
	jdff dff_B_vJYesSgQ2_1(.din(w_dff_B_wFafgjDp1_1),.dout(w_dff_B_vJYesSgQ2_1),.clk(gclk));
	jdff dff_B_1hL04zqt9_1(.din(w_dff_B_vJYesSgQ2_1),.dout(w_dff_B_1hL04zqt9_1),.clk(gclk));
	jdff dff_B_1XAG4UB94_1(.din(w_dff_B_1hL04zqt9_1),.dout(w_dff_B_1XAG4UB94_1),.clk(gclk));
	jdff dff_B_XIBLpbuT5_1(.din(w_dff_B_1XAG4UB94_1),.dout(w_dff_B_XIBLpbuT5_1),.clk(gclk));
	jdff dff_B_7xXww1s13_1(.din(w_dff_B_XIBLpbuT5_1),.dout(w_dff_B_7xXww1s13_1),.clk(gclk));
	jdff dff_B_20GffJfk8_1(.din(w_dff_B_7xXww1s13_1),.dout(w_dff_B_20GffJfk8_1),.clk(gclk));
	jdff dff_B_kOF44eMj7_1(.din(w_dff_B_20GffJfk8_1),.dout(w_dff_B_kOF44eMj7_1),.clk(gclk));
	jdff dff_B_FcE3S7Hb0_1(.din(w_dff_B_kOF44eMj7_1),.dout(w_dff_B_FcE3S7Hb0_1),.clk(gclk));
	jdff dff_B_ohPMvGva8_1(.din(w_dff_B_FcE3S7Hb0_1),.dout(w_dff_B_ohPMvGva8_1),.clk(gclk));
	jdff dff_B_kt67avJ57_1(.din(w_dff_B_ohPMvGva8_1),.dout(w_dff_B_kt67avJ57_1),.clk(gclk));
	jdff dff_B_v4LIvFRX2_1(.din(w_dff_B_kt67avJ57_1),.dout(w_dff_B_v4LIvFRX2_1),.clk(gclk));
	jdff dff_B_IAUSHcP70_1(.din(w_dff_B_v4LIvFRX2_1),.dout(w_dff_B_IAUSHcP70_1),.clk(gclk));
	jdff dff_B_rCJXoSVM0_1(.din(w_dff_B_IAUSHcP70_1),.dout(w_dff_B_rCJXoSVM0_1),.clk(gclk));
	jdff dff_B_fI3iXvtQ8_1(.din(w_dff_B_rCJXoSVM0_1),.dout(w_dff_B_fI3iXvtQ8_1),.clk(gclk));
	jdff dff_B_DRCfWsLp8_1(.din(w_dff_B_fI3iXvtQ8_1),.dout(w_dff_B_DRCfWsLp8_1),.clk(gclk));
	jdff dff_B_0eWZonhG5_1(.din(w_dff_B_DRCfWsLp8_1),.dout(w_dff_B_0eWZonhG5_1),.clk(gclk));
	jdff dff_B_SlYcJ2tf3_1(.din(w_dff_B_0eWZonhG5_1),.dout(w_dff_B_SlYcJ2tf3_1),.clk(gclk));
	jdff dff_B_cRFX9r2w7_1(.din(w_dff_B_SlYcJ2tf3_1),.dout(w_dff_B_cRFX9r2w7_1),.clk(gclk));
	jdff dff_B_mPT6U0vQ3_0(.din(n1628),.dout(w_dff_B_mPT6U0vQ3_0),.clk(gclk));
	jdff dff_B_PxBszWCK7_0(.din(w_dff_B_mPT6U0vQ3_0),.dout(w_dff_B_PxBszWCK7_0),.clk(gclk));
	jdff dff_B_GCtCjRgK1_0(.din(w_dff_B_PxBszWCK7_0),.dout(w_dff_B_GCtCjRgK1_0),.clk(gclk));
	jdff dff_B_A9LejHtE9_0(.din(w_dff_B_GCtCjRgK1_0),.dout(w_dff_B_A9LejHtE9_0),.clk(gclk));
	jdff dff_B_qgpV7zM45_0(.din(w_dff_B_A9LejHtE9_0),.dout(w_dff_B_qgpV7zM45_0),.clk(gclk));
	jdff dff_B_zcSyOTBC1_0(.din(w_dff_B_qgpV7zM45_0),.dout(w_dff_B_zcSyOTBC1_0),.clk(gclk));
	jdff dff_B_RRbwzLUp8_0(.din(w_dff_B_zcSyOTBC1_0),.dout(w_dff_B_RRbwzLUp8_0),.clk(gclk));
	jdff dff_B_pV9SSINE3_0(.din(w_dff_B_RRbwzLUp8_0),.dout(w_dff_B_pV9SSINE3_0),.clk(gclk));
	jdff dff_B_H4xIpi0f4_0(.din(w_dff_B_pV9SSINE3_0),.dout(w_dff_B_H4xIpi0f4_0),.clk(gclk));
	jdff dff_B_n41wXQkQ7_0(.din(w_dff_B_H4xIpi0f4_0),.dout(w_dff_B_n41wXQkQ7_0),.clk(gclk));
	jdff dff_B_qB89Bdb28_0(.din(w_dff_B_n41wXQkQ7_0),.dout(w_dff_B_qB89Bdb28_0),.clk(gclk));
	jdff dff_B_sRa9pirE5_0(.din(w_dff_B_qB89Bdb28_0),.dout(w_dff_B_sRa9pirE5_0),.clk(gclk));
	jdff dff_B_cZ5Z913j9_0(.din(w_dff_B_sRa9pirE5_0),.dout(w_dff_B_cZ5Z913j9_0),.clk(gclk));
	jdff dff_B_5adj63mH4_0(.din(w_dff_B_cZ5Z913j9_0),.dout(w_dff_B_5adj63mH4_0),.clk(gclk));
	jdff dff_B_raffp4Gz1_0(.din(w_dff_B_5adj63mH4_0),.dout(w_dff_B_raffp4Gz1_0),.clk(gclk));
	jdff dff_B_DStWDLom9_0(.din(w_dff_B_raffp4Gz1_0),.dout(w_dff_B_DStWDLom9_0),.clk(gclk));
	jdff dff_B_nOi1Eb6f7_0(.din(w_dff_B_DStWDLom9_0),.dout(w_dff_B_nOi1Eb6f7_0),.clk(gclk));
	jdff dff_B_LiCEL3ez6_0(.din(w_dff_B_nOi1Eb6f7_0),.dout(w_dff_B_LiCEL3ez6_0),.clk(gclk));
	jdff dff_B_ndLxsYM54_0(.din(w_dff_B_LiCEL3ez6_0),.dout(w_dff_B_ndLxsYM54_0),.clk(gclk));
	jdff dff_A_vIxuH3bn2_1(.dout(w_n1609_0[1]),.din(w_dff_A_vIxuH3bn2_1),.clk(gclk));
	jdff dff_A_ySeyDz0k8_1(.dout(w_dff_A_vIxuH3bn2_1),.din(w_dff_A_ySeyDz0k8_1),.clk(gclk));
	jdff dff_A_sYySZKhM7_1(.dout(w_dff_A_ySeyDz0k8_1),.din(w_dff_A_sYySZKhM7_1),.clk(gclk));
	jdff dff_A_iAeNujxT2_1(.dout(w_dff_A_sYySZKhM7_1),.din(w_dff_A_iAeNujxT2_1),.clk(gclk));
	jdff dff_A_GuEfVYmM7_1(.dout(w_dff_A_iAeNujxT2_1),.din(w_dff_A_GuEfVYmM7_1),.clk(gclk));
	jdff dff_A_nngtRCkn2_1(.dout(w_dff_A_GuEfVYmM7_1),.din(w_dff_A_nngtRCkn2_1),.clk(gclk));
	jdff dff_A_28AHSCOU8_1(.dout(w_dff_A_nngtRCkn2_1),.din(w_dff_A_28AHSCOU8_1),.clk(gclk));
	jdff dff_A_ljhqv3wv9_1(.dout(w_dff_A_28AHSCOU8_1),.din(w_dff_A_ljhqv3wv9_1),.clk(gclk));
	jdff dff_A_of8p1i5s4_1(.dout(w_dff_A_ljhqv3wv9_1),.din(w_dff_A_of8p1i5s4_1),.clk(gclk));
	jdff dff_A_V7FRgrat5_1(.dout(w_dff_A_of8p1i5s4_1),.din(w_dff_A_V7FRgrat5_1),.clk(gclk));
	jdff dff_A_G7nwF14k6_1(.dout(w_dff_A_V7FRgrat5_1),.din(w_dff_A_G7nwF14k6_1),.clk(gclk));
	jdff dff_A_h5shk5OM9_1(.dout(w_dff_A_G7nwF14k6_1),.din(w_dff_A_h5shk5OM9_1),.clk(gclk));
	jdff dff_A_kssqCnv77_1(.dout(w_dff_A_h5shk5OM9_1),.din(w_dff_A_kssqCnv77_1),.clk(gclk));
	jdff dff_A_Qq1Quq655_1(.dout(w_dff_A_kssqCnv77_1),.din(w_dff_A_Qq1Quq655_1),.clk(gclk));
	jdff dff_A_aEH3TtKE1_1(.dout(w_dff_A_Qq1Quq655_1),.din(w_dff_A_aEH3TtKE1_1),.clk(gclk));
	jdff dff_A_zUepeZO53_1(.dout(w_dff_A_aEH3TtKE1_1),.din(w_dff_A_zUepeZO53_1),.clk(gclk));
	jdff dff_A_Pfw3SXlD2_1(.dout(w_dff_A_zUepeZO53_1),.din(w_dff_A_Pfw3SXlD2_1),.clk(gclk));
	jdff dff_A_3XaApVro6_1(.dout(w_dff_A_Pfw3SXlD2_1),.din(w_dff_A_3XaApVro6_1),.clk(gclk));
	jdff dff_A_1waapGIX9_1(.dout(w_dff_A_3XaApVro6_1),.din(w_dff_A_1waapGIX9_1),.clk(gclk));
	jdff dff_A_iMMMSng30_1(.dout(w_dff_A_1waapGIX9_1),.din(w_dff_A_iMMMSng30_1),.clk(gclk));
	jdff dff_B_BHeKXnXZ2_1(.din(n1392),.dout(w_dff_B_BHeKXnXZ2_1),.clk(gclk));
	jdff dff_B_KVlBrTpP5_1(.din(w_dff_B_BHeKXnXZ2_1),.dout(w_dff_B_KVlBrTpP5_1),.clk(gclk));
	jdff dff_B_WefEbtTG6_1(.din(w_dff_B_KVlBrTpP5_1),.dout(w_dff_B_WefEbtTG6_1),.clk(gclk));
	jdff dff_B_jam0XCMa2_1(.din(w_dff_B_WefEbtTG6_1),.dout(w_dff_B_jam0XCMa2_1),.clk(gclk));
	jdff dff_B_5n2VQ88Z8_1(.din(w_dff_B_jam0XCMa2_1),.dout(w_dff_B_5n2VQ88Z8_1),.clk(gclk));
	jdff dff_B_jqjgnu9Y6_1(.din(w_dff_B_5n2VQ88Z8_1),.dout(w_dff_B_jqjgnu9Y6_1),.clk(gclk));
	jdff dff_A_0WWrV3Qm4_1(.dout(w_n1447_0[1]),.din(w_dff_A_0WWrV3Qm4_1),.clk(gclk));
	jdff dff_B_0IsRCJ7J0_1(.din(n1412),.dout(w_dff_B_0IsRCJ7J0_1),.clk(gclk));
	jdff dff_B_ToTGSQCL8_1(.din(w_dff_B_0IsRCJ7J0_1),.dout(w_dff_B_ToTGSQCL8_1),.clk(gclk));
	jdff dff_B_B9H9mwxN9_1(.din(w_dff_B_ToTGSQCL8_1),.dout(w_dff_B_B9H9mwxN9_1),.clk(gclk));
	jdff dff_B_5T2WGnII4_1(.din(w_dff_B_B9H9mwxN9_1),.dout(w_dff_B_5T2WGnII4_1),.clk(gclk));
	jdff dff_B_8GDfDaZf7_1(.din(w_dff_B_5T2WGnII4_1),.dout(w_dff_B_8GDfDaZf7_1),.clk(gclk));
	jdff dff_B_9VPRZAvV0_1(.din(w_dff_B_8GDfDaZf7_1),.dout(w_dff_B_9VPRZAvV0_1),.clk(gclk));
	jdff dff_B_jqkJz3wv9_1(.din(w_dff_B_9VPRZAvV0_1),.dout(w_dff_B_jqkJz3wv9_1),.clk(gclk));
	jdff dff_B_Ot29YlhJ6_1(.din(w_dff_B_jqkJz3wv9_1),.dout(w_dff_B_Ot29YlhJ6_1),.clk(gclk));
	jdff dff_B_Ot9mHkHa8_1(.din(w_dff_B_Ot29YlhJ6_1),.dout(w_dff_B_Ot9mHkHa8_1),.clk(gclk));
	jdff dff_B_tMFsKl7A6_1(.din(w_dff_B_Ot9mHkHa8_1),.dout(w_dff_B_tMFsKl7A6_1),.clk(gclk));
	jdff dff_B_eVVXfIIu3_0(.din(n1443),.dout(w_dff_B_eVVXfIIu3_0),.clk(gclk));
	jdff dff_B_kNcJBDK78_0(.din(n1440),.dout(w_dff_B_kNcJBDK78_0),.clk(gclk));
	jdff dff_A_QDCpwcuD4_1(.dout(w_n1438_0[1]),.din(w_dff_A_QDCpwcuD4_1),.clk(gclk));
	jdff dff_A_WZ674L7l1_1(.dout(w_dff_A_QDCpwcuD4_1),.din(w_dff_A_WZ674L7l1_1),.clk(gclk));
	jdff dff_A_oUO70yLF7_1(.dout(w_dff_A_WZ674L7l1_1),.din(w_dff_A_oUO70yLF7_1),.clk(gclk));
	jdff dff_B_E8ELHlzE2_0(.din(n1437),.dout(w_dff_B_E8ELHlzE2_0),.clk(gclk));
	jdff dff_B_hmBEblHa7_1(.din(n1427),.dout(w_dff_B_hmBEblHa7_1),.clk(gclk));
	jdff dff_B_IYst7Amn4_1(.din(n1428),.dout(w_dff_B_IYst7Amn4_1),.clk(gclk));
	jdff dff_B_8uPzYekn1_1(.din(w_dff_B_IYst7Amn4_1),.dout(w_dff_B_8uPzYekn1_1),.clk(gclk));
	jdff dff_B_g9ldojdN6_1(.din(w_dff_B_8uPzYekn1_1),.dout(w_dff_B_g9ldojdN6_1),.clk(gclk));
	jdff dff_B_aC24Z1dY1_1(.din(w_dff_B_g9ldojdN6_1),.dout(w_dff_B_aC24Z1dY1_1),.clk(gclk));
	jdff dff_B_BZbrv8zs5_1(.din(w_dff_B_aC24Z1dY1_1),.dout(w_dff_B_BZbrv8zs5_1),.clk(gclk));
	jdff dff_B_Tn6q7SvF2_1(.din(w_dff_B_BZbrv8zs5_1),.dout(w_dff_B_Tn6q7SvF2_1),.clk(gclk));
	jdff dff_B_42Ps8CYr7_1(.din(w_dff_B_Tn6q7SvF2_1),.dout(w_dff_B_42Ps8CYr7_1),.clk(gclk));
	jdff dff_B_WbCOkQ0C7_1(.din(w_dff_B_42Ps8CYr7_1),.dout(w_dff_B_WbCOkQ0C7_1),.clk(gclk));
	jdff dff_B_CnHwM22T6_1(.din(w_dff_B_WbCOkQ0C7_1),.dout(w_dff_B_CnHwM22T6_1),.clk(gclk));
	jdff dff_B_41ZhxqkA9_1(.din(w_dff_B_CnHwM22T6_1),.dout(w_dff_B_41ZhxqkA9_1),.clk(gclk));
	jdff dff_B_nf95VBKY2_1(.din(w_dff_B_41ZhxqkA9_1),.dout(w_dff_B_nf95VBKY2_1),.clk(gclk));
	jdff dff_B_3XZyGNpK2_1(.din(n1414),.dout(w_dff_B_3XZyGNpK2_1),.clk(gclk));
	jdff dff_B_UFy47rG22_1(.din(w_dff_B_3XZyGNpK2_1),.dout(w_dff_B_UFy47rG22_1),.clk(gclk));
	jdff dff_B_fiyu5Gxj7_1(.din(w_dff_B_UFy47rG22_1),.dout(w_dff_B_fiyu5Gxj7_1),.clk(gclk));
	jdff dff_B_y49ND7CU4_1(.din(w_dff_B_fiyu5Gxj7_1),.dout(w_dff_B_y49ND7CU4_1),.clk(gclk));
	jdff dff_B_OTErftW91_1(.din(n1423),.dout(w_dff_B_OTErftW91_1),.clk(gclk));
	jdff dff_B_1KhJuAEY4_0(.din(n1422),.dout(w_dff_B_1KhJuAEY4_0),.clk(gclk));
	jdff dff_A_4fcUXYff2_0(.dout(w_n1421_0[0]),.din(w_dff_A_4fcUXYff2_0),.clk(gclk));
	jdff dff_A_brSy7YNQ1_0(.dout(w_dff_A_4fcUXYff2_0),.din(w_dff_A_brSy7YNQ1_0),.clk(gclk));
	jdff dff_A_XpGcU9sY8_0(.dout(w_dff_A_brSy7YNQ1_0),.din(w_dff_A_XpGcU9sY8_0),.clk(gclk));
	jdff dff_B_76ZUcUfQ7_1(.din(n1415),.dout(w_dff_B_76ZUcUfQ7_1),.clk(gclk));
	jdff dff_A_FkPSMB6o6_1(.dout(w_n829_0[1]),.din(w_dff_A_FkPSMB6o6_1),.clk(gclk));
	jdff dff_A_zZCI2VO65_0(.dout(w_n614_1[0]),.din(w_dff_A_zZCI2VO65_0),.clk(gclk));
	jdff dff_A_xMc5mXMI1_0(.dout(w_dff_A_zZCI2VO65_0),.din(w_dff_A_xMc5mXMI1_0),.clk(gclk));
	jdff dff_A_QI8vLCMf4_0(.dout(w_dff_A_xMc5mXMI1_0),.din(w_dff_A_QI8vLCMf4_0),.clk(gclk));
	jdff dff_A_FdhXM2JR2_0(.dout(w_dff_A_QI8vLCMf4_0),.din(w_dff_A_FdhXM2JR2_0),.clk(gclk));
	jdff dff_A_VCistAtS2_0(.dout(w_dff_A_FdhXM2JR2_0),.din(w_dff_A_VCistAtS2_0),.clk(gclk));
	jdff dff_A_09s7L97M0_2(.dout(w_n614_1[2]),.din(w_dff_A_09s7L97M0_2),.clk(gclk));
	jdff dff_A_FTyIHLeY4_2(.dout(w_dff_A_09s7L97M0_2),.din(w_dff_A_FTyIHLeY4_2),.clk(gclk));
	jdff dff_A_qYfta7xC9_2(.dout(w_dff_A_FTyIHLeY4_2),.din(w_dff_A_qYfta7xC9_2),.clk(gclk));
	jdff dff_A_hH9bAMMd6_2(.dout(w_dff_A_qYfta7xC9_2),.din(w_dff_A_hH9bAMMd6_2),.clk(gclk));
	jdff dff_A_oyGDJ2Jt1_2(.dout(w_dff_A_hH9bAMMd6_2),.din(w_dff_A_oyGDJ2Jt1_2),.clk(gclk));
	jdff dff_A_p8xOZy5d0_2(.dout(w_dff_A_oyGDJ2Jt1_2),.din(w_dff_A_p8xOZy5d0_2),.clk(gclk));
	jdff dff_A_BCiL83yU1_1(.dout(w_n828_0[1]),.din(w_dff_A_BCiL83yU1_1),.clk(gclk));
	jdff dff_A_6d1ddAg80_1(.dout(w_dff_A_BCiL83yU1_1),.din(w_dff_A_6d1ddAg80_1),.clk(gclk));
	jdff dff_A_C3xtNIXA3_1(.dout(w_dff_A_6d1ddAg80_1),.din(w_dff_A_C3xtNIXA3_1),.clk(gclk));
	jdff dff_A_iRhT1CDt2_1(.dout(w_dff_A_C3xtNIXA3_1),.din(w_dff_A_iRhT1CDt2_1),.clk(gclk));
	jdff dff_A_7FCyCoJM5_1(.dout(w_dff_A_iRhT1CDt2_1),.din(w_dff_A_7FCyCoJM5_1),.clk(gclk));
	jdff dff_A_7jdad2lW2_1(.dout(w_dff_A_7FCyCoJM5_1),.din(w_dff_A_7jdad2lW2_1),.clk(gclk));
	jdff dff_A_T5NMb1MX1_2(.dout(w_n828_0[2]),.din(w_dff_A_T5NMb1MX1_2),.clk(gclk));
	jdff dff_A_OJIT8lba9_2(.dout(w_dff_A_T5NMb1MX1_2),.din(w_dff_A_OJIT8lba9_2),.clk(gclk));
	jdff dff_B_Mh3JndIn2_2(.din(n787),.dout(w_dff_B_Mh3JndIn2_2),.clk(gclk));
	jdff dff_B_MZQNFqqM5_2(.din(w_dff_B_Mh3JndIn2_2),.dout(w_dff_B_MZQNFqqM5_2),.clk(gclk));
	jdff dff_B_rNOq08aD8_2(.din(w_dff_B_MZQNFqqM5_2),.dout(w_dff_B_rNOq08aD8_2),.clk(gclk));
	jdff dff_B_Yd3RaHDl1_2(.din(w_dff_B_rNOq08aD8_2),.dout(w_dff_B_Yd3RaHDl1_2),.clk(gclk));
	jdff dff_B_TVIXFEki8_2(.din(w_dff_B_Yd3RaHDl1_2),.dout(w_dff_B_TVIXFEki8_2),.clk(gclk));
	jdff dff_B_phM7qrV39_2(.din(w_dff_B_TVIXFEki8_2),.dout(w_dff_B_phM7qrV39_2),.clk(gclk));
	jdff dff_B_GgWPJpw72_2(.din(w_dff_B_phM7qrV39_2),.dout(w_dff_B_GgWPJpw72_2),.clk(gclk));
	jdff dff_B_ROTYPJsD2_2(.din(w_dff_B_GgWPJpw72_2),.dout(w_dff_B_ROTYPJsD2_2),.clk(gclk));
	jdff dff_B_FSISOWg23_2(.din(w_dff_B_ROTYPJsD2_2),.dout(w_dff_B_FSISOWg23_2),.clk(gclk));
	jdff dff_A_rcpRD7dV0_1(.dout(w_n779_0[1]),.din(w_dff_A_rcpRD7dV0_1),.clk(gclk));
	jdff dff_A_nLpx2NTb8_1(.dout(w_dff_A_rcpRD7dV0_1),.din(w_dff_A_nLpx2NTb8_1),.clk(gclk));
	jdff dff_A_yCOEN5au0_1(.dout(w_dff_A_nLpx2NTb8_1),.din(w_dff_A_yCOEN5au0_1),.clk(gclk));
	jdff dff_A_Ml2bBaEz1_1(.dout(w_dff_A_yCOEN5au0_1),.din(w_dff_A_Ml2bBaEz1_1),.clk(gclk));
	jdff dff_A_67u18kr91_1(.dout(w_dff_A_Ml2bBaEz1_1),.din(w_dff_A_67u18kr91_1),.clk(gclk));
	jdff dff_A_c7oDginB8_1(.dout(w_dff_A_67u18kr91_1),.din(w_dff_A_c7oDginB8_1),.clk(gclk));
	jdff dff_A_wClsaO2M6_1(.dout(w_dff_A_c7oDginB8_1),.din(w_dff_A_wClsaO2M6_1),.clk(gclk));
	jdff dff_A_iWVUUbPu3_1(.dout(w_dff_A_wClsaO2M6_1),.din(w_dff_A_iWVUUbPu3_1),.clk(gclk));
	jdff dff_A_cYWoVSJP6_1(.dout(w_dff_A_iWVUUbPu3_1),.din(w_dff_A_cYWoVSJP6_1),.clk(gclk));
	jdff dff_A_ddv5fYwH6_1(.dout(w_dff_A_cYWoVSJP6_1),.din(w_dff_A_ddv5fYwH6_1),.clk(gclk));
	jdff dff_A_k26LsMPL1_1(.dout(w_dff_A_ddv5fYwH6_1),.din(w_dff_A_k26LsMPL1_1),.clk(gclk));
	jdff dff_A_MaU7TXpH9_1(.dout(w_dff_A_k26LsMPL1_1),.din(w_dff_A_MaU7TXpH9_1),.clk(gclk));
	jdff dff_A_ZP4UbCEf5_1(.dout(w_n636_1[1]),.din(w_dff_A_ZP4UbCEf5_1),.clk(gclk));
	jdff dff_A_l10nIiRm6_1(.dout(w_dff_A_ZP4UbCEf5_1),.din(w_dff_A_l10nIiRm6_1),.clk(gclk));
	jdff dff_A_6BEI3sAR2_2(.dout(w_n636_0[2]),.din(w_dff_A_6BEI3sAR2_2),.clk(gclk));
	jdff dff_A_4B1mheP25_0(.dout(w_n1411_0[0]),.din(w_dff_A_4B1mheP25_0),.clk(gclk));
	jdff dff_A_Gqh8Jh6F4_0(.dout(w_dff_A_4B1mheP25_0),.din(w_dff_A_Gqh8Jh6F4_0),.clk(gclk));
	jdff dff_A_fLXyLqX78_0(.dout(w_dff_A_Gqh8Jh6F4_0),.din(w_dff_A_fLXyLqX78_0),.clk(gclk));
	jdff dff_A_Of2vPbt25_0(.dout(w_dff_A_fLXyLqX78_0),.din(w_dff_A_Of2vPbt25_0),.clk(gclk));
	jdff dff_A_z6De8r066_0(.dout(w_dff_A_Of2vPbt25_0),.din(w_dff_A_z6De8r066_0),.clk(gclk));
	jdff dff_A_hVQnnvja8_0(.dout(w_dff_A_z6De8r066_0),.din(w_dff_A_hVQnnvja8_0),.clk(gclk));
	jdff dff_A_59eggMik5_0(.dout(w_dff_A_hVQnnvja8_0),.din(w_dff_A_59eggMik5_0),.clk(gclk));
	jdff dff_A_rsD7FIMN5_0(.dout(w_dff_A_59eggMik5_0),.din(w_dff_A_rsD7FIMN5_0),.clk(gclk));
	jdff dff_A_RcUXlHWv0_0(.dout(w_dff_A_rsD7FIMN5_0),.din(w_dff_A_RcUXlHWv0_0),.clk(gclk));
	jdff dff_A_WaAZAjwT5_0(.dout(w_dff_A_RcUXlHWv0_0),.din(w_dff_A_WaAZAjwT5_0),.clk(gclk));
	jdff dff_A_7HpJId9l8_0(.dout(w_dff_A_WaAZAjwT5_0),.din(w_dff_A_7HpJId9l8_0),.clk(gclk));
	jdff dff_A_nLPM3D7D0_0(.dout(w_n1409_0[0]),.din(w_dff_A_nLPM3D7D0_0),.clk(gclk));
	jdff dff_B_uCKs5HVf6_1(.din(n1405),.dout(w_dff_B_uCKs5HVf6_1),.clk(gclk));
	jdff dff_B_wtl9Oema5_0(.din(n1407),.dout(w_dff_B_wtl9Oema5_0),.clk(gclk));
	jdff dff_B_Flsaga4c0_0(.din(w_dff_B_wtl9Oema5_0),.dout(w_dff_B_Flsaga4c0_0),.clk(gclk));
	jdff dff_B_nXVhM1Rx0_0(.din(w_dff_B_Flsaga4c0_0),.dout(w_dff_B_nXVhM1Rx0_0),.clk(gclk));
	jdff dff_B_qscW8IVx3_0(.din(w_dff_B_nXVhM1Rx0_0),.dout(w_dff_B_qscW8IVx3_0),.clk(gclk));
	jdff dff_A_iLfKEUtW7_1(.dout(w_n968_0[1]),.din(w_dff_A_iLfKEUtW7_1),.clk(gclk));
	jdff dff_A_PXyvd2ks5_1(.dout(w_dff_A_iLfKEUtW7_1),.din(w_dff_A_PXyvd2ks5_1),.clk(gclk));
	jdff dff_A_9O5UXZ154_1(.dout(w_dff_A_PXyvd2ks5_1),.din(w_dff_A_9O5UXZ154_1),.clk(gclk));
	jdff dff_A_qFTtFlRi2_1(.dout(w_dff_A_9O5UXZ154_1),.din(w_dff_A_qFTtFlRi2_1),.clk(gclk));
	jdff dff_A_RjAXddZ37_1(.dout(w_dff_A_qFTtFlRi2_1),.din(w_dff_A_RjAXddZ37_1),.clk(gclk));
	jdff dff_B_kt9B0qJD9_2(.din(n968),.dout(w_dff_B_kt9B0qJD9_2),.clk(gclk));
	jdff dff_B_MOfdpE6P9_2(.din(w_dff_B_kt9B0qJD9_2),.dout(w_dff_B_MOfdpE6P9_2),.clk(gclk));
	jdff dff_B_Nj8WUajz9_2(.din(w_dff_B_MOfdpE6P9_2),.dout(w_dff_B_Nj8WUajz9_2),.clk(gclk));
	jdff dff_B_SLMTPtCs1_2(.din(w_dff_B_Nj8WUajz9_2),.dout(w_dff_B_SLMTPtCs1_2),.clk(gclk));
	jdff dff_B_BywBpOYm8_2(.din(w_dff_B_SLMTPtCs1_2),.dout(w_dff_B_BywBpOYm8_2),.clk(gclk));
	jdff dff_B_rZr6ZrTy5_0(.din(n1404),.dout(w_dff_B_rZr6ZrTy5_0),.clk(gclk));
	jdff dff_B_3RbFhSx97_0(.din(w_dff_B_rZr6ZrTy5_0),.dout(w_dff_B_3RbFhSx97_0),.clk(gclk));
	jdff dff_B_c2AMwgBo0_1(.din(n1401),.dout(w_dff_B_c2AMwgBo0_1),.clk(gclk));
	jdff dff_B_0prXEDw41_1(.din(w_dff_B_c2AMwgBo0_1),.dout(w_dff_B_0prXEDw41_1),.clk(gclk));
	jdff dff_B_ztEuUki02_1(.din(w_dff_B_0prXEDw41_1),.dout(w_dff_B_ztEuUki02_1),.clk(gclk));
	jdff dff_A_Cka2V7856_1(.dout(w_n651_0[1]),.din(w_dff_A_Cka2V7856_1),.clk(gclk));
	jdff dff_A_3wpdnrIV2_1(.dout(w_dff_A_Cka2V7856_1),.din(w_dff_A_3wpdnrIV2_1),.clk(gclk));
	jdff dff_A_tPlTKaWH6_1(.dout(w_dff_A_3wpdnrIV2_1),.din(w_dff_A_tPlTKaWH6_1),.clk(gclk));
	jdff dff_A_dhReTvlB7_2(.dout(w_n651_0[2]),.din(w_dff_A_dhReTvlB7_2),.clk(gclk));
	jdff dff_A_ePq601SJ4_2(.dout(w_dff_A_dhReTvlB7_2),.din(w_dff_A_ePq601SJ4_2),.clk(gclk));
	jdff dff_A_GxFhgmSn1_2(.dout(w_dff_A_ePq601SJ4_2),.din(w_dff_A_GxFhgmSn1_2),.clk(gclk));
	jdff dff_A_CsVBg2om0_2(.dout(w_dff_A_GxFhgmSn1_2),.din(w_dff_A_CsVBg2om0_2),.clk(gclk));
	jdff dff_A_fREJw3An9_2(.dout(w_dff_A_CsVBg2om0_2),.din(w_dff_A_fREJw3An9_2),.clk(gclk));
	jdff dff_A_U6OwVIsN2_2(.dout(w_dff_A_fREJw3An9_2),.din(w_dff_A_U6OwVIsN2_2),.clk(gclk));
	jdff dff_A_HqFGmp4m9_2(.dout(w_dff_A_U6OwVIsN2_2),.din(w_dff_A_HqFGmp4m9_2),.clk(gclk));
	jdff dff_B_HqYOc0uM0_3(.din(n651),.dout(w_dff_B_HqYOc0uM0_3),.clk(gclk));
	jdff dff_A_y7xTsVOc6_0(.dout(w_n650_0[0]),.din(w_dff_A_y7xTsVOc6_0),.clk(gclk));
	jdff dff_A_kun5VUET6_0(.dout(w_dff_A_y7xTsVOc6_0),.din(w_dff_A_kun5VUET6_0),.clk(gclk));
	jdff dff_A_tBp2Hsn68_0(.dout(w_dff_A_kun5VUET6_0),.din(w_dff_A_tBp2Hsn68_0),.clk(gclk));
	jdff dff_A_jYxV5az43_0(.dout(w_dff_A_tBp2Hsn68_0),.din(w_dff_A_jYxV5az43_0),.clk(gclk));
	jdff dff_A_ssGrBkRW2_0(.dout(w_dff_A_jYxV5az43_0),.din(w_dff_A_ssGrBkRW2_0),.clk(gclk));
	jdff dff_A_axq4HGjQ0_0(.dout(w_dff_A_ssGrBkRW2_0),.din(w_dff_A_axq4HGjQ0_0),.clk(gclk));
	jdff dff_A_Ussb0dT78_0(.dout(w_dff_A_axq4HGjQ0_0),.din(w_dff_A_Ussb0dT78_0),.clk(gclk));
	jdff dff_A_L14DxMQa2_0(.dout(w_dff_A_Ussb0dT78_0),.din(w_dff_A_L14DxMQa2_0),.clk(gclk));
	jdff dff_A_Td0FQIsI3_0(.dout(w_dff_A_L14DxMQa2_0),.din(w_dff_A_Td0FQIsI3_0),.clk(gclk));
	jdff dff_B_4M2MQAlr4_1(.din(n1395),.dout(w_dff_B_4M2MQAlr4_1),.clk(gclk));
	jdff dff_A_NgjfhL585_1(.dout(w_n740_0[1]),.din(w_dff_A_NgjfhL585_1),.clk(gclk));
	jdff dff_A_9b00a6Wm0_0(.dout(w_n739_1[0]),.din(w_dff_A_9b00a6Wm0_0),.clk(gclk));
	jdff dff_A_WM9O4aQN3_0(.dout(w_dff_A_9b00a6Wm0_0),.din(w_dff_A_WM9O4aQN3_0),.clk(gclk));
	jdff dff_A_PziGP8hv4_0(.dout(w_dff_A_WM9O4aQN3_0),.din(w_dff_A_PziGP8hv4_0),.clk(gclk));
	jdff dff_A_R3Yk2wKz5_0(.dout(w_dff_A_PziGP8hv4_0),.din(w_dff_A_R3Yk2wKz5_0),.clk(gclk));
	jdff dff_A_ZSZNXX9l0_0(.dout(w_dff_A_R3Yk2wKz5_0),.din(w_dff_A_ZSZNXX9l0_0),.clk(gclk));
	jdff dff_A_VEFizTQq6_0(.dout(w_dff_A_ZSZNXX9l0_0),.din(w_dff_A_VEFizTQq6_0),.clk(gclk));
	jdff dff_A_D3LNxEph9_0(.dout(w_dff_A_VEFizTQq6_0),.din(w_dff_A_D3LNxEph9_0),.clk(gclk));
	jdff dff_A_7OoVbUce7_0(.dout(w_dff_A_D3LNxEph9_0),.din(w_dff_A_7OoVbUce7_0),.clk(gclk));
	jdff dff_A_0Yj7e50W7_0(.dout(w_dff_A_7OoVbUce7_0),.din(w_dff_A_0Yj7e50W7_0),.clk(gclk));
	jdff dff_A_rcOAliD40_2(.dout(w_n739_0[2]),.din(w_dff_A_rcOAliD40_2),.clk(gclk));
	jdff dff_A_vuGKH9bt2_2(.dout(w_dff_A_rcOAliD40_2),.din(w_dff_A_vuGKH9bt2_2),.clk(gclk));
	jdff dff_A_3fHr742m8_2(.dout(w_dff_A_vuGKH9bt2_2),.din(w_dff_A_3fHr742m8_2),.clk(gclk));
	jdff dff_A_rjE4E3PC6_2(.dout(w_dff_A_3fHr742m8_2),.din(w_dff_A_rjE4E3PC6_2),.clk(gclk));
	jdff dff_A_ZiHBGFqw1_2(.dout(w_dff_A_rjE4E3PC6_2),.din(w_dff_A_ZiHBGFqw1_2),.clk(gclk));
	jdff dff_A_h601iIzf1_2(.dout(w_n649_0[2]),.din(w_dff_A_h601iIzf1_2),.clk(gclk));
	jdff dff_B_ajomxJhW9_0(.din(n648),.dout(w_dff_B_ajomxJhW9_0),.clk(gclk));
	jdff dff_B_OVby5Z5C3_1(.din(G323),.dout(w_dff_B_OVby5Z5C3_1),.clk(gclk));
	jdff dff_A_9Z8YzaJR0_0(.dout(w_n640_1[0]),.din(w_dff_A_9Z8YzaJR0_0),.clk(gclk));
	jdff dff_A_hoLr25wI1_0(.dout(w_dff_A_9Z8YzaJR0_0),.din(w_dff_A_hoLr25wI1_0),.clk(gclk));
	jdff dff_A_333dDAbD8_0(.dout(w_dff_A_hoLr25wI1_0),.din(w_dff_A_333dDAbD8_0),.clk(gclk));
	jdff dff_A_1Cp6KO1i0_0(.dout(w_dff_A_333dDAbD8_0),.din(w_dff_A_1Cp6KO1i0_0),.clk(gclk));
	jdff dff_A_HHnB3VB34_0(.dout(w_dff_A_1Cp6KO1i0_0),.din(w_dff_A_HHnB3VB34_0),.clk(gclk));
	jdff dff_A_neDUdMgU6_0(.dout(w_dff_A_HHnB3VB34_0),.din(w_dff_A_neDUdMgU6_0),.clk(gclk));
	jdff dff_A_VNnF3vLh9_0(.dout(w_dff_A_neDUdMgU6_0),.din(w_dff_A_VNnF3vLh9_0),.clk(gclk));
	jdff dff_A_Ucl5ZpZa5_0(.dout(w_dff_A_VNnF3vLh9_0),.din(w_dff_A_Ucl5ZpZa5_0),.clk(gclk));
	jdff dff_A_78w0CKoW7_0(.dout(w_dff_A_Ucl5ZpZa5_0),.din(w_dff_A_78w0CKoW7_0),.clk(gclk));
	jdff dff_A_Ln1P0pbx4_0(.dout(w_dff_A_78w0CKoW7_0),.din(w_dff_A_Ln1P0pbx4_0),.clk(gclk));
	jdff dff_A_D7AxmQ9P6_0(.dout(w_dff_A_Ln1P0pbx4_0),.din(w_dff_A_D7AxmQ9P6_0),.clk(gclk));
	jdff dff_A_4ZtY3t7X9_0(.dout(w_n646_0[0]),.din(w_dff_A_4ZtY3t7X9_0),.clk(gclk));
	jdff dff_A_6BIevfPr4_0(.dout(w_dff_A_4ZtY3t7X9_0),.din(w_dff_A_6BIevfPr4_0),.clk(gclk));
	jdff dff_B_UOnL0LPK6_0(.din(n644),.dout(w_dff_B_UOnL0LPK6_0),.clk(gclk));
	jdff dff_B_5Qogf0L47_1(.din(G315),.dout(w_dff_B_5Qogf0L47_1),.clk(gclk));
	jdff dff_A_1SvuEk1l6_1(.dout(w_n640_0[1]),.din(w_dff_A_1SvuEk1l6_1),.clk(gclk));
	jdff dff_A_T34XIiGr7_2(.dout(w_n640_0[2]),.din(w_dff_A_T34XIiGr7_2),.clk(gclk));
	jdff dff_A_Un4by8Su6_2(.dout(w_dff_A_T34XIiGr7_2),.din(w_dff_A_Un4by8Su6_2),.clk(gclk));
	jdff dff_A_TBuxjPfM6_2(.dout(w_dff_A_Un4by8Su6_2),.din(w_dff_A_TBuxjPfM6_2),.clk(gclk));
	jdff dff_A_PZ46vJmd6_2(.dout(w_dff_A_TBuxjPfM6_2),.din(w_dff_A_PZ46vJmd6_2),.clk(gclk));
	jdff dff_A_b6iIEez91_2(.dout(w_dff_A_PZ46vJmd6_2),.din(w_dff_A_b6iIEez91_2),.clk(gclk));
	jdff dff_A_tE1zBRHh8_2(.dout(w_dff_A_b6iIEez91_2),.din(w_dff_A_tE1zBRHh8_2),.clk(gclk));
	jdff dff_A_gpHzgrZb4_2(.dout(w_dff_A_tE1zBRHh8_2),.din(w_dff_A_gpHzgrZb4_2),.clk(gclk));
	jdff dff_A_Nj4cffsC8_2(.dout(w_dff_A_gpHzgrZb4_2),.din(w_dff_A_Nj4cffsC8_2),.clk(gclk));
	jdff dff_A_zDCSsXC69_2(.dout(w_dff_A_Nj4cffsC8_2),.din(w_dff_A_zDCSsXC69_2),.clk(gclk));
	jdff dff_A_FCeaU0Lj3_2(.dout(w_dff_A_zDCSsXC69_2),.din(w_dff_A_FCeaU0Lj3_2),.clk(gclk));
	jdff dff_A_LO8JhS1b5_2(.dout(w_dff_A_FCeaU0Lj3_2),.din(w_dff_A_LO8JhS1b5_2),.clk(gclk));
	jdff dff_B_wQ37Nmac5_1(.din(n637),.dout(w_dff_B_wQ37Nmac5_1),.clk(gclk));
	jdff dff_B_Cqd1kKUi5_1(.din(G307),.dout(w_dff_B_Cqd1kKUi5_1),.clk(gclk));
	jdff dff_B_ueR6QxYH8_0(.din(n1393),.dout(w_dff_B_ueR6QxYH8_0),.clk(gclk));
	jdff dff_B_0n2iSvza1_0(.din(w_dff_B_ueR6QxYH8_0),.dout(w_dff_B_0n2iSvza1_0),.clk(gclk));
	jdff dff_B_sTEgEJtc9_0(.din(w_dff_B_0n2iSvza1_0),.dout(w_dff_B_sTEgEJtc9_0),.clk(gclk));
	jdff dff_A_tVf5I4i34_0(.dout(w_n631_0[0]),.din(w_dff_A_tVf5I4i34_0),.clk(gclk));
	jdff dff_A_TGiwqkbc7_0(.dout(w_dff_A_tVf5I4i34_0),.din(w_dff_A_TGiwqkbc7_0),.clk(gclk));
	jdff dff_A_BHyEiyWj8_0(.dout(w_dff_A_TGiwqkbc7_0),.din(w_dff_A_BHyEiyWj8_0),.clk(gclk));
	jdff dff_A_gRJu8dra0_1(.dout(w_n629_0[1]),.din(w_dff_A_gRJu8dra0_1),.clk(gclk));
	jdff dff_A_PaftL0gZ0_1(.dout(w_dff_A_gRJu8dra0_1),.din(w_dff_A_PaftL0gZ0_1),.clk(gclk));
	jdff dff_A_t9pJYt2t9_1(.dout(w_dff_A_PaftL0gZ0_1),.din(w_dff_A_t9pJYt2t9_1),.clk(gclk));
	jdff dff_A_OuIvP6MH8_1(.dout(w_n628_0[1]),.din(w_dff_A_OuIvP6MH8_1),.clk(gclk));
	jdff dff_B_sy6KjLuo3_0(.din(n627),.dout(w_dff_B_sy6KjLuo3_0),.clk(gclk));
	jdff dff_A_6FBPsbun8_0(.dout(w_n625_0[0]),.din(w_dff_A_6FBPsbun8_0),.clk(gclk));
	jdff dff_A_zIdAlXXi9_2(.dout(w_n625_0[2]),.din(w_dff_A_zIdAlXXi9_2),.clk(gclk));
	jdff dff_A_VdAWrNPu1_0(.dout(w_n623_0[0]),.din(w_dff_A_VdAWrNPu1_0),.clk(gclk));
	jdff dff_B_rRKEK39E6_0(.din(n616),.dout(w_dff_B_rRKEK39E6_0),.clk(gclk));
	jdff dff_A_3lcgRqEX1_0(.dout(w_G2174_0[0]),.din(w_dff_A_3lcgRqEX1_0),.clk(gclk));
	jdff dff_A_Pf5VAkFP8_0(.dout(w_dff_A_3lcgRqEX1_0),.din(w_dff_A_Pf5VAkFP8_0),.clk(gclk));
	jdff dff_A_sXQc0UB34_0(.dout(w_dff_A_Pf5VAkFP8_0),.din(w_dff_A_sXQc0UB34_0),.clk(gclk));
	jdff dff_A_bGQnNttp7_0(.dout(w_dff_A_sXQc0UB34_0),.din(w_dff_A_bGQnNttp7_0),.clk(gclk));
	jdff dff_A_NTRfhQdx2_0(.dout(w_dff_A_bGQnNttp7_0),.din(w_dff_A_NTRfhQdx2_0),.clk(gclk));
	jdff dff_A_hgT2m9R40_0(.dout(w_dff_A_NTRfhQdx2_0),.din(w_dff_A_hgT2m9R40_0),.clk(gclk));
	jdff dff_A_x0rP3c8Z5_0(.dout(w_dff_A_hgT2m9R40_0),.din(w_dff_A_x0rP3c8Z5_0),.clk(gclk));
	jdff dff_A_FRltRma56_0(.dout(w_dff_A_x0rP3c8Z5_0),.din(w_dff_A_FRltRma56_0),.clk(gclk));
	jdff dff_A_Px5ZGXrK0_0(.dout(w_dff_A_FRltRma56_0),.din(w_dff_A_Px5ZGXrK0_0),.clk(gclk));
	jdff dff_A_uaJnVHqy2_0(.dout(w_dff_A_Px5ZGXrK0_0),.din(w_dff_A_uaJnVHqy2_0),.clk(gclk));
	jdff dff_A_Z08EWguM7_0(.dout(w_dff_A_uaJnVHqy2_0),.din(w_dff_A_Z08EWguM7_0),.clk(gclk));
	jdff dff_A_l5bz6pxi6_2(.dout(w_G2174_0[2]),.din(w_dff_A_l5bz6pxi6_2),.clk(gclk));
	jdff dff_A_16V4Hxzh5_2(.dout(w_dff_A_l5bz6pxi6_2),.din(w_dff_A_16V4Hxzh5_2),.clk(gclk));
	jdff dff_A_fixQuJMB8_2(.dout(w_dff_A_16V4Hxzh5_2),.din(w_dff_A_fixQuJMB8_2),.clk(gclk));
	jdff dff_A_hoAfj9jr7_2(.dout(w_dff_A_fixQuJMB8_2),.din(w_dff_A_hoAfj9jr7_2),.clk(gclk));
	jdff dff_A_4GDP5TXL1_2(.dout(w_dff_A_hoAfj9jr7_2),.din(w_dff_A_4GDP5TXL1_2),.clk(gclk));
	jdff dff_A_1wQP34qU5_2(.dout(w_dff_A_4GDP5TXL1_2),.din(w_dff_A_1wQP34qU5_2),.clk(gclk));
	jdff dff_A_LwJ5T8GU8_2(.dout(w_dff_A_1wQP34qU5_2),.din(w_dff_A_LwJ5T8GU8_2),.clk(gclk));
	jdff dff_A_5KgIyjV38_2(.dout(w_dff_A_LwJ5T8GU8_2),.din(w_dff_A_5KgIyjV38_2),.clk(gclk));
	jdff dff_B_nwTId6tV3_1(.din(n711),.dout(w_dff_B_nwTId6tV3_1),.clk(gclk));
	jdff dff_B_TNNtcrsm6_1(.din(w_dff_B_nwTId6tV3_1),.dout(w_dff_B_TNNtcrsm6_1),.clk(gclk));
	jdff dff_B_BWdDp12D4_1(.din(w_dff_B_TNNtcrsm6_1),.dout(w_dff_B_BWdDp12D4_1),.clk(gclk));
	jdff dff_B_pZXcCq6v4_1(.din(w_dff_B_BWdDp12D4_1),.dout(w_dff_B_pZXcCq6v4_1),.clk(gclk));
	jdff dff_B_j3t6z3pP4_1(.din(w_dff_B_pZXcCq6v4_1),.dout(w_dff_B_j3t6z3pP4_1),.clk(gclk));
	jdff dff_B_37SCrA0S9_1(.din(w_dff_B_j3t6z3pP4_1),.dout(w_dff_B_37SCrA0S9_1),.clk(gclk));
	jdff dff_B_3iwYDHDS5_1(.din(n712),.dout(w_dff_B_3iwYDHDS5_1),.clk(gclk));
	jdff dff_B_36KGz4ig5_1(.din(w_dff_B_3iwYDHDS5_1),.dout(w_dff_B_36KGz4ig5_1),.clk(gclk));
	jdff dff_B_N3s96bPx9_1(.din(w_dff_B_36KGz4ig5_1),.dout(w_dff_B_N3s96bPx9_1),.clk(gclk));
	jdff dff_B_wvi7Aap69_1(.din(w_dff_B_N3s96bPx9_1),.dout(w_dff_B_wvi7Aap69_1),.clk(gclk));
	jdff dff_B_s7NA25D62_1(.din(w_dff_B_wvi7Aap69_1),.dout(w_dff_B_s7NA25D62_1),.clk(gclk));
	jdff dff_B_geJVyNwW7_1(.din(n713),.dout(w_dff_B_geJVyNwW7_1),.clk(gclk));
	jdff dff_B_32HAyE5l5_1(.din(w_dff_B_geJVyNwW7_1),.dout(w_dff_B_32HAyE5l5_1),.clk(gclk));
	jdff dff_B_RUmbkIb40_1(.din(w_dff_B_32HAyE5l5_1),.dout(w_dff_B_RUmbkIb40_1),.clk(gclk));
	jdff dff_B_zFRFbdqH0_1(.din(w_dff_B_RUmbkIb40_1),.dout(w_dff_B_zFRFbdqH0_1),.clk(gclk));
	jdff dff_A_2osJTg5r6_0(.dout(w_n723_0[0]),.din(w_dff_A_2osJTg5r6_0),.clk(gclk));
	jdff dff_A_64zhRRF94_0(.dout(w_n621_2[0]),.din(w_dff_A_64zhRRF94_0),.clk(gclk));
	jdff dff_A_lKBBG9nc4_1(.dout(w_n721_0[1]),.din(w_dff_A_lKBBG9nc4_1),.clk(gclk));
	jdff dff_A_iIioO9lY3_1(.dout(w_dff_A_lKBBG9nc4_1),.din(w_dff_A_iIioO9lY3_1),.clk(gclk));
	jdff dff_A_TpbrnZoO6_1(.dout(w_dff_A_iIioO9lY3_1),.din(w_dff_A_TpbrnZoO6_1),.clk(gclk));
	jdff dff_A_0gVNNokL9_1(.dout(w_dff_A_TpbrnZoO6_1),.din(w_dff_A_0gVNNokL9_1),.clk(gclk));
	jdff dff_A_1Lie9nTu7_1(.dout(w_dff_A_0gVNNokL9_1),.din(w_dff_A_1Lie9nTu7_1),.clk(gclk));
	jdff dff_A_RRSfynhV3_1(.dout(w_dff_A_1Lie9nTu7_1),.din(w_dff_A_RRSfynhV3_1),.clk(gclk));
	jdff dff_A_EcPFPxEC7_0(.dout(w_G358_0[0]),.din(w_dff_A_EcPFPxEC7_0),.clk(gclk));
	jdff dff_A_HIVMkKha8_0(.dout(w_n388_1[0]),.din(w_dff_A_HIVMkKha8_0),.clk(gclk));
	jdff dff_A_sYehwKfj0_1(.dout(w_n388_1[1]),.din(w_dff_A_sYehwKfj0_1),.clk(gclk));
	jdff dff_A_6ITWIBCe7_1(.dout(w_n717_0[1]),.din(w_dff_A_6ITWIBCe7_1),.clk(gclk));
	jdff dff_A_41tmBw654_1(.dout(w_dff_A_6ITWIBCe7_1),.din(w_dff_A_41tmBw654_1),.clk(gclk));
	jdff dff_A_b8mN4CkN8_1(.dout(w_dff_A_41tmBw654_1),.din(w_dff_A_b8mN4CkN8_1),.clk(gclk));
	jdff dff_A_tphtfBPB4_2(.dout(w_n717_0[2]),.din(w_dff_A_tphtfBPB4_2),.clk(gclk));
	jdff dff_A_VhxFh8dI9_2(.dout(w_dff_A_tphtfBPB4_2),.din(w_dff_A_VhxFh8dI9_2),.clk(gclk));
	jdff dff_A_F1MW2BrB7_0(.dout(w_G348_0[0]),.din(w_dff_A_F1MW2BrB7_0),.clk(gclk));
	jdff dff_A_SjAokIeW6_0(.dout(w_G332_2[0]),.din(w_dff_A_SjAokIeW6_0),.clk(gclk));
	jdff dff_A_wnFGLyFC2_0(.dout(w_n437_1[0]),.din(w_dff_A_wnFGLyFC2_0),.clk(gclk));
	jdff dff_A_W8kNSJ959_1(.dout(w_n437_1[1]),.din(w_dff_A_W8kNSJ959_1),.clk(gclk));
	jdff dff_A_CrsoojyL3_0(.dout(w_G332_3[0]),.din(w_dff_A_CrsoojyL3_0),.clk(gclk));
	jdff dff_A_iDRi8Z7q6_2(.dout(w_G332_3[2]),.din(w_dff_A_iDRi8Z7q6_2),.clk(gclk));
	jdff dff_A_RHDn8gJ77_0(.dout(w_n410_1[0]),.din(w_dff_A_RHDn8gJ77_0),.clk(gclk));
	jdff dff_A_NGjVTmbe1_0(.dout(w_n614_2[0]),.din(w_dff_A_NGjVTmbe1_0),.clk(gclk));
	jdff dff_A_Vfr0JD8t2_0(.dout(w_dff_A_NGjVTmbe1_0),.din(w_dff_A_Vfr0JD8t2_0),.clk(gclk));
	jdff dff_A_sPNwFVsy2_0(.dout(w_dff_A_Vfr0JD8t2_0),.din(w_dff_A_sPNwFVsy2_0),.clk(gclk));
	jdff dff_A_qTO4q7QN5_1(.dout(w_n614_0[1]),.din(w_dff_A_qTO4q7QN5_1),.clk(gclk));
	jdff dff_A_5lRKS5Go0_1(.dout(w_dff_A_qTO4q7QN5_1),.din(w_dff_A_5lRKS5Go0_1),.clk(gclk));
	jdff dff_A_vZh9OXyE6_2(.dout(w_n614_0[2]),.din(w_dff_A_vZh9OXyE6_2),.clk(gclk));
	jdff dff_A_DThUBnis6_2(.dout(w_dff_A_vZh9OXyE6_2),.din(w_dff_A_DThUBnis6_2),.clk(gclk));
	jdff dff_A_OnmdS1oM1_2(.dout(w_dff_A_DThUBnis6_2),.din(w_dff_A_OnmdS1oM1_2),.clk(gclk));
	jdff dff_A_0LLucqvu0_2(.dout(w_dff_A_OnmdS1oM1_2),.din(w_dff_A_0LLucqvu0_2),.clk(gclk));
	jdff dff_B_Tse1RMZe5_1(.din(n610),.dout(w_dff_B_Tse1RMZe5_1),.clk(gclk));
	jdff dff_A_EeOoDiHL9_0(.dout(w_G332_4[0]),.din(w_dff_A_EeOoDiHL9_0),.clk(gclk));
	jdff dff_A_XlcVMFwu1_2(.dout(w_G332_1[2]),.din(w_dff_A_XlcVMFwu1_2),.clk(gclk));
	jdff dff_A_AvITlxYr9_1(.dout(w_G331_0[1]),.din(w_dff_A_AvITlxYr9_1),.clk(gclk));
	jdff dff_A_8snwYWZG3_0(.dout(w_n1391_0[0]),.din(w_dff_A_8snwYWZG3_0),.clk(gclk));
	jdff dff_A_j84CDqMi4_0(.dout(w_dff_A_8snwYWZG3_0),.din(w_dff_A_j84CDqMi4_0),.clk(gclk));
	jdff dff_A_sF3fyNOK1_0(.dout(w_dff_A_j84CDqMi4_0),.din(w_dff_A_sF3fyNOK1_0),.clk(gclk));
	jdff dff_A_6suxaqd71_0(.dout(w_dff_A_sF3fyNOK1_0),.din(w_dff_A_6suxaqd71_0),.clk(gclk));
	jdff dff_A_1771ZTwu0_0(.dout(w_dff_A_6suxaqd71_0),.din(w_dff_A_1771ZTwu0_0),.clk(gclk));
	jdff dff_A_miAybj3Y3_0(.dout(w_dff_A_1771ZTwu0_0),.din(w_dff_A_miAybj3Y3_0),.clk(gclk));
	jdff dff_A_EZ2RwlKo8_0(.dout(w_dff_A_miAybj3Y3_0),.din(w_dff_A_EZ2RwlKo8_0),.clk(gclk));
	jdff dff_B_CbKVzz7k2_1(.din(n1389),.dout(w_dff_B_CbKVzz7k2_1),.clk(gclk));
	jdff dff_B_r7EWpylQ1_1(.din(w_dff_B_CbKVzz7k2_1),.dout(w_dff_B_r7EWpylQ1_1),.clk(gclk));
	jdff dff_A_yTm2tt4S6_1(.dout(w_G4091_1[1]),.din(w_dff_A_yTm2tt4S6_1),.clk(gclk));
	jdff dff_A_3oiJsFeB4_1(.dout(w_dff_A_yTm2tt4S6_1),.din(w_dff_A_3oiJsFeB4_1),.clk(gclk));
	jdff dff_A_yupCMjfw9_1(.dout(w_dff_A_3oiJsFeB4_1),.din(w_dff_A_yupCMjfw9_1),.clk(gclk));
	jdff dff_A_CUzQPcYa0_1(.dout(w_dff_A_yupCMjfw9_1),.din(w_dff_A_CUzQPcYa0_1),.clk(gclk));
	jdff dff_A_82YZAv663_1(.dout(w_dff_A_CUzQPcYa0_1),.din(w_dff_A_82YZAv663_1),.clk(gclk));
	jdff dff_A_GKwyiBR81_1(.dout(w_dff_A_82YZAv663_1),.din(w_dff_A_GKwyiBR81_1),.clk(gclk));
	jdff dff_A_nIvZjjzB4_1(.dout(w_dff_A_GKwyiBR81_1),.din(w_dff_A_nIvZjjzB4_1),.clk(gclk));
	jdff dff_A_2aYNoF4G8_1(.dout(w_dff_A_nIvZjjzB4_1),.din(w_dff_A_2aYNoF4G8_1),.clk(gclk));
	jdff dff_A_FUbKw7eB0_1(.dout(w_dff_A_2aYNoF4G8_1),.din(w_dff_A_FUbKw7eB0_1),.clk(gclk));
	jdff dff_A_UBRmLcbE0_1(.dout(w_dff_A_FUbKw7eB0_1),.din(w_dff_A_UBRmLcbE0_1),.clk(gclk));
	jdff dff_A_oXLwo3uF8_1(.dout(w_dff_A_UBRmLcbE0_1),.din(w_dff_A_oXLwo3uF8_1),.clk(gclk));
	jdff dff_A_y5ZDPO9D8_1(.dout(w_dff_A_oXLwo3uF8_1),.din(w_dff_A_y5ZDPO9D8_1),.clk(gclk));
	jdff dff_A_3fzlM4684_1(.dout(w_dff_A_y5ZDPO9D8_1),.din(w_dff_A_3fzlM4684_1),.clk(gclk));
	jdff dff_A_WZaGHca36_1(.dout(w_dff_A_3fzlM4684_1),.din(w_dff_A_WZaGHca36_1),.clk(gclk));
	jdff dff_A_FVXWl3FD7_1(.dout(w_dff_A_WZaGHca36_1),.din(w_dff_A_FVXWl3FD7_1),.clk(gclk));
	jdff dff_A_kjImmVOb9_1(.dout(w_dff_A_FVXWl3FD7_1),.din(w_dff_A_kjImmVOb9_1),.clk(gclk));
	jdff dff_A_6SFRLNe67_1(.dout(w_dff_A_kjImmVOb9_1),.din(w_dff_A_6SFRLNe67_1),.clk(gclk));
	jdff dff_A_hl1WHQlu0_1(.dout(w_dff_A_6SFRLNe67_1),.din(w_dff_A_hl1WHQlu0_1),.clk(gclk));
	jdff dff_A_D3C8o9HN8_2(.dout(w_G4091_1[2]),.din(w_dff_A_D3C8o9HN8_2),.clk(gclk));
	jdff dff_A_fYMbMDMp3_2(.dout(w_dff_A_D3C8o9HN8_2),.din(w_dff_A_fYMbMDMp3_2),.clk(gclk));
	jdff dff_A_BgaD9RHb7_2(.dout(w_dff_A_fYMbMDMp3_2),.din(w_dff_A_BgaD9RHb7_2),.clk(gclk));
	jdff dff_A_2p0oSSNB8_2(.dout(w_dff_A_BgaD9RHb7_2),.din(w_dff_A_2p0oSSNB8_2),.clk(gclk));
	jdff dff_A_0e6U2DBd6_2(.dout(w_dff_A_2p0oSSNB8_2),.din(w_dff_A_0e6U2DBd6_2),.clk(gclk));
	jdff dff_A_Xuznx5uz1_2(.dout(w_dff_A_0e6U2DBd6_2),.din(w_dff_A_Xuznx5uz1_2),.clk(gclk));
	jdff dff_A_rTU8kwPP7_2(.dout(w_dff_A_Xuznx5uz1_2),.din(w_dff_A_rTU8kwPP7_2),.clk(gclk));
	jdff dff_A_d4unRuEc8_2(.dout(w_dff_A_rTU8kwPP7_2),.din(w_dff_A_d4unRuEc8_2),.clk(gclk));
	jdff dff_A_Nia2hEuS7_2(.dout(w_dff_A_d4unRuEc8_2),.din(w_dff_A_Nia2hEuS7_2),.clk(gclk));
	jdff dff_A_Dcor2tS24_2(.dout(w_dff_A_Nia2hEuS7_2),.din(w_dff_A_Dcor2tS24_2),.clk(gclk));
	jdff dff_A_om3N0AQY7_0(.dout(w_n1383_0[0]),.din(w_dff_A_om3N0AQY7_0),.clk(gclk));
	jdff dff_A_sN4mtC7W7_0(.dout(w_dff_A_om3N0AQY7_0),.din(w_dff_A_sN4mtC7W7_0),.clk(gclk));
	jdff dff_B_PByhN64L5_1(.din(n1363),.dout(w_dff_B_PByhN64L5_1),.clk(gclk));
	jdff dff_B_sPMlff716_1(.din(w_dff_B_PByhN64L5_1),.dout(w_dff_B_sPMlff716_1),.clk(gclk));
	jdff dff_B_nHvIWuat9_1(.din(n1376),.dout(w_dff_B_nHvIWuat9_1),.clk(gclk));
	jdff dff_B_MPpmLCTT3_1(.din(n1377),.dout(w_dff_B_MPpmLCTT3_1),.clk(gclk));
	jdff dff_A_t9VyOwxo3_1(.dout(w_n426_0[1]),.din(w_dff_A_t9VyOwxo3_1),.clk(gclk));
	jdff dff_A_KI74boHH4_0(.dout(w_G503_1[0]),.din(w_dff_A_KI74boHH4_0),.clk(gclk));
	jdff dff_A_JLWgZOeG5_0(.dout(w_dff_A_KI74boHH4_0),.din(w_dff_A_JLWgZOeG5_0),.clk(gclk));
	jdff dff_A_Xge3qlDa3_0(.dout(w_dff_A_JLWgZOeG5_0),.din(w_dff_A_Xge3qlDa3_0),.clk(gclk));
	jdff dff_A_FFQSG4AZ9_0(.dout(w_dff_A_Xge3qlDa3_0),.din(w_dff_A_FFQSG4AZ9_0),.clk(gclk));
	jdff dff_A_R2qompgH1_1(.dout(w_G503_1[1]),.din(w_dff_A_R2qompgH1_1),.clk(gclk));
	jdff dff_A_5HmmIuF97_1(.dout(w_G503_0[1]),.din(w_dff_A_5HmmIuF97_1),.clk(gclk));
	jdff dff_A_84OCqbd11_1(.dout(w_dff_A_5HmmIuF97_1),.din(w_dff_A_84OCqbd11_1),.clk(gclk));
	jdff dff_A_vrlvvKg91_2(.dout(w_G503_0[2]),.din(w_dff_A_vrlvvKg91_2),.clk(gclk));
	jdff dff_A_5zYvxq7W2_2(.dout(w_dff_A_vrlvvKg91_2),.din(w_dff_A_5zYvxq7W2_2),.clk(gclk));
	jdff dff_A_LGtPvX8K8_2(.dout(w_dff_A_5zYvxq7W2_2),.din(w_dff_A_LGtPvX8K8_2),.clk(gclk));
	jdff dff_A_HyLyg6kX7_2(.dout(w_dff_A_LGtPvX8K8_2),.din(w_dff_A_HyLyg6kX7_2),.clk(gclk));
	jdff dff_A_f2Bes9Bs9_1(.dout(w_G324_1[1]),.din(w_dff_A_f2Bes9Bs9_1),.clk(gclk));
	jdff dff_A_X2o6mQP26_1(.dout(w_G324_0[1]),.din(w_dff_A_X2o6mQP26_1),.clk(gclk));
	jdff dff_B_pk6zXsK44_1(.din(n1368),.dout(w_dff_B_pk6zXsK44_1),.clk(gclk));
	jdff dff_B_QKm8l0wr0_1(.din(w_dff_B_pk6zXsK44_1),.dout(w_dff_B_QKm8l0wr0_1),.clk(gclk));
	jdff dff_A_a3hhoJix0_2(.dout(w_n388_0[2]),.din(w_dff_A_a3hhoJix0_2),.clk(gclk));
	jdff dff_B_yHrQBdqF8_3(.din(n388),.dout(w_dff_B_yHrQBdqF8_3),.clk(gclk));
	jdff dff_A_xzOc3OnQ6_0(.dout(w_G534_1[0]),.din(w_dff_A_xzOc3OnQ6_0),.clk(gclk));
	jdff dff_A_Bv3pi35O0_0(.dout(w_dff_A_xzOc3OnQ6_0),.din(w_dff_A_Bv3pi35O0_0),.clk(gclk));
	jdff dff_A_FFhWWLlg1_0(.dout(w_dff_A_Bv3pi35O0_0),.din(w_dff_A_FFhWWLlg1_0),.clk(gclk));
	jdff dff_A_DX0O2Syd8_1(.dout(w_G534_1[1]),.din(w_dff_A_DX0O2Syd8_1),.clk(gclk));
	jdff dff_B_LBOSmfTe1_1(.din(n1364),.dout(w_dff_B_LBOSmfTe1_1),.clk(gclk));
	jdff dff_A_HY2aFV2P3_1(.dout(w_G351_2[1]),.din(w_dff_A_HY2aFV2P3_1),.clk(gclk));
	jdff dff_A_ELM8S4fv3_1(.dout(w_G534_0[1]),.din(w_dff_A_ELM8S4fv3_1),.clk(gclk));
	jdff dff_A_vd4oStN78_1(.dout(w_dff_A_ELM8S4fv3_1),.din(w_dff_A_vd4oStN78_1),.clk(gclk));
	jdff dff_A_JjHqfE2P8_2(.dout(w_G534_0[2]),.din(w_dff_A_JjHqfE2P8_2),.clk(gclk));
	jdff dff_A_4gOKqh2V3_2(.dout(w_dff_A_JjHqfE2P8_2),.din(w_dff_A_4gOKqh2V3_2),.clk(gclk));
	jdff dff_A_ogSajMlJ4_2(.dout(w_dff_A_4gOKqh2V3_2),.din(w_dff_A_ogSajMlJ4_2),.clk(gclk));
	jdff dff_A_hXqnvGe07_0(.dout(w_G351_1[0]),.din(w_dff_A_hXqnvGe07_0),.clk(gclk));
	jdff dff_A_tVLIpjof3_2(.dout(w_n410_0[2]),.din(w_dff_A_tVLIpjof3_2),.clk(gclk));
	jdff dff_A_tg6NZPpn6_1(.dout(w_G514_0[1]),.din(w_dff_A_tg6NZPpn6_1),.clk(gclk));
	jdff dff_A_HajIFmL30_2(.dout(w_G514_0[2]),.din(w_dff_A_HajIFmL30_2),.clk(gclk));
	jdff dff_A_Z4IRXIZx4_2(.dout(w_dff_A_HajIFmL30_2),.din(w_dff_A_Z4IRXIZx4_2),.clk(gclk));
	jdff dff_A_2gyqCwep7_1(.dout(w_G361_0[1]),.din(w_dff_A_2gyqCwep7_1),.clk(gclk));
	jdff dff_B_Q9sxPbQ39_1(.din(n1354),.dout(w_dff_B_Q9sxPbQ39_1),.clk(gclk));
	jdff dff_B_Xn8RU2f01_1(.din(w_dff_B_Q9sxPbQ39_1),.dout(w_dff_B_Xn8RU2f01_1),.clk(gclk));
	jdff dff_B_hVArdk7n8_1(.din(n1355),.dout(w_dff_B_hVArdk7n8_1),.clk(gclk));
	jdff dff_B_mR1RJ9Tk9_1(.din(n378),.dout(w_dff_B_mR1RJ9Tk9_1),.clk(gclk));
	jdff dff_B_MzvEPU5s9_1(.din(n379),.dout(w_dff_B_MzvEPU5s9_1),.clk(gclk));
	jdff dff_A_A5X5yhsF9_0(.dout(w_G490_1[0]),.din(w_dff_A_A5X5yhsF9_0),.clk(gclk));
	jdff dff_A_v7GQKGqV5_0(.dout(w_dff_A_A5X5yhsF9_0),.din(w_dff_A_v7GQKGqV5_0),.clk(gclk));
	jdff dff_A_XRPK02d44_0(.dout(w_dff_A_v7GQKGqV5_0),.din(w_dff_A_XRPK02d44_0),.clk(gclk));
	jdff dff_A_p6vRd7Fz8_1(.dout(w_G490_1[1]),.din(w_dff_A_p6vRd7Fz8_1),.clk(gclk));
	jdff dff_A_nzThzmNM3_1(.dout(w_dff_A_p6vRd7Fz8_1),.din(w_dff_A_nzThzmNM3_1),.clk(gclk));
	jdff dff_A_VpsuK4DU7_1(.dout(w_G490_0[1]),.din(w_dff_A_VpsuK4DU7_1),.clk(gclk));
	jdff dff_A_KPhwFbOo5_1(.dout(w_dff_A_VpsuK4DU7_1),.din(w_dff_A_KPhwFbOo5_1),.clk(gclk));
	jdff dff_A_wQ07uUHs9_1(.dout(w_dff_A_KPhwFbOo5_1),.din(w_dff_A_wQ07uUHs9_1),.clk(gclk));
	jdff dff_A_5b5e9Wvx1_2(.dout(w_G490_0[2]),.din(w_dff_A_5b5e9Wvx1_2),.clk(gclk));
	jdff dff_A_x4tZzhZR6_2(.dout(w_dff_A_5b5e9Wvx1_2),.din(w_dff_A_x4tZzhZR6_2),.clk(gclk));
	jdff dff_A_OJtfwC613_2(.dout(w_dff_A_x4tZzhZR6_2),.din(w_dff_A_OJtfwC613_2),.clk(gclk));
	jdff dff_A_WRca75ot1_0(.dout(w_G316_1[0]),.din(w_dff_A_WRca75ot1_0),.clk(gclk));
	jdff dff_B_65tFn0Ix8_1(.din(n365),.dout(w_dff_B_65tFn0Ix8_1),.clk(gclk));
	jdff dff_B_eBibGzSN8_1(.din(n367),.dout(w_dff_B_eBibGzSN8_1),.clk(gclk));
	jdff dff_A_AO0pwfjq9_0(.dout(w_n362_0[0]),.din(w_dff_A_AO0pwfjq9_0),.clk(gclk));
	jdff dff_A_lWn202HJ2_0(.dout(w_dff_A_AO0pwfjq9_0),.din(w_dff_A_lWn202HJ2_0),.clk(gclk));
	jdff dff_A_E50FNLHQ9_0(.dout(w_dff_A_lWn202HJ2_0),.din(w_dff_A_E50FNLHQ9_0),.clk(gclk));
	jdff dff_A_5vLUvMLA7_0(.dout(w_G479_1[0]),.din(w_dff_A_5vLUvMLA7_0),.clk(gclk));
	jdff dff_A_38xu0fvJ7_0(.dout(w_dff_A_5vLUvMLA7_0),.din(w_dff_A_38xu0fvJ7_0),.clk(gclk));
	jdff dff_A_srWn93J30_1(.dout(w_G479_0[1]),.din(w_dff_A_srWn93J30_1),.clk(gclk));
	jdff dff_A_LUrWZIuz1_1(.dout(w_dff_A_srWn93J30_1),.din(w_dff_A_LUrWZIuz1_1),.clk(gclk));
	jdff dff_A_wvmDIRuM7_1(.dout(w_dff_A_LUrWZIuz1_1),.din(w_dff_A_wvmDIRuM7_1),.clk(gclk));
	jdff dff_A_QPWzXnZF4_2(.dout(w_G479_0[2]),.din(w_dff_A_QPWzXnZF4_2),.clk(gclk));
	jdff dff_A_3IDIkQpR3_2(.dout(w_dff_A_QPWzXnZF4_2),.din(w_dff_A_3IDIkQpR3_2),.clk(gclk));
	jdff dff_A_YYBiyCFM4_2(.dout(w_dff_A_3IDIkQpR3_2),.din(w_dff_A_YYBiyCFM4_2),.clk(gclk));
	jdff dff_A_Z06Ba6Xd8_0(.dout(w_G308_1[0]),.din(w_dff_A_Z06Ba6Xd8_0),.clk(gclk));
	jdff dff_A_FTOzRZ710_0(.dout(w_G302_0[0]),.din(w_dff_A_FTOzRZ710_0),.clk(gclk));
	jdff dff_A_5EZWNJ094_1(.dout(w_G302_0[1]),.din(w_dff_A_5EZWNJ094_1),.clk(gclk));
	jdff dff_A_tYEALtjI1_0(.dout(w_n401_0[0]),.din(w_dff_A_tYEALtjI1_0),.clk(gclk));
	jdff dff_A_55YIOMal5_2(.dout(w_n401_0[2]),.din(w_dff_A_55YIOMal5_2),.clk(gclk));
	jdff dff_A_ClLpTeIE1_1(.dout(w_G293_0[1]),.din(w_dff_A_ClLpTeIE1_1),.clk(gclk));
	jdff dff_B_ZC3lkNWB4_1(.din(n1349),.dout(w_dff_B_ZC3lkNWB4_1),.clk(gclk));
	jdff dff_B_G3JSTTyC0_1(.din(n1350),.dout(w_dff_B_G3JSTTyC0_1),.clk(gclk));
	jdff dff_A_ugTUNeBj5_0(.dout(w_n437_0[0]),.din(w_dff_A_ugTUNeBj5_0),.clk(gclk));
	jdff dff_A_hiWDEWT99_2(.dout(w_n437_0[2]),.din(w_dff_A_hiWDEWT99_2),.clk(gclk));
	jdff dff_A_UKFq0IAf2_2(.dout(w_dff_A_hiWDEWT99_2),.din(w_dff_A_UKFq0IAf2_2),.clk(gclk));
	jdff dff_A_7maiGc5N3_0(.dout(w_G523_1[0]),.din(w_dff_A_7maiGc5N3_0),.clk(gclk));
	jdff dff_A_sDHb6b4O3_1(.dout(w_G523_0[1]),.din(w_dff_A_sDHb6b4O3_1),.clk(gclk));
	jdff dff_A_R93ISZ5k6_1(.dout(w_dff_A_sDHb6b4O3_1),.din(w_dff_A_R93ISZ5k6_1),.clk(gclk));
	jdff dff_A_Jk1aUJmI7_1(.dout(w_dff_A_R93ISZ5k6_1),.din(w_dff_A_Jk1aUJmI7_1),.clk(gclk));
	jdff dff_A_6jMeSYC38_2(.dout(w_G523_0[2]),.din(w_dff_A_6jMeSYC38_2),.clk(gclk));
	jdff dff_A_7dGOx6od9_2(.dout(w_dff_A_6jMeSYC38_2),.din(w_dff_A_7dGOx6od9_2),.clk(gclk));
	jdff dff_A_YGYkLDhj5_1(.dout(w_G341_2[1]),.din(w_dff_A_YGYkLDhj5_1),.clk(gclk));
	jdff dff_A_YiyeAhCF0_2(.dout(w_G341_0[2]),.din(w_dff_A_YiyeAhCF0_2),.clk(gclk));
	jdff dff_A_9Oadu2nu0_2(.dout(w_n746_0[2]),.din(w_dff_A_9Oadu2nu0_2),.clk(gclk));
	jdff dff_A_9AB4Gv7c2_2(.dout(w_dff_A_9Oadu2nu0_2),.din(w_dff_A_9AB4Gv7c2_2),.clk(gclk));
	jdff dff_A_H74xHTCF5_2(.dout(w_dff_A_9AB4Gv7c2_2),.din(w_dff_A_H74xHTCF5_2),.clk(gclk));
	jdff dff_A_5GfGXW058_2(.dout(w_dff_A_H74xHTCF5_2),.din(w_dff_A_5GfGXW058_2),.clk(gclk));
	jdff dff_A_mqFVnjb22_2(.dout(w_dff_A_5GfGXW058_2),.din(w_dff_A_mqFVnjb22_2),.clk(gclk));
	jdff dff_A_dfRVq1zI3_2(.dout(w_dff_A_mqFVnjb22_2),.din(w_dff_A_dfRVq1zI3_2),.clk(gclk));
	jdff dff_A_ej7CPOa77_2(.dout(w_dff_A_dfRVq1zI3_2),.din(w_dff_A_ej7CPOa77_2),.clk(gclk));
	jdff dff_A_zipsQr5v1_2(.dout(w_dff_A_ej7CPOa77_2),.din(w_dff_A_zipsQr5v1_2),.clk(gclk));
	jdff dff_A_YM6urWMD0_2(.dout(w_dff_A_zipsQr5v1_2),.din(w_dff_A_YM6urWMD0_2),.clk(gclk));
	jdff dff_A_BDSPxLJq6_2(.dout(w_dff_A_YM6urWMD0_2),.din(w_dff_A_BDSPxLJq6_2),.clk(gclk));
	jdff dff_A_mTgfSlbB7_2(.dout(w_dff_A_BDSPxLJq6_2),.din(w_dff_A_mTgfSlbB7_2),.clk(gclk));
	jdff dff_A_7ggp5Ux39_0(.dout(w_n1002_1[0]),.din(w_dff_A_7ggp5Ux39_0),.clk(gclk));
	jdff dff_A_nnZXttfa8_0(.dout(w_dff_A_7ggp5Ux39_0),.din(w_dff_A_nnZXttfa8_0),.clk(gclk));
	jdff dff_A_0tyBVRu23_0(.dout(w_dff_A_nnZXttfa8_0),.din(w_dff_A_0tyBVRu23_0),.clk(gclk));
	jdff dff_A_CSjwxdJN3_0(.dout(w_dff_A_0tyBVRu23_0),.din(w_dff_A_CSjwxdJN3_0),.clk(gclk));
	jdff dff_A_D1dy12dg0_0(.dout(w_dff_A_CSjwxdJN3_0),.din(w_dff_A_D1dy12dg0_0),.clk(gclk));
	jdff dff_A_966KkFoe3_0(.dout(w_dff_A_D1dy12dg0_0),.din(w_dff_A_966KkFoe3_0),.clk(gclk));
	jdff dff_A_KW6NuIfj9_2(.dout(w_n1002_1[2]),.din(w_dff_A_KW6NuIfj9_2),.clk(gclk));
	jdff dff_A_nCKZH5oX1_2(.dout(w_dff_A_KW6NuIfj9_2),.din(w_dff_A_nCKZH5oX1_2),.clk(gclk));
	jdff dff_A_lT6JCe9K1_2(.dout(w_dff_A_nCKZH5oX1_2),.din(w_dff_A_lT6JCe9K1_2),.clk(gclk));
	jdff dff_A_QGWsjoSk8_2(.dout(w_dff_A_lT6JCe9K1_2),.din(w_dff_A_QGWsjoSk8_2),.clk(gclk));
	jdff dff_A_Q1kJlyPq1_2(.dout(w_dff_A_QGWsjoSk8_2),.din(w_dff_A_Q1kJlyPq1_2),.clk(gclk));
	jdff dff_A_O5b5TPBz6_2(.dout(w_dff_A_Q1kJlyPq1_2),.din(w_dff_A_O5b5TPBz6_2),.clk(gclk));
	jdff dff_A_zVpT7JMg6_2(.dout(w_dff_A_O5b5TPBz6_2),.din(w_dff_A_zVpT7JMg6_2),.clk(gclk));
	jdff dff_A_hvbSankV7_2(.dout(w_dff_A_zVpT7JMg6_2),.din(w_dff_A_hvbSankV7_2),.clk(gclk));
	jdff dff_A_ZMoQtbfK2_2(.dout(w_dff_A_hvbSankV7_2),.din(w_dff_A_ZMoQtbfK2_2),.clk(gclk));
	jdff dff_A_cjfNjDfN8_2(.dout(w_dff_A_ZMoQtbfK2_2),.din(w_dff_A_cjfNjDfN8_2),.clk(gclk));
	jdff dff_A_5M8zWWMe8_2(.dout(w_dff_A_cjfNjDfN8_2),.din(w_dff_A_5M8zWWMe8_2),.clk(gclk));
	jdff dff_A_rANZesdT1_2(.dout(w_dff_A_5M8zWWMe8_2),.din(w_dff_A_rANZesdT1_2),.clk(gclk));
	jdff dff_A_hYVvEH8k1_2(.dout(w_dff_A_rANZesdT1_2),.din(w_dff_A_hYVvEH8k1_2),.clk(gclk));
	jdff dff_A_DRiJzPKp3_2(.dout(w_dff_A_hYVvEH8k1_2),.din(w_dff_A_DRiJzPKp3_2),.clk(gclk));
	jdff dff_A_MzHK8kA45_2(.dout(w_dff_A_DRiJzPKp3_2),.din(w_dff_A_MzHK8kA45_2),.clk(gclk));
	jdff dff_A_ovlJJ6Mc1_2(.dout(w_dff_A_MzHK8kA45_2),.din(w_dff_A_ovlJJ6Mc1_2),.clk(gclk));
	jdff dff_A_Dfx2R6WO6_2(.dout(w_dff_A_ovlJJ6Mc1_2),.din(w_dff_A_Dfx2R6WO6_2),.clk(gclk));
	jdff dff_A_q93wqV3h6_2(.dout(w_dff_A_Dfx2R6WO6_2),.din(w_dff_A_q93wqV3h6_2),.clk(gclk));
	jdff dff_A_voDyk4lD2_1(.dout(w_n1002_0[1]),.din(w_dff_A_voDyk4lD2_1),.clk(gclk));
	jdff dff_A_cIlpqCWR9_1(.dout(w_dff_A_voDyk4lD2_1),.din(w_dff_A_cIlpqCWR9_1),.clk(gclk));
	jdff dff_A_RUOoy5O83_1(.dout(w_dff_A_cIlpqCWR9_1),.din(w_dff_A_RUOoy5O83_1),.clk(gclk));
	jdff dff_A_WdZ9Phl33_1(.dout(w_dff_A_RUOoy5O83_1),.din(w_dff_A_WdZ9Phl33_1),.clk(gclk));
	jdff dff_A_MIbnbtuL8_1(.dout(w_dff_A_WdZ9Phl33_1),.din(w_dff_A_MIbnbtuL8_1),.clk(gclk));
	jdff dff_A_AF624G4h9_1(.dout(w_dff_A_MIbnbtuL8_1),.din(w_dff_A_AF624G4h9_1),.clk(gclk));
	jdff dff_A_XrkqKJF24_1(.dout(w_dff_A_AF624G4h9_1),.din(w_dff_A_XrkqKJF24_1),.clk(gclk));
	jdff dff_A_yt3tsEhN3_1(.dout(w_dff_A_XrkqKJF24_1),.din(w_dff_A_yt3tsEhN3_1),.clk(gclk));
	jdff dff_A_xHk4giye6_1(.dout(w_dff_A_yt3tsEhN3_1),.din(w_dff_A_xHk4giye6_1),.clk(gclk));
	jdff dff_A_qSiXrfL87_1(.dout(w_dff_A_xHk4giye6_1),.din(w_dff_A_qSiXrfL87_1),.clk(gclk));
	jdff dff_A_tlpMJSzr4_1(.dout(w_dff_A_qSiXrfL87_1),.din(w_dff_A_tlpMJSzr4_1),.clk(gclk));
	jdff dff_A_RQnR9Z2z7_1(.dout(w_dff_A_tlpMJSzr4_1),.din(w_dff_A_RQnR9Z2z7_1),.clk(gclk));
	jdff dff_A_8NeluTTn1_1(.dout(w_dff_A_RQnR9Z2z7_1),.din(w_dff_A_8NeluTTn1_1),.clk(gclk));
	jdff dff_A_Bz2T7az03_1(.dout(w_dff_A_8NeluTTn1_1),.din(w_dff_A_Bz2T7az03_1),.clk(gclk));
	jdff dff_A_tPdzturL8_1(.dout(w_dff_A_Bz2T7az03_1),.din(w_dff_A_tPdzturL8_1),.clk(gclk));
	jdff dff_A_IJvihPOl2_1(.dout(w_dff_A_tPdzturL8_1),.din(w_dff_A_IJvihPOl2_1),.clk(gclk));
	jdff dff_A_RVqfX0ie3_2(.dout(w_n1002_0[2]),.din(w_dff_A_RVqfX0ie3_2),.clk(gclk));
	jdff dff_A_FRwjEamb9_2(.dout(w_dff_A_RVqfX0ie3_2),.din(w_dff_A_FRwjEamb9_2),.clk(gclk));
	jdff dff_A_MMUzKkQ14_2(.dout(w_dff_A_FRwjEamb9_2),.din(w_dff_A_MMUzKkQ14_2),.clk(gclk));
	jdff dff_A_xSw0jKL40_2(.dout(w_dff_A_MMUzKkQ14_2),.din(w_dff_A_xSw0jKL40_2),.clk(gclk));
	jdff dff_A_aC7ZYpJE6_2(.dout(w_dff_A_xSw0jKL40_2),.din(w_dff_A_aC7ZYpJE6_2),.clk(gclk));
	jdff dff_A_ZpM9mmJf0_2(.dout(w_dff_A_aC7ZYpJE6_2),.din(w_dff_A_ZpM9mmJf0_2),.clk(gclk));
	jdff dff_A_Qs8lUsEQ2_2(.dout(w_dff_A_ZpM9mmJf0_2),.din(w_dff_A_Qs8lUsEQ2_2),.clk(gclk));
	jdff dff_B_liGyRj4Q1_1(.din(n1641),.dout(w_dff_B_liGyRj4Q1_1),.clk(gclk));
	jdff dff_B_OJ5HfNRL9_1(.din(w_dff_B_liGyRj4Q1_1),.dout(w_dff_B_OJ5HfNRL9_1),.clk(gclk));
	jdff dff_B_0TEmTxzM6_1(.din(w_dff_B_OJ5HfNRL9_1),.dout(w_dff_B_0TEmTxzM6_1),.clk(gclk));
	jdff dff_B_0aP2VCWM6_1(.din(w_dff_B_0TEmTxzM6_1),.dout(w_dff_B_0aP2VCWM6_1),.clk(gclk));
	jdff dff_B_08P3VPFK4_1(.din(w_dff_B_0aP2VCWM6_1),.dout(w_dff_B_08P3VPFK4_1),.clk(gclk));
	jdff dff_B_omhSyZ459_1(.din(w_dff_B_08P3VPFK4_1),.dout(w_dff_B_omhSyZ459_1),.clk(gclk));
	jdff dff_B_jckNwaR91_1(.din(w_dff_B_omhSyZ459_1),.dout(w_dff_B_jckNwaR91_1),.clk(gclk));
	jdff dff_B_MLQIsMuH8_1(.din(w_dff_B_jckNwaR91_1),.dout(w_dff_B_MLQIsMuH8_1),.clk(gclk));
	jdff dff_B_7jWKwy5r6_1(.din(w_dff_B_MLQIsMuH8_1),.dout(w_dff_B_7jWKwy5r6_1),.clk(gclk));
	jdff dff_B_UE95Re2t4_1(.din(w_dff_B_7jWKwy5r6_1),.dout(w_dff_B_UE95Re2t4_1),.clk(gclk));
	jdff dff_B_ddPsgluX1_1(.din(w_dff_B_UE95Re2t4_1),.dout(w_dff_B_ddPsgluX1_1),.clk(gclk));
	jdff dff_B_M7gHhWNt2_1(.din(w_dff_B_ddPsgluX1_1),.dout(w_dff_B_M7gHhWNt2_1),.clk(gclk));
	jdff dff_B_1JIu4NRL5_1(.din(w_dff_B_M7gHhWNt2_1),.dout(w_dff_B_1JIu4NRL5_1),.clk(gclk));
	jdff dff_B_bkC1scp71_1(.din(w_dff_B_1JIu4NRL5_1),.dout(w_dff_B_bkC1scp71_1),.clk(gclk));
	jdff dff_B_lw3J3g0N6_1(.din(w_dff_B_bkC1scp71_1),.dout(w_dff_B_lw3J3g0N6_1),.clk(gclk));
	jdff dff_B_Vss8iiPJ5_1(.din(w_dff_B_lw3J3g0N6_1),.dout(w_dff_B_Vss8iiPJ5_1),.clk(gclk));
	jdff dff_B_65m2zDPh4_1(.din(w_dff_B_Vss8iiPJ5_1),.dout(w_dff_B_65m2zDPh4_1),.clk(gclk));
	jdff dff_B_FcdK7Hcj1_1(.din(w_dff_B_65m2zDPh4_1),.dout(w_dff_B_FcdK7Hcj1_1),.clk(gclk));
	jdff dff_B_pR7GSL0Y7_1(.din(w_dff_B_FcdK7Hcj1_1),.dout(w_dff_B_pR7GSL0Y7_1),.clk(gclk));
	jdff dff_B_e0zrZFup3_0(.din(n1600),.dout(w_dff_B_e0zrZFup3_0),.clk(gclk));
	jdff dff_B_6O7fnQNo2_0(.din(w_dff_B_e0zrZFup3_0),.dout(w_dff_B_6O7fnQNo2_0),.clk(gclk));
	jdff dff_B_zWB4DmA52_0(.din(w_dff_B_6O7fnQNo2_0),.dout(w_dff_B_zWB4DmA52_0),.clk(gclk));
	jdff dff_B_XBWlxRN51_0(.din(w_dff_B_zWB4DmA52_0),.dout(w_dff_B_XBWlxRN51_0),.clk(gclk));
	jdff dff_B_dl97fqRg4_0(.din(w_dff_B_XBWlxRN51_0),.dout(w_dff_B_dl97fqRg4_0),.clk(gclk));
	jdff dff_B_lSCZGfZS8_0(.din(w_dff_B_dl97fqRg4_0),.dout(w_dff_B_lSCZGfZS8_0),.clk(gclk));
	jdff dff_B_FolDlFxt7_0(.din(w_dff_B_lSCZGfZS8_0),.dout(w_dff_B_FolDlFxt7_0),.clk(gclk));
	jdff dff_B_ovF0zvai4_0(.din(w_dff_B_FolDlFxt7_0),.dout(w_dff_B_ovF0zvai4_0),.clk(gclk));
	jdff dff_B_FUwn0LRS8_0(.din(w_dff_B_ovF0zvai4_0),.dout(w_dff_B_FUwn0LRS8_0),.clk(gclk));
	jdff dff_B_7f94zMcT0_0(.din(w_dff_B_FUwn0LRS8_0),.dout(w_dff_B_7f94zMcT0_0),.clk(gclk));
	jdff dff_B_o3gIcTf50_0(.din(w_dff_B_7f94zMcT0_0),.dout(w_dff_B_o3gIcTf50_0),.clk(gclk));
	jdff dff_B_ipHBBiCP9_0(.din(w_dff_B_o3gIcTf50_0),.dout(w_dff_B_ipHBBiCP9_0),.clk(gclk));
	jdff dff_B_JYjRxzTa0_0(.din(w_dff_B_ipHBBiCP9_0),.dout(w_dff_B_JYjRxzTa0_0),.clk(gclk));
	jdff dff_B_2f0bdyTH6_0(.din(w_dff_B_JYjRxzTa0_0),.dout(w_dff_B_2f0bdyTH6_0),.clk(gclk));
	jdff dff_B_5qGAiS8O8_0(.din(w_dff_B_2f0bdyTH6_0),.dout(w_dff_B_5qGAiS8O8_0),.clk(gclk));
	jdff dff_B_K8rmROJK2_0(.din(w_dff_B_5qGAiS8O8_0),.dout(w_dff_B_K8rmROJK2_0),.clk(gclk));
	jdff dff_B_2huLCqb88_0(.din(w_dff_B_K8rmROJK2_0),.dout(w_dff_B_2huLCqb88_0),.clk(gclk));
	jdff dff_B_NPy4TpUC3_0(.din(w_dff_B_2huLCqb88_0),.dout(w_dff_B_NPy4TpUC3_0),.clk(gclk));
	jdff dff_B_Yrygy9EL4_0(.din(w_dff_B_NPy4TpUC3_0),.dout(w_dff_B_Yrygy9EL4_0),.clk(gclk));
	jdff dff_B_yCq0ZVJN9_1(.din(n1540),.dout(w_dff_B_yCq0ZVJN9_1),.clk(gclk));
	jdff dff_B_JbFcHKGO0_1(.din(w_dff_B_yCq0ZVJN9_1),.dout(w_dff_B_JbFcHKGO0_1),.clk(gclk));
	jdff dff_B_zuUBF6Gq3_1(.din(w_dff_B_JbFcHKGO0_1),.dout(w_dff_B_zuUBF6Gq3_1),.clk(gclk));
	jdff dff_B_WhspaehD7_1(.din(w_dff_B_zuUBF6Gq3_1),.dout(w_dff_B_WhspaehD7_1),.clk(gclk));
	jdff dff_B_B2x6Xiyd7_1(.din(w_dff_B_WhspaehD7_1),.dout(w_dff_B_B2x6Xiyd7_1),.clk(gclk));
	jdff dff_B_lEtp34gp1_1(.din(w_dff_B_B2x6Xiyd7_1),.dout(w_dff_B_lEtp34gp1_1),.clk(gclk));
	jdff dff_B_tYi7udAD2_1(.din(w_dff_B_lEtp34gp1_1),.dout(w_dff_B_tYi7udAD2_1),.clk(gclk));
	jdff dff_B_QcHQcyID4_1(.din(w_dff_B_tYi7udAD2_1),.dout(w_dff_B_QcHQcyID4_1),.clk(gclk));
	jdff dff_B_s4uYJj257_0(.din(n1589),.dout(w_dff_B_s4uYJj257_0),.clk(gclk));
	jdff dff_B_iCRNtnLO0_0(.din(w_dff_B_s4uYJj257_0),.dout(w_dff_B_iCRNtnLO0_0),.clk(gclk));
	jdff dff_B_EtojTeXx9_1(.din(n1579),.dout(w_dff_B_EtojTeXx9_1),.clk(gclk));
	jdff dff_B_ohrudmbV7_0(.din(n1586),.dout(w_dff_B_ohrudmbV7_0),.clk(gclk));
	jdff dff_B_XxUMWEiy2_0(.din(w_dff_B_ohrudmbV7_0),.dout(w_dff_B_XxUMWEiy2_0),.clk(gclk));
	jdff dff_B_aWwzQuXm1_0(.din(w_dff_B_XxUMWEiy2_0),.dout(w_dff_B_aWwzQuXm1_0),.clk(gclk));
	jdff dff_B_OZLQFGTU9_0(.din(n1584),.dout(w_dff_B_OZLQFGTU9_0),.clk(gclk));
	jdff dff_B_1ugzbJt42_1(.din(n1567),.dout(w_dff_B_1ugzbJt42_1),.clk(gclk));
	jdff dff_B_yhPL1mvI4_1(.din(w_dff_B_1ugzbJt42_1),.dout(w_dff_B_yhPL1mvI4_1),.clk(gclk));
	jdff dff_B_fiXlRQhm6_1(.din(w_dff_B_yhPL1mvI4_1),.dout(w_dff_B_fiXlRQhm6_1),.clk(gclk));
	jdff dff_B_U7FZVWcd5_1(.din(w_dff_B_fiXlRQhm6_1),.dout(w_dff_B_U7FZVWcd5_1),.clk(gclk));
	jdff dff_B_bxgfQRrM6_1(.din(w_dff_B_U7FZVWcd5_1),.dout(w_dff_B_bxgfQRrM6_1),.clk(gclk));
	jdff dff_B_SUWRyUAo3_1(.din(w_dff_B_bxgfQRrM6_1),.dout(w_dff_B_SUWRyUAo3_1),.clk(gclk));
	jdff dff_B_5PhlypIg2_1(.din(w_dff_B_SUWRyUAo3_1),.dout(w_dff_B_5PhlypIg2_1),.clk(gclk));
	jdff dff_B_rYGBZQAS1_1(.din(w_dff_B_5PhlypIg2_1),.dout(w_dff_B_rYGBZQAS1_1),.clk(gclk));
	jdff dff_B_9ndrnDAh8_1(.din(w_dff_B_rYGBZQAS1_1),.dout(w_dff_B_9ndrnDAh8_1),.clk(gclk));
	jdff dff_B_nnE2UKrf0_1(.din(w_dff_B_9ndrnDAh8_1),.dout(w_dff_B_nnE2UKrf0_1),.clk(gclk));
	jdff dff_B_xgf0Q80y2_1(.din(w_dff_B_nnE2UKrf0_1),.dout(w_dff_B_xgf0Q80y2_1),.clk(gclk));
	jdff dff_B_cMf6aa0h5_1(.din(w_dff_B_xgf0Q80y2_1),.dout(w_dff_B_cMf6aa0h5_1),.clk(gclk));
	jdff dff_B_KYhvU6y66_1(.din(w_dff_B_cMf6aa0h5_1),.dout(w_dff_B_KYhvU6y66_1),.clk(gclk));
	jdff dff_B_dTFJsWoQ6_1(.din(n1570),.dout(w_dff_B_dTFJsWoQ6_1),.clk(gclk));
	jdff dff_B_8wmzcDz37_1(.din(w_dff_B_dTFJsWoQ6_1),.dout(w_dff_B_8wmzcDz37_1),.clk(gclk));
	jdff dff_B_BY6gYS6B7_1(.din(w_dff_B_8wmzcDz37_1),.dout(w_dff_B_BY6gYS6B7_1),.clk(gclk));
	jdff dff_B_s14nKBMl3_1(.din(w_dff_B_BY6gYS6B7_1),.dout(w_dff_B_s14nKBMl3_1),.clk(gclk));
	jdff dff_B_Gq9c9ON17_1(.din(n1571),.dout(w_dff_B_Gq9c9ON17_1),.clk(gclk));
	jdff dff_B_ilc10LQn9_1(.din(w_dff_B_Gq9c9ON17_1),.dout(w_dff_B_ilc10LQn9_1),.clk(gclk));
	jdff dff_B_PpbW6kti0_1(.din(w_dff_B_ilc10LQn9_1),.dout(w_dff_B_PpbW6kti0_1),.clk(gclk));
	jdff dff_B_ECree2Cn4_1(.din(w_dff_B_PpbW6kti0_1),.dout(w_dff_B_ECree2Cn4_1),.clk(gclk));
	jdff dff_B_gi6eUhAL8_1(.din(w_dff_B_ECree2Cn4_1),.dout(w_dff_B_gi6eUhAL8_1),.clk(gclk));
	jdff dff_B_KctnXjBN9_1(.din(w_dff_B_gi6eUhAL8_1),.dout(w_dff_B_KctnXjBN9_1),.clk(gclk));
	jdff dff_A_XXL0aiQW4_0(.dout(w_n855_0[0]),.din(w_dff_A_XXL0aiQW4_0),.clk(gclk));
	jdff dff_A_an92ggBv9_1(.dout(w_n853_0[1]),.din(w_dff_A_an92ggBv9_1),.clk(gclk));
	jdff dff_B_swnD9oMO4_2(.din(n853),.dout(w_dff_B_swnD9oMO4_2),.clk(gclk));
	jdff dff_B_WUOsOuwl1_2(.din(w_dff_B_swnD9oMO4_2),.dout(w_dff_B_WUOsOuwl1_2),.clk(gclk));
	jdff dff_B_t5ysg7OS6_2(.din(w_dff_B_WUOsOuwl1_2),.dout(w_dff_B_t5ysg7OS6_2),.clk(gclk));
	jdff dff_B_P1SYit4Z8_2(.din(w_dff_B_t5ysg7OS6_2),.dout(w_dff_B_P1SYit4Z8_2),.clk(gclk));
	jdff dff_A_UFU9iMn87_0(.dout(w_n681_1[0]),.din(w_dff_A_UFU9iMn87_0),.clk(gclk));
	jdff dff_A_VBWCWI629_0(.dout(w_dff_A_UFU9iMn87_0),.din(w_dff_A_VBWCWI629_0),.clk(gclk));
	jdff dff_A_3QGKgOPX4_0(.dout(w_dff_A_VBWCWI629_0),.din(w_dff_A_3QGKgOPX4_0),.clk(gclk));
	jdff dff_A_5ZnwEata7_0(.dout(w_dff_A_3QGKgOPX4_0),.din(w_dff_A_5ZnwEata7_0),.clk(gclk));
	jdff dff_A_IznMhbn49_1(.dout(w_n681_1[1]),.din(w_dff_A_IznMhbn49_1),.clk(gclk));
	jdff dff_A_QBOcDrZP2_1(.dout(w_n1568_0[1]),.din(w_dff_A_QBOcDrZP2_1),.clk(gclk));
	jdff dff_B_yPRmIuMF4_1(.din(n1562),.dout(w_dff_B_yPRmIuMF4_1),.clk(gclk));
	jdff dff_B_bPw4S0de1_0(.din(n1563),.dout(w_dff_B_bPw4S0de1_0),.clk(gclk));
	jdff dff_B_tJK6alD19_1(.din(n1557),.dout(w_dff_B_tJK6alD19_1),.clk(gclk));
	jdff dff_A_TQPcLq8Y1_0(.dout(w_n1555_0[0]),.din(w_dff_A_TQPcLq8Y1_0),.clk(gclk));
	jdff dff_A_qVskqiBq8_0(.dout(w_dff_A_TQPcLq8Y1_0),.din(w_dff_A_qVskqiBq8_0),.clk(gclk));
	jdff dff_B_5mIHG5uh0_2(.din(n1553),.dout(w_dff_B_5mIHG5uh0_2),.clk(gclk));
	jdff dff_B_dTE99gFY9_2(.din(w_dff_B_5mIHG5uh0_2),.dout(w_dff_B_dTE99gFY9_2),.clk(gclk));
	jdff dff_B_M0lIgbye8_2(.din(w_dff_B_dTE99gFY9_2),.dout(w_dff_B_M0lIgbye8_2),.clk(gclk));
	jdff dff_B_g7CoFDCG5_2(.din(w_dff_B_M0lIgbye8_2),.dout(w_dff_B_g7CoFDCG5_2),.clk(gclk));
	jdff dff_B_i2ziskj46_2(.din(w_dff_B_g7CoFDCG5_2),.dout(w_dff_B_i2ziskj46_2),.clk(gclk));
	jdff dff_B_g7uquTPI9_2(.din(w_dff_B_i2ziskj46_2),.dout(w_dff_B_g7uquTPI9_2),.clk(gclk));
	jdff dff_B_szxuXp6g0_0(.din(n1551),.dout(w_dff_B_szxuXp6g0_0),.clk(gclk));
	jdff dff_B_Bv05TyMV1_0(.din(w_dff_B_szxuXp6g0_0),.dout(w_dff_B_Bv05TyMV1_0),.clk(gclk));
	jdff dff_B_znBonFDJ3_0(.din(w_dff_B_Bv05TyMV1_0),.dout(w_dff_B_znBonFDJ3_0),.clk(gclk));
	jdff dff_B_2MSOpb3o0_0(.din(n1550),.dout(w_dff_B_2MSOpb3o0_0),.clk(gclk));
	jdff dff_B_JzQBGI5E3_0(.din(w_dff_B_2MSOpb3o0_0),.dout(w_dff_B_JzQBGI5E3_0),.clk(gclk));
	jdff dff_B_M7YL1Mkh1_0(.din(w_dff_B_JzQBGI5E3_0),.dout(w_dff_B_M7YL1Mkh1_0),.clk(gclk));
	jdff dff_B_2CZqcMtj8_0(.din(w_dff_B_M7YL1Mkh1_0),.dout(w_dff_B_2CZqcMtj8_0),.clk(gclk));
	jdff dff_B_rbzmz5CZ9_0(.din(w_dff_B_2CZqcMtj8_0),.dout(w_dff_B_rbzmz5CZ9_0),.clk(gclk));
	jdff dff_A_6UUSTrVX6_2(.dout(w_n605_1[2]),.din(w_dff_A_6UUSTrVX6_2),.clk(gclk));
	jdff dff_A_3etelolD8_2(.dout(w_dff_A_6UUSTrVX6_2),.din(w_dff_A_3etelolD8_2),.clk(gclk));
	jdff dff_A_3caDZTan3_2(.dout(w_dff_A_3etelolD8_2),.din(w_dff_A_3caDZTan3_2),.clk(gclk));
	jdff dff_A_X1Meqaci4_2(.dout(w_dff_A_3caDZTan3_2),.din(w_dff_A_X1Meqaci4_2),.clk(gclk));
	jdff dff_A_KQupukqT0_2(.dout(w_dff_A_X1Meqaci4_2),.din(w_dff_A_KQupukqT0_2),.clk(gclk));
	jdff dff_A_uIv2YcRA2_2(.dout(w_dff_A_KQupukqT0_2),.din(w_dff_A_uIv2YcRA2_2),.clk(gclk));
	jdff dff_A_yybsGvv85_2(.dout(w_dff_A_uIv2YcRA2_2),.din(w_dff_A_yybsGvv85_2),.clk(gclk));
	jdff dff_A_xsWpch2G5_2(.dout(w_dff_A_yybsGvv85_2),.din(w_dff_A_xsWpch2G5_2),.clk(gclk));
	jdff dff_A_XWtA6UuR0_2(.dout(w_dff_A_xsWpch2G5_2),.din(w_dff_A_XWtA6UuR0_2),.clk(gclk));
	jdff dff_A_sfWyFTcT3_2(.dout(w_dff_A_XWtA6UuR0_2),.din(w_dff_A_sfWyFTcT3_2),.clk(gclk));
	jdff dff_A_JVPgjwDp8_2(.dout(w_dff_A_sfWyFTcT3_2),.din(w_dff_A_JVPgjwDp8_2),.clk(gclk));
	jdff dff_A_Aw2TO8zp6_2(.dout(w_dff_A_JVPgjwDp8_2),.din(w_dff_A_Aw2TO8zp6_2),.clk(gclk));
	jdff dff_A_eEZ6ClbX2_1(.dout(w_n944_0[1]),.din(w_dff_A_eEZ6ClbX2_1),.clk(gclk));
	jdff dff_A_vPpa6Jj87_1(.dout(w_dff_A_eEZ6ClbX2_1),.din(w_dff_A_vPpa6Jj87_1),.clk(gclk));
	jdff dff_A_ZpyLbyDc0_1(.dout(w_dff_A_vPpa6Jj87_1),.din(w_dff_A_ZpyLbyDc0_1),.clk(gclk));
	jdff dff_A_8kukiMfi7_1(.dout(w_dff_A_ZpyLbyDc0_1),.din(w_dff_A_8kukiMfi7_1),.clk(gclk));
	jdff dff_A_A497m73K3_1(.dout(w_dff_A_8kukiMfi7_1),.din(w_dff_A_A497m73K3_1),.clk(gclk));
	jdff dff_A_SbvhoUPS6_1(.dout(w_dff_A_A497m73K3_1),.din(w_dff_A_SbvhoUPS6_1),.clk(gclk));
	jdff dff_A_ZFnKkMIO5_1(.dout(w_dff_A_SbvhoUPS6_1),.din(w_dff_A_ZFnKkMIO5_1),.clk(gclk));
	jdff dff_A_Wf9am40F1_1(.dout(w_dff_A_ZFnKkMIO5_1),.din(w_dff_A_Wf9am40F1_1),.clk(gclk));
	jdff dff_A_QwGW2V7L3_1(.dout(w_dff_A_Wf9am40F1_1),.din(w_dff_A_QwGW2V7L3_1),.clk(gclk));
	jdff dff_A_wYlswrCS8_2(.dout(w_n930_0[2]),.din(w_dff_A_wYlswrCS8_2),.clk(gclk));
	jdff dff_A_51KeTvav3_2(.dout(w_dff_A_wYlswrCS8_2),.din(w_dff_A_51KeTvav3_2),.clk(gclk));
	jdff dff_A_Wp43asRs1_2(.dout(w_dff_A_51KeTvav3_2),.din(w_dff_A_Wp43asRs1_2),.clk(gclk));
	jdff dff_A_23vj8eKw1_2(.dout(w_dff_A_Wp43asRs1_2),.din(w_dff_A_23vj8eKw1_2),.clk(gclk));
	jdff dff_A_1i58seqN6_2(.dout(w_dff_A_23vj8eKw1_2),.din(w_dff_A_1i58seqN6_2),.clk(gclk));
	jdff dff_A_HkAEoIV02_2(.dout(w_dff_A_1i58seqN6_2),.din(w_dff_A_HkAEoIV02_2),.clk(gclk));
	jdff dff_A_tVodmN4C5_2(.dout(w_dff_A_HkAEoIV02_2),.din(w_dff_A_tVodmN4C5_2),.clk(gclk));
	jdff dff_A_iimUTs6z2_2(.dout(w_dff_A_tVodmN4C5_2),.din(w_dff_A_iimUTs6z2_2),.clk(gclk));
	jdff dff_A_knsfbCJo1_2(.dout(w_dff_A_iimUTs6z2_2),.din(w_dff_A_knsfbCJo1_2),.clk(gclk));
	jdff dff_B_JYxjRNqs6_3(.din(n930),.dout(w_dff_B_JYxjRNqs6_3),.clk(gclk));
	jdff dff_B_3ijbnRXv9_3(.din(w_dff_B_JYxjRNqs6_3),.dout(w_dff_B_3ijbnRXv9_3),.clk(gclk));
	jdff dff_A_Hy1lOvfA7_1(.dout(w_n700_0[1]),.din(w_dff_A_Hy1lOvfA7_1),.clk(gclk));
	jdff dff_A_AAFa1FuD2_1(.dout(w_dff_A_Hy1lOvfA7_1),.din(w_dff_A_AAFa1FuD2_1),.clk(gclk));
	jdff dff_A_PPHdl43q8_1(.dout(w_dff_A_AAFa1FuD2_1),.din(w_dff_A_PPHdl43q8_1),.clk(gclk));
	jdff dff_A_Lg42zLWs3_0(.dout(w_n706_0[0]),.din(w_dff_A_Lg42zLWs3_0),.clk(gclk));
	jdff dff_B_jWVFJh3J6_1(.din(n701),.dout(w_dff_B_jWVFJh3J6_1),.clk(gclk));
	jdff dff_B_fJkWUVKm7_1(.din(w_dff_B_jWVFJh3J6_1),.dout(w_dff_B_fJkWUVKm7_1),.clk(gclk));
	jdff dff_B_k5g8YeC02_0(.din(n599),.dout(w_dff_B_k5g8YeC02_0),.clk(gclk));
	jdff dff_B_XgANFRu84_1(.din(G233),.dout(w_dff_B_XgANFRu84_1),.clk(gclk));
	jdff dff_B_rsIdIZLY8_2(.din(n702),.dout(w_dff_B_rsIdIZLY8_2),.clk(gclk));
	jdff dff_A_qxb4VXKh9_0(.dout(w_n604_0[0]),.din(w_dff_A_qxb4VXKh9_0),.clk(gclk));
	jdff dff_B_rlpoLhJZ6_0(.din(n603),.dout(w_dff_B_rlpoLhJZ6_0),.clk(gclk));
	jdff dff_B_Od3WhJOn7_1(.din(G225),.dout(w_dff_B_Od3WhJOn7_1),.clk(gclk));
	jdff dff_A_3Xzr9Mok0_1(.dout(w_n928_0[1]),.din(w_dff_A_3Xzr9Mok0_1),.clk(gclk));
	jdff dff_A_COxX6Hug9_1(.dout(w_dff_A_3Xzr9Mok0_1),.din(w_dff_A_COxX6Hug9_1),.clk(gclk));
	jdff dff_A_H5f7fWQY6_1(.dout(w_dff_A_COxX6Hug9_1),.din(w_dff_A_H5f7fWQY6_1),.clk(gclk));
	jdff dff_A_Eq4TaIX45_1(.dout(w_dff_A_H5f7fWQY6_1),.din(w_dff_A_Eq4TaIX45_1),.clk(gclk));
	jdff dff_A_V3yLGFNH1_1(.dout(w_dff_A_Eq4TaIX45_1),.din(w_dff_A_V3yLGFNH1_1),.clk(gclk));
	jdff dff_A_ZkPL7UUL6_1(.dout(w_dff_A_V3yLGFNH1_1),.din(w_dff_A_ZkPL7UUL6_1),.clk(gclk));
	jdff dff_A_459UX8bo9_1(.dout(w_dff_A_ZkPL7UUL6_1),.din(w_dff_A_459UX8bo9_1),.clk(gclk));
	jdff dff_A_xUmdKPGb9_1(.dout(w_dff_A_459UX8bo9_1),.din(w_dff_A_xUmdKPGb9_1),.clk(gclk));
	jdff dff_A_G8ZG0IOT3_1(.dout(w_dff_A_xUmdKPGb9_1),.din(w_dff_A_G8ZG0IOT3_1),.clk(gclk));
	jdff dff_B_od7BNBhR9_2(.din(n928),.dout(w_dff_B_od7BNBhR9_2),.clk(gclk));
	jdff dff_B_dPTIeqpS1_2(.din(w_dff_B_od7BNBhR9_2),.dout(w_dff_B_dPTIeqpS1_2),.clk(gclk));
	jdff dff_B_r59SndGa8_2(.din(w_dff_B_dPTIeqpS1_2),.dout(w_dff_B_r59SndGa8_2),.clk(gclk));
	jdff dff_A_vyfh7V7W4_0(.dout(w_n596_0[0]),.din(w_dff_A_vyfh7V7W4_0),.clk(gclk));
	jdff dff_A_eBUFyfDL9_0(.dout(w_dff_A_vyfh7V7W4_0),.din(w_dff_A_eBUFyfDL9_0),.clk(gclk));
	jdff dff_A_7wscXeRN4_0(.dout(w_dff_A_eBUFyfDL9_0),.din(w_dff_A_7wscXeRN4_0),.clk(gclk));
	jdff dff_A_AutBRX7P6_0(.dout(w_dff_A_7wscXeRN4_0),.din(w_dff_A_AutBRX7P6_0),.clk(gclk));
	jdff dff_A_Hgu7Ljw35_0(.dout(w_dff_A_AutBRX7P6_0),.din(w_dff_A_Hgu7Ljw35_0),.clk(gclk));
	jdff dff_B_sQt5zr0P4_1(.din(n592),.dout(w_dff_B_sQt5zr0P4_1),.clk(gclk));
	jdff dff_B_VZOWUMFk6_1(.din(G209),.dout(w_dff_B_VZOWUMFk6_1),.clk(gclk));
	jdff dff_B_j6uxmmWU0_0(.din(n1544),.dout(w_dff_B_j6uxmmWU0_0),.clk(gclk));
	jdff dff_A_oyEdJAoc4_0(.dout(w_n585_0[0]),.din(w_dff_A_oyEdJAoc4_0),.clk(gclk));
	jdff dff_B_MrI0xqPx9_0(.din(n584),.dout(w_dff_B_MrI0xqPx9_0),.clk(gclk));
	jdff dff_B_CLDgGND10_0(.din(w_dff_B_MrI0xqPx9_0),.dout(w_dff_B_CLDgGND10_0),.clk(gclk));
	jdff dff_A_srezomRw5_0(.dout(w_n583_1[0]),.din(w_dff_A_srezomRw5_0),.clk(gclk));
	jdff dff_A_LnIAdAHM9_0(.dout(w_dff_A_srezomRw5_0),.din(w_dff_A_LnIAdAHM9_0),.clk(gclk));
	jdff dff_A_mTq4iD9w4_0(.dout(w_dff_A_LnIAdAHM9_0),.din(w_dff_A_mTq4iD9w4_0),.clk(gclk));
	jdff dff_A_B2mDDxTW7_0(.dout(w_n572_0[0]),.din(w_dff_A_B2mDDxTW7_0),.clk(gclk));
	jdff dff_A_claZv6Kr0_0(.dout(w_dff_A_B2mDDxTW7_0),.din(w_dff_A_claZv6Kr0_0),.clk(gclk));
	jdff dff_A_kAGnBtDr9_0(.dout(w_dff_A_claZv6Kr0_0),.din(w_dff_A_kAGnBtDr9_0),.clk(gclk));
	jdff dff_A_vOM2tzt18_0(.dout(w_dff_A_kAGnBtDr9_0),.din(w_dff_A_vOM2tzt18_0),.clk(gclk));
	jdff dff_A_T1e90f7s3_1(.dout(w_n567_1[1]),.din(w_dff_A_T1e90f7s3_1),.clk(gclk));
	jdff dff_A_r9gdVtro5_1(.dout(w_n567_0[1]),.din(w_dff_A_r9gdVtro5_1),.clk(gclk));
	jdff dff_A_Uk9XHvCw3_1(.dout(w_dff_A_r9gdVtro5_1),.din(w_dff_A_Uk9XHvCw3_1),.clk(gclk));
	jdff dff_A_aqXlXeOX2_1(.dout(w_dff_A_Uk9XHvCw3_1),.din(w_dff_A_aqXlXeOX2_1),.clk(gclk));
	jdff dff_A_Post4hJQ0_0(.dout(w_n497_1[0]),.din(w_dff_A_Post4hJQ0_0),.clk(gclk));
	jdff dff_A_67razSdm1_0(.dout(w_n562_0[0]),.din(w_dff_A_67razSdm1_0),.clk(gclk));
	jdff dff_A_ZUyMMdJq0_0(.dout(w_dff_A_67razSdm1_0),.din(w_dff_A_ZUyMMdJq0_0),.clk(gclk));
	jdff dff_A_pnldaA2v3_0(.dout(w_dff_A_ZUyMMdJq0_0),.din(w_dff_A_pnldaA2v3_0),.clk(gclk));
	jdff dff_A_hfuoI0jo8_0(.dout(w_dff_A_pnldaA2v3_0),.din(w_dff_A_hfuoI0jo8_0),.clk(gclk));
	jdff dff_A_uQZAZQvC3_0(.dout(w_dff_A_hfuoI0jo8_0),.din(w_dff_A_uQZAZQvC3_0),.clk(gclk));
	jdff dff_B_ussOJq4x6_2(.din(n562),.dout(w_dff_B_ussOJq4x6_2),.clk(gclk));
	jdff dff_B_Al0hJv4B7_2(.din(w_dff_B_ussOJq4x6_2),.dout(w_dff_B_Al0hJv4B7_2),.clk(gclk));
	jdff dff_A_im8jegML9_0(.dout(w_n561_0[0]),.din(w_dff_A_im8jegML9_0),.clk(gclk));
	jdff dff_A_CyFevzjJ5_1(.dout(w_n561_0[1]),.din(w_dff_A_CyFevzjJ5_1),.clk(gclk));
	jdff dff_A_BZcAxFcO4_1(.dout(w_dff_A_CyFevzjJ5_1),.din(w_dff_A_BZcAxFcO4_1),.clk(gclk));
	jdff dff_A_zoXmK7Iz9_1(.dout(w_dff_A_BZcAxFcO4_1),.din(w_dff_A_zoXmK7Iz9_1),.clk(gclk));
	jdff dff_A_nvPNabXU6_0(.dout(w_G1497_0[0]),.din(w_dff_A_nvPNabXU6_0),.clk(gclk));
	jdff dff_A_sGYejoD97_0(.dout(w_dff_A_nvPNabXU6_0),.din(w_dff_A_sGYejoD97_0),.clk(gclk));
	jdff dff_A_A30FOO4l2_0(.dout(w_dff_A_sGYejoD97_0),.din(w_dff_A_A30FOO4l2_0),.clk(gclk));
	jdff dff_A_mryewm2Q4_0(.dout(w_dff_A_A30FOO4l2_0),.din(w_dff_A_mryewm2Q4_0),.clk(gclk));
	jdff dff_A_8pyzMGoY5_0(.dout(w_dff_A_mryewm2Q4_0),.din(w_dff_A_8pyzMGoY5_0),.clk(gclk));
	jdff dff_A_NgA305G65_0(.dout(w_dff_A_8pyzMGoY5_0),.din(w_dff_A_NgA305G65_0),.clk(gclk));
	jdff dff_A_DB7W0JUv0_0(.dout(w_dff_A_NgA305G65_0),.din(w_dff_A_DB7W0JUv0_0),.clk(gclk));
	jdff dff_A_gPrNeSA64_0(.dout(w_dff_A_DB7W0JUv0_0),.din(w_dff_A_gPrNeSA64_0),.clk(gclk));
	jdff dff_A_nLKpNx1b7_0(.dout(w_dff_A_gPrNeSA64_0),.din(w_dff_A_nLKpNx1b7_0),.clk(gclk));
	jdff dff_A_atBJ4bHd9_0(.dout(w_dff_A_nLKpNx1b7_0),.din(w_dff_A_atBJ4bHd9_0),.clk(gclk));
	jdff dff_A_OTWRGP8Y7_0(.dout(w_dff_A_atBJ4bHd9_0),.din(w_dff_A_OTWRGP8Y7_0),.clk(gclk));
	jdff dff_A_YEIBHXyR5_0(.dout(w_dff_A_OTWRGP8Y7_0),.din(w_dff_A_YEIBHXyR5_0),.clk(gclk));
	jdff dff_A_XXcrqkgg2_2(.dout(w_G1497_0[2]),.din(w_dff_A_XXcrqkgg2_2),.clk(gclk));
	jdff dff_A_AHaBidWx0_2(.dout(w_dff_A_XXcrqkgg2_2),.din(w_dff_A_AHaBidWx0_2),.clk(gclk));
	jdff dff_A_m2xroV9f9_2(.dout(w_dff_A_AHaBidWx0_2),.din(w_dff_A_m2xroV9f9_2),.clk(gclk));
	jdff dff_A_NdBLsNQB4_2(.dout(w_dff_A_m2xroV9f9_2),.din(w_dff_A_NdBLsNQB4_2),.clk(gclk));
	jdff dff_A_YJvAUXfQ2_2(.dout(w_dff_A_NdBLsNQB4_2),.din(w_dff_A_YJvAUXfQ2_2),.clk(gclk));
	jdff dff_A_MG58C1ah5_2(.dout(w_dff_A_YJvAUXfQ2_2),.din(w_dff_A_MG58C1ah5_2),.clk(gclk));
	jdff dff_A_Jaq0R8y90_2(.dout(w_dff_A_MG58C1ah5_2),.din(w_dff_A_Jaq0R8y90_2),.clk(gclk));
	jdff dff_A_fqtU4tWr0_2(.dout(w_dff_A_Jaq0R8y90_2),.din(w_dff_A_fqtU4tWr0_2),.clk(gclk));
	jdff dff_A_JYsk3MQM5_2(.dout(w_dff_A_fqtU4tWr0_2),.din(w_dff_A_JYsk3MQM5_2),.clk(gclk));
	jdff dff_A_dHQDRExs4_2(.dout(w_dff_A_JYsk3MQM5_2),.din(w_dff_A_dHQDRExs4_2),.clk(gclk));
	jdff dff_B_VYjxetyZ9_1(.din(n675),.dout(w_dff_B_VYjxetyZ9_1),.clk(gclk));
	jdff dff_B_l5JERaAC2_1(.din(w_dff_B_VYjxetyZ9_1),.dout(w_dff_B_l5JERaAC2_1),.clk(gclk));
	jdff dff_B_DPpmcpte9_1(.din(w_dff_B_l5JERaAC2_1),.dout(w_dff_B_DPpmcpte9_1),.clk(gclk));
	jdff dff_B_DeBgD0QU3_1(.din(w_dff_B_DPpmcpte9_1),.dout(w_dff_B_DeBgD0QU3_1),.clk(gclk));
	jdff dff_B_6tPrnNlL0_1(.din(n676),.dout(w_dff_B_6tPrnNlL0_1),.clk(gclk));
	jdff dff_B_GAskT40k0_1(.din(w_dff_B_6tPrnNlL0_1),.dout(w_dff_B_GAskT40k0_1),.clk(gclk));
	jdff dff_B_Mr5vgPFN9_1(.din(w_dff_B_GAskT40k0_1),.dout(w_dff_B_Mr5vgPFN9_1),.clk(gclk));
	jdff dff_B_lJf389oy3_1(.din(w_dff_B_Mr5vgPFN9_1),.dout(w_dff_B_lJf389oy3_1),.clk(gclk));
	jdff dff_B_Db1QQsdW2_1(.din(w_dff_B_lJf389oy3_1),.dout(w_dff_B_Db1QQsdW2_1),.clk(gclk));
	jdff dff_A_8wQEgTCA2_1(.dout(w_n691_0[1]),.din(w_dff_A_8wQEgTCA2_1),.clk(gclk));
	jdff dff_A_UIiibPO25_0(.dout(w_n689_0[0]),.din(w_dff_A_UIiibPO25_0),.clk(gclk));
	jdff dff_A_geAXsMnP2_0(.dout(w_n687_0[0]),.din(w_dff_A_geAXsMnP2_0),.clk(gclk));
	jdff dff_A_JJrjz0nd1_1(.dout(w_n687_0[1]),.din(w_dff_A_JJrjz0nd1_1),.clk(gclk));
	jdff dff_A_YuoYuwoU9_1(.dout(w_dff_A_JJrjz0nd1_1),.din(w_dff_A_YuoYuwoU9_1),.clk(gclk));
	jdff dff_A_8a6PCgz73_1(.dout(w_dff_A_YuoYuwoU9_1),.din(w_dff_A_8a6PCgz73_1),.clk(gclk));
	jdff dff_A_DcXsmqnS8_1(.dout(w_dff_A_8a6PCgz73_1),.din(w_dff_A_DcXsmqnS8_1),.clk(gclk));
	jdff dff_A_C6bAeuK52_2(.dout(w_n571_0[2]),.din(w_dff_A_C6bAeuK52_2),.clk(gclk));
	jdff dff_A_omfJLI8Y4_2(.dout(w_dff_A_C6bAeuK52_2),.din(w_dff_A_omfJLI8Y4_2),.clk(gclk));
	jdff dff_A_xmhvvj0Z8_2(.dout(w_dff_A_omfJLI8Y4_2),.din(w_dff_A_xmhvvj0Z8_2),.clk(gclk));
	jdff dff_A_MsUDDw1v4_1(.dout(w_n569_0[1]),.din(w_dff_A_MsUDDw1v4_1),.clk(gclk));
	jdff dff_A_o9qhUCMZ1_1(.dout(w_G280_0[1]),.din(w_dff_A_o9qhUCMZ1_1),.clk(gclk));
	jdff dff_A_Iw5jiIn26_0(.dout(w_n486_1[0]),.din(w_dff_A_Iw5jiIn26_0),.clk(gclk));
	jdff dff_A_zfHbfcdg1_0(.dout(w_n681_2[0]),.din(w_dff_A_zfHbfcdg1_0),.clk(gclk));
	jdff dff_A_7EVxPVdw9_0(.dout(w_dff_A_zfHbfcdg1_0),.din(w_dff_A_7EVxPVdw9_0),.clk(gclk));
	jdff dff_A_gIyESD6S9_1(.dout(w_n680_0[1]),.din(w_dff_A_gIyESD6S9_1),.clk(gclk));
	jdff dff_B_JaGxgQWT2_2(.din(n680),.dout(w_dff_B_JaGxgQWT2_2),.clk(gclk));
	jdff dff_A_yGT0P50w9_0(.dout(w_n451_1[0]),.din(w_dff_A_yGT0P50w9_0),.clk(gclk));
	jdff dff_A_EgTalk5v9_1(.dout(w_n679_0[1]),.din(w_dff_A_EgTalk5v9_1),.clk(gclk));
	jdff dff_A_4qE7KPEQ0_1(.dout(w_dff_A_EgTalk5v9_1),.din(w_dff_A_4qE7KPEQ0_1),.clk(gclk));
	jdff dff_A_iH4CnHb29_1(.dout(w_n678_0[1]),.din(w_dff_A_iH4CnHb29_1),.clk(gclk));
	jdff dff_A_o6BsNIX50_1(.dout(w_dff_A_iH4CnHb29_1),.din(w_dff_A_o6BsNIX50_1),.clk(gclk));
	jdff dff_A_8N7eNG3U7_1(.dout(w_dff_A_o6BsNIX50_1),.din(w_dff_A_8N7eNG3U7_1),.clk(gclk));
	jdff dff_B_KJPtpKsx2_1(.din(n557),.dout(w_dff_B_KJPtpKsx2_1),.clk(gclk));
	jdff dff_B_KBAynGeM1_1(.din(G241),.dout(w_dff_B_KBAynGeM1_1),.clk(gclk));
	jdff dff_B_HPOgCEnt4_2(.din(n1543),.dout(w_dff_B_HPOgCEnt4_2),.clk(gclk));
	jdff dff_B_JXXNJSkA4_2(.din(w_dff_B_HPOgCEnt4_2),.dout(w_dff_B_JXXNJSkA4_2),.clk(gclk));
	jdff dff_B_KzH9yKB38_2(.din(w_dff_B_JXXNJSkA4_2),.dout(w_dff_B_KzH9yKB38_2),.clk(gclk));
	jdff dff_B_j90GPViM9_2(.din(w_dff_B_KzH9yKB38_2),.dout(w_dff_B_j90GPViM9_2),.clk(gclk));
	jdff dff_B_W5NYCNTJ1_2(.din(w_dff_B_j90GPViM9_2),.dout(w_dff_B_W5NYCNTJ1_2),.clk(gclk));
	jdff dff_B_xf1oSZ5z0_2(.din(w_dff_B_W5NYCNTJ1_2),.dout(w_dff_B_xf1oSZ5z0_2),.clk(gclk));
	jdff dff_B_pNYRD1394_2(.din(w_dff_B_xf1oSZ5z0_2),.dout(w_dff_B_pNYRD1394_2),.clk(gclk));
	jdff dff_B_oqpHiaKM8_2(.din(w_dff_B_pNYRD1394_2),.dout(w_dff_B_oqpHiaKM8_2),.clk(gclk));
	jdff dff_B_12Zklbrq1_2(.din(w_dff_B_oqpHiaKM8_2),.dout(w_dff_B_12Zklbrq1_2),.clk(gclk));
	jdff dff_B_ev8wgKxz4_2(.din(w_dff_B_12Zklbrq1_2),.dout(w_dff_B_ev8wgKxz4_2),.clk(gclk));
	jdff dff_A_Ts12P0AV9_2(.dout(w_n583_0[2]),.din(w_dff_A_Ts12P0AV9_2),.clk(gclk));
	jdff dff_A_0qwZDuaV1_2(.dout(w_dff_A_Ts12P0AV9_2),.din(w_dff_A_0qwZDuaV1_2),.clk(gclk));
	jdff dff_A_2dhCT1Wk4_2(.dout(w_dff_A_0qwZDuaV1_2),.din(w_dff_A_2dhCT1Wk4_2),.clk(gclk));
	jdff dff_A_5TKP5dxK2_2(.dout(w_dff_A_2dhCT1Wk4_2),.din(w_dff_A_5TKP5dxK2_2),.clk(gclk));
	jdff dff_A_crk6p3iG6_2(.dout(w_dff_A_5TKP5dxK2_2),.din(w_dff_A_crk6p3iG6_2),.clk(gclk));
	jdff dff_A_kd1v6NbK6_1(.dout(w_n578_0[1]),.din(w_dff_A_kd1v6NbK6_1),.clk(gclk));
	jdff dff_A_y0pz9t1g3_1(.dout(w_dff_A_kd1v6NbK6_1),.din(w_dff_A_y0pz9t1g3_1),.clk(gclk));
	jdff dff_A_8cro9meK8_1(.dout(w_dff_A_y0pz9t1g3_1),.din(w_dff_A_8cro9meK8_1),.clk(gclk));
	jdff dff_A_Rura2hEo7_1(.dout(w_dff_A_8cro9meK8_1),.din(w_dff_A_Rura2hEo7_1),.clk(gclk));
	jdff dff_A_2VGnmVt25_1(.dout(w_dff_A_Rura2hEo7_1),.din(w_dff_A_2VGnmVt25_1),.clk(gclk));
	jdff dff_A_JOdOdnOj3_1(.dout(w_dff_A_2VGnmVt25_1),.din(w_dff_A_JOdOdnOj3_1),.clk(gclk));
	jdff dff_A_FaJwG62n8_1(.dout(w_dff_A_JOdOdnOj3_1),.din(w_dff_A_FaJwG62n8_1),.clk(gclk));
	jdff dff_B_tbhq58vP9_0(.din(n576),.dout(w_dff_B_tbhq58vP9_0),.clk(gclk));
	jdff dff_A_D4JVfPTQ7_0(.dout(w_G335_3[0]),.din(w_dff_A_D4JVfPTQ7_0),.clk(gclk));
	jdff dff_B_LFNFrl5q5_1(.din(G264),.dout(w_dff_B_LFNFrl5q5_1),.clk(gclk));
	jdff dff_A_Nf3spo5L7_0(.dout(w_n473_1[0]),.din(w_dff_A_Nf3spo5L7_0),.clk(gclk));
	jdff dff_A_M1zNiXjj5_0(.dout(w_dff_A_Nf3spo5L7_0),.din(w_dff_A_M1zNiXjj5_0),.clk(gclk));
	jdff dff_A_5qs9epFC4_1(.dout(w_n473_1[1]),.din(w_dff_A_5qs9epFC4_1),.clk(gclk));
	jdff dff_A_9nVRPNt67_1(.dout(w_n943_0[1]),.din(w_dff_A_9nVRPNt67_1),.clk(gclk));
	jdff dff_A_pdR9RIH36_1(.dout(w_dff_A_9nVRPNt67_1),.din(w_dff_A_pdR9RIH36_1),.clk(gclk));
	jdff dff_A_by5yijvO9_1(.dout(w_dff_A_pdR9RIH36_1),.din(w_dff_A_by5yijvO9_1),.clk(gclk));
	jdff dff_A_bU9h8p941_1(.dout(w_dff_A_by5yijvO9_1),.din(w_dff_A_bU9h8p941_1),.clk(gclk));
	jdff dff_A_kbQ3KtJP4_1(.dout(w_dff_A_bU9h8p941_1),.din(w_dff_A_kbQ3KtJP4_1),.clk(gclk));
	jdff dff_A_et7Eq4Wx6_1(.dout(w_dff_A_kbQ3KtJP4_1),.din(w_dff_A_et7Eq4Wx6_1),.clk(gclk));
	jdff dff_A_IreSGpQ86_1(.dout(w_dff_A_et7Eq4Wx6_1),.din(w_dff_A_IreSGpQ86_1),.clk(gclk));
	jdff dff_A_PmNSlo4L5_1(.dout(w_dff_A_IreSGpQ86_1),.din(w_dff_A_PmNSlo4L5_1),.clk(gclk));
	jdff dff_A_waBRAppj0_1(.dout(w_dff_A_PmNSlo4L5_1),.din(w_dff_A_waBRAppj0_1),.clk(gclk));
	jdff dff_A_J9WXGZ522_1(.dout(w_dff_A_waBRAppj0_1),.din(w_dff_A_J9WXGZ522_1),.clk(gclk));
	jdff dff_A_dt1Fa41b3_1(.dout(w_dff_A_J9WXGZ522_1),.din(w_dff_A_dt1Fa41b3_1),.clk(gclk));
	jdff dff_A_WZBf4SCa2_1(.dout(w_dff_A_dt1Fa41b3_1),.din(w_dff_A_WZBf4SCa2_1),.clk(gclk));
	jdff dff_A_lDjO1o2S5_1(.dout(w_n591_0[1]),.din(w_dff_A_lDjO1o2S5_1),.clk(gclk));
	jdff dff_A_f8CAGVsM8_1(.dout(w_n590_0[1]),.din(w_dff_A_f8CAGVsM8_1),.clk(gclk));
	jdff dff_A_FWYweYQo4_1(.dout(w_dff_A_f8CAGVsM8_1),.din(w_dff_A_FWYweYQo4_1),.clk(gclk));
	jdff dff_B_uFZfeLal0_0(.din(n589),.dout(w_dff_B_uFZfeLal0_0),.clk(gclk));
	jdff dff_B_hfdQdMaW8_1(.din(G217),.dout(w_dff_B_hfdQdMaW8_1),.clk(gclk));
	jdff dff_A_dINxCVap4_0(.dout(w_G335_4[0]),.din(w_dff_A_dINxCVap4_0),.clk(gclk));
	jdff dff_A_z285s69A9_2(.dout(w_G335_1[2]),.din(w_dff_A_z285s69A9_2),.clk(gclk));
	jdff dff_A_I24ibmv85_1(.dout(w_n750_0[1]),.din(w_dff_A_I24ibmv85_1),.clk(gclk));
	jdff dff_A_yEZO1IIM9_1(.dout(w_dff_A_I24ibmv85_1),.din(w_dff_A_yEZO1IIM9_1),.clk(gclk));
	jdff dff_A_DGq2Bw4E3_1(.dout(w_dff_A_yEZO1IIM9_1),.din(w_dff_A_DGq2Bw4E3_1),.clk(gclk));
	jdff dff_A_p0aJPN2Z1_1(.dout(w_dff_A_DGq2Bw4E3_1),.din(w_dff_A_p0aJPN2Z1_1),.clk(gclk));
	jdff dff_A_36lCpSwf6_1(.dout(w_dff_A_p0aJPN2Z1_1),.din(w_dff_A_36lCpSwf6_1),.clk(gclk));
	jdff dff_A_4yC9fNkP6_1(.dout(w_dff_A_36lCpSwf6_1),.din(w_dff_A_4yC9fNkP6_1),.clk(gclk));
	jdff dff_A_hPcV7d4t9_1(.dout(w_dff_A_4yC9fNkP6_1),.din(w_dff_A_hPcV7d4t9_1),.clk(gclk));
	jdff dff_A_GpGtVjMW1_1(.dout(w_dff_A_hPcV7d4t9_1),.din(w_dff_A_GpGtVjMW1_1),.clk(gclk));
	jdff dff_A_WXAGokCV2_1(.dout(w_dff_A_GpGtVjMW1_1),.din(w_dff_A_WXAGokCV2_1),.clk(gclk));
	jdff dff_A_nPYokcY65_1(.dout(w_dff_A_WXAGokCV2_1),.din(w_dff_A_nPYokcY65_1),.clk(gclk));
	jdff dff_A_zZjDeUYC9_1(.dout(w_dff_A_nPYokcY65_1),.din(w_dff_A_zZjDeUYC9_1),.clk(gclk));
	jdff dff_A_PSuEwDMR0_1(.dout(w_dff_A_zZjDeUYC9_1),.din(w_dff_A_PSuEwDMR0_1),.clk(gclk));
	jdff dff_A_4pP9wztx5_1(.dout(w_dff_A_PSuEwDMR0_1),.din(w_dff_A_4pP9wztx5_1),.clk(gclk));
	jdff dff_A_qDVqyDDb1_1(.dout(w_dff_A_4pP9wztx5_1),.din(w_dff_A_qDVqyDDb1_1),.clk(gclk));
	jdff dff_A_jTz3AAI64_1(.dout(w_dff_A_qDVqyDDb1_1),.din(w_dff_A_jTz3AAI64_1),.clk(gclk));
	jdff dff_A_7x98A8be8_1(.dout(w_dff_A_jTz3AAI64_1),.din(w_dff_A_7x98A8be8_1),.clk(gclk));
	jdff dff_A_PqAu7HDC8_1(.dout(w_dff_A_7x98A8be8_1),.din(w_dff_A_PqAu7HDC8_1),.clk(gclk));
	jdff dff_A_pJHP8ukH6_2(.dout(w_n750_0[2]),.din(w_dff_A_pJHP8ukH6_2),.clk(gclk));
	jdff dff_A_cElaUkoG5_2(.dout(w_dff_A_pJHP8ukH6_2),.din(w_dff_A_cElaUkoG5_2),.clk(gclk));
	jdff dff_A_9KbYkFrg0_2(.dout(w_dff_A_cElaUkoG5_2),.din(w_dff_A_9KbYkFrg0_2),.clk(gclk));
	jdff dff_A_W9O4aZ8K8_2(.dout(w_dff_A_9KbYkFrg0_2),.din(w_dff_A_W9O4aZ8K8_2),.clk(gclk));
	jdff dff_A_vqtsjzzj7_2(.dout(w_dff_A_W9O4aZ8K8_2),.din(w_dff_A_vqtsjzzj7_2),.clk(gclk));
	jdff dff_A_dAwaBqhc0_2(.dout(w_dff_A_vqtsjzzj7_2),.din(w_dff_A_dAwaBqhc0_2),.clk(gclk));
	jdff dff_A_MGXlMyfQ4_2(.dout(w_dff_A_dAwaBqhc0_2),.din(w_dff_A_MGXlMyfQ4_2),.clk(gclk));
	jdff dff_A_7VL5Q9WW4_2(.dout(w_dff_A_MGXlMyfQ4_2),.din(w_dff_A_7VL5Q9WW4_2),.clk(gclk));
	jdff dff_A_AAaitIOj4_2(.dout(w_G4091_2[2]),.din(w_dff_A_AAaitIOj4_2),.clk(gclk));
	jdff dff_A_Yc6PNerJ2_2(.dout(w_G4091_0[2]),.din(w_dff_A_Yc6PNerJ2_2),.clk(gclk));
	jdff dff_A_4nFkwIba8_2(.dout(w_dff_A_Yc6PNerJ2_2),.din(w_dff_A_4nFkwIba8_2),.clk(gclk));
	jdff dff_A_4C3HrD6y1_2(.dout(w_dff_A_4nFkwIba8_2),.din(w_dff_A_4C3HrD6y1_2),.clk(gclk));
	jdff dff_A_Z7fQ9pbj9_2(.dout(w_dff_A_4C3HrD6y1_2),.din(w_dff_A_Z7fQ9pbj9_2),.clk(gclk));
	jdff dff_A_ijIv27JT2_2(.dout(w_dff_A_Z7fQ9pbj9_2),.din(w_dff_A_ijIv27JT2_2),.clk(gclk));
	jdff dff_A_kksTxhOK8_2(.dout(w_dff_A_ijIv27JT2_2),.din(w_dff_A_kksTxhOK8_2),.clk(gclk));
	jdff dff_A_2SGXp0oM2_2(.dout(w_dff_A_kksTxhOK8_2),.din(w_dff_A_2SGXp0oM2_2),.clk(gclk));
	jdff dff_A_4HolBZtJ9_2(.dout(w_dff_A_2SGXp0oM2_2),.din(w_dff_A_4HolBZtJ9_2),.clk(gclk));
	jdff dff_A_edmQBWUx8_2(.dout(w_dff_A_4HolBZtJ9_2),.din(w_dff_A_edmQBWUx8_2),.clk(gclk));
	jdff dff_A_QhwQfpfa2_2(.dout(w_dff_A_edmQBWUx8_2),.din(w_dff_A_QhwQfpfa2_2),.clk(gclk));
	jdff dff_A_677S7Hut9_2(.dout(w_dff_A_QhwQfpfa2_2),.din(w_dff_A_677S7Hut9_2),.clk(gclk));
	jdff dff_A_6cJ6o5721_2(.dout(w_dff_A_677S7Hut9_2),.din(w_dff_A_6cJ6o5721_2),.clk(gclk));
	jdff dff_A_273yAYLc6_2(.dout(w_dff_A_6cJ6o5721_2),.din(w_dff_A_273yAYLc6_2),.clk(gclk));
	jdff dff_A_DUGoD5AN0_2(.dout(w_dff_A_273yAYLc6_2),.din(w_dff_A_DUGoD5AN0_2),.clk(gclk));
	jdff dff_A_xPdKTMWM8_2(.dout(w_dff_A_DUGoD5AN0_2),.din(w_dff_A_xPdKTMWM8_2),.clk(gclk));
	jdff dff_A_pqofm7Rs6_2(.dout(w_dff_A_xPdKTMWM8_2),.din(w_dff_A_pqofm7Rs6_2),.clk(gclk));
	jdff dff_A_5s3u3bZC2_2(.dout(w_dff_A_pqofm7Rs6_2),.din(w_dff_A_5s3u3bZC2_2),.clk(gclk));
	jdff dff_A_p7lWIDlr6_2(.dout(w_dff_A_5s3u3bZC2_2),.din(w_dff_A_p7lWIDlr6_2),.clk(gclk));
	jdff dff_B_8CK6fxJ17_2(.din(n1533),.dout(w_dff_B_8CK6fxJ17_2),.clk(gclk));
	jdff dff_B_ICVIfdOc7_1(.din(n1526),.dout(w_dff_B_ICVIfdOc7_1),.clk(gclk));
	jdff dff_B_wUIvTA2e6_1(.din(n1527),.dout(w_dff_B_wUIvTA2e6_1),.clk(gclk));
	jdff dff_A_MVXiMlLm6_0(.dout(w_n486_0[0]),.din(w_dff_A_MVXiMlLm6_0),.clk(gclk));
	jdff dff_A_2vz3W4HZ9_2(.dout(w_n486_0[2]),.din(w_dff_A_2vz3W4HZ9_2),.clk(gclk));
	jdff dff_A_B8oHIgWy0_2(.dout(w_dff_A_2vz3W4HZ9_2),.din(w_dff_A_B8oHIgWy0_2),.clk(gclk));
	jdff dff_A_THdHVtNs4_0(.dout(w_G411_0[0]),.din(w_dff_A_THdHVtNs4_0),.clk(gclk));
	jdff dff_A_lp8KMlFN7_0(.dout(w_dff_A_THdHVtNs4_0),.din(w_dff_A_lp8KMlFN7_0),.clk(gclk));
	jdff dff_A_jOqVUj9t0_1(.dout(w_G411_0[1]),.din(w_dff_A_jOqVUj9t0_1),.clk(gclk));
	jdff dff_A_CgprWX050_1(.dout(w_G273_2[1]),.din(w_dff_A_CgprWX050_1),.clk(gclk));
	jdff dff_A_NUBUx68D1_2(.dout(w_G273_0[2]),.din(w_dff_A_NUBUx68D1_2),.clk(gclk));
	jdff dff_B_er0lYqO62_1(.din(n1518),.dout(w_dff_B_er0lYqO62_1),.clk(gclk));
	jdff dff_B_OicV9Q9v5_1(.din(w_dff_B_er0lYqO62_1),.dout(w_dff_B_OicV9Q9v5_1),.clk(gclk));
	jdff dff_A_EGI21scW8_2(.dout(w_n473_0[2]),.din(w_dff_A_EGI21scW8_2),.clk(gclk));
	jdff dff_A_4959dTQj2_2(.dout(w_dff_A_EGI21scW8_2),.din(w_dff_A_4959dTQj2_2),.clk(gclk));
	jdff dff_B_cNjfOzIY2_3(.din(n473),.dout(w_dff_B_cNjfOzIY2_3),.clk(gclk));
	jdff dff_B_10meFRAC4_1(.din(n1514),.dout(w_dff_B_10meFRAC4_1),.clk(gclk));
	jdff dff_A_xKkvtONz0_1(.dout(w_G257_2[1]),.din(w_dff_A_xKkvtONz0_1),.clk(gclk));
	jdff dff_A_VTAY7AXp1_0(.dout(w_G389_0[0]),.din(w_dff_A_VTAY7AXp1_0),.clk(gclk));
	jdff dff_A_deWhamyq0_0(.dout(w_dff_A_VTAY7AXp1_0),.din(w_dff_A_deWhamyq0_0),.clk(gclk));
	jdff dff_A_bdsLIN204_1(.dout(w_G389_0[1]),.din(w_dff_A_bdsLIN204_1),.clk(gclk));
	jdff dff_A_bANAr1uV7_0(.dout(w_G257_1[0]),.din(w_dff_A_bANAr1uV7_0),.clk(gclk));
	jdff dff_B_cCsAviXl1_1(.din(n1507),.dout(w_dff_B_cCsAviXl1_1),.clk(gclk));
	jdff dff_B_NJxDURGC2_1(.din(n1508),.dout(w_dff_B_NJxDURGC2_1),.clk(gclk));
	jdff dff_A_gVE6PJP04_0(.dout(w_n451_0[0]),.din(w_dff_A_gVE6PJP04_0),.clk(gclk));
	jdff dff_A_cyAvUDdr7_2(.dout(w_n451_0[2]),.din(w_dff_A_cyAvUDdr7_2),.clk(gclk));
	jdff dff_A_E1z9zFPw6_2(.dout(w_dff_A_cyAvUDdr7_2),.din(w_dff_A_E1z9zFPw6_2),.clk(gclk));
	jdff dff_A_MVwIv0GP9_0(.dout(w_G400_1[0]),.din(w_dff_A_MVwIv0GP9_0),.clk(gclk));
	jdff dff_A_UwK3clxq8_1(.dout(w_G400_0[1]),.din(w_dff_A_UwK3clxq8_1),.clk(gclk));
	jdff dff_A_9GNBrGGm0_1(.dout(w_dff_A_UwK3clxq8_1),.din(w_dff_A_9GNBrGGm0_1),.clk(gclk));
	jdff dff_A_MBcWebB95_2(.dout(w_G400_0[2]),.din(w_dff_A_MBcWebB95_2),.clk(gclk));
	jdff dff_A_DefNt8va7_2(.dout(w_dff_A_MBcWebB95_2),.din(w_dff_A_DefNt8va7_2),.clk(gclk));
	jdff dff_A_cF42Pl3q4_2(.dout(w_dff_A_DefNt8va7_2),.din(w_dff_A_cF42Pl3q4_2),.clk(gclk));
	jdff dff_A_a10Qzhlk4_0(.dout(w_G265_2[0]),.din(w_dff_A_a10Qzhlk4_0),.clk(gclk));
	jdff dff_A_CWikI4PP6_2(.dout(w_G265_0[2]),.din(w_dff_A_CWikI4PP6_2),.clk(gclk));
	jdff dff_B_GixM5bZd1_1(.din(n1498),.dout(w_dff_B_GixM5bZd1_1),.clk(gclk));
	jdff dff_B_SAipD6aa6_1(.din(n1499),.dout(w_dff_B_SAipD6aa6_1),.clk(gclk));
	jdff dff_A_t8GskBuY4_0(.dout(w_n497_0[0]),.din(w_dff_A_t8GskBuY4_0),.clk(gclk));
	jdff dff_A_n8hXXRMk4_2(.dout(w_n497_0[2]),.din(w_dff_A_n8hXXRMk4_2),.clk(gclk));
	jdff dff_A_BgIz9GOx3_2(.dout(w_dff_A_n8hXXRMk4_2),.din(w_dff_A_BgIz9GOx3_2),.clk(gclk));
	jdff dff_A_0MVFq6Xk6_0(.dout(w_G374_0[0]),.din(w_dff_A_0MVFq6Xk6_0),.clk(gclk));
	jdff dff_A_EA789TRI2_0(.dout(w_dff_A_0MVFq6Xk6_0),.din(w_dff_A_EA789TRI2_0),.clk(gclk));
	jdff dff_A_iAcg0cnm8_1(.dout(w_G374_0[1]),.din(w_dff_A_iAcg0cnm8_1),.clk(gclk));
	jdff dff_A_AAuUKy352_0(.dout(w_G281_2[0]),.din(w_dff_A_AAuUKy352_0),.clk(gclk));
	jdff dff_A_3ZfCYEqE6_2(.dout(w_G281_0[2]),.din(w_dff_A_3ZfCYEqE6_2),.clk(gclk));
	jdff dff_B_DBmktnb60_1(.din(n1463),.dout(w_dff_B_DBmktnb60_1),.clk(gclk));
	jdff dff_B_TxKrL9ni2_1(.din(w_dff_B_DBmktnb60_1),.dout(w_dff_B_TxKrL9ni2_1),.clk(gclk));
	jdff dff_B_xxXRhAoH8_1(.din(n1486),.dout(w_dff_B_xxXRhAoH8_1),.clk(gclk));
	jdff dff_B_0aMwDOAT0_1(.din(n1487),.dout(w_dff_B_0aMwDOAT0_1),.clk(gclk));
	jdff dff_A_IV5zb80V7_1(.dout(w_G210_1[1]),.din(w_dff_A_IV5zb80V7_1),.clk(gclk));
	jdff dff_A_SCGFeEfB8_1(.dout(w_n543_0[1]),.din(w_dff_A_SCGFeEfB8_1),.clk(gclk));
	jdff dff_A_73sXI6kO5_0(.dout(w_G457_2[0]),.din(w_dff_A_73sXI6kO5_0),.clk(gclk));
	jdff dff_A_AePJaZQz2_0(.dout(w_G457_0[0]),.din(w_dff_A_AePJaZQz2_0),.clk(gclk));
	jdff dff_A_Xc6ft2vN3_0(.dout(w_dff_A_AePJaZQz2_0),.din(w_dff_A_Xc6ft2vN3_0),.clk(gclk));
	jdff dff_A_Jut5NXeM6_0(.dout(w_dff_A_Xc6ft2vN3_0),.din(w_dff_A_Jut5NXeM6_0),.clk(gclk));
	jdff dff_A_fejT3bwL7_2(.dout(w_G457_0[2]),.din(w_dff_A_fejT3bwL7_2),.clk(gclk));
	jdff dff_A_xZYFZW7P3_2(.dout(w_dff_A_fejT3bwL7_2),.din(w_dff_A_xZYFZW7P3_2),.clk(gclk));
	jdff dff_A_0Pys0NPO7_1(.dout(w_G210_2[1]),.din(w_dff_A_0Pys0NPO7_1),.clk(gclk));
	jdff dff_A_BgefP6GH8_2(.dout(w_G210_0[2]),.din(w_dff_A_BgefP6GH8_2),.clk(gclk));
	jdff dff_B_yoonln1B9_1(.din(n1478),.dout(w_dff_B_yoonln1B9_1),.clk(gclk));
	jdff dff_B_kkKjk15J7_1(.din(w_dff_B_yoonln1B9_1),.dout(w_dff_B_kkKjk15J7_1),.clk(gclk));
	jdff dff_B_Jr6O50Gx2_2(.din(n509),.dout(w_dff_B_Jr6O50Gx2_2),.clk(gclk));
	jdff dff_A_y3avN7Kb8_0(.dout(w_G468_1[0]),.din(w_dff_A_y3avN7Kb8_0),.clk(gclk));
	jdff dff_A_6yDkhFjs5_0(.dout(w_dff_A_y3avN7Kb8_0),.din(w_dff_A_6yDkhFjs5_0),.clk(gclk));
	jdff dff_A_3uU7QwdY8_0(.dout(w_dff_A_6yDkhFjs5_0),.din(w_dff_A_3uU7QwdY8_0),.clk(gclk));
	jdff dff_A_UkQVmX7O7_1(.dout(w_G468_1[1]),.din(w_dff_A_UkQVmX7O7_1),.clk(gclk));
	jdff dff_B_QPKBkYa50_1(.din(n1474),.dout(w_dff_B_QPKBkYa50_1),.clk(gclk));
	jdff dff_A_dhGTwRnI9_1(.dout(w_G218_2[1]),.din(w_dff_A_dhGTwRnI9_1),.clk(gclk));
	jdff dff_A_vPjgPKnP4_1(.dout(w_G468_0[1]),.din(w_dff_A_vPjgPKnP4_1),.clk(gclk));
	jdff dff_A_2Rm7Aary5_1(.dout(w_dff_A_vPjgPKnP4_1),.din(w_dff_A_2Rm7Aary5_1),.clk(gclk));
	jdff dff_A_IyTfIq1V5_2(.dout(w_G468_0[2]),.din(w_dff_A_IyTfIq1V5_2),.clk(gclk));
	jdff dff_A_pIPAGnXt1_2(.dout(w_dff_A_IyTfIq1V5_2),.din(w_dff_A_pIPAGnXt1_2),.clk(gclk));
	jdff dff_A_YXV3NzWV7_2(.dout(w_dff_A_pIPAGnXt1_2),.din(w_dff_A_YXV3NzWV7_2),.clk(gclk));
	jdff dff_A_nXUQGQHM8_0(.dout(w_G218_1[0]),.din(w_dff_A_nXUQGQHM8_0),.clk(gclk));
	jdff dff_B_gjMBR40Q7_1(.din(n1468),.dout(w_dff_B_gjMBR40Q7_1),.clk(gclk));
	jdff dff_B_A8uZyRAU6_1(.din(w_dff_B_gjMBR40Q7_1),.dout(w_dff_B_A8uZyRAU6_1),.clk(gclk));
	jdff dff_B_3kpYIH2t1_2(.din(n532),.dout(w_dff_B_3kpYIH2t1_2),.clk(gclk));
	jdff dff_A_yRJKABJA7_0(.dout(w_G422_2[0]),.din(w_dff_A_yRJKABJA7_0),.clk(gclk));
	jdff dff_B_Tu4nLu7q1_1(.din(n1464),.dout(w_dff_B_Tu4nLu7q1_1),.clk(gclk));
	jdff dff_A_kG5zjPzZ4_1(.dout(w_G226_2[1]),.din(w_dff_A_kG5zjPzZ4_1),.clk(gclk));
	jdff dff_A_NhkLcVSS1_0(.dout(w_G422_0[0]),.din(w_dff_A_NhkLcVSS1_0),.clk(gclk));
	jdff dff_A_kFFPNKen1_0(.dout(w_dff_A_NhkLcVSS1_0),.din(w_dff_A_kFFPNKen1_0),.clk(gclk));
	jdff dff_A_J4a6OJl35_0(.dout(w_dff_A_kFFPNKen1_0),.din(w_dff_A_J4a6OJl35_0),.clk(gclk));
	jdff dff_A_fI3DVBQl6_2(.dout(w_G422_0[2]),.din(w_dff_A_fI3DVBQl6_2),.clk(gclk));
	jdff dff_A_LuvEiM885_2(.dout(w_dff_A_fI3DVBQl6_2),.din(w_dff_A_LuvEiM885_2),.clk(gclk));
	jdff dff_A_OUwJ3ss06_1(.dout(w_G251_4[1]),.din(w_dff_A_OUwJ3ss06_1),.clk(gclk));
	jdff dff_A_JLvkYXd86_2(.dout(w_G251_4[2]),.din(w_dff_A_JLvkYXd86_2),.clk(gclk));
	jdff dff_A_FE7aTk4H4_1(.dout(w_G251_1[1]),.din(w_dff_A_FE7aTk4H4_1),.clk(gclk));
	jdff dff_A_5yJTXELi2_2(.dout(w_G251_1[2]),.din(w_dff_A_5yJTXELi2_2),.clk(gclk));
	jdff dff_A_OpqiR3Vc2_0(.dout(w_G226_1[0]),.din(w_dff_A_OpqiR3Vc2_0),.clk(gclk));
	jdff dff_B_DM8NHtC44_1(.din(n523),.dout(w_dff_B_DM8NHtC44_1),.clk(gclk));
	jdff dff_B_ERk43COR3_1(.din(n524),.dout(w_dff_B_ERk43COR3_1),.clk(gclk));
	jdff dff_A_csDIYLrv1_0(.dout(w_G446_1[0]),.din(w_dff_A_csDIYLrv1_0),.clk(gclk));
	jdff dff_A_V4NBYffl6_0(.dout(w_dff_A_csDIYLrv1_0),.din(w_dff_A_V4NBYffl6_0),.clk(gclk));
	jdff dff_A_uwAD3Z5m5_0(.dout(w_dff_A_V4NBYffl6_0),.din(w_dff_A_uwAD3Z5m5_0),.clk(gclk));
	jdff dff_A_bbab6R4y3_0(.dout(w_dff_A_uwAD3Z5m5_0),.din(w_dff_A_bbab6R4y3_0),.clk(gclk));
	jdff dff_A_Zv5HTxQ87_1(.dout(w_G446_1[1]),.din(w_dff_A_Zv5HTxQ87_1),.clk(gclk));
	jdff dff_A_hEVKOsBS8_1(.dout(w_dff_A_Zv5HTxQ87_1),.din(w_dff_A_hEVKOsBS8_1),.clk(gclk));
	jdff dff_A_CI9viVWJ3_1(.dout(w_G446_0[1]),.din(w_dff_A_CI9viVWJ3_1),.clk(gclk));
	jdff dff_A_jGnHbOL21_1(.dout(w_dff_A_CI9viVWJ3_1),.din(w_dff_A_jGnHbOL21_1),.clk(gclk));
	jdff dff_A_l4IzvBjI0_1(.dout(w_dff_A_jGnHbOL21_1),.din(w_dff_A_l4IzvBjI0_1),.clk(gclk));
	jdff dff_A_89vNui0Q7_1(.dout(w_dff_A_l4IzvBjI0_1),.din(w_dff_A_89vNui0Q7_1),.clk(gclk));
	jdff dff_A_W4AvdWoO1_2(.dout(w_G446_0[2]),.din(w_dff_A_W4AvdWoO1_2),.clk(gclk));
	jdff dff_A_TE3jcuxM9_2(.dout(w_dff_A_W4AvdWoO1_2),.din(w_dff_A_TE3jcuxM9_2),.clk(gclk));
	jdff dff_A_Ys9Fg2av1_2(.dout(w_dff_A_TE3jcuxM9_2),.din(w_dff_A_Ys9Fg2av1_2),.clk(gclk));
	jdff dff_A_I0myafGa7_2(.dout(w_dff_A_Ys9Fg2av1_2),.din(w_dff_A_I0myafGa7_2),.clk(gclk));
	jdff dff_A_eMdGojBb4_0(.dout(w_G206_0[0]),.din(w_dff_A_eMdGojBb4_0),.clk(gclk));
	jdff dff_B_ts6ctaUK2_1(.din(n1458),.dout(w_dff_B_ts6ctaUK2_1),.clk(gclk));
	jdff dff_B_XmZ1eiIF8_1(.din(n1459),.dout(w_dff_B_XmZ1eiIF8_1),.clk(gclk));
	jdff dff_A_1cbmMLvm9_0(.dout(w_G242_1[0]),.din(w_dff_A_1cbmMLvm9_0),.clk(gclk));
	jdff dff_A_iYvooa9B2_1(.dout(w_G242_1[1]),.din(w_dff_A_iYvooa9B2_1),.clk(gclk));
	jdff dff_A_NOh48NUa9_1(.dout(w_G242_0[1]),.din(w_dff_A_NOh48NUa9_1),.clk(gclk));
	jdff dff_A_o2DKDKw12_2(.dout(w_G242_0[2]),.din(w_dff_A_o2DKDKw12_2),.clk(gclk));
	jdff dff_A_i7B6QyWf9_2(.dout(w_G248_3[2]),.din(w_dff_A_i7B6QyWf9_2),.clk(gclk));
	jdff dff_A_zw1S1KHt6_1(.dout(w_n462_0[1]),.din(w_dff_A_zw1S1KHt6_1),.clk(gclk));
	jdff dff_A_3ks3UEbD4_1(.dout(w_dff_A_zw1S1KHt6_1),.din(w_dff_A_3ks3UEbD4_1),.clk(gclk));
	jdff dff_A_qpkDTumY8_1(.dout(w_dff_A_3ks3UEbD4_1),.din(w_dff_A_qpkDTumY8_1),.clk(gclk));
	jdff dff_A_wrTCqjNx6_1(.dout(w_dff_A_qpkDTumY8_1),.din(w_dff_A_wrTCqjNx6_1),.clk(gclk));
	jdff dff_A_Kn1bkS712_2(.dout(w_n462_0[2]),.din(w_dff_A_Kn1bkS712_2),.clk(gclk));
	jdff dff_A_iq7LmbY75_0(.dout(w_G435_1[0]),.din(w_dff_A_iq7LmbY75_0),.clk(gclk));
	jdff dff_A_s8E2cyjG5_0(.dout(w_dff_A_iq7LmbY75_0),.din(w_dff_A_s8E2cyjG5_0),.clk(gclk));
	jdff dff_A_jouJrXEr8_0(.dout(w_dff_A_s8E2cyjG5_0),.din(w_dff_A_jouJrXEr8_0),.clk(gclk));
	jdff dff_A_veECLmaf3_0(.dout(w_dff_A_jouJrXEr8_0),.din(w_dff_A_veECLmaf3_0),.clk(gclk));
	jdff dff_A_SBOE7Fke9_1(.dout(w_G435_1[1]),.din(w_dff_A_SBOE7Fke9_1),.clk(gclk));
	jdff dff_A_3V0Vm0B15_1(.dout(w_G435_0[1]),.din(w_dff_A_3V0Vm0B15_1),.clk(gclk));
	jdff dff_A_8bvJuRvx0_1(.dout(w_dff_A_3V0Vm0B15_1),.din(w_dff_A_8bvJuRvx0_1),.clk(gclk));
	jdff dff_A_LHiAelBe1_2(.dout(w_G435_0[2]),.din(w_dff_A_LHiAelBe1_2),.clk(gclk));
	jdff dff_A_sD1utwgA9_2(.dout(w_dff_A_LHiAelBe1_2),.din(w_dff_A_sD1utwgA9_2),.clk(gclk));
	jdff dff_A_w2R1iwmP6_2(.dout(w_dff_A_sD1utwgA9_2),.din(w_dff_A_w2R1iwmP6_2),.clk(gclk));
	jdff dff_A_tGhJKCd82_2(.dout(w_dff_A_w2R1iwmP6_2),.din(w_dff_A_tGhJKCd82_2),.clk(gclk));
	jdff dff_A_qJLIzwhg0_1(.dout(w_G251_0[1]),.din(w_dff_A_qJLIzwhg0_1),.clk(gclk));
	jdff dff_A_w4RxTup30_2(.dout(w_G251_0[2]),.din(w_dff_A_w4RxTup30_2),.clk(gclk));
	jdff dff_A_s2t4eMkx3_0(.dout(w_G234_2[0]),.din(w_dff_A_s2t4eMkx3_0),.clk(gclk));
	jdff dff_A_q9w38W3Z5_2(.dout(w_G234_0[2]),.din(w_dff_A_q9w38W3Z5_2),.clk(gclk));
	jdff dff_A_SssbdDsk4_0(.dout(w_G4092_1[0]),.din(w_dff_A_SssbdDsk4_0),.clk(gclk));
	jdff dff_A_UtUx6igc9_0(.dout(w_dff_A_SssbdDsk4_0),.din(w_dff_A_UtUx6igc9_0),.clk(gclk));
	jdff dff_A_RudJcVFx6_0(.dout(w_dff_A_UtUx6igc9_0),.din(w_dff_A_RudJcVFx6_0),.clk(gclk));
	jdff dff_A_mH82zFvq4_0(.dout(w_dff_A_RudJcVFx6_0),.din(w_dff_A_mH82zFvq4_0),.clk(gclk));
	jdff dff_A_MT1G3OY36_0(.dout(w_dff_A_mH82zFvq4_0),.din(w_dff_A_MT1G3OY36_0),.clk(gclk));
	jdff dff_A_GQbrbEcQ3_0(.dout(w_dff_A_MT1G3OY36_0),.din(w_dff_A_GQbrbEcQ3_0),.clk(gclk));
	jdff dff_A_Vil1QuFM0_0(.dout(w_dff_A_GQbrbEcQ3_0),.din(w_dff_A_Vil1QuFM0_0),.clk(gclk));
	jdff dff_A_Bx9SpO2Z4_0(.dout(w_dff_A_Vil1QuFM0_0),.din(w_dff_A_Bx9SpO2Z4_0),.clk(gclk));
	jdff dff_A_fGb21stF5_0(.dout(w_dff_A_Bx9SpO2Z4_0),.din(w_dff_A_fGb21stF5_0),.clk(gclk));
	jdff dff_A_UFHV60qe1_0(.dout(w_dff_A_fGb21stF5_0),.din(w_dff_A_UFHV60qe1_0),.clk(gclk));
	jdff dff_A_HioiWyno7_0(.dout(w_dff_A_UFHV60qe1_0),.din(w_dff_A_HioiWyno7_0),.clk(gclk));
	jdff dff_A_tiqr3PDH6_1(.dout(w_G4092_1[1]),.din(w_dff_A_tiqr3PDH6_1),.clk(gclk));
	jdff dff_A_aCo5Gh4Y6_0(.dout(w_n999_1[0]),.din(w_dff_A_aCo5Gh4Y6_0),.clk(gclk));
	jdff dff_A_MsqheXaF3_0(.dout(w_dff_A_aCo5Gh4Y6_0),.din(w_dff_A_MsqheXaF3_0),.clk(gclk));
	jdff dff_A_hXX5za0E7_0(.dout(w_dff_A_MsqheXaF3_0),.din(w_dff_A_hXX5za0E7_0),.clk(gclk));
	jdff dff_A_VJssQblt5_0(.dout(w_dff_A_hXX5za0E7_0),.din(w_dff_A_VJssQblt5_0),.clk(gclk));
	jdff dff_A_ARmYp1xD2_0(.dout(w_dff_A_VJssQblt5_0),.din(w_dff_A_ARmYp1xD2_0),.clk(gclk));
	jdff dff_A_kqWYIkrs0_0(.dout(w_dff_A_ARmYp1xD2_0),.din(w_dff_A_kqWYIkrs0_0),.clk(gclk));
	jdff dff_A_i8oAcA1P3_0(.dout(w_dff_A_kqWYIkrs0_0),.din(w_dff_A_i8oAcA1P3_0),.clk(gclk));
	jdff dff_A_nW5w3hZ52_2(.dout(w_n999_1[2]),.din(w_dff_A_nW5w3hZ52_2),.clk(gclk));
	jdff dff_A_Hry0ZRis6_2(.dout(w_dff_A_nW5w3hZ52_2),.din(w_dff_A_Hry0ZRis6_2),.clk(gclk));
	jdff dff_A_yTLYQhWh3_2(.dout(w_dff_A_Hry0ZRis6_2),.din(w_dff_A_yTLYQhWh3_2),.clk(gclk));
	jdff dff_A_sfrbuVF69_2(.dout(w_dff_A_yTLYQhWh3_2),.din(w_dff_A_sfrbuVF69_2),.clk(gclk));
	jdff dff_A_dGpCHngu8_2(.dout(w_dff_A_sfrbuVF69_2),.din(w_dff_A_dGpCHngu8_2),.clk(gclk));
	jdff dff_A_P2nNnnMx7_2(.dout(w_dff_A_dGpCHngu8_2),.din(w_dff_A_P2nNnnMx7_2),.clk(gclk));
	jdff dff_A_3ySoJ11v1_2(.dout(w_dff_A_P2nNnnMx7_2),.din(w_dff_A_3ySoJ11v1_2),.clk(gclk));
	jdff dff_A_fRvdGumS9_2(.dout(w_dff_A_3ySoJ11v1_2),.din(w_dff_A_fRvdGumS9_2),.clk(gclk));
	jdff dff_A_mRQKqnyj6_2(.dout(w_dff_A_fRvdGumS9_2),.din(w_dff_A_mRQKqnyj6_2),.clk(gclk));
	jdff dff_A_wVpZ0ypX9_2(.dout(w_dff_A_mRQKqnyj6_2),.din(w_dff_A_wVpZ0ypX9_2),.clk(gclk));
	jdff dff_A_yG9WEfH69_2(.dout(w_dff_A_wVpZ0ypX9_2),.din(w_dff_A_yG9WEfH69_2),.clk(gclk));
	jdff dff_A_WeqxlSju4_2(.dout(w_dff_A_yG9WEfH69_2),.din(w_dff_A_WeqxlSju4_2),.clk(gclk));
	jdff dff_A_v5LyskgL4_2(.dout(w_dff_A_WeqxlSju4_2),.din(w_dff_A_v5LyskgL4_2),.clk(gclk));
	jdff dff_A_JA6O6dTh1_2(.dout(w_dff_A_v5LyskgL4_2),.din(w_dff_A_JA6O6dTh1_2),.clk(gclk));
	jdff dff_A_sTG3Glzy5_2(.dout(w_dff_A_JA6O6dTh1_2),.din(w_dff_A_sTG3Glzy5_2),.clk(gclk));
	jdff dff_A_GjC3orH78_2(.dout(w_dff_A_sTG3Glzy5_2),.din(w_dff_A_GjC3orH78_2),.clk(gclk));
	jdff dff_A_vnnaMtET6_2(.dout(w_dff_A_GjC3orH78_2),.din(w_dff_A_vnnaMtET6_2),.clk(gclk));
	jdff dff_A_0C7rssIX6_2(.dout(w_dff_A_vnnaMtET6_2),.din(w_dff_A_0C7rssIX6_2),.clk(gclk));
	jdff dff_A_x1eHhxId0_2(.dout(w_dff_A_0C7rssIX6_2),.din(w_dff_A_x1eHhxId0_2),.clk(gclk));
	jdff dff_A_ZtLGQnYV7_1(.dout(w_n999_0[1]),.din(w_dff_A_ZtLGQnYV7_1),.clk(gclk));
	jdff dff_A_ZvDFzrbu4_1(.dout(w_dff_A_ZtLGQnYV7_1),.din(w_dff_A_ZvDFzrbu4_1),.clk(gclk));
	jdff dff_A_wiZYGcvl5_1(.dout(w_dff_A_ZvDFzrbu4_1),.din(w_dff_A_wiZYGcvl5_1),.clk(gclk));
	jdff dff_A_QU304iMb2_1(.dout(w_dff_A_wiZYGcvl5_1),.din(w_dff_A_QU304iMb2_1),.clk(gclk));
	jdff dff_A_BQyx0Emi5_1(.dout(w_dff_A_QU304iMb2_1),.din(w_dff_A_BQyx0Emi5_1),.clk(gclk));
	jdff dff_A_UoNcJO6G7_1(.dout(w_dff_A_BQyx0Emi5_1),.din(w_dff_A_UoNcJO6G7_1),.clk(gclk));
	jdff dff_A_Cybi2LeB9_1(.dout(w_dff_A_UoNcJO6G7_1),.din(w_dff_A_Cybi2LeB9_1),.clk(gclk));
	jdff dff_A_RoEvyOu82_1(.dout(w_dff_A_Cybi2LeB9_1),.din(w_dff_A_RoEvyOu82_1),.clk(gclk));
	jdff dff_A_5k0j8sKn3_1(.dout(w_dff_A_RoEvyOu82_1),.din(w_dff_A_5k0j8sKn3_1),.clk(gclk));
	jdff dff_A_gUTMHAdq3_1(.dout(w_dff_A_5k0j8sKn3_1),.din(w_dff_A_gUTMHAdq3_1),.clk(gclk));
	jdff dff_A_yoOkNbya8_1(.dout(w_dff_A_gUTMHAdq3_1),.din(w_dff_A_yoOkNbya8_1),.clk(gclk));
	jdff dff_A_9fe40RVz0_1(.dout(w_dff_A_yoOkNbya8_1),.din(w_dff_A_9fe40RVz0_1),.clk(gclk));
	jdff dff_A_zanh6Atf6_1(.dout(w_dff_A_9fe40RVz0_1),.din(w_dff_A_zanh6Atf6_1),.clk(gclk));
	jdff dff_A_c0KHvXL23_1(.dout(w_dff_A_zanh6Atf6_1),.din(w_dff_A_c0KHvXL23_1),.clk(gclk));
	jdff dff_A_L2YAXgQa0_1(.dout(w_dff_A_c0KHvXL23_1),.din(w_dff_A_L2YAXgQa0_1),.clk(gclk));
	jdff dff_A_rLVuhbm90_1(.dout(w_dff_A_L2YAXgQa0_1),.din(w_dff_A_rLVuhbm90_1),.clk(gclk));
	jdff dff_A_3K6GrN4X4_1(.dout(w_dff_A_rLVuhbm90_1),.din(w_dff_A_3K6GrN4X4_1),.clk(gclk));
	jdff dff_A_iI4S3sc08_2(.dout(w_n999_0[2]),.din(w_dff_A_iI4S3sc08_2),.clk(gclk));
	jdff dff_A_1cobA0TI7_2(.dout(w_dff_A_iI4S3sc08_2),.din(w_dff_A_1cobA0TI7_2),.clk(gclk));
	jdff dff_A_Vlr5r1QO1_2(.dout(w_dff_A_1cobA0TI7_2),.din(w_dff_A_Vlr5r1QO1_2),.clk(gclk));
	jdff dff_A_XsHFxLCG5_2(.dout(w_dff_A_Vlr5r1QO1_2),.din(w_dff_A_XsHFxLCG5_2),.clk(gclk));
	jdff dff_A_TfcDO0ZB1_2(.dout(w_dff_A_XsHFxLCG5_2),.din(w_dff_A_TfcDO0ZB1_2),.clk(gclk));
	jdff dff_A_aA9mping5_2(.dout(w_dff_A_TfcDO0ZB1_2),.din(w_dff_A_aA9mping5_2),.clk(gclk));
	jdff dff_A_dMpSaAdQ9_2(.dout(w_dff_A_aA9mping5_2),.din(w_dff_A_dMpSaAdQ9_2),.clk(gclk));
	jdff dff_A_y2qxMShh2_2(.dout(w_dff_A_dMpSaAdQ9_2),.din(w_dff_A_y2qxMShh2_2),.clk(gclk));
	jdff dff_A_yrOUtYlm7_2(.dout(w_dff_A_y2qxMShh2_2),.din(w_dff_A_yrOUtYlm7_2),.clk(gclk));
	jdff dff_A_3t3whZ2Y3_2(.dout(w_dff_A_yrOUtYlm7_2),.din(w_dff_A_3t3whZ2Y3_2),.clk(gclk));
	jdff dff_A_dahGnmyB9_2(.dout(w_dff_A_3t3whZ2Y3_2),.din(w_dff_A_dahGnmyB9_2),.clk(gclk));
	jdff dff_A_IaEcCyU10_1(.dout(w_G1694_0[1]),.din(w_dff_A_IaEcCyU10_1),.clk(gclk));
	jdff dff_A_zWSyWcJh3_2(.dout(w_G1691_0[2]),.din(w_dff_A_zWSyWcJh3_2),.clk(gclk));
	jdff dff_B_PaArHjYw6_2(.din(n1624),.dout(w_dff_B_PaArHjYw6_2),.clk(gclk));
	jdff dff_B_zdbVsq0K2_2(.din(w_dff_B_PaArHjYw6_2),.dout(w_dff_B_zdbVsq0K2_2),.clk(gclk));
	jdff dff_B_VKhCWsLv7_2(.din(w_dff_B_zdbVsq0K2_2),.dout(w_dff_B_VKhCWsLv7_2),.clk(gclk));
	jdff dff_B_MeLGRvv19_2(.din(w_dff_B_VKhCWsLv7_2),.dout(w_dff_B_MeLGRvv19_2),.clk(gclk));
	jdff dff_B_DeWhxuHb4_2(.din(w_dff_B_MeLGRvv19_2),.dout(w_dff_B_DeWhxuHb4_2),.clk(gclk));
	jdff dff_B_hyVuRBW98_2(.din(w_dff_B_DeWhxuHb4_2),.dout(w_dff_B_hyVuRBW98_2),.clk(gclk));
	jdff dff_B_a8R01oOk4_2(.din(w_dff_B_hyVuRBW98_2),.dout(w_dff_B_a8R01oOk4_2),.clk(gclk));
	jdff dff_B_ZgqPkHwa6_2(.din(w_dff_B_a8R01oOk4_2),.dout(w_dff_B_ZgqPkHwa6_2),.clk(gclk));
	jdff dff_B_0fV5U8zh0_2(.din(w_dff_B_ZgqPkHwa6_2),.dout(w_dff_B_0fV5U8zh0_2),.clk(gclk));
	jdff dff_B_IH5kUP9c2_2(.din(w_dff_B_0fV5U8zh0_2),.dout(w_dff_B_IH5kUP9c2_2),.clk(gclk));
	jdff dff_B_np9OwCyc2_2(.din(w_dff_B_IH5kUP9c2_2),.dout(w_dff_B_np9OwCyc2_2),.clk(gclk));
	jdff dff_B_lcY3qdge8_2(.din(w_dff_B_np9OwCyc2_2),.dout(w_dff_B_lcY3qdge8_2),.clk(gclk));
	jdff dff_B_j0zQEHMk1_2(.din(w_dff_B_lcY3qdge8_2),.dout(w_dff_B_j0zQEHMk1_2),.clk(gclk));
	jdff dff_B_Z66bq53k5_2(.din(w_dff_B_j0zQEHMk1_2),.dout(w_dff_B_Z66bq53k5_2),.clk(gclk));
	jdff dff_B_czvFAzS05_2(.din(w_dff_B_Z66bq53k5_2),.dout(w_dff_B_czvFAzS05_2),.clk(gclk));
	jdff dff_B_4T5ih9X59_2(.din(w_dff_B_czvFAzS05_2),.dout(w_dff_B_4T5ih9X59_2),.clk(gclk));
	jdff dff_B_0gAnX0VS6_2(.din(w_dff_B_4T5ih9X59_2),.dout(w_dff_B_0gAnX0VS6_2),.clk(gclk));
	jdff dff_B_uAU7InlV9_2(.din(w_dff_B_0gAnX0VS6_2),.dout(w_dff_B_uAU7InlV9_2),.clk(gclk));
	jdff dff_B_hDQiykh92_2(.din(w_dff_B_uAU7InlV9_2),.dout(w_dff_B_hDQiykh92_2),.clk(gclk));
	jdff dff_B_leXMfk1o1_2(.din(w_dff_B_hDQiykh92_2),.dout(w_dff_B_leXMfk1o1_2),.clk(gclk));
	jdff dff_B_4nDZVYd27_2(.din(w_dff_B_leXMfk1o1_2),.dout(w_dff_B_4nDZVYd27_2),.clk(gclk));
	jdff dff_B_z5pUiMO61_2(.din(w_dff_B_4nDZVYd27_2),.dout(w_dff_B_z5pUiMO61_2),.clk(gclk));
	jdff dff_B_FIxQMkhB5_2(.din(w_dff_B_z5pUiMO61_2),.dout(w_dff_B_FIxQMkhB5_2),.clk(gclk));
	jdff dff_B_HJ0gmp534_2(.din(w_dff_B_FIxQMkhB5_2),.dout(w_dff_B_HJ0gmp534_2),.clk(gclk));
	jdff dff_A_hWHP13Na3_2(.dout(w_G137_3[2]),.din(w_dff_A_hWHP13Na3_2),.clk(gclk));
	jdff dff_A_yWb9TyGp6_2(.dout(w_dff_A_hWHP13Na3_2),.din(w_dff_A_yWb9TyGp6_2),.clk(gclk));
	jdff dff_A_3Jn64Rcv4_2(.dout(w_dff_A_yWb9TyGp6_2),.din(w_dff_A_3Jn64Rcv4_2),.clk(gclk));
	jdff dff_A_fNDQtBoU9_2(.dout(w_dff_A_3Jn64Rcv4_2),.din(w_dff_A_fNDQtBoU9_2),.clk(gclk));
	jdff dff_A_1oiwm1U34_2(.dout(w_dff_A_fNDQtBoU9_2),.din(w_dff_A_1oiwm1U34_2),.clk(gclk));
	jdff dff_A_wmJ7KXU28_2(.dout(w_dff_A_1oiwm1U34_2),.din(w_dff_A_wmJ7KXU28_2),.clk(gclk));
	jdff dff_A_g2NadnpD6_2(.dout(w_dff_A_wmJ7KXU28_2),.din(w_dff_A_g2NadnpD6_2),.clk(gclk));
	jdff dff_A_8N7lv18q8_2(.dout(w_dff_A_g2NadnpD6_2),.din(w_dff_A_8N7lv18q8_2),.clk(gclk));
	jdff dff_A_QfF5VCWS8_2(.dout(w_dff_A_8N7lv18q8_2),.din(w_dff_A_QfF5VCWS8_2),.clk(gclk));
	jdff dff_A_QB9sNRC20_2(.dout(w_dff_A_QfF5VCWS8_2),.din(w_dff_A_QB9sNRC20_2),.clk(gclk));
	jdff dff_A_rgcB032A9_2(.dout(w_dff_A_QB9sNRC20_2),.din(w_dff_A_rgcB032A9_2),.clk(gclk));
	jdff dff_A_2kXcv5EP4_2(.dout(w_dff_A_rgcB032A9_2),.din(w_dff_A_2kXcv5EP4_2),.clk(gclk));
	jdff dff_A_ELTcECpr2_2(.dout(w_dff_A_2kXcv5EP4_2),.din(w_dff_A_ELTcECpr2_2),.clk(gclk));
	jdff dff_A_8lGAZe4P5_2(.dout(w_dff_A_ELTcECpr2_2),.din(w_dff_A_8lGAZe4P5_2),.clk(gclk));
	jdff dff_A_am4IBHpH9_2(.dout(w_dff_A_8lGAZe4P5_2),.din(w_dff_A_am4IBHpH9_2),.clk(gclk));
	jdff dff_A_Sp41L3gm8_2(.dout(w_dff_A_am4IBHpH9_2),.din(w_dff_A_Sp41L3gm8_2),.clk(gclk));
	jdff dff_A_qNgS8F394_2(.dout(w_dff_A_Sp41L3gm8_2),.din(w_dff_A_qNgS8F394_2),.clk(gclk));
	jdff dff_A_iqdgmdfO7_2(.dout(w_dff_A_qNgS8F394_2),.din(w_dff_A_iqdgmdfO7_2),.clk(gclk));
	jdff dff_A_RXfGAZfL9_2(.dout(w_dff_A_iqdgmdfO7_2),.din(w_dff_A_RXfGAZfL9_2),.clk(gclk));
	jdff dff_A_hCrS64lY0_2(.dout(w_dff_A_RXfGAZfL9_2),.din(w_dff_A_hCrS64lY0_2),.clk(gclk));
	jdff dff_A_NICqD9a91_2(.dout(w_dff_A_hCrS64lY0_2),.din(w_dff_A_NICqD9a91_2),.clk(gclk));
	jdff dff_A_KJlkTg9i7_2(.dout(w_dff_A_NICqD9a91_2),.din(w_dff_A_KJlkTg9i7_2),.clk(gclk));
	jdff dff_A_QGAAvwDb4_2(.dout(w_dff_A_KJlkTg9i7_2),.din(w_dff_A_QGAAvwDb4_2),.clk(gclk));
	jdff dff_A_tU1ov6fD1_0(.dout(w_G137_0[0]),.din(w_dff_A_tU1ov6fD1_0),.clk(gclk));
	jdff dff_A_dJhWGqua3_0(.dout(w_dff_A_tU1ov6fD1_0),.din(w_dff_A_dJhWGqua3_0),.clk(gclk));
	jdff dff_A_bISyXt4b5_0(.dout(w_dff_A_dJhWGqua3_0),.din(w_dff_A_bISyXt4b5_0),.clk(gclk));
	jdff dff_A_F6sRyIu06_0(.dout(w_dff_A_bISyXt4b5_0),.din(w_dff_A_F6sRyIu06_0),.clk(gclk));
	jdff dff_A_nKozoKNF7_0(.dout(w_dff_A_F6sRyIu06_0),.din(w_dff_A_nKozoKNF7_0),.clk(gclk));
	jdff dff_A_4g0sPfdQ3_0(.dout(w_dff_A_nKozoKNF7_0),.din(w_dff_A_4g0sPfdQ3_0),.clk(gclk));
	jdff dff_A_hMi0SqkB0_0(.dout(w_dff_A_4g0sPfdQ3_0),.din(w_dff_A_hMi0SqkB0_0),.clk(gclk));
	jdff dff_A_uom8rbJg7_0(.dout(w_dff_A_hMi0SqkB0_0),.din(w_dff_A_uom8rbJg7_0),.clk(gclk));
	jdff dff_A_i8ENp6xF8_0(.dout(w_dff_A_uom8rbJg7_0),.din(w_dff_A_i8ENp6xF8_0),.clk(gclk));
	jdff dff_A_ntJvPZ7t5_0(.dout(w_dff_A_i8ENp6xF8_0),.din(w_dff_A_ntJvPZ7t5_0),.clk(gclk));
	jdff dff_A_7w2cHXdd8_0(.dout(w_dff_A_ntJvPZ7t5_0),.din(w_dff_A_7w2cHXdd8_0),.clk(gclk));
	jdff dff_A_nTlvFufY7_0(.dout(w_dff_A_7w2cHXdd8_0),.din(w_dff_A_nTlvFufY7_0),.clk(gclk));
	jdff dff_A_7SJP1IDB0_0(.dout(w_dff_A_nTlvFufY7_0),.din(w_dff_A_7SJP1IDB0_0),.clk(gclk));
	jdff dff_A_IcvyyfZm0_0(.dout(w_dff_A_7SJP1IDB0_0),.din(w_dff_A_IcvyyfZm0_0),.clk(gclk));
	jdff dff_A_nAywAc2n6_0(.dout(w_dff_A_IcvyyfZm0_0),.din(w_dff_A_nAywAc2n6_0),.clk(gclk));
	jdff dff_A_y8EKslp71_0(.dout(w_dff_A_nAywAc2n6_0),.din(w_dff_A_y8EKslp71_0),.clk(gclk));
	jdff dff_A_7M70bVjP4_1(.dout(w_G137_0[1]),.din(w_dff_A_7M70bVjP4_1),.clk(gclk));
	jdff dff_A_6zeM2juR0_1(.dout(w_dff_A_7M70bVjP4_1),.din(w_dff_A_6zeM2juR0_1),.clk(gclk));
	jdff dff_A_W0s8m6Dw6_1(.dout(w_dff_A_6zeM2juR0_1),.din(w_dff_A_W0s8m6Dw6_1),.clk(gclk));
	jdff dff_A_J80eq6C52_1(.dout(w_dff_A_W0s8m6Dw6_1),.din(w_dff_A_J80eq6C52_1),.clk(gclk));
	jdff dff_A_M0S4rPp63_1(.dout(w_dff_A_J80eq6C52_1),.din(w_dff_A_M0S4rPp63_1),.clk(gclk));
	jdff dff_A_tD29lgOE2_1(.dout(w_dff_A_M0S4rPp63_1),.din(w_dff_A_tD29lgOE2_1),.clk(gclk));
	jdff dff_A_1ZsIH3Tu9_1(.dout(w_dff_A_tD29lgOE2_1),.din(w_dff_A_1ZsIH3Tu9_1),.clk(gclk));
	jdff dff_A_N89QNPHs4_1(.dout(w_dff_A_1ZsIH3Tu9_1),.din(w_dff_A_N89QNPHs4_1),.clk(gclk));
	jdff dff_A_BweG7lt36_1(.dout(w_dff_A_N89QNPHs4_1),.din(w_dff_A_BweG7lt36_1),.clk(gclk));
	jdff dff_A_55ArJU9c9_1(.dout(w_dff_A_BweG7lt36_1),.din(w_dff_A_55ArJU9c9_1),.clk(gclk));
	jdff dff_A_7BUQRPrB0_1(.dout(w_dff_A_55ArJU9c9_1),.din(w_dff_A_7BUQRPrB0_1),.clk(gclk));
	jdff dff_A_okV472fm6_1(.dout(w_dff_A_ogv3lNCr0_0),.din(w_dff_A_okV472fm6_1),.clk(gclk));
	jdff dff_A_ogv3lNCr0_0(.dout(w_dff_A_oV1uorzV5_0),.din(w_dff_A_ogv3lNCr0_0),.clk(gclk));
	jdff dff_A_oV1uorzV5_0(.dout(w_dff_A_6ezAHKGO0_0),.din(w_dff_A_oV1uorzV5_0),.clk(gclk));
	jdff dff_A_6ezAHKGO0_0(.dout(w_dff_A_mfQVpu4y6_0),.din(w_dff_A_6ezAHKGO0_0),.clk(gclk));
	jdff dff_A_mfQVpu4y6_0(.dout(w_dff_A_5XrMRjGZ9_0),.din(w_dff_A_mfQVpu4y6_0),.clk(gclk));
	jdff dff_A_5XrMRjGZ9_0(.dout(w_dff_A_QSIOIiXg8_0),.din(w_dff_A_5XrMRjGZ9_0),.clk(gclk));
	jdff dff_A_QSIOIiXg8_0(.dout(w_dff_A_IIrlkdnD9_0),.din(w_dff_A_QSIOIiXg8_0),.clk(gclk));
	jdff dff_A_IIrlkdnD9_0(.dout(w_dff_A_kJYYLnkk0_0),.din(w_dff_A_IIrlkdnD9_0),.clk(gclk));
	jdff dff_A_kJYYLnkk0_0(.dout(w_dff_A_2KhvLaZT1_0),.din(w_dff_A_kJYYLnkk0_0),.clk(gclk));
	jdff dff_A_2KhvLaZT1_0(.dout(w_dff_A_zknnBtXH6_0),.din(w_dff_A_2KhvLaZT1_0),.clk(gclk));
	jdff dff_A_zknnBtXH6_0(.dout(w_dff_A_163sYPsF4_0),.din(w_dff_A_zknnBtXH6_0),.clk(gclk));
	jdff dff_A_163sYPsF4_0(.dout(w_dff_A_3llhc7En7_0),.din(w_dff_A_163sYPsF4_0),.clk(gclk));
	jdff dff_A_3llhc7En7_0(.dout(w_dff_A_KXjDxkDD7_0),.din(w_dff_A_3llhc7En7_0),.clk(gclk));
	jdff dff_A_KXjDxkDD7_0(.dout(w_dff_A_XiqObUWP7_0),.din(w_dff_A_KXjDxkDD7_0),.clk(gclk));
	jdff dff_A_XiqObUWP7_0(.dout(w_dff_A_StNbPVKd8_0),.din(w_dff_A_XiqObUWP7_0),.clk(gclk));
	jdff dff_A_StNbPVKd8_0(.dout(w_dff_A_p2lsyuUi2_0),.din(w_dff_A_StNbPVKd8_0),.clk(gclk));
	jdff dff_A_p2lsyuUi2_0(.dout(w_dff_A_qM7m0ZwE3_0),.din(w_dff_A_p2lsyuUi2_0),.clk(gclk));
	jdff dff_A_qM7m0ZwE3_0(.dout(w_dff_A_asfHprWw6_0),.din(w_dff_A_qM7m0ZwE3_0),.clk(gclk));
	jdff dff_A_asfHprWw6_0(.dout(w_dff_A_rA6LTo662_0),.din(w_dff_A_asfHprWw6_0),.clk(gclk));
	jdff dff_A_rA6LTo662_0(.dout(w_dff_A_LTWHRYH73_0),.din(w_dff_A_rA6LTo662_0),.clk(gclk));
	jdff dff_A_LTWHRYH73_0(.dout(w_dff_A_hpVaIVDg6_0),.din(w_dff_A_LTWHRYH73_0),.clk(gclk));
	jdff dff_A_hpVaIVDg6_0(.dout(w_dff_A_eJ703AlT6_0),.din(w_dff_A_hpVaIVDg6_0),.clk(gclk));
	jdff dff_A_eJ703AlT6_0(.dout(w_dff_A_glrjwNps1_0),.din(w_dff_A_eJ703AlT6_0),.clk(gclk));
	jdff dff_A_glrjwNps1_0(.dout(w_dff_A_HkFzjxmf8_0),.din(w_dff_A_glrjwNps1_0),.clk(gclk));
	jdff dff_A_HkFzjxmf8_0(.dout(w_dff_A_Vfdcr69x0_0),.din(w_dff_A_HkFzjxmf8_0),.clk(gclk));
	jdff dff_A_Vfdcr69x0_0(.dout(G144),.din(w_dff_A_Vfdcr69x0_0),.clk(gclk));
	jdff dff_A_NZDPOgPm2_1(.dout(w_dff_A_ZyfyjtQ58_0),.din(w_dff_A_NZDPOgPm2_1),.clk(gclk));
	jdff dff_A_ZyfyjtQ58_0(.dout(w_dff_A_xUsn0j0M1_0),.din(w_dff_A_ZyfyjtQ58_0),.clk(gclk));
	jdff dff_A_xUsn0j0M1_0(.dout(w_dff_A_ZemeG7VO1_0),.din(w_dff_A_xUsn0j0M1_0),.clk(gclk));
	jdff dff_A_ZemeG7VO1_0(.dout(w_dff_A_8hP8GLcc6_0),.din(w_dff_A_ZemeG7VO1_0),.clk(gclk));
	jdff dff_A_8hP8GLcc6_0(.dout(w_dff_A_7IS9ToZb2_0),.din(w_dff_A_8hP8GLcc6_0),.clk(gclk));
	jdff dff_A_7IS9ToZb2_0(.dout(w_dff_A_kZamQdsq8_0),.din(w_dff_A_7IS9ToZb2_0),.clk(gclk));
	jdff dff_A_kZamQdsq8_0(.dout(w_dff_A_8wx8sm6s8_0),.din(w_dff_A_kZamQdsq8_0),.clk(gclk));
	jdff dff_A_8wx8sm6s8_0(.dout(w_dff_A_gJV0myzi1_0),.din(w_dff_A_8wx8sm6s8_0),.clk(gclk));
	jdff dff_A_gJV0myzi1_0(.dout(w_dff_A_a6epFmHE2_0),.din(w_dff_A_gJV0myzi1_0),.clk(gclk));
	jdff dff_A_a6epFmHE2_0(.dout(w_dff_A_zZxeVQxT1_0),.din(w_dff_A_a6epFmHE2_0),.clk(gclk));
	jdff dff_A_zZxeVQxT1_0(.dout(w_dff_A_uocuKcTo0_0),.din(w_dff_A_zZxeVQxT1_0),.clk(gclk));
	jdff dff_A_uocuKcTo0_0(.dout(w_dff_A_ZVEl00kN4_0),.din(w_dff_A_uocuKcTo0_0),.clk(gclk));
	jdff dff_A_ZVEl00kN4_0(.dout(w_dff_A_LHnIaVZn7_0),.din(w_dff_A_ZVEl00kN4_0),.clk(gclk));
	jdff dff_A_LHnIaVZn7_0(.dout(w_dff_A_I6zfqJfT1_0),.din(w_dff_A_LHnIaVZn7_0),.clk(gclk));
	jdff dff_A_I6zfqJfT1_0(.dout(w_dff_A_C9SvRgiR4_0),.din(w_dff_A_I6zfqJfT1_0),.clk(gclk));
	jdff dff_A_C9SvRgiR4_0(.dout(w_dff_A_krBIP1DP1_0),.din(w_dff_A_C9SvRgiR4_0),.clk(gclk));
	jdff dff_A_krBIP1DP1_0(.dout(w_dff_A_6WtM4WiY7_0),.din(w_dff_A_krBIP1DP1_0),.clk(gclk));
	jdff dff_A_6WtM4WiY7_0(.dout(w_dff_A_NnYtvDvs9_0),.din(w_dff_A_6WtM4WiY7_0),.clk(gclk));
	jdff dff_A_NnYtvDvs9_0(.dout(w_dff_A_n6teTyJa8_0),.din(w_dff_A_NnYtvDvs9_0),.clk(gclk));
	jdff dff_A_n6teTyJa8_0(.dout(w_dff_A_yztdqtqJ6_0),.din(w_dff_A_n6teTyJa8_0),.clk(gclk));
	jdff dff_A_yztdqtqJ6_0(.dout(w_dff_A_IrafUO6r5_0),.din(w_dff_A_yztdqtqJ6_0),.clk(gclk));
	jdff dff_A_IrafUO6r5_0(.dout(w_dff_A_wExJG9WZ4_0),.din(w_dff_A_IrafUO6r5_0),.clk(gclk));
	jdff dff_A_wExJG9WZ4_0(.dout(w_dff_A_YYGfBxpA6_0),.din(w_dff_A_wExJG9WZ4_0),.clk(gclk));
	jdff dff_A_YYGfBxpA6_0(.dout(w_dff_A_SMhb38CL7_0),.din(w_dff_A_YYGfBxpA6_0),.clk(gclk));
	jdff dff_A_SMhb38CL7_0(.dout(w_dff_A_BZ2jFIPl8_0),.din(w_dff_A_SMhb38CL7_0),.clk(gclk));
	jdff dff_A_BZ2jFIPl8_0(.dout(G298),.din(w_dff_A_BZ2jFIPl8_0),.clk(gclk));
	jdff dff_A_8SfPKRXf1_1(.dout(w_dff_A_LlC6qNoO9_0),.din(w_dff_A_8SfPKRXf1_1),.clk(gclk));
	jdff dff_A_LlC6qNoO9_0(.dout(w_dff_A_HqNFrRRt4_0),.din(w_dff_A_LlC6qNoO9_0),.clk(gclk));
	jdff dff_A_HqNFrRRt4_0(.dout(w_dff_A_yvZDnkZh2_0),.din(w_dff_A_HqNFrRRt4_0),.clk(gclk));
	jdff dff_A_yvZDnkZh2_0(.dout(w_dff_A_9t4xMM6Z8_0),.din(w_dff_A_yvZDnkZh2_0),.clk(gclk));
	jdff dff_A_9t4xMM6Z8_0(.dout(w_dff_A_Kt8rJOXo9_0),.din(w_dff_A_9t4xMM6Z8_0),.clk(gclk));
	jdff dff_A_Kt8rJOXo9_0(.dout(w_dff_A_Jm1bYKHC5_0),.din(w_dff_A_Kt8rJOXo9_0),.clk(gclk));
	jdff dff_A_Jm1bYKHC5_0(.dout(w_dff_A_mqLiPzgE7_0),.din(w_dff_A_Jm1bYKHC5_0),.clk(gclk));
	jdff dff_A_mqLiPzgE7_0(.dout(w_dff_A_14G34L1o0_0),.din(w_dff_A_mqLiPzgE7_0),.clk(gclk));
	jdff dff_A_14G34L1o0_0(.dout(w_dff_A_GZudCT3D3_0),.din(w_dff_A_14G34L1o0_0),.clk(gclk));
	jdff dff_A_GZudCT3D3_0(.dout(w_dff_A_c7FLgvys3_0),.din(w_dff_A_GZudCT3D3_0),.clk(gclk));
	jdff dff_A_c7FLgvys3_0(.dout(w_dff_A_uUgr2uCA1_0),.din(w_dff_A_c7FLgvys3_0),.clk(gclk));
	jdff dff_A_uUgr2uCA1_0(.dout(w_dff_A_eScK2o8I6_0),.din(w_dff_A_uUgr2uCA1_0),.clk(gclk));
	jdff dff_A_eScK2o8I6_0(.dout(w_dff_A_XRUibDmM2_0),.din(w_dff_A_eScK2o8I6_0),.clk(gclk));
	jdff dff_A_XRUibDmM2_0(.dout(w_dff_A_j7RkDJ4j3_0),.din(w_dff_A_XRUibDmM2_0),.clk(gclk));
	jdff dff_A_j7RkDJ4j3_0(.dout(w_dff_A_K3BJWmvQ8_0),.din(w_dff_A_j7RkDJ4j3_0),.clk(gclk));
	jdff dff_A_K3BJWmvQ8_0(.dout(w_dff_A_xK8qpfUj2_0),.din(w_dff_A_K3BJWmvQ8_0),.clk(gclk));
	jdff dff_A_xK8qpfUj2_0(.dout(w_dff_A_6rP5M31f8_0),.din(w_dff_A_xK8qpfUj2_0),.clk(gclk));
	jdff dff_A_6rP5M31f8_0(.dout(w_dff_A_K2sNMlaT7_0),.din(w_dff_A_6rP5M31f8_0),.clk(gclk));
	jdff dff_A_K2sNMlaT7_0(.dout(w_dff_A_E2qBVsr26_0),.din(w_dff_A_K2sNMlaT7_0),.clk(gclk));
	jdff dff_A_E2qBVsr26_0(.dout(w_dff_A_jXxYKFhQ5_0),.din(w_dff_A_E2qBVsr26_0),.clk(gclk));
	jdff dff_A_jXxYKFhQ5_0(.dout(w_dff_A_QFhRrDUe9_0),.din(w_dff_A_jXxYKFhQ5_0),.clk(gclk));
	jdff dff_A_QFhRrDUe9_0(.dout(w_dff_A_8tPwtVAx0_0),.din(w_dff_A_QFhRrDUe9_0),.clk(gclk));
	jdff dff_A_8tPwtVAx0_0(.dout(w_dff_A_0R8davIi8_0),.din(w_dff_A_8tPwtVAx0_0),.clk(gclk));
	jdff dff_A_0R8davIi8_0(.dout(w_dff_A_6WpTeIW55_0),.din(w_dff_A_0R8davIi8_0),.clk(gclk));
	jdff dff_A_6WpTeIW55_0(.dout(w_dff_A_mZUjYeH90_0),.din(w_dff_A_6WpTeIW55_0),.clk(gclk));
	jdff dff_A_mZUjYeH90_0(.dout(G973),.din(w_dff_A_mZUjYeH90_0),.clk(gclk));
	jdff dff_A_V5AYLoBR3_1(.dout(w_dff_A_cK7bFte06_0),.din(w_dff_A_V5AYLoBR3_1),.clk(gclk));
	jdff dff_A_cK7bFte06_0(.dout(w_dff_A_bEIyv3CV0_0),.din(w_dff_A_cK7bFte06_0),.clk(gclk));
	jdff dff_A_bEIyv3CV0_0(.dout(w_dff_A_SvnUPLiK5_0),.din(w_dff_A_bEIyv3CV0_0),.clk(gclk));
	jdff dff_A_SvnUPLiK5_0(.dout(w_dff_A_dIn0g7Gl1_0),.din(w_dff_A_SvnUPLiK5_0),.clk(gclk));
	jdff dff_A_dIn0g7Gl1_0(.dout(w_dff_A_y6CqniDP2_0),.din(w_dff_A_dIn0g7Gl1_0),.clk(gclk));
	jdff dff_A_y6CqniDP2_0(.dout(w_dff_A_HP5Z9x121_0),.din(w_dff_A_y6CqniDP2_0),.clk(gclk));
	jdff dff_A_HP5Z9x121_0(.dout(w_dff_A_o2wPvOQr5_0),.din(w_dff_A_HP5Z9x121_0),.clk(gclk));
	jdff dff_A_o2wPvOQr5_0(.dout(w_dff_A_vjXx6cGV7_0),.din(w_dff_A_o2wPvOQr5_0),.clk(gclk));
	jdff dff_A_vjXx6cGV7_0(.dout(w_dff_A_WC6WBIOd7_0),.din(w_dff_A_vjXx6cGV7_0),.clk(gclk));
	jdff dff_A_WC6WBIOd7_0(.dout(w_dff_A_O6BdxDHu8_0),.din(w_dff_A_WC6WBIOd7_0),.clk(gclk));
	jdff dff_A_O6BdxDHu8_0(.dout(w_dff_A_MLAbcBpK0_0),.din(w_dff_A_O6BdxDHu8_0),.clk(gclk));
	jdff dff_A_MLAbcBpK0_0(.dout(w_dff_A_JTrxyZqm5_0),.din(w_dff_A_MLAbcBpK0_0),.clk(gclk));
	jdff dff_A_JTrxyZqm5_0(.dout(w_dff_A_DMMdjmFM7_0),.din(w_dff_A_JTrxyZqm5_0),.clk(gclk));
	jdff dff_A_DMMdjmFM7_0(.dout(w_dff_A_8L68Y3DV7_0),.din(w_dff_A_DMMdjmFM7_0),.clk(gclk));
	jdff dff_A_8L68Y3DV7_0(.dout(w_dff_A_dYTMK3Rp9_0),.din(w_dff_A_8L68Y3DV7_0),.clk(gclk));
	jdff dff_A_dYTMK3Rp9_0(.dout(w_dff_A_MmXwx7mn3_0),.din(w_dff_A_dYTMK3Rp9_0),.clk(gclk));
	jdff dff_A_MmXwx7mn3_0(.dout(w_dff_A_yf4b1s9v4_0),.din(w_dff_A_MmXwx7mn3_0),.clk(gclk));
	jdff dff_A_yf4b1s9v4_0(.dout(w_dff_A_VHClbzyf3_0),.din(w_dff_A_yf4b1s9v4_0),.clk(gclk));
	jdff dff_A_VHClbzyf3_0(.dout(w_dff_A_MMnRv6694_0),.din(w_dff_A_VHClbzyf3_0),.clk(gclk));
	jdff dff_A_MMnRv6694_0(.dout(w_dff_A_pH0bz1jt6_0),.din(w_dff_A_MMnRv6694_0),.clk(gclk));
	jdff dff_A_pH0bz1jt6_0(.dout(w_dff_A_JXJiJwas5_0),.din(w_dff_A_pH0bz1jt6_0),.clk(gclk));
	jdff dff_A_JXJiJwas5_0(.dout(w_dff_A_6Z1n3bKR4_0),.din(w_dff_A_JXJiJwas5_0),.clk(gclk));
	jdff dff_A_6Z1n3bKR4_0(.dout(w_dff_A_4bxgWxj34_0),.din(w_dff_A_6Z1n3bKR4_0),.clk(gclk));
	jdff dff_A_4bxgWxj34_0(.dout(w_dff_A_hRtNzZgp9_0),.din(w_dff_A_4bxgWxj34_0),.clk(gclk));
	jdff dff_A_hRtNzZgp9_0(.dout(G594),.din(w_dff_A_hRtNzZgp9_0),.clk(gclk));
	jdff dff_A_3L9jc5wg9_1(.dout(w_dff_A_vEKKRsGd7_0),.din(w_dff_A_3L9jc5wg9_1),.clk(gclk));
	jdff dff_A_vEKKRsGd7_0(.dout(w_dff_A_Wkh1cTgd0_0),.din(w_dff_A_vEKKRsGd7_0),.clk(gclk));
	jdff dff_A_Wkh1cTgd0_0(.dout(w_dff_A_V4AD3w623_0),.din(w_dff_A_Wkh1cTgd0_0),.clk(gclk));
	jdff dff_A_V4AD3w623_0(.dout(w_dff_A_sEdITJI15_0),.din(w_dff_A_V4AD3w623_0),.clk(gclk));
	jdff dff_A_sEdITJI15_0(.dout(w_dff_A_KZojZsK95_0),.din(w_dff_A_sEdITJI15_0),.clk(gclk));
	jdff dff_A_KZojZsK95_0(.dout(w_dff_A_ME6bXSDU7_0),.din(w_dff_A_KZojZsK95_0),.clk(gclk));
	jdff dff_A_ME6bXSDU7_0(.dout(w_dff_A_372uKjDW6_0),.din(w_dff_A_ME6bXSDU7_0),.clk(gclk));
	jdff dff_A_372uKjDW6_0(.dout(w_dff_A_4ATw8BM06_0),.din(w_dff_A_372uKjDW6_0),.clk(gclk));
	jdff dff_A_4ATw8BM06_0(.dout(w_dff_A_LFNjDd318_0),.din(w_dff_A_4ATw8BM06_0),.clk(gclk));
	jdff dff_A_LFNjDd318_0(.dout(w_dff_A_dTxQpufI2_0),.din(w_dff_A_LFNjDd318_0),.clk(gclk));
	jdff dff_A_dTxQpufI2_0(.dout(w_dff_A_chJmIE7D0_0),.din(w_dff_A_dTxQpufI2_0),.clk(gclk));
	jdff dff_A_chJmIE7D0_0(.dout(w_dff_A_8BImmkCY5_0),.din(w_dff_A_chJmIE7D0_0),.clk(gclk));
	jdff dff_A_8BImmkCY5_0(.dout(w_dff_A_ORCTvjGy5_0),.din(w_dff_A_8BImmkCY5_0),.clk(gclk));
	jdff dff_A_ORCTvjGy5_0(.dout(w_dff_A_onIyKMjz1_0),.din(w_dff_A_ORCTvjGy5_0),.clk(gclk));
	jdff dff_A_onIyKMjz1_0(.dout(w_dff_A_o5ccFe7B0_0),.din(w_dff_A_onIyKMjz1_0),.clk(gclk));
	jdff dff_A_o5ccFe7B0_0(.dout(w_dff_A_IrbJFcy67_0),.din(w_dff_A_o5ccFe7B0_0),.clk(gclk));
	jdff dff_A_IrbJFcy67_0(.dout(w_dff_A_Foi1f5FH9_0),.din(w_dff_A_IrbJFcy67_0),.clk(gclk));
	jdff dff_A_Foi1f5FH9_0(.dout(w_dff_A_7hkYaTDD6_0),.din(w_dff_A_Foi1f5FH9_0),.clk(gclk));
	jdff dff_A_7hkYaTDD6_0(.dout(w_dff_A_cfovHEdE4_0),.din(w_dff_A_7hkYaTDD6_0),.clk(gclk));
	jdff dff_A_cfovHEdE4_0(.dout(w_dff_A_t7dss5vg3_0),.din(w_dff_A_cfovHEdE4_0),.clk(gclk));
	jdff dff_A_t7dss5vg3_0(.dout(w_dff_A_Q2ijlehy2_0),.din(w_dff_A_t7dss5vg3_0),.clk(gclk));
	jdff dff_A_Q2ijlehy2_0(.dout(w_dff_A_rkNQ3HYH3_0),.din(w_dff_A_Q2ijlehy2_0),.clk(gclk));
	jdff dff_A_rkNQ3HYH3_0(.dout(w_dff_A_IBfoackQ7_0),.din(w_dff_A_rkNQ3HYH3_0),.clk(gclk));
	jdff dff_A_IBfoackQ7_0(.dout(w_dff_A_jEwMu9cN4_0),.din(w_dff_A_IBfoackQ7_0),.clk(gclk));
	jdff dff_A_jEwMu9cN4_0(.dout(G599),.din(w_dff_A_jEwMu9cN4_0),.clk(gclk));
	jdff dff_A_p2Avj4Ok5_1(.dout(w_dff_A_PvkSDAGn4_0),.din(w_dff_A_p2Avj4Ok5_1),.clk(gclk));
	jdff dff_A_PvkSDAGn4_0(.dout(w_dff_A_jGTmYm5E9_0),.din(w_dff_A_PvkSDAGn4_0),.clk(gclk));
	jdff dff_A_jGTmYm5E9_0(.dout(w_dff_A_B0ncpjQE1_0),.din(w_dff_A_jGTmYm5E9_0),.clk(gclk));
	jdff dff_A_B0ncpjQE1_0(.dout(w_dff_A_nqm7mEeW9_0),.din(w_dff_A_B0ncpjQE1_0),.clk(gclk));
	jdff dff_A_nqm7mEeW9_0(.dout(w_dff_A_17ehKx0R9_0),.din(w_dff_A_nqm7mEeW9_0),.clk(gclk));
	jdff dff_A_17ehKx0R9_0(.dout(w_dff_A_Z4ZJUrZ52_0),.din(w_dff_A_17ehKx0R9_0),.clk(gclk));
	jdff dff_A_Z4ZJUrZ52_0(.dout(w_dff_A_yUxjOSnH4_0),.din(w_dff_A_Z4ZJUrZ52_0),.clk(gclk));
	jdff dff_A_yUxjOSnH4_0(.dout(w_dff_A_56DkgF726_0),.din(w_dff_A_yUxjOSnH4_0),.clk(gclk));
	jdff dff_A_56DkgF726_0(.dout(w_dff_A_LbyzknDR6_0),.din(w_dff_A_56DkgF726_0),.clk(gclk));
	jdff dff_A_LbyzknDR6_0(.dout(w_dff_A_hR7vLwDL6_0),.din(w_dff_A_LbyzknDR6_0),.clk(gclk));
	jdff dff_A_hR7vLwDL6_0(.dout(w_dff_A_xRInDINj1_0),.din(w_dff_A_hR7vLwDL6_0),.clk(gclk));
	jdff dff_A_xRInDINj1_0(.dout(w_dff_A_5A3jwpn55_0),.din(w_dff_A_xRInDINj1_0),.clk(gclk));
	jdff dff_A_5A3jwpn55_0(.dout(w_dff_A_LOftf9yg5_0),.din(w_dff_A_5A3jwpn55_0),.clk(gclk));
	jdff dff_A_LOftf9yg5_0(.dout(w_dff_A_s7wkQ6Hz1_0),.din(w_dff_A_LOftf9yg5_0),.clk(gclk));
	jdff dff_A_s7wkQ6Hz1_0(.dout(w_dff_A_T6XvvGTH9_0),.din(w_dff_A_s7wkQ6Hz1_0),.clk(gclk));
	jdff dff_A_T6XvvGTH9_0(.dout(w_dff_A_eoPN4I3c5_0),.din(w_dff_A_T6XvvGTH9_0),.clk(gclk));
	jdff dff_A_eoPN4I3c5_0(.dout(w_dff_A_TBM72KVF3_0),.din(w_dff_A_eoPN4I3c5_0),.clk(gclk));
	jdff dff_A_TBM72KVF3_0(.dout(w_dff_A_nBhgTgC88_0),.din(w_dff_A_TBM72KVF3_0),.clk(gclk));
	jdff dff_A_nBhgTgC88_0(.dout(w_dff_A_r6YHjFLu7_0),.din(w_dff_A_nBhgTgC88_0),.clk(gclk));
	jdff dff_A_r6YHjFLu7_0(.dout(w_dff_A_wpx4jmy09_0),.din(w_dff_A_r6YHjFLu7_0),.clk(gclk));
	jdff dff_A_wpx4jmy09_0(.dout(w_dff_A_HyFR7HTm2_0),.din(w_dff_A_wpx4jmy09_0),.clk(gclk));
	jdff dff_A_HyFR7HTm2_0(.dout(w_dff_A_3tnw3Zr51_0),.din(w_dff_A_HyFR7HTm2_0),.clk(gclk));
	jdff dff_A_3tnw3Zr51_0(.dout(w_dff_A_O6WhPV7G1_0),.din(w_dff_A_3tnw3Zr51_0),.clk(gclk));
	jdff dff_A_O6WhPV7G1_0(.dout(w_dff_A_WLQln4x22_0),.din(w_dff_A_O6WhPV7G1_0),.clk(gclk));
	jdff dff_A_WLQln4x22_0(.dout(G600),.din(w_dff_A_WLQln4x22_0),.clk(gclk));
	jdff dff_A_dz8Ft8Lm5_1(.dout(w_dff_A_JSDsn5kA7_0),.din(w_dff_A_dz8Ft8Lm5_1),.clk(gclk));
	jdff dff_A_JSDsn5kA7_0(.dout(w_dff_A_YLSG9GNz5_0),.din(w_dff_A_JSDsn5kA7_0),.clk(gclk));
	jdff dff_A_YLSG9GNz5_0(.dout(w_dff_A_7F0UaqCH5_0),.din(w_dff_A_YLSG9GNz5_0),.clk(gclk));
	jdff dff_A_7F0UaqCH5_0(.dout(w_dff_A_zatp2yiT1_0),.din(w_dff_A_7F0UaqCH5_0),.clk(gclk));
	jdff dff_A_zatp2yiT1_0(.dout(w_dff_A_9B6YAoJi9_0),.din(w_dff_A_zatp2yiT1_0),.clk(gclk));
	jdff dff_A_9B6YAoJi9_0(.dout(w_dff_A_czAkkZYJ4_0),.din(w_dff_A_9B6YAoJi9_0),.clk(gclk));
	jdff dff_A_czAkkZYJ4_0(.dout(w_dff_A_aVAMlb7C0_0),.din(w_dff_A_czAkkZYJ4_0),.clk(gclk));
	jdff dff_A_aVAMlb7C0_0(.dout(w_dff_A_1g9QgtAa1_0),.din(w_dff_A_aVAMlb7C0_0),.clk(gclk));
	jdff dff_A_1g9QgtAa1_0(.dout(w_dff_A_mvp3yt8P4_0),.din(w_dff_A_1g9QgtAa1_0),.clk(gclk));
	jdff dff_A_mvp3yt8P4_0(.dout(w_dff_A_5P0tR7P50_0),.din(w_dff_A_mvp3yt8P4_0),.clk(gclk));
	jdff dff_A_5P0tR7P50_0(.dout(w_dff_A_4IeFLxLt1_0),.din(w_dff_A_5P0tR7P50_0),.clk(gclk));
	jdff dff_A_4IeFLxLt1_0(.dout(w_dff_A_71tAsMEu9_0),.din(w_dff_A_4IeFLxLt1_0),.clk(gclk));
	jdff dff_A_71tAsMEu9_0(.dout(w_dff_A_CU8oE03d1_0),.din(w_dff_A_71tAsMEu9_0),.clk(gclk));
	jdff dff_A_CU8oE03d1_0(.dout(w_dff_A_U0PMj6Bc6_0),.din(w_dff_A_CU8oE03d1_0),.clk(gclk));
	jdff dff_A_U0PMj6Bc6_0(.dout(w_dff_A_fOQcQTle7_0),.din(w_dff_A_U0PMj6Bc6_0),.clk(gclk));
	jdff dff_A_fOQcQTle7_0(.dout(w_dff_A_6aSEVCcj7_0),.din(w_dff_A_fOQcQTle7_0),.clk(gclk));
	jdff dff_A_6aSEVCcj7_0(.dout(w_dff_A_1PUlN2gS0_0),.din(w_dff_A_6aSEVCcj7_0),.clk(gclk));
	jdff dff_A_1PUlN2gS0_0(.dout(w_dff_A_2oKprsdt4_0),.din(w_dff_A_1PUlN2gS0_0),.clk(gclk));
	jdff dff_A_2oKprsdt4_0(.dout(w_dff_A_Ob9qltBQ5_0),.din(w_dff_A_2oKprsdt4_0),.clk(gclk));
	jdff dff_A_Ob9qltBQ5_0(.dout(w_dff_A_bQC6ySv07_0),.din(w_dff_A_Ob9qltBQ5_0),.clk(gclk));
	jdff dff_A_bQC6ySv07_0(.dout(w_dff_A_QkI0g3Hq5_0),.din(w_dff_A_bQC6ySv07_0),.clk(gclk));
	jdff dff_A_QkI0g3Hq5_0(.dout(w_dff_A_sIJyTJWJ8_0),.din(w_dff_A_QkI0g3Hq5_0),.clk(gclk));
	jdff dff_A_sIJyTJWJ8_0(.dout(w_dff_A_UTG4Somq5_0),.din(w_dff_A_sIJyTJWJ8_0),.clk(gclk));
	jdff dff_A_UTG4Somq5_0(.dout(w_dff_A_6VZBjnF37_0),.din(w_dff_A_UTG4Somq5_0),.clk(gclk));
	jdff dff_A_6VZBjnF37_0(.dout(G601),.din(w_dff_A_6VZBjnF37_0),.clk(gclk));
	jdff dff_A_s2RVKcId6_1(.dout(w_dff_A_tATd9YJz8_0),.din(w_dff_A_s2RVKcId6_1),.clk(gclk));
	jdff dff_A_tATd9YJz8_0(.dout(w_dff_A_6NubUDHE1_0),.din(w_dff_A_tATd9YJz8_0),.clk(gclk));
	jdff dff_A_6NubUDHE1_0(.dout(w_dff_A_rUf7Mbw61_0),.din(w_dff_A_6NubUDHE1_0),.clk(gclk));
	jdff dff_A_rUf7Mbw61_0(.dout(w_dff_A_uXM7UcU86_0),.din(w_dff_A_rUf7Mbw61_0),.clk(gclk));
	jdff dff_A_uXM7UcU86_0(.dout(w_dff_A_MrQoWlc55_0),.din(w_dff_A_uXM7UcU86_0),.clk(gclk));
	jdff dff_A_MrQoWlc55_0(.dout(w_dff_A_UudJEs7V8_0),.din(w_dff_A_MrQoWlc55_0),.clk(gclk));
	jdff dff_A_UudJEs7V8_0(.dout(w_dff_A_hNPCBG3p9_0),.din(w_dff_A_UudJEs7V8_0),.clk(gclk));
	jdff dff_A_hNPCBG3p9_0(.dout(w_dff_A_VqGfESAb5_0),.din(w_dff_A_hNPCBG3p9_0),.clk(gclk));
	jdff dff_A_VqGfESAb5_0(.dout(w_dff_A_ngFzu4ba5_0),.din(w_dff_A_VqGfESAb5_0),.clk(gclk));
	jdff dff_A_ngFzu4ba5_0(.dout(w_dff_A_DmAxYJDc0_0),.din(w_dff_A_ngFzu4ba5_0),.clk(gclk));
	jdff dff_A_DmAxYJDc0_0(.dout(w_dff_A_f2DKxFer1_0),.din(w_dff_A_DmAxYJDc0_0),.clk(gclk));
	jdff dff_A_f2DKxFer1_0(.dout(w_dff_A_5oPoE5Ht3_0),.din(w_dff_A_f2DKxFer1_0),.clk(gclk));
	jdff dff_A_5oPoE5Ht3_0(.dout(w_dff_A_EaksyIGh6_0),.din(w_dff_A_5oPoE5Ht3_0),.clk(gclk));
	jdff dff_A_EaksyIGh6_0(.dout(w_dff_A_h5j7dwQU7_0),.din(w_dff_A_EaksyIGh6_0),.clk(gclk));
	jdff dff_A_h5j7dwQU7_0(.dout(w_dff_A_h1g6MR6z3_0),.din(w_dff_A_h5j7dwQU7_0),.clk(gclk));
	jdff dff_A_h1g6MR6z3_0(.dout(w_dff_A_UbL2vsxL3_0),.din(w_dff_A_h1g6MR6z3_0),.clk(gclk));
	jdff dff_A_UbL2vsxL3_0(.dout(w_dff_A_BIH5wCk30_0),.din(w_dff_A_UbL2vsxL3_0),.clk(gclk));
	jdff dff_A_BIH5wCk30_0(.dout(w_dff_A_GXcw6zQD2_0),.din(w_dff_A_BIH5wCk30_0),.clk(gclk));
	jdff dff_A_GXcw6zQD2_0(.dout(w_dff_A_uSOO17m51_0),.din(w_dff_A_GXcw6zQD2_0),.clk(gclk));
	jdff dff_A_uSOO17m51_0(.dout(w_dff_A_XpFWsEE17_0),.din(w_dff_A_uSOO17m51_0),.clk(gclk));
	jdff dff_A_XpFWsEE17_0(.dout(w_dff_A_DPFy6FRM4_0),.din(w_dff_A_XpFWsEE17_0),.clk(gclk));
	jdff dff_A_DPFy6FRM4_0(.dout(w_dff_A_tbLsQrJW9_0),.din(w_dff_A_DPFy6FRM4_0),.clk(gclk));
	jdff dff_A_tbLsQrJW9_0(.dout(w_dff_A_DAXSPrcr1_0),.din(w_dff_A_tbLsQrJW9_0),.clk(gclk));
	jdff dff_A_DAXSPrcr1_0(.dout(w_dff_A_Y1x8Pt0Y4_0),.din(w_dff_A_DAXSPrcr1_0),.clk(gclk));
	jdff dff_A_Y1x8Pt0Y4_0(.dout(G602),.din(w_dff_A_Y1x8Pt0Y4_0),.clk(gclk));
	jdff dff_A_kcOoDOTs8_1(.dout(w_dff_A_2DVT02543_0),.din(w_dff_A_kcOoDOTs8_1),.clk(gclk));
	jdff dff_A_2DVT02543_0(.dout(w_dff_A_ZQqX4Lkn5_0),.din(w_dff_A_2DVT02543_0),.clk(gclk));
	jdff dff_A_ZQqX4Lkn5_0(.dout(w_dff_A_Jq4xC4fU9_0),.din(w_dff_A_ZQqX4Lkn5_0),.clk(gclk));
	jdff dff_A_Jq4xC4fU9_0(.dout(w_dff_A_b6NtChoc4_0),.din(w_dff_A_Jq4xC4fU9_0),.clk(gclk));
	jdff dff_A_b6NtChoc4_0(.dout(w_dff_A_XHXmZc7H3_0),.din(w_dff_A_b6NtChoc4_0),.clk(gclk));
	jdff dff_A_XHXmZc7H3_0(.dout(w_dff_A_zPnjCGk42_0),.din(w_dff_A_XHXmZc7H3_0),.clk(gclk));
	jdff dff_A_zPnjCGk42_0(.dout(w_dff_A_7zeZws047_0),.din(w_dff_A_zPnjCGk42_0),.clk(gclk));
	jdff dff_A_7zeZws047_0(.dout(w_dff_A_fsXqtNpA0_0),.din(w_dff_A_7zeZws047_0),.clk(gclk));
	jdff dff_A_fsXqtNpA0_0(.dout(w_dff_A_gAnHUW3u7_0),.din(w_dff_A_fsXqtNpA0_0),.clk(gclk));
	jdff dff_A_gAnHUW3u7_0(.dout(w_dff_A_DmeUCcow5_0),.din(w_dff_A_gAnHUW3u7_0),.clk(gclk));
	jdff dff_A_DmeUCcow5_0(.dout(w_dff_A_2Mu281sQ3_0),.din(w_dff_A_DmeUCcow5_0),.clk(gclk));
	jdff dff_A_2Mu281sQ3_0(.dout(w_dff_A_DbcBmpOW3_0),.din(w_dff_A_2Mu281sQ3_0),.clk(gclk));
	jdff dff_A_DbcBmpOW3_0(.dout(w_dff_A_OjVjaU0Q9_0),.din(w_dff_A_DbcBmpOW3_0),.clk(gclk));
	jdff dff_A_OjVjaU0Q9_0(.dout(w_dff_A_jecQuqw36_0),.din(w_dff_A_OjVjaU0Q9_0),.clk(gclk));
	jdff dff_A_jecQuqw36_0(.dout(w_dff_A_HqIFvB276_0),.din(w_dff_A_jecQuqw36_0),.clk(gclk));
	jdff dff_A_HqIFvB276_0(.dout(w_dff_A_tE3NpQdt1_0),.din(w_dff_A_HqIFvB276_0),.clk(gclk));
	jdff dff_A_tE3NpQdt1_0(.dout(w_dff_A_PwQp3b3Q5_0),.din(w_dff_A_tE3NpQdt1_0),.clk(gclk));
	jdff dff_A_PwQp3b3Q5_0(.dout(w_dff_A_k9yQ1RNl7_0),.din(w_dff_A_PwQp3b3Q5_0),.clk(gclk));
	jdff dff_A_k9yQ1RNl7_0(.dout(w_dff_A_Wm0gzxWe2_0),.din(w_dff_A_k9yQ1RNl7_0),.clk(gclk));
	jdff dff_A_Wm0gzxWe2_0(.dout(w_dff_A_t2Gusbyd9_0),.din(w_dff_A_Wm0gzxWe2_0),.clk(gclk));
	jdff dff_A_t2Gusbyd9_0(.dout(w_dff_A_fwRGXway1_0),.din(w_dff_A_t2Gusbyd9_0),.clk(gclk));
	jdff dff_A_fwRGXway1_0(.dout(w_dff_A_ZH1r2eSj6_0),.din(w_dff_A_fwRGXway1_0),.clk(gclk));
	jdff dff_A_ZH1r2eSj6_0(.dout(w_dff_A_50evll2s5_0),.din(w_dff_A_ZH1r2eSj6_0),.clk(gclk));
	jdff dff_A_50evll2s5_0(.dout(w_dff_A_4LggUN8F5_0),.din(w_dff_A_50evll2s5_0),.clk(gclk));
	jdff dff_A_4LggUN8F5_0(.dout(G603),.din(w_dff_A_4LggUN8F5_0),.clk(gclk));
	jdff dff_A_hDMD60wB6_1(.dout(w_dff_A_BCtwA5XO2_0),.din(w_dff_A_hDMD60wB6_1),.clk(gclk));
	jdff dff_A_BCtwA5XO2_0(.dout(w_dff_A_L27Jgo6W3_0),.din(w_dff_A_BCtwA5XO2_0),.clk(gclk));
	jdff dff_A_L27Jgo6W3_0(.dout(w_dff_A_lKDAFeTZ4_0),.din(w_dff_A_L27Jgo6W3_0),.clk(gclk));
	jdff dff_A_lKDAFeTZ4_0(.dout(w_dff_A_B36YSzB13_0),.din(w_dff_A_lKDAFeTZ4_0),.clk(gclk));
	jdff dff_A_B36YSzB13_0(.dout(w_dff_A_lOCQ4mXJ2_0),.din(w_dff_A_B36YSzB13_0),.clk(gclk));
	jdff dff_A_lOCQ4mXJ2_0(.dout(w_dff_A_zSFbqrLS6_0),.din(w_dff_A_lOCQ4mXJ2_0),.clk(gclk));
	jdff dff_A_zSFbqrLS6_0(.dout(w_dff_A_dqrBGxKs8_0),.din(w_dff_A_zSFbqrLS6_0),.clk(gclk));
	jdff dff_A_dqrBGxKs8_0(.dout(w_dff_A_Yqw9PheB4_0),.din(w_dff_A_dqrBGxKs8_0),.clk(gclk));
	jdff dff_A_Yqw9PheB4_0(.dout(w_dff_A_Azg8u7so6_0),.din(w_dff_A_Yqw9PheB4_0),.clk(gclk));
	jdff dff_A_Azg8u7so6_0(.dout(w_dff_A_dDD3VMX70_0),.din(w_dff_A_Azg8u7so6_0),.clk(gclk));
	jdff dff_A_dDD3VMX70_0(.dout(w_dff_A_PzNrCIkj1_0),.din(w_dff_A_dDD3VMX70_0),.clk(gclk));
	jdff dff_A_PzNrCIkj1_0(.dout(w_dff_A_oAPoFMC03_0),.din(w_dff_A_PzNrCIkj1_0),.clk(gclk));
	jdff dff_A_oAPoFMC03_0(.dout(w_dff_A_UVrokZLl8_0),.din(w_dff_A_oAPoFMC03_0),.clk(gclk));
	jdff dff_A_UVrokZLl8_0(.dout(w_dff_A_HJ6gta4a1_0),.din(w_dff_A_UVrokZLl8_0),.clk(gclk));
	jdff dff_A_HJ6gta4a1_0(.dout(w_dff_A_Mn9BlPf28_0),.din(w_dff_A_HJ6gta4a1_0),.clk(gclk));
	jdff dff_A_Mn9BlPf28_0(.dout(w_dff_A_0jTRirf47_0),.din(w_dff_A_Mn9BlPf28_0),.clk(gclk));
	jdff dff_A_0jTRirf47_0(.dout(w_dff_A_PWTnVoTw6_0),.din(w_dff_A_0jTRirf47_0),.clk(gclk));
	jdff dff_A_PWTnVoTw6_0(.dout(w_dff_A_o3iDkmJj6_0),.din(w_dff_A_PWTnVoTw6_0),.clk(gclk));
	jdff dff_A_o3iDkmJj6_0(.dout(w_dff_A_pvYdX6aT8_0),.din(w_dff_A_o3iDkmJj6_0),.clk(gclk));
	jdff dff_A_pvYdX6aT8_0(.dout(w_dff_A_DwpUNVel8_0),.din(w_dff_A_pvYdX6aT8_0),.clk(gclk));
	jdff dff_A_DwpUNVel8_0(.dout(w_dff_A_leUowjKv2_0),.din(w_dff_A_DwpUNVel8_0),.clk(gclk));
	jdff dff_A_leUowjKv2_0(.dout(w_dff_A_7XJp0Tgc2_0),.din(w_dff_A_leUowjKv2_0),.clk(gclk));
	jdff dff_A_7XJp0Tgc2_0(.dout(w_dff_A_9AvTUtQC3_0),.din(w_dff_A_7XJp0Tgc2_0),.clk(gclk));
	jdff dff_A_9AvTUtQC3_0(.dout(w_dff_A_QAO211s71_0),.din(w_dff_A_9AvTUtQC3_0),.clk(gclk));
	jdff dff_A_QAO211s71_0(.dout(G604),.din(w_dff_A_QAO211s71_0),.clk(gclk));
	jdff dff_A_u0F4vmwG6_1(.dout(w_dff_A_9iV7etma1_0),.din(w_dff_A_u0F4vmwG6_1),.clk(gclk));
	jdff dff_A_9iV7etma1_0(.dout(w_dff_A_xR1CDCiH4_0),.din(w_dff_A_9iV7etma1_0),.clk(gclk));
	jdff dff_A_xR1CDCiH4_0(.dout(w_dff_A_9mkTrHY12_0),.din(w_dff_A_xR1CDCiH4_0),.clk(gclk));
	jdff dff_A_9mkTrHY12_0(.dout(w_dff_A_gWCQvCZl6_0),.din(w_dff_A_9mkTrHY12_0),.clk(gclk));
	jdff dff_A_gWCQvCZl6_0(.dout(w_dff_A_GyU4E6NA8_0),.din(w_dff_A_gWCQvCZl6_0),.clk(gclk));
	jdff dff_A_GyU4E6NA8_0(.dout(w_dff_A_w4vdD8iZ6_0),.din(w_dff_A_GyU4E6NA8_0),.clk(gclk));
	jdff dff_A_w4vdD8iZ6_0(.dout(w_dff_A_6vkkNFpX1_0),.din(w_dff_A_w4vdD8iZ6_0),.clk(gclk));
	jdff dff_A_6vkkNFpX1_0(.dout(w_dff_A_aZqO8c5F7_0),.din(w_dff_A_6vkkNFpX1_0),.clk(gclk));
	jdff dff_A_aZqO8c5F7_0(.dout(w_dff_A_XLjHdiyH6_0),.din(w_dff_A_aZqO8c5F7_0),.clk(gclk));
	jdff dff_A_XLjHdiyH6_0(.dout(w_dff_A_jGsUjMvm1_0),.din(w_dff_A_XLjHdiyH6_0),.clk(gclk));
	jdff dff_A_jGsUjMvm1_0(.dout(w_dff_A_J2f4JC6P8_0),.din(w_dff_A_jGsUjMvm1_0),.clk(gclk));
	jdff dff_A_J2f4JC6P8_0(.dout(w_dff_A_HI9stvvD5_0),.din(w_dff_A_J2f4JC6P8_0),.clk(gclk));
	jdff dff_A_HI9stvvD5_0(.dout(w_dff_A_eUrec72X5_0),.din(w_dff_A_HI9stvvD5_0),.clk(gclk));
	jdff dff_A_eUrec72X5_0(.dout(w_dff_A_g1yjhV022_0),.din(w_dff_A_eUrec72X5_0),.clk(gclk));
	jdff dff_A_g1yjhV022_0(.dout(w_dff_A_IcadDF6t1_0),.din(w_dff_A_g1yjhV022_0),.clk(gclk));
	jdff dff_A_IcadDF6t1_0(.dout(w_dff_A_Q2HGDxci3_0),.din(w_dff_A_IcadDF6t1_0),.clk(gclk));
	jdff dff_A_Q2HGDxci3_0(.dout(w_dff_A_TzHKWsDc2_0),.din(w_dff_A_Q2HGDxci3_0),.clk(gclk));
	jdff dff_A_TzHKWsDc2_0(.dout(w_dff_A_XeaXkH5p3_0),.din(w_dff_A_TzHKWsDc2_0),.clk(gclk));
	jdff dff_A_XeaXkH5p3_0(.dout(w_dff_A_1KQqB91M8_0),.din(w_dff_A_XeaXkH5p3_0),.clk(gclk));
	jdff dff_A_1KQqB91M8_0(.dout(w_dff_A_m0ZEIDAx1_0),.din(w_dff_A_1KQqB91M8_0),.clk(gclk));
	jdff dff_A_m0ZEIDAx1_0(.dout(w_dff_A_nhN7O2Om4_0),.din(w_dff_A_m0ZEIDAx1_0),.clk(gclk));
	jdff dff_A_nhN7O2Om4_0(.dout(w_dff_A_CBXEhqr40_0),.din(w_dff_A_nhN7O2Om4_0),.clk(gclk));
	jdff dff_A_CBXEhqr40_0(.dout(w_dff_A_NlbAecwD3_0),.din(w_dff_A_CBXEhqr40_0),.clk(gclk));
	jdff dff_A_NlbAecwD3_0(.dout(w_dff_A_y4uxC6nd1_0),.din(w_dff_A_NlbAecwD3_0),.clk(gclk));
	jdff dff_A_y4uxC6nd1_0(.dout(G611),.din(w_dff_A_y4uxC6nd1_0),.clk(gclk));
	jdff dff_A_vV76YNP35_1(.dout(w_dff_A_lziMPqTj0_0),.din(w_dff_A_vV76YNP35_1),.clk(gclk));
	jdff dff_A_lziMPqTj0_0(.dout(w_dff_A_5F9DPMfw0_0),.din(w_dff_A_lziMPqTj0_0),.clk(gclk));
	jdff dff_A_5F9DPMfw0_0(.dout(w_dff_A_EBWMsjJe0_0),.din(w_dff_A_5F9DPMfw0_0),.clk(gclk));
	jdff dff_A_EBWMsjJe0_0(.dout(w_dff_A_VT7EMWLc4_0),.din(w_dff_A_EBWMsjJe0_0),.clk(gclk));
	jdff dff_A_VT7EMWLc4_0(.dout(w_dff_A_O5E1qDJi2_0),.din(w_dff_A_VT7EMWLc4_0),.clk(gclk));
	jdff dff_A_O5E1qDJi2_0(.dout(w_dff_A_8qnEGAZC1_0),.din(w_dff_A_O5E1qDJi2_0),.clk(gclk));
	jdff dff_A_8qnEGAZC1_0(.dout(w_dff_A_MQsAG5lq6_0),.din(w_dff_A_8qnEGAZC1_0),.clk(gclk));
	jdff dff_A_MQsAG5lq6_0(.dout(w_dff_A_c6Vsn3OW2_0),.din(w_dff_A_MQsAG5lq6_0),.clk(gclk));
	jdff dff_A_c6Vsn3OW2_0(.dout(w_dff_A_YL86j1d33_0),.din(w_dff_A_c6Vsn3OW2_0),.clk(gclk));
	jdff dff_A_YL86j1d33_0(.dout(w_dff_A_0jrsovDC6_0),.din(w_dff_A_YL86j1d33_0),.clk(gclk));
	jdff dff_A_0jrsovDC6_0(.dout(w_dff_A_L6iIM8QM3_0),.din(w_dff_A_0jrsovDC6_0),.clk(gclk));
	jdff dff_A_L6iIM8QM3_0(.dout(w_dff_A_tKlmUtQS7_0),.din(w_dff_A_L6iIM8QM3_0),.clk(gclk));
	jdff dff_A_tKlmUtQS7_0(.dout(w_dff_A_BpTMQnj98_0),.din(w_dff_A_tKlmUtQS7_0),.clk(gclk));
	jdff dff_A_BpTMQnj98_0(.dout(w_dff_A_KHT5ooBw7_0),.din(w_dff_A_BpTMQnj98_0),.clk(gclk));
	jdff dff_A_KHT5ooBw7_0(.dout(w_dff_A_sx1oMZqH1_0),.din(w_dff_A_KHT5ooBw7_0),.clk(gclk));
	jdff dff_A_sx1oMZqH1_0(.dout(w_dff_A_fci6eniY4_0),.din(w_dff_A_sx1oMZqH1_0),.clk(gclk));
	jdff dff_A_fci6eniY4_0(.dout(w_dff_A_YU9eLELf6_0),.din(w_dff_A_fci6eniY4_0),.clk(gclk));
	jdff dff_A_YU9eLELf6_0(.dout(w_dff_A_T0WxmrKV1_0),.din(w_dff_A_YU9eLELf6_0),.clk(gclk));
	jdff dff_A_T0WxmrKV1_0(.dout(w_dff_A_XgHagHai4_0),.din(w_dff_A_T0WxmrKV1_0),.clk(gclk));
	jdff dff_A_XgHagHai4_0(.dout(w_dff_A_vuCuXbVo5_0),.din(w_dff_A_XgHagHai4_0),.clk(gclk));
	jdff dff_A_vuCuXbVo5_0(.dout(w_dff_A_Cs3hiT9K0_0),.din(w_dff_A_vuCuXbVo5_0),.clk(gclk));
	jdff dff_A_Cs3hiT9K0_0(.dout(w_dff_A_1nJyn9qk6_0),.din(w_dff_A_Cs3hiT9K0_0),.clk(gclk));
	jdff dff_A_1nJyn9qk6_0(.dout(w_dff_A_uD2KJBVk3_0),.din(w_dff_A_1nJyn9qk6_0),.clk(gclk));
	jdff dff_A_uD2KJBVk3_0(.dout(w_dff_A_UOomnUKF3_0),.din(w_dff_A_uD2KJBVk3_0),.clk(gclk));
	jdff dff_A_UOomnUKF3_0(.dout(G612),.din(w_dff_A_UOomnUKF3_0),.clk(gclk));
	jdff dff_A_GlKmi3Mx5_2(.dout(w_dff_A_FoF28rke4_0),.din(w_dff_A_GlKmi3Mx5_2),.clk(gclk));
	jdff dff_A_FoF28rke4_0(.dout(w_dff_A_kc5WQBGy2_0),.din(w_dff_A_FoF28rke4_0),.clk(gclk));
	jdff dff_A_kc5WQBGy2_0(.dout(w_dff_A_LmKqX8Mj9_0),.din(w_dff_A_kc5WQBGy2_0),.clk(gclk));
	jdff dff_A_LmKqX8Mj9_0(.dout(w_dff_A_pGUnQGn94_0),.din(w_dff_A_LmKqX8Mj9_0),.clk(gclk));
	jdff dff_A_pGUnQGn94_0(.dout(w_dff_A_EZegEoFd7_0),.din(w_dff_A_pGUnQGn94_0),.clk(gclk));
	jdff dff_A_EZegEoFd7_0(.dout(w_dff_A_GfQslj0o0_0),.din(w_dff_A_EZegEoFd7_0),.clk(gclk));
	jdff dff_A_GfQslj0o0_0(.dout(w_dff_A_XIFE8IBm9_0),.din(w_dff_A_GfQslj0o0_0),.clk(gclk));
	jdff dff_A_XIFE8IBm9_0(.dout(w_dff_A_tIPzgF7l9_0),.din(w_dff_A_XIFE8IBm9_0),.clk(gclk));
	jdff dff_A_tIPzgF7l9_0(.dout(w_dff_A_wJC5mJQg8_0),.din(w_dff_A_tIPzgF7l9_0),.clk(gclk));
	jdff dff_A_wJC5mJQg8_0(.dout(w_dff_A_b5NydUYV6_0),.din(w_dff_A_wJC5mJQg8_0),.clk(gclk));
	jdff dff_A_b5NydUYV6_0(.dout(w_dff_A_wIskXDYU2_0),.din(w_dff_A_b5NydUYV6_0),.clk(gclk));
	jdff dff_A_wIskXDYU2_0(.dout(w_dff_A_AjpMm4TS2_0),.din(w_dff_A_wIskXDYU2_0),.clk(gclk));
	jdff dff_A_AjpMm4TS2_0(.dout(w_dff_A_l9i4VvN49_0),.din(w_dff_A_AjpMm4TS2_0),.clk(gclk));
	jdff dff_A_l9i4VvN49_0(.dout(w_dff_A_85K5QOOH6_0),.din(w_dff_A_l9i4VvN49_0),.clk(gclk));
	jdff dff_A_85K5QOOH6_0(.dout(w_dff_A_fF3m1NiH2_0),.din(w_dff_A_85K5QOOH6_0),.clk(gclk));
	jdff dff_A_fF3m1NiH2_0(.dout(w_dff_A_Z7MDiG8V9_0),.din(w_dff_A_fF3m1NiH2_0),.clk(gclk));
	jdff dff_A_Z7MDiG8V9_0(.dout(w_dff_A_nR1ZUh5U2_0),.din(w_dff_A_Z7MDiG8V9_0),.clk(gclk));
	jdff dff_A_nR1ZUh5U2_0(.dout(w_dff_A_baKoa0Ig6_0),.din(w_dff_A_nR1ZUh5U2_0),.clk(gclk));
	jdff dff_A_baKoa0Ig6_0(.dout(w_dff_A_Yzmkfj7N6_0),.din(w_dff_A_baKoa0Ig6_0),.clk(gclk));
	jdff dff_A_Yzmkfj7N6_0(.dout(w_dff_A_mQCLBEtB0_0),.din(w_dff_A_Yzmkfj7N6_0),.clk(gclk));
	jdff dff_A_mQCLBEtB0_0(.dout(w_dff_A_Z5MYojyL4_0),.din(w_dff_A_mQCLBEtB0_0),.clk(gclk));
	jdff dff_A_Z5MYojyL4_0(.dout(w_dff_A_qHp9fiAq2_0),.din(w_dff_A_Z5MYojyL4_0),.clk(gclk));
	jdff dff_A_qHp9fiAq2_0(.dout(w_dff_A_ASFLD3OY1_0),.din(w_dff_A_qHp9fiAq2_0),.clk(gclk));
	jdff dff_A_ASFLD3OY1_0(.dout(w_dff_A_b2dglj631_0),.din(w_dff_A_ASFLD3OY1_0),.clk(gclk));
	jdff dff_A_b2dglj631_0(.dout(G810),.din(w_dff_A_b2dglj631_0),.clk(gclk));
	jdff dff_A_xyLwOATF7_1(.dout(w_dff_A_eNvCPr9i4_0),.din(w_dff_A_xyLwOATF7_1),.clk(gclk));
	jdff dff_A_eNvCPr9i4_0(.dout(w_dff_A_8oRD8j3h4_0),.din(w_dff_A_eNvCPr9i4_0),.clk(gclk));
	jdff dff_A_8oRD8j3h4_0(.dout(w_dff_A_ibAyT6ij0_0),.din(w_dff_A_8oRD8j3h4_0),.clk(gclk));
	jdff dff_A_ibAyT6ij0_0(.dout(w_dff_A_vxof0kK68_0),.din(w_dff_A_ibAyT6ij0_0),.clk(gclk));
	jdff dff_A_vxof0kK68_0(.dout(w_dff_A_x7g8EHZc3_0),.din(w_dff_A_vxof0kK68_0),.clk(gclk));
	jdff dff_A_x7g8EHZc3_0(.dout(w_dff_A_pKxM4MRV2_0),.din(w_dff_A_x7g8EHZc3_0),.clk(gclk));
	jdff dff_A_pKxM4MRV2_0(.dout(w_dff_A_nkl7Wo2H5_0),.din(w_dff_A_pKxM4MRV2_0),.clk(gclk));
	jdff dff_A_nkl7Wo2H5_0(.dout(w_dff_A_hpLOQV0C5_0),.din(w_dff_A_nkl7Wo2H5_0),.clk(gclk));
	jdff dff_A_hpLOQV0C5_0(.dout(w_dff_A_Nyq8fd0V1_0),.din(w_dff_A_hpLOQV0C5_0),.clk(gclk));
	jdff dff_A_Nyq8fd0V1_0(.dout(w_dff_A_WsWtyNfe4_0),.din(w_dff_A_Nyq8fd0V1_0),.clk(gclk));
	jdff dff_A_WsWtyNfe4_0(.dout(w_dff_A_10sVEysO1_0),.din(w_dff_A_WsWtyNfe4_0),.clk(gclk));
	jdff dff_A_10sVEysO1_0(.dout(w_dff_A_MKWPLyAp1_0),.din(w_dff_A_10sVEysO1_0),.clk(gclk));
	jdff dff_A_MKWPLyAp1_0(.dout(w_dff_A_WkFiKJKM7_0),.din(w_dff_A_MKWPLyAp1_0),.clk(gclk));
	jdff dff_A_WkFiKJKM7_0(.dout(w_dff_A_JhzUAlvL1_0),.din(w_dff_A_WkFiKJKM7_0),.clk(gclk));
	jdff dff_A_JhzUAlvL1_0(.dout(w_dff_A_mGg9XuzS9_0),.din(w_dff_A_JhzUAlvL1_0),.clk(gclk));
	jdff dff_A_mGg9XuzS9_0(.dout(w_dff_A_6sR7H9hy4_0),.din(w_dff_A_mGg9XuzS9_0),.clk(gclk));
	jdff dff_A_6sR7H9hy4_0(.dout(w_dff_A_CrtDy2rj8_0),.din(w_dff_A_6sR7H9hy4_0),.clk(gclk));
	jdff dff_A_CrtDy2rj8_0(.dout(w_dff_A_Ng0nP9Pz8_0),.din(w_dff_A_CrtDy2rj8_0),.clk(gclk));
	jdff dff_A_Ng0nP9Pz8_0(.dout(w_dff_A_m95qoQ9p1_0),.din(w_dff_A_Ng0nP9Pz8_0),.clk(gclk));
	jdff dff_A_m95qoQ9p1_0(.dout(w_dff_A_dh9HbEoW8_0),.din(w_dff_A_m95qoQ9p1_0),.clk(gclk));
	jdff dff_A_dh9HbEoW8_0(.dout(w_dff_A_hCYOeZJR5_0),.din(w_dff_A_dh9HbEoW8_0),.clk(gclk));
	jdff dff_A_hCYOeZJR5_0(.dout(w_dff_A_tJcdIU2f8_0),.din(w_dff_A_hCYOeZJR5_0),.clk(gclk));
	jdff dff_A_tJcdIU2f8_0(.dout(w_dff_A_RW53ZOK86_0),.din(w_dff_A_tJcdIU2f8_0),.clk(gclk));
	jdff dff_A_RW53ZOK86_0(.dout(w_dff_A_ZsI0AaUQ5_0),.din(w_dff_A_RW53ZOK86_0),.clk(gclk));
	jdff dff_A_ZsI0AaUQ5_0(.dout(G848),.din(w_dff_A_ZsI0AaUQ5_0),.clk(gclk));
	jdff dff_A_H8rH6ICZ3_1(.dout(w_dff_A_nOtMmBbK9_0),.din(w_dff_A_H8rH6ICZ3_1),.clk(gclk));
	jdff dff_A_nOtMmBbK9_0(.dout(w_dff_A_OtbwNwYB6_0),.din(w_dff_A_nOtMmBbK9_0),.clk(gclk));
	jdff dff_A_OtbwNwYB6_0(.dout(w_dff_A_2khSAweJ4_0),.din(w_dff_A_OtbwNwYB6_0),.clk(gclk));
	jdff dff_A_2khSAweJ4_0(.dout(w_dff_A_dyVsIhlv3_0),.din(w_dff_A_2khSAweJ4_0),.clk(gclk));
	jdff dff_A_dyVsIhlv3_0(.dout(w_dff_A_oDPWNfAa3_0),.din(w_dff_A_dyVsIhlv3_0),.clk(gclk));
	jdff dff_A_oDPWNfAa3_0(.dout(w_dff_A_gQMW51AI1_0),.din(w_dff_A_oDPWNfAa3_0),.clk(gclk));
	jdff dff_A_gQMW51AI1_0(.dout(w_dff_A_HPcxssCH8_0),.din(w_dff_A_gQMW51AI1_0),.clk(gclk));
	jdff dff_A_HPcxssCH8_0(.dout(w_dff_A_bMNuzee73_0),.din(w_dff_A_HPcxssCH8_0),.clk(gclk));
	jdff dff_A_bMNuzee73_0(.dout(w_dff_A_musNaZm99_0),.din(w_dff_A_bMNuzee73_0),.clk(gclk));
	jdff dff_A_musNaZm99_0(.dout(w_dff_A_I9eo0zv08_0),.din(w_dff_A_musNaZm99_0),.clk(gclk));
	jdff dff_A_I9eo0zv08_0(.dout(w_dff_A_Y9g00JQ24_0),.din(w_dff_A_I9eo0zv08_0),.clk(gclk));
	jdff dff_A_Y9g00JQ24_0(.dout(w_dff_A_z0mWXjxE3_0),.din(w_dff_A_Y9g00JQ24_0),.clk(gclk));
	jdff dff_A_z0mWXjxE3_0(.dout(w_dff_A_CImKJKok4_0),.din(w_dff_A_z0mWXjxE3_0),.clk(gclk));
	jdff dff_A_CImKJKok4_0(.dout(w_dff_A_VaSZNCj75_0),.din(w_dff_A_CImKJKok4_0),.clk(gclk));
	jdff dff_A_VaSZNCj75_0(.dout(w_dff_A_WHcI2w6f8_0),.din(w_dff_A_VaSZNCj75_0),.clk(gclk));
	jdff dff_A_WHcI2w6f8_0(.dout(w_dff_A_GqwwfeYl1_0),.din(w_dff_A_WHcI2w6f8_0),.clk(gclk));
	jdff dff_A_GqwwfeYl1_0(.dout(w_dff_A_TRjxx3Lq9_0),.din(w_dff_A_GqwwfeYl1_0),.clk(gclk));
	jdff dff_A_TRjxx3Lq9_0(.dout(w_dff_A_cZa8AnBW9_0),.din(w_dff_A_TRjxx3Lq9_0),.clk(gclk));
	jdff dff_A_cZa8AnBW9_0(.dout(w_dff_A_pqDlsAvc7_0),.din(w_dff_A_cZa8AnBW9_0),.clk(gclk));
	jdff dff_A_pqDlsAvc7_0(.dout(w_dff_A_kzcHeqM82_0),.din(w_dff_A_pqDlsAvc7_0),.clk(gclk));
	jdff dff_A_kzcHeqM82_0(.dout(w_dff_A_goHCHCuz3_0),.din(w_dff_A_kzcHeqM82_0),.clk(gclk));
	jdff dff_A_goHCHCuz3_0(.dout(w_dff_A_CdK5SyKL2_0),.din(w_dff_A_goHCHCuz3_0),.clk(gclk));
	jdff dff_A_CdK5SyKL2_0(.dout(w_dff_A_akEnMZTu2_0),.din(w_dff_A_CdK5SyKL2_0),.clk(gclk));
	jdff dff_A_akEnMZTu2_0(.dout(w_dff_A_bRKOe4wl6_0),.din(w_dff_A_akEnMZTu2_0),.clk(gclk));
	jdff dff_A_bRKOe4wl6_0(.dout(G849),.din(w_dff_A_bRKOe4wl6_0),.clk(gclk));
	jdff dff_A_Xusarkiy7_1(.dout(w_dff_A_hrBPrJ3k4_0),.din(w_dff_A_Xusarkiy7_1),.clk(gclk));
	jdff dff_A_hrBPrJ3k4_0(.dout(w_dff_A_aaPWOIIu8_0),.din(w_dff_A_hrBPrJ3k4_0),.clk(gclk));
	jdff dff_A_aaPWOIIu8_0(.dout(w_dff_A_werb8YnI4_0),.din(w_dff_A_aaPWOIIu8_0),.clk(gclk));
	jdff dff_A_werb8YnI4_0(.dout(w_dff_A_mYezHKSE6_0),.din(w_dff_A_werb8YnI4_0),.clk(gclk));
	jdff dff_A_mYezHKSE6_0(.dout(w_dff_A_vvgoF3Lp1_0),.din(w_dff_A_mYezHKSE6_0),.clk(gclk));
	jdff dff_A_vvgoF3Lp1_0(.dout(w_dff_A_S60DZFUn0_0),.din(w_dff_A_vvgoF3Lp1_0),.clk(gclk));
	jdff dff_A_S60DZFUn0_0(.dout(w_dff_A_IoM7ebW96_0),.din(w_dff_A_S60DZFUn0_0),.clk(gclk));
	jdff dff_A_IoM7ebW96_0(.dout(w_dff_A_hNOh6rtH1_0),.din(w_dff_A_IoM7ebW96_0),.clk(gclk));
	jdff dff_A_hNOh6rtH1_0(.dout(w_dff_A_YuxYtkDv0_0),.din(w_dff_A_hNOh6rtH1_0),.clk(gclk));
	jdff dff_A_YuxYtkDv0_0(.dout(w_dff_A_JmG6gYIf4_0),.din(w_dff_A_YuxYtkDv0_0),.clk(gclk));
	jdff dff_A_JmG6gYIf4_0(.dout(w_dff_A_MRP53ePZ5_0),.din(w_dff_A_JmG6gYIf4_0),.clk(gclk));
	jdff dff_A_MRP53ePZ5_0(.dout(w_dff_A_BzvS1uvv3_0),.din(w_dff_A_MRP53ePZ5_0),.clk(gclk));
	jdff dff_A_BzvS1uvv3_0(.dout(w_dff_A_icKZ0k6n3_0),.din(w_dff_A_BzvS1uvv3_0),.clk(gclk));
	jdff dff_A_icKZ0k6n3_0(.dout(w_dff_A_LNQpHKrV1_0),.din(w_dff_A_icKZ0k6n3_0),.clk(gclk));
	jdff dff_A_LNQpHKrV1_0(.dout(w_dff_A_GZAhTFVz3_0),.din(w_dff_A_LNQpHKrV1_0),.clk(gclk));
	jdff dff_A_GZAhTFVz3_0(.dout(w_dff_A_uNsXvIKA0_0),.din(w_dff_A_GZAhTFVz3_0),.clk(gclk));
	jdff dff_A_uNsXvIKA0_0(.dout(w_dff_A_8IQsyxm79_0),.din(w_dff_A_uNsXvIKA0_0),.clk(gclk));
	jdff dff_A_8IQsyxm79_0(.dout(w_dff_A_3qu5WyOD6_0),.din(w_dff_A_8IQsyxm79_0),.clk(gclk));
	jdff dff_A_3qu5WyOD6_0(.dout(w_dff_A_JcX9TJoS0_0),.din(w_dff_A_3qu5WyOD6_0),.clk(gclk));
	jdff dff_A_JcX9TJoS0_0(.dout(w_dff_A_i4BeRQuP4_0),.din(w_dff_A_JcX9TJoS0_0),.clk(gclk));
	jdff dff_A_i4BeRQuP4_0(.dout(w_dff_A_JRIPggxw5_0),.din(w_dff_A_i4BeRQuP4_0),.clk(gclk));
	jdff dff_A_JRIPggxw5_0(.dout(w_dff_A_4QOfRiWB4_0),.din(w_dff_A_JRIPggxw5_0),.clk(gclk));
	jdff dff_A_4QOfRiWB4_0(.dout(w_dff_A_X1jHTkfH9_0),.din(w_dff_A_4QOfRiWB4_0),.clk(gclk));
	jdff dff_A_X1jHTkfH9_0(.dout(w_dff_A_MxEkLznI2_0),.din(w_dff_A_X1jHTkfH9_0),.clk(gclk));
	jdff dff_A_MxEkLznI2_0(.dout(G850),.din(w_dff_A_MxEkLznI2_0),.clk(gclk));
	jdff dff_A_pmLPKsfd4_1(.dout(w_dff_A_suFphxG97_0),.din(w_dff_A_pmLPKsfd4_1),.clk(gclk));
	jdff dff_A_suFphxG97_0(.dout(w_dff_A_lOTGBhQ59_0),.din(w_dff_A_suFphxG97_0),.clk(gclk));
	jdff dff_A_lOTGBhQ59_0(.dout(w_dff_A_lgW7zxz77_0),.din(w_dff_A_lOTGBhQ59_0),.clk(gclk));
	jdff dff_A_lgW7zxz77_0(.dout(w_dff_A_1wEnSzqF5_0),.din(w_dff_A_lgW7zxz77_0),.clk(gclk));
	jdff dff_A_1wEnSzqF5_0(.dout(w_dff_A_CeNpf4TS3_0),.din(w_dff_A_1wEnSzqF5_0),.clk(gclk));
	jdff dff_A_CeNpf4TS3_0(.dout(w_dff_A_J1Bvu7ZZ0_0),.din(w_dff_A_CeNpf4TS3_0),.clk(gclk));
	jdff dff_A_J1Bvu7ZZ0_0(.dout(w_dff_A_g5njZi7L8_0),.din(w_dff_A_J1Bvu7ZZ0_0),.clk(gclk));
	jdff dff_A_g5njZi7L8_0(.dout(w_dff_A_ik80OX237_0),.din(w_dff_A_g5njZi7L8_0),.clk(gclk));
	jdff dff_A_ik80OX237_0(.dout(w_dff_A_PLfaf77S1_0),.din(w_dff_A_ik80OX237_0),.clk(gclk));
	jdff dff_A_PLfaf77S1_0(.dout(w_dff_A_9GR8uVrz7_0),.din(w_dff_A_PLfaf77S1_0),.clk(gclk));
	jdff dff_A_9GR8uVrz7_0(.dout(w_dff_A_1KyUeUtZ2_0),.din(w_dff_A_9GR8uVrz7_0),.clk(gclk));
	jdff dff_A_1KyUeUtZ2_0(.dout(w_dff_A_euXqnPdk9_0),.din(w_dff_A_1KyUeUtZ2_0),.clk(gclk));
	jdff dff_A_euXqnPdk9_0(.dout(w_dff_A_RQvKvLTV1_0),.din(w_dff_A_euXqnPdk9_0),.clk(gclk));
	jdff dff_A_RQvKvLTV1_0(.dout(w_dff_A_zEYokS6w1_0),.din(w_dff_A_RQvKvLTV1_0),.clk(gclk));
	jdff dff_A_zEYokS6w1_0(.dout(w_dff_A_iyIxatti8_0),.din(w_dff_A_zEYokS6w1_0),.clk(gclk));
	jdff dff_A_iyIxatti8_0(.dout(w_dff_A_gTrcipWg2_0),.din(w_dff_A_iyIxatti8_0),.clk(gclk));
	jdff dff_A_gTrcipWg2_0(.dout(w_dff_A_ixKCXnwZ3_0),.din(w_dff_A_gTrcipWg2_0),.clk(gclk));
	jdff dff_A_ixKCXnwZ3_0(.dout(w_dff_A_MVwL5dF71_0),.din(w_dff_A_ixKCXnwZ3_0),.clk(gclk));
	jdff dff_A_MVwL5dF71_0(.dout(w_dff_A_BjiThJyY8_0),.din(w_dff_A_MVwL5dF71_0),.clk(gclk));
	jdff dff_A_BjiThJyY8_0(.dout(w_dff_A_GyPH7zPK1_0),.din(w_dff_A_BjiThJyY8_0),.clk(gclk));
	jdff dff_A_GyPH7zPK1_0(.dout(w_dff_A_0nUYBNEz8_0),.din(w_dff_A_GyPH7zPK1_0),.clk(gclk));
	jdff dff_A_0nUYBNEz8_0(.dout(w_dff_A_D8IQuX735_0),.din(w_dff_A_0nUYBNEz8_0),.clk(gclk));
	jdff dff_A_D8IQuX735_0(.dout(w_dff_A_BnMfACOa4_0),.din(w_dff_A_D8IQuX735_0),.clk(gclk));
	jdff dff_A_BnMfACOa4_0(.dout(w_dff_A_pAd7P8mQ8_0),.din(w_dff_A_BnMfACOa4_0),.clk(gclk));
	jdff dff_A_pAd7P8mQ8_0(.dout(G851),.din(w_dff_A_pAd7P8mQ8_0),.clk(gclk));
	jdff dff_A_RYNJc9DE7_2(.dout(w_dff_A_K0Gp274N1_0),.din(w_dff_A_RYNJc9DE7_2),.clk(gclk));
	jdff dff_A_K0Gp274N1_0(.dout(w_dff_A_MPy72eiW4_0),.din(w_dff_A_K0Gp274N1_0),.clk(gclk));
	jdff dff_A_MPy72eiW4_0(.dout(w_dff_A_LvSJJ4uN7_0),.din(w_dff_A_MPy72eiW4_0),.clk(gclk));
	jdff dff_A_LvSJJ4uN7_0(.dout(w_dff_A_PicTrorG4_0),.din(w_dff_A_LvSJJ4uN7_0),.clk(gclk));
	jdff dff_A_PicTrorG4_0(.dout(w_dff_A_bJmFwyF66_0),.din(w_dff_A_PicTrorG4_0),.clk(gclk));
	jdff dff_A_bJmFwyF66_0(.dout(w_dff_A_kK0Iytzo9_0),.din(w_dff_A_bJmFwyF66_0),.clk(gclk));
	jdff dff_A_kK0Iytzo9_0(.dout(w_dff_A_7HUGsfuw3_0),.din(w_dff_A_kK0Iytzo9_0),.clk(gclk));
	jdff dff_A_7HUGsfuw3_0(.dout(w_dff_A_zoTMS6al2_0),.din(w_dff_A_7HUGsfuw3_0),.clk(gclk));
	jdff dff_A_zoTMS6al2_0(.dout(w_dff_A_5Tikg5i43_0),.din(w_dff_A_zoTMS6al2_0),.clk(gclk));
	jdff dff_A_5Tikg5i43_0(.dout(w_dff_A_eYqwXIcD6_0),.din(w_dff_A_5Tikg5i43_0),.clk(gclk));
	jdff dff_A_eYqwXIcD6_0(.dout(w_dff_A_Am5Z8qri4_0),.din(w_dff_A_eYqwXIcD6_0),.clk(gclk));
	jdff dff_A_Am5Z8qri4_0(.dout(w_dff_A_k5QkWKsX2_0),.din(w_dff_A_Am5Z8qri4_0),.clk(gclk));
	jdff dff_A_k5QkWKsX2_0(.dout(w_dff_A_nQB22ICq8_0),.din(w_dff_A_k5QkWKsX2_0),.clk(gclk));
	jdff dff_A_nQB22ICq8_0(.dout(w_dff_A_ErQaohi93_0),.din(w_dff_A_nQB22ICq8_0),.clk(gclk));
	jdff dff_A_ErQaohi93_0(.dout(w_dff_A_DF8xFxXn1_0),.din(w_dff_A_ErQaohi93_0),.clk(gclk));
	jdff dff_A_DF8xFxXn1_0(.dout(w_dff_A_PBoDfIGd6_0),.din(w_dff_A_DF8xFxXn1_0),.clk(gclk));
	jdff dff_A_PBoDfIGd6_0(.dout(w_dff_A_BuOOO1na7_0),.din(w_dff_A_PBoDfIGd6_0),.clk(gclk));
	jdff dff_A_BuOOO1na7_0(.dout(w_dff_A_V9mPnqth7_0),.din(w_dff_A_BuOOO1na7_0),.clk(gclk));
	jdff dff_A_V9mPnqth7_0(.dout(w_dff_A_44bQQigm3_0),.din(w_dff_A_V9mPnqth7_0),.clk(gclk));
	jdff dff_A_44bQQigm3_0(.dout(w_dff_A_gdzRynCj5_0),.din(w_dff_A_44bQQigm3_0),.clk(gclk));
	jdff dff_A_gdzRynCj5_0(.dout(w_dff_A_1EuwGAOE6_0),.din(w_dff_A_gdzRynCj5_0),.clk(gclk));
	jdff dff_A_1EuwGAOE6_0(.dout(w_dff_A_V2pChiko1_0),.din(w_dff_A_1EuwGAOE6_0),.clk(gclk));
	jdff dff_A_V2pChiko1_0(.dout(w_dff_A_xMavVPiU9_0),.din(w_dff_A_V2pChiko1_0),.clk(gclk));
	jdff dff_A_xMavVPiU9_0(.dout(w_dff_A_usp0TRLn9_0),.din(w_dff_A_xMavVPiU9_0),.clk(gclk));
	jdff dff_A_usp0TRLn9_0(.dout(G634),.din(w_dff_A_usp0TRLn9_0),.clk(gclk));
	jdff dff_A_yXw8OWlh0_2(.dout(w_dff_A_6jWmU8vg1_0),.din(w_dff_A_yXw8OWlh0_2),.clk(gclk));
	jdff dff_A_6jWmU8vg1_0(.dout(w_dff_A_bF6tchFU2_0),.din(w_dff_A_6jWmU8vg1_0),.clk(gclk));
	jdff dff_A_bF6tchFU2_0(.dout(w_dff_A_9iJdGgTj6_0),.din(w_dff_A_bF6tchFU2_0),.clk(gclk));
	jdff dff_A_9iJdGgTj6_0(.dout(w_dff_A_8LdQTxzS7_0),.din(w_dff_A_9iJdGgTj6_0),.clk(gclk));
	jdff dff_A_8LdQTxzS7_0(.dout(w_dff_A_0eLUeaiW9_0),.din(w_dff_A_8LdQTxzS7_0),.clk(gclk));
	jdff dff_A_0eLUeaiW9_0(.dout(w_dff_A_Ceyaryv07_0),.din(w_dff_A_0eLUeaiW9_0),.clk(gclk));
	jdff dff_A_Ceyaryv07_0(.dout(w_dff_A_Ubbj64qM5_0),.din(w_dff_A_Ceyaryv07_0),.clk(gclk));
	jdff dff_A_Ubbj64qM5_0(.dout(w_dff_A_79uyTPsg2_0),.din(w_dff_A_Ubbj64qM5_0),.clk(gclk));
	jdff dff_A_79uyTPsg2_0(.dout(w_dff_A_GZgr1Pdm2_0),.din(w_dff_A_79uyTPsg2_0),.clk(gclk));
	jdff dff_A_GZgr1Pdm2_0(.dout(w_dff_A_MYrR1AiH1_0),.din(w_dff_A_GZgr1Pdm2_0),.clk(gclk));
	jdff dff_A_MYrR1AiH1_0(.dout(w_dff_A_LYcd1Qc95_0),.din(w_dff_A_MYrR1AiH1_0),.clk(gclk));
	jdff dff_A_LYcd1Qc95_0(.dout(w_dff_A_sUhUoX0H5_0),.din(w_dff_A_LYcd1Qc95_0),.clk(gclk));
	jdff dff_A_sUhUoX0H5_0(.dout(w_dff_A_ad0N5twf0_0),.din(w_dff_A_sUhUoX0H5_0),.clk(gclk));
	jdff dff_A_ad0N5twf0_0(.dout(w_dff_A_sVhWGoNO2_0),.din(w_dff_A_ad0N5twf0_0),.clk(gclk));
	jdff dff_A_sVhWGoNO2_0(.dout(w_dff_A_QY3ozO4E2_0),.din(w_dff_A_sVhWGoNO2_0),.clk(gclk));
	jdff dff_A_QY3ozO4E2_0(.dout(w_dff_A_V66hZaVM6_0),.din(w_dff_A_QY3ozO4E2_0),.clk(gclk));
	jdff dff_A_V66hZaVM6_0(.dout(w_dff_A_r2go5Xi55_0),.din(w_dff_A_V66hZaVM6_0),.clk(gclk));
	jdff dff_A_r2go5Xi55_0(.dout(w_dff_A_2gr0sy7n1_0),.din(w_dff_A_r2go5Xi55_0),.clk(gclk));
	jdff dff_A_2gr0sy7n1_0(.dout(w_dff_A_xLR3sFmw6_0),.din(w_dff_A_2gr0sy7n1_0),.clk(gclk));
	jdff dff_A_xLR3sFmw6_0(.dout(w_dff_A_BwEWsH041_0),.din(w_dff_A_xLR3sFmw6_0),.clk(gclk));
	jdff dff_A_BwEWsH041_0(.dout(w_dff_A_H1QIBT7v8_0),.din(w_dff_A_BwEWsH041_0),.clk(gclk));
	jdff dff_A_H1QIBT7v8_0(.dout(w_dff_A_mJNNPMaw0_0),.din(w_dff_A_H1QIBT7v8_0),.clk(gclk));
	jdff dff_A_mJNNPMaw0_0(.dout(w_dff_A_ve09drHw3_0),.din(w_dff_A_mJNNPMaw0_0),.clk(gclk));
	jdff dff_A_ve09drHw3_0(.dout(G815),.din(w_dff_A_ve09drHw3_0),.clk(gclk));
	jdff dff_A_QrS0w1hc9_2(.dout(w_dff_A_v0R7cT3A2_0),.din(w_dff_A_QrS0w1hc9_2),.clk(gclk));
	jdff dff_A_v0R7cT3A2_0(.dout(w_dff_A_qnf4sQky6_0),.din(w_dff_A_v0R7cT3A2_0),.clk(gclk));
	jdff dff_A_qnf4sQky6_0(.dout(w_dff_A_Kb0UWdzr6_0),.din(w_dff_A_qnf4sQky6_0),.clk(gclk));
	jdff dff_A_Kb0UWdzr6_0(.dout(w_dff_A_fmGQrk6p4_0),.din(w_dff_A_Kb0UWdzr6_0),.clk(gclk));
	jdff dff_A_fmGQrk6p4_0(.dout(w_dff_A_v0Xaxmzn5_0),.din(w_dff_A_fmGQrk6p4_0),.clk(gclk));
	jdff dff_A_v0Xaxmzn5_0(.dout(w_dff_A_DeGVkzQk2_0),.din(w_dff_A_v0Xaxmzn5_0),.clk(gclk));
	jdff dff_A_DeGVkzQk2_0(.dout(w_dff_A_JVSjm7gC7_0),.din(w_dff_A_DeGVkzQk2_0),.clk(gclk));
	jdff dff_A_JVSjm7gC7_0(.dout(w_dff_A_wV771ojw7_0),.din(w_dff_A_JVSjm7gC7_0),.clk(gclk));
	jdff dff_A_wV771ojw7_0(.dout(w_dff_A_cauunzu24_0),.din(w_dff_A_wV771ojw7_0),.clk(gclk));
	jdff dff_A_cauunzu24_0(.dout(w_dff_A_eFetDvas1_0),.din(w_dff_A_cauunzu24_0),.clk(gclk));
	jdff dff_A_eFetDvas1_0(.dout(w_dff_A_Vf76mOl43_0),.din(w_dff_A_eFetDvas1_0),.clk(gclk));
	jdff dff_A_Vf76mOl43_0(.dout(w_dff_A_WsAz6DbW6_0),.din(w_dff_A_Vf76mOl43_0),.clk(gclk));
	jdff dff_A_WsAz6DbW6_0(.dout(w_dff_A_7XNVSPDS9_0),.din(w_dff_A_WsAz6DbW6_0),.clk(gclk));
	jdff dff_A_7XNVSPDS9_0(.dout(w_dff_A_DFSGgDvy2_0),.din(w_dff_A_7XNVSPDS9_0),.clk(gclk));
	jdff dff_A_DFSGgDvy2_0(.dout(w_dff_A_BLedsIhK0_0),.din(w_dff_A_DFSGgDvy2_0),.clk(gclk));
	jdff dff_A_BLedsIhK0_0(.dout(w_dff_A_inFCm5b98_0),.din(w_dff_A_BLedsIhK0_0),.clk(gclk));
	jdff dff_A_inFCm5b98_0(.dout(w_dff_A_L10plpC43_0),.din(w_dff_A_inFCm5b98_0),.clk(gclk));
	jdff dff_A_L10plpC43_0(.dout(w_dff_A_Xx8EgXT19_0),.din(w_dff_A_L10plpC43_0),.clk(gclk));
	jdff dff_A_Xx8EgXT19_0(.dout(w_dff_A_STM1ZcFU2_0),.din(w_dff_A_Xx8EgXT19_0),.clk(gclk));
	jdff dff_A_STM1ZcFU2_0(.dout(w_dff_A_jc5rUWe24_0),.din(w_dff_A_STM1ZcFU2_0),.clk(gclk));
	jdff dff_A_jc5rUWe24_0(.dout(w_dff_A_NiTD0wdi5_0),.din(w_dff_A_jc5rUWe24_0),.clk(gclk));
	jdff dff_A_NiTD0wdi5_0(.dout(w_dff_A_dDlBSleA7_0),.din(w_dff_A_NiTD0wdi5_0),.clk(gclk));
	jdff dff_A_dDlBSleA7_0(.dout(w_dff_A_khFgEntc2_0),.din(w_dff_A_dDlBSleA7_0),.clk(gclk));
	jdff dff_A_khFgEntc2_0(.dout(G845),.din(w_dff_A_khFgEntc2_0),.clk(gclk));
	jdff dff_A_LSvafEGP1_1(.dout(w_dff_A_YQv15aTr9_0),.din(w_dff_A_LSvafEGP1_1),.clk(gclk));
	jdff dff_A_YQv15aTr9_0(.dout(w_dff_A_8OrmuQq63_0),.din(w_dff_A_YQv15aTr9_0),.clk(gclk));
	jdff dff_A_8OrmuQq63_0(.dout(w_dff_A_hSOEr44i2_0),.din(w_dff_A_8OrmuQq63_0),.clk(gclk));
	jdff dff_A_hSOEr44i2_0(.dout(w_dff_A_yIVB93VL1_0),.din(w_dff_A_hSOEr44i2_0),.clk(gclk));
	jdff dff_A_yIVB93VL1_0(.dout(w_dff_A_SKCuxarp6_0),.din(w_dff_A_yIVB93VL1_0),.clk(gclk));
	jdff dff_A_SKCuxarp6_0(.dout(w_dff_A_1wO0lHia8_0),.din(w_dff_A_SKCuxarp6_0),.clk(gclk));
	jdff dff_A_1wO0lHia8_0(.dout(w_dff_A_BLaFsW7q7_0),.din(w_dff_A_1wO0lHia8_0),.clk(gclk));
	jdff dff_A_BLaFsW7q7_0(.dout(w_dff_A_TeVbRD8X4_0),.din(w_dff_A_BLaFsW7q7_0),.clk(gclk));
	jdff dff_A_TeVbRD8X4_0(.dout(w_dff_A_IUuOibde7_0),.din(w_dff_A_TeVbRD8X4_0),.clk(gclk));
	jdff dff_A_IUuOibde7_0(.dout(w_dff_A_mR1x8Z0y0_0),.din(w_dff_A_IUuOibde7_0),.clk(gclk));
	jdff dff_A_mR1x8Z0y0_0(.dout(w_dff_A_Au8xFoSx1_0),.din(w_dff_A_mR1x8Z0y0_0),.clk(gclk));
	jdff dff_A_Au8xFoSx1_0(.dout(w_dff_A_LnQZhrv18_0),.din(w_dff_A_Au8xFoSx1_0),.clk(gclk));
	jdff dff_A_LnQZhrv18_0(.dout(w_dff_A_5VicGoJH0_0),.din(w_dff_A_LnQZhrv18_0),.clk(gclk));
	jdff dff_A_5VicGoJH0_0(.dout(w_dff_A_tkRk2qtZ4_0),.din(w_dff_A_5VicGoJH0_0),.clk(gclk));
	jdff dff_A_tkRk2qtZ4_0(.dout(w_dff_A_Sk04FQP71_0),.din(w_dff_A_tkRk2qtZ4_0),.clk(gclk));
	jdff dff_A_Sk04FQP71_0(.dout(w_dff_A_30QA9Yde5_0),.din(w_dff_A_Sk04FQP71_0),.clk(gclk));
	jdff dff_A_30QA9Yde5_0(.dout(w_dff_A_1XokZoC53_0),.din(w_dff_A_30QA9Yde5_0),.clk(gclk));
	jdff dff_A_1XokZoC53_0(.dout(w_dff_A_WT4Cl0NM0_0),.din(w_dff_A_1XokZoC53_0),.clk(gclk));
	jdff dff_A_WT4Cl0NM0_0(.dout(w_dff_A_CcE17NJy0_0),.din(w_dff_A_WT4Cl0NM0_0),.clk(gclk));
	jdff dff_A_CcE17NJy0_0(.dout(w_dff_A_OsiQXJQo9_0),.din(w_dff_A_CcE17NJy0_0),.clk(gclk));
	jdff dff_A_OsiQXJQo9_0(.dout(w_dff_A_zXP9mh6c1_0),.din(w_dff_A_OsiQXJQo9_0),.clk(gclk));
	jdff dff_A_zXP9mh6c1_0(.dout(w_dff_A_qCE6IiTW5_0),.din(w_dff_A_zXP9mh6c1_0),.clk(gclk));
	jdff dff_A_qCE6IiTW5_0(.dout(w_dff_A_ekCsCMJB8_0),.din(w_dff_A_qCE6IiTW5_0),.clk(gclk));
	jdff dff_A_ekCsCMJB8_0(.dout(G847),.din(w_dff_A_ekCsCMJB8_0),.clk(gclk));
	jdff dff_A_01NRIr0n5_1(.dout(w_dff_A_T0KCI0Br3_0),.din(w_dff_A_01NRIr0n5_1),.clk(gclk));
	jdff dff_A_T0KCI0Br3_0(.dout(w_dff_A_JIqo6lAF5_0),.din(w_dff_A_T0KCI0Br3_0),.clk(gclk));
	jdff dff_A_JIqo6lAF5_0(.dout(w_dff_A_HAOSnCqu0_0),.din(w_dff_A_JIqo6lAF5_0),.clk(gclk));
	jdff dff_A_HAOSnCqu0_0(.dout(w_dff_A_lJbLgato8_0),.din(w_dff_A_HAOSnCqu0_0),.clk(gclk));
	jdff dff_A_lJbLgato8_0(.dout(w_dff_A_QgPb02XW2_0),.din(w_dff_A_lJbLgato8_0),.clk(gclk));
	jdff dff_A_QgPb02XW2_0(.dout(w_dff_A_bPrzDpx25_0),.din(w_dff_A_QgPb02XW2_0),.clk(gclk));
	jdff dff_A_bPrzDpx25_0(.dout(w_dff_A_HZEVDcEq9_0),.din(w_dff_A_bPrzDpx25_0),.clk(gclk));
	jdff dff_A_HZEVDcEq9_0(.dout(w_dff_A_tKnN1aix3_0),.din(w_dff_A_HZEVDcEq9_0),.clk(gclk));
	jdff dff_A_tKnN1aix3_0(.dout(w_dff_A_oJlQzsHm4_0),.din(w_dff_A_tKnN1aix3_0),.clk(gclk));
	jdff dff_A_oJlQzsHm4_0(.dout(w_dff_A_quIB8Cb39_0),.din(w_dff_A_oJlQzsHm4_0),.clk(gclk));
	jdff dff_A_quIB8Cb39_0(.dout(w_dff_A_pazK6p7m6_0),.din(w_dff_A_quIB8Cb39_0),.clk(gclk));
	jdff dff_A_pazK6p7m6_0(.dout(w_dff_A_zXBOdUVV8_0),.din(w_dff_A_pazK6p7m6_0),.clk(gclk));
	jdff dff_A_zXBOdUVV8_0(.dout(w_dff_A_y4fXJ6dx2_0),.din(w_dff_A_zXBOdUVV8_0),.clk(gclk));
	jdff dff_A_y4fXJ6dx2_0(.dout(w_dff_A_C3vpuTLt0_0),.din(w_dff_A_y4fXJ6dx2_0),.clk(gclk));
	jdff dff_A_C3vpuTLt0_0(.dout(w_dff_A_l9MOsyXH0_0),.din(w_dff_A_C3vpuTLt0_0),.clk(gclk));
	jdff dff_A_l9MOsyXH0_0(.dout(w_dff_A_mnOm5jxk3_0),.din(w_dff_A_l9MOsyXH0_0),.clk(gclk));
	jdff dff_A_mnOm5jxk3_0(.dout(w_dff_A_vDZEMzXW4_0),.din(w_dff_A_mnOm5jxk3_0),.clk(gclk));
	jdff dff_A_vDZEMzXW4_0(.dout(w_dff_A_2EtgvZrm1_0),.din(w_dff_A_vDZEMzXW4_0),.clk(gclk));
	jdff dff_A_2EtgvZrm1_0(.dout(w_dff_A_GjBOM3mV0_0),.din(w_dff_A_2EtgvZrm1_0),.clk(gclk));
	jdff dff_A_GjBOM3mV0_0(.dout(w_dff_A_2jLytp936_0),.din(w_dff_A_GjBOM3mV0_0),.clk(gclk));
	jdff dff_A_2jLytp936_0(.dout(w_dff_A_Vz8iP4Hr0_0),.din(w_dff_A_2jLytp936_0),.clk(gclk));
	jdff dff_A_Vz8iP4Hr0_0(.dout(w_dff_A_o86rQLXx9_0),.din(w_dff_A_Vz8iP4Hr0_0),.clk(gclk));
	jdff dff_A_o86rQLXx9_0(.dout(w_dff_A_UB2FYZMP8_0),.din(w_dff_A_o86rQLXx9_0),.clk(gclk));
	jdff dff_A_UB2FYZMP8_0(.dout(w_dff_A_YnJ1tJzk2_0),.din(w_dff_A_UB2FYZMP8_0),.clk(gclk));
	jdff dff_A_YnJ1tJzk2_0(.dout(w_dff_A_pRwshihh7_0),.din(w_dff_A_YnJ1tJzk2_0),.clk(gclk));
	jdff dff_A_pRwshihh7_0(.dout(G926),.din(w_dff_A_pRwshihh7_0),.clk(gclk));
	jdff dff_A_BnnZ8yRL2_1(.dout(w_dff_A_1EQsAT453_0),.din(w_dff_A_BnnZ8yRL2_1),.clk(gclk));
	jdff dff_A_1EQsAT453_0(.dout(w_dff_A_QCNTUIu25_0),.din(w_dff_A_1EQsAT453_0),.clk(gclk));
	jdff dff_A_QCNTUIu25_0(.dout(w_dff_A_oWBKiZVp8_0),.din(w_dff_A_QCNTUIu25_0),.clk(gclk));
	jdff dff_A_oWBKiZVp8_0(.dout(w_dff_A_BYFycvHY6_0),.din(w_dff_A_oWBKiZVp8_0),.clk(gclk));
	jdff dff_A_BYFycvHY6_0(.dout(w_dff_A_V0026irJ5_0),.din(w_dff_A_BYFycvHY6_0),.clk(gclk));
	jdff dff_A_V0026irJ5_0(.dout(w_dff_A_jdCPur5z9_0),.din(w_dff_A_V0026irJ5_0),.clk(gclk));
	jdff dff_A_jdCPur5z9_0(.dout(w_dff_A_XhD97bkX3_0),.din(w_dff_A_jdCPur5z9_0),.clk(gclk));
	jdff dff_A_XhD97bkX3_0(.dout(w_dff_A_piGLnmpn8_0),.din(w_dff_A_XhD97bkX3_0),.clk(gclk));
	jdff dff_A_piGLnmpn8_0(.dout(w_dff_A_Kgi0SGy95_0),.din(w_dff_A_piGLnmpn8_0),.clk(gclk));
	jdff dff_A_Kgi0SGy95_0(.dout(w_dff_A_SJYGjweE5_0),.din(w_dff_A_Kgi0SGy95_0),.clk(gclk));
	jdff dff_A_SJYGjweE5_0(.dout(w_dff_A_VYbr9uzs3_0),.din(w_dff_A_SJYGjweE5_0),.clk(gclk));
	jdff dff_A_VYbr9uzs3_0(.dout(w_dff_A_PKCIma1I4_0),.din(w_dff_A_VYbr9uzs3_0),.clk(gclk));
	jdff dff_A_PKCIma1I4_0(.dout(w_dff_A_lqCx9CMD5_0),.din(w_dff_A_PKCIma1I4_0),.clk(gclk));
	jdff dff_A_lqCx9CMD5_0(.dout(w_dff_A_bjgza2BL2_0),.din(w_dff_A_lqCx9CMD5_0),.clk(gclk));
	jdff dff_A_bjgza2BL2_0(.dout(w_dff_A_IEAjRMro8_0),.din(w_dff_A_bjgza2BL2_0),.clk(gclk));
	jdff dff_A_IEAjRMro8_0(.dout(w_dff_A_Ba2UnCps9_0),.din(w_dff_A_IEAjRMro8_0),.clk(gclk));
	jdff dff_A_Ba2UnCps9_0(.dout(w_dff_A_YElEShL60_0),.din(w_dff_A_Ba2UnCps9_0),.clk(gclk));
	jdff dff_A_YElEShL60_0(.dout(w_dff_A_dFSTVjYn2_0),.din(w_dff_A_YElEShL60_0),.clk(gclk));
	jdff dff_A_dFSTVjYn2_0(.dout(w_dff_A_AYz8fusT0_0),.din(w_dff_A_dFSTVjYn2_0),.clk(gclk));
	jdff dff_A_AYz8fusT0_0(.dout(w_dff_A_TY7K932o2_0),.din(w_dff_A_AYz8fusT0_0),.clk(gclk));
	jdff dff_A_TY7K932o2_0(.dout(w_dff_A_CPD6Efrp8_0),.din(w_dff_A_TY7K932o2_0),.clk(gclk));
	jdff dff_A_CPD6Efrp8_0(.dout(w_dff_A_hpefC9ae1_0),.din(w_dff_A_CPD6Efrp8_0),.clk(gclk));
	jdff dff_A_hpefC9ae1_0(.dout(w_dff_A_0zIeliN32_0),.din(w_dff_A_hpefC9ae1_0),.clk(gclk));
	jdff dff_A_0zIeliN32_0(.dout(w_dff_A_ZDS7IzTM6_0),.din(w_dff_A_0zIeliN32_0),.clk(gclk));
	jdff dff_A_ZDS7IzTM6_0(.dout(w_dff_A_DaHO4N7T2_0),.din(w_dff_A_ZDS7IzTM6_0),.clk(gclk));
	jdff dff_A_DaHO4N7T2_0(.dout(G923),.din(w_dff_A_DaHO4N7T2_0),.clk(gclk));
	jdff dff_A_Lh3AxbIW3_1(.dout(w_dff_A_ImlrT97C3_0),.din(w_dff_A_Lh3AxbIW3_1),.clk(gclk));
	jdff dff_A_ImlrT97C3_0(.dout(w_dff_A_SCYZ5BkE7_0),.din(w_dff_A_ImlrT97C3_0),.clk(gclk));
	jdff dff_A_SCYZ5BkE7_0(.dout(w_dff_A_qSgrRCIc4_0),.din(w_dff_A_SCYZ5BkE7_0),.clk(gclk));
	jdff dff_A_qSgrRCIc4_0(.dout(w_dff_A_a5YIGvpc7_0),.din(w_dff_A_qSgrRCIc4_0),.clk(gclk));
	jdff dff_A_a5YIGvpc7_0(.dout(w_dff_A_NxQ5Bbpb9_0),.din(w_dff_A_a5YIGvpc7_0),.clk(gclk));
	jdff dff_A_NxQ5Bbpb9_0(.dout(w_dff_A_MmIiKObK2_0),.din(w_dff_A_NxQ5Bbpb9_0),.clk(gclk));
	jdff dff_A_MmIiKObK2_0(.dout(w_dff_A_avlQfnii2_0),.din(w_dff_A_MmIiKObK2_0),.clk(gclk));
	jdff dff_A_avlQfnii2_0(.dout(w_dff_A_iAhmQvPT1_0),.din(w_dff_A_avlQfnii2_0),.clk(gclk));
	jdff dff_A_iAhmQvPT1_0(.dout(w_dff_A_Tq5F952u4_0),.din(w_dff_A_iAhmQvPT1_0),.clk(gclk));
	jdff dff_A_Tq5F952u4_0(.dout(w_dff_A_mSSI74u32_0),.din(w_dff_A_Tq5F952u4_0),.clk(gclk));
	jdff dff_A_mSSI74u32_0(.dout(w_dff_A_qF0E5Cdl7_0),.din(w_dff_A_mSSI74u32_0),.clk(gclk));
	jdff dff_A_qF0E5Cdl7_0(.dout(w_dff_A_W6LOQr1W9_0),.din(w_dff_A_qF0E5Cdl7_0),.clk(gclk));
	jdff dff_A_W6LOQr1W9_0(.dout(w_dff_A_b3VcpK2n0_0),.din(w_dff_A_W6LOQr1W9_0),.clk(gclk));
	jdff dff_A_b3VcpK2n0_0(.dout(w_dff_A_b3CdZCJ50_0),.din(w_dff_A_b3VcpK2n0_0),.clk(gclk));
	jdff dff_A_b3CdZCJ50_0(.dout(w_dff_A_mroB81Cj5_0),.din(w_dff_A_b3CdZCJ50_0),.clk(gclk));
	jdff dff_A_mroB81Cj5_0(.dout(w_dff_A_nhVwgCod1_0),.din(w_dff_A_mroB81Cj5_0),.clk(gclk));
	jdff dff_A_nhVwgCod1_0(.dout(w_dff_A_UNby12XJ2_0),.din(w_dff_A_nhVwgCod1_0),.clk(gclk));
	jdff dff_A_UNby12XJ2_0(.dout(w_dff_A_VFkGOxeG0_0),.din(w_dff_A_UNby12XJ2_0),.clk(gclk));
	jdff dff_A_VFkGOxeG0_0(.dout(w_dff_A_f71d8YOX5_0),.din(w_dff_A_VFkGOxeG0_0),.clk(gclk));
	jdff dff_A_f71d8YOX5_0(.dout(w_dff_A_d4u2VCCL9_0),.din(w_dff_A_f71d8YOX5_0),.clk(gclk));
	jdff dff_A_d4u2VCCL9_0(.dout(w_dff_A_ks86YvjL4_0),.din(w_dff_A_d4u2VCCL9_0),.clk(gclk));
	jdff dff_A_ks86YvjL4_0(.dout(w_dff_A_6ASGuWde8_0),.din(w_dff_A_ks86YvjL4_0),.clk(gclk));
	jdff dff_A_6ASGuWde8_0(.dout(w_dff_A_wugflzAV7_0),.din(w_dff_A_6ASGuWde8_0),.clk(gclk));
	jdff dff_A_wugflzAV7_0(.dout(w_dff_A_QZ6xIBF59_0),.din(w_dff_A_wugflzAV7_0),.clk(gclk));
	jdff dff_A_QZ6xIBF59_0(.dout(w_dff_A_MPSd35nE2_0),.din(w_dff_A_QZ6xIBF59_0),.clk(gclk));
	jdff dff_A_MPSd35nE2_0(.dout(G921),.din(w_dff_A_MPSd35nE2_0),.clk(gclk));
	jdff dff_A_J5XkOm3N6_1(.dout(w_dff_A_myOflQGG3_0),.din(w_dff_A_J5XkOm3N6_1),.clk(gclk));
	jdff dff_A_myOflQGG3_0(.dout(w_dff_A_FOQwnEDt2_0),.din(w_dff_A_myOflQGG3_0),.clk(gclk));
	jdff dff_A_FOQwnEDt2_0(.dout(w_dff_A_xs7nUafR2_0),.din(w_dff_A_FOQwnEDt2_0),.clk(gclk));
	jdff dff_A_xs7nUafR2_0(.dout(w_dff_A_88eakqhA7_0),.din(w_dff_A_xs7nUafR2_0),.clk(gclk));
	jdff dff_A_88eakqhA7_0(.dout(w_dff_A_lpmANb3k2_0),.din(w_dff_A_88eakqhA7_0),.clk(gclk));
	jdff dff_A_lpmANb3k2_0(.dout(w_dff_A_so9lmTyb8_0),.din(w_dff_A_lpmANb3k2_0),.clk(gclk));
	jdff dff_A_so9lmTyb8_0(.dout(w_dff_A_Z5jBZ53w8_0),.din(w_dff_A_so9lmTyb8_0),.clk(gclk));
	jdff dff_A_Z5jBZ53w8_0(.dout(w_dff_A_uT4eruv50_0),.din(w_dff_A_Z5jBZ53w8_0),.clk(gclk));
	jdff dff_A_uT4eruv50_0(.dout(w_dff_A_1EBmzuvu6_0),.din(w_dff_A_uT4eruv50_0),.clk(gclk));
	jdff dff_A_1EBmzuvu6_0(.dout(w_dff_A_Pjrjv0Rx3_0),.din(w_dff_A_1EBmzuvu6_0),.clk(gclk));
	jdff dff_A_Pjrjv0Rx3_0(.dout(w_dff_A_gDSMpamd6_0),.din(w_dff_A_Pjrjv0Rx3_0),.clk(gclk));
	jdff dff_A_gDSMpamd6_0(.dout(w_dff_A_YGtJp68q5_0),.din(w_dff_A_gDSMpamd6_0),.clk(gclk));
	jdff dff_A_YGtJp68q5_0(.dout(w_dff_A_fTe3itQ76_0),.din(w_dff_A_YGtJp68q5_0),.clk(gclk));
	jdff dff_A_fTe3itQ76_0(.dout(w_dff_A_BTTZFMKc3_0),.din(w_dff_A_fTe3itQ76_0),.clk(gclk));
	jdff dff_A_BTTZFMKc3_0(.dout(w_dff_A_BXhTVqsY9_0),.din(w_dff_A_BTTZFMKc3_0),.clk(gclk));
	jdff dff_A_BXhTVqsY9_0(.dout(w_dff_A_mMNki7lP1_0),.din(w_dff_A_BXhTVqsY9_0),.clk(gclk));
	jdff dff_A_mMNki7lP1_0(.dout(w_dff_A_MvxY6Iah0_0),.din(w_dff_A_mMNki7lP1_0),.clk(gclk));
	jdff dff_A_MvxY6Iah0_0(.dout(w_dff_A_FRRRTgtz2_0),.din(w_dff_A_MvxY6Iah0_0),.clk(gclk));
	jdff dff_A_FRRRTgtz2_0(.dout(w_dff_A_wxG9MtEi6_0),.din(w_dff_A_FRRRTgtz2_0),.clk(gclk));
	jdff dff_A_wxG9MtEi6_0(.dout(w_dff_A_y74yrhsH9_0),.din(w_dff_A_wxG9MtEi6_0),.clk(gclk));
	jdff dff_A_y74yrhsH9_0(.dout(w_dff_A_lwAAOZ8e9_0),.din(w_dff_A_y74yrhsH9_0),.clk(gclk));
	jdff dff_A_lwAAOZ8e9_0(.dout(w_dff_A_HuiI7CWG0_0),.din(w_dff_A_lwAAOZ8e9_0),.clk(gclk));
	jdff dff_A_HuiI7CWG0_0(.dout(w_dff_A_2mFCOca89_0),.din(w_dff_A_HuiI7CWG0_0),.clk(gclk));
	jdff dff_A_2mFCOca89_0(.dout(w_dff_A_ta3JEm181_0),.din(w_dff_A_2mFCOca89_0),.clk(gclk));
	jdff dff_A_ta3JEm181_0(.dout(w_dff_A_yKxRKaqF8_0),.din(w_dff_A_ta3JEm181_0),.clk(gclk));
	jdff dff_A_yKxRKaqF8_0(.dout(G892),.din(w_dff_A_yKxRKaqF8_0),.clk(gclk));
	jdff dff_A_DyvXlmRo5_1(.dout(w_dff_A_tLXdturw1_0),.din(w_dff_A_DyvXlmRo5_1),.clk(gclk));
	jdff dff_A_tLXdturw1_0(.dout(w_dff_A_3hodUwyi5_0),.din(w_dff_A_tLXdturw1_0),.clk(gclk));
	jdff dff_A_3hodUwyi5_0(.dout(w_dff_A_ZwlNl2494_0),.din(w_dff_A_3hodUwyi5_0),.clk(gclk));
	jdff dff_A_ZwlNl2494_0(.dout(w_dff_A_sn0h8oOY2_0),.din(w_dff_A_ZwlNl2494_0),.clk(gclk));
	jdff dff_A_sn0h8oOY2_0(.dout(w_dff_A_QnKjVoYS2_0),.din(w_dff_A_sn0h8oOY2_0),.clk(gclk));
	jdff dff_A_QnKjVoYS2_0(.dout(w_dff_A_ORld5hr40_0),.din(w_dff_A_QnKjVoYS2_0),.clk(gclk));
	jdff dff_A_ORld5hr40_0(.dout(w_dff_A_wffqNnzy9_0),.din(w_dff_A_ORld5hr40_0),.clk(gclk));
	jdff dff_A_wffqNnzy9_0(.dout(w_dff_A_knN7M2ZI9_0),.din(w_dff_A_wffqNnzy9_0),.clk(gclk));
	jdff dff_A_knN7M2ZI9_0(.dout(w_dff_A_h2AQVlxP7_0),.din(w_dff_A_knN7M2ZI9_0),.clk(gclk));
	jdff dff_A_h2AQVlxP7_0(.dout(w_dff_A_3EPTT3hI8_0),.din(w_dff_A_h2AQVlxP7_0),.clk(gclk));
	jdff dff_A_3EPTT3hI8_0(.dout(w_dff_A_V0VRm04v5_0),.din(w_dff_A_3EPTT3hI8_0),.clk(gclk));
	jdff dff_A_V0VRm04v5_0(.dout(w_dff_A_WyWQ5rCf3_0),.din(w_dff_A_V0VRm04v5_0),.clk(gclk));
	jdff dff_A_WyWQ5rCf3_0(.dout(w_dff_A_xFHIHZRf1_0),.din(w_dff_A_WyWQ5rCf3_0),.clk(gclk));
	jdff dff_A_xFHIHZRf1_0(.dout(w_dff_A_09qoeox29_0),.din(w_dff_A_xFHIHZRf1_0),.clk(gclk));
	jdff dff_A_09qoeox29_0(.dout(w_dff_A_6EqdFl8v8_0),.din(w_dff_A_09qoeox29_0),.clk(gclk));
	jdff dff_A_6EqdFl8v8_0(.dout(w_dff_A_qW2PdEIs8_0),.din(w_dff_A_6EqdFl8v8_0),.clk(gclk));
	jdff dff_A_qW2PdEIs8_0(.dout(w_dff_A_1b82hlNA8_0),.din(w_dff_A_qW2PdEIs8_0),.clk(gclk));
	jdff dff_A_1b82hlNA8_0(.dout(w_dff_A_tO5O59357_0),.din(w_dff_A_1b82hlNA8_0),.clk(gclk));
	jdff dff_A_tO5O59357_0(.dout(w_dff_A_ZHPBeITe7_0),.din(w_dff_A_tO5O59357_0),.clk(gclk));
	jdff dff_A_ZHPBeITe7_0(.dout(w_dff_A_h04npl922_0),.din(w_dff_A_ZHPBeITe7_0),.clk(gclk));
	jdff dff_A_h04npl922_0(.dout(w_dff_A_jfQCWTci0_0),.din(w_dff_A_h04npl922_0),.clk(gclk));
	jdff dff_A_jfQCWTci0_0(.dout(w_dff_A_Rgsvvq4d7_0),.din(w_dff_A_jfQCWTci0_0),.clk(gclk));
	jdff dff_A_Rgsvvq4d7_0(.dout(w_dff_A_fMpYah1y6_0),.din(w_dff_A_Rgsvvq4d7_0),.clk(gclk));
	jdff dff_A_fMpYah1y6_0(.dout(w_dff_A_9vSzsBJX8_0),.din(w_dff_A_fMpYah1y6_0),.clk(gclk));
	jdff dff_A_9vSzsBJX8_0(.dout(w_dff_A_bEhDIrq66_0),.din(w_dff_A_9vSzsBJX8_0),.clk(gclk));
	jdff dff_A_bEhDIrq66_0(.dout(G887),.din(w_dff_A_bEhDIrq66_0),.clk(gclk));
	jdff dff_A_nvgG7fE58_1(.dout(w_dff_A_N3hu5bC12_0),.din(w_dff_A_nvgG7fE58_1),.clk(gclk));
	jdff dff_A_N3hu5bC12_0(.dout(w_dff_A_KPOicwMq5_0),.din(w_dff_A_N3hu5bC12_0),.clk(gclk));
	jdff dff_A_KPOicwMq5_0(.dout(w_dff_A_OCKymEXB1_0),.din(w_dff_A_KPOicwMq5_0),.clk(gclk));
	jdff dff_A_OCKymEXB1_0(.dout(w_dff_A_ucdGveD86_0),.din(w_dff_A_OCKymEXB1_0),.clk(gclk));
	jdff dff_A_ucdGveD86_0(.dout(w_dff_A_bXE7E3GN4_0),.din(w_dff_A_ucdGveD86_0),.clk(gclk));
	jdff dff_A_bXE7E3GN4_0(.dout(w_dff_A_Txy0aA5D9_0),.din(w_dff_A_bXE7E3GN4_0),.clk(gclk));
	jdff dff_A_Txy0aA5D9_0(.dout(w_dff_A_2U2VnnSb3_0),.din(w_dff_A_Txy0aA5D9_0),.clk(gclk));
	jdff dff_A_2U2VnnSb3_0(.dout(w_dff_A_zFLFNVP43_0),.din(w_dff_A_2U2VnnSb3_0),.clk(gclk));
	jdff dff_A_zFLFNVP43_0(.dout(w_dff_A_452iNvR68_0),.din(w_dff_A_zFLFNVP43_0),.clk(gclk));
	jdff dff_A_452iNvR68_0(.dout(w_dff_A_Qm3VKH1a3_0),.din(w_dff_A_452iNvR68_0),.clk(gclk));
	jdff dff_A_Qm3VKH1a3_0(.dout(w_dff_A_MRj4ygRT9_0),.din(w_dff_A_Qm3VKH1a3_0),.clk(gclk));
	jdff dff_A_MRj4ygRT9_0(.dout(w_dff_A_fiZrchch4_0),.din(w_dff_A_MRj4ygRT9_0),.clk(gclk));
	jdff dff_A_fiZrchch4_0(.dout(w_dff_A_3kIM8ibh6_0),.din(w_dff_A_fiZrchch4_0),.clk(gclk));
	jdff dff_A_3kIM8ibh6_0(.dout(w_dff_A_AVLyIPyA1_0),.din(w_dff_A_3kIM8ibh6_0),.clk(gclk));
	jdff dff_A_AVLyIPyA1_0(.dout(w_dff_A_S0LhnmTs7_0),.din(w_dff_A_AVLyIPyA1_0),.clk(gclk));
	jdff dff_A_S0LhnmTs7_0(.dout(w_dff_A_3dkV0ct89_0),.din(w_dff_A_S0LhnmTs7_0),.clk(gclk));
	jdff dff_A_3dkV0ct89_0(.dout(w_dff_A_JWLLaUqB4_0),.din(w_dff_A_3dkV0ct89_0),.clk(gclk));
	jdff dff_A_JWLLaUqB4_0(.dout(w_dff_A_4JLrEYuS9_0),.din(w_dff_A_JWLLaUqB4_0),.clk(gclk));
	jdff dff_A_4JLrEYuS9_0(.dout(w_dff_A_Lrjjx16v3_0),.din(w_dff_A_4JLrEYuS9_0),.clk(gclk));
	jdff dff_A_Lrjjx16v3_0(.dout(w_dff_A_IeJ6ryVi6_0),.din(w_dff_A_Lrjjx16v3_0),.clk(gclk));
	jdff dff_A_IeJ6ryVi6_0(.dout(w_dff_A_ZJFFcWwp6_0),.din(w_dff_A_IeJ6ryVi6_0),.clk(gclk));
	jdff dff_A_ZJFFcWwp6_0(.dout(w_dff_A_SZ3yWRj41_0),.din(w_dff_A_ZJFFcWwp6_0),.clk(gclk));
	jdff dff_A_SZ3yWRj41_0(.dout(w_dff_A_J6zAg7lC5_0),.din(w_dff_A_SZ3yWRj41_0),.clk(gclk));
	jdff dff_A_J6zAg7lC5_0(.dout(w_dff_A_cNWvPRCi8_0),.din(w_dff_A_J6zAg7lC5_0),.clk(gclk));
	jdff dff_A_cNWvPRCi8_0(.dout(G606),.din(w_dff_A_cNWvPRCi8_0),.clk(gclk));
	jdff dff_A_dtpCUlzB5_2(.dout(w_dff_A_5Eh2GO9F2_0),.din(w_dff_A_dtpCUlzB5_2),.clk(gclk));
	jdff dff_A_5Eh2GO9F2_0(.dout(w_dff_A_3suHmsej5_0),.din(w_dff_A_5Eh2GO9F2_0),.clk(gclk));
	jdff dff_A_3suHmsej5_0(.dout(w_dff_A_ksBNEb8g7_0),.din(w_dff_A_3suHmsej5_0),.clk(gclk));
	jdff dff_A_ksBNEb8g7_0(.dout(w_dff_A_tJNslEAo5_0),.din(w_dff_A_ksBNEb8g7_0),.clk(gclk));
	jdff dff_A_tJNslEAo5_0(.dout(w_dff_A_niiULae75_0),.din(w_dff_A_tJNslEAo5_0),.clk(gclk));
	jdff dff_A_niiULae75_0(.dout(w_dff_A_ZexcCbco4_0),.din(w_dff_A_niiULae75_0),.clk(gclk));
	jdff dff_A_ZexcCbco4_0(.dout(w_dff_A_c8l4WoxB8_0),.din(w_dff_A_ZexcCbco4_0),.clk(gclk));
	jdff dff_A_c8l4WoxB8_0(.dout(w_dff_A_QXxPXL2C1_0),.din(w_dff_A_c8l4WoxB8_0),.clk(gclk));
	jdff dff_A_QXxPXL2C1_0(.dout(w_dff_A_1LWx9mDd8_0),.din(w_dff_A_QXxPXL2C1_0),.clk(gclk));
	jdff dff_A_1LWx9mDd8_0(.dout(w_dff_A_DfgroJEz6_0),.din(w_dff_A_1LWx9mDd8_0),.clk(gclk));
	jdff dff_A_DfgroJEz6_0(.dout(w_dff_A_OXozIfOx0_0),.din(w_dff_A_DfgroJEz6_0),.clk(gclk));
	jdff dff_A_OXozIfOx0_0(.dout(w_dff_A_DQsS3MaV7_0),.din(w_dff_A_OXozIfOx0_0),.clk(gclk));
	jdff dff_A_DQsS3MaV7_0(.dout(w_dff_A_3C9QpG8a6_0),.din(w_dff_A_DQsS3MaV7_0),.clk(gclk));
	jdff dff_A_3C9QpG8a6_0(.dout(w_dff_A_J4ZLPBDi8_0),.din(w_dff_A_3C9QpG8a6_0),.clk(gclk));
	jdff dff_A_J4ZLPBDi8_0(.dout(w_dff_A_EjPBXT596_0),.din(w_dff_A_J4ZLPBDi8_0),.clk(gclk));
	jdff dff_A_EjPBXT596_0(.dout(w_dff_A_LnaG41ak7_0),.din(w_dff_A_EjPBXT596_0),.clk(gclk));
	jdff dff_A_LnaG41ak7_0(.dout(w_dff_A_Q1XUl7WF2_0),.din(w_dff_A_LnaG41ak7_0),.clk(gclk));
	jdff dff_A_Q1XUl7WF2_0(.dout(w_dff_A_kvcSJhn63_0),.din(w_dff_A_Q1XUl7WF2_0),.clk(gclk));
	jdff dff_A_kvcSJhn63_0(.dout(w_dff_A_3YyCJeWj3_0),.din(w_dff_A_kvcSJhn63_0),.clk(gclk));
	jdff dff_A_3YyCJeWj3_0(.dout(w_dff_A_tpObOz4f2_0),.din(w_dff_A_3YyCJeWj3_0),.clk(gclk));
	jdff dff_A_tpObOz4f2_0(.dout(w_dff_A_CGMV944R3_0),.din(w_dff_A_tpObOz4f2_0),.clk(gclk));
	jdff dff_A_CGMV944R3_0(.dout(w_dff_A_akhxLudq6_0),.din(w_dff_A_CGMV944R3_0),.clk(gclk));
	jdff dff_A_akhxLudq6_0(.dout(G656),.din(w_dff_A_akhxLudq6_0),.clk(gclk));
	jdff dff_A_Wkcf8uO35_2(.dout(w_dff_A_nVQkj7KY2_0),.din(w_dff_A_Wkcf8uO35_2),.clk(gclk));
	jdff dff_A_nVQkj7KY2_0(.dout(w_dff_A_XrIZB1W39_0),.din(w_dff_A_nVQkj7KY2_0),.clk(gclk));
	jdff dff_A_XrIZB1W39_0(.dout(w_dff_A_2RAvaipf5_0),.din(w_dff_A_XrIZB1W39_0),.clk(gclk));
	jdff dff_A_2RAvaipf5_0(.dout(w_dff_A_L5qTC1Tz5_0),.din(w_dff_A_2RAvaipf5_0),.clk(gclk));
	jdff dff_A_L5qTC1Tz5_0(.dout(w_dff_A_tkrlteuN8_0),.din(w_dff_A_L5qTC1Tz5_0),.clk(gclk));
	jdff dff_A_tkrlteuN8_0(.dout(w_dff_A_PjIRoYcv5_0),.din(w_dff_A_tkrlteuN8_0),.clk(gclk));
	jdff dff_A_PjIRoYcv5_0(.dout(w_dff_A_PXAjyjue2_0),.din(w_dff_A_PjIRoYcv5_0),.clk(gclk));
	jdff dff_A_PXAjyjue2_0(.dout(w_dff_A_bQtcwnco8_0),.din(w_dff_A_PXAjyjue2_0),.clk(gclk));
	jdff dff_A_bQtcwnco8_0(.dout(w_dff_A_1xfS7pJG0_0),.din(w_dff_A_bQtcwnco8_0),.clk(gclk));
	jdff dff_A_1xfS7pJG0_0(.dout(w_dff_A_iC1qYZAI9_0),.din(w_dff_A_1xfS7pJG0_0),.clk(gclk));
	jdff dff_A_iC1qYZAI9_0(.dout(w_dff_A_RvJEUfeB5_0),.din(w_dff_A_iC1qYZAI9_0),.clk(gclk));
	jdff dff_A_RvJEUfeB5_0(.dout(w_dff_A_4ECh9uD13_0),.din(w_dff_A_RvJEUfeB5_0),.clk(gclk));
	jdff dff_A_4ECh9uD13_0(.dout(w_dff_A_i0x8pCV67_0),.din(w_dff_A_4ECh9uD13_0),.clk(gclk));
	jdff dff_A_i0x8pCV67_0(.dout(w_dff_A_azu69xyF1_0),.din(w_dff_A_i0x8pCV67_0),.clk(gclk));
	jdff dff_A_azu69xyF1_0(.dout(w_dff_A_ge2p8Y7j5_0),.din(w_dff_A_azu69xyF1_0),.clk(gclk));
	jdff dff_A_ge2p8Y7j5_0(.dout(w_dff_A_WtbNT1NZ1_0),.din(w_dff_A_ge2p8Y7j5_0),.clk(gclk));
	jdff dff_A_WtbNT1NZ1_0(.dout(w_dff_A_uRqDqbqv6_0),.din(w_dff_A_WtbNT1NZ1_0),.clk(gclk));
	jdff dff_A_uRqDqbqv6_0(.dout(w_dff_A_AmbNLimM7_0),.din(w_dff_A_uRqDqbqv6_0),.clk(gclk));
	jdff dff_A_AmbNLimM7_0(.dout(w_dff_A_7Jy3zYRO0_0),.din(w_dff_A_AmbNLimM7_0),.clk(gclk));
	jdff dff_A_7Jy3zYRO0_0(.dout(w_dff_A_H2s2XOom2_0),.din(w_dff_A_7Jy3zYRO0_0),.clk(gclk));
	jdff dff_A_H2s2XOom2_0(.dout(w_dff_A_61abACHB9_0),.din(w_dff_A_H2s2XOom2_0),.clk(gclk));
	jdff dff_A_61abACHB9_0(.dout(w_dff_A_BJ2ZWDW55_0),.din(w_dff_A_61abACHB9_0),.clk(gclk));
	jdff dff_A_BJ2ZWDW55_0(.dout(w_dff_A_4AybJTNt1_0),.din(w_dff_A_BJ2ZWDW55_0),.clk(gclk));
	jdff dff_A_4AybJTNt1_0(.dout(G809),.din(w_dff_A_4AybJTNt1_0),.clk(gclk));
	jdff dff_A_cVuHOXky3_1(.dout(w_dff_A_oNXFHuPE6_0),.din(w_dff_A_cVuHOXky3_1),.clk(gclk));
	jdff dff_A_oNXFHuPE6_0(.dout(w_dff_A_MkyAEXfM5_0),.din(w_dff_A_oNXFHuPE6_0),.clk(gclk));
	jdff dff_A_MkyAEXfM5_0(.dout(w_dff_A_wbm6SpU57_0),.din(w_dff_A_MkyAEXfM5_0),.clk(gclk));
	jdff dff_A_wbm6SpU57_0(.dout(w_dff_A_GEQHmbgQ0_0),.din(w_dff_A_wbm6SpU57_0),.clk(gclk));
	jdff dff_A_GEQHmbgQ0_0(.dout(w_dff_A_oaA25qda8_0),.din(w_dff_A_GEQHmbgQ0_0),.clk(gclk));
	jdff dff_A_oaA25qda8_0(.dout(w_dff_A_DaZs9uKh2_0),.din(w_dff_A_oaA25qda8_0),.clk(gclk));
	jdff dff_A_DaZs9uKh2_0(.dout(w_dff_A_U9NpTuD58_0),.din(w_dff_A_DaZs9uKh2_0),.clk(gclk));
	jdff dff_A_U9NpTuD58_0(.dout(w_dff_A_zK3GZtg69_0),.din(w_dff_A_U9NpTuD58_0),.clk(gclk));
	jdff dff_A_zK3GZtg69_0(.dout(w_dff_A_4WNNsVql6_0),.din(w_dff_A_zK3GZtg69_0),.clk(gclk));
	jdff dff_A_4WNNsVql6_0(.dout(w_dff_A_m5YsQizm3_0),.din(w_dff_A_4WNNsVql6_0),.clk(gclk));
	jdff dff_A_m5YsQizm3_0(.dout(w_dff_A_l7ISEKSu8_0),.din(w_dff_A_m5YsQizm3_0),.clk(gclk));
	jdff dff_A_l7ISEKSu8_0(.dout(w_dff_A_OtdfU1Pj1_0),.din(w_dff_A_l7ISEKSu8_0),.clk(gclk));
	jdff dff_A_OtdfU1Pj1_0(.dout(w_dff_A_mue8HkJW4_0),.din(w_dff_A_OtdfU1Pj1_0),.clk(gclk));
	jdff dff_A_mue8HkJW4_0(.dout(w_dff_A_yqGfCi8F5_0),.din(w_dff_A_mue8HkJW4_0),.clk(gclk));
	jdff dff_A_yqGfCi8F5_0(.dout(w_dff_A_uoUYJGq24_0),.din(w_dff_A_yqGfCi8F5_0),.clk(gclk));
	jdff dff_A_uoUYJGq24_0(.dout(w_dff_A_acO3YlaP4_0),.din(w_dff_A_uoUYJGq24_0),.clk(gclk));
	jdff dff_A_acO3YlaP4_0(.dout(w_dff_A_ctM2dYWb6_0),.din(w_dff_A_acO3YlaP4_0),.clk(gclk));
	jdff dff_A_ctM2dYWb6_0(.dout(w_dff_A_GRk5yzkq3_0),.din(w_dff_A_ctM2dYWb6_0),.clk(gclk));
	jdff dff_A_GRk5yzkq3_0(.dout(w_dff_A_pYljRpJX2_0),.din(w_dff_A_GRk5yzkq3_0),.clk(gclk));
	jdff dff_A_pYljRpJX2_0(.dout(w_dff_A_o3rCca0V4_0),.din(w_dff_A_pYljRpJX2_0),.clk(gclk));
	jdff dff_A_o3rCca0V4_0(.dout(w_dff_A_FSbSJtL34_0),.din(w_dff_A_o3rCca0V4_0),.clk(gclk));
	jdff dff_A_FSbSJtL34_0(.dout(w_dff_A_3xBXSfal7_0),.din(w_dff_A_FSbSJtL34_0),.clk(gclk));
	jdff dff_A_3xBXSfal7_0(.dout(w_dff_A_gUEw0R6k7_0),.din(w_dff_A_3xBXSfal7_0),.clk(gclk));
	jdff dff_A_gUEw0R6k7_0(.dout(w_dff_A_nFWSTKc02_0),.din(w_dff_A_gUEw0R6k7_0),.clk(gclk));
	jdff dff_A_nFWSTKc02_0(.dout(w_dff_A_MpCT5jKU2_0),.din(w_dff_A_nFWSTKc02_0),.clk(gclk));
	jdff dff_A_MpCT5jKU2_0(.dout(G993),.din(w_dff_A_MpCT5jKU2_0),.clk(gclk));
	jdff dff_A_iX0YGi3V0_1(.dout(w_dff_A_uPMFkgiK0_0),.din(w_dff_A_iX0YGi3V0_1),.clk(gclk));
	jdff dff_A_uPMFkgiK0_0(.dout(w_dff_A_Rwek7Y8j2_0),.din(w_dff_A_uPMFkgiK0_0),.clk(gclk));
	jdff dff_A_Rwek7Y8j2_0(.dout(w_dff_A_5ZD3t5XU0_0),.din(w_dff_A_Rwek7Y8j2_0),.clk(gclk));
	jdff dff_A_5ZD3t5XU0_0(.dout(w_dff_A_ZcMaCXiN7_0),.din(w_dff_A_5ZD3t5XU0_0),.clk(gclk));
	jdff dff_A_ZcMaCXiN7_0(.dout(w_dff_A_nack7WKD7_0),.din(w_dff_A_ZcMaCXiN7_0),.clk(gclk));
	jdff dff_A_nack7WKD7_0(.dout(w_dff_A_rF0C75SO9_0),.din(w_dff_A_nack7WKD7_0),.clk(gclk));
	jdff dff_A_rF0C75SO9_0(.dout(w_dff_A_CdkQSd1x3_0),.din(w_dff_A_rF0C75SO9_0),.clk(gclk));
	jdff dff_A_CdkQSd1x3_0(.dout(w_dff_A_4OuDYHoh8_0),.din(w_dff_A_CdkQSd1x3_0),.clk(gclk));
	jdff dff_A_4OuDYHoh8_0(.dout(w_dff_A_zSZ3q2jN6_0),.din(w_dff_A_4OuDYHoh8_0),.clk(gclk));
	jdff dff_A_zSZ3q2jN6_0(.dout(w_dff_A_nhVGhS5G2_0),.din(w_dff_A_zSZ3q2jN6_0),.clk(gclk));
	jdff dff_A_nhVGhS5G2_0(.dout(w_dff_A_jFQXGY4W0_0),.din(w_dff_A_nhVGhS5G2_0),.clk(gclk));
	jdff dff_A_jFQXGY4W0_0(.dout(w_dff_A_OxYy07Nz4_0),.din(w_dff_A_jFQXGY4W0_0),.clk(gclk));
	jdff dff_A_OxYy07Nz4_0(.dout(w_dff_A_TuZ54p393_0),.din(w_dff_A_OxYy07Nz4_0),.clk(gclk));
	jdff dff_A_TuZ54p393_0(.dout(w_dff_A_Q3b3frXR6_0),.din(w_dff_A_TuZ54p393_0),.clk(gclk));
	jdff dff_A_Q3b3frXR6_0(.dout(w_dff_A_73WZmY8t9_0),.din(w_dff_A_Q3b3frXR6_0),.clk(gclk));
	jdff dff_A_73WZmY8t9_0(.dout(w_dff_A_XTVnZnC67_0),.din(w_dff_A_73WZmY8t9_0),.clk(gclk));
	jdff dff_A_XTVnZnC67_0(.dout(w_dff_A_jmRj4X3v9_0),.din(w_dff_A_XTVnZnC67_0),.clk(gclk));
	jdff dff_A_jmRj4X3v9_0(.dout(w_dff_A_9OS8w7ag8_0),.din(w_dff_A_jmRj4X3v9_0),.clk(gclk));
	jdff dff_A_9OS8w7ag8_0(.dout(w_dff_A_vGK8cV1X4_0),.din(w_dff_A_9OS8w7ag8_0),.clk(gclk));
	jdff dff_A_vGK8cV1X4_0(.dout(w_dff_A_io1MLuGf8_0),.din(w_dff_A_vGK8cV1X4_0),.clk(gclk));
	jdff dff_A_io1MLuGf8_0(.dout(w_dff_A_ZT50cMaF1_0),.din(w_dff_A_io1MLuGf8_0),.clk(gclk));
	jdff dff_A_ZT50cMaF1_0(.dout(w_dff_A_KnGPUazE0_0),.din(w_dff_A_ZT50cMaF1_0),.clk(gclk));
	jdff dff_A_KnGPUazE0_0(.dout(w_dff_A_fsCTBilZ2_0),.din(w_dff_A_KnGPUazE0_0),.clk(gclk));
	jdff dff_A_fsCTBilZ2_0(.dout(w_dff_A_LRw983rV2_0),.din(w_dff_A_fsCTBilZ2_0),.clk(gclk));
	jdff dff_A_LRw983rV2_0(.dout(w_dff_A_JNJ830t24_0),.din(w_dff_A_LRw983rV2_0),.clk(gclk));
	jdff dff_A_JNJ830t24_0(.dout(G978),.din(w_dff_A_JNJ830t24_0),.clk(gclk));
	jdff dff_A_FzCJlgsD0_1(.dout(w_dff_A_dmqgJdYK4_0),.din(w_dff_A_FzCJlgsD0_1),.clk(gclk));
	jdff dff_A_dmqgJdYK4_0(.dout(w_dff_A_2QQJPzUD8_0),.din(w_dff_A_dmqgJdYK4_0),.clk(gclk));
	jdff dff_A_2QQJPzUD8_0(.dout(w_dff_A_uE8It0L95_0),.din(w_dff_A_2QQJPzUD8_0),.clk(gclk));
	jdff dff_A_uE8It0L95_0(.dout(w_dff_A_s7llUBAs4_0),.din(w_dff_A_uE8It0L95_0),.clk(gclk));
	jdff dff_A_s7llUBAs4_0(.dout(w_dff_A_AEfoKEYj8_0),.din(w_dff_A_s7llUBAs4_0),.clk(gclk));
	jdff dff_A_AEfoKEYj8_0(.dout(w_dff_A_Pr9QXGPp1_0),.din(w_dff_A_AEfoKEYj8_0),.clk(gclk));
	jdff dff_A_Pr9QXGPp1_0(.dout(w_dff_A_kRCdJWnq7_0),.din(w_dff_A_Pr9QXGPp1_0),.clk(gclk));
	jdff dff_A_kRCdJWnq7_0(.dout(w_dff_A_ajdiTEoj5_0),.din(w_dff_A_kRCdJWnq7_0),.clk(gclk));
	jdff dff_A_ajdiTEoj5_0(.dout(w_dff_A_GB3TSgUR4_0),.din(w_dff_A_ajdiTEoj5_0),.clk(gclk));
	jdff dff_A_GB3TSgUR4_0(.dout(w_dff_A_swdJ8koh8_0),.din(w_dff_A_GB3TSgUR4_0),.clk(gclk));
	jdff dff_A_swdJ8koh8_0(.dout(w_dff_A_ilnXyLGe7_0),.din(w_dff_A_swdJ8koh8_0),.clk(gclk));
	jdff dff_A_ilnXyLGe7_0(.dout(w_dff_A_gIZtQk7r6_0),.din(w_dff_A_ilnXyLGe7_0),.clk(gclk));
	jdff dff_A_gIZtQk7r6_0(.dout(w_dff_A_lWwMjQo36_0),.din(w_dff_A_gIZtQk7r6_0),.clk(gclk));
	jdff dff_A_lWwMjQo36_0(.dout(w_dff_A_O7eCQBbb2_0),.din(w_dff_A_lWwMjQo36_0),.clk(gclk));
	jdff dff_A_O7eCQBbb2_0(.dout(w_dff_A_xTEGNqlA5_0),.din(w_dff_A_O7eCQBbb2_0),.clk(gclk));
	jdff dff_A_xTEGNqlA5_0(.dout(w_dff_A_uUZh42M83_0),.din(w_dff_A_xTEGNqlA5_0),.clk(gclk));
	jdff dff_A_uUZh42M83_0(.dout(w_dff_A_AerjJxn55_0),.din(w_dff_A_uUZh42M83_0),.clk(gclk));
	jdff dff_A_AerjJxn55_0(.dout(w_dff_A_YktjNGhO8_0),.din(w_dff_A_AerjJxn55_0),.clk(gclk));
	jdff dff_A_YktjNGhO8_0(.dout(w_dff_A_68Z6taLk3_0),.din(w_dff_A_YktjNGhO8_0),.clk(gclk));
	jdff dff_A_68Z6taLk3_0(.dout(w_dff_A_A1Uvqxpg2_0),.din(w_dff_A_68Z6taLk3_0),.clk(gclk));
	jdff dff_A_A1Uvqxpg2_0(.dout(w_dff_A_fmycmVYt0_0),.din(w_dff_A_A1Uvqxpg2_0),.clk(gclk));
	jdff dff_A_fmycmVYt0_0(.dout(w_dff_A_rz93mtqB6_0),.din(w_dff_A_fmycmVYt0_0),.clk(gclk));
	jdff dff_A_rz93mtqB6_0(.dout(w_dff_A_U97nWb8Q7_0),.din(w_dff_A_rz93mtqB6_0),.clk(gclk));
	jdff dff_A_U97nWb8Q7_0(.dout(w_dff_A_DZWc4IE48_0),.din(w_dff_A_U97nWb8Q7_0),.clk(gclk));
	jdff dff_A_DZWc4IE48_0(.dout(w_dff_A_Gub68ra10_0),.din(w_dff_A_DZWc4IE48_0),.clk(gclk));
	jdff dff_A_Gub68ra10_0(.dout(G949),.din(w_dff_A_Gub68ra10_0),.clk(gclk));
	jdff dff_A_PtVtnSx29_1(.dout(w_dff_A_fkZ5MK9m3_0),.din(w_dff_A_PtVtnSx29_1),.clk(gclk));
	jdff dff_A_fkZ5MK9m3_0(.dout(w_dff_A_B0Cr4v9X6_0),.din(w_dff_A_fkZ5MK9m3_0),.clk(gclk));
	jdff dff_A_B0Cr4v9X6_0(.dout(w_dff_A_1N53pl6k6_0),.din(w_dff_A_B0Cr4v9X6_0),.clk(gclk));
	jdff dff_A_1N53pl6k6_0(.dout(w_dff_A_Gr0SZmbl3_0),.din(w_dff_A_1N53pl6k6_0),.clk(gclk));
	jdff dff_A_Gr0SZmbl3_0(.dout(w_dff_A_408Dljpk0_0),.din(w_dff_A_Gr0SZmbl3_0),.clk(gclk));
	jdff dff_A_408Dljpk0_0(.dout(w_dff_A_SPm3Y7r77_0),.din(w_dff_A_408Dljpk0_0),.clk(gclk));
	jdff dff_A_SPm3Y7r77_0(.dout(w_dff_A_1CJ1iw1z4_0),.din(w_dff_A_SPm3Y7r77_0),.clk(gclk));
	jdff dff_A_1CJ1iw1z4_0(.dout(w_dff_A_jFjpe5yW0_0),.din(w_dff_A_1CJ1iw1z4_0),.clk(gclk));
	jdff dff_A_jFjpe5yW0_0(.dout(w_dff_A_9S70EFcj0_0),.din(w_dff_A_jFjpe5yW0_0),.clk(gclk));
	jdff dff_A_9S70EFcj0_0(.dout(w_dff_A_1qU3BK194_0),.din(w_dff_A_9S70EFcj0_0),.clk(gclk));
	jdff dff_A_1qU3BK194_0(.dout(w_dff_A_uLbWhK2j7_0),.din(w_dff_A_1qU3BK194_0),.clk(gclk));
	jdff dff_A_uLbWhK2j7_0(.dout(w_dff_A_ZCHuBAbr1_0),.din(w_dff_A_uLbWhK2j7_0),.clk(gclk));
	jdff dff_A_ZCHuBAbr1_0(.dout(w_dff_A_JJOFqeDL5_0),.din(w_dff_A_ZCHuBAbr1_0),.clk(gclk));
	jdff dff_A_JJOFqeDL5_0(.dout(w_dff_A_fWbAKXRj8_0),.din(w_dff_A_JJOFqeDL5_0),.clk(gclk));
	jdff dff_A_fWbAKXRj8_0(.dout(w_dff_A_7JKVIISd5_0),.din(w_dff_A_fWbAKXRj8_0),.clk(gclk));
	jdff dff_A_7JKVIISd5_0(.dout(w_dff_A_QF20WGQF1_0),.din(w_dff_A_7JKVIISd5_0),.clk(gclk));
	jdff dff_A_QF20WGQF1_0(.dout(w_dff_A_jZt2ctxf9_0),.din(w_dff_A_QF20WGQF1_0),.clk(gclk));
	jdff dff_A_jZt2ctxf9_0(.dout(w_dff_A_BNRjKA9u5_0),.din(w_dff_A_jZt2ctxf9_0),.clk(gclk));
	jdff dff_A_BNRjKA9u5_0(.dout(w_dff_A_xUHN77XW6_0),.din(w_dff_A_BNRjKA9u5_0),.clk(gclk));
	jdff dff_A_xUHN77XW6_0(.dout(w_dff_A_NheApzMZ7_0),.din(w_dff_A_xUHN77XW6_0),.clk(gclk));
	jdff dff_A_NheApzMZ7_0(.dout(w_dff_A_5lhFs6f03_0),.din(w_dff_A_NheApzMZ7_0),.clk(gclk));
	jdff dff_A_5lhFs6f03_0(.dout(w_dff_A_A1jHp2lW7_0),.din(w_dff_A_5lhFs6f03_0),.clk(gclk));
	jdff dff_A_A1jHp2lW7_0(.dout(w_dff_A_UOzIG68G1_0),.din(w_dff_A_A1jHp2lW7_0),.clk(gclk));
	jdff dff_A_UOzIG68G1_0(.dout(w_dff_A_YBjhP92M7_0),.din(w_dff_A_UOzIG68G1_0),.clk(gclk));
	jdff dff_A_YBjhP92M7_0(.dout(w_dff_A_M83qPGpc7_0),.din(w_dff_A_YBjhP92M7_0),.clk(gclk));
	jdff dff_A_M83qPGpc7_0(.dout(G939),.din(w_dff_A_M83qPGpc7_0),.clk(gclk));
	jdff dff_A_bcmCouej6_1(.dout(w_dff_A_0jyR4lP04_0),.din(w_dff_A_bcmCouej6_1),.clk(gclk));
	jdff dff_A_0jyR4lP04_0(.dout(w_dff_A_gmKLIKev7_0),.din(w_dff_A_0jyR4lP04_0),.clk(gclk));
	jdff dff_A_gmKLIKev7_0(.dout(w_dff_A_YTLtTUxd2_0),.din(w_dff_A_gmKLIKev7_0),.clk(gclk));
	jdff dff_A_YTLtTUxd2_0(.dout(w_dff_A_Ap2Le9Ou7_0),.din(w_dff_A_YTLtTUxd2_0),.clk(gclk));
	jdff dff_A_Ap2Le9Ou7_0(.dout(w_dff_A_h6xfBR1K8_0),.din(w_dff_A_Ap2Le9Ou7_0),.clk(gclk));
	jdff dff_A_h6xfBR1K8_0(.dout(w_dff_A_Wb3ghfmV5_0),.din(w_dff_A_h6xfBR1K8_0),.clk(gclk));
	jdff dff_A_Wb3ghfmV5_0(.dout(w_dff_A_iQxqBBte5_0),.din(w_dff_A_Wb3ghfmV5_0),.clk(gclk));
	jdff dff_A_iQxqBBte5_0(.dout(w_dff_A_I7gTCGFI3_0),.din(w_dff_A_iQxqBBte5_0),.clk(gclk));
	jdff dff_A_I7gTCGFI3_0(.dout(w_dff_A_B294Nn5X4_0),.din(w_dff_A_I7gTCGFI3_0),.clk(gclk));
	jdff dff_A_B294Nn5X4_0(.dout(w_dff_A_ZZyr5BFy2_0),.din(w_dff_A_B294Nn5X4_0),.clk(gclk));
	jdff dff_A_ZZyr5BFy2_0(.dout(w_dff_A_DbAQnLHE3_0),.din(w_dff_A_ZZyr5BFy2_0),.clk(gclk));
	jdff dff_A_DbAQnLHE3_0(.dout(w_dff_A_1wRDI2Yz8_0),.din(w_dff_A_DbAQnLHE3_0),.clk(gclk));
	jdff dff_A_1wRDI2Yz8_0(.dout(w_dff_A_Y8fz1tEs0_0),.din(w_dff_A_1wRDI2Yz8_0),.clk(gclk));
	jdff dff_A_Y8fz1tEs0_0(.dout(w_dff_A_3rMu2ikH3_0),.din(w_dff_A_Y8fz1tEs0_0),.clk(gclk));
	jdff dff_A_3rMu2ikH3_0(.dout(w_dff_A_a1lF7Oo46_0),.din(w_dff_A_3rMu2ikH3_0),.clk(gclk));
	jdff dff_A_a1lF7Oo46_0(.dout(w_dff_A_hVQg70iO8_0),.din(w_dff_A_a1lF7Oo46_0),.clk(gclk));
	jdff dff_A_hVQg70iO8_0(.dout(w_dff_A_XMlaIjP11_0),.din(w_dff_A_hVQg70iO8_0),.clk(gclk));
	jdff dff_A_XMlaIjP11_0(.dout(w_dff_A_mU4Kjgeb7_0),.din(w_dff_A_XMlaIjP11_0),.clk(gclk));
	jdff dff_A_mU4Kjgeb7_0(.dout(w_dff_A_A92cHQJO4_0),.din(w_dff_A_mU4Kjgeb7_0),.clk(gclk));
	jdff dff_A_A92cHQJO4_0(.dout(w_dff_A_4PJwjazR5_0),.din(w_dff_A_A92cHQJO4_0),.clk(gclk));
	jdff dff_A_4PJwjazR5_0(.dout(w_dff_A_VcHY7LOQ3_0),.din(w_dff_A_4PJwjazR5_0),.clk(gclk));
	jdff dff_A_VcHY7LOQ3_0(.dout(w_dff_A_jYKzQ7hn3_0),.din(w_dff_A_VcHY7LOQ3_0),.clk(gclk));
	jdff dff_A_jYKzQ7hn3_0(.dout(w_dff_A_HA24eAHg9_0),.din(w_dff_A_jYKzQ7hn3_0),.clk(gclk));
	jdff dff_A_HA24eAHg9_0(.dout(w_dff_A_ndTmpEou3_0),.din(w_dff_A_HA24eAHg9_0),.clk(gclk));
	jdff dff_A_ndTmpEou3_0(.dout(w_dff_A_dFui7bHY3_0),.din(w_dff_A_ndTmpEou3_0),.clk(gclk));
	jdff dff_A_dFui7bHY3_0(.dout(G889),.din(w_dff_A_dFui7bHY3_0),.clk(gclk));
	jdff dff_A_iy5NfA8p1_1(.dout(w_dff_A_WnizSuDl5_0),.din(w_dff_A_iy5NfA8p1_1),.clk(gclk));
	jdff dff_A_WnizSuDl5_0(.dout(w_dff_A_jqAJpjmk0_0),.din(w_dff_A_WnizSuDl5_0),.clk(gclk));
	jdff dff_A_jqAJpjmk0_0(.dout(w_dff_A_5ShCLTLz2_0),.din(w_dff_A_jqAJpjmk0_0),.clk(gclk));
	jdff dff_A_5ShCLTLz2_0(.dout(w_dff_A_edl3g0y16_0),.din(w_dff_A_5ShCLTLz2_0),.clk(gclk));
	jdff dff_A_edl3g0y16_0(.dout(w_dff_A_F23wutM29_0),.din(w_dff_A_edl3g0y16_0),.clk(gclk));
	jdff dff_A_F23wutM29_0(.dout(w_dff_A_fCjuVgCk7_0),.din(w_dff_A_F23wutM29_0),.clk(gclk));
	jdff dff_A_fCjuVgCk7_0(.dout(w_dff_A_Wd3bmiyF4_0),.din(w_dff_A_fCjuVgCk7_0),.clk(gclk));
	jdff dff_A_Wd3bmiyF4_0(.dout(w_dff_A_NlFev7FY6_0),.din(w_dff_A_Wd3bmiyF4_0),.clk(gclk));
	jdff dff_A_NlFev7FY6_0(.dout(w_dff_A_r32K8gd08_0),.din(w_dff_A_NlFev7FY6_0),.clk(gclk));
	jdff dff_A_r32K8gd08_0(.dout(w_dff_A_2fj1LZui6_0),.din(w_dff_A_r32K8gd08_0),.clk(gclk));
	jdff dff_A_2fj1LZui6_0(.dout(w_dff_A_eMI39XM03_0),.din(w_dff_A_2fj1LZui6_0),.clk(gclk));
	jdff dff_A_eMI39XM03_0(.dout(w_dff_A_J7yENLvS0_0),.din(w_dff_A_eMI39XM03_0),.clk(gclk));
	jdff dff_A_J7yENLvS0_0(.dout(w_dff_A_njOTFXhz2_0),.din(w_dff_A_J7yENLvS0_0),.clk(gclk));
	jdff dff_A_njOTFXhz2_0(.dout(w_dff_A_JmBlk7qa4_0),.din(w_dff_A_njOTFXhz2_0),.clk(gclk));
	jdff dff_A_JmBlk7qa4_0(.dout(w_dff_A_xbHFW4oG3_0),.din(w_dff_A_JmBlk7qa4_0),.clk(gclk));
	jdff dff_A_xbHFW4oG3_0(.dout(w_dff_A_cXk9f2aw7_0),.din(w_dff_A_xbHFW4oG3_0),.clk(gclk));
	jdff dff_A_cXk9f2aw7_0(.dout(w_dff_A_XF12hza79_0),.din(w_dff_A_cXk9f2aw7_0),.clk(gclk));
	jdff dff_A_XF12hza79_0(.dout(w_dff_A_Pc8IWniA8_0),.din(w_dff_A_XF12hza79_0),.clk(gclk));
	jdff dff_A_Pc8IWniA8_0(.dout(w_dff_A_HvLlkRkW3_0),.din(w_dff_A_Pc8IWniA8_0),.clk(gclk));
	jdff dff_A_HvLlkRkW3_0(.dout(w_dff_A_kTiCZk2C8_0),.din(w_dff_A_HvLlkRkW3_0),.clk(gclk));
	jdff dff_A_kTiCZk2C8_0(.dout(w_dff_A_WOCNomxj0_0),.din(w_dff_A_kTiCZk2C8_0),.clk(gclk));
	jdff dff_A_WOCNomxj0_0(.dout(w_dff_A_xQE2EbN35_0),.din(w_dff_A_WOCNomxj0_0),.clk(gclk));
	jdff dff_A_xQE2EbN35_0(.dout(w_dff_A_HB62ZxmB8_0),.din(w_dff_A_xQE2EbN35_0),.clk(gclk));
	jdff dff_A_HB62ZxmB8_0(.dout(w_dff_A_QnMQBUgv3_0),.din(w_dff_A_HB62ZxmB8_0),.clk(gclk));
	jdff dff_A_QnMQBUgv3_0(.dout(G593),.din(w_dff_A_QnMQBUgv3_0),.clk(gclk));
	jdff dff_A_DH3gqMbd6_2(.dout(w_dff_A_CmMV3JTc6_0),.din(w_dff_A_DH3gqMbd6_2),.clk(gclk));
	jdff dff_A_CmMV3JTc6_0(.dout(w_dff_A_4sAg2tf42_0),.din(w_dff_A_CmMV3JTc6_0),.clk(gclk));
	jdff dff_A_4sAg2tf42_0(.dout(w_dff_A_6TuJaMJU3_0),.din(w_dff_A_4sAg2tf42_0),.clk(gclk));
	jdff dff_A_6TuJaMJU3_0(.dout(w_dff_A_SJq7rbG52_0),.din(w_dff_A_6TuJaMJU3_0),.clk(gclk));
	jdff dff_A_SJq7rbG52_0(.dout(w_dff_A_zR1ClXM12_0),.din(w_dff_A_SJq7rbG52_0),.clk(gclk));
	jdff dff_A_zR1ClXM12_0(.dout(w_dff_A_7QSNtk6c3_0),.din(w_dff_A_zR1ClXM12_0),.clk(gclk));
	jdff dff_A_7QSNtk6c3_0(.dout(w_dff_A_0RIaDIDr2_0),.din(w_dff_A_7QSNtk6c3_0),.clk(gclk));
	jdff dff_A_0RIaDIDr2_0(.dout(w_dff_A_3ye0t4pd9_0),.din(w_dff_A_0RIaDIDr2_0),.clk(gclk));
	jdff dff_A_3ye0t4pd9_0(.dout(w_dff_A_pjsRGaGO3_0),.din(w_dff_A_3ye0t4pd9_0),.clk(gclk));
	jdff dff_A_pjsRGaGO3_0(.dout(w_dff_A_0GUbYCaN5_0),.din(w_dff_A_pjsRGaGO3_0),.clk(gclk));
	jdff dff_A_0GUbYCaN5_0(.dout(w_dff_A_g5no8Ieu0_0),.din(w_dff_A_0GUbYCaN5_0),.clk(gclk));
	jdff dff_A_g5no8Ieu0_0(.dout(w_dff_A_ovphpXRL6_0),.din(w_dff_A_g5no8Ieu0_0),.clk(gclk));
	jdff dff_A_ovphpXRL6_0(.dout(w_dff_A_w0Ofdea05_0),.din(w_dff_A_ovphpXRL6_0),.clk(gclk));
	jdff dff_A_w0Ofdea05_0(.dout(w_dff_A_7O0dIBuK8_0),.din(w_dff_A_w0Ofdea05_0),.clk(gclk));
	jdff dff_A_7O0dIBuK8_0(.dout(w_dff_A_hoZIqJxi2_0),.din(w_dff_A_7O0dIBuK8_0),.clk(gclk));
	jdff dff_A_hoZIqJxi2_0(.dout(w_dff_A_BWLc6lkr4_0),.din(w_dff_A_hoZIqJxi2_0),.clk(gclk));
	jdff dff_A_BWLc6lkr4_0(.dout(w_dff_A_n32w4r7Q7_0),.din(w_dff_A_BWLc6lkr4_0),.clk(gclk));
	jdff dff_A_n32w4r7Q7_0(.dout(w_dff_A_QqrZRL7u9_0),.din(w_dff_A_n32w4r7Q7_0),.clk(gclk));
	jdff dff_A_QqrZRL7u9_0(.dout(w_dff_A_VovFy6QC9_0),.din(w_dff_A_QqrZRL7u9_0),.clk(gclk));
	jdff dff_A_VovFy6QC9_0(.dout(w_dff_A_KDKlOLjc6_0),.din(w_dff_A_VovFy6QC9_0),.clk(gclk));
	jdff dff_A_KDKlOLjc6_0(.dout(w_dff_A_eCjy2DTL6_0),.din(w_dff_A_KDKlOLjc6_0),.clk(gclk));
	jdff dff_A_eCjy2DTL6_0(.dout(G636),.din(w_dff_A_eCjy2DTL6_0),.clk(gclk));
	jdff dff_A_4mIO0Omj6_2(.dout(w_dff_A_42libba56_0),.din(w_dff_A_4mIO0Omj6_2),.clk(gclk));
	jdff dff_A_42libba56_0(.dout(w_dff_A_ICpZIEjr2_0),.din(w_dff_A_42libba56_0),.clk(gclk));
	jdff dff_A_ICpZIEjr2_0(.dout(w_dff_A_myNgd3T04_0),.din(w_dff_A_ICpZIEjr2_0),.clk(gclk));
	jdff dff_A_myNgd3T04_0(.dout(w_dff_A_LECBlswP2_0),.din(w_dff_A_myNgd3T04_0),.clk(gclk));
	jdff dff_A_LECBlswP2_0(.dout(w_dff_A_i4mh0IRK1_0),.din(w_dff_A_LECBlswP2_0),.clk(gclk));
	jdff dff_A_i4mh0IRK1_0(.dout(w_dff_A_8dB4UqgM0_0),.din(w_dff_A_i4mh0IRK1_0),.clk(gclk));
	jdff dff_A_8dB4UqgM0_0(.dout(w_dff_A_SaT244wW4_0),.din(w_dff_A_8dB4UqgM0_0),.clk(gclk));
	jdff dff_A_SaT244wW4_0(.dout(w_dff_A_d5BNXPMn3_0),.din(w_dff_A_SaT244wW4_0),.clk(gclk));
	jdff dff_A_d5BNXPMn3_0(.dout(w_dff_A_7ifcpMUb6_0),.din(w_dff_A_d5BNXPMn3_0),.clk(gclk));
	jdff dff_A_7ifcpMUb6_0(.dout(w_dff_A_7yauADEk4_0),.din(w_dff_A_7ifcpMUb6_0),.clk(gclk));
	jdff dff_A_7yauADEk4_0(.dout(w_dff_A_hFthHK0W8_0),.din(w_dff_A_7yauADEk4_0),.clk(gclk));
	jdff dff_A_hFthHK0W8_0(.dout(w_dff_A_ZqPdSjTr7_0),.din(w_dff_A_hFthHK0W8_0),.clk(gclk));
	jdff dff_A_ZqPdSjTr7_0(.dout(w_dff_A_vnJaF1wA2_0),.din(w_dff_A_ZqPdSjTr7_0),.clk(gclk));
	jdff dff_A_vnJaF1wA2_0(.dout(w_dff_A_OTwb2gWc9_0),.din(w_dff_A_vnJaF1wA2_0),.clk(gclk));
	jdff dff_A_OTwb2gWc9_0(.dout(w_dff_A_ByzumVJf7_0),.din(w_dff_A_OTwb2gWc9_0),.clk(gclk));
	jdff dff_A_ByzumVJf7_0(.dout(w_dff_A_3sFOxuGv5_0),.din(w_dff_A_ByzumVJf7_0),.clk(gclk));
	jdff dff_A_3sFOxuGv5_0(.dout(w_dff_A_eDC7b2zl8_0),.din(w_dff_A_3sFOxuGv5_0),.clk(gclk));
	jdff dff_A_eDC7b2zl8_0(.dout(w_dff_A_7mLwgt455_0),.din(w_dff_A_eDC7b2zl8_0),.clk(gclk));
	jdff dff_A_7mLwgt455_0(.dout(w_dff_A_x2eiRihv3_0),.din(w_dff_A_7mLwgt455_0),.clk(gclk));
	jdff dff_A_x2eiRihv3_0(.dout(w_dff_A_mYNzs6kq8_0),.din(w_dff_A_x2eiRihv3_0),.clk(gclk));
	jdff dff_A_mYNzs6kq8_0(.dout(w_dff_A_vw4iXDjF4_0),.din(w_dff_A_mYNzs6kq8_0),.clk(gclk));
	jdff dff_A_vw4iXDjF4_0(.dout(G704),.din(w_dff_A_vw4iXDjF4_0),.clk(gclk));
	jdff dff_A_2Em61F4H5_2(.dout(w_dff_A_xiUguW3E1_0),.din(w_dff_A_2Em61F4H5_2),.clk(gclk));
	jdff dff_A_xiUguW3E1_0(.dout(w_dff_A_40YbK28V7_0),.din(w_dff_A_xiUguW3E1_0),.clk(gclk));
	jdff dff_A_40YbK28V7_0(.dout(w_dff_A_x7HYhBMb5_0),.din(w_dff_A_40YbK28V7_0),.clk(gclk));
	jdff dff_A_x7HYhBMb5_0(.dout(w_dff_A_pgxDGr2p1_0),.din(w_dff_A_x7HYhBMb5_0),.clk(gclk));
	jdff dff_A_pgxDGr2p1_0(.dout(w_dff_A_6sFEABCs6_0),.din(w_dff_A_pgxDGr2p1_0),.clk(gclk));
	jdff dff_A_6sFEABCs6_0(.dout(w_dff_A_O85zz5Yw9_0),.din(w_dff_A_6sFEABCs6_0),.clk(gclk));
	jdff dff_A_O85zz5Yw9_0(.dout(w_dff_A_aNcka0Tf5_0),.din(w_dff_A_O85zz5Yw9_0),.clk(gclk));
	jdff dff_A_aNcka0Tf5_0(.dout(w_dff_A_FyvA1L460_0),.din(w_dff_A_aNcka0Tf5_0),.clk(gclk));
	jdff dff_A_FyvA1L460_0(.dout(w_dff_A_btOH0xby6_0),.din(w_dff_A_FyvA1L460_0),.clk(gclk));
	jdff dff_A_btOH0xby6_0(.dout(w_dff_A_tgUyvSwV0_0),.din(w_dff_A_btOH0xby6_0),.clk(gclk));
	jdff dff_A_tgUyvSwV0_0(.dout(w_dff_A_V6IfQMwu5_0),.din(w_dff_A_tgUyvSwV0_0),.clk(gclk));
	jdff dff_A_V6IfQMwu5_0(.dout(w_dff_A_DrrzWTJH3_0),.din(w_dff_A_V6IfQMwu5_0),.clk(gclk));
	jdff dff_A_DrrzWTJH3_0(.dout(w_dff_A_1Ds676rs7_0),.din(w_dff_A_DrrzWTJH3_0),.clk(gclk));
	jdff dff_A_1Ds676rs7_0(.dout(w_dff_A_8NHAdBE15_0),.din(w_dff_A_1Ds676rs7_0),.clk(gclk));
	jdff dff_A_8NHAdBE15_0(.dout(w_dff_A_9ngVJhHv1_0),.din(w_dff_A_8NHAdBE15_0),.clk(gclk));
	jdff dff_A_9ngVJhHv1_0(.dout(w_dff_A_ggvqsBZ73_0),.din(w_dff_A_9ngVJhHv1_0),.clk(gclk));
	jdff dff_A_ggvqsBZ73_0(.dout(w_dff_A_f1588PC83_0),.din(w_dff_A_ggvqsBZ73_0),.clk(gclk));
	jdff dff_A_f1588PC83_0(.dout(w_dff_A_sHuAMXua5_0),.din(w_dff_A_f1588PC83_0),.clk(gclk));
	jdff dff_A_sHuAMXua5_0(.dout(w_dff_A_iG8A7Kc61_0),.din(w_dff_A_sHuAMXua5_0),.clk(gclk));
	jdff dff_A_iG8A7Kc61_0(.dout(w_dff_A_sYQDF5Ft9_0),.din(w_dff_A_iG8A7Kc61_0),.clk(gclk));
	jdff dff_A_sYQDF5Ft9_0(.dout(w_dff_A_4jhY0ozW6_0),.din(w_dff_A_sYQDF5Ft9_0),.clk(gclk));
	jdff dff_A_4jhY0ozW6_0(.dout(G717),.din(w_dff_A_4jhY0ozW6_0),.clk(gclk));
	jdff dff_A_A5LKfscm0_2(.dout(w_dff_A_8UVu3P1o4_0),.din(w_dff_A_A5LKfscm0_2),.clk(gclk));
	jdff dff_A_8UVu3P1o4_0(.dout(w_dff_A_IgtMrHSH0_0),.din(w_dff_A_8UVu3P1o4_0),.clk(gclk));
	jdff dff_A_IgtMrHSH0_0(.dout(w_dff_A_eQ7ytHvT5_0),.din(w_dff_A_IgtMrHSH0_0),.clk(gclk));
	jdff dff_A_eQ7ytHvT5_0(.dout(w_dff_A_BvcAjru20_0),.din(w_dff_A_eQ7ytHvT5_0),.clk(gclk));
	jdff dff_A_BvcAjru20_0(.dout(w_dff_A_Tqws9Go98_0),.din(w_dff_A_BvcAjru20_0),.clk(gclk));
	jdff dff_A_Tqws9Go98_0(.dout(w_dff_A_dO9ENwZc2_0),.din(w_dff_A_Tqws9Go98_0),.clk(gclk));
	jdff dff_A_dO9ENwZc2_0(.dout(w_dff_A_BsssJlFj5_0),.din(w_dff_A_dO9ENwZc2_0),.clk(gclk));
	jdff dff_A_BsssJlFj5_0(.dout(w_dff_A_WvTHqim74_0),.din(w_dff_A_BsssJlFj5_0),.clk(gclk));
	jdff dff_A_WvTHqim74_0(.dout(w_dff_A_nvkX9kGY8_0),.din(w_dff_A_WvTHqim74_0),.clk(gclk));
	jdff dff_A_nvkX9kGY8_0(.dout(w_dff_A_Obspi6Qb8_0),.din(w_dff_A_nvkX9kGY8_0),.clk(gclk));
	jdff dff_A_Obspi6Qb8_0(.dout(w_dff_A_Nar49g3h6_0),.din(w_dff_A_Obspi6Qb8_0),.clk(gclk));
	jdff dff_A_Nar49g3h6_0(.dout(w_dff_A_zvRhIdJR3_0),.din(w_dff_A_Nar49g3h6_0),.clk(gclk));
	jdff dff_A_zvRhIdJR3_0(.dout(w_dff_A_SFGJmORD5_0),.din(w_dff_A_zvRhIdJR3_0),.clk(gclk));
	jdff dff_A_SFGJmORD5_0(.dout(w_dff_A_cJtRRpLy3_0),.din(w_dff_A_SFGJmORD5_0),.clk(gclk));
	jdff dff_A_cJtRRpLy3_0(.dout(w_dff_A_DGuOGsEF6_0),.din(w_dff_A_cJtRRpLy3_0),.clk(gclk));
	jdff dff_A_DGuOGsEF6_0(.dout(w_dff_A_zT3UutYA1_0),.din(w_dff_A_DGuOGsEF6_0),.clk(gclk));
	jdff dff_A_zT3UutYA1_0(.dout(w_dff_A_YIwsOfxn3_0),.din(w_dff_A_zT3UutYA1_0),.clk(gclk));
	jdff dff_A_YIwsOfxn3_0(.dout(w_dff_A_0ZjIJTIx7_0),.din(w_dff_A_YIwsOfxn3_0),.clk(gclk));
	jdff dff_A_0ZjIJTIx7_0(.dout(w_dff_A_wGrbOC296_0),.din(w_dff_A_0ZjIJTIx7_0),.clk(gclk));
	jdff dff_A_wGrbOC296_0(.dout(w_dff_A_xp30hxAN5_0),.din(w_dff_A_wGrbOC296_0),.clk(gclk));
	jdff dff_A_xp30hxAN5_0(.dout(w_dff_A_lIQFrxW29_0),.din(w_dff_A_xp30hxAN5_0),.clk(gclk));
	jdff dff_A_lIQFrxW29_0(.dout(w_dff_A_NbbBuFK88_0),.din(w_dff_A_lIQFrxW29_0),.clk(gclk));
	jdff dff_A_NbbBuFK88_0(.dout(G820),.din(w_dff_A_NbbBuFK88_0),.clk(gclk));
	jdff dff_A_Dmxui67i6_2(.dout(w_dff_A_x9gktYI57_0),.din(w_dff_A_Dmxui67i6_2),.clk(gclk));
	jdff dff_A_x9gktYI57_0(.dout(w_dff_A_mVo6lrbu5_0),.din(w_dff_A_x9gktYI57_0),.clk(gclk));
	jdff dff_A_mVo6lrbu5_0(.dout(w_dff_A_JkoDpI2e9_0),.din(w_dff_A_mVo6lrbu5_0),.clk(gclk));
	jdff dff_A_JkoDpI2e9_0(.dout(w_dff_A_mxCGr4qK7_0),.din(w_dff_A_JkoDpI2e9_0),.clk(gclk));
	jdff dff_A_mxCGr4qK7_0(.dout(w_dff_A_Z5KuMd7A3_0),.din(w_dff_A_mxCGr4qK7_0),.clk(gclk));
	jdff dff_A_Z5KuMd7A3_0(.dout(w_dff_A_jqUCwjqE2_0),.din(w_dff_A_Z5KuMd7A3_0),.clk(gclk));
	jdff dff_A_jqUCwjqE2_0(.dout(w_dff_A_KdDENeJl7_0),.din(w_dff_A_jqUCwjqE2_0),.clk(gclk));
	jdff dff_A_KdDENeJl7_0(.dout(w_dff_A_GrJflWi90_0),.din(w_dff_A_KdDENeJl7_0),.clk(gclk));
	jdff dff_A_GrJflWi90_0(.dout(w_dff_A_w5EN2PPQ6_0),.din(w_dff_A_GrJflWi90_0),.clk(gclk));
	jdff dff_A_w5EN2PPQ6_0(.dout(w_dff_A_fzftObhP6_0),.din(w_dff_A_w5EN2PPQ6_0),.clk(gclk));
	jdff dff_A_fzftObhP6_0(.dout(w_dff_A_2dgtgsxt5_0),.din(w_dff_A_fzftObhP6_0),.clk(gclk));
	jdff dff_A_2dgtgsxt5_0(.dout(w_dff_A_8hesfdpX0_0),.din(w_dff_A_2dgtgsxt5_0),.clk(gclk));
	jdff dff_A_8hesfdpX0_0(.dout(w_dff_A_FCsUu0T63_0),.din(w_dff_A_8hesfdpX0_0),.clk(gclk));
	jdff dff_A_FCsUu0T63_0(.dout(w_dff_A_BbL73qQO2_0),.din(w_dff_A_FCsUu0T63_0),.clk(gclk));
	jdff dff_A_BbL73qQO2_0(.dout(w_dff_A_6xhh7bEr9_0),.din(w_dff_A_BbL73qQO2_0),.clk(gclk));
	jdff dff_A_6xhh7bEr9_0(.dout(w_dff_A_o5NfWBeA1_0),.din(w_dff_A_6xhh7bEr9_0),.clk(gclk));
	jdff dff_A_o5NfWBeA1_0(.dout(w_dff_A_FZ1sBM308_0),.din(w_dff_A_o5NfWBeA1_0),.clk(gclk));
	jdff dff_A_FZ1sBM308_0(.dout(w_dff_A_rcd1sCUV5_0),.din(w_dff_A_FZ1sBM308_0),.clk(gclk));
	jdff dff_A_rcd1sCUV5_0(.dout(w_dff_A_rDNfw0bc1_0),.din(w_dff_A_rcd1sCUV5_0),.clk(gclk));
	jdff dff_A_rDNfw0bc1_0(.dout(w_dff_A_fKR6z7ZD4_0),.din(w_dff_A_rDNfw0bc1_0),.clk(gclk));
	jdff dff_A_fKR6z7ZD4_0(.dout(G639),.din(w_dff_A_fKR6z7ZD4_0),.clk(gclk));
	jdff dff_A_HfINcbMs5_2(.dout(w_dff_A_NjjlIWWp7_0),.din(w_dff_A_HfINcbMs5_2),.clk(gclk));
	jdff dff_A_NjjlIWWp7_0(.dout(w_dff_A_wLhg0KgC0_0),.din(w_dff_A_NjjlIWWp7_0),.clk(gclk));
	jdff dff_A_wLhg0KgC0_0(.dout(w_dff_A_M5ihDUVK3_0),.din(w_dff_A_wLhg0KgC0_0),.clk(gclk));
	jdff dff_A_M5ihDUVK3_0(.dout(w_dff_A_uyJTWQvZ5_0),.din(w_dff_A_M5ihDUVK3_0),.clk(gclk));
	jdff dff_A_uyJTWQvZ5_0(.dout(w_dff_A_Q6myFDG04_0),.din(w_dff_A_uyJTWQvZ5_0),.clk(gclk));
	jdff dff_A_Q6myFDG04_0(.dout(w_dff_A_J1IczByK7_0),.din(w_dff_A_Q6myFDG04_0),.clk(gclk));
	jdff dff_A_J1IczByK7_0(.dout(w_dff_A_JDQLBS9Q9_0),.din(w_dff_A_J1IczByK7_0),.clk(gclk));
	jdff dff_A_JDQLBS9Q9_0(.dout(w_dff_A_IFH4fHVJ4_0),.din(w_dff_A_JDQLBS9Q9_0),.clk(gclk));
	jdff dff_A_IFH4fHVJ4_0(.dout(w_dff_A_XdVlqxEw6_0),.din(w_dff_A_IFH4fHVJ4_0),.clk(gclk));
	jdff dff_A_XdVlqxEw6_0(.dout(w_dff_A_yPvTAhhl9_0),.din(w_dff_A_XdVlqxEw6_0),.clk(gclk));
	jdff dff_A_yPvTAhhl9_0(.dout(w_dff_A_yFrkmDoC2_0),.din(w_dff_A_yPvTAhhl9_0),.clk(gclk));
	jdff dff_A_yFrkmDoC2_0(.dout(w_dff_A_Gpofob8w1_0),.din(w_dff_A_yFrkmDoC2_0),.clk(gclk));
	jdff dff_A_Gpofob8w1_0(.dout(w_dff_A_8IqI5o9d3_0),.din(w_dff_A_Gpofob8w1_0),.clk(gclk));
	jdff dff_A_8IqI5o9d3_0(.dout(w_dff_A_JY65UEty4_0),.din(w_dff_A_8IqI5o9d3_0),.clk(gclk));
	jdff dff_A_JY65UEty4_0(.dout(w_dff_A_mWIv4CyH7_0),.din(w_dff_A_JY65UEty4_0),.clk(gclk));
	jdff dff_A_mWIv4CyH7_0(.dout(w_dff_A_JL5VW8MT2_0),.din(w_dff_A_mWIv4CyH7_0),.clk(gclk));
	jdff dff_A_JL5VW8MT2_0(.dout(w_dff_A_MajAAWAF6_0),.din(w_dff_A_JL5VW8MT2_0),.clk(gclk));
	jdff dff_A_MajAAWAF6_0(.dout(w_dff_A_zvTHwCxX2_0),.din(w_dff_A_MajAAWAF6_0),.clk(gclk));
	jdff dff_A_zvTHwCxX2_0(.dout(w_dff_A_bf9cG4Uh4_0),.din(w_dff_A_zvTHwCxX2_0),.clk(gclk));
	jdff dff_A_bf9cG4Uh4_0(.dout(w_dff_A_XBBAZAtX5_0),.din(w_dff_A_bf9cG4Uh4_0),.clk(gclk));
	jdff dff_A_XBBAZAtX5_0(.dout(G673),.din(w_dff_A_XBBAZAtX5_0),.clk(gclk));
	jdff dff_A_tqTmAX2J9_2(.dout(w_dff_A_FbKda17C0_0),.din(w_dff_A_tqTmAX2J9_2),.clk(gclk));
	jdff dff_A_FbKda17C0_0(.dout(w_dff_A_vy1dXzfE3_0),.din(w_dff_A_FbKda17C0_0),.clk(gclk));
	jdff dff_A_vy1dXzfE3_0(.dout(w_dff_A_GwgnK8Ip5_0),.din(w_dff_A_vy1dXzfE3_0),.clk(gclk));
	jdff dff_A_GwgnK8Ip5_0(.dout(w_dff_A_KBcoGBz02_0),.din(w_dff_A_GwgnK8Ip5_0),.clk(gclk));
	jdff dff_A_KBcoGBz02_0(.dout(w_dff_A_4tPiuj820_0),.din(w_dff_A_KBcoGBz02_0),.clk(gclk));
	jdff dff_A_4tPiuj820_0(.dout(w_dff_A_c38XK2fk1_0),.din(w_dff_A_4tPiuj820_0),.clk(gclk));
	jdff dff_A_c38XK2fk1_0(.dout(w_dff_A_nGzWbQt52_0),.din(w_dff_A_c38XK2fk1_0),.clk(gclk));
	jdff dff_A_nGzWbQt52_0(.dout(w_dff_A_oJAor8DH0_0),.din(w_dff_A_nGzWbQt52_0),.clk(gclk));
	jdff dff_A_oJAor8DH0_0(.dout(w_dff_A_cmJn8vqh7_0),.din(w_dff_A_oJAor8DH0_0),.clk(gclk));
	jdff dff_A_cmJn8vqh7_0(.dout(w_dff_A_dOlrK4WA8_0),.din(w_dff_A_cmJn8vqh7_0),.clk(gclk));
	jdff dff_A_dOlrK4WA8_0(.dout(w_dff_A_E9yatNKt3_0),.din(w_dff_A_dOlrK4WA8_0),.clk(gclk));
	jdff dff_A_E9yatNKt3_0(.dout(w_dff_A_3gHNAW3k5_0),.din(w_dff_A_E9yatNKt3_0),.clk(gclk));
	jdff dff_A_3gHNAW3k5_0(.dout(w_dff_A_dTjKujKg0_0),.din(w_dff_A_3gHNAW3k5_0),.clk(gclk));
	jdff dff_A_dTjKujKg0_0(.dout(w_dff_A_ZnhYaYrQ4_0),.din(w_dff_A_dTjKujKg0_0),.clk(gclk));
	jdff dff_A_ZnhYaYrQ4_0(.dout(w_dff_A_vAwl76YB2_0),.din(w_dff_A_ZnhYaYrQ4_0),.clk(gclk));
	jdff dff_A_vAwl76YB2_0(.dout(w_dff_A_V9f7g9746_0),.din(w_dff_A_vAwl76YB2_0),.clk(gclk));
	jdff dff_A_V9f7g9746_0(.dout(w_dff_A_XlSktFXb4_0),.din(w_dff_A_V9f7g9746_0),.clk(gclk));
	jdff dff_A_XlSktFXb4_0(.dout(w_dff_A_qIno74EG6_0),.din(w_dff_A_XlSktFXb4_0),.clk(gclk));
	jdff dff_A_qIno74EG6_0(.dout(w_dff_A_sPYnRjJ17_0),.din(w_dff_A_qIno74EG6_0),.clk(gclk));
	jdff dff_A_sPYnRjJ17_0(.dout(w_dff_A_1mtzjYA46_0),.din(w_dff_A_sPYnRjJ17_0),.clk(gclk));
	jdff dff_A_1mtzjYA46_0(.dout(G707),.din(w_dff_A_1mtzjYA46_0),.clk(gclk));
	jdff dff_A_q4HuDZnG7_2(.dout(w_dff_A_TWZc9Xtm3_0),.din(w_dff_A_q4HuDZnG7_2),.clk(gclk));
	jdff dff_A_TWZc9Xtm3_0(.dout(w_dff_A_Rx6lPAWf1_0),.din(w_dff_A_TWZc9Xtm3_0),.clk(gclk));
	jdff dff_A_Rx6lPAWf1_0(.dout(w_dff_A_VIBZPs6z8_0),.din(w_dff_A_Rx6lPAWf1_0),.clk(gclk));
	jdff dff_A_VIBZPs6z8_0(.dout(w_dff_A_MKzonvyp8_0),.din(w_dff_A_VIBZPs6z8_0),.clk(gclk));
	jdff dff_A_MKzonvyp8_0(.dout(w_dff_A_5MHi83Gz0_0),.din(w_dff_A_MKzonvyp8_0),.clk(gclk));
	jdff dff_A_5MHi83Gz0_0(.dout(w_dff_A_53XiVxZg0_0),.din(w_dff_A_5MHi83Gz0_0),.clk(gclk));
	jdff dff_A_53XiVxZg0_0(.dout(w_dff_A_Kmxau93S9_0),.din(w_dff_A_53XiVxZg0_0),.clk(gclk));
	jdff dff_A_Kmxau93S9_0(.dout(w_dff_A_nGzfsclY7_0),.din(w_dff_A_Kmxau93S9_0),.clk(gclk));
	jdff dff_A_nGzfsclY7_0(.dout(w_dff_A_T1cJwZ1b2_0),.din(w_dff_A_nGzfsclY7_0),.clk(gclk));
	jdff dff_A_T1cJwZ1b2_0(.dout(w_dff_A_iJIqBvhn6_0),.din(w_dff_A_T1cJwZ1b2_0),.clk(gclk));
	jdff dff_A_iJIqBvhn6_0(.dout(w_dff_A_HgjWojgE0_0),.din(w_dff_A_iJIqBvhn6_0),.clk(gclk));
	jdff dff_A_HgjWojgE0_0(.dout(w_dff_A_XwsWGQLh1_0),.din(w_dff_A_HgjWojgE0_0),.clk(gclk));
	jdff dff_A_XwsWGQLh1_0(.dout(w_dff_A_avTfQtX47_0),.din(w_dff_A_XwsWGQLh1_0),.clk(gclk));
	jdff dff_A_avTfQtX47_0(.dout(w_dff_A_CdzOsXks1_0),.din(w_dff_A_avTfQtX47_0),.clk(gclk));
	jdff dff_A_CdzOsXks1_0(.dout(w_dff_A_0pycos278_0),.din(w_dff_A_CdzOsXks1_0),.clk(gclk));
	jdff dff_A_0pycos278_0(.dout(w_dff_A_yWTR9anx7_0),.din(w_dff_A_0pycos278_0),.clk(gclk));
	jdff dff_A_yWTR9anx7_0(.dout(w_dff_A_REVqGbwf5_0),.din(w_dff_A_yWTR9anx7_0),.clk(gclk));
	jdff dff_A_REVqGbwf5_0(.dout(w_dff_A_tmagXIk38_0),.din(w_dff_A_REVqGbwf5_0),.clk(gclk));
	jdff dff_A_tmagXIk38_0(.dout(w_dff_A_LmZjFiPI6_0),.din(w_dff_A_tmagXIk38_0),.clk(gclk));
	jdff dff_A_LmZjFiPI6_0(.dout(w_dff_A_U8gfVIhp5_0),.din(w_dff_A_LmZjFiPI6_0),.clk(gclk));
	jdff dff_A_U8gfVIhp5_0(.dout(G715),.din(w_dff_A_U8gfVIhp5_0),.clk(gclk));
	jdff dff_A_heVA6OvF9_2(.dout(w_dff_A_t8mItqJ92_0),.din(w_dff_A_heVA6OvF9_2),.clk(gclk));
	jdff dff_A_t8mItqJ92_0(.dout(w_dff_A_vosmfmve7_0),.din(w_dff_A_t8mItqJ92_0),.clk(gclk));
	jdff dff_A_vosmfmve7_0(.dout(w_dff_A_mdYMnQ570_0),.din(w_dff_A_vosmfmve7_0),.clk(gclk));
	jdff dff_A_mdYMnQ570_0(.dout(w_dff_A_F6s3PHqc5_0),.din(w_dff_A_mdYMnQ570_0),.clk(gclk));
	jdff dff_A_F6s3PHqc5_0(.dout(w_dff_A_xceauyHw8_0),.din(w_dff_A_F6s3PHqc5_0),.clk(gclk));
	jdff dff_A_xceauyHw8_0(.dout(w_dff_A_3VmWHgRi8_0),.din(w_dff_A_xceauyHw8_0),.clk(gclk));
	jdff dff_A_3VmWHgRi8_0(.dout(w_dff_A_N5nTT7Wf7_0),.din(w_dff_A_3VmWHgRi8_0),.clk(gclk));
	jdff dff_A_N5nTT7Wf7_0(.dout(w_dff_A_EAuFS8nH9_0),.din(w_dff_A_N5nTT7Wf7_0),.clk(gclk));
	jdff dff_A_EAuFS8nH9_0(.dout(w_dff_A_PfbEqwEC2_0),.din(w_dff_A_EAuFS8nH9_0),.clk(gclk));
	jdff dff_A_PfbEqwEC2_0(.dout(w_dff_A_yMf15lEb7_0),.din(w_dff_A_PfbEqwEC2_0),.clk(gclk));
	jdff dff_A_yMf15lEb7_0(.dout(w_dff_A_0czaHG583_0),.din(w_dff_A_yMf15lEb7_0),.clk(gclk));
	jdff dff_A_0czaHG583_0(.dout(w_dff_A_NOk9F1RR3_0),.din(w_dff_A_0czaHG583_0),.clk(gclk));
	jdff dff_A_NOk9F1RR3_0(.dout(w_dff_A_4hbYQgSX9_0),.din(w_dff_A_NOk9F1RR3_0),.clk(gclk));
	jdff dff_A_4hbYQgSX9_0(.dout(w_dff_A_74pB983h9_0),.din(w_dff_A_4hbYQgSX9_0),.clk(gclk));
	jdff dff_A_74pB983h9_0(.dout(w_dff_A_jUnLpZRw1_0),.din(w_dff_A_74pB983h9_0),.clk(gclk));
	jdff dff_A_jUnLpZRw1_0(.dout(w_dff_A_JdlXYvSK0_0),.din(w_dff_A_jUnLpZRw1_0),.clk(gclk));
	jdff dff_A_JdlXYvSK0_0(.dout(G598),.din(w_dff_A_JdlXYvSK0_0),.clk(gclk));
	jdff dff_A_98gOsWEt3_2(.dout(w_dff_A_B0OFEQIp4_0),.din(w_dff_A_98gOsWEt3_2),.clk(gclk));
	jdff dff_A_B0OFEQIp4_0(.dout(w_dff_A_pZowCQg91_0),.din(w_dff_A_B0OFEQIp4_0),.clk(gclk));
	jdff dff_A_pZowCQg91_0(.dout(w_dff_A_JxmTd9VK4_0),.din(w_dff_A_pZowCQg91_0),.clk(gclk));
	jdff dff_A_JxmTd9VK4_0(.dout(w_dff_A_KDWIDx9X5_0),.din(w_dff_A_JxmTd9VK4_0),.clk(gclk));
	jdff dff_A_KDWIDx9X5_0(.dout(w_dff_A_NO8x4lF96_0),.din(w_dff_A_KDWIDx9X5_0),.clk(gclk));
	jdff dff_A_NO8x4lF96_0(.dout(w_dff_A_LHnw3tqh2_0),.din(w_dff_A_NO8x4lF96_0),.clk(gclk));
	jdff dff_A_LHnw3tqh2_0(.dout(w_dff_A_dFRJKTIY3_0),.din(w_dff_A_LHnw3tqh2_0),.clk(gclk));
	jdff dff_A_dFRJKTIY3_0(.dout(w_dff_A_jjWsjl0j0_0),.din(w_dff_A_dFRJKTIY3_0),.clk(gclk));
	jdff dff_A_jjWsjl0j0_0(.dout(w_dff_A_JSZIaNST4_0),.din(w_dff_A_jjWsjl0j0_0),.clk(gclk));
	jdff dff_A_JSZIaNST4_0(.dout(w_dff_A_JGkX3g258_0),.din(w_dff_A_JSZIaNST4_0),.clk(gclk));
	jdff dff_A_JGkX3g258_0(.dout(w_dff_A_p3EM4PfW2_0),.din(w_dff_A_JGkX3g258_0),.clk(gclk));
	jdff dff_A_p3EM4PfW2_0(.dout(w_dff_A_lk1kbily6_0),.din(w_dff_A_p3EM4PfW2_0),.clk(gclk));
	jdff dff_A_lk1kbily6_0(.dout(w_dff_A_fFQcJEqi8_0),.din(w_dff_A_lk1kbily6_0),.clk(gclk));
	jdff dff_A_fFQcJEqi8_0(.dout(w_dff_A_3aJOuQ8I3_0),.din(w_dff_A_fFQcJEqi8_0),.clk(gclk));
	jdff dff_A_3aJOuQ8I3_0(.dout(w_dff_A_fnbxQkNv3_0),.din(w_dff_A_3aJOuQ8I3_0),.clk(gclk));
	jdff dff_A_fnbxQkNv3_0(.dout(w_dff_A_W5jSJ4eO7_0),.din(w_dff_A_fnbxQkNv3_0),.clk(gclk));
	jdff dff_A_W5jSJ4eO7_0(.dout(G610),.din(w_dff_A_W5jSJ4eO7_0),.clk(gclk));
	jdff dff_A_a8FPstR07_2(.dout(w_dff_A_Y76EPjOu1_0),.din(w_dff_A_a8FPstR07_2),.clk(gclk));
	jdff dff_A_Y76EPjOu1_0(.dout(w_dff_A_4sK39zaX6_0),.din(w_dff_A_Y76EPjOu1_0),.clk(gclk));
	jdff dff_A_4sK39zaX6_0(.dout(w_dff_A_SmKTwjui8_0),.din(w_dff_A_4sK39zaX6_0),.clk(gclk));
	jdff dff_A_SmKTwjui8_0(.dout(w_dff_A_QCPup3ZN5_0),.din(w_dff_A_SmKTwjui8_0),.clk(gclk));
	jdff dff_A_QCPup3ZN5_0(.dout(w_dff_A_lsmNFQ1N9_0),.din(w_dff_A_QCPup3ZN5_0),.clk(gclk));
	jdff dff_A_lsmNFQ1N9_0(.dout(w_dff_A_Tf6AjAa66_0),.din(w_dff_A_lsmNFQ1N9_0),.clk(gclk));
	jdff dff_A_Tf6AjAa66_0(.dout(w_dff_A_cnKgS36D6_0),.din(w_dff_A_Tf6AjAa66_0),.clk(gclk));
	jdff dff_A_cnKgS36D6_0(.dout(w_dff_A_4qn29nex5_0),.din(w_dff_A_cnKgS36D6_0),.clk(gclk));
	jdff dff_A_4qn29nex5_0(.dout(w_dff_A_hkN3Y5US3_0),.din(w_dff_A_4qn29nex5_0),.clk(gclk));
	jdff dff_A_hkN3Y5US3_0(.dout(w_dff_A_YUuRk3Tf1_0),.din(w_dff_A_hkN3Y5US3_0),.clk(gclk));
	jdff dff_A_YUuRk3Tf1_0(.dout(w_dff_A_54INVPiv3_0),.din(w_dff_A_YUuRk3Tf1_0),.clk(gclk));
	jdff dff_A_54INVPiv3_0(.dout(w_dff_A_J4ZslZdO7_0),.din(w_dff_A_54INVPiv3_0),.clk(gclk));
	jdff dff_A_J4ZslZdO7_0(.dout(w_dff_A_TptopMkg5_0),.din(w_dff_A_J4ZslZdO7_0),.clk(gclk));
	jdff dff_A_TptopMkg5_0(.dout(w_dff_A_oXwBPp741_0),.din(w_dff_A_TptopMkg5_0),.clk(gclk));
	jdff dff_A_oXwBPp741_0(.dout(G588),.din(w_dff_A_oXwBPp741_0),.clk(gclk));
	jdff dff_A_iLCWaaL96_2(.dout(w_dff_A_0RjeCt8U2_0),.din(w_dff_A_iLCWaaL96_2),.clk(gclk));
	jdff dff_A_0RjeCt8U2_0(.dout(w_dff_A_6FaBFqCk0_0),.din(w_dff_A_0RjeCt8U2_0),.clk(gclk));
	jdff dff_A_6FaBFqCk0_0(.dout(w_dff_A_usc74RgE8_0),.din(w_dff_A_6FaBFqCk0_0),.clk(gclk));
	jdff dff_A_usc74RgE8_0(.dout(w_dff_A_4ihPoDKK8_0),.din(w_dff_A_usc74RgE8_0),.clk(gclk));
	jdff dff_A_4ihPoDKK8_0(.dout(w_dff_A_14ba03835_0),.din(w_dff_A_4ihPoDKK8_0),.clk(gclk));
	jdff dff_A_14ba03835_0(.dout(w_dff_A_KYCdHPsg0_0),.din(w_dff_A_14ba03835_0),.clk(gclk));
	jdff dff_A_KYCdHPsg0_0(.dout(w_dff_A_UBujfgeH7_0),.din(w_dff_A_KYCdHPsg0_0),.clk(gclk));
	jdff dff_A_UBujfgeH7_0(.dout(w_dff_A_pYNG3d568_0),.din(w_dff_A_UBujfgeH7_0),.clk(gclk));
	jdff dff_A_pYNG3d568_0(.dout(w_dff_A_Cv7jV60I6_0),.din(w_dff_A_pYNG3d568_0),.clk(gclk));
	jdff dff_A_Cv7jV60I6_0(.dout(w_dff_A_b6iYVehc4_0),.din(w_dff_A_Cv7jV60I6_0),.clk(gclk));
	jdff dff_A_b6iYVehc4_0(.dout(w_dff_A_N1ZFTzWl2_0),.din(w_dff_A_b6iYVehc4_0),.clk(gclk));
	jdff dff_A_N1ZFTzWl2_0(.dout(w_dff_A_IHL1tGRu8_0),.din(w_dff_A_N1ZFTzWl2_0),.clk(gclk));
	jdff dff_A_IHL1tGRu8_0(.dout(w_dff_A_0twmngdc0_0),.din(w_dff_A_IHL1tGRu8_0),.clk(gclk));
	jdff dff_A_0twmngdc0_0(.dout(w_dff_A_5zaUQwQ88_0),.din(w_dff_A_0twmngdc0_0),.clk(gclk));
	jdff dff_A_5zaUQwQ88_0(.dout(w_dff_A_9IYrsimw1_0),.din(w_dff_A_5zaUQwQ88_0),.clk(gclk));
	jdff dff_A_9IYrsimw1_0(.dout(w_dff_A_AAXedV3U9_0),.din(w_dff_A_9IYrsimw1_0),.clk(gclk));
	jdff dff_A_AAXedV3U9_0(.dout(G615),.din(w_dff_A_AAXedV3U9_0),.clk(gclk));
	jdff dff_A_Y2JNsu3g3_2(.dout(w_dff_A_vUBCUwcC5_0),.din(w_dff_A_Y2JNsu3g3_2),.clk(gclk));
	jdff dff_A_vUBCUwcC5_0(.dout(w_dff_A_QYMabMA04_0),.din(w_dff_A_vUBCUwcC5_0),.clk(gclk));
	jdff dff_A_QYMabMA04_0(.dout(w_dff_A_Fp0HoExl9_0),.din(w_dff_A_QYMabMA04_0),.clk(gclk));
	jdff dff_A_Fp0HoExl9_0(.dout(w_dff_A_jw9xzuQn0_0),.din(w_dff_A_Fp0HoExl9_0),.clk(gclk));
	jdff dff_A_jw9xzuQn0_0(.dout(w_dff_A_V9msACep6_0),.din(w_dff_A_jw9xzuQn0_0),.clk(gclk));
	jdff dff_A_V9msACep6_0(.dout(w_dff_A_s5Ti432w4_0),.din(w_dff_A_V9msACep6_0),.clk(gclk));
	jdff dff_A_s5Ti432w4_0(.dout(w_dff_A_HSgIQdQZ1_0),.din(w_dff_A_s5Ti432w4_0),.clk(gclk));
	jdff dff_A_HSgIQdQZ1_0(.dout(w_dff_A_pyUPLJAW7_0),.din(w_dff_A_HSgIQdQZ1_0),.clk(gclk));
	jdff dff_A_pyUPLJAW7_0(.dout(w_dff_A_upNVlbE39_0),.din(w_dff_A_pyUPLJAW7_0),.clk(gclk));
	jdff dff_A_upNVlbE39_0(.dout(w_dff_A_dwo7mkOJ1_0),.din(w_dff_A_upNVlbE39_0),.clk(gclk));
	jdff dff_A_dwo7mkOJ1_0(.dout(w_dff_A_WpLPLNHG7_0),.din(w_dff_A_dwo7mkOJ1_0),.clk(gclk));
	jdff dff_A_WpLPLNHG7_0(.dout(w_dff_A_rd5YAnOU5_0),.din(w_dff_A_WpLPLNHG7_0),.clk(gclk));
	jdff dff_A_rd5YAnOU5_0(.dout(w_dff_A_xV3QuAoi6_0),.din(w_dff_A_rd5YAnOU5_0),.clk(gclk));
	jdff dff_A_xV3QuAoi6_0(.dout(w_dff_A_tZrQMKIb6_0),.din(w_dff_A_xV3QuAoi6_0),.clk(gclk));
	jdff dff_A_tZrQMKIb6_0(.dout(w_dff_A_omVFdhgg0_0),.din(w_dff_A_tZrQMKIb6_0),.clk(gclk));
	jdff dff_A_omVFdhgg0_0(.dout(w_dff_A_LW7XAMXs6_0),.din(w_dff_A_omVFdhgg0_0),.clk(gclk));
	jdff dff_A_LW7XAMXs6_0(.dout(G626),.din(w_dff_A_LW7XAMXs6_0),.clk(gclk));
	jdff dff_A_ILZVgwZy8_2(.dout(w_dff_A_PQlf6GMd2_0),.din(w_dff_A_ILZVgwZy8_2),.clk(gclk));
	jdff dff_A_PQlf6GMd2_0(.dout(w_dff_A_Mwot3wa29_0),.din(w_dff_A_PQlf6GMd2_0),.clk(gclk));
	jdff dff_A_Mwot3wa29_0(.dout(w_dff_A_JRabvF5G4_0),.din(w_dff_A_Mwot3wa29_0),.clk(gclk));
	jdff dff_A_JRabvF5G4_0(.dout(w_dff_A_vW0Eyizj4_0),.din(w_dff_A_JRabvF5G4_0),.clk(gclk));
	jdff dff_A_vW0Eyizj4_0(.dout(w_dff_A_6d9O58BP4_0),.din(w_dff_A_vW0Eyizj4_0),.clk(gclk));
	jdff dff_A_6d9O58BP4_0(.dout(w_dff_A_50drFKUZ0_0),.din(w_dff_A_6d9O58BP4_0),.clk(gclk));
	jdff dff_A_50drFKUZ0_0(.dout(w_dff_A_mszFQdJs6_0),.din(w_dff_A_50drFKUZ0_0),.clk(gclk));
	jdff dff_A_mszFQdJs6_0(.dout(w_dff_A_Ew9C0ilo8_0),.din(w_dff_A_mszFQdJs6_0),.clk(gclk));
	jdff dff_A_Ew9C0ilo8_0(.dout(w_dff_A_tkIG6ZIX9_0),.din(w_dff_A_Ew9C0ilo8_0),.clk(gclk));
	jdff dff_A_tkIG6ZIX9_0(.dout(w_dff_A_DhgW0GUa4_0),.din(w_dff_A_tkIG6ZIX9_0),.clk(gclk));
	jdff dff_A_DhgW0GUa4_0(.dout(w_dff_A_SRsdwpud5_0),.din(w_dff_A_DhgW0GUa4_0),.clk(gclk));
	jdff dff_A_SRsdwpud5_0(.dout(w_dff_A_jQSc5UrE5_0),.din(w_dff_A_SRsdwpud5_0),.clk(gclk));
	jdff dff_A_jQSc5UrE5_0(.dout(w_dff_A_2YFZ3K0t2_0),.din(w_dff_A_jQSc5UrE5_0),.clk(gclk));
	jdff dff_A_2YFZ3K0t2_0(.dout(w_dff_A_OLiViglB7_0),.din(w_dff_A_2YFZ3K0t2_0),.clk(gclk));
	jdff dff_A_OLiViglB7_0(.dout(G632),.din(w_dff_A_OLiViglB7_0),.clk(gclk));
	jdff dff_A_1v2VW66l6_1(.dout(w_dff_A_Ira4mwGl4_0),.din(w_dff_A_1v2VW66l6_1),.clk(gclk));
	jdff dff_A_Ira4mwGl4_0(.dout(w_dff_A_KjHPCE8R2_0),.din(w_dff_A_Ira4mwGl4_0),.clk(gclk));
	jdff dff_A_KjHPCE8R2_0(.dout(w_dff_A_b0b7x1cQ1_0),.din(w_dff_A_KjHPCE8R2_0),.clk(gclk));
	jdff dff_A_b0b7x1cQ1_0(.dout(w_dff_A_5thJ7mpQ6_0),.din(w_dff_A_b0b7x1cQ1_0),.clk(gclk));
	jdff dff_A_5thJ7mpQ6_0(.dout(w_dff_A_nzSsYxOa7_0),.din(w_dff_A_5thJ7mpQ6_0),.clk(gclk));
	jdff dff_A_nzSsYxOa7_0(.dout(w_dff_A_wnSh4jIM9_0),.din(w_dff_A_nzSsYxOa7_0),.clk(gclk));
	jdff dff_A_wnSh4jIM9_0(.dout(w_dff_A_oIUb7XkB7_0),.din(w_dff_A_wnSh4jIM9_0),.clk(gclk));
	jdff dff_A_oIUb7XkB7_0(.dout(w_dff_A_Iy5RohBW1_0),.din(w_dff_A_oIUb7XkB7_0),.clk(gclk));
	jdff dff_A_Iy5RohBW1_0(.dout(w_dff_A_fagOtbE00_0),.din(w_dff_A_Iy5RohBW1_0),.clk(gclk));
	jdff dff_A_fagOtbE00_0(.dout(w_dff_A_gPSsUOWk0_0),.din(w_dff_A_fagOtbE00_0),.clk(gclk));
	jdff dff_A_gPSsUOWk0_0(.dout(w_dff_A_REk4iN1w1_0),.din(w_dff_A_gPSsUOWk0_0),.clk(gclk));
	jdff dff_A_REk4iN1w1_0(.dout(w_dff_A_Xgayo0G98_0),.din(w_dff_A_REk4iN1w1_0),.clk(gclk));
	jdff dff_A_Xgayo0G98_0(.dout(w_dff_A_isge7Zwi0_0),.din(w_dff_A_Xgayo0G98_0),.clk(gclk));
	jdff dff_A_isge7Zwi0_0(.dout(w_dff_A_GXS5mcUB4_0),.din(w_dff_A_isge7Zwi0_0),.clk(gclk));
	jdff dff_A_GXS5mcUB4_0(.dout(w_dff_A_SGceFbLn2_0),.din(w_dff_A_GXS5mcUB4_0),.clk(gclk));
	jdff dff_A_SGceFbLn2_0(.dout(w_dff_A_dEhmY3mf2_0),.din(w_dff_A_SGceFbLn2_0),.clk(gclk));
	jdff dff_A_dEhmY3mf2_0(.dout(w_dff_A_AXx7NQnL9_0),.din(w_dff_A_dEhmY3mf2_0),.clk(gclk));
	jdff dff_A_AXx7NQnL9_0(.dout(w_dff_A_lkZKFyOo3_0),.din(w_dff_A_AXx7NQnL9_0),.clk(gclk));
	jdff dff_A_lkZKFyOo3_0(.dout(w_dff_A_QUueERQi5_0),.din(w_dff_A_lkZKFyOo3_0),.clk(gclk));
	jdff dff_A_QUueERQi5_0(.dout(w_dff_A_aZNTGliG6_0),.din(w_dff_A_QUueERQi5_0),.clk(gclk));
	jdff dff_A_aZNTGliG6_0(.dout(G1002),.din(w_dff_A_aZNTGliG6_0),.clk(gclk));
	jdff dff_A_nMfNfIJ88_1(.dout(w_dff_A_aia6tAyR1_0),.din(w_dff_A_nMfNfIJ88_1),.clk(gclk));
	jdff dff_A_aia6tAyR1_0(.dout(w_dff_A_3ZJMfTKa0_0),.din(w_dff_A_aia6tAyR1_0),.clk(gclk));
	jdff dff_A_3ZJMfTKa0_0(.dout(w_dff_A_BqJGGqG23_0),.din(w_dff_A_3ZJMfTKa0_0),.clk(gclk));
	jdff dff_A_BqJGGqG23_0(.dout(w_dff_A_QQOReGzZ6_0),.din(w_dff_A_BqJGGqG23_0),.clk(gclk));
	jdff dff_A_QQOReGzZ6_0(.dout(w_dff_A_vTtqk7PU2_0),.din(w_dff_A_QQOReGzZ6_0),.clk(gclk));
	jdff dff_A_vTtqk7PU2_0(.dout(w_dff_A_xHaQ98584_0),.din(w_dff_A_vTtqk7PU2_0),.clk(gclk));
	jdff dff_A_xHaQ98584_0(.dout(w_dff_A_tax63zYn0_0),.din(w_dff_A_xHaQ98584_0),.clk(gclk));
	jdff dff_A_tax63zYn0_0(.dout(w_dff_A_OuQBdFaA4_0),.din(w_dff_A_tax63zYn0_0),.clk(gclk));
	jdff dff_A_OuQBdFaA4_0(.dout(w_dff_A_vAKZcCet1_0),.din(w_dff_A_OuQBdFaA4_0),.clk(gclk));
	jdff dff_A_vAKZcCet1_0(.dout(w_dff_A_iMuTPVJI2_0),.din(w_dff_A_vAKZcCet1_0),.clk(gclk));
	jdff dff_A_iMuTPVJI2_0(.dout(w_dff_A_KboyahDh7_0),.din(w_dff_A_iMuTPVJI2_0),.clk(gclk));
	jdff dff_A_KboyahDh7_0(.dout(w_dff_A_rtJ5pmdO1_0),.din(w_dff_A_KboyahDh7_0),.clk(gclk));
	jdff dff_A_rtJ5pmdO1_0(.dout(w_dff_A_gcRAxrbN8_0),.din(w_dff_A_rtJ5pmdO1_0),.clk(gclk));
	jdff dff_A_gcRAxrbN8_0(.dout(w_dff_A_g4C1Kh1p8_0),.din(w_dff_A_gcRAxrbN8_0),.clk(gclk));
	jdff dff_A_g4C1Kh1p8_0(.dout(w_dff_A_KEATrYLB3_0),.din(w_dff_A_g4C1Kh1p8_0),.clk(gclk));
	jdff dff_A_KEATrYLB3_0(.dout(w_dff_A_U7D0JHqV1_0),.din(w_dff_A_KEATrYLB3_0),.clk(gclk));
	jdff dff_A_U7D0JHqV1_0(.dout(w_dff_A_PTdGLIUt1_0),.din(w_dff_A_U7D0JHqV1_0),.clk(gclk));
	jdff dff_A_PTdGLIUt1_0(.dout(w_dff_A_dLTj28wV3_0),.din(w_dff_A_PTdGLIUt1_0),.clk(gclk));
	jdff dff_A_dLTj28wV3_0(.dout(w_dff_A_RuScc4Lg1_0),.din(w_dff_A_dLTj28wV3_0),.clk(gclk));
	jdff dff_A_RuScc4Lg1_0(.dout(w_dff_A_oLmbBiYt2_0),.din(w_dff_A_RuScc4Lg1_0),.clk(gclk));
	jdff dff_A_oLmbBiYt2_0(.dout(G1004),.din(w_dff_A_oLmbBiYt2_0),.clk(gclk));
	jdff dff_A_oGRN7NsA0_2(.dout(w_dff_A_HCSwzBOJ5_0),.din(w_dff_A_oGRN7NsA0_2),.clk(gclk));
	jdff dff_A_HCSwzBOJ5_0(.dout(w_dff_A_fN03UcI28_0),.din(w_dff_A_HCSwzBOJ5_0),.clk(gclk));
	jdff dff_A_fN03UcI28_0(.dout(w_dff_A_htbl4Arh5_0),.din(w_dff_A_fN03UcI28_0),.clk(gclk));
	jdff dff_A_htbl4Arh5_0(.dout(w_dff_A_qikab3oX8_0),.din(w_dff_A_htbl4Arh5_0),.clk(gclk));
	jdff dff_A_qikab3oX8_0(.dout(w_dff_A_WWLLOsE74_0),.din(w_dff_A_qikab3oX8_0),.clk(gclk));
	jdff dff_A_WWLLOsE74_0(.dout(w_dff_A_k5QyiATD7_0),.din(w_dff_A_WWLLOsE74_0),.clk(gclk));
	jdff dff_A_k5QyiATD7_0(.dout(w_dff_A_T3WfK5JS4_0),.din(w_dff_A_k5QyiATD7_0),.clk(gclk));
	jdff dff_A_T3WfK5JS4_0(.dout(w_dff_A_HgUm4Wfm5_0),.din(w_dff_A_T3WfK5JS4_0),.clk(gclk));
	jdff dff_A_HgUm4Wfm5_0(.dout(w_dff_A_PIB0gAmo8_0),.din(w_dff_A_HgUm4Wfm5_0),.clk(gclk));
	jdff dff_A_PIB0gAmo8_0(.dout(w_dff_A_iUmsnd2u0_0),.din(w_dff_A_PIB0gAmo8_0),.clk(gclk));
	jdff dff_A_iUmsnd2u0_0(.dout(w_dff_A_LgYyAyff6_0),.din(w_dff_A_iUmsnd2u0_0),.clk(gclk));
	jdff dff_A_LgYyAyff6_0(.dout(G591),.din(w_dff_A_LgYyAyff6_0),.clk(gclk));
	jdff dff_A_M3kaUjHO8_2(.dout(w_dff_A_od9CFQac1_0),.din(w_dff_A_M3kaUjHO8_2),.clk(gclk));
	jdff dff_A_od9CFQac1_0(.dout(w_dff_A_nX9SPcRE3_0),.din(w_dff_A_od9CFQac1_0),.clk(gclk));
	jdff dff_A_nX9SPcRE3_0(.dout(w_dff_A_2n5ueYHb8_0),.din(w_dff_A_nX9SPcRE3_0),.clk(gclk));
	jdff dff_A_2n5ueYHb8_0(.dout(w_dff_A_JBAlqqQD3_0),.din(w_dff_A_2n5ueYHb8_0),.clk(gclk));
	jdff dff_A_JBAlqqQD3_0(.dout(w_dff_A_K7Le8zQa2_0),.din(w_dff_A_JBAlqqQD3_0),.clk(gclk));
	jdff dff_A_K7Le8zQa2_0(.dout(w_dff_A_QDFoqplF2_0),.din(w_dff_A_K7Le8zQa2_0),.clk(gclk));
	jdff dff_A_QDFoqplF2_0(.dout(w_dff_A_LgqFVPYY7_0),.din(w_dff_A_QDFoqplF2_0),.clk(gclk));
	jdff dff_A_LgqFVPYY7_0(.dout(w_dff_A_xfAN4HbR0_0),.din(w_dff_A_LgqFVPYY7_0),.clk(gclk));
	jdff dff_A_xfAN4HbR0_0(.dout(w_dff_A_Pwbwltpl3_0),.din(w_dff_A_xfAN4HbR0_0),.clk(gclk));
	jdff dff_A_Pwbwltpl3_0(.dout(w_dff_A_3Lxeulcw4_0),.din(w_dff_A_Pwbwltpl3_0),.clk(gclk));
	jdff dff_A_3Lxeulcw4_0(.dout(w_dff_A_ikhfFZ2b7_0),.din(w_dff_A_3Lxeulcw4_0),.clk(gclk));
	jdff dff_A_ikhfFZ2b7_0(.dout(G618),.din(w_dff_A_ikhfFZ2b7_0),.clk(gclk));
	jdff dff_A_k90aNcvw2_2(.dout(w_dff_A_kcddZhXl0_0),.din(w_dff_A_k90aNcvw2_2),.clk(gclk));
	jdff dff_A_kcddZhXl0_0(.dout(w_dff_A_oMly865h2_0),.din(w_dff_A_kcddZhXl0_0),.clk(gclk));
	jdff dff_A_oMly865h2_0(.dout(w_dff_A_RBF4SVrQ4_0),.din(w_dff_A_oMly865h2_0),.clk(gclk));
	jdff dff_A_RBF4SVrQ4_0(.dout(w_dff_A_6lx0kjh80_0),.din(w_dff_A_RBF4SVrQ4_0),.clk(gclk));
	jdff dff_A_6lx0kjh80_0(.dout(w_dff_A_u5xUUkRd4_0),.din(w_dff_A_6lx0kjh80_0),.clk(gclk));
	jdff dff_A_u5xUUkRd4_0(.dout(w_dff_A_K4xHwNqM3_0),.din(w_dff_A_u5xUUkRd4_0),.clk(gclk));
	jdff dff_A_K4xHwNqM3_0(.dout(w_dff_A_OAC6sqxy9_0),.din(w_dff_A_K4xHwNqM3_0),.clk(gclk));
	jdff dff_A_OAC6sqxy9_0(.dout(w_dff_A_XUAquFlY9_0),.din(w_dff_A_OAC6sqxy9_0),.clk(gclk));
	jdff dff_A_XUAquFlY9_0(.dout(w_dff_A_9mtx4GaW5_0),.din(w_dff_A_XUAquFlY9_0),.clk(gclk));
	jdff dff_A_9mtx4GaW5_0(.dout(w_dff_A_zkJmKRXE4_0),.din(w_dff_A_9mtx4GaW5_0),.clk(gclk));
	jdff dff_A_zkJmKRXE4_0(.dout(w_dff_A_WfnNI6MR0_0),.din(w_dff_A_zkJmKRXE4_0),.clk(gclk));
	jdff dff_A_WfnNI6MR0_0(.dout(G621),.din(w_dff_A_WfnNI6MR0_0),.clk(gclk));
	jdff dff_A_zku3LX0f7_2(.dout(w_dff_A_JkRydBe31_0),.din(w_dff_A_zku3LX0f7_2),.clk(gclk));
	jdff dff_A_JkRydBe31_0(.dout(w_dff_A_NvZPpkuv9_0),.din(w_dff_A_JkRydBe31_0),.clk(gclk));
	jdff dff_A_NvZPpkuv9_0(.dout(w_dff_A_icD3YL3o2_0),.din(w_dff_A_NvZPpkuv9_0),.clk(gclk));
	jdff dff_A_icD3YL3o2_0(.dout(w_dff_A_sEqoTvZ97_0),.din(w_dff_A_icD3YL3o2_0),.clk(gclk));
	jdff dff_A_sEqoTvZ97_0(.dout(w_dff_A_k3vzIK5t7_0),.din(w_dff_A_sEqoTvZ97_0),.clk(gclk));
	jdff dff_A_k3vzIK5t7_0(.dout(w_dff_A_UWZkjq8E7_0),.din(w_dff_A_k3vzIK5t7_0),.clk(gclk));
	jdff dff_A_UWZkjq8E7_0(.dout(w_dff_A_9oCgsZoT0_0),.din(w_dff_A_UWZkjq8E7_0),.clk(gclk));
	jdff dff_A_9oCgsZoT0_0(.dout(w_dff_A_ibtOhAEi6_0),.din(w_dff_A_9oCgsZoT0_0),.clk(gclk));
	jdff dff_A_ibtOhAEi6_0(.dout(w_dff_A_daXPEoIA9_0),.din(w_dff_A_ibtOhAEi6_0),.clk(gclk));
	jdff dff_A_daXPEoIA9_0(.dout(w_dff_A_cPbU9v4P8_0),.din(w_dff_A_daXPEoIA9_0),.clk(gclk));
	jdff dff_A_cPbU9v4P8_0(.dout(w_dff_A_EXRv7mO53_0),.din(w_dff_A_cPbU9v4P8_0),.clk(gclk));
	jdff dff_A_EXRv7mO53_0(.dout(G629),.din(w_dff_A_EXRv7mO53_0),.clk(gclk));
	jdff dff_A_q1tFT8lp8_1(.dout(w_dff_A_P44sLowh2_0),.din(w_dff_A_q1tFT8lp8_1),.clk(gclk));
	jdff dff_A_P44sLowh2_0(.dout(w_dff_A_eOPioVdF8_0),.din(w_dff_A_P44sLowh2_0),.clk(gclk));
	jdff dff_A_eOPioVdF8_0(.dout(w_dff_A_Jlrw9ktA1_0),.din(w_dff_A_eOPioVdF8_0),.clk(gclk));
	jdff dff_A_Jlrw9ktA1_0(.dout(w_dff_A_8F5vlDrx5_0),.din(w_dff_A_Jlrw9ktA1_0),.clk(gclk));
	jdff dff_A_8F5vlDrx5_0(.dout(w_dff_A_h3laRYog9_0),.din(w_dff_A_8F5vlDrx5_0),.clk(gclk));
	jdff dff_A_h3laRYog9_0(.dout(w_dff_A_MdCieRsr0_0),.din(w_dff_A_h3laRYog9_0),.clk(gclk));
	jdff dff_A_MdCieRsr0_0(.dout(w_dff_A_r547ROxf8_0),.din(w_dff_A_MdCieRsr0_0),.clk(gclk));
	jdff dff_A_r547ROxf8_0(.dout(w_dff_A_P4DjLPsY8_0),.din(w_dff_A_r547ROxf8_0),.clk(gclk));
	jdff dff_A_P4DjLPsY8_0(.dout(w_dff_A_aO3i0XEV3_0),.din(w_dff_A_P4DjLPsY8_0),.clk(gclk));
	jdff dff_A_aO3i0XEV3_0(.dout(w_dff_A_95qOkN0M0_0),.din(w_dff_A_aO3i0XEV3_0),.clk(gclk));
	jdff dff_A_95qOkN0M0_0(.dout(w_dff_A_N84C3P9f2_0),.din(w_dff_A_95qOkN0M0_0),.clk(gclk));
	jdff dff_A_N84C3P9f2_0(.dout(w_dff_A_QkcwueYH6_0),.din(w_dff_A_N84C3P9f2_0),.clk(gclk));
	jdff dff_A_QkcwueYH6_0(.dout(w_dff_A_WrAYzFoG5_0),.din(w_dff_A_QkcwueYH6_0),.clk(gclk));
	jdff dff_A_WrAYzFoG5_0(.dout(w_dff_A_8mFoipho1_0),.din(w_dff_A_WrAYzFoG5_0),.clk(gclk));
	jdff dff_A_8mFoipho1_0(.dout(w_dff_A_wHXTGEO89_0),.din(w_dff_A_8mFoipho1_0),.clk(gclk));
	jdff dff_A_wHXTGEO89_0(.dout(w_dff_A_2zND4OGL2_0),.din(w_dff_A_wHXTGEO89_0),.clk(gclk));
	jdff dff_A_2zND4OGL2_0(.dout(w_dff_A_9PbdJEEm1_0),.din(w_dff_A_2zND4OGL2_0),.clk(gclk));
	jdff dff_A_9PbdJEEm1_0(.dout(w_dff_A_2wxje0ys9_0),.din(w_dff_A_9PbdJEEm1_0),.clk(gclk));
	jdff dff_A_2wxje0ys9_0(.dout(G822),.din(w_dff_A_2wxje0ys9_0),.clk(gclk));
	jdff dff_A_AYO72yhU1_1(.dout(w_dff_A_XywcEaJ49_0),.din(w_dff_A_AYO72yhU1_1),.clk(gclk));
	jdff dff_A_XywcEaJ49_0(.dout(w_dff_A_s3udFBJ43_0),.din(w_dff_A_XywcEaJ49_0),.clk(gclk));
	jdff dff_A_s3udFBJ43_0(.dout(w_dff_A_dLPwlqWd0_0),.din(w_dff_A_s3udFBJ43_0),.clk(gclk));
	jdff dff_A_dLPwlqWd0_0(.dout(w_dff_A_jWz8xjl01_0),.din(w_dff_A_dLPwlqWd0_0),.clk(gclk));
	jdff dff_A_jWz8xjl01_0(.dout(w_dff_A_C6ioL0HG9_0),.din(w_dff_A_jWz8xjl01_0),.clk(gclk));
	jdff dff_A_C6ioL0HG9_0(.dout(w_dff_A_hCN6uBsO0_0),.din(w_dff_A_C6ioL0HG9_0),.clk(gclk));
	jdff dff_A_hCN6uBsO0_0(.dout(w_dff_A_Uggwwmxa7_0),.din(w_dff_A_hCN6uBsO0_0),.clk(gclk));
	jdff dff_A_Uggwwmxa7_0(.dout(w_dff_A_zkIZLCHX2_0),.din(w_dff_A_Uggwwmxa7_0),.clk(gclk));
	jdff dff_A_zkIZLCHX2_0(.dout(w_dff_A_W9cNDRiU2_0),.din(w_dff_A_zkIZLCHX2_0),.clk(gclk));
	jdff dff_A_W9cNDRiU2_0(.dout(w_dff_A_yFpiiRYf5_0),.din(w_dff_A_W9cNDRiU2_0),.clk(gclk));
	jdff dff_A_yFpiiRYf5_0(.dout(w_dff_A_TxhCSyiI7_0),.din(w_dff_A_yFpiiRYf5_0),.clk(gclk));
	jdff dff_A_TxhCSyiI7_0(.dout(w_dff_A_FAHrZ0hJ6_0),.din(w_dff_A_TxhCSyiI7_0),.clk(gclk));
	jdff dff_A_FAHrZ0hJ6_0(.dout(w_dff_A_FPqdRuPV2_0),.din(w_dff_A_FAHrZ0hJ6_0),.clk(gclk));
	jdff dff_A_FPqdRuPV2_0(.dout(w_dff_A_o2HfYUVo3_0),.din(w_dff_A_FPqdRuPV2_0),.clk(gclk));
	jdff dff_A_o2HfYUVo3_0(.dout(w_dff_A_W5WvkQ2T0_0),.din(w_dff_A_o2HfYUVo3_0),.clk(gclk));
	jdff dff_A_W5WvkQ2T0_0(.dout(w_dff_A_2L03ORBx3_0),.din(w_dff_A_W5WvkQ2T0_0),.clk(gclk));
	jdff dff_A_2L03ORBx3_0(.dout(w_dff_A_zh0iCaZF6_0),.din(w_dff_A_2L03ORBx3_0),.clk(gclk));
	jdff dff_A_zh0iCaZF6_0(.dout(G838),.din(w_dff_A_zh0iCaZF6_0),.clk(gclk));
	jdff dff_A_KfJFor9N7_1(.dout(w_dff_A_NN2k55lL9_0),.din(w_dff_A_KfJFor9N7_1),.clk(gclk));
	jdff dff_A_NN2k55lL9_0(.dout(w_dff_A_86GzOnGp2_0),.din(w_dff_A_NN2k55lL9_0),.clk(gclk));
	jdff dff_A_86GzOnGp2_0(.dout(w_dff_A_DZ79gRgf2_0),.din(w_dff_A_86GzOnGp2_0),.clk(gclk));
	jdff dff_A_DZ79gRgf2_0(.dout(w_dff_A_3bLamFKY7_0),.din(w_dff_A_DZ79gRgf2_0),.clk(gclk));
	jdff dff_A_3bLamFKY7_0(.dout(w_dff_A_5tuFy5kO6_0),.din(w_dff_A_3bLamFKY7_0),.clk(gclk));
	jdff dff_A_5tuFy5kO6_0(.dout(w_dff_A_PHA3kwzM4_0),.din(w_dff_A_5tuFy5kO6_0),.clk(gclk));
	jdff dff_A_PHA3kwzM4_0(.dout(w_dff_A_wGvFnnkW3_0),.din(w_dff_A_PHA3kwzM4_0),.clk(gclk));
	jdff dff_A_wGvFnnkW3_0(.dout(w_dff_A_Tj2n1Jc63_0),.din(w_dff_A_wGvFnnkW3_0),.clk(gclk));
	jdff dff_A_Tj2n1Jc63_0(.dout(w_dff_A_r2RlglYq9_0),.din(w_dff_A_Tj2n1Jc63_0),.clk(gclk));
	jdff dff_A_r2RlglYq9_0(.dout(w_dff_A_4CCKekpJ0_0),.din(w_dff_A_r2RlglYq9_0),.clk(gclk));
	jdff dff_A_4CCKekpJ0_0(.dout(w_dff_A_FZGNVepn3_0),.din(w_dff_A_4CCKekpJ0_0),.clk(gclk));
	jdff dff_A_FZGNVepn3_0(.dout(w_dff_A_JOfdidDz0_0),.din(w_dff_A_FZGNVepn3_0),.clk(gclk));
	jdff dff_A_JOfdidDz0_0(.dout(w_dff_A_UschAx5w8_0),.din(w_dff_A_JOfdidDz0_0),.clk(gclk));
	jdff dff_A_UschAx5w8_0(.dout(w_dff_A_HOSW48Mq9_0),.din(w_dff_A_UschAx5w8_0),.clk(gclk));
	jdff dff_A_HOSW48Mq9_0(.dout(w_dff_A_wBkrJtwD1_0),.din(w_dff_A_HOSW48Mq9_0),.clk(gclk));
	jdff dff_A_wBkrJtwD1_0(.dout(w_dff_A_iAVYVYPd1_0),.din(w_dff_A_wBkrJtwD1_0),.clk(gclk));
	jdff dff_A_iAVYVYPd1_0(.dout(w_dff_A_Mhtqgaee2_0),.din(w_dff_A_iAVYVYPd1_0),.clk(gclk));
	jdff dff_A_Mhtqgaee2_0(.dout(G861),.din(w_dff_A_Mhtqgaee2_0),.clk(gclk));
	jdff dff_A_i69PVv1d1_1(.dout(w_dff_A_wOAaABEf7_0),.din(w_dff_A_i69PVv1d1_1),.clk(gclk));
	jdff dff_A_wOAaABEf7_0(.dout(w_dff_A_AktMmHI74_0),.din(w_dff_A_wOAaABEf7_0),.clk(gclk));
	jdff dff_A_AktMmHI74_0(.dout(w_dff_A_HO4H0c6d9_0),.din(w_dff_A_AktMmHI74_0),.clk(gclk));
	jdff dff_A_HO4H0c6d9_0(.dout(w_dff_A_vaiEItOd4_0),.din(w_dff_A_HO4H0c6d9_0),.clk(gclk));
	jdff dff_A_vaiEItOd4_0(.dout(w_dff_A_EIDCrBcL4_0),.din(w_dff_A_vaiEItOd4_0),.clk(gclk));
	jdff dff_A_EIDCrBcL4_0(.dout(w_dff_A_G45eVPtF1_0),.din(w_dff_A_EIDCrBcL4_0),.clk(gclk));
	jdff dff_A_G45eVPtF1_0(.dout(G623),.din(w_dff_A_G45eVPtF1_0),.clk(gclk));
	jdff dff_A_sV8pytjm1_2(.dout(w_dff_A_GTZ7yswP5_0),.din(w_dff_A_sV8pytjm1_2),.clk(gclk));
	jdff dff_A_GTZ7yswP5_0(.dout(w_dff_A_smA2jgin7_0),.din(w_dff_A_GTZ7yswP5_0),.clk(gclk));
	jdff dff_A_smA2jgin7_0(.dout(w_dff_A_hEttIOEH2_0),.din(w_dff_A_smA2jgin7_0),.clk(gclk));
	jdff dff_A_hEttIOEH2_0(.dout(w_dff_A_NoHJkvAX1_0),.din(w_dff_A_hEttIOEH2_0),.clk(gclk));
	jdff dff_A_NoHJkvAX1_0(.dout(w_dff_A_VRsR3txa9_0),.din(w_dff_A_NoHJkvAX1_0),.clk(gclk));
	jdff dff_A_VRsR3txa9_0(.dout(w_dff_A_JD23QiaJ4_0),.din(w_dff_A_VRsR3txa9_0),.clk(gclk));
	jdff dff_A_JD23QiaJ4_0(.dout(w_dff_A_gDWVLIAC8_0),.din(w_dff_A_JD23QiaJ4_0),.clk(gclk));
	jdff dff_A_gDWVLIAC8_0(.dout(w_dff_A_O4Px5IhQ0_0),.din(w_dff_A_gDWVLIAC8_0),.clk(gclk));
	jdff dff_A_O4Px5IhQ0_0(.dout(w_dff_A_Gfh6MIS83_0),.din(w_dff_A_O4Px5IhQ0_0),.clk(gclk));
	jdff dff_A_Gfh6MIS83_0(.dout(w_dff_A_yiJOh81W8_0),.din(w_dff_A_Gfh6MIS83_0),.clk(gclk));
	jdff dff_A_yiJOh81W8_0(.dout(w_dff_A_rxWA0Uww8_0),.din(w_dff_A_yiJOh81W8_0),.clk(gclk));
	jdff dff_A_rxWA0Uww8_0(.dout(w_dff_A_KXxs2KMA3_0),.din(w_dff_A_rxWA0Uww8_0),.clk(gclk));
	jdff dff_A_KXxs2KMA3_0(.dout(w_dff_A_NlauAOvK1_0),.din(w_dff_A_KXxs2KMA3_0),.clk(gclk));
	jdff dff_A_NlauAOvK1_0(.dout(w_dff_A_2PY7AmP71_0),.din(w_dff_A_NlauAOvK1_0),.clk(gclk));
	jdff dff_A_2PY7AmP71_0(.dout(G722),.din(w_dff_A_2PY7AmP71_0),.clk(gclk));
	jdff dff_A_0wXNdgG84_1(.dout(w_dff_A_Fv9CePF61_0),.din(w_dff_A_0wXNdgG84_1),.clk(gclk));
	jdff dff_A_Fv9CePF61_0(.dout(w_dff_A_9RJTjqSd6_0),.din(w_dff_A_Fv9CePF61_0),.clk(gclk));
	jdff dff_A_9RJTjqSd6_0(.dout(w_dff_A_8mtJ3sJX8_0),.din(w_dff_A_9RJTjqSd6_0),.clk(gclk));
	jdff dff_A_8mtJ3sJX8_0(.dout(w_dff_A_23Sc72Pf9_0),.din(w_dff_A_8mtJ3sJX8_0),.clk(gclk));
	jdff dff_A_23Sc72Pf9_0(.dout(w_dff_A_nKORoGTi4_0),.din(w_dff_A_23Sc72Pf9_0),.clk(gclk));
	jdff dff_A_nKORoGTi4_0(.dout(w_dff_A_Z1vwV1fg9_0),.din(w_dff_A_nKORoGTi4_0),.clk(gclk));
	jdff dff_A_Z1vwV1fg9_0(.dout(w_dff_A_6JVam7T38_0),.din(w_dff_A_Z1vwV1fg9_0),.clk(gclk));
	jdff dff_A_6JVam7T38_0(.dout(w_dff_A_kqO1J8L91_0),.din(w_dff_A_6JVam7T38_0),.clk(gclk));
	jdff dff_A_kqO1J8L91_0(.dout(w_dff_A_aC3wlJzx9_0),.din(w_dff_A_kqO1J8L91_0),.clk(gclk));
	jdff dff_A_aC3wlJzx9_0(.dout(w_dff_A_SdBkTOWy7_0),.din(w_dff_A_aC3wlJzx9_0),.clk(gclk));
	jdff dff_A_SdBkTOWy7_0(.dout(w_dff_A_1RqMgdJa1_0),.din(w_dff_A_SdBkTOWy7_0),.clk(gclk));
	jdff dff_A_1RqMgdJa1_0(.dout(G832),.din(w_dff_A_1RqMgdJa1_0),.clk(gclk));
	jdff dff_A_wKLlrNjI5_1(.dout(w_dff_A_MFK3SxBP6_0),.din(w_dff_A_wKLlrNjI5_1),.clk(gclk));
	jdff dff_A_MFK3SxBP6_0(.dout(w_dff_A_s4jXqwk55_0),.din(w_dff_A_MFK3SxBP6_0),.clk(gclk));
	jdff dff_A_s4jXqwk55_0(.dout(w_dff_A_n5q1i7FY9_0),.din(w_dff_A_s4jXqwk55_0),.clk(gclk));
	jdff dff_A_n5q1i7FY9_0(.dout(w_dff_A_ep3x9ehP5_0),.din(w_dff_A_n5q1i7FY9_0),.clk(gclk));
	jdff dff_A_ep3x9ehP5_0(.dout(w_dff_A_018dXP870_0),.din(w_dff_A_ep3x9ehP5_0),.clk(gclk));
	jdff dff_A_018dXP870_0(.dout(w_dff_A_7Ldy8DOA4_0),.din(w_dff_A_018dXP870_0),.clk(gclk));
	jdff dff_A_7Ldy8DOA4_0(.dout(w_dff_A_4OqwkNU43_0),.din(w_dff_A_7Ldy8DOA4_0),.clk(gclk));
	jdff dff_A_4OqwkNU43_0(.dout(w_dff_A_OQiNf4Hy1_0),.din(w_dff_A_4OqwkNU43_0),.clk(gclk));
	jdff dff_A_OQiNf4Hy1_0(.dout(w_dff_A_KXP7UABL8_0),.din(w_dff_A_OQiNf4Hy1_0),.clk(gclk));
	jdff dff_A_KXP7UABL8_0(.dout(w_dff_A_Gqcwnt1r2_0),.din(w_dff_A_KXP7UABL8_0),.clk(gclk));
	jdff dff_A_Gqcwnt1r2_0(.dout(w_dff_A_GJf4cJnl9_0),.din(w_dff_A_Gqcwnt1r2_0),.clk(gclk));
	jdff dff_A_GJf4cJnl9_0(.dout(w_dff_A_uhzzR6FF1_0),.din(w_dff_A_GJf4cJnl9_0),.clk(gclk));
	jdff dff_A_uhzzR6FF1_0(.dout(w_dff_A_Bv7ww4kQ5_0),.din(w_dff_A_uhzzR6FF1_0),.clk(gclk));
	jdff dff_A_Bv7ww4kQ5_0(.dout(G834),.din(w_dff_A_Bv7ww4kQ5_0),.clk(gclk));
	jdff dff_A_ScVFdJA46_1(.dout(w_dff_A_8lyBC1yo0_0),.din(w_dff_A_ScVFdJA46_1),.clk(gclk));
	jdff dff_A_8lyBC1yo0_0(.dout(w_dff_A_3rpw4Cls2_0),.din(w_dff_A_8lyBC1yo0_0),.clk(gclk));
	jdff dff_A_3rpw4Cls2_0(.dout(w_dff_A_IwlMcOzk0_0),.din(w_dff_A_3rpw4Cls2_0),.clk(gclk));
	jdff dff_A_IwlMcOzk0_0(.dout(w_dff_A_DQZ2UmjT7_0),.din(w_dff_A_IwlMcOzk0_0),.clk(gclk));
	jdff dff_A_DQZ2UmjT7_0(.dout(w_dff_A_a4mf9Bax4_0),.din(w_dff_A_DQZ2UmjT7_0),.clk(gclk));
	jdff dff_A_a4mf9Bax4_0(.dout(w_dff_A_gB1E08NY5_0),.din(w_dff_A_a4mf9Bax4_0),.clk(gclk));
	jdff dff_A_gB1E08NY5_0(.dout(w_dff_A_0PM042256_0),.din(w_dff_A_gB1E08NY5_0),.clk(gclk));
	jdff dff_A_0PM042256_0(.dout(w_dff_A_LQ7uBeoz3_0),.din(w_dff_A_0PM042256_0),.clk(gclk));
	jdff dff_A_LQ7uBeoz3_0(.dout(w_dff_A_dkVtVOUx5_0),.din(w_dff_A_LQ7uBeoz3_0),.clk(gclk));
	jdff dff_A_dkVtVOUx5_0(.dout(w_dff_A_HJzGzpIc0_0),.din(w_dff_A_dkVtVOUx5_0),.clk(gclk));
	jdff dff_A_HJzGzpIc0_0(.dout(w_dff_A_S4dd3pon7_0),.din(w_dff_A_HJzGzpIc0_0),.clk(gclk));
	jdff dff_A_S4dd3pon7_0(.dout(w_dff_A_6vceczxd9_0),.din(w_dff_A_S4dd3pon7_0),.clk(gclk));
	jdff dff_A_6vceczxd9_0(.dout(w_dff_A_uUkxmizt2_0),.din(w_dff_A_6vceczxd9_0),.clk(gclk));
	jdff dff_A_uUkxmizt2_0(.dout(w_dff_A_JD0ybVW66_0),.din(w_dff_A_uUkxmizt2_0),.clk(gclk));
	jdff dff_A_JD0ybVW66_0(.dout(w_dff_A_zo8Acg4y6_0),.din(w_dff_A_JD0ybVW66_0),.clk(gclk));
	jdff dff_A_zo8Acg4y6_0(.dout(G836),.din(w_dff_A_zo8Acg4y6_0),.clk(gclk));
	jdff dff_A_V0Jxk4lg2_2(.dout(w_dff_A_3fAq5jVR5_0),.din(w_dff_A_V0Jxk4lg2_2),.clk(gclk));
	jdff dff_A_3fAq5jVR5_0(.dout(w_dff_A_JreTsS6M8_0),.din(w_dff_A_3fAq5jVR5_0),.clk(gclk));
	jdff dff_A_JreTsS6M8_0(.dout(w_dff_A_F36WOgGT9_0),.din(w_dff_A_JreTsS6M8_0),.clk(gclk));
	jdff dff_A_F36WOgGT9_0(.dout(w_dff_A_6RaYDjH62_0),.din(w_dff_A_F36WOgGT9_0),.clk(gclk));
	jdff dff_A_6RaYDjH62_0(.dout(w_dff_A_0JSxN4jW6_0),.din(w_dff_A_6RaYDjH62_0),.clk(gclk));
	jdff dff_A_0JSxN4jW6_0(.dout(w_dff_A_NGaX2Gbd8_0),.din(w_dff_A_0JSxN4jW6_0),.clk(gclk));
	jdff dff_A_NGaX2Gbd8_0(.dout(w_dff_A_icfMg0JI1_0),.din(w_dff_A_NGaX2Gbd8_0),.clk(gclk));
	jdff dff_A_icfMg0JI1_0(.dout(w_dff_A_8rfjwdNr7_0),.din(w_dff_A_icfMg0JI1_0),.clk(gclk));
	jdff dff_A_8rfjwdNr7_0(.dout(w_dff_A_cwR4FYFA7_0),.din(w_dff_A_8rfjwdNr7_0),.clk(gclk));
	jdff dff_A_cwR4FYFA7_0(.dout(w_dff_A_VD44ma169_0),.din(w_dff_A_cwR4FYFA7_0),.clk(gclk));
	jdff dff_A_VD44ma169_0(.dout(w_dff_A_tcCrlzQ04_0),.din(w_dff_A_VD44ma169_0),.clk(gclk));
	jdff dff_A_tcCrlzQ04_0(.dout(w_dff_A_rvBYlond9_0),.din(w_dff_A_tcCrlzQ04_0),.clk(gclk));
	jdff dff_A_rvBYlond9_0(.dout(w_dff_A_kqInnoN63_0),.din(w_dff_A_rvBYlond9_0),.clk(gclk));
	jdff dff_A_kqInnoN63_0(.dout(w_dff_A_2jvwvDog9_0),.din(w_dff_A_kqInnoN63_0),.clk(gclk));
	jdff dff_A_2jvwvDog9_0(.dout(G859),.din(w_dff_A_2jvwvDog9_0),.clk(gclk));
	jdff dff_A_xqc4ukvK3_1(.dout(w_dff_A_lN3QgUuj6_0),.din(w_dff_A_xqc4ukvK3_1),.clk(gclk));
	jdff dff_A_lN3QgUuj6_0(.dout(w_dff_A_qlI3RfQY3_0),.din(w_dff_A_lN3QgUuj6_0),.clk(gclk));
	jdff dff_A_qlI3RfQY3_0(.dout(w_dff_A_OVUrvpWZ7_0),.din(w_dff_A_qlI3RfQY3_0),.clk(gclk));
	jdff dff_A_OVUrvpWZ7_0(.dout(w_dff_A_DPxXXKgb9_0),.din(w_dff_A_OVUrvpWZ7_0),.clk(gclk));
	jdff dff_A_DPxXXKgb9_0(.dout(w_dff_A_PRENhfcU9_0),.din(w_dff_A_DPxXXKgb9_0),.clk(gclk));
	jdff dff_A_PRENhfcU9_0(.dout(w_dff_A_c6EHn7EM2_0),.din(w_dff_A_PRENhfcU9_0),.clk(gclk));
	jdff dff_A_c6EHn7EM2_0(.dout(w_dff_A_9YirO3EP8_0),.din(w_dff_A_c6EHn7EM2_0),.clk(gclk));
	jdff dff_A_9YirO3EP8_0(.dout(w_dff_A_e3LLgrUR6_0),.din(w_dff_A_9YirO3EP8_0),.clk(gclk));
	jdff dff_A_e3LLgrUR6_0(.dout(w_dff_A_YdeDvYTh5_0),.din(w_dff_A_e3LLgrUR6_0),.clk(gclk));
	jdff dff_A_YdeDvYTh5_0(.dout(G871),.din(w_dff_A_YdeDvYTh5_0),.clk(gclk));
	jdff dff_A_R11IaAAo2_1(.dout(w_dff_A_34wxYVgv2_0),.din(w_dff_A_R11IaAAo2_1),.clk(gclk));
	jdff dff_A_34wxYVgv2_0(.dout(w_dff_A_aMsFzV8k2_0),.din(w_dff_A_34wxYVgv2_0),.clk(gclk));
	jdff dff_A_aMsFzV8k2_0(.dout(w_dff_A_f2iSOEjN8_0),.din(w_dff_A_aMsFzV8k2_0),.clk(gclk));
	jdff dff_A_f2iSOEjN8_0(.dout(w_dff_A_4jZyDO4a2_0),.din(w_dff_A_f2iSOEjN8_0),.clk(gclk));
	jdff dff_A_4jZyDO4a2_0(.dout(w_dff_A_6KvbrMhZ3_0),.din(w_dff_A_4jZyDO4a2_0),.clk(gclk));
	jdff dff_A_6KvbrMhZ3_0(.dout(w_dff_A_yn9p9jYD3_0),.din(w_dff_A_6KvbrMhZ3_0),.clk(gclk));
	jdff dff_A_yn9p9jYD3_0(.dout(w_dff_A_BI9Q3Wlq4_0),.din(w_dff_A_yn9p9jYD3_0),.clk(gclk));
	jdff dff_A_BI9Q3Wlq4_0(.dout(w_dff_A_iFNhOtGr8_0),.din(w_dff_A_BI9Q3Wlq4_0),.clk(gclk));
	jdff dff_A_iFNhOtGr8_0(.dout(w_dff_A_PumRsgop7_0),.din(w_dff_A_iFNhOtGr8_0),.clk(gclk));
	jdff dff_A_PumRsgop7_0(.dout(w_dff_A_pPGSV0VE7_0),.din(w_dff_A_PumRsgop7_0),.clk(gclk));
	jdff dff_A_pPGSV0VE7_0(.dout(w_dff_A_VrTxVwbE1_0),.din(w_dff_A_pPGSV0VE7_0),.clk(gclk));
	jdff dff_A_VrTxVwbE1_0(.dout(G873),.din(w_dff_A_VrTxVwbE1_0),.clk(gclk));
	jdff dff_A_UWtWUJzu5_1(.dout(w_dff_A_39IcbON36_0),.din(w_dff_A_UWtWUJzu5_1),.clk(gclk));
	jdff dff_A_39IcbON36_0(.dout(w_dff_A_FYxACZtd5_0),.din(w_dff_A_39IcbON36_0),.clk(gclk));
	jdff dff_A_FYxACZtd5_0(.dout(w_dff_A_ayPqb62j7_0),.din(w_dff_A_FYxACZtd5_0),.clk(gclk));
	jdff dff_A_ayPqb62j7_0(.dout(w_dff_A_nkWawfgl9_0),.din(w_dff_A_ayPqb62j7_0),.clk(gclk));
	jdff dff_A_nkWawfgl9_0(.dout(w_dff_A_35pPbuLW8_0),.din(w_dff_A_nkWawfgl9_0),.clk(gclk));
	jdff dff_A_35pPbuLW8_0(.dout(w_dff_A_PV0eDmLD2_0),.din(w_dff_A_35pPbuLW8_0),.clk(gclk));
	jdff dff_A_PV0eDmLD2_0(.dout(w_dff_A_Q5O5yeK04_0),.din(w_dff_A_PV0eDmLD2_0),.clk(gclk));
	jdff dff_A_Q5O5yeK04_0(.dout(w_dff_A_dPif8dpM3_0),.din(w_dff_A_Q5O5yeK04_0),.clk(gclk));
	jdff dff_A_dPif8dpM3_0(.dout(w_dff_A_lSAPL9oN3_0),.din(w_dff_A_dPif8dpM3_0),.clk(gclk));
	jdff dff_A_lSAPL9oN3_0(.dout(w_dff_A_Aptn8CNa9_0),.din(w_dff_A_lSAPL9oN3_0),.clk(gclk));
	jdff dff_A_Aptn8CNa9_0(.dout(w_dff_A_JaIYGaxb7_0),.din(w_dff_A_Aptn8CNa9_0),.clk(gclk));
	jdff dff_A_JaIYGaxb7_0(.dout(w_dff_A_NhEquGyl5_0),.din(w_dff_A_JaIYGaxb7_0),.clk(gclk));
	jdff dff_A_NhEquGyl5_0(.dout(G875),.din(w_dff_A_NhEquGyl5_0),.clk(gclk));
	jdff dff_A_cO0UkzHS2_1(.dout(w_dff_A_ip7BzEE51_0),.din(w_dff_A_cO0UkzHS2_1),.clk(gclk));
	jdff dff_A_ip7BzEE51_0(.dout(w_dff_A_BAXNnSZN6_0),.din(w_dff_A_ip7BzEE51_0),.clk(gclk));
	jdff dff_A_BAXNnSZN6_0(.dout(w_dff_A_uvL9Ps9j7_0),.din(w_dff_A_BAXNnSZN6_0),.clk(gclk));
	jdff dff_A_uvL9Ps9j7_0(.dout(w_dff_A_Niz0Sftl6_0),.din(w_dff_A_uvL9Ps9j7_0),.clk(gclk));
	jdff dff_A_Niz0Sftl6_0(.dout(w_dff_A_AbRH6wS81_0),.din(w_dff_A_Niz0Sftl6_0),.clk(gclk));
	jdff dff_A_AbRH6wS81_0(.dout(w_dff_A_52SqaebH2_0),.din(w_dff_A_AbRH6wS81_0),.clk(gclk));
	jdff dff_A_52SqaebH2_0(.dout(w_dff_A_0z11elp72_0),.din(w_dff_A_52SqaebH2_0),.clk(gclk));
	jdff dff_A_0z11elp72_0(.dout(w_dff_A_wbxJ4dX05_0),.din(w_dff_A_0z11elp72_0),.clk(gclk));
	jdff dff_A_wbxJ4dX05_0(.dout(w_dff_A_PhSOUEfc0_0),.din(w_dff_A_wbxJ4dX05_0),.clk(gclk));
	jdff dff_A_PhSOUEfc0_0(.dout(w_dff_A_bEapAac94_0),.din(w_dff_A_PhSOUEfc0_0),.clk(gclk));
	jdff dff_A_bEapAac94_0(.dout(w_dff_A_H8DrywDq1_0),.din(w_dff_A_bEapAac94_0),.clk(gclk));
	jdff dff_A_H8DrywDq1_0(.dout(w_dff_A_gGj9Yd925_0),.din(w_dff_A_H8DrywDq1_0),.clk(gclk));
	jdff dff_A_gGj9Yd925_0(.dout(w_dff_A_OiVSYWaj6_0),.din(w_dff_A_gGj9Yd925_0),.clk(gclk));
	jdff dff_A_OiVSYWaj6_0(.dout(G877),.din(w_dff_A_OiVSYWaj6_0),.clk(gclk));
	jdff dff_A_XkoNU5Q13_1(.dout(w_dff_A_RKrC5ZHB3_0),.din(w_dff_A_XkoNU5Q13_1),.clk(gclk));
	jdff dff_A_RKrC5ZHB3_0(.dout(w_dff_A_Czml2uA94_0),.din(w_dff_A_RKrC5ZHB3_0),.clk(gclk));
	jdff dff_A_Czml2uA94_0(.dout(w_dff_A_B0VxtW2z7_0),.din(w_dff_A_Czml2uA94_0),.clk(gclk));
	jdff dff_A_B0VxtW2z7_0(.dout(w_dff_A_5gFIGXCd4_0),.din(w_dff_A_B0VxtW2z7_0),.clk(gclk));
	jdff dff_A_5gFIGXCd4_0(.dout(w_dff_A_g1LOYUUf7_0),.din(w_dff_A_5gFIGXCd4_0),.clk(gclk));
	jdff dff_A_g1LOYUUf7_0(.dout(w_dff_A_zQTHNMeU9_0),.din(w_dff_A_g1LOYUUf7_0),.clk(gclk));
	jdff dff_A_zQTHNMeU9_0(.dout(w_dff_A_irAHEeFG0_0),.din(w_dff_A_zQTHNMeU9_0),.clk(gclk));
	jdff dff_A_irAHEeFG0_0(.dout(w_dff_A_n8FKUin47_0),.din(w_dff_A_irAHEeFG0_0),.clk(gclk));
	jdff dff_A_n8FKUin47_0(.dout(w_dff_A_MWSLrTf99_0),.din(w_dff_A_n8FKUin47_0),.clk(gclk));
	jdff dff_A_MWSLrTf99_0(.dout(w_dff_A_9qqlxDDT8_0),.din(w_dff_A_MWSLrTf99_0),.clk(gclk));
	jdff dff_A_9qqlxDDT8_0(.dout(w_dff_A_LCOpbfAy6_0),.din(w_dff_A_9qqlxDDT8_0),.clk(gclk));
	jdff dff_A_LCOpbfAy6_0(.dout(w_dff_A_izv6SuXY7_0),.din(w_dff_A_LCOpbfAy6_0),.clk(gclk));
	jdff dff_A_izv6SuXY7_0(.dout(w_dff_A_7KmsnVih6_0),.din(w_dff_A_izv6SuXY7_0),.clk(gclk));
	jdff dff_A_7KmsnVih6_0(.dout(w_dff_A_bvKln7vL9_0),.din(w_dff_A_7KmsnVih6_0),.clk(gclk));
	jdff dff_A_bvKln7vL9_0(.dout(w_dff_A_RphIj3Cg1_0),.din(w_dff_A_bvKln7vL9_0),.clk(gclk));
	jdff dff_A_RphIj3Cg1_0(.dout(w_dff_A_gsdpr9LF7_0),.din(w_dff_A_RphIj3Cg1_0),.clk(gclk));
	jdff dff_A_gsdpr9LF7_0(.dout(G998),.din(w_dff_A_gsdpr9LF7_0),.clk(gclk));
	jdff dff_A_yoQ7gBu71_1(.dout(w_dff_A_iSYEqmS21_0),.din(w_dff_A_yoQ7gBu71_1),.clk(gclk));
	jdff dff_A_iSYEqmS21_0(.dout(w_dff_A_uNS3x3oT3_0),.din(w_dff_A_iSYEqmS21_0),.clk(gclk));
	jdff dff_A_uNS3x3oT3_0(.dout(w_dff_A_Lx3rdpWJ6_0),.din(w_dff_A_uNS3x3oT3_0),.clk(gclk));
	jdff dff_A_Lx3rdpWJ6_0(.dout(w_dff_A_vZ4IEJ8v7_0),.din(w_dff_A_Lx3rdpWJ6_0),.clk(gclk));
	jdff dff_A_vZ4IEJ8v7_0(.dout(w_dff_A_hEIGV5SA4_0),.din(w_dff_A_vZ4IEJ8v7_0),.clk(gclk));
	jdff dff_A_hEIGV5SA4_0(.dout(w_dff_A_weId0Al02_0),.din(w_dff_A_hEIGV5SA4_0),.clk(gclk));
	jdff dff_A_weId0Al02_0(.dout(w_dff_A_D9x0JpWX4_0),.din(w_dff_A_weId0Al02_0),.clk(gclk));
	jdff dff_A_D9x0JpWX4_0(.dout(w_dff_A_S0O6gJBc6_0),.din(w_dff_A_D9x0JpWX4_0),.clk(gclk));
	jdff dff_A_S0O6gJBc6_0(.dout(w_dff_A_YAUmi3wI3_0),.din(w_dff_A_S0O6gJBc6_0),.clk(gclk));
	jdff dff_A_YAUmi3wI3_0(.dout(w_dff_A_HEe99Rb48_0),.din(w_dff_A_YAUmi3wI3_0),.clk(gclk));
	jdff dff_A_HEe99Rb48_0(.dout(w_dff_A_7YMUW1C25_0),.din(w_dff_A_HEe99Rb48_0),.clk(gclk));
	jdff dff_A_7YMUW1C25_0(.dout(w_dff_A_xZWHCZ1w7_0),.din(w_dff_A_7YMUW1C25_0),.clk(gclk));
	jdff dff_A_xZWHCZ1w7_0(.dout(w_dff_A_S2M7FuCm3_0),.din(w_dff_A_xZWHCZ1w7_0),.clk(gclk));
	jdff dff_A_S2M7FuCm3_0(.dout(w_dff_A_zfigGTY95_0),.din(w_dff_A_S2M7FuCm3_0),.clk(gclk));
	jdff dff_A_zfigGTY95_0(.dout(w_dff_A_xE6rwWB77_0),.din(w_dff_A_zfigGTY95_0),.clk(gclk));
	jdff dff_A_xE6rwWB77_0(.dout(w_dff_A_DyG2AYCJ2_0),.din(w_dff_A_xE6rwWB77_0),.clk(gclk));
	jdff dff_A_DyG2AYCJ2_0(.dout(w_dff_A_KYIcgXZK9_0),.din(w_dff_A_DyG2AYCJ2_0),.clk(gclk));
	jdff dff_A_KYIcgXZK9_0(.dout(w_dff_A_DE0qVNGK7_0),.din(w_dff_A_KYIcgXZK9_0),.clk(gclk));
	jdff dff_A_DE0qVNGK7_0(.dout(G1000),.din(w_dff_A_DE0qVNGK7_0),.clk(gclk));
	jdff dff_A_BkWFxhEB2_2(.dout(w_dff_A_LIHDGeJw9_0),.din(w_dff_A_BkWFxhEB2_2),.clk(gclk));
	jdff dff_A_LIHDGeJw9_0(.dout(w_dff_A_Q2z2mpl82_0),.din(w_dff_A_LIHDGeJw9_0),.clk(gclk));
	jdff dff_A_Q2z2mpl82_0(.dout(w_dff_A_FK5KjLBy5_0),.din(w_dff_A_Q2z2mpl82_0),.clk(gclk));
	jdff dff_A_FK5KjLBy5_0(.dout(w_dff_A_nus5Dde81_0),.din(w_dff_A_FK5KjLBy5_0),.clk(gclk));
	jdff dff_A_nus5Dde81_0(.dout(G575),.din(w_dff_A_nus5Dde81_0),.clk(gclk));
	jdff dff_A_XLGJ52ZR5_2(.dout(w_dff_A_yO4CAvnu2_0),.din(w_dff_A_XLGJ52ZR5_2),.clk(gclk));
	jdff dff_A_yO4CAvnu2_0(.dout(w_dff_A_pxA9yVPv5_0),.din(w_dff_A_yO4CAvnu2_0),.clk(gclk));
	jdff dff_A_pxA9yVPv5_0(.dout(w_dff_A_dLK0pC1x3_0),.din(w_dff_A_pxA9yVPv5_0),.clk(gclk));
	jdff dff_A_dLK0pC1x3_0(.dout(w_dff_A_o0Jw7GZ85_0),.din(w_dff_A_dLK0pC1x3_0),.clk(gclk));
	jdff dff_A_o0Jw7GZ85_0(.dout(w_dff_A_IGgCN6zc6_0),.din(w_dff_A_o0Jw7GZ85_0),.clk(gclk));
	jdff dff_A_IGgCN6zc6_0(.dout(w_dff_A_tYqxSV9P9_0),.din(w_dff_A_IGgCN6zc6_0),.clk(gclk));
	jdff dff_A_tYqxSV9P9_0(.dout(w_dff_A_Gm6tIDHY6_0),.din(w_dff_A_tYqxSV9P9_0),.clk(gclk));
	jdff dff_A_Gm6tIDHY6_0(.dout(G585),.din(w_dff_A_Gm6tIDHY6_0),.clk(gclk));
	jdff dff_A_e2padhDy3_2(.dout(w_dff_A_uBXnkbt63_0),.din(w_dff_A_e2padhDy3_2),.clk(gclk));
	jdff dff_A_uBXnkbt63_0(.dout(w_dff_A_eEPrYxCc7_0),.din(w_dff_A_uBXnkbt63_0),.clk(gclk));
	jdff dff_A_eEPrYxCc7_0(.dout(w_dff_A_FD3nYQMz1_0),.din(w_dff_A_eEPrYxCc7_0),.clk(gclk));
	jdff dff_A_FD3nYQMz1_0(.dout(w_dff_A_KoTCeSlk2_0),.din(w_dff_A_FD3nYQMz1_0),.clk(gclk));
	jdff dff_A_KoTCeSlk2_0(.dout(w_dff_A_QonrsW5u4_0),.din(w_dff_A_KoTCeSlk2_0),.clk(gclk));
	jdff dff_A_QonrsW5u4_0(.dout(w_dff_A_5T2T07X71_0),.din(w_dff_A_QonrsW5u4_0),.clk(gclk));
	jdff dff_A_5T2T07X71_0(.dout(w_dff_A_I7e5AaJw5_0),.din(w_dff_A_5T2T07X71_0),.clk(gclk));
	jdff dff_A_I7e5AaJw5_0(.dout(w_dff_A_qZnUxT0U4_0),.din(w_dff_A_I7e5AaJw5_0),.clk(gclk));
	jdff dff_A_qZnUxT0U4_0(.dout(w_dff_A_FpbqjnAy5_0),.din(w_dff_A_qZnUxT0U4_0),.clk(gclk));
	jdff dff_A_FpbqjnAy5_0(.dout(w_dff_A_feb7IkaZ7_0),.din(w_dff_A_FpbqjnAy5_0),.clk(gclk));
	jdff dff_A_feb7IkaZ7_0(.dout(w_dff_A_OxP4DydG3_0),.din(w_dff_A_feb7IkaZ7_0),.clk(gclk));
	jdff dff_A_OxP4DydG3_0(.dout(w_dff_A_F5nQuhG97_0),.din(w_dff_A_OxP4DydG3_0),.clk(gclk));
	jdff dff_A_F5nQuhG97_0(.dout(w_dff_A_cJoOyBTr8_0),.din(w_dff_A_F5nQuhG97_0),.clk(gclk));
	jdff dff_A_cJoOyBTr8_0(.dout(G661),.din(w_dff_A_cJoOyBTr8_0),.clk(gclk));
	jdff dff_A_G2chA7m48_2(.dout(w_dff_A_wVK0n5eK1_0),.din(w_dff_A_G2chA7m48_2),.clk(gclk));
	jdff dff_A_wVK0n5eK1_0(.dout(w_dff_A_W2JuKv913_0),.din(w_dff_A_wVK0n5eK1_0),.clk(gclk));
	jdff dff_A_W2JuKv913_0(.dout(w_dff_A_xoMZBcXG3_0),.din(w_dff_A_W2JuKv913_0),.clk(gclk));
	jdff dff_A_xoMZBcXG3_0(.dout(w_dff_A_JwSLsdri0_0),.din(w_dff_A_xoMZBcXG3_0),.clk(gclk));
	jdff dff_A_JwSLsdri0_0(.dout(w_dff_A_nSVnXpew0_0),.din(w_dff_A_JwSLsdri0_0),.clk(gclk));
	jdff dff_A_nSVnXpew0_0(.dout(w_dff_A_W6ZacWyL9_0),.din(w_dff_A_nSVnXpew0_0),.clk(gclk));
	jdff dff_A_W6ZacWyL9_0(.dout(w_dff_A_rYbRjz7Y4_0),.din(w_dff_A_W6ZacWyL9_0),.clk(gclk));
	jdff dff_A_rYbRjz7Y4_0(.dout(w_dff_A_Pf22BUOx2_0),.din(w_dff_A_rYbRjz7Y4_0),.clk(gclk));
	jdff dff_A_Pf22BUOx2_0(.dout(w_dff_A_aScrGtdP7_0),.din(w_dff_A_Pf22BUOx2_0),.clk(gclk));
	jdff dff_A_aScrGtdP7_0(.dout(w_dff_A_DjvQs8ro6_0),.din(w_dff_A_aScrGtdP7_0),.clk(gclk));
	jdff dff_A_DjvQs8ro6_0(.dout(w_dff_A_YNj8iHuq2_0),.din(w_dff_A_DjvQs8ro6_0),.clk(gclk));
	jdff dff_A_YNj8iHuq2_0(.dout(w_dff_A_IeYx8ogJ0_0),.din(w_dff_A_YNj8iHuq2_0),.clk(gclk));
	jdff dff_A_IeYx8ogJ0_0(.dout(w_dff_A_P0pqoz6w3_0),.din(w_dff_A_IeYx8ogJ0_0),.clk(gclk));
	jdff dff_A_P0pqoz6w3_0(.dout(G693),.din(w_dff_A_P0pqoz6w3_0),.clk(gclk));
	jdff dff_A_KfeUhVrq5_2(.dout(w_dff_A_sw9TurKs6_0),.din(w_dff_A_KfeUhVrq5_2),.clk(gclk));
	jdff dff_A_sw9TurKs6_0(.dout(w_dff_A_gdKEuIgu0_0),.din(w_dff_A_sw9TurKs6_0),.clk(gclk));
	jdff dff_A_gdKEuIgu0_0(.dout(w_dff_A_6TAhwbi33_0),.din(w_dff_A_gdKEuIgu0_0),.clk(gclk));
	jdff dff_A_6TAhwbi33_0(.dout(w_dff_A_f8wdPuSn7_0),.din(w_dff_A_6TAhwbi33_0),.clk(gclk));
	jdff dff_A_f8wdPuSn7_0(.dout(w_dff_A_PPEJbsS00_0),.din(w_dff_A_f8wdPuSn7_0),.clk(gclk));
	jdff dff_A_PPEJbsS00_0(.dout(w_dff_A_VcBBHN7L5_0),.din(w_dff_A_PPEJbsS00_0),.clk(gclk));
	jdff dff_A_VcBBHN7L5_0(.dout(G747),.din(w_dff_A_VcBBHN7L5_0),.clk(gclk));
	jdff dff_A_PcgqmF0C8_2(.dout(w_dff_A_LlYxkoFK2_0),.din(w_dff_A_PcgqmF0C8_2),.clk(gclk));
	jdff dff_A_LlYxkoFK2_0(.dout(w_dff_A_PrxaREaY1_0),.din(w_dff_A_LlYxkoFK2_0),.clk(gclk));
	jdff dff_A_PrxaREaY1_0(.dout(w_dff_A_WrM61pGw6_0),.din(w_dff_A_PrxaREaY1_0),.clk(gclk));
	jdff dff_A_WrM61pGw6_0(.dout(w_dff_A_6Agh3nae8_0),.din(w_dff_A_WrM61pGw6_0),.clk(gclk));
	jdff dff_A_6Agh3nae8_0(.dout(w_dff_A_ZDzdhXwH2_0),.din(w_dff_A_6Agh3nae8_0),.clk(gclk));
	jdff dff_A_ZDzdhXwH2_0(.dout(w_dff_A_ubzKpfvl7_0),.din(w_dff_A_ZDzdhXwH2_0),.clk(gclk));
	jdff dff_A_ubzKpfvl7_0(.dout(w_dff_A_IoZq34576_0),.din(w_dff_A_ubzKpfvl7_0),.clk(gclk));
	jdff dff_A_IoZq34576_0(.dout(w_dff_A_zt1aQIae0_0),.din(w_dff_A_IoZq34576_0),.clk(gclk));
	jdff dff_A_zt1aQIae0_0(.dout(G752),.din(w_dff_A_zt1aQIae0_0),.clk(gclk));
	jdff dff_A_m0ajpebn0_2(.dout(w_dff_A_H21ayT7A1_0),.din(w_dff_A_m0ajpebn0_2),.clk(gclk));
	jdff dff_A_H21ayT7A1_0(.dout(w_dff_A_9qftIk2h8_0),.din(w_dff_A_H21ayT7A1_0),.clk(gclk));
	jdff dff_A_9qftIk2h8_0(.dout(w_dff_A_CEZNUDmR0_0),.din(w_dff_A_9qftIk2h8_0),.clk(gclk));
	jdff dff_A_CEZNUDmR0_0(.dout(w_dff_A_LF3C5FvE0_0),.din(w_dff_A_CEZNUDmR0_0),.clk(gclk));
	jdff dff_A_LF3C5FvE0_0(.dout(w_dff_A_O2C8IRlZ2_0),.din(w_dff_A_LF3C5FvE0_0),.clk(gclk));
	jdff dff_A_O2C8IRlZ2_0(.dout(w_dff_A_MtlKiWrl1_0),.din(w_dff_A_O2C8IRlZ2_0),.clk(gclk));
	jdff dff_A_MtlKiWrl1_0(.dout(w_dff_A_Rnp7sFGs3_0),.din(w_dff_A_MtlKiWrl1_0),.clk(gclk));
	jdff dff_A_Rnp7sFGs3_0(.dout(w_dff_A_hv5YRrBr0_0),.din(w_dff_A_Rnp7sFGs3_0),.clk(gclk));
	jdff dff_A_hv5YRrBr0_0(.dout(w_dff_A_79skVkXk9_0),.din(w_dff_A_hv5YRrBr0_0),.clk(gclk));
	jdff dff_A_79skVkXk9_0(.dout(G757),.din(w_dff_A_79skVkXk9_0),.clk(gclk));
	jdff dff_A_XI6uvqqZ6_2(.dout(w_dff_A_3m7y0daf0_0),.din(w_dff_A_XI6uvqqZ6_2),.clk(gclk));
	jdff dff_A_3m7y0daf0_0(.dout(w_dff_A_cfPFmr3Q8_0),.din(w_dff_A_3m7y0daf0_0),.clk(gclk));
	jdff dff_A_cfPFmr3Q8_0(.dout(w_dff_A_AT7wuAsi5_0),.din(w_dff_A_cfPFmr3Q8_0),.clk(gclk));
	jdff dff_A_AT7wuAsi5_0(.dout(w_dff_A_d0gbtnvA0_0),.din(w_dff_A_AT7wuAsi5_0),.clk(gclk));
	jdff dff_A_d0gbtnvA0_0(.dout(w_dff_A_o4BH9woU7_0),.din(w_dff_A_d0gbtnvA0_0),.clk(gclk));
	jdff dff_A_o4BH9woU7_0(.dout(w_dff_A_IyjwKG330_0),.din(w_dff_A_o4BH9woU7_0),.clk(gclk));
	jdff dff_A_IyjwKG330_0(.dout(w_dff_A_4rkMP9574_0),.din(w_dff_A_IyjwKG330_0),.clk(gclk));
	jdff dff_A_4rkMP9574_0(.dout(w_dff_A_CGycL2bp0_0),.din(w_dff_A_4rkMP9574_0),.clk(gclk));
	jdff dff_A_CGycL2bp0_0(.dout(w_dff_A_Ekrj35rS5_0),.din(w_dff_A_CGycL2bp0_0),.clk(gclk));
	jdff dff_A_Ekrj35rS5_0(.dout(w_dff_A_YdVTRq8h2_0),.din(w_dff_A_Ekrj35rS5_0),.clk(gclk));
	jdff dff_A_YdVTRq8h2_0(.dout(G762),.din(w_dff_A_YdVTRq8h2_0),.clk(gclk));
	jdff dff_A_DLFcmILU9_2(.dout(w_dff_A_7DsRj9d82_0),.din(w_dff_A_DLFcmILU9_2),.clk(gclk));
	jdff dff_A_7DsRj9d82_0(.dout(w_dff_A_IZWbhzad0_0),.din(w_dff_A_7DsRj9d82_0),.clk(gclk));
	jdff dff_A_IZWbhzad0_0(.dout(w_dff_A_07IHCwMa5_0),.din(w_dff_A_IZWbhzad0_0),.clk(gclk));
	jdff dff_A_07IHCwMa5_0(.dout(w_dff_A_j941N7RO1_0),.din(w_dff_A_07IHCwMa5_0),.clk(gclk));
	jdff dff_A_j941N7RO1_0(.dout(w_dff_A_CQJAyi6Z7_0),.din(w_dff_A_j941N7RO1_0),.clk(gclk));
	jdff dff_A_CQJAyi6Z7_0(.dout(w_dff_A_TuKixy3M7_0),.din(w_dff_A_CQJAyi6Z7_0),.clk(gclk));
	jdff dff_A_TuKixy3M7_0(.dout(G787),.din(w_dff_A_TuKixy3M7_0),.clk(gclk));
	jdff dff_A_YktHXzVq0_2(.dout(w_dff_A_re5PmL8l6_0),.din(w_dff_A_YktHXzVq0_2),.clk(gclk));
	jdff dff_A_re5PmL8l6_0(.dout(w_dff_A_AmdGjX9a3_0),.din(w_dff_A_re5PmL8l6_0),.clk(gclk));
	jdff dff_A_AmdGjX9a3_0(.dout(w_dff_A_L8VBNfcp8_0),.din(w_dff_A_AmdGjX9a3_0),.clk(gclk));
	jdff dff_A_L8VBNfcp8_0(.dout(w_dff_A_R4aHEPUq6_0),.din(w_dff_A_L8VBNfcp8_0),.clk(gclk));
	jdff dff_A_R4aHEPUq6_0(.dout(w_dff_A_7uUWhyxP3_0),.din(w_dff_A_R4aHEPUq6_0),.clk(gclk));
	jdff dff_A_7uUWhyxP3_0(.dout(w_dff_A_IfoUIBxR7_0),.din(w_dff_A_7uUWhyxP3_0),.clk(gclk));
	jdff dff_A_IfoUIBxR7_0(.dout(w_dff_A_CmysDfHQ4_0),.din(w_dff_A_IfoUIBxR7_0),.clk(gclk));
	jdff dff_A_CmysDfHQ4_0(.dout(w_dff_A_QLxuj4PK5_0),.din(w_dff_A_CmysDfHQ4_0),.clk(gclk));
	jdff dff_A_QLxuj4PK5_0(.dout(G792),.din(w_dff_A_QLxuj4PK5_0),.clk(gclk));
	jdff dff_A_cyMtHO7V5_2(.dout(w_dff_A_sUutweHT1_0),.din(w_dff_A_cyMtHO7V5_2),.clk(gclk));
	jdff dff_A_sUutweHT1_0(.dout(w_dff_A_fBhiAi4m1_0),.din(w_dff_A_sUutweHT1_0),.clk(gclk));
	jdff dff_A_fBhiAi4m1_0(.dout(w_dff_A_yovYQJGz1_0),.din(w_dff_A_fBhiAi4m1_0),.clk(gclk));
	jdff dff_A_yovYQJGz1_0(.dout(w_dff_A_nw5VLl9K3_0),.din(w_dff_A_yovYQJGz1_0),.clk(gclk));
	jdff dff_A_nw5VLl9K3_0(.dout(w_dff_A_Nj7wgGHs1_0),.din(w_dff_A_nw5VLl9K3_0),.clk(gclk));
	jdff dff_A_Nj7wgGHs1_0(.dout(w_dff_A_JdRDKO1R0_0),.din(w_dff_A_Nj7wgGHs1_0),.clk(gclk));
	jdff dff_A_JdRDKO1R0_0(.dout(w_dff_A_N7F4nlJd9_0),.din(w_dff_A_JdRDKO1R0_0),.clk(gclk));
	jdff dff_A_N7F4nlJd9_0(.dout(w_dff_A_gforHNgk5_0),.din(w_dff_A_N7F4nlJd9_0),.clk(gclk));
	jdff dff_A_gforHNgk5_0(.dout(w_dff_A_TqNE87JS0_0),.din(w_dff_A_gforHNgk5_0),.clk(gclk));
	jdff dff_A_TqNE87JS0_0(.dout(G797),.din(w_dff_A_TqNE87JS0_0),.clk(gclk));
	jdff dff_A_UsxZO5xA4_2(.dout(w_dff_A_G4UTTrst8_0),.din(w_dff_A_UsxZO5xA4_2),.clk(gclk));
	jdff dff_A_G4UTTrst8_0(.dout(w_dff_A_1npkqYoq4_0),.din(w_dff_A_G4UTTrst8_0),.clk(gclk));
	jdff dff_A_1npkqYoq4_0(.dout(w_dff_A_ycIUmILo3_0),.din(w_dff_A_1npkqYoq4_0),.clk(gclk));
	jdff dff_A_ycIUmILo3_0(.dout(w_dff_A_RmDXIECh4_0),.din(w_dff_A_ycIUmILo3_0),.clk(gclk));
	jdff dff_A_RmDXIECh4_0(.dout(w_dff_A_z1RsAgon6_0),.din(w_dff_A_RmDXIECh4_0),.clk(gclk));
	jdff dff_A_z1RsAgon6_0(.dout(w_dff_A_10lPO5b46_0),.din(w_dff_A_z1RsAgon6_0),.clk(gclk));
	jdff dff_A_10lPO5b46_0(.dout(w_dff_A_2WgqWnaS6_0),.din(w_dff_A_10lPO5b46_0),.clk(gclk));
	jdff dff_A_2WgqWnaS6_0(.dout(w_dff_A_E6rFXZc67_0),.din(w_dff_A_2WgqWnaS6_0),.clk(gclk));
	jdff dff_A_E6rFXZc67_0(.dout(w_dff_A_SCaJMEFS6_0),.din(w_dff_A_E6rFXZc67_0),.clk(gclk));
	jdff dff_A_SCaJMEFS6_0(.dout(w_dff_A_R4zKaMHj4_0),.din(w_dff_A_SCaJMEFS6_0),.clk(gclk));
	jdff dff_A_R4zKaMHj4_0(.dout(G802),.din(w_dff_A_R4zKaMHj4_0),.clk(gclk));
	jdff dff_A_6jd38nub0_2(.dout(w_dff_A_HUUyLBEI8_0),.din(w_dff_A_6jd38nub0_2),.clk(gclk));
	jdff dff_A_HUUyLBEI8_0(.dout(w_dff_A_NJWHBOQZ2_0),.din(w_dff_A_HUUyLBEI8_0),.clk(gclk));
	jdff dff_A_NJWHBOQZ2_0(.dout(w_dff_A_8bF9mKUP4_0),.din(w_dff_A_NJWHBOQZ2_0),.clk(gclk));
	jdff dff_A_8bF9mKUP4_0(.dout(w_dff_A_IkevpuYe7_0),.din(w_dff_A_8bF9mKUP4_0),.clk(gclk));
	jdff dff_A_IkevpuYe7_0(.dout(w_dff_A_33ApNxvO6_0),.din(w_dff_A_IkevpuYe7_0),.clk(gclk));
	jdff dff_A_33ApNxvO6_0(.dout(G642),.din(w_dff_A_33ApNxvO6_0),.clk(gclk));
	jdff dff_A_OpM8B9au0_2(.dout(w_dff_A_aI0b3nHX3_0),.din(w_dff_A_OpM8B9au0_2),.clk(gclk));
	jdff dff_A_aI0b3nHX3_0(.dout(w_dff_A_eOUS4aCB5_0),.din(w_dff_A_aI0b3nHX3_0),.clk(gclk));
	jdff dff_A_eOUS4aCB5_0(.dout(w_dff_A_Movwvcct3_0),.din(w_dff_A_eOUS4aCB5_0),.clk(gclk));
	jdff dff_A_Movwvcct3_0(.dout(w_dff_A_WU3jNiUi5_0),.din(w_dff_A_Movwvcct3_0),.clk(gclk));
	jdff dff_A_WU3jNiUi5_0(.dout(w_dff_A_QBGXEpzD3_0),.din(w_dff_A_WU3jNiUi5_0),.clk(gclk));
	jdff dff_A_QBGXEpzD3_0(.dout(w_dff_A_g0GIViA89_0),.din(w_dff_A_QBGXEpzD3_0),.clk(gclk));
	jdff dff_A_g0GIViA89_0(.dout(w_dff_A_amorDON28_0),.din(w_dff_A_g0GIViA89_0),.clk(gclk));
	jdff dff_A_amorDON28_0(.dout(w_dff_A_TezhaO5U8_0),.din(w_dff_A_amorDON28_0),.clk(gclk));
	jdff dff_A_TezhaO5U8_0(.dout(w_dff_A_bMCyt9rB7_0),.din(w_dff_A_TezhaO5U8_0),.clk(gclk));
	jdff dff_A_bMCyt9rB7_0(.dout(G664),.din(w_dff_A_bMCyt9rB7_0),.clk(gclk));
	jdff dff_A_udMizoxK1_2(.dout(w_dff_A_yBkPGO3U5_0),.din(w_dff_A_udMizoxK1_2),.clk(gclk));
	jdff dff_A_yBkPGO3U5_0(.dout(w_dff_A_wEysfK7J6_0),.din(w_dff_A_yBkPGO3U5_0),.clk(gclk));
	jdff dff_A_wEysfK7J6_0(.dout(w_dff_A_zETBLhsg2_0),.din(w_dff_A_wEysfK7J6_0),.clk(gclk));
	jdff dff_A_zETBLhsg2_0(.dout(w_dff_A_3V4LSvAs7_0),.din(w_dff_A_zETBLhsg2_0),.clk(gclk));
	jdff dff_A_3V4LSvAs7_0(.dout(w_dff_A_xMKSsKJY5_0),.din(w_dff_A_3V4LSvAs7_0),.clk(gclk));
	jdff dff_A_xMKSsKJY5_0(.dout(w_dff_A_vzrUmWJS2_0),.din(w_dff_A_xMKSsKJY5_0),.clk(gclk));
	jdff dff_A_vzrUmWJS2_0(.dout(w_dff_A_92m1C4v31_0),.din(w_dff_A_vzrUmWJS2_0),.clk(gclk));
	jdff dff_A_92m1C4v31_0(.dout(w_dff_A_fy4KqLWz1_0),.din(w_dff_A_92m1C4v31_0),.clk(gclk));
	jdff dff_A_fy4KqLWz1_0(.dout(G667),.din(w_dff_A_fy4KqLWz1_0),.clk(gclk));
	jdff dff_A_TCP58EKm3_2(.dout(w_dff_A_iqqhNhl31_0),.din(w_dff_A_TCP58EKm3_2),.clk(gclk));
	jdff dff_A_iqqhNhl31_0(.dout(w_dff_A_9P5V4bFX5_0),.din(w_dff_A_iqqhNhl31_0),.clk(gclk));
	jdff dff_A_9P5V4bFX5_0(.dout(w_dff_A_DRJfTUuy4_0),.din(w_dff_A_9P5V4bFX5_0),.clk(gclk));
	jdff dff_A_DRJfTUuy4_0(.dout(w_dff_A_LQhoXsez3_0),.din(w_dff_A_DRJfTUuy4_0),.clk(gclk));
	jdff dff_A_LQhoXsez3_0(.dout(w_dff_A_27r3yQnt9_0),.din(w_dff_A_LQhoXsez3_0),.clk(gclk));
	jdff dff_A_27r3yQnt9_0(.dout(w_dff_A_jm2Pknel3_0),.din(w_dff_A_27r3yQnt9_0),.clk(gclk));
	jdff dff_A_jm2Pknel3_0(.dout(w_dff_A_aNCUmeGx3_0),.din(w_dff_A_jm2Pknel3_0),.clk(gclk));
	jdff dff_A_aNCUmeGx3_0(.dout(G670),.din(w_dff_A_aNCUmeGx3_0),.clk(gclk));
	jdff dff_A_QvBFmF6Z6_2(.dout(w_dff_A_0fdGEpoZ3_0),.din(w_dff_A_QvBFmF6Z6_2),.clk(gclk));
	jdff dff_A_0fdGEpoZ3_0(.dout(w_dff_A_O3kUIhD13_0),.din(w_dff_A_0fdGEpoZ3_0),.clk(gclk));
	jdff dff_A_O3kUIhD13_0(.dout(w_dff_A_YqtBKm4R3_0),.din(w_dff_A_O3kUIhD13_0),.clk(gclk));
	jdff dff_A_YqtBKm4R3_0(.dout(w_dff_A_nowEBGt29_0),.din(w_dff_A_YqtBKm4R3_0),.clk(gclk));
	jdff dff_A_nowEBGt29_0(.dout(w_dff_A_paLQIGTv9_0),.din(w_dff_A_nowEBGt29_0),.clk(gclk));
	jdff dff_A_paLQIGTv9_0(.dout(G676),.din(w_dff_A_paLQIGTv9_0),.clk(gclk));
	jdff dff_A_njPQMHMP1_2(.dout(w_dff_A_8caSmFim4_0),.din(w_dff_A_njPQMHMP1_2),.clk(gclk));
	jdff dff_A_8caSmFim4_0(.dout(w_dff_A_ZIDX8myp7_0),.din(w_dff_A_8caSmFim4_0),.clk(gclk));
	jdff dff_A_ZIDX8myp7_0(.dout(w_dff_A_yt2ugcf46_0),.din(w_dff_A_ZIDX8myp7_0),.clk(gclk));
	jdff dff_A_yt2ugcf46_0(.dout(w_dff_A_1hHPdofn0_0),.din(w_dff_A_yt2ugcf46_0),.clk(gclk));
	jdff dff_A_1hHPdofn0_0(.dout(w_dff_A_ABEYC4pv5_0),.din(w_dff_A_1hHPdofn0_0),.clk(gclk));
	jdff dff_A_ABEYC4pv5_0(.dout(w_dff_A_HfBsieBw1_0),.din(w_dff_A_ABEYC4pv5_0),.clk(gclk));
	jdff dff_A_HfBsieBw1_0(.dout(w_dff_A_MeHZ2idK8_0),.din(w_dff_A_HfBsieBw1_0),.clk(gclk));
	jdff dff_A_MeHZ2idK8_0(.dout(w_dff_A_BucchbI89_0),.din(w_dff_A_MeHZ2idK8_0),.clk(gclk));
	jdff dff_A_BucchbI89_0(.dout(w_dff_A_Mrg8eEnt9_0),.din(w_dff_A_BucchbI89_0),.clk(gclk));
	jdff dff_A_Mrg8eEnt9_0(.dout(G696),.din(w_dff_A_Mrg8eEnt9_0),.clk(gclk));
	jdff dff_A_ZS1XpX9r3_2(.dout(w_dff_A_zdlHojwO9_0),.din(w_dff_A_ZS1XpX9r3_2),.clk(gclk));
	jdff dff_A_zdlHojwO9_0(.dout(w_dff_A_rXAFWKTq6_0),.din(w_dff_A_zdlHojwO9_0),.clk(gclk));
	jdff dff_A_rXAFWKTq6_0(.dout(w_dff_A_NaHH3ghF9_0),.din(w_dff_A_rXAFWKTq6_0),.clk(gclk));
	jdff dff_A_NaHH3ghF9_0(.dout(w_dff_A_HGPSY1TS8_0),.din(w_dff_A_NaHH3ghF9_0),.clk(gclk));
	jdff dff_A_HGPSY1TS8_0(.dout(w_dff_A_sZZ8GS4z4_0),.din(w_dff_A_HGPSY1TS8_0),.clk(gclk));
	jdff dff_A_sZZ8GS4z4_0(.dout(w_dff_A_0TPxsssF6_0),.din(w_dff_A_sZZ8GS4z4_0),.clk(gclk));
	jdff dff_A_0TPxsssF6_0(.dout(w_dff_A_yox6R9RO2_0),.din(w_dff_A_0TPxsssF6_0),.clk(gclk));
	jdff dff_A_yox6R9RO2_0(.dout(w_dff_A_DSeg5Ow66_0),.din(w_dff_A_yox6R9RO2_0),.clk(gclk));
	jdff dff_A_DSeg5Ow66_0(.dout(G699),.din(w_dff_A_DSeg5Ow66_0),.clk(gclk));
	jdff dff_A_zWSShnYZ7_2(.dout(w_dff_A_wKc1AnBc5_0),.din(w_dff_A_zWSShnYZ7_2),.clk(gclk));
	jdff dff_A_wKc1AnBc5_0(.dout(w_dff_A_psyDHTXp7_0),.din(w_dff_A_wKc1AnBc5_0),.clk(gclk));
	jdff dff_A_psyDHTXp7_0(.dout(w_dff_A_NBLqhgg33_0),.din(w_dff_A_psyDHTXp7_0),.clk(gclk));
	jdff dff_A_NBLqhgg33_0(.dout(w_dff_A_go4tHWlx0_0),.din(w_dff_A_NBLqhgg33_0),.clk(gclk));
	jdff dff_A_go4tHWlx0_0(.dout(w_dff_A_c9CRuBSl9_0),.din(w_dff_A_go4tHWlx0_0),.clk(gclk));
	jdff dff_A_c9CRuBSl9_0(.dout(w_dff_A_Gjjnfko22_0),.din(w_dff_A_c9CRuBSl9_0),.clk(gclk));
	jdff dff_A_Gjjnfko22_0(.dout(w_dff_A_86oNSgpI9_0),.din(w_dff_A_Gjjnfko22_0),.clk(gclk));
	jdff dff_A_86oNSgpI9_0(.dout(G702),.din(w_dff_A_86oNSgpI9_0),.clk(gclk));
	jdff dff_A_l4yz9gMX7_2(.dout(w_dff_A_zkYGFyXL7_0),.din(w_dff_A_l4yz9gMX7_2),.clk(gclk));
	jdff dff_A_zkYGFyXL7_0(.dout(w_dff_A_VRRIksgD8_0),.din(w_dff_A_zkYGFyXL7_0),.clk(gclk));
	jdff dff_A_VRRIksgD8_0(.dout(w_dff_A_r3tqBjKz0_0),.din(w_dff_A_VRRIksgD8_0),.clk(gclk));
	jdff dff_A_r3tqBjKz0_0(.dout(w_dff_A_OY81yL1H5_0),.din(w_dff_A_r3tqBjKz0_0),.clk(gclk));
	jdff dff_A_OY81yL1H5_0(.dout(G818),.din(w_dff_A_OY81yL1H5_0),.clk(gclk));
	jdff dff_A_L9zsaGmQ8_2(.dout(w_dff_A_LYpe9dVu2_0),.din(w_dff_A_L9zsaGmQ8_2),.clk(gclk));
	jdff dff_A_LYpe9dVu2_0(.dout(w_dff_A_fuy1ln707_0),.din(w_dff_A_LYpe9dVu2_0),.clk(gclk));
	jdff dff_A_fuy1ln707_0(.dout(w_dff_A_qIv0wFGT5_0),.din(w_dff_A_fuy1ln707_0),.clk(gclk));
	jdff dff_A_qIv0wFGT5_0(.dout(w_dff_A_THk1K6z39_0),.din(w_dff_A_qIv0wFGT5_0),.clk(gclk));
	jdff dff_A_THk1K6z39_0(.dout(w_dff_A_9YHmGWnu8_0),.din(w_dff_A_THk1K6z39_0),.clk(gclk));
	jdff dff_A_9YHmGWnu8_0(.dout(w_dff_A_k3ttNZWg1_0),.din(w_dff_A_9YHmGWnu8_0),.clk(gclk));
	jdff dff_A_k3ttNZWg1_0(.dout(w_dff_A_USZW6DS72_0),.din(w_dff_A_k3ttNZWg1_0),.clk(gclk));
	jdff dff_A_USZW6DS72_0(.dout(w_dff_A_JzIb8vCp1_0),.din(w_dff_A_USZW6DS72_0),.clk(gclk));
	jdff dff_A_JzIb8vCp1_0(.dout(G813),.din(w_dff_A_JzIb8vCp1_0),.clk(gclk));
	jdff dff_A_9EZjqA4L7_1(.dout(w_dff_A_bQrR0xJV0_0),.din(w_dff_A_9EZjqA4L7_1),.clk(gclk));
	jdff dff_A_bQrR0xJV0_0(.dout(w_dff_A_pCvGfdx16_0),.din(w_dff_A_bQrR0xJV0_0),.clk(gclk));
	jdff dff_A_pCvGfdx16_0(.dout(w_dff_A_YYRBnywg7_0),.din(w_dff_A_pCvGfdx16_0),.clk(gclk));
	jdff dff_A_YYRBnywg7_0(.dout(w_dff_A_wj5tLXI33_0),.din(w_dff_A_YYRBnywg7_0),.clk(gclk));
	jdff dff_A_wj5tLXI33_0(.dout(G824),.din(w_dff_A_wj5tLXI33_0),.clk(gclk));
	jdff dff_A_dwolBJTY9_1(.dout(w_dff_A_BKpGG5iG4_0),.din(w_dff_A_dwolBJTY9_1),.clk(gclk));
	jdff dff_A_BKpGG5iG4_0(.dout(w_dff_A_Hpep7J3y2_0),.din(w_dff_A_BKpGG5iG4_0),.clk(gclk));
	jdff dff_A_Hpep7J3y2_0(.dout(w_dff_A_JRdwbNRh2_0),.din(w_dff_A_Hpep7J3y2_0),.clk(gclk));
	jdff dff_A_JRdwbNRh2_0(.dout(w_dff_A_vjXltcIc1_0),.din(w_dff_A_JRdwbNRh2_0),.clk(gclk));
	jdff dff_A_vjXltcIc1_0(.dout(w_dff_A_AlalE32A0_0),.din(w_dff_A_vjXltcIc1_0),.clk(gclk));
	jdff dff_A_AlalE32A0_0(.dout(w_dff_A_m8FZdKM60_0),.din(w_dff_A_AlalE32A0_0),.clk(gclk));
	jdff dff_A_m8FZdKM60_0(.dout(w_dff_A_p1awfmKN1_0),.din(w_dff_A_m8FZdKM60_0),.clk(gclk));
	jdff dff_A_p1awfmKN1_0(.dout(G826),.din(w_dff_A_p1awfmKN1_0),.clk(gclk));
	jdff dff_A_3wJHFv7k4_1(.dout(w_dff_A_VkfNnmTx6_0),.din(w_dff_A_3wJHFv7k4_1),.clk(gclk));
	jdff dff_A_VkfNnmTx6_0(.dout(w_dff_A_3XnJbGon3_0),.din(w_dff_A_VkfNnmTx6_0),.clk(gclk));
	jdff dff_A_3XnJbGon3_0(.dout(w_dff_A_VIfu4nsG8_0),.din(w_dff_A_3XnJbGon3_0),.clk(gclk));
	jdff dff_A_VIfu4nsG8_0(.dout(w_dff_A_92RiWWjv9_0),.din(w_dff_A_VIfu4nsG8_0),.clk(gclk));
	jdff dff_A_92RiWWjv9_0(.dout(w_dff_A_IGMm0hw32_0),.din(w_dff_A_92RiWWjv9_0),.clk(gclk));
	jdff dff_A_IGMm0hw32_0(.dout(w_dff_A_M8CvIGpZ2_0),.din(w_dff_A_IGMm0hw32_0),.clk(gclk));
	jdff dff_A_M8CvIGpZ2_0(.dout(w_dff_A_6fxtla8y5_0),.din(w_dff_A_M8CvIGpZ2_0),.clk(gclk));
	jdff dff_A_6fxtla8y5_0(.dout(G828),.din(w_dff_A_6fxtla8y5_0),.clk(gclk));
	jdff dff_A_MBb3kScK9_1(.dout(w_dff_A_UGF4B9OL7_0),.din(w_dff_A_MBb3kScK9_1),.clk(gclk));
	jdff dff_A_UGF4B9OL7_0(.dout(w_dff_A_5cW82O3G2_0),.din(w_dff_A_UGF4B9OL7_0),.clk(gclk));
	jdff dff_A_5cW82O3G2_0(.dout(w_dff_A_2DXE5XMF0_0),.din(w_dff_A_5cW82O3G2_0),.clk(gclk));
	jdff dff_A_2DXE5XMF0_0(.dout(w_dff_A_zGdrRZ2t6_0),.din(w_dff_A_2DXE5XMF0_0),.clk(gclk));
	jdff dff_A_zGdrRZ2t6_0(.dout(w_dff_A_7kQy0GeY2_0),.din(w_dff_A_zGdrRZ2t6_0),.clk(gclk));
	jdff dff_A_7kQy0GeY2_0(.dout(w_dff_A_i08W0axm3_0),.din(w_dff_A_7kQy0GeY2_0),.clk(gclk));
	jdff dff_A_i08W0axm3_0(.dout(w_dff_A_EsSEP6TS5_0),.din(w_dff_A_i08W0axm3_0),.clk(gclk));
	jdff dff_A_EsSEP6TS5_0(.dout(w_dff_A_fmwDIW7V4_0),.din(w_dff_A_EsSEP6TS5_0),.clk(gclk));
	jdff dff_A_fmwDIW7V4_0(.dout(G830),.din(w_dff_A_fmwDIW7V4_0),.clk(gclk));
	jdff dff_A_nqVLCUVr3_2(.dout(w_dff_A_0VfPSdb12_0),.din(w_dff_A_nqVLCUVr3_2),.clk(gclk));
	jdff dff_A_0VfPSdb12_0(.dout(w_dff_A_Iagi2dte9_0),.din(w_dff_A_0VfPSdb12_0),.clk(gclk));
	jdff dff_A_Iagi2dte9_0(.dout(w_dff_A_FlMEXxlu2_0),.din(w_dff_A_Iagi2dte9_0),.clk(gclk));
	jdff dff_A_FlMEXxlu2_0(.dout(w_dff_A_sBiLunp72_0),.din(w_dff_A_FlMEXxlu2_0),.clk(gclk));
	jdff dff_A_sBiLunp72_0(.dout(w_dff_A_A0adeJyV5_0),.din(w_dff_A_sBiLunp72_0),.clk(gclk));
	jdff dff_A_A0adeJyV5_0(.dout(w_dff_A_Od26WcvR8_0),.din(w_dff_A_A0adeJyV5_0),.clk(gclk));
	jdff dff_A_Od26WcvR8_0(.dout(w_dff_A_na0vV0mC1_0),.din(w_dff_A_Od26WcvR8_0),.clk(gclk));
	jdff dff_A_na0vV0mC1_0(.dout(w_dff_A_cfghQrmU8_0),.din(w_dff_A_na0vV0mC1_0),.clk(gclk));
	jdff dff_A_cfghQrmU8_0(.dout(w_dff_A_lU2XKDt26_0),.din(w_dff_A_cfghQrmU8_0),.clk(gclk));
	jdff dff_A_lU2XKDt26_0(.dout(w_dff_A_p1ahxHWL0_0),.din(w_dff_A_lU2XKDt26_0),.clk(gclk));
	jdff dff_A_p1ahxHWL0_0(.dout(w_dff_A_xDQ8vvcq9_0),.din(w_dff_A_p1ahxHWL0_0),.clk(gclk));
	jdff dff_A_xDQ8vvcq9_0(.dout(w_dff_A_38UsTg3g7_0),.din(w_dff_A_xDQ8vvcq9_0),.clk(gclk));
	jdff dff_A_38UsTg3g7_0(.dout(w_dff_A_PV3dgX6G1_0),.din(w_dff_A_38UsTg3g7_0),.clk(gclk));
	jdff dff_A_PV3dgX6G1_0(.dout(w_dff_A_QFuOL9ih1_0),.din(w_dff_A_PV3dgX6G1_0),.clk(gclk));
	jdff dff_A_QFuOL9ih1_0(.dout(w_dff_A_aoOEAbmr5_0),.din(w_dff_A_QFuOL9ih1_0),.clk(gclk));
	jdff dff_A_aoOEAbmr5_0(.dout(G854),.din(w_dff_A_aoOEAbmr5_0),.clk(gclk));
	jdff dff_A_O5MACyFk6_1(.dout(w_dff_A_NZNHPMkf8_0),.din(w_dff_A_O5MACyFk6_1),.clk(gclk));
	jdff dff_A_NZNHPMkf8_0(.dout(w_dff_A_nrSWo5Hn7_0),.din(w_dff_A_NZNHPMkf8_0),.clk(gclk));
	jdff dff_A_nrSWo5Hn7_0(.dout(w_dff_A_5l5XOZcE6_0),.din(w_dff_A_nrSWo5Hn7_0),.clk(gclk));
	jdff dff_A_5l5XOZcE6_0(.dout(G863),.din(w_dff_A_5l5XOZcE6_0),.clk(gclk));
	jdff dff_A_qeZz187w9_1(.dout(w_dff_A_SsNyH2IT6_0),.din(w_dff_A_qeZz187w9_1),.clk(gclk));
	jdff dff_A_SsNyH2IT6_0(.dout(w_dff_A_aRHYR99A4_0),.din(w_dff_A_SsNyH2IT6_0),.clk(gclk));
	jdff dff_A_aRHYR99A4_0(.dout(w_dff_A_5X9sX5nS6_0),.din(w_dff_A_aRHYR99A4_0),.clk(gclk));
	jdff dff_A_5X9sX5nS6_0(.dout(w_dff_A_v0mXYtEf6_0),.din(w_dff_A_5X9sX5nS6_0),.clk(gclk));
	jdff dff_A_v0mXYtEf6_0(.dout(G865),.din(w_dff_A_v0mXYtEf6_0),.clk(gclk));
	jdff dff_A_JgOw3Pju8_1(.dout(w_dff_A_sJ5zsEQo0_0),.din(w_dff_A_JgOw3Pju8_1),.clk(gclk));
	jdff dff_A_sJ5zsEQo0_0(.dout(w_dff_A_FV1ZoX9j0_0),.din(w_dff_A_sJ5zsEQo0_0),.clk(gclk));
	jdff dff_A_FV1ZoX9j0_0(.dout(w_dff_A_u57xHKBL7_0),.din(w_dff_A_FV1ZoX9j0_0),.clk(gclk));
	jdff dff_A_u57xHKBL7_0(.dout(w_dff_A_Vsy9ohhV8_0),.din(w_dff_A_u57xHKBL7_0),.clk(gclk));
	jdff dff_A_Vsy9ohhV8_0(.dout(w_dff_A_yVWuYFiZ9_0),.din(w_dff_A_Vsy9ohhV8_0),.clk(gclk));
	jdff dff_A_yVWuYFiZ9_0(.dout(w_dff_A_1POWETG96_0),.din(w_dff_A_yVWuYFiZ9_0),.clk(gclk));
	jdff dff_A_1POWETG96_0(.dout(G867),.din(w_dff_A_1POWETG96_0),.clk(gclk));
	jdff dff_A_4kASBhIa2_1(.dout(w_dff_A_ALiaipha0_0),.din(w_dff_A_4kASBhIa2_1),.clk(gclk));
	jdff dff_A_ALiaipha0_0(.dout(w_dff_A_ULjYCfey9_0),.din(w_dff_A_ALiaipha0_0),.clk(gclk));
	jdff dff_A_ULjYCfey9_0(.dout(w_dff_A_YwmtFct39_0),.din(w_dff_A_ULjYCfey9_0),.clk(gclk));
	jdff dff_A_YwmtFct39_0(.dout(w_dff_A_Ax9852qS7_0),.din(w_dff_A_YwmtFct39_0),.clk(gclk));
	jdff dff_A_Ax9852qS7_0(.dout(w_dff_A_Lv5BfZpU2_0),.din(w_dff_A_Ax9852qS7_0),.clk(gclk));
	jdff dff_A_Lv5BfZpU2_0(.dout(w_dff_A_PVNJ4laq9_0),.din(w_dff_A_Lv5BfZpU2_0),.clk(gclk));
	jdff dff_A_PVNJ4laq9_0(.dout(w_dff_A_JnOKkwIw7_0),.din(w_dff_A_PVNJ4laq9_0),.clk(gclk));
	jdff dff_A_JnOKkwIw7_0(.dout(G869),.din(w_dff_A_JnOKkwIw7_0),.clk(gclk));
	jdff dff_A_EPXAZVpy7_2(.dout(w_dff_A_U2KV2y4S7_0),.din(w_dff_A_EPXAZVpy7_2),.clk(gclk));
	jdff dff_A_U2KV2y4S7_0(.dout(w_dff_A_8rFUIk6B2_0),.din(w_dff_A_U2KV2y4S7_0),.clk(gclk));
	jdff dff_A_8rFUIk6B2_0(.dout(G712),.din(w_dff_A_8rFUIk6B2_0),.clk(gclk));
	jdff dff_A_A0bT2Z0q4_2(.dout(w_dff_A_a1LOtgJo5_0),.din(w_dff_A_A0bT2Z0q4_2),.clk(gclk));
	jdff dff_A_a1LOtgJo5_0(.dout(w_dff_A_AonfvHhS2_0),.din(w_dff_A_a1LOtgJo5_0),.clk(gclk));
	jdff dff_A_AonfvHhS2_0(.dout(G727),.din(w_dff_A_AonfvHhS2_0),.clk(gclk));
	jdff dff_A_aSx5mPAn3_2(.dout(w_dff_A_98miXHfY4_0),.din(w_dff_A_aSx5mPAn3_2),.clk(gclk));
	jdff dff_A_98miXHfY4_0(.dout(w_dff_A_N8kAfbe75_0),.din(w_dff_A_98miXHfY4_0),.clk(gclk));
	jdff dff_A_N8kAfbe75_0(.dout(w_dff_A_B9YxbKYa1_0),.din(w_dff_A_N8kAfbe75_0),.clk(gclk));
	jdff dff_A_B9YxbKYa1_0(.dout(G732),.din(w_dff_A_B9YxbKYa1_0),.clk(gclk));
	jdff dff_A_EvzIhjy47_2(.dout(w_dff_A_lE73QFUH6_0),.din(w_dff_A_EvzIhjy47_2),.clk(gclk));
	jdff dff_A_lE73QFUH6_0(.dout(w_dff_A_brAqeK2M2_0),.din(w_dff_A_lE73QFUH6_0),.clk(gclk));
	jdff dff_A_brAqeK2M2_0(.dout(w_dff_A_gmj7bXCZ4_0),.din(w_dff_A_brAqeK2M2_0),.clk(gclk));
	jdff dff_A_gmj7bXCZ4_0(.dout(G737),.din(w_dff_A_gmj7bXCZ4_0),.clk(gclk));
	jdff dff_A_5IAg5QGE8_2(.dout(w_dff_A_cczKyqNy3_0),.din(w_dff_A_5IAg5QGE8_2),.clk(gclk));
	jdff dff_A_cczKyqNy3_0(.dout(w_dff_A_6fF4pLax1_0),.din(w_dff_A_cczKyqNy3_0),.clk(gclk));
	jdff dff_A_6fF4pLax1_0(.dout(w_dff_A_IUweG6cp8_0),.din(w_dff_A_6fF4pLax1_0),.clk(gclk));
	jdff dff_A_IUweG6cp8_0(.dout(w_dff_A_YPI6aWDE5_0),.din(w_dff_A_IUweG6cp8_0),.clk(gclk));
	jdff dff_A_YPI6aWDE5_0(.dout(G742),.din(w_dff_A_YPI6aWDE5_0),.clk(gclk));
	jdff dff_A_KRUM41us5_2(.dout(w_dff_A_Z4Js1zJe9_0),.din(w_dff_A_KRUM41us5_2),.clk(gclk));
	jdff dff_A_Z4Js1zJe9_0(.dout(w_dff_A_XS2z2DUo2_0),.din(w_dff_A_Z4Js1zJe9_0),.clk(gclk));
	jdff dff_A_XS2z2DUo2_0(.dout(w_dff_A_uO8HpWfq1_0),.din(w_dff_A_XS2z2DUo2_0),.clk(gclk));
	jdff dff_A_uO8HpWfq1_0(.dout(G772),.din(w_dff_A_uO8HpWfq1_0),.clk(gclk));
	jdff dff_A_RrTJUjUs0_2(.dout(w_dff_A_uaTZb3Xr7_0),.din(w_dff_A_RrTJUjUs0_2),.clk(gclk));
	jdff dff_A_uaTZb3Xr7_0(.dout(w_dff_A_Yb1mhufn6_0),.din(w_dff_A_uaTZb3Xr7_0),.clk(gclk));
	jdff dff_A_Yb1mhufn6_0(.dout(w_dff_A_FRtqdOhg9_0),.din(w_dff_A_Yb1mhufn6_0),.clk(gclk));
	jdff dff_A_FRtqdOhg9_0(.dout(G777),.din(w_dff_A_FRtqdOhg9_0),.clk(gclk));
	jdff dff_A_sdnfD5209_2(.dout(w_dff_A_MxF9yI1R1_0),.din(w_dff_A_sdnfD5209_2),.clk(gclk));
	jdff dff_A_MxF9yI1R1_0(.dout(w_dff_A_oHh2Qmiy7_0),.din(w_dff_A_MxF9yI1R1_0),.clk(gclk));
	jdff dff_A_oHh2Qmiy7_0(.dout(w_dff_A_MnACyr4n1_0),.din(w_dff_A_oHh2Qmiy7_0),.clk(gclk));
	jdff dff_A_MnACyr4n1_0(.dout(w_dff_A_RgW3IAYd3_0),.din(w_dff_A_MnACyr4n1_0),.clk(gclk));
	jdff dff_A_RgW3IAYd3_0(.dout(G782),.din(w_dff_A_RgW3IAYd3_0),.clk(gclk));
	jdff dff_A_Gwj90k1Q2_2(.dout(w_dff_A_9ysUNOTD0_0),.din(w_dff_A_Gwj90k1Q2_2),.clk(gclk));
	jdff dff_A_9ysUNOTD0_0(.dout(w_dff_A_QHls6gRw0_0),.din(w_dff_A_9ysUNOTD0_0),.clk(gclk));
	jdff dff_A_QHls6gRw0_0(.dout(w_dff_A_0GymOqF51_0),.din(w_dff_A_QHls6gRw0_0),.clk(gclk));
	jdff dff_A_0GymOqF51_0(.dout(G645),.din(w_dff_A_0GymOqF51_0),.clk(gclk));
	jdff dff_A_G2E6wyy35_2(.dout(w_dff_A_LNUwRMhl1_0),.din(w_dff_A_G2E6wyy35_2),.clk(gclk));
	jdff dff_A_LNUwRMhl1_0(.dout(w_dff_A_7VnH1jEX5_0),.din(w_dff_A_LNUwRMhl1_0),.clk(gclk));
	jdff dff_A_7VnH1jEX5_0(.dout(G648),.din(w_dff_A_7VnH1jEX5_0),.clk(gclk));
	jdff dff_A_sGgb8Vsx5_2(.dout(w_dff_A_Ln59w4Pj7_0),.din(w_dff_A_sGgb8Vsx5_2),.clk(gclk));
	jdff dff_A_Ln59w4Pj7_0(.dout(w_dff_A_OapA63Vb1_0),.din(w_dff_A_Ln59w4Pj7_0),.clk(gclk));
	jdff dff_A_OapA63Vb1_0(.dout(G651),.din(w_dff_A_OapA63Vb1_0),.clk(gclk));
	jdff dff_A_7PhnTXaZ8_2(.dout(w_dff_A_U3jvNd3r3_0),.din(w_dff_A_7PhnTXaZ8_2),.clk(gclk));
	jdff dff_A_U3jvNd3r3_0(.dout(G654),.din(w_dff_A_U3jvNd3r3_0),.clk(gclk));
	jdff dff_A_RjIELs5s6_2(.dout(w_dff_A_lDl6L8a50_0),.din(w_dff_A_RjIELs5s6_2),.clk(gclk));
	jdff dff_A_lDl6L8a50_0(.dout(w_dff_A_G4lu5pDk8_0),.din(w_dff_A_lDl6L8a50_0),.clk(gclk));
	jdff dff_A_G4lu5pDk8_0(.dout(w_dff_A_JLHAKdxX1_0),.din(w_dff_A_G4lu5pDk8_0),.clk(gclk));
	jdff dff_A_JLHAKdxX1_0(.dout(G679),.din(w_dff_A_JLHAKdxX1_0),.clk(gclk));
	jdff dff_A_nq2iXq3a8_2(.dout(w_dff_A_AaUtWyPQ7_0),.din(w_dff_A_nq2iXq3a8_2),.clk(gclk));
	jdff dff_A_AaUtWyPQ7_0(.dout(w_dff_A_sqk5T6Ib0_0),.din(w_dff_A_AaUtWyPQ7_0),.clk(gclk));
	jdff dff_A_sqk5T6Ib0_0(.dout(G682),.din(w_dff_A_sqk5T6Ib0_0),.clk(gclk));
	jdff dff_A_LZXvWiyX4_2(.dout(w_dff_A_W7owOvbo8_0),.din(w_dff_A_LZXvWiyX4_2),.clk(gclk));
	jdff dff_A_W7owOvbo8_0(.dout(w_dff_A_rCUTpasy5_0),.din(w_dff_A_W7owOvbo8_0),.clk(gclk));
	jdff dff_A_rCUTpasy5_0(.dout(G685),.din(w_dff_A_rCUTpasy5_0),.clk(gclk));
	jdff dff_A_wCM0Ubje4_2(.dout(w_dff_A_G8P3GmPF3_0),.din(w_dff_A_wCM0Ubje4_2),.clk(gclk));
	jdff dff_A_G8P3GmPF3_0(.dout(G688),.din(w_dff_A_G8P3GmPF3_0),.clk(gclk));
	jdff dff_A_NFX8Ro7t6_2(.dout(w_dff_A_PLc1xrpK6_0),.din(w_dff_A_NFX8Ro7t6_2),.clk(gclk));
	jdff dff_A_PLc1xrpK6_0(.dout(w_dff_A_C7vfaVHx9_0),.din(w_dff_A_PLc1xrpK6_0),.clk(gclk));
	jdff dff_A_C7vfaVHx9_0(.dout(w_dff_A_CTAO9IKv4_0),.din(w_dff_A_C7vfaVHx9_0),.clk(gclk));
	jdff dff_A_CTAO9IKv4_0(.dout(G843),.din(w_dff_A_CTAO9IKv4_0),.clk(gclk));
	jdff dff_A_bDIpSuPb9_2(.dout(w_dff_A_lrlwHHYA8_0),.din(w_dff_A_bDIpSuPb9_2),.clk(gclk));
	jdff dff_A_lrlwHHYA8_0(.dout(w_dff_A_mKw851y78_0),.din(w_dff_A_lrlwHHYA8_0),.clk(gclk));
	jdff dff_A_mKw851y78_0(.dout(w_dff_A_VCgMwWwu9_0),.din(w_dff_A_mKw851y78_0),.clk(gclk));
	jdff dff_A_VCgMwWwu9_0(.dout(G882),.din(w_dff_A_VCgMwWwu9_0),.clk(gclk));
	jdff dff_A_5NIX1Iv46_2(.dout(G767),.din(w_dff_A_5NIX1Iv46_2),.clk(gclk));
	jdff dff_A_X47nM5mB6_2(.dout(G807),.din(w_dff_A_X47nM5mB6_2),.clk(gclk));
endmodule

