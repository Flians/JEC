// Benchmark "c5315" written by ABC on Wed May 27 22:07:38 2020

module rf_c5315 ( 
    G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37,
    G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79,
    G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106,
    G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122,
    G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G140,
    G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170, G173,
    G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206, G209,
    G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248, G251,
    G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292, G293,
    G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335, G338,
    G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386, G389,
    G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514, G523,
    G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691,
    G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717,
    G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115,
    G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612,
    G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921,
    G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636,
    G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626,
    G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623,
    G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000,
    G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802,
    G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826,
    G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742,
    G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843,
    G882, G767, G807, G658, G690  );
  input  G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34,
    G37, G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76,
    G79, G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103,
    G106, G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121,
    G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137,
    G140, G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170,
    G173, G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206,
    G209, G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248,
    G251, G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292,
    G293, G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335,
    G338, G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386,
    G389, G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514,
    G523, G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690,
    G1691, G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552,
    G3717, G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115;
  output G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611,
    G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923,
    G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593,
    G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615,
    G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861,
    G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998,
    G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792,
    G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813,
    G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732,
    G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685,
    G688, G843, G882, G767, G807, G658, G690;
  wire n314, n316, n318, n320, n321, n325, n326, n327, n328, n329, n330,
    n332, n333, n334, n335, n336, n338, n340, n341, n342, n343, n345, n346,
    n347, n348, n350, n351, n352, n353, n355, n356, n357, n358, n360, n361,
    n362, n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
    n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
    n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
    n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
    n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420, n421,
    n422, n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
    n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444, n445,
    n446, n447, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
    n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
    n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481, n482,
    n483, n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
    n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
    n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
    n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
    n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541, n542,
    n543, n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
    n556, n557, n558, n559, n560, n561, n562, n563, n564, n565, n566, n567,
    n568, n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
    n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
    n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602, n603,
    n604, n605, n606, n607, n609, n610, n611, n612, n613, n614, n615, n616,
    n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
    n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
    n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
    n654, n655, n656, n657, n658, n659, n660, n661, n663, n664, n665, n666,
    n667, n668, n669, n670, n671, n673, n674, n675, n676, n677, n678, n679,
    n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691,
    n692, n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
    n704, n705, n706, n707, n708, n709, n711, n712, n713, n714, n715, n716,
    n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
    n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740,
    n741, n742, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n758, n759, n760, n761, n762, n763, n764, n765, n766,
    n767, n768, n769, n771, n772, n773, n774, n775, n776, n777, n779, n780,
    n781, n782, n783, n784, n785, n786, n787, n788, n789, n791, n792, n793,
    n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n806,
    n807, n808, n809, n810, n811, n812, n813, n814, n816, n817, n818, n819,
    n820, n821, n822, n823, n824, n825, n826, n828, n829, n830, n831, n832,
    n833, n834, n835, n836, n837, n839, n840, n841, n842, n843, n844, n845,
    n846, n847, n848, n849, n850, n852, n853, n854, n855, n856, n857, n858,
    n859, n860, n861, n862, n863, n864, n865, n866, n867, n869, n870, n871,
    n872, n873, n874, n876, n877, n878, n879, n880, n881, n882, n883, n884,
    n885, n886, n887, n889, n890, n891, n892, n893, n894, n895, n896, n897,
    n898, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
    n911, n912, n913, n914, n916, n917, n918, n919, n920, n921, n922, n923,
    n924, n925, n926, n928, n929, n930, n931, n932, n933, n934, n935, n936,
    n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
    n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959, n960,
    n961, n962, n963, n964, n965, n967, n968, n969, n970, n971, n972, n973,
    n974, n975, n976, n977, n978, n979, n980, n981, n982, n984, n985, n986,
    n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1021,
    n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1030, n1031, n1032,
    n1033, n1034, n1035, n1036, n1037, n1039, n1040, n1041, n1042, n1043,
    n1044, n1045, n1046, n1048, n1049, n1050, n1051, n1052, n1053, n1055,
    n1056, n1057, n1058, n1059, n1060, n1062, n1063, n1064, n1065, n1066,
    n1067, n1069, n1070, n1071, n1072, n1073, n1074, n1076, n1077, n1078,
    n1079, n1080, n1081, n1082, n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1100, n1101,
    n1102, n1103, n1104, n1105, n1106, n1108, n1109, n1110, n1111, n1112,
    n1113, n1114, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1124,
    n1125, n1126, n1127, n1128, n1129, n1130, n1132, n1133, n1134, n1135,
    n1136, n1137, n1138, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
    n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1157,
    n1159, n1160, n1161, n1162, n1163, n1165, n1166, n1167, n1168, n1169,
    n1171, n1172, n1173, n1174, n1175, n1177, n1178, n1179, n1180, n1181,
    n1182, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1192, n1193,
    n1194, n1195, n1196, n1197, n1199, n1200, n1201, n1202, n1203, n1204,
    n1205, n1207, n1208, n1209, n1210, n1211, n1213, n1214, n1215, n1216,
    n1217, n1218, n1220, n1221, n1222, n1223, n1224, n1225, n1227, n1228,
    n1229, n1230, n1231, n1232, n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1251,
    n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1260, n1261, n1262,
    n1263, n1264, n1265, n1267, n1268, n1269, n1270, n1271, n1272, n1274,
    n1275, n1276, n1277, n1278, n1279, n1281, n1282, n1283, n1284, n1285,
    n1286, n1287, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1297,
    n1298, n1299, n1300, n1301, n1302, n1303, n1305, n1306, n1307, n1308,
    n1309, n1310, n1311, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
    n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1329, n1330, n1331,
    n1332, n1333, n1334, n1335, n1337, n1338, n1339, n1340, n1341, n1342,
    n1343, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
    n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
    n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
    n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
    n1384, n1385, n1386, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
    n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
    n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
    n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
    n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
    n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
    n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1454, n1455,
    n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
    n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
    n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
    n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
    n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
    n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
    n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
    n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
    n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
    n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
    n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
    n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
    n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
    n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
    n1596, n1597, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
    n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1617,
    n1618, n1619, n1620, n1621, n1622, n1624, n1625, n1626, n1627, n1628,
    n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
    n1639, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
    n1650, n1651;
  jnot g0000(.din(G545), .dout(G594));
  jnot g0001(.din(G348), .dout(G599));
  jnot g0002(.din(G366), .dout(G600));
  jand g0003(.dina(G562), .dinb(G552), .dout(G601));
  jnot g0004(.din(G549), .dout(G602));
  jnot g0005(.din(G338), .dout(G611));
  jnot g0006(.din(G358), .dout(G612));
  jand g0007(.dina(G145), .dinb(G141), .dout(G810));
  jnot g0008(.din(G245), .dout(G848));
  jnot g0009(.din(G552), .dout(G849));
  jnot g0010(.din(G562), .dout(G850));
  jnot g0011(.din(G559), .dout(G851));
  jand g0012(.dina(G373), .dinb(G1), .dout(G634));
  jnot g0013(.din(G3173), .dout(n314));
  jand g0014(.dina(n314), .dinb(G136), .dout(G815));
  jnot g0015(.din(G27), .dout(n316));
  jor  g0016(.dina(G2824), .dinb(n316), .dout(G845));
  jand g0017(.dina(G556), .dinb(G386), .dout(n318));
  jnot g0018(.din(n318), .dout(G847));
  jnot g0019(.din(G140), .dout(n320));
  jnot g0020(.din(G31), .dout(n321));
  jor  g0021(.dina(n321), .dinb(n316), .dout(G809));
  jor  g0022(.dina(G809), .dinb(n320), .dout(G656));
  jnot g0023(.din(G299), .dout(G593));
  jnot g0024(.din(G86), .dout(n325));
  jnot g0025(.din(G2358), .dout(n326));
  jand g0026(.dina(n326), .dinb(n325), .dout(n327));
  jnot g0027(.din(G87), .dout(n328));
  jand g0028(.dina(G2358), .dinb(n328), .dout(n329));
  jor  g0029(.dina(n329), .dinb(G809), .dout(n330));
  jor  g0030(.dina(n330), .dinb(n327), .dout(G636));
  jnot g0031(.din(G88), .dout(n332));
  jand g0032(.dina(n326), .dinb(n332), .dout(n333));
  jnot g0033(.din(G34), .dout(n334));
  jand g0034(.dina(G2358), .dinb(n334), .dout(n335));
  jor  g0035(.dina(n335), .dinb(G809), .dout(n336));
  jor  g0036(.dina(n336), .dinb(n333), .dout(G704));
  jnot g0037(.din(G83), .dout(n338));
  jor  g0038(.dina(G809), .dinb(n338), .dout(G820));
  jand g0039(.dina(n326), .dinb(G24), .dout(n340));
  jand g0040(.dina(G2358), .dinb(G25), .dout(n341));
  jor  g0041(.dina(n341), .dinb(G809), .dout(n342));
  jor  g0042(.dina(n342), .dinb(n340), .dout(n343));
  jand g0043(.dina(n343), .dinb(G141), .dout(G639));
  jand g0044(.dina(n326), .dinb(G26), .dout(n345));
  jand g0045(.dina(G2358), .dinb(G81), .dout(n346));
  jor  g0046(.dina(n346), .dinb(G809), .dout(n347));
  jor  g0047(.dina(n347), .dinb(n345), .dout(n348));
  jand g0048(.dina(n348), .dinb(G141), .dout(G673));
  jand g0049(.dina(n326), .dinb(G79), .dout(n350));
  jand g0050(.dina(G2358), .dinb(G23), .dout(n351));
  jor  g0051(.dina(n351), .dinb(G809), .dout(n352));
  jor  g0052(.dina(n352), .dinb(n350), .dout(n353));
  jand g0053(.dina(n353), .dinb(G141), .dout(G707));
  jand g0054(.dina(n326), .dinb(G82), .dout(n355));
  jand g0055(.dina(G2358), .dinb(G80), .dout(n356));
  jor  g0056(.dina(n356), .dinb(G809), .dout(n357));
  jor  g0057(.dina(n357), .dinb(n355), .dout(n358));
  jand g0058(.dina(n358), .dinb(G141), .dout(G715));
  jnot g0059(.din(G308), .dout(n360));
  jand g0060(.dina(n360), .dinb(G251), .dout(n361));
  jnot g0061(.din(G479), .dout(n362));
  jand g0062(.dina(G308), .dinb(G248), .dout(n363));
  jor  g0063(.dina(n363), .dinb(n362), .dout(n364));
  jor  g0064(.dina(n364), .dinb(n361), .dout(n365));
  jnot g0065(.din(G254), .dout(n366));
  jand g0066(.dina(n360), .dinb(n366), .dout(n367));
  jnot g0067(.din(G242), .dout(n368));
  jand g0068(.dina(G308), .dinb(n368), .dout(n369));
  jor  g0069(.dina(n369), .dinb(G479), .dout(n370));
  jor  g0070(.dina(n370), .dinb(n367), .dout(n371));
  jand g0071(.dina(n371), .dinb(n365), .dout(n372));
  jnot g0072(.din(G316), .dout(n373));
  jand g0073(.dina(n373), .dinb(G251), .dout(n374));
  jnot g0074(.din(G490), .dout(n375));
  jand g0075(.dina(G316), .dinb(G248), .dout(n376));
  jor  g0076(.dina(n376), .dinb(n375), .dout(n377));
  jor  g0077(.dina(n377), .dinb(n374), .dout(n378));
  jand g0078(.dina(n373), .dinb(n366), .dout(n379));
  jand g0079(.dina(G316), .dinb(n368), .dout(n380));
  jor  g0080(.dina(n380), .dinb(G490), .dout(n381));
  jor  g0081(.dina(n381), .dinb(n379), .dout(n382));
  jand g0082(.dina(n382), .dinb(n378), .dout(n383));
  jand g0083(.dina(n383), .dinb(n372), .dout(n384));
  jnot g0084(.din(G351), .dout(n385));
  jnot g0085(.din(G3550), .dout(n386));
  jand g0086(.dina(n386), .dinb(n385), .dout(n387));
  jnot g0087(.din(G534), .dout(n388));
  jnot g0088(.din(G3552), .dout(n389));
  jand g0089(.dina(n389), .dinb(G351), .dout(n390));
  jor  g0090(.dina(n390), .dinb(n388), .dout(n391));
  jor  g0091(.dina(n391), .dinb(n387), .dout(n392));
  jand g0092(.dina(G3548), .dinb(n385), .dout(n393));
  jand g0093(.dina(G3546), .dinb(G351), .dout(n394));
  jor  g0094(.dina(n394), .dinb(G534), .dout(n395));
  jor  g0095(.dina(n395), .dinb(n393), .dout(n396));
  jand g0096(.dina(n396), .dinb(n392), .dout(n397));
  jnot g0097(.din(G293), .dout(n398));
  jand g0098(.dina(n398), .dinb(n366), .dout(n399));
  jand g0099(.dina(G293), .dinb(n368), .dout(n400));
  jor  g0100(.dina(n400), .dinb(n399), .dout(n401));
  jnot g0101(.din(G251), .dout(n402));
  jnot g0102(.din(G302), .dout(n403));
  jand g0103(.dina(n403), .dinb(n402), .dout(n404));
  jnot g0104(.din(G248), .dout(n405));
  jand g0105(.dina(G302), .dinb(n405), .dout(n406));
  jor  g0106(.dina(n406), .dinb(n404), .dout(n407));
  jnot g0107(.din(n407), .dout(n408));
  jand g0108(.dina(n408), .dinb(n401), .dout(n409));
  jnot g0109(.din(G514), .dout(n410));
  jnot g0110(.din(G3546), .dout(n411));
  jand g0111(.dina(n411), .dinb(n410), .dout(n412));
  jand g0112(.dina(G3552), .dinb(G514), .dout(n413));
  jor  g0113(.dina(n413), .dinb(n412), .dout(n414));
  jnot g0114(.din(n414), .dout(n415));
  jnot g0115(.din(G361), .dout(n416));
  jand g0116(.dina(n416), .dinb(n402), .dout(n417));
  jand g0117(.dina(G361), .dinb(n405), .dout(n418));
  jor  g0118(.dina(n418), .dinb(n417), .dout(n419));
  jnot g0119(.din(n419), .dout(n420));
  jand g0120(.dina(n420), .dinb(n415), .dout(n421));
  jand g0121(.dina(n421), .dinb(n409), .dout(n422));
  jand g0122(.dina(n422), .dinb(n397), .dout(n423));
  jnot g0123(.din(G324), .dout(n424));
  jand g0124(.dina(n386), .dinb(n424), .dout(n425));
  jnot g0125(.din(G503), .dout(n426));
  jand g0126(.dina(n389), .dinb(G324), .dout(n427));
  jor  g0127(.dina(n427), .dinb(n426), .dout(n428));
  jor  g0128(.dina(n428), .dinb(n425), .dout(n429));
  jand g0129(.dina(G3548), .dinb(n424), .dout(n430));
  jand g0130(.dina(G3546), .dinb(G324), .dout(n431));
  jor  g0131(.dina(n431), .dinb(G503), .dout(n432));
  jor  g0132(.dina(n432), .dinb(n430), .dout(n433));
  jand g0133(.dina(n433), .dinb(n429), .dout(n434));
  jnot g0134(.din(G341), .dout(n435));
  jand g0135(.dina(n386), .dinb(n435), .dout(n436));
  jnot g0136(.din(G523), .dout(n437));
  jand g0137(.dina(n389), .dinb(G341), .dout(n438));
  jor  g0138(.dina(n438), .dinb(n437), .dout(n439));
  jor  g0139(.dina(n439), .dinb(n436), .dout(n440));
  jand g0140(.dina(G3548), .dinb(n435), .dout(n441));
  jand g0141(.dina(G3546), .dinb(G341), .dout(n442));
  jor  g0142(.dina(n442), .dinb(G523), .dout(n443));
  jor  g0143(.dina(n443), .dinb(n441), .dout(n444));
  jand g0144(.dina(n444), .dinb(n440), .dout(n445));
  jand g0145(.dina(n445), .dinb(n434), .dout(n446));
  jand g0146(.dina(n446), .dinb(n423), .dout(n447));
  jand g0147(.dina(n447), .dinb(n384), .dout(G598));
  jnot g0148(.din(G265), .dout(n449));
  jand g0149(.dina(n386), .dinb(n449), .dout(n450));
  jnot g0150(.din(G400), .dout(n451));
  jand g0151(.dina(n389), .dinb(G265), .dout(n452));
  jor  g0152(.dina(n452), .dinb(n451), .dout(n453));
  jor  g0153(.dina(n453), .dinb(n450), .dout(n454));
  jand g0154(.dina(G3548), .dinb(n449), .dout(n455));
  jand g0155(.dina(G3546), .dinb(G265), .dout(n456));
  jor  g0156(.dina(n456), .dinb(G400), .dout(n457));
  jor  g0157(.dina(n457), .dinb(n455), .dout(n458));
  jand g0158(.dina(n458), .dinb(n454), .dout(n459));
  jnot g0159(.din(G234), .dout(n460));
  jand g0160(.dina(n386), .dinb(n460), .dout(n461));
  jnot g0161(.din(G435), .dout(n462));
  jand g0162(.dina(n389), .dinb(G234), .dout(n463));
  jor  g0163(.dina(n463), .dinb(n462), .dout(n464));
  jor  g0164(.dina(n464), .dinb(n461), .dout(n465));
  jand g0165(.dina(G3548), .dinb(n460), .dout(n466));
  jand g0166(.dina(G3546), .dinb(G234), .dout(n467));
  jor  g0167(.dina(n467), .dinb(G435), .dout(n468));
  jor  g0168(.dina(n468), .dinb(n466), .dout(n469));
  jand g0169(.dina(n469), .dinb(n465), .dout(n470));
  jnot g0170(.din(G257), .dout(n471));
  jand g0171(.dina(n386), .dinb(n471), .dout(n472));
  jnot g0172(.din(G389), .dout(n473));
  jand g0173(.dina(n389), .dinb(G257), .dout(n474));
  jor  g0174(.dina(n474), .dinb(n473), .dout(n475));
  jor  g0175(.dina(n475), .dinb(n472), .dout(n476));
  jand g0176(.dina(G3548), .dinb(n471), .dout(n477));
  jand g0177(.dina(G3546), .dinb(G257), .dout(n478));
  jor  g0178(.dina(n478), .dinb(G389), .dout(n479));
  jor  g0179(.dina(n479), .dinb(n477), .dout(n480));
  jand g0180(.dina(n480), .dinb(n476), .dout(n481));
  jand g0181(.dina(n481), .dinb(n470), .dout(n482));
  jand g0182(.dina(n482), .dinb(n459), .dout(n483));
  jnot g0183(.din(G273), .dout(n484));
  jand g0184(.dina(n386), .dinb(n484), .dout(n485));
  jnot g0185(.din(G411), .dout(n486));
  jand g0186(.dina(n389), .dinb(G273), .dout(n487));
  jor  g0187(.dina(n487), .dinb(n486), .dout(n488));
  jor  g0188(.dina(n488), .dinb(n485), .dout(n489));
  jand g0189(.dina(G3548), .dinb(n484), .dout(n490));
  jand g0190(.dina(G3546), .dinb(G273), .dout(n491));
  jor  g0191(.dina(n491), .dinb(G411), .dout(n492));
  jor  g0192(.dina(n492), .dinb(n490), .dout(n493));
  jand g0193(.dina(n493), .dinb(n489), .dout(n494));
  jnot g0194(.din(G281), .dout(n495));
  jand g0195(.dina(n386), .dinb(n495), .dout(n496));
  jnot g0196(.din(G374), .dout(n497));
  jand g0197(.dina(n389), .dinb(G281), .dout(n498));
  jor  g0198(.dina(n498), .dinb(n497), .dout(n499));
  jor  g0199(.dina(n499), .dinb(n496), .dout(n500));
  jand g0200(.dina(G3548), .dinb(n495), .dout(n501));
  jand g0201(.dina(G3546), .dinb(G281), .dout(n502));
  jor  g0202(.dina(n502), .dinb(G374), .dout(n503));
  jor  g0203(.dina(n503), .dinb(n501), .dout(n504));
  jand g0204(.dina(n504), .dinb(n500), .dout(n505));
  jand g0205(.dina(n505), .dinb(n494), .dout(n506));
  jnot g0206(.din(G218), .dout(n507));
  jand g0207(.dina(n386), .dinb(n507), .dout(n508));
  jnot g0208(.din(G468), .dout(n509));
  jand g0209(.dina(n389), .dinb(G218), .dout(n510));
  jor  g0210(.dina(n510), .dinb(n509), .dout(n511));
  jor  g0211(.dina(n511), .dinb(n508), .dout(n512));
  jand g0212(.dina(G3548), .dinb(n507), .dout(n513));
  jand g0213(.dina(G3546), .dinb(G218), .dout(n514));
  jor  g0214(.dina(n514), .dinb(G468), .dout(n515));
  jor  g0215(.dina(n515), .dinb(n513), .dout(n516));
  jand g0216(.dina(n516), .dinb(n512), .dout(n517));
  jnot g0217(.din(G206), .dout(n518));
  jand g0218(.dina(G251), .dinb(n518), .dout(n519));
  jnot g0219(.din(G446), .dout(n520));
  jand g0220(.dina(G248), .dinb(G206), .dout(n521));
  jor  g0221(.dina(n521), .dinb(n520), .dout(n522));
  jor  g0222(.dina(n522), .dinb(n519), .dout(n523));
  jand g0223(.dina(n366), .dinb(n518), .dout(n524));
  jand g0224(.dina(n368), .dinb(G206), .dout(n525));
  jor  g0225(.dina(n525), .dinb(G446), .dout(n526));
  jor  g0226(.dina(n526), .dinb(n524), .dout(n527));
  jand g0227(.dina(n527), .dinb(n523), .dout(n528));
  jand g0228(.dina(n528), .dinb(n517), .dout(n529));
  jnot g0229(.din(G226), .dout(n530));
  jand g0230(.dina(n386), .dinb(n530), .dout(n531));
  jnot g0231(.din(G422), .dout(n532));
  jand g0232(.dina(n389), .dinb(G226), .dout(n533));
  jor  g0233(.dina(n533), .dinb(n532), .dout(n534));
  jor  g0234(.dina(n534), .dinb(n531), .dout(n535));
  jand g0235(.dina(G3548), .dinb(n530), .dout(n536));
  jand g0236(.dina(G3546), .dinb(G226), .dout(n537));
  jor  g0237(.dina(n537), .dinb(G422), .dout(n538));
  jor  g0238(.dina(n538), .dinb(n536), .dout(n539));
  jand g0239(.dina(n539), .dinb(n535), .dout(n540));
  jnot g0240(.din(G210), .dout(n541));
  jand g0241(.dina(n386), .dinb(n541), .dout(n542));
  jnot g0242(.din(G457), .dout(n543));
  jand g0243(.dina(n389), .dinb(G210), .dout(n544));
  jor  g0244(.dina(n544), .dinb(n543), .dout(n545));
  jor  g0245(.dina(n545), .dinb(n542), .dout(n546));
  jand g0246(.dina(G3548), .dinb(n541), .dout(n547));
  jand g0247(.dina(G3546), .dinb(G210), .dout(n548));
  jor  g0248(.dina(n548), .dinb(G457), .dout(n549));
  jor  g0249(.dina(n549), .dinb(n547), .dout(n550));
  jand g0250(.dina(n550), .dinb(n546), .dout(n551));
  jand g0251(.dina(n551), .dinb(n540), .dout(n552));
  jand g0252(.dina(n552), .dinb(n529), .dout(n553));
  jand g0253(.dina(n553), .dinb(n506), .dout(n554));
  jand g0254(.dina(n554), .dinb(n483), .dout(G610));
  jnot g0255(.din(G335), .dout(n556));
  jor  g0256(.dina(n556), .dinb(G241), .dout(n557));
  jand g0257(.dina(n556), .dinb(n460), .dout(n558));
  jnot g0258(.din(n558), .dout(n559));
  jand g0259(.dina(n559), .dinb(n557), .dout(n560));
  jxor g0260(.dina(n560), .dinb(G435), .dout(n561));
  jnot g0261(.din(n561), .dout(n562));
  jnot g0262(.din(G288), .dout(n563));
  jand g0263(.dina(G335), .dinb(n563), .dout(n564));
  jand g0264(.dina(n556), .dinb(n495), .dout(n565));
  jor  g0265(.dina(n565), .dinb(n564), .dout(n566));
  jxor g0266(.dina(n566), .dinb(n497), .dout(n567));
  jor  g0267(.dina(n556), .dinb(G280), .dout(n568));
  jor  g0268(.dina(G335), .dinb(G273), .dout(n569));
  jand g0269(.dina(n569), .dinb(n568), .dout(n570));
  jxor g0270(.dina(n570), .dinb(n486), .dout(n571));
  jnot g0271(.din(n571), .dout(n572));
  jand g0272(.dina(n572), .dinb(n567), .dout(n573));
  jnot g0273(.din(n573), .dout(n574));
  jor  g0274(.dina(n556), .dinb(G264), .dout(n575));
  jor  g0275(.dina(G335), .dinb(G257), .dout(n576));
  jand g0276(.dina(n576), .dinb(n575), .dout(n577));
  jxor g0277(.dina(n577), .dinb(n473), .dout(n578));
  jnot g0278(.din(G272), .dout(n579));
  jand g0279(.dina(G335), .dinb(n579), .dout(n580));
  jand g0280(.dina(n556), .dinb(n449), .dout(n581));
  jor  g0281(.dina(n581), .dinb(n580), .dout(n582));
  jxor g0282(.dina(n582), .dinb(G400), .dout(n583));
  jor  g0283(.dina(n583), .dinb(n578), .dout(n584));
  jor  g0284(.dina(n584), .dinb(n574), .dout(n585));
  jor  g0285(.dina(n585), .dinb(n562), .dout(n586));
  jnot g0286(.din(n586), .dout(n587));
  jor  g0287(.dina(n556), .dinb(G217), .dout(n588));
  jor  g0288(.dina(G335), .dinb(G210), .dout(n589));
  jand g0289(.dina(n589), .dinb(n588), .dout(n590));
  jxor g0290(.dina(n590), .dinb(G457), .dout(n591));
  jor  g0291(.dina(n556), .dinb(G209), .dout(n592));
  jand g0292(.dina(n556), .dinb(n518), .dout(n593));
  jnot g0293(.din(n593), .dout(n594));
  jand g0294(.dina(n594), .dinb(n592), .dout(n595));
  jxor g0295(.dina(n595), .dinb(G446), .dout(n596));
  jand g0296(.dina(n596), .dinb(n591), .dout(n597));
  jor  g0297(.dina(n556), .dinb(G233), .dout(n598));
  jor  g0298(.dina(G335), .dinb(G226), .dout(n599));
  jand g0299(.dina(n599), .dinb(n598), .dout(n600));
  jxor g0300(.dina(n600), .dinb(G422), .dout(n601));
  jor  g0301(.dina(n556), .dinb(G225), .dout(n602));
  jor  g0302(.dina(G335), .dinb(G218), .dout(n603));
  jand g0303(.dina(n603), .dinb(n602), .dout(n604));
  jxor g0304(.dina(n604), .dinb(G468), .dout(n605));
  jand g0305(.dina(n605), .dinb(n601), .dout(n606));
  jand g0306(.dina(n606), .dinb(n597), .dout(n607));
  jand g0307(.dina(n607), .dinb(n587), .dout(G588));
  jnot g0308(.din(G332), .dout(n609));
  jor  g0309(.dina(n609), .dinb(G331), .dout(n610));
  jand g0310(.dina(n609), .dinb(n424), .dout(n611));
  jnot g0311(.din(n611), .dout(n612));
  jand g0312(.dina(n612), .dinb(n610), .dout(n613));
  jxor g0313(.dina(n613), .dinb(G503), .dout(n614));
  jor  g0314(.dina(G358), .dinb(n609), .dout(n615));
  jor  g0315(.dina(G351), .dinb(G332), .dout(n616));
  jand g0316(.dina(n616), .dinb(n615), .dout(n617));
  jxor g0317(.dina(n617), .dinb(n388), .dout(n618));
  jand g0318(.dina(G600), .dinb(G332), .dout(n619));
  jand g0319(.dina(n416), .dinb(n609), .dout(n620));
  jor  g0320(.dina(n620), .dinb(n619), .dout(n621));
  jnot g0321(.din(n621), .dout(n622));
  jor  g0322(.dina(n622), .dinb(n618), .dout(n623));
  jand g0323(.dina(G611), .dinb(G332), .dout(n624));
  jxor g0324(.dina(n624), .dinb(G514), .dout(n625));
  jor  g0325(.dina(G348), .dinb(n609), .dout(n626));
  jor  g0326(.dina(G341), .dinb(G332), .dout(n627));
  jand g0327(.dina(n627), .dinb(n626), .dout(n628));
  jxor g0328(.dina(n628), .dinb(n437), .dout(n629));
  jor  g0329(.dina(n629), .dinb(n625), .dout(n630));
  jor  g0330(.dina(n630), .dinb(n623), .dout(n631));
  jnot g0331(.din(n631), .dout(n632));
  jand g0332(.dina(n632), .dinb(n614), .dout(n633));
  jand g0333(.dina(G332), .dinb(G593), .dout(n634));
  jand g0334(.dina(n609), .dinb(n398), .dout(n635));
  jor  g0335(.dina(n635), .dinb(n634), .dout(n636));
  jor  g0336(.dina(n609), .dinb(G307), .dout(n637));
  jand g0337(.dina(n609), .dinb(n403), .dout(n638));
  jnot g0338(.din(n638), .dout(n639));
  jand g0339(.dina(n639), .dinb(n637), .dout(n640));
  jnot g0340(.din(n640), .dout(n641));
  jand g0341(.dina(n641), .dinb(n636), .dout(n642));
  jor  g0342(.dina(n609), .dinb(G315), .dout(n643));
  jor  g0343(.dina(G332), .dinb(G308), .dout(n644));
  jand g0344(.dina(n644), .dinb(n643), .dout(n645));
  jxor g0345(.dina(n645), .dinb(G479), .dout(n646));
  jor  g0346(.dina(n609), .dinb(G323), .dout(n647));
  jor  g0347(.dina(G332), .dinb(G316), .dout(n648));
  jand g0348(.dina(n648), .dinb(n647), .dout(n649));
  jxor g0349(.dina(n649), .dinb(G490), .dout(n650));
  jand g0350(.dina(n650), .dinb(n646), .dout(n651));
  jand g0351(.dina(n651), .dinb(n642), .dout(n652));
  jand g0352(.dina(n652), .dinb(n633), .dout(G615));
  jxor g0353(.dina(G316), .dinb(G308), .dout(n654));
  jxor g0354(.dina(G351), .dinb(G341), .dout(n655));
  jxor g0355(.dina(n655), .dinb(n654), .dout(n656));
  jxor g0356(.dina(G369), .dinb(G361), .dout(n657));
  jxor g0357(.dina(n657), .dinb(n424), .dout(n658));
  jxor g0358(.dina(G302), .dinb(n398), .dout(n659));
  jxor g0359(.dina(n659), .dinb(n658), .dout(n660));
  jxor g0360(.dina(n660), .dinb(n656), .dout(n661));
  jnot g0361(.din(n661), .dout(G1002));
  jxor g0362(.dina(G226), .dinb(G218), .dout(n663));
  jxor g0363(.dina(G273), .dinb(G265), .dout(n664));
  jxor g0364(.dina(n664), .dinb(n663), .dout(n665));
  jxor g0365(.dina(G289), .dinb(G281), .dout(n666));
  jxor g0366(.dina(G257), .dinb(G234), .dout(n667));
  jxor g0367(.dina(n667), .dinb(n666), .dout(n668));
  jxor g0368(.dina(G210), .dinb(n518), .dout(n669));
  jxor g0369(.dina(n669), .dinb(n668), .dout(n670));
  jxor g0370(.dina(n670), .dinb(n665), .dout(n671));
  jnot g0371(.din(n671), .dout(G1004));
  jnot g0372(.din(n560), .dout(n673));
  jand g0373(.dina(n673), .dinb(n462), .dout(n674));
  jnot g0374(.din(n674), .dout(n675));
  jand g0375(.dina(n560), .dinb(G435), .dout(n676));
  jnot g0376(.din(n577), .dout(n677));
  jand g0377(.dina(n677), .dinb(n473), .dout(n678));
  jor  g0378(.dina(n677), .dinb(n473), .dout(n679));
  jand g0379(.dina(n582), .dinb(n451), .dout(n680));
  jor  g0380(.dina(n566), .dinb(n497), .dout(n681));
  jor  g0381(.dina(n571), .dinb(n681), .dout(n682));
  jnot g0382(.din(G280), .dout(n683));
  jand g0383(.dina(G335), .dinb(n683), .dout(n684));
  jnot g0384(.din(n569), .dout(n685));
  jor  g0385(.dina(n685), .dinb(n684), .dout(n686));
  jor  g0386(.dina(n686), .dinb(n486), .dout(n687));
  jor  g0387(.dina(n582), .dinb(n451), .dout(n688));
  jand g0388(.dina(n688), .dinb(n687), .dout(n689));
  jand g0389(.dina(n689), .dinb(n682), .dout(n690));
  jor  g0390(.dina(n690), .dinb(n680), .dout(n691));
  jand g0391(.dina(n691), .dinb(n679), .dout(n692));
  jor  g0392(.dina(n692), .dinb(n678), .dout(n693));
  jnot g0393(.din(n693), .dout(n694));
  jor  g0394(.dina(n694), .dinb(n676), .dout(n695));
  jand g0395(.dina(n695), .dinb(n675), .dout(n696));
  jand g0396(.dina(n696), .dinb(n607), .dout(n697));
  jand g0397(.dina(n595), .dinb(G446), .dout(n698));
  jor  g0398(.dina(n595), .dinb(G446), .dout(n699));
  jor  g0399(.dina(n590), .dinb(G457), .dout(n700));
  jand g0400(.dina(n590), .dinb(G457), .dout(n701));
  jand g0401(.dina(n604), .dinb(G468), .dout(n702));
  jand g0402(.dina(n600), .dinb(G422), .dout(n703));
  jand g0403(.dina(n605), .dinb(n703), .dout(n704));
  jor  g0404(.dina(n704), .dinb(n702), .dout(n705));
  jor  g0405(.dina(n705), .dinb(n701), .dout(n706));
  jand g0406(.dina(n706), .dinb(n700), .dout(n707));
  jand g0407(.dina(n707), .dinb(n699), .dout(n708));
  jor  g0408(.dina(n708), .dinb(n698), .dout(n709));
  jor  g0409(.dina(n709), .dinb(n697), .dout(G591));
  jand g0410(.dina(n613), .dinb(G503), .dout(n711));
  jor  g0411(.dina(n624), .dinb(n410), .dout(n712));
  jand g0412(.dina(n624), .dinb(n410), .dout(n713));
  jand g0413(.dina(G599), .dinb(G332), .dout(n714));
  jand g0414(.dina(n435), .dinb(n609), .dout(n715));
  jor  g0415(.dina(n715), .dinb(n714), .dout(n716));
  jand g0416(.dina(n716), .dinb(n437), .dout(n717));
  jand g0417(.dina(G612), .dinb(G332), .dout(n718));
  jand g0418(.dina(n385), .dinb(n609), .dout(n719));
  jor  g0419(.dina(n719), .dinb(n718), .dout(n720));
  jand g0420(.dina(n720), .dinb(n388), .dout(n721));
  jor  g0421(.dina(n621), .dinb(n721), .dout(n722));
  jor  g0422(.dina(n720), .dinb(n388), .dout(n723));
  jor  g0423(.dina(n716), .dinb(n437), .dout(n724));
  jand g0424(.dina(n724), .dinb(n723), .dout(n725));
  jand g0425(.dina(n725), .dinb(n722), .dout(n726));
  jor  g0426(.dina(n726), .dinb(n717), .dout(n727));
  jor  g0427(.dina(n727), .dinb(n713), .dout(n728));
  jand g0428(.dina(n728), .dinb(n712), .dout(n729));
  jnot g0429(.din(n729), .dout(n730));
  jand g0430(.dina(n730), .dinb(n614), .dout(n731));
  jor  g0431(.dina(n731), .dinb(n711), .dout(n732));
  jand g0432(.dina(n732), .dinb(n651), .dout(n733));
  jnot g0433(.din(n642), .dout(n734));
  jnot g0434(.din(n645), .dout(n735));
  jand g0435(.dina(n735), .dinb(n362), .dout(n736));
  jnot g0436(.din(n736), .dout(n737));
  jand g0437(.dina(n645), .dinb(G479), .dout(n738));
  jand g0438(.dina(n649), .dinb(G490), .dout(n739));
  jor  g0439(.dina(n739), .dinb(n738), .dout(n740));
  jand g0440(.dina(n740), .dinb(n737), .dout(n741));
  jor  g0441(.dina(n741), .dinb(n734), .dout(n742));
  jor  g0442(.dina(n742), .dinb(n733), .dout(G618));
  jnot g0443(.din(G54), .dout(n744));
  jxor g0444(.dina(n621), .dinb(n744), .dout(n745));
  jnot g0445(.din(G4092), .dout(n746));
  jand g0446(.dina(n746), .dinb(G4091), .dout(n747));
  jnot g0447(.din(n747), .dout(n748));
  jor  g0448(.dina(n748), .dinb(n745), .dout(n749));
  jnot g0449(.din(G4091), .dout(n750));
  jand g0450(.dina(n746), .dinb(n750), .dout(n751));
  jand g0451(.dina(n751), .dinb(n419), .dout(n752));
  jand g0452(.dina(G4092), .dinb(n750), .dout(n753));
  jand g0453(.dina(n753), .dinb(G131), .dout(n754));
  jor  g0454(.dina(n754), .dinb(n752), .dout(n755));
  jnot g0455(.din(n755), .dout(n756));
  jand g0456(.dina(n756), .dinb(n749), .dout(G822));
  jnot g0457(.din(n618), .dout(n758));
  jand g0458(.dina(n621), .dinb(n744), .dout(n759));
  jnot g0459(.din(n759), .dout(n760));
  jand g0460(.dina(n760), .dinb(n758), .dout(n761));
  jand g0461(.dina(n759), .dinb(n618), .dout(n762));
  jor  g0462(.dina(n762), .dinb(n748), .dout(n763));
  jor  g0463(.dina(n763), .dinb(n761), .dout(n764));
  jnot g0464(.din(n751), .dout(n765));
  jor  g0465(.dina(n765), .dinb(n397), .dout(n766));
  jand g0466(.dina(n753), .dinb(G129), .dout(n767));
  jnot g0467(.din(n767), .dout(n768));
  jand g0468(.dina(n768), .dinb(n766), .dout(n769));
  jand g0469(.dina(n769), .dinb(n764), .dout(G838));
  jxor g0470(.dina(n567), .dinb(G4), .dout(n771));
  jand g0471(.dina(n771), .dinb(n747), .dout(n772));
  jnot g0472(.din(n772), .dout(n773));
  jor  g0473(.dina(n765), .dinb(n505), .dout(n774));
  jand g0474(.dina(n753), .dinb(G117), .dout(n775));
  jnot g0475(.din(n775), .dout(n776));
  jand g0476(.dina(n776), .dinb(n774), .dout(n777));
  jand g0477(.dina(n777), .dinb(n773), .dout(G861));
  jnot g0478(.din(n636), .dout(n779));
  jand g0479(.dina(n633), .dinb(G54), .dout(n780));
  jor  g0480(.dina(n780), .dinb(n732), .dout(n781));
  jand g0481(.dina(n781), .dinb(n651), .dout(n782));
  jor  g0482(.dina(n782), .dinb(n741), .dout(n783));
  jnot g0483(.din(n783), .dout(n784));
  jor  g0484(.dina(n784), .dinb(n779), .dout(n785));
  jxor g0485(.dina(n640), .dinb(n779), .dout(n786));
  jnot g0486(.din(n786), .dout(n787));
  jor  g0487(.dina(n787), .dinb(n783), .dout(n788));
  jand g0488(.dina(n788), .dinb(n785), .dout(n789));
  jnot g0489(.din(n789), .dout(G623));
  jnot g0490(.din(G861), .dout(n791));
  jnot g0491(.din(G4087), .dout(n792));
  jand g0492(.dina(G4088), .dinb(n792), .dout(n793));
  jand g0493(.dina(n793), .dinb(n791), .dout(n794));
  jnot g0494(.din(G822), .dout(n795));
  jnot g0495(.din(G4088), .dout(n796));
  jand g0496(.dina(n796), .dinb(n792), .dout(n797));
  jand g0497(.dina(n797), .dinb(n795), .dout(n798));
  jand g0498(.dina(n796), .dinb(G4087), .dout(n799));
  jand g0499(.dina(n799), .dinb(G11), .dout(n800));
  jand g0500(.dina(G4088), .dinb(G4087), .dout(n801));
  jand g0501(.dina(n801), .dinb(G61), .dout(n802));
  jor  g0502(.dina(n802), .dinb(n800), .dout(n803));
  jor  g0503(.dina(n803), .dinb(n798), .dout(n804));
  jor  g0504(.dina(n804), .dinb(n794), .dout(G722));
  jand g0505(.dina(n729), .dinb(n631), .dout(n806));
  jand g0506(.dina(n729), .dinb(n744), .dout(n807));
  jor  g0507(.dina(n807), .dinb(n806), .dout(n808));
  jxor g0508(.dina(n808), .dinb(n614), .dout(n809));
  jor  g0509(.dina(n809), .dinb(n748), .dout(n810));
  jor  g0510(.dina(n765), .dinb(n434), .dout(n811));
  jand g0511(.dina(n753), .dinb(G52), .dout(n812));
  jnot g0512(.din(n812), .dout(n813));
  jand g0513(.dina(n813), .dinb(n811), .dout(n814));
  jand g0514(.dina(n814), .dinb(n810), .dout(G832));
  jnot g0515(.din(n625), .dout(n816));
  jand g0516(.dina(n727), .dinb(n744), .dout(n817));
  jand g0517(.dina(n726), .dinb(n623), .dout(n818));
  jor  g0518(.dina(n818), .dinb(n717), .dout(n819));
  jor  g0519(.dina(n819), .dinb(n817), .dout(n820));
  jxor g0520(.dina(n820), .dinb(n816), .dout(n821));
  jor  g0521(.dina(n821), .dinb(n748), .dout(n822));
  jand g0522(.dina(n751), .dinb(n414), .dout(n823));
  jand g0523(.dina(n753), .dinb(G130), .dout(n824));
  jor  g0524(.dina(n824), .dinb(n823), .dout(n825));
  jnot g0525(.din(n825), .dout(n826));
  jand g0526(.dina(n826), .dinb(n822), .dout(G834));
  jor  g0527(.dina(n617), .dinb(G534), .dout(n828));
  jand g0528(.dina(n617), .dinb(G534), .dout(n829));
  jor  g0529(.dina(n760), .dinb(n829), .dout(n830));
  jand g0530(.dina(n830), .dinb(n828), .dout(n831));
  jxor g0531(.dina(n831), .dinb(n629), .dout(n832));
  jor  g0532(.dina(n832), .dinb(n748), .dout(n833));
  jor  g0533(.dina(n765), .dinb(n445), .dout(n834));
  jand g0534(.dina(n753), .dinb(G119), .dout(n835));
  jnot g0535(.din(n835), .dout(n836));
  jand g0536(.dina(n836), .dinb(n834), .dout(n837));
  jand g0537(.dina(n837), .dinb(n833), .dout(G836));
  jnot g0538(.din(G4090), .dout(n839));
  jand g0539(.dina(n839), .dinb(G4089), .dout(n840));
  jand g0540(.dina(n840), .dinb(n791), .dout(n841));
  jnot g0541(.din(G4089), .dout(n842));
  jand g0542(.dina(n839), .dinb(n842), .dout(n843));
  jand g0543(.dina(n843), .dinb(n795), .dout(n844));
  jand g0544(.dina(G4090), .dinb(n842), .dout(n845));
  jand g0545(.dina(n845), .dinb(G11), .dout(n846));
  jand g0546(.dina(G4090), .dinb(G4089), .dout(n847));
  jand g0547(.dina(n847), .dinb(G61), .dout(n848));
  jor  g0548(.dina(n848), .dinb(n846), .dout(n849));
  jor  g0549(.dina(n849), .dinb(n844), .dout(n850));
  jor  g0550(.dina(n850), .dinb(n841), .dout(G859));
  jnot g0551(.din(n678), .dout(n852));
  jnot g0552(.din(n679), .dout(n853));
  jor  g0553(.dina(n583), .dinb(n574), .dout(n854));
  jand g0554(.dina(n854), .dinb(n691), .dout(n855));
  jnot g0555(.din(n855), .dout(n856));
  jnot g0556(.din(n691), .dout(n857));
  jor  g0557(.dina(n857), .dinb(G4), .dout(n858));
  jand g0558(.dina(n858), .dinb(n856), .dout(n859));
  jor  g0559(.dina(n859), .dinb(n853), .dout(n860));
  jand g0560(.dina(n860), .dinb(n852), .dout(n861));
  jxor g0561(.dina(n861), .dinb(n562), .dout(n862));
  jor  g0562(.dina(n862), .dinb(n748), .dout(n863));
  jor  g0563(.dina(n765), .dinb(n470), .dout(n864));
  jand g0564(.dina(n753), .dinb(G122), .dout(n865));
  jnot g0565(.din(n865), .dout(n866));
  jand g0566(.dina(n866), .dinb(n864), .dout(n867));
  jand g0567(.dina(n867), .dinb(n863), .dout(G871));
  jxor g0568(.dina(n859), .dinb(n578), .dout(n869));
  jor  g0569(.dina(n869), .dinb(n748), .dout(n870));
  jor  g0570(.dina(n765), .dinb(n481), .dout(n871));
  jand g0571(.dina(n753), .dinb(G128), .dout(n872));
  jnot g0572(.din(n872), .dout(n873));
  jand g0573(.dina(n873), .dinb(n871), .dout(n874));
  jand g0574(.dina(n874), .dinb(n870), .dout(G873));
  jand g0575(.dina(n567), .dinb(G4), .dout(n876));
  jnot g0576(.din(n876), .dout(n877));
  jand g0577(.dina(n877), .dinb(n681), .dout(n878));
  jor  g0578(.dina(n878), .dinb(n571), .dout(n879));
  jand g0579(.dina(n879), .dinb(n687), .dout(n880));
  jxor g0580(.dina(n880), .dinb(n583), .dout(n881));
  jand g0581(.dina(n881), .dinb(n747), .dout(n882));
  jnot g0582(.din(n882), .dout(n883));
  jor  g0583(.dina(n765), .dinb(n459), .dout(n884));
  jand g0584(.dina(n753), .dinb(G127), .dout(n885));
  jnot g0585(.din(n885), .dout(n886));
  jand g0586(.dina(n886), .dinb(n884), .dout(n887));
  jand g0587(.dina(n887), .dinb(n883), .dout(G875));
  jand g0588(.dina(n571), .dinb(n681), .dout(n889));
  jand g0589(.dina(n889), .dinb(n877), .dout(n890));
  jnot g0590(.din(n890), .dout(n891));
  jand g0591(.dina(n891), .dinb(n879), .dout(n892));
  jand g0592(.dina(n892), .dinb(n747), .dout(n893));
  jnot g0593(.din(n893), .dout(n894));
  jor  g0594(.dina(n765), .dinb(n494), .dout(n895));
  jand g0595(.dina(n753), .dinb(G126), .dout(n896));
  jnot g0596(.din(n896), .dout(n897));
  jand g0597(.dina(n897), .dinb(n895), .dout(n898));
  jand g0598(.dina(n898), .dinb(n894), .dout(G877));
  jxor g0599(.dina(n649), .dinb(n735), .dout(n900));
  jxor g0600(.dina(n900), .dinb(n786), .dout(n901));
  jxor g0601(.dina(n901), .dinb(n621), .dout(n902));
  jand g0602(.dina(G369), .dinb(n609), .dout(n903));
  jand g0603(.dina(G372), .dinb(G332), .dout(n904));
  jor  g0604(.dina(n904), .dinb(n903), .dout(n905));
  jxor g0605(.dina(n905), .dinb(n617), .dout(n906));
  jxor g0606(.dina(n906), .dinb(n628), .dout(n907));
  jnot g0607(.din(G331), .dout(n908));
  jand g0608(.dina(n624), .dinb(n908), .dout(n909));
  jnot g0609(.din(n624), .dout(n910));
  jand g0610(.dina(n910), .dinb(n613), .dout(n911));
  jor  g0611(.dina(n911), .dinb(n909), .dout(n912));
  jxor g0612(.dina(n912), .dinb(n907), .dout(n913));
  jxor g0613(.dina(n913), .dinb(n902), .dout(n914));
  jnot g0614(.din(n914), .dout(G998));
  jxor g0615(.dina(n577), .dinb(n566), .dout(n916));
  jxor g0616(.dina(n582), .dinb(n570), .dout(n917));
  jxor g0617(.dina(n917), .dinb(n916), .dout(n918));
  jxor g0618(.dina(n918), .dinb(n590), .dout(n919));
  jand g0619(.dina(n556), .dinb(G289), .dout(n920));
  jand g0620(.dina(G335), .dinb(G292), .dout(n921));
  jor  g0621(.dina(n921), .dinb(n920), .dout(n922));
  jxor g0622(.dina(n922), .dinb(n600), .dout(n923));
  jxor g0623(.dina(n923), .dinb(n560), .dout(n924));
  jxor g0624(.dina(n604), .dinb(n595), .dout(n925));
  jxor g0625(.dina(n925), .dinb(n924), .dout(n926));
  jxor g0626(.dina(n926), .dinb(n919), .dout(G1000));
  jnot g0627(.din(n596), .dout(n928));
  jnot g0628(.din(n707), .dout(n929));
  jnot g0629(.din(n700), .dout(n930));
  jnot g0630(.din(n605), .dout(n931));
  jnot g0631(.din(n601), .dout(n932));
  jnot g0632(.din(n696), .dout(n933));
  jand g0633(.dina(n587), .dinb(G4), .dout(n934));
  jnot g0634(.din(n934), .dout(n935));
  jand g0635(.dina(n935), .dinb(n933), .dout(n936));
  jor  g0636(.dina(n936), .dinb(n932), .dout(n937));
  jor  g0637(.dina(n937), .dinb(n931), .dout(n938));
  jor  g0638(.dina(n938), .dinb(n930), .dout(n939));
  jand g0639(.dina(n939), .dinb(n929), .dout(n940));
  jxor g0640(.dina(n940), .dinb(n928), .dout(n941));
  jnot g0641(.din(n941), .dout(n942));
  jnot g0642(.din(n591), .dout(n943));
  jnot g0643(.din(n705), .dout(n944));
  jand g0644(.dina(n938), .dinb(n944), .dout(n945));
  jxor g0645(.dina(n945), .dinb(n943), .dout(n946));
  jnot g0646(.din(n946), .dout(n947));
  jor  g0647(.dina(n600), .dinb(G422), .dout(n948));
  jnot g0648(.din(n948), .dout(n949));
  jnot g0649(.din(n703), .dout(n950));
  jand g0650(.dina(n936), .dinb(n950), .dout(n951));
  jor  g0651(.dina(n951), .dinb(n949), .dout(n952));
  jxor g0652(.dina(n952), .dinb(n605), .dout(n953));
  jxor g0653(.dina(n936), .dinb(n932), .dout(n954));
  jnot g0654(.din(n954), .dout(n955));
  jnot g0655(.din(n881), .dout(n956));
  jnot g0656(.din(n771), .dout(n957));
  jnot g0657(.din(n892), .dout(n958));
  jand g0658(.dina(n958), .dinb(n957), .dout(n959));
  jand g0659(.dina(n959), .dinb(n956), .dout(n960));
  jand g0660(.dina(n960), .dinb(n869), .dout(n961));
  jand g0661(.dina(n961), .dinb(n862), .dout(n962));
  jand g0662(.dina(n962), .dinb(n955), .dout(n963));
  jand g0663(.dina(n963), .dinb(n953), .dout(n964));
  jand g0664(.dina(n964), .dinb(n947), .dout(n965));
  jand g0665(.dina(n965), .dinb(n942), .dout(G575));
  jnot g0666(.din(n646), .dout(n967));
  jor  g0667(.dina(n649), .dinb(G490), .dout(n968));
  jor  g0668(.dina(n781), .dinb(n739), .dout(n969));
  jand g0669(.dina(n969), .dinb(n968), .dout(n970));
  jxor g0670(.dina(n970), .dinb(n967), .dout(n971));
  jxor g0671(.dina(n783), .dinb(n640), .dout(n972));
  jxor g0672(.dina(n781), .dinb(n650), .dout(n973));
  jnot g0673(.din(n973), .dout(n974));
  jor  g0674(.dina(n621), .dinb(n744), .dout(n975));
  jand g0675(.dina(n975), .dinb(n636), .dout(n976));
  jand g0676(.dina(n976), .dinb(n761), .dout(n977));
  jand g0677(.dina(n977), .dinb(n832), .dout(n978));
  jand g0678(.dina(n978), .dinb(n821), .dout(n979));
  jand g0679(.dina(n979), .dinb(n809), .dout(n980));
  jand g0680(.dina(n980), .dinb(n974), .dout(n981));
  jand g0681(.dina(n981), .dinb(n972), .dout(n982));
  jand g0682(.dina(n982), .dinb(n971), .dout(G585));
  jnot g0683(.din(G1690), .dout(n984));
  jand g0684(.dina(n984), .dinb(G1689), .dout(n985));
  jand g0685(.dina(n985), .dinb(n791), .dout(n986));
  jnot g0686(.din(G1689), .dout(n987));
  jand g0687(.dina(n984), .dinb(n987), .dout(n988));
  jand g0688(.dina(n988), .dinb(n795), .dout(n989));
  jand g0689(.dina(G1690), .dinb(n987), .dout(n990));
  jand g0690(.dina(n990), .dinb(G182), .dout(n991));
  jand g0691(.dina(G1690), .dinb(G1689), .dout(n992));
  jand g0692(.dina(n992), .dinb(G185), .dout(n993));
  jor  g0693(.dina(n993), .dinb(n991), .dout(n994));
  jor  g0694(.dina(n994), .dinb(n989), .dout(n995));
  jor  g0695(.dina(n995), .dinb(n986), .dout(n996));
  jand g0696(.dina(n996), .dinb(G137), .dout(G661));
  jnot g0697(.din(G1694), .dout(n998));
  jand g0698(.dina(n998), .dinb(G1691), .dout(n999));
  jand g0699(.dina(n999), .dinb(n791), .dout(n1000));
  jnot g0700(.din(G1691), .dout(n1001));
  jand g0701(.dina(n998), .dinb(n1001), .dout(n1002));
  jand g0702(.dina(n1002), .dinb(n795), .dout(n1003));
  jand g0703(.dina(G1694), .dinb(n1001), .dout(n1004));
  jand g0704(.dina(n1004), .dinb(G182), .dout(n1005));
  jand g0705(.dina(G1694), .dinb(G1691), .dout(n1006));
  jand g0706(.dina(n1006), .dinb(G185), .dout(n1007));
  jor  g0707(.dina(n1007), .dinb(n1005), .dout(n1008));
  jor  g0708(.dina(n1008), .dinb(n1003), .dout(n1009));
  jor  g0709(.dina(n1009), .dinb(n1000), .dout(n1010));
  jand g0710(.dina(n1010), .dinb(G137), .dout(G693));
  jnot g0711(.din(G871), .dout(n1012));
  jand g0712(.dina(n1012), .dinb(n793), .dout(n1013));
  jnot g0713(.din(G832), .dout(n1014));
  jand g0714(.dina(n1014), .dinb(n797), .dout(n1015));
  jand g0715(.dina(n799), .dinb(G43), .dout(n1016));
  jand g0716(.dina(n801), .dinb(G37), .dout(n1017));
  jor  g0717(.dina(n1017), .dinb(n1016), .dout(n1018));
  jor  g0718(.dina(n1018), .dinb(n1015), .dout(n1019));
  jor  g0719(.dina(n1019), .dinb(n1013), .dout(G747));
  jnot g0720(.din(G873), .dout(n1021));
  jand g0721(.dina(n1021), .dinb(n793), .dout(n1022));
  jnot g0722(.din(G834), .dout(n1023));
  jand g0723(.dina(n1023), .dinb(n797), .dout(n1024));
  jand g0724(.dina(n799), .dinb(G76), .dout(n1025));
  jand g0725(.dina(n801), .dinb(G20), .dout(n1026));
  jor  g0726(.dina(n1026), .dinb(n1025), .dout(n1027));
  jor  g0727(.dina(n1027), .dinb(n1024), .dout(n1028));
  jor  g0728(.dina(n1028), .dinb(n1022), .dout(G752));
  jnot g0729(.din(G875), .dout(n1030));
  jand g0730(.dina(n1030), .dinb(n793), .dout(n1031));
  jnot g0731(.din(G836), .dout(n1032));
  jand g0732(.dina(n1032), .dinb(n797), .dout(n1033));
  jand g0733(.dina(n799), .dinb(G73), .dout(n1034));
  jand g0734(.dina(n801), .dinb(G17), .dout(n1035));
  jor  g0735(.dina(n1035), .dinb(n1034), .dout(n1036));
  jor  g0736(.dina(n1036), .dinb(n1033), .dout(n1037));
  jor  g0737(.dina(n1037), .dinb(n1031), .dout(G757));
  jnot g0738(.din(G877), .dout(n1039));
  jand g0739(.dina(n1039), .dinb(n793), .dout(n1040));
  jnot g0740(.din(G838), .dout(n1041));
  jand g0741(.dina(n797), .dinb(n1041), .dout(n1042));
  jand g0742(.dina(n799), .dinb(G67), .dout(n1043));
  jand g0743(.dina(n801), .dinb(G70), .dout(n1044));
  jor  g0744(.dina(n1044), .dinb(n1043), .dout(n1045));
  jor  g0745(.dina(n1045), .dinb(n1042), .dout(n1046));
  jor  g0746(.dina(n1046), .dinb(n1040), .dout(G762));
  jand g0747(.dina(n1012), .dinb(n840), .dout(n1048));
  jand g0748(.dina(n843), .dinb(n1014), .dout(n1049));
  jand g0749(.dina(n845), .dinb(G43), .dout(n1050));
  jand g0750(.dina(n847), .dinb(G37), .dout(n1051));
  jor  g0751(.dina(n1051), .dinb(n1050), .dout(n1052));
  jor  g0752(.dina(n1052), .dinb(n1049), .dout(n1053));
  jor  g0753(.dina(n1053), .dinb(n1048), .dout(G787));
  jand g0754(.dina(n1021), .dinb(n840), .dout(n1055));
  jand g0755(.dina(n843), .dinb(n1023), .dout(n1056));
  jand g0756(.dina(n845), .dinb(G76), .dout(n1057));
  jand g0757(.dina(n847), .dinb(G20), .dout(n1058));
  jor  g0758(.dina(n1058), .dinb(n1057), .dout(n1059));
  jor  g0759(.dina(n1059), .dinb(n1056), .dout(n1060));
  jor  g0760(.dina(n1060), .dinb(n1055), .dout(G792));
  jand g0761(.dina(n1030), .dinb(n840), .dout(n1062));
  jand g0762(.dina(n843), .dinb(n1032), .dout(n1063));
  jand g0763(.dina(n845), .dinb(G73), .dout(n1064));
  jand g0764(.dina(n847), .dinb(G17), .dout(n1065));
  jor  g0765(.dina(n1065), .dinb(n1064), .dout(n1066));
  jor  g0766(.dina(n1066), .dinb(n1063), .dout(n1067));
  jor  g0767(.dina(n1067), .dinb(n1062), .dout(G797));
  jand g0768(.dina(n1039), .dinb(n840), .dout(n1069));
  jand g0769(.dina(n843), .dinb(n1041), .dout(n1070));
  jand g0770(.dina(n845), .dinb(G67), .dout(n1071));
  jand g0771(.dina(n847), .dinb(G70), .dout(n1072));
  jor  g0772(.dina(n1072), .dinb(n1071), .dout(n1073));
  jor  g0773(.dina(n1073), .dinb(n1070), .dout(n1074));
  jor  g0774(.dina(n1074), .dinb(n1069), .dout(G802));
  jand g0775(.dina(n985), .dinb(n1012), .dout(n1076));
  jand g0776(.dina(n988), .dinb(n1014), .dout(n1077));
  jand g0777(.dina(n990), .dinb(G200), .dout(n1078));
  jand g0778(.dina(n992), .dinb(G170), .dout(n1079));
  jor  g0779(.dina(n1079), .dinb(n1078), .dout(n1080));
  jor  g0780(.dina(n1080), .dinb(n1077), .dout(n1081));
  jor  g0781(.dina(n1081), .dinb(n1076), .dout(n1082));
  jand g0782(.dina(n1082), .dinb(G137), .dout(G642));
  jand g0783(.dina(n985), .dinb(n1039), .dout(n1084));
  jand g0784(.dina(n988), .dinb(n1041), .dout(n1085));
  jand g0785(.dina(n990), .dinb(G188), .dout(n1086));
  jand g0786(.dina(n992), .dinb(G158), .dout(n1087));
  jor  g0787(.dina(n1087), .dinb(n1086), .dout(n1088));
  jor  g0788(.dina(n1088), .dinb(n1085), .dout(n1089));
  jor  g0789(.dina(n1089), .dinb(n1084), .dout(n1090));
  jand g0790(.dina(n1090), .dinb(G137), .dout(G664));
  jand g0791(.dina(n985), .dinb(n1030), .dout(n1092));
  jand g0792(.dina(n988), .dinb(n1032), .dout(n1093));
  jand g0793(.dina(n990), .dinb(G155), .dout(n1094));
  jand g0794(.dina(n992), .dinb(G152), .dout(n1095));
  jor  g0795(.dina(n1095), .dinb(n1094), .dout(n1096));
  jor  g0796(.dina(n1096), .dinb(n1093), .dout(n1097));
  jor  g0797(.dina(n1097), .dinb(n1092), .dout(n1098));
  jand g0798(.dina(n1098), .dinb(G137), .dout(G667));
  jand g0799(.dina(n985), .dinb(n1021), .dout(n1100));
  jand g0800(.dina(n988), .dinb(n1023), .dout(n1101));
  jand g0801(.dina(n990), .dinb(G149), .dout(n1102));
  jand g0802(.dina(n992), .dinb(G146), .dout(n1103));
  jor  g0803(.dina(n1103), .dinb(n1102), .dout(n1104));
  jor  g0804(.dina(n1104), .dinb(n1101), .dout(n1105));
  jor  g0805(.dina(n1105), .dinb(n1100), .dout(n1106));
  jand g0806(.dina(n1106), .dinb(G137), .dout(G670));
  jand g0807(.dina(n999), .dinb(n1012), .dout(n1108));
  jand g0808(.dina(n1002), .dinb(n1014), .dout(n1109));
  jand g0809(.dina(n1004), .dinb(G200), .dout(n1110));
  jand g0810(.dina(n1006), .dinb(G170), .dout(n1111));
  jor  g0811(.dina(n1111), .dinb(n1110), .dout(n1112));
  jor  g0812(.dina(n1112), .dinb(n1109), .dout(n1113));
  jor  g0813(.dina(n1113), .dinb(n1108), .dout(n1114));
  jand g0814(.dina(n1114), .dinb(G137), .dout(G676));
  jand g0815(.dina(n999), .dinb(n1039), .dout(n1116));
  jand g0816(.dina(n1002), .dinb(n1041), .dout(n1117));
  jand g0817(.dina(n1004), .dinb(G188), .dout(n1118));
  jand g0818(.dina(n1006), .dinb(G158), .dout(n1119));
  jor  g0819(.dina(n1119), .dinb(n1118), .dout(n1120));
  jor  g0820(.dina(n1120), .dinb(n1117), .dout(n1121));
  jor  g0821(.dina(n1121), .dinb(n1116), .dout(n1122));
  jand g0822(.dina(n1122), .dinb(G137), .dout(G696));
  jand g0823(.dina(n999), .dinb(n1030), .dout(n1124));
  jand g0824(.dina(n1002), .dinb(n1032), .dout(n1125));
  jand g0825(.dina(n1004), .dinb(G155), .dout(n1126));
  jand g0826(.dina(n1006), .dinb(G152), .dout(n1127));
  jor  g0827(.dina(n1127), .dinb(n1126), .dout(n1128));
  jor  g0828(.dina(n1128), .dinb(n1125), .dout(n1129));
  jor  g0829(.dina(n1129), .dinb(n1124), .dout(n1130));
  jand g0830(.dina(n1130), .dinb(G137), .dout(G699));
  jand g0831(.dina(n999), .dinb(n1021), .dout(n1132));
  jand g0832(.dina(n1002), .dinb(n1023), .dout(n1133));
  jand g0833(.dina(n1004), .dinb(G149), .dout(n1134));
  jand g0834(.dina(n1006), .dinb(G146), .dout(n1135));
  jor  g0835(.dina(n1135), .dinb(n1134), .dout(n1136));
  jor  g0836(.dina(n1136), .dinb(n1133), .dout(n1137));
  jor  g0837(.dina(n1137), .dinb(n1132), .dout(n1138));
  jand g0838(.dina(n1138), .dinb(G137), .dout(G702));
  jand g0839(.dina(n789), .dinb(G3724), .dout(n1140));
  jnot g0840(.din(G3717), .dout(n1141));
  jnot g0841(.din(G3724), .dout(n1142));
  jand g0842(.dina(n1142), .dinb(G123), .dout(n1143));
  jor  g0843(.dina(n1143), .dinb(n1141), .dout(n1144));
  jor  g0844(.dina(n1144), .dinb(n1140), .dout(n1145));
  jnot g0845(.din(G135), .dout(n1146));
  jnot g0846(.din(G4115), .dout(n1147));
  jor  g0847(.dina(n1147), .dinb(n1146), .dout(n1148));
  jxor g0848(.dina(n636), .dinb(G132), .dout(n1149));
  jand g0849(.dina(n1149), .dinb(G3724), .dout(n1150));
  jnot g0850(.din(n401), .dout(n1151));
  jand g0851(.dina(n1151), .dinb(n1142), .dout(n1152));
  jor  g0852(.dina(n1152), .dinb(G3717), .dout(n1153));
  jor  g0853(.dina(n1153), .dinb(n1150), .dout(n1154));
  jand g0854(.dina(n1154), .dinb(n1148), .dout(n1155));
  jand g0855(.dina(n1155), .dinb(n1145), .dout(G818));
  jor  g0856(.dina(n783), .dinb(n640), .dout(n1157));
  jxor g0857(.dina(n1157), .dinb(G132), .dout(G813));
  jand g0858(.dina(n789), .dinb(n747), .dout(n1159));
  jand g0859(.dina(n753), .dinb(G123), .dout(n1160));
  jand g0860(.dina(n751), .dinb(n1151), .dout(n1161));
  jor  g0861(.dina(n1161), .dinb(n1160), .dout(n1162));
  jor  g0862(.dina(n1162), .dinb(n1159), .dout(n1163));
  jnot g0863(.din(n1163), .dout(G824));
  jor  g0864(.dina(n972), .dinb(n748), .dout(n1165));
  jand g0865(.dina(n751), .dinb(n407), .dout(n1166));
  jand g0866(.dina(n753), .dinb(G121), .dout(n1167));
  jor  g0867(.dina(n1167), .dinb(n1166), .dout(n1168));
  jnot g0868(.din(n1168), .dout(n1169));
  jand g0869(.dina(n1169), .dinb(n1165), .dout(G826));
  jor  g0870(.dina(n971), .dinb(n748), .dout(n1171));
  jor  g0871(.dina(n765), .dinb(n372), .dout(n1172));
  jand g0872(.dina(n753), .dinb(G116), .dout(n1173));
  jnot g0873(.din(n1173), .dout(n1174));
  jand g0874(.dina(n1174), .dinb(n1172), .dout(n1175));
  jand g0875(.dina(n1175), .dinb(n1171), .dout(G828));
  jand g0876(.dina(n973), .dinb(n747), .dout(n1177));
  jnot g0877(.din(n1177), .dout(n1178));
  jor  g0878(.dina(n765), .dinb(n383), .dout(n1179));
  jand g0879(.dina(n753), .dinb(G112), .dout(n1180));
  jnot g0880(.din(n1180), .dout(n1181));
  jand g0881(.dina(n1181), .dinb(n1179), .dout(n1182));
  jand g0882(.dina(n1182), .dinb(n1178), .dout(G830));
  jnot g0883(.din(G1000), .dout(n1184));
  jand g0884(.dina(G559), .dinb(G245), .dout(n1185));
  jand g0885(.dina(n1185), .dinb(n318), .dout(n1186));
  jand g0886(.dina(n1186), .dinb(G601), .dout(n1187));
  jand g0887(.dina(n1187), .dinb(n661), .dout(n1188));
  jand g0888(.dina(n1188), .dinb(n671), .dout(n1189));
  jand g0889(.dina(n1189), .dinb(n914), .dout(n1190));
  jand g0890(.dina(n1190), .dinb(n1184), .dout(G854));
  jand g0891(.dina(n941), .dinb(n747), .dout(n1192));
  jnot g0892(.din(n528), .dout(n1193));
  jand g0893(.dina(n751), .dinb(n1193), .dout(n1194));
  jand g0894(.dina(n753), .dinb(G115), .dout(n1195));
  jor  g0895(.dina(n1195), .dinb(n1194), .dout(n1196));
  jor  g0896(.dina(n1196), .dinb(n1192), .dout(n1197));
  jnot g0897(.din(n1197), .dout(G863));
  jand g0898(.dina(n946), .dinb(n747), .dout(n1199));
  jor  g0899(.dina(n765), .dinb(n551), .dout(n1200));
  jand g0900(.dina(n753), .dinb(G114), .dout(n1201));
  jnot g0901(.din(n1201), .dout(n1202));
  jand g0902(.dina(n1202), .dinb(n1200), .dout(n1203));
  jnot g0903(.din(n1203), .dout(n1204));
  jor  g0904(.dina(n1204), .dinb(n1199), .dout(n1205));
  jnot g0905(.din(n1205), .dout(G865));
  jor  g0906(.dina(n953), .dinb(n748), .dout(n1207));
  jor  g0907(.dina(n765), .dinb(n517), .dout(n1208));
  jand g0908(.dina(n753), .dinb(G53), .dout(n1209));
  jnot g0909(.din(n1209), .dout(n1210));
  jand g0910(.dina(n1210), .dinb(n1208), .dout(n1211));
  jand g0911(.dina(n1211), .dinb(n1207), .dout(G867));
  jand g0912(.dina(n954), .dinb(n747), .dout(n1213));
  jnot g0913(.din(n1213), .dout(n1214));
  jor  g0914(.dina(n765), .dinb(n540), .dout(n1215));
  jand g0915(.dina(n753), .dinb(G113), .dout(n1216));
  jnot g0916(.din(n1216), .dout(n1217));
  jand g0917(.dina(n1217), .dinb(n1215), .dout(n1218));
  jand g0918(.dina(n1218), .dinb(n1214), .dout(G869));
  jand g0919(.dina(n1197), .dinb(n840), .dout(n1220));
  jand g0920(.dina(n1163), .dinb(n843), .dout(n1221));
  jand g0921(.dina(n845), .dinb(G109), .dout(n1222));
  jand g0922(.dina(n847), .dinb(G106), .dout(n1223));
  jor  g0923(.dina(n1223), .dinb(n1222), .dout(n1224));
  jor  g0924(.dina(n1224), .dinb(n1221), .dout(n1225));
  jor  g0925(.dina(n1225), .dinb(n1220), .dout(G712));
  jand g0926(.dina(n1197), .dinb(n793), .dout(n1227));
  jand g0927(.dina(n1163), .dinb(n797), .dout(n1228));
  jand g0928(.dina(n799), .dinb(G109), .dout(n1229));
  jand g0929(.dina(n801), .dinb(G106), .dout(n1230));
  jor  g0930(.dina(n1230), .dinb(n1229), .dout(n1231));
  jor  g0931(.dina(n1231), .dinb(n1228), .dout(n1232));
  jor  g0932(.dina(n1232), .dinb(n1227), .dout(G727));
  jand g0933(.dina(n1205), .dinb(n793), .dout(n1234));
  jnot g0934(.din(G826), .dout(n1235));
  jand g0935(.dina(n1235), .dinb(n797), .dout(n1236));
  jand g0936(.dina(n799), .dinb(G46), .dout(n1237));
  jand g0937(.dina(n801), .dinb(G49), .dout(n1238));
  jor  g0938(.dina(n1238), .dinb(n1237), .dout(n1239));
  jor  g0939(.dina(n1239), .dinb(n1236), .dout(n1240));
  jor  g0940(.dina(n1240), .dinb(n1234), .dout(G732));
  jnot g0941(.din(G867), .dout(n1242));
  jand g0942(.dina(n1242), .dinb(n793), .dout(n1243));
  jnot g0943(.din(G828), .dout(n1244));
  jand g0944(.dina(n1244), .dinb(n797), .dout(n1245));
  jand g0945(.dina(n799), .dinb(G100), .dout(n1246));
  jand g0946(.dina(n801), .dinb(G103), .dout(n1247));
  jor  g0947(.dina(n1247), .dinb(n1246), .dout(n1248));
  jor  g0948(.dina(n1248), .dinb(n1245), .dout(n1249));
  jor  g0949(.dina(n1249), .dinb(n1243), .dout(G737));
  jnot g0950(.din(G869), .dout(n1251));
  jand g0951(.dina(n1251), .dinb(n793), .dout(n1252));
  jnot g0952(.din(G830), .dout(n1253));
  jand g0953(.dina(n1253), .dinb(n797), .dout(n1254));
  jand g0954(.dina(n799), .dinb(G91), .dout(n1255));
  jand g0955(.dina(n801), .dinb(G40), .dout(n1256));
  jor  g0956(.dina(n1256), .dinb(n1255), .dout(n1257));
  jor  g0957(.dina(n1257), .dinb(n1254), .dout(n1258));
  jor  g0958(.dina(n1258), .dinb(n1252), .dout(G742));
  jand g0959(.dina(n1205), .dinb(n840), .dout(n1260));
  jand g0960(.dina(n1235), .dinb(n843), .dout(n1261));
  jand g0961(.dina(n845), .dinb(G46), .dout(n1262));
  jand g0962(.dina(n847), .dinb(G49), .dout(n1263));
  jor  g0963(.dina(n1263), .dinb(n1262), .dout(n1264));
  jor  g0964(.dina(n1264), .dinb(n1261), .dout(n1265));
  jor  g0965(.dina(n1265), .dinb(n1260), .dout(G772));
  jand g0966(.dina(n1242), .dinb(n840), .dout(n1267));
  jand g0967(.dina(n1244), .dinb(n843), .dout(n1268));
  jand g0968(.dina(n845), .dinb(G100), .dout(n1269));
  jand g0969(.dina(n847), .dinb(G103), .dout(n1270));
  jor  g0970(.dina(n1270), .dinb(n1269), .dout(n1271));
  jor  g0971(.dina(n1271), .dinb(n1268), .dout(n1272));
  jor  g0972(.dina(n1272), .dinb(n1267), .dout(G777));
  jand g0973(.dina(n1251), .dinb(n840), .dout(n1274));
  jand g0974(.dina(n1253), .dinb(n843), .dout(n1275));
  jand g0975(.dina(n845), .dinb(G91), .dout(n1276));
  jand g0976(.dina(n847), .dinb(G40), .dout(n1277));
  jor  g0977(.dina(n1277), .dinb(n1276), .dout(n1278));
  jor  g0978(.dina(n1278), .dinb(n1275), .dout(n1279));
  jor  g0979(.dina(n1279), .dinb(n1274), .dout(G782));
  jand g0980(.dina(n1251), .dinb(n985), .dout(n1281));
  jand g0981(.dina(n1253), .dinb(n988), .dout(n1282));
  jand g0982(.dina(n990), .dinb(G203), .dout(n1283));
  jand g0983(.dina(n992), .dinb(G173), .dout(n1284));
  jor  g0984(.dina(n1284), .dinb(n1283), .dout(n1285));
  jor  g0985(.dina(n1285), .dinb(n1282), .dout(n1286));
  jor  g0986(.dina(n1286), .dinb(n1281), .dout(n1287));
  jand g0987(.dina(n1287), .dinb(G137), .dout(G645));
  jand g0988(.dina(n1242), .dinb(n985), .dout(n1289));
  jand g0989(.dina(n1244), .dinb(n988), .dout(n1290));
  jand g0990(.dina(n990), .dinb(G197), .dout(n1291));
  jand g0991(.dina(n992), .dinb(G167), .dout(n1292));
  jor  g0992(.dina(n1292), .dinb(n1291), .dout(n1293));
  jor  g0993(.dina(n1293), .dinb(n1290), .dout(n1294));
  jor  g0994(.dina(n1294), .dinb(n1289), .dout(n1295));
  jand g0995(.dina(n1295), .dinb(G137), .dout(G648));
  jand g0996(.dina(n1205), .dinb(n985), .dout(n1297));
  jand g0997(.dina(n1235), .dinb(n988), .dout(n1298));
  jand g0998(.dina(n990), .dinb(G194), .dout(n1299));
  jand g0999(.dina(n992), .dinb(G164), .dout(n1300));
  jor  g1000(.dina(n1300), .dinb(n1299), .dout(n1301));
  jor  g1001(.dina(n1301), .dinb(n1298), .dout(n1302));
  jor  g1002(.dina(n1302), .dinb(n1297), .dout(n1303));
  jand g1003(.dina(n1303), .dinb(G137), .dout(G651));
  jand g1004(.dina(n1197), .dinb(n985), .dout(n1305));
  jand g1005(.dina(n1163), .dinb(n988), .dout(n1306));
  jand g1006(.dina(n990), .dinb(G191), .dout(n1307));
  jand g1007(.dina(n992), .dinb(G161), .dout(n1308));
  jor  g1008(.dina(n1308), .dinb(n1307), .dout(n1309));
  jor  g1009(.dina(n1309), .dinb(n1306), .dout(n1310));
  jor  g1010(.dina(n1310), .dinb(n1305), .dout(n1311));
  jand g1011(.dina(n1311), .dinb(G137), .dout(G654));
  jand g1012(.dina(n1251), .dinb(n999), .dout(n1313));
  jand g1013(.dina(n1253), .dinb(n1002), .dout(n1314));
  jand g1014(.dina(n1004), .dinb(G203), .dout(n1315));
  jand g1015(.dina(n1006), .dinb(G173), .dout(n1316));
  jor  g1016(.dina(n1316), .dinb(n1315), .dout(n1317));
  jor  g1017(.dina(n1317), .dinb(n1314), .dout(n1318));
  jor  g1018(.dina(n1318), .dinb(n1313), .dout(n1319));
  jand g1019(.dina(n1319), .dinb(G137), .dout(G679));
  jand g1020(.dina(n1242), .dinb(n999), .dout(n1321));
  jand g1021(.dina(n1244), .dinb(n1002), .dout(n1322));
  jand g1022(.dina(n1004), .dinb(G197), .dout(n1323));
  jand g1023(.dina(n1006), .dinb(G167), .dout(n1324));
  jor  g1024(.dina(n1324), .dinb(n1323), .dout(n1325));
  jor  g1025(.dina(n1325), .dinb(n1322), .dout(n1326));
  jor  g1026(.dina(n1326), .dinb(n1321), .dout(n1327));
  jand g1027(.dina(n1327), .dinb(G137), .dout(G682));
  jand g1028(.dina(n1205), .dinb(n999), .dout(n1329));
  jand g1029(.dina(n1235), .dinb(n1002), .dout(n1330));
  jand g1030(.dina(n1004), .dinb(G194), .dout(n1331));
  jand g1031(.dina(n1006), .dinb(G164), .dout(n1332));
  jor  g1032(.dina(n1332), .dinb(n1331), .dout(n1333));
  jor  g1033(.dina(n1333), .dinb(n1330), .dout(n1334));
  jor  g1034(.dina(n1334), .dinb(n1329), .dout(n1335));
  jand g1035(.dina(n1335), .dinb(G137), .dout(G685));
  jand g1036(.dina(n1197), .dinb(n999), .dout(n1337));
  jand g1037(.dina(n1163), .dinb(n1002), .dout(n1338));
  jand g1038(.dina(n1004), .dinb(G191), .dout(n1339));
  jand g1039(.dina(n1006), .dinb(G161), .dout(n1340));
  jor  g1040(.dina(n1340), .dinb(n1339), .dout(n1341));
  jor  g1041(.dina(n1341), .dinb(n1338), .dout(n1342));
  jor  g1042(.dina(n1342), .dinb(n1337), .dout(n1343));
  jand g1043(.dina(n1343), .dinb(G137), .dout(G688));
  jor  g1044(.dina(G4091), .dinb(G120), .dout(n1345));
  jand g1045(.dina(n435), .dinb(G251), .dout(n1346));
  jand g1046(.dina(G341), .dinb(G248), .dout(n1347));
  jor  g1047(.dina(n1347), .dinb(n437), .dout(n1348));
  jor  g1048(.dina(n1348), .dinb(n1346), .dout(n1349));
  jand g1049(.dina(n435), .dinb(n366), .dout(n1350));
  jand g1050(.dina(G341), .dinb(n368), .dout(n1351));
  jor  g1051(.dina(n1351), .dinb(G523), .dout(n1352));
  jor  g1052(.dina(n1352), .dinb(n1350), .dout(n1353));
  jand g1053(.dina(n1353), .dinb(n1349), .dout(n1354));
  jxor g1054(.dina(n408), .dinb(n401), .dout(n1355));
  jxor g1055(.dina(n383), .dinb(n372), .dout(n1356));
  jxor g1056(.dina(n1356), .dinb(n1355), .dout(n1357));
  jxor g1057(.dina(n1357), .dinb(n1354), .dout(n1358));
  jnot g1058(.din(n1358), .dout(n1359));
  jor  g1059(.dina(n410), .dinb(G248), .dout(n1360));
  jor  g1060(.dina(G514), .dinb(n368), .dout(n1361));
  jand g1061(.dina(n1361), .dinb(n1360), .dout(n1362));
  jxor g1062(.dina(n1362), .dinb(n419), .dout(n1363));
  jor  g1063(.dina(G351), .dinb(n402), .dout(n1364));
  jor  g1064(.dina(n385), .dinb(n405), .dout(n1365));
  jand g1065(.dina(n1365), .dinb(G534), .dout(n1366));
  jand g1066(.dina(n1366), .dinb(n1364), .dout(n1367));
  jor  g1067(.dina(G351), .dinb(G254), .dout(n1368));
  jor  g1068(.dina(n385), .dinb(G242), .dout(n1369));
  jand g1069(.dina(n1369), .dinb(n388), .dout(n1370));
  jand g1070(.dina(n1370), .dinb(n1368), .dout(n1371));
  jor  g1071(.dina(n1371), .dinb(n1367), .dout(n1372));
  jand g1072(.dina(n424), .dinb(G251), .dout(n1373));
  jand g1073(.dina(G324), .dinb(G248), .dout(n1374));
  jor  g1074(.dina(n1374), .dinb(n426), .dout(n1375));
  jor  g1075(.dina(n1375), .dinb(n1373), .dout(n1376));
  jand g1076(.dina(n424), .dinb(n366), .dout(n1377));
  jand g1077(.dina(G324), .dinb(n368), .dout(n1378));
  jor  g1078(.dina(n1378), .dinb(G503), .dout(n1379));
  jor  g1079(.dina(n1379), .dinb(n1377), .dout(n1380));
  jand g1080(.dina(n1380), .dinb(n1376), .dout(n1381));
  jxor g1081(.dina(n1381), .dinb(n1372), .dout(n1382));
  jxor g1082(.dina(n1382), .dinb(n1363), .dout(n1383));
  jnot g1083(.din(n1383), .dout(n1384));
  jand g1084(.dina(n1383), .dinb(n1359), .dout(n1385));
  jor  g1085(.dina(n1385), .dinb(G4091), .dout(n1386));
  jor  g1086(.dina(n1345), .dinb(n746), .dout(n1388));
  jand g1087(.dina(n1384), .dinb(n1358), .dout(n1389));
  jor  g1088(.dina(n1386), .dinb(n1389), .dout(n1390));
  jand g1089(.dina(n1390), .dinb(n746), .dout(n1391));
  jnot g1090(.din(n1391), .dout(n1392));
  jand g1091(.dina(n633), .dinb(G2174), .dout(n1393));
  jor  g1092(.dina(n1393), .dinb(n732), .dout(n1394));
  jand g1093(.dina(n736), .dinb(n640), .dout(n1395));
  jor  g1094(.dina(n740), .dinb(n641), .dout(n1396));
  jand g1095(.dina(n1396), .dinb(n646), .dout(n1397));
  jor  g1096(.dina(n1397), .dinb(n1395), .dout(n1398));
  jnot g1097(.din(n1398), .dout(n1399));
  jand g1098(.dina(n1399), .dinb(n739), .dout(n1400));
  jnot g1099(.din(n739), .dout(n1401));
  jand g1100(.dina(n1398), .dinb(n1401), .dout(n1402));
  jor  g1101(.dina(n1402), .dinb(n651), .dout(n1403));
  jor  g1102(.dina(n1403), .dinb(n1400), .dout(n1404));
  jand g1103(.dina(n1404), .dinb(n1394), .dout(n1405));
  jnot g1104(.din(n1394), .dout(n1406));
  jxor g1105(.dina(n1399), .dinb(n968), .dout(n1407));
  jand g1106(.dina(n1407), .dinb(n1406), .dout(n1408));
  jor  g1107(.dina(n1408), .dinb(n1405), .dout(n1409));
  jnot g1108(.din(n1409), .dout(n1410));
  jxor g1109(.dina(n629), .dinb(n625), .dout(n1411));
  jnot g1110(.din(n1411), .dout(n1412));
  jxor g1111(.dina(n806), .dinb(n828), .dout(n1413));
  jnot g1112(.din(n614), .dout(n1414));
  jnot g1113(.din(n717), .dout(n1415));
  jand g1114(.dina(n622), .dinb(n828), .dout(n1416));
  jand g1115(.dina(n628), .dinb(G523), .dout(n1417));
  jor  g1116(.dina(n1417), .dinb(n829), .dout(n1418));
  jor  g1117(.dina(n1418), .dinb(n1416), .dout(n1419));
  jand g1118(.dina(n1419), .dinb(n1415), .dout(n1420));
  jxor g1119(.dina(n622), .dinb(n618), .dout(n1421));
  jnot g1120(.din(n1421), .dout(n1422));
  jor  g1121(.dina(n1422), .dinb(n1420), .dout(n1423));
  jor  g1122(.dina(n1421), .dinb(n819), .dout(n1424));
  jand g1123(.dina(n1424), .dinb(n1423), .dout(n1425));
  jxor g1124(.dina(n1425), .dinb(n1414), .dout(n1426));
  jand g1125(.dina(n1426), .dinb(n1413), .dout(n1427));
  jnot g1126(.din(G2174), .dout(n1428));
  jxor g1127(.dina(n806), .dinb(n721), .dout(n1429));
  jxor g1128(.dina(n1425), .dinb(n614), .dout(n1430));
  jand g1129(.dina(n1430), .dinb(n1429), .dout(n1431));
  jor  g1130(.dina(n1431), .dinb(n1428), .dout(n1432));
  jor  g1131(.dina(n1432), .dinb(n1427), .dout(n1433));
  jxor g1132(.dina(n729), .dinb(n614), .dout(n1434));
  jnot g1133(.din(n1434), .dout(n1435));
  jor  g1134(.dina(n622), .dinb(n721), .dout(n1436));
  jand g1135(.dina(n1436), .dinb(n723), .dout(n1437));
  jxor g1136(.dina(n1437), .dinb(n727), .dout(n1438));
  jand g1137(.dina(n1438), .dinb(n1435), .dout(n1439));
  jnot g1138(.din(n1438), .dout(n1440));
  jand g1139(.dina(n1440), .dinb(n1434), .dout(n1441));
  jor  g1140(.dina(n1441), .dinb(G2174), .dout(n1442));
  jor  g1141(.dina(n1442), .dinb(n1439), .dout(n1443));
  jand g1142(.dina(n1443), .dinb(n1433), .dout(n1444));
  jxor g1143(.dina(n1444), .dinb(n787), .dout(n1445));
  jxor g1144(.dina(n1445), .dinb(n1412), .dout(n1446));
  jor  g1145(.dina(n1446), .dinb(n1410), .dout(n1447));
  jxor g1146(.dina(n1445), .dinb(n1411), .dout(n1448));
  jor  g1147(.dina(n1448), .dinb(n1409), .dout(n1449));
  jand g1148(.dina(n1449), .dinb(G4091), .dout(n1450));
  jand g1149(.dina(n1450), .dinb(n1447), .dout(n1451));
  jor  g1150(.dina(n1451), .dinb(n1392), .dout(n1452));
  jand g1151(.dina(n1452), .dinb(n1388), .dout(G843));
  jor  g1152(.dina(G4091), .dinb(G118), .dout(n1454));
  jand g1153(.dina(G251), .dinb(n460), .dout(n1455));
  jand g1154(.dina(G248), .dinb(G234), .dout(n1456));
  jor  g1155(.dina(n1456), .dinb(n462), .dout(n1457));
  jor  g1156(.dina(n1457), .dinb(n1455), .dout(n1458));
  jand g1157(.dina(n366), .dinb(n460), .dout(n1459));
  jand g1158(.dina(n368), .dinb(G234), .dout(n1460));
  jor  g1159(.dina(n1460), .dinb(G435), .dout(n1461));
  jor  g1160(.dina(n1461), .dinb(n1459), .dout(n1462));
  jand g1161(.dina(n1462), .dinb(n1458), .dout(n1463));
  jor  g1162(.dina(n402), .dinb(G226), .dout(n1464));
  jor  g1163(.dina(n405), .dinb(n530), .dout(n1465));
  jand g1164(.dina(n1465), .dinb(G422), .dout(n1466));
  jand g1165(.dina(n1466), .dinb(n1464), .dout(n1467));
  jor  g1166(.dina(G254), .dinb(G226), .dout(n1468));
  jor  g1167(.dina(G242), .dinb(n530), .dout(n1469));
  jand g1168(.dina(n1469), .dinb(n532), .dout(n1470));
  jand g1169(.dina(n1470), .dinb(n1468), .dout(n1471));
  jor  g1170(.dina(n1471), .dinb(n1467), .dout(n1472));
  jxor g1171(.dina(n1472), .dinb(n528), .dout(n1473));
  jor  g1172(.dina(n402), .dinb(G218), .dout(n1474));
  jor  g1173(.dina(n405), .dinb(n507), .dout(n1475));
  jand g1174(.dina(n1475), .dinb(G468), .dout(n1476));
  jand g1175(.dina(n1476), .dinb(n1474), .dout(n1477));
  jor  g1176(.dina(G254), .dinb(G218), .dout(n1478));
  jor  g1177(.dina(G242), .dinb(n507), .dout(n1479));
  jand g1178(.dina(n1479), .dinb(n509), .dout(n1480));
  jand g1179(.dina(n1480), .dinb(n1478), .dout(n1481));
  jor  g1180(.dina(n1481), .dinb(n1477), .dout(n1482));
  jand g1181(.dina(G251), .dinb(n541), .dout(n1483));
  jand g1182(.dina(G248), .dinb(G210), .dout(n1484));
  jor  g1183(.dina(n1484), .dinb(n543), .dout(n1485));
  jor  g1184(.dina(n1485), .dinb(n1483), .dout(n1486));
  jand g1185(.dina(n366), .dinb(n541), .dout(n1487));
  jand g1186(.dina(n368), .dinb(G210), .dout(n1488));
  jor  g1187(.dina(n1488), .dinb(G457), .dout(n1489));
  jor  g1188(.dina(n1489), .dinb(n1487), .dout(n1490));
  jand g1189(.dina(n1490), .dinb(n1486), .dout(n1491));
  jxor g1190(.dina(n1491), .dinb(n1482), .dout(n1492));
  jxor g1191(.dina(n1492), .dinb(n1473), .dout(n1493));
  jxor g1192(.dina(n1493), .dinb(n1463), .dout(n1494));
  jand g1193(.dina(n495), .dinb(G251), .dout(n1495));
  jand g1194(.dina(G281), .dinb(G248), .dout(n1496));
  jor  g1195(.dina(n1496), .dinb(n497), .dout(n1497));
  jor  g1196(.dina(n1497), .dinb(n1495), .dout(n1498));
  jand g1197(.dina(n495), .dinb(n366), .dout(n1499));
  jand g1198(.dina(G281), .dinb(n368), .dout(n1500));
  jor  g1199(.dina(n1500), .dinb(G374), .dout(n1501));
  jor  g1200(.dina(n1501), .dinb(n1499), .dout(n1502));
  jand g1201(.dina(n1502), .dinb(n1498), .dout(n1503));
  jand g1202(.dina(n449), .dinb(G251), .dout(n1504));
  jand g1203(.dina(G265), .dinb(G248), .dout(n1505));
  jor  g1204(.dina(n1505), .dinb(n451), .dout(n1506));
  jor  g1205(.dina(n1506), .dinb(n1504), .dout(n1507));
  jand g1206(.dina(n449), .dinb(n366), .dout(n1508));
  jand g1207(.dina(G265), .dinb(n368), .dout(n1509));
  jor  g1208(.dina(n1509), .dinb(G400), .dout(n1510));
  jor  g1209(.dina(n1510), .dinb(n1508), .dout(n1511));
  jand g1210(.dina(n1511), .dinb(n1507), .dout(n1512));
  jxor g1211(.dina(n1512), .dinb(n1503), .dout(n1513));
  jor  g1212(.dina(G257), .dinb(n402), .dout(n1514));
  jor  g1213(.dina(n471), .dinb(n405), .dout(n1515));
  jand g1214(.dina(n1515), .dinb(G389), .dout(n1516));
  jand g1215(.dina(n1516), .dinb(n1514), .dout(n1517));
  jor  g1216(.dina(G257), .dinb(G254), .dout(n1518));
  jor  g1217(.dina(n471), .dinb(G242), .dout(n1519));
  jand g1218(.dina(n1519), .dinb(n473), .dout(n1520));
  jand g1219(.dina(n1520), .dinb(n1518), .dout(n1521));
  jor  g1220(.dina(n1521), .dinb(n1517), .dout(n1522));
  jand g1221(.dina(n484), .dinb(G251), .dout(n1523));
  jand g1222(.dina(G273), .dinb(G248), .dout(n1524));
  jor  g1223(.dina(n1524), .dinb(n486), .dout(n1525));
  jor  g1224(.dina(n1525), .dinb(n1523), .dout(n1526));
  jand g1225(.dina(n484), .dinb(n366), .dout(n1527));
  jand g1226(.dina(G273), .dinb(n368), .dout(n1528));
  jor  g1227(.dina(n1528), .dinb(G411), .dout(n1529));
  jor  g1228(.dina(n1529), .dinb(n1527), .dout(n1530));
  jand g1229(.dina(n1530), .dinb(n1526), .dout(n1531));
  jxor g1230(.dina(n1531), .dinb(n1522), .dout(n1532));
  jxor g1231(.dina(n1532), .dinb(n1513), .dout(n1533));
  jand g1232(.dina(n1533), .dinb(n1494), .dout(n1534));
  jnot g1233(.din(n1534), .dout(n1535));
  jor  g1234(.dina(n1533), .dinb(n1494), .dout(n1536));
  jand g1235(.dina(n1536), .dinb(n750), .dout(n1537));
  jand g1236(.dina(n1537), .dinb(n1535), .dout(n1538));
  jor  g1237(.dina(n1454), .dinb(n746), .dout(n1539));
  jor  g1238(.dina(n1538), .dinb(G4092), .dout(n1540));
  jxor g1239(.dina(n583), .dinb(n578), .dout(n1541));
  jxor g1240(.dina(n1541), .dinb(n943), .dout(n1542));
  jnot g1241(.din(n1542), .dout(n1543));
  jand g1242(.dina(n587), .dinb(G1497), .dout(n1544));
  jor  g1243(.dina(n1544), .dinb(n696), .dout(n1545));
  jnot g1244(.din(n1545), .dout(n1546));
  jor  g1245(.dina(n944), .dinb(n930), .dout(n1547));
  jand g1246(.dina(n1547), .dinb(n706), .dout(n1548));
  jxor g1247(.dina(n1548), .dinb(n928), .dout(n1549));
  jxor g1248(.dina(n605), .dinb(n948), .dout(n1550));
  jxor g1249(.dina(n1550), .dinb(n1549), .dout(n1551));
  jand g1250(.dina(n1551), .dinb(n1546), .dout(n1552));
  jxor g1251(.dina(n605), .dinb(n703), .dout(n1553));
  jand g1252(.dina(n605), .dinb(n948), .dout(n1554));
  jor  g1253(.dina(n1554), .dinb(n702), .dout(n1555));
  jnot g1254(.din(n1555), .dout(n1556));
  jor  g1255(.dina(n1556), .dinb(n930), .dout(n1557));
  jor  g1256(.dina(n1555), .dinb(n707), .dout(n1558));
  jand g1257(.dina(n1558), .dinb(n1557), .dout(n1559));
  jxor g1258(.dina(n1559), .dinb(n596), .dout(n1560));
  jand g1259(.dina(n1560), .dinb(n1553), .dout(n1561));
  jnot g1260(.din(n1561), .dout(n1562));
  jor  g1261(.dina(n1560), .dinb(n1553), .dout(n1563));
  jand g1262(.dina(n1563), .dinb(n1545), .dout(n1564));
  jand g1263(.dina(n1564), .dinb(n1562), .dout(n1565));
  jor  g1264(.dina(n1565), .dinb(n1552), .dout(n1566));
  jnot g1265(.din(G1497), .dout(n1567));
  jand g1266(.dina(n682), .dinb(n687), .dout(n1568));
  jand g1267(.dina(n1568), .dinb(n574), .dout(n1569));
  jxor g1268(.dina(n1569), .dinb(n561), .dout(n1570));
  jxor g1269(.dina(n572), .dinb(n681), .dout(n1571));
  jor  g1270(.dina(n856), .dinb(n853), .dout(n1572));
  jand g1271(.dina(n693), .dinb(n585), .dout(n1573));
  jor  g1272(.dina(n1573), .dinb(n855), .dout(n1574));
  jand g1273(.dina(n1574), .dinb(n1572), .dout(n1575));
  jxor g1274(.dina(n1575), .dinb(n1571), .dout(n1576));
  jxor g1275(.dina(n1576), .dinb(n1570), .dout(n1577));
  jor  g1276(.dina(n1577), .dinb(n1567), .dout(n1578));
  jxor g1277(.dina(n693), .dinb(n572), .dout(n1579));
  jor  g1278(.dina(n857), .dinb(n681), .dout(n1580));
  jnot g1279(.din(n681), .dout(n1581));
  jor  g1280(.dina(n680), .dinb(n1581), .dout(n1582));
  jor  g1281(.dina(n1582), .dinb(n689), .dout(n1583));
  jxor g1282(.dina(n1583), .dinb(n567), .dout(n1584));
  jand g1283(.dina(n1584), .dinb(n1580), .dout(n1585));
  jxor g1284(.dina(n1568), .dinb(n561), .dout(n1586));
  jxor g1285(.dina(n1586), .dinb(n1585), .dout(n1587));
  jxor g1286(.dina(n1587), .dinb(n1579), .dout(n1588));
  jor  g1287(.dina(n1588), .dinb(G1497), .dout(n1589));
  jand g1288(.dina(n1589), .dinb(n1578), .dout(n1590));
  jxor g1289(.dina(n1590), .dinb(n1566), .dout(n1591));
  jand g1290(.dina(n1591), .dinb(n1543), .dout(n1592));
  jnot g1291(.din(n1592), .dout(n1593));
  jor  g1292(.dina(n1591), .dinb(n1543), .dout(n1594));
  jand g1293(.dina(n1594), .dinb(G4091), .dout(n1595));
  jand g1294(.dina(n1595), .dinb(n1593), .dout(n1596));
  jor  g1295(.dina(n1596), .dinb(n1540), .dout(n1597));
  jand g1296(.dina(n1597), .dinb(n1539), .dout(G882));
  jand g1297(.dina(G4092), .dinb(G97), .dout(n1599));
  jnot g1298(.din(n1599), .dout(n1600));
  jand g1299(.dina(n1600), .dinb(n1597), .dout(n1601));
  jnot g1300(.din(n1601), .dout(n1602));
  jand g1301(.dina(n1602), .dinb(n793), .dout(n1603));
  jnot g1302(.din(n1447), .dout(n1604));
  jand g1303(.dina(n1446), .dinb(n1410), .dout(n1605));
  jor  g1304(.dina(n1605), .dinb(n750), .dout(n1606));
  jor  g1305(.dina(n1606), .dinb(n1604), .dout(n1607));
  jand g1306(.dina(n1607), .dinb(n1391), .dout(n1608));
  jand g1307(.dina(G4092), .dinb(G94), .dout(n1609));
  jor  g1308(.dina(n1609), .dinb(n1608), .dout(n1610));
  jand g1309(.dina(n1610), .dinb(n797), .dout(n1611));
  jand g1310(.dina(n799), .dinb(G14), .dout(n1612));
  jand g1311(.dina(n801), .dinb(G64), .dout(n1613));
  jor  g1312(.dina(n1613), .dinb(n1612), .dout(n1614));
  jor  g1313(.dina(n1614), .dinb(n1611), .dout(n1615));
  jor  g1314(.dina(n1615), .dinb(n1603), .dout(G767));
  jand g1315(.dina(n1602), .dinb(n840), .dout(n1617));
  jand g1316(.dina(n1610), .dinb(n843), .dout(n1618));
  jand g1317(.dina(n845), .dinb(G14), .dout(n1619));
  jand g1318(.dina(n847), .dinb(G64), .dout(n1620));
  jor  g1319(.dina(n1620), .dinb(n1619), .dout(n1621));
  jor  g1320(.dina(n1621), .dinb(n1618), .dout(n1622));
  jor  g1321(.dina(n1622), .dinb(n1617), .dout(G807));
  jnot g1322(.din(G137), .dout(n1624));
  jnot g1323(.din(n985), .dout(n1625));
  jor  g1324(.dina(n1601), .dinb(n1625), .dout(n1626));
  jnot g1325(.din(n988), .dout(n1627));
  jnot g1326(.din(n1609), .dout(n1628));
  jand g1327(.dina(n1628), .dinb(n1452), .dout(n1629));
  jor  g1328(.dina(n1629), .dinb(n1627), .dout(n1630));
  jnot g1329(.din(G179), .dout(n1631));
  jnot g1330(.din(n992), .dout(n1632));
  jor  g1331(.dina(n1632), .dinb(n1631), .dout(n1633));
  jnot g1332(.din(G176), .dout(n1634));
  jnot g1333(.din(n990), .dout(n1635));
  jor  g1334(.dina(n1635), .dinb(n1634), .dout(n1636));
  jand g1335(.dina(n1636), .dinb(n1633), .dout(n1637));
  jand g1336(.dina(n1637), .dinb(n1630), .dout(n1638));
  jand g1337(.dina(n1638), .dinb(n1626), .dout(n1639));
  jor  g1338(.dina(n1639), .dinb(n1624), .dout(G658));
  jnot g1339(.din(n999), .dout(n1641));
  jor  g1340(.dina(n1601), .dinb(n1641), .dout(n1642));
  jnot g1341(.din(n1002), .dout(n1643));
  jor  g1342(.dina(n1629), .dinb(n1643), .dout(n1644));
  jnot g1343(.din(n1006), .dout(n1645));
  jor  g1344(.dina(n1645), .dinb(n1631), .dout(n1646));
  jnot g1345(.din(n1004), .dout(n1647));
  jor  g1346(.dina(n1647), .dinb(n1634), .dout(n1648));
  jand g1347(.dina(n1648), .dinb(n1646), .dout(n1649));
  jand g1348(.dina(n1649), .dinb(n1644), .dout(n1650));
  jand g1349(.dina(n1650), .dinb(n1642), .dout(n1651));
  jor  g1350(.dina(n1651), .dinb(n1624), .dout(G690));
  jdff  g1351(.din(G141), .dout(G144));
  jdff  g1352(.din(G293), .dout(G298));
  jdff  g1353(.din(G3173), .dout(G973));
  jnot g1354(.din(G545), .dout(G603));
  jnot g1355(.din(G545), .dout(G604));
  jdff  g1356(.din(G137), .dout(G926));
  jdff  g1357(.din(G141), .dout(G923));
  jdff  g1358(.din(G1), .dout(G921));
  jdff  g1359(.din(G549), .dout(G892));
  jdff  g1360(.din(G299), .dout(G887));
  jnot g1361(.din(G549), .dout(G606));
  jdff  g1362(.din(G1), .dout(G993));
  jdff  g1363(.din(G1), .dout(G978));
  jdff  g1364(.din(G1), .dout(G949));
  jdff  g1365(.din(G1), .dout(G939));
  jdff  g1366(.din(G299), .dout(G889));
  jor  g1367(.dina(n336), .dinb(n333), .dout(G717));
  jand g1368(.dina(n652), .dinb(n633), .dout(G626));
  jand g1369(.dina(n607), .dinb(n587), .dout(G632));
  jor  g1370(.dina(n709), .dinb(n697), .dout(G621));
  jor  g1371(.dina(n742), .dinb(n733), .dout(G629));
endmodule


