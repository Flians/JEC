/*

c7552:
	jxor: 228
	jspl: 345
	jspl3: 346
	jnot: 270
	jdff: 4170
	jor: 395
	jand: 513

Summary:
	jxor: 228
	jspl: 345
	jspl3: 346
	jnot: 270
	jdff: 4170
	jor: 395
	jand: 513
*/

module c7552(gclk, G1, G5, G9, G12, G15, G18, G23, G26, G29, G32, G35, G38, G41, G44, G47, G50, G53, G54, G55, G56, G57, G58, G59, G60, G61, G62, G63, G64, G65, G66, G69, G70, G73, G74, G75, G76, G77, G78, G79, G80, G81, G82, G83, G84, G85, G86, G87, G88, G89, G94, G97, G100, G103, G106, G109, G110, G111, G112, G113, G114, G115, G118, G121, G124, G127, G130, G133, G134, G135, G138, G141, G144, G147, G150, G151, G152, G153, G154, G155, G156, G157, G158, G159, G160, G161, G162, G163, G164, G165, G166, G167, G168, G169, G170, G171, G172, G173, G174, G175, G176, G177, G178, G179, G180, G181, G182, G183, G184, G185, G186, G187, G188, G189, G190, G191, G192, G193, G194, G195, G196, G197, G198, G199, G200, G201, G202, G203, G204, G205, G206, G207, G208, G209, G210, G211, G212, G213, G214, G215, G216, G217, G218, G219, G220, G221, G222, G223, G224, G225, G226, G227, G228, G229, G230, G231, G232, G233, G234, G235, G236, G237, G238, G239, G240, G339, G1197, G1455, G1459, G1462, G1469, G1480, G1486, G1492, G1496, G2204, G2208, G2211, G2218, G2224, G2230, G2236, G2239, G2247, G2253, G2256, G3698, G3701, G3705, G3711, G3717, G3723, G3729, G3737, G3743, G3749, G4393, G4394, G4400, G4405, G4410, G4415, G4420, G4427, G4432, G4437, G4526, G4528, G2, G3, G450, G448, G444, G442, G440, G438, G496, G494, G492, G490, G488, G486, G484, G482, G480, G560, G542, G558, G556, G554, G552, G550, G548, G546, G544, G540, G538, G536, G534, G532, G530, G528, G526, G524, G279, G436, G478, G522, G402, G404, G406, G408, G410, G432, G446, G284, G286, G289, G292, G341, G281, G453, G278, G373, G246, G258, G264, G270, G388, G391, G394, G397, G376, G379, G382, G385, G412, G414, G416, G249, G295, G324, G252, G276, G310, G313, G316, G319, G327, G330, G333, G336, G418, G273, G298, G301, G304, G307, G344, G422, G469, G419, G471, G359, G362, G365, G368, G347, G350, G353, G356, G321, G338, G370, G399);
	input gclk;
	input G1;
	input G5;
	input G9;
	input G12;
	input G15;
	input G18;
	input G23;
	input G26;
	input G29;
	input G32;
	input G35;
	input G38;
	input G41;
	input G44;
	input G47;
	input G50;
	input G53;
	input G54;
	input G55;
	input G56;
	input G57;
	input G58;
	input G59;
	input G60;
	input G61;
	input G62;
	input G63;
	input G64;
	input G65;
	input G66;
	input G69;
	input G70;
	input G73;
	input G74;
	input G75;
	input G76;
	input G77;
	input G78;
	input G79;
	input G80;
	input G81;
	input G82;
	input G83;
	input G84;
	input G85;
	input G86;
	input G87;
	input G88;
	input G89;
	input G94;
	input G97;
	input G100;
	input G103;
	input G106;
	input G109;
	input G110;
	input G111;
	input G112;
	input G113;
	input G114;
	input G115;
	input G118;
	input G121;
	input G124;
	input G127;
	input G130;
	input G133;
	input G134;
	input G135;
	input G138;
	input G141;
	input G144;
	input G147;
	input G150;
	input G151;
	input G152;
	input G153;
	input G154;
	input G155;
	input G156;
	input G157;
	input G158;
	input G159;
	input G160;
	input G161;
	input G162;
	input G163;
	input G164;
	input G165;
	input G166;
	input G167;
	input G168;
	input G169;
	input G170;
	input G171;
	input G172;
	input G173;
	input G174;
	input G175;
	input G176;
	input G177;
	input G178;
	input G179;
	input G180;
	input G181;
	input G182;
	input G183;
	input G184;
	input G185;
	input G186;
	input G187;
	input G188;
	input G189;
	input G190;
	input G191;
	input G192;
	input G193;
	input G194;
	input G195;
	input G196;
	input G197;
	input G198;
	input G199;
	input G200;
	input G201;
	input G202;
	input G203;
	input G204;
	input G205;
	input G206;
	input G207;
	input G208;
	input G209;
	input G210;
	input G211;
	input G212;
	input G213;
	input G214;
	input G215;
	input G216;
	input G217;
	input G218;
	input G219;
	input G220;
	input G221;
	input G222;
	input G223;
	input G224;
	input G225;
	input G226;
	input G227;
	input G228;
	input G229;
	input G230;
	input G231;
	input G232;
	input G233;
	input G234;
	input G235;
	input G236;
	input G237;
	input G238;
	input G239;
	input G240;
	input G339;
	input G1197;
	input G1455;
	input G1459;
	input G1462;
	input G1469;
	input G1480;
	input G1486;
	input G1492;
	input G1496;
	input G2204;
	input G2208;
	input G2211;
	input G2218;
	input G2224;
	input G2230;
	input G2236;
	input G2239;
	input G2247;
	input G2253;
	input G2256;
	input G3698;
	input G3701;
	input G3705;
	input G3711;
	input G3717;
	input G3723;
	input G3729;
	input G3737;
	input G3743;
	input G3749;
	input G4393;
	input G4394;
	input G4400;
	input G4405;
	input G4410;
	input G4415;
	input G4420;
	input G4427;
	input G4432;
	input G4437;
	input G4526;
	input G4528;
	output G2;
	output G3;
	output G450;
	output G448;
	output G444;
	output G442;
	output G440;
	output G438;
	output G496;
	output G494;
	output G492;
	output G490;
	output G488;
	output G486;
	output G484;
	output G482;
	output G480;
	output G560;
	output G542;
	output G558;
	output G556;
	output G554;
	output G552;
	output G550;
	output G548;
	output G546;
	output G544;
	output G540;
	output G538;
	output G536;
	output G534;
	output G532;
	output G530;
	output G528;
	output G526;
	output G524;
	output G279;
	output G436;
	output G478;
	output G522;
	output G402;
	output G404;
	output G406;
	output G408;
	output G410;
	output G432;
	output G446;
	output G284;
	output G286;
	output G289;
	output G292;
	output G341;
	output G281;
	output G453;
	output G278;
	output G373;
	output G246;
	output G258;
	output G264;
	output G270;
	output G388;
	output G391;
	output G394;
	output G397;
	output G376;
	output G379;
	output G382;
	output G385;
	output G412;
	output G414;
	output G416;
	output G249;
	output G295;
	output G324;
	output G252;
	output G276;
	output G310;
	output G313;
	output G316;
	output G319;
	output G327;
	output G330;
	output G333;
	output G336;
	output G418;
	output G273;
	output G298;
	output G301;
	output G304;
	output G307;
	output G344;
	output G422;
	output G469;
	output G419;
	output G471;
	output G359;
	output G362;
	output G365;
	output G368;
	output G347;
	output G350;
	output G353;
	output G356;
	output G321;
	output G338;
	output G370;
	output G399;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n331;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n345;
	wire n347;
	wire n348;
	wire n349;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1134;
	wire n1136;
	wire n1137;
	wire n1139;
	wire n1140;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1146;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1410;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1417;
	wire n1418;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1429;
	wire n1430;
	wire n1432;
	wire n1433;
	wire n1435;
	wire n1436;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1451;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1477;
	wire n1479;
	wire n1480;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1490;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1667;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1673;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1684;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1690;
	wire n1691;
	wire n1692;
	wire n1693;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1707;
	wire n1708;
	wire[2:0] w_G1_0;
	wire[2:0] w_G1_1;
	wire[2:0] w_G5_0;
	wire[2:0] w_G5_1;
	wire[2:0] w_G15_0;
	wire[2:0] w_G18_0;
	wire[2:0] w_G18_1;
	wire[2:0] w_G18_2;
	wire[2:0] w_G18_3;
	wire[2:0] w_G18_4;
	wire[2:0] w_G18_5;
	wire[2:0] w_G18_6;
	wire[2:0] w_G18_7;
	wire[2:0] w_G18_8;
	wire[2:0] w_G18_9;
	wire[2:0] w_G18_10;
	wire[2:0] w_G18_11;
	wire[2:0] w_G18_12;
	wire[2:0] w_G18_13;
	wire[2:0] w_G18_14;
	wire[2:0] w_G18_15;
	wire[2:0] w_G18_16;
	wire[2:0] w_G18_17;
	wire[2:0] w_G18_18;
	wire[2:0] w_G18_19;
	wire[2:0] w_G18_20;
	wire[2:0] w_G18_21;
	wire[2:0] w_G18_22;
	wire[2:0] w_G18_23;
	wire[2:0] w_G18_24;
	wire[2:0] w_G18_25;
	wire[2:0] w_G18_26;
	wire[2:0] w_G18_27;
	wire[2:0] w_G18_28;
	wire[2:0] w_G18_29;
	wire[2:0] w_G18_30;
	wire[2:0] w_G18_31;
	wire[2:0] w_G18_32;
	wire[2:0] w_G18_33;
	wire[2:0] w_G18_34;
	wire[2:0] w_G18_35;
	wire[2:0] w_G18_36;
	wire[2:0] w_G18_37;
	wire[2:0] w_G18_38;
	wire[2:0] w_G18_39;
	wire[2:0] w_G18_40;
	wire[2:0] w_G18_41;
	wire[2:0] w_G18_42;
	wire[2:0] w_G18_43;
	wire[2:0] w_G18_44;
	wire[2:0] w_G18_45;
	wire[2:0] w_G18_46;
	wire[2:0] w_G18_47;
	wire[2:0] w_G18_48;
	wire[2:0] w_G18_49;
	wire[2:0] w_G18_50;
	wire[2:0] w_G18_51;
	wire[2:0] w_G18_52;
	wire[2:0] w_G18_53;
	wire[2:0] w_G18_54;
	wire[2:0] w_G18_55;
	wire[2:0] w_G18_56;
	wire[2:0] w_G18_57;
	wire[2:0] w_G18_58;
	wire[2:0] w_G38_0;
	wire[2:0] w_G38_1;
	wire[2:0] w_G41_0;
	wire[1:0] w_G69_0;
	wire[1:0] w_G70_0;
	wire[2:0] w_G106_0;
	wire[1:0] w_G106_1;
	wire[1:0] w_G229_0;
	wire[2:0] w_G1455_0;
	wire[1:0] w_G1459_0;
	wire[2:0] w_G1462_0;
	wire[2:0] w_G1469_0;
	wire[1:0] w_G1469_1;
	wire[2:0] w_G1480_0;
	wire[2:0] w_G1486_0;
	wire[2:0] w_G1492_0;
	wire[1:0] w_G1492_1;
	wire[2:0] w_G1496_0;
	wire[2:0] w_G2204_0;
	wire[1:0] w_G2208_0;
	wire[2:0] w_G2211_0;
	wire[2:0] w_G2218_0;
	wire[2:0] w_G2224_0;
	wire[1:0] w_G2224_1;
	wire[2:0] w_G2230_0;
	wire[1:0] w_G2230_1;
	wire[2:0] w_G2236_0;
	wire[1:0] w_G2236_1;
	wire[2:0] w_G2239_0;
	wire[2:0] w_G2247_0;
	wire[2:0] w_G2253_0;
	wire[1:0] w_G2253_1;
	wire[2:0] w_G2256_0;
	wire[1:0] w_G2256_1;
	wire[1:0] w_G3698_0;
	wire[2:0] w_G3701_0;
	wire[1:0] w_G3701_1;
	wire[2:0] w_G3705_0;
	wire[2:0] w_G3705_1;
	wire[1:0] w_G3705_2;
	wire[2:0] w_G3711_0;
	wire[1:0] w_G3711_1;
	wire[2:0] w_G3717_0;
	wire[2:0] w_G3717_1;
	wire[1:0] w_G3717_2;
	wire[2:0] w_G3723_0;
	wire[1:0] w_G3723_1;
	wire[2:0] w_G3729_0;
	wire[1:0] w_G3729_1;
	wire[2:0] w_G3737_0;
	wire[1:0] w_G3737_1;
	wire[2:0] w_G3743_0;
	wire[2:0] w_G3743_1;
	wire[2:0] w_G3749_0;
	wire[1:0] w_G3749_1;
	wire[1:0] w_G4393_0;
	wire[2:0] w_G4394_0;
	wire[1:0] w_G4394_1;
	wire[2:0] w_G4400_0;
	wire[2:0] w_G4405_0;
	wire[2:0] w_G4405_1;
	wire[2:0] w_G4410_0;
	wire[1:0] w_G4410_1;
	wire[2:0] w_G4415_0;
	wire[1:0] w_G4415_1;
	wire[2:0] w_G4420_0;
	wire[1:0] w_G4427_0;
	wire[2:0] w_G4432_0;
	wire[1:0] w_G4432_1;
	wire[2:0] w_G4437_0;
	wire[2:0] w_G4526_0;
	wire[1:0] w_G4526_1;
	wire[2:0] w_G4528_0;
	wire w_G404_0;
	wire G404_fa_;
	wire w_G406_0;
	wire G406_fa_;
	wire w_G408_0;
	wire G408_fa_;
	wire w_G410_0;
	wire G410_fa_;
	wire w_G412_0;
	wire G412_fa_;
	wire w_G414_0;
	wire G414_fa_;
	wire w_G416_0;
	wire G416_fa_;
	wire[1:0] w_n345_0;
	wire[1:0] w_n349_0;
	wire[2:0] w_n353_0;
	wire[2:0] w_n354_0;
	wire[2:0] w_n354_1;
	wire[2:0] w_n355_0;
	wire[2:0] w_n355_1;
	wire[2:0] w_n355_2;
	wire[2:0] w_n355_3;
	wire[2:0] w_n355_4;
	wire[2:0] w_n355_5;
	wire[2:0] w_n355_6;
	wire[2:0] w_n355_7;
	wire[2:0] w_n355_8;
	wire[2:0] w_n355_9;
	wire[2:0] w_n355_10;
	wire[2:0] w_n355_11;
	wire[2:0] w_n355_12;
	wire[2:0] w_n355_13;
	wire[2:0] w_n355_14;
	wire[2:0] w_n355_15;
	wire[2:0] w_n355_16;
	wire[2:0] w_n355_17;
	wire[2:0] w_n355_18;
	wire[2:0] w_n355_19;
	wire[2:0] w_n355_20;
	wire[2:0] w_n355_21;
	wire[2:0] w_n355_22;
	wire[2:0] w_n355_23;
	wire[2:0] w_n355_24;
	wire[2:0] w_n355_25;
	wire[1:0] w_n355_26;
	wire[2:0] w_n356_0;
	wire[1:0] w_n358_0;
	wire[1:0] w_n359_0;
	wire[2:0] w_n362_0;
	wire[1:0] w_n364_0;
	wire[1:0] w_n365_0;
	wire[1:0] w_n366_0;
	wire[1:0] w_n370_0;
	wire[2:0] w_n371_0;
	wire[1:0] w_n371_1;
	wire[2:0] w_n372_0;
	wire[2:0] w_n372_1;
	wire[1:0] w_n376_0;
	wire[2:0] w_n377_0;
	wire[2:0] w_n377_1;
	wire[2:0] w_n379_0;
	wire[1:0] w_n379_1;
	wire[2:0] w_n380_0;
	wire[1:0] w_n385_0;
	wire[2:0] w_n386_0;
	wire[2:0] w_n387_0;
	wire[2:0] w_n387_1;
	wire[2:0] w_n388_0;
	wire[1:0] w_n389_0;
	wire[2:0] w_n390_0;
	wire[1:0] w_n390_1;
	wire[2:0] w_n395_0;
	wire[1:0] w_n400_0;
	wire[2:0] w_n401_0;
	wire[2:0] w_n401_1;
	wire[2:0] w_n402_0;
	wire[1:0] w_n402_1;
	wire[1:0] w_n403_0;
	wire[1:0] w_n404_0;
	wire[2:0] w_n405_0;
	wire[2:0] w_n407_0;
	wire[1:0] w_n408_0;
	wire[1:0] w_n410_0;
	wire[2:0] w_n412_0;
	wire[2:0] w_n413_0;
	wire[1:0] w_n413_1;
	wire[2:0] w_n417_0;
	wire[1:0] w_n419_0;
	wire[2:0] w_n422_0;
	wire[2:0] w_n422_1;
	wire[1:0] w_n427_0;
	wire[2:0] w_n428_0;
	wire[2:0] w_n429_0;
	wire[2:0] w_n429_1;
	wire[1:0] w_n429_2;
	wire[1:0] w_n430_0;
	wire[1:0] w_n434_0;
	wire[2:0] w_n435_0;
	wire[1:0] w_n435_1;
	wire[1:0] w_n436_0;
	wire[1:0] w_n437_0;
	wire[1:0] w_n441_0;
	wire[2:0] w_n442_0;
	wire[1:0] w_n443_0;
	wire[1:0] w_n445_0;
	wire[2:0] w_n446_0;
	wire[1:0] w_n446_1;
	wire[1:0] w_n448_0;
	wire[2:0] w_n449_0;
	wire[2:0] w_n450_0;
	wire[1:0] w_n452_0;
	wire[1:0] w_n454_0;
	wire[1:0] w_n455_0;
	wire[2:0] w_n456_0;
	wire[1:0] w_n457_0;
	wire[2:0] w_n458_0;
	wire[2:0] w_n460_0;
	wire[1:0] w_n461_0;
	wire[2:0] w_n462_0;
	wire[1:0] w_n464_0;
	wire[2:0] w_n465_0;
	wire[1:0] w_n466_0;
	wire[1:0] w_n468_0;
	wire[2:0] w_n469_0;
	wire[1:0] w_n469_1;
	wire[2:0] w_n470_0;
	wire[2:0] w_n471_0;
	wire[1:0] w_n473_0;
	wire[2:0] w_n474_0;
	wire[1:0] w_n474_1;
	wire[2:0] w_n475_0;
	wire[1:0] w_n475_1;
	wire[1:0] w_n477_0;
	wire[1:0] w_n478_0;
	wire[1:0] w_n479_0;
	wire[2:0] w_n480_0;
	wire[1:0] w_n480_1;
	wire[2:0] w_n481_0;
	wire[1:0] w_n482_0;
	wire[1:0] w_n484_0;
	wire[2:0] w_n485_0;
	wire[2:0] w_n486_0;
	wire[1:0] w_n488_0;
	wire[1:0] w_n489_0;
	wire[2:0] w_n490_0;
	wire[2:0] w_n491_0;
	wire[1:0] w_n491_1;
	wire[1:0] w_n493_0;
	wire[1:0] w_n494_0;
	wire[1:0] w_n502_0;
	wire[1:0] w_n503_0;
	wire[1:0] w_n505_0;
	wire[2:0] w_n507_0;
	wire[2:0] w_n507_1;
	wire[1:0] w_n508_0;
	wire[1:0] w_n509_0;
	wire[1:0] w_n510_0;
	wire[1:0] w_n512_0;
	wire[2:0] w_n514_0;
	wire[2:0] w_n516_0;
	wire[1:0] w_n518_0;
	wire[1:0] w_n519_0;
	wire[2:0] w_n520_0;
	wire[1:0] w_n522_0;
	wire[2:0] w_n523_0;
	wire[2:0] w_n524_0;
	wire[2:0] w_n524_1;
	wire[1:0] w_n524_2;
	wire[2:0] w_n525_0;
	wire[1:0] w_n527_0;
	wire[2:0] w_n528_0;
	wire[1:0] w_n528_1;
	wire[1:0] w_n529_0;
	wire[1:0] w_n530_0;
	wire[2:0] w_n531_0;
	wire[1:0] w_n533_0;
	wire[2:0] w_n534_0;
	wire[1:0] w_n534_1;
	wire[2:0] w_n535_0;
	wire[1:0] w_n535_1;
	wire[1:0] w_n536_0;
	wire[1:0] w_n538_0;
	wire[2:0] w_n539_0;
	wire[1:0] w_n539_1;
	wire[2:0] w_n540_0;
	wire[1:0] w_n542_0;
	wire[1:0] w_n549_0;
	wire[1:0] w_n551_0;
	wire[1:0] w_n552_0;
	wire[1:0] w_n553_0;
	wire[2:0] w_n554_0;
	wire[2:0] w_n556_0;
	wire[1:0] w_n557_0;
	wire[2:0] w_n558_0;
	wire[1:0] w_n560_0;
	wire[2:0] w_n562_0;
	wire[1:0] w_n563_0;
	wire[2:0] w_n564_0;
	wire[2:0] w_n565_0;
	wire[2:0] w_n565_1;
	wire[2:0] w_n565_2;
	wire[2:0] w_n565_3;
	wire[2:0] w_n565_4;
	wire[2:0] w_n565_5;
	wire[2:0] w_n565_6;
	wire[2:0] w_n565_7;
	wire[2:0] w_n565_8;
	wire[2:0] w_n565_9;
	wire[1:0] w_n565_10;
	wire[2:0] w_n567_0;
	wire[1:0] w_n567_1;
	wire[2:0] w_n568_0;
	wire[2:0] w_n569_0;
	wire[1:0] w_n570_0;
	wire[2:0] w_n572_0;
	wire[1:0] w_n572_1;
	wire[2:0] w_n573_0;
	wire[1:0] w_n573_1;
	wire[1:0] w_n574_0;
	wire[1:0] w_n575_0;
	wire[2:0] w_n577_0;
	wire[2:0] w_n578_0;
	wire[1:0] w_n578_1;
	wire[2:0] w_n579_0;
	wire[1:0] w_n580_0;
	wire[1:0] w_n581_0;
	wire[2:0] w_n583_0;
	wire[1:0] w_n583_1;
	wire[2:0] w_n584_0;
	wire[1:0] w_n585_0;
	wire[1:0] w_n586_0;
	wire[2:0] w_n588_0;
	wire[1:0] w_n588_1;
	wire[2:0] w_n589_0;
	wire[1:0] w_n589_1;
	wire[1:0] w_n591_0;
	wire[1:0] w_n592_0;
	wire[1:0] w_n599_0;
	wire[1:0] w_n605_0;
	wire[2:0] w_n606_0;
	wire[2:0] w_n606_1;
	wire[1:0] w_n607_0;
	wire[2:0] w_n608_0;
	wire[1:0] w_n610_0;
	wire[1:0] w_n612_0;
	wire[2:0] w_n613_0;
	wire[2:0] w_n615_0;
	wire[1:0] w_n615_1;
	wire[1:0] w_n617_0;
	wire[2:0] w_n618_0;
	wire[1:0] w_n619_0;
	wire[1:0] w_n620_0;
	wire[2:0] w_n621_0;
	wire[2:0] w_n622_0;
	wire[1:0] w_n622_1;
	wire[2:0] w_n623_0;
	wire[1:0] w_n624_0;
	wire[2:0] w_n625_0;
	wire[1:0] w_n626_0;
	wire[1:0] w_n627_0;
	wire[1:0] w_n628_0;
	wire[1:0] w_n629_0;
	wire[2:0] w_n630_0;
	wire[1:0] w_n631_0;
	wire[1:0] w_n632_0;
	wire[1:0] w_n633_0;
	wire[2:0] w_n634_0;
	wire[2:0] w_n635_0;
	wire[1:0] w_n637_0;
	wire[1:0] w_n642_0;
	wire[1:0] w_n643_0;
	wire[2:0] w_n645_0;
	wire[1:0] w_n647_0;
	wire[2:0] w_n648_0;
	wire[1:0] w_n649_0;
	wire[1:0] w_n650_0;
	wire[1:0] w_n652_0;
	wire[2:0] w_n653_0;
	wire[1:0] w_n653_1;
	wire[1:0] w_n656_0;
	wire[2:0] w_n657_0;
	wire[1:0] w_n657_1;
	wire[2:0] w_n658_0;
	wire[1:0] w_n659_0;
	wire[2:0] w_n660_0;
	wire[1:0] w_n660_1;
	wire[1:0] w_n661_0;
	wire[2:0] w_n662_0;
	wire[1:0] w_n663_0;
	wire[2:0] w_n664_0;
	wire[1:0] w_n664_1;
	wire[2:0] w_n665_0;
	wire[1:0] w_n666_0;
	wire[1:0] w_n667_0;
	wire[2:0] w_n668_0;
	wire[2:0] w_n669_0;
	wire[1:0] w_n671_0;
	wire[1:0] w_n672_0;
	wire[2:0] w_n673_0;
	wire[2:0] w_n674_0;
	wire[1:0] w_n674_1;
	wire[2:0] w_n675_0;
	wire[1:0] w_n676_0;
	wire[2:0] w_n677_0;
	wire[2:0] w_n678_0;
	wire[2:0] w_n679_0;
	wire[1:0] w_n679_1;
	wire[1:0] w_n680_0;
	wire[1:0] w_n683_0;
	wire[1:0] w_n686_0;
	wire[1:0] w_n687_0;
	wire[1:0] w_n690_0;
	wire[1:0] w_n692_0;
	wire[1:0] w_n693_0;
	wire[2:0] w_n697_0;
	wire[2:0] w_n699_0;
	wire[1:0] w_n699_1;
	wire[2:0] w_n701_0;
	wire[1:0] w_n701_1;
	wire[1:0] w_n703_0;
	wire[1:0] w_n704_0;
	wire[1:0] w_n705_0;
	wire[2:0] w_n707_0;
	wire[1:0] w_n708_0;
	wire[2:0] w_n709_0;
	wire[1:0] w_n709_1;
	wire[1:0] w_n710_0;
	wire[1:0] w_n711_0;
	wire[1:0] w_n712_0;
	wire[2:0] w_n713_0;
	wire[1:0] w_n713_1;
	wire[1:0] w_n714_0;
	wire[2:0] w_n715_0;
	wire[2:0] w_n716_0;
	wire[1:0] w_n716_1;
	wire[2:0] w_n720_0;
	wire[1:0] w_n720_1;
	wire[2:0] w_n723_0;
	wire[2:0] w_n727_0;
	wire[1:0] w_n728_0;
	wire[2:0] w_n730_0;
	wire[2:0] w_n734_0;
	wire[1:0] w_n735_0;
	wire[2:0] w_n737_0;
	wire[2:0] w_n741_0;
	wire[1:0] w_n742_0;
	wire[2:0] w_n744_0;
	wire[2:0] w_n748_0;
	wire[1:0] w_n751_0;
	wire[1:0] w_n752_0;
	wire[2:0] w_n754_0;
	wire[2:0] w_n758_0;
	wire[1:0] w_n759_0;
	wire[1:0] w_n764_0;
	wire[1:0] w_n765_0;
	wire[1:0] w_n782_0;
	wire[2:0] w_n784_0;
	wire[2:0] w_n787_0;
	wire[2:0] w_n790_0;
	wire[1:0] w_n790_1;
	wire[2:0] w_n793_0;
	wire[1:0] w_n793_1;
	wire[1:0] w_n795_0;
	wire[2:0] w_n797_0;
	wire[1:0] w_n797_1;
	wire[2:0] w_n801_0;
	wire[1:0] w_n801_1;
	wire[1:0] w_n802_0;
	wire[2:0] w_n804_0;
	wire[2:0] w_n807_0;
	wire[2:0] w_n810_0;
	wire[2:0] w_n812_0;
	wire[2:0] w_n816_0;
	wire[1:0] w_n817_0;
	wire[2:0] w_n819_0;
	wire[2:0] w_n823_0;
	wire[1:0] w_n824_0;
	wire[2:0] w_n827_0;
	wire[2:0] w_n831_0;
	wire[1:0] w_n832_0;
	wire[1:0] w_n834_0;
	wire[1:0] w_n838_0;
	wire[2:0] w_n843_0;
	wire[2:0] w_n847_0;
	wire[1:0] w_n848_0;
	wire[2:0] w_n851_0;
	wire[2:0] w_n855_0;
	wire[1:0] w_n856_0;
	wire[2:0] w_n858_0;
	wire[1:0] w_n859_0;
	wire[1:0] w_n864_0;
	wire[1:0] w_n865_0;
	wire[2:0] w_n869_0;
	wire[2:0] w_n873_0;
	wire[1:0] w_n874_0;
	wire[2:0] w_n878_0;
	wire[2:0] w_n882_0;
	wire[1:0] w_n885_0;
	wire[1:0] w_n887_0;
	wire[1:0] w_n889_0;
	wire[2:0] w_n891_0;
	wire[1:0] w_n891_1;
	wire[2:0] w_n895_0;
	wire[1:0] w_n895_1;
	wire[1:0] w_n896_0;
	wire[2:0] w_n899_0;
	wire[2:0] w_n902_0;
	wire[2:0] w_n905_0;
	wire[2:0] w_n908_0;
	wire[2:0] w_n912_0;
	wire[1:0] w_n913_0;
	wire[2:0] w_n916_0;
	wire[2:0] w_n920_0;
	wire[1:0] w_n921_0;
	wire[1:0] w_n923_0;
	wire[2:0] w_n927_0;
	wire[2:0] w_n931_0;
	wire[1:0] w_n932_0;
	wire[1:0] w_n935_0;
	wire[1:0] w_n937_0;
	wire[1:0] w_n939_0;
	wire[2:0] w_n945_0;
	wire[1:0] w_n945_1;
	wire[2:0] w_n948_0;
	wire[1:0] w_n948_1;
	wire[1:0] w_n950_0;
	wire[1:0] w_n952_0;
	wire[1:0] w_n957_0;
	wire[1:0] w_n972_0;
	wire[1:0] w_n981_0;
	wire[1:0] w_n987_0;
	wire[2:0] w_n988_0;
	wire[2:0] w_n992_0;
	wire[1:0] w_n993_0;
	wire[1:0] w_n994_0;
	wire[2:0] w_n995_0;
	wire[2:0] w_n999_0;
	wire[1:0] w_n1000_0;
	wire[1:0] w_n1003_0;
	wire[1:0] w_n1007_0;
	wire[1:0] w_n1008_0;
	wire[2:0] w_n1009_0;
	wire[1:0] w_n1009_1;
	wire[2:0] w_n1013_0;
	wire[1:0] w_n1013_1;
	wire[1:0] w_n1014_0;
	wire[1:0] w_n1015_0;
	wire[2:0] w_n1016_0;
	wire[2:0] w_n1019_0;
	wire[1:0] w_n1022_0;
	wire[1:0] w_n1033_0;
	wire[1:0] w_n1044_0;
	wire[2:0] w_n1061_0;
	wire[1:0] w_n1062_0;
	wire[2:0] w_n1066_0;
	wire[1:0] w_n1068_0;
	wire[1:0] w_n1069_0;
	wire[2:0] w_n1073_0;
	wire[1:0] w_n1075_0;
	wire[1:0] w_n1076_0;
	wire[2:0] w_n1077_0;
	wire[2:0] w_n1081_0;
	wire[1:0] w_n1082_0;
	wire[2:0] w_n1086_0;
	wire[1:0] w_n1092_0;
	wire[1:0] w_n1095_0;
	wire[2:0] w_n1096_0;
	wire[2:0] w_n1100_0;
	wire[1:0] w_n1102_0;
	wire[1:0] w_n1104_0;
	wire[1:0] w_n1105_0;
	wire[1:0] w_n1116_0;
	wire[2:0] w_n1122_0;
	wire[2:0] w_n1125_0;
	wire[1:0] w_n1127_0;
	wire[2:0] w_n1128_0;
	wire[1:0] w_n1128_1;
	wire[1:0] w_n1130_0;
	wire[1:0] w_n1136_0;
	wire[1:0] w_n1142_0;
	wire[2:0] w_n1148_0;
	wire[1:0] w_n1156_0;
	wire[1:0] w_n1166_0;
	wire[1:0] w_n1173_0;
	wire[1:0] w_n1189_0;
	wire[1:0] w_n1205_0;
	wire[1:0] w_n1236_0;
	wire[1:0] w_n1244_0;
	wire[1:0] w_n1283_0;
	wire[1:0] w_n1301_0;
	wire[1:0] w_n1309_0;
	wire[1:0] w_n1317_0;
	wire[1:0] w_n1325_0;
	wire[2:0] w_n1359_0;
	wire[2:0] w_n1360_0;
	wire[1:0] w_n1360_1;
	wire[1:0] w_n1361_0;
	wire[1:0] w_n1362_0;
	wire[1:0] w_n1376_0;
	wire[2:0] w_n1380_0;
	wire[1:0] w_n1380_1;
	wire[2:0] w_n1383_0;
	wire[2:0] w_n1383_1;
	wire[2:0] w_n1385_0;
	wire[1:0] w_n1385_1;
	wire[2:0] w_n1389_0;
	wire[1:0] w_n1389_1;
	wire[2:0] w_n1392_0;
	wire[1:0] w_n1392_1;
	wire[1:0] w_n1401_0;
	wire[1:0] w_n1402_0;
	wire[1:0] w_n1403_0;
	wire[1:0] w_n1404_0;
	wire[1:0] w_n1405_0;
	wire[1:0] w_n1406_0;
	wire[1:0] w_n1414_0;
	wire[2:0] w_n1420_0;
	wire[1:0] w_n1421_0;
	wire[1:0] w_n1422_0;
	wire[1:0] w_n1424_0;
	wire[1:0] w_n1425_0;
	wire[2:0] w_n1444_0;
	wire[1:0] w_n1445_0;
	wire[1:0] w_n1447_0;
	wire[1:0] w_n1454_0;
	wire[2:0] w_n1463_0;
	wire[1:0] w_n1464_0;
	wire[1:0] w_n1465_0;
	wire[1:0] w_n1468_0;
	wire[1:0] w_n1469_0;
	wire[1:0] w_n1470_0;
	wire[1:0] w_n1471_0;
	wire[1:0] w_n1472_0;
	wire[1:0] w_n1473_0;
	wire[1:0] w_n1479_0;
	wire[1:0] w_n1482_0;
	wire[1:0] w_n1486_0;
	wire[2:0] w_n1494_0;
	wire[1:0] w_n1501_0;
	wire[1:0] w_n1510_0;
	wire[1:0] w_n1520_0;
	wire[1:0] w_n1536_0;
	wire[1:0] w_n1571_0;
	wire[1:0] w_n1599_0;
	wire[1:0] w_n1610_0;
	wire[1:0] w_n1611_0;
	wire[1:0] w_n1625_0;
	wire[1:0] w_n1642_0;
	wire[1:0] w_n1644_0;
	wire[1:0] w_n1651_0;
	wire[1:0] w_n1654_0;
	wire[1:0] w_n1659_0;
	wire[1:0] w_n1667_0;
	wire[1:0] w_n1670_0;
	wire[1:0] w_n1672_0;
	wire[1:0] w_n1675_0;
	wire[1:0] w_n1680_0;
	wire[1:0] w_n1687_0;
	wire[1:0] w_n1689_0;
	wire[1:0] w_n1699_0;
	wire w_dff_A_Pos9QPwV7_0;
	wire w_dff_A_XGfauPzp1_0;
	wire w_dff_A_IEvszadD0_1;
	wire w_dff_A_HjETiJKP7_1;
	wire w_dff_A_tdRIK4cs5_1;
	wire w_dff_A_QndkNCew9_2;
	wire w_dff_B_wgDSXUDG2_0;
	wire w_dff_B_fWyqtvR81_3;
	wire w_dff_B_uoINvDSa8_3;
	wire w_dff_B_WTbhWZhI7_3;
	wire w_dff_B_7QJvHfSv5_3;
	wire w_dff_B_uGCHlJxK9_3;
	wire w_dff_B_kbXJdWzf8_3;
	wire w_dff_B_gTpgSbmF2_3;
	wire w_dff_B_gsg21ktp1_3;
	wire w_dff_B_nHZK4yve1_3;
	wire w_dff_B_htnMHrbg4_3;
	wire w_dff_B_q1wIQwTM4_3;
	wire w_dff_B_NwX8w6Vb0_3;
	wire w_dff_B_dJxNXdWa0_3;
	wire w_dff_B_qfU08Cof6_3;
	wire w_dff_B_nI1NuC2F0_3;
	wire w_dff_B_0iF05mWz2_3;
	wire w_dff_B_lqJRKDNW7_1;
	wire w_dff_B_KC1varD37_0;
	wire w_dff_B_N91gti7d4_0;
	wire w_dff_B_xXyVJF5x1_0;
	wire w_dff_B_zF2G5PQf4_0;
	wire w_dff_B_3IxjCjfR7_0;
	wire w_dff_B_1glBVTOx1_0;
	wire w_dff_B_eowfTFGQ0_0;
	wire w_dff_B_TR8eBgc44_0;
	wire w_dff_B_uEgPLN9I8_0;
	wire w_dff_B_4g0KHQgb9_0;
	wire w_dff_B_UVTHnIgH5_0;
	wire w_dff_B_C5muFh6p3_0;
	wire w_dff_B_DZE264KT4_0;
	wire w_dff_B_SFE4sIHa2_0;
	wire w_dff_B_pZAfrZYo5_0;
	wire w_dff_B_mTKgg1164_0;
	wire w_dff_B_L2KMdVHu3_0;
	wire w_dff_B_ryF06tMX0_0;
	wire w_dff_B_ipbujmWF3_0;
	wire w_dff_B_RiW4jPHy1_0;
	wire w_dff_B_w1tGP8yo3_0;
	wire w_dff_B_5EDT2rnP2_1;
	wire w_dff_B_PhMNAOfy1_1;
	wire w_dff_B_V9LgDelO6_1;
	wire w_dff_A_2H7UVBdK3_1;
	wire w_dff_A_dK8hF1rC4_0;
	wire w_dff_A_XgMhCSMX3_0;
	wire w_dff_A_YNttyCCi4_0;
	wire w_dff_B_bVaJ0Cf89_0;
	wire w_dff_B_gOANsO7i2_0;
	wire w_dff_B_xeUFODug7_0;
	wire w_dff_B_xlePdhEl3_0;
	wire w_dff_B_Gc98jEYO0_0;
	wire w_dff_B_wkkZXIpM0_0;
	wire w_dff_B_ySOYDXTl2_0;
	wire w_dff_B_RKBX27OC2_0;
	wire w_dff_B_vrsafaGC8_0;
	wire w_dff_B_ApusimQ42_0;
	wire w_dff_A_bNXtfWRE3_1;
	wire w_dff_A_kAEMKNcT9_1;
	wire w_dff_A_koKZi9Uv9_1;
	wire w_dff_A_uBfCaew78_1;
	wire w_dff_A_YYyzousl5_1;
	wire w_dff_A_ReZ75tPd8_1;
	wire w_dff_B_tB2GeuHj0_2;
	wire w_dff_B_MTWo24nU6_0;
	wire w_dff_B_AMOHr3Vf6_0;
	wire w_dff_B_n58IivwY1_0;
	wire w_dff_A_EYKd06HK4_0;
	wire w_dff_A_pYjNPTOh3_0;
	wire w_dff_A_14yKmCqw2_1;
	wire w_dff_B_afESf26d0_1;
	wire w_dff_B_SC8tEvs74_1;
	wire w_dff_B_234lh4O68_1;
	wire w_dff_B_9kGRiarq1_1;
	wire w_dff_B_RDXZWQRJ4_0;
	wire w_dff_B_dJjfIWKK6_0;
	wire w_dff_A_lYcNZSyi0_1;
	wire w_dff_A_ZKFrcWGh3_1;
	wire w_dff_A_RJt6C40d5_1;
	wire w_dff_A_Q9txt8M98_1;
	wire w_dff_A_Mf0742Hd8_1;
	wire w_dff_B_MDMrVRml4_1;
	wire w_dff_B_GYqy8mHM6_0;
	wire w_dff_B_JeT5s1nr0_0;
	wire w_dff_B_lzCG9mPr6_0;
	wire w_dff_B_374cMAJc9_0;
	wire w_dff_A_SSZO0uzt5_0;
	wire w_dff_A_qkOoyJRf5_0;
	wire w_dff_A_tR9lgU7T7_1;
	wire w_dff_A_ekM6GQ1p6_1;
	wire w_dff_A_gnYb3llh5_1;
	wire w_dff_A_yzHYW8jW8_1;
	wire w_dff_B_NqZ7nwu76_2;
	wire w_dff_A_E9LU2zbd2_1;
	wire w_dff_A_4eqkkdOn0_1;
	wire w_dff_A_atfaHIcj9_1;
	wire w_dff_A_x53jfDaD6_1;
	wire w_dff_B_gdK7QGUf4_2;
	wire w_dff_B_2CyjtYCN9_1;
	wire w_dff_B_NZtnnIIa5_1;
	wire w_dff_B_tkcTmpq62_1;
	wire w_dff_B_T7vY4eHE7_1;
	wire w_dff_B_oqO2spPR1_0;
	wire w_dff_B_CNs4IfNm6_0;
	wire w_dff_B_P5WZjbkc1_0;
	wire w_dff_B_4d4R3abv3_1;
	wire w_dff_B_bSGiMxoB1_1;
	wire w_dff_B_5qNLIagO9_1;
	wire w_dff_B_Maxmj71J6_1;
	wire w_dff_B_FVzcyAbF7_1;
	wire w_dff_B_lgvf0JUe6_1;
	wire w_dff_B_qOY9c4NC0_1;
	wire w_dff_B_2JkFxvEv9_1;
	wire w_dff_B_AN0P4XMB2_1;
	wire w_dff_B_mI1w0mBq3_1;
	wire w_dff_B_Yi2ITFyq1_1;
	wire w_dff_A_7pUNrHii4_0;
	wire w_dff_B_LEyrmZNw7_1;
	wire w_dff_A_ze6hIAz33_1;
	wire w_dff_A_DrbNfpRo1_0;
	wire w_dff_B_INOoEPE86_3;
	wire w_dff_B_2p6vx4go2_0;
	wire w_dff_B_Uh0Dhd3p5_0;
	wire w_dff_A_rwP99a5q0_0;
	wire w_dff_B_kXm7rX3S9_2;
	wire w_dff_B_N1uTPie67_0;
	wire w_dff_B_wtZEieFg8_0;
	wire w_dff_B_w8MyrbaO0_0;
	wire w_dff_B_XbHFmXLl3_0;
	wire w_dff_B_0ybnmimc7_0;
	wire w_dff_B_qVKgIB5E4_2;
	wire w_dff_A_oK3vFRv77_1;
	wire w_dff_B_CJYLLkVd5_0;
	wire w_dff_A_XaL3CtiK4_0;
	wire w_dff_A_g9V4GvzL7_0;
	wire w_dff_A_RD61e9T25_0;
	wire w_dff_A_MoDIOIRi2_0;
	wire w_dff_A_tWV56WJ98_0;
	wire w_dff_A_j8FtofYP3_0;
	wire w_dff_B_HHy6QElJ5_1;
	wire w_dff_B_MLNtxgJY4_1;
	wire w_dff_B_2ir4DjU72_0;
	wire w_dff_B_C3rdXGV10_1;
	wire w_dff_A_bO3nzByT2_0;
	wire w_dff_A_ajdf93iQ9_0;
	wire w_dff_A_AgAEvzEB1_0;
	wire w_dff_A_9AfuIthu8_0;
	wire w_dff_A_Mdj67B3H9_0;
	wire w_dff_A_7YvRhIar6_0;
	wire w_dff_B_pxRVTx135_0;
	wire w_dff_A_wUpRfK0p1_0;
	wire w_dff_A_rALwFiav9_2;
	wire w_dff_A_uObGZouh4_1;
	wire w_dff_A_kvQeBA0D2_0;
	wire w_dff_A_4IEJ6hOt6_0;
	wire w_dff_A_q9dCrBA79_0;
	wire w_dff_A_vhkzGJZA8_0;
	wire w_dff_A_RJjKOlTb6_0;
	wire w_dff_A_lonv2OjE2_0;
	wire w_dff_A_BAORIDP98_0;
	wire w_dff_A_aZDu4bpW2_0;
	wire w_dff_A_sbM22p8l0_2;
	wire w_dff_B_Lt3ej8b54_3;
	wire w_dff_B_7O3vY0Tl6_3;
	wire w_dff_A_GjdtnPFR2_0;
	wire w_dff_A_OV1iY6yU0_0;
	wire w_dff_A_BPA1aUZG7_0;
	wire w_dff_A_vv33bzPQ6_0;
	wire w_dff_A_aH6FkRrb9_0;
	wire w_dff_A_vpyBiBU25_0;
	wire w_dff_A_zhxyA46L1_0;
	wire w_dff_B_sHtAJ7Vc2_2;
	wire w_dff_B_Ub74zJxg8_1;
	wire w_dff_B_3dEfFBv87_1;
	wire w_dff_B_GRMGV4p45_1;
	wire w_dff_A_sYrWn1lF6_0;
	wire w_dff_B_5UkBZUQG5_2;
	wire w_dff_B_Lx68BShZ5_2;
	wire w_dff_B_BalxW1tI9_2;
	wire w_dff_B_5uR70sS67_2;
	wire w_dff_B_r7oTZR028_2;
	wire w_dff_B_bCdNpCG38_2;
	wire w_dff_B_1606UYPJ6_2;
	wire w_dff_B_0tVqPFTC9_2;
	wire w_dff_B_3opfKOob2_2;
	wire w_dff_B_hafqao8N8_2;
	wire w_dff_B_8Nc6R9i03_2;
	wire w_dff_B_AiAGUhmX1_2;
	wire w_dff_B_AUYeWQXa8_2;
	wire w_dff_A_S1cGnyRj8_0;
	wire w_dff_B_746NndkO3_2;
	wire w_dff_B_ytwst5vl8_2;
	wire w_dff_B_x7fUxwPR6_2;
	wire w_dff_B_aB5VuoxX1_2;
	wire w_dff_B_5EYh9UZe2_2;
	wire w_dff_B_W1OiaX8U2_2;
	wire w_dff_B_CqLy1fsw5_2;
	wire w_dff_B_LGxucHPi1_2;
	wire w_dff_B_LYL7E7sq7_2;
	wire w_dff_B_np24wlFa0_2;
	wire w_dff_B_vVWifAh97_2;
	wire w_dff_B_uPWYFGOB2_2;
	wire w_dff_B_5khcQBDh4_1;
	wire w_dff_B_OcWJQwsh7_1;
	wire w_dff_B_Mkf1omzt6_1;
	wire w_dff_B_I9yQ9RFt1_1;
	wire w_dff_B_wuRRRZup3_1;
	wire w_dff_B_zAvWvozQ3_1;
	wire w_dff_B_EBsxEAGr1_1;
	wire w_dff_B_u8elYLWU8_1;
	wire w_dff_B_u1ar03Fe3_1;
	wire w_dff_B_lWOZhuri6_1;
	wire w_dff_B_vLvoP0xY1_1;
	wire w_dff_B_wHaSt9t09_1;
	wire w_dff_A_T00sBlkf8_0;
	wire w_dff_B_dAJRi7KG0_2;
	wire w_dff_B_J5IjTRTA3_2;
	wire w_dff_B_8MXUWefQ3_2;
	wire w_dff_B_BvOQF7Do1_2;
	wire w_dff_B_20Yr7Jtx5_2;
	wire w_dff_B_jRDqtOyY5_2;
	wire w_dff_B_ngA7dIag5_2;
	wire w_dff_B_jz2kvfDP2_2;
	wire w_dff_B_eDlhJ25O6_2;
	wire w_dff_B_bRoaWIUD0_2;
	wire w_dff_B_Ce5B3vS49_2;
	wire w_dff_B_QvM587fe2_2;
	wire w_dff_B_n5UtTM7n8_2;
	wire w_dff_B_4itl8JOs0_2;
	wire w_dff_B_rpvwD1GV5_2;
	wire w_dff_B_gPVNGtcT7_2;
	wire w_dff_B_RFmgFe5b7_2;
	wire w_dff_B_CtWkk8hY4_1;
	wire w_dff_B_0x2VHRbv1_1;
	wire w_dff_B_NXHes7CG4_1;
	wire w_dff_B_I7Upk33g6_1;
	wire w_dff_B_dAjkBzzb0_1;
	wire w_dff_B_iK0ZXs7J2_1;
	wire w_dff_B_3q7MxW0d0_1;
	wire w_dff_B_02u2SS0A2_1;
	wire w_dff_B_0LIEmeDZ2_1;
	wire w_dff_B_p37xndZ06_1;
	wire w_dff_B_YG5cchkR7_1;
	wire w_dff_B_BVxSmfl52_1;
	wire w_dff_B_PYxL9Co86_1;
	wire w_dff_B_XisaLX904_0;
	wire w_dff_B_q9YFTezs7_0;
	wire w_dff_B_w2up1oTz5_0;
	wire w_dff_B_wmBPS0CK8_0;
	wire w_dff_B_JVLeYO0G3_0;
	wire w_dff_B_bTJhcQWi8_0;
	wire w_dff_B_dYISN1vL1_0;
	wire w_dff_B_sDosGpL87_0;
	wire w_dff_B_YofwYuaG2_0;
	wire w_dff_B_sDdFbHZ11_0;
	wire w_dff_B_FlHUG2RS1_0;
	wire w_dff_B_CvdsZYuR1_0;
	wire w_dff_B_mt8eOiKy4_0;
	wire w_dff_B_PUHfyred4_0;
	wire w_dff_A_fzo1EyOA9_0;
	wire w_dff_B_MOoZF4NQ8_2;
	wire w_dff_B_4HTsDXSe4_2;
	wire w_dff_B_z5dpkfli4_2;
	wire w_dff_B_xWmAT5HH3_2;
	wire w_dff_B_87SFmAYK4_2;
	wire w_dff_B_hLpvyjlw0_2;
	wire w_dff_B_ix3vso725_2;
	wire w_dff_B_6gkSW4iq7_2;
	wire w_dff_B_HVV2WRDk6_2;
	wire w_dff_B_jp264nbJ3_2;
	wire w_dff_B_94YtK0fd1_2;
	wire w_dff_B_KFMkvf9j7_2;
	wire w_dff_B_ZEbX4XJv2_2;
	wire w_dff_B_CzMhrrsW6_2;
	wire w_dff_B_TsEdxkGT1_2;
	wire w_dff_B_yF9TZLdu0_2;
	wire w_dff_B_hCYdVrMU3_0;
	wire w_dff_B_zZmEURSA8_0;
	wire w_dff_B_EO7nhuqW7_0;
	wire w_dff_B_Myj1SZaj4_0;
	wire w_dff_B_Qk0SAoBB3_0;
	wire w_dff_B_pwXohnk63_0;
	wire w_dff_B_bln28hL01_0;
	wire w_dff_B_RWA6pG1u7_0;
	wire w_dff_B_PXNiVJ5t5_0;
	wire w_dff_B_MqGAPJKl8_1;
	wire w_dff_B_jid7V4CH7_1;
	wire w_dff_B_BBu6uxmD6_0;
	wire w_dff_B_7gLDT3bK5_1;
	wire w_dff_B_3eoJBKu19_1;
	wire w_dff_B_3mrAU2E69_1;
	wire w_dff_B_o2vmRTrk6_1;
	wire w_dff_B_9mCP92cT2_1;
	wire w_dff_B_kRuQ7SBN6_1;
	wire w_dff_B_h5HuSvVj9_1;
	wire w_dff_B_wiKNmkLb3_1;
	wire w_dff_B_hMQE5yCy6_1;
	wire w_dff_B_WsO6eCcY2_1;
	wire w_dff_B_1PUvQFvx8_1;
	wire w_dff_B_RLt04rw04_1;
	wire w_dff_B_KvbD5UbJ4_0;
	wire w_dff_B_DMTwZLiq9_0;
	wire w_dff_B_S8pldWix3_1;
	wire w_dff_B_zn8jTR373_1;
	wire w_dff_B_gkcq18WH8_1;
	wire w_dff_B_vpusSyN26_1;
	wire w_dff_B_S0kEqjWA1_1;
	wire w_dff_B_ffWWzdU89_1;
	wire w_dff_B_hEFGgJ5U5_1;
	wire w_dff_B_vpv4Ip8T8_1;
	wire w_dff_B_lOTosTFb6_0;
	wire w_dff_B_RolcQy8L8_0;
	wire w_dff_B_SziSQuS05_0;
	wire w_dff_B_9Wcolvdi7_0;
	wire w_dff_B_pgKwBpz86_0;
	wire w_dff_B_m95GODcv4_0;
	wire w_dff_B_kKkyU2GE6_0;
	wire w_dff_B_MNnsejKZ3_1;
	wire w_dff_B_AeVhvwdi6_1;
	wire w_dff_B_OXiC4uOZ9_1;
	wire w_dff_B_K95d2xDO4_1;
	wire w_dff_B_n5d7e1jm1_1;
	wire w_dff_B_8iWpoCgo4_1;
	wire w_dff_B_cMeKLzGs4_0;
	wire w_dff_B_geTJlya88_0;
	wire w_dff_B_2f6GBAe88_0;
	wire w_dff_B_YIasQm2p8_0;
	wire w_dff_B_L2o6AYYH5_0;
	wire w_dff_B_6oUft6vE8_0;
	wire w_dff_B_RzSElG5A5_0;
	wire w_dff_B_89KUHvEO0_0;
	wire w_dff_B_S4p4rGHS7_0;
	wire w_dff_B_QPrMLEMA6_0;
	wire w_dff_B_pSeVm3Mk5_0;
	wire w_dff_A_tL4pS8RP3_0;
	wire w_dff_B_ymWx1Ohc5_0;
	wire w_dff_B_EQiSFkrb1_1;
	wire w_dff_B_jGiJQ0wV2_1;
	wire w_dff_B_p992Tqr93_1;
	wire w_dff_B_MovuNc1j0_1;
	wire w_dff_B_dmVOihU45_1;
	wire w_dff_B_pyGI4mB35_0;
	wire w_dff_B_TQzO71He6_0;
	wire w_dff_B_yqqpsv4E3_0;
	wire w_dff_B_oaivzYWu2_0;
	wire w_dff_B_O0Vd6TmT8_0;
	wire w_dff_B_KEa91tD61_0;
	wire w_dff_B_mbOqfH1Y6_0;
	wire w_dff_B_BrXuCZOI4_0;
	wire w_dff_B_bYbZRTHw0_0;
	wire w_dff_B_l4rg2tHX6_0;
	wire w_dff_B_f4DIV2E73_1;
	wire w_dff_B_aYGp1ZGM9_1;
	wire w_dff_B_1bITEiIi8_1;
	wire w_dff_B_fbU8G7Lj5_0;
	wire w_dff_B_tmteiliS8_0;
	wire w_dff_A_cGZBiJwI7_1;
	wire w_dff_B_SoIl8LzQ8_0;
	wire w_dff_B_y2lQnTGk1_0;
	wire w_dff_B_DeWSW7nC9_0;
	wire w_dff_B_fQnMEHd96_0;
	wire w_dff_B_3kyWkG664_0;
	wire w_dff_B_dahXD1oR3_0;
	wire w_dff_B_jPTP5tlu9_0;
	wire w_dff_B_VrqhbXKF4_0;
	wire w_dff_B_HOoNpVCD2_0;
	wire w_dff_B_KyMlupGs9_0;
	wire w_dff_B_XSsA1Wql7_0;
	wire w_dff_B_lOMOsdSt8_0;
	wire w_dff_B_PWdaVupe0_0;
	wire w_dff_A_Hqdbi7JV4_1;
	wire w_dff_B_0CT38OSx1_0;
	wire w_dff_B_54cKlWns1_0;
	wire w_dff_B_PST0blmv8_0;
	wire w_dff_B_CXnBBQwP6_0;
	wire w_dff_A_48ZOUHfV8_0;
	wire w_dff_A_CwlY1HgX1_0;
	wire w_dff_B_Wf7nYgeZ5_0;
	wire w_dff_B_q7BVBUQk7_1;
	wire w_dff_B_nrWiBURo9_0;
	wire w_dff_B_EqwYgOAb4_0;
	wire w_dff_B_NZouYTI96_0;
	wire w_dff_B_sSfu5jc82_0;
	wire w_dff_A_ETdALzzl9_2;
	wire w_dff_A_jvMIQD1H6_2;
	wire w_dff_A_IHi45kUJ0_0;
	wire w_dff_A_jdynXXo00_0;
	wire w_dff_B_P7acJj6O5_0;
	wire w_dff_A_z9rFL9Qs7_0;
	wire w_dff_A_l1Fd4mzB7_0;
	wire w_dff_B_go3tZ8237_0;
	wire w_dff_A_eOGCc9MY9_0;
	wire w_dff_A_xmqyPieu1_1;
	wire w_dff_B_SaZRZ3eC7_1;
	wire w_dff_B_BBcmIffi9_0;
	wire w_dff_A_DPI265385_0;
	wire w_dff_B_wyRCCiEu4_0;
	wire w_dff_A_mVf8HqKT3_0;
	wire w_dff_A_Rudi88Ma5_0;
	wire w_dff_A_3oTeT6Q66_0;
	wire w_dff_B_MoBmqS1O8_1;
	wire w_dff_B_XgTx141R4_1;
	wire w_dff_B_eKyjidAx3_0;
	wire w_dff_B_tHgUzJFw0_0;
	wire w_dff_B_5Z0ZvisL2_0;
	wire w_dff_B_AtF61fDY2_1;
	wire w_dff_B_FCQlh5Dj1_0;
	wire w_dff_B_ImjzZV4d2_0;
	wire w_dff_A_hwfUxLGL7_1;
	wire w_dff_B_Dv298iPP6_0;
	wire w_dff_B_a2d6WJsL9_0;
	wire w_dff_B_JiLRwsqs5_0;
	wire w_dff_B_k7lL40703_0;
	wire w_dff_A_HTROHZQK8_0;
	wire w_dff_A_fbjRGt6H7_0;
	wire w_dff_B_k7AAB8Kr6_0;
	wire w_dff_B_G3fOBOAh3_1;
	wire w_dff_B_aSMhC8VD8_0;
	wire w_dff_B_MZwE7jgl3_0;
	wire w_dff_B_rcYx8yKf4_0;
	wire w_dff_A_dYIGB10U4_0;
	wire w_dff_B_0yBXJo9z0_0;
	wire w_dff_A_Uh6msUUb7_0;
	wire w_dff_B_L7t6hzka9_0;
	wire w_dff_B_H2CRhkLX8_1;
	wire w_dff_B_ji1kzFuV4_0;
	wire w_dff_B_eTd8rISp4_0;
	wire w_dff_A_xh58VgyV7_1;
	wire w_dff_B_GwnOSJim7_1;
	wire w_dff_B_1lI4iuCx7_1;
	wire w_dff_B_vQSB5hO77_1;
	wire w_dff_B_QHRDrX0e1_1;
	wire w_dff_B_ovWBiHve8_1;
	wire w_dff_A_ABytohFn0_1;
	wire w_dff_A_Voxo0vv56_2;
	wire w_dff_B_v0d9Pcq65_1;
	wire w_dff_B_RvBlhviK6_1;
	wire w_dff_A_kfTwIkQA1_1;
	wire w_dff_A_wlzDAiYg7_2;
	wire w_dff_B_O5SW7v0n6_1;
	wire w_dff_A_kZe7phSE5_1;
	wire w_dff_A_q50Fv1v73_2;
	wire w_dff_B_NDxgaqFP7_1;
	wire w_dff_A_ENCyuXag9_1;
	wire w_dff_A_2yNquiOy5_2;
	wire w_dff_B_fGFTF0XU1_1;
	wire w_dff_A_SZuNFr1P2_0;
	wire w_dff_A_4oRPwfXE4_2;
	wire w_dff_B_pi3wdSqF9_1;
	wire w_dff_A_OL2RzQCe5_1;
	wire w_dff_A_GNJJtZnm1_2;
	wire w_dff_B_NrCPywIU0_1;
	wire w_dff_A_JJ89itmx3_0;
	wire w_dff_A_iQkRFewx6_0;
	wire w_dff_A_dHpbrnif0_1;
	wire w_dff_B_iLWJF1Hp3_3;
	wire w_dff_B_NUpiunu24_1;
	wire w_dff_B_a4N3anBT4_1;
	wire w_dff_B_aLvfeHDS9_1;
	wire w_dff_B_5vCkOg337_1;
	wire w_dff_B_qk2e6yzr7_1;
	wire w_dff_B_763OWH5q8_0;
	wire w_dff_B_FXgMXwFy3_0;
	wire w_dff_A_l640jkIo4_1;
	wire w_dff_A_I9KtYtk61_1;
	wire w_dff_B_6iLd3lGi5_1;
	wire w_dff_B_9UIE7en39_1;
	wire w_dff_B_iKVVTLIe3_1;
	wire w_dff_B_gMghVbHt7_1;
	wire w_dff_B_U64D73rS2_1;
	wire w_dff_B_ME82u0P10_1;
	wire w_dff_A_CC1cSYvL9_0;
	wire w_dff_B_8ePvQrtz7_1;
	wire w_dff_B_AUOibp789_1;
	wire w_dff_B_llGRv8mi5_1;
	wire w_dff_B_IdjBLrfV7_3;
	wire w_dff_B_9BfjA4og5_3;
	wire w_dff_B_pLPjMUlg0_3;
	wire w_dff_B_XBuut1l53_3;
	wire w_dff_B_o7C5KK9Q1_3;
	wire w_dff_B_EJ1wzUhh8_3;
	wire w_dff_B_rhc9L5xJ1_3;
	wire w_dff_B_npBiyaxb7_3;
	wire w_dff_B_y0O2kR962_3;
	wire w_dff_B_MnsduYnO8_3;
	wire w_dff_B_8sbhzKj90_3;
	wire w_dff_B_O3qcBfn54_3;
	wire w_dff_B_0N8uFRUA7_3;
	wire w_dff_B_rMlRfwdG0_3;
	wire w_dff_B_0giEvvrD3_3;
	wire w_dff_B_tMqqm3EM5_3;
	wire w_dff_B_mCDgaTCp3_3;
	wire w_dff_B_Nlr6LKx27_3;
	wire w_dff_B_wwhembUv9_3;
	wire w_dff_B_bzIU7bhA5_3;
	wire w_dff_B_ZKPdG3yj8_3;
	wire w_dff_B_x019fOFD0_1;
	wire w_dff_B_DJUXuzfR5_1;
	wire w_dff_B_2NR1HArv1_1;
	wire w_dff_B_fDvnNcQc3_1;
	wire w_dff_B_x56lNv725_1;
	wire w_dff_B_RdsBE9xP4_1;
	wire w_dff_B_XO3NzWg02_1;
	wire w_dff_B_8iUwmmxU1_1;
	wire w_dff_B_8w6Ejsrg6_1;
	wire w_dff_B_8E6Si50q8_1;
	wire w_dff_B_SWHMzrLs6_1;
	wire w_dff_B_h37MDbom1_1;
	wire w_dff_B_Gwax1Gzy7_1;
	wire w_dff_B_YR4BPWLM1_1;
	wire w_dff_B_qW4ciP0a2_1;
	wire w_dff_B_hvcuFbb39_1;
	wire w_dff_A_QFVvSBXs1_0;
	wire w_dff_A_ovTq2xU49_1;
	wire w_dff_A_Ckj1AOyH1_0;
	wire w_dff_B_TOpau3XT3_2;
	wire w_dff_B_ATBd61GY6_2;
	wire w_dff_B_Mkym6Kci4_2;
	wire w_dff_B_UiM5x9MF9_2;
	wire w_dff_B_yo0imXru5_2;
	wire w_dff_B_7qFPsQRP3_2;
	wire w_dff_B_Jcbt0k3I2_2;
	wire w_dff_B_5sZLto4h2_2;
	wire w_dff_B_La9vFLI37_2;
	wire w_dff_A_cJhQqle97_0;
	wire w_dff_B_LkdWkJ8g7_2;
	wire w_dff_B_1gkzg7R10_2;
	wire w_dff_B_b4mHv3Ng6_2;
	wire w_dff_B_1Kmi0HtZ6_2;
	wire w_dff_B_1Kw8nNbx2_2;
	wire w_dff_B_llMY8War6_2;
	wire w_dff_B_KKg45cXB6_2;
	wire w_dff_B_7PTogLGb4_1;
	wire w_dff_B_jXVjhxPA7_1;
	wire w_dff_B_B0jVdQZK5_1;
	wire w_dff_B_HMC3Mo6w6_1;
	wire w_dff_B_GZoZRhPB5_1;
	wire w_dff_B_zCZ1gWyq6_1;
	wire w_dff_B_MAfprkEt8_1;
	wire w_dff_B_AzlUtPke4_1;
	wire w_dff_B_TwUTlE3B4_1;
	wire w_dff_B_tYZ2TMyR3_1;
	wire w_dff_B_PPbMZT6d2_1;
	wire w_dff_B_FLUsvZJe6_1;
	wire w_dff_B_7es6Sl7R1_1;
	wire w_dff_B_L0aE1pJH9_1;
	wire w_dff_B_mt6EQCSe3_1;
	wire w_dff_B_xkiUoI6d8_0;
	wire w_dff_B_mAKxwxqz1_0;
	wire w_dff_B_fGAAYMSZ9_0;
	wire w_dff_B_RDwCv1ed2_0;
	wire w_dff_B_eATi8HMD6_1;
	wire w_dff_B_oj7vR2wc0_1;
	wire w_dff_B_25NFH76a5_1;
	wire w_dff_B_2ZeCTHMn8_1;
	wire w_dff_B_k7HXkkHM6_1;
	wire w_dff_B_wUzjKcsA2_1;
	wire w_dff_B_XvPI7GAs4_1;
	wire w_dff_B_pnT5QBZn4_1;
	wire w_dff_B_WA4gBXwc1_1;
	wire w_dff_B_nQNILQLi0_1;
	wire w_dff_B_m54To6v88_1;
	wire w_dff_B_wa7J2Vx24_1;
	wire w_dff_B_47O9ffhk8_0;
	wire w_dff_B_H19Doc6T6_1;
	wire w_dff_B_pkJzjAA13_0;
	wire w_dff_A_0RAVFEVr1_1;
	wire w_dff_A_eOyVXiE77_1;
	wire w_dff_A_b8zTXIi13_1;
	wire w_dff_A_sRXZ4qhC5_1;
	wire w_dff_A_Kpy41kBj3_1;
	wire w_dff_A_xghiZztM6_1;
	wire w_dff_A_5uPzxucX4_1;
	wire w_dff_A_IW5KJ3Dj5_1;
	wire w_dff_A_WBXkA0S14_1;
	wire w_dff_A_mxJkPqv15_1;
	wire w_dff_B_bMdm3kIy3_1;
	wire w_dff_A_Q4G3Vr6v2_1;
	wire w_dff_A_5cF9i9ps0_1;
	wire w_dff_A_Fg0GymQ76_1;
	wire w_dff_A_jPMQ1vXE5_1;
	wire w_dff_A_20vVuD9A2_1;
	wire w_dff_A_HLu4tZgU8_1;
	wire w_dff_A_45Mf1pPl0_1;
	wire w_dff_A_LUAz2R5u7_1;
	wire w_dff_A_jOasjh7M6_1;
	wire w_dff_B_pNqP6SDG5_2;
	wire w_dff_B_vAm4i5Er2_0;
	wire w_dff_B_VZarvOZq4_0;
	wire w_dff_B_1sUUPRfg5_0;
	wire w_dff_B_OJow9Vyl2_1;
	wire w_dff_B_U1goTxm30_1;
	wire w_dff_B_QDq6Jaas7_0;
	wire w_dff_B_ordt9V3h7_0;
	wire w_dff_B_jAFUiruS4_0;
	wire w_dff_B_N6gXHevE0_1;
	wire w_dff_A_FzYkVwt71_1;
	wire w_dff_A_Xm39ijup5_1;
	wire w_dff_A_KQjVIlGn5_1;
	wire w_dff_A_4ys7vwfR2_1;
	wire w_dff_A_3TleVXER0_1;
	wire w_dff_A_Apm4yrQa9_1;
	wire w_dff_A_H1VOLBDP6_1;
	wire w_dff_A_hBqkJqjS1_1;
	wire w_dff_A_ZmUqUEXr6_1;
	wire w_dff_B_tlAcGgC34_2;
	wire w_dff_B_YXY9vh597_2;
	wire w_dff_B_uiMlzBmr5_2;
	wire w_dff_B_mBMAvR3y5_2;
	wire w_dff_B_QqnObltz0_2;
	wire w_dff_B_Ypk94iqM7_2;
	wire w_dff_A_trCzAZP81_1;
	wire w_dff_B_XX0mknTh8_0;
	wire w_dff_B_Z4uhcWtN0_0;
	wire w_dff_B_TymWwy7E5_0;
	wire w_dff_B_Qbdzpj2C1_0;
	wire w_dff_B_eiKQTK2w9_0;
	wire w_dff_B_ztIY41Q55_1;
	wire w_dff_B_rbiPKVwW4_1;
	wire w_dff_B_XiJPqNd82_1;
	wire w_dff_B_ra5xCKJj3_1;
	wire w_dff_B_whGYmxuB1_1;
	wire w_dff_B_1qVDS2KB7_1;
	wire w_dff_B_rzNwJKfw7_0;
	wire w_dff_A_RMpuFhPp5_1;
	wire w_dff_A_p5TL9DJ66_1;
	wire w_dff_A_PKoctAc01_1;
	wire w_dff_A_yukqebI99_1;
	wire w_dff_A_YQ5Y2fgs9_1;
	wire w_dff_A_ZWcRm7Km3_1;
	wire w_dff_A_IlyOiMQ73_1;
	wire w_dff_A_w4QdJfPC3_1;
	wire w_dff_A_oGuhTOFj2_1;
	wire w_dff_A_ILt6LRmd0_1;
	wire w_dff_A_sXuwNK8R4_1;
	wire w_dff_B_oKWTF6hl0_2;
	wire w_dff_B_FE7WUiIF0_0;
	wire w_dff_B_idJEKtUL7_0;
	wire w_dff_B_jtp16RiP5_0;
	wire w_dff_B_s88beJ2U6_0;
	wire w_dff_B_b5nqAN7c3_0;
	wire w_dff_B_yIW1yNUH0_0;
	wire w_dff_B_GRpJRWRw0_0;
	wire w_dff_A_OZfn1ucS1_0;
	wire w_dff_A_TA0aTwIG6_0;
	wire w_dff_A_XrdWwc4R2_2;
	wire w_dff_A_JoHABMJ87_2;
	wire w_dff_A_zWjy8oUP2_2;
	wire w_dff_A_8cwtMwTA2_2;
	wire w_dff_A_8qFpqZGO9_2;
	wire w_dff_A_HINHVoHg8_2;
	wire w_dff_A_lI3gZliT6_2;
	wire w_dff_A_bJzo3sLd7_2;
	wire w_dff_A_A17pJVNn5_2;
	wire w_dff_A_uL5Vjebj3_2;
	wire w_dff_A_RijIaEAN0_2;
	wire w_dff_A_s0GIDYHk9_2;
	wire w_dff_A_W0oVwpZc9_2;
	wire w_dff_B_qnMenjZs7_3;
	wire w_dff_B_8ItX7a3K5_3;
	wire w_dff_B_H6Ftr2x54_3;
	wire w_dff_B_nLkcjZeK0_3;
	wire w_dff_A_K8finmwX0_1;
	wire w_dff_A_fCO3Igr54_1;
	wire w_dff_A_uQPGZkEK6_1;
	wire w_dff_A_s5UHIRKd7_1;
	wire w_dff_A_YS3sKKuK9_1;
	wire w_dff_A_dLHHILYu7_1;
	wire w_dff_A_ZLOlZNlP0_1;
	wire w_dff_A_uMZQ4TGC6_1;
	wire w_dff_A_aOg9zfBa6_1;
	wire w_dff_A_Q9N2VMIL7_1;
	wire w_dff_A_tTgmfphQ8_1;
	wire w_dff_A_pHdo0g8s9_1;
	wire w_dff_B_rgXWuGbk1_2;
	wire w_dff_B_lEOwJkwd9_2;
	wire w_dff_B_HNfOPdWG3_2;
	wire w_dff_B_b60A2s786_2;
	wire w_dff_B_2QcC4uf46_2;
	wire w_dff_B_CPgWZ9vI4_0;
	wire w_dff_B_BQKshNcL9_0;
	wire w_dff_B_L9CTJBsM8_0;
	wire w_dff_B_BT1wfhvp5_1;
	wire w_dff_B_vRekUBR52_1;
	wire w_dff_B_OJFvKyQI8_1;
	wire w_dff_B_MDjvm9xl0_1;
	wire w_dff_B_BFZeTVQt1_1;
	wire w_dff_B_wbZ2kgpr0_1;
	wire w_dff_B_3e994TVL5_1;
	wire w_dff_B_o1ld9FgW2_1;
	wire w_dff_B_QwlKy81m2_1;
	wire w_dff_B_Vnhx5BuQ2_1;
	wire w_dff_B_S7UP4dzI8_1;
	wire w_dff_B_irgtnqym3_1;
	wire w_dff_B_LL0vGEG51_1;
	wire w_dff_B_KwCLLSB36_1;
	wire w_dff_B_4lppfiRp5_1;
	wire w_dff_B_GfkogCA50_1;
	wire w_dff_B_Lun4TgfG5_1;
	wire w_dff_B_0JtIXeks0_0;
	wire w_dff_B_gbAOKVfw2_0;
	wire w_dff_B_5Bwc77lF8_0;
	wire w_dff_B_gdFh1aYu1_0;
	wire w_dff_B_PV7Z3eCq6_0;
	wire w_dff_B_BApgaGwq5_0;
	wire w_dff_B_l8XTke5Z7_0;
	wire w_dff_B_OAS7MuBZ6_0;
	wire w_dff_B_B9JBJ9031_1;
	wire w_dff_B_O7xxMIBe2_1;
	wire w_dff_B_SdDV3byI7_1;
	wire w_dff_B_iEA9xJDk0_0;
	wire w_dff_B_Cta6HihX1_0;
	wire w_dff_B_2rjMd3se2_0;
	wire w_dff_B_I7zxjpBj9_0;
	wire w_dff_B_7shGJBdY2_0;
	wire w_dff_B_5J46EBdU9_0;
	wire w_dff_B_ugAVC3ph0_0;
	wire w_dff_B_kr5Q7uVQ5_0;
	wire w_dff_B_CVGMQyU47_0;
	wire w_dff_B_X2z5vmO42_0;
	wire w_dff_B_9NmeohgU2_0;
	wire w_dff_B_290SYT7O3_0;
	wire w_dff_B_IVsL0sZo9_0;
	wire w_dff_B_l8UL9uop4_0;
	wire w_dff_B_B3GFjWaI7_0;
	wire w_dff_B_JG5CIk200_0;
	wire w_dff_B_4pwTS0wB0_0;
	wire w_dff_A_nDaZdZov6_1;
	wire w_dff_A_rcujZ2oE8_1;
	wire w_dff_A_I42mvFI97_1;
	wire w_dff_A_UQBvNC652_1;
	wire w_dff_A_JuciOKGi8_2;
	wire w_dff_A_pxZtaReL0_2;
	wire w_dff_A_477LDJ4G8_2;
	wire w_dff_A_NWEkugVQ3_2;
	wire w_dff_A_wRe8lVGu0_2;
	wire w_dff_A_dVAfYEhO8_2;
	wire w_dff_A_gUPPNxoU6_2;
	wire w_dff_A_STqZxIi20_2;
	wire w_dff_A_y0JqANA15_2;
	wire w_dff_A_mtZqKfHV3_2;
	wire w_dff_A_fzW89w8z8_2;
	wire w_dff_A_57MW5ouo1_2;
	wire w_dff_A_VfDUbObf6_2;
	wire w_dff_A_su9DqBxa6_2;
	wire w_dff_A_Y7WKfHCC6_2;
	wire w_dff_A_9egDAeHd7_2;
	wire w_dff_B_m5hw7YnI1_3;
	wire w_dff_B_1enUmcj93_3;
	wire w_dff_B_jbCKAF4M3_3;
	wire w_dff_B_qbRnz3Ku9_0;
	wire w_dff_B_rdIMQoTt5_0;
	wire w_dff_B_7vykC2Sy8_0;
	wire w_dff_B_Id4qsDKp8_0;
	wire w_dff_B_0CS3cZfD4_0;
	wire w_dff_B_EP5t6Ueb1_0;
	wire w_dff_B_cyiGqZzo3_0;
	wire w_dff_B_3ZnM1Mw94_0;
	wire w_dff_B_yfGAFMFW6_0;
	wire w_dff_B_FOWnRYgm5_0;
	wire w_dff_B_UmDUmI8U8_0;
	wire w_dff_B_8aGUcFe22_0;
	wire w_dff_A_AdRreLLg7_1;
	wire w_dff_A_T4VSx2Fc3_1;
	wire w_dff_A_Os34ysUw2_1;
	wire w_dff_A_cntpAp7F7_1;
	wire w_dff_A_umttXLsx6_1;
	wire w_dff_A_78EKFMid6_1;
	wire w_dff_A_YE6unQTE1_1;
	wire w_dff_B_mE4r2VJp7_2;
	wire w_dff_B_7JCPp54f4_2;
	wire w_dff_B_TpvOAebs8_2;
	wire w_dff_B_ae0WsQPs3_2;
	wire w_dff_B_2hCUtnVv2_2;
	wire w_dff_B_7LQryvWr4_2;
	wire w_dff_B_jU9Y2Liy2_2;
	wire w_dff_B_jyPnGC367_2;
	wire w_dff_B_8kfqkchA5_2;
	wire w_dff_B_slQaUEwN2_2;
	wire w_dff_B_as9m61SM4_2;
	wire w_dff_B_TNqvWjH05_2;
	wire w_dff_B_RNFNZPNZ6_0;
	wire w_dff_B_BYgSR66Y5_0;
	wire w_dff_B_tnGwUCCF3_0;
	wire w_dff_B_h774zQpj6_0;
	wire w_dff_B_btPUfdhX8_0;
	wire w_dff_B_5wWHOG5Z8_0;
	wire w_dff_B_Ipi3dn0D4_0;
	wire w_dff_B_gtNNXPav0_0;
	wire w_dff_B_oX7W0P6n7_0;
	wire w_dff_B_aUl8IxEi7_0;
	wire w_dff_B_ZetI8zSD9_0;
	wire w_dff_B_UGxZ7lFd5_0;
	wire w_dff_B_o3Lxyyui5_3;
	wire w_dff_B_1qJbNLwG1_3;
	wire w_dff_B_PXk43iGC9_3;
	wire w_dff_B_35fkCRxo0_3;
	wire w_dff_B_VeKVQlt00_3;
	wire w_dff_B_s2NUqyJr0_3;
	wire w_dff_B_IjYFWwaV1_3;
	wire w_dff_B_A17VGGhj5_3;
	wire w_dff_B_4mU5CPv50_3;
	wire w_dff_B_nrtOx7dN6_3;
	wire w_dff_B_bfeFApFI5_3;
	wire w_dff_B_1TtCNeJd6_3;
	wire w_dff_B_vddRwIyd2_3;
	wire w_dff_B_5jMRDQqI2_3;
	wire w_dff_B_3feuBcIM0_3;
	wire w_dff_B_dX4Zthjp2_3;
	wire w_dff_B_4DpitqpM3_3;
	wire w_dff_B_h5i4nYIP8_3;
	wire w_dff_B_EQWtMFSW0_3;
	wire w_dff_A_qm3V73ow2_0;
	wire w_dff_A_Tjs7jqik5_0;
	wire w_dff_A_F9HH5xu79_0;
	wire w_dff_A_qRwU4ddM5_0;
	wire w_dff_A_uzrdb2sV6_0;
	wire w_dff_A_XTJGXc3d5_0;
	wire w_dff_A_kvAyxm348_0;
	wire w_dff_A_IP7mBN9E7_0;
	wire w_dff_A_GzFwDnGV1_0;
	wire w_dff_A_efIUWXha9_0;
	wire w_dff_A_i0n28pc09_0;
	wire w_dff_A_Ol78IyE07_0;
	wire w_dff_A_Pic31c0g9_0;
	wire w_dff_A_hFyNf2gp7_0;
	wire w_dff_A_XVbKIfHm6_1;
	wire w_dff_A_gphEXCPu7_1;
	wire w_dff_A_YtxervhW8_1;
	wire w_dff_A_0BCslKa28_1;
	wire w_dff_A_sIlKmTIk2_1;
	wire w_dff_A_UkuR83006_1;
	wire w_dff_A_MBQafO8t9_1;
	wire w_dff_A_LaJMjqf63_1;
	wire w_dff_A_1Ze5oN6V2_1;
	wire w_dff_A_CQCZnukW9_1;
	wire w_dff_B_9zmlM31z8_1;
	wire w_dff_B_K5O94ioG0_1;
	wire w_dff_B_D0HAbg2r7_1;
	wire w_dff_B_R8fjVUsO4_1;
	wire w_dff_B_zoj3t5tp7_1;
	wire w_dff_B_PGSPpr9L6_1;
	wire w_dff_B_y0AQQQ5r5_1;
	wire w_dff_B_cAueN9243_1;
	wire w_dff_B_A0nkvEoo2_1;
	wire w_dff_B_1PVp4q1H5_1;
	wire w_dff_B_vGa7ZA0O3_1;
	wire w_dff_B_TdT9F8l34_1;
	wire w_dff_B_rdUN98LT6_1;
	wire w_dff_B_7AlBMn8z4_1;
	wire w_dff_B_Fs1JxQFF8_1;
	wire w_dff_B_jzhRgWuO1_1;
	wire w_dff_B_BPk0jcx12_1;
	wire w_dff_B_5UKvz1BV5_1;
	wire w_dff_B_SvFmXFXy0_1;
	wire w_dff_A_IBNlclkX0_0;
	wire w_dff_A_mYqwX8PM9_0;
	wire w_dff_A_YnWSadld2_0;
	wire w_dff_A_J0SmL0Lz6_0;
	wire w_dff_A_NpT0gloa1_0;
	wire w_dff_A_1gR5hOrD4_0;
	wire w_dff_A_9JdlS2n67_0;
	wire w_dff_A_jVAIWxSm1_0;
	wire w_dff_A_d8remCbq1_0;
	wire w_dff_A_u4QAVovr0_0;
	wire w_dff_A_BWxM5W4l6_0;
	wire w_dff_B_scTNcYtf5_1;
	wire w_dff_B_D7KAaGaU8_1;
	wire w_dff_B_LFBeO9jF8_1;
	wire w_dff_B_u7Ko2cDu1_1;
	wire w_dff_B_X0nIvMJv5_1;
	wire w_dff_B_0VaK6qKA7_1;
	wire w_dff_B_rTyk81Ci5_1;
	wire w_dff_B_ihuTnrWi8_1;
	wire w_dff_B_Qe26gSrG6_1;
	wire w_dff_B_YznDGJU62_0;
	wire w_dff_A_GAUrzCC51_0;
	wire w_dff_A_ybOcknkA1_0;
	wire w_dff_A_8ikj3pmB8_0;
	wire w_dff_A_OB0T8kDx4_0;
	wire w_dff_A_fDdH1Y1f5_0;
	wire w_dff_A_cgqoNBhx2_0;
	wire w_dff_A_n7CHZb1D0_0;
	wire w_dff_A_yv34kAe32_0;
	wire w_dff_A_7mL1KvRt6_0;
	wire w_dff_A_NCva8RBO6_0;
	wire w_dff_A_vSbt27XT8_0;
	wire w_dff_A_hEchCG9b8_0;
	wire w_dff_A_fZs2ZWdW2_1;
	wire w_dff_A_EX1LRekP0_1;
	wire w_dff_A_cj3BLgXr6_1;
	wire w_dff_A_SajO6ibN1_1;
	wire w_dff_A_50kmlw7L5_1;
	wire w_dff_A_m6X3qeO16_1;
	wire w_dff_A_uWFW5vFM3_1;
	wire w_dff_A_6iGsjrnf4_1;
	wire w_dff_A_kPXeZyBL2_1;
	wire w_dff_A_Fd6zMXsT1_1;
	wire w_dff_A_RCqGhqE04_1;
	wire w_dff_A_roiBgEmt3_1;
	wire w_dff_A_D8HwYQTS2_1;
	wire w_dff_A_EXJ3Ihjh4_1;
	wire w_dff_A_nc8Ki9XG2_1;
	wire w_dff_A_tYqylR2b8_1;
	wire w_dff_A_uyp60RjA7_1;
	wire w_dff_A_GalQl23S9_1;
	wire w_dff_A_alPEdqvK7_1;
	wire w_dff_B_3zMMKSHN0_2;
	wire w_dff_B_YtmsBo2T0_2;
	wire w_dff_B_VTfTOa1U4_2;
	wire w_dff_B_wjvOcLtB7_2;
	wire w_dff_B_JDTa9cxO0_2;
	wire w_dff_A_ei9GWXxs3_0;
	wire w_dff_A_wQk6P4as0_0;
	wire w_dff_A_vL3DhvzU0_0;
	wire w_dff_A_WC9bGbaM2_0;
	wire w_dff_A_JtQI1AOW4_0;
	wire w_dff_B_hhmIj0YZ6_0;
	wire w_dff_B_BsDb86gk3_0;
	wire w_dff_B_M5HAi76b4_0;
	wire w_dff_B_lAstQ9Ae1_0;
	wire w_dff_B_SpmEtieD5_0;
	wire w_dff_B_bnhpgtgG5_0;
	wire w_dff_B_yzkbhmro8_0;
	wire w_dff_B_FRhg6m2f5_0;
	wire w_dff_B_qwAs0RzU0_0;
	wire w_dff_B_AGQyKOT99_0;
	wire w_dff_B_tc57UX8A4_0;
	wire w_dff_B_feVGc99K0_0;
	wire w_dff_A_9XCsPnyq0_0;
	wire w_dff_A_8eEhKBq17_0;
	wire w_dff_A_5OMXwIDe1_0;
	wire w_dff_A_Ti09UHVE7_0;
	wire w_dff_A_Daa9saj76_0;
	wire w_dff_A_8WWlmnKE4_1;
	wire w_dff_A_rbPYaqof3_1;
	wire w_dff_A_FRanbqnu6_2;
	wire w_dff_A_fvdlIUf07_0;
	wire w_dff_A_hE0veTSZ4_0;
	wire w_dff_A_V3BLaXsn7_0;
	wire w_dff_A_rD5zJ8nL4_0;
	wire w_dff_A_V3ymn84W6_0;
	wire w_dff_A_YT94TjR65_0;
	wire w_dff_A_0fGialP43_0;
	wire w_dff_A_PB3WXhFH4_0;
	wire w_dff_A_TYaNBxp94_0;
	wire w_dff_A_nP3cP89Q1_0;
	wire w_dff_A_xda0SqpW2_0;
	wire w_dff_A_tRuD1V2k2_0;
	wire w_dff_A_6oNDj94a0_0;
	wire w_dff_A_iA5BEcc10_0;
	wire w_dff_A_jdcYEks77_0;
	wire w_dff_A_TO1bcOxd6_0;
	wire w_dff_A_xiihzCYQ5_1;
	wire w_dff_A_AyQQ2bSt9_1;
	wire w_dff_A_GNBlyuSq0_1;
	wire w_dff_A_fY9xoZWJ3_1;
	wire w_dff_A_mJBtE6ap4_1;
	wire w_dff_A_s4WJXje08_1;
	wire w_dff_A_PDB5Xoln1_1;
	wire w_dff_A_VKbcsXEq2_1;
	wire w_dff_A_06HFvkNS3_1;
	wire w_dff_A_DeDgElBp2_1;
	wire w_dff_A_jMCt2khf6_1;
	wire w_dff_A_7ZCymeVj2_1;
	wire w_dff_A_aWopnpTk0_1;
	wire w_dff_A_4nmzhXjS1_1;
	wire w_dff_A_fPeRa39J5_1;
	wire w_dff_A_KLSNYSLk1_1;
	wire w_dff_B_udsJNlPp0_0;
	wire w_dff_B_WK6fjMJF0_3;
	wire w_dff_B_GUFRaQMM5_3;
	wire w_dff_A_JGRcI2k97_0;
	wire w_dff_A_bgfH7TTV2_0;
	wire w_dff_A_OTuDoVcH2_0;
	wire w_dff_A_Iv7RmCSa2_0;
	wire w_dff_A_rHVxTPQG0_0;
	wire w_dff_A_3RqUMvrE7_0;
	wire w_dff_A_vJEghP9R5_0;
	wire w_dff_A_lTbCO6GF2_0;
	wire w_dff_A_aCjbTltz9_0;
	wire w_dff_A_LE96f8vS1_0;
	wire w_dff_A_ZODp8GNB0_0;
	wire w_dff_A_3c6MWIrS9_0;
	wire w_dff_A_ZUv04b8S4_0;
	wire w_dff_A_prV4Fc1H6_0;
	wire w_dff_A_cFtqU0P68_0;
	wire w_dff_A_yJEJunf87_0;
	wire w_dff_A_HNKgZz319_0;
	wire w_dff_A_DsUS2yNh5_0;
	wire w_dff_A_xDywGDeL8_1;
	wire w_dff_A_gdaA7rRV3_1;
	wire w_dff_A_TScRDQKd7_1;
	wire w_dff_A_T5GcRxaG5_1;
	wire w_dff_A_2sHnn7nZ5_1;
	wire w_dff_A_vrYJmitD3_1;
	wire w_dff_A_iNDNhe8h1_1;
	wire w_dff_A_CM21eqFK8_1;
	wire w_dff_A_fZ7jKNA22_1;
	wire w_dff_A_3OXEH8oE9_1;
	wire w_dff_A_tTZJIxOV3_1;
	wire w_dff_A_orLETswG8_1;
	wire w_dff_A_USr6oUuH6_1;
	wire w_dff_A_jSWqxQtg4_0;
	wire w_dff_A_h8xI2N846_0;
	wire w_dff_B_weg95XQN7_0;
	wire w_dff_B_pV88N8Af2_2;
	wire w_dff_B_Eyc3M63f7_2;
	wire w_dff_A_l5zi4vCn3_0;
	wire w_dff_A_QgTKHKAo5_0;
	wire w_dff_A_fruoJbux2_0;
	wire w_dff_A_LscgSKAo6_0;
	wire w_dff_A_iaF6eQku4_0;
	wire w_dff_A_geoSaktb6_0;
	wire w_dff_B_e0zlQvZn0_0;
	wire w_dff_B_jgMXV8T65_2;
	wire w_dff_B_wObdoSbL6_2;
	wire w_dff_A_XntA4lmx0_0;
	wire w_dff_A_KMuYR9Ki9_0;
	wire w_dff_A_MkTrKxAc3_0;
	wire w_dff_A_OEopb4TV0_0;
	wire w_dff_B_5Zv08cyB5_0;
	wire w_dff_B_nVVeEWNQ7_3;
	wire w_dff_B_85BJkmhI0_3;
	wire w_dff_A_IJW7lCWL1_1;
	wire w_dff_A_jxNuVVNz2_1;
	wire w_dff_B_Fp6gxk5S3_0;
	wire w_dff_B_jHmAqFaa1_3;
	wire w_dff_B_FnI5fl3B8_3;
	wire w_dff_A_qVeOrooV1_1;
	wire w_dff_A_qSpE3dCf7_1;
	wire w_dff_A_LscvcbqR1_1;
	wire w_dff_A_3BY8umy39_1;
	wire w_dff_A_zCK0k53w2_1;
	wire w_dff_A_IkbB7Ann4_1;
	wire w_dff_A_X1PHcyRL8_1;
	wire w_dff_A_GCDSSDzN3_1;
	wire w_dff_A_KeIE0M3X6_1;
	wire w_dff_B_YgOYIF3J7_1;
	wire w_dff_B_69j5AqhJ2_1;
	wire w_dff_B_03msNVtN4_1;
	wire w_dff_B_tDOpbQM73_1;
	wire w_dff_B_435MBe004_0;
	wire w_dff_B_ckRGBXmw0_0;
	wire w_dff_A_bNteBb4o9_0;
	wire w_dff_A_eaJWVmC34_0;
	wire w_dff_A_b6OPPDXl6_0;
	wire w_dff_A_q6D6LlFW4_0;
	wire w_dff_A_awmwhBX11_0;
	wire w_dff_A_EvfdTHg96_0;
	wire w_dff_A_tH90sqyA2_0;
	wire w_dff_A_z7d9PcIj6_0;
	wire w_dff_A_OS3DCQfI6_0;
	wire w_dff_A_PdjvSOFp3_0;
	wire w_dff_A_00GPrgor6_0;
	wire w_dff_A_luDb0KQi7_0;
	wire w_dff_A_nOz2c55t1_0;
	wire w_dff_A_Mx6Eqkxj6_0;
	wire w_dff_A_b79Vmeps7_0;
	wire w_dff_A_lhQwHW589_1;
	wire w_dff_A_DJPvStd51_1;
	wire w_dff_A_KJrEFhzp3_1;
	wire w_dff_A_ugyXVVpA3_1;
	wire w_dff_A_CkolcgPb0_1;
	wire w_dff_A_SlJU4UrV7_1;
	wire w_dff_A_uQx4ckUS8_1;
	wire w_dff_A_TzXperJG2_1;
	wire w_dff_A_zM1eOZtC8_1;
	wire w_dff_A_vugQn8406_1;
	wire w_dff_A_AUAQRt9i6_1;
	wire w_dff_A_YzinDvIG0_1;
	wire w_dff_A_GDRDDe720_1;
	wire w_dff_A_5hJs1hqs3_1;
	wire w_dff_A_5EVaKySu6_1;
	wire w_dff_B_S3vLjFV19_1;
	wire w_dff_A_uEeCJ1Kd7_0;
	wire w_dff_A_QHpEqIbG6_1;
	wire w_dff_A_ZFBqdPzH8_1;
	wire w_dff_A_YECXhcwt4_1;
	wire w_dff_A_6qsqugpf0_1;
	wire w_dff_A_yzBiQcqj7_1;
	wire w_dff_A_6zVeFx6p9_1;
	wire w_dff_A_4hJKT1sK1_1;
	wire w_dff_A_XH7GOK6u1_1;
	wire w_dff_A_TAgsMGfK2_1;
	wire w_dff_A_FNk3zqNX8_1;
	wire w_dff_A_xbUZFV986_1;
	wire w_dff_A_21BPTPe51_1;
	wire w_dff_A_ANqimZD49_1;
	wire w_dff_A_2b5r9XDY0_1;
	wire w_dff_A_vbxwZFMd3_1;
	wire w_dff_A_vkydJDqY9_0;
	wire w_dff_A_4MCI9L6I6_0;
	wire w_dff_A_j5XxWvrR8_0;
	wire w_dff_A_fbr8mnGz1_0;
	wire w_dff_A_Uec39Vxm9_0;
	wire w_dff_A_XpT8h68v5_0;
	wire w_dff_A_JT7c7LVJ0_0;
	wire w_dff_A_RtbzAyDX5_0;
	wire w_dff_A_SSwrhQ8X7_0;
	wire w_dff_A_cDmOmi2l9_0;
	wire w_dff_A_SGFZ6jdn9_0;
	wire w_dff_A_jBuDZjtb2_0;
	wire w_dff_A_MDhyBYyy5_0;
	wire w_dff_A_Ai9LT4dN0_0;
	wire w_dff_B_o1O7qU5H6_2;
	wire w_dff_B_IqbrtGa19_2;
	wire w_dff_A_pQkm35fj1_0;
	wire w_dff_A_FMkZpi7v5_0;
	wire w_dff_A_cG90Depa6_0;
	wire w_dff_A_unpagc5b3_0;
	wire w_dff_A_5Zp1Rz6K0_0;
	wire w_dff_B_KqLYUZDQ6_0;
	wire w_dff_B_e7htl35A0_0;
	wire w_dff_B_F2BKuxDP9_0;
	wire w_dff_B_6j8hxfvM7_0;
	wire w_dff_B_MsCHrmr83_0;
	wire w_dff_B_X4PMTLHp7_0;
	wire w_dff_B_DOzSByfZ5_0;
	wire w_dff_B_sMzYAUte7_0;
	wire w_dff_B_QJV3MsJg7_0;
	wire w_dff_B_65m4t7KB8_0;
	wire w_dff_B_091w0Pok9_0;
	wire w_dff_A_ybfPvBur3_0;
	wire w_dff_A_pI7MVA4b9_0;
	wire w_dff_A_8EHDGjs86_0;
	wire w_dff_A_dWI06zRd7_0;
	wire w_dff_A_8MIFdefm4_0;
	wire w_dff_A_8d4m0tp26_0;
	wire w_dff_A_zFQxOV633_0;
	wire w_dff_A_Vjj4665X5_0;
	wire w_dff_A_6IeYrVai6_0;
	wire w_dff_A_AMtld9Wl3_0;
	wire w_dff_A_vDntd9NQ4_0;
	wire w_dff_A_RgGa0dKo8_0;
	wire w_dff_A_97LXNt6R5_0;
	wire w_dff_A_Ak9pEssV8_0;
	wire w_dff_A_4kuSY1976_0;
	wire w_dff_B_IaCFlZPL7_0;
	wire w_dff_B_ecKi21p28_2;
	wire w_dff_B_KBlbIcD88_2;
	wire w_dff_A_LhxZ9yvu1_0;
	wire w_dff_A_3ecQssV03_0;
	wire w_dff_A_B9TyBP2u3_0;
	wire w_dff_A_u1mi4Nci9_0;
	wire w_dff_A_ChkCkPCG1_0;
	wire w_dff_A_a1W6TsAm6_0;
	wire w_dff_B_kkY0ITpc8_0;
	wire w_dff_B_DIXkC6457_2;
	wire w_dff_B_rDypx3QF1_2;
	wire w_dff_A_jsDu7JGM6_0;
	wire w_dff_A_EQpDDZVm1_0;
	wire w_dff_A_uCDmfV8Y8_0;
	wire w_dff_A_TzYAG5a67_0;
	wire w_dff_A_QWnGeewX5_0;
	wire w_dff_A_dL7AEjMH8_0;
	wire w_dff_A_uiXOHSwA0_0;
	wire w_dff_A_OHXkGUO91_0;
	wire w_dff_A_yxnOPSmp4_0;
	wire w_dff_A_7DKIzzbP0_0;
	wire w_dff_A_84v2MvXe0_0;
	wire w_dff_A_l3ve8aSz6_0;
	wire w_dff_A_vE46GMCE9_0;
	wire w_dff_A_Zmjj8Jnz9_0;
	wire w_dff_A_v2SSRHR16_0;
	wire w_dff_A_u5ULDn1n2_0;
	wire w_dff_A_wa18ZgDf7_0;
	wire w_dff_A_bwotvWOV0_0;
	wire w_dff_A_plzIH1ja0_0;
	wire w_dff_A_7oRzPrHY1_0;
	wire w_dff_B_tR2tjaxm1_0;
	wire w_dff_A_lbBsmh1h3_1;
	wire w_dff_A_SQQVOfIU1_1;
	wire w_dff_A_EDIaxeYi4_2;
	wire w_dff_A_339cPwC63_2;
	wire w_dff_A_xedMLPzf4_1;
	wire w_dff_A_445cJRKc6_1;
	wire w_dff_A_RmpajueA3_1;
	wire w_dff_A_utSlhqib3_1;
	wire w_dff_A_O9JauSfY0_2;
	wire w_dff_A_wsX0YNC02_2;
	wire w_dff_A_r4P6cOGv4_2;
	wire w_dff_A_EQH8NnY96_2;
	wire w_dff_A_yVK7dEXE8_2;
	wire w_dff_A_BPCBrWS85_2;
	wire w_dff_A_XSDoLaRM3_2;
	wire w_dff_A_MPcsl6oq8_2;
	wire w_dff_A_SO4bQKQp2_2;
	wire w_dff_A_Dk6p4Npt7_2;
	wire w_dff_A_7d0795xP8_2;
	wire w_dff_A_EIJwjZK89_2;
	wire w_dff_A_csZHfrIq6_2;
	wire w_dff_A_nOxzqm5H3_2;
	wire w_dff_A_Qo2yRsu17_2;
	wire w_dff_A_xLohmLmE5_2;
	wire w_dff_A_H0gCuUDW9_0;
	wire w_dff_A_CCugBIQk7_0;
	wire w_dff_B_CjTSjO7E8_0;
	wire w_dff_B_ADpLKgMs9_2;
	wire w_dff_B_dndzmJYW5_2;
	wire w_dff_A_Qol9Hgyz9_1;
	wire w_dff_A_IOQKiYa81_1;
	wire w_dff_A_yPBV31yn5_1;
	wire w_dff_A_YfhzjrCU4_1;
	wire w_dff_A_blJgktoG6_1;
	wire w_dff_B_0WeHEjwT6_1;
	wire w_dff_B_UaDBvB3V8_1;
	wire w_dff_B_y5nWNQdk5_1;
	wire w_dff_B_Ua8xhl6L1_1;
	wire w_dff_B_aiMcBI5F2_1;
	wire w_dff_B_fRSBs2f97_1;
	wire w_dff_B_C4xbRZC99_1;
	wire w_dff_B_UqPa0uPt4_1;
	wire w_dff_B_jFUutsB47_1;
	wire w_dff_B_CDa1NEFu9_1;
	wire w_dff_B_MzJuDY4q3_1;
	wire w_dff_A_huNN60yY5_0;
	wire w_dff_A_TpdLIMfW3_0;
	wire w_dff_A_UDdkHcvX9_0;
	wire w_dff_A_h5SWxiMo9_0;
	wire w_dff_A_bezJG88q0_0;
	wire w_dff_A_0llaWvgg7_0;
	wire w_dff_A_8FalD9Nv6_0;
	wire w_dff_A_N7kOG1OK9_0;
	wire w_dff_A_FfUoooxR6_0;
	wire w_dff_B_ljb0zYS01_1;
	wire w_dff_B_sKZIO4Kl7_1;
	wire w_dff_B_Xl0nzo603_1;
	wire w_dff_B_AfjZREIl4_1;
	wire w_dff_B_kJRIfhOg9_1;
	wire w_dff_B_fy9JpJqG4_1;
	wire w_dff_B_eIy8GjQg9_1;
	wire w_dff_A_J4NwGS2D7_1;
	wire w_dff_A_FDiXDb1n2_1;
	wire w_dff_A_ZXnimiPQ6_1;
	wire w_dff_A_40yMJiQN1_1;
	wire w_dff_A_mtHNvLUC4_1;
	wire w_dff_A_Kl9881X80_1;
	wire w_dff_A_qjketKGe4_1;
	wire w_dff_A_J8jpYEg64_1;
	wire w_dff_A_0hSalTxC6_1;
	wire w_dff_A_NpEFCCjl2_1;
	wire w_dff_A_HHg4Rz2y6_0;
	wire w_dff_A_xXkZjEFp7_0;
	wire w_dff_A_nf5lgtpQ7_0;
	wire w_dff_A_L8Ushhu59_0;
	wire w_dff_A_bZekAmin1_0;
	wire w_dff_A_x4bIKLof6_0;
	wire w_dff_A_dhhsFBbt7_0;
	wire w_dff_A_A9i6iMN36_0;
	wire w_dff_A_kaXZPYvP4_1;
	wire w_dff_A_GkDG18xJ9_1;
	wire w_dff_A_SNKgBfrg9_1;
	wire w_dff_A_10WBB4Jz3_1;
	wire w_dff_A_yfMtXqFG7_1;
	wire w_dff_A_zmmBnKTY3_1;
	wire w_dff_A_hdKrECdf5_1;
	wire w_dff_A_DJtqrTPq6_1;
	wire w_dff_A_OC8CCdl30_1;
	wire w_dff_A_Fh8TcCSe5_1;
	wire w_dff_A_218tGpni1_1;
	wire w_dff_A_df66RkNt7_1;
	wire w_dff_A_yf1K9M6n8_1;
	wire w_dff_A_4jb3fm2h9_0;
	wire w_dff_A_PTrey4Yo3_0;
	wire w_dff_A_GphfJqkJ9_0;
	wire w_dff_A_NdxeDYtO8_0;
	wire w_dff_A_01lbMFDm6_0;
	wire w_dff_B_JUhqLK8e8_0;
	wire w_dff_B_bnaJMKkr2_0;
	wire w_dff_B_Z93NSqwa0_0;
	wire w_dff_B_ao231VoQ1_0;
	wire w_dff_B_i76IiTVh7_0;
	wire w_dff_B_yGKU4BSb7_0;
	wire w_dff_B_8bNiacfX0_0;
	wire w_dff_B_DshOYC767_0;
	wire w_dff_A_JtqXeOdU1_0;
	wire w_dff_A_xzq3fRFG5_0;
	wire w_dff_A_UINr5WXI7_0;
	wire w_dff_A_2AiPig9S6_0;
	wire w_dff_A_9lSxNiku9_0;
	wire w_dff_A_KFPKnCKc0_0;
	wire w_dff_A_91GB3Sui2_0;
	wire w_dff_A_Ev4PBiJo0_0;
	wire w_dff_A_LLjFKsmq6_0;
	wire w_dff_A_uzIPxl4Y3_1;
	wire w_dff_B_HUTl7wB53_0;
	wire w_dff_B_EydYX5KM5_0;
	wire w_dff_B_NsXq0WyH9_2;
	wire w_dff_B_UbAXsghV7_2;
	wire w_dff_A_Us4OlCG36_0;
	wire w_dff_A_6bamHLNX1_0;
	wire w_dff_A_KYOOwmgG7_0;
	wire w_dff_A_3fPnOUAI5_0;
	wire w_dff_B_3aDczcGY4_0;
	wire w_dff_B_9kVB0bVY5_0;
	wire w_dff_B_YkQHhCKw0_2;
	wire w_dff_B_4m3qZeri9_2;
	wire w_dff_A_jGDrnAcx1_0;
	wire w_dff_A_LwacJX3S2_0;
	wire w_dff_A_KWi8CPzx4_0;
	wire w_dff_A_ivVSklLk1_0;
	wire w_dff_A_U5qfBbV10_0;
	wire w_dff_A_HocFgn0q5_0;
	wire w_dff_A_NUNImgY63_0;
	wire w_dff_A_3jTbFiWp1_0;
	wire w_dff_A_EpI35P097_0;
	wire w_dff_A_SInSAymw0_0;
	wire w_dff_A_ICPYsPUf0_0;
	wire w_dff_A_0vIhUAtM6_0;
	wire w_dff_A_958fcH956_0;
	wire w_dff_A_7pKwJ1Y80_0;
	wire w_dff_A_n07Ayx659_0;
	wire w_dff_A_9gZkPiu00_0;
	wire w_dff_A_cUNyhs7f3_1;
	wire w_dff_A_sBX2iUXP2_1;
	wire w_dff_A_5n4RnWEL6_1;
	wire w_dff_A_6gxuXLXQ4_1;
	wire w_dff_A_ZevnK9nJ6_2;
	wire w_dff_A_JrS3Fiud8_2;
	wire w_dff_A_vYQiPYYA5_2;
	wire w_dff_A_PjzYXQo94_2;
	wire w_dff_A_coFkWsRA8_2;
	wire w_dff_A_CRZCnrDa6_2;
	wire w_dff_A_UA2YDocM0_2;
	wire w_dff_A_Gpzedp2Q0_2;
	wire w_dff_A_6xvmeIWB7_2;
	wire w_dff_A_TR7IL9VK4_2;
	wire w_dff_A_n0ESUz6X3_2;
	wire w_dff_A_OjqN8yyk2_2;
	wire w_dff_B_0zBk2jvP7_0;
	wire w_dff_B_8B9DvCFK8_0;
	wire w_dff_B_PXXc8GBO5_2;
	wire w_dff_B_RLctYm3i2_2;
	wire w_dff_A_BLKIIpEP7_2;
	wire w_dff_A_PVoVcUMl6_2;
	wire w_dff_A_FCQ6gevJ6_2;
	wire w_dff_A_ZvkmHsyq6_2;
	wire w_dff_A_nTbbieea2_2;
	wire w_dff_A_gKcfYQCM3_2;
	wire w_dff_A_JZJusJjl4_2;
	wire w_dff_A_0qeCP5Pi8_2;
	wire w_dff_A_Ab2DlB5i8_2;
	wire w_dff_A_B5DfgghN8_2;
	wire w_dff_A_AL7tSTXe6_2;
	wire w_dff_A_8NK7dJPs5_2;
	wire w_dff_A_7VhT2UQB1_2;
	wire w_dff_A_Gqf84gAp9_2;
	wire w_dff_A_eyU1szws7_2;
	wire w_dff_B_qkHOgTH72_0;
	wire w_dff_B_YG35GxyW3_0;
	wire w_dff_B_PEQ9VT1z2_3;
	wire w_dff_B_PQGBc40z6_3;
	wire w_dff_A_MRFqdrPo2_0;
	wire w_dff_A_krJLXUrV1_0;
	wire w_dff_A_txuTezv14_0;
	wire w_dff_A_VNCGnUvp7_0;
	wire w_dff_A_jxIX0lJ19_2;
	wire w_dff_A_aV5KfnpY0_2;
	wire w_dff_B_fEbOTJcJ7_0;
	wire w_dff_A_MNG6Rabt6_0;
	wire w_dff_A_6wKJ42DQ3_0;
	wire w_dff_A_M2g0VMm52_0;
	wire w_dff_A_pDl1u0AP0_1;
	wire w_dff_B_r5qQAagg4_2;
	wire w_dff_B_EfYlwM1z4_2;
	wire w_dff_A_vtTJ75Jn1_0;
	wire w_dff_A_jXPJP4Ul0_0;
	wire w_dff_A_jlNxoxLR6_0;
	wire w_dff_A_jLE2n0rJ9_0;
	wire w_dff_B_xQBl0tyx8_0;
	wire w_dff_B_DGXLujUx0_0;
	wire w_dff_B_EeZCxGzL1_0;
	wire w_dff_B_LlkusSHQ2_0;
	wire w_dff_A_YNiCY31p0_0;
	wire w_dff_A_5OV1dwPW1_0;
	wire w_dff_A_FBZQshe61_0;
	wire w_dff_A_ABp5S7ct5_0;
	wire w_dff_A_QUz8ApJj9_0;
	wire w_dff_B_2x7k6Izw8_1;
	wire w_dff_B_m5qLykB48_1;
	wire w_dff_B_JtxtzyDc6_1;
	wire w_dff_B_VooOvSZ25_1;
	wire w_dff_B_OzIA1lgn4_1;
	wire w_dff_B_ol73AUFQ1_1;
	wire w_dff_B_OM3RWix06_1;
	wire w_dff_B_Zg42mpPj3_0;
	wire w_dff_B_YfdNglBp5_0;
	wire w_dff_B_780b8s1n6_0;
	wire w_dff_B_ISB3JEFm3_0;
	wire w_dff_B_PYnusFwX1_0;
	wire w_dff_B_EIEfZT132_0;
	wire w_dff_B_o0PEMrjh5_0;
	wire w_dff_A_gA2jriS08_0;
	wire w_dff_A_XeLStNUO4_0;
	wire w_dff_A_7IJbK2cu0_0;
	wire w_dff_A_cox8FrSk7_0;
	wire w_dff_A_y9PMKQPI2_0;
	wire w_dff_A_0RPCVCxN5_0;
	wire w_dff_A_fbNsijmB8_0;
	wire w_dff_A_Zh6HOU566_0;
	wire w_dff_A_X6FvcRRw4_0;
	wire w_dff_A_0Evq6HH87_0;
	wire w_dff_A_HZIoMgTR1_0;
	wire w_dff_A_KNh9Uhix2_0;
	wire w_dff_A_MoaKYuRC0_0;
	wire w_dff_A_LmPmyEAH3_0;
	wire w_dff_A_NJxuuXfY2_0;
	wire w_dff_A_tg3J5Qw19_0;
	wire w_dff_A_u3O8q0dd0_0;
	wire w_dff_A_nNYgLdSa5_0;
	wire w_dff_A_SgbzgMBx0_0;
	wire w_dff_A_xZRp3sQ61_0;
	wire w_dff_A_HBeBFwuV4_0;
	wire w_dff_A_RV9OZxoL4_0;
	wire w_dff_A_cZaE98gp3_0;
	wire w_dff_A_J3trp0RF9_0;
	wire w_dff_A_Q2OfWQ9W8_0;
	wire w_dff_A_D5xr9PFH4_0;
	wire w_dff_A_sFRKSLiG5_0;
	wire w_dff_A_bV9CZwQh1_0;
	wire w_dff_A_m509t6VE6_0;
	wire w_dff_A_Khm9731N6_0;
	wire w_dff_A_t4sFYymZ0_0;
	wire w_dff_A_AOmBRrzc7_0;
	wire w_dff_A_qa52qAz58_0;
	wire w_dff_A_dZUBlL9L3_0;
	wire w_dff_A_6x7fUC5X2_0;
	wire w_dff_A_yZyCMx2o7_0;
	wire w_dff_A_d1M3wBli3_0;
	wire w_dff_A_x9XEglM08_0;
	wire w_dff_A_9LvIBP7d9_0;
	wire w_dff_A_cHaWjaGn3_0;
	wire w_dff_A_t4HvP0Lb3_0;
	wire w_dff_A_M7PvdOKY1_0;
	wire w_dff_A_Ic3AEWiT2_0;
	wire w_dff_A_JHH89ISz2_0;
	wire w_dff_A_f3vWnTh30_0;
	wire w_dff_A_5pIYaN4v3_0;
	wire w_dff_A_NEib7nIp7_0;
	wire w_dff_A_a2yjqdUT8_0;
	wire w_dff_A_lneF3gDB1_0;
	wire w_dff_A_QA9ZD07p6_0;
	wire w_dff_A_lOhW6SaF6_0;
	wire w_dff_A_Cin2kwwM7_1;
	wire w_dff_A_cbOkA64P4_1;
	wire w_dff_A_JQ0S1JPM9_1;
	wire w_dff_A_5iLq8Cye5_1;
	wire w_dff_A_SzJHuo2M9_1;
	wire w_dff_A_coXT6OT86_1;
	wire w_dff_A_z00A8m8a4_1;
	wire w_dff_A_uzKLdXwp8_1;
	wire w_dff_A_kcUFjEsL6_1;
	wire w_dff_A_H2UhE8jp1_1;
	wire w_dff_A_XAnvY1zi3_1;
	wire w_dff_A_PY4Dn2pN8_1;
	wire w_dff_A_E8pfDTvF5_1;
	wire w_dff_A_MTjSPOR93_1;
	wire w_dff_A_i6EBz8z02_1;
	wire w_dff_A_RdIulqLn6_1;
	wire w_dff_A_ce52Zyu94_1;
	wire w_dff_A_ZDgOUspn3_1;
	wire w_dff_A_s5cqszX06_1;
	wire w_dff_B_rN5cNUVh2_0;
	wire w_dff_A_yRaGuZBV6_1;
	wire w_dff_A_jCNZtjfD1_1;
	wire w_dff_A_EAf0qjq49_1;
	wire w_dff_A_HUXqwlAR4_1;
	wire w_dff_A_eufje9bP7_1;
	wire w_dff_A_zZdGEytR0_1;
	wire w_dff_A_eenzGgUX0_1;
	wire w_dff_A_jh9KSGLR7_1;
	wire w_dff_A_p99mBJgi9_1;
	wire w_dff_A_oxfc5nJO4_1;
	wire w_dff_A_2G0y3i8v0_1;
	wire w_dff_A_vR7pSnCd3_1;
	wire w_dff_A_6P8zEAdh0_1;
	wire w_dff_A_vjXGWoYN2_1;
	wire w_dff_A_SbRehflK6_1;
	wire w_dff_A_EKRQMMUG3_1;
	wire w_dff_A_5UtrnW0b2_1;
	wire w_dff_A_tYEP0C1I7_1;
	wire w_dff_A_zrpSyQ9n2_1;
	wire w_dff_A_9gAtgxeD5_1;
	wire w_dff_A_8jy4uN992_1;
	wire w_dff_A_k4RWJ9WP6_0;
	wire w_dff_A_6US0F5m16_0;
	wire w_dff_A_3uwX3wIX5_0;
	wire w_dff_A_SMU084j52_2;
	wire w_dff_A_RMHGHZKQ8_1;
	wire w_dff_A_qtVxapno2_2;
	wire w_dff_A_nW69HDsr6_2;
	wire w_dff_B_jRtvoOkf6_1;
	wire w_dff_B_3dmKPqL63_1;
	wire w_dff_B_yvlUL8yN0_1;
	wire w_dff_B_cfCD5Gl36_1;
	wire w_dff_B_16f7dWCt9_1;
	wire w_dff_B_W7q1z4qJ7_1;
	wire w_dff_B_Ckxr55D59_1;
	wire w_dff_B_mq7toIlo6_1;
	wire w_dff_B_d4AAX7vs6_1;
	wire w_dff_B_v0fKB7sD8_1;
	wire w_dff_B_JHDTJUgh7_1;
	wire w_dff_B_mcI2YI0y3_1;
	wire w_dff_B_FhF1XEca0_1;
	wire w_dff_B_VDYO2Rpt6_1;
	wire w_dff_B_dnpg8Gl39_1;
	wire w_dff_B_9R9VV1R75_1;
	wire w_dff_B_K53FRdr76_1;
	wire w_dff_B_7aDvH7Ol3_1;
	wire w_dff_B_igRn2kT56_1;
	wire w_dff_B_kIUMZ3y72_1;
	wire w_dff_B_Tk1X9D675_1;
	wire w_dff_B_MIfDYEr94_1;
	wire w_dff_B_7XUiODAV7_1;
	wire w_dff_B_H67iYjbW1_1;
	wire w_dff_B_fCfGZnj25_1;
	wire w_dff_B_GOcO4ZDS3_1;
	wire w_dff_B_YRuKFWpL5_1;
	wire w_dff_B_O32HxyCm5_1;
	wire w_dff_B_xxEQ6N0d9_1;
	wire w_dff_B_HgkmMpkq4_1;
	wire w_dff_B_t5Q83ilq6_1;
	wire w_dff_B_N9Vq1s1r7_1;
	wire w_dff_B_VeIFWBtK7_0;
	wire w_dff_B_bBJAt9h86_0;
	wire w_dff_A_sFb5TV286_1;
	wire w_dff_A_8oBhqTHT1_1;
	wire w_dff_A_QOxPP0Lv3_1;
	wire w_dff_A_lqz8PcDP1_1;
	wire w_dff_A_lkSCW3v69_1;
	wire w_dff_A_pe8t0RV05_1;
	wire w_dff_A_g9hjSyA09_1;
	wire w_dff_A_UhRr5FxT5_1;
	wire w_dff_A_xgnpDOvd9_1;
	wire w_dff_A_zPCfDnca1_1;
	wire w_dff_A_8wgZDwou2_1;
	wire w_dff_B_LIg25Xc01_1;
	wire w_dff_B_dPh0iSfw8_1;
	wire w_dff_B_NnsfubA92_1;
	wire w_dff_B_tEfZilgs7_1;
	wire w_dff_B_oosQi0KE3_1;
	wire w_dff_B_es06gPn80_1;
	wire w_dff_B_8MEA0ppJ8_0;
	wire w_dff_A_zc8s8CG83_1;
	wire w_dff_A_KvwON2zq1_1;
	wire w_dff_A_ryXHJU2R3_1;
	wire w_dff_A_pBDT5ZAl5_1;
	wire w_dff_A_HVlgAT7E0_1;
	wire w_dff_A_45qkWINe8_1;
	wire w_dff_A_iLnKSvBK5_1;
	wire w_dff_A_ALdcHJPQ8_1;
	wire w_dff_A_SxindvZG8_1;
	wire w_dff_A_q4B4tKmh9_1;
	wire w_dff_A_ImXngjWN9_1;
	wire w_dff_A_iKGJ2GEw0_1;
	wire w_dff_B_9ajlYZdr3_2;
	wire w_dff_B_invpDyNA8_2;
	wire w_dff_B_ZIXfBbNh2_2;
	wire w_dff_B_8hjx9cwO1_2;
	wire w_dff_B_SRgwEUGB7_2;
	wire w_dff_B_0LmqApjW4_2;
	wire w_dff_B_vDp3rU3n0_2;
	wire w_dff_B_dDHCOc7C7_1;
	wire w_dff_B_8lzZujin8_0;
	wire w_dff_B_alLF9ndC9_0;
	wire w_dff_B_pubdDgxt8_1;
	wire w_dff_B_aC9HYw690_1;
	wire w_dff_B_aCGE8svr5_1;
	wire w_dff_B_KOp4eg1C7_1;
	wire w_dff_B_AhLXTjoJ4_1;
	wire w_dff_B_7nAtSZzz0_0;
	wire w_dff_A_hQattbZ39_0;
	wire w_dff_A_xTaIYJsU6_1;
	wire w_dff_A_4HxMOBzB0_1;
	wire w_dff_A_oTTWZ4n12_1;
	wire w_dff_A_fSJa1hQi3_1;
	wire w_dff_A_Dfo02qTY1_1;
	wire w_dff_A_wNrVRr4m0_1;
	wire w_dff_A_HIYgWKut1_1;
	wire w_dff_A_H569RaTp6_1;
	wire w_dff_A_iC0lMWdM1_1;
	wire w_dff_A_OQdcaMSn4_1;
	wire w_dff_B_3o2Gmpu88_0;
	wire w_dff_B_U6Y7eEEh5_0;
	wire w_dff_B_ykGpgJUh3_0;
	wire w_dff_B_H1VZyRNg0_0;
	wire w_dff_B_DOyrpJvK3_0;
	wire w_dff_B_Zg1Nctpa2_0;
	wire w_dff_B_F3j65Tk89_0;
	wire w_dff_A_Z1DwoZXy7_2;
	wire w_dff_A_w5hToErj1_2;
	wire w_dff_A_WxIS492Z8_2;
	wire w_dff_A_KQi5rTxb2_2;
	wire w_dff_A_WR1umVCz7_2;
	wire w_dff_A_1NCt1dSV6_2;
	wire w_dff_A_PRTQMjPF0_2;
	wire w_dff_A_lC5KzlNe7_2;
	wire w_dff_A_78EQe3MQ0_1;
	wire w_dff_A_qBGngdX23_1;
	wire w_dff_A_2KyFx0Bm4_2;
	wire w_dff_A_8nzIWA842_2;
	wire w_dff_A_ZeZZs0dV3_2;
	wire w_dff_A_UoqdUvOb5_2;
	wire w_dff_A_1SsLvTh40_2;
	wire w_dff_A_RreyfHQB5_2;
	wire w_dff_A_e4ZBWO9m4_2;
	wire w_dff_A_Zpd9tXee3_2;
	wire w_dff_A_SHEZpuKz4_2;
	wire w_dff_A_Dy7sPzxc4_2;
	wire w_dff_A_FmolRADu2_2;
	wire w_dff_A_tLCwrIOT5_2;
	wire w_dff_B_KP4L5NZK5_1;
	wire w_dff_B_FxcGtuwp1_1;
	wire w_dff_B_zAykQ3Zi5_1;
	wire w_dff_B_0aFNqMVK8_1;
	wire w_dff_B_YoGxxV7h9_0;
	wire w_dff_A_g1ouEMrq9_1;
	wire w_dff_B_tB8FLDBO1_2;
	wire w_dff_B_Ekj3GVEX2_2;
	wire w_dff_A_dCRZ8exy4_1;
	wire w_dff_A_EAmY7fFJ8_1;
	wire w_dff_A_uzqCdOZH0_1;
	wire w_dff_A_ix5hyEg16_1;
	wire w_dff_A_I3wjzGvY9_1;
	wire w_dff_A_HVi33uRr1_1;
	wire w_dff_A_a0i57bQe4_1;
	wire w_dff_A_QnAjQ93k8_1;
	wire w_dff_A_QX6Uod323_1;
	wire w_dff_A_L5XegHHS8_1;
	wire w_dff_A_QKQ2amWD8_1;
	wire w_dff_A_tJfaK4Ju3_1;
	wire w_dff_A_FTOhM2mj4_1;
	wire w_dff_A_pdOZCc329_1;
	wire w_dff_A_Z5Ds0Uve1_1;
	wire w_dff_A_3c8LB2TV3_1;
	wire w_dff_A_k3g2QycC6_1;
	wire w_dff_A_9782IDLv3_1;
	wire w_dff_A_vqJTOoUp7_1;
	wire w_dff_A_95FZA3Zm5_1;
	wire w_dff_B_I0QzRyjh5_1;
	wire w_dff_B_F8ISny507_0;
	wire w_dff_A_sTiYDLQz0_1;
	wire w_dff_A_kwZnzYGS7_1;
	wire w_dff_A_lRoOg2Uc0_2;
	wire w_dff_A_fe8fo5r10_2;
	wire w_dff_A_fwJ1w6eR5_1;
	wire w_dff_A_WhG7ffGB8_1;
	wire w_dff_A_sBxsNhxh5_1;
	wire w_dff_A_YC2tkVlL3_1;
	wire w_dff_A_IOiWJg5o5_2;
	wire w_dff_A_8JjfnqII7_2;
	wire w_dff_A_8dfze55T3_0;
	wire w_dff_A_vv5S50hW9_0;
	wire w_dff_B_B10ySFGf6_2;
	wire w_dff_B_97p8fcFJ9_1;
	wire w_dff_B_yFaDUAMU1_0;
	wire w_dff_A_Xd8iHAHD4_1;
	wire w_dff_A_tEZvOvdz5_1;
	wire w_dff_A_lgvxJug60_2;
	wire w_dff_A_0y5Ha0Y56_2;
	wire w_dff_A_RtiSY4fQ2_0;
	wire w_dff_A_fdX7CWqp1_0;
	wire w_dff_A_zLmGukhK8_0;
	wire w_dff_A_bqpQrA9F8_0;
	wire w_dff_A_JWLxaX346_0;
	wire w_dff_A_KmUpYuOj5_0;
	wire w_dff_A_GUN2MG2N4_0;
	wire w_dff_A_EilkRqAs1_0;
	wire w_dff_A_2eLJHofx6_0;
	wire w_dff_A_9xUOQxEp4_0;
	wire w_dff_A_eYpMDjrG1_0;
	wire w_dff_A_Kx8Fz1th4_0;
	wire w_dff_A_I8x6vdEz0_1;
	wire w_dff_B_z56kjaHO9_1;
	wire w_dff_B_Wt9cimE64_0;
	wire w_dff_A_qqZdnrpo0_1;
	wire w_dff_A_YqWCkFnU9_1;
	wire w_dff_A_2TAlZ9ka6_2;
	wire w_dff_A_w0Fgt6lT0_2;
	wire w_dff_A_ex8w77Gc8_1;
	wire w_dff_A_HGDNZH0E4_1;
	wire w_dff_A_LU3hBHnd8_1;
	wire w_dff_A_qntVsXhl5_1;
	wire w_dff_A_5SfUobBg9_1;
	wire w_dff_B_wYhbOksX3_1;
	wire w_dff_B_TqirbmY73_1;
	wire w_dff_B_tteSSYUL1_1;
	wire w_dff_B_z3PaCVmp0_1;
	wire w_dff_B_Ch26jVpJ5_1;
	wire w_dff_B_2yFhqfr89_1;
	wire w_dff_B_3ABd8Tn76_1;
	wire w_dff_B_ShIWzOkd9_1;
	wire w_dff_B_m2xCqVHy2_1;
	wire w_dff_B_gl1CDZkN4_1;
	wire w_dff_B_SZj7H64q1_1;
	wire w_dff_A_yPmzw50R3_1;
	wire w_dff_A_S2mrRg5I6_1;
	wire w_dff_A_uiWlQ2a99_1;
	wire w_dff_A_Pqka6t3i7_1;
	wire w_dff_A_W7mZd8nP7_1;
	wire w_dff_B_kkbqWu3W4_1;
	wire w_dff_B_1NJpbKnL3_1;
	wire w_dff_B_fczQLOE96_1;
	wire w_dff_A_3O4irouc6_1;
	wire w_dff_A_i8KOMWV04_1;
	wire w_dff_A_R0nhVeYO9_1;
	wire w_dff_A_EtzBKUza9_1;
	wire w_dff_A_2EV3RvmL5_1;
	wire w_dff_A_HM97nvu99_1;
	wire w_dff_A_FTpluSiU1_0;
	wire w_dff_A_flRhmxis9_0;
	wire w_dff_A_sN80vvk98_0;
	wire w_dff_A_TWgdoSAu6_0;
	wire w_dff_A_qvGD8QD72_2;
	wire w_dff_A_4kQZVwXf8_2;
	wire w_dff_A_857j7mv22_2;
	wire w_dff_A_SrxoqYpU5_2;
	wire w_dff_A_yB9qZISK9_1;
	wire w_dff_B_XhCpM7G88_2;
	wire w_dff_A_JqcRgyAl8_0;
	wire w_dff_A_ia4ZqPFa5_0;
	wire w_dff_B_Xx4hh2Hp1_2;
	wire w_dff_B_Ij49NSmw6_2;
	wire w_dff_B_3nfjAfVU4_2;
	wire w_dff_B_EaTX5xwa0_2;
	wire w_dff_B_Y348e3jW9_0;
	wire w_dff_B_WV33yBBi5_0;
	wire w_dff_B_kxkwTheF8_0;
	wire w_dff_A_6xDLqePH0_0;
	wire w_dff_A_jFlnITkq0_0;
	wire w_dff_A_yaaScwek6_0;
	wire w_dff_A_7mpuZtjD6_0;
	wire w_dff_A_YgyQP05y7_0;
	wire w_dff_A_G8MzJ7MA5_0;
	wire w_dff_A_8roTyld63_0;
	wire w_dff_A_Hp7boeQl5_0;
	wire w_dff_A_khTztlvm4_0;
	wire w_dff_A_NQl7Rqat5_0;
	wire w_dff_A_qntXB8sd5_0;
	wire w_dff_A_KIFSArAG1_0;
	wire w_dff_A_uIbQgI7W1_0;
	wire w_dff_A_l8ZtE8Sn4_0;
	wire w_dff_A_VVnNbHzg0_0;
	wire w_dff_A_keEUnmVx0_1;
	wire w_dff_A_oUm0klVa5_1;
	wire w_dff_A_rFFq4SYb4_1;
	wire w_dff_A_CYHEFmLD2_2;
	wire w_dff_A_jw7BCaO68_2;
	wire w_dff_A_IywU0Cun9_2;
	wire w_dff_A_TE6sAppO1_2;
	wire w_dff_A_4cSmD5gy5_2;
	wire w_dff_A_trKnJhZs1_2;
	wire w_dff_A_nGLOxQN57_2;
	wire w_dff_B_m5PZQapt5_1;
	wire w_dff_B_COBhojxa7_0;
	wire w_dff_A_fPlEzJqL3_0;
	wire w_dff_A_AbIZFLkS2_0;
	wire w_dff_A_x7xqnppb8_0;
	wire w_dff_A_PS3VzGrE0_0;
	wire w_dff_A_yTBxxcit6_1;
	wire w_dff_A_xgz0nFoM5_1;
	wire w_dff_A_LMRh3XSK2_2;
	wire w_dff_A_4E29kbFd3_2;
	wire w_dff_A_Z7XSjzxx0_2;
	wire w_dff_A_3wCQvhAm0_2;
	wire w_dff_A_PhRHS0Mz5_2;
	wire w_dff_A_PlYYp1HR2_2;
	wire w_dff_A_b2HDrILW8_2;
	wire w_dff_A_x5GUgam20_2;
	wire w_dff_A_eu9gHB4t5_2;
	wire w_dff_A_knNpTlxh2_2;
	wire w_dff_B_ZBbtVsur2_1;
	wire w_dff_B_LQ7pEVUH6_0;
	wire w_dff_B_yjs8ziQ73_3;
	wire w_dff_B_7v6UQacD2_3;
	wire w_dff_A_cTchlEhg0_0;
	wire w_dff_A_gfkGvZBc3_0;
	wire w_dff_A_r2bCk0VM8_0;
	wire w_dff_A_RV0X8r4x8_0;
	wire w_dff_A_TxZ6rDGb9_2;
	wire w_dff_A_6jZbSEWD6_2;
	wire w_dff_A_9cGYOAGn6_2;
	wire w_dff_B_zliV9cO33_1;
	wire w_dff_B_fMrwYs659_0;
	wire w_dff_B_ZA2YkqfJ9_2;
	wire w_dff_B_Sq1hXx1k3_2;
	wire w_dff_A_I0Mqpxop7_0;
	wire w_dff_A_FaoZZSWF2_0;
	wire w_dff_A_bn8IRPe41_0;
	wire w_dff_A_X1Xekpxs6_0;
	wire w_dff_A_odcbesw53_0;
	wire w_dff_A_0gJh73xG8_0;
	wire w_dff_A_8cDr3tWy7_0;
	wire w_dff_A_WazBq6Ez1_0;
	wire w_dff_A_rX7nEYGu3_1;
	wire w_dff_A_V7MBk9M43_1;
	wire w_dff_A_jXb34jZa4_1;
	wire w_dff_A_nJ6YFvbH5_0;
	wire w_dff_A_ViGJP46Z6_0;
	wire w_dff_A_BCgUxyrU9_0;
	wire w_dff_A_44Lhg1Uy2_0;
	wire w_dff_A_hoGJtfG63_0;
	wire w_dff_A_8rzJjEAT2_0;
	wire w_dff_A_jup20k5Y2_0;
	wire w_dff_A_noX17VGj4_0;
	wire w_dff_A_YYOCxAdK6_0;
	wire w_dff_A_TLkKiRen5_0;
	wire w_dff_B_weC9zydJ4_2;
	wire w_dff_B_3rT1SpkR9_2;
	wire w_dff_A_PYzgD2YE7_0;
	wire w_dff_A_ptpoevLv0_0;
	wire w_dff_A_sBlCRa8G5_0;
	wire w_dff_A_koUiVA1f6_0;
	wire w_dff_A_G2xvfzQQ1_0;
	wire w_dff_A_lgiSVfCS8_0;
	wire w_dff_A_sA0c8zSZ7_1;
	wire w_dff_A_QIQb9Krg9_1;
	wire w_dff_A_4UNmYwgZ2_1;
	wire w_dff_B_esNCd9Ls0_1;
	wire w_dff_B_rIPQjVRj5_0;
	wire w_dff_A_f45I65Ob2_0;
	wire w_dff_A_jtVdBGyi4_0;
	wire w_dff_A_TvmN6IC27_0;
	wire w_dff_A_Q5yWBHKi1_0;
	wire w_dff_A_pd39079P7_0;
	wire w_dff_A_a1ePKEFb4_2;
	wire w_dff_B_HiEtNCOm9_1;
	wire w_dff_B_Dw4rdbuH0_0;
	wire w_dff_B_VTW1elSc5_2;
	wire w_dff_B_jCrKePCp9_2;
	wire w_dff_A_RjZ9GCLL4_0;
	wire w_dff_A_8JVjjYZ15_0;
	wire w_dff_A_kxamI6kf1_0;
	wire w_dff_A_r5O3ypv00_0;
	wire w_dff_A_WSw6kBLS3_0;
	wire w_dff_A_8WeyrEFP5_0;
	wire w_dff_A_MJ2MGH4C0_1;
	wire w_dff_A_O0D74pKg7_1;
	wire w_dff_A_XXzyaZCe2_1;
	wire w_dff_A_WF0JWylQ5_1;
	wire w_dff_A_CSxwEZoC8_1;
	wire w_dff_A_5v8rNG9A4_1;
	wire w_dff_A_TBklSHzn0_1;
	wire w_dff_A_VW0sKbXd3_1;
	wire w_dff_A_F1DFpK1S7_1;
	wire w_dff_A_Br6k1EEH0_1;
	wire w_dff_A_GVT8uyKf9_1;
	wire w_dff_A_izyj3GnA6_1;
	wire w_dff_B_dHFxbENz8_1;
	wire w_dff_B_VzS5hBIf6_0;
	wire w_dff_B_x67f0iET4_2;
	wire w_dff_B_LJ3KrJqL9_2;
	wire w_dff_A_uK3mcUtQ1_0;
	wire w_dff_A_MJoPGurE9_0;
	wire w_dff_A_xLxDpNkr2_0;
	wire w_dff_A_A9SH6JlV4_0;
	wire w_dff_B_m00CwWkB1_1;
	wire w_dff_B_lKlqVw6l0_1;
	wire w_dff_B_op9X8sWH4_1;
	wire w_dff_B_At9nBWda5_1;
	wire w_dff_B_oDjgaoxa9_1;
	wire w_dff_B_jLjsK8R24_1;
	wire w_dff_B_J3vu9VkB6_1;
	wire w_dff_B_khkA4of51_1;
	wire w_dff_B_hZAdVbBO1_1;
	wire w_dff_B_9TVi3SFO8_1;
	wire w_dff_B_jQok6wNt8_1;
	wire w_dff_B_5vbgQBOk3_1;
	wire w_dff_B_SVwCx3Jk3_1;
	wire w_dff_B_6RsXKspr8_1;
	wire w_dff_B_dhPpRk0k0_1;
	wire w_dff_B_irw7pONr3_1;
	wire w_dff_B_s4b1bcjP6_1;
	wire w_dff_B_M2fLyGP78_1;
	wire w_dff_B_IzjJuRlZ8_0;
	wire w_dff_B_BBzXyyqI9_1;
	wire w_dff_B_lFsbFdkU4_1;
	wire w_dff_B_b9J8I6ba1_0;
	wire w_dff_B_4ZB7phqf9_0;
	wire w_dff_B_BRgOB9fC5_0;
	wire w_dff_B_2PExhUiz4_0;
	wire w_dff_B_MB2iYhoR7_0;
	wire w_dff_B_9LO6AAe94_0;
	wire w_dff_B_mcHUToWf6_0;
	wire w_dff_B_gm9gynBi1_1;
	wire w_dff_B_QFJrQ7Xm1_1;
	wire w_dff_B_o4Bl01oL7_1;
	wire w_dff_B_4cJYevke8_1;
	wire w_dff_B_wOKvsKX93_1;
	wire w_dff_B_aCsvP5CA5_1;
	wire w_dff_B_YU5oIvu96_1;
	wire w_dff_B_MW7VhB9m1_1;
	wire w_dff_B_O5UXEisZ1_1;
	wire w_dff_A_huJLn5st9_1;
	wire w_dff_A_CUMEv2pZ1_1;
	wire w_dff_A_I6t17dkg8_1;
	wire w_dff_A_PJc2GGi80_1;
	wire w_dff_B_TJ6gxjLw2_1;
	wire w_dff_A_2h9RBzpc9_0;
	wire w_dff_A_Q55QeYa29_0;
	wire w_dff_A_DL60yFMg3_0;
	wire w_dff_B_urJFtoOG4_2;
	wire w_dff_B_0YojitN27_2;
	wire w_dff_B_GYOl95Xk6_2;
	wire w_dff_B_K27cHxuK1_2;
	wire w_dff_A_iNx813JT8_1;
	wire w_dff_A_1oOPgSJ67_1;
	wire w_dff_A_xRUPsRID2_1;
	wire w_dff_B_9EZizkRl8_1;
	wire w_dff_B_HpY57gf01_1;
	wire w_dff_B_n0jEM33v8_0;
	wire w_dff_B_LG4LL9yI8_0;
	wire w_dff_A_PfUyz38B3_0;
	wire w_dff_A_qPYvkuac0_0;
	wire w_dff_A_1G1L2k840_0;
	wire w_dff_A_c9mCUYb77_1;
	wire w_dff_B_ZBD1w1uZ9_1;
	wire w_dff_B_GfJ845uw0_1;
	wire w_dff_B_db5qHDMU1_1;
	wire w_dff_B_PXdKW4HM7_1;
	wire w_dff_B_X5INP1zd1_1;
	wire w_dff_B_LU6sU5v11_1;
	wire w_dff_B_jGBSEGLF8_1;
	wire w_dff_B_GhpJh8ku0_1;
	wire w_dff_B_0Gr5VV637_1;
	wire w_dff_B_ca3YkLIG2_1;
	wire w_dff_A_fKpm5dyE3_0;
	wire w_dff_A_FMnGLo105_0;
	wire w_dff_A_fYmTU2qH0_0;
	wire w_dff_A_tDZA1xRC0_0;
	wire w_dff_B_pO9vYmEx8_1;
	wire w_dff_A_jO2s0pGZ6_1;
	wire w_dff_A_VKwZtXWT9_0;
	wire w_dff_A_vMV7Up726_0;
	wire w_dff_A_OAlXRzLj4_0;
	wire w_dff_A_AMzFpknM9_1;
	wire w_dff_A_lSW5RBm45_1;
	wire w_dff_A_PSFGRNPQ9_1;
	wire w_dff_A_0t1fKIX47_0;
	wire w_dff_A_u3HAFNlj0_0;
	wire w_dff_A_aacO2efu7_0;
	wire w_dff_A_EciIcRXr9_0;
	wire w_dff_A_QVIFmCto7_0;
	wire w_dff_B_wb1SXgaB4_0;
	wire w_dff_A_BskuEaBp5_1;
	wire w_dff_A_8DGK2zaE1_1;
	wire w_dff_A_16N29usL4_1;
	wire w_dff_A_4hPMsaKX4_2;
	wire w_dff_A_pKYTFRI76_2;
	wire w_dff_B_dxIieSIK9_0;
	wire w_dff_A_2GEKLgiy4_0;
	wire w_dff_A_ue6tcNJq6_0;
	wire w_dff_A_5mFDGhUz1_0;
	wire w_dff_A_LnyQNl3O7_1;
	wire w_dff_A_pHzc0oGT9_1;
	wire w_dff_A_4OpryYFd5_1;
	wire w_dff_B_L31IHJIT9_0;
	wire w_dff_B_loaANmcM8_0;
	wire w_dff_B_K4lgHV8e3_0;
	wire w_dff_B_c83Pyh6j7_0;
	wire w_dff_A_Jhv9FVMp7_1;
	wire w_dff_A_q80ykMn44_1;
	wire w_dff_A_eGSqPnke0_1;
	wire w_dff_A_2Y9KbueZ0_1;
	wire w_dff_A_NOCwwBkH1_1;
	wire w_dff_A_TNk2zobb9_1;
	wire w_dff_A_3ashGlaE8_1;
	wire w_dff_A_s5TRwFlx1_1;
	wire w_dff_A_hMPxqBCX0_1;
	wire w_dff_A_NBGRQgba6_1;
	wire w_dff_A_NXQDkBSO4_1;
	wire w_dff_A_1oemz8iY6_1;
	wire w_dff_B_toRcHFRg4_0;
	wire w_dff_A_rLLsVKt47_1;
	wire w_dff_A_R2SucpmA7_1;
	wire w_dff_B_K4gcKoet5_1;
	wire w_dff_A_zYrrV5Nr2_0;
	wire w_dff_A_hLSbtrog4_0;
	wire w_dff_A_BUUQM5Am5_0;
	wire w_dff_A_ge3nwBvm9_0;
	wire w_dff_A_74ChuIys9_0;
	wire w_dff_A_9zZV5BU62_0;
	wire w_dff_A_xw4mA3Og7_0;
	wire w_dff_A_Lz0Uftj19_0;
	wire w_dff_A_ynFzRE1J4_1;
	wire w_dff_A_YrfkQ3QR3_1;
	wire w_dff_A_ErMpNqaH7_1;
	wire w_dff_A_GsEEhB1g8_1;
	wire w_dff_A_yo6ADf9Q9_1;
	wire w_dff_A_MXCZR0Z74_0;
	wire w_dff_A_XCnpn9aE4_0;
	wire w_dff_A_b2VlgxhT9_0;
	wire w_dff_A_tUXNCgyV3_1;
	wire w_dff_A_eb3uJuHK3_0;
	wire w_dff_A_KfyikFRM7_0;
	wire w_dff_A_1jGxRfYS0_2;
	wire w_dff_A_U16CpbZ10_2;
	wire w_dff_A_RlLKWvkN5_2;
	wire w_dff_A_S3JU1x8F2_2;
	wire w_dff_A_YpwkgRTq9_2;
	wire w_dff_A_C5QUNZM13_2;
	wire w_dff_A_JAuJ1xwf2_2;
	wire w_dff_A_vEMXFiWM5_2;
	wire w_dff_A_RBqqfmj90_2;
	wire w_dff_A_rNHh4MfQ2_2;
	wire w_dff_B_dy0x9oPk3_3;
	wire w_dff_A_wWuBBJtQ6_2;
	wire w_dff_A_0n0NhMk98_2;
	wire w_dff_A_7Qn0UCgU2_1;
	wire w_dff_A_q3xzslil1_1;
	wire w_dff_A_tGm2WAAL5_1;
	wire w_dff_A_E8O9XLfM7_1;
	wire w_dff_A_UFOubWhK7_1;
	wire w_dff_A_pVaAoIcP4_1;
	wire w_dff_A_FzS2S2zR1_1;
	wire w_dff_A_OzwzaeGN9_1;
	wire w_dff_A_kv03YZqk2_1;
	wire w_dff_A_DwwcC0kn8_1;
	wire w_dff_A_dlbfW2eX1_2;
	wire w_dff_A_fCONKPFv9_2;
	wire w_dff_A_7BZFgUcx4_2;
	wire w_dff_B_CnzNEovY4_1;
	wire w_dff_B_hZCxe38Z9_1;
	wire w_dff_A_sPVJRPqW6_0;
	wire w_dff_A_KD5l7uKl2_0;
	wire w_dff_A_tQXoU1Lv0_0;
	wire w_dff_A_my3fTdNO3_0;
	wire w_dff_A_Nbe0h9oQ0_0;
	wire w_dff_A_86X0fj5T4_1;
	wire w_dff_A_vTR1YCna4_2;
	wire w_dff_A_574BHCIW0_2;
	wire w_dff_A_Ijknd9154_2;
	wire w_dff_A_xkbWnlis2_2;
	wire w_dff_A_tq5Yg5jr0_2;
	wire w_dff_B_PjRmLE2K8_3;
	wire w_dff_A_0qBs17pA6_0;
	wire w_dff_A_KWKXI7In8_0;
	wire w_dff_A_G2VPD0zK0_0;
	wire w_dff_A_E1lKdqdn1_0;
	wire w_dff_A_1rd0G7VB5_1;
	wire w_dff_A_OMo2FIRs2_1;
	wire w_dff_A_mENYvAB70_0;
	wire w_dff_A_2JLbCXVs9_0;
	wire w_dff_A_Ad37vWO88_0;
	wire w_dff_A_iigKqD6s2_0;
	wire w_dff_A_3rHATCLF8_0;
	wire w_dff_A_BLi0UKQr9_0;
	wire w_dff_A_76LSyMpR6_0;
	wire w_dff_A_InABorcy2_0;
	wire w_dff_A_suXKcclV2_0;
	wire w_dff_A_prRyeJR16_0;
	wire w_dff_A_SWBB6UnT6_0;
	wire w_dff_A_cuIgAHEu2_0;
	wire w_dff_A_g0dGJFmc4_2;
	wire w_dff_B_FV2WavSE5_3;
	wire w_dff_B_UoKPGbX53_3;
	wire w_dff_B_QVtI5MwH7_3;
	wire w_dff_B_saPTinh99_3;
	wire w_dff_A_Kou2KRdq7_1;
	wire w_dff_A_Af6X7UU30_1;
	wire w_dff_A_eaja6E129_1;
	wire w_dff_A_Vq2ID94O4_1;
	wire w_dff_A_KWA32Iz23_1;
	wire w_dff_A_R4UfypZu6_1;
	wire w_dff_A_fk14z9ty7_1;
	wire w_dff_A_ef5Ya6w85_1;
	wire w_dff_A_EEK5FmLK4_1;
	wire w_dff_A_Rsp5iJf80_1;
	wire w_dff_A_OnJU2gOs5_1;
	wire w_dff_A_MvC8enj97_1;
	wire w_dff_A_amY1LlFT9_1;
	wire w_dff_A_DfeiJWSB7_1;
	wire w_dff_A_RvJxSXRF2_1;
	wire w_dff_A_KdKlVakS3_1;
	wire w_dff_A_JD3Ar4P25_1;
	wire w_dff_A_exvZSVku9_1;
	wire w_dff_A_h7bxFk6z9_1;
	wire w_dff_A_7vaAMfFm2_1;
	wire w_dff_A_YZVpOyPU1_2;
	wire w_dff_A_sIBlrrHb1_2;
	wire w_dff_A_SbbCDg6y1_2;
	wire w_dff_A_9mi9xNZI5_2;
	wire w_dff_A_XvbWsxkx5_2;
	wire w_dff_A_P5m2N7wQ0_2;
	wire w_dff_A_lsfaQNUV0_1;
	wire w_dff_A_8axANUzT3_2;
	wire w_dff_A_zk68B4uQ0_2;
	wire w_dff_A_S7GzmQcL3_2;
	wire w_dff_A_hLmf92Cq2_1;
	wire w_dff_A_wfjjHBUE6_2;
	wire w_dff_A_qFKh4Mwt1_2;
	wire w_dff_A_X3DDNoHb1_0;
	wire w_dff_A_l77Ob5Vl6_0;
	wire w_dff_A_k12A8vKM6_0;
	wire w_dff_A_WvRS9wm33_1;
	wire w_dff_A_E2ls2dy89_1;
	wire w_dff_A_0cVCnH8u6_1;
	wire w_dff_A_shkWyTIS3_1;
	wire w_dff_A_zhpWkmtW3_1;
	wire w_dff_A_c5Rjr2fz6_1;
	wire w_dff_A_N5OXkWGO2_1;
	wire w_dff_A_5K07dMlU0_1;
	wire w_dff_A_ifjz7Lz00_1;
	wire w_dff_A_SZ5hkSWU0_1;
	wire w_dff_A_62c1h1sh6_1;
	wire w_dff_A_6Omdyta77_1;
	wire w_dff_A_w24k1fuu7_1;
	wire w_dff_A_x0axQ3Bo1_1;
	wire w_dff_A_C3zAqD5D5_2;
	wire w_dff_A_RXw50PGt5_2;
	wire w_dff_A_SPX8CwoT2_2;
	wire w_dff_A_WLYOpdFI1_2;
	wire w_dff_A_B7jS1dD42_2;
	wire w_dff_A_RNZYMGlC6_1;
	wire w_dff_A_tmkzqfJY2_1;
	wire w_dff_A_uojVJZWA6_1;
	wire w_dff_A_1cEzrf637_1;
	wire w_dff_A_h1ttq40p0_1;
	wire w_dff_A_y3ZBwYeY9_1;
	wire w_dff_A_NgEWRMSy3_1;
	wire w_dff_A_QQ5oLMlx3_1;
	wire w_dff_A_Qti2oXgi2_1;
	wire w_dff_A_LIIwCuBS1_1;
	wire w_dff_A_IhVKzAON9_1;
	wire w_dff_A_tITEsiEi1_2;
	wire w_dff_A_a9GAOO5S5_1;
	wire w_dff_A_gfk7h11r3_1;
	wire w_dff_A_hd2Mqzaw6_1;
	wire w_dff_A_0VNCIHMr9_1;
	wire w_dff_A_347Xpci38_1;
	wire w_dff_A_qgODzEOp3_1;
	wire w_dff_A_Tn3xV7u60_2;
	wire w_dff_A_ltJ4xc1Z3_2;
	wire w_dff_A_Zrtl5PyM0_2;
	wire w_dff_A_edWdi51Q7_2;
	wire w_dff_A_7Di1SXeX2_2;
	wire w_dff_A_7iVYC6bE9_2;
	wire w_dff_A_VoH33dSh0_2;
	wire w_dff_A_n14xedSG8_2;
	wire w_dff_A_sSClofRu0_1;
	wire w_dff_A_nlsLvHub1_1;
	wire w_dff_A_2d9BXJgZ3_1;
	wire w_dff_A_cItkywVa0_0;
	wire w_dff_A_XEIQ8Suh5_0;
	wire w_dff_A_dX3Ou6of5_0;
	wire w_dff_A_UPJetWPG9_2;
	wire w_dff_A_glUjB8zC3_2;
	wire w_dff_A_AXGb06am4_2;
	wire w_dff_B_q47WmY2E4_0;
	wire w_dff_B_wwJofFRd7_0;
	wire w_dff_B_qT63xhAG7_0;
	wire w_dff_B_5utHCWxS3_0;
	wire w_dff_B_kr9fsSUC8_0;
	wire w_dff_A_KBogXAzk3_0;
	wire w_dff_A_697IDlBx8_0;
	wire w_dff_A_bxwSwk7h3_0;
	wire w_dff_A_SQ5dMzzb5_0;
	wire w_dff_A_G0ij57U76_0;
	wire w_dff_A_MFPvexyx4_2;
	wire w_dff_A_RlEgPJkJ5_2;
	wire w_dff_A_26U4zmwJ3_2;
	wire w_dff_A_rJr8v8aj7_2;
	wire w_dff_A_qqx0P7Gd4_2;
	wire w_dff_A_yMBoJk9R6_2;
	wire w_dff_A_Zq4XkfBT7_2;
	wire w_dff_A_4UnqXQDH0_2;
	wire w_dff_A_ApPtfim87_2;
	wire w_dff_A_71krTW544_2;
	wire w_dff_A_mw6XjQHc2_2;
	wire w_dff_A_maRqugNU2_2;
	wire w_dff_A_QfBOhM2q5_2;
	wire w_dff_A_bSXExciB9_2;
	wire w_dff_B_mqNpbHV58_1;
	wire w_dff_A_yll1UEar9_1;
	wire w_dff_A_YbD6cyVf2_1;
	wire w_dff_A_njaxN7py0_0;
	wire w_dff_A_EZP3UGOg6_1;
	wire w_dff_A_NexS8Rvc1_1;
	wire w_dff_A_jTTnyWji3_1;
	wire w_dff_A_hPF8mIgd4_1;
	wire w_dff_A_CwnsNRDR3_1;
	wire w_dff_A_4bpRI8ih8_1;
	wire w_dff_A_lylUlSUn6_1;
	wire w_dff_A_gUs6QCIy7_1;
	wire w_dff_A_jlRhkfG69_1;
	wire w_dff_A_5vcpByya4_1;
	wire w_dff_A_ltp8zNyl2_1;
	wire w_dff_A_AnLtE6ts9_1;
	wire w_dff_A_jgZq5uJh2_0;
	wire w_dff_A_DtAQiGrm6_0;
	wire w_dff_A_jLgSfpG66_0;
	wire w_dff_A_ReUw0QMK2_2;
	wire w_dff_A_s7wugzvr8_2;
	wire w_dff_A_5XXE8IiG8_2;
	wire w_dff_B_MBUHsfhs2_1;
	wire w_dff_B_VUCu99sn2_1;
	wire w_dff_B_aj8GmS9T1_2;
	wire w_dff_A_3oBneEWV8_0;
	wire w_dff_A_xFyGdOtk0_2;
	wire w_dff_A_FtdZB51Q5_0;
	wire w_dff_A_bh05FPEv9_0;
	wire w_dff_A_xMIJMFxM8_0;
	wire w_dff_A_mg9fQe3p8_1;
	wire w_dff_A_AywLlYws1_1;
	wire w_dff_A_7DviQrrN0_1;
	wire w_dff_A_e4k50gv77_1;
	wire w_dff_A_6tXVjXax1_1;
	wire w_dff_A_eqJec2Nj5_1;
	wire w_dff_A_TE0SQFFm2_2;
	wire w_dff_A_sLLTmDtc5_2;
	wire w_dff_A_oO3tLiTK8_2;
	wire w_dff_A_DD47hUac5_2;
	wire w_dff_A_mQdCxS0s9_0;
	wire w_dff_A_EP7Qe2SJ0_0;
	wire w_dff_A_u9uvz5bD2_0;
	wire w_dff_A_ISnzp72h4_0;
	wire w_dff_B_TuWjnrE81_2;
	wire w_dff_A_DSMDT6GG3_0;
	wire w_dff_A_KB3kCZ4T9_0;
	wire w_dff_A_iJ9qPTqX3_0;
	wire w_dff_A_JseIA2988_0;
	wire w_dff_A_Ru4qcSYj5_1;
	wire w_dff_A_WCVjazkL5_0;
	wire w_dff_A_89rg4po88_0;
	wire w_dff_A_4esZn9dF8_0;
	wire w_dff_A_bOu4PHaO3_1;
	wire w_dff_A_CC5J1EOU6_1;
	wire w_dff_A_A0qf5rob6_1;
	wire w_dff_A_frdadZpM8_1;
	wire w_dff_A_tbWG8swD2_1;
	wire w_dff_A_TDUxJksk1_1;
	wire w_dff_A_7ComxtNr4_1;
	wire w_dff_A_WGXE9GoW3_2;
	wire w_dff_B_xKIuOT5q4_3;
	wire w_dff_B_GRmSurMV5_1;
	wire w_dff_B_Xj2Too0S0_0;
	wire w_dff_A_aOnlIr1H2_2;
	wire w_dff_A_fK8Tqv5j2_1;
	wire w_dff_A_3OVEMHkP7_2;
	wire w_dff_A_FieKRVQY5_2;
	wire w_dff_A_InQBo1k44_0;
	wire w_dff_A_BeMhbzOL0_1;
	wire w_dff_A_kgFhyGZ54_0;
	wire w_dff_A_d6LidJjF0_0;
	wire w_dff_A_MoLiEjan8_0;
	wire w_dff_A_4tZotuGY6_1;
	wire w_dff_A_1PLsBlBv4_2;
	wire w_dff_A_bNf9o2zb6_2;
	wire w_dff_A_65MHYZTc6_2;
	wire w_dff_A_HIATtF3z8_2;
	wire w_dff_B_VAc8eLdj7_1;
	wire w_dff_B_Q2fH6EwX9_1;
	wire w_dff_A_VIfWgAQG6_0;
	wire w_dff_A_Cblcpy8O5_2;
	wire w_dff_A_NdfEdzRG9_0;
	wire w_dff_A_pD8Zds0M9_0;
	wire w_dff_A_W1sTOOLS3_0;
	wire w_dff_A_Jepw3d0D3_1;
	wire w_dff_A_zEiTH9Zm9_0;
	wire w_dff_A_DaHyrcul0_0;
	wire w_dff_A_0iKJLw0g1_0;
	wire w_dff_A_AV6wUJgT5_0;
	wire w_dff_A_sRT22TuU9_0;
	wire w_dff_A_Dy8rk1pJ4_0;
	wire w_dff_A_6s52Yf0B8_0;
	wire w_dff_A_uQ130t9g2_0;
	wire w_dff_A_TAJP4QAD4_0;
	wire w_dff_A_O20LuOqV8_0;
	wire w_dff_A_bXAFYU1j4_0;
	wire w_dff_A_neZh8IbH5_0;
	wire w_dff_A_JVLOdUQK4_0;
	wire w_dff_A_hUbSJeN43_0;
	wire w_dff_A_403s3Cp35_0;
	wire w_dff_A_VUTjnMhO5_0;
	wire w_dff_A_jilfT6S19_0;
	wire w_dff_A_eWWRG6EK1_0;
	wire w_dff_A_fi0SRwT30_0;
	wire w_dff_A_qgtoXBKW1_0;
	wire w_dff_A_EhaEvVca8_0;
	wire w_dff_A_BdMyEXeo0_0;
	wire w_dff_A_wJ2uW7JW4_0;
	wire w_dff_A_OtkEzkzU6_0;
	wire w_dff_A_6grC1mMW8_0;
	wire w_dff_A_03HxQqjA3_0;
	wire w_dff_A_OVoNiMA70_1;
	wire w_dff_A_QciStLOZ8_0;
	wire w_dff_A_CwhGq5X68_0;
	wire w_dff_A_ZnbdIMLO8_0;
	wire w_dff_A_23Jebp907_0;
	wire w_dff_A_DgzauxaI8_0;
	wire w_dff_A_Ral94vLK9_0;
	wire w_dff_A_XtGDoldv8_0;
	wire w_dff_A_2iokJu8B2_0;
	wire w_dff_A_FnhgHlMu6_0;
	wire w_dff_A_j8LcjXOq1_0;
	wire w_dff_A_38YiM4ev2_0;
	wire w_dff_A_T9HddJap8_0;
	wire w_dff_A_RR49LlaI2_0;
	wire w_dff_A_eRjoXH4Y1_0;
	wire w_dff_A_t3w2MgIX5_0;
	wire w_dff_A_c5tvgWyQ8_0;
	wire w_dff_A_YaHKVIjQ4_0;
	wire w_dff_A_yT5GGK2q8_0;
	wire w_dff_A_oFfxPMDC6_0;
	wire w_dff_A_eIDU1cto8_0;
	wire w_dff_A_yerG3EhD5_0;
	wire w_dff_A_DNWumpAE1_0;
	wire w_dff_A_nn5bK9qR9_0;
	wire w_dff_A_i56gBVxo8_0;
	wire w_dff_A_0AfyUwUz9_0;
	wire w_dff_A_eg1Qo7Sp4_0;
	wire w_dff_A_At8WbDNn7_1;
	wire w_dff_A_zQnPEr3a7_0;
	wire w_dff_A_6SrnGdpF8_0;
	wire w_dff_A_mAfGAQ7J3_0;
	wire w_dff_A_zqgWuKbR3_0;
	wire w_dff_A_6sVYvNCF7_0;
	wire w_dff_A_J63G1yqV1_0;
	wire w_dff_A_RL5973yj6_0;
	wire w_dff_A_Il9fFpgK9_0;
	wire w_dff_A_EYtrwJv03_0;
	wire w_dff_A_t1NbP4ef0_0;
	wire w_dff_A_MDxGcarH7_0;
	wire w_dff_A_QorPNhsu1_0;
	wire w_dff_A_y3qeqxKp2_0;
	wire w_dff_A_hQytYnNU3_0;
	wire w_dff_A_VoGp1lo68_0;
	wire w_dff_A_qoip3ETL9_0;
	wire w_dff_A_maDAORxL5_0;
	wire w_dff_A_iDZZJ2Ol4_0;
	wire w_dff_A_gIY056G84_0;
	wire w_dff_A_G8sE0S8J5_0;
	wire w_dff_A_HFisGFMX4_0;
	wire w_dff_A_6dIB8NHN8_0;
	wire w_dff_A_vj91fIyb9_0;
	wire w_dff_A_yW2bb9pu3_0;
	wire w_dff_A_ka0RPZsU3_0;
	wire w_dff_A_j8j9jEo48_0;
	wire w_dff_A_gI7ydG0x6_1;
	wire w_dff_A_G4yDRt4f5_0;
	wire w_dff_A_k1B6fnLc5_0;
	wire w_dff_A_8WK0lKBh8_0;
	wire w_dff_A_9wZfpoQ30_0;
	wire w_dff_A_bH11QFBu1_0;
	wire w_dff_A_lPuW7BpP8_0;
	wire w_dff_A_vNVSKerB0_0;
	wire w_dff_A_QIjBGaPL9_0;
	wire w_dff_A_3gUMWUZQ5_0;
	wire w_dff_A_z4SyoYGQ5_0;
	wire w_dff_A_jcbGwhXk7_0;
	wire w_dff_A_SRkM66zP5_0;
	wire w_dff_A_P5e56rgL0_0;
	wire w_dff_A_GJyUpxno1_0;
	wire w_dff_A_w2phcBaP4_0;
	wire w_dff_A_9udBX3An0_0;
	wire w_dff_A_VaNwzoIP1_0;
	wire w_dff_A_xfKS2rmf2_0;
	wire w_dff_A_pj2PDQJZ5_0;
	wire w_dff_A_5tLmyzuw0_0;
	wire w_dff_A_S4xL5rtv1_0;
	wire w_dff_A_StaLl54y4_0;
	wire w_dff_A_5ZuSJLAl0_0;
	wire w_dff_A_HaOa1EMT9_0;
	wire w_dff_A_gJ1AdJRW5_0;
	wire w_dff_A_mWcJ8sZC0_0;
	wire w_dff_A_jVuSQxh25_1;
	wire w_dff_A_zUQEsvNU9_0;
	wire w_dff_A_zl4mvXi31_0;
	wire w_dff_A_2wNEygOh1_0;
	wire w_dff_A_0swNFLFA6_0;
	wire w_dff_A_NZAlXzUr8_0;
	wire w_dff_A_NGGMxrWH5_0;
	wire w_dff_A_tvTmI1Tq3_0;
	wire w_dff_A_Pd0J3bWB7_0;
	wire w_dff_A_evCZlh8E2_0;
	wire w_dff_A_nZMUM3jn7_0;
	wire w_dff_A_Awu2sevJ3_0;
	wire w_dff_A_bKmoNKZj4_0;
	wire w_dff_A_y7o9PyG60_0;
	wire w_dff_A_1nIWNPCK1_0;
	wire w_dff_A_nwDPreT13_0;
	wire w_dff_A_vmRHQ5fn1_0;
	wire w_dff_A_snynsPTN9_0;
	wire w_dff_A_GTCf4Bjd8_0;
	wire w_dff_A_PYfdSkSZ1_0;
	wire w_dff_A_EvvD1VHe5_0;
	wire w_dff_A_ZxTN4VId9_0;
	wire w_dff_A_NKZUlvlm9_0;
	wire w_dff_A_1N6hAOFS7_0;
	wire w_dff_A_Iv6iHDMa5_0;
	wire w_dff_A_Zk10VM4i3_0;
	wire w_dff_A_V9vjuaoO2_0;
	wire w_dff_A_ACjOL8Hd5_1;
	wire w_dff_A_OsKPVMcV6_0;
	wire w_dff_A_2gfKfQHW3_0;
	wire w_dff_A_eD6EWofz2_0;
	wire w_dff_A_4VigFBum1_0;
	wire w_dff_A_quPWRA4Z3_0;
	wire w_dff_A_JyuF0Syz4_0;
	wire w_dff_A_0AG89SoL6_0;
	wire w_dff_A_Slb9vga44_0;
	wire w_dff_A_nQA2QG915_0;
	wire w_dff_A_cAJ3BJeM4_0;
	wire w_dff_A_tSEgBoEL6_0;
	wire w_dff_A_lpBuYtKj5_0;
	wire w_dff_A_14wjCRfa1_0;
	wire w_dff_A_eq92qN2f8_0;
	wire w_dff_A_GFc4KQPw7_0;
	wire w_dff_A_FWZk4rll9_0;
	wire w_dff_A_psqGVi775_0;
	wire w_dff_A_xplWFAFY2_0;
	wire w_dff_A_5CmrKyPA8_0;
	wire w_dff_A_SNhernBQ0_0;
	wire w_dff_A_aJnWPzrI3_0;
	wire w_dff_A_PzMXKrYC4_0;
	wire w_dff_A_UVS6p7Ir9_0;
	wire w_dff_A_wisXWKJy9_0;
	wire w_dff_A_1nExP96H4_0;
	wire w_dff_A_hU3KpgwW4_0;
	wire w_dff_A_6cIJftIc7_1;
	wire w_dff_A_Lh6GAcnc6_0;
	wire w_dff_A_USVsrT7K7_0;
	wire w_dff_A_0sXoFXr06_0;
	wire w_dff_A_WN6L333g9_0;
	wire w_dff_A_VPYzLF6A0_0;
	wire w_dff_A_mmpYzzaL2_0;
	wire w_dff_A_TgDvA8u84_0;
	wire w_dff_A_vdyd8aUp2_0;
	wire w_dff_A_cruvJj447_0;
	wire w_dff_A_AYSMuxkX9_0;
	wire w_dff_A_CVYaBjgn4_0;
	wire w_dff_A_VGC4STos7_0;
	wire w_dff_A_mapEkjdk6_0;
	wire w_dff_A_jhhwobVe1_0;
	wire w_dff_A_sTbIxCxx5_0;
	wire w_dff_A_BRZyLWxa4_0;
	wire w_dff_A_kGQb8RrU4_0;
	wire w_dff_A_hYViNUUV3_0;
	wire w_dff_A_U8jzsR4N0_0;
	wire w_dff_A_NqlRo4AM4_0;
	wire w_dff_A_0PrzMRwF7_0;
	wire w_dff_A_iX2JAqtC9_0;
	wire w_dff_A_vjOGv9ky3_0;
	wire w_dff_A_K8uS5mrL0_0;
	wire w_dff_A_nMzacDpw0_0;
	wire w_dff_A_b2Azpo0M9_0;
	wire w_dff_A_oLMHIQy68_1;
	wire w_dff_A_U2TGf1IM1_0;
	wire w_dff_A_PVYwONKp7_0;
	wire w_dff_A_DFrsNgQV8_0;
	wire w_dff_A_rT2n1vbr7_0;
	wire w_dff_A_VzUZMQtS0_0;
	wire w_dff_A_2n1N2GAQ2_0;
	wire w_dff_A_WzWsWerw1_0;
	wire w_dff_A_3mObb0Dn6_0;
	wire w_dff_A_mCeZDr0O2_0;
	wire w_dff_A_9tUgrR6C3_0;
	wire w_dff_A_JYSKCyf58_0;
	wire w_dff_A_7CgXu5O03_0;
	wire w_dff_A_LFZhklvn0_0;
	wire w_dff_A_HaQ5rRU27_0;
	wire w_dff_A_9EfvHjjF8_0;
	wire w_dff_A_H6kECw7M1_0;
	wire w_dff_A_MiApOLDo8_0;
	wire w_dff_A_EccW5sm02_0;
	wire w_dff_A_QNCFt2GF6_0;
	wire w_dff_A_t0SZeUVc0_0;
	wire w_dff_A_ayYtbDTE4_0;
	wire w_dff_A_fLAGXdEm5_0;
	wire w_dff_A_W7KxjQ2U3_0;
	wire w_dff_A_6GE3KT1J6_0;
	wire w_dff_A_YuAapg5j7_0;
	wire w_dff_A_NATs0cOt0_0;
	wire w_dff_A_PH2dp2Gh6_1;
	wire w_dff_A_3uBwvu5V0_0;
	wire w_dff_A_cay00hC52_0;
	wire w_dff_A_UOFRSfUm6_0;
	wire w_dff_A_YQq5HJFC9_0;
	wire w_dff_A_UF1V6TqY3_0;
	wire w_dff_A_eQLXca4z5_0;
	wire w_dff_A_I4ooIf943_0;
	wire w_dff_A_Lpth9xgc7_0;
	wire w_dff_A_irtSG1Av6_0;
	wire w_dff_A_1FuVCvfx8_0;
	wire w_dff_A_R7OBf5QS3_0;
	wire w_dff_A_52wq3IfU8_0;
	wire w_dff_A_rA4OQhkI8_0;
	wire w_dff_A_xgNM9Hm82_0;
	wire w_dff_A_1mFIJGt20_0;
	wire w_dff_A_pV8d6myB8_0;
	wire w_dff_A_fkYSKB0U2_0;
	wire w_dff_A_DBrXzvVZ9_0;
	wire w_dff_A_ZYBwbVix6_0;
	wire w_dff_A_KFSS2HHL3_0;
	wire w_dff_A_gC9Q4zzD6_0;
	wire w_dff_A_vTmF3Vgi8_0;
	wire w_dff_A_1x3LKIsn4_0;
	wire w_dff_A_Gq4r9SHf6_0;
	wire w_dff_A_rp4WfyMj0_0;
	wire w_dff_A_Kozqd2sm0_0;
	wire w_dff_A_ck3mftU05_1;
	wire w_dff_A_5QkZzppr9_0;
	wire w_dff_A_4i9L9jy14_0;
	wire w_dff_A_FbNyRffT5_0;
	wire w_dff_A_9SyphRnW5_0;
	wire w_dff_A_rfqA71EW5_0;
	wire w_dff_A_IXqBEUwM7_0;
	wire w_dff_A_uxkjaRNX6_0;
	wire w_dff_A_IZssx8BL3_0;
	wire w_dff_A_q3JCjGgB5_0;
	wire w_dff_A_fIVMpX423_0;
	wire w_dff_A_GA1ZIZGA0_0;
	wire w_dff_A_MIwtfxl14_0;
	wire w_dff_A_OM3UJLKk1_0;
	wire w_dff_A_t2oPecny4_0;
	wire w_dff_A_g1J0EXoi1_0;
	wire w_dff_A_HRSZ4uTR0_0;
	wire w_dff_A_5RS1Sbyd9_0;
	wire w_dff_A_RH4rAyJb7_0;
	wire w_dff_A_c5Xfhjm95_0;
	wire w_dff_A_mhSKdxut6_0;
	wire w_dff_A_UtoDTZYn0_0;
	wire w_dff_A_EjPZGGWJ3_0;
	wire w_dff_A_2yHgo7sQ9_0;
	wire w_dff_A_aNaLIc3A8_0;
	wire w_dff_A_WNdDMffj4_0;
	wire w_dff_A_9Te3iLBO1_0;
	wire w_dff_A_vip4ZzAz3_1;
	wire w_dff_A_AV4YQpCp2_0;
	wire w_dff_A_h8xZlgyj0_0;
	wire w_dff_A_58AbwFuW7_0;
	wire w_dff_A_hcYwSQ2s7_0;
	wire w_dff_A_yonyJIBb3_0;
	wire w_dff_A_VCdq4rgj6_0;
	wire w_dff_A_OJNR7WCi4_0;
	wire w_dff_A_BKl1XY1o9_0;
	wire w_dff_A_gaQh5O730_0;
	wire w_dff_A_X7Q2Wy8J1_0;
	wire w_dff_A_bSupoS2p8_0;
	wire w_dff_A_5V6VCIyV1_0;
	wire w_dff_A_uWqHp8hr0_0;
	wire w_dff_A_9bOX0rlD9_0;
	wire w_dff_A_WNVCM9Z43_0;
	wire w_dff_A_0L5yOjg40_0;
	wire w_dff_A_qStqOnBr0_0;
	wire w_dff_A_Jis98WqO4_0;
	wire w_dff_A_GHrDsJGs6_0;
	wire w_dff_A_8xhs9iWv1_0;
	wire w_dff_A_lemmLzko6_0;
	wire w_dff_A_3A3nZ2Ff8_0;
	wire w_dff_A_gLgzK0w67_0;
	wire w_dff_A_cNZYIumD6_0;
	wire w_dff_A_gasweF2w8_0;
	wire w_dff_A_7WSSQWkS9_0;
	wire w_dff_A_jyfYMINM3_1;
	wire w_dff_A_eI5d90CH7_0;
	wire w_dff_A_dm5rUY5J0_0;
	wire w_dff_A_5U3jWzoV9_0;
	wire w_dff_A_xG5t2Viz6_0;
	wire w_dff_A_564LMFfM6_0;
	wire w_dff_A_93efPrR40_0;
	wire w_dff_A_3QCK2Y0q2_0;
	wire w_dff_A_9cSxeKhO9_0;
	wire w_dff_A_5MRGyAFT1_0;
	wire w_dff_A_PGLlR02d9_0;
	wire w_dff_A_FtOHGXm27_0;
	wire w_dff_A_AbNKHRsZ8_0;
	wire w_dff_A_aUwouS491_0;
	wire w_dff_A_scwVVDns8_0;
	wire w_dff_A_1MRHAMBf8_0;
	wire w_dff_A_c6VPGdOW4_0;
	wire w_dff_A_ahB1yBrd7_0;
	wire w_dff_A_PAOHaUL88_0;
	wire w_dff_A_hQpXWMcN8_0;
	wire w_dff_A_4v2CthqX5_0;
	wire w_dff_A_T08au5NZ9_0;
	wire w_dff_A_yJT368vh5_0;
	wire w_dff_A_P08PhQeu8_0;
	wire w_dff_A_uisEK8NY1_0;
	wire w_dff_A_2YzGgPL20_0;
	wire w_dff_A_8HtwiNIy5_0;
	wire w_dff_A_M7WkONvQ8_1;
	wire w_dff_A_cyPCU36U8_0;
	wire w_dff_A_suqT5l4x3_0;
	wire w_dff_A_6xfY8LbF6_0;
	wire w_dff_A_uPLLNTll7_0;
	wire w_dff_A_l8lB22ox4_0;
	wire w_dff_A_DlZXrZS05_0;
	wire w_dff_A_dJTLvTv41_0;
	wire w_dff_A_POqfTGWV1_0;
	wire w_dff_A_ZooAC3JN4_0;
	wire w_dff_A_RAT5AKzx5_0;
	wire w_dff_A_zk4foa114_0;
	wire w_dff_A_OXYE1hiF0_0;
	wire w_dff_A_7AQkkkbb8_0;
	wire w_dff_A_vgw4zCMV6_0;
	wire w_dff_A_tJ8UBXPL4_0;
	wire w_dff_A_m9pQ2itu2_0;
	wire w_dff_A_Od6sMVbx0_0;
	wire w_dff_A_USI4Smfu5_0;
	wire w_dff_A_enYjavb83_0;
	wire w_dff_A_458wZoyV6_0;
	wire w_dff_A_rrKHGKDr5_0;
	wire w_dff_A_9ONo0ROf7_0;
	wire w_dff_A_aSa4X3sQ4_0;
	wire w_dff_A_PtmdTOeI8_0;
	wire w_dff_A_JsNmkiST9_0;
	wire w_dff_A_GTd40T6T8_0;
	wire w_dff_A_e0o8y8if7_1;
	wire w_dff_A_Cd4p4fpU6_0;
	wire w_dff_A_2nhgyW6M1_0;
	wire w_dff_A_nvtOrw3v2_0;
	wire w_dff_A_qsf2dGYj5_0;
	wire w_dff_A_riVGJaof1_0;
	wire w_dff_A_OHKMqvh01_0;
	wire w_dff_A_UoJBATPS9_0;
	wire w_dff_A_qxcCGIN92_0;
	wire w_dff_A_4xrl7kY22_0;
	wire w_dff_A_Mknr19478_0;
	wire w_dff_A_svA8ebz61_0;
	wire w_dff_A_kzivBmBK6_0;
	wire w_dff_A_0K3Z0x605_0;
	wire w_dff_A_QrJLNkz36_0;
	wire w_dff_A_PPdWaEfW9_0;
	wire w_dff_A_I06EFKln0_0;
	wire w_dff_A_cHBsiLY41_0;
	wire w_dff_A_B1AYvbQT0_0;
	wire w_dff_A_wW4vcGgr0_0;
	wire w_dff_A_h2wgMVTM7_0;
	wire w_dff_A_xwEIdTjY5_0;
	wire w_dff_A_Ate1bxrH2_0;
	wire w_dff_A_xWrJP4dV4_0;
	wire w_dff_A_TfHyFaw49_0;
	wire w_dff_A_t1HdQShF2_0;
	wire w_dff_A_iSfEZZln7_0;
	wire w_dff_A_XVcUMRCc4_1;
	wire w_dff_A_2XL32K5a5_0;
	wire w_dff_A_uiqhQbLz0_0;
	wire w_dff_A_I0H3EQxG6_0;
	wire w_dff_A_skrDqLjC7_0;
	wire w_dff_A_eKPiFpX24_0;
	wire w_dff_A_XS5ZKPZQ2_0;
	wire w_dff_A_d9JQBQNR5_0;
	wire w_dff_A_Qe9mA7ZK9_0;
	wire w_dff_A_H7cQi2ZZ9_0;
	wire w_dff_A_5hcZCbP67_0;
	wire w_dff_A_YYcf8xH19_0;
	wire w_dff_A_qJML1HvV1_0;
	wire w_dff_A_itBdxZap8_0;
	wire w_dff_A_q7V6uhHE9_0;
	wire w_dff_A_flJafpRa3_0;
	wire w_dff_A_7HqnoKcr9_0;
	wire w_dff_A_am6kfWTJ2_0;
	wire w_dff_A_PT97TR9n8_0;
	wire w_dff_A_nEO17RJ86_0;
	wire w_dff_A_nMXbaVKT6_0;
	wire w_dff_A_cx7gEuE66_0;
	wire w_dff_A_0ajAiqWc5_0;
	wire w_dff_A_8A9axYqh7_0;
	wire w_dff_A_XspSFBXe7_0;
	wire w_dff_A_if33SzG11_0;
	wire w_dff_A_Zc6ARDFB9_0;
	wire w_dff_A_2X5xRMEh0_1;
	wire w_dff_A_QhKLMCDo0_0;
	wire w_dff_A_xoJHySdq8_0;
	wire w_dff_A_x2EV1CAA2_0;
	wire w_dff_A_Q2FxQJNX8_0;
	wire w_dff_A_iuf1dv8M4_0;
	wire w_dff_A_K8U8DyHM7_0;
	wire w_dff_A_itkhR4eT1_0;
	wire w_dff_A_AgbtkyvS5_0;
	wire w_dff_A_ouI8tdeK2_0;
	wire w_dff_A_oBgR1p2P5_0;
	wire w_dff_A_6AUMgknj6_0;
	wire w_dff_A_TljI974m2_0;
	wire w_dff_A_rOlg9TRa1_0;
	wire w_dff_A_H6k6SU3b9_0;
	wire w_dff_A_z6eheY2D6_0;
	wire w_dff_A_D0db2zeP7_0;
	wire w_dff_A_yAmStAph0_0;
	wire w_dff_A_JCvmZCsm9_0;
	wire w_dff_A_MoXNtrmj5_0;
	wire w_dff_A_aWvnoDxi1_0;
	wire w_dff_A_WFxlR3mX4_0;
	wire w_dff_A_KVDf182v8_0;
	wire w_dff_A_VYsIQfsL2_0;
	wire w_dff_A_tWLu8ACo1_0;
	wire w_dff_A_SAREJ7FE5_0;
	wire w_dff_A_BQV1a3BO5_0;
	wire w_dff_A_UVJM26EF8_1;
	wire w_dff_A_i6TuLoRs3_0;
	wire w_dff_A_9oRqyi9l5_0;
	wire w_dff_A_6kCn5a197_0;
	wire w_dff_A_fqm05VUl5_0;
	wire w_dff_A_E9KPb7G35_0;
	wire w_dff_A_H5iiDeJ55_0;
	wire w_dff_A_QU1YMUfJ3_0;
	wire w_dff_A_xRbZXwEe4_0;
	wire w_dff_A_hwpKUmEP9_0;
	wire w_dff_A_B8SMUqDP0_0;
	wire w_dff_A_XcnpKTvR5_0;
	wire w_dff_A_dCgBkjfG5_0;
	wire w_dff_A_H9IGAGpg8_0;
	wire w_dff_A_ku4suilp2_0;
	wire w_dff_A_VD3HGzX16_0;
	wire w_dff_A_GWFkJgQs7_0;
	wire w_dff_A_q0fx0zhG4_0;
	wire w_dff_A_N3xuPTX42_0;
	wire w_dff_A_MRqUz9zT0_0;
	wire w_dff_A_4ljUYqqs2_0;
	wire w_dff_A_VVYC8VWJ8_0;
	wire w_dff_A_4KzcN3DW1_0;
	wire w_dff_A_ztYYscuJ9_0;
	wire w_dff_A_ahxJdMfr0_0;
	wire w_dff_A_NCk9sWGy3_0;
	wire w_dff_A_uXRT81rD0_0;
	wire w_dff_A_a6FX4fFz9_1;
	wire w_dff_A_eiRbZAcj3_0;
	wire w_dff_A_2NGTuXiE8_0;
	wire w_dff_A_ECqpv6Si5_0;
	wire w_dff_A_q2IyGvVA7_0;
	wire w_dff_A_OGRgURPJ6_0;
	wire w_dff_A_3WwiB7mi3_0;
	wire w_dff_A_ghmiQXIz0_0;
	wire w_dff_A_xbKUBTv07_0;
	wire w_dff_A_4XwgKWSw7_0;
	wire w_dff_A_DfPAWoO77_0;
	wire w_dff_A_1E4wGx5g0_0;
	wire w_dff_A_aJuQUz3s2_0;
	wire w_dff_A_pX7Ngyzw3_0;
	wire w_dff_A_v6Xn2vI24_0;
	wire w_dff_A_rupQpY467_0;
	wire w_dff_A_GlKq3nDu6_0;
	wire w_dff_A_I4GJ84Kh3_0;
	wire w_dff_A_MvtqI6Uu6_0;
	wire w_dff_A_1mmkwmZc5_0;
	wire w_dff_A_7zvifdWB9_0;
	wire w_dff_A_uE0b65iD8_0;
	wire w_dff_A_PlQ2456R7_0;
	wire w_dff_A_MUdrsE2A6_0;
	wire w_dff_A_CTuzU1hT1_0;
	wire w_dff_A_4xyssGQu3_0;
	wire w_dff_A_GbszCoWy4_0;
	wire w_dff_A_HMyMtu9z5_1;
	wire w_dff_A_Oda4MulR5_0;
	wire w_dff_A_02eHjLip2_0;
	wire w_dff_A_TXoHwLFK6_0;
	wire w_dff_A_TrKKGpym4_0;
	wire w_dff_A_1l0W9sy27_0;
	wire w_dff_A_1C3jH5xg4_0;
	wire w_dff_A_k4JahgB24_0;
	wire w_dff_A_npH477mu3_0;
	wire w_dff_A_QVhByDoc8_0;
	wire w_dff_A_WX0wXZdp9_0;
	wire w_dff_A_KR2LJcZ93_0;
	wire w_dff_A_ALkl92LC8_0;
	wire w_dff_A_a4x8kVNw2_0;
	wire w_dff_A_sSIPKGpG6_0;
	wire w_dff_A_rEny0QEk6_0;
	wire w_dff_A_AYL74And5_0;
	wire w_dff_A_IumQ7v2L5_0;
	wire w_dff_A_1vJbo5Dd8_0;
	wire w_dff_A_VnItcIAc9_0;
	wire w_dff_A_kUvtkle29_0;
	wire w_dff_A_iHYF3vKC0_0;
	wire w_dff_A_kHX26XH09_0;
	wire w_dff_A_XomNeiLg2_0;
	wire w_dff_A_kf7QsZNn2_0;
	wire w_dff_A_SSEskHef4_0;
	wire w_dff_A_9ScruEEl7_0;
	wire w_dff_A_OHRyQi3h5_1;
	wire w_dff_A_W2WcKkq43_0;
	wire w_dff_A_8YUjki5V6_0;
	wire w_dff_A_umkkhyZQ7_0;
	wire w_dff_A_anJuRmiT8_0;
	wire w_dff_A_IXEjX2Zj5_0;
	wire w_dff_A_TjqDjezA9_0;
	wire w_dff_A_QpdUBKOj0_0;
	wire w_dff_A_AkhbvrF87_0;
	wire w_dff_A_rD44rxAP8_0;
	wire w_dff_A_JJfsPPqT3_0;
	wire w_dff_A_YkeD6l6y2_0;
	wire w_dff_A_orUc6Xb24_0;
	wire w_dff_A_qkWj9AlW2_0;
	wire w_dff_A_zNYmYpgW6_0;
	wire w_dff_A_bCUkCvry3_0;
	wire w_dff_A_ZBcUn4h43_0;
	wire w_dff_A_Yk9Xn3tS8_0;
	wire w_dff_A_loWhWcEG5_0;
	wire w_dff_A_geT7kneF7_0;
	wire w_dff_A_Jr7JidRa7_0;
	wire w_dff_A_iaADX08z7_0;
	wire w_dff_A_6lNPjQJD2_0;
	wire w_dff_A_eDdb3zBx5_0;
	wire w_dff_A_ETV3iEVH1_0;
	wire w_dff_A_j9RR9sOp0_0;
	wire w_dff_A_dSihZrmM2_0;
	wire w_dff_A_dqNBR2IS5_1;
	wire w_dff_A_S1DAVp1q5_0;
	wire w_dff_A_zhsLltyh1_0;
	wire w_dff_A_RT9v651b1_0;
	wire w_dff_A_A13NeRXC2_0;
	wire w_dff_A_vIQoAH6w6_0;
	wire w_dff_A_uWRfxGeZ3_0;
	wire w_dff_A_Y0LhGxmk0_0;
	wire w_dff_A_xrYYrI2L2_0;
	wire w_dff_A_1UiSVUEH1_0;
	wire w_dff_A_SkN7ktfM0_0;
	wire w_dff_A_1XAxCiMS3_0;
	wire w_dff_A_CZgN9Gqr8_0;
	wire w_dff_A_7t0dQJ0K0_0;
	wire w_dff_A_UgVaJFKq7_0;
	wire w_dff_A_oj0xsLmL4_0;
	wire w_dff_A_qYB2syE41_0;
	wire w_dff_A_uBg0JGeT4_0;
	wire w_dff_A_Vi7D5nUp8_0;
	wire w_dff_A_Xq68wXmm9_0;
	wire w_dff_A_4H6abfMT1_0;
	wire w_dff_A_WEHCrI3G6_0;
	wire w_dff_A_nQTkL1FI6_0;
	wire w_dff_A_V03hrBgb5_0;
	wire w_dff_A_C94sgvYw2_0;
	wire w_dff_A_8zOvM1ON5_0;
	wire w_dff_A_Ovb05qxY2_0;
	wire w_dff_A_0ww2XJtm7_1;
	wire w_dff_A_n42dURt56_0;
	wire w_dff_A_wZgojSWX6_0;
	wire w_dff_A_XmT3ztM21_0;
	wire w_dff_A_PpBJ0wIq6_0;
	wire w_dff_A_VaOJbH567_0;
	wire w_dff_A_FWh45Sc56_0;
	wire w_dff_A_PD5Hi5G89_0;
	wire w_dff_A_jY9AWEXO9_0;
	wire w_dff_A_bUCTdUdC6_0;
	wire w_dff_A_K6j75fEW5_0;
	wire w_dff_A_0hiITqoz4_0;
	wire w_dff_A_8l5G66fv5_0;
	wire w_dff_A_MJScctTp4_0;
	wire w_dff_A_NZNle9D65_0;
	wire w_dff_A_RJU9zxHS7_0;
	wire w_dff_A_IqURtX018_0;
	wire w_dff_A_OGBoosG52_0;
	wire w_dff_A_Y3SAtFLq1_0;
	wire w_dff_A_MxI6ffKQ9_0;
	wire w_dff_A_a6yuZfwa0_0;
	wire w_dff_A_VxiBZGlw9_0;
	wire w_dff_A_M1DoU9cO0_0;
	wire w_dff_A_cc22uoNB1_0;
	wire w_dff_A_E0jpqo7z0_0;
	wire w_dff_A_pyrRYMqX5_0;
	wire w_dff_A_NC3FtzoI3_0;
	wire w_dff_A_wEixxhLY1_1;
	wire w_dff_A_iL3knU1R5_0;
	wire w_dff_A_Zw0v5R6c1_0;
	wire w_dff_A_S4i9spnq0_0;
	wire w_dff_A_T2GnmU1C6_0;
	wire w_dff_A_3h8ks7S83_0;
	wire w_dff_A_5T0ksZaP8_0;
	wire w_dff_A_940vZeEa0_0;
	wire w_dff_A_icrPN5md5_0;
	wire w_dff_A_owhbLnWn4_0;
	wire w_dff_A_EYBjuh1g9_0;
	wire w_dff_A_863N7VV51_0;
	wire w_dff_A_k8i8ZwRV2_0;
	wire w_dff_A_OUszzLtT2_0;
	wire w_dff_A_ipEg6L4a3_0;
	wire w_dff_A_Z82bfm5B6_0;
	wire w_dff_A_fmOlB9oe5_0;
	wire w_dff_A_PD7BoTEb9_0;
	wire w_dff_A_o6lqqRf64_0;
	wire w_dff_A_1aDcas5O5_0;
	wire w_dff_A_Bp9lLQnl1_0;
	wire w_dff_A_Lk1djuk33_0;
	wire w_dff_A_tIKM2B2x1_0;
	wire w_dff_A_uUAeA6aC8_0;
	wire w_dff_A_3BVRq0st5_0;
	wire w_dff_A_qx9WmvKS0_0;
	wire w_dff_A_e60Q0Gj75_0;
	wire w_dff_A_puMfuoYc7_1;
	wire w_dff_A_pmnPc5h48_0;
	wire w_dff_A_aBHWQcLr9_0;
	wire w_dff_A_C68e9Zjy5_0;
	wire w_dff_A_GTCLMMJE9_0;
	wire w_dff_A_I2vpgGa29_0;
	wire w_dff_A_tQdzbWnE9_0;
	wire w_dff_A_Llpzg4Xh7_0;
	wire w_dff_A_qZo5rroK9_0;
	wire w_dff_A_yFkLVq7c6_0;
	wire w_dff_A_ksjhtiKw1_0;
	wire w_dff_A_XJhfglIC7_0;
	wire w_dff_A_h9e6mIHC0_0;
	wire w_dff_A_x9Hqfv1A4_0;
	wire w_dff_A_hqgkOqdv3_0;
	wire w_dff_A_hnluwi503_0;
	wire w_dff_A_CjG9sA1S8_0;
	wire w_dff_A_r20o283g3_0;
	wire w_dff_A_O1KXQbKG0_0;
	wire w_dff_A_aeYwBjJS7_0;
	wire w_dff_A_Krojhl2E2_0;
	wire w_dff_A_wladRYMI2_0;
	wire w_dff_A_CdFHsTjf5_0;
	wire w_dff_A_gOVZkuNo0_0;
	wire w_dff_A_HT8prmZC8_0;
	wire w_dff_A_IDn74baS5_0;
	wire w_dff_A_UxV47m7T2_0;
	wire w_dff_A_Zq66Xln94_1;
	wire w_dff_A_k912QvlV9_0;
	wire w_dff_A_JDVWLYkO3_0;
	wire w_dff_A_UZy8oTVM4_0;
	wire w_dff_A_kFtPJFQr4_0;
	wire w_dff_A_zIMye9rk6_0;
	wire w_dff_A_mToo5dkM1_0;
	wire w_dff_A_l2BcZYmm0_0;
	wire w_dff_A_MSwxwvR52_0;
	wire w_dff_A_6l7HzzmG6_0;
	wire w_dff_A_QN0khxl39_0;
	wire w_dff_A_29wWV7m68_0;
	wire w_dff_A_MCAWVTKd1_0;
	wire w_dff_A_pDnqd1NK9_0;
	wire w_dff_A_uZDFHRXA0_0;
	wire w_dff_A_Hf6hh8u79_0;
	wire w_dff_A_e16w1sRj6_0;
	wire w_dff_A_mz0zHQ308_0;
	wire w_dff_A_mTtOyiuh8_0;
	wire w_dff_A_L4xd6kf04_0;
	wire w_dff_A_tMj5Ac5K4_0;
	wire w_dff_A_yDuHrXsz0_0;
	wire w_dff_A_D3ngKS0I9_0;
	wire w_dff_A_n3n1o1sq7_0;
	wire w_dff_A_2GW4XwH87_0;
	wire w_dff_A_aAstr5y95_0;
	wire w_dff_A_KXsfjgmM0_0;
	wire w_dff_A_DDaoXkJA6_1;
	wire w_dff_A_7uPgKn8s1_0;
	wire w_dff_A_R9PqNNcb8_0;
	wire w_dff_A_4wer1PBI5_0;
	wire w_dff_A_H9h25ZeW8_0;
	wire w_dff_A_7Yg1dQTv9_0;
	wire w_dff_A_BX4u5fLA2_0;
	wire w_dff_A_nvPrDDjS7_0;
	wire w_dff_A_RS0yCt0l4_0;
	wire w_dff_A_UozTiDTO2_0;
	wire w_dff_A_JfCAGHWD6_0;
	wire w_dff_A_mJYsnTG26_0;
	wire w_dff_A_TBI6YeTV5_0;
	wire w_dff_A_AcpUpPxQ2_0;
	wire w_dff_A_q3l5svan7_0;
	wire w_dff_A_IECtLNfC7_0;
	wire w_dff_A_m2XGcXWk1_0;
	wire w_dff_A_93thysza7_0;
	wire w_dff_A_Y0xtZ38t1_0;
	wire w_dff_A_8hYapcuP6_0;
	wire w_dff_A_24F6oHqj8_0;
	wire w_dff_A_5uo41Vol4_0;
	wire w_dff_A_JBEVRVV80_0;
	wire w_dff_A_ddrsVdYQ1_0;
	wire w_dff_A_7GF6ZAcv3_0;
	wire w_dff_A_5AwN8fNi3_0;
	wire w_dff_A_rB18fipo2_0;
	wire w_dff_A_YECV73dN5_1;
	wire w_dff_A_p6HRyqvL5_0;
	wire w_dff_A_HHLGkS7H2_0;
	wire w_dff_A_DWFMMH563_0;
	wire w_dff_A_6LUERjae3_0;
	wire w_dff_A_rdv0ugAc8_0;
	wire w_dff_A_PyidGCmK2_0;
	wire w_dff_A_cBJpMe1Z6_0;
	wire w_dff_A_Z4x7Vb2R6_0;
	wire w_dff_A_JUWoiqKm1_0;
	wire w_dff_A_7S72pRih8_0;
	wire w_dff_A_ONwUSsQr5_0;
	wire w_dff_A_60NfhBHI5_0;
	wire w_dff_A_uqwKGK1x7_0;
	wire w_dff_A_AZFr2EUz2_0;
	wire w_dff_A_kBtBVXNo6_0;
	wire w_dff_A_5tIJVuTk2_0;
	wire w_dff_A_LmQwbT5r8_0;
	wire w_dff_A_aBRXscI79_0;
	wire w_dff_A_DSjUA1kS3_0;
	wire w_dff_A_i1qy4bcu6_0;
	wire w_dff_A_XOFoBH051_0;
	wire w_dff_A_ZkXE4HVC4_0;
	wire w_dff_A_OiBHMBkw4_0;
	wire w_dff_A_vrl2u6ps1_0;
	wire w_dff_A_DJePysRw1_0;
	wire w_dff_A_PwWKa3ae2_0;
	wire w_dff_A_9XjXRFMW1_1;
	wire w_dff_A_AoUmo7h10_0;
	wire w_dff_A_FrxE5A4p6_0;
	wire w_dff_A_UdHgtBIZ3_0;
	wire w_dff_A_lHZHKMWD3_0;
	wire w_dff_A_KlvwRLCr0_0;
	wire w_dff_A_qoNARPjP1_0;
	wire w_dff_A_y4jI1la98_0;
	wire w_dff_A_f2EUylyZ9_0;
	wire w_dff_A_qhh83PyN0_0;
	wire w_dff_A_N3RzjaRJ4_0;
	wire w_dff_A_IgKW3cWW5_0;
	wire w_dff_A_lDlx0eDO9_0;
	wire w_dff_A_H6cN5fG00_0;
	wire w_dff_A_cm5z690o8_0;
	wire w_dff_A_codDEp5I4_0;
	wire w_dff_A_IAWee61O5_0;
	wire w_dff_A_OxwJpBWY7_0;
	wire w_dff_A_m6Dj9tEO0_0;
	wire w_dff_A_Xn8SI23c7_0;
	wire w_dff_A_MrwHxCFr2_0;
	wire w_dff_A_RIcbXtz61_0;
	wire w_dff_A_HCwZUYPN8_0;
	wire w_dff_A_WY14eKx50_0;
	wire w_dff_A_jKwzFe9f8_0;
	wire w_dff_A_PvlRxVMa5_0;
	wire w_dff_A_mWbi3MvK5_0;
	wire w_dff_A_oNY1Iu5k2_1;
	wire w_dff_A_3ygRFRxZ4_0;
	wire w_dff_A_J3t9Owan0_0;
	wire w_dff_A_ggriSJyQ2_0;
	wire w_dff_A_HKErTrDQ9_0;
	wire w_dff_A_nJfkujWH1_0;
	wire w_dff_A_tqaqhby31_0;
	wire w_dff_A_1xfJCtFC3_0;
	wire w_dff_A_Q3A6fB6d8_0;
	wire w_dff_A_ukLxuOnf8_0;
	wire w_dff_A_vAbD0RGV7_0;
	wire w_dff_A_6hCQc7Mr5_0;
	wire w_dff_A_J4KLCAFv7_0;
	wire w_dff_A_J8C7zaQw3_0;
	wire w_dff_A_htoNZU9T9_0;
	wire w_dff_A_Fl3z1Gvv5_0;
	wire w_dff_A_4BknDiRD4_0;
	wire w_dff_A_ct70PNLr9_0;
	wire w_dff_A_leMRrTmm6_0;
	wire w_dff_A_flGKh7kk5_0;
	wire w_dff_A_l4gcUjJS5_0;
	wire w_dff_A_rZVWJr572_0;
	wire w_dff_A_srPGCgnv0_0;
	wire w_dff_A_eMhCmY6B5_0;
	wire w_dff_A_5AnLIGkc5_0;
	wire w_dff_A_itE0S7pK2_0;
	wire w_dff_A_pBF4rZ0k0_0;
	wire w_dff_A_A7hwHenU7_1;
	wire w_dff_A_mY29OrUp4_0;
	wire w_dff_A_31r5hcBQ9_0;
	wire w_dff_A_wJIocf6w0_0;
	wire w_dff_A_MAmOy4hl2_0;
	wire w_dff_A_63qWM3Pk8_0;
	wire w_dff_A_7oNoLsoJ9_0;
	wire w_dff_A_4VE4d1ar9_0;
	wire w_dff_A_NupIPhb90_0;
	wire w_dff_A_lpVs4XQl0_0;
	wire w_dff_A_1DjMUDJ22_0;
	wire w_dff_A_K0FtxPjW5_0;
	wire w_dff_A_DB5N1ORG7_0;
	wire w_dff_A_FMxxLnl60_0;
	wire w_dff_A_bGETVDBm9_0;
	wire w_dff_A_vrQUpQ849_0;
	wire w_dff_A_nvjl7GsZ5_0;
	wire w_dff_A_2Rb93uy34_0;
	wire w_dff_A_2Bt7Ot1C7_0;
	wire w_dff_A_svUEaiP50_0;
	wire w_dff_A_dNhxAr2S8_0;
	wire w_dff_A_d1bcCcJi4_0;
	wire w_dff_A_1CZvWQSm7_0;
	wire w_dff_A_S0g7mT5z8_0;
	wire w_dff_A_PimE1lvm5_0;
	wire w_dff_A_T7SYX85T2_0;
	wire w_dff_A_M11ZEwKf4_0;
	wire w_dff_A_5NPOVR0c6_1;
	wire w_dff_A_kedJpPF42_0;
	wire w_dff_A_hXvorjZe9_0;
	wire w_dff_A_5SdqaOmZ9_0;
	wire w_dff_A_yqYBKEO11_0;
	wire w_dff_A_ErwYmcM25_0;
	wire w_dff_A_9dg5GZsc4_0;
	wire w_dff_A_nqLbCdKB5_0;
	wire w_dff_A_gAHekINO4_0;
	wire w_dff_A_AJAY8mQs6_0;
	wire w_dff_A_HTskUTgm7_0;
	wire w_dff_A_9EhZHAuz8_0;
	wire w_dff_A_AAZVSc7z6_0;
	wire w_dff_A_qgevseyZ0_0;
	wire w_dff_A_SnCrtqNN6_0;
	wire w_dff_A_K5nXN7co7_0;
	wire w_dff_A_NsCGsO2B0_0;
	wire w_dff_A_nMPmUtWn1_0;
	wire w_dff_A_60JdOhcx9_0;
	wire w_dff_A_EP2NLLMm1_0;
	wire w_dff_A_P8wM2yDM1_0;
	wire w_dff_A_xrwBTyES9_0;
	wire w_dff_A_m2AgbVBL1_0;
	wire w_dff_A_22kH0UT49_0;
	wire w_dff_A_9c6o8sG65_0;
	wire w_dff_A_IDtfuMVe4_0;
	wire w_dff_A_CldaB4NW2_0;
	wire w_dff_A_lE27KfQ80_1;
	wire w_dff_A_IbcGrrkx1_0;
	wire w_dff_A_0Silw3NH3_0;
	wire w_dff_A_8p6ceSdA9_0;
	wire w_dff_A_Z1fCUz068_0;
	wire w_dff_A_8p41aVx76_0;
	wire w_dff_A_Bnvis7W37_0;
	wire w_dff_A_kx2HdYFi5_0;
	wire w_dff_A_OxGy5Pi77_0;
	wire w_dff_A_2c0q00AJ9_0;
	wire w_dff_A_wXjsufIw8_0;
	wire w_dff_A_6yFE6mpt9_0;
	wire w_dff_A_Nm4AP3zM7_0;
	wire w_dff_A_ISCZtJ2D2_0;
	wire w_dff_A_2lZVGOtZ8_0;
	wire w_dff_A_vqQU3vVM5_0;
	wire w_dff_A_M7XmWZI61_0;
	wire w_dff_A_BSGBPpLy8_0;
	wire w_dff_A_pGYpMhT88_0;
	wire w_dff_A_hwYNBimw2_0;
	wire w_dff_A_AYZKThBq8_0;
	wire w_dff_A_E8yAJYQA3_0;
	wire w_dff_A_GXcE2zvF3_0;
	wire w_dff_A_fLdT3Ohf0_0;
	wire w_dff_A_STI1Ss9b1_0;
	wire w_dff_A_xShdlbbk2_0;
	wire w_dff_A_IDaEoSGw1_0;
	wire w_dff_A_f8Cco9ft3_1;
	wire w_dff_A_9BNqIGXe7_0;
	wire w_dff_A_BOXFVgi66_0;
	wire w_dff_A_VlNZvv7n2_0;
	wire w_dff_A_lbjgfEZc1_0;
	wire w_dff_A_dAiTvqkL4_0;
	wire w_dff_A_MIXq8aL45_0;
	wire w_dff_A_LxR7kWq03_0;
	wire w_dff_A_Lzzkozoo4_0;
	wire w_dff_A_NAuNH7fS2_0;
	wire w_dff_A_OUDpUV965_0;
	wire w_dff_A_TZAoCCV31_0;
	wire w_dff_A_O2FWET2g9_0;
	wire w_dff_A_PGVRFjAI4_0;
	wire w_dff_A_B9TB6Ra76_0;
	wire w_dff_A_g59qcJCk6_0;
	wire w_dff_A_dYkdEKo59_0;
	wire w_dff_A_DjZfWBE83_0;
	wire w_dff_A_urMTT55F8_0;
	wire w_dff_A_pcLWPbgW1_0;
	wire w_dff_A_Z3IeNUj21_0;
	wire w_dff_A_YlWRmJC72_0;
	wire w_dff_A_lM445oJ85_0;
	wire w_dff_A_XCXeeEA88_0;
	wire w_dff_A_NWhdtGAi3_0;
	wire w_dff_A_783XIXnD7_0;
	wire w_dff_A_5OphFUEH4_0;
	wire w_dff_A_k7IiztBr1_1;
	wire w_dff_A_75iqSxfi4_0;
	wire w_dff_A_C3t7ycBr1_0;
	wire w_dff_A_2KDC6p2n0_0;
	wire w_dff_A_vOW9esJO1_0;
	wire w_dff_A_zbKfCUOS9_0;
	wire w_dff_A_t9SxDMGz4_0;
	wire w_dff_A_bn23TTcZ1_0;
	wire w_dff_A_CBRDBPW60_0;
	wire w_dff_A_opfWlgAV3_0;
	wire w_dff_A_osNiFCJ52_0;
	wire w_dff_A_iay9kg3H6_0;
	wire w_dff_A_8gc3hqAk5_0;
	wire w_dff_A_CMotSE9g8_0;
	wire w_dff_A_ZXnRSZ9T4_0;
	wire w_dff_A_rCuwRK9n1_0;
	wire w_dff_A_VV41j3Yu1_0;
	wire w_dff_A_eYDKNdy51_0;
	wire w_dff_A_7jW1el0h4_0;
	wire w_dff_A_yIE63RQf3_0;
	wire w_dff_A_fHoGpDUt4_0;
	wire w_dff_A_xG7OdISr2_0;
	wire w_dff_A_zwzzsLCO1_0;
	wire w_dff_A_DLRMPsiG2_0;
	wire w_dff_A_8MD8h5AY9_0;
	wire w_dff_A_5PgaDN0w5_0;
	wire w_dff_A_8KK8V2FU1_0;
	wire w_dff_A_c5MQTItK9_1;
	wire w_dff_A_4VOsYttB2_0;
	wire w_dff_A_6vGJ4YZW7_0;
	wire w_dff_A_hetQ05u51_0;
	wire w_dff_A_6rQxUhNr3_0;
	wire w_dff_A_Ug98WgI21_0;
	wire w_dff_A_hRGOfzIj6_0;
	wire w_dff_A_xQaZ1ijH3_0;
	wire w_dff_A_p1B058RH4_0;
	wire w_dff_A_W1Uf4Nqh9_0;
	wire w_dff_A_fC8vsPNg6_0;
	wire w_dff_A_AjwKw59x1_0;
	wire w_dff_A_gWvU7Oov8_0;
	wire w_dff_A_6bx00GY61_0;
	wire w_dff_A_7NoJdSJJ4_0;
	wire w_dff_A_q2aJEgkd5_0;
	wire w_dff_A_mtWUUNXM5_0;
	wire w_dff_A_VZSXlrIl4_0;
	wire w_dff_A_Y3J4dLad2_0;
	wire w_dff_A_VHl2Qsm91_0;
	wire w_dff_A_GjB697Ok2_0;
	wire w_dff_A_O2OfC5Ja7_0;
	wire w_dff_A_IYRYfPIz5_0;
	wire w_dff_A_EuZuotvZ8_0;
	wire w_dff_A_DvThwb6U7_0;
	wire w_dff_A_oLccsbfM2_0;
	wire w_dff_A_QfuqvVLH2_0;
	wire w_dff_A_xu1agTiB2_1;
	wire w_dff_A_lrqAy2L44_0;
	wire w_dff_A_2LhSkjYI2_0;
	wire w_dff_A_KwbHDxT89_0;
	wire w_dff_A_pKmkvdXK3_0;
	wire w_dff_A_wriAhwEy3_0;
	wire w_dff_A_zjFNdKXD4_0;
	wire w_dff_A_ABPQTlRW3_0;
	wire w_dff_A_oKvp4cll4_0;
	wire w_dff_A_7t0PUetP6_0;
	wire w_dff_A_Xrrzqlz08_0;
	wire w_dff_A_B2B8eAdk1_0;
	wire w_dff_A_11t3bD4x2_0;
	wire w_dff_A_CErQ3RXZ8_0;
	wire w_dff_A_TnYSVxcW8_0;
	wire w_dff_A_ONiOXrDK7_0;
	wire w_dff_A_jGqhMNPh6_0;
	wire w_dff_A_o6qYlUTn1_0;
	wire w_dff_A_t00olKhs4_0;
	wire w_dff_A_FF481w1r1_0;
	wire w_dff_A_tpxobTtJ5_0;
	wire w_dff_A_s0QMpRhn5_0;
	wire w_dff_A_TrAEPDb11_0;
	wire w_dff_A_rMDW1a3L4_0;
	wire w_dff_A_osaNfKJg7_0;
	wire w_dff_A_ufg8Bxsy6_0;
	wire w_dff_A_kvlVS9Fw7_0;
	wire w_dff_A_7bvST8917_1;
	wire w_dff_A_8BvXaxfK7_0;
	wire w_dff_A_TWtU7c1f1_0;
	wire w_dff_A_pQyHmwTQ6_0;
	wire w_dff_A_I9iFABSc3_0;
	wire w_dff_A_vWpyJEp82_0;
	wire w_dff_A_439c9kkD0_0;
	wire w_dff_A_EsHXbldW7_0;
	wire w_dff_A_oYriIHjx0_0;
	wire w_dff_A_b07LerSg3_0;
	wire w_dff_A_pyQfw6Du5_0;
	wire w_dff_A_QNnptJA61_0;
	wire w_dff_A_UYmtoCrC7_0;
	wire w_dff_A_rbA6QmCE6_0;
	wire w_dff_A_Xz54Jsmr9_0;
	wire w_dff_A_SHKX5rW55_0;
	wire w_dff_A_WiqDAh0n7_0;
	wire w_dff_A_EILdXOk58_0;
	wire w_dff_A_gLPZjr6N7_0;
	wire w_dff_A_DRuwiEfA0_0;
	wire w_dff_A_cbqdluqx1_0;
	wire w_dff_A_bnllwroc5_0;
	wire w_dff_A_MofP6H440_0;
	wire w_dff_A_4iIdPi8J8_0;
	wire w_dff_A_L0FaI5wy3_0;
	wire w_dff_A_I1Y7i4EX3_0;
	wire w_dff_A_6UWDOWSA1_1;
	wire w_dff_A_vn8vYwO54_0;
	wire w_dff_A_5Tgf4Bdv8_0;
	wire w_dff_A_jGFbwH2A8_0;
	wire w_dff_A_FWEA7P7f1_0;
	wire w_dff_A_VTdHVwMc6_0;
	wire w_dff_A_QrAC74wH8_0;
	wire w_dff_A_vpRfzOOT8_0;
	wire w_dff_A_Lno3wbIi4_0;
	wire w_dff_A_yj41Odb64_0;
	wire w_dff_A_ChCYih8I6_0;
	wire w_dff_A_D1cZPIEM3_0;
	wire w_dff_A_D9WFSkqf7_0;
	wire w_dff_A_lN9HBeEW6_0;
	wire w_dff_A_uOqTjRE81_0;
	wire w_dff_A_wW6giJO10_0;
	wire w_dff_A_9hd2PDPw2_0;
	wire w_dff_A_Yk2Zh7iN3_0;
	wire w_dff_A_m2Ezucv33_0;
	wire w_dff_A_KBDbDuUW1_0;
	wire w_dff_A_o8uZ0s8r0_0;
	wire w_dff_A_gxUG7u9A0_0;
	wire w_dff_A_4irXiDOc8_0;
	wire w_dff_A_vgs9vWSN5_0;
	wire w_dff_A_9QLzCYgU1_0;
	wire w_dff_A_cz8UdtXi3_0;
	wire w_dff_A_0pbaQvQh7_0;
	wire w_dff_A_l4pLZDe96_1;
	wire w_dff_A_dBuom1lU3_0;
	wire w_dff_A_LP2Tqdkx4_0;
	wire w_dff_A_oLc7MfjE4_0;
	wire w_dff_A_aJAFwLE92_0;
	wire w_dff_A_cjd4Il9M2_0;
	wire w_dff_A_bglDhIb82_0;
	wire w_dff_A_Ik0JOtjQ5_0;
	wire w_dff_A_JHpvRwiM7_0;
	wire w_dff_A_Pdd57MkJ3_0;
	wire w_dff_A_zZndK0pA8_0;
	wire w_dff_A_BkKRg6jA4_0;
	wire w_dff_A_ZCeitO3o9_0;
	wire w_dff_A_cutHzJP41_0;
	wire w_dff_A_WxeP7fne2_0;
	wire w_dff_A_USYmMaZP7_0;
	wire w_dff_A_GSzvcO6H5_0;
	wire w_dff_A_XAashtOp0_0;
	wire w_dff_A_ulDPMT8X6_0;
	wire w_dff_A_eho0bCVh8_0;
	wire w_dff_A_Ey6KZK048_0;
	wire w_dff_A_MehFAZ5B4_0;
	wire w_dff_A_NUne2LM84_0;
	wire w_dff_A_HWRUraAz0_0;
	wire w_dff_A_4RCNy5d40_0;
	wire w_dff_A_Iobuwp0F1_0;
	wire w_dff_A_WiUtrs525_0;
	wire w_dff_A_eaYLuokZ0_1;
	wire w_dff_A_HzgHeKjZ5_0;
	wire w_dff_A_7HfhwGA17_0;
	wire w_dff_A_lZsVeOrI8_0;
	wire w_dff_A_O4TWv1f76_0;
	wire w_dff_A_80PdiP009_0;
	wire w_dff_A_qnNiLbsw4_0;
	wire w_dff_A_1GMG43Jq0_0;
	wire w_dff_A_rRlWRf4x4_0;
	wire w_dff_A_ZE7WKBQ35_0;
	wire w_dff_A_nD04OMSb6_0;
	wire w_dff_A_bQU9CVZf9_0;
	wire w_dff_A_G9QN4jvF3_0;
	wire w_dff_A_PnvknPpP6_0;
	wire w_dff_A_UlMEasx26_0;
	wire w_dff_A_U6ITe5oR7_0;
	wire w_dff_A_1g68nLPq2_0;
	wire w_dff_A_WjyvEmKn7_0;
	wire w_dff_A_TNuN9byB5_0;
	wire w_dff_A_81v4I8Ew4_0;
	wire w_dff_A_scxawDpb4_0;
	wire w_dff_A_2sMe1RwB0_0;
	wire w_dff_A_uTljhGQn9_0;
	wire w_dff_A_tPSQsWNp6_0;
	wire w_dff_A_zimTBsAz4_0;
	wire w_dff_A_dhJQa4vr0_0;
	wire w_dff_A_AY2UsahH4_0;
	wire w_dff_A_c5Bpdw724_2;
	wire w_dff_A_OGQmfdLx7_0;
	wire w_dff_A_jDqFtL9x1_0;
	wire w_dff_A_3VuG7dLC2_0;
	wire w_dff_A_foG3f27D3_0;
	wire w_dff_A_VdeLpShU8_0;
	wire w_dff_A_Ipx5d0C58_0;
	wire w_dff_A_GX23GRlu3_0;
	wire w_dff_A_UG2DYt5s1_0;
	wire w_dff_A_P1SrnOu53_0;
	wire w_dff_A_m554hjvt9_0;
	wire w_dff_A_oF1LMhTv4_0;
	wire w_dff_A_W24l9afA7_0;
	wire w_dff_A_G0FVvffF3_0;
	wire w_dff_A_vX7o7EMY6_0;
	wire w_dff_A_uMYkhgM23_0;
	wire w_dff_A_mdksk9u94_0;
	wire w_dff_A_U6raieEU1_0;
	wire w_dff_A_MXbUDuQv9_0;
	wire w_dff_A_uAbWB8pv4_0;
	wire w_dff_A_oszbms297_0;
	wire w_dff_A_2CkbKNXS3_0;
	wire w_dff_A_Lhg4OACg7_0;
	wire w_dff_A_Dep6pJPm6_0;
	wire w_dff_A_vgStCyCG2_0;
	wire w_dff_A_9XGX6FUe8_0;
	wire w_dff_A_JtkNZIA12_1;
	wire w_dff_A_4WY3wfai9_0;
	wire w_dff_A_GDFVRGeD1_0;
	wire w_dff_A_6OXD3BVa8_0;
	wire w_dff_A_RZv2ZpI35_0;
	wire w_dff_A_q0UzIxli6_0;
	wire w_dff_A_E8rjbMvU3_0;
	wire w_dff_A_8xyq2cwx8_0;
	wire w_dff_A_pP9XxWYx0_0;
	wire w_dff_A_qSot8xif5_0;
	wire w_dff_A_0RlWnT658_0;
	wire w_dff_A_LY4MRAap9_0;
	wire w_dff_A_gWs4m90F6_0;
	wire w_dff_A_7CZWdSKy8_0;
	wire w_dff_A_2KkwN80j9_0;
	wire w_dff_A_2nBJX9c12_0;
	wire w_dff_A_yU2NPQD99_0;
	wire w_dff_A_MIdyw7zw1_0;
	wire w_dff_A_MTaFvIEq7_0;
	wire w_dff_A_4V4E08a95_0;
	wire w_dff_A_779SVaTk8_0;
	wire w_dff_A_lQAeoPEx4_0;
	wire w_dff_A_tApUQjOd3_0;
	wire w_dff_A_F0ZFqzmZ1_0;
	wire w_dff_A_wBQV3noA7_1;
	wire w_dff_A_vI62fLtD9_0;
	wire w_dff_A_fUbbepUN5_0;
	wire w_dff_A_RX7e92Sr5_0;
	wire w_dff_A_FBYe2Uek3_0;
	wire w_dff_A_x76m5M6j0_0;
	wire w_dff_A_IhIgCuvW5_0;
	wire w_dff_A_ECE7xGUS0_0;
	wire w_dff_A_MU1A8api7_0;
	wire w_dff_A_MCRGttNN8_0;
	wire w_dff_A_ePc4h8MT0_0;
	wire w_dff_A_UupNxGsL8_0;
	wire w_dff_A_nOJxS9Jg1_0;
	wire w_dff_A_EHkxXtRZ9_0;
	wire w_dff_A_xJw1jpc66_0;
	wire w_dff_A_QNczrOVf9_0;
	wire w_dff_A_wFZ3ijgK6_0;
	wire w_dff_A_Czqn3NUB0_0;
	wire w_dff_A_3eu3AR8j4_0;
	wire w_dff_A_UewIoyYU2_0;
	wire w_dff_A_3xUuhlZG1_0;
	wire w_dff_A_gZDCfb638_0;
	wire w_dff_A_e21azBOc4_0;
	wire w_dff_A_eUfihHxS6_0;
	wire w_dff_A_QqfC4UY36_1;
	wire w_dff_A_58tDZlpT4_0;
	wire w_dff_A_gjeEsi102_0;
	wire w_dff_A_m3fq1gcI0_0;
	wire w_dff_A_687HZ5zR4_0;
	wire w_dff_A_m1WaA9nU2_0;
	wire w_dff_A_aSmhwjCD5_0;
	wire w_dff_A_iwZZDib65_0;
	wire w_dff_A_GKzRefx24_0;
	wire w_dff_A_jAb0X6Xd5_0;
	wire w_dff_A_1yitxy5p3_0;
	wire w_dff_A_3d2dIPKw5_0;
	wire w_dff_A_plu2t9V74_0;
	wire w_dff_A_zxxe1Bm74_0;
	wire w_dff_A_gTeWXvt37_0;
	wire w_dff_A_Phyk4F5i4_0;
	wire w_dff_A_tIXNc8o60_0;
	wire w_dff_A_4S4oYqpz7_0;
	wire w_dff_A_2F5jgnQF5_0;
	wire w_dff_A_DPYnJdeI3_0;
	wire w_dff_A_ekwhykXE1_0;
	wire w_dff_A_B71DuFdv2_0;
	wire w_dff_A_fpcD7gLA1_0;
	wire w_dff_A_j8DZDwYc3_0;
	wire w_dff_A_wN1COxFA1_1;
	wire w_dff_A_UXhXXOMd1_0;
	wire w_dff_A_rNbJSLRS5_0;
	wire w_dff_A_tuQKwvRI1_0;
	wire w_dff_A_bKOgxtYK9_0;
	wire w_dff_A_7UzdgSs08_0;
	wire w_dff_A_gdi3aaTK4_0;
	wire w_dff_A_1I73ylGv1_0;
	wire w_dff_A_tr8P846U6_0;
	wire w_dff_A_jGtw6X0j1_0;
	wire w_dff_A_guz3Wv0c0_0;
	wire w_dff_A_HndTTY115_0;
	wire w_dff_A_VnetsG9r8_0;
	wire w_dff_A_RW8JLp5w8_0;
	wire w_dff_A_oLWOCoJM7_0;
	wire w_dff_A_zWtNHpzM6_0;
	wire w_dff_A_Kq3F9tLn8_0;
	wire w_dff_A_YvYsigHO8_0;
	wire w_dff_A_zw8snAnD6_0;
	wire w_dff_A_tMdYx3le6_0;
	wire w_dff_A_eIxVDBlg5_0;
	wire w_dff_A_g8CsW1aQ8_0;
	wire w_dff_A_1qxbycY08_0;
	wire w_dff_A_yW9PUCHW0_0;
	wire w_dff_A_bxKrKb576_1;
	wire w_dff_A_DOvQuR2g0_0;
	wire w_dff_A_seCvDu1X3_0;
	wire w_dff_A_IhzefiQx5_0;
	wire w_dff_A_vpXS2Vdr8_0;
	wire w_dff_A_lFABJ5my6_0;
	wire w_dff_A_MQCWwP5C6_0;
	wire w_dff_A_uDIsdkRv2_0;
	wire w_dff_A_5lO8EgHw1_0;
	wire w_dff_A_BwphV7pv4_0;
	wire w_dff_A_rN8FldBp4_0;
	wire w_dff_A_722YTZtX6_0;
	wire w_dff_A_JoVputvT0_0;
	wire w_dff_A_BUy5xOgU7_0;
	wire w_dff_A_ZUSa5Pzw9_0;
	wire w_dff_A_JsUWcN0v9_0;
	wire w_dff_A_vSBQXyM61_0;
	wire w_dff_A_VoVKRvgu9_0;
	wire w_dff_A_Cpcprkzt3_0;
	wire w_dff_A_ambPSS9G6_0;
	wire w_dff_A_M3oNdF5o9_0;
	wire w_dff_A_TpENOab82_0;
	wire w_dff_A_orjNISZW6_0;
	wire w_dff_A_HLEa5dzA4_0;
	wire w_dff_A_kJQVnKHp1_0;
	wire w_dff_A_DWZLgRVD1_0;
	wire w_dff_A_DNtqkJDi5_0;
	wire w_dff_A_lXPJgvRR0_1;
	wire w_dff_A_Qwp48rKC0_0;
	wire w_dff_A_61zFQQar8_0;
	wire w_dff_A_4Hbvc1QT5_0;
	wire w_dff_A_b7OF5PqX4_0;
	wire w_dff_A_yNZ0DHT43_0;
	wire w_dff_A_3Y0UdgSe4_0;
	wire w_dff_A_D7FTGf7z9_0;
	wire w_dff_A_ihh5PTuA2_0;
	wire w_dff_A_jgk8HQXv6_0;
	wire w_dff_A_u8CbI35r0_0;
	wire w_dff_A_tb4djUUj7_0;
	wire w_dff_A_vHKDxMlm4_0;
	wire w_dff_A_DCc2tDDX9_0;
	wire w_dff_A_IJH2Brp98_0;
	wire w_dff_A_oT0rsEt19_0;
	wire w_dff_A_xhIDkBHd1_0;
	wire w_dff_A_yvbSGFRa9_0;
	wire w_dff_A_p8j8ckKQ6_0;
	wire w_dff_A_82lYXakP8_0;
	wire w_dff_A_VTJIuf3R1_0;
	wire w_dff_A_d52LjHTs3_0;
	wire w_dff_A_ZYyu616n8_0;
	wire w_dff_A_o1A1ZTF14_0;
	wire w_dff_A_5t6PR8h28_0;
	wire w_dff_A_maAE4afP8_0;
	wire w_dff_A_MdPzYG3f5_0;
	wire w_dff_A_pZTZwLvs9_2;
	wire w_dff_A_uHCJWSLz2_0;
	wire w_dff_A_kqRh5e7s2_0;
	wire w_dff_A_WHezx8f96_0;
	wire w_dff_A_SorlaUJ19_0;
	wire w_dff_A_BVxgosoN9_0;
	wire w_dff_A_mzyaUjDb2_0;
	wire w_dff_A_bdtivdEl9_0;
	wire w_dff_A_gerkpQKj0_0;
	wire w_dff_A_3eVzLDRo1_0;
	wire w_dff_A_GAoxwLYc9_0;
	wire w_dff_A_kcHwxb6m7_0;
	wire w_dff_A_Q7x3eYi17_0;
	wire w_dff_A_668Mfmxb6_0;
	wire w_dff_A_7GAbXbNd6_0;
	wire w_dff_A_UiMGESzz3_0;
	wire w_dff_A_C1Z9Z9Kw0_0;
	wire w_dff_A_EsggchHu8_0;
	wire w_dff_A_8JVdgzId5_0;
	wire w_dff_A_JffIFJ3K9_0;
	wire w_dff_A_nfffUmky5_0;
	wire w_dff_A_QUuVqL9d8_0;
	wire w_dff_A_BsbD4sss9_0;
	wire w_dff_A_YHeMACUH6_0;
	wire w_dff_A_MP5Q4Jtz3_0;
	wire w_dff_A_eCUBokED4_1;
	wire w_dff_A_RnSNRzgX1_0;
	wire w_dff_A_bqKY1ank8_0;
	wire w_dff_A_EAREiTWX9_0;
	wire w_dff_A_frUEwr0U4_0;
	wire w_dff_A_rMX5vMuu1_0;
	wire w_dff_A_C1YHji7f5_0;
	wire w_dff_A_9jxMTJDm4_0;
	wire w_dff_A_z8WbIWXs3_0;
	wire w_dff_A_giDFloJd0_0;
	wire w_dff_A_VUJrQzoM0_0;
	wire w_dff_A_Jctpfofv4_0;
	wire w_dff_A_GYEIOdVE0_0;
	wire w_dff_A_5r0YoeG36_0;
	wire w_dff_A_eZlf5nWa3_0;
	wire w_dff_A_oD6ZDMiO5_0;
	wire w_dff_A_YsrsOS6p4_0;
	wire w_dff_A_ozKdBggJ7_0;
	wire w_dff_A_daKv7Bc13_0;
	wire w_dff_A_jPAMB7SH8_0;
	wire w_dff_A_pGBm3lmP3_0;
	wire w_dff_A_Nkq8LCm59_0;
	wire w_dff_A_78VAapmA2_0;
	wire w_dff_A_uO16OH9U4_0;
	wire w_dff_A_CsoApEUQ3_0;
	wire w_dff_A_AFPm4Vdq3_0;
	wire w_dff_A_FYQc2eRh8_2;
	wire w_dff_A_KLfJguYR5_0;
	wire w_dff_A_2J5FgEL79_0;
	wire w_dff_A_ogUKhVPc4_0;
	wire w_dff_A_IW9uyKCq2_0;
	wire w_dff_A_GTEHJHr11_0;
	wire w_dff_A_P8N7C4kW6_0;
	wire w_dff_A_BS1xp1Vg2_0;
	wire w_dff_A_HtbMXH465_0;
	wire w_dff_A_2WchYrdZ4_0;
	wire w_dff_A_WM9FRa6U2_0;
	wire w_dff_A_0wkvtvXM7_0;
	wire w_dff_A_5JJVyeKX7_0;
	wire w_dff_A_5u2NkGBQ0_0;
	wire w_dff_A_HPoNnLaf9_0;
	wire w_dff_A_zjM5TtBf8_0;
	wire w_dff_A_zKCY6qMT3_0;
	wire w_dff_A_ELSFogIC5_0;
	wire w_dff_A_LE6gOCuF0_0;
	wire w_dff_A_Xzaig07Y1_0;
	wire w_dff_A_ia8NrkBF7_0;
	wire w_dff_A_wVQwyipg4_0;
	wire w_dff_A_SdCvp1Oi1_0;
	wire w_dff_A_aivzwgzo6_0;
	wire w_dff_A_SCWtELTJ2_0;
	wire w_dff_A_ykhwGoNg6_2;
	wire w_dff_A_zYKSdpIZ3_0;
	wire w_dff_A_OvmsZo7W9_0;
	wire w_dff_A_ZeGmODYM2_0;
	wire w_dff_A_MHYM4iGP5_0;
	wire w_dff_A_XH2gTiXA7_0;
	wire w_dff_A_TCn667am8_0;
	wire w_dff_A_PfiLlCQu8_0;
	wire w_dff_A_lbb4ojyu0_0;
	wire w_dff_A_MJLIf0s93_0;
	wire w_dff_A_puwKJnUy9_0;
	wire w_dff_A_yj5UMYdx5_0;
	wire w_dff_A_Nta5g0kw6_0;
	wire w_dff_A_82BdCJjf1_0;
	wire w_dff_A_l4yGPLa39_0;
	wire w_dff_A_iqME2LgY7_0;
	wire w_dff_A_l0iQdBqX3_0;
	wire w_dff_A_cp4ruuO85_0;
	wire w_dff_A_YDpNDwXu7_0;
	wire w_dff_A_PliiTkmn7_0;
	wire w_dff_A_BC2gfvBM3_0;
	wire w_dff_A_GwSdQOOu6_0;
	wire w_dff_A_nPlPe1ob8_0;
	wire w_dff_A_LmjUrBmH6_0;
	wire w_dff_A_RVsCS7MB2_1;
	wire w_dff_A_JkGYnqp37_0;
	wire w_dff_A_cfLyZ6Eo5_0;
	wire w_dff_A_SZbOLmFu6_0;
	wire w_dff_A_iDp6iamO7_0;
	wire w_dff_A_lHiyOdug9_0;
	wire w_dff_A_53a1d0Hl8_0;
	wire w_dff_A_qKM3VT7L2_0;
	wire w_dff_A_i7Bvnpz17_0;
	wire w_dff_A_MEonsgzx3_0;
	wire w_dff_A_rIlrQLfQ1_0;
	wire w_dff_A_w9Tvkphw0_0;
	wire w_dff_A_5zMHCsLt9_0;
	wire w_dff_A_3iAiTpOV0_0;
	wire w_dff_A_6xOZ2zoO4_0;
	wire w_dff_A_pW2OTON93_0;
	wire w_dff_A_FDWcwLv91_0;
	wire w_dff_A_Zt5yfqYZ8_0;
	wire w_dff_A_WvD9IXS60_0;
	wire w_dff_A_PTzSNQ7D1_0;
	wire w_dff_A_JqcPZAzv8_0;
	wire w_dff_A_YJN1uq7d8_0;
	wire w_dff_A_LEKuSqlI2_0;
	wire w_dff_A_I6qbjVjc3_0;
	wire w_dff_A_SyOqRWI99_0;
	wire w_dff_A_41YS9oF26_0;
	wire w_dff_A_waTYV5cR5_2;
	wire w_dff_A_izDvKc0i8_0;
	wire w_dff_A_C2iaPpQG5_0;
	wire w_dff_A_WuyTt3mA2_0;
	wire w_dff_A_m9gheg8O1_0;
	wire w_dff_A_uGqKwkWM7_0;
	wire w_dff_A_YLXpkA7n9_0;
	wire w_dff_A_uOEKxG5v5_0;
	wire w_dff_A_TCRqD5Xv5_0;
	wire w_dff_A_kXB3zvQ49_0;
	wire w_dff_A_x4VsyKIq4_0;
	wire w_dff_A_jT5HZZph8_0;
	wire w_dff_A_u34PkPXl5_0;
	wire w_dff_A_nJlLwVJu7_0;
	wire w_dff_A_Xl74Pygk4_0;
	wire w_dff_A_i8rVA1lx6_0;
	wire w_dff_A_AL0ZVEBo8_0;
	wire w_dff_A_8jGHLbsB9_0;
	wire w_dff_A_2JJUyQSP0_0;
	wire w_dff_A_QSZQQ8Fx5_0;
	wire w_dff_A_f6GMjrkO1_0;
	wire w_dff_A_uEYRmXI90_0;
	wire w_dff_A_q600awFH0_0;
	wire w_dff_A_stwab5bd3_0;
	wire w_dff_A_fFEFrf1N6_1;
	wire w_dff_A_ePGjtmuI1_0;
	wire w_dff_A_05KYiG352_0;
	wire w_dff_A_BHdTPs5J3_0;
	wire w_dff_A_FVSLWOXv1_0;
	wire w_dff_A_gk9Bxukh2_0;
	wire w_dff_A_qWmYEwaA2_0;
	wire w_dff_A_0TFtlHzA5_0;
	wire w_dff_A_Vd2UvW9V4_0;
	wire w_dff_A_vu7rD0D33_0;
	wire w_dff_A_L3nmsKUv4_0;
	wire w_dff_A_1BwNLuVf4_0;
	wire w_dff_A_CThb3KVb2_0;
	wire w_dff_A_8bUTNctd4_0;
	wire w_dff_A_w8uLVGec0_0;
	wire w_dff_A_ngPergAi7_0;
	wire w_dff_A_QJrkdR7R0_0;
	wire w_dff_A_ircsX5gO4_0;
	wire w_dff_A_tVAvbdUP7_0;
	wire w_dff_A_Ppvba4146_0;
	wire w_dff_A_7hflrjqg9_0;
	wire w_dff_A_4CSQxZGI3_0;
	wire w_dff_A_rVXUJMHr0_0;
	wire w_dff_A_2ezQkJns7_0;
	wire w_dff_A_dqs0LX706_0;
	wire w_dff_A_kxQ9F6iF6_0;
	wire w_dff_A_lIGWgudn4_0;
	wire w_dff_A_SPuBfask4_2;
	wire w_dff_A_rbNpX5TS7_0;
	wire w_dff_A_rrknosF80_0;
	wire w_dff_A_5629ZiVs6_0;
	wire w_dff_A_183cX33w5_0;
	wire w_dff_A_PYToVF158_0;
	wire w_dff_A_7Kh27GAg9_0;
	wire w_dff_A_OHaUO1y64_0;
	wire w_dff_A_Bo04xigm6_0;
	wire w_dff_A_H75SOTxV2_0;
	wire w_dff_A_2wzeLbk01_0;
	wire w_dff_A_bic1SOq49_0;
	wire w_dff_A_wUBKt1Ue2_0;
	wire w_dff_A_nrCKNOix1_0;
	wire w_dff_A_ocV9Ai8E3_0;
	wire w_dff_A_gnfs6vU70_0;
	wire w_dff_A_yzmGzPvZ4_0;
	wire w_dff_A_ykuUuQvB5_0;
	wire w_dff_A_HUfBXmwX9_0;
	wire w_dff_A_wYMGb9mr3_0;
	wire w_dff_A_EVOOIMjv0_0;
	wire w_dff_A_NZKV8M4g0_0;
	wire w_dff_A_pQ1BT9QM1_0;
	wire w_dff_A_67PhyOSU5_0;
	wire w_dff_A_Y1zM5GUK2_0;
	wire w_dff_A_z14xZSHc4_0;
	wire w_dff_A_suIs7AHU8_2;
	wire w_dff_A_Zl7v79IQ9_0;
	wire w_dff_A_PETjAI8f2_0;
	wire w_dff_A_l9oPxLRk8_0;
	wire w_dff_A_AVwQQI0p1_0;
	wire w_dff_A_NhV9N0yC4_0;
	wire w_dff_A_OJc5aHP87_0;
	wire w_dff_A_hlpsEyBO5_0;
	wire w_dff_A_RFjQIz3m1_0;
	wire w_dff_A_oemZXJFF6_0;
	wire w_dff_A_5mSVcpfS8_0;
	wire w_dff_A_aTFF7Bz75_0;
	wire w_dff_A_llvpSK2r4_0;
	wire w_dff_A_7P89TQuY2_0;
	wire w_dff_A_z6e0Xm7G4_0;
	wire w_dff_A_iQK2QjP91_0;
	wire w_dff_A_i8PkzgsH9_0;
	wire w_dff_A_CukQvbtM3_0;
	wire w_dff_A_zwu4hvFi6_0;
	wire w_dff_A_K9vaKYfA5_0;
	wire w_dff_A_1hd6NNdi5_0;
	wire w_dff_A_JtpzOXIh8_2;
	wire w_dff_A_W0B7nnBb3_2;
	wire w_dff_A_zlWXXEha6_0;
	wire w_dff_A_cEnFVj2R0_0;
	wire w_dff_A_PTYC8VVJ5_0;
	wire w_dff_A_IAWs3H189_0;
	wire w_dff_A_opnM4RV00_0;
	wire w_dff_A_atu7ZuN71_0;
	wire w_dff_A_5YJ3wHUN2_2;
	wire w_dff_A_8CNtwnPS2_0;
	wire w_dff_A_DueYmvrc5_0;
	wire w_dff_A_Nou3FzeV2_0;
	wire w_dff_A_BKstMjwm9_0;
	wire w_dff_A_sVr04Vhk7_0;
	wire w_dff_A_f2arjRAU3_0;
	wire w_dff_A_FnZbY9aw9_2;
	wire w_dff_A_EFX9NOPw8_2;
	wire w_dff_A_lAfW20ax2_0;
	wire w_dff_A_ZFHJvkG30_0;
	wire w_dff_A_1vOj1xHI3_0;
	wire w_dff_A_IdmYffwd3_0;
	wire w_dff_A_ZF7HLi277_0;
	wire w_dff_A_f6pOu2Od7_0;
	wire w_dff_A_I3jd4brz3_0;
	wire w_dff_A_fhRfHGXa2_0;
	wire w_dff_A_nuIUhyMq8_0;
	wire w_dff_A_zwFTOozw9_0;
	wire w_dff_A_R2BZc8dp6_0;
	wire w_dff_A_PcmfU9xn5_0;
	wire w_dff_A_L0s6fA2O4_0;
	wire w_dff_A_vvm9IkcB8_0;
	wire w_dff_A_xvoXLmi80_2;
	wire w_dff_A_t1IMydfR8_0;
	wire w_dff_A_ywwcwF1e8_0;
	wire w_dff_A_deLvbHvC9_0;
	wire w_dff_A_xn75DcLZ9_0;
	wire w_dff_A_62RcKnEW0_0;
	wire w_dff_A_FFtHcsj90_0;
	wire w_dff_A_OoHBHvrF2_0;
	wire w_dff_A_cALSsssT3_0;
	wire w_dff_A_9gzshRGi6_0;
	wire w_dff_A_mOTFYfuF1_0;
	wire w_dff_A_bEzimCrj0_0;
	wire w_dff_A_vVe9MpS49_0;
	wire w_dff_A_KicLbHz72_0;
	wire w_dff_A_JiPxb9tQ0_0;
	wire w_dff_A_wU0cGKNP1_0;
	wire w_dff_A_uWOxwEd42_0;
	wire w_dff_A_7MoqT9H23_2;
	wire w_dff_A_B46vVDxc7_0;
	wire w_dff_A_6NKRiTk75_0;
	wire w_dff_A_yOUlHH040_0;
	wire w_dff_A_CDEzwtfL8_0;
	wire w_dff_A_cBqXkpBh4_0;
	wire w_dff_A_IcxbCaoa2_0;
	wire w_dff_A_YAu1NTss0_0;
	wire w_dff_A_JEBvJAwg2_0;
	wire w_dff_A_NGIN4VwU8_0;
	wire w_dff_A_KiDmOa0U3_0;
	wire w_dff_A_ENP4IxIW6_0;
	wire w_dff_A_0YB5Jr5P4_0;
	wire w_dff_A_1qWRxIx40_0;
	wire w_dff_A_IJO3GBE61_0;
	wire w_dff_A_zw4vaEnL5_0;
	wire w_dff_A_udJWUOW08_0;
	wire w_dff_A_0LrTun7G6_0;
	wire w_dff_A_iAHGgVal8_2;
	wire w_dff_A_I74EMTpF6_0;
	wire w_dff_A_Cf6IPG4M3_0;
	wire w_dff_A_pY6MpF7n5_0;
	wire w_dff_A_vYfE49QH5_0;
	wire w_dff_A_feGpzxdt6_0;
	wire w_dff_A_8TcsxdWB7_0;
	wire w_dff_A_GOlA94eU7_0;
	wire w_dff_A_vWC0rTMe7_0;
	wire w_dff_A_U6oIQtNI3_0;
	wire w_dff_A_l9eJBuwm9_0;
	wire w_dff_A_9M2BkVY72_0;
	wire w_dff_A_zKbseXdY1_0;
	wire w_dff_A_uxJcFMq33_0;
	wire w_dff_A_Ms3374Ws4_0;
	wire w_dff_A_A4lppiT41_0;
	wire w_dff_A_2C9hefZm2_0;
	wire w_dff_A_8ys43FSg0_0;
	wire w_dff_A_X3V7BDyI1_0;
	wire w_dff_A_HM031umB3_2;
	wire w_dff_A_d0l0xFV00_0;
	wire w_dff_A_0KKg9AiX0_0;
	wire w_dff_A_EkGfxABn4_0;
	wire w_dff_A_uJ6MDq2z2_0;
	wire w_dff_A_m3TIo9fU3_0;
	wire w_dff_A_NSHg86dI9_0;
	wire w_dff_A_7CHquQjY2_0;
	wire w_dff_A_InK39cDJ2_0;
	wire w_dff_A_gp7jE4gq9_0;
	wire w_dff_A_Mzlw1Mw87_0;
	wire w_dff_A_wy3cn1jy8_0;
	wire w_dff_A_jC9Luir46_0;
	wire w_dff_A_8OItUSdo4_2;
	wire w_dff_A_3puuAy3g7_0;
	wire w_dff_A_4BsxKgGG7_0;
	wire w_dff_A_JwQwdRJd9_0;
	wire w_dff_A_6IjPNA3O8_0;
	wire w_dff_A_iiXZWytQ1_0;
	wire w_dff_A_5hYABx7c3_0;
	wire w_dff_A_vYwIJLai4_0;
	wire w_dff_A_3W1KTZyC1_0;
	wire w_dff_A_lXjAEmul2_0;
	wire w_dff_A_CqmAF5Af3_0;
	wire w_dff_A_v4aVc9Fu2_0;
	wire w_dff_A_cIDyJVvq4_0;
	wire w_dff_A_bLSFTOs08_0;
	wire w_dff_A_inYkeue56_2;
	wire w_dff_A_2QOm5tTa3_0;
	wire w_dff_A_kkFX7zbn4_0;
	wire w_dff_A_n1DQ6Hyo9_0;
	wire w_dff_A_lePGEnyB7_0;
	wire w_dff_A_UYlZJ24e4_0;
	wire w_dff_A_1gygvsue4_0;
	wire w_dff_A_7ksOeu1C5_0;
	wire w_dff_A_ZpcKkR5f0_0;
	wire w_dff_A_MUP3aR5S5_0;
	wire w_dff_A_ail1nSTa5_0;
	wire w_dff_A_KW6wmjNm7_0;
	wire w_dff_A_mZxXFjU60_0;
	wire w_dff_A_zpQ5j4nn3_0;
	wire w_dff_A_YuMbcDwy0_2;
	wire w_dff_A_zW47M1Cl9_0;
	wire w_dff_A_9TFxO4n12_0;
	wire w_dff_A_YHGaE2yP9_0;
	wire w_dff_A_rmSN70mW1_0;
	wire w_dff_A_d4LYHthq4_0;
	wire w_dff_A_MGQenSyl3_0;
	wire w_dff_A_bp9JPRAO1_0;
	wire w_dff_A_5ebaY0NB4_0;
	wire w_dff_A_q61o1CA68_0;
	wire w_dff_A_9Q0UF8CC5_0;
	wire w_dff_A_iA2GrFun9_0;
	wire w_dff_A_DiLYexTM8_0;
	wire w_dff_A_otGRFl6Z0_0;
	wire w_dff_A_jCr3aH0v0_0;
	wire w_dff_A_0u8hVAdx7_0;
	wire w_dff_A_vKTTodl25_1;
	wire w_dff_A_1SNUD7x36_0;
	wire w_dff_A_6PtWGPY90_0;
	wire w_dff_A_lQ4MsByd2_0;
	wire w_dff_A_UMCOfAL28_0;
	wire w_dff_A_1gS5BeSi5_0;
	wire w_dff_A_dFYhTuT95_0;
	wire w_dff_A_Vo3arQaY1_0;
	wire w_dff_A_Qyma0x8A6_0;
	wire w_dff_A_5pnbjrPM1_0;
	wire w_dff_A_eYGLvuyF7_0;
	wire w_dff_A_nTsDorUF7_0;
	wire w_dff_A_IncAMnTY7_0;
	wire w_dff_A_XhGGlwzN4_0;
	wire w_dff_A_xnA5D6Te8_0;
	wire w_dff_A_wSfUCgex2_0;
	wire w_dff_A_09UngzC83_1;
	wire w_dff_A_lbqh8aXs4_0;
	wire w_dff_A_Ii9eUP6J9_0;
	wire w_dff_A_VT96i3Eu1_0;
	wire w_dff_A_bgmwtF6n8_0;
	wire w_dff_A_YUXqakBE9_0;
	wire w_dff_A_RsgyrWvQ6_0;
	wire w_dff_A_jS8xAlv22_0;
	wire w_dff_A_ib4bd8ej0_0;
	wire w_dff_A_YJtMS9783_0;
	wire w_dff_A_6dxDDTUe7_0;
	wire w_dff_A_zhIstHAG6_0;
	wire w_dff_A_E5az9PlC2_0;
	wire w_dff_A_9NdZmENl4_0;
	wire w_dff_A_csKpx9Jp4_0;
	wire w_dff_A_qQQyCCo16_0;
	wire w_dff_A_43cNgcPY5_1;
	wire w_dff_A_YuP3xOfQ8_0;
	wire w_dff_A_5OBjewN68_0;
	wire w_dff_A_NG6SqmY73_0;
	wire w_dff_A_MwFGg6kr2_0;
	wire w_dff_A_c06rjhzr0_0;
	wire w_dff_A_cpUVx2x90_0;
	wire w_dff_A_G6h6vG254_0;
	wire w_dff_A_iDdVmCoa8_0;
	wire w_dff_A_vvPkSMG95_0;
	wire w_dff_A_IES5gsep5_0;
	wire w_dff_A_v6PjrZEA2_0;
	wire w_dff_A_GBKT7SiV3_0;
	wire w_dff_A_bemAgK2w3_0;
	wire w_dff_A_tocXicLV2_2;
	wire w_dff_A_WDr71kD12_0;
	wire w_dff_A_9v82n2yI3_0;
	wire w_dff_A_oXJ2JL4K5_0;
	wire w_dff_A_nLZZwu0d9_0;
	wire w_dff_A_KEUS3aF96_0;
	wire w_dff_A_bwK6dfun3_0;
	wire w_dff_A_R2mLLwKi2_2;
	wire w_dff_A_S2pIv6CO0_0;
	wire w_dff_A_42pMZg4T4_0;
	wire w_dff_A_NgHBOebl6_0;
	wire w_dff_A_tUH3328i7_0;
	wire w_dff_A_OIzph72k1_0;
	wire w_dff_A_EnKcLzSO6_0;
	wire w_dff_A_hhUqR0WX6_0;
	wire w_dff_A_ehmDPqH06_0;
	wire w_dff_A_sDXAHvYj2_0;
	wire w_dff_A_kWtpVriV9_2;
	wire w_dff_A_LwuAuHUQ8_0;
	wire w_dff_A_uNXpyo9T9_0;
	wire w_dff_A_PNdJsUEN7_0;
	wire w_dff_A_WZE92r3R6_0;
	wire w_dff_A_tWIqak8g0_0;
	wire w_dff_A_jUZ9oWmy2_2;
	wire w_dff_A_7lBMX5AL7_0;
	wire w_dff_A_zh1NqjjA8_0;
	wire w_dff_A_CaHjyrq47_0;
	wire w_dff_A_uGeCxVnY4_0;
	wire w_dff_A_EBG2ZNh52_0;
	wire w_dff_A_nlrj6dYC5_0;
	wire w_dff_A_hQqt921o4_0;
	wire w_dff_A_sJgjWK4R2_0;
	wire w_dff_A_gJEkRr062_0;
	wire w_dff_A_u65loDku7_2;
	wire w_dff_A_bs3dCZUn0_2;
	wire w_dff_A_d5I7HYBu6_0;
	wire w_dff_A_UJ8zaBR02_0;
	wire w_dff_A_rZPzMJ467_0;
	wire w_dff_A_qUejOMLH0_0;
	wire w_dff_A_HHjaTWLT9_0;
	wire w_dff_A_amWUnRaU2_2;
	wire w_dff_A_tQHjlOxl1_0;
	wire w_dff_A_5ZJs7CSk4_0;
	wire w_dff_A_ilIpNWmd5_0;
	wire w_dff_A_7TSTUoMv9_0;
	wire w_dff_A_UZYjd2Ag6_0;
	wire w_dff_A_uq0eShYm4_0;
	wire w_dff_A_hR2WjjY39_2;
	wire w_dff_A_jTTaRbyp0_0;
	wire w_dff_A_4EyhSLwu4_0;
	wire w_dff_A_KRqJ0BaK6_0;
	wire w_dff_A_WDsUy5CT6_0;
	wire w_dff_A_9aEZRltC3_0;
	wire w_dff_A_Vtb3DA6f9_0;
	wire w_dff_A_QTIIJAgD2_0;
	wire w_dff_A_DEUGBpxE4_2;
	wire w_dff_A_3LDz5kvJ5_0;
	wire w_dff_A_AiWTeekL2_0;
	wire w_dff_A_Xhs6slgQ5_0;
	wire w_dff_A_QOxPoQFD5_0;
	wire w_dff_A_m7KmafAM5_0;
	wire w_dff_A_Vhi4oWOV7_0;
	wire w_dff_A_VRC1E4O96_0;
	wire w_dff_A_AdXSab4c0_2;
	wire w_dff_A_N8ez5Be21_0;
	wire w_dff_A_tDqTzf6y5_2;
	wire w_dff_A_WQJSos3G3_0;
	wire w_dff_A_4zuOeTUn8_0;
	wire w_dff_A_pC7Cjpvr8_2;
	wire w_dff_A_OhDGTutM7_0;
	wire w_dff_A_UhHQux9E2_0;
	wire w_dff_A_UcyusA3V2_0;
	wire w_dff_A_pWEqVmr15_2;
	wire w_dff_A_5qLxu60L2_0;
	wire w_dff_A_US3dwx8F9_0;
	wire w_dff_A_8yBKoaa10_0;
	wire w_dff_A_8GhQPmXM9_2;
	wire w_dff_A_HjdfjwHP0_0;
	wire w_dff_A_h8NITfi00_0;
	wire w_dff_A_pajs5PTE8_0;
	wire w_dff_A_VtObylxT9_0;
	wire w_dff_A_AUecmcjN3_0;
	wire w_dff_A_fFNtUUEv8_0;
	wire w_dff_A_hDPW3WLJ2_0;
	wire w_dff_A_9hEZxHmz4_0;
	wire w_dff_A_ALaRuceH1_0;
	wire w_dff_A_66IERIMB8_0;
	wire w_dff_A_cXIGW9EM4_0;
	wire w_dff_A_rnuc3wek8_2;
	wire w_dff_A_BfQSCrDb1_2;
	wire w_dff_A_egvpQFI02_0;
	wire w_dff_A_5p4R2p4r9_0;
	wire w_dff_A_bVZdos4u9_0;
	wire w_dff_A_LvjRIxn72_2;
	wire w_dff_A_03OrYuA79_0;
	wire w_dff_A_kt4TUV400_0;
	wire w_dff_A_yPsxLdux3_0;
	wire w_dff_A_FCyRsOtw1_0;
	wire w_dff_A_kiqIxzv19_0;
	wire w_dff_A_9o2BrKL15_2;
	wire w_dff_A_IT05QvZ51_0;
	wire w_dff_A_Jw8QBLpY4_0;
	wire w_dff_A_OHU5xNHF9_0;
	wire w_dff_A_l9zrvFcK4_0;
	wire w_dff_A_3sHBIowx4_0;
	wire w_dff_A_TB6D4vo83_2;
	wire w_dff_A_kzXUpVAQ3_0;
	wire w_dff_A_yrSKSwGe6_0;
	wire w_dff_A_UnIAgsPA8_0;
	wire w_dff_A_8I6MWYIg6_0;
	wire w_dff_A_epUeQGpD1_0;
	wire w_dff_A_MQg6KNYn1_0;
	wire w_dff_A_TJuwzeWO2_0;
	wire w_dff_A_VdTQjnjS5_2;
	wire w_dff_A_WiKhgYf83_0;
	wire w_dff_A_KgwgZIgZ2_0;
	wire w_dff_A_QXo3CoVZ5_0;
	wire w_dff_A_GBgOnyp30_0;
	wire w_dff_A_NZOmZO4Y7_0;
	wire w_dff_A_Qb6tYkXv7_0;
	wire w_dff_A_750Ii5E99_0;
	wire w_dff_A_Wcbiwsft1_0;
	wire w_dff_A_Q1XuOow32_0;
	wire w_dff_A_fScZqcuv5_0;
	wire w_dff_A_QmWurOe12_0;
	wire w_dff_A_BCSA4pmd6_0;
	wire w_dff_A_psZAIvTZ2_0;
	wire w_dff_A_m62Wobqa2_2;
	wire w_dff_A_FCyTexHS6_2;
	wire w_dff_A_WnsCWwMe4_2;
	wire w_dff_A_McKfIN4R6_0;
	wire w_dff_A_oUNzt51x0_0;
	wire w_dff_A_n9EzxzAo3_0;
	wire w_dff_A_uZI5p8W54_2;
	wire w_dff_A_iIojHEYs1_0;
	wire w_dff_A_PRcRXwuq3_0;
	wire w_dff_A_uw64MFh48_0;
	wire w_dff_A_I98csHOR7_2;
	wire w_dff_A_6N3kyfxF4_0;
	wire w_dff_A_sKhdD7Wt2_0;
	wire w_dff_A_zJXQwMGB2_0;
	wire w_dff_A_VLNjR7jZ4_0;
	wire w_dff_A_hGJOsO0k5_0;
	wire w_dff_A_haoo7cx71_0;
	wire w_dff_A_5ZluDnGQ9_0;
	wire w_dff_A_dIxTTPXT3_0;
	wire w_dff_A_1qrQnMpl8_0;
	wire w_dff_A_4R0St17A7_2;
	wire w_dff_A_zsKJpD2c6_0;
	wire w_dff_A_35N0Fvqu8_0;
	wire w_dff_A_BtEK6LCY6_0;
	wire w_dff_A_ANvtHa8D1_0;
	wire w_dff_A_1dR5VbvT5_0;
	wire w_dff_A_elF8ijvU6_0;
	wire w_dff_A_i7NT7RgT4_0;
	wire w_dff_A_oct90Hxu0_0;
	wire w_dff_A_e7pL2a0O3_0;
	wire w_dff_A_skNQEqNp0_0;
	wire w_dff_A_y4w19iT65_2;
	wire w_dff_A_mElVkZNX0_0;
	wire w_dff_A_VayYY6z12_0;
	wire w_dff_A_AfASEeIM2_0;
	wire w_dff_A_geMncHqD5_0;
	wire w_dff_A_46QOf2457_0;
	wire w_dff_A_tGjRx1Ix5_0;
	wire w_dff_A_b5gUGwaq7_0;
	wire w_dff_A_4w5cc3Js4_0;
	wire w_dff_A_6mjS7akw2_0;
	wire w_dff_A_t7vtsbDg7_0;
	wire w_dff_A_wFzNw0zK1_0;
	wire w_dff_A_8IAwW4586_2;
	wire w_dff_A_3OD6zrLh5_0;
	wire w_dff_A_E8YGGwpI7_0;
	wire w_dff_A_ZtYm5JhM5_0;
	wire w_dff_A_NGbqTv520_0;
	wire w_dff_A_A6SPs8pl3_0;
	wire w_dff_A_mklG8sXh5_0;
	wire w_dff_A_j6samyKX8_0;
	wire w_dff_A_NXvY6m2q2_0;
	wire w_dff_A_CKV8gBZk0_0;
	wire w_dff_A_OVhqUaDg6_0;
	wire w_dff_A_NKTSE4xa0_0;
	wire w_dff_A_fT0oI7CZ9_2;
	wire w_dff_A_v6CnyEDK5_0;
	wire w_dff_A_9QchQL8X3_0;
	wire w_dff_A_dJ15G3nQ0_0;
	wire w_dff_A_2ZHnWZN29_0;
	wire w_dff_A_FBjujRKJ9_0;
	wire w_dff_A_Ws2qIQNZ8_0;
	wire w_dff_A_DW6ZtK2o2_0;
	wire w_dff_A_16NqH9lB9_0;
	wire w_dff_A_aLzr4soI2_2;
	wire w_dff_A_upe8VqZn9_0;
	wire w_dff_A_KhCUihHE5_0;
	wire w_dff_A_MiSNBpgs1_0;
	wire w_dff_A_TxCmoLst1_0;
	wire w_dff_A_CDWnwMX23_0;
	wire w_dff_A_RTY0VLuR8_0;
	wire w_dff_A_BMocbvuz7_0;
	wire w_dff_A_IEHIzVXN2_0;
	wire w_dff_A_HZ5CMwWe8_0;
	wire w_dff_A_cdExsKih7_2;
	wire w_dff_A_lpCLC8Rj2_0;
	wire w_dff_A_NvIaDVch8_0;
	wire w_dff_A_Rmpyx10o1_0;
	wire w_dff_A_3GZdn6GM6_0;
	wire w_dff_A_WPUddwiv7_0;
	wire w_dff_A_XXNZpkSH3_0;
	wire w_dff_A_p61JToQo1_0;
	wire w_dff_A_TBBlG3BN4_0;
	wire w_dff_A_jWnpwcbL9_0;
	wire w_dff_A_JyIKjTuE8_2;
	wire w_dff_A_btQS2cq52_0;
	wire w_dff_A_cR6uF9Sp4_0;
	wire w_dff_A_SYzNlNCk8_0;
	wire w_dff_A_5QVUp1sS7_0;
	wire w_dff_A_nJdlwJI62_0;
	wire w_dff_A_g0MTB0zb6_0;
	wire w_dff_A_TP4r8a0M6_0;
	wire w_dff_A_DuHT5O0J3_0;
	wire w_dff_A_eJiXW1rd9_0;
	wire w_dff_A_G24BZ6301_0;
	wire w_dff_A_nn7hbzyR8_0;
	wire w_dff_A_3t7SkkRt9_2;
	wire w_dff_A_nyzdXdNn6_0;
	wire w_dff_A_pvq4Wukz3_0;
	wire w_dff_A_JNV2UDlX4_0;
	wire w_dff_A_iYXbgv9d9_0;
	wire w_dff_A_zYe5zPoI5_2;
	wire w_dff_A_VCfA5K0z6_0;
	wire w_dff_A_m13q9lbd0_0;
	wire w_dff_A_Xlosk2MW1_0;
	wire w_dff_A_jAs2ksC12_0;
	wire w_dff_A_zEMdixAm4_0;
	wire w_dff_A_rLt5lsyh1_0;
	wire w_dff_A_QNml90eu3_2;
	wire w_dff_A_8CmAzMgN4_0;
	wire w_dff_A_VP2UI0Kb1_0;
	wire w_dff_A_ttHqGC0e8_0;
	wire w_dff_A_JI1SDc3z1_0;
	jnot g0000(.din(w_G15_0[2]),.dout(w_dff_A_7bvST8917_1),.clk(gclk));
	jor g0001(.dina(G57),.dinb(w_G5_1[2]),.dout(w_dff_A_c5Bpdw724_2),.clk(gclk));
	jnot g0002(.din(G184),.dout(n317),.clk(gclk));
	jnot g0003(.din(G228),.dout(n318),.clk(gclk));
	jor g0004(.dina(n318),.dinb(n317),.dout(n319),.clk(gclk));
	jnot g0005(.din(G150),.dout(n320),.clk(gclk));
	jnot g0006(.din(G240),.dout(n321),.clk(gclk));
	jor g0007(.dina(n321),.dinb(n320),.dout(n322),.clk(gclk));
	jor g0008(.dina(n322),.dinb(n319),.dout(G404_fa_),.clk(gclk));
	jnot g0009(.din(G210),.dout(n324),.clk(gclk));
	jnot g0010(.din(G218),.dout(n325),.clk(gclk));
	jor g0011(.dina(n325),.dinb(n324),.dout(n326),.clk(gclk));
	jnot g0012(.din(G152),.dout(n327),.clk(gclk));
	jnot g0013(.din(G230),.dout(n328),.clk(gclk));
	jor g0014(.dina(n328),.dinb(n327),.dout(n329),.clk(gclk));
	jor g0015(.dina(n329),.dinb(n326),.dout(G406_fa_),.clk(gclk));
	jnot g0016(.din(G183),.dout(n331),.clk(gclk));
	jnot g0017(.din(G185),.dout(n332),.clk(gclk));
	jor g0018(.dina(n332),.dinb(n331),.dout(n333),.clk(gclk));
	jnot g0019(.din(G182),.dout(n334),.clk(gclk));
	jnot g0020(.din(G186),.dout(n335),.clk(gclk));
	jor g0021(.dina(n335),.dinb(n334),.dout(n336),.clk(gclk));
	jor g0022(.dina(n336),.dinb(n333),.dout(G408_fa_),.clk(gclk));
	jnot g0023(.din(G172),.dout(n338),.clk(gclk));
	jnot g0024(.din(G188),.dout(n339),.clk(gclk));
	jor g0025(.dina(n339),.dinb(n338),.dout(n340),.clk(gclk));
	jnot g0026(.din(G162),.dout(n341),.clk(gclk));
	jnot g0027(.din(G199),.dout(n342),.clk(gclk));
	jor g0028(.dina(n342),.dinb(n341),.dout(n343),.clk(gclk));
	jor g0029(.dina(n343),.dinb(n340),.dout(G410_fa_),.clk(gclk));
	jnot g0030(.din(G1197),.dout(n345),.clk(gclk));
	jor g0031(.dina(w_n345_0[1]),.dinb(w_G5_1[1]),.dout(w_dff_A_pZTZwLvs9_2),.clk(gclk));
	jnot g0032(.din(G133),.dout(n347),.clk(gclk));
	jnot g0033(.din(G134),.dout(n348),.clk(gclk));
	jor g0034(.dina(n348),.dinb(n347),.dout(n349),.clk(gclk));
	jor g0035(.dina(w_n349_0[1]),.dinb(w_G5_1[0]),.dout(w_dff_A_ykhwGoNg6_2),.clk(gclk));
	jand g0036(.dina(G163),.dinb(w_G1_1[2]),.dout(w_dff_A_SPuBfask4_2),.clk(gclk));
	jnot g0037(.din(w_G41_0[2]),.dout(n352),.clk(gclk));
	jor g0038(.dina(n352),.dinb(w_G18_58[2]),.dout(n353),.clk(gclk));
	jor g0039(.dina(w_n353_0[2]),.dinb(w_G3701_1[1]),.dout(n354),.clk(gclk));
	jnot g0040(.din(w_G18_58[1]),.dout(n355),.clk(gclk));
	jand g0041(.dina(w_G41_0[1]),.dinb(w_n355_26[1]),.dout(n356),.clk(gclk));
	jand g0042(.dina(w_G229_0[1]),.dinb(w_G18_58[0]),.dout(n357),.clk(gclk));
	jor g0043(.dina(w_dff_B_wb1SXgaB4_0),.dinb(w_n356_0[2]),.dout(n358),.clk(gclk));
	jand g0044(.dina(w_G3701_1[0]),.dinb(w_n355_26[0]),.dout(n359),.clk(gclk));
	jnot g0045(.din(w_n359_0[1]),.dout(n360),.clk(gclk));
	jor g0046(.dina(n360),.dinb(w_n358_0[1]),.dout(n361),.clk(gclk));
	jand g0047(.dina(n361),.dinb(w_n354_1[2]),.dout(n362),.clk(gclk));
	jxor g0048(.dina(w_n362_0[2]),.dinb(w_G4526_1[1]),.dout(w_dff_A_suIs7AHU8_2),.clk(gclk));
	jand g0049(.dina(w_G4528_0[2]),.dinb(w_G1496_0[2]),.dout(n364),.clk(gclk));
	jxor g0050(.dina(w_n364_0[1]),.dinb(w_G38_1[2]),.dout(n365),.clk(gclk));
	jnot g0051(.din(w_G3723_1[1]),.dout(n366),.clk(gclk));
	jand g0052(.dina(G235),.dinb(w_G18_57[2]),.dout(n367),.clk(gclk));
	jnot g0053(.din(n367),.dout(n368),.clk(gclk));
	jnot g0054(.din(G103),.dout(n369),.clk(gclk));
	jor g0055(.dina(n369),.dinb(w_G18_57[1]),.dout(n370),.clk(gclk));
	jand g0056(.dina(w_n370_0[1]),.dinb(n368),.dout(n371),.clk(gclk));
	jxor g0057(.dina(w_n371_1[1]),.dinb(w_n366_0[1]),.dout(n372),.clk(gclk));
	jand g0058(.dina(G236),.dinb(w_G18_57[0]),.dout(n373),.clk(gclk));
	jnot g0059(.din(n373),.dout(n374),.clk(gclk));
	jnot g0060(.din(G23),.dout(n375),.clk(gclk));
	jor g0061(.dina(n375),.dinb(w_G18_56[2]),.dout(n376),.clk(gclk));
	jand g0062(.dina(w_n376_0[1]),.dinb(n374),.dout(n377),.clk(gclk));
	jnot g0063(.din(w_n377_1[2]),.dout(n378),.clk(gclk));
	jxor g0064(.dina(n378),.dinb(w_G3717_2[1]),.dout(n379),.clk(gclk));
	jor g0065(.dina(w_n379_1[1]),.dinb(w_n372_1[2]),.dout(n380),.clk(gclk));
	jnot g0066(.din(w_G3711_1[1]),.dout(n381),.clk(gclk));
	jand g0067(.dina(G237),.dinb(w_G18_56[1]),.dout(n382),.clk(gclk));
	jnot g0068(.din(n382),.dout(n383),.clk(gclk));
	jnot g0069(.din(G26),.dout(n384),.clk(gclk));
	jor g0070(.dina(n384),.dinb(w_G18_56[0]),.dout(n385),.clk(gclk));
	jand g0071(.dina(w_n385_0[1]),.dinb(n383),.dout(n386),.clk(gclk));
	jxor g0072(.dina(w_n386_0[2]),.dinb(w_dff_B_Q2fH6EwX9_1),.dout(n387),.clk(gclk));
	jnot g0073(.din(w_G4526_1[0]),.dout(n388),.clk(gclk));
	jnot g0074(.din(w_G3701_0[2]),.dout(n389),.clk(gclk));
	jand g0075(.dina(w_n356_0[1]),.dinb(w_n389_0[1]),.dout(n390),.clk(gclk));
	jnot g0076(.din(w_G229_0[0]),.dout(n391),.clk(gclk));
	jor g0077(.dina(n391),.dinb(w_n355_25[2]),.dout(n392),.clk(gclk));
	jand g0078(.dina(n392),.dinb(w_n353_0[1]),.dout(n393),.clk(gclk));
	jand g0079(.dina(w_n359_0[0]),.dinb(n393),.dout(n394),.clk(gclk));
	jor g0080(.dina(n394),.dinb(w_n390_1[1]),.dout(n395),.clk(gclk));
	jnot g0081(.din(w_G3705_2[1]),.dout(n396),.clk(gclk));
	jnot g0082(.din(G238),.dout(n397),.clk(gclk));
	jor g0083(.dina(n397),.dinb(w_n355_25[1]),.dout(n398),.clk(gclk));
	jnot g0084(.din(G29),.dout(n399),.clk(gclk));
	jor g0085(.dina(n399),.dinb(w_G18_55[2]),.dout(n400),.clk(gclk));
	jand g0086(.dina(w_n400_0[1]),.dinb(n398),.dout(n401),.clk(gclk));
	jxor g0087(.dina(w_n401_1[2]),.dinb(w_dff_B_hZCxe38Z9_1),.dout(n402),.clk(gclk));
	jor g0088(.dina(w_n402_1[1]),.dinb(w_n395_0[2]),.dout(n403),.clk(gclk));
	jor g0089(.dina(w_n403_0[1]),.dinb(w_n388_0[2]),.dout(n404),.clk(gclk));
	jor g0090(.dina(w_n404_0[1]),.dinb(w_n387_1[2]),.dout(n405),.clk(gclk));
	jor g0091(.dina(w_n405_0[2]),.dinb(w_n380_0[2]),.dout(n406),.clk(gclk));
	jor g0092(.dina(w_n386_0[1]),.dinb(w_G3711_1[0]),.dout(n407),.clk(gclk));
	jor g0093(.dina(w_n402_1[0]),.dinb(w_n354_1[1]),.dout(n408),.clk(gclk));
	jor g0094(.dina(w_n408_0[1]),.dinb(w_n387_1[1]),.dout(n409),.clk(gclk));
	jand g0095(.dina(n409),.dinb(w_n407_0[2]),.dout(n410),.clk(gclk));
	jor g0096(.dina(w_n410_0[1]),.dinb(w_n380_0[1]),.dout(n411),.clk(gclk));
	jor g0097(.dina(w_n401_1[1]),.dinb(w_G3705_2[0]),.dout(n412),.clk(gclk));
	jor g0098(.dina(w_n412_0[2]),.dinb(w_n387_1[0]),.dout(n413),.clk(gclk));
	jor g0099(.dina(w_n413_1[1]),.dinb(w_n380_0[0]),.dout(n414),.clk(gclk));
	jor g0100(.dina(w_n371_1[0]),.dinb(w_G3723_1[0]),.dout(n415),.clk(gclk));
	jand g0101(.dina(w_n371_0[2]),.dinb(w_G3723_0[2]),.dout(n416),.clk(gclk));
	jor g0102(.dina(w_n377_1[1]),.dinb(w_G3717_2[0]),.dout(n417),.clk(gclk));
	jor g0103(.dina(w_n417_0[2]),.dinb(n416),.dout(n418),.clk(gclk));
	jand g0104(.dina(n418),.dinb(w_dff_B_K4gcKoet5_1),.dout(n419),.clk(gclk));
	jand g0105(.dina(w_n419_0[1]),.dinb(n414),.dout(n420),.clk(gclk));
	jand g0106(.dina(n420),.dinb(n411),.dout(n421),.clk(gclk));
	jand g0107(.dina(n421),.dinb(n406),.dout(n422),.clk(gclk));
	jnot g0108(.din(w_G3737_1[1]),.dout(n423),.clk(gclk));
	jand g0109(.dina(G233),.dinb(w_G18_55[1]),.dout(n424),.clk(gclk));
	jnot g0110(.din(n424),.dout(n425),.clk(gclk));
	jnot g0111(.din(G127),.dout(n426),.clk(gclk));
	jor g0112(.dina(n426),.dinb(w_G18_55[0]),.dout(n427),.clk(gclk));
	jand g0113(.dina(w_n427_0[1]),.dinb(n425),.dout(n428),.clk(gclk));
	jxor g0114(.dina(w_n428_0[2]),.dinb(w_dff_B_VUCu99sn2_1),.dout(n429),.clk(gclk));
	jnot g0115(.din(w_G3729_1[1]),.dout(n430),.clk(gclk));
	jand g0116(.dina(G234),.dinb(w_G18_54[2]),.dout(n431),.clk(gclk));
	jnot g0117(.din(n431),.dout(n432),.clk(gclk));
	jnot g0118(.din(G130),.dout(n433),.clk(gclk));
	jor g0119(.dina(n433),.dinb(w_G18_54[1]),.dout(n434),.clk(gclk));
	jand g0120(.dina(w_n434_0[1]),.dinb(n432),.dout(n435),.clk(gclk));
	jxor g0121(.dina(w_n435_1[1]),.dinb(w_n430_0[1]),.dout(n436),.clk(gclk));
	jor g0122(.dina(w_n436_0[1]),.dinb(w_n429_2[1]),.dout(n437),.clk(gclk));
	jand g0123(.dina(G231),.dinb(w_G18_54[0]),.dout(n438),.clk(gclk));
	jnot g0124(.din(n438),.dout(n439),.clk(gclk));
	jnot g0125(.din(G100),.dout(n440),.clk(gclk));
	jor g0126(.dina(n440),.dinb(w_G18_53[2]),.dout(n441),.clk(gclk));
	jand g0127(.dina(w_n441_0[1]),.dinb(n439),.dout(n442),.clk(gclk));
	jor g0128(.dina(w_n442_0[2]),.dinb(w_G3749_1[1]),.dout(n443),.clk(gclk));
	jnot g0129(.din(w_n443_0[1]),.dout(n444),.clk(gclk));
	jand g0130(.dina(w_n442_0[1]),.dinb(w_G3749_1[0]),.dout(n445),.clk(gclk));
	jor g0131(.dina(w_n445_0[1]),.dinb(n444),.dout(n446),.clk(gclk));
	jand g0132(.dina(G232),.dinb(w_G18_53[1]),.dout(n447),.clk(gclk));
	jand g0133(.dina(w_dff_B_Xj2Too0S0_0),.dinb(w_n355_25[0]),.dout(n448),.clk(gclk));
	jor g0134(.dina(w_n448_0[1]),.dinb(w_dff_B_GRmSurMV5_1),.dout(n449),.clk(gclk));
	jxor g0135(.dina(w_n449_0[2]),.dinb(w_G3743_1[2]),.dout(n450),.clk(gclk));
	jor g0136(.dina(w_n450_0[2]),.dinb(w_n446_1[1]),.dout(n451),.clk(gclk));
	jor g0137(.dina(n451),.dinb(w_n437_0[1]),.dout(n452),.clk(gclk));
	jor g0138(.dina(w_n452_0[1]),.dinb(w_n422_1[2]),.dout(n453),.clk(gclk));
	jnot g0139(.din(w_n449_0[1]),.dout(n454),.clk(gclk));
	jor g0140(.dina(w_n454_0[1]),.dinb(w_G3743_1[1]),.dout(n455),.clk(gclk));
	jand g0141(.dina(w_n454_0[0]),.dinb(w_G3743_1[0]),.dout(n456),.clk(gclk));
	jor g0142(.dina(w_n428_0[1]),.dinb(w_G3737_1[0]),.dout(n457),.clk(gclk));
	jor g0143(.dina(w_n435_1[0]),.dinb(w_G3729_1[0]),.dout(n458),.clk(gclk));
	jor g0144(.dina(w_n458_0[2]),.dinb(w_n429_2[0]),.dout(n459),.clk(gclk));
	jand g0145(.dina(n459),.dinb(w_n457_0[1]),.dout(n460),.clk(gclk));
	jor g0146(.dina(w_n460_0[2]),.dinb(w_n456_0[2]),.dout(n461),.clk(gclk));
	jand g0147(.dina(w_n461_0[1]),.dinb(w_n455_0[1]),.dout(n462),.clk(gclk));
	jand g0148(.dina(w_n462_0[2]),.dinb(w_n443_0[0]),.dout(n463),.clk(gclk));
	jor g0149(.dina(n463),.dinb(w_n445_0[0]),.dout(n464),.clk(gclk));
	jand g0150(.dina(w_n464_0[1]),.dinb(n453),.dout(n465),.clk(gclk));
	jnot g0151(.din(w_G4415_1[1]),.dout(n466),.clk(gclk));
	jand g0152(.dina(G223),.dinb(w_G18_53[0]),.dout(n467),.clk(gclk));
	jand g0153(.dina(w_dff_B_fMrwYs659_0),.dinb(w_n355_24[2]),.dout(n468),.clk(gclk));
	jor g0154(.dina(w_n468_0[1]),.dinb(w_dff_B_zliV9cO33_1),.dout(n469),.clk(gclk));
	jxor g0155(.dina(w_n469_1[1]),.dinb(w_n466_0[1]),.dout(n470),.clk(gclk));
	jnot g0156(.din(w_G4400_0[2]),.dout(n471),.clk(gclk));
	jand g0157(.dina(G226),.dinb(w_G18_52[2]),.dout(n472),.clk(gclk));
	jand g0158(.dina(w_dff_B_LQ7pEVUH6_0),.dinb(w_n355_24[1]),.dout(n473),.clk(gclk));
	jor g0159(.dina(w_n473_0[1]),.dinb(w_dff_B_ZBbtVsur2_1),.dout(n474),.clk(gclk));
	jxor g0160(.dina(w_n474_1[1]),.dinb(w_n471_0[2]),.dout(n475),.clk(gclk));
	jand g0161(.dina(G217),.dinb(w_G18_52[1]),.dout(n476),.clk(gclk));
	jand g0162(.dina(w_dff_B_COBhojxa7_0),.dinb(w_n355_24[0]),.dout(n477),.clk(gclk));
	jor g0163(.dina(w_n477_0[1]),.dinb(w_dff_B_m5PZQapt5_1),.dout(n478),.clk(gclk));
	jnot g0164(.din(w_n478_0[1]),.dout(n479),.clk(gclk));
	jxor g0165(.dina(w_n479_0[1]),.dinb(w_G4394_1[1]),.dout(n480),.clk(gclk));
	jand g0166(.dina(w_n480_1[1]),.dinb(w_n475_1[1]),.dout(n481),.clk(gclk));
	jnot g0167(.din(w_G4410_1[1]),.dout(n482),.clk(gclk));
	jand g0168(.dina(G224),.dinb(w_G18_52[0]),.dout(n483),.clk(gclk));
	jand g0169(.dina(w_dff_B_Dw4rdbuH0_0),.dinb(w_n355_23[2]),.dout(n484),.clk(gclk));
	jor g0170(.dina(w_n484_0[1]),.dinb(w_dff_B_HiEtNCOm9_1),.dout(n485),.clk(gclk));
	jxor g0171(.dina(w_n485_0[2]),.dinb(w_n482_0[1]),.dout(n486),.clk(gclk));
	jand g0172(.dina(G225),.dinb(w_G18_51[2]),.dout(n487),.clk(gclk));
	jand g0173(.dina(w_dff_B_rIPQjVRj5_0),.dinb(w_n355_23[1]),.dout(n488),.clk(gclk));
	jor g0174(.dina(w_n488_0[1]),.dinb(w_dff_B_esNCd9Ls0_1),.dout(n489),.clk(gclk));
	jnot g0175(.din(w_n489_0[1]),.dout(n490),.clk(gclk));
	jxor g0176(.dina(w_n490_0[2]),.dinb(w_G4405_1[2]),.dout(n491),.clk(gclk));
	jand g0177(.dina(w_n491_1[1]),.dinb(w_n486_0[2]),.dout(n492),.clk(gclk));
	jand g0178(.dina(n492),.dinb(w_n481_0[2]),.dout(n493),.clk(gclk));
	jand g0179(.dina(w_n493_0[1]),.dinb(w_n470_0[2]),.dout(n494),.clk(gclk));
	jnot g0180(.din(w_n494_0[1]),.dout(n495),.clk(gclk));
	jor g0181(.dina(w_dff_B_kxkwTheF8_0),.dinb(w_n465_0[2]),.dout(n496),.clk(gclk));
	jnot g0182(.din(w_n469_1[0]),.dout(n497),.clk(gclk));
	jand g0183(.dina(n497),.dinb(w_G4415_1[0]),.dout(n498),.clk(gclk));
	jand g0184(.dina(w_n469_0[2]),.dinb(w_n466_0[0]),.dout(n499),.clk(gclk));
	jnot g0185(.din(n499),.dout(n500),.clk(gclk));
	jand g0186(.dina(w_n485_0[1]),.dinb(w_n482_0[0]),.dout(n501),.clk(gclk));
	jnot g0187(.din(n501),.dout(n502),.clk(gclk));
	jnot g0188(.din(w_n485_0[0]),.dout(n503),.clk(gclk));
	jand g0189(.dina(w_n503_0[1]),.dinb(w_G4410_1[0]),.dout(n504),.clk(gclk));
	jand g0190(.dina(w_n490_0[1]),.dinb(w_G4405_1[1]),.dout(n505),.clk(gclk));
	jnot g0191(.din(w_n475_1[0]),.dout(n506),.clk(gclk));
	jor g0192(.dina(w_n479_0[0]),.dinb(w_G4394_1[0]),.dout(n507),.clk(gclk));
	jor g0193(.dina(w_n507_1[2]),.dinb(n506),.dout(n508),.clk(gclk));
	jand g0194(.dina(w_n474_1[0]),.dinb(w_n471_0[1]),.dout(n509),.clk(gclk));
	jnot g0195(.din(w_n509_0[1]),.dout(n510),.clk(gclk));
	jor g0196(.dina(w_n490_0[0]),.dinb(w_G4405_1[0]),.dout(n511),.clk(gclk));
	jand g0197(.dina(n511),.dinb(w_n510_0[1]),.dout(n512),.clk(gclk));
	jand g0198(.dina(w_n512_0[1]),.dinb(w_n508_0[1]),.dout(n513),.clk(gclk));
	jor g0199(.dina(n513),.dinb(w_n505_0[1]),.dout(n514),.clk(gclk));
	jor g0200(.dina(w_n514_0[2]),.dinb(w_dff_B_fczQLOE96_1),.dout(n515),.clk(gclk));
	jand g0201(.dina(n515),.dinb(w_n502_0[1]),.dout(n516),.clk(gclk));
	jand g0202(.dina(w_n516_0[2]),.dinb(w_dff_B_SZj7H64q1_1),.dout(n517),.clk(gclk));
	jor g0203(.dina(n517),.dinb(w_dff_B_2yFhqfr89_1),.dout(n518),.clk(gclk));
	jand g0204(.dina(w_n518_0[1]),.dinb(n496),.dout(n519),.clk(gclk));
	jnot g0205(.din(w_G4427_0[1]),.dout(n520),.clk(gclk));
	jand g0206(.dina(G221),.dinb(w_G18_51[1]),.dout(n521),.clk(gclk));
	jand g0207(.dina(w_dff_B_yFaDUAMU1_0),.dinb(w_n355_23[0]),.dout(n522),.clk(gclk));
	jor g0208(.dina(w_n522_0[1]),.dinb(w_dff_B_97p8fcFJ9_1),.dout(n523),.clk(gclk));
	jxor g0209(.dina(w_n523_0[2]),.dinb(w_n520_0[2]),.dout(n524),.clk(gclk));
	jnot g0210(.din(w_G4420_0[2]),.dout(n525),.clk(gclk));
	jand g0211(.dina(G222),.dinb(w_G18_51[0]),.dout(n526),.clk(gclk));
	jand g0212(.dina(w_dff_B_F8ISny507_0),.dinb(w_n355_22[2]),.dout(n527),.clk(gclk));
	jor g0213(.dina(w_n527_0[1]),.dinb(w_dff_B_I0QzRyjh5_1),.dout(n528),.clk(gclk));
	jxor g0214(.dina(w_n528_1[1]),.dinb(w_n525_0[2]),.dout(n529),.clk(gclk));
	jand g0215(.dina(w_n529_0[1]),.dinb(w_n524_2[1]),.dout(n530),.clk(gclk));
	jnot g0216(.din(w_G4437_0[2]),.dout(n531),.clk(gclk));
	jand g0217(.dina(G219),.dinb(w_G18_50[2]),.dout(n532),.clk(gclk));
	jand g0218(.dina(w_dff_B_Wt9cimE64_0),.dinb(w_n355_22[1]),.dout(n533),.clk(gclk));
	jor g0219(.dina(w_n533_0[1]),.dinb(w_dff_B_z56kjaHO9_1),.dout(n534),.clk(gclk));
	jxor g0220(.dina(w_n534_1[1]),.dinb(w_n531_0[2]),.dout(n535),.clk(gclk));
	jnot g0221(.din(w_G4432_1[1]),.dout(n536),.clk(gclk));
	jand g0222(.dina(G220),.dinb(w_G18_50[1]),.dout(n537),.clk(gclk));
	jand g0223(.dina(w_dff_B_VzS5hBIf6_0),.dinb(w_n355_22[0]),.dout(n538),.clk(gclk));
	jor g0224(.dina(w_n538_0[1]),.dinb(w_dff_B_dHFxbENz8_1),.dout(n539),.clk(gclk));
	jxor g0225(.dina(w_n539_1[1]),.dinb(w_n536_0[1]),.dout(n540),.clk(gclk));
	jand g0226(.dina(w_n540_0[2]),.dinb(w_n535_1[1]),.dout(n541),.clk(gclk));
	jand g0227(.dina(n541),.dinb(w_n530_0[1]),.dout(n542),.clk(gclk));
	jnot g0228(.din(w_n542_0[1]),.dout(n543),.clk(gclk));
	jor g0229(.dina(w_dff_B_o0PEMrjh5_0),.dinb(w_n519_0[1]),.dout(n544),.clk(gclk));
	jnot g0230(.din(w_n534_1[0]),.dout(n545),.clk(gclk));
	jand g0231(.dina(n545),.dinb(w_G4437_0[1]),.dout(n546),.clk(gclk));
	jnot g0232(.din(n546),.dout(n547),.clk(gclk));
	jand g0233(.dina(w_n534_0[2]),.dinb(w_n531_0[1]),.dout(n548),.clk(gclk));
	jand g0234(.dina(w_n539_1[0]),.dinb(w_n536_0[0]),.dout(n549),.clk(gclk));
	jnot g0235(.din(w_n539_0[2]),.dout(n550),.clk(gclk));
	jand g0236(.dina(n550),.dinb(w_G4432_1[0]),.dout(n551),.clk(gclk));
	jnot g0237(.din(w_n551_0[1]),.dout(n552),.clk(gclk));
	jand g0238(.dina(w_n523_0[1]),.dinb(w_n520_0[1]),.dout(n553),.clk(gclk));
	jand g0239(.dina(w_n528_1[0]),.dinb(w_n525_0[1]),.dout(n554),.clk(gclk));
	jand g0240(.dina(w_n554_0[2]),.dinb(w_n524_2[0]),.dout(n555),.clk(gclk));
	jor g0241(.dina(n555),.dinb(w_n553_0[1]),.dout(n556),.clk(gclk));
	jand g0242(.dina(w_n556_0[2]),.dinb(w_n552_0[1]),.dout(n557),.clk(gclk));
	jor g0243(.dina(w_n557_0[1]),.dinb(w_n549_0[1]),.dout(n558),.clk(gclk));
	jor g0244(.dina(w_n558_0[2]),.dinb(w_dff_B_OM3RWix06_1),.dout(n559),.clk(gclk));
	jand g0245(.dina(n559),.dinb(w_dff_B_JtxtzyDc6_1),.dout(n560),.clk(gclk));
	jnot g0246(.din(w_n560_0[1]),.dout(n561),.clk(gclk));
	jand g0247(.dina(w_dff_B_LlkusSHQ2_0),.dinb(n544),.dout(n562),.clk(gclk));
	jnot g0248(.din(w_G2236_1[1]),.dout(n563),.clk(gclk));
	jand g0249(.dina(G12),.dinb(G9),.dout(n564),.clk(gclk));
	jnot g0250(.din(w_n564_0[2]),.dout(n565),.clk(gclk));
	jor g0251(.dina(w_dff_B_fEbOTJcJ7_0),.dinb(w_n355_21[2]),.dout(n566),.clk(gclk));
	jand g0252(.dina(n566),.dinb(w_n565_10[1]),.dout(n567),.clk(gclk));
	jxor g0253(.dina(w_n567_1[1]),.dinb(w_n563_0[1]),.dout(n568),.clk(gclk));
	jnot g0254(.din(w_G2218_0[2]),.dout(n569),.clk(gclk));
	jand g0255(.dina(w_dff_B_YG35GxyW3_0),.dinb(w_n355_21[1]),.dout(n570),.clk(gclk));
	jand g0256(.dina(G160),.dinb(w_G18_50[0]),.dout(n571),.clk(gclk));
	jor g0257(.dina(w_dff_B_qkHOgTH72_0),.dinb(w_n570_0[1]),.dout(n572),.clk(gclk));
	jxor g0258(.dina(w_n572_1[1]),.dinb(w_n569_0[2]),.dout(n573),.clk(gclk));
	jnot g0259(.din(w_G2211_0[2]),.dout(n574),.clk(gclk));
	jand g0260(.dina(w_dff_B_8B9DvCFK8_0),.dinb(w_n355_21[0]),.dout(n575),.clk(gclk));
	jand g0261(.dina(G151),.dinb(w_G18_49[2]),.dout(n576),.clk(gclk));
	jor g0262(.dina(w_dff_B_0zBk2jvP7_0),.dinb(w_n575_0[1]),.dout(n577),.clk(gclk));
	jxor g0263(.dina(w_n577_0[2]),.dinb(w_n574_0[1]),.dout(n578),.clk(gclk));
	jand g0264(.dina(w_n578_1[1]),.dinb(w_n573_1[1]),.dout(n579),.clk(gclk));
	jnot g0265(.din(w_G2230_1[1]),.dout(n580),.clk(gclk));
	jand g0266(.dina(w_dff_B_9kVB0bVY5_0),.dinb(w_n355_20[2]),.dout(n581),.clk(gclk));
	jand g0267(.dina(G158),.dinb(w_G18_49[1]),.dout(n582),.clk(gclk));
	jor g0268(.dina(w_dff_B_3aDczcGY4_0),.dinb(w_n581_0[1]),.dout(n583),.clk(gclk));
	jxor g0269(.dina(w_n583_1[1]),.dinb(w_n580_0[1]),.dout(n584),.clk(gclk));
	jnot g0270(.din(w_G2224_1[1]),.dout(n585),.clk(gclk));
	jand g0271(.dina(w_dff_B_EydYX5KM5_0),.dinb(w_n355_20[1]),.dout(n586),.clk(gclk));
	jand g0272(.dina(G159),.dinb(w_G18_49[0]),.dout(n587),.clk(gclk));
	jor g0273(.dina(w_dff_B_HUTl7wB53_0),.dinb(w_n586_0[1]),.dout(n588),.clk(gclk));
	jxor g0274(.dina(w_n588_1[1]),.dinb(w_n585_0[1]),.dout(n589),.clk(gclk));
	jand g0275(.dina(w_n589_1[1]),.dinb(w_n584_0[2]),.dout(n590),.clk(gclk));
	jand g0276(.dina(n590),.dinb(w_n579_0[2]),.dout(n591),.clk(gclk));
	jand g0277(.dina(w_n591_0[1]),.dinb(w_n568_0[2]),.dout(n592),.clk(gclk));
	jnot g0278(.din(w_n592_0[1]),.dout(n593),.clk(gclk));
	jor g0279(.dina(w_dff_B_DshOYC767_0),.dinb(w_n562_0[2]),.dout(n594),.clk(gclk));
	jand g0280(.dina(w_n567_1[0]),.dinb(w_n563_0[0]),.dout(n595),.clk(gclk));
	jnot g0281(.din(n595),.dout(n596),.clk(gclk));
	jnot g0282(.din(w_n567_0[2]),.dout(n597),.clk(gclk));
	jand g0283(.dina(n597),.dinb(w_G2236_1[0]),.dout(n598),.clk(gclk));
	jand g0284(.dina(w_n583_1[0]),.dinb(w_n580_0[0]),.dout(n599),.clk(gclk));
	jnot g0285(.din(w_n599_0[1]),.dout(n600),.clk(gclk));
	jnot g0286(.din(w_n583_0[2]),.dout(n601),.clk(gclk));
	jand g0287(.dina(n601),.dinb(w_G2230_1[0]),.dout(n602),.clk(gclk));
	jnot g0288(.din(w_n588_1[0]),.dout(n603),.clk(gclk));
	jand g0289(.dina(n603),.dinb(w_G2224_1[0]),.dout(n604),.clk(gclk));
	jnot g0290(.din(n604),.dout(n605),.clk(gclk));
	jand g0291(.dina(w_n577_0[1]),.dinb(w_n574_0[0]),.dout(n606),.clk(gclk));
	jand g0292(.dina(w_n606_1[2]),.dinb(w_n573_1[0]),.dout(n607),.clk(gclk));
	jand g0293(.dina(w_n572_1[0]),.dinb(w_n569_0[1]),.dout(n608),.clk(gclk));
	jand g0294(.dina(w_n588_0[2]),.dinb(w_n585_0[0]),.dout(n609),.clk(gclk));
	jor g0295(.dina(n609),.dinb(w_n608_0[2]),.dout(n610),.clk(gclk));
	jor g0296(.dina(w_n610_0[1]),.dinb(w_n607_0[1]),.dout(n611),.clk(gclk));
	jand g0297(.dina(n611),.dinb(w_n605_0[1]),.dout(n612),.clk(gclk));
	jnot g0298(.din(w_n612_0[1]),.dout(n613),.clk(gclk));
	jor g0299(.dina(w_n613_0[2]),.dinb(w_dff_B_eIy8GjQg9_1),.dout(n614),.clk(gclk));
	jand g0300(.dina(n614),.dinb(w_dff_B_AfjZREIl4_1),.dout(n615),.clk(gclk));
	jor g0301(.dina(w_n615_1[1]),.dinb(w_dff_B_MzJuDY4q3_1),.dout(n616),.clk(gclk));
	jand g0302(.dina(n616),.dinb(w_dff_B_fRSBs2f97_1),.dout(n617),.clk(gclk));
	jand g0303(.dina(w_n617_0[1]),.dinb(n594),.dout(n618),.clk(gclk));
	jnot g0304(.din(w_G2247_0[2]),.dout(n619),.clk(gclk));
	jor g0305(.dina(w_dff_B_CjTSjO7E8_0),.dinb(w_n355_20[0]),.dout(n620),.clk(gclk));
	jand g0306(.dina(w_n620_0[1]),.dinb(w_n565_10[0]),.dout(n621),.clk(gclk));
	jxor g0307(.dina(w_n621_0[2]),.dinb(w_n619_0[1]),.dout(n622),.clk(gclk));
	jnot g0308(.din(w_G2239_0[2]),.dout(n623),.clk(gclk));
	jor g0309(.dina(w_dff_B_tR2tjaxm1_0),.dinb(w_n355_19[2]),.dout(n624),.clk(gclk));
	jand g0310(.dina(w_n624_0[1]),.dinb(w_n565_9[2]),.dout(n625),.clk(gclk));
	jxor g0311(.dina(w_n625_0[2]),.dinb(w_n623_0[2]),.dout(n626),.clk(gclk));
	jand g0312(.dina(w_n626_0[1]),.dinb(w_n622_1[1]),.dout(n627),.clk(gclk));
	jnot g0313(.din(w_G2256_1[1]),.dout(n628),.clk(gclk));
	jor g0314(.dina(w_dff_B_kkY0ITpc8_0),.dinb(w_n355_19[1]),.dout(n629),.clk(gclk));
	jand g0315(.dina(w_n629_0[1]),.dinb(w_n565_9[1]),.dout(n630),.clk(gclk));
	jxor g0316(.dina(w_n630_0[2]),.dinb(w_n628_0[1]),.dout(n631),.clk(gclk));
	jnot g0317(.din(w_G2253_1[1]),.dout(n632),.clk(gclk));
	jor g0318(.dina(w_dff_B_IaCFlZPL7_0),.dinb(w_n355_19[0]),.dout(n633),.clk(gclk));
	jand g0319(.dina(w_n633_0[1]),.dinb(w_n565_9[0]),.dout(n634),.clk(gclk));
	jxor g0320(.dina(w_n634_0[2]),.dinb(w_n632_0[1]),.dout(n635),.clk(gclk));
	jand g0321(.dina(w_n635_0[2]),.dinb(w_n631_0[1]),.dout(n636),.clk(gclk));
	jand g0322(.dina(n636),.dinb(w_n627_0[1]),.dout(n637),.clk(gclk));
	jnot g0323(.din(w_n637_0[1]),.dout(n638),.clk(gclk));
	jor g0324(.dina(w_dff_B_091w0Pok9_0),.dinb(w_n618_0[2]),.dout(n639),.clk(gclk));
	jand g0325(.dina(w_n630_0[1]),.dinb(w_n628_0[0]),.dout(n640),.clk(gclk));
	jnot g0326(.din(n640),.dout(n641),.clk(gclk));
	jand g0327(.dina(w_n634_0[1]),.dinb(w_n632_0[0]),.dout(n642),.clk(gclk));
	jnot g0328(.din(w_n642_0[1]),.dout(n643),.clk(gclk));
	jand g0329(.dina(w_n621_0[1]),.dinb(w_n619_0[0]),.dout(n644),.clk(gclk));
	jand g0330(.dina(w_n625_0[1]),.dinb(w_n623_0[1]),.dout(n645),.clk(gclk));
	jand g0331(.dina(w_n645_0[2]),.dinb(w_n622_1[0]),.dout(n646),.clk(gclk));
	jor g0332(.dina(n646),.dinb(w_dff_B_S3vLjFV19_1),.dout(n647),.clk(gclk));
	jnot g0333(.din(w_n647_0[1]),.dout(n648),.clk(gclk));
	jand g0334(.dina(w_n648_0[2]),.dinb(w_n643_0[1]),.dout(n649),.clk(gclk));
	jnot g0335(.din(w_n630_0[0]),.dout(n650),.clk(gclk));
	jand g0336(.dina(w_n650_0[1]),.dinb(w_G2256_1[0]),.dout(n651),.clk(gclk));
	jnot g0337(.din(w_n634_0[0]),.dout(n652),.clk(gclk));
	jand g0338(.dina(w_n652_0[1]),.dinb(w_G2253_1[0]),.dout(n653),.clk(gclk));
	jor g0339(.dina(w_n653_1[1]),.dinb(n651),.dout(n654),.clk(gclk));
	jor g0340(.dina(w_dff_B_ckRGBXmw0_0),.dinb(w_n649_0[1]),.dout(n655),.clk(gclk));
	jand g0341(.dina(n655),.dinb(w_dff_B_tDOpbQM73_1),.dout(n656),.clk(gclk));
	jand g0342(.dina(w_n656_0[1]),.dinb(n639),.dout(n657),.clk(gclk));
	jnot g0343(.din(w_G1486_0[2]),.dout(n658),.clk(gclk));
	jor g0344(.dina(w_dff_B_Fp6gxk5S3_0),.dinb(w_n355_18[2]),.dout(n659),.clk(gclk));
	jand g0345(.dina(w_n659_0[1]),.dinb(w_n565_8[2]),.dout(n660),.clk(gclk));
	jxor g0346(.dina(w_n660_1[1]),.dinb(w_n658_0[2]),.dout(n661),.clk(gclk));
	jnot g0347(.din(w_G1480_0[2]),.dout(n662),.clk(gclk));
	jor g0348(.dina(w_dff_B_5Zv08cyB5_0),.dinb(w_n355_18[1]),.dout(n663),.clk(gclk));
	jand g0349(.dina(w_n663_0[1]),.dinb(w_n565_8[1]),.dout(n664),.clk(gclk));
	jxor g0350(.dina(w_n664_1[1]),.dinb(w_n662_0[2]),.dout(n665),.clk(gclk));
	jnot g0351(.din(w_G106_1[1]),.dout(n666),.clk(gclk));
	jor g0352(.dina(w_dff_B_e0zlQvZn0_0),.dinb(w_n355_18[0]),.dout(n667),.clk(gclk));
	jand g0353(.dina(w_n667_0[1]),.dinb(w_n565_8[0]),.dout(n668),.clk(gclk));
	jxor g0354(.dina(w_n668_0[2]),.dinb(w_n666_0[1]),.dout(n669),.clk(gclk));
	jand g0355(.dina(w_n669_0[2]),.dinb(w_n665_0[2]),.dout(n670),.clk(gclk));
	jnot g0356(.din(w_G1469_1[1]),.dout(n671),.clk(gclk));
	jor g0357(.dina(w_dff_B_weg95XQN7_0),.dinb(w_n355_17[2]),.dout(n672),.clk(gclk));
	jand g0358(.dina(w_n672_0[1]),.dinb(w_n565_7[2]),.dout(n673),.clk(gclk));
	jxor g0359(.dina(w_n673_0[2]),.dinb(w_n671_0[1]),.dout(n674),.clk(gclk));
	jnot g0360(.din(w_G1462_0[2]),.dout(n675),.clk(gclk));
	jor g0361(.dina(w_dff_B_udsJNlPp0_0),.dinb(w_n355_17[1]),.dout(n676),.clk(gclk));
	jand g0362(.dina(w_n676_0[1]),.dinb(w_n565_7[1]),.dout(n677),.clk(gclk));
	jxor g0363(.dina(w_n677_0[2]),.dinb(w_n675_0[2]),.dout(n678),.clk(gclk));
	jand g0364(.dina(w_n678_0[2]),.dinb(w_n674_1[1]),.dout(n679),.clk(gclk));
	jand g0365(.dina(w_n679_1[1]),.dinb(n670),.dout(n680),.clk(gclk));
	jand g0366(.dina(w_n680_0[1]),.dinb(w_n661_0[1]),.dout(n681),.clk(gclk));
	jnot g0367(.din(n681),.dout(n682),.clk(gclk));
	jor g0368(.dina(w_dff_B_feVGc99K0_0),.dinb(w_n657_1[1]),.dout(n683),.clk(gclk));
	jand g0369(.dina(w_n660_1[0]),.dinb(w_n658_0[1]),.dout(n684),.clk(gclk));
	jor g0370(.dina(w_n660_0[2]),.dinb(w_n658_0[0]),.dout(n685),.clk(gclk));
	jand g0371(.dina(w_n664_1[0]),.dinb(w_n662_0[1]),.dout(n686),.clk(gclk));
	jnot g0372(.din(w_n686_0[1]),.dout(n687),.clk(gclk));
	jor g0373(.dina(w_n664_0[2]),.dinb(w_n662_0[0]),.dout(n688),.clk(gclk));
	jand g0374(.dina(w_n668_0[1]),.dinb(w_n666_0[0]),.dout(n689),.clk(gclk));
	jnot g0375(.din(w_n668_0[0]),.dout(n690),.clk(gclk));
	jand g0376(.dina(w_n690_0[1]),.dinb(w_G106_1[0]),.dout(n691),.clk(gclk));
	jnot g0377(.din(n691),.dout(n692),.clk(gclk));
	jnot g0378(.din(w_n673_0[1]),.dout(n693),.clk(gclk));
	jand g0379(.dina(w_n693_0[1]),.dinb(w_G1469_1[0]),.dout(n694),.clk(gclk));
	jnot g0380(.din(n694),.dout(n695),.clk(gclk));
	jand g0381(.dina(w_n673_0[0]),.dinb(w_n671_0[0]),.dout(n696),.clk(gclk));
	jand g0382(.dina(w_n677_0[1]),.dinb(w_n675_0[1]),.dout(n697),.clk(gclk));
	jor g0383(.dina(w_n697_0[2]),.dinb(n696),.dout(n698),.clk(gclk));
	jand g0384(.dina(w_dff_B_YznDGJU62_0),.dinb(n695),.dout(n699),.clk(gclk));
	jand g0385(.dina(w_n699_1[1]),.dinb(w_n692_0[1]),.dout(n700),.clk(gclk));
	jor g0386(.dina(n700),.dinb(w_dff_B_Qe26gSrG6_1),.dout(n701),.clk(gclk));
	jand g0387(.dina(w_n701_1[1]),.dinb(w_dff_B_X0nIvMJv5_1),.dout(n702),.clk(gclk));
	jnot g0388(.din(n702),.dout(n703),.clk(gclk));
	jand g0389(.dina(w_n703_0[1]),.dinb(w_n687_0[1]),.dout(n704),.clk(gclk));
	jnot g0390(.din(w_n704_0[1]),.dout(n705),.clk(gclk));
	jand g0391(.dina(w_n705_0[1]),.dinb(w_dff_B_SvFmXFXy0_1),.dout(n706),.clk(gclk));
	jor g0392(.dina(n706),.dinb(w_dff_B_1PVp4q1H5_1),.dout(n707),.clk(gclk));
	jnot g0393(.din(w_n707_0[2]),.dout(n708),.clk(gclk));
	jand g0394(.dina(w_n708_0[1]),.dinb(w_n683_0[1]),.dout(n709),.clk(gclk));
	jnot g0395(.din(w_G38_1[1]),.dout(n710),.clk(gclk));
	jand g0396(.dina(w_G4528_0[1]),.dinb(w_G1492_1[1]),.dout(n711),.clk(gclk));
	jxor g0397(.dina(w_n711_0[1]),.dinb(w_n710_0[1]),.dout(n712),.clk(gclk));
	jnot g0398(.din(w_n712_0[1]),.dout(n713),.clk(gclk));
	jor g0399(.dina(w_n713_1[1]),.dinb(w_n709_1[1]),.dout(n714),.clk(gclk));
	jor g0400(.dina(w_n714_0[1]),.dinb(w_n365_0[1]),.dout(n715),.clk(gclk));
	jnot g0401(.din(w_n715_0[2]),.dout(n716),.clk(gclk));
	jnot g0402(.din(w_G1492_1[0]),.dout(n717),.clk(gclk));
	jnot g0403(.din(w_n364_0[0]),.dout(n718),.clk(gclk));
	jor g0404(.dina(n718),.dinb(w_dff_B_x019fOFD0_1),.dout(n719),.clk(gclk));
	jand g0405(.dina(n719),.dinb(w_G38_1[0]),.dout(n720),.clk(gclk));
	jor g0406(.dina(w_n720_1[1]),.dinb(w_n716_1[1]),.dout(w_dff_A_JtpzOXIh8_2),.clk(gclk));
	jor g0407(.dina(w_dff_B_S4p4rGHS7_0),.dinb(w_n355_17[0]),.dout(n722),.clk(gclk));
	jand g0408(.dina(n722),.dinb(w_n565_7[0]),.dout(n723),.clk(gclk));
	jand g0409(.dina(w_G2236_0[2]),.dinb(w_G18_48[2]),.dout(n724),.clk(gclk));
	jnot g0410(.din(n724),.dout(n725),.clk(gclk));
	jor g0411(.dina(G64),.dinb(w_G18_48[1]),.dout(n726),.clk(gclk));
	jand g0412(.dina(w_dff_B_k7AAB8Kr6_0),.dinb(n725),.dout(n727),.clk(gclk));
	jor g0413(.dina(w_n727_0[2]),.dinb(w_n723_0[2]),.dout(n728),.clk(gclk));
	jand g0414(.dina(G178),.dinb(w_G18_48[0]),.dout(n729),.clk(gclk));
	jor g0415(.dina(w_dff_B_pSeVm3Mk5_0),.dinb(w_n581_0[0]),.dout(n730),.clk(gclk));
	jand g0416(.dina(w_G2230_0[2]),.dinb(w_G18_47[2]),.dout(n731),.clk(gclk));
	jnot g0417(.din(n731),.dout(n732),.clk(gclk));
	jor g0418(.dina(G85),.dinb(w_G18_47[1]),.dout(n733),.clk(gclk));
	jand g0419(.dina(w_dff_B_5Z0ZvisL2_0),.dinb(n732),.dout(n734),.clk(gclk));
	jor g0420(.dina(w_n734_0[2]),.dinb(w_n730_0[2]),.dout(n735),.clk(gclk));
	jand g0421(.dina(G179),.dinb(w_G18_47[0]),.dout(n736),.clk(gclk));
	jor g0422(.dina(w_dff_B_ymWx1Ohc5_0),.dinb(w_n586_0[0]),.dout(n737),.clk(gclk));
	jand g0423(.dina(w_G2224_0[2]),.dinb(w_G18_46[2]),.dout(n738),.clk(gclk));
	jnot g0424(.din(n738),.dout(n739),.clk(gclk));
	jor g0425(.dina(G84),.dinb(w_G18_46[1]),.dout(n740),.clk(gclk));
	jand g0426(.dina(w_dff_B_tHgUzJFw0_0),.dinb(n739),.dout(n741),.clk(gclk));
	jand g0427(.dina(w_n741_0[2]),.dinb(w_n737_0[2]),.dout(n742),.clk(gclk));
	jand g0428(.dina(G180),.dinb(w_G18_46[0]),.dout(n743),.clk(gclk));
	jor g0429(.dina(w_dff_B_QPrMLEMA6_0),.dinb(w_n570_0[0]),.dout(n744),.clk(gclk));
	jand g0430(.dina(w_G2218_0[1]),.dinb(w_G18_45[2]),.dout(n745),.clk(gclk));
	jnot g0431(.din(n745),.dout(n746),.clk(gclk));
	jor g0432(.dina(G83),.dinb(w_G18_45[1]),.dout(n747),.clk(gclk));
	jand g0433(.dina(w_dff_B_ImjzZV4d2_0),.dinb(n746),.dout(n748),.clk(gclk));
	jor g0434(.dina(w_n748_0[2]),.dinb(w_n744_0[2]),.dout(n749),.clk(gclk));
	jor g0435(.dina(w_n741_0[1]),.dinb(w_n737_0[1]),.dout(n750),.clk(gclk));
	jand g0436(.dina(n750),.dinb(n749),.dout(n751),.clk(gclk));
	jand g0437(.dina(w_n748_0[1]),.dinb(w_n744_0[1]),.dout(n752),.clk(gclk));
	jand g0438(.dina(G171),.dinb(w_G18_45[0]),.dout(n753),.clk(gclk));
	jor g0439(.dina(w_dff_B_89KUHvEO0_0),.dinb(w_n575_0[0]),.dout(n754),.clk(gclk));
	jand g0440(.dina(w_G2211_0[1]),.dinb(w_G18_44[2]),.dout(n755),.clk(gclk));
	jnot g0441(.din(n755),.dout(n756),.clk(gclk));
	jor g0442(.dina(G65),.dinb(w_G18_44[1]),.dout(n757),.clk(gclk));
	jand g0443(.dina(w_dff_B_FCQlh5Dj1_0),.dinb(n756),.dout(n758),.clk(gclk));
	jand g0444(.dina(w_n758_0[2]),.dinb(w_n754_0[2]),.dout(n759),.clk(gclk));
	jor g0445(.dina(w_n759_0[1]),.dinb(w_n752_0[1]),.dout(n760),.clk(gclk));
	jand g0446(.dina(n760),.dinb(w_n751_0[1]),.dout(n761),.clk(gclk));
	jor g0447(.dina(n761),.dinb(w_n742_0[1]),.dout(n762),.clk(gclk));
	jand g0448(.dina(n762),.dinb(w_n735_0[1]),.dout(n763),.clk(gclk));
	jand g0449(.dina(w_n734_0[1]),.dinb(w_n730_0[1]),.dout(n764),.clk(gclk));
	jand g0450(.dina(w_n727_0[1]),.dinb(w_n723_0[1]),.dout(n765),.clk(gclk));
	jor g0451(.dina(w_n765_0[1]),.dinb(w_n764_0[1]),.dout(n766),.clk(gclk));
	jor g0452(.dina(w_dff_B_374cMAJc9_0),.dinb(n763),.dout(n767),.clk(gclk));
	jand g0453(.dina(n767),.dinb(w_n728_0[1]),.dout(n768),.clk(gclk));
	jnot g0454(.din(w_n752_0[0]),.dout(n769),.clk(gclk));
	jand g0455(.dina(n769),.dinb(w_n735_0[0]),.dout(n770),.clk(gclk));
	jnot g0456(.din(w_n742_0[0]),.dout(n771),.clk(gclk));
	jnot g0457(.din(w_n759_0[0]),.dout(n772),.clk(gclk));
	jand g0458(.dina(n772),.dinb(n771),.dout(n773),.clk(gclk));
	jand g0459(.dina(n773),.dinb(n770),.dout(n774),.clk(gclk));
	jnot g0460(.din(w_n765_0[0]),.dout(n775),.clk(gclk));
	jor g0461(.dina(w_n758_0[1]),.dinb(w_n754_0[1]),.dout(n776),.clk(gclk));
	jand g0462(.dina(w_dff_B_GYqy8mHM6_0),.dinb(n775),.dout(n777),.clk(gclk));
	jnot g0463(.din(w_n764_0[0]),.dout(n778),.clk(gclk));
	jand g0464(.dina(n778),.dinb(w_n728_0[0]),.dout(n779),.clk(gclk));
	jand g0465(.dina(n779),.dinb(n777),.dout(n780),.clk(gclk));
	jand g0466(.dina(n780),.dinb(w_n751_0[0]),.dout(n781),.clk(gclk));
	jand g0467(.dina(n781),.dinb(w_dff_B_MDMrVRml4_1),.dout(n782),.clk(gclk));
	jand g0468(.dina(G191),.dinb(w_G18_44[0]),.dout(n783),.clk(gclk));
	jor g0469(.dina(w_dff_B_CXnBBQwP6_0),.dinb(w_n522_0[0]),.dout(n784),.clk(gclk));
	jor g0470(.dina(G60),.dinb(w_G18_43[2]),.dout(n785),.clk(gclk));
	jor g0471(.dina(w_n520_0[0]),.dinb(w_n355_16[2]),.dout(n786),.clk(gclk));
	jand g0472(.dina(n786),.dinb(w_dff_B_gMghVbHt7_1),.dout(n787),.clk(gclk));
	jxor g0473(.dina(w_n787_0[2]),.dinb(w_n784_0[2]),.dout(n788),.clk(gclk));
	jand g0474(.dina(G189),.dinb(w_G18_43[1]),.dout(n789),.clk(gclk));
	jor g0475(.dina(w_dff_B_PST0blmv8_0),.dinb(w_n533_0[0]),.dout(n790),.clk(gclk));
	jor g0476(.dina(G62),.dinb(w_G18_43[0]),.dout(n791),.clk(gclk));
	jor g0477(.dina(w_n531_0[0]),.dinb(w_n355_16[1]),.dout(n792),.clk(gclk));
	jand g0478(.dina(n792),.dinb(w_dff_B_iKVVTLIe3_1),.dout(n793),.clk(gclk));
	jxor g0479(.dina(w_n793_1[1]),.dinb(w_n790_1[1]),.dout(n794),.clk(gclk));
	jand g0480(.dina(n794),.dinb(n788),.dout(n795),.clk(gclk));
	jand g0481(.dina(G190),.dinb(w_G18_42[2]),.dout(n796),.clk(gclk));
	jor g0482(.dina(w_dff_B_54cKlWns1_0),.dinb(w_n538_0[0]),.dout(n797),.clk(gclk));
	jor g0483(.dina(G61),.dinb(w_G18_42[1]),.dout(n798),.clk(gclk));
	jand g0484(.dina(w_G4432_0[2]),.dinb(w_G18_42[0]),.dout(n799),.clk(gclk));
	jnot g0485(.din(n799),.dout(n800),.clk(gclk));
	jand g0486(.dina(n800),.dinb(w_dff_B_9UIE7en39_1),.dout(n801),.clk(gclk));
	jxor g0487(.dina(w_n801_1[1]),.dinb(w_n797_1[1]),.dout(n802),.clk(gclk));
	jand g0488(.dina(G192),.dinb(w_G18_41[2]),.dout(n803),.clk(gclk));
	jor g0489(.dina(w_dff_B_0CT38OSx1_0),.dinb(w_n527_0[0]),.dout(n804),.clk(gclk));
	jor g0490(.dina(G79),.dinb(w_G18_41[1]),.dout(n805),.clk(gclk));
	jor g0491(.dina(w_n525_0[0]),.dinb(w_n355_16[0]),.dout(n806),.clk(gclk));
	jand g0492(.dina(n806),.dinb(w_dff_B_6iLd3lGi5_1),.dout(n807),.clk(gclk));
	jxor g0493(.dina(w_n807_0[2]),.dinb(w_n804_0[2]),.dout(n808),.clk(gclk));
	jand g0494(.dina(n808),.dinb(w_n802_0[1]),.dout(n809),.clk(gclk));
	jand g0495(.dina(n809),.dinb(w_n795_0[1]),.dout(n810),.clk(gclk));
	jand g0496(.dina(G196),.dinb(w_G18_41[0]),.dout(n811),.clk(gclk));
	jor g0497(.dina(w_dff_B_HOoNpVCD2_0),.dinb(w_n473_0[0]),.dout(n812),.clk(gclk));
	jor g0498(.dina(G78),.dinb(w_G18_40[2]),.dout(n813),.clk(gclk));
	jand g0499(.dina(w_G4400_0[1]),.dinb(w_G18_40[1]),.dout(n814),.clk(gclk));
	jnot g0500(.din(n814),.dout(n815),.clk(gclk));
	jand g0501(.dina(n815),.dinb(w_dff_B_ME82u0P10_1),.dout(n816),.clk(gclk));
	jor g0502(.dina(w_n816_0[2]),.dinb(w_n812_0[2]),.dout(n817),.clk(gclk));
	jand g0503(.dina(G195),.dinb(w_G18_40[0]),.dout(n818),.clk(gclk));
	jor g0504(.dina(w_dff_B_XSsA1Wql7_0),.dinb(w_n488_0[0]),.dout(n819),.clk(gclk));
	jor g0505(.dina(G59),.dinb(w_G18_39[2]),.dout(n820),.clk(gclk));
	jand g0506(.dina(w_G4405_0[2]),.dinb(w_G18_39[1]),.dout(n821),.clk(gclk));
	jnot g0507(.din(n821),.dout(n822),.clk(gclk));
	jand g0508(.dina(n822),.dinb(w_dff_B_llGRv8mi5_1),.dout(n823),.clk(gclk));
	jor g0509(.dina(w_n823_0[2]),.dinb(w_n819_0[2]),.dout(n824),.clk(gclk));
	jand g0510(.dina(w_n824_0[1]),.dinb(w_n817_0[1]),.dout(n825),.clk(gclk));
	jand g0511(.dina(G187),.dinb(w_G18_39[0]),.dout(n826),.clk(gclk));
	jor g0512(.dina(w_dff_B_KyMlupGs9_0),.dinb(w_n477_0[0]),.dout(n827),.clk(gclk));
	jor g0513(.dina(G77),.dinb(w_G18_38[2]),.dout(n828),.clk(gclk));
	jand g0514(.dina(w_G4394_0[2]),.dinb(w_G18_38[1]),.dout(n829),.clk(gclk));
	jnot g0515(.din(n829),.dout(n830),.clk(gclk));
	jand g0516(.dina(n830),.dinb(w_dff_B_AUOibp789_1),.dout(n831),.clk(gclk));
	jand g0517(.dina(w_n831_0[2]),.dinb(w_n827_0[2]),.dout(n832),.clk(gclk));
	jnot g0518(.din(w_n832_0[1]),.dout(n833),.clk(gclk));
	jand g0519(.dina(w_n823_0[1]),.dinb(w_n819_0[1]),.dout(n834),.clk(gclk));
	jnot g0520(.din(w_n834_0[1]),.dout(n835),.clk(gclk));
	jand g0521(.dina(n835),.dinb(n833),.dout(n836),.clk(gclk));
	jand g0522(.dina(n836),.dinb(w_dff_B_C3rdXGV10_1),.dout(n837),.clk(gclk));
	jand g0523(.dina(w_n816_0[1]),.dinb(w_n812_0[1]),.dout(n838),.clk(gclk));
	jnot g0524(.din(w_n838_0[1]),.dout(n839),.clk(gclk));
	jor g0525(.dina(w_n831_0[1]),.dinb(w_n827_0[1]),.dout(n840),.clk(gclk));
	jand g0526(.dina(w_dff_B_2ir4DjU72_0),.dinb(n839),.dout(n841),.clk(gclk));
	jand g0527(.dina(G193),.dinb(w_G18_38[0]),.dout(n842),.clk(gclk));
	jor g0528(.dina(w_dff_B_VrqhbXKF4_0),.dinb(w_n468_0[0]),.dout(n843),.clk(gclk));
	jor g0529(.dina(G80),.dinb(w_G18_37[2]),.dout(n844),.clk(gclk));
	jand g0530(.dina(w_G4415_0[2]),.dinb(w_G18_37[1]),.dout(n845),.clk(gclk));
	jnot g0531(.din(n845),.dout(n846),.clk(gclk));
	jand g0532(.dina(n846),.dinb(w_dff_B_U64D73rS2_1),.dout(n847),.clk(gclk));
	jand g0533(.dina(w_n847_0[2]),.dinb(w_n843_0[2]),.dout(n848),.clk(gclk));
	jnot g0534(.din(w_n848_0[1]),.dout(n849),.clk(gclk));
	jand g0535(.dina(G194),.dinb(w_G18_37[0]),.dout(n850),.clk(gclk));
	jor g0536(.dina(w_dff_B_Wf7nYgeZ5_0),.dinb(w_n484_0[0]),.dout(n851),.clk(gclk));
	jor g0537(.dina(G81),.dinb(w_G18_36[2]),.dout(n852),.clk(gclk));
	jand g0538(.dina(w_G4410_0[2]),.dinb(w_G18_36[1]),.dout(n853),.clk(gclk));
	jnot g0539(.din(n853),.dout(n854),.clk(gclk));
	jand g0540(.dina(n854),.dinb(w_dff_B_8ePvQrtz7_1),.dout(n855),.clk(gclk));
	jor g0541(.dina(w_n855_0[2]),.dinb(w_n851_0[2]),.dout(n856),.clk(gclk));
	jand g0542(.dina(w_n856_0[1]),.dinb(n849),.dout(n857),.clk(gclk));
	jor g0543(.dina(w_n847_0[1]),.dinb(w_n843_0[1]),.dout(n858),.clk(gclk));
	jand g0544(.dina(w_n855_0[1]),.dinb(w_n851_0[1]),.dout(n859),.clk(gclk));
	jnot g0545(.din(w_n859_0[1]),.dout(n860),.clk(gclk));
	jand g0546(.dina(n860),.dinb(w_n858_0[2]),.dout(n861),.clk(gclk));
	jand g0547(.dina(n861),.dinb(n857),.dout(n862),.clk(gclk));
	jand g0548(.dina(n862),.dinb(w_dff_B_MLNtxgJY4_1),.dout(n863),.clk(gclk));
	jand g0549(.dina(n863),.dinb(w_dff_B_HHy6QElJ5_1),.dout(n864),.clk(gclk));
	jand g0550(.dina(w_n864_0[1]),.dinb(w_n810_0[2]),.dout(n865),.clk(gclk));
	jand g0551(.dina(G200),.dinb(w_G18_36[0]),.dout(n866),.clk(gclk));
	jnot g0552(.din(n866),.dout(n867),.clk(gclk));
	jand g0553(.dina(n867),.dinb(w_n441_0[0]),.dout(n868),.clk(gclk));
	jnot g0554(.din(n868),.dout(n869),.clk(gclk));
	jor g0555(.dina(G56),.dinb(w_G18_35[2]),.dout(n870),.clk(gclk));
	jand g0556(.dina(w_G3749_0[2]),.dinb(w_G18_35[1]),.dout(n871),.clk(gclk));
	jnot g0557(.din(n871),.dout(n872),.clk(gclk));
	jand g0558(.dina(n872),.dinb(w_dff_B_NDxgaqFP7_1),.dout(n873),.clk(gclk));
	jand g0559(.dina(w_n873_0[2]),.dinb(w_n869_0[2]),.dout(n874),.clk(gclk));
	jnot g0560(.din(w_n874_0[1]),.dout(n875),.clk(gclk));
	jnot g0561(.din(w_n427_0[0]),.dout(n876),.clk(gclk));
	jand g0562(.dina(G202),.dinb(w_G18_35[0]),.dout(n877),.clk(gclk));
	jor g0563(.dina(w_dff_B_DeWSW7nC9_0),.dinb(n876),.dout(n878),.clk(gclk));
	jor g0564(.dina(G54),.dinb(w_G18_34[2]),.dout(n879),.clk(gclk));
	jand g0565(.dina(w_G3737_0[2]),.dinb(w_G18_34[1]),.dout(n880),.clk(gclk));
	jnot g0566(.din(n880),.dout(n881),.clk(gclk));
	jand g0567(.dina(n881),.dinb(w_dff_B_O5SW7v0n6_1),.dout(n882),.clk(gclk));
	jor g0568(.dina(w_n882_0[2]),.dinb(w_n878_0[2]),.dout(n883),.clk(gclk));
	jand g0569(.dina(w_dff_B_CJYLLkVd5_0),.dinb(n875),.dout(n884),.clk(gclk));
	jand g0570(.dina(w_n882_0[1]),.dinb(w_n878_0[1]),.dout(n885),.clk(gclk));
	jnot g0571(.din(w_n885_0[1]),.dout(n886),.clk(gclk));
	jor g0572(.dina(w_n873_0[1]),.dinb(w_n869_0[1]),.dout(n887),.clk(gclk));
	jand g0573(.dina(w_n887_0[1]),.dinb(n886),.dout(n888),.clk(gclk));
	jand g0574(.dina(n888),.dinb(n884),.dout(n889),.clk(gclk));
	jand g0575(.dina(G201),.dinb(w_G18_34[0]),.dout(n890),.clk(gclk));
	jor g0576(.dina(w_dff_B_SoIl8LzQ8_0),.dinb(w_n448_0[0]),.dout(n891),.clk(gclk));
	jor g0577(.dina(G55),.dinb(w_G18_33[2]),.dout(n892),.clk(gclk));
	jand g0578(.dina(w_G3743_0[2]),.dinb(w_G18_33[1]),.dout(n893),.clk(gclk));
	jnot g0579(.din(n893),.dout(n894),.clk(gclk));
	jand g0580(.dina(n894),.dinb(w_dff_B_RvBlhviK6_1),.dout(n895),.clk(gclk));
	jxor g0581(.dina(w_n895_1[1]),.dinb(w_n891_1[1]),.dout(n896),.clk(gclk));
	jnot g0582(.din(w_n434_0[0]),.dout(n897),.clk(gclk));
	jand g0583(.dina(G203),.dinb(w_G18_33[0]),.dout(n898),.clk(gclk));
	jor g0584(.dina(w_dff_B_tmteiliS8_0),.dinb(n897),.dout(n899),.clk(gclk));
	jor g0585(.dina(G53),.dinb(w_G18_32[2]),.dout(n900),.clk(gclk));
	jor g0586(.dina(w_n430_0[0]),.dinb(w_n355_15[2]),.dout(n901),.clk(gclk));
	jand g0587(.dina(n901),.dinb(w_dff_B_v0d9Pcq65_1),.dout(n902),.clk(gclk));
	jxor g0588(.dina(w_n902_0[2]),.dinb(w_n899_0[2]),.dout(n903),.clk(gclk));
	jand g0589(.dina(n903),.dinb(w_n896_0[1]),.dout(n904),.clk(gclk));
	jand g0590(.dina(w_dff_B_Uh0Dhd3p5_0),.dinb(w_n889_0[1]),.dout(n905),.clk(gclk));
	jnot g0591(.din(w_n400_0[0]),.dout(n906),.clk(gclk));
	jand g0592(.dina(G207),.dinb(w_G18_32[1]),.dout(n907),.clk(gclk));
	jor g0593(.dina(w_dff_B_oaivzYWu2_0),.dinb(n906),.dout(n908),.clk(gclk));
	jor g0594(.dina(G74),.dinb(w_G18_32[0]),.dout(n909),.clk(gclk));
	jand g0595(.dina(w_G3705_1[2]),.dinb(w_G18_31[2]),.dout(n910),.clk(gclk));
	jnot g0596(.din(n910),.dout(n911),.clk(gclk));
	jand g0597(.dina(n911),.dinb(w_dff_B_NUpiunu24_1),.dout(n912),.clk(gclk));
	jor g0598(.dina(w_n912_0[2]),.dinb(w_n908_0[2]),.dout(n913),.clk(gclk));
	jnot g0599(.din(w_n376_0[0]),.dout(n914),.clk(gclk));
	jand g0600(.dina(G205),.dinb(w_G18_31[1]),.dout(n915),.clk(gclk));
	jor g0601(.dina(w_dff_B_l4rg2tHX6_0),.dinb(n914),.dout(n916),.clk(gclk));
	jor g0602(.dina(G75),.dinb(w_G18_31[0]),.dout(n917),.clk(gclk));
	jand g0603(.dina(w_G3717_1[2]),.dinb(w_G18_30[2]),.dout(n918),.clk(gclk));
	jnot g0604(.din(n918),.dout(n919),.clk(gclk));
	jand g0605(.dina(n919),.dinb(w_dff_B_fGFTF0XU1_1),.dout(n920),.clk(gclk));
	jor g0606(.dina(w_n920_0[2]),.dinb(w_n916_0[2]),.dout(n921),.clk(gclk));
	jand g0607(.dina(w_n921_0[1]),.dinb(w_n913_0[1]),.dout(n922),.clk(gclk));
	jand g0608(.dina(w_n920_0[1]),.dinb(w_n916_0[1]),.dout(n923),.clk(gclk));
	jnot g0609(.din(w_n923_0[1]),.dout(n924),.clk(gclk));
	jnot g0610(.din(w_n385_0[0]),.dout(n925),.clk(gclk));
	jand g0611(.dina(G206),.dinb(w_G18_30[1]),.dout(n926),.clk(gclk));
	jor g0612(.dina(w_dff_B_BrXuCZOI4_0),.dinb(n925),.dout(n927),.clk(gclk));
	jor g0613(.dina(G76),.dinb(w_G18_30[0]),.dout(n928),.clk(gclk));
	jand g0614(.dina(w_G3711_0[2]),.dinb(w_G18_29[2]),.dout(n929),.clk(gclk));
	jnot g0615(.din(n929),.dout(n930),.clk(gclk));
	jand g0616(.dina(n930),.dinb(w_dff_B_NrCPywIU0_1),.dout(n931),.clk(gclk));
	jor g0617(.dina(w_n931_0[2]),.dinb(w_n927_0[2]),.dout(n932),.clk(gclk));
	jand g0618(.dina(w_n932_0[1]),.dinb(n924),.dout(n933),.clk(gclk));
	jand g0619(.dina(n933),.dinb(w_dff_B_LEyrmZNw7_1),.dout(n934),.clk(gclk));
	jnot g0620(.din(w_G70_0[1]),.dout(n935),.clk(gclk));
	jand g0621(.dina(w_n935_0[1]),.dinb(w_n355_15[1]),.dout(n936),.clk(gclk));
	jnot g0622(.din(n936),.dout(n937),.clk(gclk));
	jor g0623(.dina(w_n937_0[1]),.dinb(w_G41_0[0]),.dout(n938),.clk(gclk));
	jand g0624(.dina(w_n937_0[0]),.dinb(w_n356_0[0]),.dout(n939),.clk(gclk));
	jnot g0625(.din(w_n939_0[1]),.dout(n940),.clk(gclk));
	jand g0626(.dina(n940),.dinb(w_dff_B_Yi2ITFyq1_1),.dout(n941),.clk(gclk));
	jand g0627(.dina(n941),.dinb(w_dff_B_lgvf0JUe6_1),.dout(n942),.clk(gclk));
	jnot g0628(.din(w_n370_0[0]),.dout(n943),.clk(gclk));
	jand g0629(.dina(G204),.dinb(w_G18_29[1]),.dout(n944),.clk(gclk));
	jor g0630(.dina(w_dff_B_KEa91tD61_0),.dinb(n943),.dout(n945),.clk(gclk));
	jor g0631(.dina(G73),.dinb(w_G18_29[0]),.dout(n946),.clk(gclk));
	jor g0632(.dina(w_n366_0[0]),.dinb(w_n355_15[0]),.dout(n947),.clk(gclk));
	jand g0633(.dina(n947),.dinb(w_dff_B_pi3wdSqF9_1),.dout(n948),.clk(gclk));
	jxor g0634(.dina(w_n948_1[1]),.dinb(w_n945_1[1]),.dout(n949),.clk(gclk));
	jand g0635(.dina(w_n912_0[1]),.dinb(w_n908_0[1]),.dout(n950),.clk(gclk));
	jnot g0636(.din(w_n950_0[1]),.dout(n951),.clk(gclk));
	jand g0637(.dina(w_n931_0[1]),.dinb(w_n927_0[1]),.dout(n952),.clk(gclk));
	jnot g0638(.din(w_n952_0[1]),.dout(n953),.clk(gclk));
	jand g0639(.dina(n953),.dinb(n951),.dout(n954),.clk(gclk));
	jand g0640(.dina(n954),.dinb(w_dff_B_Maxmj71J6_1),.dout(n955),.clk(gclk));
	jand g0641(.dina(n955),.dinb(w_dff_B_bSGiMxoB1_1),.dout(n956),.clk(gclk));
	jand g0642(.dina(n956),.dinb(w_dff_B_4d4R3abv3_1),.dout(n957),.clk(gclk));
	jand g0643(.dina(w_n957_0[1]),.dinb(w_n905_0[2]),.dout(n958),.clk(gclk));
	jand g0644(.dina(n958),.dinb(w_n865_0[1]),.dout(n959),.clk(gclk));
	jand g0645(.dina(w_n807_0[1]),.dinb(w_n804_0[1]),.dout(n960),.clk(gclk));
	jand g0646(.dina(n960),.dinb(w_n802_0[0]),.dout(n961),.clk(gclk));
	jand g0647(.dina(n961),.dinb(w_n795_0[0]),.dout(n962),.clk(gclk));
	jand g0648(.dina(w_n793_1[0]),.dinb(w_n790_1[0]),.dout(n963),.clk(gclk));
	jand g0649(.dina(w_n787_0[1]),.dinb(w_n784_0[1]),.dout(n964),.clk(gclk));
	jand g0650(.dina(w_n801_1[0]),.dinb(w_n797_1[0]),.dout(n965),.clk(gclk));
	jor g0651(.dina(n965),.dinb(n964),.dout(n966),.clk(gclk));
	jor g0652(.dina(w_n793_0[2]),.dinb(w_n790_0[2]),.dout(n967),.clk(gclk));
	jor g0653(.dina(w_n801_0[2]),.dinb(w_n797_0[2]),.dout(n968),.clk(gclk));
	jand g0654(.dina(n968),.dinb(n967),.dout(n969),.clk(gclk));
	jand g0655(.dina(n969),.dinb(n966),.dout(n970),.clk(gclk));
	jor g0656(.dina(n970),.dinb(w_dff_B_GRMGV4p45_1),.dout(n971),.clk(gclk));
	jor g0657(.dina(n971),.dinb(w_dff_B_Ub74zJxg8_1),.dout(n972),.clk(gclk));
	jand g0658(.dina(w_n832_0[0]),.dinb(w_n817_0[0]),.dout(n973),.clk(gclk));
	jor g0659(.dina(w_n838_0[0]),.dinb(w_n834_0[0]),.dout(n974),.clk(gclk));
	jor g0660(.dina(n974),.dinb(n973),.dout(n975),.clk(gclk));
	jand g0661(.dina(w_n858_0[1]),.dinb(w_n856_0[0]),.dout(n976),.clk(gclk));
	jand g0662(.dina(n976),.dinb(w_n824_0[0]),.dout(n977),.clk(gclk));
	jand g0663(.dina(n977),.dinb(n975),.dout(n978),.clk(gclk));
	jand g0664(.dina(w_n859_0[0]),.dinb(w_n858_0[0]),.dout(n979),.clk(gclk));
	jor g0665(.dina(n979),.dinb(w_n848_0[0]),.dout(n980),.clk(gclk));
	jor g0666(.dina(w_dff_B_pxRVTx135_0),.dinb(n978),.dout(n981),.clk(gclk));
	jand g0667(.dina(w_n981_0[1]),.dinb(w_n810_0[1]),.dout(n982),.clk(gclk));
	jor g0668(.dina(n982),.dinb(w_n972_0[1]),.dout(n983),.clk(gclk));
	jor g0669(.dina(w_dff_B_dJjfIWKK6_0),.dinb(n959),.dout(n984),.clk(gclk));
	jand g0670(.dina(n984),.dinb(w_n782_0[1]),.dout(n985),.clk(gclk));
	jor g0671(.dina(n985),.dinb(w_dff_B_9kGRiarq1_1),.dout(n986),.clk(gclk));
	jor g0672(.dina(w_dff_B_L2o6AYYH5_0),.dinb(w_n355_14[2]),.dout(n987),.clk(gclk));
	jand g0673(.dina(w_n987_0[1]),.dinb(w_n565_6[2]),.dout(n988),.clk(gclk));
	jand g0674(.dina(w_G2256_0[2]),.dinb(w_G18_28[2]),.dout(n989),.clk(gclk));
	jnot g0675(.din(n989),.dout(n990),.clk(gclk));
	jor g0676(.dina(G110),.dinb(w_G18_28[1]),.dout(n991),.clk(gclk));
	jand g0677(.dina(w_dff_B_k7lL40703_0),.dinb(n990),.dout(n992),.clk(gclk));
	jor g0678(.dina(w_n992_0[2]),.dinb(w_n988_0[2]),.dout(n993),.clk(gclk));
	jor g0679(.dina(w_dff_B_RzSElG5A5_0),.dinb(w_n355_14[1]),.dout(n994),.clk(gclk));
	jand g0680(.dina(w_n994_0[1]),.dinb(w_n565_6[1]),.dout(n995),.clk(gclk));
	jand g0681(.dina(w_G2247_0[1]),.dinb(w_G18_28[0]),.dout(n996),.clk(gclk));
	jnot g0682(.din(n996),.dout(n997),.clk(gclk));
	jor g0683(.dina(G86),.dinb(w_G18_27[2]),.dout(n998),.clk(gclk));
	jand g0684(.dina(w_dff_B_JiLRwsqs5_0),.dinb(n997),.dout(n999),.clk(gclk));
	jand g0685(.dina(w_n999_0[2]),.dinb(w_n995_0[2]),.dout(n1000),.clk(gclk));
	jnot g0686(.din(w_n1000_0[1]),.dout(n1001),.clk(gclk));
	jand g0687(.dina(n1001),.dinb(w_n993_0[1]),.dout(n1002),.clk(gclk));
	jand g0688(.dina(w_n992_0[1]),.dinb(w_n988_0[1]),.dout(n1003),.clk(gclk));
	jnot g0689(.din(w_n1003_0[1]),.dout(n1004),.clk(gclk));
	jor g0690(.dina(w_n999_0[1]),.dinb(w_n995_0[1]),.dout(n1005),.clk(gclk));
	jand g0691(.dina(w_dff_B_n58IivwY1_0),.dinb(n1004),.dout(n1006),.clk(gclk));
	jand g0692(.dina(n1006),.dinb(n1002),.dout(n1007),.clk(gclk));
	jor g0693(.dina(w_dff_B_YIasQm2p8_0),.dinb(w_n355_14[0]),.dout(n1008),.clk(gclk));
	jand g0694(.dina(w_n1008_0[1]),.dinb(w_n565_6[0]),.dout(n1009),.clk(gclk));
	jand g0695(.dina(w_G2253_0[2]),.dinb(w_G18_27[1]),.dout(n1010),.clk(gclk));
	jnot g0696(.din(n1010),.dout(n1011),.clk(gclk));
	jor g0697(.dina(G109),.dinb(w_G18_27[0]),.dout(n1012),.clk(gclk));
	jand g0698(.dina(w_dff_B_a2d6WJsL9_0),.dinb(n1011),.dout(n1013),.clk(gclk));
	jxor g0699(.dina(w_n1013_1[1]),.dinb(w_n1009_1[1]),.dout(n1014),.clk(gclk));
	jor g0700(.dina(w_dff_B_6oUft6vE8_0),.dinb(w_n355_13[2]),.dout(n1015),.clk(gclk));
	jand g0701(.dina(w_n1015_0[1]),.dinb(w_n565_5[2]),.dout(n1016),.clk(gclk));
	jor g0702(.dina(w_n623_0[0]),.dinb(w_n355_13[1]),.dout(n1017),.clk(gclk));
	jor g0703(.dina(G63),.dinb(w_G18_26[2]),.dout(n1018),.clk(gclk));
	jand g0704(.dina(w_dff_B_Dv298iPP6_0),.dinb(n1017),.dout(n1019),.clk(gclk));
	jxor g0705(.dina(w_n1019_0[2]),.dinb(w_n1016_0[2]),.dout(n1020),.clk(gclk));
	jand g0706(.dina(n1020),.dinb(w_n1014_0[1]),.dout(n1021),.clk(gclk));
	jand g0707(.dina(w_dff_B_AMOHr3Vf6_0),.dinb(w_n1007_0[1]),.dout(n1022),.clk(gclk));
	jand g0708(.dina(w_n1022_0[1]),.dinb(n986),.dout(n1023),.clk(gclk));
	jand g0709(.dina(w_n948_1[0]),.dinb(w_n945_1[0]),.dout(n1024),.clk(gclk));
	jor g0710(.dina(w_n950_0[0]),.dinb(w_n939_0[0]),.dout(n1025),.clk(gclk));
	jand g0711(.dina(w_n932_0[0]),.dinb(w_n913_0[0]),.dout(n1026),.clk(gclk));
	jand g0712(.dina(n1026),.dinb(n1025),.dout(n1027),.clk(gclk));
	jor g0713(.dina(w_n952_0[0]),.dinb(w_n923_0[0]),.dout(n1028),.clk(gclk));
	jor g0714(.dina(w_dff_B_P5WZjbkc1_0),.dinb(n1027),.dout(n1029),.clk(gclk));
	jor g0715(.dina(w_n948_0[2]),.dinb(w_n945_0[2]),.dout(n1030),.clk(gclk));
	jand g0716(.dina(n1030),.dinb(w_n921_0[0]),.dout(n1031),.clk(gclk));
	jand g0717(.dina(w_dff_B_CNs4IfNm6_0),.dinb(n1029),.dout(n1032),.clk(gclk));
	jor g0718(.dina(n1032),.dinb(w_dff_B_T7vY4eHE7_1),.dout(n1033),.clk(gclk));
	jand g0719(.dina(w_n1033_0[1]),.dinb(w_n905_0[1]),.dout(n1034),.clk(gclk));
	jand g0720(.dina(w_n902_0[1]),.dinb(w_n899_0[1]),.dout(n1035),.clk(gclk));
	jand g0721(.dina(n1035),.dinb(w_n896_0[0]),.dout(n1036),.clk(gclk));
	jand g0722(.dina(w_dff_B_0ybnmimc7_0),.dinb(w_n889_0[0]),.dout(n1037),.clk(gclk));
	jand g0723(.dina(w_n895_1[0]),.dinb(w_n891_1[0]),.dout(n1038),.clk(gclk));
	jor g0724(.dina(w_dff_B_w8MyrbaO0_0),.dinb(w_n885_0[0]),.dout(n1039),.clk(gclk));
	jor g0725(.dina(w_n895_0[2]),.dinb(w_n891_0[2]),.dout(n1040),.clk(gclk));
	jand g0726(.dina(w_dff_B_wtZEieFg8_0),.dinb(w_n887_0[0]),.dout(n1041),.clk(gclk));
	jand g0727(.dina(n1041),.dinb(n1039),.dout(n1042),.clk(gclk));
	jor g0728(.dina(n1042),.dinb(w_n874_0[0]),.dout(n1043),.clk(gclk));
	jor g0729(.dina(w_dff_B_N1uTPie67_0),.dinb(n1037),.dout(n1044),.clk(gclk));
	jor g0730(.dina(w_n1044_0[1]),.dinb(n1034),.dout(n1045),.clk(gclk));
	jand g0731(.dina(w_n1022_0[0]),.dinb(w_n782_0[0]),.dout(n1046),.clk(gclk));
	jand g0732(.dina(n1046),.dinb(w_n865_0[0]),.dout(n1047),.clk(gclk));
	jand g0733(.dina(w_dff_B_ApusimQ42_0),.dinb(n1045),.dout(n1048),.clk(gclk));
	jand g0734(.dina(w_n1019_0[1]),.dinb(w_n1016_0[1]),.dout(n1049),.clk(gclk));
	jand g0735(.dina(n1049),.dinb(w_n1014_0[0]),.dout(n1050),.clk(gclk));
	jand g0736(.dina(w_dff_B_vrsafaGC8_0),.dinb(w_n1007_0[0]),.dout(n1051),.clk(gclk));
	jand g0737(.dina(w_n1013_1[0]),.dinb(w_n1009_1[0]),.dout(n1052),.clk(gclk));
	jor g0738(.dina(n1052),.dinb(w_n1000_0[0]),.dout(n1053),.clk(gclk));
	jor g0739(.dina(w_n1013_0[2]),.dinb(w_n1009_0[2]),.dout(n1054),.clk(gclk));
	jand g0740(.dina(n1054),.dinb(w_n993_0[0]),.dout(n1055),.clk(gclk));
	jand g0741(.dina(n1055),.dinb(n1053),.dout(n1056),.clk(gclk));
	jor g0742(.dina(n1056),.dinb(w_n1003_0[0]),.dout(n1057),.clk(gclk));
	jor g0743(.dina(w_dff_B_ySOYDXTl2_0),.dinb(n1051),.dout(n1058),.clk(gclk));
	jor g0744(.dina(w_dff_B_wkkZXIpM0_0),.dinb(n1048),.dout(n1059),.clk(gclk));
	jor g0745(.dina(w_dff_B_gOANsO7i2_0),.dinb(n1023),.dout(n1060),.clk(gclk));
	jor g0746(.dina(w_dff_B_wyRCCiEu4_0),.dinb(w_n355_13[0]),.dout(n1061),.clk(gclk));
	jand g0747(.dina(w_n1061_0[2]),.dinb(w_n565_5[1]),.dout(n1062),.clk(gclk));
	jand g0748(.dina(w_G1480_0[1]),.dinb(w_G18_26[1]),.dout(n1063),.clk(gclk));
	jnot g0749(.din(n1063),.dout(n1064),.clk(gclk));
	jor g0750(.dina(G112),.dinb(w_G18_26[0]),.dout(n1065),.clk(gclk));
	jand g0751(.dina(w_dff_B_L7t6hzka9_0),.dinb(n1064),.dout(n1066),.clk(gclk));
	jor g0752(.dina(w_n1066_0[2]),.dinb(w_n1062_0[1]),.dout(n1067),.clk(gclk));
	jor g0753(.dina(w_dff_B_BBcmIffi9_0),.dinb(w_n355_12[2]),.dout(n1068),.clk(gclk));
	jand g0754(.dina(w_n1068_0[1]),.dinb(w_n565_5[0]),.dout(n1069),.clk(gclk));
	jand g0755(.dina(w_G1486_0[1]),.dinb(w_G18_25[2]),.dout(n1070),.clk(gclk));
	jnot g0756(.din(n1070),.dout(n1071),.clk(gclk));
	jor g0757(.dina(G88),.dinb(w_G18_25[1]),.dout(n1072),.clk(gclk));
	jand g0758(.dina(w_dff_B_0yBXJo9z0_0),.dinb(n1071),.dout(n1073),.clk(gclk));
	jor g0759(.dina(w_n1073_0[2]),.dinb(w_n1069_0[1]),.dout(n1074),.clk(gclk));
	jand g0760(.dina(n1074),.dinb(n1067),.dout(n1075),.clk(gclk));
	jor g0761(.dina(w_dff_B_go3tZ8237_0),.dinb(w_n355_12[1]),.dout(n1076),.clk(gclk));
	jand g0762(.dina(w_n1076_0[1]),.dinb(w_n565_4[2]),.dout(n1077),.clk(gclk));
	jand g0763(.dina(w_G1469_0[2]),.dinb(w_G18_25[0]),.dout(n1078),.clk(gclk));
	jnot g0764(.din(n1078),.dout(n1079),.clk(gclk));
	jor g0765(.dina(G111),.dinb(w_G18_24[2]),.dout(n1080),.clk(gclk));
	jand g0766(.dina(w_dff_B_eTd8rISp4_0),.dinb(n1079),.dout(n1081),.clk(gclk));
	jor g0767(.dina(w_n1081_0[2]),.dinb(w_n1077_0[2]),.dout(n1082),.clk(gclk));
	jand g0768(.dina(w_G1462_0[1]),.dinb(w_G18_24[1]),.dout(n1083),.clk(gclk));
	jnot g0769(.din(n1083),.dout(n1084),.clk(gclk));
	jor g0770(.dina(G113),.dinb(w_G18_24[0]),.dout(n1085),.clk(gclk));
	jand g0771(.dina(w_dff_B_ji1kzFuV4_0),.dinb(n1084),.dout(n1086),.clk(gclk));
	jor g0772(.dina(w_n1086_0[2]),.dinb(w_n565_4[1]),.dout(n1087),.clk(gclk));
	jand g0773(.dina(n1087),.dinb(w_n1082_0[1]),.dout(n1088),.clk(gclk));
	jand g0774(.dina(n1088),.dinb(w_n1075_0[1]),.dout(n1089),.clk(gclk));
	jand g0775(.dina(w_n1081_0[1]),.dinb(w_n1077_0[1]),.dout(n1090),.clk(gclk));
	jand g0776(.dina(w_n1086_0[1]),.dinb(w_n565_4[0]),.dout(n1091),.clk(gclk));
	jor g0777(.dina(n1091),.dinb(n1090),.dout(n1092),.clk(gclk));
	jnot g0778(.din(w_n1092_0[1]),.dout(n1093),.clk(gclk));
	jand g0779(.dina(w_n1066_0[1]),.dinb(w_n1062_0[0]),.dout(n1094),.clk(gclk));
	jor g0780(.dina(w_dff_B_P7acJj6O5_0),.dinb(w_n355_12[0]),.dout(n1095),.clk(gclk));
	jand g0781(.dina(w_n1095_0[1]),.dinb(w_n565_3[2]),.dout(n1096),.clk(gclk));
	jand g0782(.dina(w_G106_0[2]),.dinb(w_G18_23[2]),.dout(n1097),.clk(gclk));
	jnot g0783(.din(n1097),.dout(n1098),.clk(gclk));
	jor g0784(.dina(G87),.dinb(w_G18_23[1]),.dout(n1099),.clk(gclk));
	jand g0785(.dina(w_dff_B_rcYx8yKf4_0),.dinb(n1098),.dout(n1100),.clk(gclk));
	jand g0786(.dina(w_n1100_0[2]),.dinb(w_n1096_0[2]),.dout(n1101),.clk(gclk));
	jor g0787(.dina(n1101),.dinb(n1094),.dout(n1102),.clk(gclk));
	jnot g0788(.din(w_n1102_0[1]),.dout(n1103),.clk(gclk));
	jor g0789(.dina(w_n1100_0[1]),.dinb(w_n1096_0[1]),.dout(n1104),.clk(gclk));
	jand g0790(.dina(w_n1073_0[1]),.dinb(w_n1069_0[0]),.dout(n1105),.clk(gclk));
	jnot g0791(.din(w_n1105_0[1]),.dout(n1106),.clk(gclk));
	jand g0792(.dina(n1106),.dinb(w_n1104_0[1]),.dout(n1107),.clk(gclk));
	jand g0793(.dina(n1107),.dinb(n1103),.dout(n1108),.clk(gclk));
	jand g0794(.dina(n1108),.dinb(w_dff_B_V9LgDelO6_1),.dout(n1109),.clk(gclk));
	jand g0795(.dina(n1109),.dinb(w_dff_B_PhMNAOfy1_1),.dout(n1110),.clk(gclk));
	jand g0796(.dina(w_dff_B_w1tGP8yo3_0),.dinb(n1060),.dout(n1111),.clk(gclk));
	jand g0797(.dina(w_n1104_0[0]),.dinb(w_n1082_0[0]),.dout(n1112),.clk(gclk));
	jand g0798(.dina(n1112),.dinb(w_n1092_0[0]),.dout(n1113),.clk(gclk));
	jor g0799(.dina(n1113),.dinb(w_n1102_0[0]),.dout(n1114),.clk(gclk));
	jand g0800(.dina(n1114),.dinb(w_n1075_0[0]),.dout(n1115),.clk(gclk));
	jnot g0801(.din(w_G4528_0[0]),.dout(n1116),.clk(gclk));
	jor g0802(.dina(w_G2204_0[2]),.dinb(w_G1455_0[2]),.dout(n1117),.clk(gclk));
	jor g0803(.dina(n1117),.dinb(w_n1116_0[1]),.dout(n1118),.clk(gclk));
	jand g0804(.dina(n1118),.dinb(w_G38_0[2]),.dout(n1119),.clk(gclk));
	jor g0805(.dina(w_dff_B_DZE264KT4_0),.dinb(w_n1105_0[0]),.dout(n1120),.clk(gclk));
	jor g0806(.dina(w_dff_B_C5muFh6p3_0),.dinb(n1115),.dout(n1121),.clk(gclk));
	jor g0807(.dina(w_dff_B_uEgPLN9I8_0),.dinb(n1111),.dout(n1122),.clk(gclk));
	jand g0808(.dina(w_G2204_0[1]),.dinb(w_G1455_0[1]),.dout(n1123),.clk(gclk));
	jor g0809(.dina(w_n1116_0[0]),.dinb(w_G38_0[1]),.dout(n1124),.clk(gclk));
	jor g0810(.dina(n1124),.dinb(w_dff_B_lqJRKDNW7_1),.dout(n1125),.clk(gclk));
	jand g0811(.dina(w_n1125_0[2]),.dinb(w_n1122_0[2]),.dout(w_dff_A_W0B7nnBb3_2),.clk(gclk));
	jand g0812(.dina(w_n377_1[0]),.dinb(w_G3717_1[1]),.dout(n1127),.clk(gclk));
	jand g0813(.dina(w_n413_1[0]),.dinb(w_n410_0[0]),.dout(n1128),.clk(gclk));
	jor g0814(.dina(w_n1128_1[1]),.dinb(w_n1127_0[1]),.dout(n1129),.clk(gclk));
	jand g0815(.dina(n1129),.dinb(w_n417_0[1]),.dout(n1130),.clk(gclk));
	jor g0816(.dina(w_n405_0[1]),.dinb(w_n379_1[0]),.dout(n1131),.clk(gclk));
	jand g0817(.dina(w_dff_B_wgDSXUDG2_0),.dinb(w_n1130_0[1]),.dout(n1132),.clk(gclk));
	jxor g0818(.dina(n1132),.dinb(w_n372_1[1]),.dout(w_dff_A_EFX9NOPw8_2),.clk(gclk));
	jand g0819(.dina(w_n1128_1[0]),.dinb(w_n405_0[0]),.dout(n1134),.clk(gclk));
	jxor g0820(.dina(n1134),.dinb(w_n379_0[2]),.dout(w_dff_A_xvoXLmi80_2),.clk(gclk));
	jand g0821(.dina(w_n408_0[0]),.dinb(w_n412_0[1]),.dout(n1136),.clk(gclk));
	jand g0822(.dina(w_n1136_0[1]),.dinb(w_n404_0[0]),.dout(n1137),.clk(gclk));
	jxor g0823(.dina(n1137),.dinb(w_n387_0[2]),.dout(w_dff_A_7MoqT9H23_2),.clk(gclk));
	jor g0824(.dina(w_n395_0[1]),.dinb(w_n388_0[1]),.dout(n1139),.clk(gclk));
	jand g0825(.dina(n1139),.dinb(w_n354_1[0]),.dout(n1140),.clk(gclk));
	jxor g0826(.dina(n1140),.dinb(w_n402_0[2]),.dout(w_dff_A_iAHGgVal8_2),.clk(gclk));
	jor g0827(.dina(w_n437_0[0]),.dinb(w_n422_1[1]),.dout(n1142),.clk(gclk));
	jor g0828(.dina(w_n1142_0[1]),.dinb(w_n456_0[1]),.dout(n1143),.clk(gclk));
	jand g0829(.dina(n1143),.dinb(w_n462_0[1]),.dout(n1144),.clk(gclk));
	jxor g0830(.dina(n1144),.dinb(w_n446_1[0]),.dout(w_dff_A_HM031umB3_2),.clk(gclk));
	jand g0831(.dina(w_n1142_0[0]),.dinb(w_n460_0[1]),.dout(n1146),.clk(gclk));
	jxor g0832(.dina(n1146),.dinb(w_n450_0[1]),.dout(w_dff_A_8OItUSdo4_2),.clk(gclk));
	jand g0833(.dina(w_n435_0[2]),.dinb(w_G3729_0[2]),.dout(n1148),.clk(gclk));
	jor g0834(.dina(w_n1148_0[2]),.dinb(w_n422_1[0]),.dout(n1149),.clk(gclk));
	jand g0835(.dina(n1149),.dinb(w_n458_0[1]),.dout(n1150),.clk(gclk));
	jxor g0836(.dina(n1150),.dinb(w_n429_1[2]),.dout(w_dff_A_inYkeue56_2),.clk(gclk));
	jxor g0837(.dina(w_n436_0[0]),.dinb(w_n422_0[2]),.dout(w_dff_A_YuMbcDwy0_2),.clk(gclk));
	jxor g0838(.dina(w_n583_0[1]),.dinb(w_n577_0[0]),.dout(n1153),.clk(gclk));
	jxor g0839(.dina(w_n588_0[1]),.dinb(w_n567_0[1]),.dout(n1154),.clk(gclk));
	jxor g0840(.dina(n1154),.dinb(w_n572_0[2]),.dout(n1155),.clk(gclk));
	jnot g0841(.din(w_n625_0[0]),.dout(n1156),.clk(gclk));
	jor g0842(.dina(w_n1156_0[1]),.dinb(w_n620_0[0]),.dout(n1157),.clk(gclk));
	jnot g0843(.din(w_n621_0[0]),.dout(n1158),.clk(gclk));
	jor g0844(.dina(w_n624_0[0]),.dinb(n1158),.dout(n1159),.clk(gclk));
	jand g0845(.dina(n1159),.dinb(n1157),.dout(n1160),.clk(gclk));
	jor g0846(.dina(w_n652_0[0]),.dinb(w_n629_0[0]),.dout(n1161),.clk(gclk));
	jor g0847(.dina(w_n633_0[0]),.dinb(w_n650_0[0]),.dout(n1162),.clk(gclk));
	jand g0848(.dina(n1162),.dinb(n1161),.dout(n1163),.clk(gclk));
	jxor g0849(.dina(n1163),.dinb(n1160),.dout(n1164),.clk(gclk));
	jnot g0850(.din(G141),.dout(n1165),.clk(gclk));
	jor g0851(.dina(n1165),.dinb(w_G18_23[0]),.dout(n1166),.clk(gclk));
	jnot g0852(.din(G161),.dout(n1167),.clk(gclk));
	jor g0853(.dina(n1167),.dinb(w_n355_11[2]),.dout(n1168),.clk(gclk));
	jand g0854(.dina(n1168),.dinb(w_n1166_0[1]),.dout(n1169),.clk(gclk));
	jxor g0855(.dina(w_dff_B_9Wcolvdi7_0),.dinb(n1164),.dout(n1170),.clk(gclk));
	jxor g0856(.dina(n1170),.dinb(w_dff_B_vpv4Ip8T8_1),.dout(n1171),.clk(gclk));
	jxor g0857(.dina(n1171),.dinb(w_dff_B_S0kEqjWA1_1),.dout(n1172),.clk(gclk));
	jand g0858(.dina(w_n565_3[1]),.dinb(w_G18_22[2]),.dout(n1173),.clk(gclk));
	jxor g0859(.dina(G212),.dinb(G211),.dout(n1174),.clk(gclk));
	jand g0860(.dina(w_dff_B_DMTwZLiq9_0),.dinb(w_n1173_0[1]),.dout(n1175),.clk(gclk));
	jor g0861(.dina(w_n676_0[0]),.dinb(w_n564_0[1]),.dout(n1176),.clk(gclk));
	jnot g0862(.din(w_n659_0[0]),.dout(n1177),.clk(gclk));
	jand g0863(.dina(w_n664_0[1]),.dinb(n1177),.dout(n1178),.clk(gclk));
	jnot g0864(.din(w_n663_0[0]),.dout(n1179),.clk(gclk));
	jand g0865(.dina(n1179),.dinb(w_n660_0[1]),.dout(n1180),.clk(gclk));
	jor g0866(.dina(n1180),.dinb(n1178),.dout(n1181),.clk(gclk));
	jor g0867(.dina(w_n693_0[0]),.dinb(w_n667_0[0]),.dout(n1182),.clk(gclk));
	jor g0868(.dina(w_n672_0[0]),.dinb(w_n690_0[0]),.dout(n1183),.clk(gclk));
	jand g0869(.dina(n1183),.dinb(n1182),.dout(n1184),.clk(gclk));
	jxor g0870(.dina(n1184),.dinb(w_dff_B_RLt04rw04_1),.dout(n1185),.clk(gclk));
	jxor g0871(.dina(n1185),.dinb(w_dff_B_1PUvQFvx8_1),.dout(n1186),.clk(gclk));
	jxor g0872(.dina(n1186),.dinb(w_dff_B_h5HuSvVj9_1),.dout(n1187),.clk(gclk));
	jand g0873(.dina(G239),.dinb(w_G18_22[1]),.dout(n1188),.clk(gclk));
	jand g0874(.dina(w_dff_B_3kyWkG664_0),.dinb(w_n355_11[1]),.dout(n1189),.clk(gclk));
	jor g0875(.dina(w_n1189_0[1]),.dinb(w_dff_B_3mrAU2E69_1),.dout(n1190),.clk(gclk));
	jxor g0876(.dina(w_n442_0[0]),.dinb(w_n428_0[0]),.dout(n1191),.clk(gclk));
	jxor g0877(.dina(w_n449_0[0]),.dinb(w_n435_0[1]),.dout(n1192),.clk(gclk));
	jxor g0878(.dina(n1192),.dinb(n1191),.dout(n1193),.clk(gclk));
	jxor g0879(.dina(n1193),.dinb(w_dff_B_3eoJBKu19_1),.dout(n1194),.clk(gclk));
	jxor g0880(.dina(w_n401_1[0]),.dinb(w_n371_0[1]),.dout(n1195),.clk(gclk));
	jxor g0881(.dina(n1195),.dinb(w_n377_0[2]),.dout(n1196),.clk(gclk));
	jxor g0882(.dina(w_n386_0[0]),.dinb(w_n358_0[0]),.dout(n1197),.clk(gclk));
	jxor g0883(.dina(w_dff_B_BBu6uxmD6_0),.dinb(n1196),.dout(n1198),.clk(gclk));
	jxor g0884(.dina(n1198),.dinb(n1194),.dout(n1199),.clk(gclk));
	jxor g0885(.dina(w_n534_0[1]),.dinb(w_n523_0[0]),.dout(n1200),.clk(gclk));
	jxor g0886(.dina(w_n539_0[1]),.dinb(w_n528_0[2]),.dout(n1201),.clk(gclk));
	jxor g0887(.dina(n1201),.dinb(n1200),.dout(n1202),.clk(gclk));
	jxor g0888(.dina(n1202),.dinb(w_n503_0[0]),.dout(n1203),.clk(gclk));
	jand g0889(.dina(G227),.dinb(w_G18_22[0]),.dout(n1204),.clk(gclk));
	jand g0890(.dina(w_dff_B_PWdaVupe0_0),.dinb(w_n355_11[0]),.dout(n1205),.clk(gclk));
	jor g0891(.dina(w_n1205_0[1]),.dinb(w_dff_B_jid7V4CH7_1),.dout(n1206),.clk(gclk));
	jxor g0892(.dina(w_n489_0[0]),.dinb(w_n478_0[0]),.dout(n1207),.clk(gclk));
	jxor g0893(.dina(n1207),.dinb(w_dff_B_MqGAPJKl8_1),.dout(n1208),.clk(gclk));
	jxor g0894(.dina(w_n474_0[2]),.dinb(w_n469_0[1]),.dout(n1209),.clk(gclk));
	jxor g0895(.dina(w_dff_B_PXNiVJ5t5_0),.dinb(n1208),.dout(n1210),.clk(gclk));
	jxor g0896(.dina(n1210),.dinb(n1203),.dout(n1211),.clk(gclk));
	jor g0897(.dina(n1211),.dinb(n1199),.dout(n1212),.clk(gclk));
	jor g0898(.dina(w_dff_B_RWA6pG1u7_0),.dinb(n1187),.dout(n1213),.clk(gclk));
	jor g0899(.dina(n1213),.dinb(n1172),.dout(G412_fa_),.clk(gclk));
	jxor g0900(.dina(w_n831_0[0]),.dinb(w_n823_0[0]),.dout(n1215),.clk(gclk));
	jxor g0901(.dina(w_n847_0[0]),.dinb(w_n816_0[0]),.dout(n1216),.clk(gclk));
	jxor g0902(.dina(n1216),.dinb(w_n855_0[0]),.dout(n1217),.clk(gclk));
	jxor g0903(.dina(w_n793_0[1]),.dinb(w_n787_0[0]),.dout(n1218),.clk(gclk));
	jxor g0904(.dina(w_n807_0[0]),.dinb(w_n801_0[1]),.dout(n1219),.clk(gclk));
	jxor g0905(.dina(n1219),.dinb(n1218),.dout(n1220),.clk(gclk));
	jor g0906(.dina(w_G4393_0[1]),.dinb(w_n355_10[2]),.dout(n1221),.clk(gclk));
	jnot g0907(.din(G58),.dout(n1222),.clk(gclk));
	jor g0908(.dina(n1222),.dinb(w_G18_21[2]),.dout(n1223),.clk(gclk));
	jand g0909(.dina(n1223),.dinb(n1221),.dout(n1224),.clk(gclk));
	jxor g0910(.dina(w_dff_B_FXgMXwFy3_0),.dinb(n1220),.dout(n1225),.clk(gclk));
	jxor g0911(.dina(n1225),.dinb(w_dff_B_qk2e6yzr7_1),.dout(n1226),.clk(gclk));
	jxor g0912(.dina(n1226),.dinb(w_dff_B_5vCkOg337_1),.dout(n1227),.clk(gclk));
	jxor g0913(.dina(w_n389_0[0]),.dinb(w_G3698_0[1]),.dout(n1228),.clk(gclk));
	jor g0914(.dina(n1228),.dinb(w_n355_10[1]),.dout(n1229),.clk(gclk));
	jnot g0915(.din(w_G69_0[1]),.dout(n1230),.clk(gclk));
	jand g0916(.dina(w_n935_0[0]),.dinb(n1230),.dout(n1231),.clk(gclk));
	jand g0917(.dina(w_G70_0[0]),.dinb(w_G69_0[0]),.dout(n1232),.clk(gclk));
	jor g0918(.dina(n1232),.dinb(w_G18_21[1]),.dout(n1233),.clk(gclk));
	jor g0919(.dina(n1233),.dinb(n1231),.dout(n1234),.clk(gclk));
	jand g0920(.dina(n1234),.dinb(n1229),.dout(n1235),.clk(gclk));
	jxor g0921(.dina(n1235),.dinb(w_n912_0[0]),.dout(n1236),.clk(gclk));
	jnot g0922(.din(w_n1236_0[1]),.dout(n1237),.clk(gclk));
	jxor g0923(.dina(w_n948_0[1]),.dinb(w_n931_0[0]),.dout(n1238),.clk(gclk));
	jnot g0924(.din(w_n920_0[0]),.dout(n1239),.clk(gclk));
	jxor g0925(.dina(w_n882_0[0]),.dinb(w_n873_0[0]),.dout(n1240),.clk(gclk));
	jxor g0926(.dina(w_n902_0[0]),.dinb(w_n895_0[1]),.dout(n1241),.clk(gclk));
	jxor g0927(.dina(n1241),.dinb(n1240),.dout(n1242),.clk(gclk));
	jxor g0928(.dina(n1242),.dinb(w_dff_B_ovWBiHve8_1),.dout(n1243),.clk(gclk));
	jxor g0929(.dina(n1243),.dinb(w_dff_B_QHRDrX0e1_1),.dout(n1244),.clk(gclk));
	jnot g0930(.din(w_n1244_0[1]),.dout(n1245),.clk(gclk));
	jand g0931(.dina(n1245),.dinb(w_dff_B_1lI4iuCx7_1),.dout(n1246),.clk(gclk));
	jand g0932(.dina(w_n1244_0[0]),.dinb(w_n1236_0[0]),.dout(n1247),.clk(gclk));
	jor g0933(.dina(w_G1459_0[1]),.dinb(w_n355_10[0]),.dout(n1248),.clk(gclk));
	jnot g0934(.din(G114),.dout(n1249),.clk(gclk));
	jor g0935(.dina(n1249),.dinb(w_G18_21[0]),.dout(n1250),.clk(gclk));
	jand g0936(.dina(n1250),.dinb(n1248),.dout(n1251),.clk(gclk));
	jxor g0937(.dina(w_n1086_0[0]),.dinb(w_n1081_0[0]),.dout(n1252),.clk(gclk));
	jxor g0938(.dina(n1252),.dinb(w_dff_B_H2CRhkLX8_1),.dout(n1253),.clk(gclk));
	jxor g0939(.dina(w_n1100_0[0]),.dinb(w_n1073_0[0]),.dout(n1254),.clk(gclk));
	jxor g0940(.dina(n1254),.dinb(w_n1066_0[0]),.dout(n1255),.clk(gclk));
	jxor g0941(.dina(w_G1496_0[1]),.dinb(w_G1492_0[2]),.dout(n1256),.clk(gclk));
	jor g0942(.dina(n1256),.dinb(w_n355_9[2]),.dout(n1257),.clk(gclk));
	jxor g0943(.dina(w_G2204_0[0]),.dinb(w_G1455_0[0]),.dout(n1258),.clk(gclk));
	jor g0944(.dina(n1258),.dinb(w_G18_20[2]),.dout(n1259),.clk(gclk));
	jand g0945(.dina(n1259),.dinb(n1257),.dout(n1260),.clk(gclk));
	jxor g0946(.dina(w_dff_B_MZwE7jgl3_0),.dinb(n1255),.dout(n1261),.clk(gclk));
	jxor g0947(.dina(n1261),.dinb(w_dff_B_G3fOBOAh3_1),.dout(n1262),.clk(gclk));
	jxor g0948(.dina(w_n999_0[0]),.dinb(w_n992_0[0]),.dout(n1263),.clk(gclk));
	jxor g0949(.dina(w_n1019_0[0]),.dinb(w_n1013_0[1]),.dout(n1264),.clk(gclk));
	jxor g0950(.dina(n1264),.dinb(n1263),.dout(n1265),.clk(gclk));
	jxor g0951(.dina(n1265),.dinb(w_n727_0[0]),.dout(n1266),.clk(gclk));
	jor g0952(.dina(w_G2208_0[1]),.dinb(w_n355_9[1]),.dout(n1267),.clk(gclk));
	jnot g0953(.din(G82),.dout(n1268),.clk(gclk));
	jor g0954(.dina(n1268),.dinb(w_G18_20[1]),.dout(n1269),.clk(gclk));
	jand g0955(.dina(n1269),.dinb(n1267),.dout(n1270),.clk(gclk));
	jxor g0956(.dina(w_n758_0[0]),.dinb(w_n748_0[0]),.dout(n1271),.clk(gclk));
	jxor g0957(.dina(n1271),.dinb(w_dff_B_AtF61fDY2_1),.dout(n1272),.clk(gclk));
	jxor g0958(.dina(w_n741_0[0]),.dinb(w_n734_0[0]),.dout(n1273),.clk(gclk));
	jxor g0959(.dina(w_dff_B_eKyjidAx3_0),.dinb(n1272),.dout(n1274),.clk(gclk));
	jxor g0960(.dina(n1274),.dinb(n1266),.dout(n1275),.clk(gclk));
	jor g0961(.dina(n1275),.dinb(n1262),.dout(n1276),.clk(gclk));
	jor g0962(.dina(n1276),.dinb(n1247),.dout(n1277),.clk(gclk));
	jor g0963(.dina(n1277),.dinb(n1246),.dout(n1278),.clk(gclk));
	jor g0964(.dina(n1278),.dinb(w_dff_B_XgTx141R4_1),.dout(G414_fa_),.clk(gclk));
	jnot g0965(.din(w_n1061_0[1]),.dout(n1280),.clk(gclk));
	jnot g0966(.din(G170),.dout(n1281),.clk(gclk));
	jand g0967(.dina(n1281),.dinb(w_G18_20[0]),.dout(n1282),.clk(gclk));
	jxor g0968(.dina(n1282),.dinb(w_n1068_0[0]),.dout(n1283),.clk(gclk));
	jnot g0969(.din(w_n1283_0[1]),.dout(n1284),.clk(gclk));
	jand g0970(.dina(n1284),.dinb(w_dff_B_SaZRZ3eC7_1),.dout(n1285),.clk(gclk));
	jand g0971(.dina(w_n1283_0[0]),.dinb(w_n1061_0[0]),.dout(n1286),.clk(gclk));
	jor g0972(.dina(n1286),.dinb(w_n564_0[0]),.dout(n1287),.clk(gclk));
	jor g0973(.dina(n1287),.dinb(n1285),.dout(n1288),.clk(gclk));
	jnot g0974(.din(w_n1077_0[0]),.dout(n1289),.clk(gclk));
	jor g0975(.dina(w_n1095_0[0]),.dinb(n1289),.dout(n1290),.clk(gclk));
	jnot g0976(.din(w_n1096_0[0]),.dout(n1291),.clk(gclk));
	jor g0977(.dina(n1291),.dinb(w_n1076_0[0]),.dout(n1292),.clk(gclk));
	jand g0978(.dina(n1292),.dinb(n1290),.dout(n1293),.clk(gclk));
	jxor g0979(.dina(G165),.dinb(G164),.dout(n1294),.clk(gclk));
	jand g0980(.dina(w_dff_B_sSfu5jc82_0),.dinb(w_n1173_0[0]),.dout(n1295),.clk(gclk));
	jxor g0981(.dina(w_dff_B_EqwYgOAb4_0),.dinb(n1293),.dout(n1296),.clk(gclk));
	jxor g0982(.dina(n1296),.dinb(w_dff_B_q7BVBUQk7_1),.dout(n1297),.clk(gclk));
	jxor g0983(.dina(w_n790_0[1]),.dinb(w_n784_0[0]),.dout(n1298),.clk(gclk));
	jxor g0984(.dina(w_n804_0[0]),.dinb(w_n797_0[1]),.dout(n1299),.clk(gclk));
	jxor g0985(.dina(n1299),.dinb(n1298),.dout(n1300),.clk(gclk));
	jxor g0986(.dina(n1300),.dinb(w_n851_0[0]),.dout(n1301),.clk(gclk));
	jand g0987(.dina(G197),.dinb(w_G18_19[2]),.dout(n1302),.clk(gclk));
	jor g0988(.dina(w_dff_B_lOMOsdSt8_0),.dinb(w_n1205_0[0]),.dout(n1303),.clk(gclk));
	jnot g0989(.din(n1303),.dout(n1304),.clk(gclk));
	jxor g0990(.dina(w_n827_0[0]),.dinb(w_n819_0[0]),.dout(n1305),.clk(gclk));
	jxor g0991(.dina(n1305),.dinb(n1304),.dout(n1306),.clk(gclk));
	jnot g0992(.din(n1306),.dout(n1307),.clk(gclk));
	jxor g0993(.dina(w_n843_0[0]),.dinb(w_n812_0[0]),.dout(n1308),.clk(gclk));
	jxor g0994(.dina(w_dff_B_jPTP5tlu9_0),.dinb(n1307),.dout(n1309),.clk(gclk));
	jand g0995(.dina(w_n1309_0[1]),.dinb(w_n1301_0[1]),.dout(n1310),.clk(gclk));
	jor g0996(.dina(n1310),.dinb(n1297),.dout(n1311),.clk(gclk));
	jand g0997(.dina(G208),.dinb(w_G18_19[1]),.dout(n1312),.clk(gclk));
	jor g0998(.dina(w_dff_B_fQnMEHd96_0),.dinb(w_n1189_0[0]),.dout(n1313),.clk(gclk));
	jxor g0999(.dina(w_n878_0[0]),.dinb(w_n869_0[0]),.dout(n1314),.clk(gclk));
	jxor g1000(.dina(w_n899_0[0]),.dinb(w_n891_0[1]),.dout(n1315),.clk(gclk));
	jxor g1001(.dina(n1315),.dinb(n1314),.dout(n1316),.clk(gclk));
	jxor g1002(.dina(n1316),.dinb(w_dff_B_1bITEiIi8_1),.dout(n1317),.clk(gclk));
	jnot g1003(.din(w_n916_0[0]),.dout(n1318),.clk(gclk));
	jxor g1004(.dina(w_n945_0[1]),.dinb(w_n927_0[0]),.dout(n1319),.clk(gclk));
	jxor g1005(.dina(n1319),.dinb(n1318),.dout(n1320),.clk(gclk));
	jnot g1006(.din(G198),.dout(n1321),.clk(gclk));
	jor g1007(.dina(n1321),.dinb(w_n355_9[0]),.dout(n1322),.clk(gclk));
	jand g1008(.dina(n1322),.dinb(w_n353_0[0]),.dout(n1323),.clk(gclk));
	jxor g1009(.dina(w_dff_B_TQzO71He6_0),.dinb(w_n908_0[0]),.dout(n1324),.clk(gclk));
	jxor g1010(.dina(w_dff_B_pyGI4mB35_0),.dinb(n1320),.dout(n1325),.clk(gclk));
	jand g1011(.dina(w_n1325_0[1]),.dinb(w_n1317_0[1]),.dout(n1326),.clk(gclk));
	jnot g1012(.din(w_n1301_0[0]),.dout(n1327),.clk(gclk));
	jnot g1013(.din(w_n1309_0[0]),.dout(n1328),.clk(gclk));
	jand g1014(.dina(n1328),.dinb(w_dff_B_dmVOihU45_1),.dout(n1329),.clk(gclk));
	jnot g1015(.din(w_n1317_0[0]),.dout(n1330),.clk(gclk));
	jnot g1016(.din(w_n1325_0[0]),.dout(n1331),.clk(gclk));
	jand g1017(.dina(n1331),.dinb(n1330),.dout(n1332),.clk(gclk));
	jor g1018(.dina(n1332),.dinb(n1329),.dout(n1333),.clk(gclk));
	jor g1019(.dina(n1333),.dinb(w_dff_B_MovuNc1j0_1),.dout(n1334),.clk(gclk));
	jor g1020(.dina(n1334),.dinb(w_dff_B_jGiJQ0wV2_1),.dout(n1335),.clk(gclk));
	jxor g1021(.dina(w_n744_0[0]),.dinb(w_n730_0[0]),.dout(n1336),.clk(gclk));
	jxor g1022(.dina(n1336),.dinb(w_n737_0[0]),.dout(n1337),.clk(gclk));
	jxor g1023(.dina(w_n754_0[0]),.dinb(w_n723_0[0]),.dout(n1338),.clk(gclk));
	jnot g1024(.din(w_n994_0[0]),.dout(n1339),.clk(gclk));
	jand g1025(.dina(w_n1016_0[0]),.dinb(n1339),.dout(n1340),.clk(gclk));
	jnot g1026(.din(w_n1015_0[0]),.dout(n1341),.clk(gclk));
	jand g1027(.dina(n1341),.dinb(w_n995_0[0]),.dout(n1342),.clk(gclk));
	jor g1028(.dina(n1342),.dinb(n1340),.dout(n1343),.clk(gclk));
	jnot g1029(.din(w_n987_0[0]),.dout(n1344),.clk(gclk));
	jand g1030(.dina(w_n1009_0[1]),.dinb(n1344),.dout(n1345),.clk(gclk));
	jnot g1031(.din(w_n1008_0[0]),.dout(n1346),.clk(gclk));
	jand g1032(.dina(n1346),.dinb(w_n988_0[0]),.dout(n1347),.clk(gclk));
	jor g1033(.dina(n1347),.dinb(n1345),.dout(n1348),.clk(gclk));
	jxor g1034(.dina(n1348),.dinb(n1343),.dout(n1349),.clk(gclk));
	jnot g1035(.din(G181),.dout(n1350),.clk(gclk));
	jor g1036(.dina(n1350),.dinb(w_n355_8[2]),.dout(n1351),.clk(gclk));
	jand g1037(.dina(n1351),.dinb(w_n1166_0[0]),.dout(n1352),.clk(gclk));
	jxor g1038(.dina(w_dff_B_2f6GBAe88_0),.dinb(n1349),.dout(n1353),.clk(gclk));
	jxor g1039(.dina(n1353),.dinb(w_dff_B_8iWpoCgo4_1),.dout(n1354),.clk(gclk));
	jxor g1040(.dina(n1354),.dinb(w_dff_B_OXiC4uOZ9_1),.dout(n1355),.clk(gclk));
	jor g1041(.dina(w_dff_B_kKkyU2GE6_0),.dinb(n1335),.dout(G416_fa_),.clk(gclk));
	jnot g1042(.din(w_n372_1[0]),.dout(n1357),.clk(gclk));
	jxor g1043(.dina(w_n377_0[1]),.dinb(w_G3717_1[0]),.dout(n1358),.clk(gclk));
	jand g1044(.dina(w_dff_B_dxIieSIK9_0),.dinb(n1357),.dout(n1359),.clk(gclk));
	jnot g1045(.din(w_n387_0[1]),.dout(n1360),.clk(gclk));
	jxor g1046(.dina(w_n401_0[2]),.dinb(w_G3705_1[1]),.dout(n1361),.clk(gclk));
	jand g1047(.dina(w_n1361_0[1]),.dinb(w_n362_0[1]),.dout(n1362),.clk(gclk));
	jand g1048(.dina(w_n1362_0[1]),.dinb(w_G4526_0[2]),.dout(n1363),.clk(gclk));
	jand g1049(.dina(n1363),.dinb(w_n1360_1[1]),.dout(n1364),.clk(gclk));
	jand g1050(.dina(n1364),.dinb(w_n1359_0[2]),.dout(n1365),.clk(gclk));
	jnot g1051(.din(w_n407_0[1]),.dout(n1366),.clk(gclk));
	jand g1052(.dina(w_n1361_0[0]),.dinb(w_n390_1[0]),.dout(n1367),.clk(gclk));
	jand g1053(.dina(n1367),.dinb(w_n1360_1[0]),.dout(n1368),.clk(gclk));
	jor g1054(.dina(n1368),.dinb(w_dff_B_pO9vYmEx8_1),.dout(n1369),.clk(gclk));
	jand g1055(.dina(n1369),.dinb(w_n1359_0[1]),.dout(n1370),.clk(gclk));
	jnot g1056(.din(w_n413_0[2]),.dout(n1371),.clk(gclk));
	jand g1057(.dina(n1371),.dinb(w_n1359_0[0]),.dout(n1372),.clk(gclk));
	jnot g1058(.din(w_n419_0[0]),.dout(n1373),.clk(gclk));
	jor g1059(.dina(n1373),.dinb(n1372),.dout(n1374),.clk(gclk));
	jor g1060(.dina(n1374),.dinb(n1370),.dout(n1375),.clk(gclk));
	jor g1061(.dina(n1375),.dinb(n1365),.dout(n1376),.clk(gclk));
	jnot g1062(.din(w_n452_0[0]),.dout(n1377),.clk(gclk));
	jand g1063(.dina(w_dff_B_3o2Gmpu88_0),.dinb(w_n1376_0[1]),.dout(n1378),.clk(gclk));
	jnot g1064(.din(w_n464_0[0]),.dout(n1379),.clk(gclk));
	jor g1065(.dina(n1379),.dinb(n1378),.dout(n1380),.clk(gclk));
	jand g1066(.dina(w_n494_0[0]),.dinb(w_n1380_1[1]),.dout(n1381),.clk(gclk));
	jnot g1067(.din(w_n518_0[0]),.dout(n1382),.clk(gclk));
	jor g1068(.dina(n1382),.dinb(n1381),.dout(n1383),.clk(gclk));
	jand g1069(.dina(w_n542_0[0]),.dinb(w_n1383_1[2]),.dout(n1384),.clk(gclk));
	jor g1070(.dina(w_n560_0[0]),.dinb(n1384),.dout(n1385),.clk(gclk));
	jxor g1071(.dina(w_n578_1[0]),.dinb(w_n1385_1[1]),.dout(w_dff_A_R2mLLwKi2_2),.clk(gclk));
	jand g1072(.dina(w_n592_0[0]),.dinb(w_n1385_1[0]),.dout(n1387),.clk(gclk));
	jnot g1073(.din(w_n617_0[0]),.dout(n1388),.clk(gclk));
	jor g1074(.dina(w_dff_B_UGxZ7lFd5_0),.dinb(n1387),.dout(n1389),.clk(gclk));
	jand g1075(.dina(w_n637_0[0]),.dinb(w_n1389_1[1]),.dout(n1390),.clk(gclk));
	jnot g1076(.din(w_n656_0[0]),.dout(n1391),.clk(gclk));
	jor g1077(.dina(w_dff_B_gtNNXPav0_0),.dinb(n1390),.dout(n1392),.clk(gclk));
	jxor g1078(.dina(w_n678_0[1]),.dinb(w_n1392_1[1]),.dout(w_dff_A_kWtpVriV9_2),.clk(gclk));
	jor g1079(.dina(w_n1033_0[0]),.dinb(w_n957_0[0]),.dout(n1394),.clk(gclk));
	jand g1080(.dina(n1394),.dinb(w_n905_0[0]),.dout(n1395),.clk(gclk));
	jor g1081(.dina(n1395),.dinb(w_n1044_0[0]),.dout(n1396),.clk(gclk));
	jand g1082(.dina(n1396),.dinb(w_n864_0[0]),.dout(n1397),.clk(gclk));
	jor g1083(.dina(n1397),.dinb(w_n981_0[0]),.dout(n1398),.clk(gclk));
	jand g1084(.dina(n1398),.dinb(w_n810_0[0]),.dout(n1399),.clk(gclk));
	jor g1085(.dina(n1399),.dinb(w_n972_0[0]),.dout(w_dff_A_jUZ9oWmy2_2),.clk(gclk));
	jnot g1086(.din(w_n568_0[1]),.dout(n1401),.clk(gclk));
	jnot g1087(.din(w_n584_0[1]),.dout(n1402),.clk(gclk));
	jnot g1088(.din(w_n589_1[0]),.dout(n1403),.clk(gclk));
	jnot g1089(.din(w_n579_0[1]),.dout(n1404),.clk(gclk));
	jor g1090(.dina(w_n1404_0[1]),.dinb(w_n562_0[1]),.dout(n1405),.clk(gclk));
	jor g1091(.dina(w_n1405_0[1]),.dinb(w_n1403_0[1]),.dout(n1406),.clk(gclk));
	jor g1092(.dina(w_n1406_0[1]),.dinb(w_n1402_0[1]),.dout(n1407),.clk(gclk));
	jand g1093(.dina(n1407),.dinb(w_n615_1[0]),.dout(n1408),.clk(gclk));
	jxor g1094(.dina(n1408),.dinb(w_n1401_0[1]),.dout(w_dff_A_bs3dCZUn0_2),.clk(gclk));
	jand g1095(.dina(w_n1406_0[0]),.dinb(w_n613_0[1]),.dout(n1410),.clk(gclk));
	jxor g1096(.dina(n1410),.dinb(w_n1402_0[0]),.dout(w_dff_A_amWUnRaU2_2),.clk(gclk));
	jnot g1097(.din(w_n608_0[1]),.dout(n1412),.clk(gclk));
	jnot g1098(.din(w_n607_0[0]),.dout(n1413),.clk(gclk));
	jand g1099(.dina(n1413),.dinb(w_dff_B_bMdm3kIy3_1),.dout(n1414),.clk(gclk));
	jand g1100(.dina(w_n1414_0[1]),.dinb(w_n1405_0[0]),.dout(n1415),.clk(gclk));
	jxor g1101(.dina(n1415),.dinb(w_n1403_0[0]),.dout(w_dff_A_hR2WjjY39_2),.clk(gclk));
	jand g1102(.dina(w_n578_0[2]),.dinb(w_n1385_0[2]),.dout(n1417),.clk(gclk));
	jor g1103(.dina(n1417),.dinb(w_n606_1[1]),.dout(n1418),.clk(gclk));
	jxor g1104(.dina(n1418),.dinb(w_n573_0[2]),.dout(w_dff_A_DEUGBpxE4_2),.clk(gclk));
	jnot g1105(.din(w_n661_0[0]),.dout(n1420),.clk(gclk));
	jnot g1106(.din(w_n665_0[1]),.dout(n1421),.clk(gclk));
	jnot g1107(.din(w_n669_0[1]),.dout(n1422),.clk(gclk));
	jnot g1108(.din(w_n679_1[0]),.dout(n1423),.clk(gclk));
	jor g1109(.dina(w_dff_B_PUHfyred4_0),.dinb(w_n657_1[0]),.dout(n1424),.clk(gclk));
	jor g1110(.dina(w_n1424_0[1]),.dinb(w_n1422_0[1]),.dout(n1425),.clk(gclk));
	jor g1111(.dina(w_n1425_0[1]),.dinb(w_n1421_0[1]),.dout(n1426),.clk(gclk));
	jand g1112(.dina(n1426),.dinb(w_n704_0[0]),.dout(n1427),.clk(gclk));
	jxor g1113(.dina(n1427),.dinb(w_n1420_0[2]),.dout(w_dff_A_AdXSab4c0_2),.clk(gclk));
	jnot g1114(.din(w_n701_1[0]),.dout(n1429),.clk(gclk));
	jand g1115(.dina(w_n1425_0[0]),.dinb(w_dff_B_wHaSt9t09_1),.dout(n1430),.clk(gclk));
	jxor g1116(.dina(n1430),.dinb(w_n1421_0[0]),.dout(w_dff_A_tDqTzf6y5_2),.clk(gclk));
	jnot g1117(.din(w_n699_1[0]),.dout(n1432),.clk(gclk));
	jand g1118(.dina(w_n1424_0[0]),.dinb(w_dff_B_PYxL9Co86_1),.dout(n1433),.clk(gclk));
	jxor g1119(.dina(n1433),.dinb(w_n1422_0[0]),.dout(w_dff_A_pC7Cjpvr8_2),.clk(gclk));
	jand g1120(.dina(w_n678_0[0]),.dinb(w_n1392_1[0]),.dout(n1435),.clk(gclk));
	jor g1121(.dina(n1435),.dinb(w_n697_0[1]),.dout(n1436),.clk(gclk));
	jxor g1122(.dina(n1436),.dinb(w_n674_1[0]),.dout(w_dff_A_pWEqVmr15_2),.clk(gclk));
	jor g1123(.dina(w_G408_0),.dinb(w_G404_0),.dout(n1438),.clk(gclk));
	jor g1124(.dina(w_G410_0),.dinb(w_G406_0),.dout(n1439),.clk(gclk));
	jor g1125(.dina(n1439),.dinb(n1438),.dout(n1440),.clk(gclk));
	jor g1126(.dina(w_dff_B_bln28hL01_0),.dinb(w_G412_0),.dout(n1441),.clk(gclk));
	jor g1127(.dina(w_dff_B_hCYdVrMU3_0),.dinb(w_G416_0),.dout(n1442),.clk(gclk));
	jor g1128(.dina(n1442),.dinb(w_G414_0),.dout(w_dff_A_8GhQPmXM9_2),.clk(gclk));
	jnot g1129(.din(w_n631_0[0]),.dout(n1444),.clk(gclk));
	jnot g1130(.din(w_n627_0[0]),.dout(n1445),.clk(gclk));
	jor g1131(.dina(w_n1445_0[1]),.dinb(w_n618_0[1]),.dout(n1446),.clk(gclk));
	jand g1132(.dina(n1446),.dinb(w_n648_0[1]),.dout(n1447),.clk(gclk));
	jor g1133(.dina(w_n1447_0[1]),.dinb(w_n653_1[0]),.dout(n1448),.clk(gclk));
	jand g1134(.dina(n1448),.dinb(w_n643_0[0]),.dout(n1449),.clk(gclk));
	jxor g1135(.dina(n1449),.dinb(w_n1444_0[2]),.dout(w_dff_A_BfQSCrDb1_2),.clk(gclk));
	jnot g1136(.din(w_n635_0[1]),.dout(n1451),.clk(gclk));
	jxor g1137(.dina(w_n1447_0[0]),.dinb(w_dff_B_hvcuFbb39_1),.dout(w_dff_A_LvjRIxn72_2),.clk(gclk));
	jand g1138(.dina(w_n1156_0[0]),.dinb(w_G2239_0[1]),.dout(n1453),.clk(gclk));
	jnot g1139(.din(n1453),.dout(n1454),.clk(gclk));
	jand g1140(.dina(w_n1454_0[1]),.dinb(w_n1389_1[0]),.dout(n1455),.clk(gclk));
	jor g1141(.dina(n1455),.dinb(w_n645_0[1]),.dout(n1456),.clk(gclk));
	jxor g1142(.dina(n1456),.dinb(w_n622_0[2]),.dout(w_dff_A_9o2BrKL15_2),.clk(gclk));
	jxor g1143(.dina(w_n626_0[0]),.dinb(w_n1389_0[2]),.dout(w_dff_A_TB6D4vo83_2),.clk(gclk));
	jxor g1144(.dina(w_n480_1[0]),.dinb(w_n1380_1[0]),.dout(w_dff_A_VdTQjnjS5_2),.clk(gclk));
	jnot g1145(.din(w_n714_0[0]),.dout(n1460),.clk(gclk));
	jnot g1146(.din(w_n365_0[0]),.dout(n1461),.clk(gclk));
	jor g1147(.dina(w_n711_0[0]),.dinb(w_n710_0[0]),.dout(n1462),.clk(gclk));
	jxor g1148(.dina(w_dff_B_rN5cNUVh2_0),.dinb(n1461),.dout(n1463),.clk(gclk));
	jnot g1149(.din(w_n1463_0[2]),.dout(n1464),.clk(gclk));
	jor g1150(.dina(w_n1464_0[1]),.dinb(n1460),.dout(n1465),.clk(gclk));
	jand g1151(.dina(w_n1465_0[1]),.dinb(w_n715_0[1]),.dout(w_dff_A_m62Wobqa2_2),.clk(gclk));
	jxor g1152(.dina(w_n713_1[0]),.dinb(w_n709_1[0]),.dout(w_dff_A_WnsCWwMe4_2),.clk(gclk));
	jnot g1153(.din(w_n470_0[1]),.dout(n1468),.clk(gclk));
	jnot g1154(.din(w_n486_0[1]),.dout(n1469),.clk(gclk));
	jnot g1155(.din(w_n491_1[0]),.dout(n1470),.clk(gclk));
	jnot g1156(.din(w_n481_0[1]),.dout(n1471),.clk(gclk));
	jor g1157(.dina(w_n1471_0[1]),.dinb(w_n465_0[1]),.dout(n1472),.clk(gclk));
	jor g1158(.dina(w_n1472_0[1]),.dinb(w_n1470_0[1]),.dout(n1473),.clk(gclk));
	jor g1159(.dina(w_n1473_0[1]),.dinb(w_n1469_0[1]),.dout(n1474),.clk(gclk));
	jand g1160(.dina(n1474),.dinb(w_n516_0[1]),.dout(n1475),.clk(gclk));
	jxor g1161(.dina(n1475),.dinb(w_n1468_0[1]),.dout(w_dff_A_I98csHOR7_2),.clk(gclk));
	jand g1162(.dina(w_n1473_0[0]),.dinb(w_n514_0[1]),.dout(n1477),.clk(gclk));
	jxor g1163(.dina(n1477),.dinb(w_n1469_0[0]),.dout(w_dff_A_4R0St17A7_2),.clk(gclk));
	jand g1164(.dina(w_n508_0[0]),.dinb(w_n510_0[0]),.dout(n1479),.clk(gclk));
	jand g1165(.dina(w_n1479_0[1]),.dinb(w_n1472_0[0]),.dout(n1480),.clk(gclk));
	jxor g1166(.dina(n1480),.dinb(w_n1470_0[0]),.dout(w_dff_A_y4w19iT65_2),.clk(gclk));
	jnot g1167(.din(w_n507_1[1]),.dout(n1482),.clk(gclk));
	jand g1168(.dina(w_n480_0[2]),.dinb(w_n1380_0[2]),.dout(n1483),.clk(gclk));
	jor g1169(.dina(n1483),.dinb(w_n1482_0[1]),.dout(n1484),.clk(gclk));
	jxor g1170(.dina(n1484),.dinb(w_n475_0[2]),.dout(w_dff_A_8IAwW4586_2),.clk(gclk));
	jand g1171(.dina(w_n530_0[0]),.dinb(w_n1383_1[1]),.dout(n1486),.clk(gclk));
	jand g1172(.dina(w_n1486_0[1]),.dinb(w_n552_0[0]),.dout(n1487),.clk(gclk));
	jor g1173(.dina(n1487),.dinb(w_n558_0[1]),.dout(n1488),.clk(gclk));
	jxor g1174(.dina(n1488),.dinb(w_n535_1[0]),.dout(w_dff_A_fT0oI7CZ9_2),.clk(gclk));
	jor g1175(.dina(w_n1486_0[0]),.dinb(w_n556_0[1]),.dout(n1490),.clk(gclk));
	jxor g1176(.dina(n1490),.dinb(w_n540_0[1]),.dout(w_dff_A_aLzr4soI2_2),.clk(gclk));
	jnot g1177(.din(w_n528_0[1]),.dout(n1492),.clk(gclk));
	jand g1178(.dina(n1492),.dinb(w_G4420_0[1]),.dout(n1493),.clk(gclk));
	jnot g1179(.din(n1493),.dout(n1494),.clk(gclk));
	jand g1180(.dina(w_n1494_0[2]),.dinb(w_n1383_1[0]),.dout(n1495),.clk(gclk));
	jor g1181(.dina(n1495),.dinb(w_n554_0[1]),.dout(n1496),.clk(gclk));
	jxor g1182(.dina(n1496),.dinb(w_n524_1[2]),.dout(w_dff_A_cdExsKih7_2),.clk(gclk));
	jxor g1183(.dina(w_n529_0[0]),.dinb(w_n1383_0[2]),.dout(w_dff_A_JyIKjTuE8_2),.clk(gclk));
	jxor g1184(.dina(w_n589_0[2]),.dinb(w_n584_0[0]),.dout(n1499),.clk(gclk));
	jxor g1185(.dina(n1499),.dinb(w_n635_0[0]),.dout(n1500),.clk(gclk));
	jnot g1186(.din(w_n622_0[1]),.dout(n1501),.clk(gclk));
	jnot g1187(.din(w_n653_0[2]),.dout(n1502),.clk(gclk));
	jand g1188(.dina(w_n647_0[0]),.dinb(n1502),.dout(n1503),.clk(gclk));
	jor g1189(.dina(w_dff_B_GRpJRWRw0_0),.dinb(w_n649_0[0]),.dout(n1504),.clk(gclk));
	jxor g1190(.dina(n1504),.dinb(w_n1444_0[1]),.dout(n1505),.clk(gclk));
	jxor g1191(.dina(n1505),.dinb(w_n1501_0[1]),.dout(n1506),.clk(gclk));
	jxor g1192(.dina(n1506),.dinb(w_n1454_0[0]),.dout(n1507),.clk(gclk));
	jand g1193(.dina(w_dff_B_yIW1yNUH0_0),.dinb(w_n618_0[0]),.dout(n1508),.clk(gclk));
	jxor g1194(.dina(w_n645_0[0]),.dinb(w_n1501_0[0]),.dout(n1509),.clk(gclk));
	jand g1195(.dina(w_n648_0[0]),.dinb(w_n1445_0[0]),.dout(n1510),.clk(gclk));
	jnot g1196(.din(w_n1510_0[1]),.dout(n1511),.clk(gclk));
	jor g1197(.dina(n1511),.dinb(w_n642_0[0]),.dout(n1512),.clk(gclk));
	jor g1198(.dina(w_n1510_0[0]),.dinb(w_n653_0[1]),.dout(n1513),.clk(gclk));
	jand g1199(.dina(w_dff_B_rzNwJKfw7_0),.dinb(n1512),.dout(n1514),.clk(gclk));
	jxor g1200(.dina(n1514),.dinb(w_n1444_0[0]),.dout(n1515),.clk(gclk));
	jxor g1201(.dina(n1515),.dinb(w_dff_B_1qVDS2KB7_1),.dout(n1516),.clk(gclk));
	jand g1202(.dina(w_dff_B_eiKQTK2w9_0),.dinb(w_n1389_0[1]),.dout(n1517),.clk(gclk));
	jor g1203(.dina(n1517),.dinb(n1508),.dout(n1518),.clk(gclk));
	jand g1204(.dina(w_n613_0[0]),.dinb(w_n606_1[0]),.dout(n1519),.clk(gclk));
	jnot g1205(.din(w_n606_0[2]),.dout(n1520),.clk(gclk));
	jand g1206(.dina(w_n605_0[0]),.dinb(w_n1520_0[1]),.dout(n1521),.clk(gclk));
	jand g1207(.dina(n1521),.dinb(w_n610_0[0]),.dout(n1522),.clk(gclk));
	jxor g1208(.dina(n1522),.dinb(w_n578_0[1]),.dout(n1523),.clk(gclk));
	jor g1209(.dina(n1523),.dinb(n1519),.dout(n1524),.clk(gclk));
	jor g1210(.dina(w_n572_0[1]),.dinb(w_n569_0[0]),.dout(n1525),.clk(gclk));
	jand g1211(.dina(w_n1520_0[0]),.dinb(w_dff_B_N6gXHevE0_1),.dout(n1526),.clk(gclk));
	jor g1212(.dina(n1526),.dinb(w_n608_0[0]),.dout(n1527),.clk(gclk));
	jxor g1213(.dina(w_dff_B_jAFUiruS4_0),.dinb(w_n615_0[2]),.dout(n1528),.clk(gclk));
	jxor g1214(.dina(n1528),.dinb(w_n1401_0[0]),.dout(n1529),.clk(gclk));
	jxor g1215(.dina(n1529),.dinb(w_dff_B_U1goTxm30_1),.dout(n1530),.clk(gclk));
	jor g1216(.dina(w_dff_B_1sUUPRfg5_0),.dinb(w_n1385_0[1]),.dout(n1531),.clk(gclk));
	jand g1217(.dina(w_n1414_0[0]),.dinb(w_n1404_0[0]),.dout(n1532),.clk(gclk));
	jxor g1218(.dina(n1532),.dinb(w_n568_0[0]),.dout(n1533),.clk(gclk));
	jxor g1219(.dina(w_n606_0[1]),.dinb(w_n573_0[1]),.dout(n1534),.clk(gclk));
	jand g1220(.dina(w_n589_0[1]),.dinb(w_n579_0[0]),.dout(n1535),.clk(gclk));
	jor g1221(.dina(w_dff_B_pkJzjAA13_0),.dinb(w_n612_0[0]),.dout(n1536),.clk(gclk));
	jnot g1222(.din(w_n1536_0[1]),.dout(n1537),.clk(gclk));
	jand g1223(.dina(n1537),.dinb(w_n599_0[0]),.dout(n1538),.clk(gclk));
	jnot g1224(.din(w_n591_0[0]),.dout(n1539),.clk(gclk));
	jand g1225(.dina(w_n1536_0[0]),.dinb(w_dff_B_H19Doc6T6_1),.dout(n1540),.clk(gclk));
	jand g1226(.dina(w_dff_B_47O9ffhk8_0),.dinb(w_n615_0[1]),.dout(n1541),.clk(gclk));
	jor g1227(.dina(n1541),.dinb(w_dff_B_wa7J2Vx24_1),.dout(n1542),.clk(gclk));
	jxor g1228(.dina(n1542),.dinb(w_dff_B_m54To6v88_1),.dout(n1543),.clk(gclk));
	jxor g1229(.dina(n1543),.dinb(w_dff_B_2ZeCTHMn8_1),.dout(n1544),.clk(gclk));
	jor g1230(.dina(w_dff_B_RDwCv1ed2_0),.dinb(w_n562_0[0]),.dout(n1545),.clk(gclk));
	jand g1231(.dina(n1545),.dinb(n1531),.dout(n1546),.clk(gclk));
	jxor g1232(.dina(w_dff_B_mAKxwxqz1_0),.dinb(n1518),.dout(n1547),.clk(gclk));
	jxor g1233(.dina(n1547),.dinb(w_dff_B_mt6EQCSe3_1),.dout(w_dff_A_3t7SkkRt9_2),.clk(gclk));
	jand g1234(.dina(w_n713_0[2]),.dinb(w_n709_0[2]),.dout(n1549),.clk(gclk));
	jor g1235(.dina(n1549),.dinb(w_n1463_0[1]),.dout(n1550),.clk(gclk));
	jnot g1236(.din(w_n683_0[0]),.dout(n1551),.clk(gclk));
	jand g1237(.dina(w_n707_0[1]),.dinb(w_n1392_0[2]),.dout(n1552),.clk(gclk));
	jand g1238(.dina(w_n712_0[0]),.dinb(w_n708_0[0]),.dout(n1553),.clk(gclk));
	jor g1239(.dina(n1553),.dinb(w_n1464_0[0]),.dout(n1554),.clk(gclk));
	jor g1240(.dina(w_dff_B_8aGUcFe22_0),.dinb(n1552),.dout(n1555),.clk(gclk));
	jor g1241(.dina(n1555),.dinb(n1551),.dout(n1556),.clk(gclk));
	jand g1242(.dina(w_dff_B_yfGAFMFW6_0),.dinb(n1550),.dout(n1557),.clk(gclk));
	jand g1243(.dina(w_n1463_0[0]),.dinb(w_n707_0[0]),.dout(n1558),.clk(gclk));
	jand g1244(.dina(w_dff_B_3ZnM1Mw94_0),.dinb(w_n657_0[2]),.dout(n1559),.clk(gclk));
	jor g1245(.dina(w_dff_B_Id4qsDKp8_0),.dinb(n1557),.dout(n1560),.clk(gclk));
	jxor g1246(.dina(w_n669_0[0]),.dinb(w_n665_0[0]),.dout(n1561),.clk(gclk));
	jor g1247(.dina(w_n701_0[2]),.dinb(w_n686_0[0]),.dout(n1562),.clk(gclk));
	jand g1248(.dina(w_dff_B_4pwTS0wB0_0),.dinb(w_n703_0[0]),.dout(n1563),.clk(gclk));
	jxor g1249(.dina(n1563),.dinb(w_n1420_0[1]),.dout(n1564),.clk(gclk));
	jor g1250(.dina(w_n677_0[0]),.dinb(w_n675_0[0]),.dout(n1565),.clk(gclk));
	jxor g1251(.dina(n1565),.dinb(w_n674_0[2]),.dout(n1566),.clk(gclk));
	jxor g1252(.dina(w_dff_B_JG5CIk200_0),.dinb(w_n699_0[2]),.dout(n1567),.clk(gclk));
	jxor g1253(.dina(w_dff_B_l8UL9uop4_0),.dinb(n1564),.dout(n1568),.clk(gclk));
	jand g1254(.dina(w_dff_B_CVGMQyU47_0),.dinb(w_n657_0[1]),.dout(n1569),.clk(gclk));
	jand g1255(.dina(w_n679_0[2]),.dinb(w_n692_0[0]),.dout(n1570),.clk(gclk));
	jor g1256(.dina(w_dff_B_2rjMd3se2_0),.dinb(w_n701_0[1]),.dout(n1571),.clk(gclk));
	jor g1257(.dina(w_n1571_0[1]),.dinb(w_n687_0[0]),.dout(n1572),.clk(gclk));
	jnot g1258(.din(w_n1571_0[0]),.dout(n1573),.clk(gclk));
	jor g1259(.dina(n1573),.dinb(w_n680_0[0]),.dout(n1574),.clk(gclk));
	jor g1260(.dina(w_dff_B_iEA9xJDk0_0),.dinb(w_n705_0[0]),.dout(n1575),.clk(gclk));
	jand g1261(.dina(n1575),.dinb(w_dff_B_SdDV3byI7_1),.dout(n1576),.clk(gclk));
	jor g1262(.dina(w_n699_0[1]),.dinb(w_n679_0[1]),.dout(n1577),.clk(gclk));
	jxor g1263(.dina(n1577),.dinb(w_n1420_0[0]),.dout(n1578),.clk(gclk));
	jxor g1264(.dina(w_dff_B_OAS7MuBZ6_0),.dinb(n1576),.dout(n1579),.clk(gclk));
	jxor g1265(.dina(n1579),.dinb(w_n697_0[0]),.dout(n1580),.clk(gclk));
	jxor g1266(.dina(n1580),.dinb(w_n674_0[1]),.dout(n1581),.clk(gclk));
	jand g1267(.dina(w_dff_B_gbAOKVfw2_0),.dinb(w_n1392_0[1]),.dout(n1582),.clk(gclk));
	jor g1268(.dina(n1582),.dinb(n1569),.dout(n1583),.clk(gclk));
	jxor g1269(.dina(n1583),.dinb(w_dff_B_Lun4TgfG5_1),.dout(n1584),.clk(gclk));
	jxor g1270(.dina(w_dff_B_L9CTJBsM8_0),.dinb(n1560),.dout(G338),.clk(gclk));
	jxor g1271(.dina(w_n491_0[2]),.dinb(w_n486_0[0]),.dout(n1586),.clk(gclk));
	jxor g1272(.dina(n1586),.dinb(w_n540_0[0]),.dout(n1587),.clk(gclk));
	jnot g1273(.din(w_n535_0[2]),.dout(n1588),.clk(gclk));
	jnot g1274(.din(w_n557_0[0]),.dout(n1589),.clk(gclk));
	jor g1275(.dina(w_n556_0[0]),.dinb(w_n549_0[0]),.dout(n1590),.clk(gclk));
	jand g1276(.dina(w_dff_B_YoGxxV7h9_0),.dinb(n1589),.dout(n1591),.clk(gclk));
	jxor g1277(.dina(n1591),.dinb(w_dff_B_0aFNqMVK8_1),.dout(n1592),.clk(gclk));
	jxor g1278(.dina(w_n1494_0[1]),.dinb(w_n524_1[1]),.dout(n1593),.clk(gclk));
	jxor g1279(.dina(w_dff_B_F3j65Tk89_0),.dinb(n1592),.dout(n1594),.clk(gclk));
	jand g1280(.dina(w_dff_B_H1VZyRNg0_0),.dinb(w_n519_0[0]),.dout(n1595),.clk(gclk));
	jxor g1281(.dina(w_n554_0[0]),.dinb(w_n524_1[0]),.dout(n1596),.clk(gclk));
	jxor g1282(.dina(n1596),.dinb(w_n535_0[1]),.dout(n1597),.clk(gclk));
	jand g1283(.dina(w_n1494_0[0]),.dinb(w_n524_0[2]),.dout(n1598),.clk(gclk));
	jor g1284(.dina(n1598),.dinb(w_n553_0[0]),.dout(n1599),.clk(gclk));
	jnot g1285(.din(w_n1599_0[1]),.dout(n1600),.clk(gclk));
	jand g1286(.dina(n1600),.dinb(w_n558_0[0]),.dout(n1601),.clk(gclk));
	jand g1287(.dina(w_n1599_0[0]),.dinb(w_n551_0[0]),.dout(n1602),.clk(gclk));
	jor g1288(.dina(w_dff_B_7nAtSZzz0_0),.dinb(n1601),.dout(n1603),.clk(gclk));
	jxor g1289(.dina(n1603),.dinb(w_dff_B_AhLXTjoJ4_1),.dout(n1604),.clk(gclk));
	jand g1290(.dina(w_dff_B_alLF9ndC9_0),.dinb(w_n1383_0[1]),.dout(n1605),.clk(gclk));
	jor g1291(.dina(n1605),.dinb(n1595),.dout(n1606),.clk(gclk));
	jor g1292(.dina(w_n474_0[1]),.dinb(w_n471_0[0]),.dout(n1607),.clk(gclk));
	jand g1293(.dina(w_n507_1[0]),.dinb(w_dff_B_dDHCOc7C7_1),.dout(n1608),.clk(gclk));
	jor g1294(.dina(n1608),.dinb(w_n509_0[0]),.dout(n1609),.clk(gclk));
	jnot g1295(.din(w_n516_0[0]),.dout(n1610),.clk(gclk));
	jnot g1296(.din(w_n514_0[0]),.dout(n1611),.clk(gclk));
	jor g1297(.dina(w_n1611_0[1]),.dinb(w_n507_0[2]),.dout(n1612),.clk(gclk));
	jor g1298(.dina(w_n505_0[0]),.dinb(w_n1482_0[0]),.dout(n1613),.clk(gclk));
	jor g1299(.dina(n1613),.dinb(w_n512_0[0]),.dout(n1614),.clk(gclk));
	jxor g1300(.dina(n1614),.dinb(w_n480_0[1]),.dout(n1615),.clk(gclk));
	jand g1301(.dina(w_dff_B_8MEA0ppJ8_0),.dinb(n1612),.dout(n1616),.clk(gclk));
	jxor g1302(.dina(n1616),.dinb(w_n1468_0[0]),.dout(n1617),.clk(gclk));
	jxor g1303(.dina(n1617),.dinb(w_n1610_0[1]),.dout(n1618),.clk(gclk));
	jxor g1304(.dina(n1618),.dinb(w_dff_B_es06gPn80_1),.dout(n1619),.clk(gclk));
	jor g1305(.dina(n1619),.dinb(w_n1380_0[1]),.dout(n1620),.clk(gclk));
	jand g1306(.dina(w_n1479_0[0]),.dinb(w_n1471_0[0]),.dout(n1621),.clk(gclk));
	jxor g1307(.dina(n1621),.dinb(w_n470_0[0]),.dout(n1622),.clk(gclk));
	jxor g1308(.dina(w_n507_0[1]),.dinb(w_n475_0[1]),.dout(n1623),.clk(gclk));
	jand g1309(.dina(w_n491_0[1]),.dinb(w_n481_0[0]),.dout(n1624),.clk(gclk));
	jor g1310(.dina(w_dff_B_bBJAt9h86_0),.dinb(w_n1611_0[0]),.dout(n1625),.clk(gclk));
	jor g1311(.dina(w_n1625_0[1]),.dinb(w_n502_0[0]),.dout(n1626),.clk(gclk));
	jnot g1312(.din(w_n1625_0[0]),.dout(n1627),.clk(gclk));
	jor g1313(.dina(n1627),.dinb(w_n493_0[0]),.dout(n1628),.clk(gclk));
	jor g1314(.dina(n1628),.dinb(w_n1610_0[0]),.dout(n1629),.clk(gclk));
	jand g1315(.dina(n1629),.dinb(w_dff_B_N9Vq1s1r7_1),.dout(n1630),.clk(gclk));
	jxor g1316(.dina(n1630),.dinb(w_dff_B_HgkmMpkq4_1),.dout(n1631),.clk(gclk));
	jxor g1317(.dina(n1631),.dinb(w_dff_B_MIfDYEr94_1),.dout(n1632),.clk(gclk));
	jor g1318(.dina(n1632),.dinb(w_n465_0[0]),.dout(n1633),.clk(gclk));
	jand g1319(.dina(n1633),.dinb(w_dff_B_9R9VV1R75_1),.dout(n1634),.clk(gclk));
	jxor g1320(.dina(n1634),.dinb(w_dff_B_VDYO2Rpt6_1),.dout(n1635),.clk(gclk));
	jxor g1321(.dina(n1635),.dinb(w_dff_B_mcI2YI0y3_1),.dout(w_dff_A_zYe5zPoI5_2),.clk(gclk));
	jxor g1322(.dina(w_n450_0[0]),.dinb(w_n1360_0[2]),.dout(n1637),.clk(gclk));
	jnot g1323(.din(w_n455_0[0]),.dout(n1638),.clk(gclk));
	jnot g1324(.din(w_n460_0[0]),.dout(n1639),.clk(gclk));
	jor g1325(.dina(n1639),.dinb(w_dff_B_mqNpbHV58_1),.dout(n1640),.clk(gclk));
	jand g1326(.dina(n1640),.dinb(w_n461_0[0]),.dout(n1641),.clk(gclk));
	jxor g1327(.dina(n1641),.dinb(w_n446_0[2]),.dout(n1642),.clk(gclk));
	jnot g1328(.din(w_n1642_0[1]),.dout(n1643),.clk(gclk));
	jxor g1329(.dina(w_n1148_0[1]),.dinb(w_n429_1[1]),.dout(n1644),.clk(gclk));
	jnot g1330(.din(w_n1644_0[1]),.dout(n1645),.clk(gclk));
	jor g1331(.dina(w_dff_B_kr9fsSUC8_0),.dinb(n1643),.dout(n1646),.clk(gclk));
	jor g1332(.dina(w_n1644_0[0]),.dinb(w_n1642_0[0]),.dout(n1647),.clk(gclk));
	jand g1333(.dina(n1647),.dinb(w_n422_0[1]),.dout(n1648),.clk(gclk));
	jand g1334(.dina(n1648),.dinb(n1646),.dout(n1649),.clk(gclk));
	jxor g1335(.dina(w_n458_0[0]),.dinb(w_n429_1[0]),.dout(n1650),.clk(gclk));
	jxor g1336(.dina(w_dff_B_toRcHFRg4_0),.dinb(w_n446_0[1]),.dout(n1651),.clk(gclk));
	jnot g1337(.din(w_n462_0[0]),.dout(n1652),.clk(gclk));
	jor g1338(.dina(w_n1148_0[0]),.dinb(w_n429_0[2]),.dout(n1653),.clk(gclk));
	jand g1339(.dina(n1653),.dinb(w_n457_0[0]),.dout(n1654),.clk(gclk));
	jand g1340(.dina(w_n1654_0[1]),.dinb(n1652),.dout(n1655),.clk(gclk));
	jnot g1341(.din(n1655),.dout(n1656),.clk(gclk));
	jnot g1342(.din(w_n456_0[0]),.dout(n1657),.clk(gclk));
	jor g1343(.dina(w_n1654_0[0]),.dinb(n1657),.dout(n1658),.clk(gclk));
	jand g1344(.dina(w_dff_B_c83Pyh6j7_0),.dinb(n1656),.dout(n1659),.clk(gclk));
	jor g1345(.dina(w_n1659_0[1]),.dinb(w_n1651_0[1]),.dout(n1660),.clk(gclk));
	jnot g1346(.din(w_n1651_0[0]),.dout(n1661),.clk(gclk));
	jnot g1347(.din(w_n1659_0[0]),.dout(n1662),.clk(gclk));
	jor g1348(.dina(n1662),.dinb(w_dff_B_ca3YkLIG2_1),.dout(n1663),.clk(gclk));
	jand g1349(.dina(n1663),.dinb(w_n1376_0[0]),.dout(n1664),.clk(gclk));
	jand g1350(.dina(n1664),.dinb(w_dff_B_X5INP1zd1_1),.dout(n1665),.clk(gclk));
	jor g1351(.dina(n1665),.dinb(w_dff_B_db5qHDMU1_1),.dout(n1666),.clk(gclk));
	jand g1352(.dina(w_n1136_0[0]),.dinb(w_n403_0[0]),.dout(n1667),.clk(gclk));
	jnot g1353(.din(w_n1667_0[1]),.dout(n1668),.clk(gclk));
	jor g1354(.dina(n1668),.dinb(w_n1128_0[2]),.dout(n1669),.clk(gclk));
	jnot g1355(.din(w_n1128_0[1]),.dout(n1670),.clk(gclk));
	jand g1356(.dina(w_n1362_0[0]),.dinb(w_n1360_0[1]),.dout(n1671),.clk(gclk));
	jor g1357(.dina(w_dff_B_LG4LL9yI8_0),.dinb(w_n1670_0[1]),.dout(n1672),.clk(gclk));
	jor g1358(.dina(w_n1672_0[1]),.dinb(w_n1667_0[0]),.dout(n1673),.clk(gclk));
	jand g1359(.dina(n1673),.dinb(w_dff_B_HpY57gf01_1),.dout(n1674),.clk(gclk));
	jxor g1360(.dina(n1674),.dinb(w_n372_0[2]),.dout(n1675),.clk(gclk));
	jnot g1361(.din(w_n1672_0[0]),.dout(n1676),.clk(gclk));
	jor g1362(.dina(n1676),.dinb(w_n1127_0[0]),.dout(n1677),.clk(gclk));
	jand g1363(.dina(n1677),.dinb(w_n417_0[0]),.dout(n1678),.clk(gclk));
	jxor g1364(.dina(n1678),.dinb(w_n402_0[1]),.dout(n1679),.clk(gclk));
	jxor g1365(.dina(n1679),.dinb(w_n354_0[2]),.dout(n1680),.clk(gclk));
	jnot g1366(.din(w_n1680_0[1]),.dout(n1681),.clk(gclk));
	jand g1367(.dina(n1681),.dinb(w_n1675_0[1]),.dout(n1682),.clk(gclk));
	jnot g1368(.din(w_n1675_0[0]),.dout(n1683),.clk(gclk));
	jand g1369(.dina(w_n1680_0[0]),.dinb(w_dff_B_TJ6gxjLw2_1),.dout(n1684),.clk(gclk));
	jor g1370(.dina(n1684),.dinb(w_n388_0[0]),.dout(n1685),.clk(gclk));
	jor g1371(.dina(n1685),.dinb(n1682),.dout(n1686),.clk(gclk));
	jxor g1372(.dina(w_n1130_0[0]),.dinb(w_n372_0[1]),.dout(n1687),.clk(gclk));
	jand g1373(.dina(w_n407_0[0]),.dinb(w_n354_0[1]),.dout(n1688),.clk(gclk));
	jand g1374(.dina(n1688),.dinb(w_n413_0[1]),.dout(n1689),.clk(gclk));
	jand g1375(.dina(w_n1689_0[1]),.dinb(w_n395_0[0]),.dout(n1690),.clk(gclk));
	jnot g1376(.din(w_n1689_0[0]),.dout(n1691),.clk(gclk));
	jand g1377(.dina(w_n1670_0[0]),.dinb(w_n390_0[2]),.dout(n1692),.clk(gclk));
	jor g1378(.dina(n1692),.dinb(w_n362_0[0]),.dout(n1693),.clk(gclk));
	jand g1379(.dina(n1693),.dinb(w_dff_B_O5UXEisZ1_1),.dout(n1694),.clk(gclk));
	jor g1380(.dina(n1694),.dinb(w_dff_B_wOKvsKX93_1),.dout(n1695),.clk(gclk));
	jand g1381(.dina(w_n401_0[1]),.dinb(w_G3705_1[0]),.dout(n1696),.clk(gclk));
	jor g1382(.dina(n1696),.dinb(w_n390_0[1]),.dout(n1697),.clk(gclk));
	jand g1383(.dina(n1697),.dinb(w_n412_0[0]),.dout(n1698),.clk(gclk));
	jxor g1384(.dina(w_dff_B_mcHUToWf6_0),.dinb(n1695),.dout(n1699),.clk(gclk));
	jnot g1385(.din(w_n1699_0[1]),.dout(n1700),.clk(gclk));
	jand g1386(.dina(n1700),.dinb(w_n1687_0[1]),.dout(n1701),.clk(gclk));
	jnot g1387(.din(w_n1687_0[0]),.dout(n1702),.clk(gclk));
	jand g1388(.dina(w_n1699_0[0]),.dinb(w_dff_B_lFsbFdkU4_1),.dout(n1703),.clk(gclk));
	jor g1389(.dina(n1703),.dinb(w_G4526_0[1]),.dout(n1704),.clk(gclk));
	jor g1390(.dina(n1704),.dinb(n1701),.dout(n1705),.clk(gclk));
	jand g1391(.dina(w_dff_B_IzjJuRlZ8_0),.dinb(n1686),.dout(n1706),.clk(gclk));
	jxor g1392(.dina(n1706),.dinb(w_n379_0[1]),.dout(n1707),.clk(gclk));
	jxor g1393(.dina(n1707),.dinb(w_dff_B_M2fLyGP78_1),.dout(n1708),.clk(gclk));
	jxor g1394(.dina(n1708),.dinb(w_dff_B_dhPpRk0k0_1),.dout(w_dff_A_QNml90eu3_2),.clk(gclk));
	buf g1395(.din(w_G1_1[1]),.dout(w_dff_A_Jepw3d0D3_1));
	buf g1396(.din(w_G1_1[0]),.dout(w_dff_A_OVoNiMA70_1));
	buf g1397(.din(w_G1459_0[0]),.dout(w_dff_A_At8WbDNn7_1));
	buf g1398(.din(w_G1469_0[1]),.dout(w_dff_A_gI7ydG0x6_1));
	buf g1399(.din(w_G1480_0[0]),.dout(w_dff_A_jVuSQxh25_1));
	buf g1400(.din(w_G1486_0[0]),.dout(w_dff_A_ACjOL8Hd5_1));
	buf g1401(.din(w_G1492_0[1]),.dout(w_dff_A_6cIJftIc7_1));
	buf g1402(.din(w_G1496_0[0]),.dout(w_dff_A_oLMHIQy68_1));
	buf g1403(.din(w_G2208_0[0]),.dout(w_dff_A_PH2dp2Gh6_1));
	buf g1404(.din(w_G2218_0[0]),.dout(w_dff_A_ck3mftU05_1));
	buf g1405(.din(w_G2224_0[1]),.dout(w_dff_A_vip4ZzAz3_1));
	buf g1406(.din(w_G2230_0[1]),.dout(w_dff_A_jyfYMINM3_1));
	buf g1407(.din(w_G2236_0[1]),.dout(w_dff_A_M7WkONvQ8_1));
	buf g1408(.din(w_G2239_0[0]),.dout(w_dff_A_e0o8y8if7_1));
	buf g1409(.din(w_G2247_0[0]),.dout(w_dff_A_XVcUMRCc4_1));
	buf g1410(.din(w_G2253_0[1]),.dout(w_dff_A_2X5xRMEh0_1));
	buf g1411(.din(w_G2256_0[1]),.dout(w_dff_A_UVJM26EF8_1));
	buf g1412(.din(w_G3698_0[0]),.dout(w_dff_A_a6FX4fFz9_1));
	buf g1413(.din(w_G3701_0[1]),.dout(w_dff_A_HMyMtu9z5_1));
	buf g1414(.din(w_G3705_0[2]),.dout(w_dff_A_OHRyQi3h5_1));
	buf g1415(.din(w_G3711_0[1]),.dout(w_dff_A_dqNBR2IS5_1));
	buf g1416(.din(w_G3717_0[2]),.dout(w_dff_A_0ww2XJtm7_1));
	buf g1417(.din(w_G3723_0[1]),.dout(w_dff_A_wEixxhLY1_1));
	buf g1418(.din(w_G3729_0[1]),.dout(w_dff_A_puMfuoYc7_1));
	buf g1419(.din(w_G3737_0[1]),.dout(w_dff_A_Zq66Xln94_1));
	buf g1420(.din(w_G3743_0[1]),.dout(w_dff_A_DDaoXkJA6_1));
	buf g1421(.din(w_G3749_0[1]),.dout(w_dff_A_YECV73dN5_1));
	buf g1422(.din(w_G4393_0[0]),.dout(w_dff_A_9XjXRFMW1_1));
	buf g1423(.din(w_G4400_0[0]),.dout(w_dff_A_oNY1Iu5k2_1));
	buf g1424(.din(w_G4405_0[1]),.dout(w_dff_A_A7hwHenU7_1));
	buf g1425(.din(w_G4410_0[1]),.dout(w_dff_A_5NPOVR0c6_1));
	buf g1426(.din(w_G4415_0[1]),.dout(w_dff_A_lE27KfQ80_1));
	buf g1427(.din(w_G4420_0[0]),.dout(w_dff_A_f8Cco9ft3_1));
	buf g1428(.din(w_G4427_0[0]),.dout(w_dff_A_k7IiztBr1_1));
	buf g1429(.din(w_G4432_0[1]),.dout(w_dff_A_c5MQTItK9_1));
	buf g1430(.din(w_G4437_0[0]),.dout(w_dff_A_xu1agTiB2_1));
	buf g1431(.din(w_G1462_0[0]),.dout(w_dff_A_6UWDOWSA1_1));
	buf g1432(.din(w_G2211_0[0]),.dout(w_dff_A_l4pLZDe96_1));
	buf g1433(.din(w_G4394_0[1]),.dout(w_dff_A_eaYLuokZ0_1));
	buf g1434(.din(w_G1_0[2]),.dout(w_dff_A_bxKrKb576_1));
	buf g1435(.din(w_G106_0[1]),.dout(w_dff_A_lXPJgvRR0_1));
	jnot g1436(.din(w_G15_0[1]),.dout(w_dff_A_eCUBokED4_1),.clk(gclk));
	jor g1437(.dina(w_n345_0[0]),.dinb(w_G5_0[2]),.dout(w_dff_A_FYQc2eRh8_2),.clk(gclk));
	jnot g1438(.din(w_G15_0[0]),.dout(w_dff_A_RVsCS7MB2_1),.clk(gclk));
	jor g1439(.dina(w_n349_0[0]),.dinb(w_G5_0[1]),.dout(w_dff_A_waTYV5cR5_2),.clk(gclk));
	buf g1440(.din(w_G1_0[1]),.dout(w_dff_A_fFEFrf1N6_1));
	jand g1441(.dina(w_n1125_0[1]),.dinb(w_n1122_0[1]),.dout(w_dff_A_5YJ3wHUN2_2),.clk(gclk));
	jor g1442(.dina(w_n720_1[0]),.dinb(w_n716_1[0]),.dout(w_dff_A_FnZbY9aw9_2),.clk(gclk));
	jand g1443(.dina(w_n1125_0[0]),.dinb(w_n1122_0[0]),.dout(w_dff_A_tocXicLV2_2),.clk(gclk));
	jor g1444(.dina(w_n720_0[2]),.dinb(w_n716_0[2]),.dout(w_dff_A_u65loDku7_2),.clk(gclk));
	jor g1445(.dina(w_n720_0[1]),.dinb(w_n716_0[1]),.dout(w_dff_A_rnuc3wek8_2),.clk(gclk));
	jand g1446(.dina(w_n1465_0[0]),.dinb(w_n715_0[0]),.dout(w_dff_A_FCyTexHS6_2),.clk(gclk));
	jxor g1447(.dina(w_n713_0[1]),.dinb(w_n709_0[1]),.dout(w_dff_A_uZI5p8W54_2),.clk(gclk));
	jspl3 jspl3_w_G1_0(.douta(w_G1_0[0]),.doutb(w_G1_0[1]),.doutc(w_G1_0[2]),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_G1_1[0]),.doutb(w_G1_1[1]),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl3 jspl3_w_G5_0(.douta(w_G5_0[0]),.doutb(w_dff_A_tdRIK4cs5_1),.doutc(w_dff_A_QndkNCew9_2),.din(G5));
	jspl3 jspl3_w_G5_1(.douta(w_dff_A_XGfauPzp1_0),.doutb(w_dff_A_IEvszadD0_1),.doutc(w_G5_1[2]),.din(w_G5_0[0]));
	jspl3 jspl3_w_G15_0(.douta(w_G15_0[0]),.doutb(w_G15_0[1]),.doutc(w_G15_0[2]),.din(G15));
	jspl3 jspl3_w_G18_0(.douta(w_G18_0[0]),.doutb(w_G18_0[1]),.doutc(w_G18_0[2]),.din(G18));
	jspl3 jspl3_w_G18_1(.douta(w_G18_1[0]),.doutb(w_G18_1[1]),.doutc(w_G18_1[2]),.din(w_G18_0[0]));
	jspl3 jspl3_w_G18_2(.douta(w_G18_2[0]),.doutb(w_G18_2[1]),.doutc(w_G18_2[2]),.din(w_G18_0[1]));
	jspl3 jspl3_w_G18_3(.douta(w_G18_3[0]),.doutb(w_G18_3[1]),.doutc(w_G18_3[2]),.din(w_G18_0[2]));
	jspl3 jspl3_w_G18_4(.douta(w_G18_4[0]),.doutb(w_G18_4[1]),.doutc(w_G18_4[2]),.din(w_G18_1[0]));
	jspl3 jspl3_w_G18_5(.douta(w_G18_5[0]),.doutb(w_G18_5[1]),.doutc(w_G18_5[2]),.din(w_G18_1[1]));
	jspl3 jspl3_w_G18_6(.douta(w_G18_6[0]),.doutb(w_dff_A_fK8Tqv5j2_1),.doutc(w_dff_A_3OVEMHkP7_2),.din(w_G18_1[2]));
	jspl3 jspl3_w_G18_7(.douta(w_G18_7[0]),.doutb(w_G18_7[1]),.doutc(w_G18_7[2]),.din(w_G18_2[0]));
	jspl3 jspl3_w_G18_8(.douta(w_G18_8[0]),.doutb(w_G18_8[1]),.doutc(w_G18_8[2]),.din(w_G18_2[1]));
	jspl3 jspl3_w_G18_9(.douta(w_G18_9[0]),.doutb(w_G18_9[1]),.doutc(w_G18_9[2]),.din(w_G18_2[2]));
	jspl3 jspl3_w_G18_10(.douta(w_G18_10[0]),.doutb(w_G18_10[1]),.doutc(w_G18_10[2]),.din(w_G18_3[0]));
	jspl3 jspl3_w_G18_11(.douta(w_G18_11[0]),.doutb(w_G18_11[1]),.doutc(w_G18_11[2]),.din(w_G18_3[1]));
	jspl3 jspl3_w_G18_12(.douta(w_G18_12[0]),.doutb(w_G18_12[1]),.doutc(w_G18_12[2]),.din(w_G18_3[2]));
	jspl3 jspl3_w_G18_13(.douta(w_G18_13[0]),.doutb(w_G18_13[1]),.doutc(w_G18_13[2]),.din(w_G18_4[0]));
	jspl3 jspl3_w_G18_14(.douta(w_G18_14[0]),.doutb(w_G18_14[1]),.doutc(w_G18_14[2]),.din(w_G18_4[1]));
	jspl3 jspl3_w_G18_15(.douta(w_G18_15[0]),.doutb(w_G18_15[1]),.doutc(w_G18_15[2]),.din(w_G18_4[2]));
	jspl3 jspl3_w_G18_16(.douta(w_G18_16[0]),.doutb(w_G18_16[1]),.doutc(w_G18_16[2]),.din(w_G18_5[0]));
	jspl3 jspl3_w_G18_17(.douta(w_G18_17[0]),.doutb(w_G18_17[1]),.doutc(w_G18_17[2]),.din(w_G18_5[1]));
	jspl3 jspl3_w_G18_18(.douta(w_G18_18[0]),.doutb(w_G18_18[1]),.doutc(w_G18_18[2]),.din(w_G18_5[2]));
	jspl3 jspl3_w_G18_19(.douta(w_G18_19[0]),.doutb(w_G18_19[1]),.doutc(w_G18_19[2]),.din(w_G18_6[0]));
	jspl3 jspl3_w_G18_20(.douta(w_G18_20[0]),.doutb(w_G18_20[1]),.doutc(w_G18_20[2]),.din(w_G18_6[1]));
	jspl3 jspl3_w_G18_21(.douta(w_G18_21[0]),.doutb(w_G18_21[1]),.doutc(w_G18_21[2]),.din(w_G18_6[2]));
	jspl3 jspl3_w_G18_22(.douta(w_G18_22[0]),.doutb(w_G18_22[1]),.doutc(w_dff_A_jvMIQD1H6_2),.din(w_G18_7[0]));
	jspl3 jspl3_w_G18_23(.douta(w_dff_A_dYIGB10U4_0),.doutb(w_G18_23[1]),.doutc(w_G18_23[2]),.din(w_G18_7[1]));
	jspl3 jspl3_w_G18_24(.douta(w_G18_24[0]),.doutb(w_G18_24[1]),.doutc(w_G18_24[2]),.din(w_G18_7[2]));
	jspl3 jspl3_w_G18_25(.douta(w_G18_25[0]),.doutb(w_G18_25[1]),.doutc(w_G18_25[2]),.din(w_G18_8[0]));
	jspl3 jspl3_w_G18_26(.douta(w_G18_26[0]),.doutb(w_G18_26[1]),.doutc(w_G18_26[2]),.din(w_G18_8[1]));
	jspl3 jspl3_w_G18_27(.douta(w_G18_27[0]),.doutb(w_G18_27[1]),.doutc(w_G18_27[2]),.din(w_G18_8[2]));
	jspl3 jspl3_w_G18_28(.douta(w_G18_28[0]),.doutb(w_G18_28[1]),.doutc(w_G18_28[2]),.din(w_G18_9[0]));
	jspl3 jspl3_w_G18_29(.douta(w_G18_29[0]),.doutb(w_G18_29[1]),.doutc(w_G18_29[2]),.din(w_G18_9[1]));
	jspl3 jspl3_w_G18_30(.douta(w_G18_30[0]),.doutb(w_G18_30[1]),.doutc(w_G18_30[2]),.din(w_G18_9[2]));
	jspl3 jspl3_w_G18_31(.douta(w_G18_31[0]),.doutb(w_G18_31[1]),.doutc(w_G18_31[2]),.din(w_G18_10[0]));
	jspl3 jspl3_w_G18_32(.douta(w_G18_32[0]),.doutb(w_G18_32[1]),.doutc(w_G18_32[2]),.din(w_G18_10[1]));
	jspl3 jspl3_w_G18_33(.douta(w_G18_33[0]),.doutb(w_G18_33[1]),.doutc(w_G18_33[2]),.din(w_G18_10[2]));
	jspl3 jspl3_w_G18_34(.douta(w_G18_34[0]),.doutb(w_G18_34[1]),.doutc(w_G18_34[2]),.din(w_G18_11[0]));
	jspl3 jspl3_w_G18_35(.douta(w_G18_35[0]),.doutb(w_G18_35[1]),.doutc(w_G18_35[2]),.din(w_G18_11[1]));
	jspl3 jspl3_w_G18_36(.douta(w_G18_36[0]),.doutb(w_G18_36[1]),.doutc(w_G18_36[2]),.din(w_G18_11[2]));
	jspl3 jspl3_w_G18_37(.douta(w_G18_37[0]),.doutb(w_G18_37[1]),.doutc(w_G18_37[2]),.din(w_G18_12[0]));
	jspl3 jspl3_w_G18_38(.douta(w_G18_38[0]),.doutb(w_G18_38[1]),.doutc(w_G18_38[2]),.din(w_G18_12[1]));
	jspl3 jspl3_w_G18_39(.douta(w_G18_39[0]),.doutb(w_G18_39[1]),.doutc(w_G18_39[2]),.din(w_G18_12[2]));
	jspl3 jspl3_w_G18_40(.douta(w_G18_40[0]),.doutb(w_G18_40[1]),.doutc(w_G18_40[2]),.din(w_G18_13[0]));
	jspl3 jspl3_w_G18_41(.douta(w_G18_41[0]),.doutb(w_G18_41[1]),.doutc(w_G18_41[2]),.din(w_G18_13[1]));
	jspl3 jspl3_w_G18_42(.douta(w_G18_42[0]),.doutb(w_G18_42[1]),.doutc(w_G18_42[2]),.din(w_G18_13[2]));
	jspl3 jspl3_w_G18_43(.douta(w_G18_43[0]),.doutb(w_G18_43[1]),.doutc(w_G18_43[2]),.din(w_G18_14[0]));
	jspl3 jspl3_w_G18_44(.douta(w_G18_44[0]),.doutb(w_G18_44[1]),.doutc(w_G18_44[2]),.din(w_G18_14[1]));
	jspl3 jspl3_w_G18_45(.douta(w_G18_45[0]),.doutb(w_G18_45[1]),.doutc(w_G18_45[2]),.din(w_G18_14[2]));
	jspl3 jspl3_w_G18_46(.douta(w_G18_46[0]),.doutb(w_G18_46[1]),.doutc(w_G18_46[2]),.din(w_G18_15[0]));
	jspl3 jspl3_w_G18_47(.douta(w_G18_47[0]),.doutb(w_G18_47[1]),.doutc(w_G18_47[2]),.din(w_G18_15[1]));
	jspl3 jspl3_w_G18_48(.douta(w_G18_48[0]),.doutb(w_G18_48[1]),.doutc(w_G18_48[2]),.din(w_G18_15[2]));
	jspl3 jspl3_w_G18_49(.douta(w_G18_49[0]),.doutb(w_G18_49[1]),.doutc(w_G18_49[2]),.din(w_G18_16[0]));
	jspl3 jspl3_w_G18_50(.douta(w_G18_50[0]),.doutb(w_G18_50[1]),.doutc(w_G18_50[2]),.din(w_G18_16[1]));
	jspl3 jspl3_w_G18_51(.douta(w_G18_51[0]),.doutb(w_G18_51[1]),.doutc(w_G18_51[2]),.din(w_G18_16[2]));
	jspl3 jspl3_w_G18_52(.douta(w_G18_52[0]),.doutb(w_G18_52[1]),.doutc(w_G18_52[2]),.din(w_G18_17[0]));
	jspl3 jspl3_w_G18_53(.douta(w_G18_53[0]),.doutb(w_G18_53[1]),.doutc(w_dff_A_FieKRVQY5_2),.din(w_G18_17[1]));
	jspl3 jspl3_w_G18_54(.douta(w_G18_54[0]),.doutb(w_dff_A_Ru4qcSYj5_1),.doutc(w_G18_54[2]),.din(w_G18_17[2]));
	jspl3 jspl3_w_G18_55(.douta(w_dff_A_3oBneEWV8_0),.doutb(w_G18_55[1]),.doutc(w_dff_A_xFyGdOtk0_2),.din(w_G18_18[0]));
	jspl3 jspl3_w_G18_56(.douta(w_dff_A_VIfWgAQG6_0),.doutb(w_G18_56[1]),.doutc(w_dff_A_Cblcpy8O5_2),.din(w_G18_18[1]));
	jspl3 jspl3_w_G18_57(.douta(w_G18_57[0]),.doutb(w_dff_A_sSClofRu0_1),.doutc(w_G18_57[2]),.din(w_G18_18[2]));
	jspl3 jspl3_w_G18_58(.douta(w_G18_58[0]),.doutb(w_G18_58[1]),.doutc(w_dff_A_aOnlIr1H2_2),.din(w_G18_19[0]));
	jspl3 jspl3_w_G38_0(.douta(w_G38_0[0]),.doutb(w_dff_A_RMHGHZKQ8_1),.doutc(w_dff_A_nW69HDsr6_2),.din(G38));
	jspl3 jspl3_w_G38_1(.douta(w_dff_A_3uwX3wIX5_0),.doutb(w_G38_1[1]),.doutc(w_dff_A_SMU084j52_2),.din(w_G38_0[0]));
	jspl3 jspl3_w_G41_0(.douta(w_dff_A_E1lKdqdn1_0),.doutb(w_dff_A_1rd0G7VB5_1),.doutc(w_G41_0[2]),.din(G41));
	jspl jspl_w_G69_0(.douta(w_G69_0[0]),.doutb(w_G69_0[1]),.din(G69));
	jspl jspl_w_G70_0(.douta(w_G70_0[0]),.doutb(w_G70_0[1]),.din(G70));
	jspl3 jspl3_w_G106_0(.douta(w_G106_0[0]),.doutb(w_G106_0[1]),.doutc(w_G106_0[2]),.din(G106));
	jspl jspl_w_G106_1(.douta(w_dff_A_OEopb4TV0_0),.doutb(w_G106_1[1]),.din(w_G106_0[0]));
	jspl jspl_w_G229_0(.douta(w_G229_0[0]),.doutb(w_G229_0[1]),.din(G229));
	jspl3 jspl3_w_G1455_0(.douta(w_G1455_0[0]),.doutb(w_G1455_0[1]),.doutc(w_G1455_0[2]),.din(G1455));
	jspl jspl_w_G1459_0(.douta(w_G1459_0[0]),.doutb(w_dff_A_xh58VgyV7_1),.din(G1459));
	jspl3 jspl3_w_G1462_0(.douta(w_G1462_0[0]),.doutb(w_G1462_0[1]),.doutc(w_G1462_0[2]),.din(G1462));
	jspl3 jspl3_w_G1469_0(.douta(w_G1469_0[0]),.doutb(w_G1469_0[1]),.doutc(w_G1469_0[2]),.din(G1469));
	jspl jspl_w_G1469_1(.douta(w_dff_A_LscgSKAo6_0),.doutb(w_G1469_1[1]),.din(w_G1469_0[0]));
	jspl3 jspl3_w_G1480_0(.douta(w_G1480_0[0]),.doutb(w_G1480_0[1]),.doutc(w_G1480_0[2]),.din(G1480));
	jspl3 jspl3_w_G1486_0(.douta(w_G1486_0[0]),.doutb(w_G1486_0[1]),.doutc(w_G1486_0[2]),.din(G1486));
	jspl3 jspl3_w_G1492_0(.douta(w_G1492_0[0]),.doutb(w_G1492_0[1]),.doutc(w_G1492_0[2]),.din(G1492));
	jspl jspl_w_G1492_1(.douta(w_G1492_1[0]),.doutb(w_G1492_1[1]),.din(w_G1492_0[0]));
	jspl3 jspl3_w_G1496_0(.douta(w_G1496_0[0]),.doutb(w_G1496_0[1]),.doutc(w_G1496_0[2]),.din(G1496));
	jspl3 jspl3_w_G2204_0(.douta(w_G2204_0[0]),.doutb(w_G2204_0[1]),.doutc(w_G2204_0[2]),.din(G2204));
	jspl jspl_w_G2208_0(.douta(w_G2208_0[0]),.doutb(w_dff_A_hwfUxLGL7_1),.din(G2208));
	jspl3 jspl3_w_G2211_0(.douta(w_G2211_0[0]),.doutb(w_G2211_0[1]),.doutc(w_G2211_0[2]),.din(G2211));
	jspl3 jspl3_w_G2218_0(.douta(w_G2218_0[0]),.doutb(w_G2218_0[1]),.doutc(w_G2218_0[2]),.din(G2218));
	jspl3 jspl3_w_G2224_0(.douta(w_G2224_0[0]),.doutb(w_G2224_0[1]),.doutc(w_G2224_0[2]),.din(G2224));
	jspl jspl_w_G2224_1(.douta(w_dff_A_3fPnOUAI5_0),.doutb(w_G2224_1[1]),.din(w_G2224_0[0]));
	jspl3 jspl3_w_G2230_0(.douta(w_G2230_0[0]),.doutb(w_G2230_0[1]),.doutc(w_G2230_0[2]),.din(G2230));
	jspl jspl_w_G2230_1(.douta(w_dff_A_ivVSklLk1_0),.doutb(w_G2230_1[1]),.din(w_G2230_0[0]));
	jspl3 jspl3_w_G2236_0(.douta(w_G2236_0[0]),.doutb(w_G2236_0[1]),.doutc(w_G2236_0[2]),.din(G2236));
	jspl jspl_w_G2236_1(.douta(w_dff_A_jLE2n0rJ9_0),.doutb(w_G2236_1[1]),.din(w_G2236_0[0]));
	jspl3 jspl3_w_G2239_0(.douta(w_G2239_0[0]),.doutb(w_dff_A_utSlhqib3_1),.doutc(w_G2239_0[2]),.din(G2239));
	jspl3 jspl3_w_G2247_0(.douta(w_G2247_0[0]),.doutb(w_G2247_0[1]),.doutc(w_G2247_0[2]),.din(G2247));
	jspl3 jspl3_w_G2253_0(.douta(w_G2253_0[0]),.doutb(w_G2253_0[1]),.doutc(w_G2253_0[2]),.din(G2253));
	jspl jspl_w_G2253_1(.douta(w_dff_A_u1mi4Nci9_0),.doutb(w_G2253_1[1]),.din(w_G2253_0[0]));
	jspl3 jspl3_w_G2256_0(.douta(w_G2256_0[0]),.doutb(w_G2256_0[1]),.doutc(w_G2256_0[2]),.din(G2256));
	jspl jspl_w_G2256_1(.douta(w_dff_A_TzYAG5a67_0),.doutb(w_G2256_1[1]),.din(w_G2256_0[0]));
	jspl jspl_w_G3698_0(.douta(w_G3698_0[0]),.doutb(w_dff_A_dHpbrnif0_1),.din(G3698));
	jspl3 jspl3_w_G3701_0(.douta(w_dff_A_mENYvAB70_0),.doutb(w_G3701_0[1]),.doutc(w_G3701_0[2]),.din(G3701));
	jspl jspl_w_G3701_1(.douta(w_G3701_1[0]),.doutb(w_dff_A_86X0fj5T4_1),.din(w_G3701_0[0]));
	jspl3 jspl3_w_G3705_0(.douta(w_G3705_0[0]),.doutb(w_G3705_0[1]),.doutc(w_G3705_0[2]),.din(G3705));
	jspl3 jspl3_w_G3705_1(.douta(w_dff_A_OAlXRzLj4_0),.doutb(w_dff_A_PSFGRNPQ9_1),.doutc(w_G3705_1[2]),.din(w_G3705_0[0]));
	jspl jspl_w_G3705_2(.douta(w_dff_A_tQXoU1Lv0_0),.doutb(w_G3705_2[1]),.din(w_G3705_0[1]));
	jspl3 jspl3_w_G3711_0(.douta(w_G3711_0[0]),.doutb(w_G3711_0[1]),.doutc(w_G3711_0[2]),.din(G3711));
	jspl jspl_w_G3711_1(.douta(w_dff_A_W1sTOOLS3_0),.doutb(w_G3711_1[1]),.din(w_G3711_0[0]));
	jspl3 jspl3_w_G3717_0(.douta(w_G3717_0[0]),.doutb(w_dff_A_1cEzrf637_1),.doutc(w_G3717_0[2]),.din(G3717));
	jspl3 jspl3_w_G3717_1(.douta(w_dff_A_5mFDGhUz1_0),.doutb(w_dff_A_4OpryYFd5_1),.doutc(w_G3717_1[2]),.din(w_G3717_0[0]));
	jspl jspl_w_G3717_2(.douta(w_G3717_2[0]),.doutb(w_dff_A_RNZYMGlC6_1),.din(w_G3717_0[1]));
	jspl3 jspl3_w_G3723_0(.douta(w_G3723_0[0]),.doutb(w_G3723_0[1]),.doutc(w_dff_A_AXGb06am4_2),.din(G3723));
	jspl jspl_w_G3723_1(.douta(w_dff_A_dX3Ou6of5_0),.doutb(w_G3723_1[1]),.din(w_G3723_0[0]));
	jspl3 jspl3_w_G3729_0(.douta(w_G3729_0[0]),.doutb(w_G3729_0[1]),.doutc(w_dff_A_5XXE8IiG8_2),.din(G3729));
	jspl jspl_w_G3729_1(.douta(w_dff_A_jLgSfpG66_0),.doutb(w_G3729_1[1]),.din(w_G3729_0[0]));
	jspl3 jspl3_w_G3737_0(.douta(w_G3737_0[0]),.doutb(w_G3737_0[1]),.doutc(w_G3737_0[2]),.din(G3737));
	jspl jspl_w_G3737_1(.douta(w_dff_A_xMIJMFxM8_0),.doutb(w_G3737_1[1]),.din(w_G3737_0[0]));
	jspl3 jspl3_w_G3743_0(.douta(w_dff_A_MoLiEjan8_0),.doutb(w_G3743_0[1]),.doutc(w_G3743_0[2]),.din(G3743));
	jspl3 jspl3_w_G3743_1(.douta(w_dff_A_InQBo1k44_0),.doutb(w_dff_A_BeMhbzOL0_1),.doutc(w_G3743_1[2]),.din(w_G3743_0[0]));
	jspl3 jspl3_w_G3749_0(.douta(w_dff_A_4esZn9dF8_0),.doutb(w_G3749_0[1]),.doutc(w_G3749_0[2]),.din(G3749));
	jspl jspl_w_G3749_1(.douta(w_G3749_1[0]),.doutb(w_G3749_1[1]),.din(w_G3749_0[0]));
	jspl jspl_w_G4393_0(.douta(w_G4393_0[0]),.doutb(w_dff_A_l640jkIo4_1),.din(G4393));
	jspl3 jspl3_w_G4394_0(.douta(w_dff_A_PS3VzGrE0_0),.doutb(w_G4394_0[1]),.doutc(w_G4394_0[2]),.din(G4394));
	jspl jspl_w_G4394_1(.douta(w_G4394_1[0]),.doutb(w_G4394_1[1]),.din(w_G4394_0[0]));
	jspl3 jspl3_w_G4400_0(.douta(w_G4400_0[0]),.doutb(w_G4400_0[1]),.doutc(w_G4400_0[2]),.din(G4400));
	jspl3 jspl3_w_G4405_0(.douta(w_dff_A_Q5yWBHKi1_0),.doutb(w_G4405_0[1]),.doutc(w_G4405_0[2]),.din(G4405));
	jspl3 jspl3_w_G4405_1(.douta(w_G4405_1[0]),.doutb(w_G4405_1[1]),.doutc(w_G4405_1[2]),.din(w_G4405_0[0]));
	jspl3 jspl3_w_G4410_0(.douta(w_G4410_0[0]),.doutb(w_G4410_0[1]),.doutc(w_G4410_0[2]),.din(G4410));
	jspl jspl_w_G4410_1(.douta(w_dff_A_r5O3ypv00_0),.doutb(w_G4410_1[1]),.din(w_G4410_0[0]));
	jspl3 jspl3_w_G4415_0(.douta(w_G4415_0[0]),.doutb(w_G4415_0[1]),.doutc(w_G4415_0[2]),.din(G4415));
	jspl jspl_w_G4415_1(.douta(w_dff_A_X1Xekpxs6_0),.doutb(w_G4415_1[1]),.din(w_G4415_0[0]));
	jspl3 jspl3_w_G4420_0(.douta(w_G4420_0[0]),.doutb(w_dff_A_YC2tkVlL3_1),.doutc(w_G4420_0[2]),.din(G4420));
	jspl jspl_w_G4427_0(.douta(w_G4427_0[0]),.doutb(w_G4427_0[1]),.din(G4427));
	jspl3 jspl3_w_G4432_0(.douta(w_G4432_0[0]),.doutb(w_G4432_0[1]),.doutc(w_G4432_0[2]),.din(G4432));
	jspl jspl_w_G4432_1(.douta(w_dff_A_A9SH6JlV4_0),.doutb(w_G4432_1[1]),.din(w_G4432_0[0]));
	jspl3 jspl3_w_G4437_0(.douta(w_G4437_0[0]),.doutb(w_dff_A_qntVsXhl5_1),.doutc(w_G4437_0[2]),.din(G4437));
	jspl3 jspl3_w_G4526_0(.douta(w_G4526_0[0]),.doutb(w_dff_A_7vaAMfFm2_1),.doutc(w_dff_A_P5m2N7wQ0_2),.din(G4526));
	jspl jspl_w_G4526_1(.douta(w_G4526_1[0]),.doutb(w_dff_A_KWA32Iz23_1),.din(w_G4526_0[0]));
	jspl3 jspl3_w_G4528_0(.douta(w_G4528_0[0]),.doutb(w_G4528_0[1]),.doutc(w_G4528_0[2]),.din(G4528));
	jspl jspl_w_G404_0(.douta(w_G404_0),.doutb(w_dff_A_JtkNZIA12_1),.din(G404_fa_));
	jspl jspl_w_G406_0(.douta(w_G406_0),.doutb(w_dff_A_wBQV3noA7_1),.din(G406_fa_));
	jspl jspl_w_G408_0(.douta(w_G408_0),.doutb(w_dff_A_QqfC4UY36_1),.din(G408_fa_));
	jspl jspl_w_G410_0(.douta(w_G410_0),.doutb(w_dff_A_wN1COxFA1_1),.din(G410_fa_));
	jspl jspl_w_G412_0(.douta(w_G412_0),.doutb(w_dff_A_vKTTodl25_1),.din(G412_fa_));
	jspl jspl_w_G414_0(.douta(w_dff_A_3oTeT6Q66_0),.doutb(w_dff_A_09UngzC83_1),.din(G414_fa_));
	jspl jspl_w_G416_0(.douta(w_G416_0),.doutb(w_dff_A_43cNgcPY5_1),.din(G416_fa_));
	jspl jspl_w_n345_0(.douta(w_n345_0[0]),.doutb(w_n345_0[1]),.din(n345));
	jspl jspl_w_n349_0(.douta(w_n349_0[0]),.doutb(w_n349_0[1]),.din(n349));
	jspl3 jspl3_w_n353_0(.douta(w_n353_0[0]),.doutb(w_n353_0[1]),.doutc(w_n353_0[2]),.din(n353));
	jspl3 jspl3_w_n354_0(.douta(w_n354_0[0]),.doutb(w_n354_0[1]),.doutc(w_dff_A_rNHh4MfQ2_2),.din(w_dff_B_dy0x9oPk3_3));
	jspl3 jspl3_w_n354_1(.douta(w_dff_A_KfyikFRM7_0),.doutb(w_n354_1[1]),.doutc(w_n354_1[2]),.din(w_n354_0[0]));
	jspl3 jspl3_w_n355_0(.douta(w_n355_0[0]),.doutb(w_n355_0[1]),.doutc(w_n355_0[2]),.din(n355));
	jspl3 jspl3_w_n355_1(.douta(w_n355_1[0]),.doutb(w_n355_1[1]),.doutc(w_n355_1[2]),.din(w_n355_0[0]));
	jspl3 jspl3_w_n355_2(.douta(w_n355_2[0]),.doutb(w_n355_2[1]),.doutc(w_n355_2[2]),.din(w_n355_0[1]));
	jspl3 jspl3_w_n355_3(.douta(w_n355_3[0]),.doutb(w_n355_3[1]),.doutc(w_n355_3[2]),.din(w_n355_0[2]));
	jspl3 jspl3_w_n355_4(.douta(w_n355_4[0]),.doutb(w_n355_4[1]),.doutc(w_n355_4[2]),.din(w_n355_1[0]));
	jspl3 jspl3_w_n355_5(.douta(w_n355_5[0]),.doutb(w_n355_5[1]),.doutc(w_n355_5[2]),.din(w_n355_1[1]));
	jspl3 jspl3_w_n355_6(.douta(w_n355_6[0]),.doutb(w_n355_6[1]),.doutc(w_n355_6[2]),.din(w_n355_1[2]));
	jspl3 jspl3_w_n355_7(.douta(w_n355_7[0]),.doutb(w_n355_7[1]),.doutc(w_n355_7[2]),.din(w_n355_2[0]));
	jspl3 jspl3_w_n355_8(.douta(w_n355_8[0]),.doutb(w_n355_8[1]),.doutc(w_n355_8[2]),.din(w_n355_2[1]));
	jspl3 jspl3_w_n355_9(.douta(w_n355_9[0]),.doutb(w_n355_9[1]),.doutc(w_n355_9[2]),.din(w_n355_2[2]));
	jspl3 jspl3_w_n355_10(.douta(w_n355_10[0]),.doutb(w_dff_A_I9KtYtk61_1),.doutc(w_n355_10[2]),.din(w_n355_3[0]));
	jspl3 jspl3_w_n355_11(.douta(w_n355_11[0]),.doutb(w_n355_11[1]),.doutc(w_n355_11[2]),.din(w_n355_3[1]));
	jspl3 jspl3_w_n355_12(.douta(w_n355_12[0]),.doutb(w_n355_12[1]),.doutc(w_n355_12[2]),.din(w_n355_3[2]));
	jspl3 jspl3_w_n355_13(.douta(w_n355_13[0]),.doutb(w_n355_13[1]),.doutc(w_n355_13[2]),.din(w_n355_4[0]));
	jspl3 jspl3_w_n355_14(.douta(w_n355_14[0]),.doutb(w_n355_14[1]),.doutc(w_n355_14[2]),.din(w_n355_4[1]));
	jspl3 jspl3_w_n355_15(.douta(w_n355_15[0]),.doutb(w_n355_15[1]),.doutc(w_n355_15[2]),.din(w_n355_4[2]));
	jspl3 jspl3_w_n355_16(.douta(w_n355_16[0]),.doutb(w_n355_16[1]),.doutc(w_n355_16[2]),.din(w_n355_5[0]));
	jspl3 jspl3_w_n355_17(.douta(w_n355_17[0]),.doutb(w_n355_17[1]),.doutc(w_n355_17[2]),.din(w_n355_5[1]));
	jspl3 jspl3_w_n355_18(.douta(w_n355_18[0]),.doutb(w_n355_18[1]),.doutc(w_n355_18[2]),.din(w_n355_5[2]));
	jspl3 jspl3_w_n355_19(.douta(w_n355_19[0]),.doutb(w_n355_19[1]),.doutc(w_n355_19[2]),.din(w_n355_6[0]));
	jspl3 jspl3_w_n355_20(.douta(w_n355_20[0]),.doutb(w_n355_20[1]),.doutc(w_n355_20[2]),.din(w_n355_6[1]));
	jspl3 jspl3_w_n355_21(.douta(w_n355_21[0]),.doutb(w_n355_21[1]),.doutc(w_n355_21[2]),.din(w_n355_6[2]));
	jspl3 jspl3_w_n355_22(.douta(w_n355_22[0]),.doutb(w_n355_22[1]),.doutc(w_n355_22[2]),.din(w_n355_7[0]));
	jspl3 jspl3_w_n355_23(.douta(w_n355_23[0]),.doutb(w_n355_23[1]),.doutc(w_n355_23[2]),.din(w_n355_7[1]));
	jspl3 jspl3_w_n355_24(.douta(w_n355_24[0]),.doutb(w_n355_24[1]),.doutc(w_n355_24[2]),.din(w_n355_7[2]));
	jspl3 jspl3_w_n355_25(.douta(w_n355_25[0]),.doutb(w_n355_25[1]),.doutc(w_n355_25[2]),.din(w_n355_8[0]));
	jspl jspl_w_n355_26(.douta(w_n355_26[0]),.doutb(w_n355_26[1]),.din(w_n355_8[1]));
	jspl3 jspl3_w_n356_0(.douta(w_dff_A_0qBs17pA6_0),.doutb(w_n356_0[1]),.doutc(w_n356_0[2]),.din(n356));
	jspl jspl_w_n358_0(.douta(w_n358_0[0]),.doutb(w_n358_0[1]),.din(n358));
	jspl jspl_w_n359_0(.douta(w_dff_A_Nbe0h9oQ0_0),.doutb(w_n359_0[1]),.din(n359));
	jspl3 jspl3_w_n362_0(.douta(w_dff_A_QVIFmCto7_0),.doutb(w_n362_0[1]),.doutc(w_n362_0[2]),.din(n362));
	jspl jspl_w_n364_0(.douta(w_n364_0[0]),.doutb(w_n364_0[1]),.din(n364));
	jspl jspl_w_n365_0(.douta(w_n365_0[0]),.doutb(w_dff_A_8jy4uN992_1),.din(n365));
	jspl jspl_w_n366_0(.douta(w_n366_0[0]),.doutb(w_dff_A_2d9BXJgZ3_1),.din(n366));
	jspl jspl_w_n370_0(.douta(w_n370_0[0]),.doutb(w_n370_0[1]),.din(n370));
	jspl3 jspl3_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.doutc(w_n371_0[2]),.din(n371));
	jspl jspl_w_n371_1(.douta(w_n371_1[0]),.doutb(w_n371_1[1]),.din(w_n371_0[0]));
	jspl3 jspl3_w_n372_0(.douta(w_n372_0[0]),.doutb(w_dff_A_qgODzEOp3_1),.doutc(w_dff_A_n14xedSG8_2),.din(n372));
	jspl3 jspl3_w_n372_1(.douta(w_n372_1[0]),.doutb(w_dff_A_IhVKzAON9_1),.doutc(w_dff_A_tITEsiEi1_2),.din(w_n372_0[0]));
	jspl jspl_w_n376_0(.douta(w_n376_0[0]),.doutb(w_n376_0[1]),.din(n376));
	jspl3 jspl3_w_n377_0(.douta(w_n377_0[0]),.doutb(w_n377_0[1]),.doutc(w_dff_A_B7jS1dD42_2),.din(n377));
	jspl3 jspl3_w_n377_1(.douta(w_n377_1[0]),.doutb(w_n377_1[1]),.doutc(w_n377_1[2]),.din(w_n377_0[0]));
	jspl3 jspl3_w_n379_0(.douta(w_n379_0[0]),.doutb(w_dff_A_x0axQ3Bo1_1),.doutc(w_dff_A_WLYOpdFI1_2),.din(n379));
	jspl jspl_w_n379_1(.douta(w_dff_A_k12A8vKM6_0),.doutb(w_n379_1[1]),.din(w_n379_0[0]));
	jspl3 jspl3_w_n380_0(.douta(w_n380_0[0]),.doutb(w_dff_A_hLmf92Cq2_1),.doutc(w_dff_A_qFKh4Mwt1_2),.din(n380));
	jspl jspl_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.din(n385));
	jspl3 jspl3_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.doutc(w_n386_0[2]),.din(n386));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_dff_A_HIATtF3z8_2),.din(n387));
	jspl3 jspl3_w_n387_1(.douta(w_n387_1[0]),.doutb(w_dff_A_lsfaQNUV0_1),.doutc(w_dff_A_S7GzmQcL3_2),.din(w_n387_0[0]));
	jspl3 jspl3_w_n388_0(.douta(w_dff_A_cuIgAHEu2_0),.doutb(w_n388_0[1]),.doutc(w_dff_A_g0dGJFmc4_2),.din(w_dff_B_saPTinh99_3));
	jspl jspl_w_n389_0(.douta(w_n389_0[0]),.doutb(w_dff_A_OMo2FIRs2_1),.din(n389));
	jspl3 jspl3_w_n390_0(.douta(w_n390_0[0]),.doutb(w_n390_0[1]),.doutc(w_dff_A_tq5Yg5jr0_2),.din(w_dff_B_PjRmLE2K8_3));
	jspl jspl_w_n390_1(.douta(w_n390_1[0]),.doutb(w_n390_1[1]),.din(w_n390_0[0]));
	jspl3 jspl3_w_n395_0(.douta(w_dff_A_my3fTdNO3_0),.doutb(w_n395_0[1]),.doutc(w_n395_0[2]),.din(n395));
	jspl jspl_w_n400_0(.douta(w_n400_0[0]),.doutb(w_n400_0[1]),.din(n400));
	jspl3 jspl3_w_n401_0(.douta(w_n401_0[0]),.doutb(w_n401_0[1]),.doutc(w_n401_0[2]),.din(n401));
	jspl3 jspl3_w_n401_1(.douta(w_n401_1[0]),.doutb(w_n401_1[1]),.doutc(w_n401_1[2]),.din(w_n401_0[0]));
	jspl3 jspl3_w_n402_0(.douta(w_n402_0[0]),.doutb(w_dff_A_DwwcC0kn8_1),.doutc(w_dff_A_7BZFgUcx4_2),.din(n402));
	jspl jspl_w_n402_1(.douta(w_n402_1[0]),.doutb(w_dff_A_7Qn0UCgU2_1),.din(w_n402_0[0]));
	jspl jspl_w_n403_0(.douta(w_n403_0[0]),.doutb(w_n403_0[1]),.din(n403));
	jspl jspl_w_n404_0(.douta(w_n404_0[0]),.doutb(w_n404_0[1]),.din(n404));
	jspl3 jspl3_w_n405_0(.douta(w_n405_0[0]),.doutb(w_n405_0[1]),.doutc(w_n405_0[2]),.din(n405));
	jspl3 jspl3_w_n407_0(.douta(w_n407_0[0]),.doutb(w_n407_0[1]),.doutc(w_dff_A_0n0NhMk98_2),.din(n407));
	jspl jspl_w_n408_0(.douta(w_n408_0[0]),.doutb(w_n408_0[1]),.din(n408));
	jspl jspl_w_n410_0(.douta(w_n410_0[0]),.doutb(w_n410_0[1]),.din(n410));
	jspl3 jspl3_w_n412_0(.douta(w_dff_A_b2VlgxhT9_0),.doutb(w_dff_A_tUXNCgyV3_1),.doutc(w_n412_0[2]),.din(n412));
	jspl3 jspl3_w_n413_0(.douta(w_dff_A_XCnpn9aE4_0),.doutb(w_n413_0[1]),.doutc(w_n413_0[2]),.din(n413));
	jspl jspl_w_n413_1(.douta(w_dff_A_MXCZR0Z74_0),.doutb(w_n413_1[1]),.din(w_n413_0[0]));
	jspl3 jspl3_w_n417_0(.douta(w_dff_A_Lz0Uftj19_0),.doutb(w_dff_A_yo6ADf9Q9_1),.doutc(w_n417_0[2]),.din(n417));
	jspl jspl_w_n419_0(.douta(w_n419_0[0]),.doutb(w_dff_A_R2SucpmA7_1),.din(n419));
	jspl3 jspl3_w_n422_0(.douta(w_n422_0[0]),.doutb(w_dff_A_rLLsVKt47_1),.doutc(w_n422_0[2]),.din(n422));
	jspl3 jspl3_w_n422_1(.douta(w_n422_1[0]),.doutb(w_n422_1[1]),.doutc(w_n422_1[2]),.din(w_n422_0[0]));
	jspl jspl_w_n427_0(.douta(w_n427_0[0]),.doutb(w_n427_0[1]),.din(n427));
	jspl3 jspl3_w_n428_0(.douta(w_n428_0[0]),.doutb(w_n428_0[1]),.doutc(w_n428_0[2]),.din(n428));
	jspl3 jspl3_w_n429_0(.douta(w_n429_0[0]),.doutb(w_n429_0[1]),.doutc(w_n429_0[2]),.din(n429));
	jspl3 jspl3_w_n429_1(.douta(w_n429_1[0]),.doutb(w_n429_1[1]),.doutc(w_dff_A_bSXExciB9_2),.din(w_n429_0[0]));
	jspl jspl_w_n429_2(.douta(w_n429_2[0]),.doutb(w_n429_2[1]),.din(w_n429_0[1]));
	jspl jspl_w_n430_0(.douta(w_n430_0[0]),.doutb(w_dff_A_QIQb9Krg9_1),.din(n430));
	jspl jspl_w_n434_0(.douta(w_n434_0[0]),.doutb(w_n434_0[1]),.din(n434));
	jspl3 jspl3_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.doutc(w_n435_0[2]),.din(n435));
	jspl jspl_w_n435_1(.douta(w_n435_1[0]),.doutb(w_n435_1[1]),.din(w_n435_0[0]));
	jspl jspl_w_n436_0(.douta(w_dff_A_lgiSVfCS8_0),.doutb(w_n436_0[1]),.din(n436));
	jspl jspl_w_n437_0(.douta(w_dff_A_TLkKiRen5_0),.doutb(w_n437_0[1]),.din(w_dff_B_3rT1SpkR9_2));
	jspl jspl_w_n441_0(.douta(w_n441_0[0]),.doutb(w_n441_0[1]),.din(n441));
	jspl3 jspl3_w_n442_0(.douta(w_n442_0[0]),.doutb(w_n442_0[1]),.doutc(w_n442_0[2]),.din(n442));
	jspl jspl_w_n443_0(.douta(w_dff_A_JseIA2988_0),.doutb(w_n443_0[1]),.din(n443));
	jspl jspl_w_n445_0(.douta(w_dff_A_ISnzp72h4_0),.doutb(w_n445_0[1]),.din(w_dff_B_TuWjnrE81_2));
	jspl3 jspl3_w_n446_0(.douta(w_n446_0[0]),.doutb(w_n446_0[1]),.doutc(w_dff_A_DD47hUac5_2),.din(n446));
	jspl jspl_w_n446_1(.douta(w_dff_A_jup20k5Y2_0),.doutb(w_n446_1[1]),.din(w_n446_0[0]));
	jspl jspl_w_n448_0(.douta(w_n448_0[0]),.doutb(w_n448_0[1]),.din(n448));
	jspl3 jspl3_w_n449_0(.douta(w_n449_0[0]),.doutb(w_n449_0[1]),.doutc(w_n449_0[2]),.din(n449));
	jspl3 jspl3_w_n450_0(.douta(w_n450_0[0]),.doutb(w_dff_A_7ComxtNr4_1),.doutc(w_dff_A_WGXE9GoW3_2),.din(w_dff_B_xKIuOT5q4_3));
	jspl jspl_w_n452_0(.douta(w_n452_0[0]),.doutb(w_dff_A_jXb34jZa4_1),.din(n452));
	jspl jspl_w_n454_0(.douta(w_n454_0[0]),.doutb(w_n454_0[1]),.din(n454));
	jspl jspl_w_n455_0(.douta(w_n455_0[0]),.doutb(w_dff_A_YbD6cyVf2_1),.din(n455));
	jspl3 jspl3_w_n456_0(.douta(w_n456_0[0]),.doutb(w_dff_A_eqJec2Nj5_1),.doutc(w_dff_A_TE0SQFFm2_2),.din(n456));
	jspl jspl_w_n457_0(.douta(w_n457_0[0]),.doutb(w_n457_0[1]),.din(w_dff_B_aj8GmS9T1_2));
	jspl3 jspl3_w_n458_0(.douta(w_n458_0[0]),.doutb(w_dff_A_AnLtE6ts9_1),.doutc(w_n458_0[2]),.din(n458));
	jspl3 jspl3_w_n460_0(.douta(w_n460_0[0]),.doutb(w_dff_A_CwnsNRDR3_1),.doutc(w_n460_0[2]),.din(n460));
	jspl jspl_w_n461_0(.douta(w_dff_A_njaxN7py0_0),.doutb(w_n461_0[1]),.din(n461));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_dff_A_3ashGlaE8_1),.doutc(w_n462_0[2]),.din(n462));
	jspl jspl_w_n464_0(.douta(w_n464_0[0]),.doutb(w_dff_A_rX7nEYGu3_1),.din(n464));
	jspl3 jspl3_w_n465_0(.douta(w_dff_A_WazBq6Ez1_0),.doutb(w_n465_0[1]),.doutc(w_n465_0[2]),.din(n465));
	jspl jspl_w_n466_0(.douta(w_n466_0[0]),.doutb(w_n466_0[1]),.din(w_dff_B_Sq1hXx1k3_2));
	jspl jspl_w_n468_0(.douta(w_n468_0[0]),.doutb(w_n468_0[1]),.din(n468));
	jspl3 jspl3_w_n469_0(.douta(w_n469_0[0]),.doutb(w_n469_0[1]),.doutc(w_n469_0[2]),.din(n469));
	jspl jspl_w_n469_1(.douta(w_n469_1[0]),.doutb(w_n469_1[1]),.din(w_n469_0[0]));
	jspl3 jspl3_w_n470_0(.douta(w_dff_A_RV0X8r4x8_0),.doutb(w_n470_0[1]),.doutc(w_dff_A_9cGYOAGn6_2),.din(n470));
	jspl3 jspl3_w_n471_0(.douta(w_n471_0[0]),.doutb(w_n471_0[1]),.doutc(w_n471_0[2]),.din(w_dff_B_7v6UQacD2_3));
	jspl jspl_w_n473_0(.douta(w_n473_0[0]),.doutb(w_n473_0[1]),.din(n473));
	jspl3 jspl3_w_n474_0(.douta(w_n474_0[0]),.doutb(w_n474_0[1]),.doutc(w_n474_0[2]),.din(n474));
	jspl jspl_w_n474_1(.douta(w_n474_1[0]),.doutb(w_n474_1[1]),.din(w_n474_0[0]));
	jspl3 jspl3_w_n475_0(.douta(w_n475_0[0]),.doutb(w_dff_A_xgz0nFoM5_1),.doutc(w_dff_A_knNpTlxh2_2),.din(n475));
	jspl jspl_w_n475_1(.douta(w_n475_1[0]),.doutb(w_dff_A_yTBxxcit6_1),.din(w_n475_0[0]));
	jspl jspl_w_n477_0(.douta(w_n477_0[0]),.doutb(w_n477_0[1]),.din(n477));
	jspl jspl_w_n478_0(.douta(w_n478_0[0]),.doutb(w_n478_0[1]),.din(n478));
	jspl jspl_w_n479_0(.douta(w_n479_0[0]),.doutb(w_n479_0[1]),.din(n479));
	jspl3 jspl3_w_n480_0(.douta(w_n480_0[0]),.doutb(w_dff_A_rFFq4SYb4_1),.doutc(w_dff_A_nGLOxQN57_2),.din(n480));
	jspl jspl_w_n480_1(.douta(w_dff_A_VVnNbHzg0_0),.doutb(w_n480_1[1]),.din(w_n480_0[0]));
	jspl3 jspl3_w_n481_0(.douta(w_n481_0[0]),.doutb(w_n481_0[1]),.doutc(w_n481_0[2]),.din(n481));
	jspl jspl_w_n482_0(.douta(w_n482_0[0]),.doutb(w_n482_0[1]),.din(w_dff_B_jCrKePCp9_2));
	jspl jspl_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.din(n484));
	jspl3 jspl3_w_n485_0(.douta(w_n485_0[0]),.doutb(w_n485_0[1]),.doutc(w_n485_0[2]),.din(n485));
	jspl3 jspl3_w_n486_0(.douta(w_dff_A_pd39079P7_0),.doutb(w_n486_0[1]),.doutc(w_dff_A_a1ePKEFb4_2),.din(n486));
	jspl jspl_w_n488_0(.douta(w_n488_0[0]),.doutb(w_n488_0[1]),.din(n488));
	jspl jspl_w_n489_0(.douta(w_n489_0[0]),.doutb(w_n489_0[1]),.din(n489));
	jspl3 jspl3_w_n490_0(.douta(w_n490_0[0]),.doutb(w_n490_0[1]),.doutc(w_n490_0[2]),.din(n490));
	jspl3 jspl3_w_n491_0(.douta(w_n491_0[0]),.doutb(w_dff_A_4UNmYwgZ2_1),.doutc(w_n491_0[2]),.din(n491));
	jspl jspl_w_n491_1(.douta(w_n491_1[0]),.doutb(w_n491_1[1]),.din(w_n491_0[0]));
	jspl jspl_w_n493_0(.douta(w_dff_A_Hp7boeQl5_0),.doutb(w_n493_0[1]),.din(n493));
	jspl jspl_w_n494_0(.douta(w_dff_A_7mpuZtjD6_0),.doutb(w_n494_0[1]),.din(n494));
	jspl jspl_w_n502_0(.douta(w_dff_A_ia4ZqPFa5_0),.doutb(w_n502_0[1]),.din(w_dff_B_EaTX5xwa0_2));
	jspl jspl_w_n503_0(.douta(w_dff_A_JqcRgyAl8_0),.doutb(w_n503_0[1]),.din(n503));
	jspl jspl_w_n505_0(.douta(w_n505_0[0]),.doutb(w_dff_A_yB9qZISK9_1),.din(w_dff_B_XhCpM7G88_2));
	jspl3 jspl3_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.doutc(w_dff_A_SrxoqYpU5_2),.din(n507));
	jspl3 jspl3_w_n507_1(.douta(w_n507_1[0]),.doutb(w_n507_1[1]),.doutc(w_n507_1[2]),.din(w_n507_0[0]));
	jspl jspl_w_n508_0(.douta(w_n508_0[0]),.doutb(w_n508_0[1]),.din(n508));
	jspl jspl_w_n509_0(.douta(w_dff_A_TWgdoSAu6_0),.doutb(w_n509_0[1]),.din(n509));
	jspl jspl_w_n510_0(.douta(w_dff_A_flRhmxis9_0),.doutb(w_n510_0[1]),.din(n510));
	jspl jspl_w_n512_0(.douta(w_dff_A_FTpluSiU1_0),.doutb(w_n512_0[1]),.din(n512));
	jspl3 jspl3_w_n514_0(.douta(w_n514_0[0]),.doutb(w_dff_A_HM97nvu99_1),.doutc(w_n514_0[2]),.din(n514));
	jspl3 jspl3_w_n516_0(.douta(w_n516_0[0]),.doutb(w_dff_A_W7mZd8nP7_1),.doutc(w_n516_0[2]),.din(n516));
	jspl jspl_w_n518_0(.douta(w_n518_0[0]),.doutb(w_dff_A_5SfUobBg9_1),.din(n518));
	jspl jspl_w_n519_0(.douta(w_n519_0[0]),.doutb(w_n519_0[1]),.din(n519));
	jspl3 jspl3_w_n520_0(.douta(w_n520_0[0]),.doutb(w_dff_A_tEZvOvdz5_1),.doutc(w_dff_A_0y5Ha0Y56_2),.din(n520));
	jspl jspl_w_n522_0(.douta(w_n522_0[0]),.doutb(w_n522_0[1]),.din(n522));
	jspl3 jspl3_w_n523_0(.douta(w_n523_0[0]),.doutb(w_n523_0[1]),.doutc(w_n523_0[2]),.din(n523));
	jspl3 jspl3_w_n524_0(.douta(w_n524_0[0]),.doutb(w_n524_0[1]),.doutc(w_dff_A_8JjfnqII7_2),.din(n524));
	jspl3 jspl3_w_n524_1(.douta(w_n524_1[0]),.doutb(w_dff_A_qBGngdX23_1),.doutc(w_dff_A_tLCwrIOT5_2),.din(w_n524_0[0]));
	jspl jspl_w_n524_2(.douta(w_n524_2[0]),.doutb(w_n524_2[1]),.din(w_n524_0[1]));
	jspl3 jspl3_w_n525_0(.douta(w_n525_0[0]),.doutb(w_dff_A_kwZnzYGS7_1),.doutc(w_dff_A_fe8fo5r10_2),.din(n525));
	jspl jspl_w_n527_0(.douta(w_n527_0[0]),.doutb(w_n527_0[1]),.din(n527));
	jspl3 jspl3_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.doutc(w_n528_0[2]),.din(n528));
	jspl jspl_w_n528_1(.douta(w_n528_1[0]),.doutb(w_n528_1[1]),.din(w_n528_0[0]));
	jspl jspl_w_n529_0(.douta(w_dff_A_cHaWjaGn3_0),.doutb(w_n529_0[1]),.din(n529));
	jspl jspl_w_n530_0(.douta(w_dff_A_Khm9731N6_0),.doutb(w_n530_0[1]),.din(n530));
	jspl3 jspl3_w_n531_0(.douta(w_n531_0[0]),.doutb(w_dff_A_YqWCkFnU9_1),.doutc(w_dff_A_w0Fgt6lT0_2),.din(n531));
	jspl jspl_w_n533_0(.douta(w_n533_0[0]),.doutb(w_n533_0[1]),.din(n533));
	jspl3 jspl3_w_n534_0(.douta(w_n534_0[0]),.doutb(w_n534_0[1]),.doutc(w_n534_0[2]),.din(n534));
	jspl jspl_w_n534_1(.douta(w_n534_1[0]),.doutb(w_n534_1[1]),.din(w_n534_0[0]));
	jspl3 jspl3_w_n535_0(.douta(w_n535_0[0]),.doutb(w_dff_A_I8x6vdEz0_1),.doutc(w_n535_0[2]),.din(n535));
	jspl jspl_w_n535_1(.douta(w_dff_A_HBeBFwuV4_0),.doutb(w_n535_1[1]),.din(w_n535_0[0]));
	jspl jspl_w_n536_0(.douta(w_n536_0[0]),.doutb(w_n536_0[1]),.din(w_dff_B_LJ3KrJqL9_2));
	jspl jspl_w_n538_0(.douta(w_n538_0[0]),.doutb(w_n538_0[1]),.din(n538));
	jspl3 jspl3_w_n539_0(.douta(w_n539_0[0]),.doutb(w_n539_0[1]),.doutc(w_n539_0[2]),.din(n539));
	jspl jspl_w_n539_1(.douta(w_n539_1[0]),.doutb(w_n539_1[1]),.din(w_n539_0[0]));
	jspl3 jspl3_w_n540_0(.douta(w_dff_A_8WeyrEFP5_0),.doutb(w_dff_A_izyj3GnA6_1),.doutc(w_n540_0[2]),.din(n540));
	jspl jspl_w_n542_0(.douta(w_dff_A_Zh6HOU566_0),.doutb(w_n542_0[1]),.din(n542));
	jspl jspl_w_n549_0(.douta(w_n549_0[0]),.doutb(w_dff_A_g1ouEMrq9_1),.din(w_dff_B_Ekj3GVEX2_2));
	jspl jspl_w_n551_0(.douta(w_dff_A_Kx8Fz1th4_0),.doutb(w_n551_0[1]),.din(n551));
	jspl jspl_w_n552_0(.douta(w_dff_A_2eLJHofx6_0),.doutb(w_n552_0[1]),.din(n552));
	jspl jspl_w_n553_0(.douta(w_dff_A_vv5S50hW9_0),.doutb(w_n553_0[1]),.din(w_dff_B_B10ySFGf6_2));
	jspl3 jspl3_w_n554_0(.douta(w_n554_0[0]),.doutb(w_dff_A_95FZA3Zm5_1),.doutc(w_n554_0[2]),.din(n554));
	jspl3 jspl3_w_n556_0(.douta(w_n556_0[0]),.doutb(w_dff_A_QX6Uod323_1),.doutc(w_n556_0[2]),.din(n556));
	jspl jspl_w_n557_0(.douta(w_n557_0[0]),.doutb(w_n557_0[1]),.din(n557));
	jspl3 jspl3_w_n558_0(.douta(w_dff_A_hQattbZ39_0),.doutb(w_dff_A_H569RaTp6_1),.doutc(w_n558_0[2]),.din(n558));
	jspl jspl_w_n560_0(.douta(w_dff_A_QUz8ApJj9_0),.doutb(w_n560_0[1]),.din(n560));
	jspl3 jspl3_w_n562_0(.douta(w_n562_0[0]),.doutb(w_n562_0[1]),.doutc(w_n562_0[2]),.din(n562));
	jspl jspl_w_n563_0(.douta(w_n563_0[0]),.doutb(w_n563_0[1]),.din(w_dff_B_EfYlwM1z4_2));
	jspl3 jspl3_w_n564_0(.douta(w_dff_A_M2g0VMm52_0),.doutb(w_dff_A_pDl1u0AP0_1),.doutc(w_n564_0[2]),.din(n564));
	jspl3 jspl3_w_n565_0(.douta(w_n565_0[0]),.doutb(w_n565_0[1]),.doutc(w_n565_0[2]),.din(n565));
	jspl3 jspl3_w_n565_1(.douta(w_n565_1[0]),.doutb(w_n565_1[1]),.doutc(w_n565_1[2]),.din(w_n565_0[0]));
	jspl3 jspl3_w_n565_2(.douta(w_n565_2[0]),.doutb(w_n565_2[1]),.doutc(w_n565_2[2]),.din(w_n565_0[1]));
	jspl3 jspl3_w_n565_3(.douta(w_n565_3[0]),.doutb(w_n565_3[1]),.doutc(w_n565_3[2]),.din(w_n565_0[2]));
	jspl3 jspl3_w_n565_4(.douta(w_dff_A_eOGCc9MY9_0),.doutb(w_dff_A_xmqyPieu1_1),.doutc(w_n565_4[2]),.din(w_n565_1[0]));
	jspl3 jspl3_w_n565_5(.douta(w_n565_5[0]),.doutb(w_n565_5[1]),.doutc(w_n565_5[2]),.din(w_n565_1[1]));
	jspl3 jspl3_w_n565_6(.douta(w_n565_6[0]),.doutb(w_n565_6[1]),.doutc(w_n565_6[2]),.din(w_n565_1[2]));
	jspl3 jspl3_w_n565_7(.douta(w_n565_7[0]),.doutb(w_n565_7[1]),.doutc(w_n565_7[2]),.din(w_n565_2[0]));
	jspl3 jspl3_w_n565_8(.douta(w_n565_8[0]),.doutb(w_n565_8[1]),.doutc(w_n565_8[2]),.din(w_n565_2[1]));
	jspl3 jspl3_w_n565_9(.douta(w_n565_9[0]),.doutb(w_n565_9[1]),.doutc(w_n565_9[2]),.din(w_n565_2[2]));
	jspl jspl_w_n565_10(.douta(w_n565_10[0]),.doutb(w_n565_10[1]),.din(w_n565_3[0]));
	jspl3 jspl3_w_n567_0(.douta(w_n567_0[0]),.doutb(w_n567_0[1]),.doutc(w_n567_0[2]),.din(n567));
	jspl jspl_w_n567_1(.douta(w_n567_1[0]),.doutb(w_n567_1[1]),.din(w_n567_0[0]));
	jspl3 jspl3_w_n568_0(.douta(w_dff_A_VNCGnUvp7_0),.doutb(w_n568_0[1]),.doutc(w_dff_A_aV5KfnpY0_2),.din(n568));
	jspl3 jspl3_w_n569_0(.douta(w_n569_0[0]),.doutb(w_n569_0[1]),.doutc(w_n569_0[2]),.din(w_dff_B_PQGBc40z6_3));
	jspl jspl_w_n570_0(.douta(w_n570_0[0]),.doutb(w_n570_0[1]),.din(n570));
	jspl3 jspl3_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.doutc(w_dff_A_eyU1szws7_2),.din(n572));
	jspl jspl_w_n572_1(.douta(w_n572_1[0]),.doutb(w_n572_1[1]),.din(w_n572_0[0]));
	jspl3 jspl3_w_n573_0(.douta(w_n573_0[0]),.doutb(w_n573_0[1]),.doutc(w_dff_A_Gqf84gAp9_2),.din(n573));
	jspl jspl_w_n573_1(.douta(w_n573_1[0]),.doutb(w_n573_1[1]),.din(w_n573_0[0]));
	jspl jspl_w_n574_0(.douta(w_n574_0[0]),.doutb(w_n574_0[1]),.din(w_dff_B_RLctYm3i2_2));
	jspl jspl_w_n575_0(.douta(w_n575_0[0]),.doutb(w_n575_0[1]),.din(n575));
	jspl3 jspl3_w_n577_0(.douta(w_n577_0[0]),.doutb(w_n577_0[1]),.doutc(w_n577_0[2]),.din(n577));
	jspl3 jspl3_w_n578_0(.douta(w_n578_0[0]),.doutb(w_dff_A_6gxuXLXQ4_1),.doutc(w_dff_A_OjqN8yyk2_2),.din(n578));
	jspl jspl_w_n578_1(.douta(w_dff_A_9gZkPiu00_0),.doutb(w_n578_1[1]),.din(w_n578_0[0]));
	jspl3 jspl3_w_n579_0(.douta(w_n579_0[0]),.doutb(w_n579_0[1]),.doutc(w_n579_0[2]),.din(n579));
	jspl jspl_w_n580_0(.douta(w_n580_0[0]),.doutb(w_n580_0[1]),.din(w_dff_B_4m3qZeri9_2));
	jspl jspl_w_n581_0(.douta(w_n581_0[0]),.doutb(w_n581_0[1]),.din(n581));
	jspl3 jspl3_w_n583_0(.douta(w_n583_0[0]),.doutb(w_n583_0[1]),.doutc(w_n583_0[2]),.din(n583));
	jspl jspl_w_n583_1(.douta(w_n583_1[0]),.doutb(w_n583_1[1]),.din(w_n583_0[0]));
	jspl3 jspl3_w_n584_0(.douta(w_n584_0[0]),.doutb(w_n584_0[1]),.doutc(w_n584_0[2]),.din(n584));
	jspl jspl_w_n585_0(.douta(w_n585_0[0]),.doutb(w_n585_0[1]),.din(w_dff_B_UbAXsghV7_2));
	jspl jspl_w_n586_0(.douta(w_n586_0[0]),.doutb(w_n586_0[1]),.din(n586));
	jspl3 jspl3_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.doutc(w_n588_0[2]),.din(n588));
	jspl jspl_w_n588_1(.douta(w_n588_1[0]),.doutb(w_n588_1[1]),.din(w_n588_0[0]));
	jspl3 jspl3_w_n589_0(.douta(w_n589_0[0]),.doutb(w_dff_A_uzIPxl4Y3_1),.doutc(w_n589_0[2]),.din(n589));
	jspl jspl_w_n589_1(.douta(w_n589_1[0]),.doutb(w_n589_1[1]),.din(w_n589_0[0]));
	jspl jspl_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.din(n591));
	jspl jspl_w_n592_0(.douta(w_dff_A_LLjFKsmq6_0),.doutb(w_n592_0[1]),.din(n592));
	jspl jspl_w_n599_0(.douta(w_dff_A_01lbMFDm6_0),.doutb(w_n599_0[1]),.din(n599));
	jspl jspl_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.din(n605));
	jspl3 jspl3_w_n606_0(.douta(w_n606_0[0]),.doutb(w_n606_0[1]),.doutc(w_n606_0[2]),.din(n606));
	jspl3 jspl3_w_n606_1(.douta(w_dff_A_A9i6iMN36_0),.doutb(w_dff_A_yf1K9M6n8_1),.doutc(w_n606_1[2]),.din(w_n606_0[0]));
	jspl jspl_w_n607_0(.douta(w_n607_0[0]),.doutb(w_n607_0[1]),.din(n607));
	jspl3 jspl3_w_n608_0(.douta(w_dff_A_L8Ushhu59_0),.doutb(w_n608_0[1]),.doutc(w_n608_0[2]),.din(n608));
	jspl jspl_w_n610_0(.douta(w_dff_A_xXkZjEFp7_0),.doutb(w_n610_0[1]),.din(n610));
	jspl jspl_w_n612_0(.douta(w_n612_0[0]),.doutb(w_n612_0[1]),.din(n612));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_dff_A_NpEFCCjl2_1),.doutc(w_n613_0[2]),.din(n613));
	jspl3 jspl3_w_n615_0(.douta(w_n615_0[0]),.doutb(w_n615_0[1]),.doutc(w_n615_0[2]),.din(n615));
	jspl jspl_w_n615_1(.douta(w_dff_A_FfUoooxR6_0),.doutb(w_n615_1[1]),.din(w_n615_0[0]));
	jspl jspl_w_n617_0(.douta(w_n617_0[0]),.doutb(w_dff_A_blJgktoG6_1),.din(n617));
	jspl3 jspl3_w_n618_0(.douta(w_n618_0[0]),.doutb(w_n618_0[1]),.doutc(w_n618_0[2]),.din(n618));
	jspl jspl_w_n619_0(.douta(w_n619_0[0]),.doutb(w_n619_0[1]),.din(w_dff_B_dndzmJYW5_2));
	jspl jspl_w_n620_0(.douta(w_dff_A_CCugBIQk7_0),.doutb(w_n620_0[1]),.din(n620));
	jspl3 jspl3_w_n621_0(.douta(w_n621_0[0]),.doutb(w_n621_0[1]),.doutc(w_n621_0[2]),.din(n621));
	jspl3 jspl3_w_n622_0(.douta(w_n622_0[0]),.doutb(w_n622_0[1]),.doutc(w_dff_A_xLohmLmE5_2),.din(n622));
	jspl jspl_w_n622_1(.douta(w_n622_1[0]),.doutb(w_n622_1[1]),.din(w_n622_0[0]));
	jspl3 jspl3_w_n623_0(.douta(w_n623_0[0]),.doutb(w_dff_A_SQQVOfIU1_1),.doutc(w_dff_A_339cPwC63_2),.din(n623));
	jspl jspl_w_n624_0(.douta(w_dff_A_7oRzPrHY1_0),.doutb(w_n624_0[1]),.din(n624));
	jspl3 jspl3_w_n625_0(.douta(w_n625_0[0]),.doutb(w_n625_0[1]),.doutc(w_n625_0[2]),.din(n625));
	jspl jspl_w_n626_0(.douta(w_dff_A_bwotvWOV0_0),.doutb(w_n626_0[1]),.din(n626));
	jspl jspl_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.din(n627));
	jspl jspl_w_n628_0(.douta(w_n628_0[0]),.doutb(w_n628_0[1]),.din(w_dff_B_rDypx3QF1_2));
	jspl jspl_w_n629_0(.douta(w_dff_A_a1W6TsAm6_0),.doutb(w_n629_0[1]),.din(n629));
	jspl3 jspl3_w_n630_0(.douta(w_n630_0[0]),.doutb(w_n630_0[1]),.doutc(w_n630_0[2]),.din(n630));
	jspl jspl_w_n631_0(.douta(w_n631_0[0]),.doutb(w_n631_0[1]),.din(n631));
	jspl jspl_w_n632_0(.douta(w_n632_0[0]),.doutb(w_n632_0[1]),.din(w_dff_B_KBlbIcD88_2));
	jspl jspl_w_n633_0(.douta(w_dff_A_4kuSY1976_0),.doutb(w_n633_0[1]),.din(n633));
	jspl3 jspl3_w_n634_0(.douta(w_n634_0[0]),.doutb(w_n634_0[1]),.doutc(w_n634_0[2]),.din(n634));
	jspl3 jspl3_w_n635_0(.douta(w_dff_A_97LXNt6R5_0),.doutb(w_n635_0[1]),.doutc(w_n635_0[2]),.din(n635));
	jspl jspl_w_n637_0(.douta(w_dff_A_RgGa0dKo8_0),.doutb(w_n637_0[1]),.din(n637));
	jspl jspl_w_n642_0(.douta(w_dff_A_5Zp1Rz6K0_0),.doutb(w_n642_0[1]),.din(n642));
	jspl jspl_w_n643_0(.douta(w_dff_A_Ai9LT4dN0_0),.doutb(w_n643_0[1]),.din(w_dff_B_IqbrtGa19_2));
	jspl3 jspl3_w_n645_0(.douta(w_dff_A_uEeCJ1Kd7_0),.doutb(w_dff_A_vbxwZFMd3_1),.doutc(w_n645_0[2]),.din(n645));
	jspl jspl_w_n647_0(.douta(w_n647_0[0]),.doutb(w_n647_0[1]),.din(n647));
	jspl3 jspl3_w_n648_0(.douta(w_n648_0[0]),.doutb(w_dff_A_5EVaKySu6_1),.doutc(w_n648_0[2]),.din(n648));
	jspl jspl_w_n649_0(.douta(w_n649_0[0]),.doutb(w_n649_0[1]),.din(n649));
	jspl jspl_w_n650_0(.douta(w_n650_0[0]),.doutb(w_n650_0[1]),.din(n650));
	jspl jspl_w_n652_0(.douta(w_n652_0[0]),.doutb(w_n652_0[1]),.din(n652));
	jspl3 jspl3_w_n653_0(.douta(w_n653_0[0]),.doutb(w_dff_A_KJrEFhzp3_1),.doutc(w_n653_0[2]),.din(n653));
	jspl jspl_w_n653_1(.douta(w_dff_A_b79Vmeps7_0),.doutb(w_n653_1[1]),.din(w_n653_0[0]));
	jspl jspl_w_n656_0(.douta(w_n656_0[0]),.doutb(w_dff_A_KeIE0M3X6_1),.din(n656));
	jspl3 jspl3_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.doutc(w_n657_0[2]),.din(n657));
	jspl jspl_w_n657_1(.douta(w_n657_1[0]),.doutb(w_n657_1[1]),.din(w_n657_0[0]));
	jspl3 jspl3_w_n658_0(.douta(w_n658_0[0]),.doutb(w_n658_0[1]),.doutc(w_n658_0[2]),.din(w_dff_B_FnI5fl3B8_3));
	jspl jspl_w_n659_0(.douta(w_n659_0[0]),.doutb(w_n659_0[1]),.din(n659));
	jspl3 jspl3_w_n660_0(.douta(w_n660_0[0]),.doutb(w_n660_0[1]),.doutc(w_n660_0[2]),.din(n660));
	jspl jspl_w_n660_1(.douta(w_n660_1[0]),.doutb(w_n660_1[1]),.din(w_n660_0[0]));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_dff_A_jxNuVVNz2_1),.din(n661));
	jspl3 jspl3_w_n662_0(.douta(w_n662_0[0]),.doutb(w_n662_0[1]),.doutc(w_n662_0[2]),.din(w_dff_B_85BJkmhI0_3));
	jspl jspl_w_n663_0(.douta(w_n663_0[0]),.doutb(w_n663_0[1]),.din(n663));
	jspl3 jspl3_w_n664_0(.douta(w_n664_0[0]),.doutb(w_n664_0[1]),.doutc(w_n664_0[2]),.din(n664));
	jspl jspl_w_n664_1(.douta(w_n664_1[0]),.doutb(w_n664_1[1]),.din(w_n664_0[0]));
	jspl3 jspl3_w_n665_0(.douta(w_n665_0[0]),.doutb(w_n665_0[1]),.doutc(w_n665_0[2]),.din(n665));
	jspl jspl_w_n666_0(.douta(w_n666_0[0]),.doutb(w_n666_0[1]),.din(w_dff_B_wObdoSbL6_2));
	jspl jspl_w_n667_0(.douta(w_dff_A_geoSaktb6_0),.doutb(w_n667_0[1]),.din(n667));
	jspl3 jspl3_w_n668_0(.douta(w_n668_0[0]),.doutb(w_n668_0[1]),.doutc(w_n668_0[2]),.din(n668));
	jspl3 jspl3_w_n669_0(.douta(w_n669_0[0]),.doutb(w_n669_0[1]),.doutc(w_n669_0[2]),.din(n669));
	jspl jspl_w_n671_0(.douta(w_n671_0[0]),.doutb(w_n671_0[1]),.din(w_dff_B_Eyc3M63f7_2));
	jspl jspl_w_n672_0(.douta(w_dff_A_h8xI2N846_0),.doutb(w_n672_0[1]),.din(n672));
	jspl3 jspl3_w_n673_0(.douta(w_n673_0[0]),.doutb(w_n673_0[1]),.doutc(w_n673_0[2]),.din(n673));
	jspl3 jspl3_w_n674_0(.douta(w_n674_0[0]),.doutb(w_dff_A_USr6oUuH6_1),.doutc(w_n674_0[2]),.din(n674));
	jspl jspl_w_n674_1(.douta(w_dff_A_DsUS2yNh5_0),.doutb(w_n674_1[1]),.din(w_n674_0[0]));
	jspl3 jspl3_w_n675_0(.douta(w_n675_0[0]),.doutb(w_n675_0[1]),.doutc(w_n675_0[2]),.din(w_dff_B_GUFRaQMM5_3));
	jspl jspl_w_n676_0(.douta(w_n676_0[0]),.doutb(w_n676_0[1]),.din(n676));
	jspl3 jspl3_w_n677_0(.douta(w_n677_0[0]),.doutb(w_n677_0[1]),.doutc(w_n677_0[2]),.din(n677));
	jspl3 jspl3_w_n678_0(.douta(w_dff_A_TO1bcOxd6_0),.doutb(w_dff_A_KLSNYSLk1_1),.doutc(w_n678_0[2]),.din(n678));
	jspl3 jspl3_w_n679_0(.douta(w_n679_0[0]),.doutb(w_dff_A_rbPYaqof3_1),.doutc(w_dff_A_FRanbqnu6_2),.din(n679));
	jspl jspl_w_n679_1(.douta(w_n679_1[0]),.doutb(w_n679_1[1]),.din(w_n679_0[0]));
	jspl jspl_w_n680_0(.douta(w_dff_A_Daa9saj76_0),.doutb(w_n680_0[1]),.din(n680));
	jspl jspl_w_n683_0(.douta(w_n683_0[0]),.doutb(w_n683_0[1]),.din(n683));
	jspl jspl_w_n686_0(.douta(w_dff_A_JtQI1AOW4_0),.doutb(w_n686_0[1]),.din(n686));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_dff_A_alPEdqvK7_1),.din(w_dff_B_JDTa9cxO0_2));
	jspl jspl_w_n690_0(.douta(w_n690_0[0]),.doutb(w_n690_0[1]),.din(n690));
	jspl jspl_w_n692_0(.douta(w_n692_0[0]),.doutb(w_dff_A_GalQl23S9_1),.din(n692));
	jspl jspl_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.din(n693));
	jspl3 jspl3_w_n697_0(.douta(w_dff_A_hEchCG9b8_0),.doutb(w_dff_A_uyp60RjA7_1),.doutc(w_n697_0[2]),.din(n697));
	jspl3 jspl3_w_n699_0(.douta(w_n699_0[0]),.doutb(w_n699_0[1]),.doutc(w_n699_0[2]),.din(n699));
	jspl jspl_w_n699_1(.douta(w_n699_1[0]),.doutb(w_n699_1[1]),.din(w_n699_0[0]));
	jspl3 jspl3_w_n701_0(.douta(w_n701_0[0]),.doutb(w_n701_0[1]),.doutc(w_n701_0[2]),.din(n701));
	jspl jspl_w_n701_1(.douta(w_n701_1[0]),.doutb(w_n701_1[1]),.din(w_n701_0[0]));
	jspl jspl_w_n703_0(.douta(w_n703_0[0]),.doutb(w_n703_0[1]),.din(n703));
	jspl jspl_w_n704_0(.douta(w_dff_A_BWxM5W4l6_0),.doutb(w_n704_0[1]),.din(n704));
	jspl jspl_w_n705_0(.douta(w_n705_0[0]),.doutb(w_n705_0[1]),.din(n705));
	jspl3 jspl3_w_n707_0(.douta(w_n707_0[0]),.doutb(w_dff_A_CQCZnukW9_1),.doutc(w_n707_0[2]),.din(n707));
	jspl jspl_w_n708_0(.douta(w_n708_0[0]),.doutb(w_dff_A_sIlKmTIk2_1),.din(n708));
	jspl3 jspl3_w_n709_0(.douta(w_n709_0[0]),.doutb(w_n709_0[1]),.doutc(w_n709_0[2]),.din(n709));
	jspl jspl_w_n709_1(.douta(w_n709_1[0]),.doutb(w_n709_1[1]),.din(w_n709_0[0]));
	jspl jspl_w_n710_0(.douta(w_n710_0[0]),.doutb(w_n710_0[1]),.din(n710));
	jspl jspl_w_n711_0(.douta(w_n711_0[0]),.doutb(w_n711_0[1]),.din(n711));
	jspl jspl_w_n712_0(.douta(w_dff_A_hFyNf2gp7_0),.doutb(w_n712_0[1]),.din(n712));
	jspl3 jspl3_w_n713_0(.douta(w_n713_0[0]),.doutb(w_n713_0[1]),.doutc(w_n713_0[2]),.din(w_dff_B_EQWtMFSW0_3));
	jspl jspl_w_n713_1(.douta(w_n713_1[0]),.doutb(w_n713_1[1]),.din(w_n713_0[0]));
	jspl jspl_w_n714_0(.douta(w_n714_0[0]),.doutb(w_n714_0[1]),.din(n714));
	jspl3 jspl3_w_n715_0(.douta(w_dff_A_QFVvSBXs1_0),.doutb(w_dff_A_ovTq2xU49_1),.doutc(w_n715_0[2]),.din(n715));
	jspl3 jspl3_w_n716_0(.douta(w_n716_0[0]),.doutb(w_n716_0[1]),.doutc(w_n716_0[2]),.din(n716));
	jspl jspl_w_n716_1(.douta(w_n716_1[0]),.doutb(w_n716_1[1]),.din(w_n716_0[0]));
	jspl3 jspl3_w_n720_0(.douta(w_n720_0[0]),.doutb(w_n720_0[1]),.doutc(w_n720_0[2]),.din(w_dff_B_ZKPdG3yj8_3));
	jspl jspl_w_n720_1(.douta(w_n720_1[0]),.doutb(w_n720_1[1]),.din(w_n720_0[0]));
	jspl3 jspl3_w_n723_0(.douta(w_n723_0[0]),.doutb(w_n723_0[1]),.doutc(w_n723_0[2]),.din(n723));
	jspl3 jspl3_w_n727_0(.douta(w_dff_A_fbjRGt6H7_0),.doutb(w_n727_0[1]),.doutc(w_n727_0[2]),.din(n727));
	jspl jspl_w_n728_0(.douta(w_n728_0[0]),.doutb(w_dff_A_x53jfDaD6_1),.din(w_dff_B_gdK7QGUf4_2));
	jspl3 jspl3_w_n730_0(.douta(w_n730_0[0]),.doutb(w_n730_0[1]),.doutc(w_n730_0[2]),.din(n730));
	jspl3 jspl3_w_n734_0(.douta(w_n734_0[0]),.doutb(w_n734_0[1]),.doutc(w_n734_0[2]),.din(n734));
	jspl jspl_w_n735_0(.douta(w_n735_0[0]),.doutb(w_dff_A_yzHYW8jW8_1),.din(w_dff_B_NqZ7nwu76_2));
	jspl3 jspl3_w_n737_0(.douta(w_dff_A_tL4pS8RP3_0),.doutb(w_n737_0[1]),.doutc(w_n737_0[2]),.din(n737));
	jspl3 jspl3_w_n741_0(.douta(w_n741_0[0]),.doutb(w_n741_0[1]),.doutc(w_n741_0[2]),.din(n741));
	jspl jspl_w_n742_0(.douta(w_n742_0[0]),.doutb(w_dff_A_ekM6GQ1p6_1),.din(n742));
	jspl3 jspl3_w_n744_0(.douta(w_n744_0[0]),.doutb(w_n744_0[1]),.doutc(w_n744_0[2]),.din(n744));
	jspl3 jspl3_w_n748_0(.douta(w_n748_0[0]),.doutb(w_n748_0[1]),.doutc(w_n748_0[2]),.din(n748));
	jspl jspl_w_n751_0(.douta(w_dff_A_qkOoyJRf5_0),.doutb(w_n751_0[1]),.din(n751));
	jspl jspl_w_n752_0(.douta(w_n752_0[0]),.doutb(w_n752_0[1]),.din(n752));
	jspl3 jspl3_w_n754_0(.douta(w_n754_0[0]),.doutb(w_n754_0[1]),.doutc(w_n754_0[2]),.din(n754));
	jspl3 jspl3_w_n758_0(.douta(w_n758_0[0]),.doutb(w_n758_0[1]),.doutc(w_n758_0[2]),.din(n758));
	jspl jspl_w_n759_0(.douta(w_n759_0[0]),.doutb(w_n759_0[1]),.din(n759));
	jspl jspl_w_n764_0(.douta(w_n764_0[0]),.doutb(w_n764_0[1]),.din(n764));
	jspl jspl_w_n765_0(.douta(w_n765_0[0]),.doutb(w_n765_0[1]),.din(n765));
	jspl jspl_w_n782_0(.douta(w_n782_0[0]),.doutb(w_dff_A_Mf0742Hd8_1),.din(n782));
	jspl3 jspl3_w_n784_0(.douta(w_n784_0[0]),.doutb(w_n784_0[1]),.doutc(w_n784_0[2]),.din(n784));
	jspl3 jspl3_w_n787_0(.douta(w_n787_0[0]),.doutb(w_n787_0[1]),.doutc(w_n787_0[2]),.din(n787));
	jspl3 jspl3_w_n790_0(.douta(w_n790_0[0]),.doutb(w_n790_0[1]),.doutc(w_n790_0[2]),.din(n790));
	jspl jspl_w_n790_1(.douta(w_n790_1[0]),.doutb(w_n790_1[1]),.din(w_n790_0[0]));
	jspl3 jspl3_w_n793_0(.douta(w_n793_0[0]),.doutb(w_n793_0[1]),.doutc(w_n793_0[2]),.din(n793));
	jspl jspl_w_n793_1(.douta(w_n793_1[0]),.doutb(w_n793_1[1]),.din(w_n793_0[0]));
	jspl jspl_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.din(n795));
	jspl3 jspl3_w_n797_0(.douta(w_n797_0[0]),.doutb(w_n797_0[1]),.doutc(w_n797_0[2]),.din(n797));
	jspl jspl_w_n797_1(.douta(w_n797_1[0]),.doutb(w_n797_1[1]),.din(w_n797_0[0]));
	jspl3 jspl3_w_n801_0(.douta(w_n801_0[0]),.doutb(w_n801_0[1]),.doutc(w_n801_0[2]),.din(n801));
	jspl jspl_w_n801_1(.douta(w_n801_1[0]),.doutb(w_n801_1[1]),.din(w_n801_0[0]));
	jspl jspl_w_n802_0(.douta(w_n802_0[0]),.doutb(w_n802_0[1]),.din(n802));
	jspl3 jspl3_w_n804_0(.douta(w_n804_0[0]),.doutb(w_n804_0[1]),.doutc(w_n804_0[2]),.din(n804));
	jspl3 jspl3_w_n807_0(.douta(w_n807_0[0]),.doutb(w_n807_0[1]),.doutc(w_n807_0[2]),.din(n807));
	jspl3 jspl3_w_n810_0(.douta(w_dff_A_aZDu4bpW2_0),.doutb(w_n810_0[1]),.doutc(w_dff_A_sbM22p8l0_2),.din(w_dff_B_7O3vY0Tl6_3));
	jspl3 jspl3_w_n812_0(.douta(w_n812_0[0]),.doutb(w_n812_0[1]),.doutc(w_n812_0[2]),.din(n812));
	jspl3 jspl3_w_n816_0(.douta(w_n816_0[0]),.doutb(w_n816_0[1]),.doutc(w_n816_0[2]),.din(n816));
	jspl jspl_w_n817_0(.douta(w_n817_0[0]),.doutb(w_n817_0[1]),.din(n817));
	jspl3 jspl3_w_n819_0(.douta(w_n819_0[0]),.doutb(w_n819_0[1]),.doutc(w_n819_0[2]),.din(n819));
	jspl3 jspl3_w_n823_0(.douta(w_n823_0[0]),.doutb(w_n823_0[1]),.doutc(w_n823_0[2]),.din(n823));
	jspl jspl_w_n824_0(.douta(w_dff_A_kvQeBA0D2_0),.doutb(w_n824_0[1]),.din(n824));
	jspl3 jspl3_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.doutc(w_n827_0[2]),.din(n827));
	jspl3 jspl3_w_n831_0(.douta(w_n831_0[0]),.doutb(w_n831_0[1]),.doutc(w_n831_0[2]),.din(n831));
	jspl jspl_w_n832_0(.douta(w_n832_0[0]),.doutb(w_n832_0[1]),.din(n832));
	jspl jspl_w_n834_0(.douta(w_n834_0[0]),.doutb(w_n834_0[1]),.din(n834));
	jspl jspl_w_n838_0(.douta(w_n838_0[0]),.doutb(w_n838_0[1]),.din(n838));
	jspl3 jspl3_w_n843_0(.douta(w_n843_0[0]),.doutb(w_n843_0[1]),.doutc(w_n843_0[2]),.din(n843));
	jspl3 jspl3_w_n847_0(.douta(w_n847_0[0]),.doutb(w_n847_0[1]),.doutc(w_n847_0[2]),.din(n847));
	jspl jspl_w_n848_0(.douta(w_dff_A_wUpRfK0p1_0),.doutb(w_n848_0[1]),.din(n848));
	jspl3 jspl3_w_n851_0(.douta(w_dff_A_CwlY1HgX1_0),.doutb(w_n851_0[1]),.doutc(w_n851_0[2]),.din(n851));
	jspl3 jspl3_w_n855_0(.douta(w_dff_A_CC1cSYvL9_0),.doutb(w_n855_0[1]),.doutc(w_n855_0[2]),.din(n855));
	jspl jspl_w_n856_0(.douta(w_n856_0[0]),.doutb(w_dff_A_uObGZouh4_1),.din(n856));
	jspl3 jspl3_w_n858_0(.douta(w_n858_0[0]),.doutb(w_n858_0[1]),.doutc(w_dff_A_rALwFiav9_2),.din(n858));
	jspl jspl_w_n859_0(.douta(w_n859_0[0]),.doutb(w_n859_0[1]),.din(n859));
	jspl jspl_w_n864_0(.douta(w_dff_A_j8FtofYP3_0),.doutb(w_n864_0[1]),.din(n864));
	jspl jspl_w_n865_0(.douta(w_n865_0[0]),.doutb(w_dff_A_lYcNZSyi0_1),.din(n865));
	jspl3 jspl3_w_n869_0(.douta(w_n869_0[0]),.doutb(w_n869_0[1]),.doutc(w_n869_0[2]),.din(n869));
	jspl3 jspl3_w_n873_0(.douta(w_n873_0[0]),.doutb(w_dff_A_kZe7phSE5_1),.doutc(w_dff_A_q50Fv1v73_2),.din(n873));
	jspl jspl_w_n874_0(.douta(w_dff_A_g9V4GvzL7_0),.doutb(w_n874_0[1]),.din(n874));
	jspl3 jspl3_w_n878_0(.douta(w_n878_0[0]),.doutb(w_n878_0[1]),.doutc(w_n878_0[2]),.din(n878));
	jspl3 jspl3_w_n882_0(.douta(w_n882_0[0]),.doutb(w_dff_A_kfTwIkQA1_1),.doutc(w_dff_A_wlzDAiYg7_2),.din(n882));
	jspl jspl_w_n885_0(.douta(w_n885_0[0]),.doutb(w_n885_0[1]),.din(n885));
	jspl jspl_w_n887_0(.douta(w_n887_0[0]),.doutb(w_dff_A_oK3vFRv77_1),.din(n887));
	jspl jspl_w_n889_0(.douta(w_n889_0[0]),.doutb(w_n889_0[1]),.din(n889));
	jspl3 jspl3_w_n891_0(.douta(w_n891_0[0]),.doutb(w_dff_A_cGZBiJwI7_1),.doutc(w_n891_0[2]),.din(n891));
	jspl jspl_w_n891_1(.douta(w_n891_1[0]),.doutb(w_n891_1[1]),.din(w_n891_0[0]));
	jspl3 jspl3_w_n895_0(.douta(w_n895_0[0]),.doutb(w_n895_0[1]),.doutc(w_n895_0[2]),.din(n895));
	jspl jspl_w_n895_1(.douta(w_n895_1[0]),.doutb(w_n895_1[1]),.din(w_n895_0[0]));
	jspl jspl_w_n896_0(.douta(w_n896_0[0]),.doutb(w_n896_0[1]),.din(w_dff_B_qVKgIB5E4_2));
	jspl3 jspl3_w_n899_0(.douta(w_n899_0[0]),.doutb(w_n899_0[1]),.doutc(w_n899_0[2]),.din(n899));
	jspl3 jspl3_w_n902_0(.douta(w_n902_0[0]),.doutb(w_dff_A_ABytohFn0_1),.doutc(w_dff_A_Voxo0vv56_2),.din(n902));
	jspl3 jspl3_w_n905_0(.douta(w_dff_A_DrbNfpRo1_0),.doutb(w_n905_0[1]),.doutc(w_n905_0[2]),.din(w_dff_B_INOoEPE86_3));
	jspl3 jspl3_w_n908_0(.douta(w_n908_0[0]),.doutb(w_n908_0[1]),.doutc(w_n908_0[2]),.din(n908));
	jspl3 jspl3_w_n912_0(.douta(w_n912_0[0]),.doutb(w_n912_0[1]),.doutc(w_n912_0[2]),.din(w_dff_B_iLWJF1Hp3_3));
	jspl jspl_w_n913_0(.douta(w_n913_0[0]),.doutb(w_n913_0[1]),.din(n913));
	jspl3 jspl3_w_n916_0(.douta(w_n916_0[0]),.doutb(w_n916_0[1]),.doutc(w_n916_0[2]),.din(n916));
	jspl3 jspl3_w_n920_0(.douta(w_n920_0[0]),.doutb(w_dff_A_ENCyuXag9_1),.doutc(w_dff_A_2yNquiOy5_2),.din(n920));
	jspl jspl_w_n921_0(.douta(w_n921_0[0]),.doutb(w_n921_0[1]),.din(n921));
	jspl jspl_w_n923_0(.douta(w_n923_0[0]),.doutb(w_n923_0[1]),.din(n923));
	jspl3 jspl3_w_n927_0(.douta(w_n927_0[0]),.doutb(w_n927_0[1]),.doutc(w_n927_0[2]),.din(n927));
	jspl3 jspl3_w_n931_0(.douta(w_n931_0[0]),.doutb(w_dff_A_OL2RzQCe5_1),.doutc(w_dff_A_GNJJtZnm1_2),.din(n931));
	jspl jspl_w_n932_0(.douta(w_n932_0[0]),.doutb(w_dff_A_ze6hIAz33_1),.din(n932));
	jspl jspl_w_n935_0(.douta(w_n935_0[0]),.doutb(w_n935_0[1]),.din(n935));
	jspl jspl_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.din(n937));
	jspl jspl_w_n939_0(.douta(w_dff_A_7pUNrHii4_0),.doutb(w_n939_0[1]),.din(n939));
	jspl3 jspl3_w_n945_0(.douta(w_n945_0[0]),.doutb(w_n945_0[1]),.doutc(w_n945_0[2]),.din(n945));
	jspl jspl_w_n945_1(.douta(w_n945_1[0]),.doutb(w_n945_1[1]),.din(w_n945_0[0]));
	jspl3 jspl3_w_n948_0(.douta(w_dff_A_SZuNFr1P2_0),.doutb(w_n948_0[1]),.doutc(w_dff_A_4oRPwfXE4_2),.din(n948));
	jspl jspl_w_n948_1(.douta(w_n948_1[0]),.doutb(w_n948_1[1]),.din(w_n948_0[0]));
	jspl jspl_w_n950_0(.douta(w_n950_0[0]),.doutb(w_n950_0[1]),.din(n950));
	jspl jspl_w_n952_0(.douta(w_n952_0[0]),.doutb(w_n952_0[1]),.din(n952));
	jspl jspl_w_n957_0(.douta(w_n957_0[0]),.doutb(w_n957_0[1]),.din(n957));
	jspl jspl_w_n972_0(.douta(w_dff_A_zhxyA46L1_0),.doutb(w_n972_0[1]),.din(w_dff_B_sHtAJ7Vc2_2));
	jspl jspl_w_n981_0(.douta(w_dff_A_7YvRhIar6_0),.doutb(w_n981_0[1]),.din(n981));
	jspl jspl_w_n987_0(.douta(w_n987_0[0]),.doutb(w_n987_0[1]),.din(n987));
	jspl3 jspl3_w_n988_0(.douta(w_n988_0[0]),.doutb(w_n988_0[1]),.doutc(w_n988_0[2]),.din(n988));
	jspl3 jspl3_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.doutc(w_n992_0[2]),.din(n992));
	jspl jspl_w_n993_0(.douta(w_n993_0[0]),.doutb(w_dff_A_14yKmCqw2_1),.din(n993));
	jspl jspl_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.din(n994));
	jspl3 jspl3_w_n995_0(.douta(w_n995_0[0]),.doutb(w_n995_0[1]),.doutc(w_n995_0[2]),.din(n995));
	jspl3 jspl3_w_n999_0(.douta(w_n999_0[0]),.doutb(w_n999_0[1]),.doutc(w_n999_0[2]),.din(n999));
	jspl jspl_w_n1000_0(.douta(w_n1000_0[0]),.doutb(w_n1000_0[1]),.din(n1000));
	jspl jspl_w_n1003_0(.douta(w_dff_A_pYjNPTOh3_0),.doutb(w_n1003_0[1]),.din(n1003));
	jspl jspl_w_n1007_0(.douta(w_n1007_0[0]),.doutb(w_n1007_0[1]),.din(n1007));
	jspl jspl_w_n1008_0(.douta(w_n1008_0[0]),.doutb(w_n1008_0[1]),.din(n1008));
	jspl3 jspl3_w_n1009_0(.douta(w_n1009_0[0]),.doutb(w_n1009_0[1]),.doutc(w_n1009_0[2]),.din(n1009));
	jspl jspl_w_n1009_1(.douta(w_n1009_1[0]),.doutb(w_n1009_1[1]),.din(w_n1009_0[0]));
	jspl3 jspl3_w_n1013_0(.douta(w_n1013_0[0]),.doutb(w_n1013_0[1]),.doutc(w_n1013_0[2]),.din(n1013));
	jspl jspl_w_n1013_1(.douta(w_n1013_1[0]),.doutb(w_n1013_1[1]),.din(w_n1013_0[0]));
	jspl jspl_w_n1014_0(.douta(w_n1014_0[0]),.doutb(w_n1014_0[1]),.din(n1014));
	jspl jspl_w_n1015_0(.douta(w_n1015_0[0]),.doutb(w_n1015_0[1]),.din(n1015));
	jspl3 jspl3_w_n1016_0(.douta(w_n1016_0[0]),.doutb(w_n1016_0[1]),.doutc(w_n1016_0[2]),.din(n1016));
	jspl3 jspl3_w_n1019_0(.douta(w_n1019_0[0]),.doutb(w_n1019_0[1]),.doutc(w_n1019_0[2]),.din(n1019));
	jspl jspl_w_n1022_0(.douta(w_n1022_0[0]),.doutb(w_dff_A_ReZ75tPd8_1),.din(w_dff_B_tB2GeuHj0_2));
	jspl jspl_w_n1033_0(.douta(w_n1033_0[0]),.doutb(w_n1033_0[1]),.din(n1033));
	jspl jspl_w_n1044_0(.douta(w_dff_A_rwP99a5q0_0),.doutb(w_n1044_0[1]),.din(w_dff_B_kXm7rX3S9_2));
	jspl3 jspl3_w_n1061_0(.douta(w_dff_A_DPI265385_0),.doutb(w_n1061_0[1]),.doutc(w_n1061_0[2]),.din(n1061));
	jspl jspl_w_n1062_0(.douta(w_n1062_0[0]),.doutb(w_n1062_0[1]),.din(n1062));
	jspl3 jspl3_w_n1066_0(.douta(w_dff_A_Uh6msUUb7_0),.doutb(w_n1066_0[1]),.doutc(w_n1066_0[2]),.din(n1066));
	jspl jspl_w_n1068_0(.douta(w_n1068_0[0]),.doutb(w_n1068_0[1]),.din(n1068));
	jspl jspl_w_n1069_0(.douta(w_n1069_0[0]),.doutb(w_n1069_0[1]),.din(n1069));
	jspl3 jspl3_w_n1073_0(.douta(w_n1073_0[0]),.doutb(w_n1073_0[1]),.doutc(w_n1073_0[2]),.din(n1073));
	jspl jspl_w_n1075_0(.douta(w_dff_A_YNttyCCi4_0),.doutb(w_n1075_0[1]),.din(n1075));
	jspl jspl_w_n1076_0(.douta(w_dff_A_l1Fd4mzB7_0),.doutb(w_n1076_0[1]),.din(n1076));
	jspl3 jspl3_w_n1077_0(.douta(w_n1077_0[0]),.doutb(w_n1077_0[1]),.doutc(w_n1077_0[2]),.din(n1077));
	jspl3 jspl3_w_n1081_0(.douta(w_n1081_0[0]),.doutb(w_n1081_0[1]),.doutc(w_n1081_0[2]),.din(n1081));
	jspl jspl_w_n1082_0(.douta(w_n1082_0[0]),.doutb(w_n1082_0[1]),.din(n1082));
	jspl3 jspl3_w_n1086_0(.douta(w_n1086_0[0]),.doutb(w_n1086_0[1]),.doutc(w_n1086_0[2]),.din(n1086));
	jspl jspl_w_n1092_0(.douta(w_n1092_0[0]),.doutb(w_n1092_0[1]),.din(n1092));
	jspl jspl_w_n1095_0(.douta(w_dff_A_jdynXXo00_0),.doutb(w_n1095_0[1]),.din(n1095));
	jspl3 jspl3_w_n1096_0(.douta(w_n1096_0[0]),.doutb(w_n1096_0[1]),.doutc(w_n1096_0[2]),.din(n1096));
	jspl3 jspl3_w_n1100_0(.douta(w_n1100_0[0]),.doutb(w_n1100_0[1]),.doutc(w_n1100_0[2]),.din(n1100));
	jspl jspl_w_n1102_0(.douta(w_dff_A_dK8hF1rC4_0),.doutb(w_n1102_0[1]),.din(n1102));
	jspl jspl_w_n1104_0(.douta(w_n1104_0[0]),.doutb(w_dff_A_2H7UVBdK3_1),.din(n1104));
	jspl jspl_w_n1105_0(.douta(w_n1105_0[0]),.doutb(w_n1105_0[1]),.din(n1105));
	jspl jspl_w_n1116_0(.douta(w_n1116_0[0]),.doutb(w_n1116_0[1]),.din(n1116));
	jspl3 jspl3_w_n1122_0(.douta(w_n1122_0[0]),.doutb(w_n1122_0[1]),.doutc(w_n1122_0[2]),.din(n1122));
	jspl3 jspl3_w_n1125_0(.douta(w_n1125_0[0]),.doutb(w_n1125_0[1]),.doutc(w_n1125_0[2]),.din(w_dff_B_0iF05mWz2_3));
	jspl jspl_w_n1127_0(.douta(w_dff_A_DL60yFMg3_0),.doutb(w_n1127_0[1]),.din(w_dff_B_K27cHxuK1_2));
	jspl3 jspl3_w_n1128_0(.douta(w_n1128_0[0]),.doutb(w_n1128_0[1]),.doutc(w_n1128_0[2]),.din(n1128));
	jspl jspl_w_n1128_1(.douta(w_n1128_1[0]),.doutb(w_n1128_1[1]),.din(w_n1128_0[0]));
	jspl jspl_w_n1130_0(.douta(w_n1130_0[0]),.doutb(w_n1130_0[1]),.din(n1130));
	jspl jspl_w_n1136_0(.douta(w_n1136_0[0]),.doutb(w_dff_A_c9mCUYb77_1),.din(n1136));
	jspl jspl_w_n1142_0(.douta(w_n1142_0[0]),.doutb(w_n1142_0[1]),.din(n1142));
	jspl3 jspl3_w_n1148_0(.douta(w_n1148_0[0]),.doutb(w_n1148_0[1]),.doutc(w_dff_A_yMBoJk9R6_2),.din(n1148));
	jspl jspl_w_n1156_0(.douta(w_n1156_0[0]),.doutb(w_n1156_0[1]),.din(n1156));
	jspl jspl_w_n1166_0(.douta(w_n1166_0[0]),.doutb(w_n1166_0[1]),.din(n1166));
	jspl jspl_w_n1173_0(.douta(w_n1173_0[0]),.doutb(w_n1173_0[1]),.din(n1173));
	jspl jspl_w_n1189_0(.douta(w_n1189_0[0]),.doutb(w_n1189_0[1]),.din(n1189));
	jspl jspl_w_n1205_0(.douta(w_n1205_0[0]),.doutb(w_n1205_0[1]),.din(n1205));
	jspl jspl_w_n1236_0(.douta(w_dff_A_iQkRFewx6_0),.doutb(w_n1236_0[1]),.din(n1236));
	jspl jspl_w_n1244_0(.douta(w_n1244_0[0]),.doutb(w_n1244_0[1]),.din(n1244));
	jspl jspl_w_n1283_0(.douta(w_n1283_0[0]),.doutb(w_n1283_0[1]),.din(n1283));
	jspl jspl_w_n1301_0(.douta(w_n1301_0[0]),.doutb(w_dff_A_Hqdbi7JV4_1),.din(n1301));
	jspl jspl_w_n1309_0(.douta(w_n1309_0[0]),.doutb(w_n1309_0[1]),.din(n1309));
	jspl jspl_w_n1317_0(.douta(w_n1317_0[0]),.doutb(w_n1317_0[1]),.din(n1317));
	jspl jspl_w_n1325_0(.douta(w_n1325_0[0]),.doutb(w_n1325_0[1]),.din(n1325));
	jspl3 jspl3_w_n1359_0(.douta(w_n1359_0[0]),.doutb(w_dff_A_16N29usL4_1),.doutc(w_dff_A_pKYTFRI76_2),.din(n1359));
	jspl3 jspl3_w_n1360_0(.douta(w_n1360_0[0]),.doutb(w_dff_A_4tZotuGY6_1),.doutc(w_n1360_0[2]),.din(n1360));
	jspl jspl_w_n1360_1(.douta(w_n1360_1[0]),.doutb(w_dff_A_8DGK2zaE1_1),.din(w_n1360_0[0]));
	jspl jspl_w_n1361_0(.douta(w_n1361_0[0]),.doutb(w_dff_A_jO2s0pGZ6_1),.din(n1361));
	jspl jspl_w_n1362_0(.douta(w_n1362_0[0]),.doutb(w_n1362_0[1]),.din(n1362));
	jspl jspl_w_n1376_0(.douta(w_dff_A_tDZA1xRC0_0),.doutb(w_n1376_0[1]),.din(n1376));
	jspl3 jspl3_w_n1380_0(.douta(w_n1380_0[0]),.doutb(w_dff_A_OQdcaMSn4_1),.doutc(w_n1380_0[2]),.din(n1380));
	jspl jspl_w_n1380_1(.douta(w_n1380_1[0]),.doutb(w_n1380_1[1]),.din(w_n1380_0[0]));
	jspl3 jspl3_w_n1383_0(.douta(w_n1383_0[0]),.doutb(w_n1383_0[1]),.doutc(w_n1383_0[2]),.din(n1383));
	jspl3 jspl3_w_n1383_1(.douta(w_n1383_1[0]),.doutb(w_n1383_1[1]),.doutc(w_n1383_1[2]),.din(w_n1383_0[0]));
	jspl3 jspl3_w_n1385_0(.douta(w_n1385_0[0]),.doutb(w_n1385_0[1]),.doutc(w_n1385_0[2]),.din(n1385));
	jspl jspl_w_n1385_1(.douta(w_n1385_1[0]),.doutb(w_n1385_1[1]),.din(w_n1385_0[0]));
	jspl3 jspl3_w_n1389_0(.douta(w_n1389_0[0]),.doutb(w_n1389_0[1]),.doutc(w_n1389_0[2]),.din(n1389));
	jspl jspl_w_n1389_1(.douta(w_n1389_1[0]),.doutb(w_n1389_1[1]),.din(w_n1389_0[0]));
	jspl3 jspl3_w_n1392_0(.douta(w_n1392_0[0]),.doutb(w_n1392_0[1]),.doutc(w_n1392_0[2]),.din(n1392));
	jspl jspl_w_n1392_1(.douta(w_n1392_1[0]),.doutb(w_n1392_1[1]),.din(w_n1392_0[0]));
	jspl jspl_w_n1401_0(.douta(w_n1401_0[0]),.doutb(w_dff_A_ZmUqUEXr6_1),.din(w_dff_B_Ypk94iqM7_2));
	jspl jspl_w_n1402_0(.douta(w_dff_A_sYrWn1lF6_0),.doutb(w_n1402_0[1]),.din(w_dff_B_AUYeWQXa8_2));
	jspl jspl_w_n1403_0(.douta(w_dff_A_S1cGnyRj8_0),.doutb(w_n1403_0[1]),.din(w_dff_B_uPWYFGOB2_2));
	jspl jspl_w_n1404_0(.douta(w_n1404_0[0]),.doutb(w_dff_A_jOasjh7M6_1),.din(w_dff_B_pNqP6SDG5_2));
	jspl jspl_w_n1405_0(.douta(w_n1405_0[0]),.doutb(w_n1405_0[1]),.din(n1405));
	jspl jspl_w_n1406_0(.douta(w_n1406_0[0]),.doutb(w_n1406_0[1]),.din(n1406));
	jspl jspl_w_n1414_0(.douta(w_n1414_0[0]),.doutb(w_dff_A_mxJkPqv15_1),.din(n1414));
	jspl3 jspl3_w_n1420_0(.douta(w_n1420_0[0]),.doutb(w_dff_A_UQBvNC652_1),.doutc(w_dff_A_9egDAeHd7_2),.din(w_dff_B_jbCKAF4M3_3));
	jspl jspl_w_n1421_0(.douta(w_dff_A_T00sBlkf8_0),.doutb(w_n1421_0[1]),.din(w_dff_B_RFmgFe5b7_2));
	jspl jspl_w_n1422_0(.douta(w_dff_A_fzo1EyOA9_0),.doutb(w_n1422_0[1]),.din(w_dff_B_yF9TZLdu0_2));
	jspl jspl_w_n1424_0(.douta(w_n1424_0[0]),.doutb(w_n1424_0[1]),.din(n1424));
	jspl jspl_w_n1425_0(.douta(w_n1425_0[0]),.doutb(w_n1425_0[1]),.din(n1425));
	jspl3 jspl3_w_n1444_0(.douta(w_dff_A_TA0aTwIG6_0),.doutb(w_n1444_0[1]),.doutc(w_dff_A_W0oVwpZc9_2),.din(w_dff_B_nLkcjZeK0_3));
	jspl jspl_w_n1445_0(.douta(w_n1445_0[0]),.doutb(w_dff_A_sXuwNK8R4_1),.din(w_dff_B_oKWTF6hl0_2));
	jspl jspl_w_n1447_0(.douta(w_n1447_0[0]),.doutb(w_n1447_0[1]),.din(n1447));
	jspl jspl_w_n1454_0(.douta(w_n1454_0[0]),.doutb(w_dff_A_pHdo0g8s9_1),.din(w_dff_B_2QcC4uf46_2));
	jspl3 jspl3_w_n1463_0(.douta(w_dff_A_lOhW6SaF6_0),.doutb(w_dff_A_s5cqszX06_1),.doutc(w_n1463_0[2]),.din(n1463));
	jspl jspl_w_n1464_0(.douta(w_n1464_0[0]),.doutb(w_dff_A_YE6unQTE1_1),.din(w_dff_B_TNqvWjH05_2));
	jspl jspl_w_n1465_0(.douta(w_n1465_0[0]),.doutb(w_n1465_0[1]),.din(n1465));
	jspl jspl_w_n1468_0(.douta(w_n1468_0[0]),.doutb(w_dff_A_iKGJ2GEw0_1),.din(w_dff_B_0LmqApjW4_2));
	jspl jspl_w_n1469_0(.douta(w_dff_A_Ckj1AOyH1_0),.doutb(w_n1469_0[1]),.din(w_dff_B_La9vFLI37_2));
	jspl jspl_w_n1470_0(.douta(w_dff_A_cJhQqle97_0),.doutb(w_n1470_0[1]),.din(w_dff_B_KKg45cXB6_2));
	jspl jspl_w_n1471_0(.douta(w_n1471_0[0]),.doutb(w_dff_A_8wgZDwou2_1),.din(n1471));
	jspl jspl_w_n1472_0(.douta(w_n1472_0[0]),.doutb(w_n1472_0[1]),.din(n1472));
	jspl jspl_w_n1473_0(.douta(w_n1473_0[0]),.doutb(w_n1473_0[1]),.din(n1473));
	jspl jspl_w_n1479_0(.douta(w_n1479_0[0]),.doutb(w_dff_A_pe8t0RV05_1),.din(n1479));
	jspl jspl_w_n1482_0(.douta(w_n1482_0[0]),.doutb(w_dff_A_iLnKSvBK5_1),.din(n1482));
	jspl jspl_w_n1486_0(.douta(w_n1486_0[0]),.doutb(w_n1486_0[1]),.din(n1486));
	jspl3 jspl3_w_n1494_0(.douta(w_n1494_0[0]),.doutb(w_n1494_0[1]),.doutc(w_dff_A_lC5KzlNe7_2),.din(n1494));
	jspl jspl_w_n1501_0(.douta(w_n1501_0[0]),.doutb(w_dff_A_YS3sKKuK9_1),.din(n1501));
	jspl jspl_w_n1510_0(.douta(w_n1510_0[0]),.doutb(w_n1510_0[1]),.din(n1510));
	jspl jspl_w_n1520_0(.douta(w_n1520_0[0]),.doutb(w_dff_A_trCzAZP81_1),.din(n1520));
	jspl jspl_w_n1536_0(.douta(w_n1536_0[0]),.doutb(w_n1536_0[1]),.din(n1536));
	jspl jspl_w_n1571_0(.douta(w_n1571_0[0]),.doutb(w_n1571_0[1]),.din(n1571));
	jspl jspl_w_n1599_0(.douta(w_n1599_0[0]),.doutb(w_n1599_0[1]),.din(n1599));
	jspl jspl_w_n1610_0(.douta(w_n1610_0[0]),.doutb(w_n1610_0[1]),.din(w_dff_B_vDp3rU3n0_2));
	jspl jspl_w_n1611_0(.douta(w_n1611_0[0]),.doutb(w_n1611_0[1]),.din(n1611));
	jspl jspl_w_n1625_0(.douta(w_n1625_0[0]),.doutb(w_n1625_0[1]),.din(n1625));
	jspl jspl_w_n1642_0(.douta(w_n1642_0[0]),.doutb(w_n1642_0[1]),.din(n1642));
	jspl jspl_w_n1644_0(.douta(w_dff_A_G0ij57U76_0),.doutb(w_n1644_0[1]),.din(n1644));
	jspl jspl_w_n1651_0(.douta(w_n1651_0[0]),.doutb(w_dff_A_1oemz8iY6_1),.din(n1651));
	jspl jspl_w_n1654_0(.douta(w_n1654_0[0]),.doutb(w_dff_A_eGSqPnke0_1),.din(n1654));
	jspl jspl_w_n1659_0(.douta(w_n1659_0[0]),.doutb(w_n1659_0[1]),.din(n1659));
	jspl jspl_w_n1667_0(.douta(w_dff_A_1G1L2k840_0),.doutb(w_n1667_0[1]),.din(n1667));
	jspl jspl_w_n1670_0(.douta(w_n1670_0[0]),.doutb(w_n1670_0[1]),.din(n1670));
	jspl jspl_w_n1672_0(.douta(w_n1672_0[0]),.doutb(w_n1672_0[1]),.din(n1672));
	jspl jspl_w_n1675_0(.douta(w_n1675_0[0]),.doutb(w_dff_A_xRUPsRID2_1),.din(n1675));
	jspl jspl_w_n1680_0(.douta(w_n1680_0[0]),.doutb(w_n1680_0[1]),.din(n1680));
	jspl jspl_w_n1687_0(.douta(w_n1687_0[0]),.doutb(w_dff_A_PJc2GGi80_1),.din(n1687));
	jspl jspl_w_n1689_0(.douta(w_n1689_0[0]),.doutb(w_n1689_0[1]),.din(n1689));
	jspl jspl_w_n1699_0(.douta(w_n1699_0[0]),.doutb(w_n1699_0[1]),.din(n1699));
	jdff dff_A_Pos9QPwV7_0(.dout(w_G5_1[0]),.din(w_dff_A_Pos9QPwV7_0),.clk(gclk));
	jdff dff_A_XGfauPzp1_0(.dout(w_dff_A_Pos9QPwV7_0),.din(w_dff_A_XGfauPzp1_0),.clk(gclk));
	jdff dff_A_IEvszadD0_1(.dout(w_G5_1[1]),.din(w_dff_A_IEvszadD0_1),.clk(gclk));
	jdff dff_A_HjETiJKP7_1(.dout(w_G5_0[1]),.din(w_dff_A_HjETiJKP7_1),.clk(gclk));
	jdff dff_A_tdRIK4cs5_1(.dout(w_dff_A_HjETiJKP7_1),.din(w_dff_A_tdRIK4cs5_1),.clk(gclk));
	jdff dff_A_QndkNCew9_2(.dout(w_G5_0[2]),.din(w_dff_A_QndkNCew9_2),.clk(gclk));
	jdff dff_B_wgDSXUDG2_0(.din(n1131),.dout(w_dff_B_wgDSXUDG2_0),.clk(gclk));
	jdff dff_B_fWyqtvR81_3(.din(n1125),.dout(w_dff_B_fWyqtvR81_3),.clk(gclk));
	jdff dff_B_uoINvDSa8_3(.din(w_dff_B_fWyqtvR81_3),.dout(w_dff_B_uoINvDSa8_3),.clk(gclk));
	jdff dff_B_WTbhWZhI7_3(.din(w_dff_B_uoINvDSa8_3),.dout(w_dff_B_WTbhWZhI7_3),.clk(gclk));
	jdff dff_B_7QJvHfSv5_3(.din(w_dff_B_WTbhWZhI7_3),.dout(w_dff_B_7QJvHfSv5_3),.clk(gclk));
	jdff dff_B_uGCHlJxK9_3(.din(w_dff_B_7QJvHfSv5_3),.dout(w_dff_B_uGCHlJxK9_3),.clk(gclk));
	jdff dff_B_kbXJdWzf8_3(.din(w_dff_B_uGCHlJxK9_3),.dout(w_dff_B_kbXJdWzf8_3),.clk(gclk));
	jdff dff_B_gTpgSbmF2_3(.din(w_dff_B_kbXJdWzf8_3),.dout(w_dff_B_gTpgSbmF2_3),.clk(gclk));
	jdff dff_B_gsg21ktp1_3(.din(w_dff_B_gTpgSbmF2_3),.dout(w_dff_B_gsg21ktp1_3),.clk(gclk));
	jdff dff_B_nHZK4yve1_3(.din(w_dff_B_gsg21ktp1_3),.dout(w_dff_B_nHZK4yve1_3),.clk(gclk));
	jdff dff_B_htnMHrbg4_3(.din(w_dff_B_nHZK4yve1_3),.dout(w_dff_B_htnMHrbg4_3),.clk(gclk));
	jdff dff_B_q1wIQwTM4_3(.din(w_dff_B_htnMHrbg4_3),.dout(w_dff_B_q1wIQwTM4_3),.clk(gclk));
	jdff dff_B_NwX8w6Vb0_3(.din(w_dff_B_q1wIQwTM4_3),.dout(w_dff_B_NwX8w6Vb0_3),.clk(gclk));
	jdff dff_B_dJxNXdWa0_3(.din(w_dff_B_NwX8w6Vb0_3),.dout(w_dff_B_dJxNXdWa0_3),.clk(gclk));
	jdff dff_B_qfU08Cof6_3(.din(w_dff_B_dJxNXdWa0_3),.dout(w_dff_B_qfU08Cof6_3),.clk(gclk));
	jdff dff_B_nI1NuC2F0_3(.din(w_dff_B_qfU08Cof6_3),.dout(w_dff_B_nI1NuC2F0_3),.clk(gclk));
	jdff dff_B_0iF05mWz2_3(.din(w_dff_B_nI1NuC2F0_3),.dout(w_dff_B_0iF05mWz2_3),.clk(gclk));
	jdff dff_B_lqJRKDNW7_1(.din(n1123),.dout(w_dff_B_lqJRKDNW7_1),.clk(gclk));
	jdff dff_B_KC1varD37_0(.din(n1121),.dout(w_dff_B_KC1varD37_0),.clk(gclk));
	jdff dff_B_N91gti7d4_0(.din(w_dff_B_KC1varD37_0),.dout(w_dff_B_N91gti7d4_0),.clk(gclk));
	jdff dff_B_xXyVJF5x1_0(.din(w_dff_B_N91gti7d4_0),.dout(w_dff_B_xXyVJF5x1_0),.clk(gclk));
	jdff dff_B_zF2G5PQf4_0(.din(w_dff_B_xXyVJF5x1_0),.dout(w_dff_B_zF2G5PQf4_0),.clk(gclk));
	jdff dff_B_3IxjCjfR7_0(.din(w_dff_B_zF2G5PQf4_0),.dout(w_dff_B_3IxjCjfR7_0),.clk(gclk));
	jdff dff_B_1glBVTOx1_0(.din(w_dff_B_3IxjCjfR7_0),.dout(w_dff_B_1glBVTOx1_0),.clk(gclk));
	jdff dff_B_eowfTFGQ0_0(.din(w_dff_B_1glBVTOx1_0),.dout(w_dff_B_eowfTFGQ0_0),.clk(gclk));
	jdff dff_B_TR8eBgc44_0(.din(w_dff_B_eowfTFGQ0_0),.dout(w_dff_B_TR8eBgc44_0),.clk(gclk));
	jdff dff_B_uEgPLN9I8_0(.din(w_dff_B_TR8eBgc44_0),.dout(w_dff_B_uEgPLN9I8_0),.clk(gclk));
	jdff dff_B_4g0KHQgb9_0(.din(n1120),.dout(w_dff_B_4g0KHQgb9_0),.clk(gclk));
	jdff dff_B_UVTHnIgH5_0(.din(w_dff_B_4g0KHQgb9_0),.dout(w_dff_B_UVTHnIgH5_0),.clk(gclk));
	jdff dff_B_C5muFh6p3_0(.din(w_dff_B_UVTHnIgH5_0),.dout(w_dff_B_C5muFh6p3_0),.clk(gclk));
	jdff dff_B_DZE264KT4_0(.din(n1119),.dout(w_dff_B_DZE264KT4_0),.clk(gclk));
	jdff dff_B_SFE4sIHa2_0(.din(n1110),.dout(w_dff_B_SFE4sIHa2_0),.clk(gclk));
	jdff dff_B_pZAfrZYo5_0(.din(w_dff_B_SFE4sIHa2_0),.dout(w_dff_B_pZAfrZYo5_0),.clk(gclk));
	jdff dff_B_mTKgg1164_0(.din(w_dff_B_pZAfrZYo5_0),.dout(w_dff_B_mTKgg1164_0),.clk(gclk));
	jdff dff_B_L2KMdVHu3_0(.din(w_dff_B_mTKgg1164_0),.dout(w_dff_B_L2KMdVHu3_0),.clk(gclk));
	jdff dff_B_ryF06tMX0_0(.din(w_dff_B_L2KMdVHu3_0),.dout(w_dff_B_ryF06tMX0_0),.clk(gclk));
	jdff dff_B_ipbujmWF3_0(.din(w_dff_B_ryF06tMX0_0),.dout(w_dff_B_ipbujmWF3_0),.clk(gclk));
	jdff dff_B_RiW4jPHy1_0(.din(w_dff_B_ipbujmWF3_0),.dout(w_dff_B_RiW4jPHy1_0),.clk(gclk));
	jdff dff_B_w1tGP8yo3_0(.din(w_dff_B_RiW4jPHy1_0),.dout(w_dff_B_w1tGP8yo3_0),.clk(gclk));
	jdff dff_B_5EDT2rnP2_1(.din(n1089),.dout(w_dff_B_5EDT2rnP2_1),.clk(gclk));
	jdff dff_B_PhMNAOfy1_1(.din(w_dff_B_5EDT2rnP2_1),.dout(w_dff_B_PhMNAOfy1_1),.clk(gclk));
	jdff dff_B_V9LgDelO6_1(.din(n1093),.dout(w_dff_B_V9LgDelO6_1),.clk(gclk));
	jdff dff_A_2H7UVBdK3_1(.dout(w_n1104_0[1]),.din(w_dff_A_2H7UVBdK3_1),.clk(gclk));
	jdff dff_A_dK8hF1rC4_0(.dout(w_n1102_0[0]),.din(w_dff_A_dK8hF1rC4_0),.clk(gclk));
	jdff dff_A_XgMhCSMX3_0(.dout(w_n1075_0[0]),.din(w_dff_A_XgMhCSMX3_0),.clk(gclk));
	jdff dff_A_YNttyCCi4_0(.dout(w_dff_A_XgMhCSMX3_0),.din(w_dff_A_YNttyCCi4_0),.clk(gclk));
	jdff dff_B_bVaJ0Cf89_0(.din(n1059),.dout(w_dff_B_bVaJ0Cf89_0),.clk(gclk));
	jdff dff_B_gOANsO7i2_0(.din(w_dff_B_bVaJ0Cf89_0),.dout(w_dff_B_gOANsO7i2_0),.clk(gclk));
	jdff dff_B_xeUFODug7_0(.din(n1058),.dout(w_dff_B_xeUFODug7_0),.clk(gclk));
	jdff dff_B_xlePdhEl3_0(.din(w_dff_B_xeUFODug7_0),.dout(w_dff_B_xlePdhEl3_0),.clk(gclk));
	jdff dff_B_Gc98jEYO0_0(.din(w_dff_B_xlePdhEl3_0),.dout(w_dff_B_Gc98jEYO0_0),.clk(gclk));
	jdff dff_B_wkkZXIpM0_0(.din(w_dff_B_Gc98jEYO0_0),.dout(w_dff_B_wkkZXIpM0_0),.clk(gclk));
	jdff dff_B_ySOYDXTl2_0(.din(n1057),.dout(w_dff_B_ySOYDXTl2_0),.clk(gclk));
	jdff dff_B_RKBX27OC2_0(.din(n1050),.dout(w_dff_B_RKBX27OC2_0),.clk(gclk));
	jdff dff_B_vrsafaGC8_0(.din(w_dff_B_RKBX27OC2_0),.dout(w_dff_B_vrsafaGC8_0),.clk(gclk));
	jdff dff_B_ApusimQ42_0(.din(n1047),.dout(w_dff_B_ApusimQ42_0),.clk(gclk));
	jdff dff_A_bNXtfWRE3_1(.dout(w_n1022_0[1]),.din(w_dff_A_bNXtfWRE3_1),.clk(gclk));
	jdff dff_A_kAEMKNcT9_1(.dout(w_dff_A_bNXtfWRE3_1),.din(w_dff_A_kAEMKNcT9_1),.clk(gclk));
	jdff dff_A_koKZi9Uv9_1(.dout(w_dff_A_kAEMKNcT9_1),.din(w_dff_A_koKZi9Uv9_1),.clk(gclk));
	jdff dff_A_uBfCaew78_1(.dout(w_dff_A_koKZi9Uv9_1),.din(w_dff_A_uBfCaew78_1),.clk(gclk));
	jdff dff_A_YYyzousl5_1(.dout(w_dff_A_uBfCaew78_1),.din(w_dff_A_YYyzousl5_1),.clk(gclk));
	jdff dff_A_ReZ75tPd8_1(.dout(w_dff_A_YYyzousl5_1),.din(w_dff_A_ReZ75tPd8_1),.clk(gclk));
	jdff dff_B_tB2GeuHj0_2(.din(n1022),.dout(w_dff_B_tB2GeuHj0_2),.clk(gclk));
	jdff dff_B_MTWo24nU6_0(.din(n1021),.dout(w_dff_B_MTWo24nU6_0),.clk(gclk));
	jdff dff_B_AMOHr3Vf6_0(.din(w_dff_B_MTWo24nU6_0),.dout(w_dff_B_AMOHr3Vf6_0),.clk(gclk));
	jdff dff_B_n58IivwY1_0(.din(n1005),.dout(w_dff_B_n58IivwY1_0),.clk(gclk));
	jdff dff_A_EYKd06HK4_0(.dout(w_n1003_0[0]),.din(w_dff_A_EYKd06HK4_0),.clk(gclk));
	jdff dff_A_pYjNPTOh3_0(.dout(w_dff_A_EYKd06HK4_0),.din(w_dff_A_pYjNPTOh3_0),.clk(gclk));
	jdff dff_A_14yKmCqw2_1(.dout(w_n993_0[1]),.din(w_dff_A_14yKmCqw2_1),.clk(gclk));
	jdff dff_B_afESf26d0_1(.din(n768),.dout(w_dff_B_afESf26d0_1),.clk(gclk));
	jdff dff_B_SC8tEvs74_1(.din(w_dff_B_afESf26d0_1),.dout(w_dff_B_SC8tEvs74_1),.clk(gclk));
	jdff dff_B_234lh4O68_1(.din(w_dff_B_SC8tEvs74_1),.dout(w_dff_B_234lh4O68_1),.clk(gclk));
	jdff dff_B_9kGRiarq1_1(.din(w_dff_B_234lh4O68_1),.dout(w_dff_B_9kGRiarq1_1),.clk(gclk));
	jdff dff_B_RDXZWQRJ4_0(.din(n983),.dout(w_dff_B_RDXZWQRJ4_0),.clk(gclk));
	jdff dff_B_dJjfIWKK6_0(.din(w_dff_B_RDXZWQRJ4_0),.dout(w_dff_B_dJjfIWKK6_0),.clk(gclk));
	jdff dff_A_lYcNZSyi0_1(.dout(w_n865_0[1]),.din(w_dff_A_lYcNZSyi0_1),.clk(gclk));
	jdff dff_A_ZKFrcWGh3_1(.dout(w_n782_0[1]),.din(w_dff_A_ZKFrcWGh3_1),.clk(gclk));
	jdff dff_A_RJt6C40d5_1(.dout(w_dff_A_ZKFrcWGh3_1),.din(w_dff_A_RJt6C40d5_1),.clk(gclk));
	jdff dff_A_Q9txt8M98_1(.dout(w_dff_A_RJt6C40d5_1),.din(w_dff_A_Q9txt8M98_1),.clk(gclk));
	jdff dff_A_Mf0742Hd8_1(.dout(w_dff_A_Q9txt8M98_1),.din(w_dff_A_Mf0742Hd8_1),.clk(gclk));
	jdff dff_B_MDMrVRml4_1(.din(n774),.dout(w_dff_B_MDMrVRml4_1),.clk(gclk));
	jdff dff_B_GYqy8mHM6_0(.din(n776),.dout(w_dff_B_GYqy8mHM6_0),.clk(gclk));
	jdff dff_B_JeT5s1nr0_0(.din(n766),.dout(w_dff_B_JeT5s1nr0_0),.clk(gclk));
	jdff dff_B_lzCG9mPr6_0(.din(w_dff_B_JeT5s1nr0_0),.dout(w_dff_B_lzCG9mPr6_0),.clk(gclk));
	jdff dff_B_374cMAJc9_0(.din(w_dff_B_lzCG9mPr6_0),.dout(w_dff_B_374cMAJc9_0),.clk(gclk));
	jdff dff_A_SSZO0uzt5_0(.dout(w_n751_0[0]),.din(w_dff_A_SSZO0uzt5_0),.clk(gclk));
	jdff dff_A_qkOoyJRf5_0(.dout(w_dff_A_SSZO0uzt5_0),.din(w_dff_A_qkOoyJRf5_0),.clk(gclk));
	jdff dff_A_tR9lgU7T7_1(.dout(w_n742_0[1]),.din(w_dff_A_tR9lgU7T7_1),.clk(gclk));
	jdff dff_A_ekM6GQ1p6_1(.dout(w_dff_A_tR9lgU7T7_1),.din(w_dff_A_ekM6GQ1p6_1),.clk(gclk));
	jdff dff_A_gnYb3llh5_1(.dout(w_n735_0[1]),.din(w_dff_A_gnYb3llh5_1),.clk(gclk));
	jdff dff_A_yzHYW8jW8_1(.dout(w_dff_A_gnYb3llh5_1),.din(w_dff_A_yzHYW8jW8_1),.clk(gclk));
	jdff dff_B_NqZ7nwu76_2(.din(n735),.dout(w_dff_B_NqZ7nwu76_2),.clk(gclk));
	jdff dff_A_E9LU2zbd2_1(.dout(w_n728_0[1]),.din(w_dff_A_E9LU2zbd2_1),.clk(gclk));
	jdff dff_A_4eqkkdOn0_1(.dout(w_dff_A_E9LU2zbd2_1),.din(w_dff_A_4eqkkdOn0_1),.clk(gclk));
	jdff dff_A_atfaHIcj9_1(.dout(w_dff_A_4eqkkdOn0_1),.din(w_dff_A_atfaHIcj9_1),.clk(gclk));
	jdff dff_A_x53jfDaD6_1(.dout(w_dff_A_atfaHIcj9_1),.din(w_dff_A_x53jfDaD6_1),.clk(gclk));
	jdff dff_B_gdK7QGUf4_2(.din(n728),.dout(w_dff_B_gdK7QGUf4_2),.clk(gclk));
	jdff dff_B_2CyjtYCN9_1(.din(n1024),.dout(w_dff_B_2CyjtYCN9_1),.clk(gclk));
	jdff dff_B_NZtnnIIa5_1(.din(w_dff_B_2CyjtYCN9_1),.dout(w_dff_B_NZtnnIIa5_1),.clk(gclk));
	jdff dff_B_tkcTmpq62_1(.din(w_dff_B_NZtnnIIa5_1),.dout(w_dff_B_tkcTmpq62_1),.clk(gclk));
	jdff dff_B_T7vY4eHE7_1(.din(w_dff_B_tkcTmpq62_1),.dout(w_dff_B_T7vY4eHE7_1),.clk(gclk));
	jdff dff_B_oqO2spPR1_0(.din(n1031),.dout(w_dff_B_oqO2spPR1_0),.clk(gclk));
	jdff dff_B_CNs4IfNm6_0(.din(w_dff_B_oqO2spPR1_0),.dout(w_dff_B_CNs4IfNm6_0),.clk(gclk));
	jdff dff_B_P5WZjbkc1_0(.din(n1028),.dout(w_dff_B_P5WZjbkc1_0),.clk(gclk));
	jdff dff_B_4d4R3abv3_1(.din(n934),.dout(w_dff_B_4d4R3abv3_1),.clk(gclk));
	jdff dff_B_bSGiMxoB1_1(.din(n942),.dout(w_dff_B_bSGiMxoB1_1),.clk(gclk));
	jdff dff_B_5qNLIagO9_1(.din(n949),.dout(w_dff_B_5qNLIagO9_1),.clk(gclk));
	jdff dff_B_Maxmj71J6_1(.din(w_dff_B_5qNLIagO9_1),.dout(w_dff_B_Maxmj71J6_1),.clk(gclk));
	jdff dff_B_FVzcyAbF7_1(.din(n938),.dout(w_dff_B_FVzcyAbF7_1),.clk(gclk));
	jdff dff_B_lgvf0JUe6_1(.din(w_dff_B_FVzcyAbF7_1),.dout(w_dff_B_lgvf0JUe6_1),.clk(gclk));
	jdff dff_B_qOY9c4NC0_1(.din(G89),.dout(w_dff_B_qOY9c4NC0_1),.clk(gclk));
	jdff dff_B_2JkFxvEv9_1(.din(w_dff_B_qOY9c4NC0_1),.dout(w_dff_B_2JkFxvEv9_1),.clk(gclk));
	jdff dff_B_AN0P4XMB2_1(.din(w_dff_B_2JkFxvEv9_1),.dout(w_dff_B_AN0P4XMB2_1),.clk(gclk));
	jdff dff_B_mI1w0mBq3_1(.din(w_dff_B_AN0P4XMB2_1),.dout(w_dff_B_mI1w0mBq3_1),.clk(gclk));
	jdff dff_B_Yi2ITFyq1_1(.din(w_dff_B_mI1w0mBq3_1),.dout(w_dff_B_Yi2ITFyq1_1),.clk(gclk));
	jdff dff_A_7pUNrHii4_0(.dout(w_n939_0[0]),.din(w_dff_A_7pUNrHii4_0),.clk(gclk));
	jdff dff_B_LEyrmZNw7_1(.din(n922),.dout(w_dff_B_LEyrmZNw7_1),.clk(gclk));
	jdff dff_A_ze6hIAz33_1(.dout(w_n932_0[1]),.din(w_dff_A_ze6hIAz33_1),.clk(gclk));
	jdff dff_A_DrbNfpRo1_0(.dout(w_n905_0[0]),.din(w_dff_A_DrbNfpRo1_0),.clk(gclk));
	jdff dff_B_INOoEPE86_3(.din(n905),.dout(w_dff_B_INOoEPE86_3),.clk(gclk));
	jdff dff_B_2p6vx4go2_0(.din(n904),.dout(w_dff_B_2p6vx4go2_0),.clk(gclk));
	jdff dff_B_Uh0Dhd3p5_0(.din(w_dff_B_2p6vx4go2_0),.dout(w_dff_B_Uh0Dhd3p5_0),.clk(gclk));
	jdff dff_A_rwP99a5q0_0(.dout(w_n1044_0[0]),.din(w_dff_A_rwP99a5q0_0),.clk(gclk));
	jdff dff_B_kXm7rX3S9_2(.din(n1044),.dout(w_dff_B_kXm7rX3S9_2),.clk(gclk));
	jdff dff_B_N1uTPie67_0(.din(n1043),.dout(w_dff_B_N1uTPie67_0),.clk(gclk));
	jdff dff_B_wtZEieFg8_0(.din(n1040),.dout(w_dff_B_wtZEieFg8_0),.clk(gclk));
	jdff dff_B_w8MyrbaO0_0(.din(n1038),.dout(w_dff_B_w8MyrbaO0_0),.clk(gclk));
	jdff dff_B_XbHFmXLl3_0(.din(n1036),.dout(w_dff_B_XbHFmXLl3_0),.clk(gclk));
	jdff dff_B_0ybnmimc7_0(.din(w_dff_B_XbHFmXLl3_0),.dout(w_dff_B_0ybnmimc7_0),.clk(gclk));
	jdff dff_B_qVKgIB5E4_2(.din(n896),.dout(w_dff_B_qVKgIB5E4_2),.clk(gclk));
	jdff dff_A_oK3vFRv77_1(.dout(w_n887_0[1]),.din(w_dff_A_oK3vFRv77_1),.clk(gclk));
	jdff dff_B_CJYLLkVd5_0(.din(n883),.dout(w_dff_B_CJYLLkVd5_0),.clk(gclk));
	jdff dff_A_XaL3CtiK4_0(.dout(w_n874_0[0]),.din(w_dff_A_XaL3CtiK4_0),.clk(gclk));
	jdff dff_A_g9V4GvzL7_0(.dout(w_dff_A_XaL3CtiK4_0),.din(w_dff_A_g9V4GvzL7_0),.clk(gclk));
	jdff dff_A_RD61e9T25_0(.dout(w_n864_0[0]),.din(w_dff_A_RD61e9T25_0),.clk(gclk));
	jdff dff_A_MoDIOIRi2_0(.dout(w_dff_A_RD61e9T25_0),.din(w_dff_A_MoDIOIRi2_0),.clk(gclk));
	jdff dff_A_tWV56WJ98_0(.dout(w_dff_A_MoDIOIRi2_0),.din(w_dff_A_tWV56WJ98_0),.clk(gclk));
	jdff dff_A_j8FtofYP3_0(.dout(w_dff_A_tWV56WJ98_0),.din(w_dff_A_j8FtofYP3_0),.clk(gclk));
	jdff dff_B_HHy6QElJ5_1(.din(n837),.dout(w_dff_B_HHy6QElJ5_1),.clk(gclk));
	jdff dff_B_MLNtxgJY4_1(.din(n841),.dout(w_dff_B_MLNtxgJY4_1),.clk(gclk));
	jdff dff_B_2ir4DjU72_0(.din(n840),.dout(w_dff_B_2ir4DjU72_0),.clk(gclk));
	jdff dff_B_C3rdXGV10_1(.din(n825),.dout(w_dff_B_C3rdXGV10_1),.clk(gclk));
	jdff dff_A_bO3nzByT2_0(.dout(w_n981_0[0]),.din(w_dff_A_bO3nzByT2_0),.clk(gclk));
	jdff dff_A_ajdf93iQ9_0(.dout(w_dff_A_bO3nzByT2_0),.din(w_dff_A_ajdf93iQ9_0),.clk(gclk));
	jdff dff_A_AgAEvzEB1_0(.dout(w_dff_A_ajdf93iQ9_0),.din(w_dff_A_AgAEvzEB1_0),.clk(gclk));
	jdff dff_A_9AfuIthu8_0(.dout(w_dff_A_AgAEvzEB1_0),.din(w_dff_A_9AfuIthu8_0),.clk(gclk));
	jdff dff_A_Mdj67B3H9_0(.dout(w_dff_A_9AfuIthu8_0),.din(w_dff_A_Mdj67B3H9_0),.clk(gclk));
	jdff dff_A_7YvRhIar6_0(.dout(w_dff_A_Mdj67B3H9_0),.din(w_dff_A_7YvRhIar6_0),.clk(gclk));
	jdff dff_B_pxRVTx135_0(.din(n980),.dout(w_dff_B_pxRVTx135_0),.clk(gclk));
	jdff dff_A_wUpRfK0p1_0(.dout(w_n848_0[0]),.din(w_dff_A_wUpRfK0p1_0),.clk(gclk));
	jdff dff_A_rALwFiav9_2(.dout(w_n858_0[2]),.din(w_dff_A_rALwFiav9_2),.clk(gclk));
	jdff dff_A_uObGZouh4_1(.dout(w_n856_0[1]),.din(w_dff_A_uObGZouh4_1),.clk(gclk));
	jdff dff_A_kvQeBA0D2_0(.dout(w_n824_0[0]),.din(w_dff_A_kvQeBA0D2_0),.clk(gclk));
	jdff dff_A_4IEJ6hOt6_0(.dout(w_n810_0[0]),.din(w_dff_A_4IEJ6hOt6_0),.clk(gclk));
	jdff dff_A_q9dCrBA79_0(.dout(w_dff_A_4IEJ6hOt6_0),.din(w_dff_A_q9dCrBA79_0),.clk(gclk));
	jdff dff_A_vhkzGJZA8_0(.dout(w_dff_A_q9dCrBA79_0),.din(w_dff_A_vhkzGJZA8_0),.clk(gclk));
	jdff dff_A_RJjKOlTb6_0(.dout(w_dff_A_vhkzGJZA8_0),.din(w_dff_A_RJjKOlTb6_0),.clk(gclk));
	jdff dff_A_lonv2OjE2_0(.dout(w_dff_A_RJjKOlTb6_0),.din(w_dff_A_lonv2OjE2_0),.clk(gclk));
	jdff dff_A_BAORIDP98_0(.dout(w_dff_A_lonv2OjE2_0),.din(w_dff_A_BAORIDP98_0),.clk(gclk));
	jdff dff_A_aZDu4bpW2_0(.dout(w_dff_A_BAORIDP98_0),.din(w_dff_A_aZDu4bpW2_0),.clk(gclk));
	jdff dff_A_sbM22p8l0_2(.dout(w_n810_0[2]),.din(w_dff_A_sbM22p8l0_2),.clk(gclk));
	jdff dff_B_Lt3ej8b54_3(.din(n810),.dout(w_dff_B_Lt3ej8b54_3),.clk(gclk));
	jdff dff_B_7O3vY0Tl6_3(.din(w_dff_B_Lt3ej8b54_3),.dout(w_dff_B_7O3vY0Tl6_3),.clk(gclk));
	jdff dff_A_GjdtnPFR2_0(.dout(w_n972_0[0]),.din(w_dff_A_GjdtnPFR2_0),.clk(gclk));
	jdff dff_A_OV1iY6yU0_0(.dout(w_dff_A_GjdtnPFR2_0),.din(w_dff_A_OV1iY6yU0_0),.clk(gclk));
	jdff dff_A_BPA1aUZG7_0(.dout(w_dff_A_OV1iY6yU0_0),.din(w_dff_A_BPA1aUZG7_0),.clk(gclk));
	jdff dff_A_vv33bzPQ6_0(.dout(w_dff_A_BPA1aUZG7_0),.din(w_dff_A_vv33bzPQ6_0),.clk(gclk));
	jdff dff_A_aH6FkRrb9_0(.dout(w_dff_A_vv33bzPQ6_0),.din(w_dff_A_aH6FkRrb9_0),.clk(gclk));
	jdff dff_A_vpyBiBU25_0(.dout(w_dff_A_aH6FkRrb9_0),.din(w_dff_A_vpyBiBU25_0),.clk(gclk));
	jdff dff_A_zhxyA46L1_0(.dout(w_dff_A_vpyBiBU25_0),.din(w_dff_A_zhxyA46L1_0),.clk(gclk));
	jdff dff_B_sHtAJ7Vc2_2(.din(n972),.dout(w_dff_B_sHtAJ7Vc2_2),.clk(gclk));
	jdff dff_B_Ub74zJxg8_1(.din(n962),.dout(w_dff_B_Ub74zJxg8_1),.clk(gclk));
	jdff dff_B_3dEfFBv87_1(.din(n963),.dout(w_dff_B_3dEfFBv87_1),.clk(gclk));
	jdff dff_B_GRMGV4p45_1(.din(w_dff_B_3dEfFBv87_1),.dout(w_dff_B_GRMGV4p45_1),.clk(gclk));
	jdff dff_A_sYrWn1lF6_0(.dout(w_n1402_0[0]),.din(w_dff_A_sYrWn1lF6_0),.clk(gclk));
	jdff dff_B_5UkBZUQG5_2(.din(n1402),.dout(w_dff_B_5UkBZUQG5_2),.clk(gclk));
	jdff dff_B_Lx68BShZ5_2(.din(w_dff_B_5UkBZUQG5_2),.dout(w_dff_B_Lx68BShZ5_2),.clk(gclk));
	jdff dff_B_BalxW1tI9_2(.din(w_dff_B_Lx68BShZ5_2),.dout(w_dff_B_BalxW1tI9_2),.clk(gclk));
	jdff dff_B_5uR70sS67_2(.din(w_dff_B_BalxW1tI9_2),.dout(w_dff_B_5uR70sS67_2),.clk(gclk));
	jdff dff_B_r7oTZR028_2(.din(w_dff_B_5uR70sS67_2),.dout(w_dff_B_r7oTZR028_2),.clk(gclk));
	jdff dff_B_bCdNpCG38_2(.din(w_dff_B_r7oTZR028_2),.dout(w_dff_B_bCdNpCG38_2),.clk(gclk));
	jdff dff_B_1606UYPJ6_2(.din(w_dff_B_bCdNpCG38_2),.dout(w_dff_B_1606UYPJ6_2),.clk(gclk));
	jdff dff_B_0tVqPFTC9_2(.din(w_dff_B_1606UYPJ6_2),.dout(w_dff_B_0tVqPFTC9_2),.clk(gclk));
	jdff dff_B_3opfKOob2_2(.din(w_dff_B_0tVqPFTC9_2),.dout(w_dff_B_3opfKOob2_2),.clk(gclk));
	jdff dff_B_hafqao8N8_2(.din(w_dff_B_3opfKOob2_2),.dout(w_dff_B_hafqao8N8_2),.clk(gclk));
	jdff dff_B_8Nc6R9i03_2(.din(w_dff_B_hafqao8N8_2),.dout(w_dff_B_8Nc6R9i03_2),.clk(gclk));
	jdff dff_B_AiAGUhmX1_2(.din(w_dff_B_8Nc6R9i03_2),.dout(w_dff_B_AiAGUhmX1_2),.clk(gclk));
	jdff dff_B_AUYeWQXa8_2(.din(w_dff_B_AiAGUhmX1_2),.dout(w_dff_B_AUYeWQXa8_2),.clk(gclk));
	jdff dff_A_S1cGnyRj8_0(.dout(w_n1403_0[0]),.din(w_dff_A_S1cGnyRj8_0),.clk(gclk));
	jdff dff_B_746NndkO3_2(.din(n1403),.dout(w_dff_B_746NndkO3_2),.clk(gclk));
	jdff dff_B_ytwst5vl8_2(.din(w_dff_B_746NndkO3_2),.dout(w_dff_B_ytwst5vl8_2),.clk(gclk));
	jdff dff_B_x7fUxwPR6_2(.din(w_dff_B_ytwst5vl8_2),.dout(w_dff_B_x7fUxwPR6_2),.clk(gclk));
	jdff dff_B_aB5VuoxX1_2(.din(w_dff_B_x7fUxwPR6_2),.dout(w_dff_B_aB5VuoxX1_2),.clk(gclk));
	jdff dff_B_5EYh9UZe2_2(.din(w_dff_B_aB5VuoxX1_2),.dout(w_dff_B_5EYh9UZe2_2),.clk(gclk));
	jdff dff_B_W1OiaX8U2_2(.din(w_dff_B_5EYh9UZe2_2),.dout(w_dff_B_W1OiaX8U2_2),.clk(gclk));
	jdff dff_B_CqLy1fsw5_2(.din(w_dff_B_W1OiaX8U2_2),.dout(w_dff_B_CqLy1fsw5_2),.clk(gclk));
	jdff dff_B_LGxucHPi1_2(.din(w_dff_B_CqLy1fsw5_2),.dout(w_dff_B_LGxucHPi1_2),.clk(gclk));
	jdff dff_B_LYL7E7sq7_2(.din(w_dff_B_LGxucHPi1_2),.dout(w_dff_B_LYL7E7sq7_2),.clk(gclk));
	jdff dff_B_np24wlFa0_2(.din(w_dff_B_LYL7E7sq7_2),.dout(w_dff_B_np24wlFa0_2),.clk(gclk));
	jdff dff_B_vVWifAh97_2(.din(w_dff_B_np24wlFa0_2),.dout(w_dff_B_vVWifAh97_2),.clk(gclk));
	jdff dff_B_uPWYFGOB2_2(.din(w_dff_B_vVWifAh97_2),.dout(w_dff_B_uPWYFGOB2_2),.clk(gclk));
	jdff dff_B_5khcQBDh4_1(.din(n1429),.dout(w_dff_B_5khcQBDh4_1),.clk(gclk));
	jdff dff_B_OcWJQwsh7_1(.din(w_dff_B_5khcQBDh4_1),.dout(w_dff_B_OcWJQwsh7_1),.clk(gclk));
	jdff dff_B_Mkf1omzt6_1(.din(w_dff_B_OcWJQwsh7_1),.dout(w_dff_B_Mkf1omzt6_1),.clk(gclk));
	jdff dff_B_I9yQ9RFt1_1(.din(w_dff_B_Mkf1omzt6_1),.dout(w_dff_B_I9yQ9RFt1_1),.clk(gclk));
	jdff dff_B_wuRRRZup3_1(.din(w_dff_B_I9yQ9RFt1_1),.dout(w_dff_B_wuRRRZup3_1),.clk(gclk));
	jdff dff_B_zAvWvozQ3_1(.din(w_dff_B_wuRRRZup3_1),.dout(w_dff_B_zAvWvozQ3_1),.clk(gclk));
	jdff dff_B_EBsxEAGr1_1(.din(w_dff_B_zAvWvozQ3_1),.dout(w_dff_B_EBsxEAGr1_1),.clk(gclk));
	jdff dff_B_u8elYLWU8_1(.din(w_dff_B_EBsxEAGr1_1),.dout(w_dff_B_u8elYLWU8_1),.clk(gclk));
	jdff dff_B_u1ar03Fe3_1(.din(w_dff_B_u8elYLWU8_1),.dout(w_dff_B_u1ar03Fe3_1),.clk(gclk));
	jdff dff_B_lWOZhuri6_1(.din(w_dff_B_u1ar03Fe3_1),.dout(w_dff_B_lWOZhuri6_1),.clk(gclk));
	jdff dff_B_vLvoP0xY1_1(.din(w_dff_B_lWOZhuri6_1),.dout(w_dff_B_vLvoP0xY1_1),.clk(gclk));
	jdff dff_B_wHaSt9t09_1(.din(w_dff_B_vLvoP0xY1_1),.dout(w_dff_B_wHaSt9t09_1),.clk(gclk));
	jdff dff_A_T00sBlkf8_0(.dout(w_n1421_0[0]),.din(w_dff_A_T00sBlkf8_0),.clk(gclk));
	jdff dff_B_dAJRi7KG0_2(.din(n1421),.dout(w_dff_B_dAJRi7KG0_2),.clk(gclk));
	jdff dff_B_J5IjTRTA3_2(.din(w_dff_B_dAJRi7KG0_2),.dout(w_dff_B_J5IjTRTA3_2),.clk(gclk));
	jdff dff_B_8MXUWefQ3_2(.din(w_dff_B_J5IjTRTA3_2),.dout(w_dff_B_8MXUWefQ3_2),.clk(gclk));
	jdff dff_B_BvOQF7Do1_2(.din(w_dff_B_8MXUWefQ3_2),.dout(w_dff_B_BvOQF7Do1_2),.clk(gclk));
	jdff dff_B_20Yr7Jtx5_2(.din(w_dff_B_BvOQF7Do1_2),.dout(w_dff_B_20Yr7Jtx5_2),.clk(gclk));
	jdff dff_B_jRDqtOyY5_2(.din(w_dff_B_20Yr7Jtx5_2),.dout(w_dff_B_jRDqtOyY5_2),.clk(gclk));
	jdff dff_B_ngA7dIag5_2(.din(w_dff_B_jRDqtOyY5_2),.dout(w_dff_B_ngA7dIag5_2),.clk(gclk));
	jdff dff_B_jz2kvfDP2_2(.din(w_dff_B_ngA7dIag5_2),.dout(w_dff_B_jz2kvfDP2_2),.clk(gclk));
	jdff dff_B_eDlhJ25O6_2(.din(w_dff_B_jz2kvfDP2_2),.dout(w_dff_B_eDlhJ25O6_2),.clk(gclk));
	jdff dff_B_bRoaWIUD0_2(.din(w_dff_B_eDlhJ25O6_2),.dout(w_dff_B_bRoaWIUD0_2),.clk(gclk));
	jdff dff_B_Ce5B3vS49_2(.din(w_dff_B_bRoaWIUD0_2),.dout(w_dff_B_Ce5B3vS49_2),.clk(gclk));
	jdff dff_B_QvM587fe2_2(.din(w_dff_B_Ce5B3vS49_2),.dout(w_dff_B_QvM587fe2_2),.clk(gclk));
	jdff dff_B_n5UtTM7n8_2(.din(w_dff_B_QvM587fe2_2),.dout(w_dff_B_n5UtTM7n8_2),.clk(gclk));
	jdff dff_B_4itl8JOs0_2(.din(w_dff_B_n5UtTM7n8_2),.dout(w_dff_B_4itl8JOs0_2),.clk(gclk));
	jdff dff_B_rpvwD1GV5_2(.din(w_dff_B_4itl8JOs0_2),.dout(w_dff_B_rpvwD1GV5_2),.clk(gclk));
	jdff dff_B_gPVNGtcT7_2(.din(w_dff_B_rpvwD1GV5_2),.dout(w_dff_B_gPVNGtcT7_2),.clk(gclk));
	jdff dff_B_RFmgFe5b7_2(.din(w_dff_B_gPVNGtcT7_2),.dout(w_dff_B_RFmgFe5b7_2),.clk(gclk));
	jdff dff_B_CtWkk8hY4_1(.din(n1432),.dout(w_dff_B_CtWkk8hY4_1),.clk(gclk));
	jdff dff_B_0x2VHRbv1_1(.din(w_dff_B_CtWkk8hY4_1),.dout(w_dff_B_0x2VHRbv1_1),.clk(gclk));
	jdff dff_B_NXHes7CG4_1(.din(w_dff_B_0x2VHRbv1_1),.dout(w_dff_B_NXHes7CG4_1),.clk(gclk));
	jdff dff_B_I7Upk33g6_1(.din(w_dff_B_NXHes7CG4_1),.dout(w_dff_B_I7Upk33g6_1),.clk(gclk));
	jdff dff_B_dAjkBzzb0_1(.din(w_dff_B_I7Upk33g6_1),.dout(w_dff_B_dAjkBzzb0_1),.clk(gclk));
	jdff dff_B_iK0ZXs7J2_1(.din(w_dff_B_dAjkBzzb0_1),.dout(w_dff_B_iK0ZXs7J2_1),.clk(gclk));
	jdff dff_B_3q7MxW0d0_1(.din(w_dff_B_iK0ZXs7J2_1),.dout(w_dff_B_3q7MxW0d0_1),.clk(gclk));
	jdff dff_B_02u2SS0A2_1(.din(w_dff_B_3q7MxW0d0_1),.dout(w_dff_B_02u2SS0A2_1),.clk(gclk));
	jdff dff_B_0LIEmeDZ2_1(.din(w_dff_B_02u2SS0A2_1),.dout(w_dff_B_0LIEmeDZ2_1),.clk(gclk));
	jdff dff_B_p37xndZ06_1(.din(w_dff_B_0LIEmeDZ2_1),.dout(w_dff_B_p37xndZ06_1),.clk(gclk));
	jdff dff_B_YG5cchkR7_1(.din(w_dff_B_p37xndZ06_1),.dout(w_dff_B_YG5cchkR7_1),.clk(gclk));
	jdff dff_B_BVxSmfl52_1(.din(w_dff_B_YG5cchkR7_1),.dout(w_dff_B_BVxSmfl52_1),.clk(gclk));
	jdff dff_B_PYxL9Co86_1(.din(w_dff_B_BVxSmfl52_1),.dout(w_dff_B_PYxL9Co86_1),.clk(gclk));
	jdff dff_B_XisaLX904_0(.din(n1423),.dout(w_dff_B_XisaLX904_0),.clk(gclk));
	jdff dff_B_q9YFTezs7_0(.din(w_dff_B_XisaLX904_0),.dout(w_dff_B_q9YFTezs7_0),.clk(gclk));
	jdff dff_B_w2up1oTz5_0(.din(w_dff_B_q9YFTezs7_0),.dout(w_dff_B_w2up1oTz5_0),.clk(gclk));
	jdff dff_B_wmBPS0CK8_0(.din(w_dff_B_w2up1oTz5_0),.dout(w_dff_B_wmBPS0CK8_0),.clk(gclk));
	jdff dff_B_JVLeYO0G3_0(.din(w_dff_B_wmBPS0CK8_0),.dout(w_dff_B_JVLeYO0G3_0),.clk(gclk));
	jdff dff_B_bTJhcQWi8_0(.din(w_dff_B_JVLeYO0G3_0),.dout(w_dff_B_bTJhcQWi8_0),.clk(gclk));
	jdff dff_B_dYISN1vL1_0(.din(w_dff_B_bTJhcQWi8_0),.dout(w_dff_B_dYISN1vL1_0),.clk(gclk));
	jdff dff_B_sDosGpL87_0(.din(w_dff_B_dYISN1vL1_0),.dout(w_dff_B_sDosGpL87_0),.clk(gclk));
	jdff dff_B_YofwYuaG2_0(.din(w_dff_B_sDosGpL87_0),.dout(w_dff_B_YofwYuaG2_0),.clk(gclk));
	jdff dff_B_sDdFbHZ11_0(.din(w_dff_B_YofwYuaG2_0),.dout(w_dff_B_sDdFbHZ11_0),.clk(gclk));
	jdff dff_B_FlHUG2RS1_0(.din(w_dff_B_sDdFbHZ11_0),.dout(w_dff_B_FlHUG2RS1_0),.clk(gclk));
	jdff dff_B_CvdsZYuR1_0(.din(w_dff_B_FlHUG2RS1_0),.dout(w_dff_B_CvdsZYuR1_0),.clk(gclk));
	jdff dff_B_mt8eOiKy4_0(.din(w_dff_B_CvdsZYuR1_0),.dout(w_dff_B_mt8eOiKy4_0),.clk(gclk));
	jdff dff_B_PUHfyred4_0(.din(w_dff_B_mt8eOiKy4_0),.dout(w_dff_B_PUHfyred4_0),.clk(gclk));
	jdff dff_A_fzo1EyOA9_0(.dout(w_n1422_0[0]),.din(w_dff_A_fzo1EyOA9_0),.clk(gclk));
	jdff dff_B_MOoZF4NQ8_2(.din(n1422),.dout(w_dff_B_MOoZF4NQ8_2),.clk(gclk));
	jdff dff_B_4HTsDXSe4_2(.din(w_dff_B_MOoZF4NQ8_2),.dout(w_dff_B_4HTsDXSe4_2),.clk(gclk));
	jdff dff_B_z5dpkfli4_2(.din(w_dff_B_4HTsDXSe4_2),.dout(w_dff_B_z5dpkfli4_2),.clk(gclk));
	jdff dff_B_xWmAT5HH3_2(.din(w_dff_B_z5dpkfli4_2),.dout(w_dff_B_xWmAT5HH3_2),.clk(gclk));
	jdff dff_B_87SFmAYK4_2(.din(w_dff_B_xWmAT5HH3_2),.dout(w_dff_B_87SFmAYK4_2),.clk(gclk));
	jdff dff_B_hLpvyjlw0_2(.din(w_dff_B_87SFmAYK4_2),.dout(w_dff_B_hLpvyjlw0_2),.clk(gclk));
	jdff dff_B_ix3vso725_2(.din(w_dff_B_hLpvyjlw0_2),.dout(w_dff_B_ix3vso725_2),.clk(gclk));
	jdff dff_B_6gkSW4iq7_2(.din(w_dff_B_ix3vso725_2),.dout(w_dff_B_6gkSW4iq7_2),.clk(gclk));
	jdff dff_B_HVV2WRDk6_2(.din(w_dff_B_6gkSW4iq7_2),.dout(w_dff_B_HVV2WRDk6_2),.clk(gclk));
	jdff dff_B_jp264nbJ3_2(.din(w_dff_B_HVV2WRDk6_2),.dout(w_dff_B_jp264nbJ3_2),.clk(gclk));
	jdff dff_B_94YtK0fd1_2(.din(w_dff_B_jp264nbJ3_2),.dout(w_dff_B_94YtK0fd1_2),.clk(gclk));
	jdff dff_B_KFMkvf9j7_2(.din(w_dff_B_94YtK0fd1_2),.dout(w_dff_B_KFMkvf9j7_2),.clk(gclk));
	jdff dff_B_ZEbX4XJv2_2(.din(w_dff_B_KFMkvf9j7_2),.dout(w_dff_B_ZEbX4XJv2_2),.clk(gclk));
	jdff dff_B_CzMhrrsW6_2(.din(w_dff_B_ZEbX4XJv2_2),.dout(w_dff_B_CzMhrrsW6_2),.clk(gclk));
	jdff dff_B_TsEdxkGT1_2(.din(w_dff_B_CzMhrrsW6_2),.dout(w_dff_B_TsEdxkGT1_2),.clk(gclk));
	jdff dff_B_yF9TZLdu0_2(.din(w_dff_B_TsEdxkGT1_2),.dout(w_dff_B_yF9TZLdu0_2),.clk(gclk));
	jdff dff_B_hCYdVrMU3_0(.din(n1441),.dout(w_dff_B_hCYdVrMU3_0),.clk(gclk));
	jdff dff_B_zZmEURSA8_0(.din(n1440),.dout(w_dff_B_zZmEURSA8_0),.clk(gclk));
	jdff dff_B_EO7nhuqW7_0(.din(w_dff_B_zZmEURSA8_0),.dout(w_dff_B_EO7nhuqW7_0),.clk(gclk));
	jdff dff_B_Myj1SZaj4_0(.din(w_dff_B_EO7nhuqW7_0),.dout(w_dff_B_Myj1SZaj4_0),.clk(gclk));
	jdff dff_B_Qk0SAoBB3_0(.din(w_dff_B_Myj1SZaj4_0),.dout(w_dff_B_Qk0SAoBB3_0),.clk(gclk));
	jdff dff_B_pwXohnk63_0(.din(w_dff_B_Qk0SAoBB3_0),.dout(w_dff_B_pwXohnk63_0),.clk(gclk));
	jdff dff_B_bln28hL01_0(.din(w_dff_B_pwXohnk63_0),.dout(w_dff_B_bln28hL01_0),.clk(gclk));
	jdff dff_B_RWA6pG1u7_0(.din(n1212),.dout(w_dff_B_RWA6pG1u7_0),.clk(gclk));
	jdff dff_B_PXNiVJ5t5_0(.din(n1209),.dout(w_dff_B_PXNiVJ5t5_0),.clk(gclk));
	jdff dff_B_MqGAPJKl8_1(.din(n1206),.dout(w_dff_B_MqGAPJKl8_1),.clk(gclk));
	jdff dff_B_jid7V4CH7_1(.din(n1204),.dout(w_dff_B_jid7V4CH7_1),.clk(gclk));
	jdff dff_B_BBu6uxmD6_0(.din(n1197),.dout(w_dff_B_BBu6uxmD6_0),.clk(gclk));
	jdff dff_B_7gLDT3bK5_1(.din(n1190),.dout(w_dff_B_7gLDT3bK5_1),.clk(gclk));
	jdff dff_B_3eoJBKu19_1(.din(w_dff_B_7gLDT3bK5_1),.dout(w_dff_B_3eoJBKu19_1),.clk(gclk));
	jdff dff_B_3mrAU2E69_1(.din(n1188),.dout(w_dff_B_3mrAU2E69_1),.clk(gclk));
	jdff dff_B_o2vmRTrk6_1(.din(n1175),.dout(w_dff_B_o2vmRTrk6_1),.clk(gclk));
	jdff dff_B_9mCP92cT2_1(.din(w_dff_B_o2vmRTrk6_1),.dout(w_dff_B_9mCP92cT2_1),.clk(gclk));
	jdff dff_B_kRuQ7SBN6_1(.din(w_dff_B_9mCP92cT2_1),.dout(w_dff_B_kRuQ7SBN6_1),.clk(gclk));
	jdff dff_B_h5HuSvVj9_1(.din(w_dff_B_kRuQ7SBN6_1),.dout(w_dff_B_h5HuSvVj9_1),.clk(gclk));
	jdff dff_B_wiKNmkLb3_1(.din(n1176),.dout(w_dff_B_wiKNmkLb3_1),.clk(gclk));
	jdff dff_B_hMQE5yCy6_1(.din(w_dff_B_wiKNmkLb3_1),.dout(w_dff_B_hMQE5yCy6_1),.clk(gclk));
	jdff dff_B_WsO6eCcY2_1(.din(w_dff_B_hMQE5yCy6_1),.dout(w_dff_B_WsO6eCcY2_1),.clk(gclk));
	jdff dff_B_1PUvQFvx8_1(.din(w_dff_B_WsO6eCcY2_1),.dout(w_dff_B_1PUvQFvx8_1),.clk(gclk));
	jdff dff_B_RLt04rw04_1(.din(n1181),.dout(w_dff_B_RLt04rw04_1),.clk(gclk));
	jdff dff_B_KvbD5UbJ4_0(.din(n1174),.dout(w_dff_B_KvbD5UbJ4_0),.clk(gclk));
	jdff dff_B_DMTwZLiq9_0(.din(w_dff_B_KvbD5UbJ4_0),.dout(w_dff_B_DMTwZLiq9_0),.clk(gclk));
	jdff dff_B_S8pldWix3_1(.din(n1153),.dout(w_dff_B_S8pldWix3_1),.clk(gclk));
	jdff dff_B_zn8jTR373_1(.din(w_dff_B_S8pldWix3_1),.dout(w_dff_B_zn8jTR373_1),.clk(gclk));
	jdff dff_B_gkcq18WH8_1(.din(w_dff_B_zn8jTR373_1),.dout(w_dff_B_gkcq18WH8_1),.clk(gclk));
	jdff dff_B_vpusSyN26_1(.din(w_dff_B_gkcq18WH8_1),.dout(w_dff_B_vpusSyN26_1),.clk(gclk));
	jdff dff_B_S0kEqjWA1_1(.din(w_dff_B_vpusSyN26_1),.dout(w_dff_B_S0kEqjWA1_1),.clk(gclk));
	jdff dff_B_ffWWzdU89_1(.din(n1155),.dout(w_dff_B_ffWWzdU89_1),.clk(gclk));
	jdff dff_B_hEFGgJ5U5_1(.din(w_dff_B_ffWWzdU89_1),.dout(w_dff_B_hEFGgJ5U5_1),.clk(gclk));
	jdff dff_B_vpv4Ip8T8_1(.din(w_dff_B_hEFGgJ5U5_1),.dout(w_dff_B_vpv4Ip8T8_1),.clk(gclk));
	jdff dff_B_lOTosTFb6_0(.din(n1169),.dout(w_dff_B_lOTosTFb6_0),.clk(gclk));
	jdff dff_B_RolcQy8L8_0(.din(w_dff_B_lOTosTFb6_0),.dout(w_dff_B_RolcQy8L8_0),.clk(gclk));
	jdff dff_B_SziSQuS05_0(.din(w_dff_B_RolcQy8L8_0),.dout(w_dff_B_SziSQuS05_0),.clk(gclk));
	jdff dff_B_9Wcolvdi7_0(.din(w_dff_B_SziSQuS05_0),.dout(w_dff_B_9Wcolvdi7_0),.clk(gclk));
	jdff dff_B_pgKwBpz86_0(.din(n1355),.dout(w_dff_B_pgKwBpz86_0),.clk(gclk));
	jdff dff_B_m95GODcv4_0(.din(w_dff_B_pgKwBpz86_0),.dout(w_dff_B_m95GODcv4_0),.clk(gclk));
	jdff dff_B_kKkyU2GE6_0(.din(w_dff_B_m95GODcv4_0),.dout(w_dff_B_kKkyU2GE6_0),.clk(gclk));
	jdff dff_B_MNnsejKZ3_1(.din(n1337),.dout(w_dff_B_MNnsejKZ3_1),.clk(gclk));
	jdff dff_B_AeVhvwdi6_1(.din(w_dff_B_MNnsejKZ3_1),.dout(w_dff_B_AeVhvwdi6_1),.clk(gclk));
	jdff dff_B_OXiC4uOZ9_1(.din(w_dff_B_AeVhvwdi6_1),.dout(w_dff_B_OXiC4uOZ9_1),.clk(gclk));
	jdff dff_B_K95d2xDO4_1(.din(n1338),.dout(w_dff_B_K95d2xDO4_1),.clk(gclk));
	jdff dff_B_n5d7e1jm1_1(.din(w_dff_B_K95d2xDO4_1),.dout(w_dff_B_n5d7e1jm1_1),.clk(gclk));
	jdff dff_B_8iWpoCgo4_1(.din(w_dff_B_n5d7e1jm1_1),.dout(w_dff_B_8iWpoCgo4_1),.clk(gclk));
	jdff dff_B_cMeKLzGs4_0(.din(n1352),.dout(w_dff_B_cMeKLzGs4_0),.clk(gclk));
	jdff dff_B_geTJlya88_0(.din(w_dff_B_cMeKLzGs4_0),.dout(w_dff_B_geTJlya88_0),.clk(gclk));
	jdff dff_B_2f6GBAe88_0(.din(w_dff_B_geTJlya88_0),.dout(w_dff_B_2f6GBAe88_0),.clk(gclk));
	jdff dff_B_YIasQm2p8_0(.din(G174),.dout(w_dff_B_YIasQm2p8_0),.clk(gclk));
	jdff dff_B_L2o6AYYH5_0(.din(G173),.dout(w_dff_B_L2o6AYYH5_0),.clk(gclk));
	jdff dff_B_6oUft6vE8_0(.din(G176),.dout(w_dff_B_6oUft6vE8_0),.clk(gclk));
	jdff dff_B_RzSElG5A5_0(.din(G175),.dout(w_dff_B_RzSElG5A5_0),.clk(gclk));
	jdff dff_B_89KUHvEO0_0(.din(n753),.dout(w_dff_B_89KUHvEO0_0),.clk(gclk));
	jdff dff_B_S4p4rGHS7_0(.din(G177),.dout(w_dff_B_S4p4rGHS7_0),.clk(gclk));
	jdff dff_B_QPrMLEMA6_0(.din(n743),.dout(w_dff_B_QPrMLEMA6_0),.clk(gclk));
	jdff dff_B_pSeVm3Mk5_0(.din(n729),.dout(w_dff_B_pSeVm3Mk5_0),.clk(gclk));
	jdff dff_A_tL4pS8RP3_0(.dout(w_n737_0[0]),.din(w_dff_A_tL4pS8RP3_0),.clk(gclk));
	jdff dff_B_ymWx1Ohc5_0(.din(n736),.dout(w_dff_B_ymWx1Ohc5_0),.clk(gclk));
	jdff dff_B_EQiSFkrb1_1(.din(n1311),.dout(w_dff_B_EQiSFkrb1_1),.clk(gclk));
	jdff dff_B_jGiJQ0wV2_1(.din(w_dff_B_EQiSFkrb1_1),.dout(w_dff_B_jGiJQ0wV2_1),.clk(gclk));
	jdff dff_B_p992Tqr93_1(.din(n1326),.dout(w_dff_B_p992Tqr93_1),.clk(gclk));
	jdff dff_B_MovuNc1j0_1(.din(w_dff_B_p992Tqr93_1),.dout(w_dff_B_MovuNc1j0_1),.clk(gclk));
	jdff dff_B_dmVOihU45_1(.din(n1327),.dout(w_dff_B_dmVOihU45_1),.clk(gclk));
	jdff dff_B_pyGI4mB35_0(.din(n1324),.dout(w_dff_B_pyGI4mB35_0),.clk(gclk));
	jdff dff_B_TQzO71He6_0(.din(n1323),.dout(w_dff_B_TQzO71He6_0),.clk(gclk));
	jdff dff_B_yqqpsv4E3_0(.din(n907),.dout(w_dff_B_yqqpsv4E3_0),.clk(gclk));
	jdff dff_B_oaivzYWu2_0(.din(w_dff_B_yqqpsv4E3_0),.dout(w_dff_B_oaivzYWu2_0),.clk(gclk));
	jdff dff_B_O0Vd6TmT8_0(.din(n944),.dout(w_dff_B_O0Vd6TmT8_0),.clk(gclk));
	jdff dff_B_KEa91tD61_0(.din(w_dff_B_O0Vd6TmT8_0),.dout(w_dff_B_KEa91tD61_0),.clk(gclk));
	jdff dff_B_mbOqfH1Y6_0(.din(n926),.dout(w_dff_B_mbOqfH1Y6_0),.clk(gclk));
	jdff dff_B_BrXuCZOI4_0(.din(w_dff_B_mbOqfH1Y6_0),.dout(w_dff_B_BrXuCZOI4_0),.clk(gclk));
	jdff dff_B_bYbZRTHw0_0(.din(n915),.dout(w_dff_B_bYbZRTHw0_0),.clk(gclk));
	jdff dff_B_l4rg2tHX6_0(.din(w_dff_B_bYbZRTHw0_0),.dout(w_dff_B_l4rg2tHX6_0),.clk(gclk));
	jdff dff_B_f4DIV2E73_1(.din(n1313),.dout(w_dff_B_f4DIV2E73_1),.clk(gclk));
	jdff dff_B_aYGp1ZGM9_1(.din(w_dff_B_f4DIV2E73_1),.dout(w_dff_B_aYGp1ZGM9_1),.clk(gclk));
	jdff dff_B_1bITEiIi8_1(.din(w_dff_B_aYGp1ZGM9_1),.dout(w_dff_B_1bITEiIi8_1),.clk(gclk));
	jdff dff_B_fbU8G7Lj5_0(.din(n898),.dout(w_dff_B_fbU8G7Lj5_0),.clk(gclk));
	jdff dff_B_tmteiliS8_0(.din(w_dff_B_fbU8G7Lj5_0),.dout(w_dff_B_tmteiliS8_0),.clk(gclk));
	jdff dff_A_cGZBiJwI7_1(.dout(w_n891_0[1]),.din(w_dff_A_cGZBiJwI7_1),.clk(gclk));
	jdff dff_B_SoIl8LzQ8_0(.din(n890),.dout(w_dff_B_SoIl8LzQ8_0),.clk(gclk));
	jdff dff_B_y2lQnTGk1_0(.din(n877),.dout(w_dff_B_y2lQnTGk1_0),.clk(gclk));
	jdff dff_B_DeWSW7nC9_0(.din(w_dff_B_y2lQnTGk1_0),.dout(w_dff_B_DeWSW7nC9_0),.clk(gclk));
	jdff dff_B_fQnMEHd96_0(.din(n1312),.dout(w_dff_B_fQnMEHd96_0),.clk(gclk));
	jdff dff_B_3kyWkG664_0(.din(G44),.dout(w_dff_B_3kyWkG664_0),.clk(gclk));
	jdff dff_B_dahXD1oR3_0(.din(n1308),.dout(w_dff_B_dahXD1oR3_0),.clk(gclk));
	jdff dff_B_jPTP5tlu9_0(.din(w_dff_B_dahXD1oR3_0),.dout(w_dff_B_jPTP5tlu9_0),.clk(gclk));
	jdff dff_B_VrqhbXKF4_0(.din(n842),.dout(w_dff_B_VrqhbXKF4_0),.clk(gclk));
	jdff dff_B_HOoNpVCD2_0(.din(n811),.dout(w_dff_B_HOoNpVCD2_0),.clk(gclk));
	jdff dff_B_KyMlupGs9_0(.din(n826),.dout(w_dff_B_KyMlupGs9_0),.clk(gclk));
	jdff dff_B_XSsA1Wql7_0(.din(n818),.dout(w_dff_B_XSsA1Wql7_0),.clk(gclk));
	jdff dff_B_lOMOsdSt8_0(.din(n1302),.dout(w_dff_B_lOMOsdSt8_0),.clk(gclk));
	jdff dff_B_PWdaVupe0_0(.din(G115),.dout(w_dff_B_PWdaVupe0_0),.clk(gclk));
	jdff dff_A_Hqdbi7JV4_1(.dout(w_n1301_0[1]),.din(w_dff_A_Hqdbi7JV4_1),.clk(gclk));
	jdff dff_B_0CT38OSx1_0(.din(n803),.dout(w_dff_B_0CT38OSx1_0),.clk(gclk));
	jdff dff_B_54cKlWns1_0(.din(n796),.dout(w_dff_B_54cKlWns1_0),.clk(gclk));
	jdff dff_B_PST0blmv8_0(.din(n789),.dout(w_dff_B_PST0blmv8_0),.clk(gclk));
	jdff dff_B_CXnBBQwP6_0(.din(n783),.dout(w_dff_B_CXnBBQwP6_0),.clk(gclk));
	jdff dff_A_48ZOUHfV8_0(.dout(w_n851_0[0]),.din(w_dff_A_48ZOUHfV8_0),.clk(gclk));
	jdff dff_A_CwlY1HgX1_0(.dout(w_dff_A_48ZOUHfV8_0),.din(w_dff_A_CwlY1HgX1_0),.clk(gclk));
	jdff dff_B_Wf7nYgeZ5_0(.din(n850),.dout(w_dff_B_Wf7nYgeZ5_0),.clk(gclk));
	jdff dff_B_q7BVBUQk7_1(.din(n1288),.dout(w_dff_B_q7BVBUQk7_1),.clk(gclk));
	jdff dff_B_nrWiBURo9_0(.din(n1295),.dout(w_dff_B_nrWiBURo9_0),.clk(gclk));
	jdff dff_B_EqwYgOAb4_0(.din(w_dff_B_nrWiBURo9_0),.dout(w_dff_B_EqwYgOAb4_0),.clk(gclk));
	jdff dff_B_NZouYTI96_0(.din(n1294),.dout(w_dff_B_NZouYTI96_0),.clk(gclk));
	jdff dff_B_sSfu5jc82_0(.din(w_dff_B_NZouYTI96_0),.dout(w_dff_B_sSfu5jc82_0),.clk(gclk));
	jdff dff_A_ETdALzzl9_2(.dout(w_G18_22[2]),.din(w_dff_A_ETdALzzl9_2),.clk(gclk));
	jdff dff_A_jvMIQD1H6_2(.dout(w_dff_A_ETdALzzl9_2),.din(w_dff_A_jvMIQD1H6_2),.clk(gclk));
	jdff dff_A_IHi45kUJ0_0(.dout(w_n1095_0[0]),.din(w_dff_A_IHi45kUJ0_0),.clk(gclk));
	jdff dff_A_jdynXXo00_0(.dout(w_dff_A_IHi45kUJ0_0),.din(w_dff_A_jdynXXo00_0),.clk(gclk));
	jdff dff_B_P7acJj6O5_0(.din(G168),.dout(w_dff_B_P7acJj6O5_0),.clk(gclk));
	jdff dff_A_z9rFL9Qs7_0(.dout(w_n1076_0[0]),.din(w_dff_A_z9rFL9Qs7_0),.clk(gclk));
	jdff dff_A_l1Fd4mzB7_0(.dout(w_dff_A_z9rFL9Qs7_0),.din(w_dff_A_l1Fd4mzB7_0),.clk(gclk));
	jdff dff_B_go3tZ8237_0(.din(G169),.dout(w_dff_B_go3tZ8237_0),.clk(gclk));
	jdff dff_A_eOGCc9MY9_0(.dout(w_n565_4[0]),.din(w_dff_A_eOGCc9MY9_0),.clk(gclk));
	jdff dff_A_xmqyPieu1_1(.dout(w_n565_4[1]),.din(w_dff_A_xmqyPieu1_1),.clk(gclk));
	jdff dff_B_SaZRZ3eC7_1(.din(n1280),.dout(w_dff_B_SaZRZ3eC7_1),.clk(gclk));
	jdff dff_B_BBcmIffi9_0(.din(G166),.dout(w_dff_B_BBcmIffi9_0),.clk(gclk));
	jdff dff_A_DPI265385_0(.dout(w_n1061_0[0]),.din(w_dff_A_DPI265385_0),.clk(gclk));
	jdff dff_B_wyRCCiEu4_0(.din(G167),.dout(w_dff_B_wyRCCiEu4_0),.clk(gclk));
	jdff dff_A_mVf8HqKT3_0(.dout(w_G414_0),.din(w_dff_A_mVf8HqKT3_0),.clk(gclk));
	jdff dff_A_Rudi88Ma5_0(.dout(w_dff_A_mVf8HqKT3_0),.din(w_dff_A_Rudi88Ma5_0),.clk(gclk));
	jdff dff_A_3oTeT6Q66_0(.dout(w_dff_A_Rudi88Ma5_0),.din(w_dff_A_3oTeT6Q66_0),.clk(gclk));
	jdff dff_B_MoBmqS1O8_1(.din(n1227),.dout(w_dff_B_MoBmqS1O8_1),.clk(gclk));
	jdff dff_B_XgTx141R4_1(.din(w_dff_B_MoBmqS1O8_1),.dout(w_dff_B_XgTx141R4_1),.clk(gclk));
	jdff dff_B_eKyjidAx3_0(.din(n1273),.dout(w_dff_B_eKyjidAx3_0),.clk(gclk));
	jdff dff_B_tHgUzJFw0_0(.din(n740),.dout(w_dff_B_tHgUzJFw0_0),.clk(gclk));
	jdff dff_B_5Z0ZvisL2_0(.din(n733),.dout(w_dff_B_5Z0ZvisL2_0),.clk(gclk));
	jdff dff_B_AtF61fDY2_1(.din(n1270),.dout(w_dff_B_AtF61fDY2_1),.clk(gclk));
	jdff dff_B_FCQlh5Dj1_0(.din(n757),.dout(w_dff_B_FCQlh5Dj1_0),.clk(gclk));
	jdff dff_B_ImjzZV4d2_0(.din(n747),.dout(w_dff_B_ImjzZV4d2_0),.clk(gclk));
	jdff dff_A_hwfUxLGL7_1(.dout(w_G2208_0[1]),.din(w_dff_A_hwfUxLGL7_1),.clk(gclk));
	jdff dff_B_Dv298iPP6_0(.din(n1018),.dout(w_dff_B_Dv298iPP6_0),.clk(gclk));
	jdff dff_B_a2d6WJsL9_0(.din(n1012),.dout(w_dff_B_a2d6WJsL9_0),.clk(gclk));
	jdff dff_B_JiLRwsqs5_0(.din(n998),.dout(w_dff_B_JiLRwsqs5_0),.clk(gclk));
	jdff dff_B_k7lL40703_0(.din(n991),.dout(w_dff_B_k7lL40703_0),.clk(gclk));
	jdff dff_A_HTROHZQK8_0(.dout(w_n727_0[0]),.din(w_dff_A_HTROHZQK8_0),.clk(gclk));
	jdff dff_A_fbjRGt6H7_0(.dout(w_dff_A_HTROHZQK8_0),.din(w_dff_A_fbjRGt6H7_0),.clk(gclk));
	jdff dff_B_k7AAB8Kr6_0(.din(n726),.dout(w_dff_B_k7AAB8Kr6_0),.clk(gclk));
	jdff dff_B_G3fOBOAh3_1(.din(n1253),.dout(w_dff_B_G3fOBOAh3_1),.clk(gclk));
	jdff dff_B_aSMhC8VD8_0(.din(n1260),.dout(w_dff_B_aSMhC8VD8_0),.clk(gclk));
	jdff dff_B_MZwE7jgl3_0(.din(w_dff_B_aSMhC8VD8_0),.dout(w_dff_B_MZwE7jgl3_0),.clk(gclk));
	jdff dff_B_rcYx8yKf4_0(.din(n1099),.dout(w_dff_B_rcYx8yKf4_0),.clk(gclk));
	jdff dff_A_dYIGB10U4_0(.dout(w_G18_23[0]),.din(w_dff_A_dYIGB10U4_0),.clk(gclk));
	jdff dff_B_0yBXJo9z0_0(.din(n1072),.dout(w_dff_B_0yBXJo9z0_0),.clk(gclk));
	jdff dff_A_Uh6msUUb7_0(.dout(w_n1066_0[0]),.din(w_dff_A_Uh6msUUb7_0),.clk(gclk));
	jdff dff_B_L7t6hzka9_0(.din(n1065),.dout(w_dff_B_L7t6hzka9_0),.clk(gclk));
	jdff dff_B_H2CRhkLX8_1(.din(n1251),.dout(w_dff_B_H2CRhkLX8_1),.clk(gclk));
	jdff dff_B_ji1kzFuV4_0(.din(n1085),.dout(w_dff_B_ji1kzFuV4_0),.clk(gclk));
	jdff dff_B_eTd8rISp4_0(.din(n1080),.dout(w_dff_B_eTd8rISp4_0),.clk(gclk));
	jdff dff_A_xh58VgyV7_1(.dout(w_G1459_0[1]),.din(w_dff_A_xh58VgyV7_1),.clk(gclk));
	jdff dff_B_GwnOSJim7_1(.din(n1237),.dout(w_dff_B_GwnOSJim7_1),.clk(gclk));
	jdff dff_B_1lI4iuCx7_1(.din(w_dff_B_GwnOSJim7_1),.dout(w_dff_B_1lI4iuCx7_1),.clk(gclk));
	jdff dff_B_vQSB5hO77_1(.din(n1238),.dout(w_dff_B_vQSB5hO77_1),.clk(gclk));
	jdff dff_B_QHRDrX0e1_1(.din(w_dff_B_vQSB5hO77_1),.dout(w_dff_B_QHRDrX0e1_1),.clk(gclk));
	jdff dff_B_ovWBiHve8_1(.din(n1239),.dout(w_dff_B_ovWBiHve8_1),.clk(gclk));
	jdff dff_A_ABytohFn0_1(.dout(w_n902_0[1]),.din(w_dff_A_ABytohFn0_1),.clk(gclk));
	jdff dff_A_Voxo0vv56_2(.dout(w_n902_0[2]),.din(w_dff_A_Voxo0vv56_2),.clk(gclk));
	jdff dff_B_v0d9Pcq65_1(.din(n900),.dout(w_dff_B_v0d9Pcq65_1),.clk(gclk));
	jdff dff_B_RvBlhviK6_1(.din(n892),.dout(w_dff_B_RvBlhviK6_1),.clk(gclk));
	jdff dff_A_kfTwIkQA1_1(.dout(w_n882_0[1]),.din(w_dff_A_kfTwIkQA1_1),.clk(gclk));
	jdff dff_A_wlzDAiYg7_2(.dout(w_n882_0[2]),.din(w_dff_A_wlzDAiYg7_2),.clk(gclk));
	jdff dff_B_O5SW7v0n6_1(.din(n879),.dout(w_dff_B_O5SW7v0n6_1),.clk(gclk));
	jdff dff_A_kZe7phSE5_1(.dout(w_n873_0[1]),.din(w_dff_A_kZe7phSE5_1),.clk(gclk));
	jdff dff_A_q50Fv1v73_2(.dout(w_n873_0[2]),.din(w_dff_A_q50Fv1v73_2),.clk(gclk));
	jdff dff_B_NDxgaqFP7_1(.din(n870),.dout(w_dff_B_NDxgaqFP7_1),.clk(gclk));
	jdff dff_A_ENCyuXag9_1(.dout(w_n920_0[1]),.din(w_dff_A_ENCyuXag9_1),.clk(gclk));
	jdff dff_A_2yNquiOy5_2(.dout(w_n920_0[2]),.din(w_dff_A_2yNquiOy5_2),.clk(gclk));
	jdff dff_B_fGFTF0XU1_1(.din(n917),.dout(w_dff_B_fGFTF0XU1_1),.clk(gclk));
	jdff dff_A_SZuNFr1P2_0(.dout(w_n948_0[0]),.din(w_dff_A_SZuNFr1P2_0),.clk(gclk));
	jdff dff_A_4oRPwfXE4_2(.dout(w_n948_0[2]),.din(w_dff_A_4oRPwfXE4_2),.clk(gclk));
	jdff dff_B_pi3wdSqF9_1(.din(n946),.dout(w_dff_B_pi3wdSqF9_1),.clk(gclk));
	jdff dff_A_OL2RzQCe5_1(.dout(w_n931_0[1]),.din(w_dff_A_OL2RzQCe5_1),.clk(gclk));
	jdff dff_A_GNJJtZnm1_2(.dout(w_n931_0[2]),.din(w_dff_A_GNJJtZnm1_2),.clk(gclk));
	jdff dff_B_NrCPywIU0_1(.din(n928),.dout(w_dff_B_NrCPywIU0_1),.clk(gclk));
	jdff dff_A_JJ89itmx3_0(.dout(w_n1236_0[0]),.din(w_dff_A_JJ89itmx3_0),.clk(gclk));
	jdff dff_A_iQkRFewx6_0(.dout(w_dff_A_JJ89itmx3_0),.din(w_dff_A_iQkRFewx6_0),.clk(gclk));
	jdff dff_A_dHpbrnif0_1(.dout(w_G3698_0[1]),.din(w_dff_A_dHpbrnif0_1),.clk(gclk));
	jdff dff_B_iLWJF1Hp3_3(.din(n912),.dout(w_dff_B_iLWJF1Hp3_3),.clk(gclk));
	jdff dff_B_NUpiunu24_1(.din(n909),.dout(w_dff_B_NUpiunu24_1),.clk(gclk));
	jdff dff_B_a4N3anBT4_1(.din(n1215),.dout(w_dff_B_a4N3anBT4_1),.clk(gclk));
	jdff dff_B_aLvfeHDS9_1(.din(w_dff_B_a4N3anBT4_1),.dout(w_dff_B_aLvfeHDS9_1),.clk(gclk));
	jdff dff_B_5vCkOg337_1(.din(w_dff_B_aLvfeHDS9_1),.dout(w_dff_B_5vCkOg337_1),.clk(gclk));
	jdff dff_B_qk2e6yzr7_1(.din(n1217),.dout(w_dff_B_qk2e6yzr7_1),.clk(gclk));
	jdff dff_B_763OWH5q8_0(.din(n1224),.dout(w_dff_B_763OWH5q8_0),.clk(gclk));
	jdff dff_B_FXgMXwFy3_0(.din(w_dff_B_763OWH5q8_0),.dout(w_dff_B_FXgMXwFy3_0),.clk(gclk));
	jdff dff_A_l640jkIo4_1(.dout(w_G4393_0[1]),.din(w_dff_A_l640jkIo4_1),.clk(gclk));
	jdff dff_A_I9KtYtk61_1(.dout(w_n355_10[1]),.din(w_dff_A_I9KtYtk61_1),.clk(gclk));
	jdff dff_B_6iLd3lGi5_1(.din(n805),.dout(w_dff_B_6iLd3lGi5_1),.clk(gclk));
	jdff dff_B_9UIE7en39_1(.din(n798),.dout(w_dff_B_9UIE7en39_1),.clk(gclk));
	jdff dff_B_iKVVTLIe3_1(.din(n791),.dout(w_dff_B_iKVVTLIe3_1),.clk(gclk));
	jdff dff_B_gMghVbHt7_1(.din(n785),.dout(w_dff_B_gMghVbHt7_1),.clk(gclk));
	jdff dff_B_U64D73rS2_1(.din(n844),.dout(w_dff_B_U64D73rS2_1),.clk(gclk));
	jdff dff_B_ME82u0P10_1(.din(n813),.dout(w_dff_B_ME82u0P10_1),.clk(gclk));
	jdff dff_A_CC1cSYvL9_0(.dout(w_n855_0[0]),.din(w_dff_A_CC1cSYvL9_0),.clk(gclk));
	jdff dff_B_8ePvQrtz7_1(.din(n852),.dout(w_dff_B_8ePvQrtz7_1),.clk(gclk));
	jdff dff_B_AUOibp789_1(.din(n828),.dout(w_dff_B_AUOibp789_1),.clk(gclk));
	jdff dff_B_llGRv8mi5_1(.din(n820),.dout(w_dff_B_llGRv8mi5_1),.clk(gclk));
	jdff dff_B_IdjBLrfV7_3(.din(n720),.dout(w_dff_B_IdjBLrfV7_3),.clk(gclk));
	jdff dff_B_9BfjA4og5_3(.din(w_dff_B_IdjBLrfV7_3),.dout(w_dff_B_9BfjA4og5_3),.clk(gclk));
	jdff dff_B_pLPjMUlg0_3(.din(w_dff_B_9BfjA4og5_3),.dout(w_dff_B_pLPjMUlg0_3),.clk(gclk));
	jdff dff_B_XBuut1l53_3(.din(w_dff_B_pLPjMUlg0_3),.dout(w_dff_B_XBuut1l53_3),.clk(gclk));
	jdff dff_B_o7C5KK9Q1_3(.din(w_dff_B_XBuut1l53_3),.dout(w_dff_B_o7C5KK9Q1_3),.clk(gclk));
	jdff dff_B_EJ1wzUhh8_3(.din(w_dff_B_o7C5KK9Q1_3),.dout(w_dff_B_EJ1wzUhh8_3),.clk(gclk));
	jdff dff_B_rhc9L5xJ1_3(.din(w_dff_B_EJ1wzUhh8_3),.dout(w_dff_B_rhc9L5xJ1_3),.clk(gclk));
	jdff dff_B_npBiyaxb7_3(.din(w_dff_B_rhc9L5xJ1_3),.dout(w_dff_B_npBiyaxb7_3),.clk(gclk));
	jdff dff_B_y0O2kR962_3(.din(w_dff_B_npBiyaxb7_3),.dout(w_dff_B_y0O2kR962_3),.clk(gclk));
	jdff dff_B_MnsduYnO8_3(.din(w_dff_B_y0O2kR962_3),.dout(w_dff_B_MnsduYnO8_3),.clk(gclk));
	jdff dff_B_8sbhzKj90_3(.din(w_dff_B_MnsduYnO8_3),.dout(w_dff_B_8sbhzKj90_3),.clk(gclk));
	jdff dff_B_O3qcBfn54_3(.din(w_dff_B_8sbhzKj90_3),.dout(w_dff_B_O3qcBfn54_3),.clk(gclk));
	jdff dff_B_0N8uFRUA7_3(.din(w_dff_B_O3qcBfn54_3),.dout(w_dff_B_0N8uFRUA7_3),.clk(gclk));
	jdff dff_B_rMlRfwdG0_3(.din(w_dff_B_0N8uFRUA7_3),.dout(w_dff_B_rMlRfwdG0_3),.clk(gclk));
	jdff dff_B_0giEvvrD3_3(.din(w_dff_B_rMlRfwdG0_3),.dout(w_dff_B_0giEvvrD3_3),.clk(gclk));
	jdff dff_B_tMqqm3EM5_3(.din(w_dff_B_0giEvvrD3_3),.dout(w_dff_B_tMqqm3EM5_3),.clk(gclk));
	jdff dff_B_mCDgaTCp3_3(.din(w_dff_B_tMqqm3EM5_3),.dout(w_dff_B_mCDgaTCp3_3),.clk(gclk));
	jdff dff_B_Nlr6LKx27_3(.din(w_dff_B_mCDgaTCp3_3),.dout(w_dff_B_Nlr6LKx27_3),.clk(gclk));
	jdff dff_B_wwhembUv9_3(.din(w_dff_B_Nlr6LKx27_3),.dout(w_dff_B_wwhembUv9_3),.clk(gclk));
	jdff dff_B_bzIU7bhA5_3(.din(w_dff_B_wwhembUv9_3),.dout(w_dff_B_bzIU7bhA5_3),.clk(gclk));
	jdff dff_B_ZKPdG3yj8_3(.din(w_dff_B_bzIU7bhA5_3),.dout(w_dff_B_ZKPdG3yj8_3),.clk(gclk));
	jdff dff_B_x019fOFD0_1(.din(n717),.dout(w_dff_B_x019fOFD0_1),.clk(gclk));
	jdff dff_B_DJUXuzfR5_1(.din(n1451),.dout(w_dff_B_DJUXuzfR5_1),.clk(gclk));
	jdff dff_B_2NR1HArv1_1(.din(w_dff_B_DJUXuzfR5_1),.dout(w_dff_B_2NR1HArv1_1),.clk(gclk));
	jdff dff_B_fDvnNcQc3_1(.din(w_dff_B_2NR1HArv1_1),.dout(w_dff_B_fDvnNcQc3_1),.clk(gclk));
	jdff dff_B_x56lNv725_1(.din(w_dff_B_fDvnNcQc3_1),.dout(w_dff_B_x56lNv725_1),.clk(gclk));
	jdff dff_B_RdsBE9xP4_1(.din(w_dff_B_x56lNv725_1),.dout(w_dff_B_RdsBE9xP4_1),.clk(gclk));
	jdff dff_B_XO3NzWg02_1(.din(w_dff_B_RdsBE9xP4_1),.dout(w_dff_B_XO3NzWg02_1),.clk(gclk));
	jdff dff_B_8iUwmmxU1_1(.din(w_dff_B_XO3NzWg02_1),.dout(w_dff_B_8iUwmmxU1_1),.clk(gclk));
	jdff dff_B_8w6Ejsrg6_1(.din(w_dff_B_8iUwmmxU1_1),.dout(w_dff_B_8w6Ejsrg6_1),.clk(gclk));
	jdff dff_B_8E6Si50q8_1(.din(w_dff_B_8w6Ejsrg6_1),.dout(w_dff_B_8E6Si50q8_1),.clk(gclk));
	jdff dff_B_SWHMzrLs6_1(.din(w_dff_B_8E6Si50q8_1),.dout(w_dff_B_SWHMzrLs6_1),.clk(gclk));
	jdff dff_B_h37MDbom1_1(.din(w_dff_B_SWHMzrLs6_1),.dout(w_dff_B_h37MDbom1_1),.clk(gclk));
	jdff dff_B_Gwax1Gzy7_1(.din(w_dff_B_h37MDbom1_1),.dout(w_dff_B_Gwax1Gzy7_1),.clk(gclk));
	jdff dff_B_YR4BPWLM1_1(.din(w_dff_B_Gwax1Gzy7_1),.dout(w_dff_B_YR4BPWLM1_1),.clk(gclk));
	jdff dff_B_qW4ciP0a2_1(.din(w_dff_B_YR4BPWLM1_1),.dout(w_dff_B_qW4ciP0a2_1),.clk(gclk));
	jdff dff_B_hvcuFbb39_1(.din(w_dff_B_qW4ciP0a2_1),.dout(w_dff_B_hvcuFbb39_1),.clk(gclk));
	jdff dff_A_QFVvSBXs1_0(.dout(w_n715_0[0]),.din(w_dff_A_QFVvSBXs1_0),.clk(gclk));
	jdff dff_A_ovTq2xU49_1(.dout(w_n715_0[1]),.din(w_dff_A_ovTq2xU49_1),.clk(gclk));
	jdff dff_A_Ckj1AOyH1_0(.dout(w_n1469_0[0]),.din(w_dff_A_Ckj1AOyH1_0),.clk(gclk));
	jdff dff_B_TOpau3XT3_2(.din(n1469),.dout(w_dff_B_TOpau3XT3_2),.clk(gclk));
	jdff dff_B_ATBd61GY6_2(.din(w_dff_B_TOpau3XT3_2),.dout(w_dff_B_ATBd61GY6_2),.clk(gclk));
	jdff dff_B_Mkym6Kci4_2(.din(w_dff_B_ATBd61GY6_2),.dout(w_dff_B_Mkym6Kci4_2),.clk(gclk));
	jdff dff_B_UiM5x9MF9_2(.din(w_dff_B_Mkym6Kci4_2),.dout(w_dff_B_UiM5x9MF9_2),.clk(gclk));
	jdff dff_B_yo0imXru5_2(.din(w_dff_B_UiM5x9MF9_2),.dout(w_dff_B_yo0imXru5_2),.clk(gclk));
	jdff dff_B_7qFPsQRP3_2(.din(w_dff_B_yo0imXru5_2),.dout(w_dff_B_7qFPsQRP3_2),.clk(gclk));
	jdff dff_B_Jcbt0k3I2_2(.din(w_dff_B_7qFPsQRP3_2),.dout(w_dff_B_Jcbt0k3I2_2),.clk(gclk));
	jdff dff_B_5sZLto4h2_2(.din(w_dff_B_Jcbt0k3I2_2),.dout(w_dff_B_5sZLto4h2_2),.clk(gclk));
	jdff dff_B_La9vFLI37_2(.din(w_dff_B_5sZLto4h2_2),.dout(w_dff_B_La9vFLI37_2),.clk(gclk));
	jdff dff_A_cJhQqle97_0(.dout(w_n1470_0[0]),.din(w_dff_A_cJhQqle97_0),.clk(gclk));
	jdff dff_B_LkdWkJ8g7_2(.din(n1470),.dout(w_dff_B_LkdWkJ8g7_2),.clk(gclk));
	jdff dff_B_1gkzg7R10_2(.din(w_dff_B_LkdWkJ8g7_2),.dout(w_dff_B_1gkzg7R10_2),.clk(gclk));
	jdff dff_B_b4mHv3Ng6_2(.din(w_dff_B_1gkzg7R10_2),.dout(w_dff_B_b4mHv3Ng6_2),.clk(gclk));
	jdff dff_B_1Kmi0HtZ6_2(.din(w_dff_B_b4mHv3Ng6_2),.dout(w_dff_B_1Kmi0HtZ6_2),.clk(gclk));
	jdff dff_B_1Kw8nNbx2_2(.din(w_dff_B_1Kmi0HtZ6_2),.dout(w_dff_B_1Kw8nNbx2_2),.clk(gclk));
	jdff dff_B_llMY8War6_2(.din(w_dff_B_1Kw8nNbx2_2),.dout(w_dff_B_llMY8War6_2),.clk(gclk));
	jdff dff_B_KKg45cXB6_2(.din(w_dff_B_llMY8War6_2),.dout(w_dff_B_KKg45cXB6_2),.clk(gclk));
	jdff dff_B_7PTogLGb4_1(.din(n1500),.dout(w_dff_B_7PTogLGb4_1),.clk(gclk));
	jdff dff_B_jXVjhxPA7_1(.din(w_dff_B_7PTogLGb4_1),.dout(w_dff_B_jXVjhxPA7_1),.clk(gclk));
	jdff dff_B_B0jVdQZK5_1(.din(w_dff_B_jXVjhxPA7_1),.dout(w_dff_B_B0jVdQZK5_1),.clk(gclk));
	jdff dff_B_HMC3Mo6w6_1(.din(w_dff_B_B0jVdQZK5_1),.dout(w_dff_B_HMC3Mo6w6_1),.clk(gclk));
	jdff dff_B_GZoZRhPB5_1(.din(w_dff_B_HMC3Mo6w6_1),.dout(w_dff_B_GZoZRhPB5_1),.clk(gclk));
	jdff dff_B_zCZ1gWyq6_1(.din(w_dff_B_GZoZRhPB5_1),.dout(w_dff_B_zCZ1gWyq6_1),.clk(gclk));
	jdff dff_B_MAfprkEt8_1(.din(w_dff_B_zCZ1gWyq6_1),.dout(w_dff_B_MAfprkEt8_1),.clk(gclk));
	jdff dff_B_AzlUtPke4_1(.din(w_dff_B_MAfprkEt8_1),.dout(w_dff_B_AzlUtPke4_1),.clk(gclk));
	jdff dff_B_TwUTlE3B4_1(.din(w_dff_B_AzlUtPke4_1),.dout(w_dff_B_TwUTlE3B4_1),.clk(gclk));
	jdff dff_B_tYZ2TMyR3_1(.din(w_dff_B_TwUTlE3B4_1),.dout(w_dff_B_tYZ2TMyR3_1),.clk(gclk));
	jdff dff_B_PPbMZT6d2_1(.din(w_dff_B_tYZ2TMyR3_1),.dout(w_dff_B_PPbMZT6d2_1),.clk(gclk));
	jdff dff_B_FLUsvZJe6_1(.din(w_dff_B_PPbMZT6d2_1),.dout(w_dff_B_FLUsvZJe6_1),.clk(gclk));
	jdff dff_B_7es6Sl7R1_1(.din(w_dff_B_FLUsvZJe6_1),.dout(w_dff_B_7es6Sl7R1_1),.clk(gclk));
	jdff dff_B_L0aE1pJH9_1(.din(w_dff_B_7es6Sl7R1_1),.dout(w_dff_B_L0aE1pJH9_1),.clk(gclk));
	jdff dff_B_mt6EQCSe3_1(.din(w_dff_B_L0aE1pJH9_1),.dout(w_dff_B_mt6EQCSe3_1),.clk(gclk));
	jdff dff_B_xkiUoI6d8_0(.din(n1546),.dout(w_dff_B_xkiUoI6d8_0),.clk(gclk));
	jdff dff_B_mAKxwxqz1_0(.din(w_dff_B_xkiUoI6d8_0),.dout(w_dff_B_mAKxwxqz1_0),.clk(gclk));
	jdff dff_B_fGAAYMSZ9_0(.din(n1544),.dout(w_dff_B_fGAAYMSZ9_0),.clk(gclk));
	jdff dff_B_RDwCv1ed2_0(.din(w_dff_B_fGAAYMSZ9_0),.dout(w_dff_B_RDwCv1ed2_0),.clk(gclk));
	jdff dff_B_eATi8HMD6_1(.din(n1533),.dout(w_dff_B_eATi8HMD6_1),.clk(gclk));
	jdff dff_B_oj7vR2wc0_1(.din(w_dff_B_eATi8HMD6_1),.dout(w_dff_B_oj7vR2wc0_1),.clk(gclk));
	jdff dff_B_25NFH76a5_1(.din(w_dff_B_oj7vR2wc0_1),.dout(w_dff_B_25NFH76a5_1),.clk(gclk));
	jdff dff_B_2ZeCTHMn8_1(.din(w_dff_B_25NFH76a5_1),.dout(w_dff_B_2ZeCTHMn8_1),.clk(gclk));
	jdff dff_B_k7HXkkHM6_1(.din(n1534),.dout(w_dff_B_k7HXkkHM6_1),.clk(gclk));
	jdff dff_B_wUzjKcsA2_1(.din(w_dff_B_k7HXkkHM6_1),.dout(w_dff_B_wUzjKcsA2_1),.clk(gclk));
	jdff dff_B_XvPI7GAs4_1(.din(w_dff_B_wUzjKcsA2_1),.dout(w_dff_B_XvPI7GAs4_1),.clk(gclk));
	jdff dff_B_pnT5QBZn4_1(.din(w_dff_B_XvPI7GAs4_1),.dout(w_dff_B_pnT5QBZn4_1),.clk(gclk));
	jdff dff_B_WA4gBXwc1_1(.din(w_dff_B_pnT5QBZn4_1),.dout(w_dff_B_WA4gBXwc1_1),.clk(gclk));
	jdff dff_B_nQNILQLi0_1(.din(w_dff_B_WA4gBXwc1_1),.dout(w_dff_B_nQNILQLi0_1),.clk(gclk));
	jdff dff_B_m54To6v88_1(.din(w_dff_B_nQNILQLi0_1),.dout(w_dff_B_m54To6v88_1),.clk(gclk));
	jdff dff_B_wa7J2Vx24_1(.din(n1538),.dout(w_dff_B_wa7J2Vx24_1),.clk(gclk));
	jdff dff_B_47O9ffhk8_0(.din(n1540),.dout(w_dff_B_47O9ffhk8_0),.clk(gclk));
	jdff dff_B_H19Doc6T6_1(.din(n1539),.dout(w_dff_B_H19Doc6T6_1),.clk(gclk));
	jdff dff_B_pkJzjAA13_0(.din(n1535),.dout(w_dff_B_pkJzjAA13_0),.clk(gclk));
	jdff dff_A_0RAVFEVr1_1(.dout(w_n1414_0[1]),.din(w_dff_A_0RAVFEVr1_1),.clk(gclk));
	jdff dff_A_eOyVXiE77_1(.dout(w_dff_A_0RAVFEVr1_1),.din(w_dff_A_eOyVXiE77_1),.clk(gclk));
	jdff dff_A_b8zTXIi13_1(.dout(w_dff_A_eOyVXiE77_1),.din(w_dff_A_b8zTXIi13_1),.clk(gclk));
	jdff dff_A_sRXZ4qhC5_1(.dout(w_dff_A_b8zTXIi13_1),.din(w_dff_A_sRXZ4qhC5_1),.clk(gclk));
	jdff dff_A_Kpy41kBj3_1(.dout(w_dff_A_sRXZ4qhC5_1),.din(w_dff_A_Kpy41kBj3_1),.clk(gclk));
	jdff dff_A_xghiZztM6_1(.dout(w_dff_A_Kpy41kBj3_1),.din(w_dff_A_xghiZztM6_1),.clk(gclk));
	jdff dff_A_5uPzxucX4_1(.dout(w_dff_A_xghiZztM6_1),.din(w_dff_A_5uPzxucX4_1),.clk(gclk));
	jdff dff_A_IW5KJ3Dj5_1(.dout(w_dff_A_5uPzxucX4_1),.din(w_dff_A_IW5KJ3Dj5_1),.clk(gclk));
	jdff dff_A_WBXkA0S14_1(.dout(w_dff_A_IW5KJ3Dj5_1),.din(w_dff_A_WBXkA0S14_1),.clk(gclk));
	jdff dff_A_mxJkPqv15_1(.dout(w_dff_A_WBXkA0S14_1),.din(w_dff_A_mxJkPqv15_1),.clk(gclk));
	jdff dff_B_bMdm3kIy3_1(.din(n1412),.dout(w_dff_B_bMdm3kIy3_1),.clk(gclk));
	jdff dff_A_Q4G3Vr6v2_1(.dout(w_n1404_0[1]),.din(w_dff_A_Q4G3Vr6v2_1),.clk(gclk));
	jdff dff_A_5cF9i9ps0_1(.dout(w_dff_A_Q4G3Vr6v2_1),.din(w_dff_A_5cF9i9ps0_1),.clk(gclk));
	jdff dff_A_Fg0GymQ76_1(.dout(w_dff_A_5cF9i9ps0_1),.din(w_dff_A_Fg0GymQ76_1),.clk(gclk));
	jdff dff_A_jPMQ1vXE5_1(.dout(w_dff_A_Fg0GymQ76_1),.din(w_dff_A_jPMQ1vXE5_1),.clk(gclk));
	jdff dff_A_20vVuD9A2_1(.dout(w_dff_A_jPMQ1vXE5_1),.din(w_dff_A_20vVuD9A2_1),.clk(gclk));
	jdff dff_A_HLu4tZgU8_1(.dout(w_dff_A_20vVuD9A2_1),.din(w_dff_A_HLu4tZgU8_1),.clk(gclk));
	jdff dff_A_45Mf1pPl0_1(.dout(w_dff_A_HLu4tZgU8_1),.din(w_dff_A_45Mf1pPl0_1),.clk(gclk));
	jdff dff_A_LUAz2R5u7_1(.dout(w_dff_A_45Mf1pPl0_1),.din(w_dff_A_LUAz2R5u7_1),.clk(gclk));
	jdff dff_A_jOasjh7M6_1(.dout(w_dff_A_LUAz2R5u7_1),.din(w_dff_A_jOasjh7M6_1),.clk(gclk));
	jdff dff_B_pNqP6SDG5_2(.din(n1404),.dout(w_dff_B_pNqP6SDG5_2),.clk(gclk));
	jdff dff_B_vAm4i5Er2_0(.din(n1530),.dout(w_dff_B_vAm4i5Er2_0),.clk(gclk));
	jdff dff_B_VZarvOZq4_0(.din(w_dff_B_vAm4i5Er2_0),.dout(w_dff_B_VZarvOZq4_0),.clk(gclk));
	jdff dff_B_1sUUPRfg5_0(.din(w_dff_B_VZarvOZq4_0),.dout(w_dff_B_1sUUPRfg5_0),.clk(gclk));
	jdff dff_B_OJow9Vyl2_1(.din(n1524),.dout(w_dff_B_OJow9Vyl2_1),.clk(gclk));
	jdff dff_B_U1goTxm30_1(.din(w_dff_B_OJow9Vyl2_1),.dout(w_dff_B_U1goTxm30_1),.clk(gclk));
	jdff dff_B_QDq6Jaas7_0(.din(n1527),.dout(w_dff_B_QDq6Jaas7_0),.clk(gclk));
	jdff dff_B_ordt9V3h7_0(.din(w_dff_B_QDq6Jaas7_0),.dout(w_dff_B_ordt9V3h7_0),.clk(gclk));
	jdff dff_B_jAFUiruS4_0(.din(w_dff_B_ordt9V3h7_0),.dout(w_dff_B_jAFUiruS4_0),.clk(gclk));
	jdff dff_B_N6gXHevE0_1(.din(n1525),.dout(w_dff_B_N6gXHevE0_1),.clk(gclk));
	jdff dff_A_FzYkVwt71_1(.dout(w_n1401_0[1]),.din(w_dff_A_FzYkVwt71_1),.clk(gclk));
	jdff dff_A_Xm39ijup5_1(.dout(w_dff_A_FzYkVwt71_1),.din(w_dff_A_Xm39ijup5_1),.clk(gclk));
	jdff dff_A_KQjVIlGn5_1(.dout(w_dff_A_Xm39ijup5_1),.din(w_dff_A_KQjVIlGn5_1),.clk(gclk));
	jdff dff_A_4ys7vwfR2_1(.dout(w_dff_A_KQjVIlGn5_1),.din(w_dff_A_4ys7vwfR2_1),.clk(gclk));
	jdff dff_A_3TleVXER0_1(.dout(w_dff_A_4ys7vwfR2_1),.din(w_dff_A_3TleVXER0_1),.clk(gclk));
	jdff dff_A_Apm4yrQa9_1(.dout(w_dff_A_3TleVXER0_1),.din(w_dff_A_Apm4yrQa9_1),.clk(gclk));
	jdff dff_A_H1VOLBDP6_1(.dout(w_dff_A_Apm4yrQa9_1),.din(w_dff_A_H1VOLBDP6_1),.clk(gclk));
	jdff dff_A_hBqkJqjS1_1(.dout(w_dff_A_H1VOLBDP6_1),.din(w_dff_A_hBqkJqjS1_1),.clk(gclk));
	jdff dff_A_ZmUqUEXr6_1(.dout(w_dff_A_hBqkJqjS1_1),.din(w_dff_A_ZmUqUEXr6_1),.clk(gclk));
	jdff dff_B_tlAcGgC34_2(.din(n1401),.dout(w_dff_B_tlAcGgC34_2),.clk(gclk));
	jdff dff_B_YXY9vh597_2(.din(w_dff_B_tlAcGgC34_2),.dout(w_dff_B_YXY9vh597_2),.clk(gclk));
	jdff dff_B_uiMlzBmr5_2(.din(w_dff_B_YXY9vh597_2),.dout(w_dff_B_uiMlzBmr5_2),.clk(gclk));
	jdff dff_B_mBMAvR3y5_2(.din(w_dff_B_uiMlzBmr5_2),.dout(w_dff_B_mBMAvR3y5_2),.clk(gclk));
	jdff dff_B_QqnObltz0_2(.din(w_dff_B_mBMAvR3y5_2),.dout(w_dff_B_QqnObltz0_2),.clk(gclk));
	jdff dff_B_Ypk94iqM7_2(.din(w_dff_B_QqnObltz0_2),.dout(w_dff_B_Ypk94iqM7_2),.clk(gclk));
	jdff dff_A_trCzAZP81_1(.dout(w_n1520_0[1]),.din(w_dff_A_trCzAZP81_1),.clk(gclk));
	jdff dff_B_XX0mknTh8_0(.din(n1516),.dout(w_dff_B_XX0mknTh8_0),.clk(gclk));
	jdff dff_B_Z4uhcWtN0_0(.din(w_dff_B_XX0mknTh8_0),.dout(w_dff_B_Z4uhcWtN0_0),.clk(gclk));
	jdff dff_B_TymWwy7E5_0(.din(w_dff_B_Z4uhcWtN0_0),.dout(w_dff_B_TymWwy7E5_0),.clk(gclk));
	jdff dff_B_Qbdzpj2C1_0(.din(w_dff_B_TymWwy7E5_0),.dout(w_dff_B_Qbdzpj2C1_0),.clk(gclk));
	jdff dff_B_eiKQTK2w9_0(.din(w_dff_B_Qbdzpj2C1_0),.dout(w_dff_B_eiKQTK2w9_0),.clk(gclk));
	jdff dff_B_ztIY41Q55_1(.din(n1509),.dout(w_dff_B_ztIY41Q55_1),.clk(gclk));
	jdff dff_B_rbiPKVwW4_1(.din(w_dff_B_ztIY41Q55_1),.dout(w_dff_B_rbiPKVwW4_1),.clk(gclk));
	jdff dff_B_XiJPqNd82_1(.din(w_dff_B_rbiPKVwW4_1),.dout(w_dff_B_XiJPqNd82_1),.clk(gclk));
	jdff dff_B_ra5xCKJj3_1(.din(w_dff_B_XiJPqNd82_1),.dout(w_dff_B_ra5xCKJj3_1),.clk(gclk));
	jdff dff_B_whGYmxuB1_1(.din(w_dff_B_ra5xCKJj3_1),.dout(w_dff_B_whGYmxuB1_1),.clk(gclk));
	jdff dff_B_1qVDS2KB7_1(.din(w_dff_B_whGYmxuB1_1),.dout(w_dff_B_1qVDS2KB7_1),.clk(gclk));
	jdff dff_B_rzNwJKfw7_0(.din(n1513),.dout(w_dff_B_rzNwJKfw7_0),.clk(gclk));
	jdff dff_A_RMpuFhPp5_1(.dout(w_n1445_0[1]),.din(w_dff_A_RMpuFhPp5_1),.clk(gclk));
	jdff dff_A_p5TL9DJ66_1(.dout(w_dff_A_RMpuFhPp5_1),.din(w_dff_A_p5TL9DJ66_1),.clk(gclk));
	jdff dff_A_PKoctAc01_1(.dout(w_dff_A_p5TL9DJ66_1),.din(w_dff_A_PKoctAc01_1),.clk(gclk));
	jdff dff_A_yukqebI99_1(.dout(w_dff_A_PKoctAc01_1),.din(w_dff_A_yukqebI99_1),.clk(gclk));
	jdff dff_A_YQ5Y2fgs9_1(.dout(w_dff_A_yukqebI99_1),.din(w_dff_A_YQ5Y2fgs9_1),.clk(gclk));
	jdff dff_A_ZWcRm7Km3_1(.dout(w_dff_A_YQ5Y2fgs9_1),.din(w_dff_A_ZWcRm7Km3_1),.clk(gclk));
	jdff dff_A_IlyOiMQ73_1(.dout(w_dff_A_ZWcRm7Km3_1),.din(w_dff_A_IlyOiMQ73_1),.clk(gclk));
	jdff dff_A_w4QdJfPC3_1(.dout(w_dff_A_IlyOiMQ73_1),.din(w_dff_A_w4QdJfPC3_1),.clk(gclk));
	jdff dff_A_oGuhTOFj2_1(.dout(w_dff_A_w4QdJfPC3_1),.din(w_dff_A_oGuhTOFj2_1),.clk(gclk));
	jdff dff_A_ILt6LRmd0_1(.dout(w_dff_A_oGuhTOFj2_1),.din(w_dff_A_ILt6LRmd0_1),.clk(gclk));
	jdff dff_A_sXuwNK8R4_1(.dout(w_dff_A_ILt6LRmd0_1),.din(w_dff_A_sXuwNK8R4_1),.clk(gclk));
	jdff dff_B_oKWTF6hl0_2(.din(n1445),.dout(w_dff_B_oKWTF6hl0_2),.clk(gclk));
	jdff dff_B_FE7WUiIF0_0(.din(n1507),.dout(w_dff_B_FE7WUiIF0_0),.clk(gclk));
	jdff dff_B_idJEKtUL7_0(.din(w_dff_B_FE7WUiIF0_0),.dout(w_dff_B_idJEKtUL7_0),.clk(gclk));
	jdff dff_B_jtp16RiP5_0(.din(w_dff_B_idJEKtUL7_0),.dout(w_dff_B_jtp16RiP5_0),.clk(gclk));
	jdff dff_B_s88beJ2U6_0(.din(w_dff_B_jtp16RiP5_0),.dout(w_dff_B_s88beJ2U6_0),.clk(gclk));
	jdff dff_B_b5nqAN7c3_0(.din(w_dff_B_s88beJ2U6_0),.dout(w_dff_B_b5nqAN7c3_0),.clk(gclk));
	jdff dff_B_yIW1yNUH0_0(.din(w_dff_B_b5nqAN7c3_0),.dout(w_dff_B_yIW1yNUH0_0),.clk(gclk));
	jdff dff_B_GRpJRWRw0_0(.din(n1503),.dout(w_dff_B_GRpJRWRw0_0),.clk(gclk));
	jdff dff_A_OZfn1ucS1_0(.dout(w_n1444_0[0]),.din(w_dff_A_OZfn1ucS1_0),.clk(gclk));
	jdff dff_A_TA0aTwIG6_0(.dout(w_dff_A_OZfn1ucS1_0),.din(w_dff_A_TA0aTwIG6_0),.clk(gclk));
	jdff dff_A_XrdWwc4R2_2(.dout(w_n1444_0[2]),.din(w_dff_A_XrdWwc4R2_2),.clk(gclk));
	jdff dff_A_JoHABMJ87_2(.dout(w_dff_A_XrdWwc4R2_2),.din(w_dff_A_JoHABMJ87_2),.clk(gclk));
	jdff dff_A_zWjy8oUP2_2(.dout(w_dff_A_JoHABMJ87_2),.din(w_dff_A_zWjy8oUP2_2),.clk(gclk));
	jdff dff_A_8cwtMwTA2_2(.dout(w_dff_A_zWjy8oUP2_2),.din(w_dff_A_8cwtMwTA2_2),.clk(gclk));
	jdff dff_A_8qFpqZGO9_2(.dout(w_dff_A_8cwtMwTA2_2),.din(w_dff_A_8qFpqZGO9_2),.clk(gclk));
	jdff dff_A_HINHVoHg8_2(.dout(w_dff_A_8qFpqZGO9_2),.din(w_dff_A_HINHVoHg8_2),.clk(gclk));
	jdff dff_A_lI3gZliT6_2(.dout(w_dff_A_HINHVoHg8_2),.din(w_dff_A_lI3gZliT6_2),.clk(gclk));
	jdff dff_A_bJzo3sLd7_2(.dout(w_dff_A_lI3gZliT6_2),.din(w_dff_A_bJzo3sLd7_2),.clk(gclk));
	jdff dff_A_A17pJVNn5_2(.dout(w_dff_A_bJzo3sLd7_2),.din(w_dff_A_A17pJVNn5_2),.clk(gclk));
	jdff dff_A_uL5Vjebj3_2(.dout(w_dff_A_A17pJVNn5_2),.din(w_dff_A_uL5Vjebj3_2),.clk(gclk));
	jdff dff_A_RijIaEAN0_2(.dout(w_dff_A_uL5Vjebj3_2),.din(w_dff_A_RijIaEAN0_2),.clk(gclk));
	jdff dff_A_s0GIDYHk9_2(.dout(w_dff_A_RijIaEAN0_2),.din(w_dff_A_s0GIDYHk9_2),.clk(gclk));
	jdff dff_A_W0oVwpZc9_2(.dout(w_dff_A_s0GIDYHk9_2),.din(w_dff_A_W0oVwpZc9_2),.clk(gclk));
	jdff dff_B_qnMenjZs7_3(.din(n1444),.dout(w_dff_B_qnMenjZs7_3),.clk(gclk));
	jdff dff_B_8ItX7a3K5_3(.din(w_dff_B_qnMenjZs7_3),.dout(w_dff_B_8ItX7a3K5_3),.clk(gclk));
	jdff dff_B_H6Ftr2x54_3(.din(w_dff_B_8ItX7a3K5_3),.dout(w_dff_B_H6Ftr2x54_3),.clk(gclk));
	jdff dff_B_nLkcjZeK0_3(.din(w_dff_B_H6Ftr2x54_3),.dout(w_dff_B_nLkcjZeK0_3),.clk(gclk));
	jdff dff_A_K8finmwX0_1(.dout(w_n1501_0[1]),.din(w_dff_A_K8finmwX0_1),.clk(gclk));
	jdff dff_A_fCO3Igr54_1(.dout(w_dff_A_K8finmwX0_1),.din(w_dff_A_fCO3Igr54_1),.clk(gclk));
	jdff dff_A_uQPGZkEK6_1(.dout(w_dff_A_fCO3Igr54_1),.din(w_dff_A_uQPGZkEK6_1),.clk(gclk));
	jdff dff_A_s5UHIRKd7_1(.dout(w_dff_A_uQPGZkEK6_1),.din(w_dff_A_s5UHIRKd7_1),.clk(gclk));
	jdff dff_A_YS3sKKuK9_1(.dout(w_dff_A_s5UHIRKd7_1),.din(w_dff_A_YS3sKKuK9_1),.clk(gclk));
	jdff dff_A_dLHHILYu7_1(.dout(w_n1454_0[1]),.din(w_dff_A_dLHHILYu7_1),.clk(gclk));
	jdff dff_A_ZLOlZNlP0_1(.dout(w_dff_A_dLHHILYu7_1),.din(w_dff_A_ZLOlZNlP0_1),.clk(gclk));
	jdff dff_A_uMZQ4TGC6_1(.dout(w_dff_A_ZLOlZNlP0_1),.din(w_dff_A_uMZQ4TGC6_1),.clk(gclk));
	jdff dff_A_aOg9zfBa6_1(.dout(w_dff_A_uMZQ4TGC6_1),.din(w_dff_A_aOg9zfBa6_1),.clk(gclk));
	jdff dff_A_Q9N2VMIL7_1(.dout(w_dff_A_aOg9zfBa6_1),.din(w_dff_A_Q9N2VMIL7_1),.clk(gclk));
	jdff dff_A_tTgmfphQ8_1(.dout(w_dff_A_Q9N2VMIL7_1),.din(w_dff_A_tTgmfphQ8_1),.clk(gclk));
	jdff dff_A_pHdo0g8s9_1(.dout(w_dff_A_tTgmfphQ8_1),.din(w_dff_A_pHdo0g8s9_1),.clk(gclk));
	jdff dff_B_rgXWuGbk1_2(.din(n1454),.dout(w_dff_B_rgXWuGbk1_2),.clk(gclk));
	jdff dff_B_lEOwJkwd9_2(.din(w_dff_B_rgXWuGbk1_2),.dout(w_dff_B_lEOwJkwd9_2),.clk(gclk));
	jdff dff_B_HNfOPdWG3_2(.din(w_dff_B_lEOwJkwd9_2),.dout(w_dff_B_HNfOPdWG3_2),.clk(gclk));
	jdff dff_B_b60A2s786_2(.din(w_dff_B_HNfOPdWG3_2),.dout(w_dff_B_b60A2s786_2),.clk(gclk));
	jdff dff_B_2QcC4uf46_2(.din(w_dff_B_b60A2s786_2),.dout(w_dff_B_2QcC4uf46_2),.clk(gclk));
	jdff dff_B_CPgWZ9vI4_0(.din(n1584),.dout(w_dff_B_CPgWZ9vI4_0),.clk(gclk));
	jdff dff_B_BQKshNcL9_0(.din(w_dff_B_CPgWZ9vI4_0),.dout(w_dff_B_BQKshNcL9_0),.clk(gclk));
	jdff dff_B_L9CTJBsM8_0(.din(w_dff_B_BQKshNcL9_0),.dout(w_dff_B_L9CTJBsM8_0),.clk(gclk));
	jdff dff_B_BT1wfhvp5_1(.din(n1561),.dout(w_dff_B_BT1wfhvp5_1),.clk(gclk));
	jdff dff_B_vRekUBR52_1(.din(w_dff_B_BT1wfhvp5_1),.dout(w_dff_B_vRekUBR52_1),.clk(gclk));
	jdff dff_B_OJFvKyQI8_1(.din(w_dff_B_vRekUBR52_1),.dout(w_dff_B_OJFvKyQI8_1),.clk(gclk));
	jdff dff_B_MDjvm9xl0_1(.din(w_dff_B_OJFvKyQI8_1),.dout(w_dff_B_MDjvm9xl0_1),.clk(gclk));
	jdff dff_B_BFZeTVQt1_1(.din(w_dff_B_MDjvm9xl0_1),.dout(w_dff_B_BFZeTVQt1_1),.clk(gclk));
	jdff dff_B_wbZ2kgpr0_1(.din(w_dff_B_BFZeTVQt1_1),.dout(w_dff_B_wbZ2kgpr0_1),.clk(gclk));
	jdff dff_B_3e994TVL5_1(.din(w_dff_B_wbZ2kgpr0_1),.dout(w_dff_B_3e994TVL5_1),.clk(gclk));
	jdff dff_B_o1ld9FgW2_1(.din(w_dff_B_3e994TVL5_1),.dout(w_dff_B_o1ld9FgW2_1),.clk(gclk));
	jdff dff_B_QwlKy81m2_1(.din(w_dff_B_o1ld9FgW2_1),.dout(w_dff_B_QwlKy81m2_1),.clk(gclk));
	jdff dff_B_Vnhx5BuQ2_1(.din(w_dff_B_QwlKy81m2_1),.dout(w_dff_B_Vnhx5BuQ2_1),.clk(gclk));
	jdff dff_B_S7UP4dzI8_1(.din(w_dff_B_Vnhx5BuQ2_1),.dout(w_dff_B_S7UP4dzI8_1),.clk(gclk));
	jdff dff_B_irgtnqym3_1(.din(w_dff_B_S7UP4dzI8_1),.dout(w_dff_B_irgtnqym3_1),.clk(gclk));
	jdff dff_B_LL0vGEG51_1(.din(w_dff_B_irgtnqym3_1),.dout(w_dff_B_LL0vGEG51_1),.clk(gclk));
	jdff dff_B_KwCLLSB36_1(.din(w_dff_B_LL0vGEG51_1),.dout(w_dff_B_KwCLLSB36_1),.clk(gclk));
	jdff dff_B_4lppfiRp5_1(.din(w_dff_B_KwCLLSB36_1),.dout(w_dff_B_4lppfiRp5_1),.clk(gclk));
	jdff dff_B_GfkogCA50_1(.din(w_dff_B_4lppfiRp5_1),.dout(w_dff_B_GfkogCA50_1),.clk(gclk));
	jdff dff_B_Lun4TgfG5_1(.din(w_dff_B_GfkogCA50_1),.dout(w_dff_B_Lun4TgfG5_1),.clk(gclk));
	jdff dff_B_0JtIXeks0_0(.din(n1581),.dout(w_dff_B_0JtIXeks0_0),.clk(gclk));
	jdff dff_B_gbAOKVfw2_0(.din(w_dff_B_0JtIXeks0_0),.dout(w_dff_B_gbAOKVfw2_0),.clk(gclk));
	jdff dff_B_5Bwc77lF8_0(.din(n1578),.dout(w_dff_B_5Bwc77lF8_0),.clk(gclk));
	jdff dff_B_gdFh1aYu1_0(.din(w_dff_B_5Bwc77lF8_0),.dout(w_dff_B_gdFh1aYu1_0),.clk(gclk));
	jdff dff_B_PV7Z3eCq6_0(.din(w_dff_B_gdFh1aYu1_0),.dout(w_dff_B_PV7Z3eCq6_0),.clk(gclk));
	jdff dff_B_BApgaGwq5_0(.din(w_dff_B_PV7Z3eCq6_0),.dout(w_dff_B_BApgaGwq5_0),.clk(gclk));
	jdff dff_B_l8XTke5Z7_0(.din(w_dff_B_BApgaGwq5_0),.dout(w_dff_B_l8XTke5Z7_0),.clk(gclk));
	jdff dff_B_OAS7MuBZ6_0(.din(w_dff_B_l8XTke5Z7_0),.dout(w_dff_B_OAS7MuBZ6_0),.clk(gclk));
	jdff dff_B_B9JBJ9031_1(.din(n1572),.dout(w_dff_B_B9JBJ9031_1),.clk(gclk));
	jdff dff_B_O7xxMIBe2_1(.din(w_dff_B_B9JBJ9031_1),.dout(w_dff_B_O7xxMIBe2_1),.clk(gclk));
	jdff dff_B_SdDV3byI7_1(.din(w_dff_B_O7xxMIBe2_1),.dout(w_dff_B_SdDV3byI7_1),.clk(gclk));
	jdff dff_B_iEA9xJDk0_0(.din(n1574),.dout(w_dff_B_iEA9xJDk0_0),.clk(gclk));
	jdff dff_B_Cta6HihX1_0(.din(n1570),.dout(w_dff_B_Cta6HihX1_0),.clk(gclk));
	jdff dff_B_2rjMd3se2_0(.din(w_dff_B_Cta6HihX1_0),.dout(w_dff_B_2rjMd3se2_0),.clk(gclk));
	jdff dff_B_I7zxjpBj9_0(.din(n1568),.dout(w_dff_B_I7zxjpBj9_0),.clk(gclk));
	jdff dff_B_7shGJBdY2_0(.din(w_dff_B_I7zxjpBj9_0),.dout(w_dff_B_7shGJBdY2_0),.clk(gclk));
	jdff dff_B_5J46EBdU9_0(.din(w_dff_B_7shGJBdY2_0),.dout(w_dff_B_5J46EBdU9_0),.clk(gclk));
	jdff dff_B_ugAVC3ph0_0(.din(w_dff_B_5J46EBdU9_0),.dout(w_dff_B_ugAVC3ph0_0),.clk(gclk));
	jdff dff_B_kr5Q7uVQ5_0(.din(w_dff_B_ugAVC3ph0_0),.dout(w_dff_B_kr5Q7uVQ5_0),.clk(gclk));
	jdff dff_B_CVGMQyU47_0(.din(w_dff_B_kr5Q7uVQ5_0),.dout(w_dff_B_CVGMQyU47_0),.clk(gclk));
	jdff dff_B_X2z5vmO42_0(.din(n1567),.dout(w_dff_B_X2z5vmO42_0),.clk(gclk));
	jdff dff_B_9NmeohgU2_0(.din(w_dff_B_X2z5vmO42_0),.dout(w_dff_B_9NmeohgU2_0),.clk(gclk));
	jdff dff_B_290SYT7O3_0(.din(w_dff_B_9NmeohgU2_0),.dout(w_dff_B_290SYT7O3_0),.clk(gclk));
	jdff dff_B_IVsL0sZo9_0(.din(w_dff_B_290SYT7O3_0),.dout(w_dff_B_IVsL0sZo9_0),.clk(gclk));
	jdff dff_B_l8UL9uop4_0(.din(w_dff_B_IVsL0sZo9_0),.dout(w_dff_B_l8UL9uop4_0),.clk(gclk));
	jdff dff_B_B3GFjWaI7_0(.din(n1566),.dout(w_dff_B_B3GFjWaI7_0),.clk(gclk));
	jdff dff_B_JG5CIk200_0(.din(w_dff_B_B3GFjWaI7_0),.dout(w_dff_B_JG5CIk200_0),.clk(gclk));
	jdff dff_B_4pwTS0wB0_0(.din(n1562),.dout(w_dff_B_4pwTS0wB0_0),.clk(gclk));
	jdff dff_A_nDaZdZov6_1(.dout(w_n1420_0[1]),.din(w_dff_A_nDaZdZov6_1),.clk(gclk));
	jdff dff_A_rcujZ2oE8_1(.dout(w_dff_A_nDaZdZov6_1),.din(w_dff_A_rcujZ2oE8_1),.clk(gclk));
	jdff dff_A_I42mvFI97_1(.dout(w_dff_A_rcujZ2oE8_1),.din(w_dff_A_I42mvFI97_1),.clk(gclk));
	jdff dff_A_UQBvNC652_1(.dout(w_dff_A_I42mvFI97_1),.din(w_dff_A_UQBvNC652_1),.clk(gclk));
	jdff dff_A_JuciOKGi8_2(.dout(w_n1420_0[2]),.din(w_dff_A_JuciOKGi8_2),.clk(gclk));
	jdff dff_A_pxZtaReL0_2(.dout(w_dff_A_JuciOKGi8_2),.din(w_dff_A_pxZtaReL0_2),.clk(gclk));
	jdff dff_A_477LDJ4G8_2(.dout(w_dff_A_pxZtaReL0_2),.din(w_dff_A_477LDJ4G8_2),.clk(gclk));
	jdff dff_A_NWEkugVQ3_2(.dout(w_dff_A_477LDJ4G8_2),.din(w_dff_A_NWEkugVQ3_2),.clk(gclk));
	jdff dff_A_wRe8lVGu0_2(.dout(w_dff_A_NWEkugVQ3_2),.din(w_dff_A_wRe8lVGu0_2),.clk(gclk));
	jdff dff_A_dVAfYEhO8_2(.dout(w_dff_A_wRe8lVGu0_2),.din(w_dff_A_dVAfYEhO8_2),.clk(gclk));
	jdff dff_A_gUPPNxoU6_2(.dout(w_dff_A_dVAfYEhO8_2),.din(w_dff_A_gUPPNxoU6_2),.clk(gclk));
	jdff dff_A_STqZxIi20_2(.dout(w_dff_A_gUPPNxoU6_2),.din(w_dff_A_STqZxIi20_2),.clk(gclk));
	jdff dff_A_y0JqANA15_2(.dout(w_dff_A_STqZxIi20_2),.din(w_dff_A_y0JqANA15_2),.clk(gclk));
	jdff dff_A_mtZqKfHV3_2(.dout(w_dff_A_y0JqANA15_2),.din(w_dff_A_mtZqKfHV3_2),.clk(gclk));
	jdff dff_A_fzW89w8z8_2(.dout(w_dff_A_mtZqKfHV3_2),.din(w_dff_A_fzW89w8z8_2),.clk(gclk));
	jdff dff_A_57MW5ouo1_2(.dout(w_dff_A_fzW89w8z8_2),.din(w_dff_A_57MW5ouo1_2),.clk(gclk));
	jdff dff_A_VfDUbObf6_2(.dout(w_dff_A_57MW5ouo1_2),.din(w_dff_A_VfDUbObf6_2),.clk(gclk));
	jdff dff_A_su9DqBxa6_2(.dout(w_dff_A_VfDUbObf6_2),.din(w_dff_A_su9DqBxa6_2),.clk(gclk));
	jdff dff_A_Y7WKfHCC6_2(.dout(w_dff_A_su9DqBxa6_2),.din(w_dff_A_Y7WKfHCC6_2),.clk(gclk));
	jdff dff_A_9egDAeHd7_2(.dout(w_dff_A_Y7WKfHCC6_2),.din(w_dff_A_9egDAeHd7_2),.clk(gclk));
	jdff dff_B_m5hw7YnI1_3(.din(n1420),.dout(w_dff_B_m5hw7YnI1_3),.clk(gclk));
	jdff dff_B_1enUmcj93_3(.din(w_dff_B_m5hw7YnI1_3),.dout(w_dff_B_1enUmcj93_3),.clk(gclk));
	jdff dff_B_jbCKAF4M3_3(.din(w_dff_B_1enUmcj93_3),.dout(w_dff_B_jbCKAF4M3_3),.clk(gclk));
	jdff dff_B_qbRnz3Ku9_0(.din(n1559),.dout(w_dff_B_qbRnz3Ku9_0),.clk(gclk));
	jdff dff_B_rdIMQoTt5_0(.din(w_dff_B_qbRnz3Ku9_0),.dout(w_dff_B_rdIMQoTt5_0),.clk(gclk));
	jdff dff_B_7vykC2Sy8_0(.din(w_dff_B_rdIMQoTt5_0),.dout(w_dff_B_7vykC2Sy8_0),.clk(gclk));
	jdff dff_B_Id4qsDKp8_0(.din(w_dff_B_7vykC2Sy8_0),.dout(w_dff_B_Id4qsDKp8_0),.clk(gclk));
	jdff dff_B_0CS3cZfD4_0(.din(n1558),.dout(w_dff_B_0CS3cZfD4_0),.clk(gclk));
	jdff dff_B_EP5t6Ueb1_0(.din(w_dff_B_0CS3cZfD4_0),.dout(w_dff_B_EP5t6Ueb1_0),.clk(gclk));
	jdff dff_B_cyiGqZzo3_0(.din(w_dff_B_EP5t6Ueb1_0),.dout(w_dff_B_cyiGqZzo3_0),.clk(gclk));
	jdff dff_B_3ZnM1Mw94_0(.din(w_dff_B_cyiGqZzo3_0),.dout(w_dff_B_3ZnM1Mw94_0),.clk(gclk));
	jdff dff_B_yfGAFMFW6_0(.din(n1556),.dout(w_dff_B_yfGAFMFW6_0),.clk(gclk));
	jdff dff_B_FOWnRYgm5_0(.din(n1554),.dout(w_dff_B_FOWnRYgm5_0),.clk(gclk));
	jdff dff_B_UmDUmI8U8_0(.din(w_dff_B_FOWnRYgm5_0),.dout(w_dff_B_UmDUmI8U8_0),.clk(gclk));
	jdff dff_B_8aGUcFe22_0(.din(w_dff_B_UmDUmI8U8_0),.dout(w_dff_B_8aGUcFe22_0),.clk(gclk));
	jdff dff_A_AdRreLLg7_1(.dout(w_n1464_0[1]),.din(w_dff_A_AdRreLLg7_1),.clk(gclk));
	jdff dff_A_T4VSx2Fc3_1(.dout(w_dff_A_AdRreLLg7_1),.din(w_dff_A_T4VSx2Fc3_1),.clk(gclk));
	jdff dff_A_Os34ysUw2_1(.dout(w_dff_A_T4VSx2Fc3_1),.din(w_dff_A_Os34ysUw2_1),.clk(gclk));
	jdff dff_A_cntpAp7F7_1(.dout(w_dff_A_Os34ysUw2_1),.din(w_dff_A_cntpAp7F7_1),.clk(gclk));
	jdff dff_A_umttXLsx6_1(.dout(w_dff_A_cntpAp7F7_1),.din(w_dff_A_umttXLsx6_1),.clk(gclk));
	jdff dff_A_78EKFMid6_1(.dout(w_dff_A_umttXLsx6_1),.din(w_dff_A_78EKFMid6_1),.clk(gclk));
	jdff dff_A_YE6unQTE1_1(.dout(w_dff_A_78EKFMid6_1),.din(w_dff_A_YE6unQTE1_1),.clk(gclk));
	jdff dff_B_mE4r2VJp7_2(.din(n1464),.dout(w_dff_B_mE4r2VJp7_2),.clk(gclk));
	jdff dff_B_7JCPp54f4_2(.din(w_dff_B_mE4r2VJp7_2),.dout(w_dff_B_7JCPp54f4_2),.clk(gclk));
	jdff dff_B_TpvOAebs8_2(.din(w_dff_B_7JCPp54f4_2),.dout(w_dff_B_TpvOAebs8_2),.clk(gclk));
	jdff dff_B_ae0WsQPs3_2(.din(w_dff_B_TpvOAebs8_2),.dout(w_dff_B_ae0WsQPs3_2),.clk(gclk));
	jdff dff_B_2hCUtnVv2_2(.din(w_dff_B_ae0WsQPs3_2),.dout(w_dff_B_2hCUtnVv2_2),.clk(gclk));
	jdff dff_B_7LQryvWr4_2(.din(w_dff_B_2hCUtnVv2_2),.dout(w_dff_B_7LQryvWr4_2),.clk(gclk));
	jdff dff_B_jU9Y2Liy2_2(.din(w_dff_B_7LQryvWr4_2),.dout(w_dff_B_jU9Y2Liy2_2),.clk(gclk));
	jdff dff_B_jyPnGC367_2(.din(w_dff_B_jU9Y2Liy2_2),.dout(w_dff_B_jyPnGC367_2),.clk(gclk));
	jdff dff_B_8kfqkchA5_2(.din(w_dff_B_jyPnGC367_2),.dout(w_dff_B_8kfqkchA5_2),.clk(gclk));
	jdff dff_B_slQaUEwN2_2(.din(w_dff_B_8kfqkchA5_2),.dout(w_dff_B_slQaUEwN2_2),.clk(gclk));
	jdff dff_B_as9m61SM4_2(.din(w_dff_B_slQaUEwN2_2),.dout(w_dff_B_as9m61SM4_2),.clk(gclk));
	jdff dff_B_TNqvWjH05_2(.din(w_dff_B_as9m61SM4_2),.dout(w_dff_B_TNqvWjH05_2),.clk(gclk));
	jdff dff_B_RNFNZPNZ6_0(.din(n1391),.dout(w_dff_B_RNFNZPNZ6_0),.clk(gclk));
	jdff dff_B_BYgSR66Y5_0(.din(w_dff_B_RNFNZPNZ6_0),.dout(w_dff_B_BYgSR66Y5_0),.clk(gclk));
	jdff dff_B_tnGwUCCF3_0(.din(w_dff_B_BYgSR66Y5_0),.dout(w_dff_B_tnGwUCCF3_0),.clk(gclk));
	jdff dff_B_h774zQpj6_0(.din(w_dff_B_tnGwUCCF3_0),.dout(w_dff_B_h774zQpj6_0),.clk(gclk));
	jdff dff_B_btPUfdhX8_0(.din(w_dff_B_h774zQpj6_0),.dout(w_dff_B_btPUfdhX8_0),.clk(gclk));
	jdff dff_B_5wWHOG5Z8_0(.din(w_dff_B_btPUfdhX8_0),.dout(w_dff_B_5wWHOG5Z8_0),.clk(gclk));
	jdff dff_B_Ipi3dn0D4_0(.din(w_dff_B_5wWHOG5Z8_0),.dout(w_dff_B_Ipi3dn0D4_0),.clk(gclk));
	jdff dff_B_gtNNXPav0_0(.din(w_dff_B_Ipi3dn0D4_0),.dout(w_dff_B_gtNNXPav0_0),.clk(gclk));
	jdff dff_B_oX7W0P6n7_0(.din(n1388),.dout(w_dff_B_oX7W0P6n7_0),.clk(gclk));
	jdff dff_B_aUl8IxEi7_0(.din(w_dff_B_oX7W0P6n7_0),.dout(w_dff_B_aUl8IxEi7_0),.clk(gclk));
	jdff dff_B_ZetI8zSD9_0(.din(w_dff_B_aUl8IxEi7_0),.dout(w_dff_B_ZetI8zSD9_0),.clk(gclk));
	jdff dff_B_UGxZ7lFd5_0(.din(w_dff_B_ZetI8zSD9_0),.dout(w_dff_B_UGxZ7lFd5_0),.clk(gclk));
	jdff dff_B_o3Lxyyui5_3(.din(n713),.dout(w_dff_B_o3Lxyyui5_3),.clk(gclk));
	jdff dff_B_1qJbNLwG1_3(.din(w_dff_B_o3Lxyyui5_3),.dout(w_dff_B_1qJbNLwG1_3),.clk(gclk));
	jdff dff_B_PXk43iGC9_3(.din(w_dff_B_1qJbNLwG1_3),.dout(w_dff_B_PXk43iGC9_3),.clk(gclk));
	jdff dff_B_35fkCRxo0_3(.din(w_dff_B_PXk43iGC9_3),.dout(w_dff_B_35fkCRxo0_3),.clk(gclk));
	jdff dff_B_VeKVQlt00_3(.din(w_dff_B_35fkCRxo0_3),.dout(w_dff_B_VeKVQlt00_3),.clk(gclk));
	jdff dff_B_s2NUqyJr0_3(.din(w_dff_B_VeKVQlt00_3),.dout(w_dff_B_s2NUqyJr0_3),.clk(gclk));
	jdff dff_B_IjYFWwaV1_3(.din(w_dff_B_s2NUqyJr0_3),.dout(w_dff_B_IjYFWwaV1_3),.clk(gclk));
	jdff dff_B_A17VGGhj5_3(.din(w_dff_B_IjYFWwaV1_3),.dout(w_dff_B_A17VGGhj5_3),.clk(gclk));
	jdff dff_B_4mU5CPv50_3(.din(w_dff_B_A17VGGhj5_3),.dout(w_dff_B_4mU5CPv50_3),.clk(gclk));
	jdff dff_B_nrtOx7dN6_3(.din(w_dff_B_4mU5CPv50_3),.dout(w_dff_B_nrtOx7dN6_3),.clk(gclk));
	jdff dff_B_bfeFApFI5_3(.din(w_dff_B_nrtOx7dN6_3),.dout(w_dff_B_bfeFApFI5_3),.clk(gclk));
	jdff dff_B_1TtCNeJd6_3(.din(w_dff_B_bfeFApFI5_3),.dout(w_dff_B_1TtCNeJd6_3),.clk(gclk));
	jdff dff_B_vddRwIyd2_3(.din(w_dff_B_1TtCNeJd6_3),.dout(w_dff_B_vddRwIyd2_3),.clk(gclk));
	jdff dff_B_5jMRDQqI2_3(.din(w_dff_B_vddRwIyd2_3),.dout(w_dff_B_5jMRDQqI2_3),.clk(gclk));
	jdff dff_B_3feuBcIM0_3(.din(w_dff_B_5jMRDQqI2_3),.dout(w_dff_B_3feuBcIM0_3),.clk(gclk));
	jdff dff_B_dX4Zthjp2_3(.din(w_dff_B_3feuBcIM0_3),.dout(w_dff_B_dX4Zthjp2_3),.clk(gclk));
	jdff dff_B_4DpitqpM3_3(.din(w_dff_B_dX4Zthjp2_3),.dout(w_dff_B_4DpitqpM3_3),.clk(gclk));
	jdff dff_B_h5i4nYIP8_3(.din(w_dff_B_4DpitqpM3_3),.dout(w_dff_B_h5i4nYIP8_3),.clk(gclk));
	jdff dff_B_EQWtMFSW0_3(.din(w_dff_B_h5i4nYIP8_3),.dout(w_dff_B_EQWtMFSW0_3),.clk(gclk));
	jdff dff_A_qm3V73ow2_0(.dout(w_n712_0[0]),.din(w_dff_A_qm3V73ow2_0),.clk(gclk));
	jdff dff_A_Tjs7jqik5_0(.dout(w_dff_A_qm3V73ow2_0),.din(w_dff_A_Tjs7jqik5_0),.clk(gclk));
	jdff dff_A_F9HH5xu79_0(.dout(w_dff_A_Tjs7jqik5_0),.din(w_dff_A_F9HH5xu79_0),.clk(gclk));
	jdff dff_A_qRwU4ddM5_0(.dout(w_dff_A_F9HH5xu79_0),.din(w_dff_A_qRwU4ddM5_0),.clk(gclk));
	jdff dff_A_uzrdb2sV6_0(.dout(w_dff_A_qRwU4ddM5_0),.din(w_dff_A_uzrdb2sV6_0),.clk(gclk));
	jdff dff_A_XTJGXc3d5_0(.dout(w_dff_A_uzrdb2sV6_0),.din(w_dff_A_XTJGXc3d5_0),.clk(gclk));
	jdff dff_A_kvAyxm348_0(.dout(w_dff_A_XTJGXc3d5_0),.din(w_dff_A_kvAyxm348_0),.clk(gclk));
	jdff dff_A_IP7mBN9E7_0(.dout(w_dff_A_kvAyxm348_0),.din(w_dff_A_IP7mBN9E7_0),.clk(gclk));
	jdff dff_A_GzFwDnGV1_0(.dout(w_dff_A_IP7mBN9E7_0),.din(w_dff_A_GzFwDnGV1_0),.clk(gclk));
	jdff dff_A_efIUWXha9_0(.dout(w_dff_A_GzFwDnGV1_0),.din(w_dff_A_efIUWXha9_0),.clk(gclk));
	jdff dff_A_i0n28pc09_0(.dout(w_dff_A_efIUWXha9_0),.din(w_dff_A_i0n28pc09_0),.clk(gclk));
	jdff dff_A_Ol78IyE07_0(.dout(w_dff_A_i0n28pc09_0),.din(w_dff_A_Ol78IyE07_0),.clk(gclk));
	jdff dff_A_Pic31c0g9_0(.dout(w_dff_A_Ol78IyE07_0),.din(w_dff_A_Pic31c0g9_0),.clk(gclk));
	jdff dff_A_hFyNf2gp7_0(.dout(w_dff_A_Pic31c0g9_0),.din(w_dff_A_hFyNf2gp7_0),.clk(gclk));
	jdff dff_A_XVbKIfHm6_1(.dout(w_n708_0[1]),.din(w_dff_A_XVbKIfHm6_1),.clk(gclk));
	jdff dff_A_gphEXCPu7_1(.dout(w_dff_A_XVbKIfHm6_1),.din(w_dff_A_gphEXCPu7_1),.clk(gclk));
	jdff dff_A_YtxervhW8_1(.dout(w_dff_A_gphEXCPu7_1),.din(w_dff_A_YtxervhW8_1),.clk(gclk));
	jdff dff_A_0BCslKa28_1(.dout(w_dff_A_YtxervhW8_1),.din(w_dff_A_0BCslKa28_1),.clk(gclk));
	jdff dff_A_sIlKmTIk2_1(.dout(w_dff_A_0BCslKa28_1),.din(w_dff_A_sIlKmTIk2_1),.clk(gclk));
	jdff dff_A_UkuR83006_1(.dout(w_n707_0[1]),.din(w_dff_A_UkuR83006_1),.clk(gclk));
	jdff dff_A_MBQafO8t9_1(.dout(w_dff_A_UkuR83006_1),.din(w_dff_A_MBQafO8t9_1),.clk(gclk));
	jdff dff_A_LaJMjqf63_1(.dout(w_dff_A_MBQafO8t9_1),.din(w_dff_A_LaJMjqf63_1),.clk(gclk));
	jdff dff_A_1Ze5oN6V2_1(.dout(w_dff_A_LaJMjqf63_1),.din(w_dff_A_1Ze5oN6V2_1),.clk(gclk));
	jdff dff_A_CQCZnukW9_1(.dout(w_dff_A_1Ze5oN6V2_1),.din(w_dff_A_CQCZnukW9_1),.clk(gclk));
	jdff dff_B_9zmlM31z8_1(.din(n684),.dout(w_dff_B_9zmlM31z8_1),.clk(gclk));
	jdff dff_B_K5O94ioG0_1(.din(w_dff_B_9zmlM31z8_1),.dout(w_dff_B_K5O94ioG0_1),.clk(gclk));
	jdff dff_B_D0HAbg2r7_1(.din(w_dff_B_K5O94ioG0_1),.dout(w_dff_B_D0HAbg2r7_1),.clk(gclk));
	jdff dff_B_R8fjVUsO4_1(.din(w_dff_B_D0HAbg2r7_1),.dout(w_dff_B_R8fjVUsO4_1),.clk(gclk));
	jdff dff_B_zoj3t5tp7_1(.din(w_dff_B_R8fjVUsO4_1),.dout(w_dff_B_zoj3t5tp7_1),.clk(gclk));
	jdff dff_B_PGSPpr9L6_1(.din(w_dff_B_zoj3t5tp7_1),.dout(w_dff_B_PGSPpr9L6_1),.clk(gclk));
	jdff dff_B_y0AQQQ5r5_1(.din(w_dff_B_PGSPpr9L6_1),.dout(w_dff_B_y0AQQQ5r5_1),.clk(gclk));
	jdff dff_B_cAueN9243_1(.din(w_dff_B_y0AQQQ5r5_1),.dout(w_dff_B_cAueN9243_1),.clk(gclk));
	jdff dff_B_A0nkvEoo2_1(.din(w_dff_B_cAueN9243_1),.dout(w_dff_B_A0nkvEoo2_1),.clk(gclk));
	jdff dff_B_1PVp4q1H5_1(.din(w_dff_B_A0nkvEoo2_1),.dout(w_dff_B_1PVp4q1H5_1),.clk(gclk));
	jdff dff_B_vGa7ZA0O3_1(.din(n685),.dout(w_dff_B_vGa7ZA0O3_1),.clk(gclk));
	jdff dff_B_TdT9F8l34_1(.din(w_dff_B_vGa7ZA0O3_1),.dout(w_dff_B_TdT9F8l34_1),.clk(gclk));
	jdff dff_B_rdUN98LT6_1(.din(w_dff_B_TdT9F8l34_1),.dout(w_dff_B_rdUN98LT6_1),.clk(gclk));
	jdff dff_B_7AlBMn8z4_1(.din(w_dff_B_rdUN98LT6_1),.dout(w_dff_B_7AlBMn8z4_1),.clk(gclk));
	jdff dff_B_Fs1JxQFF8_1(.din(w_dff_B_7AlBMn8z4_1),.dout(w_dff_B_Fs1JxQFF8_1),.clk(gclk));
	jdff dff_B_jzhRgWuO1_1(.din(w_dff_B_Fs1JxQFF8_1),.dout(w_dff_B_jzhRgWuO1_1),.clk(gclk));
	jdff dff_B_BPk0jcx12_1(.din(w_dff_B_jzhRgWuO1_1),.dout(w_dff_B_BPk0jcx12_1),.clk(gclk));
	jdff dff_B_5UKvz1BV5_1(.din(w_dff_B_BPk0jcx12_1),.dout(w_dff_B_5UKvz1BV5_1),.clk(gclk));
	jdff dff_B_SvFmXFXy0_1(.din(w_dff_B_5UKvz1BV5_1),.dout(w_dff_B_SvFmXFXy0_1),.clk(gclk));
	jdff dff_A_IBNlclkX0_0(.dout(w_n704_0[0]),.din(w_dff_A_IBNlclkX0_0),.clk(gclk));
	jdff dff_A_mYqwX8PM9_0(.dout(w_dff_A_IBNlclkX0_0),.din(w_dff_A_mYqwX8PM9_0),.clk(gclk));
	jdff dff_A_YnWSadld2_0(.dout(w_dff_A_mYqwX8PM9_0),.din(w_dff_A_YnWSadld2_0),.clk(gclk));
	jdff dff_A_J0SmL0Lz6_0(.dout(w_dff_A_YnWSadld2_0),.din(w_dff_A_J0SmL0Lz6_0),.clk(gclk));
	jdff dff_A_NpT0gloa1_0(.dout(w_dff_A_J0SmL0Lz6_0),.din(w_dff_A_NpT0gloa1_0),.clk(gclk));
	jdff dff_A_1gR5hOrD4_0(.dout(w_dff_A_NpT0gloa1_0),.din(w_dff_A_1gR5hOrD4_0),.clk(gclk));
	jdff dff_A_9JdlS2n67_0(.dout(w_dff_A_1gR5hOrD4_0),.din(w_dff_A_9JdlS2n67_0),.clk(gclk));
	jdff dff_A_jVAIWxSm1_0(.dout(w_dff_A_9JdlS2n67_0),.din(w_dff_A_jVAIWxSm1_0),.clk(gclk));
	jdff dff_A_d8remCbq1_0(.dout(w_dff_A_jVAIWxSm1_0),.din(w_dff_A_d8remCbq1_0),.clk(gclk));
	jdff dff_A_u4QAVovr0_0(.dout(w_dff_A_d8remCbq1_0),.din(w_dff_A_u4QAVovr0_0),.clk(gclk));
	jdff dff_A_BWxM5W4l6_0(.dout(w_dff_A_u4QAVovr0_0),.din(w_dff_A_BWxM5W4l6_0),.clk(gclk));
	jdff dff_B_scTNcYtf5_1(.din(n688),.dout(w_dff_B_scTNcYtf5_1),.clk(gclk));
	jdff dff_B_D7KAaGaU8_1(.din(w_dff_B_scTNcYtf5_1),.dout(w_dff_B_D7KAaGaU8_1),.clk(gclk));
	jdff dff_B_LFBeO9jF8_1(.din(w_dff_B_D7KAaGaU8_1),.dout(w_dff_B_LFBeO9jF8_1),.clk(gclk));
	jdff dff_B_u7Ko2cDu1_1(.din(w_dff_B_LFBeO9jF8_1),.dout(w_dff_B_u7Ko2cDu1_1),.clk(gclk));
	jdff dff_B_X0nIvMJv5_1(.din(w_dff_B_u7Ko2cDu1_1),.dout(w_dff_B_X0nIvMJv5_1),.clk(gclk));
	jdff dff_B_0VaK6qKA7_1(.din(n689),.dout(w_dff_B_0VaK6qKA7_1),.clk(gclk));
	jdff dff_B_rTyk81Ci5_1(.din(w_dff_B_0VaK6qKA7_1),.dout(w_dff_B_rTyk81Ci5_1),.clk(gclk));
	jdff dff_B_ihuTnrWi8_1(.din(w_dff_B_rTyk81Ci5_1),.dout(w_dff_B_ihuTnrWi8_1),.clk(gclk));
	jdff dff_B_Qe26gSrG6_1(.din(w_dff_B_ihuTnrWi8_1),.dout(w_dff_B_Qe26gSrG6_1),.clk(gclk));
	jdff dff_B_YznDGJU62_0(.din(n698),.dout(w_dff_B_YznDGJU62_0),.clk(gclk));
	jdff dff_A_GAUrzCC51_0(.dout(w_n697_0[0]),.din(w_dff_A_GAUrzCC51_0),.clk(gclk));
	jdff dff_A_ybOcknkA1_0(.dout(w_dff_A_GAUrzCC51_0),.din(w_dff_A_ybOcknkA1_0),.clk(gclk));
	jdff dff_A_8ikj3pmB8_0(.dout(w_dff_A_ybOcknkA1_0),.din(w_dff_A_8ikj3pmB8_0),.clk(gclk));
	jdff dff_A_OB0T8kDx4_0(.dout(w_dff_A_8ikj3pmB8_0),.din(w_dff_A_OB0T8kDx4_0),.clk(gclk));
	jdff dff_A_fDdH1Y1f5_0(.dout(w_dff_A_OB0T8kDx4_0),.din(w_dff_A_fDdH1Y1f5_0),.clk(gclk));
	jdff dff_A_cgqoNBhx2_0(.dout(w_dff_A_fDdH1Y1f5_0),.din(w_dff_A_cgqoNBhx2_0),.clk(gclk));
	jdff dff_A_n7CHZb1D0_0(.dout(w_dff_A_cgqoNBhx2_0),.din(w_dff_A_n7CHZb1D0_0),.clk(gclk));
	jdff dff_A_yv34kAe32_0(.dout(w_dff_A_n7CHZb1D0_0),.din(w_dff_A_yv34kAe32_0),.clk(gclk));
	jdff dff_A_7mL1KvRt6_0(.dout(w_dff_A_yv34kAe32_0),.din(w_dff_A_7mL1KvRt6_0),.clk(gclk));
	jdff dff_A_NCva8RBO6_0(.dout(w_dff_A_7mL1KvRt6_0),.din(w_dff_A_NCva8RBO6_0),.clk(gclk));
	jdff dff_A_vSbt27XT8_0(.dout(w_dff_A_NCva8RBO6_0),.din(w_dff_A_vSbt27XT8_0),.clk(gclk));
	jdff dff_A_hEchCG9b8_0(.dout(w_dff_A_vSbt27XT8_0),.din(w_dff_A_hEchCG9b8_0),.clk(gclk));
	jdff dff_A_fZs2ZWdW2_1(.dout(w_n697_0[1]),.din(w_dff_A_fZs2ZWdW2_1),.clk(gclk));
	jdff dff_A_EX1LRekP0_1(.dout(w_dff_A_fZs2ZWdW2_1),.din(w_dff_A_EX1LRekP0_1),.clk(gclk));
	jdff dff_A_cj3BLgXr6_1(.dout(w_dff_A_EX1LRekP0_1),.din(w_dff_A_cj3BLgXr6_1),.clk(gclk));
	jdff dff_A_SajO6ibN1_1(.dout(w_dff_A_cj3BLgXr6_1),.din(w_dff_A_SajO6ibN1_1),.clk(gclk));
	jdff dff_A_50kmlw7L5_1(.dout(w_dff_A_SajO6ibN1_1),.din(w_dff_A_50kmlw7L5_1),.clk(gclk));
	jdff dff_A_m6X3qeO16_1(.dout(w_dff_A_50kmlw7L5_1),.din(w_dff_A_m6X3qeO16_1),.clk(gclk));
	jdff dff_A_uWFW5vFM3_1(.dout(w_dff_A_m6X3qeO16_1),.din(w_dff_A_uWFW5vFM3_1),.clk(gclk));
	jdff dff_A_6iGsjrnf4_1(.dout(w_dff_A_uWFW5vFM3_1),.din(w_dff_A_6iGsjrnf4_1),.clk(gclk));
	jdff dff_A_kPXeZyBL2_1(.dout(w_dff_A_6iGsjrnf4_1),.din(w_dff_A_kPXeZyBL2_1),.clk(gclk));
	jdff dff_A_Fd6zMXsT1_1(.dout(w_dff_A_kPXeZyBL2_1),.din(w_dff_A_Fd6zMXsT1_1),.clk(gclk));
	jdff dff_A_RCqGhqE04_1(.dout(w_dff_A_Fd6zMXsT1_1),.din(w_dff_A_RCqGhqE04_1),.clk(gclk));
	jdff dff_A_roiBgEmt3_1(.dout(w_dff_A_RCqGhqE04_1),.din(w_dff_A_roiBgEmt3_1),.clk(gclk));
	jdff dff_A_D8HwYQTS2_1(.dout(w_dff_A_roiBgEmt3_1),.din(w_dff_A_D8HwYQTS2_1),.clk(gclk));
	jdff dff_A_EXJ3Ihjh4_1(.dout(w_dff_A_D8HwYQTS2_1),.din(w_dff_A_EXJ3Ihjh4_1),.clk(gclk));
	jdff dff_A_nc8Ki9XG2_1(.dout(w_dff_A_EXJ3Ihjh4_1),.din(w_dff_A_nc8Ki9XG2_1),.clk(gclk));
	jdff dff_A_tYqylR2b8_1(.dout(w_dff_A_nc8Ki9XG2_1),.din(w_dff_A_tYqylR2b8_1),.clk(gclk));
	jdff dff_A_uyp60RjA7_1(.dout(w_dff_A_tYqylR2b8_1),.din(w_dff_A_uyp60RjA7_1),.clk(gclk));
	jdff dff_A_GalQl23S9_1(.dout(w_n692_0[1]),.din(w_dff_A_GalQl23S9_1),.clk(gclk));
	jdff dff_A_alPEdqvK7_1(.dout(w_n687_0[1]),.din(w_dff_A_alPEdqvK7_1),.clk(gclk));
	jdff dff_B_3zMMKSHN0_2(.din(n687),.dout(w_dff_B_3zMMKSHN0_2),.clk(gclk));
	jdff dff_B_YtmsBo2T0_2(.din(w_dff_B_3zMMKSHN0_2),.dout(w_dff_B_YtmsBo2T0_2),.clk(gclk));
	jdff dff_B_VTfTOa1U4_2(.din(w_dff_B_YtmsBo2T0_2),.dout(w_dff_B_VTfTOa1U4_2),.clk(gclk));
	jdff dff_B_wjvOcLtB7_2(.din(w_dff_B_VTfTOa1U4_2),.dout(w_dff_B_wjvOcLtB7_2),.clk(gclk));
	jdff dff_B_JDTa9cxO0_2(.din(w_dff_B_wjvOcLtB7_2),.dout(w_dff_B_JDTa9cxO0_2),.clk(gclk));
	jdff dff_A_ei9GWXxs3_0(.dout(w_n686_0[0]),.din(w_dff_A_ei9GWXxs3_0),.clk(gclk));
	jdff dff_A_wQk6P4as0_0(.dout(w_dff_A_ei9GWXxs3_0),.din(w_dff_A_wQk6P4as0_0),.clk(gclk));
	jdff dff_A_vL3DhvzU0_0(.dout(w_dff_A_wQk6P4as0_0),.din(w_dff_A_vL3DhvzU0_0),.clk(gclk));
	jdff dff_A_WC9bGbaM2_0(.dout(w_dff_A_vL3DhvzU0_0),.din(w_dff_A_WC9bGbaM2_0),.clk(gclk));
	jdff dff_A_JtQI1AOW4_0(.dout(w_dff_A_WC9bGbaM2_0),.din(w_dff_A_JtQI1AOW4_0),.clk(gclk));
	jdff dff_B_hhmIj0YZ6_0(.din(n682),.dout(w_dff_B_hhmIj0YZ6_0),.clk(gclk));
	jdff dff_B_BsDb86gk3_0(.din(w_dff_B_hhmIj0YZ6_0),.dout(w_dff_B_BsDb86gk3_0),.clk(gclk));
	jdff dff_B_M5HAi76b4_0(.din(w_dff_B_BsDb86gk3_0),.dout(w_dff_B_M5HAi76b4_0),.clk(gclk));
	jdff dff_B_lAstQ9Ae1_0(.din(w_dff_B_M5HAi76b4_0),.dout(w_dff_B_lAstQ9Ae1_0),.clk(gclk));
	jdff dff_B_SpmEtieD5_0(.din(w_dff_B_lAstQ9Ae1_0),.dout(w_dff_B_SpmEtieD5_0),.clk(gclk));
	jdff dff_B_bnhpgtgG5_0(.din(w_dff_B_SpmEtieD5_0),.dout(w_dff_B_bnhpgtgG5_0),.clk(gclk));
	jdff dff_B_yzkbhmro8_0(.din(w_dff_B_bnhpgtgG5_0),.dout(w_dff_B_yzkbhmro8_0),.clk(gclk));
	jdff dff_B_FRhg6m2f5_0(.din(w_dff_B_yzkbhmro8_0),.dout(w_dff_B_FRhg6m2f5_0),.clk(gclk));
	jdff dff_B_qwAs0RzU0_0(.din(w_dff_B_FRhg6m2f5_0),.dout(w_dff_B_qwAs0RzU0_0),.clk(gclk));
	jdff dff_B_AGQyKOT99_0(.din(w_dff_B_qwAs0RzU0_0),.dout(w_dff_B_AGQyKOT99_0),.clk(gclk));
	jdff dff_B_tc57UX8A4_0(.din(w_dff_B_AGQyKOT99_0),.dout(w_dff_B_tc57UX8A4_0),.clk(gclk));
	jdff dff_B_feVGc99K0_0(.din(w_dff_B_tc57UX8A4_0),.dout(w_dff_B_feVGc99K0_0),.clk(gclk));
	jdff dff_A_9XCsPnyq0_0(.dout(w_n680_0[0]),.din(w_dff_A_9XCsPnyq0_0),.clk(gclk));
	jdff dff_A_8eEhKBq17_0(.dout(w_dff_A_9XCsPnyq0_0),.din(w_dff_A_8eEhKBq17_0),.clk(gclk));
	jdff dff_A_5OMXwIDe1_0(.dout(w_dff_A_8eEhKBq17_0),.din(w_dff_A_5OMXwIDe1_0),.clk(gclk));
	jdff dff_A_Ti09UHVE7_0(.dout(w_dff_A_5OMXwIDe1_0),.din(w_dff_A_Ti09UHVE7_0),.clk(gclk));
	jdff dff_A_Daa9saj76_0(.dout(w_dff_A_Ti09UHVE7_0),.din(w_dff_A_Daa9saj76_0),.clk(gclk));
	jdff dff_A_8WWlmnKE4_1(.dout(w_n679_0[1]),.din(w_dff_A_8WWlmnKE4_1),.clk(gclk));
	jdff dff_A_rbPYaqof3_1(.dout(w_dff_A_8WWlmnKE4_1),.din(w_dff_A_rbPYaqof3_1),.clk(gclk));
	jdff dff_A_FRanbqnu6_2(.dout(w_n679_0[2]),.din(w_dff_A_FRanbqnu6_2),.clk(gclk));
	jdff dff_A_fvdlIUf07_0(.dout(w_n678_0[0]),.din(w_dff_A_fvdlIUf07_0),.clk(gclk));
	jdff dff_A_hE0veTSZ4_0(.dout(w_dff_A_fvdlIUf07_0),.din(w_dff_A_hE0veTSZ4_0),.clk(gclk));
	jdff dff_A_V3BLaXsn7_0(.dout(w_dff_A_hE0veTSZ4_0),.din(w_dff_A_V3BLaXsn7_0),.clk(gclk));
	jdff dff_A_rD5zJ8nL4_0(.dout(w_dff_A_V3BLaXsn7_0),.din(w_dff_A_rD5zJ8nL4_0),.clk(gclk));
	jdff dff_A_V3ymn84W6_0(.dout(w_dff_A_rD5zJ8nL4_0),.din(w_dff_A_V3ymn84W6_0),.clk(gclk));
	jdff dff_A_YT94TjR65_0(.dout(w_dff_A_V3ymn84W6_0),.din(w_dff_A_YT94TjR65_0),.clk(gclk));
	jdff dff_A_0fGialP43_0(.dout(w_dff_A_YT94TjR65_0),.din(w_dff_A_0fGialP43_0),.clk(gclk));
	jdff dff_A_PB3WXhFH4_0(.dout(w_dff_A_0fGialP43_0),.din(w_dff_A_PB3WXhFH4_0),.clk(gclk));
	jdff dff_A_TYaNBxp94_0(.dout(w_dff_A_PB3WXhFH4_0),.din(w_dff_A_TYaNBxp94_0),.clk(gclk));
	jdff dff_A_nP3cP89Q1_0(.dout(w_dff_A_TYaNBxp94_0),.din(w_dff_A_nP3cP89Q1_0),.clk(gclk));
	jdff dff_A_xda0SqpW2_0(.dout(w_dff_A_nP3cP89Q1_0),.din(w_dff_A_xda0SqpW2_0),.clk(gclk));
	jdff dff_A_tRuD1V2k2_0(.dout(w_dff_A_xda0SqpW2_0),.din(w_dff_A_tRuD1V2k2_0),.clk(gclk));
	jdff dff_A_6oNDj94a0_0(.dout(w_dff_A_tRuD1V2k2_0),.din(w_dff_A_6oNDj94a0_0),.clk(gclk));
	jdff dff_A_iA5BEcc10_0(.dout(w_dff_A_6oNDj94a0_0),.din(w_dff_A_iA5BEcc10_0),.clk(gclk));
	jdff dff_A_jdcYEks77_0(.dout(w_dff_A_iA5BEcc10_0),.din(w_dff_A_jdcYEks77_0),.clk(gclk));
	jdff dff_A_TO1bcOxd6_0(.dout(w_dff_A_jdcYEks77_0),.din(w_dff_A_TO1bcOxd6_0),.clk(gclk));
	jdff dff_A_xiihzCYQ5_1(.dout(w_n678_0[1]),.din(w_dff_A_xiihzCYQ5_1),.clk(gclk));
	jdff dff_A_AyQQ2bSt9_1(.dout(w_dff_A_xiihzCYQ5_1),.din(w_dff_A_AyQQ2bSt9_1),.clk(gclk));
	jdff dff_A_GNBlyuSq0_1(.dout(w_dff_A_AyQQ2bSt9_1),.din(w_dff_A_GNBlyuSq0_1),.clk(gclk));
	jdff dff_A_fY9xoZWJ3_1(.dout(w_dff_A_GNBlyuSq0_1),.din(w_dff_A_fY9xoZWJ3_1),.clk(gclk));
	jdff dff_A_mJBtE6ap4_1(.dout(w_dff_A_fY9xoZWJ3_1),.din(w_dff_A_mJBtE6ap4_1),.clk(gclk));
	jdff dff_A_s4WJXje08_1(.dout(w_dff_A_mJBtE6ap4_1),.din(w_dff_A_s4WJXje08_1),.clk(gclk));
	jdff dff_A_PDB5Xoln1_1(.dout(w_dff_A_s4WJXje08_1),.din(w_dff_A_PDB5Xoln1_1),.clk(gclk));
	jdff dff_A_VKbcsXEq2_1(.dout(w_dff_A_PDB5Xoln1_1),.din(w_dff_A_VKbcsXEq2_1),.clk(gclk));
	jdff dff_A_06HFvkNS3_1(.dout(w_dff_A_VKbcsXEq2_1),.din(w_dff_A_06HFvkNS3_1),.clk(gclk));
	jdff dff_A_DeDgElBp2_1(.dout(w_dff_A_06HFvkNS3_1),.din(w_dff_A_DeDgElBp2_1),.clk(gclk));
	jdff dff_A_jMCt2khf6_1(.dout(w_dff_A_DeDgElBp2_1),.din(w_dff_A_jMCt2khf6_1),.clk(gclk));
	jdff dff_A_7ZCymeVj2_1(.dout(w_dff_A_jMCt2khf6_1),.din(w_dff_A_7ZCymeVj2_1),.clk(gclk));
	jdff dff_A_aWopnpTk0_1(.dout(w_dff_A_7ZCymeVj2_1),.din(w_dff_A_aWopnpTk0_1),.clk(gclk));
	jdff dff_A_4nmzhXjS1_1(.dout(w_dff_A_aWopnpTk0_1),.din(w_dff_A_4nmzhXjS1_1),.clk(gclk));
	jdff dff_A_fPeRa39J5_1(.dout(w_dff_A_4nmzhXjS1_1),.din(w_dff_A_fPeRa39J5_1),.clk(gclk));
	jdff dff_A_KLSNYSLk1_1(.dout(w_dff_A_fPeRa39J5_1),.din(w_dff_A_KLSNYSLk1_1),.clk(gclk));
	jdff dff_B_udsJNlPp0_0(.din(G209),.dout(w_dff_B_udsJNlPp0_0),.clk(gclk));
	jdff dff_B_WK6fjMJF0_3(.din(n675),.dout(w_dff_B_WK6fjMJF0_3),.clk(gclk));
	jdff dff_B_GUFRaQMM5_3(.din(w_dff_B_WK6fjMJF0_3),.dout(w_dff_B_GUFRaQMM5_3),.clk(gclk));
	jdff dff_A_JGRcI2k97_0(.dout(w_n674_1[0]),.din(w_dff_A_JGRcI2k97_0),.clk(gclk));
	jdff dff_A_bgfH7TTV2_0(.dout(w_dff_A_JGRcI2k97_0),.din(w_dff_A_bgfH7TTV2_0),.clk(gclk));
	jdff dff_A_OTuDoVcH2_0(.dout(w_dff_A_bgfH7TTV2_0),.din(w_dff_A_OTuDoVcH2_0),.clk(gclk));
	jdff dff_A_Iv7RmCSa2_0(.dout(w_dff_A_OTuDoVcH2_0),.din(w_dff_A_Iv7RmCSa2_0),.clk(gclk));
	jdff dff_A_rHVxTPQG0_0(.dout(w_dff_A_Iv7RmCSa2_0),.din(w_dff_A_rHVxTPQG0_0),.clk(gclk));
	jdff dff_A_3RqUMvrE7_0(.dout(w_dff_A_rHVxTPQG0_0),.din(w_dff_A_3RqUMvrE7_0),.clk(gclk));
	jdff dff_A_vJEghP9R5_0(.dout(w_dff_A_3RqUMvrE7_0),.din(w_dff_A_vJEghP9R5_0),.clk(gclk));
	jdff dff_A_lTbCO6GF2_0(.dout(w_dff_A_vJEghP9R5_0),.din(w_dff_A_lTbCO6GF2_0),.clk(gclk));
	jdff dff_A_aCjbTltz9_0(.dout(w_dff_A_lTbCO6GF2_0),.din(w_dff_A_aCjbTltz9_0),.clk(gclk));
	jdff dff_A_LE96f8vS1_0(.dout(w_dff_A_aCjbTltz9_0),.din(w_dff_A_LE96f8vS1_0),.clk(gclk));
	jdff dff_A_ZODp8GNB0_0(.dout(w_dff_A_LE96f8vS1_0),.din(w_dff_A_ZODp8GNB0_0),.clk(gclk));
	jdff dff_A_3c6MWIrS9_0(.dout(w_dff_A_ZODp8GNB0_0),.din(w_dff_A_3c6MWIrS9_0),.clk(gclk));
	jdff dff_A_ZUv04b8S4_0(.dout(w_dff_A_3c6MWIrS9_0),.din(w_dff_A_ZUv04b8S4_0),.clk(gclk));
	jdff dff_A_prV4Fc1H6_0(.dout(w_dff_A_ZUv04b8S4_0),.din(w_dff_A_prV4Fc1H6_0),.clk(gclk));
	jdff dff_A_cFtqU0P68_0(.dout(w_dff_A_prV4Fc1H6_0),.din(w_dff_A_cFtqU0P68_0),.clk(gclk));
	jdff dff_A_yJEJunf87_0(.dout(w_dff_A_cFtqU0P68_0),.din(w_dff_A_yJEJunf87_0),.clk(gclk));
	jdff dff_A_HNKgZz319_0(.dout(w_dff_A_yJEJunf87_0),.din(w_dff_A_HNKgZz319_0),.clk(gclk));
	jdff dff_A_DsUS2yNh5_0(.dout(w_dff_A_HNKgZz319_0),.din(w_dff_A_DsUS2yNh5_0),.clk(gclk));
	jdff dff_A_xDywGDeL8_1(.dout(w_n674_0[1]),.din(w_dff_A_xDywGDeL8_1),.clk(gclk));
	jdff dff_A_gdaA7rRV3_1(.dout(w_dff_A_xDywGDeL8_1),.din(w_dff_A_gdaA7rRV3_1),.clk(gclk));
	jdff dff_A_TScRDQKd7_1(.dout(w_dff_A_gdaA7rRV3_1),.din(w_dff_A_TScRDQKd7_1),.clk(gclk));
	jdff dff_A_T5GcRxaG5_1(.dout(w_dff_A_TScRDQKd7_1),.din(w_dff_A_T5GcRxaG5_1),.clk(gclk));
	jdff dff_A_2sHnn7nZ5_1(.dout(w_dff_A_T5GcRxaG5_1),.din(w_dff_A_2sHnn7nZ5_1),.clk(gclk));
	jdff dff_A_vrYJmitD3_1(.dout(w_dff_A_2sHnn7nZ5_1),.din(w_dff_A_vrYJmitD3_1),.clk(gclk));
	jdff dff_A_iNDNhe8h1_1(.dout(w_dff_A_vrYJmitD3_1),.din(w_dff_A_iNDNhe8h1_1),.clk(gclk));
	jdff dff_A_CM21eqFK8_1(.dout(w_dff_A_iNDNhe8h1_1),.din(w_dff_A_CM21eqFK8_1),.clk(gclk));
	jdff dff_A_fZ7jKNA22_1(.dout(w_dff_A_CM21eqFK8_1),.din(w_dff_A_fZ7jKNA22_1),.clk(gclk));
	jdff dff_A_3OXEH8oE9_1(.dout(w_dff_A_fZ7jKNA22_1),.din(w_dff_A_3OXEH8oE9_1),.clk(gclk));
	jdff dff_A_tTZJIxOV3_1(.dout(w_dff_A_3OXEH8oE9_1),.din(w_dff_A_tTZJIxOV3_1),.clk(gclk));
	jdff dff_A_orLETswG8_1(.dout(w_dff_A_tTZJIxOV3_1),.din(w_dff_A_orLETswG8_1),.clk(gclk));
	jdff dff_A_USr6oUuH6_1(.dout(w_dff_A_orLETswG8_1),.din(w_dff_A_USr6oUuH6_1),.clk(gclk));
	jdff dff_A_jSWqxQtg4_0(.dout(w_n672_0[0]),.din(w_dff_A_jSWqxQtg4_0),.clk(gclk));
	jdff dff_A_h8xI2N846_0(.dout(w_dff_A_jSWqxQtg4_0),.din(w_dff_A_h8xI2N846_0),.clk(gclk));
	jdff dff_B_weg95XQN7_0(.din(G216),.dout(w_dff_B_weg95XQN7_0),.clk(gclk));
	jdff dff_B_pV88N8Af2_2(.din(n671),.dout(w_dff_B_pV88N8Af2_2),.clk(gclk));
	jdff dff_B_Eyc3M63f7_2(.din(w_dff_B_pV88N8Af2_2),.dout(w_dff_B_Eyc3M63f7_2),.clk(gclk));
	jdff dff_A_l5zi4vCn3_0(.dout(w_G1469_1[0]),.din(w_dff_A_l5zi4vCn3_0),.clk(gclk));
	jdff dff_A_QgTKHKAo5_0(.dout(w_dff_A_l5zi4vCn3_0),.din(w_dff_A_QgTKHKAo5_0),.clk(gclk));
	jdff dff_A_fruoJbux2_0(.dout(w_dff_A_QgTKHKAo5_0),.din(w_dff_A_fruoJbux2_0),.clk(gclk));
	jdff dff_A_LscgSKAo6_0(.dout(w_dff_A_fruoJbux2_0),.din(w_dff_A_LscgSKAo6_0),.clk(gclk));
	jdff dff_A_iaF6eQku4_0(.dout(w_n667_0[0]),.din(w_dff_A_iaF6eQku4_0),.clk(gclk));
	jdff dff_A_geoSaktb6_0(.dout(w_dff_A_iaF6eQku4_0),.din(w_dff_A_geoSaktb6_0),.clk(gclk));
	jdff dff_B_e0zlQvZn0_0(.din(G215),.dout(w_dff_B_e0zlQvZn0_0),.clk(gclk));
	jdff dff_B_jgMXV8T65_2(.din(n666),.dout(w_dff_B_jgMXV8T65_2),.clk(gclk));
	jdff dff_B_wObdoSbL6_2(.din(w_dff_B_jgMXV8T65_2),.dout(w_dff_B_wObdoSbL6_2),.clk(gclk));
	jdff dff_A_XntA4lmx0_0(.dout(w_G106_1[0]),.din(w_dff_A_XntA4lmx0_0),.clk(gclk));
	jdff dff_A_KMuYR9Ki9_0(.dout(w_dff_A_XntA4lmx0_0),.din(w_dff_A_KMuYR9Ki9_0),.clk(gclk));
	jdff dff_A_MkTrKxAc3_0(.dout(w_dff_A_KMuYR9Ki9_0),.din(w_dff_A_MkTrKxAc3_0),.clk(gclk));
	jdff dff_A_OEopb4TV0_0(.dout(w_dff_A_MkTrKxAc3_0),.din(w_dff_A_OEopb4TV0_0),.clk(gclk));
	jdff dff_B_5Zv08cyB5_0(.din(G214),.dout(w_dff_B_5Zv08cyB5_0),.clk(gclk));
	jdff dff_B_nVVeEWNQ7_3(.din(n662),.dout(w_dff_B_nVVeEWNQ7_3),.clk(gclk));
	jdff dff_B_85BJkmhI0_3(.din(w_dff_B_nVVeEWNQ7_3),.dout(w_dff_B_85BJkmhI0_3),.clk(gclk));
	jdff dff_A_IJW7lCWL1_1(.dout(w_n661_0[1]),.din(w_dff_A_IJW7lCWL1_1),.clk(gclk));
	jdff dff_A_jxNuVVNz2_1(.dout(w_dff_A_IJW7lCWL1_1),.din(w_dff_A_jxNuVVNz2_1),.clk(gclk));
	jdff dff_B_Fp6gxk5S3_0(.din(G213),.dout(w_dff_B_Fp6gxk5S3_0),.clk(gclk));
	jdff dff_B_jHmAqFaa1_3(.din(n658),.dout(w_dff_B_jHmAqFaa1_3),.clk(gclk));
	jdff dff_B_FnI5fl3B8_3(.din(w_dff_B_jHmAqFaa1_3),.dout(w_dff_B_FnI5fl3B8_3),.clk(gclk));
	jdff dff_A_qVeOrooV1_1(.dout(w_n656_0[1]),.din(w_dff_A_qVeOrooV1_1),.clk(gclk));
	jdff dff_A_qSpE3dCf7_1(.dout(w_dff_A_qVeOrooV1_1),.din(w_dff_A_qSpE3dCf7_1),.clk(gclk));
	jdff dff_A_LscvcbqR1_1(.dout(w_dff_A_qSpE3dCf7_1),.din(w_dff_A_LscvcbqR1_1),.clk(gclk));
	jdff dff_A_3BY8umy39_1(.dout(w_dff_A_LscvcbqR1_1),.din(w_dff_A_3BY8umy39_1),.clk(gclk));
	jdff dff_A_zCK0k53w2_1(.dout(w_dff_A_3BY8umy39_1),.din(w_dff_A_zCK0k53w2_1),.clk(gclk));
	jdff dff_A_IkbB7Ann4_1(.dout(w_dff_A_zCK0k53w2_1),.din(w_dff_A_IkbB7Ann4_1),.clk(gclk));
	jdff dff_A_X1PHcyRL8_1(.dout(w_dff_A_IkbB7Ann4_1),.din(w_dff_A_X1PHcyRL8_1),.clk(gclk));
	jdff dff_A_GCDSSDzN3_1(.dout(w_dff_A_X1PHcyRL8_1),.din(w_dff_A_GCDSSDzN3_1),.clk(gclk));
	jdff dff_A_KeIE0M3X6_1(.dout(w_dff_A_GCDSSDzN3_1),.din(w_dff_A_KeIE0M3X6_1),.clk(gclk));
	jdff dff_B_YgOYIF3J7_1(.din(n641),.dout(w_dff_B_YgOYIF3J7_1),.clk(gclk));
	jdff dff_B_69j5AqhJ2_1(.din(w_dff_B_YgOYIF3J7_1),.dout(w_dff_B_69j5AqhJ2_1),.clk(gclk));
	jdff dff_B_03msNVtN4_1(.din(w_dff_B_69j5AqhJ2_1),.dout(w_dff_B_03msNVtN4_1),.clk(gclk));
	jdff dff_B_tDOpbQM73_1(.din(w_dff_B_03msNVtN4_1),.dout(w_dff_B_tDOpbQM73_1),.clk(gclk));
	jdff dff_B_435MBe004_0(.din(n654),.dout(w_dff_B_435MBe004_0),.clk(gclk));
	jdff dff_B_ckRGBXmw0_0(.din(w_dff_B_435MBe004_0),.dout(w_dff_B_ckRGBXmw0_0),.clk(gclk));
	jdff dff_A_bNteBb4o9_0(.dout(w_n653_1[0]),.din(w_dff_A_bNteBb4o9_0),.clk(gclk));
	jdff dff_A_eaJWVmC34_0(.dout(w_dff_A_bNteBb4o9_0),.din(w_dff_A_eaJWVmC34_0),.clk(gclk));
	jdff dff_A_b6OPPDXl6_0(.dout(w_dff_A_eaJWVmC34_0),.din(w_dff_A_b6OPPDXl6_0),.clk(gclk));
	jdff dff_A_q6D6LlFW4_0(.dout(w_dff_A_b6OPPDXl6_0),.din(w_dff_A_q6D6LlFW4_0),.clk(gclk));
	jdff dff_A_awmwhBX11_0(.dout(w_dff_A_q6D6LlFW4_0),.din(w_dff_A_awmwhBX11_0),.clk(gclk));
	jdff dff_A_EvfdTHg96_0(.dout(w_dff_A_awmwhBX11_0),.din(w_dff_A_EvfdTHg96_0),.clk(gclk));
	jdff dff_A_tH90sqyA2_0(.dout(w_dff_A_EvfdTHg96_0),.din(w_dff_A_tH90sqyA2_0),.clk(gclk));
	jdff dff_A_z7d9PcIj6_0(.dout(w_dff_A_tH90sqyA2_0),.din(w_dff_A_z7d9PcIj6_0),.clk(gclk));
	jdff dff_A_OS3DCQfI6_0(.dout(w_dff_A_z7d9PcIj6_0),.din(w_dff_A_OS3DCQfI6_0),.clk(gclk));
	jdff dff_A_PdjvSOFp3_0(.dout(w_dff_A_OS3DCQfI6_0),.din(w_dff_A_PdjvSOFp3_0),.clk(gclk));
	jdff dff_A_00GPrgor6_0(.dout(w_dff_A_PdjvSOFp3_0),.din(w_dff_A_00GPrgor6_0),.clk(gclk));
	jdff dff_A_luDb0KQi7_0(.dout(w_dff_A_00GPrgor6_0),.din(w_dff_A_luDb0KQi7_0),.clk(gclk));
	jdff dff_A_nOz2c55t1_0(.dout(w_dff_A_luDb0KQi7_0),.din(w_dff_A_nOz2c55t1_0),.clk(gclk));
	jdff dff_A_Mx6Eqkxj6_0(.dout(w_dff_A_nOz2c55t1_0),.din(w_dff_A_Mx6Eqkxj6_0),.clk(gclk));
	jdff dff_A_b79Vmeps7_0(.dout(w_dff_A_Mx6Eqkxj6_0),.din(w_dff_A_b79Vmeps7_0),.clk(gclk));
	jdff dff_A_lhQwHW589_1(.dout(w_n653_0[1]),.din(w_dff_A_lhQwHW589_1),.clk(gclk));
	jdff dff_A_DJPvStd51_1(.dout(w_dff_A_lhQwHW589_1),.din(w_dff_A_DJPvStd51_1),.clk(gclk));
	jdff dff_A_KJrEFhzp3_1(.dout(w_dff_A_DJPvStd51_1),.din(w_dff_A_KJrEFhzp3_1),.clk(gclk));
	jdff dff_A_ugyXVVpA3_1(.dout(w_n648_0[1]),.din(w_dff_A_ugyXVVpA3_1),.clk(gclk));
	jdff dff_A_CkolcgPb0_1(.dout(w_dff_A_ugyXVVpA3_1),.din(w_dff_A_CkolcgPb0_1),.clk(gclk));
	jdff dff_A_SlJU4UrV7_1(.dout(w_dff_A_CkolcgPb0_1),.din(w_dff_A_SlJU4UrV7_1),.clk(gclk));
	jdff dff_A_uQx4ckUS8_1(.dout(w_dff_A_SlJU4UrV7_1),.din(w_dff_A_uQx4ckUS8_1),.clk(gclk));
	jdff dff_A_TzXperJG2_1(.dout(w_dff_A_uQx4ckUS8_1),.din(w_dff_A_TzXperJG2_1),.clk(gclk));
	jdff dff_A_zM1eOZtC8_1(.dout(w_dff_A_TzXperJG2_1),.din(w_dff_A_zM1eOZtC8_1),.clk(gclk));
	jdff dff_A_vugQn8406_1(.dout(w_dff_A_zM1eOZtC8_1),.din(w_dff_A_vugQn8406_1),.clk(gclk));
	jdff dff_A_AUAQRt9i6_1(.dout(w_dff_A_vugQn8406_1),.din(w_dff_A_AUAQRt9i6_1),.clk(gclk));
	jdff dff_A_YzinDvIG0_1(.dout(w_dff_A_AUAQRt9i6_1),.din(w_dff_A_YzinDvIG0_1),.clk(gclk));
	jdff dff_A_GDRDDe720_1(.dout(w_dff_A_YzinDvIG0_1),.din(w_dff_A_GDRDDe720_1),.clk(gclk));
	jdff dff_A_5hJs1hqs3_1(.dout(w_dff_A_GDRDDe720_1),.din(w_dff_A_5hJs1hqs3_1),.clk(gclk));
	jdff dff_A_5EVaKySu6_1(.dout(w_dff_A_5hJs1hqs3_1),.din(w_dff_A_5EVaKySu6_1),.clk(gclk));
	jdff dff_B_S3vLjFV19_1(.din(n644),.dout(w_dff_B_S3vLjFV19_1),.clk(gclk));
	jdff dff_A_uEeCJ1Kd7_0(.dout(w_n645_0[0]),.din(w_dff_A_uEeCJ1Kd7_0),.clk(gclk));
	jdff dff_A_QHpEqIbG6_1(.dout(w_n645_0[1]),.din(w_dff_A_QHpEqIbG6_1),.clk(gclk));
	jdff dff_A_ZFBqdPzH8_1(.dout(w_dff_A_QHpEqIbG6_1),.din(w_dff_A_ZFBqdPzH8_1),.clk(gclk));
	jdff dff_A_YECXhcwt4_1(.dout(w_dff_A_ZFBqdPzH8_1),.din(w_dff_A_YECXhcwt4_1),.clk(gclk));
	jdff dff_A_6qsqugpf0_1(.dout(w_dff_A_YECXhcwt4_1),.din(w_dff_A_6qsqugpf0_1),.clk(gclk));
	jdff dff_A_yzBiQcqj7_1(.dout(w_dff_A_6qsqugpf0_1),.din(w_dff_A_yzBiQcqj7_1),.clk(gclk));
	jdff dff_A_6zVeFx6p9_1(.dout(w_dff_A_yzBiQcqj7_1),.din(w_dff_A_6zVeFx6p9_1),.clk(gclk));
	jdff dff_A_4hJKT1sK1_1(.dout(w_dff_A_6zVeFx6p9_1),.din(w_dff_A_4hJKT1sK1_1),.clk(gclk));
	jdff dff_A_XH7GOK6u1_1(.dout(w_dff_A_4hJKT1sK1_1),.din(w_dff_A_XH7GOK6u1_1),.clk(gclk));
	jdff dff_A_TAgsMGfK2_1(.dout(w_dff_A_XH7GOK6u1_1),.din(w_dff_A_TAgsMGfK2_1),.clk(gclk));
	jdff dff_A_FNk3zqNX8_1(.dout(w_dff_A_TAgsMGfK2_1),.din(w_dff_A_FNk3zqNX8_1),.clk(gclk));
	jdff dff_A_xbUZFV986_1(.dout(w_dff_A_FNk3zqNX8_1),.din(w_dff_A_xbUZFV986_1),.clk(gclk));
	jdff dff_A_21BPTPe51_1(.dout(w_dff_A_xbUZFV986_1),.din(w_dff_A_21BPTPe51_1),.clk(gclk));
	jdff dff_A_ANqimZD49_1(.dout(w_dff_A_21BPTPe51_1),.din(w_dff_A_ANqimZD49_1),.clk(gclk));
	jdff dff_A_2b5r9XDY0_1(.dout(w_dff_A_ANqimZD49_1),.din(w_dff_A_2b5r9XDY0_1),.clk(gclk));
	jdff dff_A_vbxwZFMd3_1(.dout(w_dff_A_2b5r9XDY0_1),.din(w_dff_A_vbxwZFMd3_1),.clk(gclk));
	jdff dff_A_vkydJDqY9_0(.dout(w_n643_0[0]),.din(w_dff_A_vkydJDqY9_0),.clk(gclk));
	jdff dff_A_4MCI9L6I6_0(.dout(w_dff_A_vkydJDqY9_0),.din(w_dff_A_4MCI9L6I6_0),.clk(gclk));
	jdff dff_A_j5XxWvrR8_0(.dout(w_dff_A_4MCI9L6I6_0),.din(w_dff_A_j5XxWvrR8_0),.clk(gclk));
	jdff dff_A_fbr8mnGz1_0(.dout(w_dff_A_j5XxWvrR8_0),.din(w_dff_A_fbr8mnGz1_0),.clk(gclk));
	jdff dff_A_Uec39Vxm9_0(.dout(w_dff_A_fbr8mnGz1_0),.din(w_dff_A_Uec39Vxm9_0),.clk(gclk));
	jdff dff_A_XpT8h68v5_0(.dout(w_dff_A_Uec39Vxm9_0),.din(w_dff_A_XpT8h68v5_0),.clk(gclk));
	jdff dff_A_JT7c7LVJ0_0(.dout(w_dff_A_XpT8h68v5_0),.din(w_dff_A_JT7c7LVJ0_0),.clk(gclk));
	jdff dff_A_RtbzAyDX5_0(.dout(w_dff_A_JT7c7LVJ0_0),.din(w_dff_A_RtbzAyDX5_0),.clk(gclk));
	jdff dff_A_SSwrhQ8X7_0(.dout(w_dff_A_RtbzAyDX5_0),.din(w_dff_A_SSwrhQ8X7_0),.clk(gclk));
	jdff dff_A_cDmOmi2l9_0(.dout(w_dff_A_SSwrhQ8X7_0),.din(w_dff_A_cDmOmi2l9_0),.clk(gclk));
	jdff dff_A_SGFZ6jdn9_0(.dout(w_dff_A_cDmOmi2l9_0),.din(w_dff_A_SGFZ6jdn9_0),.clk(gclk));
	jdff dff_A_jBuDZjtb2_0(.dout(w_dff_A_SGFZ6jdn9_0),.din(w_dff_A_jBuDZjtb2_0),.clk(gclk));
	jdff dff_A_MDhyBYyy5_0(.dout(w_dff_A_jBuDZjtb2_0),.din(w_dff_A_MDhyBYyy5_0),.clk(gclk));
	jdff dff_A_Ai9LT4dN0_0(.dout(w_dff_A_MDhyBYyy5_0),.din(w_dff_A_Ai9LT4dN0_0),.clk(gclk));
	jdff dff_B_o1O7qU5H6_2(.din(n643),.dout(w_dff_B_o1O7qU5H6_2),.clk(gclk));
	jdff dff_B_IqbrtGa19_2(.din(w_dff_B_o1O7qU5H6_2),.dout(w_dff_B_IqbrtGa19_2),.clk(gclk));
	jdff dff_A_pQkm35fj1_0(.dout(w_n642_0[0]),.din(w_dff_A_pQkm35fj1_0),.clk(gclk));
	jdff dff_A_FMkZpi7v5_0(.dout(w_dff_A_pQkm35fj1_0),.din(w_dff_A_FMkZpi7v5_0),.clk(gclk));
	jdff dff_A_cG90Depa6_0(.dout(w_dff_A_FMkZpi7v5_0),.din(w_dff_A_cG90Depa6_0),.clk(gclk));
	jdff dff_A_unpagc5b3_0(.dout(w_dff_A_cG90Depa6_0),.din(w_dff_A_unpagc5b3_0),.clk(gclk));
	jdff dff_A_5Zp1Rz6K0_0(.dout(w_dff_A_unpagc5b3_0),.din(w_dff_A_5Zp1Rz6K0_0),.clk(gclk));
	jdff dff_B_KqLYUZDQ6_0(.din(n638),.dout(w_dff_B_KqLYUZDQ6_0),.clk(gclk));
	jdff dff_B_e7htl35A0_0(.din(w_dff_B_KqLYUZDQ6_0),.dout(w_dff_B_e7htl35A0_0),.clk(gclk));
	jdff dff_B_F2BKuxDP9_0(.din(w_dff_B_e7htl35A0_0),.dout(w_dff_B_F2BKuxDP9_0),.clk(gclk));
	jdff dff_B_6j8hxfvM7_0(.din(w_dff_B_F2BKuxDP9_0),.dout(w_dff_B_6j8hxfvM7_0),.clk(gclk));
	jdff dff_B_MsCHrmr83_0(.din(w_dff_B_6j8hxfvM7_0),.dout(w_dff_B_MsCHrmr83_0),.clk(gclk));
	jdff dff_B_X4PMTLHp7_0(.din(w_dff_B_MsCHrmr83_0),.dout(w_dff_B_X4PMTLHp7_0),.clk(gclk));
	jdff dff_B_DOzSByfZ5_0(.din(w_dff_B_X4PMTLHp7_0),.dout(w_dff_B_DOzSByfZ5_0),.clk(gclk));
	jdff dff_B_sMzYAUte7_0(.din(w_dff_B_DOzSByfZ5_0),.dout(w_dff_B_sMzYAUte7_0),.clk(gclk));
	jdff dff_B_QJV3MsJg7_0(.din(w_dff_B_sMzYAUte7_0),.dout(w_dff_B_QJV3MsJg7_0),.clk(gclk));
	jdff dff_B_65m4t7KB8_0(.din(w_dff_B_QJV3MsJg7_0),.dout(w_dff_B_65m4t7KB8_0),.clk(gclk));
	jdff dff_B_091w0Pok9_0(.din(w_dff_B_65m4t7KB8_0),.dout(w_dff_B_091w0Pok9_0),.clk(gclk));
	jdff dff_A_ybfPvBur3_0(.dout(w_n637_0[0]),.din(w_dff_A_ybfPvBur3_0),.clk(gclk));
	jdff dff_A_pI7MVA4b9_0(.dout(w_dff_A_ybfPvBur3_0),.din(w_dff_A_pI7MVA4b9_0),.clk(gclk));
	jdff dff_A_8EHDGjs86_0(.dout(w_dff_A_pI7MVA4b9_0),.din(w_dff_A_8EHDGjs86_0),.clk(gclk));
	jdff dff_A_dWI06zRd7_0(.dout(w_dff_A_8EHDGjs86_0),.din(w_dff_A_dWI06zRd7_0),.clk(gclk));
	jdff dff_A_8MIFdefm4_0(.dout(w_dff_A_dWI06zRd7_0),.din(w_dff_A_8MIFdefm4_0),.clk(gclk));
	jdff dff_A_8d4m0tp26_0(.dout(w_dff_A_8MIFdefm4_0),.din(w_dff_A_8d4m0tp26_0),.clk(gclk));
	jdff dff_A_zFQxOV633_0(.dout(w_dff_A_8d4m0tp26_0),.din(w_dff_A_zFQxOV633_0),.clk(gclk));
	jdff dff_A_Vjj4665X5_0(.dout(w_dff_A_zFQxOV633_0),.din(w_dff_A_Vjj4665X5_0),.clk(gclk));
	jdff dff_A_6IeYrVai6_0(.dout(w_dff_A_Vjj4665X5_0),.din(w_dff_A_6IeYrVai6_0),.clk(gclk));
	jdff dff_A_AMtld9Wl3_0(.dout(w_dff_A_6IeYrVai6_0),.din(w_dff_A_AMtld9Wl3_0),.clk(gclk));
	jdff dff_A_vDntd9NQ4_0(.dout(w_dff_A_AMtld9Wl3_0),.din(w_dff_A_vDntd9NQ4_0),.clk(gclk));
	jdff dff_A_RgGa0dKo8_0(.dout(w_dff_A_vDntd9NQ4_0),.din(w_dff_A_RgGa0dKo8_0),.clk(gclk));
	jdff dff_A_97LXNt6R5_0(.dout(w_n635_0[0]),.din(w_dff_A_97LXNt6R5_0),.clk(gclk));
	jdff dff_A_Ak9pEssV8_0(.dout(w_n633_0[0]),.din(w_dff_A_Ak9pEssV8_0),.clk(gclk));
	jdff dff_A_4kuSY1976_0(.dout(w_dff_A_Ak9pEssV8_0),.din(w_dff_A_4kuSY1976_0),.clk(gclk));
	jdff dff_B_IaCFlZPL7_0(.din(G154),.dout(w_dff_B_IaCFlZPL7_0),.clk(gclk));
	jdff dff_B_ecKi21p28_2(.din(n632),.dout(w_dff_B_ecKi21p28_2),.clk(gclk));
	jdff dff_B_KBlbIcD88_2(.din(w_dff_B_ecKi21p28_2),.dout(w_dff_B_KBlbIcD88_2),.clk(gclk));
	jdff dff_A_LhxZ9yvu1_0(.dout(w_G2253_1[0]),.din(w_dff_A_LhxZ9yvu1_0),.clk(gclk));
	jdff dff_A_3ecQssV03_0(.dout(w_dff_A_LhxZ9yvu1_0),.din(w_dff_A_3ecQssV03_0),.clk(gclk));
	jdff dff_A_B9TyBP2u3_0(.dout(w_dff_A_3ecQssV03_0),.din(w_dff_A_B9TyBP2u3_0),.clk(gclk));
	jdff dff_A_u1mi4Nci9_0(.dout(w_dff_A_B9TyBP2u3_0),.din(w_dff_A_u1mi4Nci9_0),.clk(gclk));
	jdff dff_A_ChkCkPCG1_0(.dout(w_n629_0[0]),.din(w_dff_A_ChkCkPCG1_0),.clk(gclk));
	jdff dff_A_a1W6TsAm6_0(.dout(w_dff_A_ChkCkPCG1_0),.din(w_dff_A_a1W6TsAm6_0),.clk(gclk));
	jdff dff_B_kkY0ITpc8_0(.din(G153),.dout(w_dff_B_kkY0ITpc8_0),.clk(gclk));
	jdff dff_B_DIXkC6457_2(.din(n628),.dout(w_dff_B_DIXkC6457_2),.clk(gclk));
	jdff dff_B_rDypx3QF1_2(.din(w_dff_B_DIXkC6457_2),.dout(w_dff_B_rDypx3QF1_2),.clk(gclk));
	jdff dff_A_jsDu7JGM6_0(.dout(w_G2256_1[0]),.din(w_dff_A_jsDu7JGM6_0),.clk(gclk));
	jdff dff_A_EQpDDZVm1_0(.dout(w_dff_A_jsDu7JGM6_0),.din(w_dff_A_EQpDDZVm1_0),.clk(gclk));
	jdff dff_A_uCDmfV8Y8_0(.dout(w_dff_A_EQpDDZVm1_0),.din(w_dff_A_uCDmfV8Y8_0),.clk(gclk));
	jdff dff_A_TzYAG5a67_0(.dout(w_dff_A_uCDmfV8Y8_0),.din(w_dff_A_TzYAG5a67_0),.clk(gclk));
	jdff dff_A_QWnGeewX5_0(.dout(w_n626_0[0]),.din(w_dff_A_QWnGeewX5_0),.clk(gclk));
	jdff dff_A_dL7AEjMH8_0(.dout(w_dff_A_QWnGeewX5_0),.din(w_dff_A_dL7AEjMH8_0),.clk(gclk));
	jdff dff_A_uiXOHSwA0_0(.dout(w_dff_A_dL7AEjMH8_0),.din(w_dff_A_uiXOHSwA0_0),.clk(gclk));
	jdff dff_A_OHXkGUO91_0(.dout(w_dff_A_uiXOHSwA0_0),.din(w_dff_A_OHXkGUO91_0),.clk(gclk));
	jdff dff_A_yxnOPSmp4_0(.dout(w_dff_A_OHXkGUO91_0),.din(w_dff_A_yxnOPSmp4_0),.clk(gclk));
	jdff dff_A_7DKIzzbP0_0(.dout(w_dff_A_yxnOPSmp4_0),.din(w_dff_A_7DKIzzbP0_0),.clk(gclk));
	jdff dff_A_84v2MvXe0_0(.dout(w_dff_A_7DKIzzbP0_0),.din(w_dff_A_84v2MvXe0_0),.clk(gclk));
	jdff dff_A_l3ve8aSz6_0(.dout(w_dff_A_84v2MvXe0_0),.din(w_dff_A_l3ve8aSz6_0),.clk(gclk));
	jdff dff_A_vE46GMCE9_0(.dout(w_dff_A_l3ve8aSz6_0),.din(w_dff_A_vE46GMCE9_0),.clk(gclk));
	jdff dff_A_Zmjj8Jnz9_0(.dout(w_dff_A_vE46GMCE9_0),.din(w_dff_A_Zmjj8Jnz9_0),.clk(gclk));
	jdff dff_A_v2SSRHR16_0(.dout(w_dff_A_Zmjj8Jnz9_0),.din(w_dff_A_v2SSRHR16_0),.clk(gclk));
	jdff dff_A_u5ULDn1n2_0(.dout(w_dff_A_v2SSRHR16_0),.din(w_dff_A_u5ULDn1n2_0),.clk(gclk));
	jdff dff_A_wa18ZgDf7_0(.dout(w_dff_A_u5ULDn1n2_0),.din(w_dff_A_wa18ZgDf7_0),.clk(gclk));
	jdff dff_A_bwotvWOV0_0(.dout(w_dff_A_wa18ZgDf7_0),.din(w_dff_A_bwotvWOV0_0),.clk(gclk));
	jdff dff_A_plzIH1ja0_0(.dout(w_n624_0[0]),.din(w_dff_A_plzIH1ja0_0),.clk(gclk));
	jdff dff_A_7oRzPrHY1_0(.dout(w_dff_A_plzIH1ja0_0),.din(w_dff_A_7oRzPrHY1_0),.clk(gclk));
	jdff dff_B_tR2tjaxm1_0(.din(G156),.dout(w_dff_B_tR2tjaxm1_0),.clk(gclk));
	jdff dff_A_lbBsmh1h3_1(.dout(w_n623_0[1]),.din(w_dff_A_lbBsmh1h3_1),.clk(gclk));
	jdff dff_A_SQQVOfIU1_1(.dout(w_dff_A_lbBsmh1h3_1),.din(w_dff_A_SQQVOfIU1_1),.clk(gclk));
	jdff dff_A_EDIaxeYi4_2(.dout(w_n623_0[2]),.din(w_dff_A_EDIaxeYi4_2),.clk(gclk));
	jdff dff_A_339cPwC63_2(.dout(w_dff_A_EDIaxeYi4_2),.din(w_dff_A_339cPwC63_2),.clk(gclk));
	jdff dff_A_xedMLPzf4_1(.dout(w_G2239_0[1]),.din(w_dff_A_xedMLPzf4_1),.clk(gclk));
	jdff dff_A_445cJRKc6_1(.dout(w_dff_A_xedMLPzf4_1),.din(w_dff_A_445cJRKc6_1),.clk(gclk));
	jdff dff_A_RmpajueA3_1(.dout(w_dff_A_445cJRKc6_1),.din(w_dff_A_RmpajueA3_1),.clk(gclk));
	jdff dff_A_utSlhqib3_1(.dout(w_dff_A_RmpajueA3_1),.din(w_dff_A_utSlhqib3_1),.clk(gclk));
	jdff dff_A_O9JauSfY0_2(.dout(w_n622_0[2]),.din(w_dff_A_O9JauSfY0_2),.clk(gclk));
	jdff dff_A_wsX0YNC02_2(.dout(w_dff_A_O9JauSfY0_2),.din(w_dff_A_wsX0YNC02_2),.clk(gclk));
	jdff dff_A_r4P6cOGv4_2(.dout(w_dff_A_wsX0YNC02_2),.din(w_dff_A_r4P6cOGv4_2),.clk(gclk));
	jdff dff_A_EQH8NnY96_2(.dout(w_dff_A_r4P6cOGv4_2),.din(w_dff_A_EQH8NnY96_2),.clk(gclk));
	jdff dff_A_yVK7dEXE8_2(.dout(w_dff_A_EQH8NnY96_2),.din(w_dff_A_yVK7dEXE8_2),.clk(gclk));
	jdff dff_A_BPCBrWS85_2(.dout(w_dff_A_yVK7dEXE8_2),.din(w_dff_A_BPCBrWS85_2),.clk(gclk));
	jdff dff_A_XSDoLaRM3_2(.dout(w_dff_A_BPCBrWS85_2),.din(w_dff_A_XSDoLaRM3_2),.clk(gclk));
	jdff dff_A_MPcsl6oq8_2(.dout(w_dff_A_XSDoLaRM3_2),.din(w_dff_A_MPcsl6oq8_2),.clk(gclk));
	jdff dff_A_SO4bQKQp2_2(.dout(w_dff_A_MPcsl6oq8_2),.din(w_dff_A_SO4bQKQp2_2),.clk(gclk));
	jdff dff_A_Dk6p4Npt7_2(.dout(w_dff_A_SO4bQKQp2_2),.din(w_dff_A_Dk6p4Npt7_2),.clk(gclk));
	jdff dff_A_7d0795xP8_2(.dout(w_dff_A_Dk6p4Npt7_2),.din(w_dff_A_7d0795xP8_2),.clk(gclk));
	jdff dff_A_EIJwjZK89_2(.dout(w_dff_A_7d0795xP8_2),.din(w_dff_A_EIJwjZK89_2),.clk(gclk));
	jdff dff_A_csZHfrIq6_2(.dout(w_dff_A_EIJwjZK89_2),.din(w_dff_A_csZHfrIq6_2),.clk(gclk));
	jdff dff_A_nOxzqm5H3_2(.dout(w_dff_A_csZHfrIq6_2),.din(w_dff_A_nOxzqm5H3_2),.clk(gclk));
	jdff dff_A_Qo2yRsu17_2(.dout(w_dff_A_nOxzqm5H3_2),.din(w_dff_A_Qo2yRsu17_2),.clk(gclk));
	jdff dff_A_xLohmLmE5_2(.dout(w_dff_A_Qo2yRsu17_2),.din(w_dff_A_xLohmLmE5_2),.clk(gclk));
	jdff dff_A_H0gCuUDW9_0(.dout(w_n620_0[0]),.din(w_dff_A_H0gCuUDW9_0),.clk(gclk));
	jdff dff_A_CCugBIQk7_0(.dout(w_dff_A_H0gCuUDW9_0),.din(w_dff_A_CCugBIQk7_0),.clk(gclk));
	jdff dff_B_CjTSjO7E8_0(.din(G155),.dout(w_dff_B_CjTSjO7E8_0),.clk(gclk));
	jdff dff_B_ADpLKgMs9_2(.din(n619),.dout(w_dff_B_ADpLKgMs9_2),.clk(gclk));
	jdff dff_B_dndzmJYW5_2(.din(w_dff_B_ADpLKgMs9_2),.dout(w_dff_B_dndzmJYW5_2),.clk(gclk));
	jdff dff_A_Qol9Hgyz9_1(.dout(w_n617_0[1]),.din(w_dff_A_Qol9Hgyz9_1),.clk(gclk));
	jdff dff_A_IOQKiYa81_1(.dout(w_dff_A_Qol9Hgyz9_1),.din(w_dff_A_IOQKiYa81_1),.clk(gclk));
	jdff dff_A_yPBV31yn5_1(.dout(w_dff_A_IOQKiYa81_1),.din(w_dff_A_yPBV31yn5_1),.clk(gclk));
	jdff dff_A_YfhzjrCU4_1(.dout(w_dff_A_yPBV31yn5_1),.din(w_dff_A_YfhzjrCU4_1),.clk(gclk));
	jdff dff_A_blJgktoG6_1(.dout(w_dff_A_YfhzjrCU4_1),.din(w_dff_A_blJgktoG6_1),.clk(gclk));
	jdff dff_B_0WeHEjwT6_1(.din(n596),.dout(w_dff_B_0WeHEjwT6_1),.clk(gclk));
	jdff dff_B_UaDBvB3V8_1(.din(w_dff_B_0WeHEjwT6_1),.dout(w_dff_B_UaDBvB3V8_1),.clk(gclk));
	jdff dff_B_y5nWNQdk5_1(.din(w_dff_B_UaDBvB3V8_1),.dout(w_dff_B_y5nWNQdk5_1),.clk(gclk));
	jdff dff_B_Ua8xhl6L1_1(.din(w_dff_B_y5nWNQdk5_1),.dout(w_dff_B_Ua8xhl6L1_1),.clk(gclk));
	jdff dff_B_aiMcBI5F2_1(.din(w_dff_B_Ua8xhl6L1_1),.dout(w_dff_B_aiMcBI5F2_1),.clk(gclk));
	jdff dff_B_fRSBs2f97_1(.din(w_dff_B_aiMcBI5F2_1),.dout(w_dff_B_fRSBs2f97_1),.clk(gclk));
	jdff dff_B_C4xbRZC99_1(.din(n598),.dout(w_dff_B_C4xbRZC99_1),.clk(gclk));
	jdff dff_B_UqPa0uPt4_1(.din(w_dff_B_C4xbRZC99_1),.dout(w_dff_B_UqPa0uPt4_1),.clk(gclk));
	jdff dff_B_jFUutsB47_1(.din(w_dff_B_UqPa0uPt4_1),.dout(w_dff_B_jFUutsB47_1),.clk(gclk));
	jdff dff_B_CDa1NEFu9_1(.din(w_dff_B_jFUutsB47_1),.dout(w_dff_B_CDa1NEFu9_1),.clk(gclk));
	jdff dff_B_MzJuDY4q3_1(.din(w_dff_B_CDa1NEFu9_1),.dout(w_dff_B_MzJuDY4q3_1),.clk(gclk));
	jdff dff_A_huNN60yY5_0(.dout(w_n615_1[0]),.din(w_dff_A_huNN60yY5_0),.clk(gclk));
	jdff dff_A_TpdLIMfW3_0(.dout(w_dff_A_huNN60yY5_0),.din(w_dff_A_TpdLIMfW3_0),.clk(gclk));
	jdff dff_A_UDdkHcvX9_0(.dout(w_dff_A_TpdLIMfW3_0),.din(w_dff_A_UDdkHcvX9_0),.clk(gclk));
	jdff dff_A_h5SWxiMo9_0(.dout(w_dff_A_UDdkHcvX9_0),.din(w_dff_A_h5SWxiMo9_0),.clk(gclk));
	jdff dff_A_bezJG88q0_0(.dout(w_dff_A_h5SWxiMo9_0),.din(w_dff_A_bezJG88q0_0),.clk(gclk));
	jdff dff_A_0llaWvgg7_0(.dout(w_dff_A_bezJG88q0_0),.din(w_dff_A_0llaWvgg7_0),.clk(gclk));
	jdff dff_A_8FalD9Nv6_0(.dout(w_dff_A_0llaWvgg7_0),.din(w_dff_A_8FalD9Nv6_0),.clk(gclk));
	jdff dff_A_N7kOG1OK9_0(.dout(w_dff_A_8FalD9Nv6_0),.din(w_dff_A_N7kOG1OK9_0),.clk(gclk));
	jdff dff_A_FfUoooxR6_0(.dout(w_dff_A_N7kOG1OK9_0),.din(w_dff_A_FfUoooxR6_0),.clk(gclk));
	jdff dff_B_ljb0zYS01_1(.din(n600),.dout(w_dff_B_ljb0zYS01_1),.clk(gclk));
	jdff dff_B_sKZIO4Kl7_1(.din(w_dff_B_ljb0zYS01_1),.dout(w_dff_B_sKZIO4Kl7_1),.clk(gclk));
	jdff dff_B_Xl0nzo603_1(.din(w_dff_B_sKZIO4Kl7_1),.dout(w_dff_B_Xl0nzo603_1),.clk(gclk));
	jdff dff_B_AfjZREIl4_1(.din(w_dff_B_Xl0nzo603_1),.dout(w_dff_B_AfjZREIl4_1),.clk(gclk));
	jdff dff_B_kJRIfhOg9_1(.din(n602),.dout(w_dff_B_kJRIfhOg9_1),.clk(gclk));
	jdff dff_B_fy9JpJqG4_1(.din(w_dff_B_kJRIfhOg9_1),.dout(w_dff_B_fy9JpJqG4_1),.clk(gclk));
	jdff dff_B_eIy8GjQg9_1(.din(w_dff_B_fy9JpJqG4_1),.dout(w_dff_B_eIy8GjQg9_1),.clk(gclk));
	jdff dff_A_J4NwGS2D7_1(.dout(w_n613_0[1]),.din(w_dff_A_J4NwGS2D7_1),.clk(gclk));
	jdff dff_A_FDiXDb1n2_1(.dout(w_dff_A_J4NwGS2D7_1),.din(w_dff_A_FDiXDb1n2_1),.clk(gclk));
	jdff dff_A_ZXnimiPQ6_1(.dout(w_dff_A_FDiXDb1n2_1),.din(w_dff_A_ZXnimiPQ6_1),.clk(gclk));
	jdff dff_A_40yMJiQN1_1(.dout(w_dff_A_ZXnimiPQ6_1),.din(w_dff_A_40yMJiQN1_1),.clk(gclk));
	jdff dff_A_mtHNvLUC4_1(.dout(w_dff_A_40yMJiQN1_1),.din(w_dff_A_mtHNvLUC4_1),.clk(gclk));
	jdff dff_A_Kl9881X80_1(.dout(w_dff_A_mtHNvLUC4_1),.din(w_dff_A_Kl9881X80_1),.clk(gclk));
	jdff dff_A_qjketKGe4_1(.dout(w_dff_A_Kl9881X80_1),.din(w_dff_A_qjketKGe4_1),.clk(gclk));
	jdff dff_A_J8jpYEg64_1(.dout(w_dff_A_qjketKGe4_1),.din(w_dff_A_J8jpYEg64_1),.clk(gclk));
	jdff dff_A_0hSalTxC6_1(.dout(w_dff_A_J8jpYEg64_1),.din(w_dff_A_0hSalTxC6_1),.clk(gclk));
	jdff dff_A_NpEFCCjl2_1(.dout(w_dff_A_0hSalTxC6_1),.din(w_dff_A_NpEFCCjl2_1),.clk(gclk));
	jdff dff_A_HHg4Rz2y6_0(.dout(w_n610_0[0]),.din(w_dff_A_HHg4Rz2y6_0),.clk(gclk));
	jdff dff_A_xXkZjEFp7_0(.dout(w_dff_A_HHg4Rz2y6_0),.din(w_dff_A_xXkZjEFp7_0),.clk(gclk));
	jdff dff_A_nf5lgtpQ7_0(.dout(w_n608_0[0]),.din(w_dff_A_nf5lgtpQ7_0),.clk(gclk));
	jdff dff_A_L8Ushhu59_0(.dout(w_dff_A_nf5lgtpQ7_0),.din(w_dff_A_L8Ushhu59_0),.clk(gclk));
	jdff dff_A_bZekAmin1_0(.dout(w_n606_1[0]),.din(w_dff_A_bZekAmin1_0),.clk(gclk));
	jdff dff_A_x4bIKLof6_0(.dout(w_dff_A_bZekAmin1_0),.din(w_dff_A_x4bIKLof6_0),.clk(gclk));
	jdff dff_A_dhhsFBbt7_0(.dout(w_dff_A_x4bIKLof6_0),.din(w_dff_A_dhhsFBbt7_0),.clk(gclk));
	jdff dff_A_A9i6iMN36_0(.dout(w_dff_A_dhhsFBbt7_0),.din(w_dff_A_A9i6iMN36_0),.clk(gclk));
	jdff dff_A_kaXZPYvP4_1(.dout(w_n606_1[1]),.din(w_dff_A_kaXZPYvP4_1),.clk(gclk));
	jdff dff_A_GkDG18xJ9_1(.dout(w_dff_A_kaXZPYvP4_1),.din(w_dff_A_GkDG18xJ9_1),.clk(gclk));
	jdff dff_A_SNKgBfrg9_1(.dout(w_dff_A_GkDG18xJ9_1),.din(w_dff_A_SNKgBfrg9_1),.clk(gclk));
	jdff dff_A_10WBB4Jz3_1(.dout(w_dff_A_SNKgBfrg9_1),.din(w_dff_A_10WBB4Jz3_1),.clk(gclk));
	jdff dff_A_yfMtXqFG7_1(.dout(w_dff_A_10WBB4Jz3_1),.din(w_dff_A_yfMtXqFG7_1),.clk(gclk));
	jdff dff_A_zmmBnKTY3_1(.dout(w_dff_A_yfMtXqFG7_1),.din(w_dff_A_zmmBnKTY3_1),.clk(gclk));
	jdff dff_A_hdKrECdf5_1(.dout(w_dff_A_zmmBnKTY3_1),.din(w_dff_A_hdKrECdf5_1),.clk(gclk));
	jdff dff_A_DJtqrTPq6_1(.dout(w_dff_A_hdKrECdf5_1),.din(w_dff_A_DJtqrTPq6_1),.clk(gclk));
	jdff dff_A_OC8CCdl30_1(.dout(w_dff_A_DJtqrTPq6_1),.din(w_dff_A_OC8CCdl30_1),.clk(gclk));
	jdff dff_A_Fh8TcCSe5_1(.dout(w_dff_A_OC8CCdl30_1),.din(w_dff_A_Fh8TcCSe5_1),.clk(gclk));
	jdff dff_A_218tGpni1_1(.dout(w_dff_A_Fh8TcCSe5_1),.din(w_dff_A_218tGpni1_1),.clk(gclk));
	jdff dff_A_df66RkNt7_1(.dout(w_dff_A_218tGpni1_1),.din(w_dff_A_df66RkNt7_1),.clk(gclk));
	jdff dff_A_yf1K9M6n8_1(.dout(w_dff_A_df66RkNt7_1),.din(w_dff_A_yf1K9M6n8_1),.clk(gclk));
	jdff dff_A_4jb3fm2h9_0(.dout(w_n599_0[0]),.din(w_dff_A_4jb3fm2h9_0),.clk(gclk));
	jdff dff_A_PTrey4Yo3_0(.dout(w_dff_A_4jb3fm2h9_0),.din(w_dff_A_PTrey4Yo3_0),.clk(gclk));
	jdff dff_A_GphfJqkJ9_0(.dout(w_dff_A_PTrey4Yo3_0),.din(w_dff_A_GphfJqkJ9_0),.clk(gclk));
	jdff dff_A_NdxeDYtO8_0(.dout(w_dff_A_GphfJqkJ9_0),.din(w_dff_A_NdxeDYtO8_0),.clk(gclk));
	jdff dff_A_01lbMFDm6_0(.dout(w_dff_A_NdxeDYtO8_0),.din(w_dff_A_01lbMFDm6_0),.clk(gclk));
	jdff dff_B_JUhqLK8e8_0(.din(n593),.dout(w_dff_B_JUhqLK8e8_0),.clk(gclk));
	jdff dff_B_bnaJMKkr2_0(.din(w_dff_B_JUhqLK8e8_0),.dout(w_dff_B_bnaJMKkr2_0),.clk(gclk));
	jdff dff_B_Z93NSqwa0_0(.din(w_dff_B_bnaJMKkr2_0),.dout(w_dff_B_Z93NSqwa0_0),.clk(gclk));
	jdff dff_B_ao231VoQ1_0(.din(w_dff_B_Z93NSqwa0_0),.dout(w_dff_B_ao231VoQ1_0),.clk(gclk));
	jdff dff_B_i76IiTVh7_0(.din(w_dff_B_ao231VoQ1_0),.dout(w_dff_B_i76IiTVh7_0),.clk(gclk));
	jdff dff_B_yGKU4BSb7_0(.din(w_dff_B_i76IiTVh7_0),.dout(w_dff_B_yGKU4BSb7_0),.clk(gclk));
	jdff dff_B_8bNiacfX0_0(.din(w_dff_B_yGKU4BSb7_0),.dout(w_dff_B_8bNiacfX0_0),.clk(gclk));
	jdff dff_B_DshOYC767_0(.din(w_dff_B_8bNiacfX0_0),.dout(w_dff_B_DshOYC767_0),.clk(gclk));
	jdff dff_A_JtqXeOdU1_0(.dout(w_n592_0[0]),.din(w_dff_A_JtqXeOdU1_0),.clk(gclk));
	jdff dff_A_xzq3fRFG5_0(.dout(w_dff_A_JtqXeOdU1_0),.din(w_dff_A_xzq3fRFG5_0),.clk(gclk));
	jdff dff_A_UINr5WXI7_0(.dout(w_dff_A_xzq3fRFG5_0),.din(w_dff_A_UINr5WXI7_0),.clk(gclk));
	jdff dff_A_2AiPig9S6_0(.dout(w_dff_A_UINr5WXI7_0),.din(w_dff_A_2AiPig9S6_0),.clk(gclk));
	jdff dff_A_9lSxNiku9_0(.dout(w_dff_A_2AiPig9S6_0),.din(w_dff_A_9lSxNiku9_0),.clk(gclk));
	jdff dff_A_KFPKnCKc0_0(.dout(w_dff_A_9lSxNiku9_0),.din(w_dff_A_KFPKnCKc0_0),.clk(gclk));
	jdff dff_A_91GB3Sui2_0(.dout(w_dff_A_KFPKnCKc0_0),.din(w_dff_A_91GB3Sui2_0),.clk(gclk));
	jdff dff_A_Ev4PBiJo0_0(.dout(w_dff_A_91GB3Sui2_0),.din(w_dff_A_Ev4PBiJo0_0),.clk(gclk));
	jdff dff_A_LLjFKsmq6_0(.dout(w_dff_A_Ev4PBiJo0_0),.din(w_dff_A_LLjFKsmq6_0),.clk(gclk));
	jdff dff_A_uzIPxl4Y3_1(.dout(w_n589_0[1]),.din(w_dff_A_uzIPxl4Y3_1),.clk(gclk));
	jdff dff_B_HUTl7wB53_0(.din(n587),.dout(w_dff_B_HUTl7wB53_0),.clk(gclk));
	jdff dff_B_EydYX5KM5_0(.din(G144),.dout(w_dff_B_EydYX5KM5_0),.clk(gclk));
	jdff dff_B_NsXq0WyH9_2(.din(n585),.dout(w_dff_B_NsXq0WyH9_2),.clk(gclk));
	jdff dff_B_UbAXsghV7_2(.din(w_dff_B_NsXq0WyH9_2),.dout(w_dff_B_UbAXsghV7_2),.clk(gclk));
	jdff dff_A_Us4OlCG36_0(.dout(w_G2224_1[0]),.din(w_dff_A_Us4OlCG36_0),.clk(gclk));
	jdff dff_A_6bamHLNX1_0(.dout(w_dff_A_Us4OlCG36_0),.din(w_dff_A_6bamHLNX1_0),.clk(gclk));
	jdff dff_A_KYOOwmgG7_0(.dout(w_dff_A_6bamHLNX1_0),.din(w_dff_A_KYOOwmgG7_0),.clk(gclk));
	jdff dff_A_3fPnOUAI5_0(.dout(w_dff_A_KYOOwmgG7_0),.din(w_dff_A_3fPnOUAI5_0),.clk(gclk));
	jdff dff_B_3aDczcGY4_0(.din(n582),.dout(w_dff_B_3aDczcGY4_0),.clk(gclk));
	jdff dff_B_9kVB0bVY5_0(.din(G135),.dout(w_dff_B_9kVB0bVY5_0),.clk(gclk));
	jdff dff_B_YkQHhCKw0_2(.din(n580),.dout(w_dff_B_YkQHhCKw0_2),.clk(gclk));
	jdff dff_B_4m3qZeri9_2(.din(w_dff_B_YkQHhCKw0_2),.dout(w_dff_B_4m3qZeri9_2),.clk(gclk));
	jdff dff_A_jGDrnAcx1_0(.dout(w_G2230_1[0]),.din(w_dff_A_jGDrnAcx1_0),.clk(gclk));
	jdff dff_A_LwacJX3S2_0(.dout(w_dff_A_jGDrnAcx1_0),.din(w_dff_A_LwacJX3S2_0),.clk(gclk));
	jdff dff_A_KWi8CPzx4_0(.dout(w_dff_A_LwacJX3S2_0),.din(w_dff_A_KWi8CPzx4_0),.clk(gclk));
	jdff dff_A_ivVSklLk1_0(.dout(w_dff_A_KWi8CPzx4_0),.din(w_dff_A_ivVSklLk1_0),.clk(gclk));
	jdff dff_A_U5qfBbV10_0(.dout(w_n578_1[0]),.din(w_dff_A_U5qfBbV10_0),.clk(gclk));
	jdff dff_A_HocFgn0q5_0(.dout(w_dff_A_U5qfBbV10_0),.din(w_dff_A_HocFgn0q5_0),.clk(gclk));
	jdff dff_A_NUNImgY63_0(.dout(w_dff_A_HocFgn0q5_0),.din(w_dff_A_NUNImgY63_0),.clk(gclk));
	jdff dff_A_3jTbFiWp1_0(.dout(w_dff_A_NUNImgY63_0),.din(w_dff_A_3jTbFiWp1_0),.clk(gclk));
	jdff dff_A_EpI35P097_0(.dout(w_dff_A_3jTbFiWp1_0),.din(w_dff_A_EpI35P097_0),.clk(gclk));
	jdff dff_A_SInSAymw0_0(.dout(w_dff_A_EpI35P097_0),.din(w_dff_A_SInSAymw0_0),.clk(gclk));
	jdff dff_A_ICPYsPUf0_0(.dout(w_dff_A_SInSAymw0_0),.din(w_dff_A_ICPYsPUf0_0),.clk(gclk));
	jdff dff_A_0vIhUAtM6_0(.dout(w_dff_A_ICPYsPUf0_0),.din(w_dff_A_0vIhUAtM6_0),.clk(gclk));
	jdff dff_A_958fcH956_0(.dout(w_dff_A_0vIhUAtM6_0),.din(w_dff_A_958fcH956_0),.clk(gclk));
	jdff dff_A_7pKwJ1Y80_0(.dout(w_dff_A_958fcH956_0),.din(w_dff_A_7pKwJ1Y80_0),.clk(gclk));
	jdff dff_A_n07Ayx659_0(.dout(w_dff_A_7pKwJ1Y80_0),.din(w_dff_A_n07Ayx659_0),.clk(gclk));
	jdff dff_A_9gZkPiu00_0(.dout(w_dff_A_n07Ayx659_0),.din(w_dff_A_9gZkPiu00_0),.clk(gclk));
	jdff dff_A_cUNyhs7f3_1(.dout(w_n578_0[1]),.din(w_dff_A_cUNyhs7f3_1),.clk(gclk));
	jdff dff_A_sBX2iUXP2_1(.dout(w_dff_A_cUNyhs7f3_1),.din(w_dff_A_sBX2iUXP2_1),.clk(gclk));
	jdff dff_A_5n4RnWEL6_1(.dout(w_dff_A_sBX2iUXP2_1),.din(w_dff_A_5n4RnWEL6_1),.clk(gclk));
	jdff dff_A_6gxuXLXQ4_1(.dout(w_dff_A_5n4RnWEL6_1),.din(w_dff_A_6gxuXLXQ4_1),.clk(gclk));
	jdff dff_A_ZevnK9nJ6_2(.dout(w_n578_0[2]),.din(w_dff_A_ZevnK9nJ6_2),.clk(gclk));
	jdff dff_A_JrS3Fiud8_2(.dout(w_dff_A_ZevnK9nJ6_2),.din(w_dff_A_JrS3Fiud8_2),.clk(gclk));
	jdff dff_A_vYQiPYYA5_2(.dout(w_dff_A_JrS3Fiud8_2),.din(w_dff_A_vYQiPYYA5_2),.clk(gclk));
	jdff dff_A_PjzYXQo94_2(.dout(w_dff_A_vYQiPYYA5_2),.din(w_dff_A_PjzYXQo94_2),.clk(gclk));
	jdff dff_A_coFkWsRA8_2(.dout(w_dff_A_PjzYXQo94_2),.din(w_dff_A_coFkWsRA8_2),.clk(gclk));
	jdff dff_A_CRZCnrDa6_2(.dout(w_dff_A_coFkWsRA8_2),.din(w_dff_A_CRZCnrDa6_2),.clk(gclk));
	jdff dff_A_UA2YDocM0_2(.dout(w_dff_A_CRZCnrDa6_2),.din(w_dff_A_UA2YDocM0_2),.clk(gclk));
	jdff dff_A_Gpzedp2Q0_2(.dout(w_dff_A_UA2YDocM0_2),.din(w_dff_A_Gpzedp2Q0_2),.clk(gclk));
	jdff dff_A_6xvmeIWB7_2(.dout(w_dff_A_Gpzedp2Q0_2),.din(w_dff_A_6xvmeIWB7_2),.clk(gclk));
	jdff dff_A_TR7IL9VK4_2(.dout(w_dff_A_6xvmeIWB7_2),.din(w_dff_A_TR7IL9VK4_2),.clk(gclk));
	jdff dff_A_n0ESUz6X3_2(.dout(w_dff_A_TR7IL9VK4_2),.din(w_dff_A_n0ESUz6X3_2),.clk(gclk));
	jdff dff_A_OjqN8yyk2_2(.dout(w_dff_A_n0ESUz6X3_2),.din(w_dff_A_OjqN8yyk2_2),.clk(gclk));
	jdff dff_B_0zBk2jvP7_0(.din(n576),.dout(w_dff_B_0zBk2jvP7_0),.clk(gclk));
	jdff dff_B_8B9DvCFK8_0(.din(G147),.dout(w_dff_B_8B9DvCFK8_0),.clk(gclk));
	jdff dff_B_PXXc8GBO5_2(.din(n574),.dout(w_dff_B_PXXc8GBO5_2),.clk(gclk));
	jdff dff_B_RLctYm3i2_2(.din(w_dff_B_PXXc8GBO5_2),.dout(w_dff_B_RLctYm3i2_2),.clk(gclk));
	jdff dff_A_BLKIIpEP7_2(.dout(w_n573_0[2]),.din(w_dff_A_BLKIIpEP7_2),.clk(gclk));
	jdff dff_A_PVoVcUMl6_2(.dout(w_dff_A_BLKIIpEP7_2),.din(w_dff_A_PVoVcUMl6_2),.clk(gclk));
	jdff dff_A_FCQ6gevJ6_2(.dout(w_dff_A_PVoVcUMl6_2),.din(w_dff_A_FCQ6gevJ6_2),.clk(gclk));
	jdff dff_A_ZvkmHsyq6_2(.dout(w_dff_A_FCQ6gevJ6_2),.din(w_dff_A_ZvkmHsyq6_2),.clk(gclk));
	jdff dff_A_nTbbieea2_2(.dout(w_dff_A_ZvkmHsyq6_2),.din(w_dff_A_nTbbieea2_2),.clk(gclk));
	jdff dff_A_gKcfYQCM3_2(.dout(w_dff_A_nTbbieea2_2),.din(w_dff_A_gKcfYQCM3_2),.clk(gclk));
	jdff dff_A_JZJusJjl4_2(.dout(w_dff_A_gKcfYQCM3_2),.din(w_dff_A_JZJusJjl4_2),.clk(gclk));
	jdff dff_A_0qeCP5Pi8_2(.dout(w_dff_A_JZJusJjl4_2),.din(w_dff_A_0qeCP5Pi8_2),.clk(gclk));
	jdff dff_A_Ab2DlB5i8_2(.dout(w_dff_A_0qeCP5Pi8_2),.din(w_dff_A_Ab2DlB5i8_2),.clk(gclk));
	jdff dff_A_B5DfgghN8_2(.dout(w_dff_A_Ab2DlB5i8_2),.din(w_dff_A_B5DfgghN8_2),.clk(gclk));
	jdff dff_A_AL7tSTXe6_2(.dout(w_dff_A_B5DfgghN8_2),.din(w_dff_A_AL7tSTXe6_2),.clk(gclk));
	jdff dff_A_8NK7dJPs5_2(.dout(w_dff_A_AL7tSTXe6_2),.din(w_dff_A_8NK7dJPs5_2),.clk(gclk));
	jdff dff_A_7VhT2UQB1_2(.dout(w_dff_A_8NK7dJPs5_2),.din(w_dff_A_7VhT2UQB1_2),.clk(gclk));
	jdff dff_A_Gqf84gAp9_2(.dout(w_dff_A_7VhT2UQB1_2),.din(w_dff_A_Gqf84gAp9_2),.clk(gclk));
	jdff dff_A_eyU1szws7_2(.dout(w_n572_0[2]),.din(w_dff_A_eyU1szws7_2),.clk(gclk));
	jdff dff_B_qkHOgTH72_0(.din(n571),.dout(w_dff_B_qkHOgTH72_0),.clk(gclk));
	jdff dff_B_YG35GxyW3_0(.din(G138),.dout(w_dff_B_YG35GxyW3_0),.clk(gclk));
	jdff dff_B_PEQ9VT1z2_3(.din(n569),.dout(w_dff_B_PEQ9VT1z2_3),.clk(gclk));
	jdff dff_B_PQGBc40z6_3(.din(w_dff_B_PEQ9VT1z2_3),.dout(w_dff_B_PQGBc40z6_3),.clk(gclk));
	jdff dff_A_MRFqdrPo2_0(.dout(w_n568_0[0]),.din(w_dff_A_MRFqdrPo2_0),.clk(gclk));
	jdff dff_A_krJLXUrV1_0(.dout(w_dff_A_MRFqdrPo2_0),.din(w_dff_A_krJLXUrV1_0),.clk(gclk));
	jdff dff_A_txuTezv14_0(.dout(w_dff_A_krJLXUrV1_0),.din(w_dff_A_txuTezv14_0),.clk(gclk));
	jdff dff_A_VNCGnUvp7_0(.dout(w_dff_A_txuTezv14_0),.din(w_dff_A_VNCGnUvp7_0),.clk(gclk));
	jdff dff_A_jxIX0lJ19_2(.dout(w_n568_0[2]),.din(w_dff_A_jxIX0lJ19_2),.clk(gclk));
	jdff dff_A_aV5KfnpY0_2(.dout(w_dff_A_jxIX0lJ19_2),.din(w_dff_A_aV5KfnpY0_2),.clk(gclk));
	jdff dff_B_fEbOTJcJ7_0(.din(G157),.dout(w_dff_B_fEbOTJcJ7_0),.clk(gclk));
	jdff dff_A_MNG6Rabt6_0(.dout(w_n564_0[0]),.din(w_dff_A_MNG6Rabt6_0),.clk(gclk));
	jdff dff_A_6wKJ42DQ3_0(.dout(w_dff_A_MNG6Rabt6_0),.din(w_dff_A_6wKJ42DQ3_0),.clk(gclk));
	jdff dff_A_M2g0VMm52_0(.dout(w_dff_A_6wKJ42DQ3_0),.din(w_dff_A_M2g0VMm52_0),.clk(gclk));
	jdff dff_A_pDl1u0AP0_1(.dout(w_n564_0[1]),.din(w_dff_A_pDl1u0AP0_1),.clk(gclk));
	jdff dff_B_r5qQAagg4_2(.din(n563),.dout(w_dff_B_r5qQAagg4_2),.clk(gclk));
	jdff dff_B_EfYlwM1z4_2(.din(w_dff_B_r5qQAagg4_2),.dout(w_dff_B_EfYlwM1z4_2),.clk(gclk));
	jdff dff_A_vtTJ75Jn1_0(.dout(w_G2236_1[0]),.din(w_dff_A_vtTJ75Jn1_0),.clk(gclk));
	jdff dff_A_jXPJP4Ul0_0(.dout(w_dff_A_vtTJ75Jn1_0),.din(w_dff_A_jXPJP4Ul0_0),.clk(gclk));
	jdff dff_A_jlNxoxLR6_0(.dout(w_dff_A_jXPJP4Ul0_0),.din(w_dff_A_jlNxoxLR6_0),.clk(gclk));
	jdff dff_A_jLE2n0rJ9_0(.dout(w_dff_A_jlNxoxLR6_0),.din(w_dff_A_jLE2n0rJ9_0),.clk(gclk));
	jdff dff_B_xQBl0tyx8_0(.din(n561),.dout(w_dff_B_xQBl0tyx8_0),.clk(gclk));
	jdff dff_B_DGXLujUx0_0(.din(w_dff_B_xQBl0tyx8_0),.dout(w_dff_B_DGXLujUx0_0),.clk(gclk));
	jdff dff_B_EeZCxGzL1_0(.din(w_dff_B_DGXLujUx0_0),.dout(w_dff_B_EeZCxGzL1_0),.clk(gclk));
	jdff dff_B_LlkusSHQ2_0(.din(w_dff_B_EeZCxGzL1_0),.dout(w_dff_B_LlkusSHQ2_0),.clk(gclk));
	jdff dff_A_YNiCY31p0_0(.dout(w_n560_0[0]),.din(w_dff_A_YNiCY31p0_0),.clk(gclk));
	jdff dff_A_5OV1dwPW1_0(.dout(w_dff_A_YNiCY31p0_0),.din(w_dff_A_5OV1dwPW1_0),.clk(gclk));
	jdff dff_A_FBZQshe61_0(.dout(w_dff_A_5OV1dwPW1_0),.din(w_dff_A_FBZQshe61_0),.clk(gclk));
	jdff dff_A_ABp5S7ct5_0(.dout(w_dff_A_FBZQshe61_0),.din(w_dff_A_ABp5S7ct5_0),.clk(gclk));
	jdff dff_A_QUz8ApJj9_0(.dout(w_dff_A_ABp5S7ct5_0),.din(w_dff_A_QUz8ApJj9_0),.clk(gclk));
	jdff dff_B_2x7k6Izw8_1(.din(n547),.dout(w_dff_B_2x7k6Izw8_1),.clk(gclk));
	jdff dff_B_m5qLykB48_1(.din(w_dff_B_2x7k6Izw8_1),.dout(w_dff_B_m5qLykB48_1),.clk(gclk));
	jdff dff_B_JtxtzyDc6_1(.din(w_dff_B_m5qLykB48_1),.dout(w_dff_B_JtxtzyDc6_1),.clk(gclk));
	jdff dff_B_VooOvSZ25_1(.din(n548),.dout(w_dff_B_VooOvSZ25_1),.clk(gclk));
	jdff dff_B_OzIA1lgn4_1(.din(w_dff_B_VooOvSZ25_1),.dout(w_dff_B_OzIA1lgn4_1),.clk(gclk));
	jdff dff_B_ol73AUFQ1_1(.din(w_dff_B_OzIA1lgn4_1),.dout(w_dff_B_ol73AUFQ1_1),.clk(gclk));
	jdff dff_B_OM3RWix06_1(.din(w_dff_B_ol73AUFQ1_1),.dout(w_dff_B_OM3RWix06_1),.clk(gclk));
	jdff dff_B_Zg42mpPj3_0(.din(n543),.dout(w_dff_B_Zg42mpPj3_0),.clk(gclk));
	jdff dff_B_YfdNglBp5_0(.din(w_dff_B_Zg42mpPj3_0),.dout(w_dff_B_YfdNglBp5_0),.clk(gclk));
	jdff dff_B_780b8s1n6_0(.din(w_dff_B_YfdNglBp5_0),.dout(w_dff_B_780b8s1n6_0),.clk(gclk));
	jdff dff_B_ISB3JEFm3_0(.din(w_dff_B_780b8s1n6_0),.dout(w_dff_B_ISB3JEFm3_0),.clk(gclk));
	jdff dff_B_PYnusFwX1_0(.din(w_dff_B_ISB3JEFm3_0),.dout(w_dff_B_PYnusFwX1_0),.clk(gclk));
	jdff dff_B_EIEfZT132_0(.din(w_dff_B_PYnusFwX1_0),.dout(w_dff_B_EIEfZT132_0),.clk(gclk));
	jdff dff_B_o0PEMrjh5_0(.din(w_dff_B_EIEfZT132_0),.dout(w_dff_B_o0PEMrjh5_0),.clk(gclk));
	jdff dff_A_gA2jriS08_0(.dout(w_n542_0[0]),.din(w_dff_A_gA2jriS08_0),.clk(gclk));
	jdff dff_A_XeLStNUO4_0(.dout(w_dff_A_gA2jriS08_0),.din(w_dff_A_XeLStNUO4_0),.clk(gclk));
	jdff dff_A_7IJbK2cu0_0(.dout(w_dff_A_XeLStNUO4_0),.din(w_dff_A_7IJbK2cu0_0),.clk(gclk));
	jdff dff_A_cox8FrSk7_0(.dout(w_dff_A_7IJbK2cu0_0),.din(w_dff_A_cox8FrSk7_0),.clk(gclk));
	jdff dff_A_y9PMKQPI2_0(.dout(w_dff_A_cox8FrSk7_0),.din(w_dff_A_y9PMKQPI2_0),.clk(gclk));
	jdff dff_A_0RPCVCxN5_0(.dout(w_dff_A_y9PMKQPI2_0),.din(w_dff_A_0RPCVCxN5_0),.clk(gclk));
	jdff dff_A_fbNsijmB8_0(.dout(w_dff_A_0RPCVCxN5_0),.din(w_dff_A_fbNsijmB8_0),.clk(gclk));
	jdff dff_A_Zh6HOU566_0(.dout(w_dff_A_fbNsijmB8_0),.din(w_dff_A_Zh6HOU566_0),.clk(gclk));
	jdff dff_A_X6FvcRRw4_0(.dout(w_n535_1[0]),.din(w_dff_A_X6FvcRRw4_0),.clk(gclk));
	jdff dff_A_0Evq6HH87_0(.dout(w_dff_A_X6FvcRRw4_0),.din(w_dff_A_0Evq6HH87_0),.clk(gclk));
	jdff dff_A_HZIoMgTR1_0(.dout(w_dff_A_0Evq6HH87_0),.din(w_dff_A_HZIoMgTR1_0),.clk(gclk));
	jdff dff_A_KNh9Uhix2_0(.dout(w_dff_A_HZIoMgTR1_0),.din(w_dff_A_KNh9Uhix2_0),.clk(gclk));
	jdff dff_A_MoaKYuRC0_0(.dout(w_dff_A_KNh9Uhix2_0),.din(w_dff_A_MoaKYuRC0_0),.clk(gclk));
	jdff dff_A_LmPmyEAH3_0(.dout(w_dff_A_MoaKYuRC0_0),.din(w_dff_A_LmPmyEAH3_0),.clk(gclk));
	jdff dff_A_NJxuuXfY2_0(.dout(w_dff_A_LmPmyEAH3_0),.din(w_dff_A_NJxuuXfY2_0),.clk(gclk));
	jdff dff_A_tg3J5Qw19_0(.dout(w_dff_A_NJxuuXfY2_0),.din(w_dff_A_tg3J5Qw19_0),.clk(gclk));
	jdff dff_A_u3O8q0dd0_0(.dout(w_dff_A_tg3J5Qw19_0),.din(w_dff_A_u3O8q0dd0_0),.clk(gclk));
	jdff dff_A_nNYgLdSa5_0(.dout(w_dff_A_u3O8q0dd0_0),.din(w_dff_A_nNYgLdSa5_0),.clk(gclk));
	jdff dff_A_SgbzgMBx0_0(.dout(w_dff_A_nNYgLdSa5_0),.din(w_dff_A_SgbzgMBx0_0),.clk(gclk));
	jdff dff_A_xZRp3sQ61_0(.dout(w_dff_A_SgbzgMBx0_0),.din(w_dff_A_xZRp3sQ61_0),.clk(gclk));
	jdff dff_A_HBeBFwuV4_0(.dout(w_dff_A_xZRp3sQ61_0),.din(w_dff_A_HBeBFwuV4_0),.clk(gclk));
	jdff dff_A_RV9OZxoL4_0(.dout(w_n530_0[0]),.din(w_dff_A_RV9OZxoL4_0),.clk(gclk));
	jdff dff_A_cZaE98gp3_0(.dout(w_dff_A_RV9OZxoL4_0),.din(w_dff_A_cZaE98gp3_0),.clk(gclk));
	jdff dff_A_J3trp0RF9_0(.dout(w_dff_A_cZaE98gp3_0),.din(w_dff_A_J3trp0RF9_0),.clk(gclk));
	jdff dff_A_Q2OfWQ9W8_0(.dout(w_dff_A_J3trp0RF9_0),.din(w_dff_A_Q2OfWQ9W8_0),.clk(gclk));
	jdff dff_A_D5xr9PFH4_0(.dout(w_dff_A_Q2OfWQ9W8_0),.din(w_dff_A_D5xr9PFH4_0),.clk(gclk));
	jdff dff_A_sFRKSLiG5_0(.dout(w_dff_A_D5xr9PFH4_0),.din(w_dff_A_sFRKSLiG5_0),.clk(gclk));
	jdff dff_A_bV9CZwQh1_0(.dout(w_dff_A_sFRKSLiG5_0),.din(w_dff_A_bV9CZwQh1_0),.clk(gclk));
	jdff dff_A_m509t6VE6_0(.dout(w_dff_A_bV9CZwQh1_0),.din(w_dff_A_m509t6VE6_0),.clk(gclk));
	jdff dff_A_Khm9731N6_0(.dout(w_dff_A_m509t6VE6_0),.din(w_dff_A_Khm9731N6_0),.clk(gclk));
	jdff dff_A_t4sFYymZ0_0(.dout(w_n529_0[0]),.din(w_dff_A_t4sFYymZ0_0),.clk(gclk));
	jdff dff_A_AOmBRrzc7_0(.dout(w_dff_A_t4sFYymZ0_0),.din(w_dff_A_AOmBRrzc7_0),.clk(gclk));
	jdff dff_A_qa52qAz58_0(.dout(w_dff_A_AOmBRrzc7_0),.din(w_dff_A_qa52qAz58_0),.clk(gclk));
	jdff dff_A_dZUBlL9L3_0(.dout(w_dff_A_qa52qAz58_0),.din(w_dff_A_dZUBlL9L3_0),.clk(gclk));
	jdff dff_A_6x7fUC5X2_0(.dout(w_dff_A_dZUBlL9L3_0),.din(w_dff_A_6x7fUC5X2_0),.clk(gclk));
	jdff dff_A_yZyCMx2o7_0(.dout(w_dff_A_6x7fUC5X2_0),.din(w_dff_A_yZyCMx2o7_0),.clk(gclk));
	jdff dff_A_d1M3wBli3_0(.dout(w_dff_A_yZyCMx2o7_0),.din(w_dff_A_d1M3wBli3_0),.clk(gclk));
	jdff dff_A_x9XEglM08_0(.dout(w_dff_A_d1M3wBli3_0),.din(w_dff_A_x9XEglM08_0),.clk(gclk));
	jdff dff_A_9LvIBP7d9_0(.dout(w_dff_A_x9XEglM08_0),.din(w_dff_A_9LvIBP7d9_0),.clk(gclk));
	jdff dff_A_cHaWjaGn3_0(.dout(w_dff_A_9LvIBP7d9_0),.din(w_dff_A_cHaWjaGn3_0),.clk(gclk));
	jdff dff_A_t4HvP0Lb3_0(.dout(w_n1463_0[0]),.din(w_dff_A_t4HvP0Lb3_0),.clk(gclk));
	jdff dff_A_M7PvdOKY1_0(.dout(w_dff_A_t4HvP0Lb3_0),.din(w_dff_A_M7PvdOKY1_0),.clk(gclk));
	jdff dff_A_Ic3AEWiT2_0(.dout(w_dff_A_M7PvdOKY1_0),.din(w_dff_A_Ic3AEWiT2_0),.clk(gclk));
	jdff dff_A_JHH89ISz2_0(.dout(w_dff_A_Ic3AEWiT2_0),.din(w_dff_A_JHH89ISz2_0),.clk(gclk));
	jdff dff_A_f3vWnTh30_0(.dout(w_dff_A_JHH89ISz2_0),.din(w_dff_A_f3vWnTh30_0),.clk(gclk));
	jdff dff_A_5pIYaN4v3_0(.dout(w_dff_A_f3vWnTh30_0),.din(w_dff_A_5pIYaN4v3_0),.clk(gclk));
	jdff dff_A_NEib7nIp7_0(.dout(w_dff_A_5pIYaN4v3_0),.din(w_dff_A_NEib7nIp7_0),.clk(gclk));
	jdff dff_A_a2yjqdUT8_0(.dout(w_dff_A_NEib7nIp7_0),.din(w_dff_A_a2yjqdUT8_0),.clk(gclk));
	jdff dff_A_lneF3gDB1_0(.dout(w_dff_A_a2yjqdUT8_0),.din(w_dff_A_lneF3gDB1_0),.clk(gclk));
	jdff dff_A_QA9ZD07p6_0(.dout(w_dff_A_lneF3gDB1_0),.din(w_dff_A_QA9ZD07p6_0),.clk(gclk));
	jdff dff_A_lOhW6SaF6_0(.dout(w_dff_A_QA9ZD07p6_0),.din(w_dff_A_lOhW6SaF6_0),.clk(gclk));
	jdff dff_A_Cin2kwwM7_1(.dout(w_n1463_0[1]),.din(w_dff_A_Cin2kwwM7_1),.clk(gclk));
	jdff dff_A_cbOkA64P4_1(.dout(w_dff_A_Cin2kwwM7_1),.din(w_dff_A_cbOkA64P4_1),.clk(gclk));
	jdff dff_A_JQ0S1JPM9_1(.dout(w_dff_A_cbOkA64P4_1),.din(w_dff_A_JQ0S1JPM9_1),.clk(gclk));
	jdff dff_A_5iLq8Cye5_1(.dout(w_dff_A_JQ0S1JPM9_1),.din(w_dff_A_5iLq8Cye5_1),.clk(gclk));
	jdff dff_A_SzJHuo2M9_1(.dout(w_dff_A_5iLq8Cye5_1),.din(w_dff_A_SzJHuo2M9_1),.clk(gclk));
	jdff dff_A_coXT6OT86_1(.dout(w_dff_A_SzJHuo2M9_1),.din(w_dff_A_coXT6OT86_1),.clk(gclk));
	jdff dff_A_z00A8m8a4_1(.dout(w_dff_A_coXT6OT86_1),.din(w_dff_A_z00A8m8a4_1),.clk(gclk));
	jdff dff_A_uzKLdXwp8_1(.dout(w_dff_A_z00A8m8a4_1),.din(w_dff_A_uzKLdXwp8_1),.clk(gclk));
	jdff dff_A_kcUFjEsL6_1(.dout(w_dff_A_uzKLdXwp8_1),.din(w_dff_A_kcUFjEsL6_1),.clk(gclk));
	jdff dff_A_H2UhE8jp1_1(.dout(w_dff_A_kcUFjEsL6_1),.din(w_dff_A_H2UhE8jp1_1),.clk(gclk));
	jdff dff_A_XAnvY1zi3_1(.dout(w_dff_A_H2UhE8jp1_1),.din(w_dff_A_XAnvY1zi3_1),.clk(gclk));
	jdff dff_A_PY4Dn2pN8_1(.dout(w_dff_A_XAnvY1zi3_1),.din(w_dff_A_PY4Dn2pN8_1),.clk(gclk));
	jdff dff_A_E8pfDTvF5_1(.dout(w_dff_A_PY4Dn2pN8_1),.din(w_dff_A_E8pfDTvF5_1),.clk(gclk));
	jdff dff_A_MTjSPOR93_1(.dout(w_dff_A_E8pfDTvF5_1),.din(w_dff_A_MTjSPOR93_1),.clk(gclk));
	jdff dff_A_i6EBz8z02_1(.dout(w_dff_A_MTjSPOR93_1),.din(w_dff_A_i6EBz8z02_1),.clk(gclk));
	jdff dff_A_RdIulqLn6_1(.dout(w_dff_A_i6EBz8z02_1),.din(w_dff_A_RdIulqLn6_1),.clk(gclk));
	jdff dff_A_ce52Zyu94_1(.dout(w_dff_A_RdIulqLn6_1),.din(w_dff_A_ce52Zyu94_1),.clk(gclk));
	jdff dff_A_ZDgOUspn3_1(.dout(w_dff_A_ce52Zyu94_1),.din(w_dff_A_ZDgOUspn3_1),.clk(gclk));
	jdff dff_A_s5cqszX06_1(.dout(w_dff_A_ZDgOUspn3_1),.din(w_dff_A_s5cqszX06_1),.clk(gclk));
	jdff dff_B_rN5cNUVh2_0(.din(n1462),.dout(w_dff_B_rN5cNUVh2_0),.clk(gclk));
	jdff dff_A_yRaGuZBV6_1(.dout(w_n365_0[1]),.din(w_dff_A_yRaGuZBV6_1),.clk(gclk));
	jdff dff_A_jCNZtjfD1_1(.dout(w_dff_A_yRaGuZBV6_1),.din(w_dff_A_jCNZtjfD1_1),.clk(gclk));
	jdff dff_A_EAf0qjq49_1(.dout(w_dff_A_jCNZtjfD1_1),.din(w_dff_A_EAf0qjq49_1),.clk(gclk));
	jdff dff_A_HUXqwlAR4_1(.dout(w_dff_A_EAf0qjq49_1),.din(w_dff_A_HUXqwlAR4_1),.clk(gclk));
	jdff dff_A_eufje9bP7_1(.dout(w_dff_A_HUXqwlAR4_1),.din(w_dff_A_eufje9bP7_1),.clk(gclk));
	jdff dff_A_zZdGEytR0_1(.dout(w_dff_A_eufje9bP7_1),.din(w_dff_A_zZdGEytR0_1),.clk(gclk));
	jdff dff_A_eenzGgUX0_1(.dout(w_dff_A_zZdGEytR0_1),.din(w_dff_A_eenzGgUX0_1),.clk(gclk));
	jdff dff_A_jh9KSGLR7_1(.dout(w_dff_A_eenzGgUX0_1),.din(w_dff_A_jh9KSGLR7_1),.clk(gclk));
	jdff dff_A_p99mBJgi9_1(.dout(w_dff_A_jh9KSGLR7_1),.din(w_dff_A_p99mBJgi9_1),.clk(gclk));
	jdff dff_A_oxfc5nJO4_1(.dout(w_dff_A_p99mBJgi9_1),.din(w_dff_A_oxfc5nJO4_1),.clk(gclk));
	jdff dff_A_2G0y3i8v0_1(.dout(w_dff_A_oxfc5nJO4_1),.din(w_dff_A_2G0y3i8v0_1),.clk(gclk));
	jdff dff_A_vR7pSnCd3_1(.dout(w_dff_A_2G0y3i8v0_1),.din(w_dff_A_vR7pSnCd3_1),.clk(gclk));
	jdff dff_A_6P8zEAdh0_1(.dout(w_dff_A_vR7pSnCd3_1),.din(w_dff_A_6P8zEAdh0_1),.clk(gclk));
	jdff dff_A_vjXGWoYN2_1(.dout(w_dff_A_6P8zEAdh0_1),.din(w_dff_A_vjXGWoYN2_1),.clk(gclk));
	jdff dff_A_SbRehflK6_1(.dout(w_dff_A_vjXGWoYN2_1),.din(w_dff_A_SbRehflK6_1),.clk(gclk));
	jdff dff_A_EKRQMMUG3_1(.dout(w_dff_A_SbRehflK6_1),.din(w_dff_A_EKRQMMUG3_1),.clk(gclk));
	jdff dff_A_5UtrnW0b2_1(.dout(w_dff_A_EKRQMMUG3_1),.din(w_dff_A_5UtrnW0b2_1),.clk(gclk));
	jdff dff_A_tYEP0C1I7_1(.dout(w_dff_A_5UtrnW0b2_1),.din(w_dff_A_tYEP0C1I7_1),.clk(gclk));
	jdff dff_A_zrpSyQ9n2_1(.dout(w_dff_A_tYEP0C1I7_1),.din(w_dff_A_zrpSyQ9n2_1),.clk(gclk));
	jdff dff_A_9gAtgxeD5_1(.dout(w_dff_A_zrpSyQ9n2_1),.din(w_dff_A_9gAtgxeD5_1),.clk(gclk));
	jdff dff_A_8jy4uN992_1(.dout(w_dff_A_9gAtgxeD5_1),.din(w_dff_A_8jy4uN992_1),.clk(gclk));
	jdff dff_A_k4RWJ9WP6_0(.dout(w_G38_1[0]),.din(w_dff_A_k4RWJ9WP6_0),.clk(gclk));
	jdff dff_A_6US0F5m16_0(.dout(w_dff_A_k4RWJ9WP6_0),.din(w_dff_A_6US0F5m16_0),.clk(gclk));
	jdff dff_A_3uwX3wIX5_0(.dout(w_dff_A_6US0F5m16_0),.din(w_dff_A_3uwX3wIX5_0),.clk(gclk));
	jdff dff_A_SMU084j52_2(.dout(w_G38_1[2]),.din(w_dff_A_SMU084j52_2),.clk(gclk));
	jdff dff_A_RMHGHZKQ8_1(.dout(w_G38_0[1]),.din(w_dff_A_RMHGHZKQ8_1),.clk(gclk));
	jdff dff_A_qtVxapno2_2(.dout(w_G38_0[2]),.din(w_dff_A_qtVxapno2_2),.clk(gclk));
	jdff dff_A_nW69HDsr6_2(.dout(w_dff_A_qtVxapno2_2),.din(w_dff_A_nW69HDsr6_2),.clk(gclk));
	jdff dff_B_jRtvoOkf6_1(.din(n1587),.dout(w_dff_B_jRtvoOkf6_1),.clk(gclk));
	jdff dff_B_3dmKPqL63_1(.din(w_dff_B_jRtvoOkf6_1),.dout(w_dff_B_3dmKPqL63_1),.clk(gclk));
	jdff dff_B_yvlUL8yN0_1(.din(w_dff_B_3dmKPqL63_1),.dout(w_dff_B_yvlUL8yN0_1),.clk(gclk));
	jdff dff_B_cfCD5Gl36_1(.din(w_dff_B_yvlUL8yN0_1),.dout(w_dff_B_cfCD5Gl36_1),.clk(gclk));
	jdff dff_B_16f7dWCt9_1(.din(w_dff_B_cfCD5Gl36_1),.dout(w_dff_B_16f7dWCt9_1),.clk(gclk));
	jdff dff_B_W7q1z4qJ7_1(.din(w_dff_B_16f7dWCt9_1),.dout(w_dff_B_W7q1z4qJ7_1),.clk(gclk));
	jdff dff_B_Ckxr55D59_1(.din(w_dff_B_W7q1z4qJ7_1),.dout(w_dff_B_Ckxr55D59_1),.clk(gclk));
	jdff dff_B_mq7toIlo6_1(.din(w_dff_B_Ckxr55D59_1),.dout(w_dff_B_mq7toIlo6_1),.clk(gclk));
	jdff dff_B_d4AAX7vs6_1(.din(w_dff_B_mq7toIlo6_1),.dout(w_dff_B_d4AAX7vs6_1),.clk(gclk));
	jdff dff_B_v0fKB7sD8_1(.din(w_dff_B_d4AAX7vs6_1),.dout(w_dff_B_v0fKB7sD8_1),.clk(gclk));
	jdff dff_B_JHDTJUgh7_1(.din(w_dff_B_v0fKB7sD8_1),.dout(w_dff_B_JHDTJUgh7_1),.clk(gclk));
	jdff dff_B_mcI2YI0y3_1(.din(w_dff_B_JHDTJUgh7_1),.dout(w_dff_B_mcI2YI0y3_1),.clk(gclk));
	jdff dff_B_FhF1XEca0_1(.din(n1606),.dout(w_dff_B_FhF1XEca0_1),.clk(gclk));
	jdff dff_B_VDYO2Rpt6_1(.din(w_dff_B_FhF1XEca0_1),.dout(w_dff_B_VDYO2Rpt6_1),.clk(gclk));
	jdff dff_B_dnpg8Gl39_1(.din(n1620),.dout(w_dff_B_dnpg8Gl39_1),.clk(gclk));
	jdff dff_B_9R9VV1R75_1(.din(w_dff_B_dnpg8Gl39_1),.dout(w_dff_B_9R9VV1R75_1),.clk(gclk));
	jdff dff_B_K53FRdr76_1(.din(n1622),.dout(w_dff_B_K53FRdr76_1),.clk(gclk));
	jdff dff_B_7aDvH7Ol3_1(.din(w_dff_B_K53FRdr76_1),.dout(w_dff_B_7aDvH7Ol3_1),.clk(gclk));
	jdff dff_B_igRn2kT56_1(.din(w_dff_B_7aDvH7Ol3_1),.dout(w_dff_B_igRn2kT56_1),.clk(gclk));
	jdff dff_B_kIUMZ3y72_1(.din(w_dff_B_igRn2kT56_1),.dout(w_dff_B_kIUMZ3y72_1),.clk(gclk));
	jdff dff_B_Tk1X9D675_1(.din(w_dff_B_kIUMZ3y72_1),.dout(w_dff_B_Tk1X9D675_1),.clk(gclk));
	jdff dff_B_MIfDYEr94_1(.din(w_dff_B_Tk1X9D675_1),.dout(w_dff_B_MIfDYEr94_1),.clk(gclk));
	jdff dff_B_7XUiODAV7_1(.din(n1623),.dout(w_dff_B_7XUiODAV7_1),.clk(gclk));
	jdff dff_B_H67iYjbW1_1(.din(w_dff_B_7XUiODAV7_1),.dout(w_dff_B_H67iYjbW1_1),.clk(gclk));
	jdff dff_B_fCfGZnj25_1(.din(w_dff_B_H67iYjbW1_1),.dout(w_dff_B_fCfGZnj25_1),.clk(gclk));
	jdff dff_B_GOcO4ZDS3_1(.din(w_dff_B_fCfGZnj25_1),.dout(w_dff_B_GOcO4ZDS3_1),.clk(gclk));
	jdff dff_B_YRuKFWpL5_1(.din(w_dff_B_GOcO4ZDS3_1),.dout(w_dff_B_YRuKFWpL5_1),.clk(gclk));
	jdff dff_B_O32HxyCm5_1(.din(w_dff_B_YRuKFWpL5_1),.dout(w_dff_B_O32HxyCm5_1),.clk(gclk));
	jdff dff_B_xxEQ6N0d9_1(.din(w_dff_B_O32HxyCm5_1),.dout(w_dff_B_xxEQ6N0d9_1),.clk(gclk));
	jdff dff_B_HgkmMpkq4_1(.din(w_dff_B_xxEQ6N0d9_1),.dout(w_dff_B_HgkmMpkq4_1),.clk(gclk));
	jdff dff_B_t5Q83ilq6_1(.din(n1626),.dout(w_dff_B_t5Q83ilq6_1),.clk(gclk));
	jdff dff_B_N9Vq1s1r7_1(.din(w_dff_B_t5Q83ilq6_1),.dout(w_dff_B_N9Vq1s1r7_1),.clk(gclk));
	jdff dff_B_VeIFWBtK7_0(.din(n1624),.dout(w_dff_B_VeIFWBtK7_0),.clk(gclk));
	jdff dff_B_bBJAt9h86_0(.din(w_dff_B_VeIFWBtK7_0),.dout(w_dff_B_bBJAt9h86_0),.clk(gclk));
	jdff dff_A_sFb5TV286_1(.dout(w_n1479_0[1]),.din(w_dff_A_sFb5TV286_1),.clk(gclk));
	jdff dff_A_8oBhqTHT1_1(.dout(w_dff_A_sFb5TV286_1),.din(w_dff_A_8oBhqTHT1_1),.clk(gclk));
	jdff dff_A_QOxPP0Lv3_1(.dout(w_dff_A_8oBhqTHT1_1),.din(w_dff_A_QOxPP0Lv3_1),.clk(gclk));
	jdff dff_A_lqz8PcDP1_1(.dout(w_dff_A_QOxPP0Lv3_1),.din(w_dff_A_lqz8PcDP1_1),.clk(gclk));
	jdff dff_A_lkSCW3v69_1(.dout(w_dff_A_lqz8PcDP1_1),.din(w_dff_A_lkSCW3v69_1),.clk(gclk));
	jdff dff_A_pe8t0RV05_1(.dout(w_dff_A_lkSCW3v69_1),.din(w_dff_A_pe8t0RV05_1),.clk(gclk));
	jdff dff_A_g9hjSyA09_1(.dout(w_n1471_0[1]),.din(w_dff_A_g9hjSyA09_1),.clk(gclk));
	jdff dff_A_UhRr5FxT5_1(.dout(w_dff_A_g9hjSyA09_1),.din(w_dff_A_UhRr5FxT5_1),.clk(gclk));
	jdff dff_A_xgnpDOvd9_1(.dout(w_dff_A_UhRr5FxT5_1),.din(w_dff_A_xgnpDOvd9_1),.clk(gclk));
	jdff dff_A_zPCfDnca1_1(.dout(w_dff_A_xgnpDOvd9_1),.din(w_dff_A_zPCfDnca1_1),.clk(gclk));
	jdff dff_A_8wgZDwou2_1(.dout(w_dff_A_zPCfDnca1_1),.din(w_dff_A_8wgZDwou2_1),.clk(gclk));
	jdff dff_B_LIg25Xc01_1(.din(n1609),.dout(w_dff_B_LIg25Xc01_1),.clk(gclk));
	jdff dff_B_dPh0iSfw8_1(.din(w_dff_B_LIg25Xc01_1),.dout(w_dff_B_dPh0iSfw8_1),.clk(gclk));
	jdff dff_B_NnsfubA92_1(.din(w_dff_B_dPh0iSfw8_1),.dout(w_dff_B_NnsfubA92_1),.clk(gclk));
	jdff dff_B_tEfZilgs7_1(.din(w_dff_B_NnsfubA92_1),.dout(w_dff_B_tEfZilgs7_1),.clk(gclk));
	jdff dff_B_oosQi0KE3_1(.din(w_dff_B_tEfZilgs7_1),.dout(w_dff_B_oosQi0KE3_1),.clk(gclk));
	jdff dff_B_es06gPn80_1(.din(w_dff_B_oosQi0KE3_1),.dout(w_dff_B_es06gPn80_1),.clk(gclk));
	jdff dff_B_8MEA0ppJ8_0(.din(n1615),.dout(w_dff_B_8MEA0ppJ8_0),.clk(gclk));
	jdff dff_A_zc8s8CG83_1(.dout(w_n1482_0[1]),.din(w_dff_A_zc8s8CG83_1),.clk(gclk));
	jdff dff_A_KvwON2zq1_1(.dout(w_dff_A_zc8s8CG83_1),.din(w_dff_A_KvwON2zq1_1),.clk(gclk));
	jdff dff_A_ryXHJU2R3_1(.dout(w_dff_A_KvwON2zq1_1),.din(w_dff_A_ryXHJU2R3_1),.clk(gclk));
	jdff dff_A_pBDT5ZAl5_1(.dout(w_dff_A_ryXHJU2R3_1),.din(w_dff_A_pBDT5ZAl5_1),.clk(gclk));
	jdff dff_A_HVlgAT7E0_1(.dout(w_dff_A_pBDT5ZAl5_1),.din(w_dff_A_HVlgAT7E0_1),.clk(gclk));
	jdff dff_A_45qkWINe8_1(.dout(w_dff_A_HVlgAT7E0_1),.din(w_dff_A_45qkWINe8_1),.clk(gclk));
	jdff dff_A_iLnKSvBK5_1(.dout(w_dff_A_45qkWINe8_1),.din(w_dff_A_iLnKSvBK5_1),.clk(gclk));
	jdff dff_A_ALdcHJPQ8_1(.dout(w_n1468_0[1]),.din(w_dff_A_ALdcHJPQ8_1),.clk(gclk));
	jdff dff_A_SxindvZG8_1(.dout(w_dff_A_ALdcHJPQ8_1),.din(w_dff_A_SxindvZG8_1),.clk(gclk));
	jdff dff_A_q4B4tKmh9_1(.dout(w_dff_A_SxindvZG8_1),.din(w_dff_A_q4B4tKmh9_1),.clk(gclk));
	jdff dff_A_ImXngjWN9_1(.dout(w_dff_A_q4B4tKmh9_1),.din(w_dff_A_ImXngjWN9_1),.clk(gclk));
	jdff dff_A_iKGJ2GEw0_1(.dout(w_dff_A_ImXngjWN9_1),.din(w_dff_A_iKGJ2GEw0_1),.clk(gclk));
	jdff dff_B_9ajlYZdr3_2(.din(n1468),.dout(w_dff_B_9ajlYZdr3_2),.clk(gclk));
	jdff dff_B_invpDyNA8_2(.din(w_dff_B_9ajlYZdr3_2),.dout(w_dff_B_invpDyNA8_2),.clk(gclk));
	jdff dff_B_ZIXfBbNh2_2(.din(w_dff_B_invpDyNA8_2),.dout(w_dff_B_ZIXfBbNh2_2),.clk(gclk));
	jdff dff_B_8hjx9cwO1_2(.din(w_dff_B_ZIXfBbNh2_2),.dout(w_dff_B_8hjx9cwO1_2),.clk(gclk));
	jdff dff_B_SRgwEUGB7_2(.din(w_dff_B_8hjx9cwO1_2),.dout(w_dff_B_SRgwEUGB7_2),.clk(gclk));
	jdff dff_B_0LmqApjW4_2(.din(w_dff_B_SRgwEUGB7_2),.dout(w_dff_B_0LmqApjW4_2),.clk(gclk));
	jdff dff_B_vDp3rU3n0_2(.din(n1610),.dout(w_dff_B_vDp3rU3n0_2),.clk(gclk));
	jdff dff_B_dDHCOc7C7_1(.din(n1607),.dout(w_dff_B_dDHCOc7C7_1),.clk(gclk));
	jdff dff_B_8lzZujin8_0(.din(n1604),.dout(w_dff_B_8lzZujin8_0),.clk(gclk));
	jdff dff_B_alLF9ndC9_0(.din(w_dff_B_8lzZujin8_0),.dout(w_dff_B_alLF9ndC9_0),.clk(gclk));
	jdff dff_B_pubdDgxt8_1(.din(n1597),.dout(w_dff_B_pubdDgxt8_1),.clk(gclk));
	jdff dff_B_aC9HYw690_1(.din(w_dff_B_pubdDgxt8_1),.dout(w_dff_B_aC9HYw690_1),.clk(gclk));
	jdff dff_B_aCGE8svr5_1(.din(w_dff_B_aC9HYw690_1),.dout(w_dff_B_aCGE8svr5_1),.clk(gclk));
	jdff dff_B_KOp4eg1C7_1(.din(w_dff_B_aCGE8svr5_1),.dout(w_dff_B_KOp4eg1C7_1),.clk(gclk));
	jdff dff_B_AhLXTjoJ4_1(.din(w_dff_B_KOp4eg1C7_1),.dout(w_dff_B_AhLXTjoJ4_1),.clk(gclk));
	jdff dff_B_7nAtSZzz0_0(.din(n1602),.dout(w_dff_B_7nAtSZzz0_0),.clk(gclk));
	jdff dff_A_hQattbZ39_0(.dout(w_n558_0[0]),.din(w_dff_A_hQattbZ39_0),.clk(gclk));
	jdff dff_A_xTaIYJsU6_1(.dout(w_n558_0[1]),.din(w_dff_A_xTaIYJsU6_1),.clk(gclk));
	jdff dff_A_4HxMOBzB0_1(.dout(w_dff_A_xTaIYJsU6_1),.din(w_dff_A_4HxMOBzB0_1),.clk(gclk));
	jdff dff_A_oTTWZ4n12_1(.dout(w_dff_A_4HxMOBzB0_1),.din(w_dff_A_oTTWZ4n12_1),.clk(gclk));
	jdff dff_A_fSJa1hQi3_1(.dout(w_dff_A_oTTWZ4n12_1),.din(w_dff_A_fSJa1hQi3_1),.clk(gclk));
	jdff dff_A_Dfo02qTY1_1(.dout(w_dff_A_fSJa1hQi3_1),.din(w_dff_A_Dfo02qTY1_1),.clk(gclk));
	jdff dff_A_wNrVRr4m0_1(.dout(w_dff_A_Dfo02qTY1_1),.din(w_dff_A_wNrVRr4m0_1),.clk(gclk));
	jdff dff_A_HIYgWKut1_1(.dout(w_dff_A_wNrVRr4m0_1),.din(w_dff_A_HIYgWKut1_1),.clk(gclk));
	jdff dff_A_H569RaTp6_1(.dout(w_dff_A_HIYgWKut1_1),.din(w_dff_A_H569RaTp6_1),.clk(gclk));
	jdff dff_A_iC0lMWdM1_1(.dout(w_n1380_0[1]),.din(w_dff_A_iC0lMWdM1_1),.clk(gclk));
	jdff dff_A_OQdcaMSn4_1(.dout(w_dff_A_iC0lMWdM1_1),.din(w_dff_A_OQdcaMSn4_1),.clk(gclk));
	jdff dff_B_3o2Gmpu88_0(.din(n1377),.dout(w_dff_B_3o2Gmpu88_0),.clk(gclk));
	jdff dff_B_U6Y7eEEh5_0(.din(n1594),.dout(w_dff_B_U6Y7eEEh5_0),.clk(gclk));
	jdff dff_B_ykGpgJUh3_0(.din(w_dff_B_U6Y7eEEh5_0),.dout(w_dff_B_ykGpgJUh3_0),.clk(gclk));
	jdff dff_B_H1VZyRNg0_0(.din(w_dff_B_ykGpgJUh3_0),.dout(w_dff_B_H1VZyRNg0_0),.clk(gclk));
	jdff dff_B_DOyrpJvK3_0(.din(n1593),.dout(w_dff_B_DOyrpJvK3_0),.clk(gclk));
	jdff dff_B_Zg1Nctpa2_0(.din(w_dff_B_DOyrpJvK3_0),.dout(w_dff_B_Zg1Nctpa2_0),.clk(gclk));
	jdff dff_B_F3j65Tk89_0(.din(w_dff_B_Zg1Nctpa2_0),.dout(w_dff_B_F3j65Tk89_0),.clk(gclk));
	jdff dff_A_Z1DwoZXy7_2(.dout(w_n1494_0[2]),.din(w_dff_A_Z1DwoZXy7_2),.clk(gclk));
	jdff dff_A_w5hToErj1_2(.dout(w_dff_A_Z1DwoZXy7_2),.din(w_dff_A_w5hToErj1_2),.clk(gclk));
	jdff dff_A_WxIS492Z8_2(.dout(w_dff_A_w5hToErj1_2),.din(w_dff_A_WxIS492Z8_2),.clk(gclk));
	jdff dff_A_KQi5rTxb2_2(.dout(w_dff_A_WxIS492Z8_2),.din(w_dff_A_KQi5rTxb2_2),.clk(gclk));
	jdff dff_A_WR1umVCz7_2(.dout(w_dff_A_KQi5rTxb2_2),.din(w_dff_A_WR1umVCz7_2),.clk(gclk));
	jdff dff_A_1NCt1dSV6_2(.dout(w_dff_A_WR1umVCz7_2),.din(w_dff_A_1NCt1dSV6_2),.clk(gclk));
	jdff dff_A_PRTQMjPF0_2(.dout(w_dff_A_1NCt1dSV6_2),.din(w_dff_A_PRTQMjPF0_2),.clk(gclk));
	jdff dff_A_lC5KzlNe7_2(.dout(w_dff_A_PRTQMjPF0_2),.din(w_dff_A_lC5KzlNe7_2),.clk(gclk));
	jdff dff_A_78EQe3MQ0_1(.dout(w_n524_1[1]),.din(w_dff_A_78EQe3MQ0_1),.clk(gclk));
	jdff dff_A_qBGngdX23_1(.dout(w_dff_A_78EQe3MQ0_1),.din(w_dff_A_qBGngdX23_1),.clk(gclk));
	jdff dff_A_2KyFx0Bm4_2(.dout(w_n524_1[2]),.din(w_dff_A_2KyFx0Bm4_2),.clk(gclk));
	jdff dff_A_8nzIWA842_2(.dout(w_dff_A_2KyFx0Bm4_2),.din(w_dff_A_8nzIWA842_2),.clk(gclk));
	jdff dff_A_ZeZZs0dV3_2(.dout(w_dff_A_8nzIWA842_2),.din(w_dff_A_ZeZZs0dV3_2),.clk(gclk));
	jdff dff_A_UoqdUvOb5_2(.dout(w_dff_A_ZeZZs0dV3_2),.din(w_dff_A_UoqdUvOb5_2),.clk(gclk));
	jdff dff_A_1SsLvTh40_2(.dout(w_dff_A_UoqdUvOb5_2),.din(w_dff_A_1SsLvTh40_2),.clk(gclk));
	jdff dff_A_RreyfHQB5_2(.dout(w_dff_A_1SsLvTh40_2),.din(w_dff_A_RreyfHQB5_2),.clk(gclk));
	jdff dff_A_e4ZBWO9m4_2(.dout(w_dff_A_RreyfHQB5_2),.din(w_dff_A_e4ZBWO9m4_2),.clk(gclk));
	jdff dff_A_Zpd9tXee3_2(.dout(w_dff_A_e4ZBWO9m4_2),.din(w_dff_A_Zpd9tXee3_2),.clk(gclk));
	jdff dff_A_SHEZpuKz4_2(.dout(w_dff_A_Zpd9tXee3_2),.din(w_dff_A_SHEZpuKz4_2),.clk(gclk));
	jdff dff_A_Dy7sPzxc4_2(.dout(w_dff_A_SHEZpuKz4_2),.din(w_dff_A_Dy7sPzxc4_2),.clk(gclk));
	jdff dff_A_FmolRADu2_2(.dout(w_dff_A_Dy7sPzxc4_2),.din(w_dff_A_FmolRADu2_2),.clk(gclk));
	jdff dff_A_tLCwrIOT5_2(.dout(w_dff_A_FmolRADu2_2),.din(w_dff_A_tLCwrIOT5_2),.clk(gclk));
	jdff dff_B_KP4L5NZK5_1(.din(n1588),.dout(w_dff_B_KP4L5NZK5_1),.clk(gclk));
	jdff dff_B_FxcGtuwp1_1(.din(w_dff_B_KP4L5NZK5_1),.dout(w_dff_B_FxcGtuwp1_1),.clk(gclk));
	jdff dff_B_zAykQ3Zi5_1(.din(w_dff_B_FxcGtuwp1_1),.dout(w_dff_B_zAykQ3Zi5_1),.clk(gclk));
	jdff dff_B_0aFNqMVK8_1(.din(w_dff_B_zAykQ3Zi5_1),.dout(w_dff_B_0aFNqMVK8_1),.clk(gclk));
	jdff dff_B_YoGxxV7h9_0(.din(n1590),.dout(w_dff_B_YoGxxV7h9_0),.clk(gclk));
	jdff dff_A_g1ouEMrq9_1(.dout(w_n549_0[1]),.din(w_dff_A_g1ouEMrq9_1),.clk(gclk));
	jdff dff_B_tB8FLDBO1_2(.din(n549),.dout(w_dff_B_tB8FLDBO1_2),.clk(gclk));
	jdff dff_B_Ekj3GVEX2_2(.din(w_dff_B_tB8FLDBO1_2),.dout(w_dff_B_Ekj3GVEX2_2),.clk(gclk));
	jdff dff_A_dCRZ8exy4_1(.dout(w_n556_0[1]),.din(w_dff_A_dCRZ8exy4_1),.clk(gclk));
	jdff dff_A_EAmY7fFJ8_1(.dout(w_dff_A_dCRZ8exy4_1),.din(w_dff_A_EAmY7fFJ8_1),.clk(gclk));
	jdff dff_A_uzqCdOZH0_1(.dout(w_dff_A_EAmY7fFJ8_1),.din(w_dff_A_uzqCdOZH0_1),.clk(gclk));
	jdff dff_A_ix5hyEg16_1(.dout(w_dff_A_uzqCdOZH0_1),.din(w_dff_A_ix5hyEg16_1),.clk(gclk));
	jdff dff_A_I3wjzGvY9_1(.dout(w_dff_A_ix5hyEg16_1),.din(w_dff_A_I3wjzGvY9_1),.clk(gclk));
	jdff dff_A_HVi33uRr1_1(.dout(w_dff_A_I3wjzGvY9_1),.din(w_dff_A_HVi33uRr1_1),.clk(gclk));
	jdff dff_A_a0i57bQe4_1(.dout(w_dff_A_HVi33uRr1_1),.din(w_dff_A_a0i57bQe4_1),.clk(gclk));
	jdff dff_A_QnAjQ93k8_1(.dout(w_dff_A_a0i57bQe4_1),.din(w_dff_A_QnAjQ93k8_1),.clk(gclk));
	jdff dff_A_QX6Uod323_1(.dout(w_dff_A_QnAjQ93k8_1),.din(w_dff_A_QX6Uod323_1),.clk(gclk));
	jdff dff_A_L5XegHHS8_1(.dout(w_n554_0[1]),.din(w_dff_A_L5XegHHS8_1),.clk(gclk));
	jdff dff_A_QKQ2amWD8_1(.dout(w_dff_A_L5XegHHS8_1),.din(w_dff_A_QKQ2amWD8_1),.clk(gclk));
	jdff dff_A_tJfaK4Ju3_1(.dout(w_dff_A_QKQ2amWD8_1),.din(w_dff_A_tJfaK4Ju3_1),.clk(gclk));
	jdff dff_A_FTOhM2mj4_1(.dout(w_dff_A_tJfaK4Ju3_1),.din(w_dff_A_FTOhM2mj4_1),.clk(gclk));
	jdff dff_A_pdOZCc329_1(.dout(w_dff_A_FTOhM2mj4_1),.din(w_dff_A_pdOZCc329_1),.clk(gclk));
	jdff dff_A_Z5Ds0Uve1_1(.dout(w_dff_A_pdOZCc329_1),.din(w_dff_A_Z5Ds0Uve1_1),.clk(gclk));
	jdff dff_A_3c8LB2TV3_1(.dout(w_dff_A_Z5Ds0Uve1_1),.din(w_dff_A_3c8LB2TV3_1),.clk(gclk));
	jdff dff_A_k3g2QycC6_1(.dout(w_dff_A_3c8LB2TV3_1),.din(w_dff_A_k3g2QycC6_1),.clk(gclk));
	jdff dff_A_9782IDLv3_1(.dout(w_dff_A_k3g2QycC6_1),.din(w_dff_A_9782IDLv3_1),.clk(gclk));
	jdff dff_A_vqJTOoUp7_1(.dout(w_dff_A_9782IDLv3_1),.din(w_dff_A_vqJTOoUp7_1),.clk(gclk));
	jdff dff_A_95FZA3Zm5_1(.dout(w_dff_A_vqJTOoUp7_1),.din(w_dff_A_95FZA3Zm5_1),.clk(gclk));
	jdff dff_B_I0QzRyjh5_1(.din(n526),.dout(w_dff_B_I0QzRyjh5_1),.clk(gclk));
	jdff dff_B_F8ISny507_0(.din(G35),.dout(w_dff_B_F8ISny507_0),.clk(gclk));
	jdff dff_A_sTiYDLQz0_1(.dout(w_n525_0[1]),.din(w_dff_A_sTiYDLQz0_1),.clk(gclk));
	jdff dff_A_kwZnzYGS7_1(.dout(w_dff_A_sTiYDLQz0_1),.din(w_dff_A_kwZnzYGS7_1),.clk(gclk));
	jdff dff_A_lRoOg2Uc0_2(.dout(w_n525_0[2]),.din(w_dff_A_lRoOg2Uc0_2),.clk(gclk));
	jdff dff_A_fe8fo5r10_2(.dout(w_dff_A_lRoOg2Uc0_2),.din(w_dff_A_fe8fo5r10_2),.clk(gclk));
	jdff dff_A_fwJ1w6eR5_1(.dout(w_G4420_0[1]),.din(w_dff_A_fwJ1w6eR5_1),.clk(gclk));
	jdff dff_A_WhG7ffGB8_1(.dout(w_dff_A_fwJ1w6eR5_1),.din(w_dff_A_WhG7ffGB8_1),.clk(gclk));
	jdff dff_A_sBxsNhxh5_1(.dout(w_dff_A_WhG7ffGB8_1),.din(w_dff_A_sBxsNhxh5_1),.clk(gclk));
	jdff dff_A_YC2tkVlL3_1(.dout(w_dff_A_sBxsNhxh5_1),.din(w_dff_A_YC2tkVlL3_1),.clk(gclk));
	jdff dff_A_IOiWJg5o5_2(.dout(w_n524_0[2]),.din(w_dff_A_IOiWJg5o5_2),.clk(gclk));
	jdff dff_A_8JjfnqII7_2(.dout(w_dff_A_IOiWJg5o5_2),.din(w_dff_A_8JjfnqII7_2),.clk(gclk));
	jdff dff_A_8dfze55T3_0(.dout(w_n553_0[0]),.din(w_dff_A_8dfze55T3_0),.clk(gclk));
	jdff dff_A_vv5S50hW9_0(.dout(w_dff_A_8dfze55T3_0),.din(w_dff_A_vv5S50hW9_0),.clk(gclk));
	jdff dff_B_B10ySFGf6_2(.din(n553),.dout(w_dff_B_B10ySFGf6_2),.clk(gclk));
	jdff dff_B_97p8fcFJ9_1(.din(n521),.dout(w_dff_B_97p8fcFJ9_1),.clk(gclk));
	jdff dff_B_yFaDUAMU1_0(.din(G32),.dout(w_dff_B_yFaDUAMU1_0),.clk(gclk));
	jdff dff_A_Xd8iHAHD4_1(.dout(w_n520_0[1]),.din(w_dff_A_Xd8iHAHD4_1),.clk(gclk));
	jdff dff_A_tEZvOvdz5_1(.dout(w_dff_A_Xd8iHAHD4_1),.din(w_dff_A_tEZvOvdz5_1),.clk(gclk));
	jdff dff_A_lgvxJug60_2(.dout(w_n520_0[2]),.din(w_dff_A_lgvxJug60_2),.clk(gclk));
	jdff dff_A_0y5Ha0Y56_2(.dout(w_dff_A_lgvxJug60_2),.din(w_dff_A_0y5Ha0Y56_2),.clk(gclk));
	jdff dff_A_RtiSY4fQ2_0(.dout(w_n552_0[0]),.din(w_dff_A_RtiSY4fQ2_0),.clk(gclk));
	jdff dff_A_fdX7CWqp1_0(.dout(w_dff_A_RtiSY4fQ2_0),.din(w_dff_A_fdX7CWqp1_0),.clk(gclk));
	jdff dff_A_zLmGukhK8_0(.dout(w_dff_A_fdX7CWqp1_0),.din(w_dff_A_zLmGukhK8_0),.clk(gclk));
	jdff dff_A_bqpQrA9F8_0(.dout(w_dff_A_zLmGukhK8_0),.din(w_dff_A_bqpQrA9F8_0),.clk(gclk));
	jdff dff_A_JWLxaX346_0(.dout(w_dff_A_bqpQrA9F8_0),.din(w_dff_A_JWLxaX346_0),.clk(gclk));
	jdff dff_A_KmUpYuOj5_0(.dout(w_dff_A_JWLxaX346_0),.din(w_dff_A_KmUpYuOj5_0),.clk(gclk));
	jdff dff_A_GUN2MG2N4_0(.dout(w_dff_A_KmUpYuOj5_0),.din(w_dff_A_GUN2MG2N4_0),.clk(gclk));
	jdff dff_A_EilkRqAs1_0(.dout(w_dff_A_GUN2MG2N4_0),.din(w_dff_A_EilkRqAs1_0),.clk(gclk));
	jdff dff_A_2eLJHofx6_0(.dout(w_dff_A_EilkRqAs1_0),.din(w_dff_A_2eLJHofx6_0),.clk(gclk));
	jdff dff_A_9xUOQxEp4_0(.dout(w_n551_0[0]),.din(w_dff_A_9xUOQxEp4_0),.clk(gclk));
	jdff dff_A_eYpMDjrG1_0(.dout(w_dff_A_9xUOQxEp4_0),.din(w_dff_A_eYpMDjrG1_0),.clk(gclk));
	jdff dff_A_Kx8Fz1th4_0(.dout(w_dff_A_eYpMDjrG1_0),.din(w_dff_A_Kx8Fz1th4_0),.clk(gclk));
	jdff dff_A_I8x6vdEz0_1(.dout(w_n535_0[1]),.din(w_dff_A_I8x6vdEz0_1),.clk(gclk));
	jdff dff_B_z56kjaHO9_1(.din(n532),.dout(w_dff_B_z56kjaHO9_1),.clk(gclk));
	jdff dff_B_Wt9cimE64_0(.din(G66),.dout(w_dff_B_Wt9cimE64_0),.clk(gclk));
	jdff dff_A_qqZdnrpo0_1(.dout(w_n531_0[1]),.din(w_dff_A_qqZdnrpo0_1),.clk(gclk));
	jdff dff_A_YqWCkFnU9_1(.dout(w_dff_A_qqZdnrpo0_1),.din(w_dff_A_YqWCkFnU9_1),.clk(gclk));
	jdff dff_A_2TAlZ9ka6_2(.dout(w_n531_0[2]),.din(w_dff_A_2TAlZ9ka6_2),.clk(gclk));
	jdff dff_A_w0Fgt6lT0_2(.dout(w_dff_A_2TAlZ9ka6_2),.din(w_dff_A_w0Fgt6lT0_2),.clk(gclk));
	jdff dff_A_ex8w77Gc8_1(.dout(w_G4437_0[1]),.din(w_dff_A_ex8w77Gc8_1),.clk(gclk));
	jdff dff_A_HGDNZH0E4_1(.dout(w_dff_A_ex8w77Gc8_1),.din(w_dff_A_HGDNZH0E4_1),.clk(gclk));
	jdff dff_A_LU3hBHnd8_1(.dout(w_dff_A_HGDNZH0E4_1),.din(w_dff_A_LU3hBHnd8_1),.clk(gclk));
	jdff dff_A_qntVsXhl5_1(.dout(w_dff_A_LU3hBHnd8_1),.din(w_dff_A_qntVsXhl5_1),.clk(gclk));
	jdff dff_A_5SfUobBg9_1(.dout(w_n518_0[1]),.din(w_dff_A_5SfUobBg9_1),.clk(gclk));
	jdff dff_B_wYhbOksX3_1(.din(n498),.dout(w_dff_B_wYhbOksX3_1),.clk(gclk));
	jdff dff_B_TqirbmY73_1(.din(w_dff_B_wYhbOksX3_1),.dout(w_dff_B_TqirbmY73_1),.clk(gclk));
	jdff dff_B_tteSSYUL1_1(.din(w_dff_B_TqirbmY73_1),.dout(w_dff_B_tteSSYUL1_1),.clk(gclk));
	jdff dff_B_z3PaCVmp0_1(.din(w_dff_B_tteSSYUL1_1),.dout(w_dff_B_z3PaCVmp0_1),.clk(gclk));
	jdff dff_B_Ch26jVpJ5_1(.din(w_dff_B_z3PaCVmp0_1),.dout(w_dff_B_Ch26jVpJ5_1),.clk(gclk));
	jdff dff_B_2yFhqfr89_1(.din(w_dff_B_Ch26jVpJ5_1),.dout(w_dff_B_2yFhqfr89_1),.clk(gclk));
	jdff dff_B_3ABd8Tn76_1(.din(n500),.dout(w_dff_B_3ABd8Tn76_1),.clk(gclk));
	jdff dff_B_ShIWzOkd9_1(.din(w_dff_B_3ABd8Tn76_1),.dout(w_dff_B_ShIWzOkd9_1),.clk(gclk));
	jdff dff_B_m2xCqVHy2_1(.din(w_dff_B_ShIWzOkd9_1),.dout(w_dff_B_m2xCqVHy2_1),.clk(gclk));
	jdff dff_B_gl1CDZkN4_1(.din(w_dff_B_m2xCqVHy2_1),.dout(w_dff_B_gl1CDZkN4_1),.clk(gclk));
	jdff dff_B_SZj7H64q1_1(.din(w_dff_B_gl1CDZkN4_1),.dout(w_dff_B_SZj7H64q1_1),.clk(gclk));
	jdff dff_A_yPmzw50R3_1(.dout(w_n516_0[1]),.din(w_dff_A_yPmzw50R3_1),.clk(gclk));
	jdff dff_A_S2mrRg5I6_1(.dout(w_dff_A_yPmzw50R3_1),.din(w_dff_A_S2mrRg5I6_1),.clk(gclk));
	jdff dff_A_uiWlQ2a99_1(.dout(w_dff_A_S2mrRg5I6_1),.din(w_dff_A_uiWlQ2a99_1),.clk(gclk));
	jdff dff_A_Pqka6t3i7_1(.dout(w_dff_A_uiWlQ2a99_1),.din(w_dff_A_Pqka6t3i7_1),.clk(gclk));
	jdff dff_A_W7mZd8nP7_1(.dout(w_dff_A_Pqka6t3i7_1),.din(w_dff_A_W7mZd8nP7_1),.clk(gclk));
	jdff dff_B_kkbqWu3W4_1(.din(n504),.dout(w_dff_B_kkbqWu3W4_1),.clk(gclk));
	jdff dff_B_1NJpbKnL3_1(.din(w_dff_B_kkbqWu3W4_1),.dout(w_dff_B_1NJpbKnL3_1),.clk(gclk));
	jdff dff_B_fczQLOE96_1(.din(w_dff_B_1NJpbKnL3_1),.dout(w_dff_B_fczQLOE96_1),.clk(gclk));
	jdff dff_A_3O4irouc6_1(.dout(w_n514_0[1]),.din(w_dff_A_3O4irouc6_1),.clk(gclk));
	jdff dff_A_i8KOMWV04_1(.dout(w_dff_A_3O4irouc6_1),.din(w_dff_A_i8KOMWV04_1),.clk(gclk));
	jdff dff_A_R0nhVeYO9_1(.dout(w_dff_A_i8KOMWV04_1),.din(w_dff_A_R0nhVeYO9_1),.clk(gclk));
	jdff dff_A_EtzBKUza9_1(.dout(w_dff_A_R0nhVeYO9_1),.din(w_dff_A_EtzBKUza9_1),.clk(gclk));
	jdff dff_A_2EV3RvmL5_1(.dout(w_dff_A_EtzBKUza9_1),.din(w_dff_A_2EV3RvmL5_1),.clk(gclk));
	jdff dff_A_HM97nvu99_1(.dout(w_dff_A_2EV3RvmL5_1),.din(w_dff_A_HM97nvu99_1),.clk(gclk));
	jdff dff_A_FTpluSiU1_0(.dout(w_n512_0[0]),.din(w_dff_A_FTpluSiU1_0),.clk(gclk));
	jdff dff_A_flRhmxis9_0(.dout(w_n510_0[0]),.din(w_dff_A_flRhmxis9_0),.clk(gclk));
	jdff dff_A_sN80vvk98_0(.dout(w_n509_0[0]),.din(w_dff_A_sN80vvk98_0),.clk(gclk));
	jdff dff_A_TWgdoSAu6_0(.dout(w_dff_A_sN80vvk98_0),.din(w_dff_A_TWgdoSAu6_0),.clk(gclk));
	jdff dff_A_qvGD8QD72_2(.dout(w_n507_0[2]),.din(w_dff_A_qvGD8QD72_2),.clk(gclk));
	jdff dff_A_4kQZVwXf8_2(.dout(w_dff_A_qvGD8QD72_2),.din(w_dff_A_4kQZVwXf8_2),.clk(gclk));
	jdff dff_A_857j7mv22_2(.dout(w_dff_A_4kQZVwXf8_2),.din(w_dff_A_857j7mv22_2),.clk(gclk));
	jdff dff_A_SrxoqYpU5_2(.dout(w_dff_A_857j7mv22_2),.din(w_dff_A_SrxoqYpU5_2),.clk(gclk));
	jdff dff_A_yB9qZISK9_1(.dout(w_n505_0[1]),.din(w_dff_A_yB9qZISK9_1),.clk(gclk));
	jdff dff_B_XhCpM7G88_2(.din(n505),.dout(w_dff_B_XhCpM7G88_2),.clk(gclk));
	jdff dff_A_JqcRgyAl8_0(.dout(w_n503_0[0]),.din(w_dff_A_JqcRgyAl8_0),.clk(gclk));
	jdff dff_A_ia4ZqPFa5_0(.dout(w_n502_0[0]),.din(w_dff_A_ia4ZqPFa5_0),.clk(gclk));
	jdff dff_B_Xx4hh2Hp1_2(.din(n502),.dout(w_dff_B_Xx4hh2Hp1_2),.clk(gclk));
	jdff dff_B_Ij49NSmw6_2(.din(w_dff_B_Xx4hh2Hp1_2),.dout(w_dff_B_Ij49NSmw6_2),.clk(gclk));
	jdff dff_B_3nfjAfVU4_2(.din(w_dff_B_Ij49NSmw6_2),.dout(w_dff_B_3nfjAfVU4_2),.clk(gclk));
	jdff dff_B_EaTX5xwa0_2(.din(w_dff_B_3nfjAfVU4_2),.dout(w_dff_B_EaTX5xwa0_2),.clk(gclk));
	jdff dff_B_Y348e3jW9_0(.din(n495),.dout(w_dff_B_Y348e3jW9_0),.clk(gclk));
	jdff dff_B_WV33yBBi5_0(.din(w_dff_B_Y348e3jW9_0),.dout(w_dff_B_WV33yBBi5_0),.clk(gclk));
	jdff dff_B_kxkwTheF8_0(.din(w_dff_B_WV33yBBi5_0),.dout(w_dff_B_kxkwTheF8_0),.clk(gclk));
	jdff dff_A_6xDLqePH0_0(.dout(w_n494_0[0]),.din(w_dff_A_6xDLqePH0_0),.clk(gclk));
	jdff dff_A_jFlnITkq0_0(.dout(w_dff_A_6xDLqePH0_0),.din(w_dff_A_jFlnITkq0_0),.clk(gclk));
	jdff dff_A_yaaScwek6_0(.dout(w_dff_A_jFlnITkq0_0),.din(w_dff_A_yaaScwek6_0),.clk(gclk));
	jdff dff_A_7mpuZtjD6_0(.dout(w_dff_A_yaaScwek6_0),.din(w_dff_A_7mpuZtjD6_0),.clk(gclk));
	jdff dff_A_YgyQP05y7_0(.dout(w_n493_0[0]),.din(w_dff_A_YgyQP05y7_0),.clk(gclk));
	jdff dff_A_G8MzJ7MA5_0(.dout(w_dff_A_YgyQP05y7_0),.din(w_dff_A_G8MzJ7MA5_0),.clk(gclk));
	jdff dff_A_8roTyld63_0(.dout(w_dff_A_G8MzJ7MA5_0),.din(w_dff_A_8roTyld63_0),.clk(gclk));
	jdff dff_A_Hp7boeQl5_0(.dout(w_dff_A_8roTyld63_0),.din(w_dff_A_Hp7boeQl5_0),.clk(gclk));
	jdff dff_A_khTztlvm4_0(.dout(w_n480_1[0]),.din(w_dff_A_khTztlvm4_0),.clk(gclk));
	jdff dff_A_NQl7Rqat5_0(.dout(w_dff_A_khTztlvm4_0),.din(w_dff_A_NQl7Rqat5_0),.clk(gclk));
	jdff dff_A_qntXB8sd5_0(.dout(w_dff_A_NQl7Rqat5_0),.din(w_dff_A_qntXB8sd5_0),.clk(gclk));
	jdff dff_A_KIFSArAG1_0(.dout(w_dff_A_qntXB8sd5_0),.din(w_dff_A_KIFSArAG1_0),.clk(gclk));
	jdff dff_A_uIbQgI7W1_0(.dout(w_dff_A_KIFSArAG1_0),.din(w_dff_A_uIbQgI7W1_0),.clk(gclk));
	jdff dff_A_l8ZtE8Sn4_0(.dout(w_dff_A_uIbQgI7W1_0),.din(w_dff_A_l8ZtE8Sn4_0),.clk(gclk));
	jdff dff_A_VVnNbHzg0_0(.dout(w_dff_A_l8ZtE8Sn4_0),.din(w_dff_A_VVnNbHzg0_0),.clk(gclk));
	jdff dff_A_keEUnmVx0_1(.dout(w_n480_0[1]),.din(w_dff_A_keEUnmVx0_1),.clk(gclk));
	jdff dff_A_oUm0klVa5_1(.dout(w_dff_A_keEUnmVx0_1),.din(w_dff_A_oUm0klVa5_1),.clk(gclk));
	jdff dff_A_rFFq4SYb4_1(.dout(w_dff_A_oUm0klVa5_1),.din(w_dff_A_rFFq4SYb4_1),.clk(gclk));
	jdff dff_A_CYHEFmLD2_2(.dout(w_n480_0[2]),.din(w_dff_A_CYHEFmLD2_2),.clk(gclk));
	jdff dff_A_jw7BCaO68_2(.dout(w_dff_A_CYHEFmLD2_2),.din(w_dff_A_jw7BCaO68_2),.clk(gclk));
	jdff dff_A_IywU0Cun9_2(.dout(w_dff_A_jw7BCaO68_2),.din(w_dff_A_IywU0Cun9_2),.clk(gclk));
	jdff dff_A_TE6sAppO1_2(.dout(w_dff_A_IywU0Cun9_2),.din(w_dff_A_TE6sAppO1_2),.clk(gclk));
	jdff dff_A_4cSmD5gy5_2(.dout(w_dff_A_TE6sAppO1_2),.din(w_dff_A_4cSmD5gy5_2),.clk(gclk));
	jdff dff_A_trKnJhZs1_2(.dout(w_dff_A_4cSmD5gy5_2),.din(w_dff_A_trKnJhZs1_2),.clk(gclk));
	jdff dff_A_nGLOxQN57_2(.dout(w_dff_A_trKnJhZs1_2),.din(w_dff_A_nGLOxQN57_2),.clk(gclk));
	jdff dff_B_m5PZQapt5_1(.din(n476),.dout(w_dff_B_m5PZQapt5_1),.clk(gclk));
	jdff dff_B_COBhojxa7_0(.din(G118),.dout(w_dff_B_COBhojxa7_0),.clk(gclk));
	jdff dff_A_fPlEzJqL3_0(.dout(w_G4394_0[0]),.din(w_dff_A_fPlEzJqL3_0),.clk(gclk));
	jdff dff_A_AbIZFLkS2_0(.dout(w_dff_A_fPlEzJqL3_0),.din(w_dff_A_AbIZFLkS2_0),.clk(gclk));
	jdff dff_A_x7xqnppb8_0(.dout(w_dff_A_AbIZFLkS2_0),.din(w_dff_A_x7xqnppb8_0),.clk(gclk));
	jdff dff_A_PS3VzGrE0_0(.dout(w_dff_A_x7xqnppb8_0),.din(w_dff_A_PS3VzGrE0_0),.clk(gclk));
	jdff dff_A_yTBxxcit6_1(.dout(w_n475_1[1]),.din(w_dff_A_yTBxxcit6_1),.clk(gclk));
	jdff dff_A_xgz0nFoM5_1(.dout(w_n475_0[1]),.din(w_dff_A_xgz0nFoM5_1),.clk(gclk));
	jdff dff_A_LMRh3XSK2_2(.dout(w_n475_0[2]),.din(w_dff_A_LMRh3XSK2_2),.clk(gclk));
	jdff dff_A_4E29kbFd3_2(.dout(w_dff_A_LMRh3XSK2_2),.din(w_dff_A_4E29kbFd3_2),.clk(gclk));
	jdff dff_A_Z7XSjzxx0_2(.dout(w_dff_A_4E29kbFd3_2),.din(w_dff_A_Z7XSjzxx0_2),.clk(gclk));
	jdff dff_A_3wCQvhAm0_2(.dout(w_dff_A_Z7XSjzxx0_2),.din(w_dff_A_3wCQvhAm0_2),.clk(gclk));
	jdff dff_A_PhRHS0Mz5_2(.dout(w_dff_A_3wCQvhAm0_2),.din(w_dff_A_PhRHS0Mz5_2),.clk(gclk));
	jdff dff_A_PlYYp1HR2_2(.dout(w_dff_A_PhRHS0Mz5_2),.din(w_dff_A_PlYYp1HR2_2),.clk(gclk));
	jdff dff_A_b2HDrILW8_2(.dout(w_dff_A_PlYYp1HR2_2),.din(w_dff_A_b2HDrILW8_2),.clk(gclk));
	jdff dff_A_x5GUgam20_2(.dout(w_dff_A_b2HDrILW8_2),.din(w_dff_A_x5GUgam20_2),.clk(gclk));
	jdff dff_A_eu9gHB4t5_2(.dout(w_dff_A_x5GUgam20_2),.din(w_dff_A_eu9gHB4t5_2),.clk(gclk));
	jdff dff_A_knNpTlxh2_2(.dout(w_dff_A_eu9gHB4t5_2),.din(w_dff_A_knNpTlxh2_2),.clk(gclk));
	jdff dff_B_ZBbtVsur2_1(.din(n472),.dout(w_dff_B_ZBbtVsur2_1),.clk(gclk));
	jdff dff_B_LQ7pEVUH6_0(.din(G97),.dout(w_dff_B_LQ7pEVUH6_0),.clk(gclk));
	jdff dff_B_yjs8ziQ73_3(.din(n471),.dout(w_dff_B_yjs8ziQ73_3),.clk(gclk));
	jdff dff_B_7v6UQacD2_3(.din(w_dff_B_yjs8ziQ73_3),.dout(w_dff_B_7v6UQacD2_3),.clk(gclk));
	jdff dff_A_cTchlEhg0_0(.dout(w_n470_0[0]),.din(w_dff_A_cTchlEhg0_0),.clk(gclk));
	jdff dff_A_gfkGvZBc3_0(.dout(w_dff_A_cTchlEhg0_0),.din(w_dff_A_gfkGvZBc3_0),.clk(gclk));
	jdff dff_A_r2bCk0VM8_0(.dout(w_dff_A_gfkGvZBc3_0),.din(w_dff_A_r2bCk0VM8_0),.clk(gclk));
	jdff dff_A_RV0X8r4x8_0(.dout(w_dff_A_r2bCk0VM8_0),.din(w_dff_A_RV0X8r4x8_0),.clk(gclk));
	jdff dff_A_TxZ6rDGb9_2(.dout(w_n470_0[2]),.din(w_dff_A_TxZ6rDGb9_2),.clk(gclk));
	jdff dff_A_6jZbSEWD6_2(.dout(w_dff_A_TxZ6rDGb9_2),.din(w_dff_A_6jZbSEWD6_2),.clk(gclk));
	jdff dff_A_9cGYOAGn6_2(.dout(w_dff_A_6jZbSEWD6_2),.din(w_dff_A_9cGYOAGn6_2),.clk(gclk));
	jdff dff_B_zliV9cO33_1(.din(n467),.dout(w_dff_B_zliV9cO33_1),.clk(gclk));
	jdff dff_B_fMrwYs659_0(.din(G47),.dout(w_dff_B_fMrwYs659_0),.clk(gclk));
	jdff dff_B_ZA2YkqfJ9_2(.din(n466),.dout(w_dff_B_ZA2YkqfJ9_2),.clk(gclk));
	jdff dff_B_Sq1hXx1k3_2(.din(w_dff_B_ZA2YkqfJ9_2),.dout(w_dff_B_Sq1hXx1k3_2),.clk(gclk));
	jdff dff_A_I0Mqpxop7_0(.dout(w_G4415_1[0]),.din(w_dff_A_I0Mqpxop7_0),.clk(gclk));
	jdff dff_A_FaoZZSWF2_0(.dout(w_dff_A_I0Mqpxop7_0),.din(w_dff_A_FaoZZSWF2_0),.clk(gclk));
	jdff dff_A_bn8IRPe41_0(.dout(w_dff_A_FaoZZSWF2_0),.din(w_dff_A_bn8IRPe41_0),.clk(gclk));
	jdff dff_A_X1Xekpxs6_0(.dout(w_dff_A_bn8IRPe41_0),.din(w_dff_A_X1Xekpxs6_0),.clk(gclk));
	jdff dff_A_odcbesw53_0(.dout(w_n465_0[0]),.din(w_dff_A_odcbesw53_0),.clk(gclk));
	jdff dff_A_0gJh73xG8_0(.dout(w_dff_A_odcbesw53_0),.din(w_dff_A_0gJh73xG8_0),.clk(gclk));
	jdff dff_A_8cDr3tWy7_0(.dout(w_dff_A_0gJh73xG8_0),.din(w_dff_A_8cDr3tWy7_0),.clk(gclk));
	jdff dff_A_WazBq6Ez1_0(.dout(w_dff_A_8cDr3tWy7_0),.din(w_dff_A_WazBq6Ez1_0),.clk(gclk));
	jdff dff_A_rX7nEYGu3_1(.dout(w_n464_0[1]),.din(w_dff_A_rX7nEYGu3_1),.clk(gclk));
	jdff dff_A_V7MBk9M43_1(.dout(w_n452_0[1]),.din(w_dff_A_V7MBk9M43_1),.clk(gclk));
	jdff dff_A_jXb34jZa4_1(.dout(w_dff_A_V7MBk9M43_1),.din(w_dff_A_jXb34jZa4_1),.clk(gclk));
	jdff dff_A_nJ6YFvbH5_0(.dout(w_n446_1[0]),.din(w_dff_A_nJ6YFvbH5_0),.clk(gclk));
	jdff dff_A_ViGJP46Z6_0(.dout(w_dff_A_nJ6YFvbH5_0),.din(w_dff_A_ViGJP46Z6_0),.clk(gclk));
	jdff dff_A_BCgUxyrU9_0(.dout(w_dff_A_ViGJP46Z6_0),.din(w_dff_A_BCgUxyrU9_0),.clk(gclk));
	jdff dff_A_44Lhg1Uy2_0(.dout(w_dff_A_BCgUxyrU9_0),.din(w_dff_A_44Lhg1Uy2_0),.clk(gclk));
	jdff dff_A_hoGJtfG63_0(.dout(w_dff_A_44Lhg1Uy2_0),.din(w_dff_A_hoGJtfG63_0),.clk(gclk));
	jdff dff_A_8rzJjEAT2_0(.dout(w_dff_A_hoGJtfG63_0),.din(w_dff_A_8rzJjEAT2_0),.clk(gclk));
	jdff dff_A_jup20k5Y2_0(.dout(w_dff_A_8rzJjEAT2_0),.din(w_dff_A_jup20k5Y2_0),.clk(gclk));
	jdff dff_A_noX17VGj4_0(.dout(w_n437_0[0]),.din(w_dff_A_noX17VGj4_0),.clk(gclk));
	jdff dff_A_YYOCxAdK6_0(.dout(w_dff_A_noX17VGj4_0),.din(w_dff_A_YYOCxAdK6_0),.clk(gclk));
	jdff dff_A_TLkKiRen5_0(.dout(w_dff_A_YYOCxAdK6_0),.din(w_dff_A_TLkKiRen5_0),.clk(gclk));
	jdff dff_B_weC9zydJ4_2(.din(n437),.dout(w_dff_B_weC9zydJ4_2),.clk(gclk));
	jdff dff_B_3rT1SpkR9_2(.din(w_dff_B_weC9zydJ4_2),.dout(w_dff_B_3rT1SpkR9_2),.clk(gclk));
	jdff dff_A_PYzgD2YE7_0(.dout(w_n436_0[0]),.din(w_dff_A_PYzgD2YE7_0),.clk(gclk));
	jdff dff_A_ptpoevLv0_0(.dout(w_dff_A_PYzgD2YE7_0),.din(w_dff_A_ptpoevLv0_0),.clk(gclk));
	jdff dff_A_sBlCRa8G5_0(.dout(w_dff_A_ptpoevLv0_0),.din(w_dff_A_sBlCRa8G5_0),.clk(gclk));
	jdff dff_A_koUiVA1f6_0(.dout(w_dff_A_sBlCRa8G5_0),.din(w_dff_A_koUiVA1f6_0),.clk(gclk));
	jdff dff_A_G2xvfzQQ1_0(.dout(w_dff_A_koUiVA1f6_0),.din(w_dff_A_G2xvfzQQ1_0),.clk(gclk));
	jdff dff_A_lgiSVfCS8_0(.dout(w_dff_A_G2xvfzQQ1_0),.din(w_dff_A_lgiSVfCS8_0),.clk(gclk));
	jdff dff_A_sA0c8zSZ7_1(.dout(w_n430_0[1]),.din(w_dff_A_sA0c8zSZ7_1),.clk(gclk));
	jdff dff_A_QIQb9Krg9_1(.dout(w_dff_A_sA0c8zSZ7_1),.din(w_dff_A_QIQb9Krg9_1),.clk(gclk));
	jdff dff_A_4UNmYwgZ2_1(.dout(w_n491_0[1]),.din(w_dff_A_4UNmYwgZ2_1),.clk(gclk));
	jdff dff_B_esNCd9Ls0_1(.din(n487),.dout(w_dff_B_esNCd9Ls0_1),.clk(gclk));
	jdff dff_B_rIPQjVRj5_0(.din(G94),.dout(w_dff_B_rIPQjVRj5_0),.clk(gclk));
	jdff dff_A_f45I65Ob2_0(.dout(w_G4405_0[0]),.din(w_dff_A_f45I65Ob2_0),.clk(gclk));
	jdff dff_A_jtVdBGyi4_0(.dout(w_dff_A_f45I65Ob2_0),.din(w_dff_A_jtVdBGyi4_0),.clk(gclk));
	jdff dff_A_TvmN6IC27_0(.dout(w_dff_A_jtVdBGyi4_0),.din(w_dff_A_TvmN6IC27_0),.clk(gclk));
	jdff dff_A_Q5yWBHKi1_0(.dout(w_dff_A_TvmN6IC27_0),.din(w_dff_A_Q5yWBHKi1_0),.clk(gclk));
	jdff dff_A_pd39079P7_0(.dout(w_n486_0[0]),.din(w_dff_A_pd39079P7_0),.clk(gclk));
	jdff dff_A_a1ePKEFb4_2(.dout(w_n486_0[2]),.din(w_dff_A_a1ePKEFb4_2),.clk(gclk));
	jdff dff_B_HiEtNCOm9_1(.din(n483),.dout(w_dff_B_HiEtNCOm9_1),.clk(gclk));
	jdff dff_B_Dw4rdbuH0_0(.din(G121),.dout(w_dff_B_Dw4rdbuH0_0),.clk(gclk));
	jdff dff_B_VTW1elSc5_2(.din(n482),.dout(w_dff_B_VTW1elSc5_2),.clk(gclk));
	jdff dff_B_jCrKePCp9_2(.din(w_dff_B_VTW1elSc5_2),.dout(w_dff_B_jCrKePCp9_2),.clk(gclk));
	jdff dff_A_RjZ9GCLL4_0(.dout(w_G4410_1[0]),.din(w_dff_A_RjZ9GCLL4_0),.clk(gclk));
	jdff dff_A_8JVjjYZ15_0(.dout(w_dff_A_RjZ9GCLL4_0),.din(w_dff_A_8JVjjYZ15_0),.clk(gclk));
	jdff dff_A_kxamI6kf1_0(.dout(w_dff_A_8JVjjYZ15_0),.din(w_dff_A_kxamI6kf1_0),.clk(gclk));
	jdff dff_A_r5O3ypv00_0(.dout(w_dff_A_kxamI6kf1_0),.din(w_dff_A_r5O3ypv00_0),.clk(gclk));
	jdff dff_A_WSw6kBLS3_0(.dout(w_n540_0[0]),.din(w_dff_A_WSw6kBLS3_0),.clk(gclk));
	jdff dff_A_8WeyrEFP5_0(.dout(w_dff_A_WSw6kBLS3_0),.din(w_dff_A_8WeyrEFP5_0),.clk(gclk));
	jdff dff_A_MJ2MGH4C0_1(.dout(w_n540_0[1]),.din(w_dff_A_MJ2MGH4C0_1),.clk(gclk));
	jdff dff_A_O0D74pKg7_1(.dout(w_dff_A_MJ2MGH4C0_1),.din(w_dff_A_O0D74pKg7_1),.clk(gclk));
	jdff dff_A_XXzyaZCe2_1(.dout(w_dff_A_O0D74pKg7_1),.din(w_dff_A_XXzyaZCe2_1),.clk(gclk));
	jdff dff_A_WF0JWylQ5_1(.dout(w_dff_A_XXzyaZCe2_1),.din(w_dff_A_WF0JWylQ5_1),.clk(gclk));
	jdff dff_A_CSxwEZoC8_1(.dout(w_dff_A_WF0JWylQ5_1),.din(w_dff_A_CSxwEZoC8_1),.clk(gclk));
	jdff dff_A_5v8rNG9A4_1(.dout(w_dff_A_CSxwEZoC8_1),.din(w_dff_A_5v8rNG9A4_1),.clk(gclk));
	jdff dff_A_TBklSHzn0_1(.dout(w_dff_A_5v8rNG9A4_1),.din(w_dff_A_TBklSHzn0_1),.clk(gclk));
	jdff dff_A_VW0sKbXd3_1(.dout(w_dff_A_TBklSHzn0_1),.din(w_dff_A_VW0sKbXd3_1),.clk(gclk));
	jdff dff_A_F1DFpK1S7_1(.dout(w_dff_A_VW0sKbXd3_1),.din(w_dff_A_F1DFpK1S7_1),.clk(gclk));
	jdff dff_A_Br6k1EEH0_1(.dout(w_dff_A_F1DFpK1S7_1),.din(w_dff_A_Br6k1EEH0_1),.clk(gclk));
	jdff dff_A_GVT8uyKf9_1(.dout(w_dff_A_Br6k1EEH0_1),.din(w_dff_A_GVT8uyKf9_1),.clk(gclk));
	jdff dff_A_izyj3GnA6_1(.dout(w_dff_A_GVT8uyKf9_1),.din(w_dff_A_izyj3GnA6_1),.clk(gclk));
	jdff dff_B_dHFxbENz8_1(.din(n537),.dout(w_dff_B_dHFxbENz8_1),.clk(gclk));
	jdff dff_B_VzS5hBIf6_0(.din(G50),.dout(w_dff_B_VzS5hBIf6_0),.clk(gclk));
	jdff dff_B_x67f0iET4_2(.din(n536),.dout(w_dff_B_x67f0iET4_2),.clk(gclk));
	jdff dff_B_LJ3KrJqL9_2(.din(w_dff_B_x67f0iET4_2),.dout(w_dff_B_LJ3KrJqL9_2),.clk(gclk));
	jdff dff_A_uK3mcUtQ1_0(.dout(w_G4432_1[0]),.din(w_dff_A_uK3mcUtQ1_0),.clk(gclk));
	jdff dff_A_MJoPGurE9_0(.dout(w_dff_A_uK3mcUtQ1_0),.din(w_dff_A_MJoPGurE9_0),.clk(gclk));
	jdff dff_A_xLxDpNkr2_0(.dout(w_dff_A_MJoPGurE9_0),.din(w_dff_A_xLxDpNkr2_0),.clk(gclk));
	jdff dff_A_A9SH6JlV4_0(.dout(w_dff_A_xLxDpNkr2_0),.din(w_dff_A_A9SH6JlV4_0),.clk(gclk));
	jdff dff_B_m00CwWkB1_1(.din(n1637),.dout(w_dff_B_m00CwWkB1_1),.clk(gclk));
	jdff dff_B_lKlqVw6l0_1(.din(w_dff_B_m00CwWkB1_1),.dout(w_dff_B_lKlqVw6l0_1),.clk(gclk));
	jdff dff_B_op9X8sWH4_1(.din(w_dff_B_lKlqVw6l0_1),.dout(w_dff_B_op9X8sWH4_1),.clk(gclk));
	jdff dff_B_At9nBWda5_1(.din(w_dff_B_op9X8sWH4_1),.dout(w_dff_B_At9nBWda5_1),.clk(gclk));
	jdff dff_B_oDjgaoxa9_1(.din(w_dff_B_At9nBWda5_1),.dout(w_dff_B_oDjgaoxa9_1),.clk(gclk));
	jdff dff_B_jLjsK8R24_1(.din(w_dff_B_oDjgaoxa9_1),.dout(w_dff_B_jLjsK8R24_1),.clk(gclk));
	jdff dff_B_J3vu9VkB6_1(.din(w_dff_B_jLjsK8R24_1),.dout(w_dff_B_J3vu9VkB6_1),.clk(gclk));
	jdff dff_B_khkA4of51_1(.din(w_dff_B_J3vu9VkB6_1),.dout(w_dff_B_khkA4of51_1),.clk(gclk));
	jdff dff_B_hZAdVbBO1_1(.din(w_dff_B_khkA4of51_1),.dout(w_dff_B_hZAdVbBO1_1),.clk(gclk));
	jdff dff_B_9TVi3SFO8_1(.din(w_dff_B_hZAdVbBO1_1),.dout(w_dff_B_9TVi3SFO8_1),.clk(gclk));
	jdff dff_B_jQok6wNt8_1(.din(w_dff_B_9TVi3SFO8_1),.dout(w_dff_B_jQok6wNt8_1),.clk(gclk));
	jdff dff_B_5vbgQBOk3_1(.din(w_dff_B_jQok6wNt8_1),.dout(w_dff_B_5vbgQBOk3_1),.clk(gclk));
	jdff dff_B_SVwCx3Jk3_1(.din(w_dff_B_5vbgQBOk3_1),.dout(w_dff_B_SVwCx3Jk3_1),.clk(gclk));
	jdff dff_B_6RsXKspr8_1(.din(w_dff_B_SVwCx3Jk3_1),.dout(w_dff_B_6RsXKspr8_1),.clk(gclk));
	jdff dff_B_dhPpRk0k0_1(.din(w_dff_B_6RsXKspr8_1),.dout(w_dff_B_dhPpRk0k0_1),.clk(gclk));
	jdff dff_B_irw7pONr3_1(.din(n1666),.dout(w_dff_B_irw7pONr3_1),.clk(gclk));
	jdff dff_B_s4b1bcjP6_1(.din(w_dff_B_irw7pONr3_1),.dout(w_dff_B_s4b1bcjP6_1),.clk(gclk));
	jdff dff_B_M2fLyGP78_1(.din(w_dff_B_s4b1bcjP6_1),.dout(w_dff_B_M2fLyGP78_1),.clk(gclk));
	jdff dff_B_IzjJuRlZ8_0(.din(n1705),.dout(w_dff_B_IzjJuRlZ8_0),.clk(gclk));
	jdff dff_B_BBzXyyqI9_1(.din(n1702),.dout(w_dff_B_BBzXyyqI9_1),.clk(gclk));
	jdff dff_B_lFsbFdkU4_1(.din(w_dff_B_BBzXyyqI9_1),.dout(w_dff_B_lFsbFdkU4_1),.clk(gclk));
	jdff dff_B_b9J8I6ba1_0(.din(n1698),.dout(w_dff_B_b9J8I6ba1_0),.clk(gclk));
	jdff dff_B_4ZB7phqf9_0(.din(w_dff_B_b9J8I6ba1_0),.dout(w_dff_B_4ZB7phqf9_0),.clk(gclk));
	jdff dff_B_BRgOB9fC5_0(.din(w_dff_B_4ZB7phqf9_0),.dout(w_dff_B_BRgOB9fC5_0),.clk(gclk));
	jdff dff_B_2PExhUiz4_0(.din(w_dff_B_BRgOB9fC5_0),.dout(w_dff_B_2PExhUiz4_0),.clk(gclk));
	jdff dff_B_MB2iYhoR7_0(.din(w_dff_B_2PExhUiz4_0),.dout(w_dff_B_MB2iYhoR7_0),.clk(gclk));
	jdff dff_B_9LO6AAe94_0(.din(w_dff_B_MB2iYhoR7_0),.dout(w_dff_B_9LO6AAe94_0),.clk(gclk));
	jdff dff_B_mcHUToWf6_0(.din(w_dff_B_9LO6AAe94_0),.dout(w_dff_B_mcHUToWf6_0),.clk(gclk));
	jdff dff_B_gm9gynBi1_1(.din(n1690),.dout(w_dff_B_gm9gynBi1_1),.clk(gclk));
	jdff dff_B_QFJrQ7Xm1_1(.din(w_dff_B_gm9gynBi1_1),.dout(w_dff_B_QFJrQ7Xm1_1),.clk(gclk));
	jdff dff_B_o4Bl01oL7_1(.din(w_dff_B_QFJrQ7Xm1_1),.dout(w_dff_B_o4Bl01oL7_1),.clk(gclk));
	jdff dff_B_4cJYevke8_1(.din(w_dff_B_o4Bl01oL7_1),.dout(w_dff_B_4cJYevke8_1),.clk(gclk));
	jdff dff_B_wOKvsKX93_1(.din(w_dff_B_4cJYevke8_1),.dout(w_dff_B_wOKvsKX93_1),.clk(gclk));
	jdff dff_B_aCsvP5CA5_1(.din(n1691),.dout(w_dff_B_aCsvP5CA5_1),.clk(gclk));
	jdff dff_B_YU5oIvu96_1(.din(w_dff_B_aCsvP5CA5_1),.dout(w_dff_B_YU5oIvu96_1),.clk(gclk));
	jdff dff_B_MW7VhB9m1_1(.din(w_dff_B_YU5oIvu96_1),.dout(w_dff_B_MW7VhB9m1_1),.clk(gclk));
	jdff dff_B_O5UXEisZ1_1(.din(w_dff_B_MW7VhB9m1_1),.dout(w_dff_B_O5UXEisZ1_1),.clk(gclk));
	jdff dff_A_huJLn5st9_1(.dout(w_n1687_0[1]),.din(w_dff_A_huJLn5st9_1),.clk(gclk));
	jdff dff_A_CUMEv2pZ1_1(.dout(w_dff_A_huJLn5st9_1),.din(w_dff_A_CUMEv2pZ1_1),.clk(gclk));
	jdff dff_A_I6t17dkg8_1(.dout(w_dff_A_CUMEv2pZ1_1),.din(w_dff_A_I6t17dkg8_1),.clk(gclk));
	jdff dff_A_PJc2GGi80_1(.dout(w_dff_A_I6t17dkg8_1),.din(w_dff_A_PJc2GGi80_1),.clk(gclk));
	jdff dff_B_TJ6gxjLw2_1(.din(n1683),.dout(w_dff_B_TJ6gxjLw2_1),.clk(gclk));
	jdff dff_A_2h9RBzpc9_0(.dout(w_n1127_0[0]),.din(w_dff_A_2h9RBzpc9_0),.clk(gclk));
	jdff dff_A_Q55QeYa29_0(.dout(w_dff_A_2h9RBzpc9_0),.din(w_dff_A_Q55QeYa29_0),.clk(gclk));
	jdff dff_A_DL60yFMg3_0(.dout(w_dff_A_Q55QeYa29_0),.din(w_dff_A_DL60yFMg3_0),.clk(gclk));
	jdff dff_B_urJFtoOG4_2(.din(n1127),.dout(w_dff_B_urJFtoOG4_2),.clk(gclk));
	jdff dff_B_0YojitN27_2(.din(w_dff_B_urJFtoOG4_2),.dout(w_dff_B_0YojitN27_2),.clk(gclk));
	jdff dff_B_GYOl95Xk6_2(.din(w_dff_B_0YojitN27_2),.dout(w_dff_B_GYOl95Xk6_2),.clk(gclk));
	jdff dff_B_K27cHxuK1_2(.din(w_dff_B_GYOl95Xk6_2),.dout(w_dff_B_K27cHxuK1_2),.clk(gclk));
	jdff dff_A_iNx813JT8_1(.dout(w_n1675_0[1]),.din(w_dff_A_iNx813JT8_1),.clk(gclk));
	jdff dff_A_1oOPgSJ67_1(.dout(w_dff_A_iNx813JT8_1),.din(w_dff_A_1oOPgSJ67_1),.clk(gclk));
	jdff dff_A_xRUPsRID2_1(.dout(w_dff_A_1oOPgSJ67_1),.din(w_dff_A_xRUPsRID2_1),.clk(gclk));
	jdff dff_B_9EZizkRl8_1(.din(n1669),.dout(w_dff_B_9EZizkRl8_1),.clk(gclk));
	jdff dff_B_HpY57gf01_1(.din(w_dff_B_9EZizkRl8_1),.dout(w_dff_B_HpY57gf01_1),.clk(gclk));
	jdff dff_B_n0jEM33v8_0(.din(n1671),.dout(w_dff_B_n0jEM33v8_0),.clk(gclk));
	jdff dff_B_LG4LL9yI8_0(.din(w_dff_B_n0jEM33v8_0),.dout(w_dff_B_LG4LL9yI8_0),.clk(gclk));
	jdff dff_A_PfUyz38B3_0(.dout(w_n1667_0[0]),.din(w_dff_A_PfUyz38B3_0),.clk(gclk));
	jdff dff_A_qPYvkuac0_0(.dout(w_dff_A_PfUyz38B3_0),.din(w_dff_A_qPYvkuac0_0),.clk(gclk));
	jdff dff_A_1G1L2k840_0(.dout(w_dff_A_qPYvkuac0_0),.din(w_dff_A_1G1L2k840_0),.clk(gclk));
	jdff dff_A_c9mCUYb77_1(.dout(w_n1136_0[1]),.din(w_dff_A_c9mCUYb77_1),.clk(gclk));
	jdff dff_B_ZBD1w1uZ9_1(.din(n1649),.dout(w_dff_B_ZBD1w1uZ9_1),.clk(gclk));
	jdff dff_B_GfJ845uw0_1(.din(w_dff_B_ZBD1w1uZ9_1),.dout(w_dff_B_GfJ845uw0_1),.clk(gclk));
	jdff dff_B_db5qHDMU1_1(.din(w_dff_B_GfJ845uw0_1),.dout(w_dff_B_db5qHDMU1_1),.clk(gclk));
	jdff dff_B_PXdKW4HM7_1(.din(n1660),.dout(w_dff_B_PXdKW4HM7_1),.clk(gclk));
	jdff dff_B_X5INP1zd1_1(.din(w_dff_B_PXdKW4HM7_1),.dout(w_dff_B_X5INP1zd1_1),.clk(gclk));
	jdff dff_B_LU6sU5v11_1(.din(n1661),.dout(w_dff_B_LU6sU5v11_1),.clk(gclk));
	jdff dff_B_jGBSEGLF8_1(.din(w_dff_B_LU6sU5v11_1),.dout(w_dff_B_jGBSEGLF8_1),.clk(gclk));
	jdff dff_B_GhpJh8ku0_1(.din(w_dff_B_jGBSEGLF8_1),.dout(w_dff_B_GhpJh8ku0_1),.clk(gclk));
	jdff dff_B_0Gr5VV637_1(.din(w_dff_B_GhpJh8ku0_1),.dout(w_dff_B_0Gr5VV637_1),.clk(gclk));
	jdff dff_B_ca3YkLIG2_1(.din(w_dff_B_0Gr5VV637_1),.dout(w_dff_B_ca3YkLIG2_1),.clk(gclk));
	jdff dff_A_fKpm5dyE3_0(.dout(w_n1376_0[0]),.din(w_dff_A_fKpm5dyE3_0),.clk(gclk));
	jdff dff_A_FMnGLo105_0(.dout(w_dff_A_fKpm5dyE3_0),.din(w_dff_A_FMnGLo105_0),.clk(gclk));
	jdff dff_A_fYmTU2qH0_0(.dout(w_dff_A_FMnGLo105_0),.din(w_dff_A_fYmTU2qH0_0),.clk(gclk));
	jdff dff_A_tDZA1xRC0_0(.dout(w_dff_A_fYmTU2qH0_0),.din(w_dff_A_tDZA1xRC0_0),.clk(gclk));
	jdff dff_B_pO9vYmEx8_1(.din(n1366),.dout(w_dff_B_pO9vYmEx8_1),.clk(gclk));
	jdff dff_A_jO2s0pGZ6_1(.dout(w_n1361_0[1]),.din(w_dff_A_jO2s0pGZ6_1),.clk(gclk));
	jdff dff_A_VKwZtXWT9_0(.dout(w_G3705_1[0]),.din(w_dff_A_VKwZtXWT9_0),.clk(gclk));
	jdff dff_A_vMV7Up726_0(.dout(w_dff_A_VKwZtXWT9_0),.din(w_dff_A_vMV7Up726_0),.clk(gclk));
	jdff dff_A_OAlXRzLj4_0(.dout(w_dff_A_vMV7Up726_0),.din(w_dff_A_OAlXRzLj4_0),.clk(gclk));
	jdff dff_A_AMzFpknM9_1(.dout(w_G3705_1[1]),.din(w_dff_A_AMzFpknM9_1),.clk(gclk));
	jdff dff_A_lSW5RBm45_1(.dout(w_dff_A_AMzFpknM9_1),.din(w_dff_A_lSW5RBm45_1),.clk(gclk));
	jdff dff_A_PSFGRNPQ9_1(.dout(w_dff_A_lSW5RBm45_1),.din(w_dff_A_PSFGRNPQ9_1),.clk(gclk));
	jdff dff_A_0t1fKIX47_0(.dout(w_n362_0[0]),.din(w_dff_A_0t1fKIX47_0),.clk(gclk));
	jdff dff_A_u3HAFNlj0_0(.dout(w_dff_A_0t1fKIX47_0),.din(w_dff_A_u3HAFNlj0_0),.clk(gclk));
	jdff dff_A_aacO2efu7_0(.dout(w_dff_A_u3HAFNlj0_0),.din(w_dff_A_aacO2efu7_0),.clk(gclk));
	jdff dff_A_EciIcRXr9_0(.dout(w_dff_A_aacO2efu7_0),.din(w_dff_A_EciIcRXr9_0),.clk(gclk));
	jdff dff_A_QVIFmCto7_0(.dout(w_dff_A_EciIcRXr9_0),.din(w_dff_A_QVIFmCto7_0),.clk(gclk));
	jdff dff_B_wb1SXgaB4_0(.din(n357),.dout(w_dff_B_wb1SXgaB4_0),.clk(gclk));
	jdff dff_A_BskuEaBp5_1(.dout(w_n1360_1[1]),.din(w_dff_A_BskuEaBp5_1),.clk(gclk));
	jdff dff_A_8DGK2zaE1_1(.dout(w_dff_A_BskuEaBp5_1),.din(w_dff_A_8DGK2zaE1_1),.clk(gclk));
	jdff dff_A_16N29usL4_1(.dout(w_n1359_0[1]),.din(w_dff_A_16N29usL4_1),.clk(gclk));
	jdff dff_A_4hPMsaKX4_2(.dout(w_n1359_0[2]),.din(w_dff_A_4hPMsaKX4_2),.clk(gclk));
	jdff dff_A_pKYTFRI76_2(.dout(w_dff_A_4hPMsaKX4_2),.din(w_dff_A_pKYTFRI76_2),.clk(gclk));
	jdff dff_B_dxIieSIK9_0(.din(n1358),.dout(w_dff_B_dxIieSIK9_0),.clk(gclk));
	jdff dff_A_2GEKLgiy4_0(.dout(w_G3717_1[0]),.din(w_dff_A_2GEKLgiy4_0),.clk(gclk));
	jdff dff_A_ue6tcNJq6_0(.dout(w_dff_A_2GEKLgiy4_0),.din(w_dff_A_ue6tcNJq6_0),.clk(gclk));
	jdff dff_A_5mFDGhUz1_0(.dout(w_dff_A_ue6tcNJq6_0),.din(w_dff_A_5mFDGhUz1_0),.clk(gclk));
	jdff dff_A_LnyQNl3O7_1(.dout(w_G3717_1[1]),.din(w_dff_A_LnyQNl3O7_1),.clk(gclk));
	jdff dff_A_pHzc0oGT9_1(.dout(w_dff_A_LnyQNl3O7_1),.din(w_dff_A_pHzc0oGT9_1),.clk(gclk));
	jdff dff_A_4OpryYFd5_1(.dout(w_dff_A_pHzc0oGT9_1),.din(w_dff_A_4OpryYFd5_1),.clk(gclk));
	jdff dff_B_L31IHJIT9_0(.din(n1658),.dout(w_dff_B_L31IHJIT9_0),.clk(gclk));
	jdff dff_B_loaANmcM8_0(.din(w_dff_B_L31IHJIT9_0),.dout(w_dff_B_loaANmcM8_0),.clk(gclk));
	jdff dff_B_K4lgHV8e3_0(.din(w_dff_B_loaANmcM8_0),.dout(w_dff_B_K4lgHV8e3_0),.clk(gclk));
	jdff dff_B_c83Pyh6j7_0(.din(w_dff_B_K4lgHV8e3_0),.dout(w_dff_B_c83Pyh6j7_0),.clk(gclk));
	jdff dff_A_Jhv9FVMp7_1(.dout(w_n1654_0[1]),.din(w_dff_A_Jhv9FVMp7_1),.clk(gclk));
	jdff dff_A_q80ykMn44_1(.dout(w_dff_A_Jhv9FVMp7_1),.din(w_dff_A_q80ykMn44_1),.clk(gclk));
	jdff dff_A_eGSqPnke0_1(.dout(w_dff_A_q80ykMn44_1),.din(w_dff_A_eGSqPnke0_1),.clk(gclk));
	jdff dff_A_2Y9KbueZ0_1(.dout(w_n462_0[1]),.din(w_dff_A_2Y9KbueZ0_1),.clk(gclk));
	jdff dff_A_NOCwwBkH1_1(.dout(w_dff_A_2Y9KbueZ0_1),.din(w_dff_A_NOCwwBkH1_1),.clk(gclk));
	jdff dff_A_TNk2zobb9_1(.dout(w_dff_A_NOCwwBkH1_1),.din(w_dff_A_TNk2zobb9_1),.clk(gclk));
	jdff dff_A_3ashGlaE8_1(.dout(w_dff_A_TNk2zobb9_1),.din(w_dff_A_3ashGlaE8_1),.clk(gclk));
	jdff dff_A_s5TRwFlx1_1(.dout(w_n1651_0[1]),.din(w_dff_A_s5TRwFlx1_1),.clk(gclk));
	jdff dff_A_hMPxqBCX0_1(.dout(w_dff_A_s5TRwFlx1_1),.din(w_dff_A_hMPxqBCX0_1),.clk(gclk));
	jdff dff_A_NBGRQgba6_1(.dout(w_dff_A_hMPxqBCX0_1),.din(w_dff_A_NBGRQgba6_1),.clk(gclk));
	jdff dff_A_NXQDkBSO4_1(.dout(w_dff_A_NBGRQgba6_1),.din(w_dff_A_NXQDkBSO4_1),.clk(gclk));
	jdff dff_A_1oemz8iY6_1(.dout(w_dff_A_NXQDkBSO4_1),.din(w_dff_A_1oemz8iY6_1),.clk(gclk));
	jdff dff_B_toRcHFRg4_0(.din(n1650),.dout(w_dff_B_toRcHFRg4_0),.clk(gclk));
	jdff dff_A_rLLsVKt47_1(.dout(w_n422_0[1]),.din(w_dff_A_rLLsVKt47_1),.clk(gclk));
	jdff dff_A_R2SucpmA7_1(.dout(w_n419_0[1]),.din(w_dff_A_R2SucpmA7_1),.clk(gclk));
	jdff dff_B_K4gcKoet5_1(.din(n415),.dout(w_dff_B_K4gcKoet5_1),.clk(gclk));
	jdff dff_A_zYrrV5Nr2_0(.dout(w_n417_0[0]),.din(w_dff_A_zYrrV5Nr2_0),.clk(gclk));
	jdff dff_A_hLSbtrog4_0(.dout(w_dff_A_zYrrV5Nr2_0),.din(w_dff_A_hLSbtrog4_0),.clk(gclk));
	jdff dff_A_BUUQM5Am5_0(.dout(w_dff_A_hLSbtrog4_0),.din(w_dff_A_BUUQM5Am5_0),.clk(gclk));
	jdff dff_A_ge3nwBvm9_0(.dout(w_dff_A_BUUQM5Am5_0),.din(w_dff_A_ge3nwBvm9_0),.clk(gclk));
	jdff dff_A_74ChuIys9_0(.dout(w_dff_A_ge3nwBvm9_0),.din(w_dff_A_74ChuIys9_0),.clk(gclk));
	jdff dff_A_9zZV5BU62_0(.dout(w_dff_A_74ChuIys9_0),.din(w_dff_A_9zZV5BU62_0),.clk(gclk));
	jdff dff_A_xw4mA3Og7_0(.dout(w_dff_A_9zZV5BU62_0),.din(w_dff_A_xw4mA3Og7_0),.clk(gclk));
	jdff dff_A_Lz0Uftj19_0(.dout(w_dff_A_xw4mA3Og7_0),.din(w_dff_A_Lz0Uftj19_0),.clk(gclk));
	jdff dff_A_ynFzRE1J4_1(.dout(w_n417_0[1]),.din(w_dff_A_ynFzRE1J4_1),.clk(gclk));
	jdff dff_A_YrfkQ3QR3_1(.dout(w_dff_A_ynFzRE1J4_1),.din(w_dff_A_YrfkQ3QR3_1),.clk(gclk));
	jdff dff_A_ErMpNqaH7_1(.dout(w_dff_A_YrfkQ3QR3_1),.din(w_dff_A_ErMpNqaH7_1),.clk(gclk));
	jdff dff_A_GsEEhB1g8_1(.dout(w_dff_A_ErMpNqaH7_1),.din(w_dff_A_GsEEhB1g8_1),.clk(gclk));
	jdff dff_A_yo6ADf9Q9_1(.dout(w_dff_A_GsEEhB1g8_1),.din(w_dff_A_yo6ADf9Q9_1),.clk(gclk));
	jdff dff_A_MXCZR0Z74_0(.dout(w_n413_1[0]),.din(w_dff_A_MXCZR0Z74_0),.clk(gclk));
	jdff dff_A_XCnpn9aE4_0(.dout(w_n413_0[0]),.din(w_dff_A_XCnpn9aE4_0),.clk(gclk));
	jdff dff_A_b2VlgxhT9_0(.dout(w_n412_0[0]),.din(w_dff_A_b2VlgxhT9_0),.clk(gclk));
	jdff dff_A_tUXNCgyV3_1(.dout(w_n412_0[1]),.din(w_dff_A_tUXNCgyV3_1),.clk(gclk));
	jdff dff_A_eb3uJuHK3_0(.dout(w_n354_1[0]),.din(w_dff_A_eb3uJuHK3_0),.clk(gclk));
	jdff dff_A_KfyikFRM7_0(.dout(w_dff_A_eb3uJuHK3_0),.din(w_dff_A_KfyikFRM7_0),.clk(gclk));
	jdff dff_A_1jGxRfYS0_2(.dout(w_n354_0[2]),.din(w_dff_A_1jGxRfYS0_2),.clk(gclk));
	jdff dff_A_U16CpbZ10_2(.dout(w_dff_A_1jGxRfYS0_2),.din(w_dff_A_U16CpbZ10_2),.clk(gclk));
	jdff dff_A_RlLKWvkN5_2(.dout(w_dff_A_U16CpbZ10_2),.din(w_dff_A_RlLKWvkN5_2),.clk(gclk));
	jdff dff_A_S3JU1x8F2_2(.dout(w_dff_A_RlLKWvkN5_2),.din(w_dff_A_S3JU1x8F2_2),.clk(gclk));
	jdff dff_A_YpwkgRTq9_2(.dout(w_dff_A_S3JU1x8F2_2),.din(w_dff_A_YpwkgRTq9_2),.clk(gclk));
	jdff dff_A_C5QUNZM13_2(.dout(w_dff_A_YpwkgRTq9_2),.din(w_dff_A_C5QUNZM13_2),.clk(gclk));
	jdff dff_A_JAuJ1xwf2_2(.dout(w_dff_A_C5QUNZM13_2),.din(w_dff_A_JAuJ1xwf2_2),.clk(gclk));
	jdff dff_A_vEMXFiWM5_2(.dout(w_dff_A_JAuJ1xwf2_2),.din(w_dff_A_vEMXFiWM5_2),.clk(gclk));
	jdff dff_A_RBqqfmj90_2(.dout(w_dff_A_vEMXFiWM5_2),.din(w_dff_A_RBqqfmj90_2),.clk(gclk));
	jdff dff_A_rNHh4MfQ2_2(.dout(w_dff_A_RBqqfmj90_2),.din(w_dff_A_rNHh4MfQ2_2),.clk(gclk));
	jdff dff_B_dy0x9oPk3_3(.din(n354),.dout(w_dff_B_dy0x9oPk3_3),.clk(gclk));
	jdff dff_A_wWuBBJtQ6_2(.dout(w_n407_0[2]),.din(w_dff_A_wWuBBJtQ6_2),.clk(gclk));
	jdff dff_A_0n0NhMk98_2(.dout(w_dff_A_wWuBBJtQ6_2),.din(w_dff_A_0n0NhMk98_2),.clk(gclk));
	jdff dff_A_7Qn0UCgU2_1(.dout(w_n402_1[1]),.din(w_dff_A_7Qn0UCgU2_1),.clk(gclk));
	jdff dff_A_q3xzslil1_1(.dout(w_n402_0[1]),.din(w_dff_A_q3xzslil1_1),.clk(gclk));
	jdff dff_A_tGm2WAAL5_1(.dout(w_dff_A_q3xzslil1_1),.din(w_dff_A_tGm2WAAL5_1),.clk(gclk));
	jdff dff_A_E8O9XLfM7_1(.dout(w_dff_A_tGm2WAAL5_1),.din(w_dff_A_E8O9XLfM7_1),.clk(gclk));
	jdff dff_A_UFOubWhK7_1(.dout(w_dff_A_E8O9XLfM7_1),.din(w_dff_A_UFOubWhK7_1),.clk(gclk));
	jdff dff_A_pVaAoIcP4_1(.dout(w_dff_A_UFOubWhK7_1),.din(w_dff_A_pVaAoIcP4_1),.clk(gclk));
	jdff dff_A_FzS2S2zR1_1(.dout(w_dff_A_pVaAoIcP4_1),.din(w_dff_A_FzS2S2zR1_1),.clk(gclk));
	jdff dff_A_OzwzaeGN9_1(.dout(w_dff_A_FzS2S2zR1_1),.din(w_dff_A_OzwzaeGN9_1),.clk(gclk));
	jdff dff_A_kv03YZqk2_1(.dout(w_dff_A_OzwzaeGN9_1),.din(w_dff_A_kv03YZqk2_1),.clk(gclk));
	jdff dff_A_DwwcC0kn8_1(.dout(w_dff_A_kv03YZqk2_1),.din(w_dff_A_DwwcC0kn8_1),.clk(gclk));
	jdff dff_A_dlbfW2eX1_2(.dout(w_n402_0[2]),.din(w_dff_A_dlbfW2eX1_2),.clk(gclk));
	jdff dff_A_fCONKPFv9_2(.dout(w_dff_A_dlbfW2eX1_2),.din(w_dff_A_fCONKPFv9_2),.clk(gclk));
	jdff dff_A_7BZFgUcx4_2(.dout(w_dff_A_fCONKPFv9_2),.din(w_dff_A_7BZFgUcx4_2),.clk(gclk));
	jdff dff_B_CnzNEovY4_1(.din(n396),.dout(w_dff_B_CnzNEovY4_1),.clk(gclk));
	jdff dff_B_hZCxe38Z9_1(.din(w_dff_B_CnzNEovY4_1),.dout(w_dff_B_hZCxe38Z9_1),.clk(gclk));
	jdff dff_A_sPVJRPqW6_0(.dout(w_G3705_2[0]),.din(w_dff_A_sPVJRPqW6_0),.clk(gclk));
	jdff dff_A_KD5l7uKl2_0(.dout(w_dff_A_sPVJRPqW6_0),.din(w_dff_A_KD5l7uKl2_0),.clk(gclk));
	jdff dff_A_tQXoU1Lv0_0(.dout(w_dff_A_KD5l7uKl2_0),.din(w_dff_A_tQXoU1Lv0_0),.clk(gclk));
	jdff dff_A_my3fTdNO3_0(.dout(w_n395_0[0]),.din(w_dff_A_my3fTdNO3_0),.clk(gclk));
	jdff dff_A_Nbe0h9oQ0_0(.dout(w_n359_0[0]),.din(w_dff_A_Nbe0h9oQ0_0),.clk(gclk));
	jdff dff_A_86X0fj5T4_1(.dout(w_G3701_1[1]),.din(w_dff_A_86X0fj5T4_1),.clk(gclk));
	jdff dff_A_vTR1YCna4_2(.dout(w_n390_0[2]),.din(w_dff_A_vTR1YCna4_2),.clk(gclk));
	jdff dff_A_574BHCIW0_2(.dout(w_dff_A_vTR1YCna4_2),.din(w_dff_A_574BHCIW0_2),.clk(gclk));
	jdff dff_A_Ijknd9154_2(.dout(w_dff_A_574BHCIW0_2),.din(w_dff_A_Ijknd9154_2),.clk(gclk));
	jdff dff_A_xkbWnlis2_2(.dout(w_dff_A_Ijknd9154_2),.din(w_dff_A_xkbWnlis2_2),.clk(gclk));
	jdff dff_A_tq5Yg5jr0_2(.dout(w_dff_A_xkbWnlis2_2),.din(w_dff_A_tq5Yg5jr0_2),.clk(gclk));
	jdff dff_B_PjRmLE2K8_3(.din(n390),.dout(w_dff_B_PjRmLE2K8_3),.clk(gclk));
	jdff dff_A_0qBs17pA6_0(.dout(w_n356_0[0]),.din(w_dff_A_0qBs17pA6_0),.clk(gclk));
	jdff dff_A_KWKXI7In8_0(.dout(w_G41_0[0]),.din(w_dff_A_KWKXI7In8_0),.clk(gclk));
	jdff dff_A_G2VPD0zK0_0(.dout(w_dff_A_KWKXI7In8_0),.din(w_dff_A_G2VPD0zK0_0),.clk(gclk));
	jdff dff_A_E1lKdqdn1_0(.dout(w_dff_A_G2VPD0zK0_0),.din(w_dff_A_E1lKdqdn1_0),.clk(gclk));
	jdff dff_A_1rd0G7VB5_1(.dout(w_G41_0[1]),.din(w_dff_A_1rd0G7VB5_1),.clk(gclk));
	jdff dff_A_OMo2FIRs2_1(.dout(w_n389_0[1]),.din(w_dff_A_OMo2FIRs2_1),.clk(gclk));
	jdff dff_A_mENYvAB70_0(.dout(w_G3701_0[0]),.din(w_dff_A_mENYvAB70_0),.clk(gclk));
	jdff dff_A_2JLbCXVs9_0(.dout(w_n388_0[0]),.din(w_dff_A_2JLbCXVs9_0),.clk(gclk));
	jdff dff_A_Ad37vWO88_0(.dout(w_dff_A_2JLbCXVs9_0),.din(w_dff_A_Ad37vWO88_0),.clk(gclk));
	jdff dff_A_iigKqD6s2_0(.dout(w_dff_A_Ad37vWO88_0),.din(w_dff_A_iigKqD6s2_0),.clk(gclk));
	jdff dff_A_3rHATCLF8_0(.dout(w_dff_A_iigKqD6s2_0),.din(w_dff_A_3rHATCLF8_0),.clk(gclk));
	jdff dff_A_BLi0UKQr9_0(.dout(w_dff_A_3rHATCLF8_0),.din(w_dff_A_BLi0UKQr9_0),.clk(gclk));
	jdff dff_A_76LSyMpR6_0(.dout(w_dff_A_BLi0UKQr9_0),.din(w_dff_A_76LSyMpR6_0),.clk(gclk));
	jdff dff_A_InABorcy2_0(.dout(w_dff_A_76LSyMpR6_0),.din(w_dff_A_InABorcy2_0),.clk(gclk));
	jdff dff_A_suXKcclV2_0(.dout(w_dff_A_InABorcy2_0),.din(w_dff_A_suXKcclV2_0),.clk(gclk));
	jdff dff_A_prRyeJR16_0(.dout(w_dff_A_suXKcclV2_0),.din(w_dff_A_prRyeJR16_0),.clk(gclk));
	jdff dff_A_SWBB6UnT6_0(.dout(w_dff_A_prRyeJR16_0),.din(w_dff_A_SWBB6UnT6_0),.clk(gclk));
	jdff dff_A_cuIgAHEu2_0(.dout(w_dff_A_SWBB6UnT6_0),.din(w_dff_A_cuIgAHEu2_0),.clk(gclk));
	jdff dff_A_g0dGJFmc4_2(.dout(w_n388_0[2]),.din(w_dff_A_g0dGJFmc4_2),.clk(gclk));
	jdff dff_B_FV2WavSE5_3(.din(n388),.dout(w_dff_B_FV2WavSE5_3),.clk(gclk));
	jdff dff_B_UoKPGbX53_3(.din(w_dff_B_FV2WavSE5_3),.dout(w_dff_B_UoKPGbX53_3),.clk(gclk));
	jdff dff_B_QVtI5MwH7_3(.din(w_dff_B_UoKPGbX53_3),.dout(w_dff_B_QVtI5MwH7_3),.clk(gclk));
	jdff dff_B_saPTinh99_3(.din(w_dff_B_QVtI5MwH7_3),.dout(w_dff_B_saPTinh99_3),.clk(gclk));
	jdff dff_A_Kou2KRdq7_1(.dout(w_G4526_1[1]),.din(w_dff_A_Kou2KRdq7_1),.clk(gclk));
	jdff dff_A_Af6X7UU30_1(.dout(w_dff_A_Kou2KRdq7_1),.din(w_dff_A_Af6X7UU30_1),.clk(gclk));
	jdff dff_A_eaja6E129_1(.dout(w_dff_A_Af6X7UU30_1),.din(w_dff_A_eaja6E129_1),.clk(gclk));
	jdff dff_A_Vq2ID94O4_1(.dout(w_dff_A_eaja6E129_1),.din(w_dff_A_Vq2ID94O4_1),.clk(gclk));
	jdff dff_A_KWA32Iz23_1(.dout(w_dff_A_Vq2ID94O4_1),.din(w_dff_A_KWA32Iz23_1),.clk(gclk));
	jdff dff_A_R4UfypZu6_1(.dout(w_G4526_0[1]),.din(w_dff_A_R4UfypZu6_1),.clk(gclk));
	jdff dff_A_fk14z9ty7_1(.dout(w_dff_A_R4UfypZu6_1),.din(w_dff_A_fk14z9ty7_1),.clk(gclk));
	jdff dff_A_ef5Ya6w85_1(.dout(w_dff_A_fk14z9ty7_1),.din(w_dff_A_ef5Ya6w85_1),.clk(gclk));
	jdff dff_A_EEK5FmLK4_1(.dout(w_dff_A_ef5Ya6w85_1),.din(w_dff_A_EEK5FmLK4_1),.clk(gclk));
	jdff dff_A_Rsp5iJf80_1(.dout(w_dff_A_EEK5FmLK4_1),.din(w_dff_A_Rsp5iJf80_1),.clk(gclk));
	jdff dff_A_OnJU2gOs5_1(.dout(w_dff_A_Rsp5iJf80_1),.din(w_dff_A_OnJU2gOs5_1),.clk(gclk));
	jdff dff_A_MvC8enj97_1(.dout(w_dff_A_OnJU2gOs5_1),.din(w_dff_A_MvC8enj97_1),.clk(gclk));
	jdff dff_A_amY1LlFT9_1(.dout(w_dff_A_MvC8enj97_1),.din(w_dff_A_amY1LlFT9_1),.clk(gclk));
	jdff dff_A_DfeiJWSB7_1(.dout(w_dff_A_amY1LlFT9_1),.din(w_dff_A_DfeiJWSB7_1),.clk(gclk));
	jdff dff_A_RvJxSXRF2_1(.dout(w_dff_A_DfeiJWSB7_1),.din(w_dff_A_RvJxSXRF2_1),.clk(gclk));
	jdff dff_A_KdKlVakS3_1(.dout(w_dff_A_RvJxSXRF2_1),.din(w_dff_A_KdKlVakS3_1),.clk(gclk));
	jdff dff_A_JD3Ar4P25_1(.dout(w_dff_A_KdKlVakS3_1),.din(w_dff_A_JD3Ar4P25_1),.clk(gclk));
	jdff dff_A_exvZSVku9_1(.dout(w_dff_A_JD3Ar4P25_1),.din(w_dff_A_exvZSVku9_1),.clk(gclk));
	jdff dff_A_h7bxFk6z9_1(.dout(w_dff_A_exvZSVku9_1),.din(w_dff_A_h7bxFk6z9_1),.clk(gclk));
	jdff dff_A_7vaAMfFm2_1(.dout(w_dff_A_h7bxFk6z9_1),.din(w_dff_A_7vaAMfFm2_1),.clk(gclk));
	jdff dff_A_YZVpOyPU1_2(.dout(w_G4526_0[2]),.din(w_dff_A_YZVpOyPU1_2),.clk(gclk));
	jdff dff_A_sIBlrrHb1_2(.dout(w_dff_A_YZVpOyPU1_2),.din(w_dff_A_sIBlrrHb1_2),.clk(gclk));
	jdff dff_A_SbbCDg6y1_2(.dout(w_dff_A_sIBlrrHb1_2),.din(w_dff_A_SbbCDg6y1_2),.clk(gclk));
	jdff dff_A_9mi9xNZI5_2(.dout(w_dff_A_SbbCDg6y1_2),.din(w_dff_A_9mi9xNZI5_2),.clk(gclk));
	jdff dff_A_XvbWsxkx5_2(.dout(w_dff_A_9mi9xNZI5_2),.din(w_dff_A_XvbWsxkx5_2),.clk(gclk));
	jdff dff_A_P5m2N7wQ0_2(.dout(w_dff_A_XvbWsxkx5_2),.din(w_dff_A_P5m2N7wQ0_2),.clk(gclk));
	jdff dff_A_lsfaQNUV0_1(.dout(w_n387_1[1]),.din(w_dff_A_lsfaQNUV0_1),.clk(gclk));
	jdff dff_A_8axANUzT3_2(.dout(w_n387_1[2]),.din(w_dff_A_8axANUzT3_2),.clk(gclk));
	jdff dff_A_zk68B4uQ0_2(.dout(w_dff_A_8axANUzT3_2),.din(w_dff_A_zk68B4uQ0_2),.clk(gclk));
	jdff dff_A_S7GzmQcL3_2(.dout(w_dff_A_zk68B4uQ0_2),.din(w_dff_A_S7GzmQcL3_2),.clk(gclk));
	jdff dff_A_hLmf92Cq2_1(.dout(w_n380_0[1]),.din(w_dff_A_hLmf92Cq2_1),.clk(gclk));
	jdff dff_A_wfjjHBUE6_2(.dout(w_n380_0[2]),.din(w_dff_A_wfjjHBUE6_2),.clk(gclk));
	jdff dff_A_qFKh4Mwt1_2(.dout(w_dff_A_wfjjHBUE6_2),.din(w_dff_A_qFKh4Mwt1_2),.clk(gclk));
	jdff dff_A_X3DDNoHb1_0(.dout(w_n379_1[0]),.din(w_dff_A_X3DDNoHb1_0),.clk(gclk));
	jdff dff_A_l77Ob5Vl6_0(.dout(w_dff_A_X3DDNoHb1_0),.din(w_dff_A_l77Ob5Vl6_0),.clk(gclk));
	jdff dff_A_k12A8vKM6_0(.dout(w_dff_A_l77Ob5Vl6_0),.din(w_dff_A_k12A8vKM6_0),.clk(gclk));
	jdff dff_A_WvRS9wm33_1(.dout(w_n379_0[1]),.din(w_dff_A_WvRS9wm33_1),.clk(gclk));
	jdff dff_A_E2ls2dy89_1(.dout(w_dff_A_WvRS9wm33_1),.din(w_dff_A_E2ls2dy89_1),.clk(gclk));
	jdff dff_A_0cVCnH8u6_1(.dout(w_dff_A_E2ls2dy89_1),.din(w_dff_A_0cVCnH8u6_1),.clk(gclk));
	jdff dff_A_shkWyTIS3_1(.dout(w_dff_A_0cVCnH8u6_1),.din(w_dff_A_shkWyTIS3_1),.clk(gclk));
	jdff dff_A_zhpWkmtW3_1(.dout(w_dff_A_shkWyTIS3_1),.din(w_dff_A_zhpWkmtW3_1),.clk(gclk));
	jdff dff_A_c5Rjr2fz6_1(.dout(w_dff_A_zhpWkmtW3_1),.din(w_dff_A_c5Rjr2fz6_1),.clk(gclk));
	jdff dff_A_N5OXkWGO2_1(.dout(w_dff_A_c5Rjr2fz6_1),.din(w_dff_A_N5OXkWGO2_1),.clk(gclk));
	jdff dff_A_5K07dMlU0_1(.dout(w_dff_A_N5OXkWGO2_1),.din(w_dff_A_5K07dMlU0_1),.clk(gclk));
	jdff dff_A_ifjz7Lz00_1(.dout(w_dff_A_5K07dMlU0_1),.din(w_dff_A_ifjz7Lz00_1),.clk(gclk));
	jdff dff_A_SZ5hkSWU0_1(.dout(w_dff_A_ifjz7Lz00_1),.din(w_dff_A_SZ5hkSWU0_1),.clk(gclk));
	jdff dff_A_62c1h1sh6_1(.dout(w_dff_A_SZ5hkSWU0_1),.din(w_dff_A_62c1h1sh6_1),.clk(gclk));
	jdff dff_A_6Omdyta77_1(.dout(w_dff_A_62c1h1sh6_1),.din(w_dff_A_6Omdyta77_1),.clk(gclk));
	jdff dff_A_w24k1fuu7_1(.dout(w_dff_A_6Omdyta77_1),.din(w_dff_A_w24k1fuu7_1),.clk(gclk));
	jdff dff_A_x0axQ3Bo1_1(.dout(w_dff_A_w24k1fuu7_1),.din(w_dff_A_x0axQ3Bo1_1),.clk(gclk));
	jdff dff_A_C3zAqD5D5_2(.dout(w_n379_0[2]),.din(w_dff_A_C3zAqD5D5_2),.clk(gclk));
	jdff dff_A_RXw50PGt5_2(.dout(w_dff_A_C3zAqD5D5_2),.din(w_dff_A_RXw50PGt5_2),.clk(gclk));
	jdff dff_A_SPX8CwoT2_2(.dout(w_dff_A_RXw50PGt5_2),.din(w_dff_A_SPX8CwoT2_2),.clk(gclk));
	jdff dff_A_WLYOpdFI1_2(.dout(w_dff_A_SPX8CwoT2_2),.din(w_dff_A_WLYOpdFI1_2),.clk(gclk));
	jdff dff_A_B7jS1dD42_2(.dout(w_n377_0[2]),.din(w_dff_A_B7jS1dD42_2),.clk(gclk));
	jdff dff_A_RNZYMGlC6_1(.dout(w_G3717_2[1]),.din(w_dff_A_RNZYMGlC6_1),.clk(gclk));
	jdff dff_A_tmkzqfJY2_1(.dout(w_G3717_0[1]),.din(w_dff_A_tmkzqfJY2_1),.clk(gclk));
	jdff dff_A_uojVJZWA6_1(.dout(w_dff_A_tmkzqfJY2_1),.din(w_dff_A_uojVJZWA6_1),.clk(gclk));
	jdff dff_A_1cEzrf637_1(.dout(w_dff_A_uojVJZWA6_1),.din(w_dff_A_1cEzrf637_1),.clk(gclk));
	jdff dff_A_h1ttq40p0_1(.dout(w_n372_1[1]),.din(w_dff_A_h1ttq40p0_1),.clk(gclk));
	jdff dff_A_y3ZBwYeY9_1(.dout(w_dff_A_h1ttq40p0_1),.din(w_dff_A_y3ZBwYeY9_1),.clk(gclk));
	jdff dff_A_NgEWRMSy3_1(.dout(w_dff_A_y3ZBwYeY9_1),.din(w_dff_A_NgEWRMSy3_1),.clk(gclk));
	jdff dff_A_QQ5oLMlx3_1(.dout(w_dff_A_NgEWRMSy3_1),.din(w_dff_A_QQ5oLMlx3_1),.clk(gclk));
	jdff dff_A_Qti2oXgi2_1(.dout(w_dff_A_QQ5oLMlx3_1),.din(w_dff_A_Qti2oXgi2_1),.clk(gclk));
	jdff dff_A_LIIwCuBS1_1(.dout(w_dff_A_Qti2oXgi2_1),.din(w_dff_A_LIIwCuBS1_1),.clk(gclk));
	jdff dff_A_IhVKzAON9_1(.dout(w_dff_A_LIIwCuBS1_1),.din(w_dff_A_IhVKzAON9_1),.clk(gclk));
	jdff dff_A_tITEsiEi1_2(.dout(w_n372_1[2]),.din(w_dff_A_tITEsiEi1_2),.clk(gclk));
	jdff dff_A_a9GAOO5S5_1(.dout(w_n372_0[1]),.din(w_dff_A_a9GAOO5S5_1),.clk(gclk));
	jdff dff_A_gfk7h11r3_1(.dout(w_dff_A_a9GAOO5S5_1),.din(w_dff_A_gfk7h11r3_1),.clk(gclk));
	jdff dff_A_hd2Mqzaw6_1(.dout(w_dff_A_gfk7h11r3_1),.din(w_dff_A_hd2Mqzaw6_1),.clk(gclk));
	jdff dff_A_0VNCIHMr9_1(.dout(w_dff_A_hd2Mqzaw6_1),.din(w_dff_A_0VNCIHMr9_1),.clk(gclk));
	jdff dff_A_347Xpci38_1(.dout(w_dff_A_0VNCIHMr9_1),.din(w_dff_A_347Xpci38_1),.clk(gclk));
	jdff dff_A_qgODzEOp3_1(.dout(w_dff_A_347Xpci38_1),.din(w_dff_A_qgODzEOp3_1),.clk(gclk));
	jdff dff_A_Tn3xV7u60_2(.dout(w_n372_0[2]),.din(w_dff_A_Tn3xV7u60_2),.clk(gclk));
	jdff dff_A_ltJ4xc1Z3_2(.dout(w_dff_A_Tn3xV7u60_2),.din(w_dff_A_ltJ4xc1Z3_2),.clk(gclk));
	jdff dff_A_Zrtl5PyM0_2(.dout(w_dff_A_ltJ4xc1Z3_2),.din(w_dff_A_Zrtl5PyM0_2),.clk(gclk));
	jdff dff_A_edWdi51Q7_2(.dout(w_dff_A_Zrtl5PyM0_2),.din(w_dff_A_edWdi51Q7_2),.clk(gclk));
	jdff dff_A_7Di1SXeX2_2(.dout(w_dff_A_edWdi51Q7_2),.din(w_dff_A_7Di1SXeX2_2),.clk(gclk));
	jdff dff_A_7iVYC6bE9_2(.dout(w_dff_A_7Di1SXeX2_2),.din(w_dff_A_7iVYC6bE9_2),.clk(gclk));
	jdff dff_A_VoH33dSh0_2(.dout(w_dff_A_7iVYC6bE9_2),.din(w_dff_A_VoH33dSh0_2),.clk(gclk));
	jdff dff_A_n14xedSG8_2(.dout(w_dff_A_VoH33dSh0_2),.din(w_dff_A_n14xedSG8_2),.clk(gclk));
	jdff dff_A_sSClofRu0_1(.dout(w_G18_57[1]),.din(w_dff_A_sSClofRu0_1),.clk(gclk));
	jdff dff_A_nlsLvHub1_1(.dout(w_n366_0[1]),.din(w_dff_A_nlsLvHub1_1),.clk(gclk));
	jdff dff_A_2d9BXJgZ3_1(.dout(w_dff_A_nlsLvHub1_1),.din(w_dff_A_2d9BXJgZ3_1),.clk(gclk));
	jdff dff_A_cItkywVa0_0(.dout(w_G3723_1[0]),.din(w_dff_A_cItkywVa0_0),.clk(gclk));
	jdff dff_A_XEIQ8Suh5_0(.dout(w_dff_A_cItkywVa0_0),.din(w_dff_A_XEIQ8Suh5_0),.clk(gclk));
	jdff dff_A_dX3Ou6of5_0(.dout(w_dff_A_XEIQ8Suh5_0),.din(w_dff_A_dX3Ou6of5_0),.clk(gclk));
	jdff dff_A_UPJetWPG9_2(.dout(w_G3723_0[2]),.din(w_dff_A_UPJetWPG9_2),.clk(gclk));
	jdff dff_A_glUjB8zC3_2(.dout(w_dff_A_UPJetWPG9_2),.din(w_dff_A_glUjB8zC3_2),.clk(gclk));
	jdff dff_A_AXGb06am4_2(.dout(w_dff_A_glUjB8zC3_2),.din(w_dff_A_AXGb06am4_2),.clk(gclk));
	jdff dff_B_q47WmY2E4_0(.din(n1645),.dout(w_dff_B_q47WmY2E4_0),.clk(gclk));
	jdff dff_B_wwJofFRd7_0(.din(w_dff_B_q47WmY2E4_0),.dout(w_dff_B_wwJofFRd7_0),.clk(gclk));
	jdff dff_B_qT63xhAG7_0(.din(w_dff_B_wwJofFRd7_0),.dout(w_dff_B_qT63xhAG7_0),.clk(gclk));
	jdff dff_B_5utHCWxS3_0(.din(w_dff_B_qT63xhAG7_0),.dout(w_dff_B_5utHCWxS3_0),.clk(gclk));
	jdff dff_B_kr9fsSUC8_0(.din(w_dff_B_5utHCWxS3_0),.dout(w_dff_B_kr9fsSUC8_0),.clk(gclk));
	jdff dff_A_KBogXAzk3_0(.dout(w_n1644_0[0]),.din(w_dff_A_KBogXAzk3_0),.clk(gclk));
	jdff dff_A_697IDlBx8_0(.dout(w_dff_A_KBogXAzk3_0),.din(w_dff_A_697IDlBx8_0),.clk(gclk));
	jdff dff_A_bxwSwk7h3_0(.dout(w_dff_A_697IDlBx8_0),.din(w_dff_A_bxwSwk7h3_0),.clk(gclk));
	jdff dff_A_SQ5dMzzb5_0(.dout(w_dff_A_bxwSwk7h3_0),.din(w_dff_A_SQ5dMzzb5_0),.clk(gclk));
	jdff dff_A_G0ij57U76_0(.dout(w_dff_A_SQ5dMzzb5_0),.din(w_dff_A_G0ij57U76_0),.clk(gclk));
	jdff dff_A_MFPvexyx4_2(.dout(w_n1148_0[2]),.din(w_dff_A_MFPvexyx4_2),.clk(gclk));
	jdff dff_A_RlEgPJkJ5_2(.dout(w_dff_A_MFPvexyx4_2),.din(w_dff_A_RlEgPJkJ5_2),.clk(gclk));
	jdff dff_A_26U4zmwJ3_2(.dout(w_dff_A_RlEgPJkJ5_2),.din(w_dff_A_26U4zmwJ3_2),.clk(gclk));
	jdff dff_A_rJr8v8aj7_2(.dout(w_dff_A_26U4zmwJ3_2),.din(w_dff_A_rJr8v8aj7_2),.clk(gclk));
	jdff dff_A_qqx0P7Gd4_2(.dout(w_dff_A_rJr8v8aj7_2),.din(w_dff_A_qqx0P7Gd4_2),.clk(gclk));
	jdff dff_A_yMBoJk9R6_2(.dout(w_dff_A_qqx0P7Gd4_2),.din(w_dff_A_yMBoJk9R6_2),.clk(gclk));
	jdff dff_A_Zq4XkfBT7_2(.dout(w_n429_1[2]),.din(w_dff_A_Zq4XkfBT7_2),.clk(gclk));
	jdff dff_A_4UnqXQDH0_2(.dout(w_dff_A_Zq4XkfBT7_2),.din(w_dff_A_4UnqXQDH0_2),.clk(gclk));
	jdff dff_A_ApPtfim87_2(.dout(w_dff_A_4UnqXQDH0_2),.din(w_dff_A_ApPtfim87_2),.clk(gclk));
	jdff dff_A_71krTW544_2(.dout(w_dff_A_ApPtfim87_2),.din(w_dff_A_71krTW544_2),.clk(gclk));
	jdff dff_A_mw6XjQHc2_2(.dout(w_dff_A_71krTW544_2),.din(w_dff_A_mw6XjQHc2_2),.clk(gclk));
	jdff dff_A_maRqugNU2_2(.dout(w_dff_A_mw6XjQHc2_2),.din(w_dff_A_maRqugNU2_2),.clk(gclk));
	jdff dff_A_QfBOhM2q5_2(.dout(w_dff_A_maRqugNU2_2),.din(w_dff_A_QfBOhM2q5_2),.clk(gclk));
	jdff dff_A_bSXExciB9_2(.dout(w_dff_A_QfBOhM2q5_2),.din(w_dff_A_bSXExciB9_2),.clk(gclk));
	jdff dff_B_mqNpbHV58_1(.din(n1638),.dout(w_dff_B_mqNpbHV58_1),.clk(gclk));
	jdff dff_A_yll1UEar9_1(.dout(w_n455_0[1]),.din(w_dff_A_yll1UEar9_1),.clk(gclk));
	jdff dff_A_YbD6cyVf2_1(.dout(w_dff_A_yll1UEar9_1),.din(w_dff_A_YbD6cyVf2_1),.clk(gclk));
	jdff dff_A_njaxN7py0_0(.dout(w_n461_0[0]),.din(w_dff_A_njaxN7py0_0),.clk(gclk));
	jdff dff_A_EZP3UGOg6_1(.dout(w_n460_0[1]),.din(w_dff_A_EZP3UGOg6_1),.clk(gclk));
	jdff dff_A_NexS8Rvc1_1(.dout(w_dff_A_EZP3UGOg6_1),.din(w_dff_A_NexS8Rvc1_1),.clk(gclk));
	jdff dff_A_jTTnyWji3_1(.dout(w_dff_A_NexS8Rvc1_1),.din(w_dff_A_jTTnyWji3_1),.clk(gclk));
	jdff dff_A_hPF8mIgd4_1(.dout(w_dff_A_jTTnyWji3_1),.din(w_dff_A_hPF8mIgd4_1),.clk(gclk));
	jdff dff_A_CwnsNRDR3_1(.dout(w_dff_A_hPF8mIgd4_1),.din(w_dff_A_CwnsNRDR3_1),.clk(gclk));
	jdff dff_A_4bpRI8ih8_1(.dout(w_n458_0[1]),.din(w_dff_A_4bpRI8ih8_1),.clk(gclk));
	jdff dff_A_lylUlSUn6_1(.dout(w_dff_A_4bpRI8ih8_1),.din(w_dff_A_lylUlSUn6_1),.clk(gclk));
	jdff dff_A_gUs6QCIy7_1(.dout(w_dff_A_lylUlSUn6_1),.din(w_dff_A_gUs6QCIy7_1),.clk(gclk));
	jdff dff_A_jlRhkfG69_1(.dout(w_dff_A_gUs6QCIy7_1),.din(w_dff_A_jlRhkfG69_1),.clk(gclk));
	jdff dff_A_5vcpByya4_1(.dout(w_dff_A_jlRhkfG69_1),.din(w_dff_A_5vcpByya4_1),.clk(gclk));
	jdff dff_A_ltp8zNyl2_1(.dout(w_dff_A_5vcpByya4_1),.din(w_dff_A_ltp8zNyl2_1),.clk(gclk));
	jdff dff_A_AnLtE6ts9_1(.dout(w_dff_A_ltp8zNyl2_1),.din(w_dff_A_AnLtE6ts9_1),.clk(gclk));
	jdff dff_A_jgZq5uJh2_0(.dout(w_G3729_1[0]),.din(w_dff_A_jgZq5uJh2_0),.clk(gclk));
	jdff dff_A_DtAQiGrm6_0(.dout(w_dff_A_jgZq5uJh2_0),.din(w_dff_A_DtAQiGrm6_0),.clk(gclk));
	jdff dff_A_jLgSfpG66_0(.dout(w_dff_A_DtAQiGrm6_0),.din(w_dff_A_jLgSfpG66_0),.clk(gclk));
	jdff dff_A_ReUw0QMK2_2(.dout(w_G3729_0[2]),.din(w_dff_A_ReUw0QMK2_2),.clk(gclk));
	jdff dff_A_s7wugzvr8_2(.dout(w_dff_A_ReUw0QMK2_2),.din(w_dff_A_s7wugzvr8_2),.clk(gclk));
	jdff dff_A_5XXE8IiG8_2(.dout(w_dff_A_s7wugzvr8_2),.din(w_dff_A_5XXE8IiG8_2),.clk(gclk));
	jdff dff_B_MBUHsfhs2_1(.din(n423),.dout(w_dff_B_MBUHsfhs2_1),.clk(gclk));
	jdff dff_B_VUCu99sn2_1(.din(w_dff_B_MBUHsfhs2_1),.dout(w_dff_B_VUCu99sn2_1),.clk(gclk));
	jdff dff_B_aj8GmS9T1_2(.din(n457),.dout(w_dff_B_aj8GmS9T1_2),.clk(gclk));
	jdff dff_A_3oBneEWV8_0(.dout(w_G18_55[0]),.din(w_dff_A_3oBneEWV8_0),.clk(gclk));
	jdff dff_A_xFyGdOtk0_2(.dout(w_G18_55[2]),.din(w_dff_A_xFyGdOtk0_2),.clk(gclk));
	jdff dff_A_FtdZB51Q5_0(.dout(w_G3737_1[0]),.din(w_dff_A_FtdZB51Q5_0),.clk(gclk));
	jdff dff_A_bh05FPEv9_0(.dout(w_dff_A_FtdZB51Q5_0),.din(w_dff_A_bh05FPEv9_0),.clk(gclk));
	jdff dff_A_xMIJMFxM8_0(.dout(w_dff_A_bh05FPEv9_0),.din(w_dff_A_xMIJMFxM8_0),.clk(gclk));
	jdff dff_A_mg9fQe3p8_1(.dout(w_n456_0[1]),.din(w_dff_A_mg9fQe3p8_1),.clk(gclk));
	jdff dff_A_AywLlYws1_1(.dout(w_dff_A_mg9fQe3p8_1),.din(w_dff_A_AywLlYws1_1),.clk(gclk));
	jdff dff_A_7DviQrrN0_1(.dout(w_dff_A_AywLlYws1_1),.din(w_dff_A_7DviQrrN0_1),.clk(gclk));
	jdff dff_A_e4k50gv77_1(.dout(w_dff_A_7DviQrrN0_1),.din(w_dff_A_e4k50gv77_1),.clk(gclk));
	jdff dff_A_6tXVjXax1_1(.dout(w_dff_A_e4k50gv77_1),.din(w_dff_A_6tXVjXax1_1),.clk(gclk));
	jdff dff_A_eqJec2Nj5_1(.dout(w_dff_A_6tXVjXax1_1),.din(w_dff_A_eqJec2Nj5_1),.clk(gclk));
	jdff dff_A_TE0SQFFm2_2(.dout(w_n456_0[2]),.din(w_dff_A_TE0SQFFm2_2),.clk(gclk));
	jdff dff_A_sLLTmDtc5_2(.dout(w_n446_0[2]),.din(w_dff_A_sLLTmDtc5_2),.clk(gclk));
	jdff dff_A_oO3tLiTK8_2(.dout(w_dff_A_sLLTmDtc5_2),.din(w_dff_A_oO3tLiTK8_2),.clk(gclk));
	jdff dff_A_DD47hUac5_2(.dout(w_dff_A_oO3tLiTK8_2),.din(w_dff_A_DD47hUac5_2),.clk(gclk));
	jdff dff_A_mQdCxS0s9_0(.dout(w_n445_0[0]),.din(w_dff_A_mQdCxS0s9_0),.clk(gclk));
	jdff dff_A_EP7Qe2SJ0_0(.dout(w_dff_A_mQdCxS0s9_0),.din(w_dff_A_EP7Qe2SJ0_0),.clk(gclk));
	jdff dff_A_u9uvz5bD2_0(.dout(w_dff_A_EP7Qe2SJ0_0),.din(w_dff_A_u9uvz5bD2_0),.clk(gclk));
	jdff dff_A_ISnzp72h4_0(.dout(w_dff_A_u9uvz5bD2_0),.din(w_dff_A_ISnzp72h4_0),.clk(gclk));
	jdff dff_B_TuWjnrE81_2(.din(n445),.dout(w_dff_B_TuWjnrE81_2),.clk(gclk));
	jdff dff_A_DSMDT6GG3_0(.dout(w_n443_0[0]),.din(w_dff_A_DSMDT6GG3_0),.clk(gclk));
	jdff dff_A_KB3kCZ4T9_0(.dout(w_dff_A_DSMDT6GG3_0),.din(w_dff_A_KB3kCZ4T9_0),.clk(gclk));
	jdff dff_A_iJ9qPTqX3_0(.dout(w_dff_A_KB3kCZ4T9_0),.din(w_dff_A_iJ9qPTqX3_0),.clk(gclk));
	jdff dff_A_JseIA2988_0(.dout(w_dff_A_iJ9qPTqX3_0),.din(w_dff_A_JseIA2988_0),.clk(gclk));
	jdff dff_A_Ru4qcSYj5_1(.dout(w_G18_54[1]),.din(w_dff_A_Ru4qcSYj5_1),.clk(gclk));
	jdff dff_A_WCVjazkL5_0(.dout(w_G3749_0[0]),.din(w_dff_A_WCVjazkL5_0),.clk(gclk));
	jdff dff_A_89rg4po88_0(.dout(w_dff_A_WCVjazkL5_0),.din(w_dff_A_89rg4po88_0),.clk(gclk));
	jdff dff_A_4esZn9dF8_0(.dout(w_dff_A_89rg4po88_0),.din(w_dff_A_4esZn9dF8_0),.clk(gclk));
	jdff dff_A_bOu4PHaO3_1(.dout(w_n450_0[1]),.din(w_dff_A_bOu4PHaO3_1),.clk(gclk));
	jdff dff_A_CC5J1EOU6_1(.dout(w_dff_A_bOu4PHaO3_1),.din(w_dff_A_CC5J1EOU6_1),.clk(gclk));
	jdff dff_A_A0qf5rob6_1(.dout(w_dff_A_CC5J1EOU6_1),.din(w_dff_A_A0qf5rob6_1),.clk(gclk));
	jdff dff_A_frdadZpM8_1(.dout(w_dff_A_A0qf5rob6_1),.din(w_dff_A_frdadZpM8_1),.clk(gclk));
	jdff dff_A_tbWG8swD2_1(.dout(w_dff_A_frdadZpM8_1),.din(w_dff_A_tbWG8swD2_1),.clk(gclk));
	jdff dff_A_TDUxJksk1_1(.dout(w_dff_A_tbWG8swD2_1),.din(w_dff_A_TDUxJksk1_1),.clk(gclk));
	jdff dff_A_7ComxtNr4_1(.dout(w_dff_A_TDUxJksk1_1),.din(w_dff_A_7ComxtNr4_1),.clk(gclk));
	jdff dff_A_WGXE9GoW3_2(.dout(w_n450_0[2]),.din(w_dff_A_WGXE9GoW3_2),.clk(gclk));
	jdff dff_B_xKIuOT5q4_3(.din(n450),.dout(w_dff_B_xKIuOT5q4_3),.clk(gclk));
	jdff dff_B_GRmSurMV5_1(.din(n447),.dout(w_dff_B_GRmSurMV5_1),.clk(gclk));
	jdff dff_B_Xj2Too0S0_0(.din(G124),.dout(w_dff_B_Xj2Too0S0_0),.clk(gclk));
	jdff dff_A_aOnlIr1H2_2(.dout(w_G18_58[2]),.din(w_dff_A_aOnlIr1H2_2),.clk(gclk));
	jdff dff_A_fK8Tqv5j2_1(.dout(w_G18_6[1]),.din(w_dff_A_fK8Tqv5j2_1),.clk(gclk));
	jdff dff_A_3OVEMHkP7_2(.dout(w_G18_6[2]),.din(w_dff_A_3OVEMHkP7_2),.clk(gclk));
	jdff dff_A_FieKRVQY5_2(.dout(w_G18_53[2]),.din(w_dff_A_FieKRVQY5_2),.clk(gclk));
	jdff dff_A_InQBo1k44_0(.dout(w_G3743_1[0]),.din(w_dff_A_InQBo1k44_0),.clk(gclk));
	jdff dff_A_BeMhbzOL0_1(.dout(w_G3743_1[1]),.din(w_dff_A_BeMhbzOL0_1),.clk(gclk));
	jdff dff_A_kgFhyGZ54_0(.dout(w_G3743_0[0]),.din(w_dff_A_kgFhyGZ54_0),.clk(gclk));
	jdff dff_A_d6LidJjF0_0(.dout(w_dff_A_kgFhyGZ54_0),.din(w_dff_A_d6LidJjF0_0),.clk(gclk));
	jdff dff_A_MoLiEjan8_0(.dout(w_dff_A_d6LidJjF0_0),.din(w_dff_A_MoLiEjan8_0),.clk(gclk));
	jdff dff_A_4tZotuGY6_1(.dout(w_n1360_0[1]),.din(w_dff_A_4tZotuGY6_1),.clk(gclk));
	jdff dff_A_1PLsBlBv4_2(.dout(w_n387_0[2]),.din(w_dff_A_1PLsBlBv4_2),.clk(gclk));
	jdff dff_A_bNf9o2zb6_2(.dout(w_dff_A_1PLsBlBv4_2),.din(w_dff_A_bNf9o2zb6_2),.clk(gclk));
	jdff dff_A_65MHYZTc6_2(.dout(w_dff_A_bNf9o2zb6_2),.din(w_dff_A_65MHYZTc6_2),.clk(gclk));
	jdff dff_A_HIATtF3z8_2(.dout(w_dff_A_65MHYZTc6_2),.din(w_dff_A_HIATtF3z8_2),.clk(gclk));
	jdff dff_B_VAc8eLdj7_1(.din(n381),.dout(w_dff_B_VAc8eLdj7_1),.clk(gclk));
	jdff dff_B_Q2fH6EwX9_1(.din(w_dff_B_VAc8eLdj7_1),.dout(w_dff_B_Q2fH6EwX9_1),.clk(gclk));
	jdff dff_A_VIfWgAQG6_0(.dout(w_G18_56[0]),.din(w_dff_A_VIfWgAQG6_0),.clk(gclk));
	jdff dff_A_Cblcpy8O5_2(.dout(w_G18_56[2]),.din(w_dff_A_Cblcpy8O5_2),.clk(gclk));
	jdff dff_A_NdfEdzRG9_0(.dout(w_G3711_1[0]),.din(w_dff_A_NdfEdzRG9_0),.clk(gclk));
	jdff dff_A_pD8Zds0M9_0(.dout(w_dff_A_NdfEdzRG9_0),.din(w_dff_A_pD8Zds0M9_0),.clk(gclk));
	jdff dff_A_W1sTOOLS3_0(.dout(w_dff_A_pD8Zds0M9_0),.din(w_dff_A_W1sTOOLS3_0),.clk(gclk));
	jdff dff_A_Jepw3d0D3_1(.dout(w_dff_A_zEiTH9Zm9_0),.din(w_dff_A_Jepw3d0D3_1),.clk(gclk));
	jdff dff_A_zEiTH9Zm9_0(.dout(w_dff_A_DaHyrcul0_0),.din(w_dff_A_zEiTH9Zm9_0),.clk(gclk));
	jdff dff_A_DaHyrcul0_0(.dout(w_dff_A_0iKJLw0g1_0),.din(w_dff_A_DaHyrcul0_0),.clk(gclk));
	jdff dff_A_0iKJLw0g1_0(.dout(w_dff_A_AV6wUJgT5_0),.din(w_dff_A_0iKJLw0g1_0),.clk(gclk));
	jdff dff_A_AV6wUJgT5_0(.dout(w_dff_A_sRT22TuU9_0),.din(w_dff_A_AV6wUJgT5_0),.clk(gclk));
	jdff dff_A_sRT22TuU9_0(.dout(w_dff_A_Dy8rk1pJ4_0),.din(w_dff_A_sRT22TuU9_0),.clk(gclk));
	jdff dff_A_Dy8rk1pJ4_0(.dout(w_dff_A_6s52Yf0B8_0),.din(w_dff_A_Dy8rk1pJ4_0),.clk(gclk));
	jdff dff_A_6s52Yf0B8_0(.dout(w_dff_A_uQ130t9g2_0),.din(w_dff_A_6s52Yf0B8_0),.clk(gclk));
	jdff dff_A_uQ130t9g2_0(.dout(w_dff_A_TAJP4QAD4_0),.din(w_dff_A_uQ130t9g2_0),.clk(gclk));
	jdff dff_A_TAJP4QAD4_0(.dout(w_dff_A_O20LuOqV8_0),.din(w_dff_A_TAJP4QAD4_0),.clk(gclk));
	jdff dff_A_O20LuOqV8_0(.dout(w_dff_A_bXAFYU1j4_0),.din(w_dff_A_O20LuOqV8_0),.clk(gclk));
	jdff dff_A_bXAFYU1j4_0(.dout(w_dff_A_neZh8IbH5_0),.din(w_dff_A_bXAFYU1j4_0),.clk(gclk));
	jdff dff_A_neZh8IbH5_0(.dout(w_dff_A_JVLOdUQK4_0),.din(w_dff_A_neZh8IbH5_0),.clk(gclk));
	jdff dff_A_JVLOdUQK4_0(.dout(w_dff_A_hUbSJeN43_0),.din(w_dff_A_JVLOdUQK4_0),.clk(gclk));
	jdff dff_A_hUbSJeN43_0(.dout(w_dff_A_403s3Cp35_0),.din(w_dff_A_hUbSJeN43_0),.clk(gclk));
	jdff dff_A_403s3Cp35_0(.dout(w_dff_A_VUTjnMhO5_0),.din(w_dff_A_403s3Cp35_0),.clk(gclk));
	jdff dff_A_VUTjnMhO5_0(.dout(w_dff_A_jilfT6S19_0),.din(w_dff_A_VUTjnMhO5_0),.clk(gclk));
	jdff dff_A_jilfT6S19_0(.dout(w_dff_A_eWWRG6EK1_0),.din(w_dff_A_jilfT6S19_0),.clk(gclk));
	jdff dff_A_eWWRG6EK1_0(.dout(w_dff_A_fi0SRwT30_0),.din(w_dff_A_eWWRG6EK1_0),.clk(gclk));
	jdff dff_A_fi0SRwT30_0(.dout(w_dff_A_qgtoXBKW1_0),.din(w_dff_A_fi0SRwT30_0),.clk(gclk));
	jdff dff_A_qgtoXBKW1_0(.dout(w_dff_A_EhaEvVca8_0),.din(w_dff_A_qgtoXBKW1_0),.clk(gclk));
	jdff dff_A_EhaEvVca8_0(.dout(w_dff_A_BdMyEXeo0_0),.din(w_dff_A_EhaEvVca8_0),.clk(gclk));
	jdff dff_A_BdMyEXeo0_0(.dout(w_dff_A_wJ2uW7JW4_0),.din(w_dff_A_BdMyEXeo0_0),.clk(gclk));
	jdff dff_A_wJ2uW7JW4_0(.dout(w_dff_A_OtkEzkzU6_0),.din(w_dff_A_wJ2uW7JW4_0),.clk(gclk));
	jdff dff_A_OtkEzkzU6_0(.dout(w_dff_A_6grC1mMW8_0),.din(w_dff_A_OtkEzkzU6_0),.clk(gclk));
	jdff dff_A_6grC1mMW8_0(.dout(w_dff_A_03HxQqjA3_0),.din(w_dff_A_6grC1mMW8_0),.clk(gclk));
	jdff dff_A_03HxQqjA3_0(.dout(G2),.din(w_dff_A_03HxQqjA3_0),.clk(gclk));
	jdff dff_A_OVoNiMA70_1(.dout(w_dff_A_QciStLOZ8_0),.din(w_dff_A_OVoNiMA70_1),.clk(gclk));
	jdff dff_A_QciStLOZ8_0(.dout(w_dff_A_CwhGq5X68_0),.din(w_dff_A_QciStLOZ8_0),.clk(gclk));
	jdff dff_A_CwhGq5X68_0(.dout(w_dff_A_ZnbdIMLO8_0),.din(w_dff_A_CwhGq5X68_0),.clk(gclk));
	jdff dff_A_ZnbdIMLO8_0(.dout(w_dff_A_23Jebp907_0),.din(w_dff_A_ZnbdIMLO8_0),.clk(gclk));
	jdff dff_A_23Jebp907_0(.dout(w_dff_A_DgzauxaI8_0),.din(w_dff_A_23Jebp907_0),.clk(gclk));
	jdff dff_A_DgzauxaI8_0(.dout(w_dff_A_Ral94vLK9_0),.din(w_dff_A_DgzauxaI8_0),.clk(gclk));
	jdff dff_A_Ral94vLK9_0(.dout(w_dff_A_XtGDoldv8_0),.din(w_dff_A_Ral94vLK9_0),.clk(gclk));
	jdff dff_A_XtGDoldv8_0(.dout(w_dff_A_2iokJu8B2_0),.din(w_dff_A_XtGDoldv8_0),.clk(gclk));
	jdff dff_A_2iokJu8B2_0(.dout(w_dff_A_FnhgHlMu6_0),.din(w_dff_A_2iokJu8B2_0),.clk(gclk));
	jdff dff_A_FnhgHlMu6_0(.dout(w_dff_A_j8LcjXOq1_0),.din(w_dff_A_FnhgHlMu6_0),.clk(gclk));
	jdff dff_A_j8LcjXOq1_0(.dout(w_dff_A_38YiM4ev2_0),.din(w_dff_A_j8LcjXOq1_0),.clk(gclk));
	jdff dff_A_38YiM4ev2_0(.dout(w_dff_A_T9HddJap8_0),.din(w_dff_A_38YiM4ev2_0),.clk(gclk));
	jdff dff_A_T9HddJap8_0(.dout(w_dff_A_RR49LlaI2_0),.din(w_dff_A_T9HddJap8_0),.clk(gclk));
	jdff dff_A_RR49LlaI2_0(.dout(w_dff_A_eRjoXH4Y1_0),.din(w_dff_A_RR49LlaI2_0),.clk(gclk));
	jdff dff_A_eRjoXH4Y1_0(.dout(w_dff_A_t3w2MgIX5_0),.din(w_dff_A_eRjoXH4Y1_0),.clk(gclk));
	jdff dff_A_t3w2MgIX5_0(.dout(w_dff_A_c5tvgWyQ8_0),.din(w_dff_A_t3w2MgIX5_0),.clk(gclk));
	jdff dff_A_c5tvgWyQ8_0(.dout(w_dff_A_YaHKVIjQ4_0),.din(w_dff_A_c5tvgWyQ8_0),.clk(gclk));
	jdff dff_A_YaHKVIjQ4_0(.dout(w_dff_A_yT5GGK2q8_0),.din(w_dff_A_YaHKVIjQ4_0),.clk(gclk));
	jdff dff_A_yT5GGK2q8_0(.dout(w_dff_A_oFfxPMDC6_0),.din(w_dff_A_yT5GGK2q8_0),.clk(gclk));
	jdff dff_A_oFfxPMDC6_0(.dout(w_dff_A_eIDU1cto8_0),.din(w_dff_A_oFfxPMDC6_0),.clk(gclk));
	jdff dff_A_eIDU1cto8_0(.dout(w_dff_A_yerG3EhD5_0),.din(w_dff_A_eIDU1cto8_0),.clk(gclk));
	jdff dff_A_yerG3EhD5_0(.dout(w_dff_A_DNWumpAE1_0),.din(w_dff_A_yerG3EhD5_0),.clk(gclk));
	jdff dff_A_DNWumpAE1_0(.dout(w_dff_A_nn5bK9qR9_0),.din(w_dff_A_DNWumpAE1_0),.clk(gclk));
	jdff dff_A_nn5bK9qR9_0(.dout(w_dff_A_i56gBVxo8_0),.din(w_dff_A_nn5bK9qR9_0),.clk(gclk));
	jdff dff_A_i56gBVxo8_0(.dout(w_dff_A_0AfyUwUz9_0),.din(w_dff_A_i56gBVxo8_0),.clk(gclk));
	jdff dff_A_0AfyUwUz9_0(.dout(w_dff_A_eg1Qo7Sp4_0),.din(w_dff_A_0AfyUwUz9_0),.clk(gclk));
	jdff dff_A_eg1Qo7Sp4_0(.dout(G3),.din(w_dff_A_eg1Qo7Sp4_0),.clk(gclk));
	jdff dff_A_At8WbDNn7_1(.dout(w_dff_A_zQnPEr3a7_0),.din(w_dff_A_At8WbDNn7_1),.clk(gclk));
	jdff dff_A_zQnPEr3a7_0(.dout(w_dff_A_6SrnGdpF8_0),.din(w_dff_A_zQnPEr3a7_0),.clk(gclk));
	jdff dff_A_6SrnGdpF8_0(.dout(w_dff_A_mAfGAQ7J3_0),.din(w_dff_A_6SrnGdpF8_0),.clk(gclk));
	jdff dff_A_mAfGAQ7J3_0(.dout(w_dff_A_zqgWuKbR3_0),.din(w_dff_A_mAfGAQ7J3_0),.clk(gclk));
	jdff dff_A_zqgWuKbR3_0(.dout(w_dff_A_6sVYvNCF7_0),.din(w_dff_A_zqgWuKbR3_0),.clk(gclk));
	jdff dff_A_6sVYvNCF7_0(.dout(w_dff_A_J63G1yqV1_0),.din(w_dff_A_6sVYvNCF7_0),.clk(gclk));
	jdff dff_A_J63G1yqV1_0(.dout(w_dff_A_RL5973yj6_0),.din(w_dff_A_J63G1yqV1_0),.clk(gclk));
	jdff dff_A_RL5973yj6_0(.dout(w_dff_A_Il9fFpgK9_0),.din(w_dff_A_RL5973yj6_0),.clk(gclk));
	jdff dff_A_Il9fFpgK9_0(.dout(w_dff_A_EYtrwJv03_0),.din(w_dff_A_Il9fFpgK9_0),.clk(gclk));
	jdff dff_A_EYtrwJv03_0(.dout(w_dff_A_t1NbP4ef0_0),.din(w_dff_A_EYtrwJv03_0),.clk(gclk));
	jdff dff_A_t1NbP4ef0_0(.dout(w_dff_A_MDxGcarH7_0),.din(w_dff_A_t1NbP4ef0_0),.clk(gclk));
	jdff dff_A_MDxGcarH7_0(.dout(w_dff_A_QorPNhsu1_0),.din(w_dff_A_MDxGcarH7_0),.clk(gclk));
	jdff dff_A_QorPNhsu1_0(.dout(w_dff_A_y3qeqxKp2_0),.din(w_dff_A_QorPNhsu1_0),.clk(gclk));
	jdff dff_A_y3qeqxKp2_0(.dout(w_dff_A_hQytYnNU3_0),.din(w_dff_A_y3qeqxKp2_0),.clk(gclk));
	jdff dff_A_hQytYnNU3_0(.dout(w_dff_A_VoGp1lo68_0),.din(w_dff_A_hQytYnNU3_0),.clk(gclk));
	jdff dff_A_VoGp1lo68_0(.dout(w_dff_A_qoip3ETL9_0),.din(w_dff_A_VoGp1lo68_0),.clk(gclk));
	jdff dff_A_qoip3ETL9_0(.dout(w_dff_A_maDAORxL5_0),.din(w_dff_A_qoip3ETL9_0),.clk(gclk));
	jdff dff_A_maDAORxL5_0(.dout(w_dff_A_iDZZJ2Ol4_0),.din(w_dff_A_maDAORxL5_0),.clk(gclk));
	jdff dff_A_iDZZJ2Ol4_0(.dout(w_dff_A_gIY056G84_0),.din(w_dff_A_iDZZJ2Ol4_0),.clk(gclk));
	jdff dff_A_gIY056G84_0(.dout(w_dff_A_G8sE0S8J5_0),.din(w_dff_A_gIY056G84_0),.clk(gclk));
	jdff dff_A_G8sE0S8J5_0(.dout(w_dff_A_HFisGFMX4_0),.din(w_dff_A_G8sE0S8J5_0),.clk(gclk));
	jdff dff_A_HFisGFMX4_0(.dout(w_dff_A_6dIB8NHN8_0),.din(w_dff_A_HFisGFMX4_0),.clk(gclk));
	jdff dff_A_6dIB8NHN8_0(.dout(w_dff_A_vj91fIyb9_0),.din(w_dff_A_6dIB8NHN8_0),.clk(gclk));
	jdff dff_A_vj91fIyb9_0(.dout(w_dff_A_yW2bb9pu3_0),.din(w_dff_A_vj91fIyb9_0),.clk(gclk));
	jdff dff_A_yW2bb9pu3_0(.dout(w_dff_A_ka0RPZsU3_0),.din(w_dff_A_yW2bb9pu3_0),.clk(gclk));
	jdff dff_A_ka0RPZsU3_0(.dout(w_dff_A_j8j9jEo48_0),.din(w_dff_A_ka0RPZsU3_0),.clk(gclk));
	jdff dff_A_j8j9jEo48_0(.dout(G450),.din(w_dff_A_j8j9jEo48_0),.clk(gclk));
	jdff dff_A_gI7ydG0x6_1(.dout(w_dff_A_G4yDRt4f5_0),.din(w_dff_A_gI7ydG0x6_1),.clk(gclk));
	jdff dff_A_G4yDRt4f5_0(.dout(w_dff_A_k1B6fnLc5_0),.din(w_dff_A_G4yDRt4f5_0),.clk(gclk));
	jdff dff_A_k1B6fnLc5_0(.dout(w_dff_A_8WK0lKBh8_0),.din(w_dff_A_k1B6fnLc5_0),.clk(gclk));
	jdff dff_A_8WK0lKBh8_0(.dout(w_dff_A_9wZfpoQ30_0),.din(w_dff_A_8WK0lKBh8_0),.clk(gclk));
	jdff dff_A_9wZfpoQ30_0(.dout(w_dff_A_bH11QFBu1_0),.din(w_dff_A_9wZfpoQ30_0),.clk(gclk));
	jdff dff_A_bH11QFBu1_0(.dout(w_dff_A_lPuW7BpP8_0),.din(w_dff_A_bH11QFBu1_0),.clk(gclk));
	jdff dff_A_lPuW7BpP8_0(.dout(w_dff_A_vNVSKerB0_0),.din(w_dff_A_lPuW7BpP8_0),.clk(gclk));
	jdff dff_A_vNVSKerB0_0(.dout(w_dff_A_QIjBGaPL9_0),.din(w_dff_A_vNVSKerB0_0),.clk(gclk));
	jdff dff_A_QIjBGaPL9_0(.dout(w_dff_A_3gUMWUZQ5_0),.din(w_dff_A_QIjBGaPL9_0),.clk(gclk));
	jdff dff_A_3gUMWUZQ5_0(.dout(w_dff_A_z4SyoYGQ5_0),.din(w_dff_A_3gUMWUZQ5_0),.clk(gclk));
	jdff dff_A_z4SyoYGQ5_0(.dout(w_dff_A_jcbGwhXk7_0),.din(w_dff_A_z4SyoYGQ5_0),.clk(gclk));
	jdff dff_A_jcbGwhXk7_0(.dout(w_dff_A_SRkM66zP5_0),.din(w_dff_A_jcbGwhXk7_0),.clk(gclk));
	jdff dff_A_SRkM66zP5_0(.dout(w_dff_A_P5e56rgL0_0),.din(w_dff_A_SRkM66zP5_0),.clk(gclk));
	jdff dff_A_P5e56rgL0_0(.dout(w_dff_A_GJyUpxno1_0),.din(w_dff_A_P5e56rgL0_0),.clk(gclk));
	jdff dff_A_GJyUpxno1_0(.dout(w_dff_A_w2phcBaP4_0),.din(w_dff_A_GJyUpxno1_0),.clk(gclk));
	jdff dff_A_w2phcBaP4_0(.dout(w_dff_A_9udBX3An0_0),.din(w_dff_A_w2phcBaP4_0),.clk(gclk));
	jdff dff_A_9udBX3An0_0(.dout(w_dff_A_VaNwzoIP1_0),.din(w_dff_A_9udBX3An0_0),.clk(gclk));
	jdff dff_A_VaNwzoIP1_0(.dout(w_dff_A_xfKS2rmf2_0),.din(w_dff_A_VaNwzoIP1_0),.clk(gclk));
	jdff dff_A_xfKS2rmf2_0(.dout(w_dff_A_pj2PDQJZ5_0),.din(w_dff_A_xfKS2rmf2_0),.clk(gclk));
	jdff dff_A_pj2PDQJZ5_0(.dout(w_dff_A_5tLmyzuw0_0),.din(w_dff_A_pj2PDQJZ5_0),.clk(gclk));
	jdff dff_A_5tLmyzuw0_0(.dout(w_dff_A_S4xL5rtv1_0),.din(w_dff_A_5tLmyzuw0_0),.clk(gclk));
	jdff dff_A_S4xL5rtv1_0(.dout(w_dff_A_StaLl54y4_0),.din(w_dff_A_S4xL5rtv1_0),.clk(gclk));
	jdff dff_A_StaLl54y4_0(.dout(w_dff_A_5ZuSJLAl0_0),.din(w_dff_A_StaLl54y4_0),.clk(gclk));
	jdff dff_A_5ZuSJLAl0_0(.dout(w_dff_A_HaOa1EMT9_0),.din(w_dff_A_5ZuSJLAl0_0),.clk(gclk));
	jdff dff_A_HaOa1EMT9_0(.dout(w_dff_A_gJ1AdJRW5_0),.din(w_dff_A_HaOa1EMT9_0),.clk(gclk));
	jdff dff_A_gJ1AdJRW5_0(.dout(w_dff_A_mWcJ8sZC0_0),.din(w_dff_A_gJ1AdJRW5_0),.clk(gclk));
	jdff dff_A_mWcJ8sZC0_0(.dout(G448),.din(w_dff_A_mWcJ8sZC0_0),.clk(gclk));
	jdff dff_A_jVuSQxh25_1(.dout(w_dff_A_zUQEsvNU9_0),.din(w_dff_A_jVuSQxh25_1),.clk(gclk));
	jdff dff_A_zUQEsvNU9_0(.dout(w_dff_A_zl4mvXi31_0),.din(w_dff_A_zUQEsvNU9_0),.clk(gclk));
	jdff dff_A_zl4mvXi31_0(.dout(w_dff_A_2wNEygOh1_0),.din(w_dff_A_zl4mvXi31_0),.clk(gclk));
	jdff dff_A_2wNEygOh1_0(.dout(w_dff_A_0swNFLFA6_0),.din(w_dff_A_2wNEygOh1_0),.clk(gclk));
	jdff dff_A_0swNFLFA6_0(.dout(w_dff_A_NZAlXzUr8_0),.din(w_dff_A_0swNFLFA6_0),.clk(gclk));
	jdff dff_A_NZAlXzUr8_0(.dout(w_dff_A_NGGMxrWH5_0),.din(w_dff_A_NZAlXzUr8_0),.clk(gclk));
	jdff dff_A_NGGMxrWH5_0(.dout(w_dff_A_tvTmI1Tq3_0),.din(w_dff_A_NGGMxrWH5_0),.clk(gclk));
	jdff dff_A_tvTmI1Tq3_0(.dout(w_dff_A_Pd0J3bWB7_0),.din(w_dff_A_tvTmI1Tq3_0),.clk(gclk));
	jdff dff_A_Pd0J3bWB7_0(.dout(w_dff_A_evCZlh8E2_0),.din(w_dff_A_Pd0J3bWB7_0),.clk(gclk));
	jdff dff_A_evCZlh8E2_0(.dout(w_dff_A_nZMUM3jn7_0),.din(w_dff_A_evCZlh8E2_0),.clk(gclk));
	jdff dff_A_nZMUM3jn7_0(.dout(w_dff_A_Awu2sevJ3_0),.din(w_dff_A_nZMUM3jn7_0),.clk(gclk));
	jdff dff_A_Awu2sevJ3_0(.dout(w_dff_A_bKmoNKZj4_0),.din(w_dff_A_Awu2sevJ3_0),.clk(gclk));
	jdff dff_A_bKmoNKZj4_0(.dout(w_dff_A_y7o9PyG60_0),.din(w_dff_A_bKmoNKZj4_0),.clk(gclk));
	jdff dff_A_y7o9PyG60_0(.dout(w_dff_A_1nIWNPCK1_0),.din(w_dff_A_y7o9PyG60_0),.clk(gclk));
	jdff dff_A_1nIWNPCK1_0(.dout(w_dff_A_nwDPreT13_0),.din(w_dff_A_1nIWNPCK1_0),.clk(gclk));
	jdff dff_A_nwDPreT13_0(.dout(w_dff_A_vmRHQ5fn1_0),.din(w_dff_A_nwDPreT13_0),.clk(gclk));
	jdff dff_A_vmRHQ5fn1_0(.dout(w_dff_A_snynsPTN9_0),.din(w_dff_A_vmRHQ5fn1_0),.clk(gclk));
	jdff dff_A_snynsPTN9_0(.dout(w_dff_A_GTCf4Bjd8_0),.din(w_dff_A_snynsPTN9_0),.clk(gclk));
	jdff dff_A_GTCf4Bjd8_0(.dout(w_dff_A_PYfdSkSZ1_0),.din(w_dff_A_GTCf4Bjd8_0),.clk(gclk));
	jdff dff_A_PYfdSkSZ1_0(.dout(w_dff_A_EvvD1VHe5_0),.din(w_dff_A_PYfdSkSZ1_0),.clk(gclk));
	jdff dff_A_EvvD1VHe5_0(.dout(w_dff_A_ZxTN4VId9_0),.din(w_dff_A_EvvD1VHe5_0),.clk(gclk));
	jdff dff_A_ZxTN4VId9_0(.dout(w_dff_A_NKZUlvlm9_0),.din(w_dff_A_ZxTN4VId9_0),.clk(gclk));
	jdff dff_A_NKZUlvlm9_0(.dout(w_dff_A_1N6hAOFS7_0),.din(w_dff_A_NKZUlvlm9_0),.clk(gclk));
	jdff dff_A_1N6hAOFS7_0(.dout(w_dff_A_Iv6iHDMa5_0),.din(w_dff_A_1N6hAOFS7_0),.clk(gclk));
	jdff dff_A_Iv6iHDMa5_0(.dout(w_dff_A_Zk10VM4i3_0),.din(w_dff_A_Iv6iHDMa5_0),.clk(gclk));
	jdff dff_A_Zk10VM4i3_0(.dout(w_dff_A_V9vjuaoO2_0),.din(w_dff_A_Zk10VM4i3_0),.clk(gclk));
	jdff dff_A_V9vjuaoO2_0(.dout(G444),.din(w_dff_A_V9vjuaoO2_0),.clk(gclk));
	jdff dff_A_ACjOL8Hd5_1(.dout(w_dff_A_OsKPVMcV6_0),.din(w_dff_A_ACjOL8Hd5_1),.clk(gclk));
	jdff dff_A_OsKPVMcV6_0(.dout(w_dff_A_2gfKfQHW3_0),.din(w_dff_A_OsKPVMcV6_0),.clk(gclk));
	jdff dff_A_2gfKfQHW3_0(.dout(w_dff_A_eD6EWofz2_0),.din(w_dff_A_2gfKfQHW3_0),.clk(gclk));
	jdff dff_A_eD6EWofz2_0(.dout(w_dff_A_4VigFBum1_0),.din(w_dff_A_eD6EWofz2_0),.clk(gclk));
	jdff dff_A_4VigFBum1_0(.dout(w_dff_A_quPWRA4Z3_0),.din(w_dff_A_4VigFBum1_0),.clk(gclk));
	jdff dff_A_quPWRA4Z3_0(.dout(w_dff_A_JyuF0Syz4_0),.din(w_dff_A_quPWRA4Z3_0),.clk(gclk));
	jdff dff_A_JyuF0Syz4_0(.dout(w_dff_A_0AG89SoL6_0),.din(w_dff_A_JyuF0Syz4_0),.clk(gclk));
	jdff dff_A_0AG89SoL6_0(.dout(w_dff_A_Slb9vga44_0),.din(w_dff_A_0AG89SoL6_0),.clk(gclk));
	jdff dff_A_Slb9vga44_0(.dout(w_dff_A_nQA2QG915_0),.din(w_dff_A_Slb9vga44_0),.clk(gclk));
	jdff dff_A_nQA2QG915_0(.dout(w_dff_A_cAJ3BJeM4_0),.din(w_dff_A_nQA2QG915_0),.clk(gclk));
	jdff dff_A_cAJ3BJeM4_0(.dout(w_dff_A_tSEgBoEL6_0),.din(w_dff_A_cAJ3BJeM4_0),.clk(gclk));
	jdff dff_A_tSEgBoEL6_0(.dout(w_dff_A_lpBuYtKj5_0),.din(w_dff_A_tSEgBoEL6_0),.clk(gclk));
	jdff dff_A_lpBuYtKj5_0(.dout(w_dff_A_14wjCRfa1_0),.din(w_dff_A_lpBuYtKj5_0),.clk(gclk));
	jdff dff_A_14wjCRfa1_0(.dout(w_dff_A_eq92qN2f8_0),.din(w_dff_A_14wjCRfa1_0),.clk(gclk));
	jdff dff_A_eq92qN2f8_0(.dout(w_dff_A_GFc4KQPw7_0),.din(w_dff_A_eq92qN2f8_0),.clk(gclk));
	jdff dff_A_GFc4KQPw7_0(.dout(w_dff_A_FWZk4rll9_0),.din(w_dff_A_GFc4KQPw7_0),.clk(gclk));
	jdff dff_A_FWZk4rll9_0(.dout(w_dff_A_psqGVi775_0),.din(w_dff_A_FWZk4rll9_0),.clk(gclk));
	jdff dff_A_psqGVi775_0(.dout(w_dff_A_xplWFAFY2_0),.din(w_dff_A_psqGVi775_0),.clk(gclk));
	jdff dff_A_xplWFAFY2_0(.dout(w_dff_A_5CmrKyPA8_0),.din(w_dff_A_xplWFAFY2_0),.clk(gclk));
	jdff dff_A_5CmrKyPA8_0(.dout(w_dff_A_SNhernBQ0_0),.din(w_dff_A_5CmrKyPA8_0),.clk(gclk));
	jdff dff_A_SNhernBQ0_0(.dout(w_dff_A_aJnWPzrI3_0),.din(w_dff_A_SNhernBQ0_0),.clk(gclk));
	jdff dff_A_aJnWPzrI3_0(.dout(w_dff_A_PzMXKrYC4_0),.din(w_dff_A_aJnWPzrI3_0),.clk(gclk));
	jdff dff_A_PzMXKrYC4_0(.dout(w_dff_A_UVS6p7Ir9_0),.din(w_dff_A_PzMXKrYC4_0),.clk(gclk));
	jdff dff_A_UVS6p7Ir9_0(.dout(w_dff_A_wisXWKJy9_0),.din(w_dff_A_UVS6p7Ir9_0),.clk(gclk));
	jdff dff_A_wisXWKJy9_0(.dout(w_dff_A_1nExP96H4_0),.din(w_dff_A_wisXWKJy9_0),.clk(gclk));
	jdff dff_A_1nExP96H4_0(.dout(w_dff_A_hU3KpgwW4_0),.din(w_dff_A_1nExP96H4_0),.clk(gclk));
	jdff dff_A_hU3KpgwW4_0(.dout(G442),.din(w_dff_A_hU3KpgwW4_0),.clk(gclk));
	jdff dff_A_6cIJftIc7_1(.dout(w_dff_A_Lh6GAcnc6_0),.din(w_dff_A_6cIJftIc7_1),.clk(gclk));
	jdff dff_A_Lh6GAcnc6_0(.dout(w_dff_A_USVsrT7K7_0),.din(w_dff_A_Lh6GAcnc6_0),.clk(gclk));
	jdff dff_A_USVsrT7K7_0(.dout(w_dff_A_0sXoFXr06_0),.din(w_dff_A_USVsrT7K7_0),.clk(gclk));
	jdff dff_A_0sXoFXr06_0(.dout(w_dff_A_WN6L333g9_0),.din(w_dff_A_0sXoFXr06_0),.clk(gclk));
	jdff dff_A_WN6L333g9_0(.dout(w_dff_A_VPYzLF6A0_0),.din(w_dff_A_WN6L333g9_0),.clk(gclk));
	jdff dff_A_VPYzLF6A0_0(.dout(w_dff_A_mmpYzzaL2_0),.din(w_dff_A_VPYzLF6A0_0),.clk(gclk));
	jdff dff_A_mmpYzzaL2_0(.dout(w_dff_A_TgDvA8u84_0),.din(w_dff_A_mmpYzzaL2_0),.clk(gclk));
	jdff dff_A_TgDvA8u84_0(.dout(w_dff_A_vdyd8aUp2_0),.din(w_dff_A_TgDvA8u84_0),.clk(gclk));
	jdff dff_A_vdyd8aUp2_0(.dout(w_dff_A_cruvJj447_0),.din(w_dff_A_vdyd8aUp2_0),.clk(gclk));
	jdff dff_A_cruvJj447_0(.dout(w_dff_A_AYSMuxkX9_0),.din(w_dff_A_cruvJj447_0),.clk(gclk));
	jdff dff_A_AYSMuxkX9_0(.dout(w_dff_A_CVYaBjgn4_0),.din(w_dff_A_AYSMuxkX9_0),.clk(gclk));
	jdff dff_A_CVYaBjgn4_0(.dout(w_dff_A_VGC4STos7_0),.din(w_dff_A_CVYaBjgn4_0),.clk(gclk));
	jdff dff_A_VGC4STos7_0(.dout(w_dff_A_mapEkjdk6_0),.din(w_dff_A_VGC4STos7_0),.clk(gclk));
	jdff dff_A_mapEkjdk6_0(.dout(w_dff_A_jhhwobVe1_0),.din(w_dff_A_mapEkjdk6_0),.clk(gclk));
	jdff dff_A_jhhwobVe1_0(.dout(w_dff_A_sTbIxCxx5_0),.din(w_dff_A_jhhwobVe1_0),.clk(gclk));
	jdff dff_A_sTbIxCxx5_0(.dout(w_dff_A_BRZyLWxa4_0),.din(w_dff_A_sTbIxCxx5_0),.clk(gclk));
	jdff dff_A_BRZyLWxa4_0(.dout(w_dff_A_kGQb8RrU4_0),.din(w_dff_A_BRZyLWxa4_0),.clk(gclk));
	jdff dff_A_kGQb8RrU4_0(.dout(w_dff_A_hYViNUUV3_0),.din(w_dff_A_kGQb8RrU4_0),.clk(gclk));
	jdff dff_A_hYViNUUV3_0(.dout(w_dff_A_U8jzsR4N0_0),.din(w_dff_A_hYViNUUV3_0),.clk(gclk));
	jdff dff_A_U8jzsR4N0_0(.dout(w_dff_A_NqlRo4AM4_0),.din(w_dff_A_U8jzsR4N0_0),.clk(gclk));
	jdff dff_A_NqlRo4AM4_0(.dout(w_dff_A_0PrzMRwF7_0),.din(w_dff_A_NqlRo4AM4_0),.clk(gclk));
	jdff dff_A_0PrzMRwF7_0(.dout(w_dff_A_iX2JAqtC9_0),.din(w_dff_A_0PrzMRwF7_0),.clk(gclk));
	jdff dff_A_iX2JAqtC9_0(.dout(w_dff_A_vjOGv9ky3_0),.din(w_dff_A_iX2JAqtC9_0),.clk(gclk));
	jdff dff_A_vjOGv9ky3_0(.dout(w_dff_A_K8uS5mrL0_0),.din(w_dff_A_vjOGv9ky3_0),.clk(gclk));
	jdff dff_A_K8uS5mrL0_0(.dout(w_dff_A_nMzacDpw0_0),.din(w_dff_A_K8uS5mrL0_0),.clk(gclk));
	jdff dff_A_nMzacDpw0_0(.dout(w_dff_A_b2Azpo0M9_0),.din(w_dff_A_nMzacDpw0_0),.clk(gclk));
	jdff dff_A_b2Azpo0M9_0(.dout(G440),.din(w_dff_A_b2Azpo0M9_0),.clk(gclk));
	jdff dff_A_oLMHIQy68_1(.dout(w_dff_A_U2TGf1IM1_0),.din(w_dff_A_oLMHIQy68_1),.clk(gclk));
	jdff dff_A_U2TGf1IM1_0(.dout(w_dff_A_PVYwONKp7_0),.din(w_dff_A_U2TGf1IM1_0),.clk(gclk));
	jdff dff_A_PVYwONKp7_0(.dout(w_dff_A_DFrsNgQV8_0),.din(w_dff_A_PVYwONKp7_0),.clk(gclk));
	jdff dff_A_DFrsNgQV8_0(.dout(w_dff_A_rT2n1vbr7_0),.din(w_dff_A_DFrsNgQV8_0),.clk(gclk));
	jdff dff_A_rT2n1vbr7_0(.dout(w_dff_A_VzUZMQtS0_0),.din(w_dff_A_rT2n1vbr7_0),.clk(gclk));
	jdff dff_A_VzUZMQtS0_0(.dout(w_dff_A_2n1N2GAQ2_0),.din(w_dff_A_VzUZMQtS0_0),.clk(gclk));
	jdff dff_A_2n1N2GAQ2_0(.dout(w_dff_A_WzWsWerw1_0),.din(w_dff_A_2n1N2GAQ2_0),.clk(gclk));
	jdff dff_A_WzWsWerw1_0(.dout(w_dff_A_3mObb0Dn6_0),.din(w_dff_A_WzWsWerw1_0),.clk(gclk));
	jdff dff_A_3mObb0Dn6_0(.dout(w_dff_A_mCeZDr0O2_0),.din(w_dff_A_3mObb0Dn6_0),.clk(gclk));
	jdff dff_A_mCeZDr0O2_0(.dout(w_dff_A_9tUgrR6C3_0),.din(w_dff_A_mCeZDr0O2_0),.clk(gclk));
	jdff dff_A_9tUgrR6C3_0(.dout(w_dff_A_JYSKCyf58_0),.din(w_dff_A_9tUgrR6C3_0),.clk(gclk));
	jdff dff_A_JYSKCyf58_0(.dout(w_dff_A_7CgXu5O03_0),.din(w_dff_A_JYSKCyf58_0),.clk(gclk));
	jdff dff_A_7CgXu5O03_0(.dout(w_dff_A_LFZhklvn0_0),.din(w_dff_A_7CgXu5O03_0),.clk(gclk));
	jdff dff_A_LFZhklvn0_0(.dout(w_dff_A_HaQ5rRU27_0),.din(w_dff_A_LFZhklvn0_0),.clk(gclk));
	jdff dff_A_HaQ5rRU27_0(.dout(w_dff_A_9EfvHjjF8_0),.din(w_dff_A_HaQ5rRU27_0),.clk(gclk));
	jdff dff_A_9EfvHjjF8_0(.dout(w_dff_A_H6kECw7M1_0),.din(w_dff_A_9EfvHjjF8_0),.clk(gclk));
	jdff dff_A_H6kECw7M1_0(.dout(w_dff_A_MiApOLDo8_0),.din(w_dff_A_H6kECw7M1_0),.clk(gclk));
	jdff dff_A_MiApOLDo8_0(.dout(w_dff_A_EccW5sm02_0),.din(w_dff_A_MiApOLDo8_0),.clk(gclk));
	jdff dff_A_EccW5sm02_0(.dout(w_dff_A_QNCFt2GF6_0),.din(w_dff_A_EccW5sm02_0),.clk(gclk));
	jdff dff_A_QNCFt2GF6_0(.dout(w_dff_A_t0SZeUVc0_0),.din(w_dff_A_QNCFt2GF6_0),.clk(gclk));
	jdff dff_A_t0SZeUVc0_0(.dout(w_dff_A_ayYtbDTE4_0),.din(w_dff_A_t0SZeUVc0_0),.clk(gclk));
	jdff dff_A_ayYtbDTE4_0(.dout(w_dff_A_fLAGXdEm5_0),.din(w_dff_A_ayYtbDTE4_0),.clk(gclk));
	jdff dff_A_fLAGXdEm5_0(.dout(w_dff_A_W7KxjQ2U3_0),.din(w_dff_A_fLAGXdEm5_0),.clk(gclk));
	jdff dff_A_W7KxjQ2U3_0(.dout(w_dff_A_6GE3KT1J6_0),.din(w_dff_A_W7KxjQ2U3_0),.clk(gclk));
	jdff dff_A_6GE3KT1J6_0(.dout(w_dff_A_YuAapg5j7_0),.din(w_dff_A_6GE3KT1J6_0),.clk(gclk));
	jdff dff_A_YuAapg5j7_0(.dout(w_dff_A_NATs0cOt0_0),.din(w_dff_A_YuAapg5j7_0),.clk(gclk));
	jdff dff_A_NATs0cOt0_0(.dout(G438),.din(w_dff_A_NATs0cOt0_0),.clk(gclk));
	jdff dff_A_PH2dp2Gh6_1(.dout(w_dff_A_3uBwvu5V0_0),.din(w_dff_A_PH2dp2Gh6_1),.clk(gclk));
	jdff dff_A_3uBwvu5V0_0(.dout(w_dff_A_cay00hC52_0),.din(w_dff_A_3uBwvu5V0_0),.clk(gclk));
	jdff dff_A_cay00hC52_0(.dout(w_dff_A_UOFRSfUm6_0),.din(w_dff_A_cay00hC52_0),.clk(gclk));
	jdff dff_A_UOFRSfUm6_0(.dout(w_dff_A_YQq5HJFC9_0),.din(w_dff_A_UOFRSfUm6_0),.clk(gclk));
	jdff dff_A_YQq5HJFC9_0(.dout(w_dff_A_UF1V6TqY3_0),.din(w_dff_A_YQq5HJFC9_0),.clk(gclk));
	jdff dff_A_UF1V6TqY3_0(.dout(w_dff_A_eQLXca4z5_0),.din(w_dff_A_UF1V6TqY3_0),.clk(gclk));
	jdff dff_A_eQLXca4z5_0(.dout(w_dff_A_I4ooIf943_0),.din(w_dff_A_eQLXca4z5_0),.clk(gclk));
	jdff dff_A_I4ooIf943_0(.dout(w_dff_A_Lpth9xgc7_0),.din(w_dff_A_I4ooIf943_0),.clk(gclk));
	jdff dff_A_Lpth9xgc7_0(.dout(w_dff_A_irtSG1Av6_0),.din(w_dff_A_Lpth9xgc7_0),.clk(gclk));
	jdff dff_A_irtSG1Av6_0(.dout(w_dff_A_1FuVCvfx8_0),.din(w_dff_A_irtSG1Av6_0),.clk(gclk));
	jdff dff_A_1FuVCvfx8_0(.dout(w_dff_A_R7OBf5QS3_0),.din(w_dff_A_1FuVCvfx8_0),.clk(gclk));
	jdff dff_A_R7OBf5QS3_0(.dout(w_dff_A_52wq3IfU8_0),.din(w_dff_A_R7OBf5QS3_0),.clk(gclk));
	jdff dff_A_52wq3IfU8_0(.dout(w_dff_A_rA4OQhkI8_0),.din(w_dff_A_52wq3IfU8_0),.clk(gclk));
	jdff dff_A_rA4OQhkI8_0(.dout(w_dff_A_xgNM9Hm82_0),.din(w_dff_A_rA4OQhkI8_0),.clk(gclk));
	jdff dff_A_xgNM9Hm82_0(.dout(w_dff_A_1mFIJGt20_0),.din(w_dff_A_xgNM9Hm82_0),.clk(gclk));
	jdff dff_A_1mFIJGt20_0(.dout(w_dff_A_pV8d6myB8_0),.din(w_dff_A_1mFIJGt20_0),.clk(gclk));
	jdff dff_A_pV8d6myB8_0(.dout(w_dff_A_fkYSKB0U2_0),.din(w_dff_A_pV8d6myB8_0),.clk(gclk));
	jdff dff_A_fkYSKB0U2_0(.dout(w_dff_A_DBrXzvVZ9_0),.din(w_dff_A_fkYSKB0U2_0),.clk(gclk));
	jdff dff_A_DBrXzvVZ9_0(.dout(w_dff_A_ZYBwbVix6_0),.din(w_dff_A_DBrXzvVZ9_0),.clk(gclk));
	jdff dff_A_ZYBwbVix6_0(.dout(w_dff_A_KFSS2HHL3_0),.din(w_dff_A_ZYBwbVix6_0),.clk(gclk));
	jdff dff_A_KFSS2HHL3_0(.dout(w_dff_A_gC9Q4zzD6_0),.din(w_dff_A_KFSS2HHL3_0),.clk(gclk));
	jdff dff_A_gC9Q4zzD6_0(.dout(w_dff_A_vTmF3Vgi8_0),.din(w_dff_A_gC9Q4zzD6_0),.clk(gclk));
	jdff dff_A_vTmF3Vgi8_0(.dout(w_dff_A_1x3LKIsn4_0),.din(w_dff_A_vTmF3Vgi8_0),.clk(gclk));
	jdff dff_A_1x3LKIsn4_0(.dout(w_dff_A_Gq4r9SHf6_0),.din(w_dff_A_1x3LKIsn4_0),.clk(gclk));
	jdff dff_A_Gq4r9SHf6_0(.dout(w_dff_A_rp4WfyMj0_0),.din(w_dff_A_Gq4r9SHf6_0),.clk(gclk));
	jdff dff_A_rp4WfyMj0_0(.dout(w_dff_A_Kozqd2sm0_0),.din(w_dff_A_rp4WfyMj0_0),.clk(gclk));
	jdff dff_A_Kozqd2sm0_0(.dout(G496),.din(w_dff_A_Kozqd2sm0_0),.clk(gclk));
	jdff dff_A_ck3mftU05_1(.dout(w_dff_A_5QkZzppr9_0),.din(w_dff_A_ck3mftU05_1),.clk(gclk));
	jdff dff_A_5QkZzppr9_0(.dout(w_dff_A_4i9L9jy14_0),.din(w_dff_A_5QkZzppr9_0),.clk(gclk));
	jdff dff_A_4i9L9jy14_0(.dout(w_dff_A_FbNyRffT5_0),.din(w_dff_A_4i9L9jy14_0),.clk(gclk));
	jdff dff_A_FbNyRffT5_0(.dout(w_dff_A_9SyphRnW5_0),.din(w_dff_A_FbNyRffT5_0),.clk(gclk));
	jdff dff_A_9SyphRnW5_0(.dout(w_dff_A_rfqA71EW5_0),.din(w_dff_A_9SyphRnW5_0),.clk(gclk));
	jdff dff_A_rfqA71EW5_0(.dout(w_dff_A_IXqBEUwM7_0),.din(w_dff_A_rfqA71EW5_0),.clk(gclk));
	jdff dff_A_IXqBEUwM7_0(.dout(w_dff_A_uxkjaRNX6_0),.din(w_dff_A_IXqBEUwM7_0),.clk(gclk));
	jdff dff_A_uxkjaRNX6_0(.dout(w_dff_A_IZssx8BL3_0),.din(w_dff_A_uxkjaRNX6_0),.clk(gclk));
	jdff dff_A_IZssx8BL3_0(.dout(w_dff_A_q3JCjGgB5_0),.din(w_dff_A_IZssx8BL3_0),.clk(gclk));
	jdff dff_A_q3JCjGgB5_0(.dout(w_dff_A_fIVMpX423_0),.din(w_dff_A_q3JCjGgB5_0),.clk(gclk));
	jdff dff_A_fIVMpX423_0(.dout(w_dff_A_GA1ZIZGA0_0),.din(w_dff_A_fIVMpX423_0),.clk(gclk));
	jdff dff_A_GA1ZIZGA0_0(.dout(w_dff_A_MIwtfxl14_0),.din(w_dff_A_GA1ZIZGA0_0),.clk(gclk));
	jdff dff_A_MIwtfxl14_0(.dout(w_dff_A_OM3UJLKk1_0),.din(w_dff_A_MIwtfxl14_0),.clk(gclk));
	jdff dff_A_OM3UJLKk1_0(.dout(w_dff_A_t2oPecny4_0),.din(w_dff_A_OM3UJLKk1_0),.clk(gclk));
	jdff dff_A_t2oPecny4_0(.dout(w_dff_A_g1J0EXoi1_0),.din(w_dff_A_t2oPecny4_0),.clk(gclk));
	jdff dff_A_g1J0EXoi1_0(.dout(w_dff_A_HRSZ4uTR0_0),.din(w_dff_A_g1J0EXoi1_0),.clk(gclk));
	jdff dff_A_HRSZ4uTR0_0(.dout(w_dff_A_5RS1Sbyd9_0),.din(w_dff_A_HRSZ4uTR0_0),.clk(gclk));
	jdff dff_A_5RS1Sbyd9_0(.dout(w_dff_A_RH4rAyJb7_0),.din(w_dff_A_5RS1Sbyd9_0),.clk(gclk));
	jdff dff_A_RH4rAyJb7_0(.dout(w_dff_A_c5Xfhjm95_0),.din(w_dff_A_RH4rAyJb7_0),.clk(gclk));
	jdff dff_A_c5Xfhjm95_0(.dout(w_dff_A_mhSKdxut6_0),.din(w_dff_A_c5Xfhjm95_0),.clk(gclk));
	jdff dff_A_mhSKdxut6_0(.dout(w_dff_A_UtoDTZYn0_0),.din(w_dff_A_mhSKdxut6_0),.clk(gclk));
	jdff dff_A_UtoDTZYn0_0(.dout(w_dff_A_EjPZGGWJ3_0),.din(w_dff_A_UtoDTZYn0_0),.clk(gclk));
	jdff dff_A_EjPZGGWJ3_0(.dout(w_dff_A_2yHgo7sQ9_0),.din(w_dff_A_EjPZGGWJ3_0),.clk(gclk));
	jdff dff_A_2yHgo7sQ9_0(.dout(w_dff_A_aNaLIc3A8_0),.din(w_dff_A_2yHgo7sQ9_0),.clk(gclk));
	jdff dff_A_aNaLIc3A8_0(.dout(w_dff_A_WNdDMffj4_0),.din(w_dff_A_aNaLIc3A8_0),.clk(gclk));
	jdff dff_A_WNdDMffj4_0(.dout(w_dff_A_9Te3iLBO1_0),.din(w_dff_A_WNdDMffj4_0),.clk(gclk));
	jdff dff_A_9Te3iLBO1_0(.dout(G494),.din(w_dff_A_9Te3iLBO1_0),.clk(gclk));
	jdff dff_A_vip4ZzAz3_1(.dout(w_dff_A_AV4YQpCp2_0),.din(w_dff_A_vip4ZzAz3_1),.clk(gclk));
	jdff dff_A_AV4YQpCp2_0(.dout(w_dff_A_h8xZlgyj0_0),.din(w_dff_A_AV4YQpCp2_0),.clk(gclk));
	jdff dff_A_h8xZlgyj0_0(.dout(w_dff_A_58AbwFuW7_0),.din(w_dff_A_h8xZlgyj0_0),.clk(gclk));
	jdff dff_A_58AbwFuW7_0(.dout(w_dff_A_hcYwSQ2s7_0),.din(w_dff_A_58AbwFuW7_0),.clk(gclk));
	jdff dff_A_hcYwSQ2s7_0(.dout(w_dff_A_yonyJIBb3_0),.din(w_dff_A_hcYwSQ2s7_0),.clk(gclk));
	jdff dff_A_yonyJIBb3_0(.dout(w_dff_A_VCdq4rgj6_0),.din(w_dff_A_yonyJIBb3_0),.clk(gclk));
	jdff dff_A_VCdq4rgj6_0(.dout(w_dff_A_OJNR7WCi4_0),.din(w_dff_A_VCdq4rgj6_0),.clk(gclk));
	jdff dff_A_OJNR7WCi4_0(.dout(w_dff_A_BKl1XY1o9_0),.din(w_dff_A_OJNR7WCi4_0),.clk(gclk));
	jdff dff_A_BKl1XY1o9_0(.dout(w_dff_A_gaQh5O730_0),.din(w_dff_A_BKl1XY1o9_0),.clk(gclk));
	jdff dff_A_gaQh5O730_0(.dout(w_dff_A_X7Q2Wy8J1_0),.din(w_dff_A_gaQh5O730_0),.clk(gclk));
	jdff dff_A_X7Q2Wy8J1_0(.dout(w_dff_A_bSupoS2p8_0),.din(w_dff_A_X7Q2Wy8J1_0),.clk(gclk));
	jdff dff_A_bSupoS2p8_0(.dout(w_dff_A_5V6VCIyV1_0),.din(w_dff_A_bSupoS2p8_0),.clk(gclk));
	jdff dff_A_5V6VCIyV1_0(.dout(w_dff_A_uWqHp8hr0_0),.din(w_dff_A_5V6VCIyV1_0),.clk(gclk));
	jdff dff_A_uWqHp8hr0_0(.dout(w_dff_A_9bOX0rlD9_0),.din(w_dff_A_uWqHp8hr0_0),.clk(gclk));
	jdff dff_A_9bOX0rlD9_0(.dout(w_dff_A_WNVCM9Z43_0),.din(w_dff_A_9bOX0rlD9_0),.clk(gclk));
	jdff dff_A_WNVCM9Z43_0(.dout(w_dff_A_0L5yOjg40_0),.din(w_dff_A_WNVCM9Z43_0),.clk(gclk));
	jdff dff_A_0L5yOjg40_0(.dout(w_dff_A_qStqOnBr0_0),.din(w_dff_A_0L5yOjg40_0),.clk(gclk));
	jdff dff_A_qStqOnBr0_0(.dout(w_dff_A_Jis98WqO4_0),.din(w_dff_A_qStqOnBr0_0),.clk(gclk));
	jdff dff_A_Jis98WqO4_0(.dout(w_dff_A_GHrDsJGs6_0),.din(w_dff_A_Jis98WqO4_0),.clk(gclk));
	jdff dff_A_GHrDsJGs6_0(.dout(w_dff_A_8xhs9iWv1_0),.din(w_dff_A_GHrDsJGs6_0),.clk(gclk));
	jdff dff_A_8xhs9iWv1_0(.dout(w_dff_A_lemmLzko6_0),.din(w_dff_A_8xhs9iWv1_0),.clk(gclk));
	jdff dff_A_lemmLzko6_0(.dout(w_dff_A_3A3nZ2Ff8_0),.din(w_dff_A_lemmLzko6_0),.clk(gclk));
	jdff dff_A_3A3nZ2Ff8_0(.dout(w_dff_A_gLgzK0w67_0),.din(w_dff_A_3A3nZ2Ff8_0),.clk(gclk));
	jdff dff_A_gLgzK0w67_0(.dout(w_dff_A_cNZYIumD6_0),.din(w_dff_A_gLgzK0w67_0),.clk(gclk));
	jdff dff_A_cNZYIumD6_0(.dout(w_dff_A_gasweF2w8_0),.din(w_dff_A_cNZYIumD6_0),.clk(gclk));
	jdff dff_A_gasweF2w8_0(.dout(w_dff_A_7WSSQWkS9_0),.din(w_dff_A_gasweF2w8_0),.clk(gclk));
	jdff dff_A_7WSSQWkS9_0(.dout(G492),.din(w_dff_A_7WSSQWkS9_0),.clk(gclk));
	jdff dff_A_jyfYMINM3_1(.dout(w_dff_A_eI5d90CH7_0),.din(w_dff_A_jyfYMINM3_1),.clk(gclk));
	jdff dff_A_eI5d90CH7_0(.dout(w_dff_A_dm5rUY5J0_0),.din(w_dff_A_eI5d90CH7_0),.clk(gclk));
	jdff dff_A_dm5rUY5J0_0(.dout(w_dff_A_5U3jWzoV9_0),.din(w_dff_A_dm5rUY5J0_0),.clk(gclk));
	jdff dff_A_5U3jWzoV9_0(.dout(w_dff_A_xG5t2Viz6_0),.din(w_dff_A_5U3jWzoV9_0),.clk(gclk));
	jdff dff_A_xG5t2Viz6_0(.dout(w_dff_A_564LMFfM6_0),.din(w_dff_A_xG5t2Viz6_0),.clk(gclk));
	jdff dff_A_564LMFfM6_0(.dout(w_dff_A_93efPrR40_0),.din(w_dff_A_564LMFfM6_0),.clk(gclk));
	jdff dff_A_93efPrR40_0(.dout(w_dff_A_3QCK2Y0q2_0),.din(w_dff_A_93efPrR40_0),.clk(gclk));
	jdff dff_A_3QCK2Y0q2_0(.dout(w_dff_A_9cSxeKhO9_0),.din(w_dff_A_3QCK2Y0q2_0),.clk(gclk));
	jdff dff_A_9cSxeKhO9_0(.dout(w_dff_A_5MRGyAFT1_0),.din(w_dff_A_9cSxeKhO9_0),.clk(gclk));
	jdff dff_A_5MRGyAFT1_0(.dout(w_dff_A_PGLlR02d9_0),.din(w_dff_A_5MRGyAFT1_0),.clk(gclk));
	jdff dff_A_PGLlR02d9_0(.dout(w_dff_A_FtOHGXm27_0),.din(w_dff_A_PGLlR02d9_0),.clk(gclk));
	jdff dff_A_FtOHGXm27_0(.dout(w_dff_A_AbNKHRsZ8_0),.din(w_dff_A_FtOHGXm27_0),.clk(gclk));
	jdff dff_A_AbNKHRsZ8_0(.dout(w_dff_A_aUwouS491_0),.din(w_dff_A_AbNKHRsZ8_0),.clk(gclk));
	jdff dff_A_aUwouS491_0(.dout(w_dff_A_scwVVDns8_0),.din(w_dff_A_aUwouS491_0),.clk(gclk));
	jdff dff_A_scwVVDns8_0(.dout(w_dff_A_1MRHAMBf8_0),.din(w_dff_A_scwVVDns8_0),.clk(gclk));
	jdff dff_A_1MRHAMBf8_0(.dout(w_dff_A_c6VPGdOW4_0),.din(w_dff_A_1MRHAMBf8_0),.clk(gclk));
	jdff dff_A_c6VPGdOW4_0(.dout(w_dff_A_ahB1yBrd7_0),.din(w_dff_A_c6VPGdOW4_0),.clk(gclk));
	jdff dff_A_ahB1yBrd7_0(.dout(w_dff_A_PAOHaUL88_0),.din(w_dff_A_ahB1yBrd7_0),.clk(gclk));
	jdff dff_A_PAOHaUL88_0(.dout(w_dff_A_hQpXWMcN8_0),.din(w_dff_A_PAOHaUL88_0),.clk(gclk));
	jdff dff_A_hQpXWMcN8_0(.dout(w_dff_A_4v2CthqX5_0),.din(w_dff_A_hQpXWMcN8_0),.clk(gclk));
	jdff dff_A_4v2CthqX5_0(.dout(w_dff_A_T08au5NZ9_0),.din(w_dff_A_4v2CthqX5_0),.clk(gclk));
	jdff dff_A_T08au5NZ9_0(.dout(w_dff_A_yJT368vh5_0),.din(w_dff_A_T08au5NZ9_0),.clk(gclk));
	jdff dff_A_yJT368vh5_0(.dout(w_dff_A_P08PhQeu8_0),.din(w_dff_A_yJT368vh5_0),.clk(gclk));
	jdff dff_A_P08PhQeu8_0(.dout(w_dff_A_uisEK8NY1_0),.din(w_dff_A_P08PhQeu8_0),.clk(gclk));
	jdff dff_A_uisEK8NY1_0(.dout(w_dff_A_2YzGgPL20_0),.din(w_dff_A_uisEK8NY1_0),.clk(gclk));
	jdff dff_A_2YzGgPL20_0(.dout(w_dff_A_8HtwiNIy5_0),.din(w_dff_A_2YzGgPL20_0),.clk(gclk));
	jdff dff_A_8HtwiNIy5_0(.dout(G490),.din(w_dff_A_8HtwiNIy5_0),.clk(gclk));
	jdff dff_A_M7WkONvQ8_1(.dout(w_dff_A_cyPCU36U8_0),.din(w_dff_A_M7WkONvQ8_1),.clk(gclk));
	jdff dff_A_cyPCU36U8_0(.dout(w_dff_A_suqT5l4x3_0),.din(w_dff_A_cyPCU36U8_0),.clk(gclk));
	jdff dff_A_suqT5l4x3_0(.dout(w_dff_A_6xfY8LbF6_0),.din(w_dff_A_suqT5l4x3_0),.clk(gclk));
	jdff dff_A_6xfY8LbF6_0(.dout(w_dff_A_uPLLNTll7_0),.din(w_dff_A_6xfY8LbF6_0),.clk(gclk));
	jdff dff_A_uPLLNTll7_0(.dout(w_dff_A_l8lB22ox4_0),.din(w_dff_A_uPLLNTll7_0),.clk(gclk));
	jdff dff_A_l8lB22ox4_0(.dout(w_dff_A_DlZXrZS05_0),.din(w_dff_A_l8lB22ox4_0),.clk(gclk));
	jdff dff_A_DlZXrZS05_0(.dout(w_dff_A_dJTLvTv41_0),.din(w_dff_A_DlZXrZS05_0),.clk(gclk));
	jdff dff_A_dJTLvTv41_0(.dout(w_dff_A_POqfTGWV1_0),.din(w_dff_A_dJTLvTv41_0),.clk(gclk));
	jdff dff_A_POqfTGWV1_0(.dout(w_dff_A_ZooAC3JN4_0),.din(w_dff_A_POqfTGWV1_0),.clk(gclk));
	jdff dff_A_ZooAC3JN4_0(.dout(w_dff_A_RAT5AKzx5_0),.din(w_dff_A_ZooAC3JN4_0),.clk(gclk));
	jdff dff_A_RAT5AKzx5_0(.dout(w_dff_A_zk4foa114_0),.din(w_dff_A_RAT5AKzx5_0),.clk(gclk));
	jdff dff_A_zk4foa114_0(.dout(w_dff_A_OXYE1hiF0_0),.din(w_dff_A_zk4foa114_0),.clk(gclk));
	jdff dff_A_OXYE1hiF0_0(.dout(w_dff_A_7AQkkkbb8_0),.din(w_dff_A_OXYE1hiF0_0),.clk(gclk));
	jdff dff_A_7AQkkkbb8_0(.dout(w_dff_A_vgw4zCMV6_0),.din(w_dff_A_7AQkkkbb8_0),.clk(gclk));
	jdff dff_A_vgw4zCMV6_0(.dout(w_dff_A_tJ8UBXPL4_0),.din(w_dff_A_vgw4zCMV6_0),.clk(gclk));
	jdff dff_A_tJ8UBXPL4_0(.dout(w_dff_A_m9pQ2itu2_0),.din(w_dff_A_tJ8UBXPL4_0),.clk(gclk));
	jdff dff_A_m9pQ2itu2_0(.dout(w_dff_A_Od6sMVbx0_0),.din(w_dff_A_m9pQ2itu2_0),.clk(gclk));
	jdff dff_A_Od6sMVbx0_0(.dout(w_dff_A_USI4Smfu5_0),.din(w_dff_A_Od6sMVbx0_0),.clk(gclk));
	jdff dff_A_USI4Smfu5_0(.dout(w_dff_A_enYjavb83_0),.din(w_dff_A_USI4Smfu5_0),.clk(gclk));
	jdff dff_A_enYjavb83_0(.dout(w_dff_A_458wZoyV6_0),.din(w_dff_A_enYjavb83_0),.clk(gclk));
	jdff dff_A_458wZoyV6_0(.dout(w_dff_A_rrKHGKDr5_0),.din(w_dff_A_458wZoyV6_0),.clk(gclk));
	jdff dff_A_rrKHGKDr5_0(.dout(w_dff_A_9ONo0ROf7_0),.din(w_dff_A_rrKHGKDr5_0),.clk(gclk));
	jdff dff_A_9ONo0ROf7_0(.dout(w_dff_A_aSa4X3sQ4_0),.din(w_dff_A_9ONo0ROf7_0),.clk(gclk));
	jdff dff_A_aSa4X3sQ4_0(.dout(w_dff_A_PtmdTOeI8_0),.din(w_dff_A_aSa4X3sQ4_0),.clk(gclk));
	jdff dff_A_PtmdTOeI8_0(.dout(w_dff_A_JsNmkiST9_0),.din(w_dff_A_PtmdTOeI8_0),.clk(gclk));
	jdff dff_A_JsNmkiST9_0(.dout(w_dff_A_GTd40T6T8_0),.din(w_dff_A_JsNmkiST9_0),.clk(gclk));
	jdff dff_A_GTd40T6T8_0(.dout(G488),.din(w_dff_A_GTd40T6T8_0),.clk(gclk));
	jdff dff_A_e0o8y8if7_1(.dout(w_dff_A_Cd4p4fpU6_0),.din(w_dff_A_e0o8y8if7_1),.clk(gclk));
	jdff dff_A_Cd4p4fpU6_0(.dout(w_dff_A_2nhgyW6M1_0),.din(w_dff_A_Cd4p4fpU6_0),.clk(gclk));
	jdff dff_A_2nhgyW6M1_0(.dout(w_dff_A_nvtOrw3v2_0),.din(w_dff_A_2nhgyW6M1_0),.clk(gclk));
	jdff dff_A_nvtOrw3v2_0(.dout(w_dff_A_qsf2dGYj5_0),.din(w_dff_A_nvtOrw3v2_0),.clk(gclk));
	jdff dff_A_qsf2dGYj5_0(.dout(w_dff_A_riVGJaof1_0),.din(w_dff_A_qsf2dGYj5_0),.clk(gclk));
	jdff dff_A_riVGJaof1_0(.dout(w_dff_A_OHKMqvh01_0),.din(w_dff_A_riVGJaof1_0),.clk(gclk));
	jdff dff_A_OHKMqvh01_0(.dout(w_dff_A_UoJBATPS9_0),.din(w_dff_A_OHKMqvh01_0),.clk(gclk));
	jdff dff_A_UoJBATPS9_0(.dout(w_dff_A_qxcCGIN92_0),.din(w_dff_A_UoJBATPS9_0),.clk(gclk));
	jdff dff_A_qxcCGIN92_0(.dout(w_dff_A_4xrl7kY22_0),.din(w_dff_A_qxcCGIN92_0),.clk(gclk));
	jdff dff_A_4xrl7kY22_0(.dout(w_dff_A_Mknr19478_0),.din(w_dff_A_4xrl7kY22_0),.clk(gclk));
	jdff dff_A_Mknr19478_0(.dout(w_dff_A_svA8ebz61_0),.din(w_dff_A_Mknr19478_0),.clk(gclk));
	jdff dff_A_svA8ebz61_0(.dout(w_dff_A_kzivBmBK6_0),.din(w_dff_A_svA8ebz61_0),.clk(gclk));
	jdff dff_A_kzivBmBK6_0(.dout(w_dff_A_0K3Z0x605_0),.din(w_dff_A_kzivBmBK6_0),.clk(gclk));
	jdff dff_A_0K3Z0x605_0(.dout(w_dff_A_QrJLNkz36_0),.din(w_dff_A_0K3Z0x605_0),.clk(gclk));
	jdff dff_A_QrJLNkz36_0(.dout(w_dff_A_PPdWaEfW9_0),.din(w_dff_A_QrJLNkz36_0),.clk(gclk));
	jdff dff_A_PPdWaEfW9_0(.dout(w_dff_A_I06EFKln0_0),.din(w_dff_A_PPdWaEfW9_0),.clk(gclk));
	jdff dff_A_I06EFKln0_0(.dout(w_dff_A_cHBsiLY41_0),.din(w_dff_A_I06EFKln0_0),.clk(gclk));
	jdff dff_A_cHBsiLY41_0(.dout(w_dff_A_B1AYvbQT0_0),.din(w_dff_A_cHBsiLY41_0),.clk(gclk));
	jdff dff_A_B1AYvbQT0_0(.dout(w_dff_A_wW4vcGgr0_0),.din(w_dff_A_B1AYvbQT0_0),.clk(gclk));
	jdff dff_A_wW4vcGgr0_0(.dout(w_dff_A_h2wgMVTM7_0),.din(w_dff_A_wW4vcGgr0_0),.clk(gclk));
	jdff dff_A_h2wgMVTM7_0(.dout(w_dff_A_xwEIdTjY5_0),.din(w_dff_A_h2wgMVTM7_0),.clk(gclk));
	jdff dff_A_xwEIdTjY5_0(.dout(w_dff_A_Ate1bxrH2_0),.din(w_dff_A_xwEIdTjY5_0),.clk(gclk));
	jdff dff_A_Ate1bxrH2_0(.dout(w_dff_A_xWrJP4dV4_0),.din(w_dff_A_Ate1bxrH2_0),.clk(gclk));
	jdff dff_A_xWrJP4dV4_0(.dout(w_dff_A_TfHyFaw49_0),.din(w_dff_A_xWrJP4dV4_0),.clk(gclk));
	jdff dff_A_TfHyFaw49_0(.dout(w_dff_A_t1HdQShF2_0),.din(w_dff_A_TfHyFaw49_0),.clk(gclk));
	jdff dff_A_t1HdQShF2_0(.dout(w_dff_A_iSfEZZln7_0),.din(w_dff_A_t1HdQShF2_0),.clk(gclk));
	jdff dff_A_iSfEZZln7_0(.dout(G486),.din(w_dff_A_iSfEZZln7_0),.clk(gclk));
	jdff dff_A_XVcUMRCc4_1(.dout(w_dff_A_2XL32K5a5_0),.din(w_dff_A_XVcUMRCc4_1),.clk(gclk));
	jdff dff_A_2XL32K5a5_0(.dout(w_dff_A_uiqhQbLz0_0),.din(w_dff_A_2XL32K5a5_0),.clk(gclk));
	jdff dff_A_uiqhQbLz0_0(.dout(w_dff_A_I0H3EQxG6_0),.din(w_dff_A_uiqhQbLz0_0),.clk(gclk));
	jdff dff_A_I0H3EQxG6_0(.dout(w_dff_A_skrDqLjC7_0),.din(w_dff_A_I0H3EQxG6_0),.clk(gclk));
	jdff dff_A_skrDqLjC7_0(.dout(w_dff_A_eKPiFpX24_0),.din(w_dff_A_skrDqLjC7_0),.clk(gclk));
	jdff dff_A_eKPiFpX24_0(.dout(w_dff_A_XS5ZKPZQ2_0),.din(w_dff_A_eKPiFpX24_0),.clk(gclk));
	jdff dff_A_XS5ZKPZQ2_0(.dout(w_dff_A_d9JQBQNR5_0),.din(w_dff_A_XS5ZKPZQ2_0),.clk(gclk));
	jdff dff_A_d9JQBQNR5_0(.dout(w_dff_A_Qe9mA7ZK9_0),.din(w_dff_A_d9JQBQNR5_0),.clk(gclk));
	jdff dff_A_Qe9mA7ZK9_0(.dout(w_dff_A_H7cQi2ZZ9_0),.din(w_dff_A_Qe9mA7ZK9_0),.clk(gclk));
	jdff dff_A_H7cQi2ZZ9_0(.dout(w_dff_A_5hcZCbP67_0),.din(w_dff_A_H7cQi2ZZ9_0),.clk(gclk));
	jdff dff_A_5hcZCbP67_0(.dout(w_dff_A_YYcf8xH19_0),.din(w_dff_A_5hcZCbP67_0),.clk(gclk));
	jdff dff_A_YYcf8xH19_0(.dout(w_dff_A_qJML1HvV1_0),.din(w_dff_A_YYcf8xH19_0),.clk(gclk));
	jdff dff_A_qJML1HvV1_0(.dout(w_dff_A_itBdxZap8_0),.din(w_dff_A_qJML1HvV1_0),.clk(gclk));
	jdff dff_A_itBdxZap8_0(.dout(w_dff_A_q7V6uhHE9_0),.din(w_dff_A_itBdxZap8_0),.clk(gclk));
	jdff dff_A_q7V6uhHE9_0(.dout(w_dff_A_flJafpRa3_0),.din(w_dff_A_q7V6uhHE9_0),.clk(gclk));
	jdff dff_A_flJafpRa3_0(.dout(w_dff_A_7HqnoKcr9_0),.din(w_dff_A_flJafpRa3_0),.clk(gclk));
	jdff dff_A_7HqnoKcr9_0(.dout(w_dff_A_am6kfWTJ2_0),.din(w_dff_A_7HqnoKcr9_0),.clk(gclk));
	jdff dff_A_am6kfWTJ2_0(.dout(w_dff_A_PT97TR9n8_0),.din(w_dff_A_am6kfWTJ2_0),.clk(gclk));
	jdff dff_A_PT97TR9n8_0(.dout(w_dff_A_nEO17RJ86_0),.din(w_dff_A_PT97TR9n8_0),.clk(gclk));
	jdff dff_A_nEO17RJ86_0(.dout(w_dff_A_nMXbaVKT6_0),.din(w_dff_A_nEO17RJ86_0),.clk(gclk));
	jdff dff_A_nMXbaVKT6_0(.dout(w_dff_A_cx7gEuE66_0),.din(w_dff_A_nMXbaVKT6_0),.clk(gclk));
	jdff dff_A_cx7gEuE66_0(.dout(w_dff_A_0ajAiqWc5_0),.din(w_dff_A_cx7gEuE66_0),.clk(gclk));
	jdff dff_A_0ajAiqWc5_0(.dout(w_dff_A_8A9axYqh7_0),.din(w_dff_A_0ajAiqWc5_0),.clk(gclk));
	jdff dff_A_8A9axYqh7_0(.dout(w_dff_A_XspSFBXe7_0),.din(w_dff_A_8A9axYqh7_0),.clk(gclk));
	jdff dff_A_XspSFBXe7_0(.dout(w_dff_A_if33SzG11_0),.din(w_dff_A_XspSFBXe7_0),.clk(gclk));
	jdff dff_A_if33SzG11_0(.dout(w_dff_A_Zc6ARDFB9_0),.din(w_dff_A_if33SzG11_0),.clk(gclk));
	jdff dff_A_Zc6ARDFB9_0(.dout(G484),.din(w_dff_A_Zc6ARDFB9_0),.clk(gclk));
	jdff dff_A_2X5xRMEh0_1(.dout(w_dff_A_QhKLMCDo0_0),.din(w_dff_A_2X5xRMEh0_1),.clk(gclk));
	jdff dff_A_QhKLMCDo0_0(.dout(w_dff_A_xoJHySdq8_0),.din(w_dff_A_QhKLMCDo0_0),.clk(gclk));
	jdff dff_A_xoJHySdq8_0(.dout(w_dff_A_x2EV1CAA2_0),.din(w_dff_A_xoJHySdq8_0),.clk(gclk));
	jdff dff_A_x2EV1CAA2_0(.dout(w_dff_A_Q2FxQJNX8_0),.din(w_dff_A_x2EV1CAA2_0),.clk(gclk));
	jdff dff_A_Q2FxQJNX8_0(.dout(w_dff_A_iuf1dv8M4_0),.din(w_dff_A_Q2FxQJNX8_0),.clk(gclk));
	jdff dff_A_iuf1dv8M4_0(.dout(w_dff_A_K8U8DyHM7_0),.din(w_dff_A_iuf1dv8M4_0),.clk(gclk));
	jdff dff_A_K8U8DyHM7_0(.dout(w_dff_A_itkhR4eT1_0),.din(w_dff_A_K8U8DyHM7_0),.clk(gclk));
	jdff dff_A_itkhR4eT1_0(.dout(w_dff_A_AgbtkyvS5_0),.din(w_dff_A_itkhR4eT1_0),.clk(gclk));
	jdff dff_A_AgbtkyvS5_0(.dout(w_dff_A_ouI8tdeK2_0),.din(w_dff_A_AgbtkyvS5_0),.clk(gclk));
	jdff dff_A_ouI8tdeK2_0(.dout(w_dff_A_oBgR1p2P5_0),.din(w_dff_A_ouI8tdeK2_0),.clk(gclk));
	jdff dff_A_oBgR1p2P5_0(.dout(w_dff_A_6AUMgknj6_0),.din(w_dff_A_oBgR1p2P5_0),.clk(gclk));
	jdff dff_A_6AUMgknj6_0(.dout(w_dff_A_TljI974m2_0),.din(w_dff_A_6AUMgknj6_0),.clk(gclk));
	jdff dff_A_TljI974m2_0(.dout(w_dff_A_rOlg9TRa1_0),.din(w_dff_A_TljI974m2_0),.clk(gclk));
	jdff dff_A_rOlg9TRa1_0(.dout(w_dff_A_H6k6SU3b9_0),.din(w_dff_A_rOlg9TRa1_0),.clk(gclk));
	jdff dff_A_H6k6SU3b9_0(.dout(w_dff_A_z6eheY2D6_0),.din(w_dff_A_H6k6SU3b9_0),.clk(gclk));
	jdff dff_A_z6eheY2D6_0(.dout(w_dff_A_D0db2zeP7_0),.din(w_dff_A_z6eheY2D6_0),.clk(gclk));
	jdff dff_A_D0db2zeP7_0(.dout(w_dff_A_yAmStAph0_0),.din(w_dff_A_D0db2zeP7_0),.clk(gclk));
	jdff dff_A_yAmStAph0_0(.dout(w_dff_A_JCvmZCsm9_0),.din(w_dff_A_yAmStAph0_0),.clk(gclk));
	jdff dff_A_JCvmZCsm9_0(.dout(w_dff_A_MoXNtrmj5_0),.din(w_dff_A_JCvmZCsm9_0),.clk(gclk));
	jdff dff_A_MoXNtrmj5_0(.dout(w_dff_A_aWvnoDxi1_0),.din(w_dff_A_MoXNtrmj5_0),.clk(gclk));
	jdff dff_A_aWvnoDxi1_0(.dout(w_dff_A_WFxlR3mX4_0),.din(w_dff_A_aWvnoDxi1_0),.clk(gclk));
	jdff dff_A_WFxlR3mX4_0(.dout(w_dff_A_KVDf182v8_0),.din(w_dff_A_WFxlR3mX4_0),.clk(gclk));
	jdff dff_A_KVDf182v8_0(.dout(w_dff_A_VYsIQfsL2_0),.din(w_dff_A_KVDf182v8_0),.clk(gclk));
	jdff dff_A_VYsIQfsL2_0(.dout(w_dff_A_tWLu8ACo1_0),.din(w_dff_A_VYsIQfsL2_0),.clk(gclk));
	jdff dff_A_tWLu8ACo1_0(.dout(w_dff_A_SAREJ7FE5_0),.din(w_dff_A_tWLu8ACo1_0),.clk(gclk));
	jdff dff_A_SAREJ7FE5_0(.dout(w_dff_A_BQV1a3BO5_0),.din(w_dff_A_SAREJ7FE5_0),.clk(gclk));
	jdff dff_A_BQV1a3BO5_0(.dout(G482),.din(w_dff_A_BQV1a3BO5_0),.clk(gclk));
	jdff dff_A_UVJM26EF8_1(.dout(w_dff_A_i6TuLoRs3_0),.din(w_dff_A_UVJM26EF8_1),.clk(gclk));
	jdff dff_A_i6TuLoRs3_0(.dout(w_dff_A_9oRqyi9l5_0),.din(w_dff_A_i6TuLoRs3_0),.clk(gclk));
	jdff dff_A_9oRqyi9l5_0(.dout(w_dff_A_6kCn5a197_0),.din(w_dff_A_9oRqyi9l5_0),.clk(gclk));
	jdff dff_A_6kCn5a197_0(.dout(w_dff_A_fqm05VUl5_0),.din(w_dff_A_6kCn5a197_0),.clk(gclk));
	jdff dff_A_fqm05VUl5_0(.dout(w_dff_A_E9KPb7G35_0),.din(w_dff_A_fqm05VUl5_0),.clk(gclk));
	jdff dff_A_E9KPb7G35_0(.dout(w_dff_A_H5iiDeJ55_0),.din(w_dff_A_E9KPb7G35_0),.clk(gclk));
	jdff dff_A_H5iiDeJ55_0(.dout(w_dff_A_QU1YMUfJ3_0),.din(w_dff_A_H5iiDeJ55_0),.clk(gclk));
	jdff dff_A_QU1YMUfJ3_0(.dout(w_dff_A_xRbZXwEe4_0),.din(w_dff_A_QU1YMUfJ3_0),.clk(gclk));
	jdff dff_A_xRbZXwEe4_0(.dout(w_dff_A_hwpKUmEP9_0),.din(w_dff_A_xRbZXwEe4_0),.clk(gclk));
	jdff dff_A_hwpKUmEP9_0(.dout(w_dff_A_B8SMUqDP0_0),.din(w_dff_A_hwpKUmEP9_0),.clk(gclk));
	jdff dff_A_B8SMUqDP0_0(.dout(w_dff_A_XcnpKTvR5_0),.din(w_dff_A_B8SMUqDP0_0),.clk(gclk));
	jdff dff_A_XcnpKTvR5_0(.dout(w_dff_A_dCgBkjfG5_0),.din(w_dff_A_XcnpKTvR5_0),.clk(gclk));
	jdff dff_A_dCgBkjfG5_0(.dout(w_dff_A_H9IGAGpg8_0),.din(w_dff_A_dCgBkjfG5_0),.clk(gclk));
	jdff dff_A_H9IGAGpg8_0(.dout(w_dff_A_ku4suilp2_0),.din(w_dff_A_H9IGAGpg8_0),.clk(gclk));
	jdff dff_A_ku4suilp2_0(.dout(w_dff_A_VD3HGzX16_0),.din(w_dff_A_ku4suilp2_0),.clk(gclk));
	jdff dff_A_VD3HGzX16_0(.dout(w_dff_A_GWFkJgQs7_0),.din(w_dff_A_VD3HGzX16_0),.clk(gclk));
	jdff dff_A_GWFkJgQs7_0(.dout(w_dff_A_q0fx0zhG4_0),.din(w_dff_A_GWFkJgQs7_0),.clk(gclk));
	jdff dff_A_q0fx0zhG4_0(.dout(w_dff_A_N3xuPTX42_0),.din(w_dff_A_q0fx0zhG4_0),.clk(gclk));
	jdff dff_A_N3xuPTX42_0(.dout(w_dff_A_MRqUz9zT0_0),.din(w_dff_A_N3xuPTX42_0),.clk(gclk));
	jdff dff_A_MRqUz9zT0_0(.dout(w_dff_A_4ljUYqqs2_0),.din(w_dff_A_MRqUz9zT0_0),.clk(gclk));
	jdff dff_A_4ljUYqqs2_0(.dout(w_dff_A_VVYC8VWJ8_0),.din(w_dff_A_4ljUYqqs2_0),.clk(gclk));
	jdff dff_A_VVYC8VWJ8_0(.dout(w_dff_A_4KzcN3DW1_0),.din(w_dff_A_VVYC8VWJ8_0),.clk(gclk));
	jdff dff_A_4KzcN3DW1_0(.dout(w_dff_A_ztYYscuJ9_0),.din(w_dff_A_4KzcN3DW1_0),.clk(gclk));
	jdff dff_A_ztYYscuJ9_0(.dout(w_dff_A_ahxJdMfr0_0),.din(w_dff_A_ztYYscuJ9_0),.clk(gclk));
	jdff dff_A_ahxJdMfr0_0(.dout(w_dff_A_NCk9sWGy3_0),.din(w_dff_A_ahxJdMfr0_0),.clk(gclk));
	jdff dff_A_NCk9sWGy3_0(.dout(w_dff_A_uXRT81rD0_0),.din(w_dff_A_NCk9sWGy3_0),.clk(gclk));
	jdff dff_A_uXRT81rD0_0(.dout(G480),.din(w_dff_A_uXRT81rD0_0),.clk(gclk));
	jdff dff_A_a6FX4fFz9_1(.dout(w_dff_A_eiRbZAcj3_0),.din(w_dff_A_a6FX4fFz9_1),.clk(gclk));
	jdff dff_A_eiRbZAcj3_0(.dout(w_dff_A_2NGTuXiE8_0),.din(w_dff_A_eiRbZAcj3_0),.clk(gclk));
	jdff dff_A_2NGTuXiE8_0(.dout(w_dff_A_ECqpv6Si5_0),.din(w_dff_A_2NGTuXiE8_0),.clk(gclk));
	jdff dff_A_ECqpv6Si5_0(.dout(w_dff_A_q2IyGvVA7_0),.din(w_dff_A_ECqpv6Si5_0),.clk(gclk));
	jdff dff_A_q2IyGvVA7_0(.dout(w_dff_A_OGRgURPJ6_0),.din(w_dff_A_q2IyGvVA7_0),.clk(gclk));
	jdff dff_A_OGRgURPJ6_0(.dout(w_dff_A_3WwiB7mi3_0),.din(w_dff_A_OGRgURPJ6_0),.clk(gclk));
	jdff dff_A_3WwiB7mi3_0(.dout(w_dff_A_ghmiQXIz0_0),.din(w_dff_A_3WwiB7mi3_0),.clk(gclk));
	jdff dff_A_ghmiQXIz0_0(.dout(w_dff_A_xbKUBTv07_0),.din(w_dff_A_ghmiQXIz0_0),.clk(gclk));
	jdff dff_A_xbKUBTv07_0(.dout(w_dff_A_4XwgKWSw7_0),.din(w_dff_A_xbKUBTv07_0),.clk(gclk));
	jdff dff_A_4XwgKWSw7_0(.dout(w_dff_A_DfPAWoO77_0),.din(w_dff_A_4XwgKWSw7_0),.clk(gclk));
	jdff dff_A_DfPAWoO77_0(.dout(w_dff_A_1E4wGx5g0_0),.din(w_dff_A_DfPAWoO77_0),.clk(gclk));
	jdff dff_A_1E4wGx5g0_0(.dout(w_dff_A_aJuQUz3s2_0),.din(w_dff_A_1E4wGx5g0_0),.clk(gclk));
	jdff dff_A_aJuQUz3s2_0(.dout(w_dff_A_pX7Ngyzw3_0),.din(w_dff_A_aJuQUz3s2_0),.clk(gclk));
	jdff dff_A_pX7Ngyzw3_0(.dout(w_dff_A_v6Xn2vI24_0),.din(w_dff_A_pX7Ngyzw3_0),.clk(gclk));
	jdff dff_A_v6Xn2vI24_0(.dout(w_dff_A_rupQpY467_0),.din(w_dff_A_v6Xn2vI24_0),.clk(gclk));
	jdff dff_A_rupQpY467_0(.dout(w_dff_A_GlKq3nDu6_0),.din(w_dff_A_rupQpY467_0),.clk(gclk));
	jdff dff_A_GlKq3nDu6_0(.dout(w_dff_A_I4GJ84Kh3_0),.din(w_dff_A_GlKq3nDu6_0),.clk(gclk));
	jdff dff_A_I4GJ84Kh3_0(.dout(w_dff_A_MvtqI6Uu6_0),.din(w_dff_A_I4GJ84Kh3_0),.clk(gclk));
	jdff dff_A_MvtqI6Uu6_0(.dout(w_dff_A_1mmkwmZc5_0),.din(w_dff_A_MvtqI6Uu6_0),.clk(gclk));
	jdff dff_A_1mmkwmZc5_0(.dout(w_dff_A_7zvifdWB9_0),.din(w_dff_A_1mmkwmZc5_0),.clk(gclk));
	jdff dff_A_7zvifdWB9_0(.dout(w_dff_A_uE0b65iD8_0),.din(w_dff_A_7zvifdWB9_0),.clk(gclk));
	jdff dff_A_uE0b65iD8_0(.dout(w_dff_A_PlQ2456R7_0),.din(w_dff_A_uE0b65iD8_0),.clk(gclk));
	jdff dff_A_PlQ2456R7_0(.dout(w_dff_A_MUdrsE2A6_0),.din(w_dff_A_PlQ2456R7_0),.clk(gclk));
	jdff dff_A_MUdrsE2A6_0(.dout(w_dff_A_CTuzU1hT1_0),.din(w_dff_A_MUdrsE2A6_0),.clk(gclk));
	jdff dff_A_CTuzU1hT1_0(.dout(w_dff_A_4xyssGQu3_0),.din(w_dff_A_CTuzU1hT1_0),.clk(gclk));
	jdff dff_A_4xyssGQu3_0(.dout(w_dff_A_GbszCoWy4_0),.din(w_dff_A_4xyssGQu3_0),.clk(gclk));
	jdff dff_A_GbszCoWy4_0(.dout(G560),.din(w_dff_A_GbszCoWy4_0),.clk(gclk));
	jdff dff_A_HMyMtu9z5_1(.dout(w_dff_A_Oda4MulR5_0),.din(w_dff_A_HMyMtu9z5_1),.clk(gclk));
	jdff dff_A_Oda4MulR5_0(.dout(w_dff_A_02eHjLip2_0),.din(w_dff_A_Oda4MulR5_0),.clk(gclk));
	jdff dff_A_02eHjLip2_0(.dout(w_dff_A_TXoHwLFK6_0),.din(w_dff_A_02eHjLip2_0),.clk(gclk));
	jdff dff_A_TXoHwLFK6_0(.dout(w_dff_A_TrKKGpym4_0),.din(w_dff_A_TXoHwLFK6_0),.clk(gclk));
	jdff dff_A_TrKKGpym4_0(.dout(w_dff_A_1l0W9sy27_0),.din(w_dff_A_TrKKGpym4_0),.clk(gclk));
	jdff dff_A_1l0W9sy27_0(.dout(w_dff_A_1C3jH5xg4_0),.din(w_dff_A_1l0W9sy27_0),.clk(gclk));
	jdff dff_A_1C3jH5xg4_0(.dout(w_dff_A_k4JahgB24_0),.din(w_dff_A_1C3jH5xg4_0),.clk(gclk));
	jdff dff_A_k4JahgB24_0(.dout(w_dff_A_npH477mu3_0),.din(w_dff_A_k4JahgB24_0),.clk(gclk));
	jdff dff_A_npH477mu3_0(.dout(w_dff_A_QVhByDoc8_0),.din(w_dff_A_npH477mu3_0),.clk(gclk));
	jdff dff_A_QVhByDoc8_0(.dout(w_dff_A_WX0wXZdp9_0),.din(w_dff_A_QVhByDoc8_0),.clk(gclk));
	jdff dff_A_WX0wXZdp9_0(.dout(w_dff_A_KR2LJcZ93_0),.din(w_dff_A_WX0wXZdp9_0),.clk(gclk));
	jdff dff_A_KR2LJcZ93_0(.dout(w_dff_A_ALkl92LC8_0),.din(w_dff_A_KR2LJcZ93_0),.clk(gclk));
	jdff dff_A_ALkl92LC8_0(.dout(w_dff_A_a4x8kVNw2_0),.din(w_dff_A_ALkl92LC8_0),.clk(gclk));
	jdff dff_A_a4x8kVNw2_0(.dout(w_dff_A_sSIPKGpG6_0),.din(w_dff_A_a4x8kVNw2_0),.clk(gclk));
	jdff dff_A_sSIPKGpG6_0(.dout(w_dff_A_rEny0QEk6_0),.din(w_dff_A_sSIPKGpG6_0),.clk(gclk));
	jdff dff_A_rEny0QEk6_0(.dout(w_dff_A_AYL74And5_0),.din(w_dff_A_rEny0QEk6_0),.clk(gclk));
	jdff dff_A_AYL74And5_0(.dout(w_dff_A_IumQ7v2L5_0),.din(w_dff_A_AYL74And5_0),.clk(gclk));
	jdff dff_A_IumQ7v2L5_0(.dout(w_dff_A_1vJbo5Dd8_0),.din(w_dff_A_IumQ7v2L5_0),.clk(gclk));
	jdff dff_A_1vJbo5Dd8_0(.dout(w_dff_A_VnItcIAc9_0),.din(w_dff_A_1vJbo5Dd8_0),.clk(gclk));
	jdff dff_A_VnItcIAc9_0(.dout(w_dff_A_kUvtkle29_0),.din(w_dff_A_VnItcIAc9_0),.clk(gclk));
	jdff dff_A_kUvtkle29_0(.dout(w_dff_A_iHYF3vKC0_0),.din(w_dff_A_kUvtkle29_0),.clk(gclk));
	jdff dff_A_iHYF3vKC0_0(.dout(w_dff_A_kHX26XH09_0),.din(w_dff_A_iHYF3vKC0_0),.clk(gclk));
	jdff dff_A_kHX26XH09_0(.dout(w_dff_A_XomNeiLg2_0),.din(w_dff_A_kHX26XH09_0),.clk(gclk));
	jdff dff_A_XomNeiLg2_0(.dout(w_dff_A_kf7QsZNn2_0),.din(w_dff_A_XomNeiLg2_0),.clk(gclk));
	jdff dff_A_kf7QsZNn2_0(.dout(w_dff_A_SSEskHef4_0),.din(w_dff_A_kf7QsZNn2_0),.clk(gclk));
	jdff dff_A_SSEskHef4_0(.dout(w_dff_A_9ScruEEl7_0),.din(w_dff_A_SSEskHef4_0),.clk(gclk));
	jdff dff_A_9ScruEEl7_0(.dout(G542),.din(w_dff_A_9ScruEEl7_0),.clk(gclk));
	jdff dff_A_OHRyQi3h5_1(.dout(w_dff_A_W2WcKkq43_0),.din(w_dff_A_OHRyQi3h5_1),.clk(gclk));
	jdff dff_A_W2WcKkq43_0(.dout(w_dff_A_8YUjki5V6_0),.din(w_dff_A_W2WcKkq43_0),.clk(gclk));
	jdff dff_A_8YUjki5V6_0(.dout(w_dff_A_umkkhyZQ7_0),.din(w_dff_A_8YUjki5V6_0),.clk(gclk));
	jdff dff_A_umkkhyZQ7_0(.dout(w_dff_A_anJuRmiT8_0),.din(w_dff_A_umkkhyZQ7_0),.clk(gclk));
	jdff dff_A_anJuRmiT8_0(.dout(w_dff_A_IXEjX2Zj5_0),.din(w_dff_A_anJuRmiT8_0),.clk(gclk));
	jdff dff_A_IXEjX2Zj5_0(.dout(w_dff_A_TjqDjezA9_0),.din(w_dff_A_IXEjX2Zj5_0),.clk(gclk));
	jdff dff_A_TjqDjezA9_0(.dout(w_dff_A_QpdUBKOj0_0),.din(w_dff_A_TjqDjezA9_0),.clk(gclk));
	jdff dff_A_QpdUBKOj0_0(.dout(w_dff_A_AkhbvrF87_0),.din(w_dff_A_QpdUBKOj0_0),.clk(gclk));
	jdff dff_A_AkhbvrF87_0(.dout(w_dff_A_rD44rxAP8_0),.din(w_dff_A_AkhbvrF87_0),.clk(gclk));
	jdff dff_A_rD44rxAP8_0(.dout(w_dff_A_JJfsPPqT3_0),.din(w_dff_A_rD44rxAP8_0),.clk(gclk));
	jdff dff_A_JJfsPPqT3_0(.dout(w_dff_A_YkeD6l6y2_0),.din(w_dff_A_JJfsPPqT3_0),.clk(gclk));
	jdff dff_A_YkeD6l6y2_0(.dout(w_dff_A_orUc6Xb24_0),.din(w_dff_A_YkeD6l6y2_0),.clk(gclk));
	jdff dff_A_orUc6Xb24_0(.dout(w_dff_A_qkWj9AlW2_0),.din(w_dff_A_orUc6Xb24_0),.clk(gclk));
	jdff dff_A_qkWj9AlW2_0(.dout(w_dff_A_zNYmYpgW6_0),.din(w_dff_A_qkWj9AlW2_0),.clk(gclk));
	jdff dff_A_zNYmYpgW6_0(.dout(w_dff_A_bCUkCvry3_0),.din(w_dff_A_zNYmYpgW6_0),.clk(gclk));
	jdff dff_A_bCUkCvry3_0(.dout(w_dff_A_ZBcUn4h43_0),.din(w_dff_A_bCUkCvry3_0),.clk(gclk));
	jdff dff_A_ZBcUn4h43_0(.dout(w_dff_A_Yk9Xn3tS8_0),.din(w_dff_A_ZBcUn4h43_0),.clk(gclk));
	jdff dff_A_Yk9Xn3tS8_0(.dout(w_dff_A_loWhWcEG5_0),.din(w_dff_A_Yk9Xn3tS8_0),.clk(gclk));
	jdff dff_A_loWhWcEG5_0(.dout(w_dff_A_geT7kneF7_0),.din(w_dff_A_loWhWcEG5_0),.clk(gclk));
	jdff dff_A_geT7kneF7_0(.dout(w_dff_A_Jr7JidRa7_0),.din(w_dff_A_geT7kneF7_0),.clk(gclk));
	jdff dff_A_Jr7JidRa7_0(.dout(w_dff_A_iaADX08z7_0),.din(w_dff_A_Jr7JidRa7_0),.clk(gclk));
	jdff dff_A_iaADX08z7_0(.dout(w_dff_A_6lNPjQJD2_0),.din(w_dff_A_iaADX08z7_0),.clk(gclk));
	jdff dff_A_6lNPjQJD2_0(.dout(w_dff_A_eDdb3zBx5_0),.din(w_dff_A_6lNPjQJD2_0),.clk(gclk));
	jdff dff_A_eDdb3zBx5_0(.dout(w_dff_A_ETV3iEVH1_0),.din(w_dff_A_eDdb3zBx5_0),.clk(gclk));
	jdff dff_A_ETV3iEVH1_0(.dout(w_dff_A_j9RR9sOp0_0),.din(w_dff_A_ETV3iEVH1_0),.clk(gclk));
	jdff dff_A_j9RR9sOp0_0(.dout(w_dff_A_dSihZrmM2_0),.din(w_dff_A_j9RR9sOp0_0),.clk(gclk));
	jdff dff_A_dSihZrmM2_0(.dout(G558),.din(w_dff_A_dSihZrmM2_0),.clk(gclk));
	jdff dff_A_dqNBR2IS5_1(.dout(w_dff_A_S1DAVp1q5_0),.din(w_dff_A_dqNBR2IS5_1),.clk(gclk));
	jdff dff_A_S1DAVp1q5_0(.dout(w_dff_A_zhsLltyh1_0),.din(w_dff_A_S1DAVp1q5_0),.clk(gclk));
	jdff dff_A_zhsLltyh1_0(.dout(w_dff_A_RT9v651b1_0),.din(w_dff_A_zhsLltyh1_0),.clk(gclk));
	jdff dff_A_RT9v651b1_0(.dout(w_dff_A_A13NeRXC2_0),.din(w_dff_A_RT9v651b1_0),.clk(gclk));
	jdff dff_A_A13NeRXC2_0(.dout(w_dff_A_vIQoAH6w6_0),.din(w_dff_A_A13NeRXC2_0),.clk(gclk));
	jdff dff_A_vIQoAH6w6_0(.dout(w_dff_A_uWRfxGeZ3_0),.din(w_dff_A_vIQoAH6w6_0),.clk(gclk));
	jdff dff_A_uWRfxGeZ3_0(.dout(w_dff_A_Y0LhGxmk0_0),.din(w_dff_A_uWRfxGeZ3_0),.clk(gclk));
	jdff dff_A_Y0LhGxmk0_0(.dout(w_dff_A_xrYYrI2L2_0),.din(w_dff_A_Y0LhGxmk0_0),.clk(gclk));
	jdff dff_A_xrYYrI2L2_0(.dout(w_dff_A_1UiSVUEH1_0),.din(w_dff_A_xrYYrI2L2_0),.clk(gclk));
	jdff dff_A_1UiSVUEH1_0(.dout(w_dff_A_SkN7ktfM0_0),.din(w_dff_A_1UiSVUEH1_0),.clk(gclk));
	jdff dff_A_SkN7ktfM0_0(.dout(w_dff_A_1XAxCiMS3_0),.din(w_dff_A_SkN7ktfM0_0),.clk(gclk));
	jdff dff_A_1XAxCiMS3_0(.dout(w_dff_A_CZgN9Gqr8_0),.din(w_dff_A_1XAxCiMS3_0),.clk(gclk));
	jdff dff_A_CZgN9Gqr8_0(.dout(w_dff_A_7t0dQJ0K0_0),.din(w_dff_A_CZgN9Gqr8_0),.clk(gclk));
	jdff dff_A_7t0dQJ0K0_0(.dout(w_dff_A_UgVaJFKq7_0),.din(w_dff_A_7t0dQJ0K0_0),.clk(gclk));
	jdff dff_A_UgVaJFKq7_0(.dout(w_dff_A_oj0xsLmL4_0),.din(w_dff_A_UgVaJFKq7_0),.clk(gclk));
	jdff dff_A_oj0xsLmL4_0(.dout(w_dff_A_qYB2syE41_0),.din(w_dff_A_oj0xsLmL4_0),.clk(gclk));
	jdff dff_A_qYB2syE41_0(.dout(w_dff_A_uBg0JGeT4_0),.din(w_dff_A_qYB2syE41_0),.clk(gclk));
	jdff dff_A_uBg0JGeT4_0(.dout(w_dff_A_Vi7D5nUp8_0),.din(w_dff_A_uBg0JGeT4_0),.clk(gclk));
	jdff dff_A_Vi7D5nUp8_0(.dout(w_dff_A_Xq68wXmm9_0),.din(w_dff_A_Vi7D5nUp8_0),.clk(gclk));
	jdff dff_A_Xq68wXmm9_0(.dout(w_dff_A_4H6abfMT1_0),.din(w_dff_A_Xq68wXmm9_0),.clk(gclk));
	jdff dff_A_4H6abfMT1_0(.dout(w_dff_A_WEHCrI3G6_0),.din(w_dff_A_4H6abfMT1_0),.clk(gclk));
	jdff dff_A_WEHCrI3G6_0(.dout(w_dff_A_nQTkL1FI6_0),.din(w_dff_A_WEHCrI3G6_0),.clk(gclk));
	jdff dff_A_nQTkL1FI6_0(.dout(w_dff_A_V03hrBgb5_0),.din(w_dff_A_nQTkL1FI6_0),.clk(gclk));
	jdff dff_A_V03hrBgb5_0(.dout(w_dff_A_C94sgvYw2_0),.din(w_dff_A_V03hrBgb5_0),.clk(gclk));
	jdff dff_A_C94sgvYw2_0(.dout(w_dff_A_8zOvM1ON5_0),.din(w_dff_A_C94sgvYw2_0),.clk(gclk));
	jdff dff_A_8zOvM1ON5_0(.dout(w_dff_A_Ovb05qxY2_0),.din(w_dff_A_8zOvM1ON5_0),.clk(gclk));
	jdff dff_A_Ovb05qxY2_0(.dout(G556),.din(w_dff_A_Ovb05qxY2_0),.clk(gclk));
	jdff dff_A_0ww2XJtm7_1(.dout(w_dff_A_n42dURt56_0),.din(w_dff_A_0ww2XJtm7_1),.clk(gclk));
	jdff dff_A_n42dURt56_0(.dout(w_dff_A_wZgojSWX6_0),.din(w_dff_A_n42dURt56_0),.clk(gclk));
	jdff dff_A_wZgojSWX6_0(.dout(w_dff_A_XmT3ztM21_0),.din(w_dff_A_wZgojSWX6_0),.clk(gclk));
	jdff dff_A_XmT3ztM21_0(.dout(w_dff_A_PpBJ0wIq6_0),.din(w_dff_A_XmT3ztM21_0),.clk(gclk));
	jdff dff_A_PpBJ0wIq6_0(.dout(w_dff_A_VaOJbH567_0),.din(w_dff_A_PpBJ0wIq6_0),.clk(gclk));
	jdff dff_A_VaOJbH567_0(.dout(w_dff_A_FWh45Sc56_0),.din(w_dff_A_VaOJbH567_0),.clk(gclk));
	jdff dff_A_FWh45Sc56_0(.dout(w_dff_A_PD5Hi5G89_0),.din(w_dff_A_FWh45Sc56_0),.clk(gclk));
	jdff dff_A_PD5Hi5G89_0(.dout(w_dff_A_jY9AWEXO9_0),.din(w_dff_A_PD5Hi5G89_0),.clk(gclk));
	jdff dff_A_jY9AWEXO9_0(.dout(w_dff_A_bUCTdUdC6_0),.din(w_dff_A_jY9AWEXO9_0),.clk(gclk));
	jdff dff_A_bUCTdUdC6_0(.dout(w_dff_A_K6j75fEW5_0),.din(w_dff_A_bUCTdUdC6_0),.clk(gclk));
	jdff dff_A_K6j75fEW5_0(.dout(w_dff_A_0hiITqoz4_0),.din(w_dff_A_K6j75fEW5_0),.clk(gclk));
	jdff dff_A_0hiITqoz4_0(.dout(w_dff_A_8l5G66fv5_0),.din(w_dff_A_0hiITqoz4_0),.clk(gclk));
	jdff dff_A_8l5G66fv5_0(.dout(w_dff_A_MJScctTp4_0),.din(w_dff_A_8l5G66fv5_0),.clk(gclk));
	jdff dff_A_MJScctTp4_0(.dout(w_dff_A_NZNle9D65_0),.din(w_dff_A_MJScctTp4_0),.clk(gclk));
	jdff dff_A_NZNle9D65_0(.dout(w_dff_A_RJU9zxHS7_0),.din(w_dff_A_NZNle9D65_0),.clk(gclk));
	jdff dff_A_RJU9zxHS7_0(.dout(w_dff_A_IqURtX018_0),.din(w_dff_A_RJU9zxHS7_0),.clk(gclk));
	jdff dff_A_IqURtX018_0(.dout(w_dff_A_OGBoosG52_0),.din(w_dff_A_IqURtX018_0),.clk(gclk));
	jdff dff_A_OGBoosG52_0(.dout(w_dff_A_Y3SAtFLq1_0),.din(w_dff_A_OGBoosG52_0),.clk(gclk));
	jdff dff_A_Y3SAtFLq1_0(.dout(w_dff_A_MxI6ffKQ9_0),.din(w_dff_A_Y3SAtFLq1_0),.clk(gclk));
	jdff dff_A_MxI6ffKQ9_0(.dout(w_dff_A_a6yuZfwa0_0),.din(w_dff_A_MxI6ffKQ9_0),.clk(gclk));
	jdff dff_A_a6yuZfwa0_0(.dout(w_dff_A_VxiBZGlw9_0),.din(w_dff_A_a6yuZfwa0_0),.clk(gclk));
	jdff dff_A_VxiBZGlw9_0(.dout(w_dff_A_M1DoU9cO0_0),.din(w_dff_A_VxiBZGlw9_0),.clk(gclk));
	jdff dff_A_M1DoU9cO0_0(.dout(w_dff_A_cc22uoNB1_0),.din(w_dff_A_M1DoU9cO0_0),.clk(gclk));
	jdff dff_A_cc22uoNB1_0(.dout(w_dff_A_E0jpqo7z0_0),.din(w_dff_A_cc22uoNB1_0),.clk(gclk));
	jdff dff_A_E0jpqo7z0_0(.dout(w_dff_A_pyrRYMqX5_0),.din(w_dff_A_E0jpqo7z0_0),.clk(gclk));
	jdff dff_A_pyrRYMqX5_0(.dout(w_dff_A_NC3FtzoI3_0),.din(w_dff_A_pyrRYMqX5_0),.clk(gclk));
	jdff dff_A_NC3FtzoI3_0(.dout(G554),.din(w_dff_A_NC3FtzoI3_0),.clk(gclk));
	jdff dff_A_wEixxhLY1_1(.dout(w_dff_A_iL3knU1R5_0),.din(w_dff_A_wEixxhLY1_1),.clk(gclk));
	jdff dff_A_iL3knU1R5_0(.dout(w_dff_A_Zw0v5R6c1_0),.din(w_dff_A_iL3knU1R5_0),.clk(gclk));
	jdff dff_A_Zw0v5R6c1_0(.dout(w_dff_A_S4i9spnq0_0),.din(w_dff_A_Zw0v5R6c1_0),.clk(gclk));
	jdff dff_A_S4i9spnq0_0(.dout(w_dff_A_T2GnmU1C6_0),.din(w_dff_A_S4i9spnq0_0),.clk(gclk));
	jdff dff_A_T2GnmU1C6_0(.dout(w_dff_A_3h8ks7S83_0),.din(w_dff_A_T2GnmU1C6_0),.clk(gclk));
	jdff dff_A_3h8ks7S83_0(.dout(w_dff_A_5T0ksZaP8_0),.din(w_dff_A_3h8ks7S83_0),.clk(gclk));
	jdff dff_A_5T0ksZaP8_0(.dout(w_dff_A_940vZeEa0_0),.din(w_dff_A_5T0ksZaP8_0),.clk(gclk));
	jdff dff_A_940vZeEa0_0(.dout(w_dff_A_icrPN5md5_0),.din(w_dff_A_940vZeEa0_0),.clk(gclk));
	jdff dff_A_icrPN5md5_0(.dout(w_dff_A_owhbLnWn4_0),.din(w_dff_A_icrPN5md5_0),.clk(gclk));
	jdff dff_A_owhbLnWn4_0(.dout(w_dff_A_EYBjuh1g9_0),.din(w_dff_A_owhbLnWn4_0),.clk(gclk));
	jdff dff_A_EYBjuh1g9_0(.dout(w_dff_A_863N7VV51_0),.din(w_dff_A_EYBjuh1g9_0),.clk(gclk));
	jdff dff_A_863N7VV51_0(.dout(w_dff_A_k8i8ZwRV2_0),.din(w_dff_A_863N7VV51_0),.clk(gclk));
	jdff dff_A_k8i8ZwRV2_0(.dout(w_dff_A_OUszzLtT2_0),.din(w_dff_A_k8i8ZwRV2_0),.clk(gclk));
	jdff dff_A_OUszzLtT2_0(.dout(w_dff_A_ipEg6L4a3_0),.din(w_dff_A_OUszzLtT2_0),.clk(gclk));
	jdff dff_A_ipEg6L4a3_0(.dout(w_dff_A_Z82bfm5B6_0),.din(w_dff_A_ipEg6L4a3_0),.clk(gclk));
	jdff dff_A_Z82bfm5B6_0(.dout(w_dff_A_fmOlB9oe5_0),.din(w_dff_A_Z82bfm5B6_0),.clk(gclk));
	jdff dff_A_fmOlB9oe5_0(.dout(w_dff_A_PD7BoTEb9_0),.din(w_dff_A_fmOlB9oe5_0),.clk(gclk));
	jdff dff_A_PD7BoTEb9_0(.dout(w_dff_A_o6lqqRf64_0),.din(w_dff_A_PD7BoTEb9_0),.clk(gclk));
	jdff dff_A_o6lqqRf64_0(.dout(w_dff_A_1aDcas5O5_0),.din(w_dff_A_o6lqqRf64_0),.clk(gclk));
	jdff dff_A_1aDcas5O5_0(.dout(w_dff_A_Bp9lLQnl1_0),.din(w_dff_A_1aDcas5O5_0),.clk(gclk));
	jdff dff_A_Bp9lLQnl1_0(.dout(w_dff_A_Lk1djuk33_0),.din(w_dff_A_Bp9lLQnl1_0),.clk(gclk));
	jdff dff_A_Lk1djuk33_0(.dout(w_dff_A_tIKM2B2x1_0),.din(w_dff_A_Lk1djuk33_0),.clk(gclk));
	jdff dff_A_tIKM2B2x1_0(.dout(w_dff_A_uUAeA6aC8_0),.din(w_dff_A_tIKM2B2x1_0),.clk(gclk));
	jdff dff_A_uUAeA6aC8_0(.dout(w_dff_A_3BVRq0st5_0),.din(w_dff_A_uUAeA6aC8_0),.clk(gclk));
	jdff dff_A_3BVRq0st5_0(.dout(w_dff_A_qx9WmvKS0_0),.din(w_dff_A_3BVRq0st5_0),.clk(gclk));
	jdff dff_A_qx9WmvKS0_0(.dout(w_dff_A_e60Q0Gj75_0),.din(w_dff_A_qx9WmvKS0_0),.clk(gclk));
	jdff dff_A_e60Q0Gj75_0(.dout(G552),.din(w_dff_A_e60Q0Gj75_0),.clk(gclk));
	jdff dff_A_puMfuoYc7_1(.dout(w_dff_A_pmnPc5h48_0),.din(w_dff_A_puMfuoYc7_1),.clk(gclk));
	jdff dff_A_pmnPc5h48_0(.dout(w_dff_A_aBHWQcLr9_0),.din(w_dff_A_pmnPc5h48_0),.clk(gclk));
	jdff dff_A_aBHWQcLr9_0(.dout(w_dff_A_C68e9Zjy5_0),.din(w_dff_A_aBHWQcLr9_0),.clk(gclk));
	jdff dff_A_C68e9Zjy5_0(.dout(w_dff_A_GTCLMMJE9_0),.din(w_dff_A_C68e9Zjy5_0),.clk(gclk));
	jdff dff_A_GTCLMMJE9_0(.dout(w_dff_A_I2vpgGa29_0),.din(w_dff_A_GTCLMMJE9_0),.clk(gclk));
	jdff dff_A_I2vpgGa29_0(.dout(w_dff_A_tQdzbWnE9_0),.din(w_dff_A_I2vpgGa29_0),.clk(gclk));
	jdff dff_A_tQdzbWnE9_0(.dout(w_dff_A_Llpzg4Xh7_0),.din(w_dff_A_tQdzbWnE9_0),.clk(gclk));
	jdff dff_A_Llpzg4Xh7_0(.dout(w_dff_A_qZo5rroK9_0),.din(w_dff_A_Llpzg4Xh7_0),.clk(gclk));
	jdff dff_A_qZo5rroK9_0(.dout(w_dff_A_yFkLVq7c6_0),.din(w_dff_A_qZo5rroK9_0),.clk(gclk));
	jdff dff_A_yFkLVq7c6_0(.dout(w_dff_A_ksjhtiKw1_0),.din(w_dff_A_yFkLVq7c6_0),.clk(gclk));
	jdff dff_A_ksjhtiKw1_0(.dout(w_dff_A_XJhfglIC7_0),.din(w_dff_A_ksjhtiKw1_0),.clk(gclk));
	jdff dff_A_XJhfglIC7_0(.dout(w_dff_A_h9e6mIHC0_0),.din(w_dff_A_XJhfglIC7_0),.clk(gclk));
	jdff dff_A_h9e6mIHC0_0(.dout(w_dff_A_x9Hqfv1A4_0),.din(w_dff_A_h9e6mIHC0_0),.clk(gclk));
	jdff dff_A_x9Hqfv1A4_0(.dout(w_dff_A_hqgkOqdv3_0),.din(w_dff_A_x9Hqfv1A4_0),.clk(gclk));
	jdff dff_A_hqgkOqdv3_0(.dout(w_dff_A_hnluwi503_0),.din(w_dff_A_hqgkOqdv3_0),.clk(gclk));
	jdff dff_A_hnluwi503_0(.dout(w_dff_A_CjG9sA1S8_0),.din(w_dff_A_hnluwi503_0),.clk(gclk));
	jdff dff_A_CjG9sA1S8_0(.dout(w_dff_A_r20o283g3_0),.din(w_dff_A_CjG9sA1S8_0),.clk(gclk));
	jdff dff_A_r20o283g3_0(.dout(w_dff_A_O1KXQbKG0_0),.din(w_dff_A_r20o283g3_0),.clk(gclk));
	jdff dff_A_O1KXQbKG0_0(.dout(w_dff_A_aeYwBjJS7_0),.din(w_dff_A_O1KXQbKG0_0),.clk(gclk));
	jdff dff_A_aeYwBjJS7_0(.dout(w_dff_A_Krojhl2E2_0),.din(w_dff_A_aeYwBjJS7_0),.clk(gclk));
	jdff dff_A_Krojhl2E2_0(.dout(w_dff_A_wladRYMI2_0),.din(w_dff_A_Krojhl2E2_0),.clk(gclk));
	jdff dff_A_wladRYMI2_0(.dout(w_dff_A_CdFHsTjf5_0),.din(w_dff_A_wladRYMI2_0),.clk(gclk));
	jdff dff_A_CdFHsTjf5_0(.dout(w_dff_A_gOVZkuNo0_0),.din(w_dff_A_CdFHsTjf5_0),.clk(gclk));
	jdff dff_A_gOVZkuNo0_0(.dout(w_dff_A_HT8prmZC8_0),.din(w_dff_A_gOVZkuNo0_0),.clk(gclk));
	jdff dff_A_HT8prmZC8_0(.dout(w_dff_A_IDn74baS5_0),.din(w_dff_A_HT8prmZC8_0),.clk(gclk));
	jdff dff_A_IDn74baS5_0(.dout(w_dff_A_UxV47m7T2_0),.din(w_dff_A_IDn74baS5_0),.clk(gclk));
	jdff dff_A_UxV47m7T2_0(.dout(G550),.din(w_dff_A_UxV47m7T2_0),.clk(gclk));
	jdff dff_A_Zq66Xln94_1(.dout(w_dff_A_k912QvlV9_0),.din(w_dff_A_Zq66Xln94_1),.clk(gclk));
	jdff dff_A_k912QvlV9_0(.dout(w_dff_A_JDVWLYkO3_0),.din(w_dff_A_k912QvlV9_0),.clk(gclk));
	jdff dff_A_JDVWLYkO3_0(.dout(w_dff_A_UZy8oTVM4_0),.din(w_dff_A_JDVWLYkO3_0),.clk(gclk));
	jdff dff_A_UZy8oTVM4_0(.dout(w_dff_A_kFtPJFQr4_0),.din(w_dff_A_UZy8oTVM4_0),.clk(gclk));
	jdff dff_A_kFtPJFQr4_0(.dout(w_dff_A_zIMye9rk6_0),.din(w_dff_A_kFtPJFQr4_0),.clk(gclk));
	jdff dff_A_zIMye9rk6_0(.dout(w_dff_A_mToo5dkM1_0),.din(w_dff_A_zIMye9rk6_0),.clk(gclk));
	jdff dff_A_mToo5dkM1_0(.dout(w_dff_A_l2BcZYmm0_0),.din(w_dff_A_mToo5dkM1_0),.clk(gclk));
	jdff dff_A_l2BcZYmm0_0(.dout(w_dff_A_MSwxwvR52_0),.din(w_dff_A_l2BcZYmm0_0),.clk(gclk));
	jdff dff_A_MSwxwvR52_0(.dout(w_dff_A_6l7HzzmG6_0),.din(w_dff_A_MSwxwvR52_0),.clk(gclk));
	jdff dff_A_6l7HzzmG6_0(.dout(w_dff_A_QN0khxl39_0),.din(w_dff_A_6l7HzzmG6_0),.clk(gclk));
	jdff dff_A_QN0khxl39_0(.dout(w_dff_A_29wWV7m68_0),.din(w_dff_A_QN0khxl39_0),.clk(gclk));
	jdff dff_A_29wWV7m68_0(.dout(w_dff_A_MCAWVTKd1_0),.din(w_dff_A_29wWV7m68_0),.clk(gclk));
	jdff dff_A_MCAWVTKd1_0(.dout(w_dff_A_pDnqd1NK9_0),.din(w_dff_A_MCAWVTKd1_0),.clk(gclk));
	jdff dff_A_pDnqd1NK9_0(.dout(w_dff_A_uZDFHRXA0_0),.din(w_dff_A_pDnqd1NK9_0),.clk(gclk));
	jdff dff_A_uZDFHRXA0_0(.dout(w_dff_A_Hf6hh8u79_0),.din(w_dff_A_uZDFHRXA0_0),.clk(gclk));
	jdff dff_A_Hf6hh8u79_0(.dout(w_dff_A_e16w1sRj6_0),.din(w_dff_A_Hf6hh8u79_0),.clk(gclk));
	jdff dff_A_e16w1sRj6_0(.dout(w_dff_A_mz0zHQ308_0),.din(w_dff_A_e16w1sRj6_0),.clk(gclk));
	jdff dff_A_mz0zHQ308_0(.dout(w_dff_A_mTtOyiuh8_0),.din(w_dff_A_mz0zHQ308_0),.clk(gclk));
	jdff dff_A_mTtOyiuh8_0(.dout(w_dff_A_L4xd6kf04_0),.din(w_dff_A_mTtOyiuh8_0),.clk(gclk));
	jdff dff_A_L4xd6kf04_0(.dout(w_dff_A_tMj5Ac5K4_0),.din(w_dff_A_L4xd6kf04_0),.clk(gclk));
	jdff dff_A_tMj5Ac5K4_0(.dout(w_dff_A_yDuHrXsz0_0),.din(w_dff_A_tMj5Ac5K4_0),.clk(gclk));
	jdff dff_A_yDuHrXsz0_0(.dout(w_dff_A_D3ngKS0I9_0),.din(w_dff_A_yDuHrXsz0_0),.clk(gclk));
	jdff dff_A_D3ngKS0I9_0(.dout(w_dff_A_n3n1o1sq7_0),.din(w_dff_A_D3ngKS0I9_0),.clk(gclk));
	jdff dff_A_n3n1o1sq7_0(.dout(w_dff_A_2GW4XwH87_0),.din(w_dff_A_n3n1o1sq7_0),.clk(gclk));
	jdff dff_A_2GW4XwH87_0(.dout(w_dff_A_aAstr5y95_0),.din(w_dff_A_2GW4XwH87_0),.clk(gclk));
	jdff dff_A_aAstr5y95_0(.dout(w_dff_A_KXsfjgmM0_0),.din(w_dff_A_aAstr5y95_0),.clk(gclk));
	jdff dff_A_KXsfjgmM0_0(.dout(G548),.din(w_dff_A_KXsfjgmM0_0),.clk(gclk));
	jdff dff_A_DDaoXkJA6_1(.dout(w_dff_A_7uPgKn8s1_0),.din(w_dff_A_DDaoXkJA6_1),.clk(gclk));
	jdff dff_A_7uPgKn8s1_0(.dout(w_dff_A_R9PqNNcb8_0),.din(w_dff_A_7uPgKn8s1_0),.clk(gclk));
	jdff dff_A_R9PqNNcb8_0(.dout(w_dff_A_4wer1PBI5_0),.din(w_dff_A_R9PqNNcb8_0),.clk(gclk));
	jdff dff_A_4wer1PBI5_0(.dout(w_dff_A_H9h25ZeW8_0),.din(w_dff_A_4wer1PBI5_0),.clk(gclk));
	jdff dff_A_H9h25ZeW8_0(.dout(w_dff_A_7Yg1dQTv9_0),.din(w_dff_A_H9h25ZeW8_0),.clk(gclk));
	jdff dff_A_7Yg1dQTv9_0(.dout(w_dff_A_BX4u5fLA2_0),.din(w_dff_A_7Yg1dQTv9_0),.clk(gclk));
	jdff dff_A_BX4u5fLA2_0(.dout(w_dff_A_nvPrDDjS7_0),.din(w_dff_A_BX4u5fLA2_0),.clk(gclk));
	jdff dff_A_nvPrDDjS7_0(.dout(w_dff_A_RS0yCt0l4_0),.din(w_dff_A_nvPrDDjS7_0),.clk(gclk));
	jdff dff_A_RS0yCt0l4_0(.dout(w_dff_A_UozTiDTO2_0),.din(w_dff_A_RS0yCt0l4_0),.clk(gclk));
	jdff dff_A_UozTiDTO2_0(.dout(w_dff_A_JfCAGHWD6_0),.din(w_dff_A_UozTiDTO2_0),.clk(gclk));
	jdff dff_A_JfCAGHWD6_0(.dout(w_dff_A_mJYsnTG26_0),.din(w_dff_A_JfCAGHWD6_0),.clk(gclk));
	jdff dff_A_mJYsnTG26_0(.dout(w_dff_A_TBI6YeTV5_0),.din(w_dff_A_mJYsnTG26_0),.clk(gclk));
	jdff dff_A_TBI6YeTV5_0(.dout(w_dff_A_AcpUpPxQ2_0),.din(w_dff_A_TBI6YeTV5_0),.clk(gclk));
	jdff dff_A_AcpUpPxQ2_0(.dout(w_dff_A_q3l5svan7_0),.din(w_dff_A_AcpUpPxQ2_0),.clk(gclk));
	jdff dff_A_q3l5svan7_0(.dout(w_dff_A_IECtLNfC7_0),.din(w_dff_A_q3l5svan7_0),.clk(gclk));
	jdff dff_A_IECtLNfC7_0(.dout(w_dff_A_m2XGcXWk1_0),.din(w_dff_A_IECtLNfC7_0),.clk(gclk));
	jdff dff_A_m2XGcXWk1_0(.dout(w_dff_A_93thysza7_0),.din(w_dff_A_m2XGcXWk1_0),.clk(gclk));
	jdff dff_A_93thysza7_0(.dout(w_dff_A_Y0xtZ38t1_0),.din(w_dff_A_93thysza7_0),.clk(gclk));
	jdff dff_A_Y0xtZ38t1_0(.dout(w_dff_A_8hYapcuP6_0),.din(w_dff_A_Y0xtZ38t1_0),.clk(gclk));
	jdff dff_A_8hYapcuP6_0(.dout(w_dff_A_24F6oHqj8_0),.din(w_dff_A_8hYapcuP6_0),.clk(gclk));
	jdff dff_A_24F6oHqj8_0(.dout(w_dff_A_5uo41Vol4_0),.din(w_dff_A_24F6oHqj8_0),.clk(gclk));
	jdff dff_A_5uo41Vol4_0(.dout(w_dff_A_JBEVRVV80_0),.din(w_dff_A_5uo41Vol4_0),.clk(gclk));
	jdff dff_A_JBEVRVV80_0(.dout(w_dff_A_ddrsVdYQ1_0),.din(w_dff_A_JBEVRVV80_0),.clk(gclk));
	jdff dff_A_ddrsVdYQ1_0(.dout(w_dff_A_7GF6ZAcv3_0),.din(w_dff_A_ddrsVdYQ1_0),.clk(gclk));
	jdff dff_A_7GF6ZAcv3_0(.dout(w_dff_A_5AwN8fNi3_0),.din(w_dff_A_7GF6ZAcv3_0),.clk(gclk));
	jdff dff_A_5AwN8fNi3_0(.dout(w_dff_A_rB18fipo2_0),.din(w_dff_A_5AwN8fNi3_0),.clk(gclk));
	jdff dff_A_rB18fipo2_0(.dout(G546),.din(w_dff_A_rB18fipo2_0),.clk(gclk));
	jdff dff_A_YECV73dN5_1(.dout(w_dff_A_p6HRyqvL5_0),.din(w_dff_A_YECV73dN5_1),.clk(gclk));
	jdff dff_A_p6HRyqvL5_0(.dout(w_dff_A_HHLGkS7H2_0),.din(w_dff_A_p6HRyqvL5_0),.clk(gclk));
	jdff dff_A_HHLGkS7H2_0(.dout(w_dff_A_DWFMMH563_0),.din(w_dff_A_HHLGkS7H2_0),.clk(gclk));
	jdff dff_A_DWFMMH563_0(.dout(w_dff_A_6LUERjae3_0),.din(w_dff_A_DWFMMH563_0),.clk(gclk));
	jdff dff_A_6LUERjae3_0(.dout(w_dff_A_rdv0ugAc8_0),.din(w_dff_A_6LUERjae3_0),.clk(gclk));
	jdff dff_A_rdv0ugAc8_0(.dout(w_dff_A_PyidGCmK2_0),.din(w_dff_A_rdv0ugAc8_0),.clk(gclk));
	jdff dff_A_PyidGCmK2_0(.dout(w_dff_A_cBJpMe1Z6_0),.din(w_dff_A_PyidGCmK2_0),.clk(gclk));
	jdff dff_A_cBJpMe1Z6_0(.dout(w_dff_A_Z4x7Vb2R6_0),.din(w_dff_A_cBJpMe1Z6_0),.clk(gclk));
	jdff dff_A_Z4x7Vb2R6_0(.dout(w_dff_A_JUWoiqKm1_0),.din(w_dff_A_Z4x7Vb2R6_0),.clk(gclk));
	jdff dff_A_JUWoiqKm1_0(.dout(w_dff_A_7S72pRih8_0),.din(w_dff_A_JUWoiqKm1_0),.clk(gclk));
	jdff dff_A_7S72pRih8_0(.dout(w_dff_A_ONwUSsQr5_0),.din(w_dff_A_7S72pRih8_0),.clk(gclk));
	jdff dff_A_ONwUSsQr5_0(.dout(w_dff_A_60NfhBHI5_0),.din(w_dff_A_ONwUSsQr5_0),.clk(gclk));
	jdff dff_A_60NfhBHI5_0(.dout(w_dff_A_uqwKGK1x7_0),.din(w_dff_A_60NfhBHI5_0),.clk(gclk));
	jdff dff_A_uqwKGK1x7_0(.dout(w_dff_A_AZFr2EUz2_0),.din(w_dff_A_uqwKGK1x7_0),.clk(gclk));
	jdff dff_A_AZFr2EUz2_0(.dout(w_dff_A_kBtBVXNo6_0),.din(w_dff_A_AZFr2EUz2_0),.clk(gclk));
	jdff dff_A_kBtBVXNo6_0(.dout(w_dff_A_5tIJVuTk2_0),.din(w_dff_A_kBtBVXNo6_0),.clk(gclk));
	jdff dff_A_5tIJVuTk2_0(.dout(w_dff_A_LmQwbT5r8_0),.din(w_dff_A_5tIJVuTk2_0),.clk(gclk));
	jdff dff_A_LmQwbT5r8_0(.dout(w_dff_A_aBRXscI79_0),.din(w_dff_A_LmQwbT5r8_0),.clk(gclk));
	jdff dff_A_aBRXscI79_0(.dout(w_dff_A_DSjUA1kS3_0),.din(w_dff_A_aBRXscI79_0),.clk(gclk));
	jdff dff_A_DSjUA1kS3_0(.dout(w_dff_A_i1qy4bcu6_0),.din(w_dff_A_DSjUA1kS3_0),.clk(gclk));
	jdff dff_A_i1qy4bcu6_0(.dout(w_dff_A_XOFoBH051_0),.din(w_dff_A_i1qy4bcu6_0),.clk(gclk));
	jdff dff_A_XOFoBH051_0(.dout(w_dff_A_ZkXE4HVC4_0),.din(w_dff_A_XOFoBH051_0),.clk(gclk));
	jdff dff_A_ZkXE4HVC4_0(.dout(w_dff_A_OiBHMBkw4_0),.din(w_dff_A_ZkXE4HVC4_0),.clk(gclk));
	jdff dff_A_OiBHMBkw4_0(.dout(w_dff_A_vrl2u6ps1_0),.din(w_dff_A_OiBHMBkw4_0),.clk(gclk));
	jdff dff_A_vrl2u6ps1_0(.dout(w_dff_A_DJePysRw1_0),.din(w_dff_A_vrl2u6ps1_0),.clk(gclk));
	jdff dff_A_DJePysRw1_0(.dout(w_dff_A_PwWKa3ae2_0),.din(w_dff_A_DJePysRw1_0),.clk(gclk));
	jdff dff_A_PwWKa3ae2_0(.dout(G544),.din(w_dff_A_PwWKa3ae2_0),.clk(gclk));
	jdff dff_A_9XjXRFMW1_1(.dout(w_dff_A_AoUmo7h10_0),.din(w_dff_A_9XjXRFMW1_1),.clk(gclk));
	jdff dff_A_AoUmo7h10_0(.dout(w_dff_A_FrxE5A4p6_0),.din(w_dff_A_AoUmo7h10_0),.clk(gclk));
	jdff dff_A_FrxE5A4p6_0(.dout(w_dff_A_UdHgtBIZ3_0),.din(w_dff_A_FrxE5A4p6_0),.clk(gclk));
	jdff dff_A_UdHgtBIZ3_0(.dout(w_dff_A_lHZHKMWD3_0),.din(w_dff_A_UdHgtBIZ3_0),.clk(gclk));
	jdff dff_A_lHZHKMWD3_0(.dout(w_dff_A_KlvwRLCr0_0),.din(w_dff_A_lHZHKMWD3_0),.clk(gclk));
	jdff dff_A_KlvwRLCr0_0(.dout(w_dff_A_qoNARPjP1_0),.din(w_dff_A_KlvwRLCr0_0),.clk(gclk));
	jdff dff_A_qoNARPjP1_0(.dout(w_dff_A_y4jI1la98_0),.din(w_dff_A_qoNARPjP1_0),.clk(gclk));
	jdff dff_A_y4jI1la98_0(.dout(w_dff_A_f2EUylyZ9_0),.din(w_dff_A_y4jI1la98_0),.clk(gclk));
	jdff dff_A_f2EUylyZ9_0(.dout(w_dff_A_qhh83PyN0_0),.din(w_dff_A_f2EUylyZ9_0),.clk(gclk));
	jdff dff_A_qhh83PyN0_0(.dout(w_dff_A_N3RzjaRJ4_0),.din(w_dff_A_qhh83PyN0_0),.clk(gclk));
	jdff dff_A_N3RzjaRJ4_0(.dout(w_dff_A_IgKW3cWW5_0),.din(w_dff_A_N3RzjaRJ4_0),.clk(gclk));
	jdff dff_A_IgKW3cWW5_0(.dout(w_dff_A_lDlx0eDO9_0),.din(w_dff_A_IgKW3cWW5_0),.clk(gclk));
	jdff dff_A_lDlx0eDO9_0(.dout(w_dff_A_H6cN5fG00_0),.din(w_dff_A_lDlx0eDO9_0),.clk(gclk));
	jdff dff_A_H6cN5fG00_0(.dout(w_dff_A_cm5z690o8_0),.din(w_dff_A_H6cN5fG00_0),.clk(gclk));
	jdff dff_A_cm5z690o8_0(.dout(w_dff_A_codDEp5I4_0),.din(w_dff_A_cm5z690o8_0),.clk(gclk));
	jdff dff_A_codDEp5I4_0(.dout(w_dff_A_IAWee61O5_0),.din(w_dff_A_codDEp5I4_0),.clk(gclk));
	jdff dff_A_IAWee61O5_0(.dout(w_dff_A_OxwJpBWY7_0),.din(w_dff_A_IAWee61O5_0),.clk(gclk));
	jdff dff_A_OxwJpBWY7_0(.dout(w_dff_A_m6Dj9tEO0_0),.din(w_dff_A_OxwJpBWY7_0),.clk(gclk));
	jdff dff_A_m6Dj9tEO0_0(.dout(w_dff_A_Xn8SI23c7_0),.din(w_dff_A_m6Dj9tEO0_0),.clk(gclk));
	jdff dff_A_Xn8SI23c7_0(.dout(w_dff_A_MrwHxCFr2_0),.din(w_dff_A_Xn8SI23c7_0),.clk(gclk));
	jdff dff_A_MrwHxCFr2_0(.dout(w_dff_A_RIcbXtz61_0),.din(w_dff_A_MrwHxCFr2_0),.clk(gclk));
	jdff dff_A_RIcbXtz61_0(.dout(w_dff_A_HCwZUYPN8_0),.din(w_dff_A_RIcbXtz61_0),.clk(gclk));
	jdff dff_A_HCwZUYPN8_0(.dout(w_dff_A_WY14eKx50_0),.din(w_dff_A_HCwZUYPN8_0),.clk(gclk));
	jdff dff_A_WY14eKx50_0(.dout(w_dff_A_jKwzFe9f8_0),.din(w_dff_A_WY14eKx50_0),.clk(gclk));
	jdff dff_A_jKwzFe9f8_0(.dout(w_dff_A_PvlRxVMa5_0),.din(w_dff_A_jKwzFe9f8_0),.clk(gclk));
	jdff dff_A_PvlRxVMa5_0(.dout(w_dff_A_mWbi3MvK5_0),.din(w_dff_A_PvlRxVMa5_0),.clk(gclk));
	jdff dff_A_mWbi3MvK5_0(.dout(G540),.din(w_dff_A_mWbi3MvK5_0),.clk(gclk));
	jdff dff_A_oNY1Iu5k2_1(.dout(w_dff_A_3ygRFRxZ4_0),.din(w_dff_A_oNY1Iu5k2_1),.clk(gclk));
	jdff dff_A_3ygRFRxZ4_0(.dout(w_dff_A_J3t9Owan0_0),.din(w_dff_A_3ygRFRxZ4_0),.clk(gclk));
	jdff dff_A_J3t9Owan0_0(.dout(w_dff_A_ggriSJyQ2_0),.din(w_dff_A_J3t9Owan0_0),.clk(gclk));
	jdff dff_A_ggriSJyQ2_0(.dout(w_dff_A_HKErTrDQ9_0),.din(w_dff_A_ggriSJyQ2_0),.clk(gclk));
	jdff dff_A_HKErTrDQ9_0(.dout(w_dff_A_nJfkujWH1_0),.din(w_dff_A_HKErTrDQ9_0),.clk(gclk));
	jdff dff_A_nJfkujWH1_0(.dout(w_dff_A_tqaqhby31_0),.din(w_dff_A_nJfkujWH1_0),.clk(gclk));
	jdff dff_A_tqaqhby31_0(.dout(w_dff_A_1xfJCtFC3_0),.din(w_dff_A_tqaqhby31_0),.clk(gclk));
	jdff dff_A_1xfJCtFC3_0(.dout(w_dff_A_Q3A6fB6d8_0),.din(w_dff_A_1xfJCtFC3_0),.clk(gclk));
	jdff dff_A_Q3A6fB6d8_0(.dout(w_dff_A_ukLxuOnf8_0),.din(w_dff_A_Q3A6fB6d8_0),.clk(gclk));
	jdff dff_A_ukLxuOnf8_0(.dout(w_dff_A_vAbD0RGV7_0),.din(w_dff_A_ukLxuOnf8_0),.clk(gclk));
	jdff dff_A_vAbD0RGV7_0(.dout(w_dff_A_6hCQc7Mr5_0),.din(w_dff_A_vAbD0RGV7_0),.clk(gclk));
	jdff dff_A_6hCQc7Mr5_0(.dout(w_dff_A_J4KLCAFv7_0),.din(w_dff_A_6hCQc7Mr5_0),.clk(gclk));
	jdff dff_A_J4KLCAFv7_0(.dout(w_dff_A_J8C7zaQw3_0),.din(w_dff_A_J4KLCAFv7_0),.clk(gclk));
	jdff dff_A_J8C7zaQw3_0(.dout(w_dff_A_htoNZU9T9_0),.din(w_dff_A_J8C7zaQw3_0),.clk(gclk));
	jdff dff_A_htoNZU9T9_0(.dout(w_dff_A_Fl3z1Gvv5_0),.din(w_dff_A_htoNZU9T9_0),.clk(gclk));
	jdff dff_A_Fl3z1Gvv5_0(.dout(w_dff_A_4BknDiRD4_0),.din(w_dff_A_Fl3z1Gvv5_0),.clk(gclk));
	jdff dff_A_4BknDiRD4_0(.dout(w_dff_A_ct70PNLr9_0),.din(w_dff_A_4BknDiRD4_0),.clk(gclk));
	jdff dff_A_ct70PNLr9_0(.dout(w_dff_A_leMRrTmm6_0),.din(w_dff_A_ct70PNLr9_0),.clk(gclk));
	jdff dff_A_leMRrTmm6_0(.dout(w_dff_A_flGKh7kk5_0),.din(w_dff_A_leMRrTmm6_0),.clk(gclk));
	jdff dff_A_flGKh7kk5_0(.dout(w_dff_A_l4gcUjJS5_0),.din(w_dff_A_flGKh7kk5_0),.clk(gclk));
	jdff dff_A_l4gcUjJS5_0(.dout(w_dff_A_rZVWJr572_0),.din(w_dff_A_l4gcUjJS5_0),.clk(gclk));
	jdff dff_A_rZVWJr572_0(.dout(w_dff_A_srPGCgnv0_0),.din(w_dff_A_rZVWJr572_0),.clk(gclk));
	jdff dff_A_srPGCgnv0_0(.dout(w_dff_A_eMhCmY6B5_0),.din(w_dff_A_srPGCgnv0_0),.clk(gclk));
	jdff dff_A_eMhCmY6B5_0(.dout(w_dff_A_5AnLIGkc5_0),.din(w_dff_A_eMhCmY6B5_0),.clk(gclk));
	jdff dff_A_5AnLIGkc5_0(.dout(w_dff_A_itE0S7pK2_0),.din(w_dff_A_5AnLIGkc5_0),.clk(gclk));
	jdff dff_A_itE0S7pK2_0(.dout(w_dff_A_pBF4rZ0k0_0),.din(w_dff_A_itE0S7pK2_0),.clk(gclk));
	jdff dff_A_pBF4rZ0k0_0(.dout(G538),.din(w_dff_A_pBF4rZ0k0_0),.clk(gclk));
	jdff dff_A_A7hwHenU7_1(.dout(w_dff_A_mY29OrUp4_0),.din(w_dff_A_A7hwHenU7_1),.clk(gclk));
	jdff dff_A_mY29OrUp4_0(.dout(w_dff_A_31r5hcBQ9_0),.din(w_dff_A_mY29OrUp4_0),.clk(gclk));
	jdff dff_A_31r5hcBQ9_0(.dout(w_dff_A_wJIocf6w0_0),.din(w_dff_A_31r5hcBQ9_0),.clk(gclk));
	jdff dff_A_wJIocf6w0_0(.dout(w_dff_A_MAmOy4hl2_0),.din(w_dff_A_wJIocf6w0_0),.clk(gclk));
	jdff dff_A_MAmOy4hl2_0(.dout(w_dff_A_63qWM3Pk8_0),.din(w_dff_A_MAmOy4hl2_0),.clk(gclk));
	jdff dff_A_63qWM3Pk8_0(.dout(w_dff_A_7oNoLsoJ9_0),.din(w_dff_A_63qWM3Pk8_0),.clk(gclk));
	jdff dff_A_7oNoLsoJ9_0(.dout(w_dff_A_4VE4d1ar9_0),.din(w_dff_A_7oNoLsoJ9_0),.clk(gclk));
	jdff dff_A_4VE4d1ar9_0(.dout(w_dff_A_NupIPhb90_0),.din(w_dff_A_4VE4d1ar9_0),.clk(gclk));
	jdff dff_A_NupIPhb90_0(.dout(w_dff_A_lpVs4XQl0_0),.din(w_dff_A_NupIPhb90_0),.clk(gclk));
	jdff dff_A_lpVs4XQl0_0(.dout(w_dff_A_1DjMUDJ22_0),.din(w_dff_A_lpVs4XQl0_0),.clk(gclk));
	jdff dff_A_1DjMUDJ22_0(.dout(w_dff_A_K0FtxPjW5_0),.din(w_dff_A_1DjMUDJ22_0),.clk(gclk));
	jdff dff_A_K0FtxPjW5_0(.dout(w_dff_A_DB5N1ORG7_0),.din(w_dff_A_K0FtxPjW5_0),.clk(gclk));
	jdff dff_A_DB5N1ORG7_0(.dout(w_dff_A_FMxxLnl60_0),.din(w_dff_A_DB5N1ORG7_0),.clk(gclk));
	jdff dff_A_FMxxLnl60_0(.dout(w_dff_A_bGETVDBm9_0),.din(w_dff_A_FMxxLnl60_0),.clk(gclk));
	jdff dff_A_bGETVDBm9_0(.dout(w_dff_A_vrQUpQ849_0),.din(w_dff_A_bGETVDBm9_0),.clk(gclk));
	jdff dff_A_vrQUpQ849_0(.dout(w_dff_A_nvjl7GsZ5_0),.din(w_dff_A_vrQUpQ849_0),.clk(gclk));
	jdff dff_A_nvjl7GsZ5_0(.dout(w_dff_A_2Rb93uy34_0),.din(w_dff_A_nvjl7GsZ5_0),.clk(gclk));
	jdff dff_A_2Rb93uy34_0(.dout(w_dff_A_2Bt7Ot1C7_0),.din(w_dff_A_2Rb93uy34_0),.clk(gclk));
	jdff dff_A_2Bt7Ot1C7_0(.dout(w_dff_A_svUEaiP50_0),.din(w_dff_A_2Bt7Ot1C7_0),.clk(gclk));
	jdff dff_A_svUEaiP50_0(.dout(w_dff_A_dNhxAr2S8_0),.din(w_dff_A_svUEaiP50_0),.clk(gclk));
	jdff dff_A_dNhxAr2S8_0(.dout(w_dff_A_d1bcCcJi4_0),.din(w_dff_A_dNhxAr2S8_0),.clk(gclk));
	jdff dff_A_d1bcCcJi4_0(.dout(w_dff_A_1CZvWQSm7_0),.din(w_dff_A_d1bcCcJi4_0),.clk(gclk));
	jdff dff_A_1CZvWQSm7_0(.dout(w_dff_A_S0g7mT5z8_0),.din(w_dff_A_1CZvWQSm7_0),.clk(gclk));
	jdff dff_A_S0g7mT5z8_0(.dout(w_dff_A_PimE1lvm5_0),.din(w_dff_A_S0g7mT5z8_0),.clk(gclk));
	jdff dff_A_PimE1lvm5_0(.dout(w_dff_A_T7SYX85T2_0),.din(w_dff_A_PimE1lvm5_0),.clk(gclk));
	jdff dff_A_T7SYX85T2_0(.dout(w_dff_A_M11ZEwKf4_0),.din(w_dff_A_T7SYX85T2_0),.clk(gclk));
	jdff dff_A_M11ZEwKf4_0(.dout(G536),.din(w_dff_A_M11ZEwKf4_0),.clk(gclk));
	jdff dff_A_5NPOVR0c6_1(.dout(w_dff_A_kedJpPF42_0),.din(w_dff_A_5NPOVR0c6_1),.clk(gclk));
	jdff dff_A_kedJpPF42_0(.dout(w_dff_A_hXvorjZe9_0),.din(w_dff_A_kedJpPF42_0),.clk(gclk));
	jdff dff_A_hXvorjZe9_0(.dout(w_dff_A_5SdqaOmZ9_0),.din(w_dff_A_hXvorjZe9_0),.clk(gclk));
	jdff dff_A_5SdqaOmZ9_0(.dout(w_dff_A_yqYBKEO11_0),.din(w_dff_A_5SdqaOmZ9_0),.clk(gclk));
	jdff dff_A_yqYBKEO11_0(.dout(w_dff_A_ErwYmcM25_0),.din(w_dff_A_yqYBKEO11_0),.clk(gclk));
	jdff dff_A_ErwYmcM25_0(.dout(w_dff_A_9dg5GZsc4_0),.din(w_dff_A_ErwYmcM25_0),.clk(gclk));
	jdff dff_A_9dg5GZsc4_0(.dout(w_dff_A_nqLbCdKB5_0),.din(w_dff_A_9dg5GZsc4_0),.clk(gclk));
	jdff dff_A_nqLbCdKB5_0(.dout(w_dff_A_gAHekINO4_0),.din(w_dff_A_nqLbCdKB5_0),.clk(gclk));
	jdff dff_A_gAHekINO4_0(.dout(w_dff_A_AJAY8mQs6_0),.din(w_dff_A_gAHekINO4_0),.clk(gclk));
	jdff dff_A_AJAY8mQs6_0(.dout(w_dff_A_HTskUTgm7_0),.din(w_dff_A_AJAY8mQs6_0),.clk(gclk));
	jdff dff_A_HTskUTgm7_0(.dout(w_dff_A_9EhZHAuz8_0),.din(w_dff_A_HTskUTgm7_0),.clk(gclk));
	jdff dff_A_9EhZHAuz8_0(.dout(w_dff_A_AAZVSc7z6_0),.din(w_dff_A_9EhZHAuz8_0),.clk(gclk));
	jdff dff_A_AAZVSc7z6_0(.dout(w_dff_A_qgevseyZ0_0),.din(w_dff_A_AAZVSc7z6_0),.clk(gclk));
	jdff dff_A_qgevseyZ0_0(.dout(w_dff_A_SnCrtqNN6_0),.din(w_dff_A_qgevseyZ0_0),.clk(gclk));
	jdff dff_A_SnCrtqNN6_0(.dout(w_dff_A_K5nXN7co7_0),.din(w_dff_A_SnCrtqNN6_0),.clk(gclk));
	jdff dff_A_K5nXN7co7_0(.dout(w_dff_A_NsCGsO2B0_0),.din(w_dff_A_K5nXN7co7_0),.clk(gclk));
	jdff dff_A_NsCGsO2B0_0(.dout(w_dff_A_nMPmUtWn1_0),.din(w_dff_A_NsCGsO2B0_0),.clk(gclk));
	jdff dff_A_nMPmUtWn1_0(.dout(w_dff_A_60JdOhcx9_0),.din(w_dff_A_nMPmUtWn1_0),.clk(gclk));
	jdff dff_A_60JdOhcx9_0(.dout(w_dff_A_EP2NLLMm1_0),.din(w_dff_A_60JdOhcx9_0),.clk(gclk));
	jdff dff_A_EP2NLLMm1_0(.dout(w_dff_A_P8wM2yDM1_0),.din(w_dff_A_EP2NLLMm1_0),.clk(gclk));
	jdff dff_A_P8wM2yDM1_0(.dout(w_dff_A_xrwBTyES9_0),.din(w_dff_A_P8wM2yDM1_0),.clk(gclk));
	jdff dff_A_xrwBTyES9_0(.dout(w_dff_A_m2AgbVBL1_0),.din(w_dff_A_xrwBTyES9_0),.clk(gclk));
	jdff dff_A_m2AgbVBL1_0(.dout(w_dff_A_22kH0UT49_0),.din(w_dff_A_m2AgbVBL1_0),.clk(gclk));
	jdff dff_A_22kH0UT49_0(.dout(w_dff_A_9c6o8sG65_0),.din(w_dff_A_22kH0UT49_0),.clk(gclk));
	jdff dff_A_9c6o8sG65_0(.dout(w_dff_A_IDtfuMVe4_0),.din(w_dff_A_9c6o8sG65_0),.clk(gclk));
	jdff dff_A_IDtfuMVe4_0(.dout(w_dff_A_CldaB4NW2_0),.din(w_dff_A_IDtfuMVe4_0),.clk(gclk));
	jdff dff_A_CldaB4NW2_0(.dout(G534),.din(w_dff_A_CldaB4NW2_0),.clk(gclk));
	jdff dff_A_lE27KfQ80_1(.dout(w_dff_A_IbcGrrkx1_0),.din(w_dff_A_lE27KfQ80_1),.clk(gclk));
	jdff dff_A_IbcGrrkx1_0(.dout(w_dff_A_0Silw3NH3_0),.din(w_dff_A_IbcGrrkx1_0),.clk(gclk));
	jdff dff_A_0Silw3NH3_0(.dout(w_dff_A_8p6ceSdA9_0),.din(w_dff_A_0Silw3NH3_0),.clk(gclk));
	jdff dff_A_8p6ceSdA9_0(.dout(w_dff_A_Z1fCUz068_0),.din(w_dff_A_8p6ceSdA9_0),.clk(gclk));
	jdff dff_A_Z1fCUz068_0(.dout(w_dff_A_8p41aVx76_0),.din(w_dff_A_Z1fCUz068_0),.clk(gclk));
	jdff dff_A_8p41aVx76_0(.dout(w_dff_A_Bnvis7W37_0),.din(w_dff_A_8p41aVx76_0),.clk(gclk));
	jdff dff_A_Bnvis7W37_0(.dout(w_dff_A_kx2HdYFi5_0),.din(w_dff_A_Bnvis7W37_0),.clk(gclk));
	jdff dff_A_kx2HdYFi5_0(.dout(w_dff_A_OxGy5Pi77_0),.din(w_dff_A_kx2HdYFi5_0),.clk(gclk));
	jdff dff_A_OxGy5Pi77_0(.dout(w_dff_A_2c0q00AJ9_0),.din(w_dff_A_OxGy5Pi77_0),.clk(gclk));
	jdff dff_A_2c0q00AJ9_0(.dout(w_dff_A_wXjsufIw8_0),.din(w_dff_A_2c0q00AJ9_0),.clk(gclk));
	jdff dff_A_wXjsufIw8_0(.dout(w_dff_A_6yFE6mpt9_0),.din(w_dff_A_wXjsufIw8_0),.clk(gclk));
	jdff dff_A_6yFE6mpt9_0(.dout(w_dff_A_Nm4AP3zM7_0),.din(w_dff_A_6yFE6mpt9_0),.clk(gclk));
	jdff dff_A_Nm4AP3zM7_0(.dout(w_dff_A_ISCZtJ2D2_0),.din(w_dff_A_Nm4AP3zM7_0),.clk(gclk));
	jdff dff_A_ISCZtJ2D2_0(.dout(w_dff_A_2lZVGOtZ8_0),.din(w_dff_A_ISCZtJ2D2_0),.clk(gclk));
	jdff dff_A_2lZVGOtZ8_0(.dout(w_dff_A_vqQU3vVM5_0),.din(w_dff_A_2lZVGOtZ8_0),.clk(gclk));
	jdff dff_A_vqQU3vVM5_0(.dout(w_dff_A_M7XmWZI61_0),.din(w_dff_A_vqQU3vVM5_0),.clk(gclk));
	jdff dff_A_M7XmWZI61_0(.dout(w_dff_A_BSGBPpLy8_0),.din(w_dff_A_M7XmWZI61_0),.clk(gclk));
	jdff dff_A_BSGBPpLy8_0(.dout(w_dff_A_pGYpMhT88_0),.din(w_dff_A_BSGBPpLy8_0),.clk(gclk));
	jdff dff_A_pGYpMhT88_0(.dout(w_dff_A_hwYNBimw2_0),.din(w_dff_A_pGYpMhT88_0),.clk(gclk));
	jdff dff_A_hwYNBimw2_0(.dout(w_dff_A_AYZKThBq8_0),.din(w_dff_A_hwYNBimw2_0),.clk(gclk));
	jdff dff_A_AYZKThBq8_0(.dout(w_dff_A_E8yAJYQA3_0),.din(w_dff_A_AYZKThBq8_0),.clk(gclk));
	jdff dff_A_E8yAJYQA3_0(.dout(w_dff_A_GXcE2zvF3_0),.din(w_dff_A_E8yAJYQA3_0),.clk(gclk));
	jdff dff_A_GXcE2zvF3_0(.dout(w_dff_A_fLdT3Ohf0_0),.din(w_dff_A_GXcE2zvF3_0),.clk(gclk));
	jdff dff_A_fLdT3Ohf0_0(.dout(w_dff_A_STI1Ss9b1_0),.din(w_dff_A_fLdT3Ohf0_0),.clk(gclk));
	jdff dff_A_STI1Ss9b1_0(.dout(w_dff_A_xShdlbbk2_0),.din(w_dff_A_STI1Ss9b1_0),.clk(gclk));
	jdff dff_A_xShdlbbk2_0(.dout(w_dff_A_IDaEoSGw1_0),.din(w_dff_A_xShdlbbk2_0),.clk(gclk));
	jdff dff_A_IDaEoSGw1_0(.dout(G532),.din(w_dff_A_IDaEoSGw1_0),.clk(gclk));
	jdff dff_A_f8Cco9ft3_1(.dout(w_dff_A_9BNqIGXe7_0),.din(w_dff_A_f8Cco9ft3_1),.clk(gclk));
	jdff dff_A_9BNqIGXe7_0(.dout(w_dff_A_BOXFVgi66_0),.din(w_dff_A_9BNqIGXe7_0),.clk(gclk));
	jdff dff_A_BOXFVgi66_0(.dout(w_dff_A_VlNZvv7n2_0),.din(w_dff_A_BOXFVgi66_0),.clk(gclk));
	jdff dff_A_VlNZvv7n2_0(.dout(w_dff_A_lbjgfEZc1_0),.din(w_dff_A_VlNZvv7n2_0),.clk(gclk));
	jdff dff_A_lbjgfEZc1_0(.dout(w_dff_A_dAiTvqkL4_0),.din(w_dff_A_lbjgfEZc1_0),.clk(gclk));
	jdff dff_A_dAiTvqkL4_0(.dout(w_dff_A_MIXq8aL45_0),.din(w_dff_A_dAiTvqkL4_0),.clk(gclk));
	jdff dff_A_MIXq8aL45_0(.dout(w_dff_A_LxR7kWq03_0),.din(w_dff_A_MIXq8aL45_0),.clk(gclk));
	jdff dff_A_LxR7kWq03_0(.dout(w_dff_A_Lzzkozoo4_0),.din(w_dff_A_LxR7kWq03_0),.clk(gclk));
	jdff dff_A_Lzzkozoo4_0(.dout(w_dff_A_NAuNH7fS2_0),.din(w_dff_A_Lzzkozoo4_0),.clk(gclk));
	jdff dff_A_NAuNH7fS2_0(.dout(w_dff_A_OUDpUV965_0),.din(w_dff_A_NAuNH7fS2_0),.clk(gclk));
	jdff dff_A_OUDpUV965_0(.dout(w_dff_A_TZAoCCV31_0),.din(w_dff_A_OUDpUV965_0),.clk(gclk));
	jdff dff_A_TZAoCCV31_0(.dout(w_dff_A_O2FWET2g9_0),.din(w_dff_A_TZAoCCV31_0),.clk(gclk));
	jdff dff_A_O2FWET2g9_0(.dout(w_dff_A_PGVRFjAI4_0),.din(w_dff_A_O2FWET2g9_0),.clk(gclk));
	jdff dff_A_PGVRFjAI4_0(.dout(w_dff_A_B9TB6Ra76_0),.din(w_dff_A_PGVRFjAI4_0),.clk(gclk));
	jdff dff_A_B9TB6Ra76_0(.dout(w_dff_A_g59qcJCk6_0),.din(w_dff_A_B9TB6Ra76_0),.clk(gclk));
	jdff dff_A_g59qcJCk6_0(.dout(w_dff_A_dYkdEKo59_0),.din(w_dff_A_g59qcJCk6_0),.clk(gclk));
	jdff dff_A_dYkdEKo59_0(.dout(w_dff_A_DjZfWBE83_0),.din(w_dff_A_dYkdEKo59_0),.clk(gclk));
	jdff dff_A_DjZfWBE83_0(.dout(w_dff_A_urMTT55F8_0),.din(w_dff_A_DjZfWBE83_0),.clk(gclk));
	jdff dff_A_urMTT55F8_0(.dout(w_dff_A_pcLWPbgW1_0),.din(w_dff_A_urMTT55F8_0),.clk(gclk));
	jdff dff_A_pcLWPbgW1_0(.dout(w_dff_A_Z3IeNUj21_0),.din(w_dff_A_pcLWPbgW1_0),.clk(gclk));
	jdff dff_A_Z3IeNUj21_0(.dout(w_dff_A_YlWRmJC72_0),.din(w_dff_A_Z3IeNUj21_0),.clk(gclk));
	jdff dff_A_YlWRmJC72_0(.dout(w_dff_A_lM445oJ85_0),.din(w_dff_A_YlWRmJC72_0),.clk(gclk));
	jdff dff_A_lM445oJ85_0(.dout(w_dff_A_XCXeeEA88_0),.din(w_dff_A_lM445oJ85_0),.clk(gclk));
	jdff dff_A_XCXeeEA88_0(.dout(w_dff_A_NWhdtGAi3_0),.din(w_dff_A_XCXeeEA88_0),.clk(gclk));
	jdff dff_A_NWhdtGAi3_0(.dout(w_dff_A_783XIXnD7_0),.din(w_dff_A_NWhdtGAi3_0),.clk(gclk));
	jdff dff_A_783XIXnD7_0(.dout(w_dff_A_5OphFUEH4_0),.din(w_dff_A_783XIXnD7_0),.clk(gclk));
	jdff dff_A_5OphFUEH4_0(.dout(G530),.din(w_dff_A_5OphFUEH4_0),.clk(gclk));
	jdff dff_A_k7IiztBr1_1(.dout(w_dff_A_75iqSxfi4_0),.din(w_dff_A_k7IiztBr1_1),.clk(gclk));
	jdff dff_A_75iqSxfi4_0(.dout(w_dff_A_C3t7ycBr1_0),.din(w_dff_A_75iqSxfi4_0),.clk(gclk));
	jdff dff_A_C3t7ycBr1_0(.dout(w_dff_A_2KDC6p2n0_0),.din(w_dff_A_C3t7ycBr1_0),.clk(gclk));
	jdff dff_A_2KDC6p2n0_0(.dout(w_dff_A_vOW9esJO1_0),.din(w_dff_A_2KDC6p2n0_0),.clk(gclk));
	jdff dff_A_vOW9esJO1_0(.dout(w_dff_A_zbKfCUOS9_0),.din(w_dff_A_vOW9esJO1_0),.clk(gclk));
	jdff dff_A_zbKfCUOS9_0(.dout(w_dff_A_t9SxDMGz4_0),.din(w_dff_A_zbKfCUOS9_0),.clk(gclk));
	jdff dff_A_t9SxDMGz4_0(.dout(w_dff_A_bn23TTcZ1_0),.din(w_dff_A_t9SxDMGz4_0),.clk(gclk));
	jdff dff_A_bn23TTcZ1_0(.dout(w_dff_A_CBRDBPW60_0),.din(w_dff_A_bn23TTcZ1_0),.clk(gclk));
	jdff dff_A_CBRDBPW60_0(.dout(w_dff_A_opfWlgAV3_0),.din(w_dff_A_CBRDBPW60_0),.clk(gclk));
	jdff dff_A_opfWlgAV3_0(.dout(w_dff_A_osNiFCJ52_0),.din(w_dff_A_opfWlgAV3_0),.clk(gclk));
	jdff dff_A_osNiFCJ52_0(.dout(w_dff_A_iay9kg3H6_0),.din(w_dff_A_osNiFCJ52_0),.clk(gclk));
	jdff dff_A_iay9kg3H6_0(.dout(w_dff_A_8gc3hqAk5_0),.din(w_dff_A_iay9kg3H6_0),.clk(gclk));
	jdff dff_A_8gc3hqAk5_0(.dout(w_dff_A_CMotSE9g8_0),.din(w_dff_A_8gc3hqAk5_0),.clk(gclk));
	jdff dff_A_CMotSE9g8_0(.dout(w_dff_A_ZXnRSZ9T4_0),.din(w_dff_A_CMotSE9g8_0),.clk(gclk));
	jdff dff_A_ZXnRSZ9T4_0(.dout(w_dff_A_rCuwRK9n1_0),.din(w_dff_A_ZXnRSZ9T4_0),.clk(gclk));
	jdff dff_A_rCuwRK9n1_0(.dout(w_dff_A_VV41j3Yu1_0),.din(w_dff_A_rCuwRK9n1_0),.clk(gclk));
	jdff dff_A_VV41j3Yu1_0(.dout(w_dff_A_eYDKNdy51_0),.din(w_dff_A_VV41j3Yu1_0),.clk(gclk));
	jdff dff_A_eYDKNdy51_0(.dout(w_dff_A_7jW1el0h4_0),.din(w_dff_A_eYDKNdy51_0),.clk(gclk));
	jdff dff_A_7jW1el0h4_0(.dout(w_dff_A_yIE63RQf3_0),.din(w_dff_A_7jW1el0h4_0),.clk(gclk));
	jdff dff_A_yIE63RQf3_0(.dout(w_dff_A_fHoGpDUt4_0),.din(w_dff_A_yIE63RQf3_0),.clk(gclk));
	jdff dff_A_fHoGpDUt4_0(.dout(w_dff_A_xG7OdISr2_0),.din(w_dff_A_fHoGpDUt4_0),.clk(gclk));
	jdff dff_A_xG7OdISr2_0(.dout(w_dff_A_zwzzsLCO1_0),.din(w_dff_A_xG7OdISr2_0),.clk(gclk));
	jdff dff_A_zwzzsLCO1_0(.dout(w_dff_A_DLRMPsiG2_0),.din(w_dff_A_zwzzsLCO1_0),.clk(gclk));
	jdff dff_A_DLRMPsiG2_0(.dout(w_dff_A_8MD8h5AY9_0),.din(w_dff_A_DLRMPsiG2_0),.clk(gclk));
	jdff dff_A_8MD8h5AY9_0(.dout(w_dff_A_5PgaDN0w5_0),.din(w_dff_A_8MD8h5AY9_0),.clk(gclk));
	jdff dff_A_5PgaDN0w5_0(.dout(w_dff_A_8KK8V2FU1_0),.din(w_dff_A_5PgaDN0w5_0),.clk(gclk));
	jdff dff_A_8KK8V2FU1_0(.dout(G528),.din(w_dff_A_8KK8V2FU1_0),.clk(gclk));
	jdff dff_A_c5MQTItK9_1(.dout(w_dff_A_4VOsYttB2_0),.din(w_dff_A_c5MQTItK9_1),.clk(gclk));
	jdff dff_A_4VOsYttB2_0(.dout(w_dff_A_6vGJ4YZW7_0),.din(w_dff_A_4VOsYttB2_0),.clk(gclk));
	jdff dff_A_6vGJ4YZW7_0(.dout(w_dff_A_hetQ05u51_0),.din(w_dff_A_6vGJ4YZW7_0),.clk(gclk));
	jdff dff_A_hetQ05u51_0(.dout(w_dff_A_6rQxUhNr3_0),.din(w_dff_A_hetQ05u51_0),.clk(gclk));
	jdff dff_A_6rQxUhNr3_0(.dout(w_dff_A_Ug98WgI21_0),.din(w_dff_A_6rQxUhNr3_0),.clk(gclk));
	jdff dff_A_Ug98WgI21_0(.dout(w_dff_A_hRGOfzIj6_0),.din(w_dff_A_Ug98WgI21_0),.clk(gclk));
	jdff dff_A_hRGOfzIj6_0(.dout(w_dff_A_xQaZ1ijH3_0),.din(w_dff_A_hRGOfzIj6_0),.clk(gclk));
	jdff dff_A_xQaZ1ijH3_0(.dout(w_dff_A_p1B058RH4_0),.din(w_dff_A_xQaZ1ijH3_0),.clk(gclk));
	jdff dff_A_p1B058RH4_0(.dout(w_dff_A_W1Uf4Nqh9_0),.din(w_dff_A_p1B058RH4_0),.clk(gclk));
	jdff dff_A_W1Uf4Nqh9_0(.dout(w_dff_A_fC8vsPNg6_0),.din(w_dff_A_W1Uf4Nqh9_0),.clk(gclk));
	jdff dff_A_fC8vsPNg6_0(.dout(w_dff_A_AjwKw59x1_0),.din(w_dff_A_fC8vsPNg6_0),.clk(gclk));
	jdff dff_A_AjwKw59x1_0(.dout(w_dff_A_gWvU7Oov8_0),.din(w_dff_A_AjwKw59x1_0),.clk(gclk));
	jdff dff_A_gWvU7Oov8_0(.dout(w_dff_A_6bx00GY61_0),.din(w_dff_A_gWvU7Oov8_0),.clk(gclk));
	jdff dff_A_6bx00GY61_0(.dout(w_dff_A_7NoJdSJJ4_0),.din(w_dff_A_6bx00GY61_0),.clk(gclk));
	jdff dff_A_7NoJdSJJ4_0(.dout(w_dff_A_q2aJEgkd5_0),.din(w_dff_A_7NoJdSJJ4_0),.clk(gclk));
	jdff dff_A_q2aJEgkd5_0(.dout(w_dff_A_mtWUUNXM5_0),.din(w_dff_A_q2aJEgkd5_0),.clk(gclk));
	jdff dff_A_mtWUUNXM5_0(.dout(w_dff_A_VZSXlrIl4_0),.din(w_dff_A_mtWUUNXM5_0),.clk(gclk));
	jdff dff_A_VZSXlrIl4_0(.dout(w_dff_A_Y3J4dLad2_0),.din(w_dff_A_VZSXlrIl4_0),.clk(gclk));
	jdff dff_A_Y3J4dLad2_0(.dout(w_dff_A_VHl2Qsm91_0),.din(w_dff_A_Y3J4dLad2_0),.clk(gclk));
	jdff dff_A_VHl2Qsm91_0(.dout(w_dff_A_GjB697Ok2_0),.din(w_dff_A_VHl2Qsm91_0),.clk(gclk));
	jdff dff_A_GjB697Ok2_0(.dout(w_dff_A_O2OfC5Ja7_0),.din(w_dff_A_GjB697Ok2_0),.clk(gclk));
	jdff dff_A_O2OfC5Ja7_0(.dout(w_dff_A_IYRYfPIz5_0),.din(w_dff_A_O2OfC5Ja7_0),.clk(gclk));
	jdff dff_A_IYRYfPIz5_0(.dout(w_dff_A_EuZuotvZ8_0),.din(w_dff_A_IYRYfPIz5_0),.clk(gclk));
	jdff dff_A_EuZuotvZ8_0(.dout(w_dff_A_DvThwb6U7_0),.din(w_dff_A_EuZuotvZ8_0),.clk(gclk));
	jdff dff_A_DvThwb6U7_0(.dout(w_dff_A_oLccsbfM2_0),.din(w_dff_A_DvThwb6U7_0),.clk(gclk));
	jdff dff_A_oLccsbfM2_0(.dout(w_dff_A_QfuqvVLH2_0),.din(w_dff_A_oLccsbfM2_0),.clk(gclk));
	jdff dff_A_QfuqvVLH2_0(.dout(G526),.din(w_dff_A_QfuqvVLH2_0),.clk(gclk));
	jdff dff_A_xu1agTiB2_1(.dout(w_dff_A_lrqAy2L44_0),.din(w_dff_A_xu1agTiB2_1),.clk(gclk));
	jdff dff_A_lrqAy2L44_0(.dout(w_dff_A_2LhSkjYI2_0),.din(w_dff_A_lrqAy2L44_0),.clk(gclk));
	jdff dff_A_2LhSkjYI2_0(.dout(w_dff_A_KwbHDxT89_0),.din(w_dff_A_2LhSkjYI2_0),.clk(gclk));
	jdff dff_A_KwbHDxT89_0(.dout(w_dff_A_pKmkvdXK3_0),.din(w_dff_A_KwbHDxT89_0),.clk(gclk));
	jdff dff_A_pKmkvdXK3_0(.dout(w_dff_A_wriAhwEy3_0),.din(w_dff_A_pKmkvdXK3_0),.clk(gclk));
	jdff dff_A_wriAhwEy3_0(.dout(w_dff_A_zjFNdKXD4_0),.din(w_dff_A_wriAhwEy3_0),.clk(gclk));
	jdff dff_A_zjFNdKXD4_0(.dout(w_dff_A_ABPQTlRW3_0),.din(w_dff_A_zjFNdKXD4_0),.clk(gclk));
	jdff dff_A_ABPQTlRW3_0(.dout(w_dff_A_oKvp4cll4_0),.din(w_dff_A_ABPQTlRW3_0),.clk(gclk));
	jdff dff_A_oKvp4cll4_0(.dout(w_dff_A_7t0PUetP6_0),.din(w_dff_A_oKvp4cll4_0),.clk(gclk));
	jdff dff_A_7t0PUetP6_0(.dout(w_dff_A_Xrrzqlz08_0),.din(w_dff_A_7t0PUetP6_0),.clk(gclk));
	jdff dff_A_Xrrzqlz08_0(.dout(w_dff_A_B2B8eAdk1_0),.din(w_dff_A_Xrrzqlz08_0),.clk(gclk));
	jdff dff_A_B2B8eAdk1_0(.dout(w_dff_A_11t3bD4x2_0),.din(w_dff_A_B2B8eAdk1_0),.clk(gclk));
	jdff dff_A_11t3bD4x2_0(.dout(w_dff_A_CErQ3RXZ8_0),.din(w_dff_A_11t3bD4x2_0),.clk(gclk));
	jdff dff_A_CErQ3RXZ8_0(.dout(w_dff_A_TnYSVxcW8_0),.din(w_dff_A_CErQ3RXZ8_0),.clk(gclk));
	jdff dff_A_TnYSVxcW8_0(.dout(w_dff_A_ONiOXrDK7_0),.din(w_dff_A_TnYSVxcW8_0),.clk(gclk));
	jdff dff_A_ONiOXrDK7_0(.dout(w_dff_A_jGqhMNPh6_0),.din(w_dff_A_ONiOXrDK7_0),.clk(gclk));
	jdff dff_A_jGqhMNPh6_0(.dout(w_dff_A_o6qYlUTn1_0),.din(w_dff_A_jGqhMNPh6_0),.clk(gclk));
	jdff dff_A_o6qYlUTn1_0(.dout(w_dff_A_t00olKhs4_0),.din(w_dff_A_o6qYlUTn1_0),.clk(gclk));
	jdff dff_A_t00olKhs4_0(.dout(w_dff_A_FF481w1r1_0),.din(w_dff_A_t00olKhs4_0),.clk(gclk));
	jdff dff_A_FF481w1r1_0(.dout(w_dff_A_tpxobTtJ5_0),.din(w_dff_A_FF481w1r1_0),.clk(gclk));
	jdff dff_A_tpxobTtJ5_0(.dout(w_dff_A_s0QMpRhn5_0),.din(w_dff_A_tpxobTtJ5_0),.clk(gclk));
	jdff dff_A_s0QMpRhn5_0(.dout(w_dff_A_TrAEPDb11_0),.din(w_dff_A_s0QMpRhn5_0),.clk(gclk));
	jdff dff_A_TrAEPDb11_0(.dout(w_dff_A_rMDW1a3L4_0),.din(w_dff_A_TrAEPDb11_0),.clk(gclk));
	jdff dff_A_rMDW1a3L4_0(.dout(w_dff_A_osaNfKJg7_0),.din(w_dff_A_rMDW1a3L4_0),.clk(gclk));
	jdff dff_A_osaNfKJg7_0(.dout(w_dff_A_ufg8Bxsy6_0),.din(w_dff_A_osaNfKJg7_0),.clk(gclk));
	jdff dff_A_ufg8Bxsy6_0(.dout(w_dff_A_kvlVS9Fw7_0),.din(w_dff_A_ufg8Bxsy6_0),.clk(gclk));
	jdff dff_A_kvlVS9Fw7_0(.dout(G524),.din(w_dff_A_kvlVS9Fw7_0),.clk(gclk));
	jdff dff_A_7bvST8917_1(.dout(w_dff_A_8BvXaxfK7_0),.din(w_dff_A_7bvST8917_1),.clk(gclk));
	jdff dff_A_8BvXaxfK7_0(.dout(w_dff_A_TWtU7c1f1_0),.din(w_dff_A_8BvXaxfK7_0),.clk(gclk));
	jdff dff_A_TWtU7c1f1_0(.dout(w_dff_A_pQyHmwTQ6_0),.din(w_dff_A_TWtU7c1f1_0),.clk(gclk));
	jdff dff_A_pQyHmwTQ6_0(.dout(w_dff_A_I9iFABSc3_0),.din(w_dff_A_pQyHmwTQ6_0),.clk(gclk));
	jdff dff_A_I9iFABSc3_0(.dout(w_dff_A_vWpyJEp82_0),.din(w_dff_A_I9iFABSc3_0),.clk(gclk));
	jdff dff_A_vWpyJEp82_0(.dout(w_dff_A_439c9kkD0_0),.din(w_dff_A_vWpyJEp82_0),.clk(gclk));
	jdff dff_A_439c9kkD0_0(.dout(w_dff_A_EsHXbldW7_0),.din(w_dff_A_439c9kkD0_0),.clk(gclk));
	jdff dff_A_EsHXbldW7_0(.dout(w_dff_A_oYriIHjx0_0),.din(w_dff_A_EsHXbldW7_0),.clk(gclk));
	jdff dff_A_oYriIHjx0_0(.dout(w_dff_A_b07LerSg3_0),.din(w_dff_A_oYriIHjx0_0),.clk(gclk));
	jdff dff_A_b07LerSg3_0(.dout(w_dff_A_pyQfw6Du5_0),.din(w_dff_A_b07LerSg3_0),.clk(gclk));
	jdff dff_A_pyQfw6Du5_0(.dout(w_dff_A_QNnptJA61_0),.din(w_dff_A_pyQfw6Du5_0),.clk(gclk));
	jdff dff_A_QNnptJA61_0(.dout(w_dff_A_UYmtoCrC7_0),.din(w_dff_A_QNnptJA61_0),.clk(gclk));
	jdff dff_A_UYmtoCrC7_0(.dout(w_dff_A_rbA6QmCE6_0),.din(w_dff_A_UYmtoCrC7_0),.clk(gclk));
	jdff dff_A_rbA6QmCE6_0(.dout(w_dff_A_Xz54Jsmr9_0),.din(w_dff_A_rbA6QmCE6_0),.clk(gclk));
	jdff dff_A_Xz54Jsmr9_0(.dout(w_dff_A_SHKX5rW55_0),.din(w_dff_A_Xz54Jsmr9_0),.clk(gclk));
	jdff dff_A_SHKX5rW55_0(.dout(w_dff_A_WiqDAh0n7_0),.din(w_dff_A_SHKX5rW55_0),.clk(gclk));
	jdff dff_A_WiqDAh0n7_0(.dout(w_dff_A_EILdXOk58_0),.din(w_dff_A_WiqDAh0n7_0),.clk(gclk));
	jdff dff_A_EILdXOk58_0(.dout(w_dff_A_gLPZjr6N7_0),.din(w_dff_A_EILdXOk58_0),.clk(gclk));
	jdff dff_A_gLPZjr6N7_0(.dout(w_dff_A_DRuwiEfA0_0),.din(w_dff_A_gLPZjr6N7_0),.clk(gclk));
	jdff dff_A_DRuwiEfA0_0(.dout(w_dff_A_cbqdluqx1_0),.din(w_dff_A_DRuwiEfA0_0),.clk(gclk));
	jdff dff_A_cbqdluqx1_0(.dout(w_dff_A_bnllwroc5_0),.din(w_dff_A_cbqdluqx1_0),.clk(gclk));
	jdff dff_A_bnllwroc5_0(.dout(w_dff_A_MofP6H440_0),.din(w_dff_A_bnllwroc5_0),.clk(gclk));
	jdff dff_A_MofP6H440_0(.dout(w_dff_A_4iIdPi8J8_0),.din(w_dff_A_MofP6H440_0),.clk(gclk));
	jdff dff_A_4iIdPi8J8_0(.dout(w_dff_A_L0FaI5wy3_0),.din(w_dff_A_4iIdPi8J8_0),.clk(gclk));
	jdff dff_A_L0FaI5wy3_0(.dout(w_dff_A_I1Y7i4EX3_0),.din(w_dff_A_L0FaI5wy3_0),.clk(gclk));
	jdff dff_A_I1Y7i4EX3_0(.dout(G279),.din(w_dff_A_I1Y7i4EX3_0),.clk(gclk));
	jdff dff_A_6UWDOWSA1_1(.dout(w_dff_A_vn8vYwO54_0),.din(w_dff_A_6UWDOWSA1_1),.clk(gclk));
	jdff dff_A_vn8vYwO54_0(.dout(w_dff_A_5Tgf4Bdv8_0),.din(w_dff_A_vn8vYwO54_0),.clk(gclk));
	jdff dff_A_5Tgf4Bdv8_0(.dout(w_dff_A_jGFbwH2A8_0),.din(w_dff_A_5Tgf4Bdv8_0),.clk(gclk));
	jdff dff_A_jGFbwH2A8_0(.dout(w_dff_A_FWEA7P7f1_0),.din(w_dff_A_jGFbwH2A8_0),.clk(gclk));
	jdff dff_A_FWEA7P7f1_0(.dout(w_dff_A_VTdHVwMc6_0),.din(w_dff_A_FWEA7P7f1_0),.clk(gclk));
	jdff dff_A_VTdHVwMc6_0(.dout(w_dff_A_QrAC74wH8_0),.din(w_dff_A_VTdHVwMc6_0),.clk(gclk));
	jdff dff_A_QrAC74wH8_0(.dout(w_dff_A_vpRfzOOT8_0),.din(w_dff_A_QrAC74wH8_0),.clk(gclk));
	jdff dff_A_vpRfzOOT8_0(.dout(w_dff_A_Lno3wbIi4_0),.din(w_dff_A_vpRfzOOT8_0),.clk(gclk));
	jdff dff_A_Lno3wbIi4_0(.dout(w_dff_A_yj41Odb64_0),.din(w_dff_A_Lno3wbIi4_0),.clk(gclk));
	jdff dff_A_yj41Odb64_0(.dout(w_dff_A_ChCYih8I6_0),.din(w_dff_A_yj41Odb64_0),.clk(gclk));
	jdff dff_A_ChCYih8I6_0(.dout(w_dff_A_D1cZPIEM3_0),.din(w_dff_A_ChCYih8I6_0),.clk(gclk));
	jdff dff_A_D1cZPIEM3_0(.dout(w_dff_A_D9WFSkqf7_0),.din(w_dff_A_D1cZPIEM3_0),.clk(gclk));
	jdff dff_A_D9WFSkqf7_0(.dout(w_dff_A_lN9HBeEW6_0),.din(w_dff_A_D9WFSkqf7_0),.clk(gclk));
	jdff dff_A_lN9HBeEW6_0(.dout(w_dff_A_uOqTjRE81_0),.din(w_dff_A_lN9HBeEW6_0),.clk(gclk));
	jdff dff_A_uOqTjRE81_0(.dout(w_dff_A_wW6giJO10_0),.din(w_dff_A_uOqTjRE81_0),.clk(gclk));
	jdff dff_A_wW6giJO10_0(.dout(w_dff_A_9hd2PDPw2_0),.din(w_dff_A_wW6giJO10_0),.clk(gclk));
	jdff dff_A_9hd2PDPw2_0(.dout(w_dff_A_Yk2Zh7iN3_0),.din(w_dff_A_9hd2PDPw2_0),.clk(gclk));
	jdff dff_A_Yk2Zh7iN3_0(.dout(w_dff_A_m2Ezucv33_0),.din(w_dff_A_Yk2Zh7iN3_0),.clk(gclk));
	jdff dff_A_m2Ezucv33_0(.dout(w_dff_A_KBDbDuUW1_0),.din(w_dff_A_m2Ezucv33_0),.clk(gclk));
	jdff dff_A_KBDbDuUW1_0(.dout(w_dff_A_o8uZ0s8r0_0),.din(w_dff_A_KBDbDuUW1_0),.clk(gclk));
	jdff dff_A_o8uZ0s8r0_0(.dout(w_dff_A_gxUG7u9A0_0),.din(w_dff_A_o8uZ0s8r0_0),.clk(gclk));
	jdff dff_A_gxUG7u9A0_0(.dout(w_dff_A_4irXiDOc8_0),.din(w_dff_A_gxUG7u9A0_0),.clk(gclk));
	jdff dff_A_4irXiDOc8_0(.dout(w_dff_A_vgs9vWSN5_0),.din(w_dff_A_4irXiDOc8_0),.clk(gclk));
	jdff dff_A_vgs9vWSN5_0(.dout(w_dff_A_9QLzCYgU1_0),.din(w_dff_A_vgs9vWSN5_0),.clk(gclk));
	jdff dff_A_9QLzCYgU1_0(.dout(w_dff_A_cz8UdtXi3_0),.din(w_dff_A_9QLzCYgU1_0),.clk(gclk));
	jdff dff_A_cz8UdtXi3_0(.dout(w_dff_A_0pbaQvQh7_0),.din(w_dff_A_cz8UdtXi3_0),.clk(gclk));
	jdff dff_A_0pbaQvQh7_0(.dout(G436),.din(w_dff_A_0pbaQvQh7_0),.clk(gclk));
	jdff dff_A_l4pLZDe96_1(.dout(w_dff_A_dBuom1lU3_0),.din(w_dff_A_l4pLZDe96_1),.clk(gclk));
	jdff dff_A_dBuom1lU3_0(.dout(w_dff_A_LP2Tqdkx4_0),.din(w_dff_A_dBuom1lU3_0),.clk(gclk));
	jdff dff_A_LP2Tqdkx4_0(.dout(w_dff_A_oLc7MfjE4_0),.din(w_dff_A_LP2Tqdkx4_0),.clk(gclk));
	jdff dff_A_oLc7MfjE4_0(.dout(w_dff_A_aJAFwLE92_0),.din(w_dff_A_oLc7MfjE4_0),.clk(gclk));
	jdff dff_A_aJAFwLE92_0(.dout(w_dff_A_cjd4Il9M2_0),.din(w_dff_A_aJAFwLE92_0),.clk(gclk));
	jdff dff_A_cjd4Il9M2_0(.dout(w_dff_A_bglDhIb82_0),.din(w_dff_A_cjd4Il9M2_0),.clk(gclk));
	jdff dff_A_bglDhIb82_0(.dout(w_dff_A_Ik0JOtjQ5_0),.din(w_dff_A_bglDhIb82_0),.clk(gclk));
	jdff dff_A_Ik0JOtjQ5_0(.dout(w_dff_A_JHpvRwiM7_0),.din(w_dff_A_Ik0JOtjQ5_0),.clk(gclk));
	jdff dff_A_JHpvRwiM7_0(.dout(w_dff_A_Pdd57MkJ3_0),.din(w_dff_A_JHpvRwiM7_0),.clk(gclk));
	jdff dff_A_Pdd57MkJ3_0(.dout(w_dff_A_zZndK0pA8_0),.din(w_dff_A_Pdd57MkJ3_0),.clk(gclk));
	jdff dff_A_zZndK0pA8_0(.dout(w_dff_A_BkKRg6jA4_0),.din(w_dff_A_zZndK0pA8_0),.clk(gclk));
	jdff dff_A_BkKRg6jA4_0(.dout(w_dff_A_ZCeitO3o9_0),.din(w_dff_A_BkKRg6jA4_0),.clk(gclk));
	jdff dff_A_ZCeitO3o9_0(.dout(w_dff_A_cutHzJP41_0),.din(w_dff_A_ZCeitO3o9_0),.clk(gclk));
	jdff dff_A_cutHzJP41_0(.dout(w_dff_A_WxeP7fne2_0),.din(w_dff_A_cutHzJP41_0),.clk(gclk));
	jdff dff_A_WxeP7fne2_0(.dout(w_dff_A_USYmMaZP7_0),.din(w_dff_A_WxeP7fne2_0),.clk(gclk));
	jdff dff_A_USYmMaZP7_0(.dout(w_dff_A_GSzvcO6H5_0),.din(w_dff_A_USYmMaZP7_0),.clk(gclk));
	jdff dff_A_GSzvcO6H5_0(.dout(w_dff_A_XAashtOp0_0),.din(w_dff_A_GSzvcO6H5_0),.clk(gclk));
	jdff dff_A_XAashtOp0_0(.dout(w_dff_A_ulDPMT8X6_0),.din(w_dff_A_XAashtOp0_0),.clk(gclk));
	jdff dff_A_ulDPMT8X6_0(.dout(w_dff_A_eho0bCVh8_0),.din(w_dff_A_ulDPMT8X6_0),.clk(gclk));
	jdff dff_A_eho0bCVh8_0(.dout(w_dff_A_Ey6KZK048_0),.din(w_dff_A_eho0bCVh8_0),.clk(gclk));
	jdff dff_A_Ey6KZK048_0(.dout(w_dff_A_MehFAZ5B4_0),.din(w_dff_A_Ey6KZK048_0),.clk(gclk));
	jdff dff_A_MehFAZ5B4_0(.dout(w_dff_A_NUne2LM84_0),.din(w_dff_A_MehFAZ5B4_0),.clk(gclk));
	jdff dff_A_NUne2LM84_0(.dout(w_dff_A_HWRUraAz0_0),.din(w_dff_A_NUne2LM84_0),.clk(gclk));
	jdff dff_A_HWRUraAz0_0(.dout(w_dff_A_4RCNy5d40_0),.din(w_dff_A_HWRUraAz0_0),.clk(gclk));
	jdff dff_A_4RCNy5d40_0(.dout(w_dff_A_Iobuwp0F1_0),.din(w_dff_A_4RCNy5d40_0),.clk(gclk));
	jdff dff_A_Iobuwp0F1_0(.dout(w_dff_A_WiUtrs525_0),.din(w_dff_A_Iobuwp0F1_0),.clk(gclk));
	jdff dff_A_WiUtrs525_0(.dout(G478),.din(w_dff_A_WiUtrs525_0),.clk(gclk));
	jdff dff_A_eaYLuokZ0_1(.dout(w_dff_A_HzgHeKjZ5_0),.din(w_dff_A_eaYLuokZ0_1),.clk(gclk));
	jdff dff_A_HzgHeKjZ5_0(.dout(w_dff_A_7HfhwGA17_0),.din(w_dff_A_HzgHeKjZ5_0),.clk(gclk));
	jdff dff_A_7HfhwGA17_0(.dout(w_dff_A_lZsVeOrI8_0),.din(w_dff_A_7HfhwGA17_0),.clk(gclk));
	jdff dff_A_lZsVeOrI8_0(.dout(w_dff_A_O4TWv1f76_0),.din(w_dff_A_lZsVeOrI8_0),.clk(gclk));
	jdff dff_A_O4TWv1f76_0(.dout(w_dff_A_80PdiP009_0),.din(w_dff_A_O4TWv1f76_0),.clk(gclk));
	jdff dff_A_80PdiP009_0(.dout(w_dff_A_qnNiLbsw4_0),.din(w_dff_A_80PdiP009_0),.clk(gclk));
	jdff dff_A_qnNiLbsw4_0(.dout(w_dff_A_1GMG43Jq0_0),.din(w_dff_A_qnNiLbsw4_0),.clk(gclk));
	jdff dff_A_1GMG43Jq0_0(.dout(w_dff_A_rRlWRf4x4_0),.din(w_dff_A_1GMG43Jq0_0),.clk(gclk));
	jdff dff_A_rRlWRf4x4_0(.dout(w_dff_A_ZE7WKBQ35_0),.din(w_dff_A_rRlWRf4x4_0),.clk(gclk));
	jdff dff_A_ZE7WKBQ35_0(.dout(w_dff_A_nD04OMSb6_0),.din(w_dff_A_ZE7WKBQ35_0),.clk(gclk));
	jdff dff_A_nD04OMSb6_0(.dout(w_dff_A_bQU9CVZf9_0),.din(w_dff_A_nD04OMSb6_0),.clk(gclk));
	jdff dff_A_bQU9CVZf9_0(.dout(w_dff_A_G9QN4jvF3_0),.din(w_dff_A_bQU9CVZf9_0),.clk(gclk));
	jdff dff_A_G9QN4jvF3_0(.dout(w_dff_A_PnvknPpP6_0),.din(w_dff_A_G9QN4jvF3_0),.clk(gclk));
	jdff dff_A_PnvknPpP6_0(.dout(w_dff_A_UlMEasx26_0),.din(w_dff_A_PnvknPpP6_0),.clk(gclk));
	jdff dff_A_UlMEasx26_0(.dout(w_dff_A_U6ITe5oR7_0),.din(w_dff_A_UlMEasx26_0),.clk(gclk));
	jdff dff_A_U6ITe5oR7_0(.dout(w_dff_A_1g68nLPq2_0),.din(w_dff_A_U6ITe5oR7_0),.clk(gclk));
	jdff dff_A_1g68nLPq2_0(.dout(w_dff_A_WjyvEmKn7_0),.din(w_dff_A_1g68nLPq2_0),.clk(gclk));
	jdff dff_A_WjyvEmKn7_0(.dout(w_dff_A_TNuN9byB5_0),.din(w_dff_A_WjyvEmKn7_0),.clk(gclk));
	jdff dff_A_TNuN9byB5_0(.dout(w_dff_A_81v4I8Ew4_0),.din(w_dff_A_TNuN9byB5_0),.clk(gclk));
	jdff dff_A_81v4I8Ew4_0(.dout(w_dff_A_scxawDpb4_0),.din(w_dff_A_81v4I8Ew4_0),.clk(gclk));
	jdff dff_A_scxawDpb4_0(.dout(w_dff_A_2sMe1RwB0_0),.din(w_dff_A_scxawDpb4_0),.clk(gclk));
	jdff dff_A_2sMe1RwB0_0(.dout(w_dff_A_uTljhGQn9_0),.din(w_dff_A_2sMe1RwB0_0),.clk(gclk));
	jdff dff_A_uTljhGQn9_0(.dout(w_dff_A_tPSQsWNp6_0),.din(w_dff_A_uTljhGQn9_0),.clk(gclk));
	jdff dff_A_tPSQsWNp6_0(.dout(w_dff_A_zimTBsAz4_0),.din(w_dff_A_tPSQsWNp6_0),.clk(gclk));
	jdff dff_A_zimTBsAz4_0(.dout(w_dff_A_dhJQa4vr0_0),.din(w_dff_A_zimTBsAz4_0),.clk(gclk));
	jdff dff_A_dhJQa4vr0_0(.dout(w_dff_A_AY2UsahH4_0),.din(w_dff_A_dhJQa4vr0_0),.clk(gclk));
	jdff dff_A_AY2UsahH4_0(.dout(G522),.din(w_dff_A_AY2UsahH4_0),.clk(gclk));
	jdff dff_A_c5Bpdw724_2(.dout(w_dff_A_OGQmfdLx7_0),.din(w_dff_A_c5Bpdw724_2),.clk(gclk));
	jdff dff_A_OGQmfdLx7_0(.dout(w_dff_A_jDqFtL9x1_0),.din(w_dff_A_OGQmfdLx7_0),.clk(gclk));
	jdff dff_A_jDqFtL9x1_0(.dout(w_dff_A_3VuG7dLC2_0),.din(w_dff_A_jDqFtL9x1_0),.clk(gclk));
	jdff dff_A_3VuG7dLC2_0(.dout(w_dff_A_foG3f27D3_0),.din(w_dff_A_3VuG7dLC2_0),.clk(gclk));
	jdff dff_A_foG3f27D3_0(.dout(w_dff_A_VdeLpShU8_0),.din(w_dff_A_foG3f27D3_0),.clk(gclk));
	jdff dff_A_VdeLpShU8_0(.dout(w_dff_A_Ipx5d0C58_0),.din(w_dff_A_VdeLpShU8_0),.clk(gclk));
	jdff dff_A_Ipx5d0C58_0(.dout(w_dff_A_GX23GRlu3_0),.din(w_dff_A_Ipx5d0C58_0),.clk(gclk));
	jdff dff_A_GX23GRlu3_0(.dout(w_dff_A_UG2DYt5s1_0),.din(w_dff_A_GX23GRlu3_0),.clk(gclk));
	jdff dff_A_UG2DYt5s1_0(.dout(w_dff_A_P1SrnOu53_0),.din(w_dff_A_UG2DYt5s1_0),.clk(gclk));
	jdff dff_A_P1SrnOu53_0(.dout(w_dff_A_m554hjvt9_0),.din(w_dff_A_P1SrnOu53_0),.clk(gclk));
	jdff dff_A_m554hjvt9_0(.dout(w_dff_A_oF1LMhTv4_0),.din(w_dff_A_m554hjvt9_0),.clk(gclk));
	jdff dff_A_oF1LMhTv4_0(.dout(w_dff_A_W24l9afA7_0),.din(w_dff_A_oF1LMhTv4_0),.clk(gclk));
	jdff dff_A_W24l9afA7_0(.dout(w_dff_A_G0FVvffF3_0),.din(w_dff_A_W24l9afA7_0),.clk(gclk));
	jdff dff_A_G0FVvffF3_0(.dout(w_dff_A_vX7o7EMY6_0),.din(w_dff_A_G0FVvffF3_0),.clk(gclk));
	jdff dff_A_vX7o7EMY6_0(.dout(w_dff_A_uMYkhgM23_0),.din(w_dff_A_vX7o7EMY6_0),.clk(gclk));
	jdff dff_A_uMYkhgM23_0(.dout(w_dff_A_mdksk9u94_0),.din(w_dff_A_uMYkhgM23_0),.clk(gclk));
	jdff dff_A_mdksk9u94_0(.dout(w_dff_A_U6raieEU1_0),.din(w_dff_A_mdksk9u94_0),.clk(gclk));
	jdff dff_A_U6raieEU1_0(.dout(w_dff_A_MXbUDuQv9_0),.din(w_dff_A_U6raieEU1_0),.clk(gclk));
	jdff dff_A_MXbUDuQv9_0(.dout(w_dff_A_uAbWB8pv4_0),.din(w_dff_A_MXbUDuQv9_0),.clk(gclk));
	jdff dff_A_uAbWB8pv4_0(.dout(w_dff_A_oszbms297_0),.din(w_dff_A_uAbWB8pv4_0),.clk(gclk));
	jdff dff_A_oszbms297_0(.dout(w_dff_A_2CkbKNXS3_0),.din(w_dff_A_oszbms297_0),.clk(gclk));
	jdff dff_A_2CkbKNXS3_0(.dout(w_dff_A_Lhg4OACg7_0),.din(w_dff_A_2CkbKNXS3_0),.clk(gclk));
	jdff dff_A_Lhg4OACg7_0(.dout(w_dff_A_Dep6pJPm6_0),.din(w_dff_A_Lhg4OACg7_0),.clk(gclk));
	jdff dff_A_Dep6pJPm6_0(.dout(w_dff_A_vgStCyCG2_0),.din(w_dff_A_Dep6pJPm6_0),.clk(gclk));
	jdff dff_A_vgStCyCG2_0(.dout(w_dff_A_9XGX6FUe8_0),.din(w_dff_A_vgStCyCG2_0),.clk(gclk));
	jdff dff_A_9XGX6FUe8_0(.dout(G402),.din(w_dff_A_9XGX6FUe8_0),.clk(gclk));
	jdff dff_A_JtkNZIA12_1(.dout(w_dff_A_4WY3wfai9_0),.din(w_dff_A_JtkNZIA12_1),.clk(gclk));
	jdff dff_A_4WY3wfai9_0(.dout(w_dff_A_GDFVRGeD1_0),.din(w_dff_A_4WY3wfai9_0),.clk(gclk));
	jdff dff_A_GDFVRGeD1_0(.dout(w_dff_A_6OXD3BVa8_0),.din(w_dff_A_GDFVRGeD1_0),.clk(gclk));
	jdff dff_A_6OXD3BVa8_0(.dout(w_dff_A_RZv2ZpI35_0),.din(w_dff_A_6OXD3BVa8_0),.clk(gclk));
	jdff dff_A_RZv2ZpI35_0(.dout(w_dff_A_q0UzIxli6_0),.din(w_dff_A_RZv2ZpI35_0),.clk(gclk));
	jdff dff_A_q0UzIxli6_0(.dout(w_dff_A_E8rjbMvU3_0),.din(w_dff_A_q0UzIxli6_0),.clk(gclk));
	jdff dff_A_E8rjbMvU3_0(.dout(w_dff_A_8xyq2cwx8_0),.din(w_dff_A_E8rjbMvU3_0),.clk(gclk));
	jdff dff_A_8xyq2cwx8_0(.dout(w_dff_A_pP9XxWYx0_0),.din(w_dff_A_8xyq2cwx8_0),.clk(gclk));
	jdff dff_A_pP9XxWYx0_0(.dout(w_dff_A_qSot8xif5_0),.din(w_dff_A_pP9XxWYx0_0),.clk(gclk));
	jdff dff_A_qSot8xif5_0(.dout(w_dff_A_0RlWnT658_0),.din(w_dff_A_qSot8xif5_0),.clk(gclk));
	jdff dff_A_0RlWnT658_0(.dout(w_dff_A_LY4MRAap9_0),.din(w_dff_A_0RlWnT658_0),.clk(gclk));
	jdff dff_A_LY4MRAap9_0(.dout(w_dff_A_gWs4m90F6_0),.din(w_dff_A_LY4MRAap9_0),.clk(gclk));
	jdff dff_A_gWs4m90F6_0(.dout(w_dff_A_7CZWdSKy8_0),.din(w_dff_A_gWs4m90F6_0),.clk(gclk));
	jdff dff_A_7CZWdSKy8_0(.dout(w_dff_A_2KkwN80j9_0),.din(w_dff_A_7CZWdSKy8_0),.clk(gclk));
	jdff dff_A_2KkwN80j9_0(.dout(w_dff_A_2nBJX9c12_0),.din(w_dff_A_2KkwN80j9_0),.clk(gclk));
	jdff dff_A_2nBJX9c12_0(.dout(w_dff_A_yU2NPQD99_0),.din(w_dff_A_2nBJX9c12_0),.clk(gclk));
	jdff dff_A_yU2NPQD99_0(.dout(w_dff_A_MIdyw7zw1_0),.din(w_dff_A_yU2NPQD99_0),.clk(gclk));
	jdff dff_A_MIdyw7zw1_0(.dout(w_dff_A_MTaFvIEq7_0),.din(w_dff_A_MIdyw7zw1_0),.clk(gclk));
	jdff dff_A_MTaFvIEq7_0(.dout(w_dff_A_4V4E08a95_0),.din(w_dff_A_MTaFvIEq7_0),.clk(gclk));
	jdff dff_A_4V4E08a95_0(.dout(w_dff_A_779SVaTk8_0),.din(w_dff_A_4V4E08a95_0),.clk(gclk));
	jdff dff_A_779SVaTk8_0(.dout(w_dff_A_lQAeoPEx4_0),.din(w_dff_A_779SVaTk8_0),.clk(gclk));
	jdff dff_A_lQAeoPEx4_0(.dout(w_dff_A_tApUQjOd3_0),.din(w_dff_A_lQAeoPEx4_0),.clk(gclk));
	jdff dff_A_tApUQjOd3_0(.dout(w_dff_A_F0ZFqzmZ1_0),.din(w_dff_A_tApUQjOd3_0),.clk(gclk));
	jdff dff_A_F0ZFqzmZ1_0(.dout(G404),.din(w_dff_A_F0ZFqzmZ1_0),.clk(gclk));
	jdff dff_A_wBQV3noA7_1(.dout(w_dff_A_vI62fLtD9_0),.din(w_dff_A_wBQV3noA7_1),.clk(gclk));
	jdff dff_A_vI62fLtD9_0(.dout(w_dff_A_fUbbepUN5_0),.din(w_dff_A_vI62fLtD9_0),.clk(gclk));
	jdff dff_A_fUbbepUN5_0(.dout(w_dff_A_RX7e92Sr5_0),.din(w_dff_A_fUbbepUN5_0),.clk(gclk));
	jdff dff_A_RX7e92Sr5_0(.dout(w_dff_A_FBYe2Uek3_0),.din(w_dff_A_RX7e92Sr5_0),.clk(gclk));
	jdff dff_A_FBYe2Uek3_0(.dout(w_dff_A_x76m5M6j0_0),.din(w_dff_A_FBYe2Uek3_0),.clk(gclk));
	jdff dff_A_x76m5M6j0_0(.dout(w_dff_A_IhIgCuvW5_0),.din(w_dff_A_x76m5M6j0_0),.clk(gclk));
	jdff dff_A_IhIgCuvW5_0(.dout(w_dff_A_ECE7xGUS0_0),.din(w_dff_A_IhIgCuvW5_0),.clk(gclk));
	jdff dff_A_ECE7xGUS0_0(.dout(w_dff_A_MU1A8api7_0),.din(w_dff_A_ECE7xGUS0_0),.clk(gclk));
	jdff dff_A_MU1A8api7_0(.dout(w_dff_A_MCRGttNN8_0),.din(w_dff_A_MU1A8api7_0),.clk(gclk));
	jdff dff_A_MCRGttNN8_0(.dout(w_dff_A_ePc4h8MT0_0),.din(w_dff_A_MCRGttNN8_0),.clk(gclk));
	jdff dff_A_ePc4h8MT0_0(.dout(w_dff_A_UupNxGsL8_0),.din(w_dff_A_ePc4h8MT0_0),.clk(gclk));
	jdff dff_A_UupNxGsL8_0(.dout(w_dff_A_nOJxS9Jg1_0),.din(w_dff_A_UupNxGsL8_0),.clk(gclk));
	jdff dff_A_nOJxS9Jg1_0(.dout(w_dff_A_EHkxXtRZ9_0),.din(w_dff_A_nOJxS9Jg1_0),.clk(gclk));
	jdff dff_A_EHkxXtRZ9_0(.dout(w_dff_A_xJw1jpc66_0),.din(w_dff_A_EHkxXtRZ9_0),.clk(gclk));
	jdff dff_A_xJw1jpc66_0(.dout(w_dff_A_QNczrOVf9_0),.din(w_dff_A_xJw1jpc66_0),.clk(gclk));
	jdff dff_A_QNczrOVf9_0(.dout(w_dff_A_wFZ3ijgK6_0),.din(w_dff_A_QNczrOVf9_0),.clk(gclk));
	jdff dff_A_wFZ3ijgK6_0(.dout(w_dff_A_Czqn3NUB0_0),.din(w_dff_A_wFZ3ijgK6_0),.clk(gclk));
	jdff dff_A_Czqn3NUB0_0(.dout(w_dff_A_3eu3AR8j4_0),.din(w_dff_A_Czqn3NUB0_0),.clk(gclk));
	jdff dff_A_3eu3AR8j4_0(.dout(w_dff_A_UewIoyYU2_0),.din(w_dff_A_3eu3AR8j4_0),.clk(gclk));
	jdff dff_A_UewIoyYU2_0(.dout(w_dff_A_3xUuhlZG1_0),.din(w_dff_A_UewIoyYU2_0),.clk(gclk));
	jdff dff_A_3xUuhlZG1_0(.dout(w_dff_A_gZDCfb638_0),.din(w_dff_A_3xUuhlZG1_0),.clk(gclk));
	jdff dff_A_gZDCfb638_0(.dout(w_dff_A_e21azBOc4_0),.din(w_dff_A_gZDCfb638_0),.clk(gclk));
	jdff dff_A_e21azBOc4_0(.dout(w_dff_A_eUfihHxS6_0),.din(w_dff_A_e21azBOc4_0),.clk(gclk));
	jdff dff_A_eUfihHxS6_0(.dout(G406),.din(w_dff_A_eUfihHxS6_0),.clk(gclk));
	jdff dff_A_QqfC4UY36_1(.dout(w_dff_A_58tDZlpT4_0),.din(w_dff_A_QqfC4UY36_1),.clk(gclk));
	jdff dff_A_58tDZlpT4_0(.dout(w_dff_A_gjeEsi102_0),.din(w_dff_A_58tDZlpT4_0),.clk(gclk));
	jdff dff_A_gjeEsi102_0(.dout(w_dff_A_m3fq1gcI0_0),.din(w_dff_A_gjeEsi102_0),.clk(gclk));
	jdff dff_A_m3fq1gcI0_0(.dout(w_dff_A_687HZ5zR4_0),.din(w_dff_A_m3fq1gcI0_0),.clk(gclk));
	jdff dff_A_687HZ5zR4_0(.dout(w_dff_A_m1WaA9nU2_0),.din(w_dff_A_687HZ5zR4_0),.clk(gclk));
	jdff dff_A_m1WaA9nU2_0(.dout(w_dff_A_aSmhwjCD5_0),.din(w_dff_A_m1WaA9nU2_0),.clk(gclk));
	jdff dff_A_aSmhwjCD5_0(.dout(w_dff_A_iwZZDib65_0),.din(w_dff_A_aSmhwjCD5_0),.clk(gclk));
	jdff dff_A_iwZZDib65_0(.dout(w_dff_A_GKzRefx24_0),.din(w_dff_A_iwZZDib65_0),.clk(gclk));
	jdff dff_A_GKzRefx24_0(.dout(w_dff_A_jAb0X6Xd5_0),.din(w_dff_A_GKzRefx24_0),.clk(gclk));
	jdff dff_A_jAb0X6Xd5_0(.dout(w_dff_A_1yitxy5p3_0),.din(w_dff_A_jAb0X6Xd5_0),.clk(gclk));
	jdff dff_A_1yitxy5p3_0(.dout(w_dff_A_3d2dIPKw5_0),.din(w_dff_A_1yitxy5p3_0),.clk(gclk));
	jdff dff_A_3d2dIPKw5_0(.dout(w_dff_A_plu2t9V74_0),.din(w_dff_A_3d2dIPKw5_0),.clk(gclk));
	jdff dff_A_plu2t9V74_0(.dout(w_dff_A_zxxe1Bm74_0),.din(w_dff_A_plu2t9V74_0),.clk(gclk));
	jdff dff_A_zxxe1Bm74_0(.dout(w_dff_A_gTeWXvt37_0),.din(w_dff_A_zxxe1Bm74_0),.clk(gclk));
	jdff dff_A_gTeWXvt37_0(.dout(w_dff_A_Phyk4F5i4_0),.din(w_dff_A_gTeWXvt37_0),.clk(gclk));
	jdff dff_A_Phyk4F5i4_0(.dout(w_dff_A_tIXNc8o60_0),.din(w_dff_A_Phyk4F5i4_0),.clk(gclk));
	jdff dff_A_tIXNc8o60_0(.dout(w_dff_A_4S4oYqpz7_0),.din(w_dff_A_tIXNc8o60_0),.clk(gclk));
	jdff dff_A_4S4oYqpz7_0(.dout(w_dff_A_2F5jgnQF5_0),.din(w_dff_A_4S4oYqpz7_0),.clk(gclk));
	jdff dff_A_2F5jgnQF5_0(.dout(w_dff_A_DPYnJdeI3_0),.din(w_dff_A_2F5jgnQF5_0),.clk(gclk));
	jdff dff_A_DPYnJdeI3_0(.dout(w_dff_A_ekwhykXE1_0),.din(w_dff_A_DPYnJdeI3_0),.clk(gclk));
	jdff dff_A_ekwhykXE1_0(.dout(w_dff_A_B71DuFdv2_0),.din(w_dff_A_ekwhykXE1_0),.clk(gclk));
	jdff dff_A_B71DuFdv2_0(.dout(w_dff_A_fpcD7gLA1_0),.din(w_dff_A_B71DuFdv2_0),.clk(gclk));
	jdff dff_A_fpcD7gLA1_0(.dout(w_dff_A_j8DZDwYc3_0),.din(w_dff_A_fpcD7gLA1_0),.clk(gclk));
	jdff dff_A_j8DZDwYc3_0(.dout(G408),.din(w_dff_A_j8DZDwYc3_0),.clk(gclk));
	jdff dff_A_wN1COxFA1_1(.dout(w_dff_A_UXhXXOMd1_0),.din(w_dff_A_wN1COxFA1_1),.clk(gclk));
	jdff dff_A_UXhXXOMd1_0(.dout(w_dff_A_rNbJSLRS5_0),.din(w_dff_A_UXhXXOMd1_0),.clk(gclk));
	jdff dff_A_rNbJSLRS5_0(.dout(w_dff_A_tuQKwvRI1_0),.din(w_dff_A_rNbJSLRS5_0),.clk(gclk));
	jdff dff_A_tuQKwvRI1_0(.dout(w_dff_A_bKOgxtYK9_0),.din(w_dff_A_tuQKwvRI1_0),.clk(gclk));
	jdff dff_A_bKOgxtYK9_0(.dout(w_dff_A_7UzdgSs08_0),.din(w_dff_A_bKOgxtYK9_0),.clk(gclk));
	jdff dff_A_7UzdgSs08_0(.dout(w_dff_A_gdi3aaTK4_0),.din(w_dff_A_7UzdgSs08_0),.clk(gclk));
	jdff dff_A_gdi3aaTK4_0(.dout(w_dff_A_1I73ylGv1_0),.din(w_dff_A_gdi3aaTK4_0),.clk(gclk));
	jdff dff_A_1I73ylGv1_0(.dout(w_dff_A_tr8P846U6_0),.din(w_dff_A_1I73ylGv1_0),.clk(gclk));
	jdff dff_A_tr8P846U6_0(.dout(w_dff_A_jGtw6X0j1_0),.din(w_dff_A_tr8P846U6_0),.clk(gclk));
	jdff dff_A_jGtw6X0j1_0(.dout(w_dff_A_guz3Wv0c0_0),.din(w_dff_A_jGtw6X0j1_0),.clk(gclk));
	jdff dff_A_guz3Wv0c0_0(.dout(w_dff_A_HndTTY115_0),.din(w_dff_A_guz3Wv0c0_0),.clk(gclk));
	jdff dff_A_HndTTY115_0(.dout(w_dff_A_VnetsG9r8_0),.din(w_dff_A_HndTTY115_0),.clk(gclk));
	jdff dff_A_VnetsG9r8_0(.dout(w_dff_A_RW8JLp5w8_0),.din(w_dff_A_VnetsG9r8_0),.clk(gclk));
	jdff dff_A_RW8JLp5w8_0(.dout(w_dff_A_oLWOCoJM7_0),.din(w_dff_A_RW8JLp5w8_0),.clk(gclk));
	jdff dff_A_oLWOCoJM7_0(.dout(w_dff_A_zWtNHpzM6_0),.din(w_dff_A_oLWOCoJM7_0),.clk(gclk));
	jdff dff_A_zWtNHpzM6_0(.dout(w_dff_A_Kq3F9tLn8_0),.din(w_dff_A_zWtNHpzM6_0),.clk(gclk));
	jdff dff_A_Kq3F9tLn8_0(.dout(w_dff_A_YvYsigHO8_0),.din(w_dff_A_Kq3F9tLn8_0),.clk(gclk));
	jdff dff_A_YvYsigHO8_0(.dout(w_dff_A_zw8snAnD6_0),.din(w_dff_A_YvYsigHO8_0),.clk(gclk));
	jdff dff_A_zw8snAnD6_0(.dout(w_dff_A_tMdYx3le6_0),.din(w_dff_A_zw8snAnD6_0),.clk(gclk));
	jdff dff_A_tMdYx3le6_0(.dout(w_dff_A_eIxVDBlg5_0),.din(w_dff_A_tMdYx3le6_0),.clk(gclk));
	jdff dff_A_eIxVDBlg5_0(.dout(w_dff_A_g8CsW1aQ8_0),.din(w_dff_A_eIxVDBlg5_0),.clk(gclk));
	jdff dff_A_g8CsW1aQ8_0(.dout(w_dff_A_1qxbycY08_0),.din(w_dff_A_g8CsW1aQ8_0),.clk(gclk));
	jdff dff_A_1qxbycY08_0(.dout(w_dff_A_yW9PUCHW0_0),.din(w_dff_A_1qxbycY08_0),.clk(gclk));
	jdff dff_A_yW9PUCHW0_0(.dout(G410),.din(w_dff_A_yW9PUCHW0_0),.clk(gclk));
	jdff dff_A_bxKrKb576_1(.dout(w_dff_A_DOvQuR2g0_0),.din(w_dff_A_bxKrKb576_1),.clk(gclk));
	jdff dff_A_DOvQuR2g0_0(.dout(w_dff_A_seCvDu1X3_0),.din(w_dff_A_DOvQuR2g0_0),.clk(gclk));
	jdff dff_A_seCvDu1X3_0(.dout(w_dff_A_IhzefiQx5_0),.din(w_dff_A_seCvDu1X3_0),.clk(gclk));
	jdff dff_A_IhzefiQx5_0(.dout(w_dff_A_vpXS2Vdr8_0),.din(w_dff_A_IhzefiQx5_0),.clk(gclk));
	jdff dff_A_vpXS2Vdr8_0(.dout(w_dff_A_lFABJ5my6_0),.din(w_dff_A_vpXS2Vdr8_0),.clk(gclk));
	jdff dff_A_lFABJ5my6_0(.dout(w_dff_A_MQCWwP5C6_0),.din(w_dff_A_lFABJ5my6_0),.clk(gclk));
	jdff dff_A_MQCWwP5C6_0(.dout(w_dff_A_uDIsdkRv2_0),.din(w_dff_A_MQCWwP5C6_0),.clk(gclk));
	jdff dff_A_uDIsdkRv2_0(.dout(w_dff_A_5lO8EgHw1_0),.din(w_dff_A_uDIsdkRv2_0),.clk(gclk));
	jdff dff_A_5lO8EgHw1_0(.dout(w_dff_A_BwphV7pv4_0),.din(w_dff_A_5lO8EgHw1_0),.clk(gclk));
	jdff dff_A_BwphV7pv4_0(.dout(w_dff_A_rN8FldBp4_0),.din(w_dff_A_BwphV7pv4_0),.clk(gclk));
	jdff dff_A_rN8FldBp4_0(.dout(w_dff_A_722YTZtX6_0),.din(w_dff_A_rN8FldBp4_0),.clk(gclk));
	jdff dff_A_722YTZtX6_0(.dout(w_dff_A_JoVputvT0_0),.din(w_dff_A_722YTZtX6_0),.clk(gclk));
	jdff dff_A_JoVputvT0_0(.dout(w_dff_A_BUy5xOgU7_0),.din(w_dff_A_JoVputvT0_0),.clk(gclk));
	jdff dff_A_BUy5xOgU7_0(.dout(w_dff_A_ZUSa5Pzw9_0),.din(w_dff_A_BUy5xOgU7_0),.clk(gclk));
	jdff dff_A_ZUSa5Pzw9_0(.dout(w_dff_A_JsUWcN0v9_0),.din(w_dff_A_ZUSa5Pzw9_0),.clk(gclk));
	jdff dff_A_JsUWcN0v9_0(.dout(w_dff_A_vSBQXyM61_0),.din(w_dff_A_JsUWcN0v9_0),.clk(gclk));
	jdff dff_A_vSBQXyM61_0(.dout(w_dff_A_VoVKRvgu9_0),.din(w_dff_A_vSBQXyM61_0),.clk(gclk));
	jdff dff_A_VoVKRvgu9_0(.dout(w_dff_A_Cpcprkzt3_0),.din(w_dff_A_VoVKRvgu9_0),.clk(gclk));
	jdff dff_A_Cpcprkzt3_0(.dout(w_dff_A_ambPSS9G6_0),.din(w_dff_A_Cpcprkzt3_0),.clk(gclk));
	jdff dff_A_ambPSS9G6_0(.dout(w_dff_A_M3oNdF5o9_0),.din(w_dff_A_ambPSS9G6_0),.clk(gclk));
	jdff dff_A_M3oNdF5o9_0(.dout(w_dff_A_TpENOab82_0),.din(w_dff_A_M3oNdF5o9_0),.clk(gclk));
	jdff dff_A_TpENOab82_0(.dout(w_dff_A_orjNISZW6_0),.din(w_dff_A_TpENOab82_0),.clk(gclk));
	jdff dff_A_orjNISZW6_0(.dout(w_dff_A_HLEa5dzA4_0),.din(w_dff_A_orjNISZW6_0),.clk(gclk));
	jdff dff_A_HLEa5dzA4_0(.dout(w_dff_A_kJQVnKHp1_0),.din(w_dff_A_HLEa5dzA4_0),.clk(gclk));
	jdff dff_A_kJQVnKHp1_0(.dout(w_dff_A_DWZLgRVD1_0),.din(w_dff_A_kJQVnKHp1_0),.clk(gclk));
	jdff dff_A_DWZLgRVD1_0(.dout(w_dff_A_DNtqkJDi5_0),.din(w_dff_A_DWZLgRVD1_0),.clk(gclk));
	jdff dff_A_DNtqkJDi5_0(.dout(G432),.din(w_dff_A_DNtqkJDi5_0),.clk(gclk));
	jdff dff_A_lXPJgvRR0_1(.dout(w_dff_A_Qwp48rKC0_0),.din(w_dff_A_lXPJgvRR0_1),.clk(gclk));
	jdff dff_A_Qwp48rKC0_0(.dout(w_dff_A_61zFQQar8_0),.din(w_dff_A_Qwp48rKC0_0),.clk(gclk));
	jdff dff_A_61zFQQar8_0(.dout(w_dff_A_4Hbvc1QT5_0),.din(w_dff_A_61zFQQar8_0),.clk(gclk));
	jdff dff_A_4Hbvc1QT5_0(.dout(w_dff_A_b7OF5PqX4_0),.din(w_dff_A_4Hbvc1QT5_0),.clk(gclk));
	jdff dff_A_b7OF5PqX4_0(.dout(w_dff_A_yNZ0DHT43_0),.din(w_dff_A_b7OF5PqX4_0),.clk(gclk));
	jdff dff_A_yNZ0DHT43_0(.dout(w_dff_A_3Y0UdgSe4_0),.din(w_dff_A_yNZ0DHT43_0),.clk(gclk));
	jdff dff_A_3Y0UdgSe4_0(.dout(w_dff_A_D7FTGf7z9_0),.din(w_dff_A_3Y0UdgSe4_0),.clk(gclk));
	jdff dff_A_D7FTGf7z9_0(.dout(w_dff_A_ihh5PTuA2_0),.din(w_dff_A_D7FTGf7z9_0),.clk(gclk));
	jdff dff_A_ihh5PTuA2_0(.dout(w_dff_A_jgk8HQXv6_0),.din(w_dff_A_ihh5PTuA2_0),.clk(gclk));
	jdff dff_A_jgk8HQXv6_0(.dout(w_dff_A_u8CbI35r0_0),.din(w_dff_A_jgk8HQXv6_0),.clk(gclk));
	jdff dff_A_u8CbI35r0_0(.dout(w_dff_A_tb4djUUj7_0),.din(w_dff_A_u8CbI35r0_0),.clk(gclk));
	jdff dff_A_tb4djUUj7_0(.dout(w_dff_A_vHKDxMlm4_0),.din(w_dff_A_tb4djUUj7_0),.clk(gclk));
	jdff dff_A_vHKDxMlm4_0(.dout(w_dff_A_DCc2tDDX9_0),.din(w_dff_A_vHKDxMlm4_0),.clk(gclk));
	jdff dff_A_DCc2tDDX9_0(.dout(w_dff_A_IJH2Brp98_0),.din(w_dff_A_DCc2tDDX9_0),.clk(gclk));
	jdff dff_A_IJH2Brp98_0(.dout(w_dff_A_oT0rsEt19_0),.din(w_dff_A_IJH2Brp98_0),.clk(gclk));
	jdff dff_A_oT0rsEt19_0(.dout(w_dff_A_xhIDkBHd1_0),.din(w_dff_A_oT0rsEt19_0),.clk(gclk));
	jdff dff_A_xhIDkBHd1_0(.dout(w_dff_A_yvbSGFRa9_0),.din(w_dff_A_xhIDkBHd1_0),.clk(gclk));
	jdff dff_A_yvbSGFRa9_0(.dout(w_dff_A_p8j8ckKQ6_0),.din(w_dff_A_yvbSGFRa9_0),.clk(gclk));
	jdff dff_A_p8j8ckKQ6_0(.dout(w_dff_A_82lYXakP8_0),.din(w_dff_A_p8j8ckKQ6_0),.clk(gclk));
	jdff dff_A_82lYXakP8_0(.dout(w_dff_A_VTJIuf3R1_0),.din(w_dff_A_82lYXakP8_0),.clk(gclk));
	jdff dff_A_VTJIuf3R1_0(.dout(w_dff_A_d52LjHTs3_0),.din(w_dff_A_VTJIuf3R1_0),.clk(gclk));
	jdff dff_A_d52LjHTs3_0(.dout(w_dff_A_ZYyu616n8_0),.din(w_dff_A_d52LjHTs3_0),.clk(gclk));
	jdff dff_A_ZYyu616n8_0(.dout(w_dff_A_o1A1ZTF14_0),.din(w_dff_A_ZYyu616n8_0),.clk(gclk));
	jdff dff_A_o1A1ZTF14_0(.dout(w_dff_A_5t6PR8h28_0),.din(w_dff_A_o1A1ZTF14_0),.clk(gclk));
	jdff dff_A_5t6PR8h28_0(.dout(w_dff_A_maAE4afP8_0),.din(w_dff_A_5t6PR8h28_0),.clk(gclk));
	jdff dff_A_maAE4afP8_0(.dout(w_dff_A_MdPzYG3f5_0),.din(w_dff_A_maAE4afP8_0),.clk(gclk));
	jdff dff_A_MdPzYG3f5_0(.dout(G446),.din(w_dff_A_MdPzYG3f5_0),.clk(gclk));
	jdff dff_A_pZTZwLvs9_2(.dout(w_dff_A_uHCJWSLz2_0),.din(w_dff_A_pZTZwLvs9_2),.clk(gclk));
	jdff dff_A_uHCJWSLz2_0(.dout(w_dff_A_kqRh5e7s2_0),.din(w_dff_A_uHCJWSLz2_0),.clk(gclk));
	jdff dff_A_kqRh5e7s2_0(.dout(w_dff_A_WHezx8f96_0),.din(w_dff_A_kqRh5e7s2_0),.clk(gclk));
	jdff dff_A_WHezx8f96_0(.dout(w_dff_A_SorlaUJ19_0),.din(w_dff_A_WHezx8f96_0),.clk(gclk));
	jdff dff_A_SorlaUJ19_0(.dout(w_dff_A_BVxgosoN9_0),.din(w_dff_A_SorlaUJ19_0),.clk(gclk));
	jdff dff_A_BVxgosoN9_0(.dout(w_dff_A_mzyaUjDb2_0),.din(w_dff_A_BVxgosoN9_0),.clk(gclk));
	jdff dff_A_mzyaUjDb2_0(.dout(w_dff_A_bdtivdEl9_0),.din(w_dff_A_mzyaUjDb2_0),.clk(gclk));
	jdff dff_A_bdtivdEl9_0(.dout(w_dff_A_gerkpQKj0_0),.din(w_dff_A_bdtivdEl9_0),.clk(gclk));
	jdff dff_A_gerkpQKj0_0(.dout(w_dff_A_3eVzLDRo1_0),.din(w_dff_A_gerkpQKj0_0),.clk(gclk));
	jdff dff_A_3eVzLDRo1_0(.dout(w_dff_A_GAoxwLYc9_0),.din(w_dff_A_3eVzLDRo1_0),.clk(gclk));
	jdff dff_A_GAoxwLYc9_0(.dout(w_dff_A_kcHwxb6m7_0),.din(w_dff_A_GAoxwLYc9_0),.clk(gclk));
	jdff dff_A_kcHwxb6m7_0(.dout(w_dff_A_Q7x3eYi17_0),.din(w_dff_A_kcHwxb6m7_0),.clk(gclk));
	jdff dff_A_Q7x3eYi17_0(.dout(w_dff_A_668Mfmxb6_0),.din(w_dff_A_Q7x3eYi17_0),.clk(gclk));
	jdff dff_A_668Mfmxb6_0(.dout(w_dff_A_7GAbXbNd6_0),.din(w_dff_A_668Mfmxb6_0),.clk(gclk));
	jdff dff_A_7GAbXbNd6_0(.dout(w_dff_A_UiMGESzz3_0),.din(w_dff_A_7GAbXbNd6_0),.clk(gclk));
	jdff dff_A_UiMGESzz3_0(.dout(w_dff_A_C1Z9Z9Kw0_0),.din(w_dff_A_UiMGESzz3_0),.clk(gclk));
	jdff dff_A_C1Z9Z9Kw0_0(.dout(w_dff_A_EsggchHu8_0),.din(w_dff_A_C1Z9Z9Kw0_0),.clk(gclk));
	jdff dff_A_EsggchHu8_0(.dout(w_dff_A_8JVdgzId5_0),.din(w_dff_A_EsggchHu8_0),.clk(gclk));
	jdff dff_A_8JVdgzId5_0(.dout(w_dff_A_JffIFJ3K9_0),.din(w_dff_A_8JVdgzId5_0),.clk(gclk));
	jdff dff_A_JffIFJ3K9_0(.dout(w_dff_A_nfffUmky5_0),.din(w_dff_A_JffIFJ3K9_0),.clk(gclk));
	jdff dff_A_nfffUmky5_0(.dout(w_dff_A_QUuVqL9d8_0),.din(w_dff_A_nfffUmky5_0),.clk(gclk));
	jdff dff_A_QUuVqL9d8_0(.dout(w_dff_A_BsbD4sss9_0),.din(w_dff_A_QUuVqL9d8_0),.clk(gclk));
	jdff dff_A_BsbD4sss9_0(.dout(w_dff_A_YHeMACUH6_0),.din(w_dff_A_BsbD4sss9_0),.clk(gclk));
	jdff dff_A_YHeMACUH6_0(.dout(w_dff_A_MP5Q4Jtz3_0),.din(w_dff_A_YHeMACUH6_0),.clk(gclk));
	jdff dff_A_MP5Q4Jtz3_0(.dout(G284),.din(w_dff_A_MP5Q4Jtz3_0),.clk(gclk));
	jdff dff_A_eCUBokED4_1(.dout(w_dff_A_RnSNRzgX1_0),.din(w_dff_A_eCUBokED4_1),.clk(gclk));
	jdff dff_A_RnSNRzgX1_0(.dout(w_dff_A_bqKY1ank8_0),.din(w_dff_A_RnSNRzgX1_0),.clk(gclk));
	jdff dff_A_bqKY1ank8_0(.dout(w_dff_A_EAREiTWX9_0),.din(w_dff_A_bqKY1ank8_0),.clk(gclk));
	jdff dff_A_EAREiTWX9_0(.dout(w_dff_A_frUEwr0U4_0),.din(w_dff_A_EAREiTWX9_0),.clk(gclk));
	jdff dff_A_frUEwr0U4_0(.dout(w_dff_A_rMX5vMuu1_0),.din(w_dff_A_frUEwr0U4_0),.clk(gclk));
	jdff dff_A_rMX5vMuu1_0(.dout(w_dff_A_C1YHji7f5_0),.din(w_dff_A_rMX5vMuu1_0),.clk(gclk));
	jdff dff_A_C1YHji7f5_0(.dout(w_dff_A_9jxMTJDm4_0),.din(w_dff_A_C1YHji7f5_0),.clk(gclk));
	jdff dff_A_9jxMTJDm4_0(.dout(w_dff_A_z8WbIWXs3_0),.din(w_dff_A_9jxMTJDm4_0),.clk(gclk));
	jdff dff_A_z8WbIWXs3_0(.dout(w_dff_A_giDFloJd0_0),.din(w_dff_A_z8WbIWXs3_0),.clk(gclk));
	jdff dff_A_giDFloJd0_0(.dout(w_dff_A_VUJrQzoM0_0),.din(w_dff_A_giDFloJd0_0),.clk(gclk));
	jdff dff_A_VUJrQzoM0_0(.dout(w_dff_A_Jctpfofv4_0),.din(w_dff_A_VUJrQzoM0_0),.clk(gclk));
	jdff dff_A_Jctpfofv4_0(.dout(w_dff_A_GYEIOdVE0_0),.din(w_dff_A_Jctpfofv4_0),.clk(gclk));
	jdff dff_A_GYEIOdVE0_0(.dout(w_dff_A_5r0YoeG36_0),.din(w_dff_A_GYEIOdVE0_0),.clk(gclk));
	jdff dff_A_5r0YoeG36_0(.dout(w_dff_A_eZlf5nWa3_0),.din(w_dff_A_5r0YoeG36_0),.clk(gclk));
	jdff dff_A_eZlf5nWa3_0(.dout(w_dff_A_oD6ZDMiO5_0),.din(w_dff_A_eZlf5nWa3_0),.clk(gclk));
	jdff dff_A_oD6ZDMiO5_0(.dout(w_dff_A_YsrsOS6p4_0),.din(w_dff_A_oD6ZDMiO5_0),.clk(gclk));
	jdff dff_A_YsrsOS6p4_0(.dout(w_dff_A_ozKdBggJ7_0),.din(w_dff_A_YsrsOS6p4_0),.clk(gclk));
	jdff dff_A_ozKdBggJ7_0(.dout(w_dff_A_daKv7Bc13_0),.din(w_dff_A_ozKdBggJ7_0),.clk(gclk));
	jdff dff_A_daKv7Bc13_0(.dout(w_dff_A_jPAMB7SH8_0),.din(w_dff_A_daKv7Bc13_0),.clk(gclk));
	jdff dff_A_jPAMB7SH8_0(.dout(w_dff_A_pGBm3lmP3_0),.din(w_dff_A_jPAMB7SH8_0),.clk(gclk));
	jdff dff_A_pGBm3lmP3_0(.dout(w_dff_A_Nkq8LCm59_0),.din(w_dff_A_pGBm3lmP3_0),.clk(gclk));
	jdff dff_A_Nkq8LCm59_0(.dout(w_dff_A_78VAapmA2_0),.din(w_dff_A_Nkq8LCm59_0),.clk(gclk));
	jdff dff_A_78VAapmA2_0(.dout(w_dff_A_uO16OH9U4_0),.din(w_dff_A_78VAapmA2_0),.clk(gclk));
	jdff dff_A_uO16OH9U4_0(.dout(w_dff_A_CsoApEUQ3_0),.din(w_dff_A_uO16OH9U4_0),.clk(gclk));
	jdff dff_A_CsoApEUQ3_0(.dout(w_dff_A_AFPm4Vdq3_0),.din(w_dff_A_CsoApEUQ3_0),.clk(gclk));
	jdff dff_A_AFPm4Vdq3_0(.dout(G286),.din(w_dff_A_AFPm4Vdq3_0),.clk(gclk));
	jdff dff_A_FYQc2eRh8_2(.dout(w_dff_A_KLfJguYR5_0),.din(w_dff_A_FYQc2eRh8_2),.clk(gclk));
	jdff dff_A_KLfJguYR5_0(.dout(w_dff_A_2J5FgEL79_0),.din(w_dff_A_KLfJguYR5_0),.clk(gclk));
	jdff dff_A_2J5FgEL79_0(.dout(w_dff_A_ogUKhVPc4_0),.din(w_dff_A_2J5FgEL79_0),.clk(gclk));
	jdff dff_A_ogUKhVPc4_0(.dout(w_dff_A_IW9uyKCq2_0),.din(w_dff_A_ogUKhVPc4_0),.clk(gclk));
	jdff dff_A_IW9uyKCq2_0(.dout(w_dff_A_GTEHJHr11_0),.din(w_dff_A_IW9uyKCq2_0),.clk(gclk));
	jdff dff_A_GTEHJHr11_0(.dout(w_dff_A_P8N7C4kW6_0),.din(w_dff_A_GTEHJHr11_0),.clk(gclk));
	jdff dff_A_P8N7C4kW6_0(.dout(w_dff_A_BS1xp1Vg2_0),.din(w_dff_A_P8N7C4kW6_0),.clk(gclk));
	jdff dff_A_BS1xp1Vg2_0(.dout(w_dff_A_HtbMXH465_0),.din(w_dff_A_BS1xp1Vg2_0),.clk(gclk));
	jdff dff_A_HtbMXH465_0(.dout(w_dff_A_2WchYrdZ4_0),.din(w_dff_A_HtbMXH465_0),.clk(gclk));
	jdff dff_A_2WchYrdZ4_0(.dout(w_dff_A_WM9FRa6U2_0),.din(w_dff_A_2WchYrdZ4_0),.clk(gclk));
	jdff dff_A_WM9FRa6U2_0(.dout(w_dff_A_0wkvtvXM7_0),.din(w_dff_A_WM9FRa6U2_0),.clk(gclk));
	jdff dff_A_0wkvtvXM7_0(.dout(w_dff_A_5JJVyeKX7_0),.din(w_dff_A_0wkvtvXM7_0),.clk(gclk));
	jdff dff_A_5JJVyeKX7_0(.dout(w_dff_A_5u2NkGBQ0_0),.din(w_dff_A_5JJVyeKX7_0),.clk(gclk));
	jdff dff_A_5u2NkGBQ0_0(.dout(w_dff_A_HPoNnLaf9_0),.din(w_dff_A_5u2NkGBQ0_0),.clk(gclk));
	jdff dff_A_HPoNnLaf9_0(.dout(w_dff_A_zjM5TtBf8_0),.din(w_dff_A_HPoNnLaf9_0),.clk(gclk));
	jdff dff_A_zjM5TtBf8_0(.dout(w_dff_A_zKCY6qMT3_0),.din(w_dff_A_zjM5TtBf8_0),.clk(gclk));
	jdff dff_A_zKCY6qMT3_0(.dout(w_dff_A_ELSFogIC5_0),.din(w_dff_A_zKCY6qMT3_0),.clk(gclk));
	jdff dff_A_ELSFogIC5_0(.dout(w_dff_A_LE6gOCuF0_0),.din(w_dff_A_ELSFogIC5_0),.clk(gclk));
	jdff dff_A_LE6gOCuF0_0(.dout(w_dff_A_Xzaig07Y1_0),.din(w_dff_A_LE6gOCuF0_0),.clk(gclk));
	jdff dff_A_Xzaig07Y1_0(.dout(w_dff_A_ia8NrkBF7_0),.din(w_dff_A_Xzaig07Y1_0),.clk(gclk));
	jdff dff_A_ia8NrkBF7_0(.dout(w_dff_A_wVQwyipg4_0),.din(w_dff_A_ia8NrkBF7_0),.clk(gclk));
	jdff dff_A_wVQwyipg4_0(.dout(w_dff_A_SdCvp1Oi1_0),.din(w_dff_A_wVQwyipg4_0),.clk(gclk));
	jdff dff_A_SdCvp1Oi1_0(.dout(w_dff_A_aivzwgzo6_0),.din(w_dff_A_SdCvp1Oi1_0),.clk(gclk));
	jdff dff_A_aivzwgzo6_0(.dout(w_dff_A_SCWtELTJ2_0),.din(w_dff_A_aivzwgzo6_0),.clk(gclk));
	jdff dff_A_SCWtELTJ2_0(.dout(G289),.din(w_dff_A_SCWtELTJ2_0),.clk(gclk));
	jdff dff_A_ykhwGoNg6_2(.dout(w_dff_A_zYKSdpIZ3_0),.din(w_dff_A_ykhwGoNg6_2),.clk(gclk));
	jdff dff_A_zYKSdpIZ3_0(.dout(w_dff_A_OvmsZo7W9_0),.din(w_dff_A_zYKSdpIZ3_0),.clk(gclk));
	jdff dff_A_OvmsZo7W9_0(.dout(w_dff_A_ZeGmODYM2_0),.din(w_dff_A_OvmsZo7W9_0),.clk(gclk));
	jdff dff_A_ZeGmODYM2_0(.dout(w_dff_A_MHYM4iGP5_0),.din(w_dff_A_ZeGmODYM2_0),.clk(gclk));
	jdff dff_A_MHYM4iGP5_0(.dout(w_dff_A_XH2gTiXA7_0),.din(w_dff_A_MHYM4iGP5_0),.clk(gclk));
	jdff dff_A_XH2gTiXA7_0(.dout(w_dff_A_TCn667am8_0),.din(w_dff_A_XH2gTiXA7_0),.clk(gclk));
	jdff dff_A_TCn667am8_0(.dout(w_dff_A_PfiLlCQu8_0),.din(w_dff_A_TCn667am8_0),.clk(gclk));
	jdff dff_A_PfiLlCQu8_0(.dout(w_dff_A_lbb4ojyu0_0),.din(w_dff_A_PfiLlCQu8_0),.clk(gclk));
	jdff dff_A_lbb4ojyu0_0(.dout(w_dff_A_MJLIf0s93_0),.din(w_dff_A_lbb4ojyu0_0),.clk(gclk));
	jdff dff_A_MJLIf0s93_0(.dout(w_dff_A_puwKJnUy9_0),.din(w_dff_A_MJLIf0s93_0),.clk(gclk));
	jdff dff_A_puwKJnUy9_0(.dout(w_dff_A_yj5UMYdx5_0),.din(w_dff_A_puwKJnUy9_0),.clk(gclk));
	jdff dff_A_yj5UMYdx5_0(.dout(w_dff_A_Nta5g0kw6_0),.din(w_dff_A_yj5UMYdx5_0),.clk(gclk));
	jdff dff_A_Nta5g0kw6_0(.dout(w_dff_A_82BdCJjf1_0),.din(w_dff_A_Nta5g0kw6_0),.clk(gclk));
	jdff dff_A_82BdCJjf1_0(.dout(w_dff_A_l4yGPLa39_0),.din(w_dff_A_82BdCJjf1_0),.clk(gclk));
	jdff dff_A_l4yGPLa39_0(.dout(w_dff_A_iqME2LgY7_0),.din(w_dff_A_l4yGPLa39_0),.clk(gclk));
	jdff dff_A_iqME2LgY7_0(.dout(w_dff_A_l0iQdBqX3_0),.din(w_dff_A_iqME2LgY7_0),.clk(gclk));
	jdff dff_A_l0iQdBqX3_0(.dout(w_dff_A_cp4ruuO85_0),.din(w_dff_A_l0iQdBqX3_0),.clk(gclk));
	jdff dff_A_cp4ruuO85_0(.dout(w_dff_A_YDpNDwXu7_0),.din(w_dff_A_cp4ruuO85_0),.clk(gclk));
	jdff dff_A_YDpNDwXu7_0(.dout(w_dff_A_PliiTkmn7_0),.din(w_dff_A_YDpNDwXu7_0),.clk(gclk));
	jdff dff_A_PliiTkmn7_0(.dout(w_dff_A_BC2gfvBM3_0),.din(w_dff_A_PliiTkmn7_0),.clk(gclk));
	jdff dff_A_BC2gfvBM3_0(.dout(w_dff_A_GwSdQOOu6_0),.din(w_dff_A_BC2gfvBM3_0),.clk(gclk));
	jdff dff_A_GwSdQOOu6_0(.dout(w_dff_A_nPlPe1ob8_0),.din(w_dff_A_GwSdQOOu6_0),.clk(gclk));
	jdff dff_A_nPlPe1ob8_0(.dout(w_dff_A_LmjUrBmH6_0),.din(w_dff_A_nPlPe1ob8_0),.clk(gclk));
	jdff dff_A_LmjUrBmH6_0(.dout(G292),.din(w_dff_A_LmjUrBmH6_0),.clk(gclk));
	jdff dff_A_RVsCS7MB2_1(.dout(w_dff_A_JkGYnqp37_0),.din(w_dff_A_RVsCS7MB2_1),.clk(gclk));
	jdff dff_A_JkGYnqp37_0(.dout(w_dff_A_cfLyZ6Eo5_0),.din(w_dff_A_JkGYnqp37_0),.clk(gclk));
	jdff dff_A_cfLyZ6Eo5_0(.dout(w_dff_A_SZbOLmFu6_0),.din(w_dff_A_cfLyZ6Eo5_0),.clk(gclk));
	jdff dff_A_SZbOLmFu6_0(.dout(w_dff_A_iDp6iamO7_0),.din(w_dff_A_SZbOLmFu6_0),.clk(gclk));
	jdff dff_A_iDp6iamO7_0(.dout(w_dff_A_lHiyOdug9_0),.din(w_dff_A_iDp6iamO7_0),.clk(gclk));
	jdff dff_A_lHiyOdug9_0(.dout(w_dff_A_53a1d0Hl8_0),.din(w_dff_A_lHiyOdug9_0),.clk(gclk));
	jdff dff_A_53a1d0Hl8_0(.dout(w_dff_A_qKM3VT7L2_0),.din(w_dff_A_53a1d0Hl8_0),.clk(gclk));
	jdff dff_A_qKM3VT7L2_0(.dout(w_dff_A_i7Bvnpz17_0),.din(w_dff_A_qKM3VT7L2_0),.clk(gclk));
	jdff dff_A_i7Bvnpz17_0(.dout(w_dff_A_MEonsgzx3_0),.din(w_dff_A_i7Bvnpz17_0),.clk(gclk));
	jdff dff_A_MEonsgzx3_0(.dout(w_dff_A_rIlrQLfQ1_0),.din(w_dff_A_MEonsgzx3_0),.clk(gclk));
	jdff dff_A_rIlrQLfQ1_0(.dout(w_dff_A_w9Tvkphw0_0),.din(w_dff_A_rIlrQLfQ1_0),.clk(gclk));
	jdff dff_A_w9Tvkphw0_0(.dout(w_dff_A_5zMHCsLt9_0),.din(w_dff_A_w9Tvkphw0_0),.clk(gclk));
	jdff dff_A_5zMHCsLt9_0(.dout(w_dff_A_3iAiTpOV0_0),.din(w_dff_A_5zMHCsLt9_0),.clk(gclk));
	jdff dff_A_3iAiTpOV0_0(.dout(w_dff_A_6xOZ2zoO4_0),.din(w_dff_A_3iAiTpOV0_0),.clk(gclk));
	jdff dff_A_6xOZ2zoO4_0(.dout(w_dff_A_pW2OTON93_0),.din(w_dff_A_6xOZ2zoO4_0),.clk(gclk));
	jdff dff_A_pW2OTON93_0(.dout(w_dff_A_FDWcwLv91_0),.din(w_dff_A_pW2OTON93_0),.clk(gclk));
	jdff dff_A_FDWcwLv91_0(.dout(w_dff_A_Zt5yfqYZ8_0),.din(w_dff_A_FDWcwLv91_0),.clk(gclk));
	jdff dff_A_Zt5yfqYZ8_0(.dout(w_dff_A_WvD9IXS60_0),.din(w_dff_A_Zt5yfqYZ8_0),.clk(gclk));
	jdff dff_A_WvD9IXS60_0(.dout(w_dff_A_PTzSNQ7D1_0),.din(w_dff_A_WvD9IXS60_0),.clk(gclk));
	jdff dff_A_PTzSNQ7D1_0(.dout(w_dff_A_JqcPZAzv8_0),.din(w_dff_A_PTzSNQ7D1_0),.clk(gclk));
	jdff dff_A_JqcPZAzv8_0(.dout(w_dff_A_YJN1uq7d8_0),.din(w_dff_A_JqcPZAzv8_0),.clk(gclk));
	jdff dff_A_YJN1uq7d8_0(.dout(w_dff_A_LEKuSqlI2_0),.din(w_dff_A_YJN1uq7d8_0),.clk(gclk));
	jdff dff_A_LEKuSqlI2_0(.dout(w_dff_A_I6qbjVjc3_0),.din(w_dff_A_LEKuSqlI2_0),.clk(gclk));
	jdff dff_A_I6qbjVjc3_0(.dout(w_dff_A_SyOqRWI99_0),.din(w_dff_A_I6qbjVjc3_0),.clk(gclk));
	jdff dff_A_SyOqRWI99_0(.dout(w_dff_A_41YS9oF26_0),.din(w_dff_A_SyOqRWI99_0),.clk(gclk));
	jdff dff_A_41YS9oF26_0(.dout(G341),.din(w_dff_A_41YS9oF26_0),.clk(gclk));
	jdff dff_A_waTYV5cR5_2(.dout(w_dff_A_izDvKc0i8_0),.din(w_dff_A_waTYV5cR5_2),.clk(gclk));
	jdff dff_A_izDvKc0i8_0(.dout(w_dff_A_C2iaPpQG5_0),.din(w_dff_A_izDvKc0i8_0),.clk(gclk));
	jdff dff_A_C2iaPpQG5_0(.dout(w_dff_A_WuyTt3mA2_0),.din(w_dff_A_C2iaPpQG5_0),.clk(gclk));
	jdff dff_A_WuyTt3mA2_0(.dout(w_dff_A_m9gheg8O1_0),.din(w_dff_A_WuyTt3mA2_0),.clk(gclk));
	jdff dff_A_m9gheg8O1_0(.dout(w_dff_A_uGqKwkWM7_0),.din(w_dff_A_m9gheg8O1_0),.clk(gclk));
	jdff dff_A_uGqKwkWM7_0(.dout(w_dff_A_YLXpkA7n9_0),.din(w_dff_A_uGqKwkWM7_0),.clk(gclk));
	jdff dff_A_YLXpkA7n9_0(.dout(w_dff_A_uOEKxG5v5_0),.din(w_dff_A_YLXpkA7n9_0),.clk(gclk));
	jdff dff_A_uOEKxG5v5_0(.dout(w_dff_A_TCRqD5Xv5_0),.din(w_dff_A_uOEKxG5v5_0),.clk(gclk));
	jdff dff_A_TCRqD5Xv5_0(.dout(w_dff_A_kXB3zvQ49_0),.din(w_dff_A_TCRqD5Xv5_0),.clk(gclk));
	jdff dff_A_kXB3zvQ49_0(.dout(w_dff_A_x4VsyKIq4_0),.din(w_dff_A_kXB3zvQ49_0),.clk(gclk));
	jdff dff_A_x4VsyKIq4_0(.dout(w_dff_A_jT5HZZph8_0),.din(w_dff_A_x4VsyKIq4_0),.clk(gclk));
	jdff dff_A_jT5HZZph8_0(.dout(w_dff_A_u34PkPXl5_0),.din(w_dff_A_jT5HZZph8_0),.clk(gclk));
	jdff dff_A_u34PkPXl5_0(.dout(w_dff_A_nJlLwVJu7_0),.din(w_dff_A_u34PkPXl5_0),.clk(gclk));
	jdff dff_A_nJlLwVJu7_0(.dout(w_dff_A_Xl74Pygk4_0),.din(w_dff_A_nJlLwVJu7_0),.clk(gclk));
	jdff dff_A_Xl74Pygk4_0(.dout(w_dff_A_i8rVA1lx6_0),.din(w_dff_A_Xl74Pygk4_0),.clk(gclk));
	jdff dff_A_i8rVA1lx6_0(.dout(w_dff_A_AL0ZVEBo8_0),.din(w_dff_A_i8rVA1lx6_0),.clk(gclk));
	jdff dff_A_AL0ZVEBo8_0(.dout(w_dff_A_8jGHLbsB9_0),.din(w_dff_A_AL0ZVEBo8_0),.clk(gclk));
	jdff dff_A_8jGHLbsB9_0(.dout(w_dff_A_2JJUyQSP0_0),.din(w_dff_A_8jGHLbsB9_0),.clk(gclk));
	jdff dff_A_2JJUyQSP0_0(.dout(w_dff_A_QSZQQ8Fx5_0),.din(w_dff_A_2JJUyQSP0_0),.clk(gclk));
	jdff dff_A_QSZQQ8Fx5_0(.dout(w_dff_A_f6GMjrkO1_0),.din(w_dff_A_QSZQQ8Fx5_0),.clk(gclk));
	jdff dff_A_f6GMjrkO1_0(.dout(w_dff_A_uEYRmXI90_0),.din(w_dff_A_f6GMjrkO1_0),.clk(gclk));
	jdff dff_A_uEYRmXI90_0(.dout(w_dff_A_q600awFH0_0),.din(w_dff_A_uEYRmXI90_0),.clk(gclk));
	jdff dff_A_q600awFH0_0(.dout(w_dff_A_stwab5bd3_0),.din(w_dff_A_q600awFH0_0),.clk(gclk));
	jdff dff_A_stwab5bd3_0(.dout(G281),.din(w_dff_A_stwab5bd3_0),.clk(gclk));
	jdff dff_A_fFEFrf1N6_1(.dout(w_dff_A_ePGjtmuI1_0),.din(w_dff_A_fFEFrf1N6_1),.clk(gclk));
	jdff dff_A_ePGjtmuI1_0(.dout(w_dff_A_05KYiG352_0),.din(w_dff_A_ePGjtmuI1_0),.clk(gclk));
	jdff dff_A_05KYiG352_0(.dout(w_dff_A_BHdTPs5J3_0),.din(w_dff_A_05KYiG352_0),.clk(gclk));
	jdff dff_A_BHdTPs5J3_0(.dout(w_dff_A_FVSLWOXv1_0),.din(w_dff_A_BHdTPs5J3_0),.clk(gclk));
	jdff dff_A_FVSLWOXv1_0(.dout(w_dff_A_gk9Bxukh2_0),.din(w_dff_A_FVSLWOXv1_0),.clk(gclk));
	jdff dff_A_gk9Bxukh2_0(.dout(w_dff_A_qWmYEwaA2_0),.din(w_dff_A_gk9Bxukh2_0),.clk(gclk));
	jdff dff_A_qWmYEwaA2_0(.dout(w_dff_A_0TFtlHzA5_0),.din(w_dff_A_qWmYEwaA2_0),.clk(gclk));
	jdff dff_A_0TFtlHzA5_0(.dout(w_dff_A_Vd2UvW9V4_0),.din(w_dff_A_0TFtlHzA5_0),.clk(gclk));
	jdff dff_A_Vd2UvW9V4_0(.dout(w_dff_A_vu7rD0D33_0),.din(w_dff_A_Vd2UvW9V4_0),.clk(gclk));
	jdff dff_A_vu7rD0D33_0(.dout(w_dff_A_L3nmsKUv4_0),.din(w_dff_A_vu7rD0D33_0),.clk(gclk));
	jdff dff_A_L3nmsKUv4_0(.dout(w_dff_A_1BwNLuVf4_0),.din(w_dff_A_L3nmsKUv4_0),.clk(gclk));
	jdff dff_A_1BwNLuVf4_0(.dout(w_dff_A_CThb3KVb2_0),.din(w_dff_A_1BwNLuVf4_0),.clk(gclk));
	jdff dff_A_CThb3KVb2_0(.dout(w_dff_A_8bUTNctd4_0),.din(w_dff_A_CThb3KVb2_0),.clk(gclk));
	jdff dff_A_8bUTNctd4_0(.dout(w_dff_A_w8uLVGec0_0),.din(w_dff_A_8bUTNctd4_0),.clk(gclk));
	jdff dff_A_w8uLVGec0_0(.dout(w_dff_A_ngPergAi7_0),.din(w_dff_A_w8uLVGec0_0),.clk(gclk));
	jdff dff_A_ngPergAi7_0(.dout(w_dff_A_QJrkdR7R0_0),.din(w_dff_A_ngPergAi7_0),.clk(gclk));
	jdff dff_A_QJrkdR7R0_0(.dout(w_dff_A_ircsX5gO4_0),.din(w_dff_A_QJrkdR7R0_0),.clk(gclk));
	jdff dff_A_ircsX5gO4_0(.dout(w_dff_A_tVAvbdUP7_0),.din(w_dff_A_ircsX5gO4_0),.clk(gclk));
	jdff dff_A_tVAvbdUP7_0(.dout(w_dff_A_Ppvba4146_0),.din(w_dff_A_tVAvbdUP7_0),.clk(gclk));
	jdff dff_A_Ppvba4146_0(.dout(w_dff_A_7hflrjqg9_0),.din(w_dff_A_Ppvba4146_0),.clk(gclk));
	jdff dff_A_7hflrjqg9_0(.dout(w_dff_A_4CSQxZGI3_0),.din(w_dff_A_7hflrjqg9_0),.clk(gclk));
	jdff dff_A_4CSQxZGI3_0(.dout(w_dff_A_rVXUJMHr0_0),.din(w_dff_A_4CSQxZGI3_0),.clk(gclk));
	jdff dff_A_rVXUJMHr0_0(.dout(w_dff_A_2ezQkJns7_0),.din(w_dff_A_rVXUJMHr0_0),.clk(gclk));
	jdff dff_A_2ezQkJns7_0(.dout(w_dff_A_dqs0LX706_0),.din(w_dff_A_2ezQkJns7_0),.clk(gclk));
	jdff dff_A_dqs0LX706_0(.dout(w_dff_A_kxQ9F6iF6_0),.din(w_dff_A_dqs0LX706_0),.clk(gclk));
	jdff dff_A_kxQ9F6iF6_0(.dout(w_dff_A_lIGWgudn4_0),.din(w_dff_A_kxQ9F6iF6_0),.clk(gclk));
	jdff dff_A_lIGWgudn4_0(.dout(G453),.din(w_dff_A_lIGWgudn4_0),.clk(gclk));
	jdff dff_A_SPuBfask4_2(.dout(w_dff_A_rbNpX5TS7_0),.din(w_dff_A_SPuBfask4_2),.clk(gclk));
	jdff dff_A_rbNpX5TS7_0(.dout(w_dff_A_rrknosF80_0),.din(w_dff_A_rbNpX5TS7_0),.clk(gclk));
	jdff dff_A_rrknosF80_0(.dout(w_dff_A_5629ZiVs6_0),.din(w_dff_A_rrknosF80_0),.clk(gclk));
	jdff dff_A_5629ZiVs6_0(.dout(w_dff_A_183cX33w5_0),.din(w_dff_A_5629ZiVs6_0),.clk(gclk));
	jdff dff_A_183cX33w5_0(.dout(w_dff_A_PYToVF158_0),.din(w_dff_A_183cX33w5_0),.clk(gclk));
	jdff dff_A_PYToVF158_0(.dout(w_dff_A_7Kh27GAg9_0),.din(w_dff_A_PYToVF158_0),.clk(gclk));
	jdff dff_A_7Kh27GAg9_0(.dout(w_dff_A_OHaUO1y64_0),.din(w_dff_A_7Kh27GAg9_0),.clk(gclk));
	jdff dff_A_OHaUO1y64_0(.dout(w_dff_A_Bo04xigm6_0),.din(w_dff_A_OHaUO1y64_0),.clk(gclk));
	jdff dff_A_Bo04xigm6_0(.dout(w_dff_A_H75SOTxV2_0),.din(w_dff_A_Bo04xigm6_0),.clk(gclk));
	jdff dff_A_H75SOTxV2_0(.dout(w_dff_A_2wzeLbk01_0),.din(w_dff_A_H75SOTxV2_0),.clk(gclk));
	jdff dff_A_2wzeLbk01_0(.dout(w_dff_A_bic1SOq49_0),.din(w_dff_A_2wzeLbk01_0),.clk(gclk));
	jdff dff_A_bic1SOq49_0(.dout(w_dff_A_wUBKt1Ue2_0),.din(w_dff_A_bic1SOq49_0),.clk(gclk));
	jdff dff_A_wUBKt1Ue2_0(.dout(w_dff_A_nrCKNOix1_0),.din(w_dff_A_wUBKt1Ue2_0),.clk(gclk));
	jdff dff_A_nrCKNOix1_0(.dout(w_dff_A_ocV9Ai8E3_0),.din(w_dff_A_nrCKNOix1_0),.clk(gclk));
	jdff dff_A_ocV9Ai8E3_0(.dout(w_dff_A_gnfs6vU70_0),.din(w_dff_A_ocV9Ai8E3_0),.clk(gclk));
	jdff dff_A_gnfs6vU70_0(.dout(w_dff_A_yzmGzPvZ4_0),.din(w_dff_A_gnfs6vU70_0),.clk(gclk));
	jdff dff_A_yzmGzPvZ4_0(.dout(w_dff_A_ykuUuQvB5_0),.din(w_dff_A_yzmGzPvZ4_0),.clk(gclk));
	jdff dff_A_ykuUuQvB5_0(.dout(w_dff_A_HUfBXmwX9_0),.din(w_dff_A_ykuUuQvB5_0),.clk(gclk));
	jdff dff_A_HUfBXmwX9_0(.dout(w_dff_A_wYMGb9mr3_0),.din(w_dff_A_HUfBXmwX9_0),.clk(gclk));
	jdff dff_A_wYMGb9mr3_0(.dout(w_dff_A_EVOOIMjv0_0),.din(w_dff_A_wYMGb9mr3_0),.clk(gclk));
	jdff dff_A_EVOOIMjv0_0(.dout(w_dff_A_NZKV8M4g0_0),.din(w_dff_A_EVOOIMjv0_0),.clk(gclk));
	jdff dff_A_NZKV8M4g0_0(.dout(w_dff_A_pQ1BT9QM1_0),.din(w_dff_A_NZKV8M4g0_0),.clk(gclk));
	jdff dff_A_pQ1BT9QM1_0(.dout(w_dff_A_67PhyOSU5_0),.din(w_dff_A_pQ1BT9QM1_0),.clk(gclk));
	jdff dff_A_67PhyOSU5_0(.dout(w_dff_A_Y1zM5GUK2_0),.din(w_dff_A_67PhyOSU5_0),.clk(gclk));
	jdff dff_A_Y1zM5GUK2_0(.dout(w_dff_A_z14xZSHc4_0),.din(w_dff_A_Y1zM5GUK2_0),.clk(gclk));
	jdff dff_A_z14xZSHc4_0(.dout(G278),.din(w_dff_A_z14xZSHc4_0),.clk(gclk));
	jdff dff_A_suIs7AHU8_2(.dout(w_dff_A_Zl7v79IQ9_0),.din(w_dff_A_suIs7AHU8_2),.clk(gclk));
	jdff dff_A_Zl7v79IQ9_0(.dout(w_dff_A_PETjAI8f2_0),.din(w_dff_A_Zl7v79IQ9_0),.clk(gclk));
	jdff dff_A_PETjAI8f2_0(.dout(w_dff_A_l9oPxLRk8_0),.din(w_dff_A_PETjAI8f2_0),.clk(gclk));
	jdff dff_A_l9oPxLRk8_0(.dout(w_dff_A_AVwQQI0p1_0),.din(w_dff_A_l9oPxLRk8_0),.clk(gclk));
	jdff dff_A_AVwQQI0p1_0(.dout(w_dff_A_NhV9N0yC4_0),.din(w_dff_A_AVwQQI0p1_0),.clk(gclk));
	jdff dff_A_NhV9N0yC4_0(.dout(w_dff_A_OJc5aHP87_0),.din(w_dff_A_NhV9N0yC4_0),.clk(gclk));
	jdff dff_A_OJc5aHP87_0(.dout(w_dff_A_hlpsEyBO5_0),.din(w_dff_A_OJc5aHP87_0),.clk(gclk));
	jdff dff_A_hlpsEyBO5_0(.dout(w_dff_A_RFjQIz3m1_0),.din(w_dff_A_hlpsEyBO5_0),.clk(gclk));
	jdff dff_A_RFjQIz3m1_0(.dout(w_dff_A_oemZXJFF6_0),.din(w_dff_A_RFjQIz3m1_0),.clk(gclk));
	jdff dff_A_oemZXJFF6_0(.dout(w_dff_A_5mSVcpfS8_0),.din(w_dff_A_oemZXJFF6_0),.clk(gclk));
	jdff dff_A_5mSVcpfS8_0(.dout(w_dff_A_aTFF7Bz75_0),.din(w_dff_A_5mSVcpfS8_0),.clk(gclk));
	jdff dff_A_aTFF7Bz75_0(.dout(w_dff_A_llvpSK2r4_0),.din(w_dff_A_aTFF7Bz75_0),.clk(gclk));
	jdff dff_A_llvpSK2r4_0(.dout(w_dff_A_7P89TQuY2_0),.din(w_dff_A_llvpSK2r4_0),.clk(gclk));
	jdff dff_A_7P89TQuY2_0(.dout(w_dff_A_z6e0Xm7G4_0),.din(w_dff_A_7P89TQuY2_0),.clk(gclk));
	jdff dff_A_z6e0Xm7G4_0(.dout(w_dff_A_iQK2QjP91_0),.din(w_dff_A_z6e0Xm7G4_0),.clk(gclk));
	jdff dff_A_iQK2QjP91_0(.dout(w_dff_A_i8PkzgsH9_0),.din(w_dff_A_iQK2QjP91_0),.clk(gclk));
	jdff dff_A_i8PkzgsH9_0(.dout(w_dff_A_CukQvbtM3_0),.din(w_dff_A_i8PkzgsH9_0),.clk(gclk));
	jdff dff_A_CukQvbtM3_0(.dout(w_dff_A_zwu4hvFi6_0),.din(w_dff_A_CukQvbtM3_0),.clk(gclk));
	jdff dff_A_zwu4hvFi6_0(.dout(w_dff_A_K9vaKYfA5_0),.din(w_dff_A_zwu4hvFi6_0),.clk(gclk));
	jdff dff_A_K9vaKYfA5_0(.dout(w_dff_A_1hd6NNdi5_0),.din(w_dff_A_K9vaKYfA5_0),.clk(gclk));
	jdff dff_A_1hd6NNdi5_0(.dout(G373),.din(w_dff_A_1hd6NNdi5_0),.clk(gclk));
	jdff dff_A_JtpzOXIh8_2(.dout(G246),.din(w_dff_A_JtpzOXIh8_2),.clk(gclk));
	jdff dff_A_W0B7nnBb3_2(.dout(w_dff_A_zlWXXEha6_0),.din(w_dff_A_W0B7nnBb3_2),.clk(gclk));
	jdff dff_A_zlWXXEha6_0(.dout(w_dff_A_cEnFVj2R0_0),.din(w_dff_A_zlWXXEha6_0),.clk(gclk));
	jdff dff_A_cEnFVj2R0_0(.dout(w_dff_A_PTYC8VVJ5_0),.din(w_dff_A_cEnFVj2R0_0),.clk(gclk));
	jdff dff_A_PTYC8VVJ5_0(.dout(w_dff_A_IAWs3H189_0),.din(w_dff_A_PTYC8VVJ5_0),.clk(gclk));
	jdff dff_A_IAWs3H189_0(.dout(w_dff_A_opnM4RV00_0),.din(w_dff_A_IAWs3H189_0),.clk(gclk));
	jdff dff_A_opnM4RV00_0(.dout(w_dff_A_atu7ZuN71_0),.din(w_dff_A_opnM4RV00_0),.clk(gclk));
	jdff dff_A_atu7ZuN71_0(.dout(G258),.din(w_dff_A_atu7ZuN71_0),.clk(gclk));
	jdff dff_A_5YJ3wHUN2_2(.dout(w_dff_A_8CNtwnPS2_0),.din(w_dff_A_5YJ3wHUN2_2),.clk(gclk));
	jdff dff_A_8CNtwnPS2_0(.dout(w_dff_A_DueYmvrc5_0),.din(w_dff_A_8CNtwnPS2_0),.clk(gclk));
	jdff dff_A_DueYmvrc5_0(.dout(w_dff_A_Nou3FzeV2_0),.din(w_dff_A_DueYmvrc5_0),.clk(gclk));
	jdff dff_A_Nou3FzeV2_0(.dout(w_dff_A_BKstMjwm9_0),.din(w_dff_A_Nou3FzeV2_0),.clk(gclk));
	jdff dff_A_BKstMjwm9_0(.dout(w_dff_A_sVr04Vhk7_0),.din(w_dff_A_BKstMjwm9_0),.clk(gclk));
	jdff dff_A_sVr04Vhk7_0(.dout(w_dff_A_f2arjRAU3_0),.din(w_dff_A_sVr04Vhk7_0),.clk(gclk));
	jdff dff_A_f2arjRAU3_0(.dout(G264),.din(w_dff_A_f2arjRAU3_0),.clk(gclk));
	jdff dff_A_FnZbY9aw9_2(.dout(G270),.din(w_dff_A_FnZbY9aw9_2),.clk(gclk));
	jdff dff_A_EFX9NOPw8_2(.dout(w_dff_A_lAfW20ax2_0),.din(w_dff_A_EFX9NOPw8_2),.clk(gclk));
	jdff dff_A_lAfW20ax2_0(.dout(w_dff_A_ZFHJvkG30_0),.din(w_dff_A_lAfW20ax2_0),.clk(gclk));
	jdff dff_A_ZFHJvkG30_0(.dout(w_dff_A_1vOj1xHI3_0),.din(w_dff_A_ZFHJvkG30_0),.clk(gclk));
	jdff dff_A_1vOj1xHI3_0(.dout(w_dff_A_IdmYffwd3_0),.din(w_dff_A_1vOj1xHI3_0),.clk(gclk));
	jdff dff_A_IdmYffwd3_0(.dout(w_dff_A_ZF7HLi277_0),.din(w_dff_A_IdmYffwd3_0),.clk(gclk));
	jdff dff_A_ZF7HLi277_0(.dout(w_dff_A_f6pOu2Od7_0),.din(w_dff_A_ZF7HLi277_0),.clk(gclk));
	jdff dff_A_f6pOu2Od7_0(.dout(w_dff_A_I3jd4brz3_0),.din(w_dff_A_f6pOu2Od7_0),.clk(gclk));
	jdff dff_A_I3jd4brz3_0(.dout(w_dff_A_fhRfHGXa2_0),.din(w_dff_A_I3jd4brz3_0),.clk(gclk));
	jdff dff_A_fhRfHGXa2_0(.dout(w_dff_A_nuIUhyMq8_0),.din(w_dff_A_fhRfHGXa2_0),.clk(gclk));
	jdff dff_A_nuIUhyMq8_0(.dout(w_dff_A_zwFTOozw9_0),.din(w_dff_A_nuIUhyMq8_0),.clk(gclk));
	jdff dff_A_zwFTOozw9_0(.dout(w_dff_A_R2BZc8dp6_0),.din(w_dff_A_zwFTOozw9_0),.clk(gclk));
	jdff dff_A_R2BZc8dp6_0(.dout(w_dff_A_PcmfU9xn5_0),.din(w_dff_A_R2BZc8dp6_0),.clk(gclk));
	jdff dff_A_PcmfU9xn5_0(.dout(w_dff_A_L0s6fA2O4_0),.din(w_dff_A_PcmfU9xn5_0),.clk(gclk));
	jdff dff_A_L0s6fA2O4_0(.dout(w_dff_A_vvm9IkcB8_0),.din(w_dff_A_L0s6fA2O4_0),.clk(gclk));
	jdff dff_A_vvm9IkcB8_0(.dout(G388),.din(w_dff_A_vvm9IkcB8_0),.clk(gclk));
	jdff dff_A_xvoXLmi80_2(.dout(w_dff_A_t1IMydfR8_0),.din(w_dff_A_xvoXLmi80_2),.clk(gclk));
	jdff dff_A_t1IMydfR8_0(.dout(w_dff_A_ywwcwF1e8_0),.din(w_dff_A_t1IMydfR8_0),.clk(gclk));
	jdff dff_A_ywwcwF1e8_0(.dout(w_dff_A_deLvbHvC9_0),.din(w_dff_A_ywwcwF1e8_0),.clk(gclk));
	jdff dff_A_deLvbHvC9_0(.dout(w_dff_A_xn75DcLZ9_0),.din(w_dff_A_deLvbHvC9_0),.clk(gclk));
	jdff dff_A_xn75DcLZ9_0(.dout(w_dff_A_62RcKnEW0_0),.din(w_dff_A_xn75DcLZ9_0),.clk(gclk));
	jdff dff_A_62RcKnEW0_0(.dout(w_dff_A_FFtHcsj90_0),.din(w_dff_A_62RcKnEW0_0),.clk(gclk));
	jdff dff_A_FFtHcsj90_0(.dout(w_dff_A_OoHBHvrF2_0),.din(w_dff_A_FFtHcsj90_0),.clk(gclk));
	jdff dff_A_OoHBHvrF2_0(.dout(w_dff_A_cALSsssT3_0),.din(w_dff_A_OoHBHvrF2_0),.clk(gclk));
	jdff dff_A_cALSsssT3_0(.dout(w_dff_A_9gzshRGi6_0),.din(w_dff_A_cALSsssT3_0),.clk(gclk));
	jdff dff_A_9gzshRGi6_0(.dout(w_dff_A_mOTFYfuF1_0),.din(w_dff_A_9gzshRGi6_0),.clk(gclk));
	jdff dff_A_mOTFYfuF1_0(.dout(w_dff_A_bEzimCrj0_0),.din(w_dff_A_mOTFYfuF1_0),.clk(gclk));
	jdff dff_A_bEzimCrj0_0(.dout(w_dff_A_vVe9MpS49_0),.din(w_dff_A_bEzimCrj0_0),.clk(gclk));
	jdff dff_A_vVe9MpS49_0(.dout(w_dff_A_KicLbHz72_0),.din(w_dff_A_vVe9MpS49_0),.clk(gclk));
	jdff dff_A_KicLbHz72_0(.dout(w_dff_A_JiPxb9tQ0_0),.din(w_dff_A_KicLbHz72_0),.clk(gclk));
	jdff dff_A_JiPxb9tQ0_0(.dout(w_dff_A_wU0cGKNP1_0),.din(w_dff_A_JiPxb9tQ0_0),.clk(gclk));
	jdff dff_A_wU0cGKNP1_0(.dout(w_dff_A_uWOxwEd42_0),.din(w_dff_A_wU0cGKNP1_0),.clk(gclk));
	jdff dff_A_uWOxwEd42_0(.dout(G391),.din(w_dff_A_uWOxwEd42_0),.clk(gclk));
	jdff dff_A_7MoqT9H23_2(.dout(w_dff_A_B46vVDxc7_0),.din(w_dff_A_7MoqT9H23_2),.clk(gclk));
	jdff dff_A_B46vVDxc7_0(.dout(w_dff_A_6NKRiTk75_0),.din(w_dff_A_B46vVDxc7_0),.clk(gclk));
	jdff dff_A_6NKRiTk75_0(.dout(w_dff_A_yOUlHH040_0),.din(w_dff_A_6NKRiTk75_0),.clk(gclk));
	jdff dff_A_yOUlHH040_0(.dout(w_dff_A_CDEzwtfL8_0),.din(w_dff_A_yOUlHH040_0),.clk(gclk));
	jdff dff_A_CDEzwtfL8_0(.dout(w_dff_A_cBqXkpBh4_0),.din(w_dff_A_CDEzwtfL8_0),.clk(gclk));
	jdff dff_A_cBqXkpBh4_0(.dout(w_dff_A_IcxbCaoa2_0),.din(w_dff_A_cBqXkpBh4_0),.clk(gclk));
	jdff dff_A_IcxbCaoa2_0(.dout(w_dff_A_YAu1NTss0_0),.din(w_dff_A_IcxbCaoa2_0),.clk(gclk));
	jdff dff_A_YAu1NTss0_0(.dout(w_dff_A_JEBvJAwg2_0),.din(w_dff_A_YAu1NTss0_0),.clk(gclk));
	jdff dff_A_JEBvJAwg2_0(.dout(w_dff_A_NGIN4VwU8_0),.din(w_dff_A_JEBvJAwg2_0),.clk(gclk));
	jdff dff_A_NGIN4VwU8_0(.dout(w_dff_A_KiDmOa0U3_0),.din(w_dff_A_NGIN4VwU8_0),.clk(gclk));
	jdff dff_A_KiDmOa0U3_0(.dout(w_dff_A_ENP4IxIW6_0),.din(w_dff_A_KiDmOa0U3_0),.clk(gclk));
	jdff dff_A_ENP4IxIW6_0(.dout(w_dff_A_0YB5Jr5P4_0),.din(w_dff_A_ENP4IxIW6_0),.clk(gclk));
	jdff dff_A_0YB5Jr5P4_0(.dout(w_dff_A_1qWRxIx40_0),.din(w_dff_A_0YB5Jr5P4_0),.clk(gclk));
	jdff dff_A_1qWRxIx40_0(.dout(w_dff_A_IJO3GBE61_0),.din(w_dff_A_1qWRxIx40_0),.clk(gclk));
	jdff dff_A_IJO3GBE61_0(.dout(w_dff_A_zw4vaEnL5_0),.din(w_dff_A_IJO3GBE61_0),.clk(gclk));
	jdff dff_A_zw4vaEnL5_0(.dout(w_dff_A_udJWUOW08_0),.din(w_dff_A_zw4vaEnL5_0),.clk(gclk));
	jdff dff_A_udJWUOW08_0(.dout(w_dff_A_0LrTun7G6_0),.din(w_dff_A_udJWUOW08_0),.clk(gclk));
	jdff dff_A_0LrTun7G6_0(.dout(G394),.din(w_dff_A_0LrTun7G6_0),.clk(gclk));
	jdff dff_A_iAHGgVal8_2(.dout(w_dff_A_I74EMTpF6_0),.din(w_dff_A_iAHGgVal8_2),.clk(gclk));
	jdff dff_A_I74EMTpF6_0(.dout(w_dff_A_Cf6IPG4M3_0),.din(w_dff_A_I74EMTpF6_0),.clk(gclk));
	jdff dff_A_Cf6IPG4M3_0(.dout(w_dff_A_pY6MpF7n5_0),.din(w_dff_A_Cf6IPG4M3_0),.clk(gclk));
	jdff dff_A_pY6MpF7n5_0(.dout(w_dff_A_vYfE49QH5_0),.din(w_dff_A_pY6MpF7n5_0),.clk(gclk));
	jdff dff_A_vYfE49QH5_0(.dout(w_dff_A_feGpzxdt6_0),.din(w_dff_A_vYfE49QH5_0),.clk(gclk));
	jdff dff_A_feGpzxdt6_0(.dout(w_dff_A_8TcsxdWB7_0),.din(w_dff_A_feGpzxdt6_0),.clk(gclk));
	jdff dff_A_8TcsxdWB7_0(.dout(w_dff_A_GOlA94eU7_0),.din(w_dff_A_8TcsxdWB7_0),.clk(gclk));
	jdff dff_A_GOlA94eU7_0(.dout(w_dff_A_vWC0rTMe7_0),.din(w_dff_A_GOlA94eU7_0),.clk(gclk));
	jdff dff_A_vWC0rTMe7_0(.dout(w_dff_A_U6oIQtNI3_0),.din(w_dff_A_vWC0rTMe7_0),.clk(gclk));
	jdff dff_A_U6oIQtNI3_0(.dout(w_dff_A_l9eJBuwm9_0),.din(w_dff_A_U6oIQtNI3_0),.clk(gclk));
	jdff dff_A_l9eJBuwm9_0(.dout(w_dff_A_9M2BkVY72_0),.din(w_dff_A_l9eJBuwm9_0),.clk(gclk));
	jdff dff_A_9M2BkVY72_0(.dout(w_dff_A_zKbseXdY1_0),.din(w_dff_A_9M2BkVY72_0),.clk(gclk));
	jdff dff_A_zKbseXdY1_0(.dout(w_dff_A_uxJcFMq33_0),.din(w_dff_A_zKbseXdY1_0),.clk(gclk));
	jdff dff_A_uxJcFMq33_0(.dout(w_dff_A_Ms3374Ws4_0),.din(w_dff_A_uxJcFMq33_0),.clk(gclk));
	jdff dff_A_Ms3374Ws4_0(.dout(w_dff_A_A4lppiT41_0),.din(w_dff_A_Ms3374Ws4_0),.clk(gclk));
	jdff dff_A_A4lppiT41_0(.dout(w_dff_A_2C9hefZm2_0),.din(w_dff_A_A4lppiT41_0),.clk(gclk));
	jdff dff_A_2C9hefZm2_0(.dout(w_dff_A_8ys43FSg0_0),.din(w_dff_A_2C9hefZm2_0),.clk(gclk));
	jdff dff_A_8ys43FSg0_0(.dout(w_dff_A_X3V7BDyI1_0),.din(w_dff_A_8ys43FSg0_0),.clk(gclk));
	jdff dff_A_X3V7BDyI1_0(.dout(G397),.din(w_dff_A_X3V7BDyI1_0),.clk(gclk));
	jdff dff_A_HM031umB3_2(.dout(w_dff_A_d0l0xFV00_0),.din(w_dff_A_HM031umB3_2),.clk(gclk));
	jdff dff_A_d0l0xFV00_0(.dout(w_dff_A_0KKg9AiX0_0),.din(w_dff_A_d0l0xFV00_0),.clk(gclk));
	jdff dff_A_0KKg9AiX0_0(.dout(w_dff_A_EkGfxABn4_0),.din(w_dff_A_0KKg9AiX0_0),.clk(gclk));
	jdff dff_A_EkGfxABn4_0(.dout(w_dff_A_uJ6MDq2z2_0),.din(w_dff_A_EkGfxABn4_0),.clk(gclk));
	jdff dff_A_uJ6MDq2z2_0(.dout(w_dff_A_m3TIo9fU3_0),.din(w_dff_A_uJ6MDq2z2_0),.clk(gclk));
	jdff dff_A_m3TIo9fU3_0(.dout(w_dff_A_NSHg86dI9_0),.din(w_dff_A_m3TIo9fU3_0),.clk(gclk));
	jdff dff_A_NSHg86dI9_0(.dout(w_dff_A_7CHquQjY2_0),.din(w_dff_A_NSHg86dI9_0),.clk(gclk));
	jdff dff_A_7CHquQjY2_0(.dout(w_dff_A_InK39cDJ2_0),.din(w_dff_A_7CHquQjY2_0),.clk(gclk));
	jdff dff_A_InK39cDJ2_0(.dout(w_dff_A_gp7jE4gq9_0),.din(w_dff_A_InK39cDJ2_0),.clk(gclk));
	jdff dff_A_gp7jE4gq9_0(.dout(w_dff_A_Mzlw1Mw87_0),.din(w_dff_A_gp7jE4gq9_0),.clk(gclk));
	jdff dff_A_Mzlw1Mw87_0(.dout(w_dff_A_wy3cn1jy8_0),.din(w_dff_A_Mzlw1Mw87_0),.clk(gclk));
	jdff dff_A_wy3cn1jy8_0(.dout(w_dff_A_jC9Luir46_0),.din(w_dff_A_wy3cn1jy8_0),.clk(gclk));
	jdff dff_A_jC9Luir46_0(.dout(G376),.din(w_dff_A_jC9Luir46_0),.clk(gclk));
	jdff dff_A_8OItUSdo4_2(.dout(w_dff_A_3puuAy3g7_0),.din(w_dff_A_8OItUSdo4_2),.clk(gclk));
	jdff dff_A_3puuAy3g7_0(.dout(w_dff_A_4BsxKgGG7_0),.din(w_dff_A_3puuAy3g7_0),.clk(gclk));
	jdff dff_A_4BsxKgGG7_0(.dout(w_dff_A_JwQwdRJd9_0),.din(w_dff_A_4BsxKgGG7_0),.clk(gclk));
	jdff dff_A_JwQwdRJd9_0(.dout(w_dff_A_6IjPNA3O8_0),.din(w_dff_A_JwQwdRJd9_0),.clk(gclk));
	jdff dff_A_6IjPNA3O8_0(.dout(w_dff_A_iiXZWytQ1_0),.din(w_dff_A_6IjPNA3O8_0),.clk(gclk));
	jdff dff_A_iiXZWytQ1_0(.dout(w_dff_A_5hYABx7c3_0),.din(w_dff_A_iiXZWytQ1_0),.clk(gclk));
	jdff dff_A_5hYABx7c3_0(.dout(w_dff_A_vYwIJLai4_0),.din(w_dff_A_5hYABx7c3_0),.clk(gclk));
	jdff dff_A_vYwIJLai4_0(.dout(w_dff_A_3W1KTZyC1_0),.din(w_dff_A_vYwIJLai4_0),.clk(gclk));
	jdff dff_A_3W1KTZyC1_0(.dout(w_dff_A_lXjAEmul2_0),.din(w_dff_A_3W1KTZyC1_0),.clk(gclk));
	jdff dff_A_lXjAEmul2_0(.dout(w_dff_A_CqmAF5Af3_0),.din(w_dff_A_lXjAEmul2_0),.clk(gclk));
	jdff dff_A_CqmAF5Af3_0(.dout(w_dff_A_v4aVc9Fu2_0),.din(w_dff_A_CqmAF5Af3_0),.clk(gclk));
	jdff dff_A_v4aVc9Fu2_0(.dout(w_dff_A_cIDyJVvq4_0),.din(w_dff_A_v4aVc9Fu2_0),.clk(gclk));
	jdff dff_A_cIDyJVvq4_0(.dout(w_dff_A_bLSFTOs08_0),.din(w_dff_A_cIDyJVvq4_0),.clk(gclk));
	jdff dff_A_bLSFTOs08_0(.dout(G379),.din(w_dff_A_bLSFTOs08_0),.clk(gclk));
	jdff dff_A_inYkeue56_2(.dout(w_dff_A_2QOm5tTa3_0),.din(w_dff_A_inYkeue56_2),.clk(gclk));
	jdff dff_A_2QOm5tTa3_0(.dout(w_dff_A_kkFX7zbn4_0),.din(w_dff_A_2QOm5tTa3_0),.clk(gclk));
	jdff dff_A_kkFX7zbn4_0(.dout(w_dff_A_n1DQ6Hyo9_0),.din(w_dff_A_kkFX7zbn4_0),.clk(gclk));
	jdff dff_A_n1DQ6Hyo9_0(.dout(w_dff_A_lePGEnyB7_0),.din(w_dff_A_n1DQ6Hyo9_0),.clk(gclk));
	jdff dff_A_lePGEnyB7_0(.dout(w_dff_A_UYlZJ24e4_0),.din(w_dff_A_lePGEnyB7_0),.clk(gclk));
	jdff dff_A_UYlZJ24e4_0(.dout(w_dff_A_1gygvsue4_0),.din(w_dff_A_UYlZJ24e4_0),.clk(gclk));
	jdff dff_A_1gygvsue4_0(.dout(w_dff_A_7ksOeu1C5_0),.din(w_dff_A_1gygvsue4_0),.clk(gclk));
	jdff dff_A_7ksOeu1C5_0(.dout(w_dff_A_ZpcKkR5f0_0),.din(w_dff_A_7ksOeu1C5_0),.clk(gclk));
	jdff dff_A_ZpcKkR5f0_0(.dout(w_dff_A_MUP3aR5S5_0),.din(w_dff_A_ZpcKkR5f0_0),.clk(gclk));
	jdff dff_A_MUP3aR5S5_0(.dout(w_dff_A_ail1nSTa5_0),.din(w_dff_A_MUP3aR5S5_0),.clk(gclk));
	jdff dff_A_ail1nSTa5_0(.dout(w_dff_A_KW6wmjNm7_0),.din(w_dff_A_ail1nSTa5_0),.clk(gclk));
	jdff dff_A_KW6wmjNm7_0(.dout(w_dff_A_mZxXFjU60_0),.din(w_dff_A_KW6wmjNm7_0),.clk(gclk));
	jdff dff_A_mZxXFjU60_0(.dout(w_dff_A_zpQ5j4nn3_0),.din(w_dff_A_mZxXFjU60_0),.clk(gclk));
	jdff dff_A_zpQ5j4nn3_0(.dout(G382),.din(w_dff_A_zpQ5j4nn3_0),.clk(gclk));
	jdff dff_A_YuMbcDwy0_2(.dout(w_dff_A_zW47M1Cl9_0),.din(w_dff_A_YuMbcDwy0_2),.clk(gclk));
	jdff dff_A_zW47M1Cl9_0(.dout(w_dff_A_9TFxO4n12_0),.din(w_dff_A_zW47M1Cl9_0),.clk(gclk));
	jdff dff_A_9TFxO4n12_0(.dout(w_dff_A_YHGaE2yP9_0),.din(w_dff_A_9TFxO4n12_0),.clk(gclk));
	jdff dff_A_YHGaE2yP9_0(.dout(w_dff_A_rmSN70mW1_0),.din(w_dff_A_YHGaE2yP9_0),.clk(gclk));
	jdff dff_A_rmSN70mW1_0(.dout(w_dff_A_d4LYHthq4_0),.din(w_dff_A_rmSN70mW1_0),.clk(gclk));
	jdff dff_A_d4LYHthq4_0(.dout(w_dff_A_MGQenSyl3_0),.din(w_dff_A_d4LYHthq4_0),.clk(gclk));
	jdff dff_A_MGQenSyl3_0(.dout(w_dff_A_bp9JPRAO1_0),.din(w_dff_A_MGQenSyl3_0),.clk(gclk));
	jdff dff_A_bp9JPRAO1_0(.dout(w_dff_A_5ebaY0NB4_0),.din(w_dff_A_bp9JPRAO1_0),.clk(gclk));
	jdff dff_A_5ebaY0NB4_0(.dout(w_dff_A_q61o1CA68_0),.din(w_dff_A_5ebaY0NB4_0),.clk(gclk));
	jdff dff_A_q61o1CA68_0(.dout(w_dff_A_9Q0UF8CC5_0),.din(w_dff_A_q61o1CA68_0),.clk(gclk));
	jdff dff_A_9Q0UF8CC5_0(.dout(w_dff_A_iA2GrFun9_0),.din(w_dff_A_9Q0UF8CC5_0),.clk(gclk));
	jdff dff_A_iA2GrFun9_0(.dout(w_dff_A_DiLYexTM8_0),.din(w_dff_A_iA2GrFun9_0),.clk(gclk));
	jdff dff_A_DiLYexTM8_0(.dout(w_dff_A_otGRFl6Z0_0),.din(w_dff_A_DiLYexTM8_0),.clk(gclk));
	jdff dff_A_otGRFl6Z0_0(.dout(w_dff_A_jCr3aH0v0_0),.din(w_dff_A_otGRFl6Z0_0),.clk(gclk));
	jdff dff_A_jCr3aH0v0_0(.dout(w_dff_A_0u8hVAdx7_0),.din(w_dff_A_jCr3aH0v0_0),.clk(gclk));
	jdff dff_A_0u8hVAdx7_0(.dout(G385),.din(w_dff_A_0u8hVAdx7_0),.clk(gclk));
	jdff dff_A_vKTTodl25_1(.dout(w_dff_A_1SNUD7x36_0),.din(w_dff_A_vKTTodl25_1),.clk(gclk));
	jdff dff_A_1SNUD7x36_0(.dout(w_dff_A_6PtWGPY90_0),.din(w_dff_A_1SNUD7x36_0),.clk(gclk));
	jdff dff_A_6PtWGPY90_0(.dout(w_dff_A_lQ4MsByd2_0),.din(w_dff_A_6PtWGPY90_0),.clk(gclk));
	jdff dff_A_lQ4MsByd2_0(.dout(w_dff_A_UMCOfAL28_0),.din(w_dff_A_lQ4MsByd2_0),.clk(gclk));
	jdff dff_A_UMCOfAL28_0(.dout(w_dff_A_1gS5BeSi5_0),.din(w_dff_A_UMCOfAL28_0),.clk(gclk));
	jdff dff_A_1gS5BeSi5_0(.dout(w_dff_A_dFYhTuT95_0),.din(w_dff_A_1gS5BeSi5_0),.clk(gclk));
	jdff dff_A_dFYhTuT95_0(.dout(w_dff_A_Vo3arQaY1_0),.din(w_dff_A_dFYhTuT95_0),.clk(gclk));
	jdff dff_A_Vo3arQaY1_0(.dout(w_dff_A_Qyma0x8A6_0),.din(w_dff_A_Vo3arQaY1_0),.clk(gclk));
	jdff dff_A_Qyma0x8A6_0(.dout(w_dff_A_5pnbjrPM1_0),.din(w_dff_A_Qyma0x8A6_0),.clk(gclk));
	jdff dff_A_5pnbjrPM1_0(.dout(w_dff_A_eYGLvuyF7_0),.din(w_dff_A_5pnbjrPM1_0),.clk(gclk));
	jdff dff_A_eYGLvuyF7_0(.dout(w_dff_A_nTsDorUF7_0),.din(w_dff_A_eYGLvuyF7_0),.clk(gclk));
	jdff dff_A_nTsDorUF7_0(.dout(w_dff_A_IncAMnTY7_0),.din(w_dff_A_nTsDorUF7_0),.clk(gclk));
	jdff dff_A_IncAMnTY7_0(.dout(w_dff_A_XhGGlwzN4_0),.din(w_dff_A_IncAMnTY7_0),.clk(gclk));
	jdff dff_A_XhGGlwzN4_0(.dout(w_dff_A_xnA5D6Te8_0),.din(w_dff_A_XhGGlwzN4_0),.clk(gclk));
	jdff dff_A_xnA5D6Te8_0(.dout(w_dff_A_wSfUCgex2_0),.din(w_dff_A_xnA5D6Te8_0),.clk(gclk));
	jdff dff_A_wSfUCgex2_0(.dout(G412),.din(w_dff_A_wSfUCgex2_0),.clk(gclk));
	jdff dff_A_09UngzC83_1(.dout(w_dff_A_lbqh8aXs4_0),.din(w_dff_A_09UngzC83_1),.clk(gclk));
	jdff dff_A_lbqh8aXs4_0(.dout(w_dff_A_Ii9eUP6J9_0),.din(w_dff_A_lbqh8aXs4_0),.clk(gclk));
	jdff dff_A_Ii9eUP6J9_0(.dout(w_dff_A_VT96i3Eu1_0),.din(w_dff_A_Ii9eUP6J9_0),.clk(gclk));
	jdff dff_A_VT96i3Eu1_0(.dout(w_dff_A_bgmwtF6n8_0),.din(w_dff_A_VT96i3Eu1_0),.clk(gclk));
	jdff dff_A_bgmwtF6n8_0(.dout(w_dff_A_YUXqakBE9_0),.din(w_dff_A_bgmwtF6n8_0),.clk(gclk));
	jdff dff_A_YUXqakBE9_0(.dout(w_dff_A_RsgyrWvQ6_0),.din(w_dff_A_YUXqakBE9_0),.clk(gclk));
	jdff dff_A_RsgyrWvQ6_0(.dout(w_dff_A_jS8xAlv22_0),.din(w_dff_A_RsgyrWvQ6_0),.clk(gclk));
	jdff dff_A_jS8xAlv22_0(.dout(w_dff_A_ib4bd8ej0_0),.din(w_dff_A_jS8xAlv22_0),.clk(gclk));
	jdff dff_A_ib4bd8ej0_0(.dout(w_dff_A_YJtMS9783_0),.din(w_dff_A_ib4bd8ej0_0),.clk(gclk));
	jdff dff_A_YJtMS9783_0(.dout(w_dff_A_6dxDDTUe7_0),.din(w_dff_A_YJtMS9783_0),.clk(gclk));
	jdff dff_A_6dxDDTUe7_0(.dout(w_dff_A_zhIstHAG6_0),.din(w_dff_A_6dxDDTUe7_0),.clk(gclk));
	jdff dff_A_zhIstHAG6_0(.dout(w_dff_A_E5az9PlC2_0),.din(w_dff_A_zhIstHAG6_0),.clk(gclk));
	jdff dff_A_E5az9PlC2_0(.dout(w_dff_A_9NdZmENl4_0),.din(w_dff_A_E5az9PlC2_0),.clk(gclk));
	jdff dff_A_9NdZmENl4_0(.dout(w_dff_A_csKpx9Jp4_0),.din(w_dff_A_9NdZmENl4_0),.clk(gclk));
	jdff dff_A_csKpx9Jp4_0(.dout(w_dff_A_qQQyCCo16_0),.din(w_dff_A_csKpx9Jp4_0),.clk(gclk));
	jdff dff_A_qQQyCCo16_0(.dout(G414),.din(w_dff_A_qQQyCCo16_0),.clk(gclk));
	jdff dff_A_43cNgcPY5_1(.dout(w_dff_A_YuP3xOfQ8_0),.din(w_dff_A_43cNgcPY5_1),.clk(gclk));
	jdff dff_A_YuP3xOfQ8_0(.dout(w_dff_A_5OBjewN68_0),.din(w_dff_A_YuP3xOfQ8_0),.clk(gclk));
	jdff dff_A_5OBjewN68_0(.dout(w_dff_A_NG6SqmY73_0),.din(w_dff_A_5OBjewN68_0),.clk(gclk));
	jdff dff_A_NG6SqmY73_0(.dout(w_dff_A_MwFGg6kr2_0),.din(w_dff_A_NG6SqmY73_0),.clk(gclk));
	jdff dff_A_MwFGg6kr2_0(.dout(w_dff_A_c06rjhzr0_0),.din(w_dff_A_MwFGg6kr2_0),.clk(gclk));
	jdff dff_A_c06rjhzr0_0(.dout(w_dff_A_cpUVx2x90_0),.din(w_dff_A_c06rjhzr0_0),.clk(gclk));
	jdff dff_A_cpUVx2x90_0(.dout(w_dff_A_G6h6vG254_0),.din(w_dff_A_cpUVx2x90_0),.clk(gclk));
	jdff dff_A_G6h6vG254_0(.dout(w_dff_A_iDdVmCoa8_0),.din(w_dff_A_G6h6vG254_0),.clk(gclk));
	jdff dff_A_iDdVmCoa8_0(.dout(w_dff_A_vvPkSMG95_0),.din(w_dff_A_iDdVmCoa8_0),.clk(gclk));
	jdff dff_A_vvPkSMG95_0(.dout(w_dff_A_IES5gsep5_0),.din(w_dff_A_vvPkSMG95_0),.clk(gclk));
	jdff dff_A_IES5gsep5_0(.dout(w_dff_A_v6PjrZEA2_0),.din(w_dff_A_IES5gsep5_0),.clk(gclk));
	jdff dff_A_v6PjrZEA2_0(.dout(w_dff_A_GBKT7SiV3_0),.din(w_dff_A_v6PjrZEA2_0),.clk(gclk));
	jdff dff_A_GBKT7SiV3_0(.dout(w_dff_A_bemAgK2w3_0),.din(w_dff_A_GBKT7SiV3_0),.clk(gclk));
	jdff dff_A_bemAgK2w3_0(.dout(G416),.din(w_dff_A_bemAgK2w3_0),.clk(gclk));
	jdff dff_A_tocXicLV2_2(.dout(w_dff_A_WDr71kD12_0),.din(w_dff_A_tocXicLV2_2),.clk(gclk));
	jdff dff_A_WDr71kD12_0(.dout(w_dff_A_9v82n2yI3_0),.din(w_dff_A_WDr71kD12_0),.clk(gclk));
	jdff dff_A_9v82n2yI3_0(.dout(w_dff_A_oXJ2JL4K5_0),.din(w_dff_A_9v82n2yI3_0),.clk(gclk));
	jdff dff_A_oXJ2JL4K5_0(.dout(w_dff_A_nLZZwu0d9_0),.din(w_dff_A_oXJ2JL4K5_0),.clk(gclk));
	jdff dff_A_nLZZwu0d9_0(.dout(w_dff_A_KEUS3aF96_0),.din(w_dff_A_nLZZwu0d9_0),.clk(gclk));
	jdff dff_A_KEUS3aF96_0(.dout(w_dff_A_bwK6dfun3_0),.din(w_dff_A_KEUS3aF96_0),.clk(gclk));
	jdff dff_A_bwK6dfun3_0(.dout(G249),.din(w_dff_A_bwK6dfun3_0),.clk(gclk));
	jdff dff_A_R2mLLwKi2_2(.dout(w_dff_A_S2pIv6CO0_0),.din(w_dff_A_R2mLLwKi2_2),.clk(gclk));
	jdff dff_A_S2pIv6CO0_0(.dout(w_dff_A_42pMZg4T4_0),.din(w_dff_A_S2pIv6CO0_0),.clk(gclk));
	jdff dff_A_42pMZg4T4_0(.dout(w_dff_A_NgHBOebl6_0),.din(w_dff_A_42pMZg4T4_0),.clk(gclk));
	jdff dff_A_NgHBOebl6_0(.dout(w_dff_A_tUH3328i7_0),.din(w_dff_A_NgHBOebl6_0),.clk(gclk));
	jdff dff_A_tUH3328i7_0(.dout(w_dff_A_OIzph72k1_0),.din(w_dff_A_tUH3328i7_0),.clk(gclk));
	jdff dff_A_OIzph72k1_0(.dout(w_dff_A_EnKcLzSO6_0),.din(w_dff_A_OIzph72k1_0),.clk(gclk));
	jdff dff_A_EnKcLzSO6_0(.dout(w_dff_A_hhUqR0WX6_0),.din(w_dff_A_EnKcLzSO6_0),.clk(gclk));
	jdff dff_A_hhUqR0WX6_0(.dout(w_dff_A_ehmDPqH06_0),.din(w_dff_A_hhUqR0WX6_0),.clk(gclk));
	jdff dff_A_ehmDPqH06_0(.dout(w_dff_A_sDXAHvYj2_0),.din(w_dff_A_ehmDPqH06_0),.clk(gclk));
	jdff dff_A_sDXAHvYj2_0(.dout(G295),.din(w_dff_A_sDXAHvYj2_0),.clk(gclk));
	jdff dff_A_kWtpVriV9_2(.dout(w_dff_A_LwuAuHUQ8_0),.din(w_dff_A_kWtpVriV9_2),.clk(gclk));
	jdff dff_A_LwuAuHUQ8_0(.dout(w_dff_A_uNXpyo9T9_0),.din(w_dff_A_LwuAuHUQ8_0),.clk(gclk));
	jdff dff_A_uNXpyo9T9_0(.dout(w_dff_A_PNdJsUEN7_0),.din(w_dff_A_uNXpyo9T9_0),.clk(gclk));
	jdff dff_A_PNdJsUEN7_0(.dout(w_dff_A_WZE92r3R6_0),.din(w_dff_A_PNdJsUEN7_0),.clk(gclk));
	jdff dff_A_WZE92r3R6_0(.dout(w_dff_A_tWIqak8g0_0),.din(w_dff_A_WZE92r3R6_0),.clk(gclk));
	jdff dff_A_tWIqak8g0_0(.dout(G324),.din(w_dff_A_tWIqak8g0_0),.clk(gclk));
	jdff dff_A_jUZ9oWmy2_2(.dout(w_dff_A_7lBMX5AL7_0),.din(w_dff_A_jUZ9oWmy2_2),.clk(gclk));
	jdff dff_A_7lBMX5AL7_0(.dout(w_dff_A_zh1NqjjA8_0),.din(w_dff_A_7lBMX5AL7_0),.clk(gclk));
	jdff dff_A_zh1NqjjA8_0(.dout(w_dff_A_CaHjyrq47_0),.din(w_dff_A_zh1NqjjA8_0),.clk(gclk));
	jdff dff_A_CaHjyrq47_0(.dout(w_dff_A_uGeCxVnY4_0),.din(w_dff_A_CaHjyrq47_0),.clk(gclk));
	jdff dff_A_uGeCxVnY4_0(.dout(w_dff_A_EBG2ZNh52_0),.din(w_dff_A_uGeCxVnY4_0),.clk(gclk));
	jdff dff_A_EBG2ZNh52_0(.dout(w_dff_A_nlrj6dYC5_0),.din(w_dff_A_EBG2ZNh52_0),.clk(gclk));
	jdff dff_A_nlrj6dYC5_0(.dout(w_dff_A_hQqt921o4_0),.din(w_dff_A_nlrj6dYC5_0),.clk(gclk));
	jdff dff_A_hQqt921o4_0(.dout(w_dff_A_sJgjWK4R2_0),.din(w_dff_A_hQqt921o4_0),.clk(gclk));
	jdff dff_A_sJgjWK4R2_0(.dout(w_dff_A_gJEkRr062_0),.din(w_dff_A_sJgjWK4R2_0),.clk(gclk));
	jdff dff_A_gJEkRr062_0(.dout(G252),.din(w_dff_A_gJEkRr062_0),.clk(gclk));
	jdff dff_A_u65loDku7_2(.dout(G276),.din(w_dff_A_u65loDku7_2),.clk(gclk));
	jdff dff_A_bs3dCZUn0_2(.dout(w_dff_A_d5I7HYBu6_0),.din(w_dff_A_bs3dCZUn0_2),.clk(gclk));
	jdff dff_A_d5I7HYBu6_0(.dout(w_dff_A_UJ8zaBR02_0),.din(w_dff_A_d5I7HYBu6_0),.clk(gclk));
	jdff dff_A_UJ8zaBR02_0(.dout(w_dff_A_rZPzMJ467_0),.din(w_dff_A_UJ8zaBR02_0),.clk(gclk));
	jdff dff_A_rZPzMJ467_0(.dout(w_dff_A_qUejOMLH0_0),.din(w_dff_A_rZPzMJ467_0),.clk(gclk));
	jdff dff_A_qUejOMLH0_0(.dout(w_dff_A_HHjaTWLT9_0),.din(w_dff_A_qUejOMLH0_0),.clk(gclk));
	jdff dff_A_HHjaTWLT9_0(.dout(G310),.din(w_dff_A_HHjaTWLT9_0),.clk(gclk));
	jdff dff_A_amWUnRaU2_2(.dout(w_dff_A_tQHjlOxl1_0),.din(w_dff_A_amWUnRaU2_2),.clk(gclk));
	jdff dff_A_tQHjlOxl1_0(.dout(w_dff_A_5ZJs7CSk4_0),.din(w_dff_A_tQHjlOxl1_0),.clk(gclk));
	jdff dff_A_5ZJs7CSk4_0(.dout(w_dff_A_ilIpNWmd5_0),.din(w_dff_A_5ZJs7CSk4_0),.clk(gclk));
	jdff dff_A_ilIpNWmd5_0(.dout(w_dff_A_7TSTUoMv9_0),.din(w_dff_A_ilIpNWmd5_0),.clk(gclk));
	jdff dff_A_7TSTUoMv9_0(.dout(w_dff_A_UZYjd2Ag6_0),.din(w_dff_A_7TSTUoMv9_0),.clk(gclk));
	jdff dff_A_UZYjd2Ag6_0(.dout(w_dff_A_uq0eShYm4_0),.din(w_dff_A_UZYjd2Ag6_0),.clk(gclk));
	jdff dff_A_uq0eShYm4_0(.dout(G313),.din(w_dff_A_uq0eShYm4_0),.clk(gclk));
	jdff dff_A_hR2WjjY39_2(.dout(w_dff_A_jTTaRbyp0_0),.din(w_dff_A_hR2WjjY39_2),.clk(gclk));
	jdff dff_A_jTTaRbyp0_0(.dout(w_dff_A_4EyhSLwu4_0),.din(w_dff_A_jTTaRbyp0_0),.clk(gclk));
	jdff dff_A_4EyhSLwu4_0(.dout(w_dff_A_KRqJ0BaK6_0),.din(w_dff_A_4EyhSLwu4_0),.clk(gclk));
	jdff dff_A_KRqJ0BaK6_0(.dout(w_dff_A_WDsUy5CT6_0),.din(w_dff_A_KRqJ0BaK6_0),.clk(gclk));
	jdff dff_A_WDsUy5CT6_0(.dout(w_dff_A_9aEZRltC3_0),.din(w_dff_A_WDsUy5CT6_0),.clk(gclk));
	jdff dff_A_9aEZRltC3_0(.dout(w_dff_A_Vtb3DA6f9_0),.din(w_dff_A_9aEZRltC3_0),.clk(gclk));
	jdff dff_A_Vtb3DA6f9_0(.dout(w_dff_A_QTIIJAgD2_0),.din(w_dff_A_Vtb3DA6f9_0),.clk(gclk));
	jdff dff_A_QTIIJAgD2_0(.dout(G316),.din(w_dff_A_QTIIJAgD2_0),.clk(gclk));
	jdff dff_A_DEUGBpxE4_2(.dout(w_dff_A_3LDz5kvJ5_0),.din(w_dff_A_DEUGBpxE4_2),.clk(gclk));
	jdff dff_A_3LDz5kvJ5_0(.dout(w_dff_A_AiWTeekL2_0),.din(w_dff_A_3LDz5kvJ5_0),.clk(gclk));
	jdff dff_A_AiWTeekL2_0(.dout(w_dff_A_Xhs6slgQ5_0),.din(w_dff_A_AiWTeekL2_0),.clk(gclk));
	jdff dff_A_Xhs6slgQ5_0(.dout(w_dff_A_QOxPoQFD5_0),.din(w_dff_A_Xhs6slgQ5_0),.clk(gclk));
	jdff dff_A_QOxPoQFD5_0(.dout(w_dff_A_m7KmafAM5_0),.din(w_dff_A_QOxPoQFD5_0),.clk(gclk));
	jdff dff_A_m7KmafAM5_0(.dout(w_dff_A_Vhi4oWOV7_0),.din(w_dff_A_m7KmafAM5_0),.clk(gclk));
	jdff dff_A_Vhi4oWOV7_0(.dout(w_dff_A_VRC1E4O96_0),.din(w_dff_A_Vhi4oWOV7_0),.clk(gclk));
	jdff dff_A_VRC1E4O96_0(.dout(G319),.din(w_dff_A_VRC1E4O96_0),.clk(gclk));
	jdff dff_A_AdXSab4c0_2(.dout(w_dff_A_N8ez5Be21_0),.din(w_dff_A_AdXSab4c0_2),.clk(gclk));
	jdff dff_A_N8ez5Be21_0(.dout(G327),.din(w_dff_A_N8ez5Be21_0),.clk(gclk));
	jdff dff_A_tDqTzf6y5_2(.dout(w_dff_A_WQJSos3G3_0),.din(w_dff_A_tDqTzf6y5_2),.clk(gclk));
	jdff dff_A_WQJSos3G3_0(.dout(w_dff_A_4zuOeTUn8_0),.din(w_dff_A_WQJSos3G3_0),.clk(gclk));
	jdff dff_A_4zuOeTUn8_0(.dout(G330),.din(w_dff_A_4zuOeTUn8_0),.clk(gclk));
	jdff dff_A_pC7Cjpvr8_2(.dout(w_dff_A_OhDGTutM7_0),.din(w_dff_A_pC7Cjpvr8_2),.clk(gclk));
	jdff dff_A_OhDGTutM7_0(.dout(w_dff_A_UhHQux9E2_0),.din(w_dff_A_OhDGTutM7_0),.clk(gclk));
	jdff dff_A_UhHQux9E2_0(.dout(w_dff_A_UcyusA3V2_0),.din(w_dff_A_UhHQux9E2_0),.clk(gclk));
	jdff dff_A_UcyusA3V2_0(.dout(G333),.din(w_dff_A_UcyusA3V2_0),.clk(gclk));
	jdff dff_A_pWEqVmr15_2(.dout(w_dff_A_5qLxu60L2_0),.din(w_dff_A_pWEqVmr15_2),.clk(gclk));
	jdff dff_A_5qLxu60L2_0(.dout(w_dff_A_US3dwx8F9_0),.din(w_dff_A_5qLxu60L2_0),.clk(gclk));
	jdff dff_A_US3dwx8F9_0(.dout(w_dff_A_8yBKoaa10_0),.din(w_dff_A_US3dwx8F9_0),.clk(gclk));
	jdff dff_A_8yBKoaa10_0(.dout(G336),.din(w_dff_A_8yBKoaa10_0),.clk(gclk));
	jdff dff_A_8GhQPmXM9_2(.dout(w_dff_A_HjdfjwHP0_0),.din(w_dff_A_8GhQPmXM9_2),.clk(gclk));
	jdff dff_A_HjdfjwHP0_0(.dout(w_dff_A_h8NITfi00_0),.din(w_dff_A_HjdfjwHP0_0),.clk(gclk));
	jdff dff_A_h8NITfi00_0(.dout(w_dff_A_pajs5PTE8_0),.din(w_dff_A_h8NITfi00_0),.clk(gclk));
	jdff dff_A_pajs5PTE8_0(.dout(w_dff_A_VtObylxT9_0),.din(w_dff_A_pajs5PTE8_0),.clk(gclk));
	jdff dff_A_VtObylxT9_0(.dout(w_dff_A_AUecmcjN3_0),.din(w_dff_A_VtObylxT9_0),.clk(gclk));
	jdff dff_A_AUecmcjN3_0(.dout(w_dff_A_fFNtUUEv8_0),.din(w_dff_A_AUecmcjN3_0),.clk(gclk));
	jdff dff_A_fFNtUUEv8_0(.dout(w_dff_A_hDPW3WLJ2_0),.din(w_dff_A_fFNtUUEv8_0),.clk(gclk));
	jdff dff_A_hDPW3WLJ2_0(.dout(w_dff_A_9hEZxHmz4_0),.din(w_dff_A_hDPW3WLJ2_0),.clk(gclk));
	jdff dff_A_9hEZxHmz4_0(.dout(w_dff_A_ALaRuceH1_0),.din(w_dff_A_9hEZxHmz4_0),.clk(gclk));
	jdff dff_A_ALaRuceH1_0(.dout(w_dff_A_66IERIMB8_0),.din(w_dff_A_ALaRuceH1_0),.clk(gclk));
	jdff dff_A_66IERIMB8_0(.dout(w_dff_A_cXIGW9EM4_0),.din(w_dff_A_66IERIMB8_0),.clk(gclk));
	jdff dff_A_cXIGW9EM4_0(.dout(G418),.din(w_dff_A_cXIGW9EM4_0),.clk(gclk));
	jdff dff_A_rnuc3wek8_2(.dout(G273),.din(w_dff_A_rnuc3wek8_2),.clk(gclk));
	jdff dff_A_BfQSCrDb1_2(.dout(w_dff_A_egvpQFI02_0),.din(w_dff_A_BfQSCrDb1_2),.clk(gclk));
	jdff dff_A_egvpQFI02_0(.dout(w_dff_A_5p4R2p4r9_0),.din(w_dff_A_egvpQFI02_0),.clk(gclk));
	jdff dff_A_5p4R2p4r9_0(.dout(w_dff_A_bVZdos4u9_0),.din(w_dff_A_5p4R2p4r9_0),.clk(gclk));
	jdff dff_A_bVZdos4u9_0(.dout(G298),.din(w_dff_A_bVZdos4u9_0),.clk(gclk));
	jdff dff_A_LvjRIxn72_2(.dout(w_dff_A_03OrYuA79_0),.din(w_dff_A_LvjRIxn72_2),.clk(gclk));
	jdff dff_A_03OrYuA79_0(.dout(w_dff_A_kt4TUV400_0),.din(w_dff_A_03OrYuA79_0),.clk(gclk));
	jdff dff_A_kt4TUV400_0(.dout(w_dff_A_yPsxLdux3_0),.din(w_dff_A_kt4TUV400_0),.clk(gclk));
	jdff dff_A_yPsxLdux3_0(.dout(w_dff_A_FCyRsOtw1_0),.din(w_dff_A_yPsxLdux3_0),.clk(gclk));
	jdff dff_A_FCyRsOtw1_0(.dout(w_dff_A_kiqIxzv19_0),.din(w_dff_A_FCyRsOtw1_0),.clk(gclk));
	jdff dff_A_kiqIxzv19_0(.dout(G301),.din(w_dff_A_kiqIxzv19_0),.clk(gclk));
	jdff dff_A_9o2BrKL15_2(.dout(w_dff_A_IT05QvZ51_0),.din(w_dff_A_9o2BrKL15_2),.clk(gclk));
	jdff dff_A_IT05QvZ51_0(.dout(w_dff_A_Jw8QBLpY4_0),.din(w_dff_A_IT05QvZ51_0),.clk(gclk));
	jdff dff_A_Jw8QBLpY4_0(.dout(w_dff_A_OHU5xNHF9_0),.din(w_dff_A_Jw8QBLpY4_0),.clk(gclk));
	jdff dff_A_OHU5xNHF9_0(.dout(w_dff_A_l9zrvFcK4_0),.din(w_dff_A_OHU5xNHF9_0),.clk(gclk));
	jdff dff_A_l9zrvFcK4_0(.dout(w_dff_A_3sHBIowx4_0),.din(w_dff_A_l9zrvFcK4_0),.clk(gclk));
	jdff dff_A_3sHBIowx4_0(.dout(G304),.din(w_dff_A_3sHBIowx4_0),.clk(gclk));
	jdff dff_A_TB6D4vo83_2(.dout(w_dff_A_kzXUpVAQ3_0),.din(w_dff_A_TB6D4vo83_2),.clk(gclk));
	jdff dff_A_kzXUpVAQ3_0(.dout(w_dff_A_yrSKSwGe6_0),.din(w_dff_A_kzXUpVAQ3_0),.clk(gclk));
	jdff dff_A_yrSKSwGe6_0(.dout(w_dff_A_UnIAgsPA8_0),.din(w_dff_A_yrSKSwGe6_0),.clk(gclk));
	jdff dff_A_UnIAgsPA8_0(.dout(w_dff_A_8I6MWYIg6_0),.din(w_dff_A_UnIAgsPA8_0),.clk(gclk));
	jdff dff_A_8I6MWYIg6_0(.dout(w_dff_A_epUeQGpD1_0),.din(w_dff_A_8I6MWYIg6_0),.clk(gclk));
	jdff dff_A_epUeQGpD1_0(.dout(w_dff_A_MQg6KNYn1_0),.din(w_dff_A_epUeQGpD1_0),.clk(gclk));
	jdff dff_A_MQg6KNYn1_0(.dout(w_dff_A_TJuwzeWO2_0),.din(w_dff_A_MQg6KNYn1_0),.clk(gclk));
	jdff dff_A_TJuwzeWO2_0(.dout(G307),.din(w_dff_A_TJuwzeWO2_0),.clk(gclk));
	jdff dff_A_VdTQjnjS5_2(.dout(w_dff_A_WiKhgYf83_0),.din(w_dff_A_VdTQjnjS5_2),.clk(gclk));
	jdff dff_A_WiKhgYf83_0(.dout(w_dff_A_KgwgZIgZ2_0),.din(w_dff_A_WiKhgYf83_0),.clk(gclk));
	jdff dff_A_KgwgZIgZ2_0(.dout(w_dff_A_QXo3CoVZ5_0),.din(w_dff_A_KgwgZIgZ2_0),.clk(gclk));
	jdff dff_A_QXo3CoVZ5_0(.dout(w_dff_A_GBgOnyp30_0),.din(w_dff_A_QXo3CoVZ5_0),.clk(gclk));
	jdff dff_A_GBgOnyp30_0(.dout(w_dff_A_NZOmZO4Y7_0),.din(w_dff_A_GBgOnyp30_0),.clk(gclk));
	jdff dff_A_NZOmZO4Y7_0(.dout(w_dff_A_Qb6tYkXv7_0),.din(w_dff_A_NZOmZO4Y7_0),.clk(gclk));
	jdff dff_A_Qb6tYkXv7_0(.dout(w_dff_A_750Ii5E99_0),.din(w_dff_A_Qb6tYkXv7_0),.clk(gclk));
	jdff dff_A_750Ii5E99_0(.dout(w_dff_A_Wcbiwsft1_0),.din(w_dff_A_750Ii5E99_0),.clk(gclk));
	jdff dff_A_Wcbiwsft1_0(.dout(w_dff_A_Q1XuOow32_0),.din(w_dff_A_Wcbiwsft1_0),.clk(gclk));
	jdff dff_A_Q1XuOow32_0(.dout(w_dff_A_fScZqcuv5_0),.din(w_dff_A_Q1XuOow32_0),.clk(gclk));
	jdff dff_A_fScZqcuv5_0(.dout(w_dff_A_QmWurOe12_0),.din(w_dff_A_fScZqcuv5_0),.clk(gclk));
	jdff dff_A_QmWurOe12_0(.dout(w_dff_A_BCSA4pmd6_0),.din(w_dff_A_QmWurOe12_0),.clk(gclk));
	jdff dff_A_BCSA4pmd6_0(.dout(w_dff_A_psZAIvTZ2_0),.din(w_dff_A_BCSA4pmd6_0),.clk(gclk));
	jdff dff_A_psZAIvTZ2_0(.dout(G344),.din(w_dff_A_psZAIvTZ2_0),.clk(gclk));
	jdff dff_A_m62Wobqa2_2(.dout(G422),.din(w_dff_A_m62Wobqa2_2),.clk(gclk));
	jdff dff_A_FCyTexHS6_2(.dout(G469),.din(w_dff_A_FCyTexHS6_2),.clk(gclk));
	jdff dff_A_WnsCWwMe4_2(.dout(w_dff_A_McKfIN4R6_0),.din(w_dff_A_WnsCWwMe4_2),.clk(gclk));
	jdff dff_A_McKfIN4R6_0(.dout(w_dff_A_oUNzt51x0_0),.din(w_dff_A_McKfIN4R6_0),.clk(gclk));
	jdff dff_A_oUNzt51x0_0(.dout(w_dff_A_n9EzxzAo3_0),.din(w_dff_A_oUNzt51x0_0),.clk(gclk));
	jdff dff_A_n9EzxzAo3_0(.dout(G419),.din(w_dff_A_n9EzxzAo3_0),.clk(gclk));
	jdff dff_A_uZI5p8W54_2(.dout(w_dff_A_iIojHEYs1_0),.din(w_dff_A_uZI5p8W54_2),.clk(gclk));
	jdff dff_A_iIojHEYs1_0(.dout(w_dff_A_PRcRXwuq3_0),.din(w_dff_A_iIojHEYs1_0),.clk(gclk));
	jdff dff_A_PRcRXwuq3_0(.dout(w_dff_A_uw64MFh48_0),.din(w_dff_A_PRcRXwuq3_0),.clk(gclk));
	jdff dff_A_uw64MFh48_0(.dout(G471),.din(w_dff_A_uw64MFh48_0),.clk(gclk));
	jdff dff_A_I98csHOR7_2(.dout(w_dff_A_6N3kyfxF4_0),.din(w_dff_A_I98csHOR7_2),.clk(gclk));
	jdff dff_A_6N3kyfxF4_0(.dout(w_dff_A_sKhdD7Wt2_0),.din(w_dff_A_6N3kyfxF4_0),.clk(gclk));
	jdff dff_A_sKhdD7Wt2_0(.dout(w_dff_A_zJXQwMGB2_0),.din(w_dff_A_sKhdD7Wt2_0),.clk(gclk));
	jdff dff_A_zJXQwMGB2_0(.dout(w_dff_A_VLNjR7jZ4_0),.din(w_dff_A_zJXQwMGB2_0),.clk(gclk));
	jdff dff_A_VLNjR7jZ4_0(.dout(w_dff_A_hGJOsO0k5_0),.din(w_dff_A_VLNjR7jZ4_0),.clk(gclk));
	jdff dff_A_hGJOsO0k5_0(.dout(w_dff_A_haoo7cx71_0),.din(w_dff_A_hGJOsO0k5_0),.clk(gclk));
	jdff dff_A_haoo7cx71_0(.dout(w_dff_A_5ZluDnGQ9_0),.din(w_dff_A_haoo7cx71_0),.clk(gclk));
	jdff dff_A_5ZluDnGQ9_0(.dout(w_dff_A_dIxTTPXT3_0),.din(w_dff_A_5ZluDnGQ9_0),.clk(gclk));
	jdff dff_A_dIxTTPXT3_0(.dout(w_dff_A_1qrQnMpl8_0),.din(w_dff_A_dIxTTPXT3_0),.clk(gclk));
	jdff dff_A_1qrQnMpl8_0(.dout(G359),.din(w_dff_A_1qrQnMpl8_0),.clk(gclk));
	jdff dff_A_4R0St17A7_2(.dout(w_dff_A_zsKJpD2c6_0),.din(w_dff_A_4R0St17A7_2),.clk(gclk));
	jdff dff_A_zsKJpD2c6_0(.dout(w_dff_A_35N0Fvqu8_0),.din(w_dff_A_zsKJpD2c6_0),.clk(gclk));
	jdff dff_A_35N0Fvqu8_0(.dout(w_dff_A_BtEK6LCY6_0),.din(w_dff_A_35N0Fvqu8_0),.clk(gclk));
	jdff dff_A_BtEK6LCY6_0(.dout(w_dff_A_ANvtHa8D1_0),.din(w_dff_A_BtEK6LCY6_0),.clk(gclk));
	jdff dff_A_ANvtHa8D1_0(.dout(w_dff_A_1dR5VbvT5_0),.din(w_dff_A_ANvtHa8D1_0),.clk(gclk));
	jdff dff_A_1dR5VbvT5_0(.dout(w_dff_A_elF8ijvU6_0),.din(w_dff_A_1dR5VbvT5_0),.clk(gclk));
	jdff dff_A_elF8ijvU6_0(.dout(w_dff_A_i7NT7RgT4_0),.din(w_dff_A_elF8ijvU6_0),.clk(gclk));
	jdff dff_A_i7NT7RgT4_0(.dout(w_dff_A_oct90Hxu0_0),.din(w_dff_A_i7NT7RgT4_0),.clk(gclk));
	jdff dff_A_oct90Hxu0_0(.dout(w_dff_A_e7pL2a0O3_0),.din(w_dff_A_oct90Hxu0_0),.clk(gclk));
	jdff dff_A_e7pL2a0O3_0(.dout(w_dff_A_skNQEqNp0_0),.din(w_dff_A_e7pL2a0O3_0),.clk(gclk));
	jdff dff_A_skNQEqNp0_0(.dout(G362),.din(w_dff_A_skNQEqNp0_0),.clk(gclk));
	jdff dff_A_y4w19iT65_2(.dout(w_dff_A_mElVkZNX0_0),.din(w_dff_A_y4w19iT65_2),.clk(gclk));
	jdff dff_A_mElVkZNX0_0(.dout(w_dff_A_VayYY6z12_0),.din(w_dff_A_mElVkZNX0_0),.clk(gclk));
	jdff dff_A_VayYY6z12_0(.dout(w_dff_A_AfASEeIM2_0),.din(w_dff_A_VayYY6z12_0),.clk(gclk));
	jdff dff_A_AfASEeIM2_0(.dout(w_dff_A_geMncHqD5_0),.din(w_dff_A_AfASEeIM2_0),.clk(gclk));
	jdff dff_A_geMncHqD5_0(.dout(w_dff_A_46QOf2457_0),.din(w_dff_A_geMncHqD5_0),.clk(gclk));
	jdff dff_A_46QOf2457_0(.dout(w_dff_A_tGjRx1Ix5_0),.din(w_dff_A_46QOf2457_0),.clk(gclk));
	jdff dff_A_tGjRx1Ix5_0(.dout(w_dff_A_b5gUGwaq7_0),.din(w_dff_A_tGjRx1Ix5_0),.clk(gclk));
	jdff dff_A_b5gUGwaq7_0(.dout(w_dff_A_4w5cc3Js4_0),.din(w_dff_A_b5gUGwaq7_0),.clk(gclk));
	jdff dff_A_4w5cc3Js4_0(.dout(w_dff_A_6mjS7akw2_0),.din(w_dff_A_4w5cc3Js4_0),.clk(gclk));
	jdff dff_A_6mjS7akw2_0(.dout(w_dff_A_t7vtsbDg7_0),.din(w_dff_A_6mjS7akw2_0),.clk(gclk));
	jdff dff_A_t7vtsbDg7_0(.dout(w_dff_A_wFzNw0zK1_0),.din(w_dff_A_t7vtsbDg7_0),.clk(gclk));
	jdff dff_A_wFzNw0zK1_0(.dout(G365),.din(w_dff_A_wFzNw0zK1_0),.clk(gclk));
	jdff dff_A_8IAwW4586_2(.dout(w_dff_A_3OD6zrLh5_0),.din(w_dff_A_8IAwW4586_2),.clk(gclk));
	jdff dff_A_3OD6zrLh5_0(.dout(w_dff_A_E8YGGwpI7_0),.din(w_dff_A_3OD6zrLh5_0),.clk(gclk));
	jdff dff_A_E8YGGwpI7_0(.dout(w_dff_A_ZtYm5JhM5_0),.din(w_dff_A_E8YGGwpI7_0),.clk(gclk));
	jdff dff_A_ZtYm5JhM5_0(.dout(w_dff_A_NGbqTv520_0),.din(w_dff_A_ZtYm5JhM5_0),.clk(gclk));
	jdff dff_A_NGbqTv520_0(.dout(w_dff_A_A6SPs8pl3_0),.din(w_dff_A_NGbqTv520_0),.clk(gclk));
	jdff dff_A_A6SPs8pl3_0(.dout(w_dff_A_mklG8sXh5_0),.din(w_dff_A_A6SPs8pl3_0),.clk(gclk));
	jdff dff_A_mklG8sXh5_0(.dout(w_dff_A_j6samyKX8_0),.din(w_dff_A_mklG8sXh5_0),.clk(gclk));
	jdff dff_A_j6samyKX8_0(.dout(w_dff_A_NXvY6m2q2_0),.din(w_dff_A_j6samyKX8_0),.clk(gclk));
	jdff dff_A_NXvY6m2q2_0(.dout(w_dff_A_CKV8gBZk0_0),.din(w_dff_A_NXvY6m2q2_0),.clk(gclk));
	jdff dff_A_CKV8gBZk0_0(.dout(w_dff_A_OVhqUaDg6_0),.din(w_dff_A_CKV8gBZk0_0),.clk(gclk));
	jdff dff_A_OVhqUaDg6_0(.dout(w_dff_A_NKTSE4xa0_0),.din(w_dff_A_OVhqUaDg6_0),.clk(gclk));
	jdff dff_A_NKTSE4xa0_0(.dout(G368),.din(w_dff_A_NKTSE4xa0_0),.clk(gclk));
	jdff dff_A_fT0oI7CZ9_2(.dout(w_dff_A_v6CnyEDK5_0),.din(w_dff_A_fT0oI7CZ9_2),.clk(gclk));
	jdff dff_A_v6CnyEDK5_0(.dout(w_dff_A_9QchQL8X3_0),.din(w_dff_A_v6CnyEDK5_0),.clk(gclk));
	jdff dff_A_9QchQL8X3_0(.dout(w_dff_A_dJ15G3nQ0_0),.din(w_dff_A_9QchQL8X3_0),.clk(gclk));
	jdff dff_A_dJ15G3nQ0_0(.dout(w_dff_A_2ZHnWZN29_0),.din(w_dff_A_dJ15G3nQ0_0),.clk(gclk));
	jdff dff_A_2ZHnWZN29_0(.dout(w_dff_A_FBjujRKJ9_0),.din(w_dff_A_2ZHnWZN29_0),.clk(gclk));
	jdff dff_A_FBjujRKJ9_0(.dout(w_dff_A_Ws2qIQNZ8_0),.din(w_dff_A_FBjujRKJ9_0),.clk(gclk));
	jdff dff_A_Ws2qIQNZ8_0(.dout(w_dff_A_DW6ZtK2o2_0),.din(w_dff_A_Ws2qIQNZ8_0),.clk(gclk));
	jdff dff_A_DW6ZtK2o2_0(.dout(w_dff_A_16NqH9lB9_0),.din(w_dff_A_DW6ZtK2o2_0),.clk(gclk));
	jdff dff_A_16NqH9lB9_0(.dout(G347),.din(w_dff_A_16NqH9lB9_0),.clk(gclk));
	jdff dff_A_aLzr4soI2_2(.dout(w_dff_A_upe8VqZn9_0),.din(w_dff_A_aLzr4soI2_2),.clk(gclk));
	jdff dff_A_upe8VqZn9_0(.dout(w_dff_A_KhCUihHE5_0),.din(w_dff_A_upe8VqZn9_0),.clk(gclk));
	jdff dff_A_KhCUihHE5_0(.dout(w_dff_A_MiSNBpgs1_0),.din(w_dff_A_KhCUihHE5_0),.clk(gclk));
	jdff dff_A_MiSNBpgs1_0(.dout(w_dff_A_TxCmoLst1_0),.din(w_dff_A_MiSNBpgs1_0),.clk(gclk));
	jdff dff_A_TxCmoLst1_0(.dout(w_dff_A_CDWnwMX23_0),.din(w_dff_A_TxCmoLst1_0),.clk(gclk));
	jdff dff_A_CDWnwMX23_0(.dout(w_dff_A_RTY0VLuR8_0),.din(w_dff_A_CDWnwMX23_0),.clk(gclk));
	jdff dff_A_RTY0VLuR8_0(.dout(w_dff_A_BMocbvuz7_0),.din(w_dff_A_RTY0VLuR8_0),.clk(gclk));
	jdff dff_A_BMocbvuz7_0(.dout(w_dff_A_IEHIzVXN2_0),.din(w_dff_A_BMocbvuz7_0),.clk(gclk));
	jdff dff_A_IEHIzVXN2_0(.dout(w_dff_A_HZ5CMwWe8_0),.din(w_dff_A_IEHIzVXN2_0),.clk(gclk));
	jdff dff_A_HZ5CMwWe8_0(.dout(G350),.din(w_dff_A_HZ5CMwWe8_0),.clk(gclk));
	jdff dff_A_cdExsKih7_2(.dout(w_dff_A_lpCLC8Rj2_0),.din(w_dff_A_cdExsKih7_2),.clk(gclk));
	jdff dff_A_lpCLC8Rj2_0(.dout(w_dff_A_NvIaDVch8_0),.din(w_dff_A_lpCLC8Rj2_0),.clk(gclk));
	jdff dff_A_NvIaDVch8_0(.dout(w_dff_A_Rmpyx10o1_0),.din(w_dff_A_NvIaDVch8_0),.clk(gclk));
	jdff dff_A_Rmpyx10o1_0(.dout(w_dff_A_3GZdn6GM6_0),.din(w_dff_A_Rmpyx10o1_0),.clk(gclk));
	jdff dff_A_3GZdn6GM6_0(.dout(w_dff_A_WPUddwiv7_0),.din(w_dff_A_3GZdn6GM6_0),.clk(gclk));
	jdff dff_A_WPUddwiv7_0(.dout(w_dff_A_XXNZpkSH3_0),.din(w_dff_A_WPUddwiv7_0),.clk(gclk));
	jdff dff_A_XXNZpkSH3_0(.dout(w_dff_A_p61JToQo1_0),.din(w_dff_A_XXNZpkSH3_0),.clk(gclk));
	jdff dff_A_p61JToQo1_0(.dout(w_dff_A_TBBlG3BN4_0),.din(w_dff_A_p61JToQo1_0),.clk(gclk));
	jdff dff_A_TBBlG3BN4_0(.dout(w_dff_A_jWnpwcbL9_0),.din(w_dff_A_TBBlG3BN4_0),.clk(gclk));
	jdff dff_A_jWnpwcbL9_0(.dout(G353),.din(w_dff_A_jWnpwcbL9_0),.clk(gclk));
	jdff dff_A_JyIKjTuE8_2(.dout(w_dff_A_btQS2cq52_0),.din(w_dff_A_JyIKjTuE8_2),.clk(gclk));
	jdff dff_A_btQS2cq52_0(.dout(w_dff_A_cR6uF9Sp4_0),.din(w_dff_A_btQS2cq52_0),.clk(gclk));
	jdff dff_A_cR6uF9Sp4_0(.dout(w_dff_A_SYzNlNCk8_0),.din(w_dff_A_cR6uF9Sp4_0),.clk(gclk));
	jdff dff_A_SYzNlNCk8_0(.dout(w_dff_A_5QVUp1sS7_0),.din(w_dff_A_SYzNlNCk8_0),.clk(gclk));
	jdff dff_A_5QVUp1sS7_0(.dout(w_dff_A_nJdlwJI62_0),.din(w_dff_A_5QVUp1sS7_0),.clk(gclk));
	jdff dff_A_nJdlwJI62_0(.dout(w_dff_A_g0MTB0zb6_0),.din(w_dff_A_nJdlwJI62_0),.clk(gclk));
	jdff dff_A_g0MTB0zb6_0(.dout(w_dff_A_TP4r8a0M6_0),.din(w_dff_A_g0MTB0zb6_0),.clk(gclk));
	jdff dff_A_TP4r8a0M6_0(.dout(w_dff_A_DuHT5O0J3_0),.din(w_dff_A_TP4r8a0M6_0),.clk(gclk));
	jdff dff_A_DuHT5O0J3_0(.dout(w_dff_A_eJiXW1rd9_0),.din(w_dff_A_DuHT5O0J3_0),.clk(gclk));
	jdff dff_A_eJiXW1rd9_0(.dout(w_dff_A_G24BZ6301_0),.din(w_dff_A_eJiXW1rd9_0),.clk(gclk));
	jdff dff_A_G24BZ6301_0(.dout(w_dff_A_nn7hbzyR8_0),.din(w_dff_A_G24BZ6301_0),.clk(gclk));
	jdff dff_A_nn7hbzyR8_0(.dout(G356),.din(w_dff_A_nn7hbzyR8_0),.clk(gclk));
	jdff dff_A_3t7SkkRt9_2(.dout(w_dff_A_nyzdXdNn6_0),.din(w_dff_A_3t7SkkRt9_2),.clk(gclk));
	jdff dff_A_nyzdXdNn6_0(.dout(w_dff_A_pvq4Wukz3_0),.din(w_dff_A_nyzdXdNn6_0),.clk(gclk));
	jdff dff_A_pvq4Wukz3_0(.dout(w_dff_A_JNV2UDlX4_0),.din(w_dff_A_pvq4Wukz3_0),.clk(gclk));
	jdff dff_A_JNV2UDlX4_0(.dout(w_dff_A_iYXbgv9d9_0),.din(w_dff_A_JNV2UDlX4_0),.clk(gclk));
	jdff dff_A_iYXbgv9d9_0(.dout(G321),.din(w_dff_A_iYXbgv9d9_0),.clk(gclk));
	jdff dff_A_zYe5zPoI5_2(.dout(w_dff_A_VCfA5K0z6_0),.din(w_dff_A_zYe5zPoI5_2),.clk(gclk));
	jdff dff_A_VCfA5K0z6_0(.dout(w_dff_A_m13q9lbd0_0),.din(w_dff_A_VCfA5K0z6_0),.clk(gclk));
	jdff dff_A_m13q9lbd0_0(.dout(w_dff_A_Xlosk2MW1_0),.din(w_dff_A_m13q9lbd0_0),.clk(gclk));
	jdff dff_A_Xlosk2MW1_0(.dout(w_dff_A_jAs2ksC12_0),.din(w_dff_A_Xlosk2MW1_0),.clk(gclk));
	jdff dff_A_jAs2ksC12_0(.dout(w_dff_A_zEMdixAm4_0),.din(w_dff_A_jAs2ksC12_0),.clk(gclk));
	jdff dff_A_zEMdixAm4_0(.dout(w_dff_A_rLt5lsyh1_0),.din(w_dff_A_zEMdixAm4_0),.clk(gclk));
	jdff dff_A_rLt5lsyh1_0(.dout(G370),.din(w_dff_A_rLt5lsyh1_0),.clk(gclk));
	jdff dff_A_QNml90eu3_2(.dout(w_dff_A_8CmAzMgN4_0),.din(w_dff_A_QNml90eu3_2),.clk(gclk));
	jdff dff_A_8CmAzMgN4_0(.dout(w_dff_A_VP2UI0Kb1_0),.din(w_dff_A_8CmAzMgN4_0),.clk(gclk));
	jdff dff_A_VP2UI0Kb1_0(.dout(w_dff_A_ttHqGC0e8_0),.din(w_dff_A_VP2UI0Kb1_0),.clk(gclk));
	jdff dff_A_ttHqGC0e8_0(.dout(w_dff_A_JI1SDc3z1_0),.din(w_dff_A_ttHqGC0e8_0),.clk(gclk));
	jdff dff_A_JI1SDc3z1_0(.dout(G399),.din(w_dff_A_JI1SDc3z1_0),.clk(gclk));
endmodule

