// Benchmark "top" written by ABC on Thu May 28 22:00:38 2020

module top ( 
    \in0[0] , \in0[1] , \in0[2] , \in0[3] , \in0[4] , \in0[5] , \in0[6] ,
    \in0[7] , \in0[8] , \in0[9] , \in0[10] , \in0[11] , \in0[12] ,
    \in0[13] , \in0[14] , \in0[15] , \in0[16] , \in0[17] , \in0[18] ,
    \in0[19] , \in0[20] , \in0[21] , \in0[22] , \in0[23] , \in0[24] ,
    \in0[25] , \in0[26] , \in0[27] , \in0[28] , \in0[29] , \in0[30] ,
    \in0[31] , \in0[32] , \in0[33] , \in0[34] , \in0[35] , \in0[36] ,
    \in0[37] , \in0[38] , \in0[39] , \in0[40] , \in0[41] , \in0[42] ,
    \in0[43] , \in0[44] , \in0[45] , \in0[46] , \in0[47] , \in0[48] ,
    \in0[49] , \in0[50] , \in0[51] , \in0[52] , \in0[53] , \in0[54] ,
    \in0[55] , \in0[56] , \in0[57] , \in0[58] , \in0[59] , \in0[60] ,
    \in0[61] , \in0[62] , \in0[63] , \in0[64] , \in0[65] , \in0[66] ,
    \in0[67] , \in0[68] , \in0[69] , \in0[70] , \in0[71] , \in0[72] ,
    \in0[73] , \in0[74] , \in0[75] , \in0[76] , \in0[77] , \in0[78] ,
    \in0[79] , \in0[80] , \in0[81] , \in0[82] , \in0[83] , \in0[84] ,
    \in0[85] , \in0[86] , \in0[87] , \in0[88] , \in0[89] , \in0[90] ,
    \in0[91] , \in0[92] , \in0[93] , \in0[94] , \in0[95] , \in0[96] ,
    \in0[97] , \in0[98] , \in0[99] , \in0[100] , \in0[101] , \in0[102] ,
    \in0[103] , \in0[104] , \in0[105] , \in0[106] , \in0[107] , \in0[108] ,
    \in0[109] , \in0[110] , \in0[111] , \in0[112] , \in0[113] , \in0[114] ,
    \in0[115] , \in0[116] , \in0[117] , \in0[118] , \in0[119] , \in0[120] ,
    \in0[121] , \in0[122] , \in0[123] , \in0[124] , \in0[125] , \in0[126] ,
    \in0[127] , \in1[0] , \in1[1] , \in1[2] , \in1[3] , \in1[4] , \in1[5] ,
    \in1[6] , \in1[7] , \in1[8] , \in1[9] , \in1[10] , \in1[11] ,
    \in1[12] , \in1[13] , \in1[14] , \in1[15] , \in1[16] , \in1[17] ,
    \in1[18] , \in1[19] , \in1[20] , \in1[21] , \in1[22] , \in1[23] ,
    \in1[24] , \in1[25] , \in1[26] , \in1[27] , \in1[28] , \in1[29] ,
    \in1[30] , \in1[31] , \in1[32] , \in1[33] , \in1[34] , \in1[35] ,
    \in1[36] , \in1[37] , \in1[38] , \in1[39] , \in1[40] , \in1[41] ,
    \in1[42] , \in1[43] , \in1[44] , \in1[45] , \in1[46] , \in1[47] ,
    \in1[48] , \in1[49] , \in1[50] , \in1[51] , \in1[52] , \in1[53] ,
    \in1[54] , \in1[55] , \in1[56] , \in1[57] , \in1[58] , \in1[59] ,
    \in1[60] , \in1[61] , \in1[62] , \in1[63] , \in1[64] , \in1[65] ,
    \in1[66] , \in1[67] , \in1[68] , \in1[69] , \in1[70] , \in1[71] ,
    \in1[72] , \in1[73] , \in1[74] , \in1[75] , \in1[76] , \in1[77] ,
    \in1[78] , \in1[79] , \in1[80] , \in1[81] , \in1[82] , \in1[83] ,
    \in1[84] , \in1[85] , \in1[86] , \in1[87] , \in1[88] , \in1[89] ,
    \in1[90] , \in1[91] , \in1[92] , \in1[93] , \in1[94] , \in1[95] ,
    \in1[96] , \in1[97] , \in1[98] , \in1[99] , \in1[100] , \in1[101] ,
    \in1[102] , \in1[103] , \in1[104] , \in1[105] , \in1[106] , \in1[107] ,
    \in1[108] , \in1[109] , \in1[110] , \in1[111] , \in1[112] , \in1[113] ,
    \in1[114] , \in1[115] , \in1[116] , \in1[117] , \in1[118] , \in1[119] ,
    \in1[120] , \in1[121] , \in1[122] , \in1[123] , \in1[124] , \in1[125] ,
    \in1[126] , \in1[127] , \in2[0] , \in2[1] , \in2[2] , \in2[3] ,
    \in2[4] , \in2[5] , \in2[6] , \in2[7] , \in2[8] , \in2[9] , \in2[10] ,
    \in2[11] , \in2[12] , \in2[13] , \in2[14] , \in2[15] , \in2[16] ,
    \in2[17] , \in2[18] , \in2[19] , \in2[20] , \in2[21] , \in2[22] ,
    \in2[23] , \in2[24] , \in2[25] , \in2[26] , \in2[27] , \in2[28] ,
    \in2[29] , \in2[30] , \in2[31] , \in2[32] , \in2[33] , \in2[34] ,
    \in2[35] , \in2[36] , \in2[37] , \in2[38] , \in2[39] , \in2[40] ,
    \in2[41] , \in2[42] , \in2[43] , \in2[44] , \in2[45] , \in2[46] ,
    \in2[47] , \in2[48] , \in2[49] , \in2[50] , \in2[51] , \in2[52] ,
    \in2[53] , \in2[54] , \in2[55] , \in2[56] , \in2[57] , \in2[58] ,
    \in2[59] , \in2[60] , \in2[61] , \in2[62] , \in2[63] , \in2[64] ,
    \in2[65] , \in2[66] , \in2[67] , \in2[68] , \in2[69] , \in2[70] ,
    \in2[71] , \in2[72] , \in2[73] , \in2[74] , \in2[75] , \in2[76] ,
    \in2[77] , \in2[78] , \in2[79] , \in2[80] , \in2[81] , \in2[82] ,
    \in2[83] , \in2[84] , \in2[85] , \in2[86] , \in2[87] , \in2[88] ,
    \in2[89] , \in2[90] , \in2[91] , \in2[92] , \in2[93] , \in2[94] ,
    \in2[95] , \in2[96] , \in2[97] , \in2[98] , \in2[99] , \in2[100] ,
    \in2[101] , \in2[102] , \in2[103] , \in2[104] , \in2[105] , \in2[106] ,
    \in2[107] , \in2[108] , \in2[109] , \in2[110] , \in2[111] , \in2[112] ,
    \in2[113] , \in2[114] , \in2[115] , \in2[116] , \in2[117] , \in2[118] ,
    \in2[119] , \in2[120] , \in2[121] , \in2[122] , \in2[123] , \in2[124] ,
    \in2[125] , \in2[126] , \in2[127] , \in3[0] , \in3[1] , \in3[2] ,
    \in3[3] , \in3[4] , \in3[5] , \in3[6] , \in3[7] , \in3[8] , \in3[9] ,
    \in3[10] , \in3[11] , \in3[12] , \in3[13] , \in3[14] , \in3[15] ,
    \in3[16] , \in3[17] , \in3[18] , \in3[19] , \in3[20] , \in3[21] ,
    \in3[22] , \in3[23] , \in3[24] , \in3[25] , \in3[26] , \in3[27] ,
    \in3[28] , \in3[29] , \in3[30] , \in3[31] , \in3[32] , \in3[33] ,
    \in3[34] , \in3[35] , \in3[36] , \in3[37] , \in3[38] , \in3[39] ,
    \in3[40] , \in3[41] , \in3[42] , \in3[43] , \in3[44] , \in3[45] ,
    \in3[46] , \in3[47] , \in3[48] , \in3[49] , \in3[50] , \in3[51] ,
    \in3[52] , \in3[53] , \in3[54] , \in3[55] , \in3[56] , \in3[57] ,
    \in3[58] , \in3[59] , \in3[60] , \in3[61] , \in3[62] , \in3[63] ,
    \in3[64] , \in3[65] , \in3[66] , \in3[67] , \in3[68] , \in3[69] ,
    \in3[70] , \in3[71] , \in3[72] , \in3[73] , \in3[74] , \in3[75] ,
    \in3[76] , \in3[77] , \in3[78] , \in3[79] , \in3[80] , \in3[81] ,
    \in3[82] , \in3[83] , \in3[84] , \in3[85] , \in3[86] , \in3[87] ,
    \in3[88] , \in3[89] , \in3[90] , \in3[91] , \in3[92] , \in3[93] ,
    \in3[94] , \in3[95] , \in3[96] , \in3[97] , \in3[98] , \in3[99] ,
    \in3[100] , \in3[101] , \in3[102] , \in3[103] , \in3[104] , \in3[105] ,
    \in3[106] , \in3[107] , \in3[108] , \in3[109] , \in3[110] , \in3[111] ,
    \in3[112] , \in3[113] , \in3[114] , \in3[115] , \in3[116] , \in3[117] ,
    \in3[118] , \in3[119] , \in3[120] , \in3[121] , \in3[122] , \in3[123] ,
    \in3[124] , \in3[125] , \in3[126] , \in3[127] ,
    \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ,
    \address[0] , \address[1]   );
  input  \in0[0] , \in0[1] , \in0[2] , \in0[3] , \in0[4] , \in0[5] ,
    \in0[6] , \in0[7] , \in0[8] , \in0[9] , \in0[10] , \in0[11] ,
    \in0[12] , \in0[13] , \in0[14] , \in0[15] , \in0[16] , \in0[17] ,
    \in0[18] , \in0[19] , \in0[20] , \in0[21] , \in0[22] , \in0[23] ,
    \in0[24] , \in0[25] , \in0[26] , \in0[27] , \in0[28] , \in0[29] ,
    \in0[30] , \in0[31] , \in0[32] , \in0[33] , \in0[34] , \in0[35] ,
    \in0[36] , \in0[37] , \in0[38] , \in0[39] , \in0[40] , \in0[41] ,
    \in0[42] , \in0[43] , \in0[44] , \in0[45] , \in0[46] , \in0[47] ,
    \in0[48] , \in0[49] , \in0[50] , \in0[51] , \in0[52] , \in0[53] ,
    \in0[54] , \in0[55] , \in0[56] , \in0[57] , \in0[58] , \in0[59] ,
    \in0[60] , \in0[61] , \in0[62] , \in0[63] , \in0[64] , \in0[65] ,
    \in0[66] , \in0[67] , \in0[68] , \in0[69] , \in0[70] , \in0[71] ,
    \in0[72] , \in0[73] , \in0[74] , \in0[75] , \in0[76] , \in0[77] ,
    \in0[78] , \in0[79] , \in0[80] , \in0[81] , \in0[82] , \in0[83] ,
    \in0[84] , \in0[85] , \in0[86] , \in0[87] , \in0[88] , \in0[89] ,
    \in0[90] , \in0[91] , \in0[92] , \in0[93] , \in0[94] , \in0[95] ,
    \in0[96] , \in0[97] , \in0[98] , \in0[99] , \in0[100] , \in0[101] ,
    \in0[102] , \in0[103] , \in0[104] , \in0[105] , \in0[106] , \in0[107] ,
    \in0[108] , \in0[109] , \in0[110] , \in0[111] , \in0[112] , \in0[113] ,
    \in0[114] , \in0[115] , \in0[116] , \in0[117] , \in0[118] , \in0[119] ,
    \in0[120] , \in0[121] , \in0[122] , \in0[123] , \in0[124] , \in0[125] ,
    \in0[126] , \in0[127] , \in1[0] , \in1[1] , \in1[2] , \in1[3] ,
    \in1[4] , \in1[5] , \in1[6] , \in1[7] , \in1[8] , \in1[9] , \in1[10] ,
    \in1[11] , \in1[12] , \in1[13] , \in1[14] , \in1[15] , \in1[16] ,
    \in1[17] , \in1[18] , \in1[19] , \in1[20] , \in1[21] , \in1[22] ,
    \in1[23] , \in1[24] , \in1[25] , \in1[26] , \in1[27] , \in1[28] ,
    \in1[29] , \in1[30] , \in1[31] , \in1[32] , \in1[33] , \in1[34] ,
    \in1[35] , \in1[36] , \in1[37] , \in1[38] , \in1[39] , \in1[40] ,
    \in1[41] , \in1[42] , \in1[43] , \in1[44] , \in1[45] , \in1[46] ,
    \in1[47] , \in1[48] , \in1[49] , \in1[50] , \in1[51] , \in1[52] ,
    \in1[53] , \in1[54] , \in1[55] , \in1[56] , \in1[57] , \in1[58] ,
    \in1[59] , \in1[60] , \in1[61] , \in1[62] , \in1[63] , \in1[64] ,
    \in1[65] , \in1[66] , \in1[67] , \in1[68] , \in1[69] , \in1[70] ,
    \in1[71] , \in1[72] , \in1[73] , \in1[74] , \in1[75] , \in1[76] ,
    \in1[77] , \in1[78] , \in1[79] , \in1[80] , \in1[81] , \in1[82] ,
    \in1[83] , \in1[84] , \in1[85] , \in1[86] , \in1[87] , \in1[88] ,
    \in1[89] , \in1[90] , \in1[91] , \in1[92] , \in1[93] , \in1[94] ,
    \in1[95] , \in1[96] , \in1[97] , \in1[98] , \in1[99] , \in1[100] ,
    \in1[101] , \in1[102] , \in1[103] , \in1[104] , \in1[105] , \in1[106] ,
    \in1[107] , \in1[108] , \in1[109] , \in1[110] , \in1[111] , \in1[112] ,
    \in1[113] , \in1[114] , \in1[115] , \in1[116] , \in1[117] , \in1[118] ,
    \in1[119] , \in1[120] , \in1[121] , \in1[122] , \in1[123] , \in1[124] ,
    \in1[125] , \in1[126] , \in1[127] , \in2[0] , \in2[1] , \in2[2] ,
    \in2[3] , \in2[4] , \in2[5] , \in2[6] , \in2[7] , \in2[8] , \in2[9] ,
    \in2[10] , \in2[11] , \in2[12] , \in2[13] , \in2[14] , \in2[15] ,
    \in2[16] , \in2[17] , \in2[18] , \in2[19] , \in2[20] , \in2[21] ,
    \in2[22] , \in2[23] , \in2[24] , \in2[25] , \in2[26] , \in2[27] ,
    \in2[28] , \in2[29] , \in2[30] , \in2[31] , \in2[32] , \in2[33] ,
    \in2[34] , \in2[35] , \in2[36] , \in2[37] , \in2[38] , \in2[39] ,
    \in2[40] , \in2[41] , \in2[42] , \in2[43] , \in2[44] , \in2[45] ,
    \in2[46] , \in2[47] , \in2[48] , \in2[49] , \in2[50] , \in2[51] ,
    \in2[52] , \in2[53] , \in2[54] , \in2[55] , \in2[56] , \in2[57] ,
    \in2[58] , \in2[59] , \in2[60] , \in2[61] , \in2[62] , \in2[63] ,
    \in2[64] , \in2[65] , \in2[66] , \in2[67] , \in2[68] , \in2[69] ,
    \in2[70] , \in2[71] , \in2[72] , \in2[73] , \in2[74] , \in2[75] ,
    \in2[76] , \in2[77] , \in2[78] , \in2[79] , \in2[80] , \in2[81] ,
    \in2[82] , \in2[83] , \in2[84] , \in2[85] , \in2[86] , \in2[87] ,
    \in2[88] , \in2[89] , \in2[90] , \in2[91] , \in2[92] , \in2[93] ,
    \in2[94] , \in2[95] , \in2[96] , \in2[97] , \in2[98] , \in2[99] ,
    \in2[100] , \in2[101] , \in2[102] , \in2[103] , \in2[104] , \in2[105] ,
    \in2[106] , \in2[107] , \in2[108] , \in2[109] , \in2[110] , \in2[111] ,
    \in2[112] , \in2[113] , \in2[114] , \in2[115] , \in2[116] , \in2[117] ,
    \in2[118] , \in2[119] , \in2[120] , \in2[121] , \in2[122] , \in2[123] ,
    \in2[124] , \in2[125] , \in2[126] , \in2[127] , \in3[0] , \in3[1] ,
    \in3[2] , \in3[3] , \in3[4] , \in3[5] , \in3[6] , \in3[7] , \in3[8] ,
    \in3[9] , \in3[10] , \in3[11] , \in3[12] , \in3[13] , \in3[14] ,
    \in3[15] , \in3[16] , \in3[17] , \in3[18] , \in3[19] , \in3[20] ,
    \in3[21] , \in3[22] , \in3[23] , \in3[24] , \in3[25] , \in3[26] ,
    \in3[27] , \in3[28] , \in3[29] , \in3[30] , \in3[31] , \in3[32] ,
    \in3[33] , \in3[34] , \in3[35] , \in3[36] , \in3[37] , \in3[38] ,
    \in3[39] , \in3[40] , \in3[41] , \in3[42] , \in3[43] , \in3[44] ,
    \in3[45] , \in3[46] , \in3[47] , \in3[48] , \in3[49] , \in3[50] ,
    \in3[51] , \in3[52] , \in3[53] , \in3[54] , \in3[55] , \in3[56] ,
    \in3[57] , \in3[58] , \in3[59] , \in3[60] , \in3[61] , \in3[62] ,
    \in3[63] , \in3[64] , \in3[65] , \in3[66] , \in3[67] , \in3[68] ,
    \in3[69] , \in3[70] , \in3[71] , \in3[72] , \in3[73] , \in3[74] ,
    \in3[75] , \in3[76] , \in3[77] , \in3[78] , \in3[79] , \in3[80] ,
    \in3[81] , \in3[82] , \in3[83] , \in3[84] , \in3[85] , \in3[86] ,
    \in3[87] , \in3[88] , \in3[89] , \in3[90] , \in3[91] , \in3[92] ,
    \in3[93] , \in3[94] , \in3[95] , \in3[96] , \in3[97] , \in3[98] ,
    \in3[99] , \in3[100] , \in3[101] , \in3[102] , \in3[103] , \in3[104] ,
    \in3[105] , \in3[106] , \in3[107] , \in3[108] , \in3[109] , \in3[110] ,
    \in3[111] , \in3[112] , \in3[113] , \in3[114] , \in3[115] , \in3[116] ,
    \in3[117] , \in3[118] , \in3[119] , \in3[120] , \in3[121] , \in3[122] ,
    \in3[123] , \in3[124] , \in3[125] , \in3[126] , \in3[127] ;
  output \result[0] , \result[1] , \result[2] , \result[3] , \result[4] ,
    \result[5] , \result[6] , \result[7] , \result[8] , \result[9] ,
    \result[10] , \result[11] , \result[12] , \result[13] , \result[14] ,
    \result[15] , \result[16] , \result[17] , \result[18] , \result[19] ,
    \result[20] , \result[21] , \result[22] , \result[23] , \result[24] ,
    \result[25] , \result[26] , \result[27] , \result[28] , \result[29] ,
    \result[30] , \result[31] , \result[32] , \result[33] , \result[34] ,
    \result[35] , \result[36] , \result[37] , \result[38] , \result[39] ,
    \result[40] , \result[41] , \result[42] , \result[43] , \result[44] ,
    \result[45] , \result[46] , \result[47] , \result[48] , \result[49] ,
    \result[50] , \result[51] , \result[52] , \result[53] , \result[54] ,
    \result[55] , \result[56] , \result[57] , \result[58] , \result[59] ,
    \result[60] , \result[61] , \result[62] , \result[63] , \result[64] ,
    \result[65] , \result[66] , \result[67] , \result[68] , \result[69] ,
    \result[70] , \result[71] , \result[72] , \result[73] , \result[74] ,
    \result[75] , \result[76] , \result[77] , \result[78] , \result[79] ,
    \result[80] , \result[81] , \result[82] , \result[83] , \result[84] ,
    \result[85] , \result[86] , \result[87] , \result[88] , \result[89] ,
    \result[90] , \result[91] , \result[92] , \result[93] , \result[94] ,
    \result[95] , \result[96] , \result[97] , \result[98] , \result[99] ,
    \result[100] , \result[101] , \result[102] , \result[103] ,
    \result[104] , \result[105] , \result[106] , \result[107] ,
    \result[108] , \result[109] , \result[110] , \result[111] ,
    \result[112] , \result[113] , \result[114] , \result[115] ,
    \result[116] , \result[117] , \result[118] , \result[119] ,
    \result[120] , \result[121] , \result[122] , \result[123] ,
    \result[124] , \result[125] , \result[126] , \result[127] ,
    \address[0] , \address[1] ;
  wire n642, n643, n644, n645, n646, n647, n648, n649, n650, n651, n652,
    n653, n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
    n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675, n676,
    n677, n678, n679, n680, n681, n682, n683, n684, n685, n686, n687, n688,
    n689, n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
    n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
    n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723, n724,
    n725, n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
    n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
    n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
    n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
    n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783, n784,
    n785, n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
    n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
    n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819, n820,
    n821, n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
    n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
    n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855, n856,
    n857, n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
    n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
    n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
    n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
    n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915, n916,
    n917, n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
    n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
    n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951, n952,
    n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
    n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
    n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987, n988,
    n989, n990, n991, n992, n993, n994, n995, n996, n997, n998, n999,
    n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009,
    n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019,
    n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029,
    n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039,
    n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049,
    n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059,
    n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069,
    n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079,
    n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089,
    n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099,
    n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109,
    n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119,
    n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129,
    n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139,
    n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149,
    n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159,
    n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169,
    n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179,
    n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189,
    n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199,
    n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209,
    n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219,
    n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229,
    n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239,
    n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249,
    n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
    n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
    n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
    n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
    n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
    n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
    n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
    n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
    n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
    n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
    n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
    n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
    n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
    n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
    n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
    n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
    n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
    n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
    n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
    n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
    n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
    n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
    n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
    n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
    n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
    n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
    n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
    n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
    n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
    n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
    n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
    n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
    n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
    n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
    n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
    n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
    n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
    n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
    n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
    n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
    n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
    n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
    n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
    n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
    n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
    n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
    n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
    n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
    n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
    n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
    n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
    n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
    n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
    n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
    n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
    n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
    n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
    n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
    n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
    n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
    n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
    n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
    n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
    n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
    n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
    n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
    n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
    n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
    n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
    n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
    n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
    n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
    n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
    n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
    n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
    n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
    n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
    n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
    n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
    n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
    n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
    n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
    n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
    n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
    n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
    n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
    n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
    n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
    n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
    n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
    n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
    n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
    n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
    n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
    n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
    n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
    n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
    n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
    n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
    n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
    n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
    n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
    n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
    n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
    n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
    n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
    n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
    n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
    n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
    n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
    n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
    n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
    n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
    n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
    n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
    n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
    n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
    n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
    n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
    n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
    n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
    n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
    n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
    n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
    n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
    n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
    n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
    n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
    n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
    n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
    n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
    n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
    n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
    n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
    n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
    n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
    n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
    n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
    n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
    n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
    n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
    n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
    n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
    n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
    n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
    n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
    n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
    n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
    n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
    n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
    n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
    n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
    n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
    n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
    n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
    n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
    n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
    n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
    n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
    n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
    n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
    n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
    n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
    n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
    n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
    n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
    n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
    n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
    n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
    n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
    n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
    n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
    n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009,
    n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019,
    n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029,
    n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039,
    n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
    n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
    n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
    n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079,
    n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089,
    n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099,
    n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109,
    n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119,
    n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129,
    n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139,
    n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
    n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159,
    n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169,
    n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179,
    n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189,
    n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199,
    n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209,
    n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219,
    n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229,
    n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239,
    n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249,
    n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259,
    n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269,
    n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279,
    n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289,
    n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299,
    n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309,
    n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319,
    n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329,
    n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339,
    n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349,
    n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359,
    n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369,
    n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379,
    n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389,
    n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399,
    n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409,
    n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419,
    n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429,
    n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439,
    n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
    n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459,
    n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469,
    n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479,
    n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489,
    n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499,
    n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509,
    n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519,
    n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529,
    n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539,
    n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549,
    n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559,
    n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569,
    n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579,
    n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589,
    n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599,
    n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609,
    n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619,
    n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629,
    n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639,
    n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649,
    n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659,
    n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669,
    n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679,
    n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
    n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
    n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
    n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
    n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
    n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
    n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
    n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
    n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
    n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
    n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
    n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799,
    n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809,
    n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819,
    n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829,
    n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839,
    n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849,
    n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859,
    n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869,
    n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879,
    n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889,
    n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899,
    n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909,
    n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919,
    n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929,
    n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939,
    n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949,
    n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
    n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
    n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
    n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
    n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
    n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009,
    n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019,
    n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029,
    n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
    n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049,
    n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059,
    n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069,
    n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079,
    n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089,
    n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099,
    n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109,
    n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119,
    n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129,
    n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139,
    n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149,
    n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159,
    n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169,
    n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179,
    n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189,
    n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199,
    n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209,
    n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219,
    n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229,
    n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239,
    n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249,
    n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259,
    n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269,
    n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279,
    n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289,
    n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299,
    n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309,
    n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319,
    n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
    n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
    n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
    n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359,
    n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369,
    n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379,
    n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389,
    n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399,
    n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409,
    n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419,
    n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429,
    n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439,
    n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449,
    n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459,
    n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469,
    n4470, n4471, n4472, n4473, n4474, n4475, n4477, n4478, n4479, n4480,
    n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
    n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
    n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
    n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
    n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
    n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
    n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
    n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
    n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
    n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
    n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
    n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
    n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
    n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
    n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
    n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
    n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4651,
    n4652, n4654, n4655, n4657, n4658, n4660, n4661, n4663, n4664, n4666,
    n4667, n4669, n4670, n4672, n4673, n4675, n4676, n4678, n4679, n4681,
    n4682, n4684, n4685, n4687, n4688, n4690, n4691, n4693, n4694, n4696,
    n4697, n4699, n4700, n4702, n4703, n4705, n4706, n4708, n4709, n4711,
    n4712, n4714, n4715, n4717, n4718, n4720, n4721, n4723, n4724, n4726,
    n4727, n4729, n4730, n4732, n4733, n4735, n4736, n4738, n4739, n4741,
    n4742, n4744, n4745, n4747, n4748, n4750, n4751, n4753, n4754, n4756,
    n4757, n4759, n4760, n4762, n4763, n4765, n4766, n4768, n4769, n4771,
    n4772, n4774, n4775, n4777, n4778, n4779, n4781, n4782, n4784, n4785,
    n4787, n4788, n4790, n4791, n4793, n4794, n4796, n4797, n4799, n4800,
    n4802, n4803, n4805, n4806, n4808, n4809, n4811, n4812, n4814, n4815,
    n4817, n4818, n4820, n4821, n4823, n4824, n4826, n4827, n4829, n4830,
    n4832, n4833, n4835, n4836, n4838, n4839, n4841, n4842, n4844, n4845,
    n4847, n4848, n4850, n4851, n4853, n4854, n4856, n4857, n4859, n4860,
    n4862, n4863, n4865, n4866, n4868, n4869, n4871, n4872, n4874, n4875,
    n4877, n4878, n4880, n4881, n4883, n4884, n4886, n4887, n4889, n4890,
    n4892, n4893, n4895, n4896, n4898, n4899, n4901, n4902, n4904, n4905,
    n4907, n4908, n4910, n4911, n4913, n4914, n4916, n4917, n4919, n4920,
    n4922, n4923, n4925, n4926, n4928, n4929, n4931, n4932, n4934, n4935,
    n4937, n4938, n4940, n4941, n4943, n4944, n4946, n4947, n4949, n4950,
    n4952, n4953, n4955, n4956, n4958, n4959, n4961, n4962, n4964, n4965,
    n4967, n4968, n4970, n4971, n4973, n4974, n4976, n4977, n4979, n4980,
    n4982, n4983, n4985, n4986, n4988, n4989, n4991, n4992, n4994, n4995,
    n4997, n4998, n5000, n5001, n5003, n5004, n5006, n5007, n5009, n5010,
    n5012, n5013, n5015, n5016, n5018, n5019, n5021, n5022, n5024, n5025,
    n5027, n5028, n5031, n5032;
  jnot g0000(.din(\in1[123] ), .dout(n642));
  jand g0001(.dina(n642), .dinb(\in0[123] ), .dout(n643));
  jnot g0002(.din(n643), .dout(n644));
  jnot g0003(.din(\in0[120] ), .dout(n645));
  jand g0004(.dina(\in1[120] ), .dinb(n645), .dout(n646));
  jnot g0005(.din(\in0[121] ), .dout(n647));
  jand g0006(.dina(\in1[121] ), .dinb(n647), .dout(n648));
  jor  g0007(.dina(n648), .dinb(n646), .dout(n649));
  jnot g0008(.din(\in0[118] ), .dout(n650));
  jand g0009(.dina(\in1[118] ), .dinb(n650), .dout(n651));
  jnot g0010(.din(\in0[119] ), .dout(n652));
  jand g0011(.dina(\in1[119] ), .dinb(n652), .dout(n653));
  jnot g0012(.din(\in0[117] ), .dout(n654));
  jand g0013(.dina(\in1[117] ), .dinb(n654), .dout(n655));
  jor  g0014(.dina(n655), .dinb(n653), .dout(n656));
  jor  g0015(.dina(n656), .dinb(n651), .dout(n657));
  jnot g0016(.din(n657), .dout(n658));
  jnot g0017(.din(\in1[117] ), .dout(n659));
  jand g0018(.dina(n659), .dinb(\in0[117] ), .dout(n660));
  jnot g0019(.din(\in1[116] ), .dout(n661));
  jand g0020(.dina(n661), .dinb(\in0[116] ), .dout(n662));
  jor  g0021(.dina(n662), .dinb(n660), .dout(n663));
  jand g0022(.dina(n663), .dinb(n658), .dout(n664));
  jnot g0023(.din(n653), .dout(n665));
  jnot g0024(.din(\in1[119] ), .dout(n666));
  jand g0025(.dina(n666), .dinb(\in0[119] ), .dout(n667));
  jnot g0026(.din(\in1[118] ), .dout(n668));
  jand g0027(.dina(n668), .dinb(\in0[118] ), .dout(n669));
  jor  g0028(.dina(n669), .dinb(n667), .dout(n670));
  jand g0029(.dina(n670), .dinb(n665), .dout(n671));
  jor  g0030(.dina(n671), .dinb(n664), .dout(n672));
  jnot g0031(.din(n672), .dout(n673));
  jnot g0032(.din(\in1[115] ), .dout(n674));
  jand g0033(.dina(n674), .dinb(\in0[115] ), .dout(n675));
  jnot g0034(.din(n675), .dout(n676));
  jnot g0035(.din(\in0[113] ), .dout(n677));
  jand g0036(.dina(\in1[113] ), .dinb(n677), .dout(n678));
  jnot g0037(.din(\in0[112] ), .dout(n679));
  jand g0038(.dina(\in1[112] ), .dinb(n679), .dout(n680));
  jor  g0039(.dina(n680), .dinb(n678), .dout(n681));
  jnot g0040(.din(\in0[110] ), .dout(n682));
  jand g0041(.dina(\in1[110] ), .dinb(n682), .dout(n683));
  jnot g0042(.din(\in0[111] ), .dout(n684));
  jand g0043(.dina(\in1[111] ), .dinb(n684), .dout(n685));
  jnot g0044(.din(\in0[109] ), .dout(n686));
  jand g0045(.dina(\in1[109] ), .dinb(n686), .dout(n687));
  jor  g0046(.dina(n687), .dinb(n685), .dout(n688));
  jor  g0047(.dina(n688), .dinb(n683), .dout(n689));
  jnot g0048(.din(n689), .dout(n690));
  jnot g0049(.din(\in1[109] ), .dout(n691));
  jand g0050(.dina(n691), .dinb(\in0[109] ), .dout(n692));
  jnot g0051(.din(\in1[108] ), .dout(n693));
  jand g0052(.dina(n693), .dinb(\in0[108] ), .dout(n694));
  jor  g0053(.dina(n694), .dinb(n692), .dout(n695));
  jand g0054(.dina(n695), .dinb(n690), .dout(n696));
  jnot g0055(.din(n685), .dout(n697));
  jnot g0056(.din(\in1[111] ), .dout(n698));
  jand g0057(.dina(n698), .dinb(\in0[111] ), .dout(n699));
  jnot g0058(.din(\in1[110] ), .dout(n700));
  jand g0059(.dina(n700), .dinb(\in0[110] ), .dout(n701));
  jor  g0060(.dina(n701), .dinb(n699), .dout(n702));
  jand g0061(.dina(n702), .dinb(n697), .dout(n703));
  jor  g0062(.dina(n703), .dinb(n696), .dout(n704));
  jnot g0063(.din(n704), .dout(n705));
  jnot g0064(.din(\in1[107] ), .dout(n706));
  jand g0065(.dina(n706), .dinb(\in0[107] ), .dout(n707));
  jnot g0066(.din(n707), .dout(n708));
  jnot g0067(.din(\in0[104] ), .dout(n709));
  jand g0068(.dina(\in1[104] ), .dinb(n709), .dout(n710));
  jnot g0069(.din(\in0[105] ), .dout(n711));
  jand g0070(.dina(\in1[105] ), .dinb(n711), .dout(n712));
  jor  g0071(.dina(n712), .dinb(n710), .dout(n713));
  jnot g0072(.din(\in0[102] ), .dout(n714));
  jand g0073(.dina(\in1[102] ), .dinb(n714), .dout(n715));
  jnot g0074(.din(\in0[103] ), .dout(n716));
  jand g0075(.dina(\in1[103] ), .dinb(n716), .dout(n717));
  jnot g0076(.din(\in0[101] ), .dout(n718));
  jand g0077(.dina(\in1[101] ), .dinb(n718), .dout(n719));
  jor  g0078(.dina(n719), .dinb(n717), .dout(n720));
  jor  g0079(.dina(n720), .dinb(n715), .dout(n721));
  jnot g0080(.din(n721), .dout(n722));
  jnot g0081(.din(\in1[101] ), .dout(n723));
  jand g0082(.dina(n723), .dinb(\in0[101] ), .dout(n724));
  jnot g0083(.din(\in1[100] ), .dout(n725));
  jand g0084(.dina(n725), .dinb(\in0[100] ), .dout(n726));
  jor  g0085(.dina(n726), .dinb(n724), .dout(n727));
  jand g0086(.dina(n727), .dinb(n722), .dout(n728));
  jnot g0087(.din(n717), .dout(n729));
  jnot g0088(.din(\in1[103] ), .dout(n730));
  jand g0089(.dina(n730), .dinb(\in0[103] ), .dout(n731));
  jnot g0090(.din(\in1[102] ), .dout(n732));
  jand g0091(.dina(n732), .dinb(\in0[102] ), .dout(n733));
  jor  g0092(.dina(n733), .dinb(n731), .dout(n734));
  jand g0093(.dina(n734), .dinb(n729), .dout(n735));
  jor  g0094(.dina(n735), .dinb(n728), .dout(n736));
  jnot g0095(.din(n736), .dout(n737));
  jnot g0096(.din(\in1[99] ), .dout(n738));
  jand g0097(.dina(n738), .dinb(\in0[99] ), .dout(n739));
  jnot g0098(.din(n739), .dout(n740));
  jnot g0099(.din(\in0[97] ), .dout(n741));
  jand g0100(.dina(\in1[97] ), .dinb(n741), .dout(n742));
  jnot g0101(.din(\in0[96] ), .dout(n743));
  jand g0102(.dina(\in1[96] ), .dinb(n743), .dout(n744));
  jor  g0103(.dina(n744), .dinb(n742), .dout(n745));
  jnot g0104(.din(\in0[94] ), .dout(n746));
  jand g0105(.dina(\in1[94] ), .dinb(n746), .dout(n747));
  jnot g0106(.din(\in0[95] ), .dout(n748));
  jand g0107(.dina(\in1[95] ), .dinb(n748), .dout(n749));
  jnot g0108(.din(\in0[93] ), .dout(n750));
  jand g0109(.dina(\in1[93] ), .dinb(n750), .dout(n751));
  jor  g0110(.dina(n751), .dinb(n749), .dout(n752));
  jor  g0111(.dina(n752), .dinb(n747), .dout(n753));
  jnot g0112(.din(n753), .dout(n754));
  jnot g0113(.din(\in1[93] ), .dout(n755));
  jand g0114(.dina(n755), .dinb(\in0[93] ), .dout(n756));
  jnot g0115(.din(\in1[92] ), .dout(n757));
  jand g0116(.dina(n757), .dinb(\in0[92] ), .dout(n758));
  jor  g0117(.dina(n758), .dinb(n756), .dout(n759));
  jand g0118(.dina(n759), .dinb(n754), .dout(n760));
  jnot g0119(.din(n749), .dout(n761));
  jnot g0120(.din(\in1[95] ), .dout(n762));
  jand g0121(.dina(n762), .dinb(\in0[95] ), .dout(n763));
  jnot g0122(.din(\in1[94] ), .dout(n764));
  jand g0123(.dina(n764), .dinb(\in0[94] ), .dout(n765));
  jor  g0124(.dina(n765), .dinb(n763), .dout(n766));
  jand g0125(.dina(n766), .dinb(n761), .dout(n767));
  jor  g0126(.dina(n767), .dinb(n760), .dout(n768));
  jnot g0127(.din(n768), .dout(n769));
  jnot g0128(.din(\in1[91] ), .dout(n770));
  jand g0129(.dina(n770), .dinb(\in0[91] ), .dout(n771));
  jnot g0130(.din(n771), .dout(n772));
  jnot g0131(.din(\in0[86] ), .dout(n773));
  jand g0132(.dina(\in1[86] ), .dinb(n773), .dout(n774));
  jnot g0133(.din(\in0[87] ), .dout(n775));
  jand g0134(.dina(\in1[87] ), .dinb(n775), .dout(n776));
  jnot g0135(.din(\in0[85] ), .dout(n777));
  jand g0136(.dina(\in1[85] ), .dinb(n777), .dout(n778));
  jor  g0137(.dina(n778), .dinb(n776), .dout(n779));
  jor  g0138(.dina(n779), .dinb(n774), .dout(n780));
  jnot g0139(.din(n780), .dout(n781));
  jnot g0140(.din(\in1[85] ), .dout(n782));
  jand g0141(.dina(n782), .dinb(\in0[85] ), .dout(n783));
  jnot g0142(.din(\in1[84] ), .dout(n784));
  jand g0143(.dina(n784), .dinb(\in0[84] ), .dout(n785));
  jor  g0144(.dina(n785), .dinb(n783), .dout(n786));
  jand g0145(.dina(n786), .dinb(n781), .dout(n787));
  jnot g0146(.din(n776), .dout(n788));
  jnot g0147(.din(\in1[87] ), .dout(n789));
  jand g0148(.dina(n789), .dinb(\in0[87] ), .dout(n790));
  jnot g0149(.din(\in1[86] ), .dout(n791));
  jand g0150(.dina(n791), .dinb(\in0[86] ), .dout(n792));
  jor  g0151(.dina(n792), .dinb(n790), .dout(n793));
  jand g0152(.dina(n793), .dinb(n788), .dout(n794));
  jor  g0153(.dina(n794), .dinb(n787), .dout(n795));
  jnot g0154(.din(n795), .dout(n796));
  jnot g0155(.din(\in1[83] ), .dout(n797));
  jand g0156(.dina(n797), .dinb(\in0[83] ), .dout(n798));
  jnot g0157(.din(n798), .dout(n799));
  jnot g0158(.din(\in0[81] ), .dout(n800));
  jand g0159(.dina(\in1[81] ), .dinb(n800), .dout(n801));
  jnot g0160(.din(\in0[80] ), .dout(n802));
  jand g0161(.dina(\in1[80] ), .dinb(n802), .dout(n803));
  jor  g0162(.dina(n803), .dinb(n801), .dout(n804));
  jnot g0163(.din(\in0[78] ), .dout(n805));
  jand g0164(.dina(\in1[78] ), .dinb(n805), .dout(n806));
  jnot g0165(.din(\in0[79] ), .dout(n807));
  jand g0166(.dina(\in1[79] ), .dinb(n807), .dout(n808));
  jnot g0167(.din(\in0[77] ), .dout(n809));
  jand g0168(.dina(\in1[77] ), .dinb(n809), .dout(n810));
  jor  g0169(.dina(n810), .dinb(n808), .dout(n811));
  jor  g0170(.dina(n811), .dinb(n806), .dout(n812));
  jnot g0171(.din(n812), .dout(n813));
  jnot g0172(.din(\in1[77] ), .dout(n814));
  jand g0173(.dina(n814), .dinb(\in0[77] ), .dout(n815));
  jnot g0174(.din(\in1[76] ), .dout(n816));
  jand g0175(.dina(n816), .dinb(\in0[76] ), .dout(n817));
  jor  g0176(.dina(n817), .dinb(n815), .dout(n818));
  jand g0177(.dina(n818), .dinb(n813), .dout(n819));
  jnot g0178(.din(n808), .dout(n820));
  jnot g0179(.din(\in1[79] ), .dout(n821));
  jand g0180(.dina(n821), .dinb(\in0[79] ), .dout(n822));
  jnot g0181(.din(\in1[78] ), .dout(n823));
  jand g0182(.dina(n823), .dinb(\in0[78] ), .dout(n824));
  jor  g0183(.dina(n824), .dinb(n822), .dout(n825));
  jand g0184(.dina(n825), .dinb(n820), .dout(n826));
  jor  g0185(.dina(n826), .dinb(n819), .dout(n827));
  jnot g0186(.din(n827), .dout(n828));
  jnot g0187(.din(\in1[75] ), .dout(n829));
  jand g0188(.dina(n829), .dinb(\in0[75] ), .dout(n830));
  jnot g0189(.din(n830), .dout(n831));
  jnot g0190(.din(\in0[72] ), .dout(n832));
  jand g0191(.dina(\in1[72] ), .dinb(n832), .dout(n833));
  jnot g0192(.din(\in0[73] ), .dout(n834));
  jand g0193(.dina(\in1[73] ), .dinb(n834), .dout(n835));
  jor  g0194(.dina(n835), .dinb(n833), .dout(n836));
  jnot g0195(.din(\in0[70] ), .dout(n837));
  jand g0196(.dina(\in1[70] ), .dinb(n837), .dout(n838));
  jnot g0197(.din(\in0[71] ), .dout(n839));
  jand g0198(.dina(\in1[71] ), .dinb(n839), .dout(n840));
  jnot g0199(.din(\in0[69] ), .dout(n841));
  jand g0200(.dina(\in1[69] ), .dinb(n841), .dout(n842));
  jor  g0201(.dina(n842), .dinb(n840), .dout(n843));
  jor  g0202(.dina(n843), .dinb(n838), .dout(n844));
  jnot g0203(.din(n844), .dout(n845));
  jnot g0204(.din(\in1[69] ), .dout(n846));
  jand g0205(.dina(n846), .dinb(\in0[69] ), .dout(n847));
  jnot g0206(.din(\in1[68] ), .dout(n848));
  jand g0207(.dina(n848), .dinb(\in0[68] ), .dout(n849));
  jor  g0208(.dina(n849), .dinb(n847), .dout(n850));
  jand g0209(.dina(n850), .dinb(n845), .dout(n851));
  jnot g0210(.din(n840), .dout(n852));
  jnot g0211(.din(\in1[71] ), .dout(n853));
  jand g0212(.dina(n853), .dinb(\in0[71] ), .dout(n854));
  jnot g0213(.din(\in1[70] ), .dout(n855));
  jand g0214(.dina(n855), .dinb(\in0[70] ), .dout(n856));
  jor  g0215(.dina(n856), .dinb(n854), .dout(n857));
  jand g0216(.dina(n857), .dinb(n852), .dout(n858));
  jor  g0217(.dina(n858), .dinb(n851), .dout(n859));
  jnot g0218(.din(n859), .dout(n860));
  jnot g0219(.din(\in1[67] ), .dout(n861));
  jand g0220(.dina(n861), .dinb(\in0[67] ), .dout(n862));
  jnot g0221(.din(n862), .dout(n863));
  jnot g0222(.din(\in0[65] ), .dout(n864));
  jand g0223(.dina(\in1[65] ), .dinb(n864), .dout(n865));
  jnot g0224(.din(n865), .dout(n866));
  jnot g0225(.din(\in1[64] ), .dout(n867));
  jand g0226(.dina(n867), .dinb(\in0[64] ), .dout(n868));
  jand g0227(.dina(n868), .dinb(n866), .dout(n869));
  jnot g0228(.din(\in1[66] ), .dout(n870));
  jand g0229(.dina(n870), .dinb(\in0[66] ), .dout(n871));
  jnot g0230(.din(\in1[65] ), .dout(n872));
  jand g0231(.dina(n872), .dinb(\in0[65] ), .dout(n873));
  jor  g0232(.dina(n873), .dinb(n871), .dout(n874));
  jor  g0233(.dina(n874), .dinb(n869), .dout(n875));
  jnot g0234(.din(n875), .dout(n876));
  jnot g0235(.din(\in1[59] ), .dout(n877));
  jnot g0236(.din(\in0[60] ), .dout(n878));
  jand g0237(.dina(\in1[60] ), .dinb(n878), .dout(n879));
  jnot g0238(.din(\in0[63] ), .dout(n880));
  jand g0239(.dina(\in1[63] ), .dinb(n880), .dout(n881));
  jnot g0240(.din(\in0[61] ), .dout(n882));
  jand g0241(.dina(\in1[61] ), .dinb(n882), .dout(n883));
  jnot g0242(.din(\in0[62] ), .dout(n884));
  jand g0243(.dina(\in1[62] ), .dinb(n884), .dout(n885));
  jor  g0244(.dina(n885), .dinb(n883), .dout(n886));
  jor  g0245(.dina(n886), .dinb(n881), .dout(n887));
  jor  g0246(.dina(n887), .dinb(n879), .dout(n888));
  jnot g0247(.din(n888), .dout(n889));
  jand g0248(.dina(n889), .dinb(\in0[59] ), .dout(n890));
  jand g0249(.dina(n890), .dinb(n877), .dout(n891));
  jnot g0250(.din(n891), .dout(n892));
  jnot g0251(.din(\in1[51] ), .dout(n893));
  jnot g0252(.din(\in0[53] ), .dout(n894));
  jand g0253(.dina(\in1[53] ), .dinb(n894), .dout(n895));
  jnot g0254(.din(\in0[55] ), .dout(n896));
  jand g0255(.dina(\in1[55] ), .dinb(n896), .dout(n897));
  jnot g0256(.din(\in0[54] ), .dout(n898));
  jand g0257(.dina(\in1[54] ), .dinb(n898), .dout(n899));
  jor  g0258(.dina(n899), .dinb(n897), .dout(n900));
  jnot g0259(.din(\in0[52] ), .dout(n901));
  jand g0260(.dina(\in1[52] ), .dinb(n901), .dout(n902));
  jor  g0261(.dina(n902), .dinb(n900), .dout(n903));
  jor  g0262(.dina(n903), .dinb(n895), .dout(n904));
  jnot g0263(.din(n904), .dout(n905));
  jand g0264(.dina(n905), .dinb(\in0[51] ), .dout(n906));
  jand g0265(.dina(n906), .dinb(n893), .dout(n907));
  jnot g0266(.din(n907), .dout(n908));
  jnot g0267(.din(\in0[44] ), .dout(n909));
  jand g0268(.dina(\in1[44] ), .dinb(n909), .dout(n910));
  jnot g0269(.din(\in0[47] ), .dout(n911));
  jand g0270(.dina(\in1[47] ), .dinb(n911), .dout(n912));
  jnot g0271(.din(\in0[45] ), .dout(n913));
  jand g0272(.dina(\in1[45] ), .dinb(n913), .dout(n914));
  jnot g0273(.din(\in0[46] ), .dout(n915));
  jand g0274(.dina(\in1[46] ), .dinb(n915), .dout(n916));
  jor  g0275(.dina(n916), .dinb(n914), .dout(n917));
  jor  g0276(.dina(n917), .dinb(n912), .dout(n918));
  jor  g0277(.dina(n918), .dinb(n910), .dout(n919));
  jnot g0278(.din(\in0[42] ), .dout(n920));
  jand g0279(.dina(\in1[42] ), .dinb(n920), .dout(n921));
  jnot g0280(.din(\in0[43] ), .dout(n922));
  jand g0281(.dina(\in1[43] ), .dinb(n922), .dout(n923));
  jor  g0282(.dina(n923), .dinb(n921), .dout(n924));
  jor  g0283(.dina(n924), .dinb(n919), .dout(n925));
  jnot g0284(.din(n925), .dout(n926));
  jnot g0285(.din(\in1[42] ), .dout(n927));
  jand g0286(.dina(n927), .dinb(\in0[42] ), .dout(n928));
  jnot g0287(.din(\in1[41] ), .dout(n929));
  jand g0288(.dina(n929), .dinb(\in0[41] ), .dout(n930));
  jnot g0289(.din(\in0[41] ), .dout(n931));
  jand g0290(.dina(\in1[41] ), .dinb(n931), .dout(n932));
  jnot g0291(.din(n932), .dout(n933));
  jnot g0292(.din(\in1[40] ), .dout(n934));
  jand g0293(.dina(n934), .dinb(\in0[40] ), .dout(n935));
  jand g0294(.dina(n935), .dinb(n933), .dout(n936));
  jor  g0295(.dina(n936), .dinb(n930), .dout(n937));
  jor  g0296(.dina(n937), .dinb(n928), .dout(n938));
  jand g0297(.dina(n938), .dinb(n926), .dout(n939));
  jnot g0298(.din(n939), .dout(n940));
  jnot g0299(.din(\in1[33] ), .dout(n941));
  jand g0300(.dina(n941), .dinb(\in0[33] ), .dout(n942));
  jnot g0301(.din(\in1[34] ), .dout(n943));
  jand g0302(.dina(n943), .dinb(\in0[34] ), .dout(n944));
  jor  g0303(.dina(n944), .dinb(n942), .dout(n945));
  jnot g0304(.din(\in0[33] ), .dout(n946));
  jand g0305(.dina(\in1[33] ), .dinb(n946), .dout(n947));
  jnot g0306(.din(n947), .dout(n948));
  jnot g0307(.din(\in1[32] ), .dout(n949));
  jand g0308(.dina(n949), .dinb(\in0[32] ), .dout(n950));
  jand g0309(.dina(n950), .dinb(n948), .dout(n951));
  jor  g0310(.dina(n951), .dinb(n945), .dout(n952));
  jnot g0311(.din(\in0[35] ), .dout(n953));
  jand g0312(.dina(\in1[35] ), .dinb(n953), .dout(n954));
  jnot g0313(.din(\in0[34] ), .dout(n955));
  jand g0314(.dina(\in1[34] ), .dinb(n955), .dout(n956));
  jor  g0315(.dina(n956), .dinb(n954), .dout(n957));
  jnot g0316(.din(\in0[36] ), .dout(n958));
  jand g0317(.dina(\in1[36] ), .dinb(n958), .dout(n959));
  jnot g0318(.din(\in0[38] ), .dout(n960));
  jand g0319(.dina(\in1[38] ), .dinb(n960), .dout(n961));
  jnot g0320(.din(\in0[39] ), .dout(n962));
  jand g0321(.dina(\in1[39] ), .dinb(n962), .dout(n963));
  jnot g0322(.din(\in0[37] ), .dout(n964));
  jand g0323(.dina(\in1[37] ), .dinb(n964), .dout(n965));
  jor  g0324(.dina(n965), .dinb(n963), .dout(n966));
  jor  g0325(.dina(n966), .dinb(n961), .dout(n967));
  jor  g0326(.dina(n967), .dinb(n959), .dout(n968));
  jor  g0327(.dina(n968), .dinb(n957), .dout(n969));
  jnot g0328(.din(n969), .dout(n970));
  jand g0329(.dina(n970), .dinb(n952), .dout(n971));
  jnot g0330(.din(n971), .dout(n972));
  jnot g0331(.din(\in0[30] ), .dout(n973));
  jand g0332(.dina(\in1[30] ), .dinb(n973), .dout(n974));
  jnot g0333(.din(\in1[29] ), .dout(n975));
  jand g0334(.dina(n975), .dinb(\in0[29] ), .dout(n976));
  jnot g0335(.din(n976), .dout(n977));
  jnot g0336(.din(\in0[29] ), .dout(n978));
  jand g0337(.dina(\in1[29] ), .dinb(n978), .dout(n979));
  jnot g0338(.din(\in1[28] ), .dout(n980));
  jand g0339(.dina(n980), .dinb(\in0[28] ), .dout(n981));
  jnot g0340(.din(n981), .dout(n982));
  jnot g0341(.din(\in0[28] ), .dout(n983));
  jand g0342(.dina(\in1[28] ), .dinb(n983), .dout(n984));
  jnot g0343(.din(\in1[27] ), .dout(n985));
  jand g0344(.dina(n985), .dinb(\in0[27] ), .dout(n986));
  jnot g0345(.din(n986), .dout(n987));
  jnot g0346(.din(\in0[27] ), .dout(n988));
  jand g0347(.dina(\in1[27] ), .dinb(n988), .dout(n989));
  jnot g0348(.din(\in1[26] ), .dout(n990));
  jand g0349(.dina(n990), .dinb(\in0[26] ), .dout(n991));
  jnot g0350(.din(n991), .dout(n992));
  jnot g0351(.din(\in0[23] ), .dout(n993));
  jand g0352(.dina(\in1[23] ), .dinb(n993), .dout(n994));
  jnot g0353(.din(\in0[22] ), .dout(n995));
  jand g0354(.dina(\in1[22] ), .dinb(n995), .dout(n996));
  jnot g0355(.din(\in1[21] ), .dout(n997));
  jand g0356(.dina(n997), .dinb(\in0[21] ), .dout(n998));
  jnot g0357(.din(n998), .dout(n999));
  jnot g0358(.din(\in0[21] ), .dout(n1000));
  jand g0359(.dina(\in1[21] ), .dinb(n1000), .dout(n1001));
  jnot g0360(.din(\in1[20] ), .dout(n1002));
  jand g0361(.dina(n1002), .dinb(\in0[20] ), .dout(n1003));
  jnot g0362(.din(n1003), .dout(n1004));
  jnot g0363(.din(\in0[20] ), .dout(n1005));
  jand g0364(.dina(\in1[20] ), .dinb(n1005), .dout(n1006));
  jnot g0365(.din(\in1[19] ), .dout(n1007));
  jand g0366(.dina(n1007), .dinb(\in0[19] ), .dout(n1008));
  jnot g0367(.din(n1008), .dout(n1009));
  jnot g0368(.din(\in0[19] ), .dout(n1010));
  jand g0369(.dina(\in1[19] ), .dinb(n1010), .dout(n1011));
  jnot g0370(.din(\in1[18] ), .dout(n1012));
  jand g0371(.dina(n1012), .dinb(\in0[18] ), .dout(n1013));
  jnot g0372(.din(n1013), .dout(n1014));
  jnot g0373(.din(\in0[15] ), .dout(n1015));
  jand g0374(.dina(\in1[15] ), .dinb(n1015), .dout(n1016));
  jnot g0375(.din(\in0[14] ), .dout(n1017));
  jand g0376(.dina(\in1[14] ), .dinb(n1017), .dout(n1018));
  jnot g0377(.din(\in1[13] ), .dout(n1019));
  jand g0378(.dina(n1019), .dinb(\in0[13] ), .dout(n1020));
  jnot g0379(.din(n1020), .dout(n1021));
  jnot g0380(.din(\in0[13] ), .dout(n1022));
  jand g0381(.dina(\in1[13] ), .dinb(n1022), .dout(n1023));
  jnot g0382(.din(\in1[12] ), .dout(n1024));
  jand g0383(.dina(n1024), .dinb(\in0[12] ), .dout(n1025));
  jnot g0384(.din(n1025), .dout(n1026));
  jnot g0385(.din(\in0[12] ), .dout(n1027));
  jand g0386(.dina(\in1[12] ), .dinb(n1027), .dout(n1028));
  jnot g0387(.din(\in1[11] ), .dout(n1029));
  jand g0388(.dina(n1029), .dinb(\in0[11] ), .dout(n1030));
  jnot g0389(.din(n1030), .dout(n1031));
  jnot g0390(.din(\in0[11] ), .dout(n1032));
  jand g0391(.dina(\in1[11] ), .dinb(n1032), .dout(n1033));
  jnot g0392(.din(\in1[10] ), .dout(n1034));
  jand g0393(.dina(n1034), .dinb(\in0[10] ), .dout(n1035));
  jnot g0394(.din(n1035), .dout(n1036));
  jnot g0395(.din(\in0[7] ), .dout(n1037));
  jand g0396(.dina(\in1[7] ), .dinb(n1037), .dout(n1038));
  jnot g0397(.din(\in0[3] ), .dout(n1039));
  jand g0398(.dina(\in1[3] ), .dinb(n1039), .dout(n1040));
  jnot g0399(.din(\in1[2] ), .dout(n1041));
  jand g0400(.dina(n1041), .dinb(\in0[2] ), .dout(n1042));
  jnot g0401(.din(n1042), .dout(n1043));
  jnot g0402(.din(\in0[1] ), .dout(n1044));
  jor  g0403(.dina(\in1[1] ), .dinb(n1044), .dout(n1045));
  jnot g0404(.din(\in0[0] ), .dout(n1046));
  jor  g0405(.dina(\in1[0] ), .dinb(n1046), .dout(n1047));
  jand g0406(.dina(n1047), .dinb(n1045), .dout(n1048));
  jnot g0407(.din(\in0[2] ), .dout(n1049));
  jand g0408(.dina(\in1[2] ), .dinb(n1049), .dout(n1050));
  jand g0409(.dina(\in1[1] ), .dinb(n1044), .dout(n1051));
  jor  g0410(.dina(n1051), .dinb(n1050), .dout(n1052));
  jor  g0411(.dina(n1052), .dinb(n1048), .dout(n1053));
  jnot g0412(.din(\in1[3] ), .dout(n1054));
  jand g0413(.dina(n1054), .dinb(\in0[3] ), .dout(n1055));
  jnot g0414(.din(n1055), .dout(n1056));
  jand g0415(.dina(n1056), .dinb(n1053), .dout(n1057));
  jand g0416(.dina(n1057), .dinb(n1043), .dout(n1058));
  jnot g0417(.din(\in0[4] ), .dout(n1059));
  jand g0418(.dina(\in1[4] ), .dinb(n1059), .dout(n1060));
  jor  g0419(.dina(n1060), .dinb(n1058), .dout(n1061));
  jor  g0420(.dina(n1061), .dinb(n1040), .dout(n1062));
  jnot g0421(.din(\in1[4] ), .dout(n1063));
  jand g0422(.dina(n1063), .dinb(\in0[4] ), .dout(n1064));
  jnot g0423(.din(\in1[5] ), .dout(n1065));
  jand g0424(.dina(n1065), .dinb(\in0[5] ), .dout(n1066));
  jor  g0425(.dina(n1066), .dinb(n1064), .dout(n1067));
  jnot g0426(.din(n1067), .dout(n1068));
  jand g0427(.dina(n1068), .dinb(n1062), .dout(n1069));
  jnot g0428(.din(\in0[6] ), .dout(n1070));
  jand g0429(.dina(\in1[6] ), .dinb(n1070), .dout(n1071));
  jnot g0430(.din(\in0[5] ), .dout(n1072));
  jand g0431(.dina(\in1[5] ), .dinb(n1072), .dout(n1073));
  jor  g0432(.dina(n1073), .dinb(n1071), .dout(n1074));
  jor  g0433(.dina(n1074), .dinb(n1069), .dout(n1075));
  jnot g0434(.din(\in1[7] ), .dout(n1076));
  jand g0435(.dina(n1076), .dinb(\in0[7] ), .dout(n1077));
  jnot g0436(.din(\in1[6] ), .dout(n1078));
  jand g0437(.dina(n1078), .dinb(\in0[6] ), .dout(n1079));
  jor  g0438(.dina(n1079), .dinb(n1077), .dout(n1080));
  jnot g0439(.din(n1080), .dout(n1081));
  jand g0440(.dina(n1081), .dinb(n1075), .dout(n1082));
  jnot g0441(.din(\in0[8] ), .dout(n1083));
  jand g0442(.dina(\in1[8] ), .dinb(n1083), .dout(n1084));
  jor  g0443(.dina(n1084), .dinb(n1082), .dout(n1085));
  jor  g0444(.dina(n1085), .dinb(n1038), .dout(n1086));
  jnot g0445(.din(\in1[8] ), .dout(n1087));
  jand g0446(.dina(n1087), .dinb(\in0[8] ), .dout(n1088));
  jnot g0447(.din(\in1[9] ), .dout(n1089));
  jand g0448(.dina(n1089), .dinb(\in0[9] ), .dout(n1090));
  jor  g0449(.dina(n1090), .dinb(n1088), .dout(n1091));
  jnot g0450(.din(n1091), .dout(n1092));
  jand g0451(.dina(n1092), .dinb(n1086), .dout(n1093));
  jnot g0452(.din(\in0[10] ), .dout(n1094));
  jand g0453(.dina(\in1[10] ), .dinb(n1094), .dout(n1095));
  jnot g0454(.din(\in0[9] ), .dout(n1096));
  jand g0455(.dina(\in1[9] ), .dinb(n1096), .dout(n1097));
  jor  g0456(.dina(n1097), .dinb(n1095), .dout(n1098));
  jor  g0457(.dina(n1098), .dinb(n1093), .dout(n1099));
  jand g0458(.dina(n1099), .dinb(n1036), .dout(n1100));
  jor  g0459(.dina(n1100), .dinb(n1033), .dout(n1101));
  jand g0460(.dina(n1101), .dinb(n1031), .dout(n1102));
  jor  g0461(.dina(n1102), .dinb(n1028), .dout(n1103));
  jand g0462(.dina(n1103), .dinb(n1026), .dout(n1104));
  jor  g0463(.dina(n1104), .dinb(n1023), .dout(n1105));
  jand g0464(.dina(n1105), .dinb(n1021), .dout(n1106));
  jor  g0465(.dina(n1106), .dinb(n1018), .dout(n1107));
  jnot g0466(.din(\in1[15] ), .dout(n1108));
  jand g0467(.dina(n1108), .dinb(\in0[15] ), .dout(n1109));
  jnot g0468(.din(\in1[14] ), .dout(n1110));
  jand g0469(.dina(n1110), .dinb(\in0[14] ), .dout(n1111));
  jor  g0470(.dina(n1111), .dinb(n1109), .dout(n1112));
  jnot g0471(.din(n1112), .dout(n1113));
  jand g0472(.dina(n1113), .dinb(n1107), .dout(n1114));
  jnot g0473(.din(\in0[16] ), .dout(n1115));
  jand g0474(.dina(\in1[16] ), .dinb(n1115), .dout(n1116));
  jor  g0475(.dina(n1116), .dinb(n1114), .dout(n1117));
  jor  g0476(.dina(n1117), .dinb(n1016), .dout(n1118));
  jnot g0477(.din(\in1[16] ), .dout(n1119));
  jand g0478(.dina(n1119), .dinb(\in0[16] ), .dout(n1120));
  jnot g0479(.din(\in1[17] ), .dout(n1121));
  jand g0480(.dina(n1121), .dinb(\in0[17] ), .dout(n1122));
  jor  g0481(.dina(n1122), .dinb(n1120), .dout(n1123));
  jnot g0482(.din(n1123), .dout(n1124));
  jand g0483(.dina(n1124), .dinb(n1118), .dout(n1125));
  jnot g0484(.din(\in0[18] ), .dout(n1126));
  jand g0485(.dina(\in1[18] ), .dinb(n1126), .dout(n1127));
  jnot g0486(.din(\in0[17] ), .dout(n1128));
  jand g0487(.dina(\in1[17] ), .dinb(n1128), .dout(n1129));
  jor  g0488(.dina(n1129), .dinb(n1127), .dout(n1130));
  jor  g0489(.dina(n1130), .dinb(n1125), .dout(n1131));
  jand g0490(.dina(n1131), .dinb(n1014), .dout(n1132));
  jor  g0491(.dina(n1132), .dinb(n1011), .dout(n1133));
  jand g0492(.dina(n1133), .dinb(n1009), .dout(n1134));
  jor  g0493(.dina(n1134), .dinb(n1006), .dout(n1135));
  jand g0494(.dina(n1135), .dinb(n1004), .dout(n1136));
  jor  g0495(.dina(n1136), .dinb(n1001), .dout(n1137));
  jand g0496(.dina(n1137), .dinb(n999), .dout(n1138));
  jor  g0497(.dina(n1138), .dinb(n996), .dout(n1139));
  jnot g0498(.din(\in1[23] ), .dout(n1140));
  jand g0499(.dina(n1140), .dinb(\in0[23] ), .dout(n1141));
  jnot g0500(.din(\in1[22] ), .dout(n1142));
  jand g0501(.dina(n1142), .dinb(\in0[22] ), .dout(n1143));
  jor  g0502(.dina(n1143), .dinb(n1141), .dout(n1144));
  jnot g0503(.din(n1144), .dout(n1145));
  jand g0504(.dina(n1145), .dinb(n1139), .dout(n1146));
  jnot g0505(.din(\in0[24] ), .dout(n1147));
  jand g0506(.dina(\in1[24] ), .dinb(n1147), .dout(n1148));
  jor  g0507(.dina(n1148), .dinb(n1146), .dout(n1149));
  jor  g0508(.dina(n1149), .dinb(n994), .dout(n1150));
  jnot g0509(.din(\in1[24] ), .dout(n1151));
  jand g0510(.dina(n1151), .dinb(\in0[24] ), .dout(n1152));
  jnot g0511(.din(\in1[25] ), .dout(n1153));
  jand g0512(.dina(n1153), .dinb(\in0[25] ), .dout(n1154));
  jor  g0513(.dina(n1154), .dinb(n1152), .dout(n1155));
  jnot g0514(.din(n1155), .dout(n1156));
  jand g0515(.dina(n1156), .dinb(n1150), .dout(n1157));
  jnot g0516(.din(\in0[26] ), .dout(n1158));
  jand g0517(.dina(\in1[26] ), .dinb(n1158), .dout(n1159));
  jnot g0518(.din(\in0[25] ), .dout(n1160));
  jand g0519(.dina(\in1[25] ), .dinb(n1160), .dout(n1161));
  jor  g0520(.dina(n1161), .dinb(n1159), .dout(n1162));
  jor  g0521(.dina(n1162), .dinb(n1157), .dout(n1163));
  jand g0522(.dina(n1163), .dinb(n992), .dout(n1164));
  jor  g0523(.dina(n1164), .dinb(n989), .dout(n1165));
  jand g0524(.dina(n1165), .dinb(n987), .dout(n1166));
  jor  g0525(.dina(n1166), .dinb(n984), .dout(n1167));
  jand g0526(.dina(n1167), .dinb(n982), .dout(n1168));
  jor  g0527(.dina(n1168), .dinb(n979), .dout(n1169));
  jand g0528(.dina(n1169), .dinb(n977), .dout(n1170));
  jor  g0529(.dina(n1170), .dinb(n974), .dout(n1171));
  jnot g0530(.din(\in1[31] ), .dout(n1172));
  jand g0531(.dina(n1172), .dinb(\in0[31] ), .dout(n1173));
  jnot g0532(.din(\in1[30] ), .dout(n1174));
  jand g0533(.dina(n1174), .dinb(\in0[30] ), .dout(n1175));
  jor  g0534(.dina(n1175), .dinb(n1173), .dout(n1176));
  jnot g0535(.din(n1176), .dout(n1177));
  jand g0536(.dina(n1177), .dinb(n1171), .dout(n1178));
  jnot g0537(.din(\in0[31] ), .dout(n1179));
  jand g0538(.dina(\in1[31] ), .dinb(n1179), .dout(n1180));
  jnot g0539(.din(\in0[32] ), .dout(n1181));
  jand g0540(.dina(\in1[32] ), .dinb(n1181), .dout(n1182));
  jor  g0541(.dina(n1182), .dinb(n1180), .dout(n1183));
  jor  g0542(.dina(n1183), .dinb(n947), .dout(n1184));
  jor  g0543(.dina(n1184), .dinb(n969), .dout(n1185));
  jor  g0544(.dina(n1185), .dinb(n1178), .dout(n1186));
  jnot g0545(.din(n967), .dout(n1187));
  jnot g0546(.din(\in1[37] ), .dout(n1188));
  jand g0547(.dina(n1188), .dinb(\in0[37] ), .dout(n1189));
  jnot g0548(.din(\in1[36] ), .dout(n1190));
  jand g0549(.dina(n1190), .dinb(\in0[36] ), .dout(n1191));
  jor  g0550(.dina(n1191), .dinb(n1189), .dout(n1192));
  jand g0551(.dina(n1192), .dinb(n1187), .dout(n1193));
  jnot g0552(.din(n968), .dout(n1194));
  jnot g0553(.din(\in1[35] ), .dout(n1195));
  jand g0554(.dina(n1195), .dinb(\in0[35] ), .dout(n1196));
  jand g0555(.dina(n1196), .dinb(n1194), .dout(n1197));
  jnot g0556(.din(\in1[39] ), .dout(n1198));
  jand g0557(.dina(n1198), .dinb(\in0[39] ), .dout(n1199));
  jnot g0558(.din(n963), .dout(n1200));
  jnot g0559(.din(\in1[38] ), .dout(n1201));
  jand g0560(.dina(n1201), .dinb(\in0[38] ), .dout(n1202));
  jand g0561(.dina(n1202), .dinb(n1200), .dout(n1203));
  jor  g0562(.dina(n1203), .dinb(n1199), .dout(n1204));
  jor  g0563(.dina(n1204), .dinb(n1197), .dout(n1205));
  jor  g0564(.dina(n1205), .dinb(n1193), .dout(n1206));
  jnot g0565(.din(n1206), .dout(n1207));
  jand g0566(.dina(n1207), .dinb(n1186), .dout(n1208));
  jand g0567(.dina(n1208), .dinb(n972), .dout(n1209));
  jnot g0568(.din(\in0[40] ), .dout(n1210));
  jand g0569(.dina(\in1[40] ), .dinb(n1210), .dout(n1211));
  jor  g0570(.dina(n1211), .dinb(n925), .dout(n1212));
  jor  g0571(.dina(n1212), .dinb(n932), .dout(n1213));
  jor  g0572(.dina(n1213), .dinb(n1209), .dout(n1214));
  jnot g0573(.din(n918), .dout(n1215));
  jnot g0574(.din(\in1[45] ), .dout(n1216));
  jand g0575(.dina(n1216), .dinb(\in0[45] ), .dout(n1217));
  jnot g0576(.din(\in1[44] ), .dout(n1218));
  jand g0577(.dina(n1218), .dinb(\in0[44] ), .dout(n1219));
  jor  g0578(.dina(n1219), .dinb(n1217), .dout(n1220));
  jand g0579(.dina(n1220), .dinb(n1215), .dout(n1221));
  jnot g0580(.din(n912), .dout(n1222));
  jnot g0581(.din(\in1[47] ), .dout(n1223));
  jand g0582(.dina(n1223), .dinb(\in0[47] ), .dout(n1224));
  jnot g0583(.din(\in1[46] ), .dout(n1225));
  jand g0584(.dina(n1225), .dinb(\in0[46] ), .dout(n1226));
  jor  g0585(.dina(n1226), .dinb(n1224), .dout(n1227));
  jand g0586(.dina(n1227), .dinb(n1222), .dout(n1228));
  jor  g0587(.dina(n1228), .dinb(n1221), .dout(n1229));
  jnot g0588(.din(n1229), .dout(n1230));
  jor  g0589(.dina(n919), .dinb(\in1[43] ), .dout(n1231));
  jor  g0590(.dina(n1231), .dinb(n922), .dout(n1232));
  jand g0591(.dina(n1232), .dinb(n1230), .dout(n1233));
  jand g0592(.dina(n1233), .dinb(n1214), .dout(n1234));
  jand g0593(.dina(n1234), .dinb(n940), .dout(n1235));
  jnot g0594(.din(\in0[48] ), .dout(n1236));
  jand g0595(.dina(\in1[48] ), .dinb(n1236), .dout(n1237));
  jnot g0596(.din(n1237), .dout(n1238));
  jnot g0597(.din(\in0[49] ), .dout(n1239));
  jand g0598(.dina(\in1[49] ), .dinb(n1239), .dout(n1240));
  jnot g0599(.din(n1240), .dout(n1241));
  jnot g0600(.din(\in0[50] ), .dout(n1242));
  jand g0601(.dina(\in1[50] ), .dinb(n1242), .dout(n1243));
  jnot g0602(.din(\in0[51] ), .dout(n1244));
  jand g0603(.dina(\in1[51] ), .dinb(n1244), .dout(n1245));
  jor  g0604(.dina(n1245), .dinb(n1243), .dout(n1246));
  jor  g0605(.dina(n1246), .dinb(n904), .dout(n1247));
  jnot g0606(.din(n1247), .dout(n1248));
  jand g0607(.dina(n1248), .dinb(n1241), .dout(n1249));
  jand g0608(.dina(n1249), .dinb(n1238), .dout(n1250));
  jnot g0609(.din(n1250), .dout(n1251));
  jor  g0610(.dina(n1251), .dinb(n1235), .dout(n1252));
  jnot g0611(.din(\in1[49] ), .dout(n1253));
  jand g0612(.dina(n1253), .dinb(\in0[49] ), .dout(n1254));
  jnot g0613(.din(\in1[50] ), .dout(n1255));
  jand g0614(.dina(n1255), .dinb(\in0[50] ), .dout(n1256));
  jor  g0615(.dina(n1256), .dinb(n1254), .dout(n1257));
  jnot g0616(.din(\in1[48] ), .dout(n1258));
  jand g0617(.dina(n1258), .dinb(\in0[48] ), .dout(n1259));
  jand g0618(.dina(n1259), .dinb(n1241), .dout(n1260));
  jor  g0619(.dina(n1260), .dinb(n1257), .dout(n1261));
  jand g0620(.dina(n1261), .dinb(n1248), .dout(n1262));
  jnot g0621(.din(\in1[55] ), .dout(n1263));
  jand g0622(.dina(n1263), .dinb(\in0[55] ), .dout(n1264));
  jnot g0623(.din(n900), .dout(n1265));
  jnot g0624(.din(n895), .dout(n1266));
  jnot g0625(.din(\in1[52] ), .dout(n1267));
  jand g0626(.dina(n1267), .dinb(\in0[52] ), .dout(n1268));
  jand g0627(.dina(n1268), .dinb(n1266), .dout(n1269));
  jnot g0628(.din(\in1[54] ), .dout(n1270));
  jand g0629(.dina(n1270), .dinb(\in0[54] ), .dout(n1271));
  jnot g0630(.din(\in1[53] ), .dout(n1272));
  jand g0631(.dina(n1272), .dinb(\in0[53] ), .dout(n1273));
  jor  g0632(.dina(n1273), .dinb(n1271), .dout(n1274));
  jor  g0633(.dina(n1274), .dinb(n1269), .dout(n1275));
  jand g0634(.dina(n1275), .dinb(n1265), .dout(n1276));
  jor  g0635(.dina(n1276), .dinb(n1264), .dout(n1277));
  jor  g0636(.dina(n1277), .dinb(n1262), .dout(n1278));
  jnot g0637(.din(n1278), .dout(n1279));
  jand g0638(.dina(n1279), .dinb(n1252), .dout(n1280));
  jand g0639(.dina(n1280), .dinb(n908), .dout(n1281));
  jnot g0640(.din(\in0[56] ), .dout(n1282));
  jand g0641(.dina(\in1[56] ), .dinb(n1282), .dout(n1283));
  jnot g0642(.din(n1283), .dout(n1284));
  jnot g0643(.din(\in0[57] ), .dout(n1285));
  jand g0644(.dina(\in1[57] ), .dinb(n1285), .dout(n1286));
  jnot g0645(.din(n1286), .dout(n1287));
  jnot g0646(.din(\in0[58] ), .dout(n1288));
  jand g0647(.dina(\in1[58] ), .dinb(n1288), .dout(n1289));
  jnot g0648(.din(\in0[59] ), .dout(n1290));
  jand g0649(.dina(\in1[59] ), .dinb(n1290), .dout(n1291));
  jor  g0650(.dina(n1291), .dinb(n1289), .dout(n1292));
  jor  g0651(.dina(n1292), .dinb(n888), .dout(n1293));
  jnot g0652(.din(n1293), .dout(n1294));
  jand g0653(.dina(n1294), .dinb(n1287), .dout(n1295));
  jand g0654(.dina(n1295), .dinb(n1284), .dout(n1296));
  jnot g0655(.din(n1296), .dout(n1297));
  jor  g0656(.dina(n1297), .dinb(n1281), .dout(n1298));
  jnot g0657(.din(\in1[57] ), .dout(n1299));
  jand g0658(.dina(n1299), .dinb(\in0[57] ), .dout(n1300));
  jnot g0659(.din(\in1[58] ), .dout(n1301));
  jand g0660(.dina(n1301), .dinb(\in0[58] ), .dout(n1302));
  jor  g0661(.dina(n1302), .dinb(n1300), .dout(n1303));
  jnot g0662(.din(\in1[56] ), .dout(n1304));
  jand g0663(.dina(n1304), .dinb(\in0[56] ), .dout(n1305));
  jand g0664(.dina(n1305), .dinb(n1287), .dout(n1306));
  jor  g0665(.dina(n1306), .dinb(n1303), .dout(n1307));
  jand g0666(.dina(n1307), .dinb(n1294), .dout(n1308));
  jnot g0667(.din(n887), .dout(n1309));
  jnot g0668(.din(\in1[61] ), .dout(n1310));
  jand g0669(.dina(n1310), .dinb(\in0[61] ), .dout(n1311));
  jnot g0670(.din(\in1[60] ), .dout(n1312));
  jand g0671(.dina(n1312), .dinb(\in0[60] ), .dout(n1313));
  jor  g0672(.dina(n1313), .dinb(n1311), .dout(n1314));
  jand g0673(.dina(n1314), .dinb(n1309), .dout(n1315));
  jnot g0674(.din(n881), .dout(n1316));
  jnot g0675(.din(\in1[63] ), .dout(n1317));
  jand g0676(.dina(n1317), .dinb(\in0[63] ), .dout(n1318));
  jnot g0677(.din(\in1[62] ), .dout(n1319));
  jand g0678(.dina(n1319), .dinb(\in0[62] ), .dout(n1320));
  jor  g0679(.dina(n1320), .dinb(n1318), .dout(n1321));
  jand g0680(.dina(n1321), .dinb(n1316), .dout(n1322));
  jor  g0681(.dina(n1322), .dinb(n1315), .dout(n1323));
  jor  g0682(.dina(n1323), .dinb(n1308), .dout(n1324));
  jnot g0683(.din(n1324), .dout(n1325));
  jand g0684(.dina(n1325), .dinb(n1298), .dout(n1326));
  jand g0685(.dina(n1326), .dinb(n892), .dout(n1327));
  jnot g0686(.din(\in0[64] ), .dout(n1328));
  jand g0687(.dina(\in1[64] ), .dinb(n1328), .dout(n1329));
  jor  g0688(.dina(n1329), .dinb(n865), .dout(n1330));
  jor  g0689(.dina(n1330), .dinb(n1327), .dout(n1331));
  jand g0690(.dina(n1331), .dinb(n876), .dout(n1332));
  jnot g0691(.din(\in0[67] ), .dout(n1333));
  jand g0692(.dina(\in1[67] ), .dinb(n1333), .dout(n1334));
  jnot g0693(.din(\in0[66] ), .dout(n1335));
  jand g0694(.dina(\in1[66] ), .dinb(n1335), .dout(n1336));
  jor  g0695(.dina(n1336), .dinb(n1334), .dout(n1337));
  jor  g0696(.dina(n1337), .dinb(n1332), .dout(n1338));
  jand g0697(.dina(n1338), .dinb(n863), .dout(n1339));
  jnot g0698(.din(\in0[68] ), .dout(n1340));
  jand g0699(.dina(\in1[68] ), .dinb(n1340), .dout(n1341));
  jor  g0700(.dina(n1341), .dinb(n844), .dout(n1342));
  jor  g0701(.dina(n1342), .dinb(n1339), .dout(n1343));
  jand g0702(.dina(n1343), .dinb(n860), .dout(n1344));
  jnot g0703(.din(\in0[75] ), .dout(n1345));
  jand g0704(.dina(\in1[75] ), .dinb(n1345), .dout(n1346));
  jnot g0705(.din(\in0[74] ), .dout(n1347));
  jand g0706(.dina(\in1[74] ), .dinb(n1347), .dout(n1348));
  jor  g0707(.dina(n1348), .dinb(n1346), .dout(n1349));
  jor  g0708(.dina(n1349), .dinb(n1344), .dout(n1350));
  jor  g0709(.dina(n1350), .dinb(n836), .dout(n1351));
  jnot g0710(.din(n1349), .dout(n1352));
  jnot g0711(.din(\in1[73] ), .dout(n1353));
  jand g0712(.dina(n1353), .dinb(\in0[73] ), .dout(n1354));
  jnot g0713(.din(\in1[74] ), .dout(n1355));
  jand g0714(.dina(n1355), .dinb(\in0[74] ), .dout(n1356));
  jor  g0715(.dina(n1356), .dinb(n1354), .dout(n1357));
  jnot g0716(.din(n835), .dout(n1358));
  jnot g0717(.din(\in1[72] ), .dout(n1359));
  jand g0718(.dina(n1359), .dinb(\in0[72] ), .dout(n1360));
  jand g0719(.dina(n1360), .dinb(n1358), .dout(n1361));
  jor  g0720(.dina(n1361), .dinb(n1357), .dout(n1362));
  jand g0721(.dina(n1362), .dinb(n1352), .dout(n1363));
  jnot g0722(.din(n1363), .dout(n1364));
  jand g0723(.dina(n1364), .dinb(n1351), .dout(n1365));
  jand g0724(.dina(n1365), .dinb(n831), .dout(n1366));
  jnot g0725(.din(\in0[76] ), .dout(n1367));
  jand g0726(.dina(\in1[76] ), .dinb(n1367), .dout(n1368));
  jor  g0727(.dina(n1368), .dinb(n812), .dout(n1369));
  jor  g0728(.dina(n1369), .dinb(n1366), .dout(n1370));
  jand g0729(.dina(n1370), .dinb(n828), .dout(n1371));
  jnot g0730(.din(\in0[83] ), .dout(n1372));
  jand g0731(.dina(\in1[83] ), .dinb(n1372), .dout(n1373));
  jnot g0732(.din(\in0[82] ), .dout(n1374));
  jand g0733(.dina(\in1[82] ), .dinb(n1374), .dout(n1375));
  jor  g0734(.dina(n1375), .dinb(n1373), .dout(n1376));
  jor  g0735(.dina(n1376), .dinb(n1371), .dout(n1377));
  jor  g0736(.dina(n1377), .dinb(n804), .dout(n1378));
  jnot g0737(.din(n1376), .dout(n1379));
  jnot g0738(.din(\in1[81] ), .dout(n1380));
  jand g0739(.dina(n1380), .dinb(\in0[81] ), .dout(n1381));
  jnot g0740(.din(\in1[82] ), .dout(n1382));
  jand g0741(.dina(n1382), .dinb(\in0[82] ), .dout(n1383));
  jor  g0742(.dina(n1383), .dinb(n1381), .dout(n1384));
  jnot g0743(.din(n801), .dout(n1385));
  jnot g0744(.din(\in1[80] ), .dout(n1386));
  jand g0745(.dina(n1386), .dinb(\in0[80] ), .dout(n1387));
  jand g0746(.dina(n1387), .dinb(n1385), .dout(n1388));
  jor  g0747(.dina(n1388), .dinb(n1384), .dout(n1389));
  jand g0748(.dina(n1389), .dinb(n1379), .dout(n1390));
  jnot g0749(.din(n1390), .dout(n1391));
  jand g0750(.dina(n1391), .dinb(n1378), .dout(n1392));
  jand g0751(.dina(n1392), .dinb(n799), .dout(n1393));
  jnot g0752(.din(\in0[84] ), .dout(n1394));
  jand g0753(.dina(\in1[84] ), .dinb(n1394), .dout(n1395));
  jor  g0754(.dina(n1395), .dinb(n780), .dout(n1396));
  jor  g0755(.dina(n1396), .dinb(n1393), .dout(n1397));
  jand g0756(.dina(n1397), .dinb(n796), .dout(n1398));
  jnot g0757(.din(\in0[91] ), .dout(n1399));
  jand g0758(.dina(\in1[91] ), .dinb(n1399), .dout(n1400));
  jnot g0759(.din(\in0[90] ), .dout(n1401));
  jand g0760(.dina(\in1[90] ), .dinb(n1401), .dout(n1402));
  jor  g0761(.dina(n1402), .dinb(n1400), .dout(n1403));
  jnot g0762(.din(\in0[88] ), .dout(n1404));
  jand g0763(.dina(\in1[88] ), .dinb(n1404), .dout(n1405));
  jnot g0764(.din(\in0[89] ), .dout(n1406));
  jand g0765(.dina(\in1[89] ), .dinb(n1406), .dout(n1407));
  jor  g0766(.dina(n1407), .dinb(n1405), .dout(n1408));
  jor  g0767(.dina(n1408), .dinb(n1403), .dout(n1409));
  jor  g0768(.dina(n1409), .dinb(n1398), .dout(n1410));
  jnot g0769(.din(n1403), .dout(n1411));
  jnot g0770(.din(\in1[89] ), .dout(n1412));
  jand g0771(.dina(n1412), .dinb(\in0[89] ), .dout(n1413));
  jnot g0772(.din(\in1[90] ), .dout(n1414));
  jand g0773(.dina(n1414), .dinb(\in0[90] ), .dout(n1415));
  jor  g0774(.dina(n1415), .dinb(n1413), .dout(n1416));
  jnot g0775(.din(n1407), .dout(n1417));
  jnot g0776(.din(\in1[88] ), .dout(n1418));
  jand g0777(.dina(n1418), .dinb(\in0[88] ), .dout(n1419));
  jand g0778(.dina(n1419), .dinb(n1417), .dout(n1420));
  jor  g0779(.dina(n1420), .dinb(n1416), .dout(n1421));
  jand g0780(.dina(n1421), .dinb(n1411), .dout(n1422));
  jnot g0781(.din(n1422), .dout(n1423));
  jand g0782(.dina(n1423), .dinb(n1410), .dout(n1424));
  jand g0783(.dina(n1424), .dinb(n772), .dout(n1425));
  jnot g0784(.din(\in0[92] ), .dout(n1426));
  jand g0785(.dina(\in1[92] ), .dinb(n1426), .dout(n1427));
  jor  g0786(.dina(n1427), .dinb(n753), .dout(n1428));
  jor  g0787(.dina(n1428), .dinb(n1425), .dout(n1429));
  jand g0788(.dina(n1429), .dinb(n769), .dout(n1430));
  jnot g0789(.din(\in0[99] ), .dout(n1431));
  jand g0790(.dina(\in1[99] ), .dinb(n1431), .dout(n1432));
  jnot g0791(.din(\in0[98] ), .dout(n1433));
  jand g0792(.dina(\in1[98] ), .dinb(n1433), .dout(n1434));
  jor  g0793(.dina(n1434), .dinb(n1432), .dout(n1435));
  jor  g0794(.dina(n1435), .dinb(n1430), .dout(n1436));
  jor  g0795(.dina(n1436), .dinb(n745), .dout(n1437));
  jnot g0796(.din(n1435), .dout(n1438));
  jnot g0797(.din(\in1[97] ), .dout(n1439));
  jand g0798(.dina(n1439), .dinb(\in0[97] ), .dout(n1440));
  jnot g0799(.din(\in1[98] ), .dout(n1441));
  jand g0800(.dina(n1441), .dinb(\in0[98] ), .dout(n1442));
  jor  g0801(.dina(n1442), .dinb(n1440), .dout(n1443));
  jnot g0802(.din(n742), .dout(n1444));
  jnot g0803(.din(\in1[96] ), .dout(n1445));
  jand g0804(.dina(n1445), .dinb(\in0[96] ), .dout(n1446));
  jand g0805(.dina(n1446), .dinb(n1444), .dout(n1447));
  jor  g0806(.dina(n1447), .dinb(n1443), .dout(n1448));
  jand g0807(.dina(n1448), .dinb(n1438), .dout(n1449));
  jnot g0808(.din(n1449), .dout(n1450));
  jand g0809(.dina(n1450), .dinb(n1437), .dout(n1451));
  jand g0810(.dina(n1451), .dinb(n740), .dout(n1452));
  jnot g0811(.din(\in0[100] ), .dout(n1453));
  jand g0812(.dina(\in1[100] ), .dinb(n1453), .dout(n1454));
  jor  g0813(.dina(n1454), .dinb(n721), .dout(n1455));
  jor  g0814(.dina(n1455), .dinb(n1452), .dout(n1456));
  jand g0815(.dina(n1456), .dinb(n737), .dout(n1457));
  jnot g0816(.din(\in0[107] ), .dout(n1458));
  jand g0817(.dina(\in1[107] ), .dinb(n1458), .dout(n1459));
  jnot g0818(.din(\in0[106] ), .dout(n1460));
  jand g0819(.dina(\in1[106] ), .dinb(n1460), .dout(n1461));
  jor  g0820(.dina(n1461), .dinb(n1459), .dout(n1462));
  jor  g0821(.dina(n1462), .dinb(n1457), .dout(n1463));
  jor  g0822(.dina(n1463), .dinb(n713), .dout(n1464));
  jnot g0823(.din(n1462), .dout(n1465));
  jnot g0824(.din(\in1[105] ), .dout(n1466));
  jand g0825(.dina(n1466), .dinb(\in0[105] ), .dout(n1467));
  jnot g0826(.din(\in1[106] ), .dout(n1468));
  jand g0827(.dina(n1468), .dinb(\in0[106] ), .dout(n1469));
  jor  g0828(.dina(n1469), .dinb(n1467), .dout(n1470));
  jnot g0829(.din(n712), .dout(n1471));
  jnot g0830(.din(\in1[104] ), .dout(n1472));
  jand g0831(.dina(n1472), .dinb(\in0[104] ), .dout(n1473));
  jand g0832(.dina(n1473), .dinb(n1471), .dout(n1474));
  jor  g0833(.dina(n1474), .dinb(n1470), .dout(n1475));
  jand g0834(.dina(n1475), .dinb(n1465), .dout(n1476));
  jnot g0835(.din(n1476), .dout(n1477));
  jand g0836(.dina(n1477), .dinb(n1464), .dout(n1478));
  jand g0837(.dina(n1478), .dinb(n708), .dout(n1479));
  jnot g0838(.din(\in0[108] ), .dout(n1480));
  jand g0839(.dina(\in1[108] ), .dinb(n1480), .dout(n1481));
  jor  g0840(.dina(n1481), .dinb(n689), .dout(n1482));
  jor  g0841(.dina(n1482), .dinb(n1479), .dout(n1483));
  jand g0842(.dina(n1483), .dinb(n705), .dout(n1484));
  jnot g0843(.din(\in0[115] ), .dout(n1485));
  jand g0844(.dina(\in1[115] ), .dinb(n1485), .dout(n1486));
  jnot g0845(.din(\in0[114] ), .dout(n1487));
  jand g0846(.dina(\in1[114] ), .dinb(n1487), .dout(n1488));
  jor  g0847(.dina(n1488), .dinb(n1486), .dout(n1489));
  jor  g0848(.dina(n1489), .dinb(n1484), .dout(n1490));
  jor  g0849(.dina(n1490), .dinb(n681), .dout(n1491));
  jnot g0850(.din(n1489), .dout(n1492));
  jnot g0851(.din(\in1[113] ), .dout(n1493));
  jand g0852(.dina(n1493), .dinb(\in0[113] ), .dout(n1494));
  jnot g0853(.din(\in1[114] ), .dout(n1495));
  jand g0854(.dina(n1495), .dinb(\in0[114] ), .dout(n1496));
  jor  g0855(.dina(n1496), .dinb(n1494), .dout(n1497));
  jnot g0856(.din(n678), .dout(n1498));
  jnot g0857(.din(\in1[112] ), .dout(n1499));
  jand g0858(.dina(n1499), .dinb(\in0[112] ), .dout(n1500));
  jand g0859(.dina(n1500), .dinb(n1498), .dout(n1501));
  jor  g0860(.dina(n1501), .dinb(n1497), .dout(n1502));
  jand g0861(.dina(n1502), .dinb(n1492), .dout(n1503));
  jnot g0862(.din(n1503), .dout(n1504));
  jand g0863(.dina(n1504), .dinb(n1491), .dout(n1505));
  jand g0864(.dina(n1505), .dinb(n676), .dout(n1506));
  jnot g0865(.din(\in0[116] ), .dout(n1507));
  jand g0866(.dina(\in1[116] ), .dinb(n1507), .dout(n1508));
  jor  g0867(.dina(n1508), .dinb(n657), .dout(n1509));
  jor  g0868(.dina(n1509), .dinb(n1506), .dout(n1510));
  jand g0869(.dina(n1510), .dinb(n673), .dout(n1511));
  jnot g0870(.din(\in0[123] ), .dout(n1512));
  jand g0871(.dina(\in1[123] ), .dinb(n1512), .dout(n1513));
  jnot g0872(.din(\in0[122] ), .dout(n1514));
  jand g0873(.dina(\in1[122] ), .dinb(n1514), .dout(n1515));
  jor  g0874(.dina(n1515), .dinb(n1513), .dout(n1516));
  jor  g0875(.dina(n1516), .dinb(n1511), .dout(n1517));
  jor  g0876(.dina(n1517), .dinb(n649), .dout(n1518));
  jnot g0877(.din(n1516), .dout(n1519));
  jnot g0878(.din(\in1[121] ), .dout(n1520));
  jand g0879(.dina(n1520), .dinb(\in0[121] ), .dout(n1521));
  jnot g0880(.din(\in1[122] ), .dout(n1522));
  jand g0881(.dina(n1522), .dinb(\in0[122] ), .dout(n1523));
  jor  g0882(.dina(n1523), .dinb(n1521), .dout(n1524));
  jnot g0883(.din(n648), .dout(n1525));
  jnot g0884(.din(\in1[120] ), .dout(n1526));
  jand g0885(.dina(n1526), .dinb(\in0[120] ), .dout(n1527));
  jand g0886(.dina(n1527), .dinb(n1525), .dout(n1528));
  jor  g0887(.dina(n1528), .dinb(n1524), .dout(n1529));
  jand g0888(.dina(n1529), .dinb(n1519), .dout(n1530));
  jnot g0889(.din(n1530), .dout(n1531));
  jand g0890(.dina(n1531), .dinb(n1518), .dout(n1532));
  jand g0891(.dina(n1532), .dinb(n644), .dout(n1533));
  jnot g0892(.din(\in0[126] ), .dout(n1534));
  jand g0893(.dina(\in1[126] ), .dinb(n1534), .dout(n1535));
  jnot g0894(.din(\in0[125] ), .dout(n1536));
  jand g0895(.dina(\in1[125] ), .dinb(n1536), .dout(n1537));
  jor  g0896(.dina(n1537), .dinb(n1535), .dout(n1538));
  jnot g0897(.din(\in0[124] ), .dout(n1539));
  jand g0898(.dina(\in1[124] ), .dinb(n1539), .dout(n1540));
  jnot g0899(.din(\in1[127] ), .dout(n1541));
  jand g0900(.dina(n1541), .dinb(\in0[127] ), .dout(n1542));
  jor  g0901(.dina(n1542), .dinb(n1540), .dout(n1543));
  jor  g0902(.dina(n1543), .dinb(n1538), .dout(n1544));
  jor  g0903(.dina(n1544), .dinb(n1533), .dout(n1545));
  jnot g0904(.din(n1542), .dout(n1546));
  jnot g0905(.din(n1538), .dout(n1547));
  jnot g0906(.din(\in1[124] ), .dout(n1548));
  jand g0907(.dina(n1548), .dinb(\in0[124] ), .dout(n1549));
  jnot g0908(.din(\in1[125] ), .dout(n1550));
  jand g0909(.dina(n1550), .dinb(\in0[125] ), .dout(n1551));
  jor  g0910(.dina(n1551), .dinb(n1549), .dout(n1552));
  jand g0911(.dina(n1552), .dinb(n1547), .dout(n1553));
  jnot g0912(.din(\in1[126] ), .dout(n1554));
  jand g0913(.dina(n1554), .dinb(\in0[126] ), .dout(n1555));
  jnot g0914(.din(\in0[127] ), .dout(n1556));
  jand g0915(.dina(\in1[127] ), .dinb(n1556), .dout(n1557));
  jor  g0916(.dina(n1557), .dinb(n1555), .dout(n1558));
  jor  g0917(.dina(n1558), .dinb(n1553), .dout(n1559));
  jand g0918(.dina(n1559), .dinb(n1546), .dout(n1560));
  jnot g0919(.din(n1560), .dout(n1561));
  jand g0920(.dina(n1561), .dinb(n1545), .dout(n1562));
  jor  g0921(.dina(n1562), .dinb(\in0[0] ), .dout(n1563));
  jnot g0922(.din(n649), .dout(n1564));
  jnot g0923(.din(n681), .dout(n1565));
  jnot g0924(.din(n713), .dout(n1566));
  jnot g0925(.din(n745), .dout(n1567));
  jnot g0926(.din(n804), .dout(n1568));
  jnot g0927(.din(n836), .dout(n1569));
  jnot g0928(.din(n974), .dout(n1570));
  jnot g0929(.din(n979), .dout(n1571));
  jnot g0930(.din(n984), .dout(n1572));
  jnot g0931(.din(n989), .dout(n1573));
  jnot g0932(.din(n994), .dout(n1574));
  jnot g0933(.din(n996), .dout(n1575));
  jnot g0934(.din(n1001), .dout(n1576));
  jnot g0935(.din(n1006), .dout(n1577));
  jnot g0936(.din(n1011), .dout(n1578));
  jnot g0937(.din(n1016), .dout(n1579));
  jnot g0938(.din(n1018), .dout(n1580));
  jnot g0939(.din(n1023), .dout(n1581));
  jnot g0940(.din(n1028), .dout(n1582));
  jnot g0941(.din(n1033), .dout(n1583));
  jnot g0942(.din(n1038), .dout(n1584));
  jnot g0943(.din(n1040), .dout(n1585));
  jnot g0944(.din(\in1[1] ), .dout(n1586));
  jand g0945(.dina(n1586), .dinb(\in0[1] ), .dout(n1587));
  jnot g0946(.din(\in1[0] ), .dout(n1588));
  jand g0947(.dina(n1588), .dinb(\in0[0] ), .dout(n1589));
  jor  g0948(.dina(n1589), .dinb(n1587), .dout(n1590));
  jor  g0949(.dina(n1041), .dinb(\in0[2] ), .dout(n1591));
  jor  g0950(.dina(n1586), .dinb(\in0[1] ), .dout(n1592));
  jand g0951(.dina(n1592), .dinb(n1591), .dout(n1593));
  jand g0952(.dina(n1593), .dinb(n1590), .dout(n1594));
  jor  g0953(.dina(n1055), .dinb(n1594), .dout(n1595));
  jor  g0954(.dina(n1595), .dinb(n1042), .dout(n1596));
  jnot g0955(.din(n1060), .dout(n1597));
  jand g0956(.dina(n1597), .dinb(n1596), .dout(n1598));
  jand g0957(.dina(n1598), .dinb(n1585), .dout(n1599));
  jor  g0958(.dina(n1067), .dinb(n1599), .dout(n1600));
  jnot g0959(.din(n1074), .dout(n1601));
  jand g0960(.dina(n1601), .dinb(n1600), .dout(n1602));
  jor  g0961(.dina(n1080), .dinb(n1602), .dout(n1603));
  jnot g0962(.din(n1084), .dout(n1604));
  jand g0963(.dina(n1604), .dinb(n1603), .dout(n1605));
  jand g0964(.dina(n1605), .dinb(n1584), .dout(n1606));
  jor  g0965(.dina(n1091), .dinb(n1606), .dout(n1607));
  jnot g0966(.din(n1098), .dout(n1608));
  jand g0967(.dina(n1608), .dinb(n1607), .dout(n1609));
  jor  g0968(.dina(n1609), .dinb(n1035), .dout(n1610));
  jand g0969(.dina(n1610), .dinb(n1583), .dout(n1611));
  jor  g0970(.dina(n1611), .dinb(n1030), .dout(n1612));
  jand g0971(.dina(n1612), .dinb(n1582), .dout(n1613));
  jor  g0972(.dina(n1613), .dinb(n1025), .dout(n1614));
  jand g0973(.dina(n1614), .dinb(n1581), .dout(n1615));
  jor  g0974(.dina(n1615), .dinb(n1020), .dout(n1616));
  jand g0975(.dina(n1616), .dinb(n1580), .dout(n1617));
  jor  g0976(.dina(n1112), .dinb(n1617), .dout(n1618));
  jnot g0977(.din(n1116), .dout(n1619));
  jand g0978(.dina(n1619), .dinb(n1618), .dout(n1620));
  jand g0979(.dina(n1620), .dinb(n1579), .dout(n1621));
  jor  g0980(.dina(n1123), .dinb(n1621), .dout(n1622));
  jnot g0981(.din(n1130), .dout(n1623));
  jand g0982(.dina(n1623), .dinb(n1622), .dout(n1624));
  jor  g0983(.dina(n1624), .dinb(n1013), .dout(n1625));
  jand g0984(.dina(n1625), .dinb(n1578), .dout(n1626));
  jor  g0985(.dina(n1626), .dinb(n1008), .dout(n1627));
  jand g0986(.dina(n1627), .dinb(n1577), .dout(n1628));
  jor  g0987(.dina(n1628), .dinb(n1003), .dout(n1629));
  jand g0988(.dina(n1629), .dinb(n1576), .dout(n1630));
  jor  g0989(.dina(n1630), .dinb(n998), .dout(n1631));
  jand g0990(.dina(n1631), .dinb(n1575), .dout(n1632));
  jor  g0991(.dina(n1144), .dinb(n1632), .dout(n1633));
  jnot g0992(.din(n1148), .dout(n1634));
  jand g0993(.dina(n1634), .dinb(n1633), .dout(n1635));
  jand g0994(.dina(n1635), .dinb(n1574), .dout(n1636));
  jor  g0995(.dina(n1155), .dinb(n1636), .dout(n1637));
  jnot g0996(.din(n1162), .dout(n1638));
  jand g0997(.dina(n1638), .dinb(n1637), .dout(n1639));
  jor  g0998(.dina(n1639), .dinb(n991), .dout(n1640));
  jand g0999(.dina(n1640), .dinb(n1573), .dout(n1641));
  jor  g1000(.dina(n1641), .dinb(n986), .dout(n1642));
  jand g1001(.dina(n1642), .dinb(n1572), .dout(n1643));
  jor  g1002(.dina(n1643), .dinb(n981), .dout(n1644));
  jand g1003(.dina(n1644), .dinb(n1571), .dout(n1645));
  jor  g1004(.dina(n1645), .dinb(n976), .dout(n1646));
  jand g1005(.dina(n1646), .dinb(n1570), .dout(n1647));
  jor  g1006(.dina(n1176), .dinb(n1647), .dout(n1648));
  jnot g1007(.din(n1185), .dout(n1649));
  jand g1008(.dina(n1649), .dinb(n1648), .dout(n1650));
  jor  g1009(.dina(n1206), .dinb(n1650), .dout(n1651));
  jor  g1010(.dina(n1651), .dinb(n971), .dout(n1652));
  jnot g1011(.din(n1213), .dout(n1653));
  jand g1012(.dina(n1653), .dinb(n1652), .dout(n1654));
  jnot g1013(.din(n1233), .dout(n1655));
  jor  g1014(.dina(n1655), .dinb(n1654), .dout(n1656));
  jor  g1015(.dina(n1656), .dinb(n939), .dout(n1657));
  jand g1016(.dina(n1250), .dinb(n1657), .dout(n1658));
  jor  g1017(.dina(n1278), .dinb(n1658), .dout(n1659));
  jor  g1018(.dina(n1659), .dinb(n907), .dout(n1660));
  jand g1019(.dina(n1296), .dinb(n1660), .dout(n1661));
  jor  g1020(.dina(n1324), .dinb(n1661), .dout(n1662));
  jor  g1021(.dina(n1662), .dinb(n891), .dout(n1663));
  jnot g1022(.din(n1330), .dout(n1664));
  jand g1023(.dina(n1664), .dinb(n1663), .dout(n1665));
  jor  g1024(.dina(n1665), .dinb(n875), .dout(n1666));
  jnot g1025(.din(n1337), .dout(n1667));
  jand g1026(.dina(n1667), .dinb(n1666), .dout(n1668));
  jor  g1027(.dina(n1668), .dinb(n862), .dout(n1669));
  jnot g1028(.din(n1342), .dout(n1670));
  jand g1029(.dina(n1670), .dinb(n1669), .dout(n1671));
  jor  g1030(.dina(n1671), .dinb(n859), .dout(n1672));
  jand g1031(.dina(n1352), .dinb(n1672), .dout(n1673));
  jand g1032(.dina(n1673), .dinb(n1569), .dout(n1674));
  jor  g1033(.dina(n1363), .dinb(n1674), .dout(n1675));
  jor  g1034(.dina(n1675), .dinb(n830), .dout(n1676));
  jnot g1035(.din(n1369), .dout(n1677));
  jand g1036(.dina(n1677), .dinb(n1676), .dout(n1678));
  jor  g1037(.dina(n1678), .dinb(n827), .dout(n1679));
  jand g1038(.dina(n1379), .dinb(n1679), .dout(n1680));
  jand g1039(.dina(n1680), .dinb(n1568), .dout(n1681));
  jor  g1040(.dina(n1390), .dinb(n1681), .dout(n1682));
  jor  g1041(.dina(n1682), .dinb(n798), .dout(n1683));
  jnot g1042(.din(n1396), .dout(n1684));
  jand g1043(.dina(n1684), .dinb(n1683), .dout(n1685));
  jor  g1044(.dina(n1685), .dinb(n795), .dout(n1686));
  jnot g1045(.din(n1409), .dout(n1687));
  jand g1046(.dina(n1687), .dinb(n1686), .dout(n1688));
  jor  g1047(.dina(n1422), .dinb(n1688), .dout(n1689));
  jor  g1048(.dina(n1689), .dinb(n771), .dout(n1690));
  jnot g1049(.din(n1428), .dout(n1691));
  jand g1050(.dina(n1691), .dinb(n1690), .dout(n1692));
  jor  g1051(.dina(n1692), .dinb(n768), .dout(n1693));
  jand g1052(.dina(n1438), .dinb(n1693), .dout(n1694));
  jand g1053(.dina(n1694), .dinb(n1567), .dout(n1695));
  jor  g1054(.dina(n1449), .dinb(n1695), .dout(n1696));
  jor  g1055(.dina(n1696), .dinb(n739), .dout(n1697));
  jnot g1056(.din(n1455), .dout(n1698));
  jand g1057(.dina(n1698), .dinb(n1697), .dout(n1699));
  jor  g1058(.dina(n1699), .dinb(n736), .dout(n1700));
  jand g1059(.dina(n1465), .dinb(n1700), .dout(n1701));
  jand g1060(.dina(n1701), .dinb(n1566), .dout(n1702));
  jor  g1061(.dina(n1476), .dinb(n1702), .dout(n1703));
  jor  g1062(.dina(n1703), .dinb(n707), .dout(n1704));
  jnot g1063(.din(n1482), .dout(n1705));
  jand g1064(.dina(n1705), .dinb(n1704), .dout(n1706));
  jor  g1065(.dina(n1706), .dinb(n704), .dout(n1707));
  jand g1066(.dina(n1492), .dinb(n1707), .dout(n1708));
  jand g1067(.dina(n1708), .dinb(n1565), .dout(n1709));
  jor  g1068(.dina(n1503), .dinb(n1709), .dout(n1710));
  jor  g1069(.dina(n1710), .dinb(n675), .dout(n1711));
  jnot g1070(.din(n1509), .dout(n1712));
  jand g1071(.dina(n1712), .dinb(n1711), .dout(n1713));
  jor  g1072(.dina(n1713), .dinb(n672), .dout(n1714));
  jand g1073(.dina(n1519), .dinb(n1714), .dout(n1715));
  jand g1074(.dina(n1715), .dinb(n1564), .dout(n1716));
  jor  g1075(.dina(n1530), .dinb(n1716), .dout(n1717));
  jor  g1076(.dina(n1717), .dinb(n643), .dout(n1718));
  jnot g1077(.din(n1544), .dout(n1719));
  jand g1078(.dina(n1719), .dinb(n1718), .dout(n1720));
  jor  g1079(.dina(n1560), .dinb(n1720), .dout(n1721));
  jor  g1080(.dina(n1721), .dinb(\in1[0] ), .dout(n1722));
  jand g1081(.dina(n1722), .dinb(n1563), .dout(n1723));
  jnot g1082(.din(\in2[126] ), .dout(n1724));
  jand g1083(.dina(\in3[126] ), .dinb(n1724), .dout(n1725));
  jnot g1084(.din(\in2[125] ), .dout(n1726));
  jand g1085(.dina(\in3[125] ), .dinb(n1726), .dout(n1727));
  jor  g1086(.dina(n1727), .dinb(n1725), .dout(n1728));
  jnot g1087(.din(n1728), .dout(n1729));
  jnot g1088(.din(\in3[124] ), .dout(n1730));
  jand g1089(.dina(n1730), .dinb(\in2[124] ), .dout(n1731));
  jnot g1090(.din(\in3[125] ), .dout(n1732));
  jand g1091(.dina(n1732), .dinb(\in2[125] ), .dout(n1733));
  jor  g1092(.dina(n1733), .dinb(n1731), .dout(n1734));
  jand g1093(.dina(n1734), .dinb(n1729), .dout(n1735));
  jnot g1094(.din(\in3[126] ), .dout(n1736));
  jand g1095(.dina(n1736), .dinb(\in2[126] ), .dout(n1737));
  jor  g1096(.dina(n1737), .dinb(n1735), .dout(n1738));
  jnot g1097(.din(n1738), .dout(n1739));
  jnot g1098(.din(\in3[123] ), .dout(n1740));
  jand g1099(.dina(n1740), .dinb(\in2[123] ), .dout(n1741));
  jnot g1100(.din(n1741), .dout(n1742));
  jnot g1101(.din(\in2[118] ), .dout(n1743));
  jand g1102(.dina(\in3[118] ), .dinb(n1743), .dout(n1744));
  jnot g1103(.din(\in2[119] ), .dout(n1745));
  jand g1104(.dina(\in3[119] ), .dinb(n1745), .dout(n1746));
  jnot g1105(.din(\in2[117] ), .dout(n1747));
  jand g1106(.dina(\in3[117] ), .dinb(n1747), .dout(n1748));
  jor  g1107(.dina(n1748), .dinb(n1746), .dout(n1749));
  jor  g1108(.dina(n1749), .dinb(n1744), .dout(n1750));
  jnot g1109(.din(n1750), .dout(n1751));
  jnot g1110(.din(\in3[117] ), .dout(n1752));
  jand g1111(.dina(n1752), .dinb(\in2[117] ), .dout(n1753));
  jnot g1112(.din(\in3[116] ), .dout(n1754));
  jand g1113(.dina(n1754), .dinb(\in2[116] ), .dout(n1755));
  jor  g1114(.dina(n1755), .dinb(n1753), .dout(n1756));
  jand g1115(.dina(n1756), .dinb(n1751), .dout(n1757));
  jnot g1116(.din(n1746), .dout(n1758));
  jnot g1117(.din(\in3[119] ), .dout(n1759));
  jand g1118(.dina(n1759), .dinb(\in2[119] ), .dout(n1760));
  jnot g1119(.din(\in3[118] ), .dout(n1761));
  jand g1120(.dina(n1761), .dinb(\in2[118] ), .dout(n1762));
  jor  g1121(.dina(n1762), .dinb(n1760), .dout(n1763));
  jand g1122(.dina(n1763), .dinb(n1758), .dout(n1764));
  jor  g1123(.dina(n1764), .dinb(n1757), .dout(n1765));
  jnot g1124(.din(n1765), .dout(n1766));
  jnot g1125(.din(\in3[115] ), .dout(n1767));
  jand g1126(.dina(n1767), .dinb(\in2[115] ), .dout(n1768));
  jnot g1127(.din(n1768), .dout(n1769));
  jnot g1128(.din(\in2[113] ), .dout(n1770));
  jand g1129(.dina(\in3[113] ), .dinb(n1770), .dout(n1771));
  jnot g1130(.din(\in2[112] ), .dout(n1772));
  jand g1131(.dina(\in3[112] ), .dinb(n1772), .dout(n1773));
  jor  g1132(.dina(n1773), .dinb(n1771), .dout(n1774));
  jnot g1133(.din(\in2[110] ), .dout(n1775));
  jand g1134(.dina(\in3[110] ), .dinb(n1775), .dout(n1776));
  jnot g1135(.din(\in2[111] ), .dout(n1777));
  jand g1136(.dina(\in3[111] ), .dinb(n1777), .dout(n1778));
  jnot g1137(.din(\in2[109] ), .dout(n1779));
  jand g1138(.dina(\in3[109] ), .dinb(n1779), .dout(n1780));
  jor  g1139(.dina(n1780), .dinb(n1778), .dout(n1781));
  jor  g1140(.dina(n1781), .dinb(n1776), .dout(n1782));
  jnot g1141(.din(n1782), .dout(n1783));
  jnot g1142(.din(\in3[109] ), .dout(n1784));
  jand g1143(.dina(n1784), .dinb(\in2[109] ), .dout(n1785));
  jnot g1144(.din(\in3[108] ), .dout(n1786));
  jand g1145(.dina(n1786), .dinb(\in2[108] ), .dout(n1787));
  jor  g1146(.dina(n1787), .dinb(n1785), .dout(n1788));
  jand g1147(.dina(n1788), .dinb(n1783), .dout(n1789));
  jnot g1148(.din(n1778), .dout(n1790));
  jnot g1149(.din(\in3[111] ), .dout(n1791));
  jand g1150(.dina(n1791), .dinb(\in2[111] ), .dout(n1792));
  jnot g1151(.din(\in3[110] ), .dout(n1793));
  jand g1152(.dina(n1793), .dinb(\in2[110] ), .dout(n1794));
  jor  g1153(.dina(n1794), .dinb(n1792), .dout(n1795));
  jand g1154(.dina(n1795), .dinb(n1790), .dout(n1796));
  jor  g1155(.dina(n1796), .dinb(n1789), .dout(n1797));
  jnot g1156(.din(n1797), .dout(n1798));
  jnot g1157(.din(\in3[107] ), .dout(n1799));
  jand g1158(.dina(n1799), .dinb(\in2[107] ), .dout(n1800));
  jnot g1159(.din(n1800), .dout(n1801));
  jnot g1160(.din(\in2[102] ), .dout(n1802));
  jand g1161(.dina(\in3[102] ), .dinb(n1802), .dout(n1803));
  jnot g1162(.din(\in2[103] ), .dout(n1804));
  jand g1163(.dina(\in3[103] ), .dinb(n1804), .dout(n1805));
  jnot g1164(.din(\in2[101] ), .dout(n1806));
  jand g1165(.dina(\in3[101] ), .dinb(n1806), .dout(n1807));
  jor  g1166(.dina(n1807), .dinb(n1805), .dout(n1808));
  jor  g1167(.dina(n1808), .dinb(n1803), .dout(n1809));
  jnot g1168(.din(n1809), .dout(n1810));
  jnot g1169(.din(\in3[101] ), .dout(n1811));
  jand g1170(.dina(n1811), .dinb(\in2[101] ), .dout(n1812));
  jnot g1171(.din(\in3[100] ), .dout(n1813));
  jand g1172(.dina(n1813), .dinb(\in2[100] ), .dout(n1814));
  jor  g1173(.dina(n1814), .dinb(n1812), .dout(n1815));
  jand g1174(.dina(n1815), .dinb(n1810), .dout(n1816));
  jnot g1175(.din(n1805), .dout(n1817));
  jnot g1176(.din(\in3[103] ), .dout(n1818));
  jand g1177(.dina(n1818), .dinb(\in2[103] ), .dout(n1819));
  jnot g1178(.din(\in3[102] ), .dout(n1820));
  jand g1179(.dina(n1820), .dinb(\in2[102] ), .dout(n1821));
  jor  g1180(.dina(n1821), .dinb(n1819), .dout(n1822));
  jand g1181(.dina(n1822), .dinb(n1817), .dout(n1823));
  jor  g1182(.dina(n1823), .dinb(n1816), .dout(n1824));
  jnot g1183(.din(n1824), .dout(n1825));
  jnot g1184(.din(\in3[99] ), .dout(n1826));
  jand g1185(.dina(n1826), .dinb(\in2[99] ), .dout(n1827));
  jnot g1186(.din(n1827), .dout(n1828));
  jnot g1187(.din(\in2[97] ), .dout(n1829));
  jand g1188(.dina(\in3[97] ), .dinb(n1829), .dout(n1830));
  jnot g1189(.din(\in2[96] ), .dout(n1831));
  jand g1190(.dina(\in3[96] ), .dinb(n1831), .dout(n1832));
  jor  g1191(.dina(n1832), .dinb(n1830), .dout(n1833));
  jnot g1192(.din(\in2[94] ), .dout(n1834));
  jand g1193(.dina(\in3[94] ), .dinb(n1834), .dout(n1835));
  jnot g1194(.din(\in2[95] ), .dout(n1836));
  jand g1195(.dina(\in3[95] ), .dinb(n1836), .dout(n1837));
  jnot g1196(.din(\in2[93] ), .dout(n1838));
  jand g1197(.dina(\in3[93] ), .dinb(n1838), .dout(n1839));
  jor  g1198(.dina(n1839), .dinb(n1837), .dout(n1840));
  jor  g1199(.dina(n1840), .dinb(n1835), .dout(n1841));
  jnot g1200(.din(n1841), .dout(n1842));
  jnot g1201(.din(\in3[93] ), .dout(n1843));
  jand g1202(.dina(n1843), .dinb(\in2[93] ), .dout(n1844));
  jnot g1203(.din(\in3[92] ), .dout(n1845));
  jand g1204(.dina(n1845), .dinb(\in2[92] ), .dout(n1846));
  jor  g1205(.dina(n1846), .dinb(n1844), .dout(n1847));
  jand g1206(.dina(n1847), .dinb(n1842), .dout(n1848));
  jnot g1207(.din(n1837), .dout(n1849));
  jnot g1208(.din(\in3[95] ), .dout(n1850));
  jand g1209(.dina(n1850), .dinb(\in2[95] ), .dout(n1851));
  jnot g1210(.din(\in3[94] ), .dout(n1852));
  jand g1211(.dina(n1852), .dinb(\in2[94] ), .dout(n1853));
  jor  g1212(.dina(n1853), .dinb(n1851), .dout(n1854));
  jand g1213(.dina(n1854), .dinb(n1849), .dout(n1855));
  jor  g1214(.dina(n1855), .dinb(n1848), .dout(n1856));
  jnot g1215(.din(n1856), .dout(n1857));
  jnot g1216(.din(\in3[91] ), .dout(n1858));
  jand g1217(.dina(n1858), .dinb(\in2[91] ), .dout(n1859));
  jnot g1218(.din(n1859), .dout(n1860));
  jnot g1219(.din(\in2[86] ), .dout(n1861));
  jand g1220(.dina(\in3[86] ), .dinb(n1861), .dout(n1862));
  jnot g1221(.din(\in2[87] ), .dout(n1863));
  jand g1222(.dina(\in3[87] ), .dinb(n1863), .dout(n1864));
  jnot g1223(.din(\in2[85] ), .dout(n1865));
  jand g1224(.dina(\in3[85] ), .dinb(n1865), .dout(n1866));
  jor  g1225(.dina(n1866), .dinb(n1864), .dout(n1867));
  jor  g1226(.dina(n1867), .dinb(n1862), .dout(n1868));
  jnot g1227(.din(n1868), .dout(n1869));
  jnot g1228(.din(\in3[85] ), .dout(n1870));
  jand g1229(.dina(n1870), .dinb(\in2[85] ), .dout(n1871));
  jnot g1230(.din(\in3[84] ), .dout(n1872));
  jand g1231(.dina(n1872), .dinb(\in2[84] ), .dout(n1873));
  jor  g1232(.dina(n1873), .dinb(n1871), .dout(n1874));
  jand g1233(.dina(n1874), .dinb(n1869), .dout(n1875));
  jnot g1234(.din(n1864), .dout(n1876));
  jnot g1235(.din(\in3[87] ), .dout(n1877));
  jand g1236(.dina(n1877), .dinb(\in2[87] ), .dout(n1878));
  jnot g1237(.din(\in3[86] ), .dout(n1879));
  jand g1238(.dina(n1879), .dinb(\in2[86] ), .dout(n1880));
  jor  g1239(.dina(n1880), .dinb(n1878), .dout(n1881));
  jand g1240(.dina(n1881), .dinb(n1876), .dout(n1882));
  jor  g1241(.dina(n1882), .dinb(n1875), .dout(n1883));
  jnot g1242(.din(n1883), .dout(n1884));
  jnot g1243(.din(\in3[83] ), .dout(n1885));
  jand g1244(.dina(n1885), .dinb(\in2[83] ), .dout(n1886));
  jnot g1245(.din(n1886), .dout(n1887));
  jnot g1246(.din(\in2[81] ), .dout(n1888));
  jand g1247(.dina(\in3[81] ), .dinb(n1888), .dout(n1889));
  jnot g1248(.din(\in2[80] ), .dout(n1890));
  jand g1249(.dina(\in3[80] ), .dinb(n1890), .dout(n1891));
  jor  g1250(.dina(n1891), .dinb(n1889), .dout(n1892));
  jnot g1251(.din(\in2[78] ), .dout(n1893));
  jand g1252(.dina(\in3[78] ), .dinb(n1893), .dout(n1894));
  jnot g1253(.din(\in2[79] ), .dout(n1895));
  jand g1254(.dina(\in3[79] ), .dinb(n1895), .dout(n1896));
  jnot g1255(.din(\in2[77] ), .dout(n1897));
  jand g1256(.dina(\in3[77] ), .dinb(n1897), .dout(n1898));
  jor  g1257(.dina(n1898), .dinb(n1896), .dout(n1899));
  jor  g1258(.dina(n1899), .dinb(n1894), .dout(n1900));
  jnot g1259(.din(n1900), .dout(n1901));
  jnot g1260(.din(\in3[77] ), .dout(n1902));
  jand g1261(.dina(n1902), .dinb(\in2[77] ), .dout(n1903));
  jnot g1262(.din(\in3[76] ), .dout(n1904));
  jand g1263(.dina(n1904), .dinb(\in2[76] ), .dout(n1905));
  jor  g1264(.dina(n1905), .dinb(n1903), .dout(n1906));
  jand g1265(.dina(n1906), .dinb(n1901), .dout(n1907));
  jnot g1266(.din(n1896), .dout(n1908));
  jnot g1267(.din(\in3[79] ), .dout(n1909));
  jand g1268(.dina(n1909), .dinb(\in2[79] ), .dout(n1910));
  jnot g1269(.din(\in3[78] ), .dout(n1911));
  jand g1270(.dina(n1911), .dinb(\in2[78] ), .dout(n1912));
  jor  g1271(.dina(n1912), .dinb(n1910), .dout(n1913));
  jand g1272(.dina(n1913), .dinb(n1908), .dout(n1914));
  jor  g1273(.dina(n1914), .dinb(n1907), .dout(n1915));
  jnot g1274(.din(n1915), .dout(n1916));
  jnot g1275(.din(\in3[75] ), .dout(n1917));
  jand g1276(.dina(n1917), .dinb(\in2[75] ), .dout(n1918));
  jnot g1277(.din(n1918), .dout(n1919));
  jnot g1278(.din(\in2[70] ), .dout(n1920));
  jand g1279(.dina(\in3[70] ), .dinb(n1920), .dout(n1921));
  jnot g1280(.din(\in2[71] ), .dout(n1922));
  jand g1281(.dina(\in3[71] ), .dinb(n1922), .dout(n1923));
  jnot g1282(.din(\in2[69] ), .dout(n1924));
  jand g1283(.dina(\in3[69] ), .dinb(n1924), .dout(n1925));
  jor  g1284(.dina(n1925), .dinb(n1923), .dout(n1926));
  jor  g1285(.dina(n1926), .dinb(n1921), .dout(n1927));
  jnot g1286(.din(n1927), .dout(n1928));
  jnot g1287(.din(\in3[69] ), .dout(n1929));
  jand g1288(.dina(n1929), .dinb(\in2[69] ), .dout(n1930));
  jnot g1289(.din(\in3[68] ), .dout(n1931));
  jand g1290(.dina(n1931), .dinb(\in2[68] ), .dout(n1932));
  jor  g1291(.dina(n1932), .dinb(n1930), .dout(n1933));
  jand g1292(.dina(n1933), .dinb(n1928), .dout(n1934));
  jnot g1293(.din(n1923), .dout(n1935));
  jnot g1294(.din(\in3[71] ), .dout(n1936));
  jand g1295(.dina(n1936), .dinb(\in2[71] ), .dout(n1937));
  jnot g1296(.din(\in3[70] ), .dout(n1938));
  jand g1297(.dina(n1938), .dinb(\in2[70] ), .dout(n1939));
  jor  g1298(.dina(n1939), .dinb(n1937), .dout(n1940));
  jand g1299(.dina(n1940), .dinb(n1935), .dout(n1941));
  jor  g1300(.dina(n1941), .dinb(n1934), .dout(n1942));
  jnot g1301(.din(n1942), .dout(n1943));
  jnot g1302(.din(\in3[67] ), .dout(n1944));
  jand g1303(.dina(n1944), .dinb(\in2[67] ), .dout(n1945));
  jnot g1304(.din(n1945), .dout(n1946));
  jnot g1305(.din(\in2[65] ), .dout(n1947));
  jand g1306(.dina(\in3[65] ), .dinb(n1947), .dout(n1948));
  jnot g1307(.din(n1948), .dout(n1949));
  jnot g1308(.din(\in3[64] ), .dout(n1950));
  jand g1309(.dina(n1950), .dinb(\in2[64] ), .dout(n1951));
  jand g1310(.dina(n1951), .dinb(n1949), .dout(n1952));
  jnot g1311(.din(\in3[66] ), .dout(n1953));
  jand g1312(.dina(n1953), .dinb(\in2[66] ), .dout(n1954));
  jnot g1313(.din(\in3[65] ), .dout(n1955));
  jand g1314(.dina(n1955), .dinb(\in2[65] ), .dout(n1956));
  jor  g1315(.dina(n1956), .dinb(n1954), .dout(n1957));
  jor  g1316(.dina(n1957), .dinb(n1952), .dout(n1958));
  jnot g1317(.din(n1958), .dout(n1959));
  jnot g1318(.din(\in3[59] ), .dout(n1960));
  jnot g1319(.din(\in2[60] ), .dout(n1961));
  jand g1320(.dina(\in3[60] ), .dinb(n1961), .dout(n1962));
  jnot g1321(.din(\in2[63] ), .dout(n1963));
  jand g1322(.dina(\in3[63] ), .dinb(n1963), .dout(n1964));
  jnot g1323(.din(\in2[61] ), .dout(n1965));
  jand g1324(.dina(\in3[61] ), .dinb(n1965), .dout(n1966));
  jnot g1325(.din(\in2[62] ), .dout(n1967));
  jand g1326(.dina(\in3[62] ), .dinb(n1967), .dout(n1968));
  jor  g1327(.dina(n1968), .dinb(n1966), .dout(n1969));
  jor  g1328(.dina(n1969), .dinb(n1964), .dout(n1970));
  jor  g1329(.dina(n1970), .dinb(n1962), .dout(n1971));
  jnot g1330(.din(n1971), .dout(n1972));
  jand g1331(.dina(n1972), .dinb(\in2[59] ), .dout(n1973));
  jand g1332(.dina(n1973), .dinb(n1960), .dout(n1974));
  jnot g1333(.din(n1974), .dout(n1975));
  jnot g1334(.din(\in3[51] ), .dout(n1976));
  jnot g1335(.din(\in2[53] ), .dout(n1977));
  jand g1336(.dina(\in3[53] ), .dinb(n1977), .dout(n1978));
  jnot g1337(.din(\in2[55] ), .dout(n1979));
  jand g1338(.dina(\in3[55] ), .dinb(n1979), .dout(n1980));
  jnot g1339(.din(\in2[54] ), .dout(n1981));
  jand g1340(.dina(\in3[54] ), .dinb(n1981), .dout(n1982));
  jor  g1341(.dina(n1982), .dinb(n1980), .dout(n1983));
  jnot g1342(.din(\in2[52] ), .dout(n1984));
  jand g1343(.dina(\in3[52] ), .dinb(n1984), .dout(n1985));
  jor  g1344(.dina(n1985), .dinb(n1983), .dout(n1986));
  jor  g1345(.dina(n1986), .dinb(n1978), .dout(n1987));
  jnot g1346(.din(n1987), .dout(n1988));
  jand g1347(.dina(n1988), .dinb(\in2[51] ), .dout(n1989));
  jand g1348(.dina(n1989), .dinb(n1976), .dout(n1990));
  jnot g1349(.din(n1990), .dout(n1991));
  jnot g1350(.din(\in3[43] ), .dout(n1992));
  jnot g1351(.din(\in2[44] ), .dout(n1993));
  jand g1352(.dina(\in3[44] ), .dinb(n1993), .dout(n1994));
  jnot g1353(.din(\in2[47] ), .dout(n1995));
  jand g1354(.dina(\in3[47] ), .dinb(n1995), .dout(n1996));
  jnot g1355(.din(\in2[45] ), .dout(n1997));
  jand g1356(.dina(\in3[45] ), .dinb(n1997), .dout(n1998));
  jnot g1357(.din(\in2[46] ), .dout(n1999));
  jand g1358(.dina(\in3[46] ), .dinb(n1999), .dout(n2000));
  jor  g1359(.dina(n2000), .dinb(n1998), .dout(n2001));
  jor  g1360(.dina(n2001), .dinb(n1996), .dout(n2002));
  jor  g1361(.dina(n2002), .dinb(n1994), .dout(n2003));
  jnot g1362(.din(n2003), .dout(n2004));
  jand g1363(.dina(n2004), .dinb(\in2[43] ), .dout(n2005));
  jand g1364(.dina(n2005), .dinb(n1992), .dout(n2006));
  jnot g1365(.din(n2006), .dout(n2007));
  jnot g1366(.din(\in3[33] ), .dout(n2008));
  jand g1367(.dina(n2008), .dinb(\in2[33] ), .dout(n2009));
  jnot g1368(.din(\in3[34] ), .dout(n2010));
  jand g1369(.dina(n2010), .dinb(\in2[34] ), .dout(n2011));
  jor  g1370(.dina(n2011), .dinb(n2009), .dout(n2012));
  jnot g1371(.din(\in2[33] ), .dout(n2013));
  jand g1372(.dina(\in3[33] ), .dinb(n2013), .dout(n2014));
  jnot g1373(.din(n2014), .dout(n2015));
  jnot g1374(.din(\in3[32] ), .dout(n2016));
  jand g1375(.dina(n2016), .dinb(\in2[32] ), .dout(n2017));
  jand g1376(.dina(n2017), .dinb(n2015), .dout(n2018));
  jor  g1377(.dina(n2018), .dinb(n2012), .dout(n2019));
  jnot g1378(.din(\in2[35] ), .dout(n2020));
  jand g1379(.dina(\in3[35] ), .dinb(n2020), .dout(n2021));
  jnot g1380(.din(\in2[34] ), .dout(n2022));
  jand g1381(.dina(\in3[34] ), .dinb(n2022), .dout(n2023));
  jor  g1382(.dina(n2023), .dinb(n2021), .dout(n2024));
  jnot g1383(.din(\in2[36] ), .dout(n2025));
  jand g1384(.dina(\in3[36] ), .dinb(n2025), .dout(n2026));
  jnot g1385(.din(\in2[38] ), .dout(n2027));
  jand g1386(.dina(\in3[38] ), .dinb(n2027), .dout(n2028));
  jnot g1387(.din(\in2[39] ), .dout(n2029));
  jand g1388(.dina(\in3[39] ), .dinb(n2029), .dout(n2030));
  jnot g1389(.din(\in2[37] ), .dout(n2031));
  jand g1390(.dina(\in3[37] ), .dinb(n2031), .dout(n2032));
  jor  g1391(.dina(n2032), .dinb(n2030), .dout(n2033));
  jor  g1392(.dina(n2033), .dinb(n2028), .dout(n2034));
  jor  g1393(.dina(n2034), .dinb(n2026), .dout(n2035));
  jor  g1394(.dina(n2035), .dinb(n2024), .dout(n2036));
  jnot g1395(.din(n2036), .dout(n2037));
  jand g1396(.dina(n2037), .dinb(n2019), .dout(n2038));
  jnot g1397(.din(n2038), .dout(n2039));
  jnot g1398(.din(\in2[30] ), .dout(n2040));
  jand g1399(.dina(\in3[30] ), .dinb(n2040), .dout(n2041));
  jnot g1400(.din(\in3[29] ), .dout(n2042));
  jand g1401(.dina(n2042), .dinb(\in2[29] ), .dout(n2043));
  jnot g1402(.din(n2043), .dout(n2044));
  jnot g1403(.din(\in2[29] ), .dout(n2045));
  jand g1404(.dina(\in3[29] ), .dinb(n2045), .dout(n2046));
  jnot g1405(.din(\in3[28] ), .dout(n2047));
  jand g1406(.dina(n2047), .dinb(\in2[28] ), .dout(n2048));
  jnot g1407(.din(n2048), .dout(n2049));
  jnot g1408(.din(\in2[28] ), .dout(n2050));
  jand g1409(.dina(\in3[28] ), .dinb(n2050), .dout(n2051));
  jnot g1410(.din(\in3[27] ), .dout(n2052));
  jand g1411(.dina(n2052), .dinb(\in2[27] ), .dout(n2053));
  jnot g1412(.din(n2053), .dout(n2054));
  jnot g1413(.din(\in2[27] ), .dout(n2055));
  jand g1414(.dina(\in3[27] ), .dinb(n2055), .dout(n2056));
  jnot g1415(.din(\in3[26] ), .dout(n2057));
  jand g1416(.dina(n2057), .dinb(\in2[26] ), .dout(n2058));
  jnot g1417(.din(n2058), .dout(n2059));
  jnot g1418(.din(\in2[23] ), .dout(n2060));
  jand g1419(.dina(\in3[23] ), .dinb(n2060), .dout(n2061));
  jnot g1420(.din(\in2[22] ), .dout(n2062));
  jand g1421(.dina(\in3[22] ), .dinb(n2062), .dout(n2063));
  jnot g1422(.din(\in3[21] ), .dout(n2064));
  jand g1423(.dina(n2064), .dinb(\in2[21] ), .dout(n2065));
  jnot g1424(.din(n2065), .dout(n2066));
  jnot g1425(.din(\in2[21] ), .dout(n2067));
  jand g1426(.dina(\in3[21] ), .dinb(n2067), .dout(n2068));
  jnot g1427(.din(\in3[20] ), .dout(n2069));
  jand g1428(.dina(n2069), .dinb(\in2[20] ), .dout(n2070));
  jnot g1429(.din(n2070), .dout(n2071));
  jnot g1430(.din(\in2[20] ), .dout(n2072));
  jand g1431(.dina(\in3[20] ), .dinb(n2072), .dout(n2073));
  jnot g1432(.din(\in3[19] ), .dout(n2074));
  jand g1433(.dina(n2074), .dinb(\in2[19] ), .dout(n2075));
  jnot g1434(.din(n2075), .dout(n2076));
  jnot g1435(.din(\in2[19] ), .dout(n2077));
  jand g1436(.dina(\in3[19] ), .dinb(n2077), .dout(n2078));
  jnot g1437(.din(\in3[18] ), .dout(n2079));
  jand g1438(.dina(n2079), .dinb(\in2[18] ), .dout(n2080));
  jnot g1439(.din(n2080), .dout(n2081));
  jnot g1440(.din(\in2[15] ), .dout(n2082));
  jand g1441(.dina(\in3[15] ), .dinb(n2082), .dout(n2083));
  jnot g1442(.din(\in2[14] ), .dout(n2084));
  jand g1443(.dina(\in3[14] ), .dinb(n2084), .dout(n2085));
  jnot g1444(.din(\in3[13] ), .dout(n2086));
  jand g1445(.dina(n2086), .dinb(\in2[13] ), .dout(n2087));
  jnot g1446(.din(n2087), .dout(n2088));
  jnot g1447(.din(\in2[13] ), .dout(n2089));
  jand g1448(.dina(\in3[13] ), .dinb(n2089), .dout(n2090));
  jnot g1449(.din(\in3[12] ), .dout(n2091));
  jand g1450(.dina(n2091), .dinb(\in2[12] ), .dout(n2092));
  jnot g1451(.din(n2092), .dout(n2093));
  jnot g1452(.din(\in2[12] ), .dout(n2094));
  jand g1453(.dina(\in3[12] ), .dinb(n2094), .dout(n2095));
  jnot g1454(.din(\in3[11] ), .dout(n2096));
  jand g1455(.dina(n2096), .dinb(\in2[11] ), .dout(n2097));
  jnot g1456(.din(n2097), .dout(n2098));
  jnot g1457(.din(\in2[11] ), .dout(n2099));
  jand g1458(.dina(\in3[11] ), .dinb(n2099), .dout(n2100));
  jnot g1459(.din(\in3[10] ), .dout(n2101));
  jand g1460(.dina(n2101), .dinb(\in2[10] ), .dout(n2102));
  jnot g1461(.din(n2102), .dout(n2103));
  jnot g1462(.din(\in2[7] ), .dout(n2104));
  jand g1463(.dina(\in3[7] ), .dinb(n2104), .dout(n2105));
  jnot g1464(.din(\in2[3] ), .dout(n2106));
  jand g1465(.dina(\in3[3] ), .dinb(n2106), .dout(n2107));
  jnot g1466(.din(\in2[2] ), .dout(n2108));
  jand g1467(.dina(\in3[2] ), .dinb(n2108), .dout(n2109));
  jnot g1468(.din(\in3[1] ), .dout(n2110));
  jand g1469(.dina(n2110), .dinb(\in2[1] ), .dout(n2111));
  jnot g1470(.din(n2111), .dout(n2112));
  jnot g1471(.din(\in2[1] ), .dout(n2113));
  jand g1472(.dina(\in3[1] ), .dinb(n2113), .dout(n2114));
  jnot g1473(.din(\in2[0] ), .dout(n2115));
  jor  g1474(.dina(\in3[0] ), .dinb(n2115), .dout(n2116));
  jor  g1475(.dina(n2116), .dinb(n2114), .dout(n2117));
  jand g1476(.dina(n2117), .dinb(n2112), .dout(n2118));
  jor  g1477(.dina(n2118), .dinb(n2109), .dout(n2119));
  jnot g1478(.din(\in3[3] ), .dout(n2120));
  jand g1479(.dina(n2120), .dinb(\in2[3] ), .dout(n2121));
  jnot g1480(.din(\in3[2] ), .dout(n2122));
  jand g1481(.dina(n2122), .dinb(\in2[2] ), .dout(n2123));
  jor  g1482(.dina(n2123), .dinb(n2121), .dout(n2124));
  jnot g1483(.din(n2124), .dout(n2125));
  jand g1484(.dina(n2125), .dinb(n2119), .dout(n2126));
  jnot g1485(.din(\in2[4] ), .dout(n2127));
  jand g1486(.dina(\in3[4] ), .dinb(n2127), .dout(n2128));
  jor  g1487(.dina(n2128), .dinb(n2126), .dout(n2129));
  jor  g1488(.dina(n2129), .dinb(n2107), .dout(n2130));
  jnot g1489(.din(\in3[4] ), .dout(n2131));
  jand g1490(.dina(n2131), .dinb(\in2[4] ), .dout(n2132));
  jnot g1491(.din(\in3[5] ), .dout(n2133));
  jand g1492(.dina(n2133), .dinb(\in2[5] ), .dout(n2134));
  jor  g1493(.dina(n2134), .dinb(n2132), .dout(n2135));
  jnot g1494(.din(n2135), .dout(n2136));
  jand g1495(.dina(n2136), .dinb(n2130), .dout(n2137));
  jnot g1496(.din(\in2[6] ), .dout(n2138));
  jand g1497(.dina(\in3[6] ), .dinb(n2138), .dout(n2139));
  jnot g1498(.din(\in2[5] ), .dout(n2140));
  jand g1499(.dina(\in3[5] ), .dinb(n2140), .dout(n2141));
  jor  g1500(.dina(n2141), .dinb(n2139), .dout(n2142));
  jor  g1501(.dina(n2142), .dinb(n2137), .dout(n2143));
  jnot g1502(.din(\in3[7] ), .dout(n2144));
  jand g1503(.dina(n2144), .dinb(\in2[7] ), .dout(n2145));
  jnot g1504(.din(\in3[6] ), .dout(n2146));
  jand g1505(.dina(n2146), .dinb(\in2[6] ), .dout(n2147));
  jor  g1506(.dina(n2147), .dinb(n2145), .dout(n2148));
  jnot g1507(.din(n2148), .dout(n2149));
  jand g1508(.dina(n2149), .dinb(n2143), .dout(n2150));
  jnot g1509(.din(\in2[8] ), .dout(n2151));
  jand g1510(.dina(\in3[8] ), .dinb(n2151), .dout(n2152));
  jor  g1511(.dina(n2152), .dinb(n2150), .dout(n2153));
  jor  g1512(.dina(n2153), .dinb(n2105), .dout(n2154));
  jnot g1513(.din(\in3[8] ), .dout(n2155));
  jand g1514(.dina(n2155), .dinb(\in2[8] ), .dout(n2156));
  jnot g1515(.din(\in3[9] ), .dout(n2157));
  jand g1516(.dina(n2157), .dinb(\in2[9] ), .dout(n2158));
  jor  g1517(.dina(n2158), .dinb(n2156), .dout(n2159));
  jnot g1518(.din(n2159), .dout(n2160));
  jand g1519(.dina(n2160), .dinb(n2154), .dout(n2161));
  jnot g1520(.din(\in2[10] ), .dout(n2162));
  jand g1521(.dina(\in3[10] ), .dinb(n2162), .dout(n2163));
  jnot g1522(.din(\in2[9] ), .dout(n2164));
  jand g1523(.dina(\in3[9] ), .dinb(n2164), .dout(n2165));
  jor  g1524(.dina(n2165), .dinb(n2163), .dout(n2166));
  jor  g1525(.dina(n2166), .dinb(n2161), .dout(n2167));
  jand g1526(.dina(n2167), .dinb(n2103), .dout(n2168));
  jor  g1527(.dina(n2168), .dinb(n2100), .dout(n2169));
  jand g1528(.dina(n2169), .dinb(n2098), .dout(n2170));
  jor  g1529(.dina(n2170), .dinb(n2095), .dout(n2171));
  jand g1530(.dina(n2171), .dinb(n2093), .dout(n2172));
  jor  g1531(.dina(n2172), .dinb(n2090), .dout(n2173));
  jand g1532(.dina(n2173), .dinb(n2088), .dout(n2174));
  jor  g1533(.dina(n2174), .dinb(n2085), .dout(n2175));
  jnot g1534(.din(\in3[15] ), .dout(n2176));
  jand g1535(.dina(n2176), .dinb(\in2[15] ), .dout(n2177));
  jnot g1536(.din(\in3[14] ), .dout(n2178));
  jand g1537(.dina(n2178), .dinb(\in2[14] ), .dout(n2179));
  jor  g1538(.dina(n2179), .dinb(n2177), .dout(n2180));
  jnot g1539(.din(n2180), .dout(n2181));
  jand g1540(.dina(n2181), .dinb(n2175), .dout(n2182));
  jnot g1541(.din(\in2[16] ), .dout(n2183));
  jand g1542(.dina(\in3[16] ), .dinb(n2183), .dout(n2184));
  jor  g1543(.dina(n2184), .dinb(n2182), .dout(n2185));
  jor  g1544(.dina(n2185), .dinb(n2083), .dout(n2186));
  jnot g1545(.din(\in3[16] ), .dout(n2187));
  jand g1546(.dina(n2187), .dinb(\in2[16] ), .dout(n2188));
  jnot g1547(.din(\in3[17] ), .dout(n2189));
  jand g1548(.dina(n2189), .dinb(\in2[17] ), .dout(n2190));
  jor  g1549(.dina(n2190), .dinb(n2188), .dout(n2191));
  jnot g1550(.din(n2191), .dout(n2192));
  jand g1551(.dina(n2192), .dinb(n2186), .dout(n2193));
  jnot g1552(.din(\in2[18] ), .dout(n2194));
  jand g1553(.dina(\in3[18] ), .dinb(n2194), .dout(n2195));
  jnot g1554(.din(\in2[17] ), .dout(n2196));
  jand g1555(.dina(\in3[17] ), .dinb(n2196), .dout(n2197));
  jor  g1556(.dina(n2197), .dinb(n2195), .dout(n2198));
  jor  g1557(.dina(n2198), .dinb(n2193), .dout(n2199));
  jand g1558(.dina(n2199), .dinb(n2081), .dout(n2200));
  jor  g1559(.dina(n2200), .dinb(n2078), .dout(n2201));
  jand g1560(.dina(n2201), .dinb(n2076), .dout(n2202));
  jor  g1561(.dina(n2202), .dinb(n2073), .dout(n2203));
  jand g1562(.dina(n2203), .dinb(n2071), .dout(n2204));
  jor  g1563(.dina(n2204), .dinb(n2068), .dout(n2205));
  jand g1564(.dina(n2205), .dinb(n2066), .dout(n2206));
  jor  g1565(.dina(n2206), .dinb(n2063), .dout(n2207));
  jnot g1566(.din(\in3[23] ), .dout(n2208));
  jand g1567(.dina(n2208), .dinb(\in2[23] ), .dout(n2209));
  jnot g1568(.din(\in3[22] ), .dout(n2210));
  jand g1569(.dina(n2210), .dinb(\in2[22] ), .dout(n2211));
  jor  g1570(.dina(n2211), .dinb(n2209), .dout(n2212));
  jnot g1571(.din(n2212), .dout(n2213));
  jand g1572(.dina(n2213), .dinb(n2207), .dout(n2214));
  jnot g1573(.din(\in2[24] ), .dout(n2215));
  jand g1574(.dina(\in3[24] ), .dinb(n2215), .dout(n2216));
  jor  g1575(.dina(n2216), .dinb(n2214), .dout(n2217));
  jor  g1576(.dina(n2217), .dinb(n2061), .dout(n2218));
  jnot g1577(.din(\in3[24] ), .dout(n2219));
  jand g1578(.dina(n2219), .dinb(\in2[24] ), .dout(n2220));
  jnot g1579(.din(\in3[25] ), .dout(n2221));
  jand g1580(.dina(n2221), .dinb(\in2[25] ), .dout(n2222));
  jor  g1581(.dina(n2222), .dinb(n2220), .dout(n2223));
  jnot g1582(.din(n2223), .dout(n2224));
  jand g1583(.dina(n2224), .dinb(n2218), .dout(n2225));
  jnot g1584(.din(\in2[26] ), .dout(n2226));
  jand g1585(.dina(\in3[26] ), .dinb(n2226), .dout(n2227));
  jnot g1586(.din(\in2[25] ), .dout(n2228));
  jand g1587(.dina(\in3[25] ), .dinb(n2228), .dout(n2229));
  jor  g1588(.dina(n2229), .dinb(n2227), .dout(n2230));
  jor  g1589(.dina(n2230), .dinb(n2225), .dout(n2231));
  jand g1590(.dina(n2231), .dinb(n2059), .dout(n2232));
  jor  g1591(.dina(n2232), .dinb(n2056), .dout(n2233));
  jand g1592(.dina(n2233), .dinb(n2054), .dout(n2234));
  jor  g1593(.dina(n2234), .dinb(n2051), .dout(n2235));
  jand g1594(.dina(n2235), .dinb(n2049), .dout(n2236));
  jor  g1595(.dina(n2236), .dinb(n2046), .dout(n2237));
  jand g1596(.dina(n2237), .dinb(n2044), .dout(n2238));
  jor  g1597(.dina(n2238), .dinb(n2041), .dout(n2239));
  jnot g1598(.din(\in3[31] ), .dout(n2240));
  jand g1599(.dina(n2240), .dinb(\in2[31] ), .dout(n2241));
  jnot g1600(.din(\in3[30] ), .dout(n2242));
  jand g1601(.dina(n2242), .dinb(\in2[30] ), .dout(n2243));
  jor  g1602(.dina(n2243), .dinb(n2241), .dout(n2244));
  jnot g1603(.din(n2244), .dout(n2245));
  jand g1604(.dina(n2245), .dinb(n2239), .dout(n2246));
  jnot g1605(.din(\in2[31] ), .dout(n2247));
  jand g1606(.dina(\in3[31] ), .dinb(n2247), .dout(n2248));
  jnot g1607(.din(\in2[32] ), .dout(n2249));
  jand g1608(.dina(\in3[32] ), .dinb(n2249), .dout(n2250));
  jor  g1609(.dina(n2250), .dinb(n2248), .dout(n2251));
  jor  g1610(.dina(n2251), .dinb(n2014), .dout(n2252));
  jor  g1611(.dina(n2252), .dinb(n2036), .dout(n2253));
  jor  g1612(.dina(n2253), .dinb(n2246), .dout(n2254));
  jnot g1613(.din(n2034), .dout(n2255));
  jnot g1614(.din(\in3[37] ), .dout(n2256));
  jand g1615(.dina(n2256), .dinb(\in2[37] ), .dout(n2257));
  jnot g1616(.din(\in3[36] ), .dout(n2258));
  jand g1617(.dina(n2258), .dinb(\in2[36] ), .dout(n2259));
  jor  g1618(.dina(n2259), .dinb(n2257), .dout(n2260));
  jand g1619(.dina(n2260), .dinb(n2255), .dout(n2261));
  jnot g1620(.din(n2035), .dout(n2262));
  jnot g1621(.din(\in3[35] ), .dout(n2263));
  jand g1622(.dina(n2263), .dinb(\in2[35] ), .dout(n2264));
  jand g1623(.dina(n2264), .dinb(n2262), .dout(n2265));
  jnot g1624(.din(\in3[39] ), .dout(n2266));
  jand g1625(.dina(n2266), .dinb(\in2[39] ), .dout(n2267));
  jnot g1626(.din(n2030), .dout(n2268));
  jnot g1627(.din(\in3[38] ), .dout(n2269));
  jand g1628(.dina(n2269), .dinb(\in2[38] ), .dout(n2270));
  jand g1629(.dina(n2270), .dinb(n2268), .dout(n2271));
  jor  g1630(.dina(n2271), .dinb(n2267), .dout(n2272));
  jor  g1631(.dina(n2272), .dinb(n2265), .dout(n2273));
  jor  g1632(.dina(n2273), .dinb(n2261), .dout(n2274));
  jnot g1633(.din(n2274), .dout(n2275));
  jand g1634(.dina(n2275), .dinb(n2254), .dout(n2276));
  jand g1635(.dina(n2276), .dinb(n2039), .dout(n2277));
  jnot g1636(.din(\in2[40] ), .dout(n2278));
  jand g1637(.dina(\in3[40] ), .dinb(n2278), .dout(n2279));
  jnot g1638(.din(n2279), .dout(n2280));
  jnot g1639(.din(\in2[41] ), .dout(n2281));
  jand g1640(.dina(\in3[41] ), .dinb(n2281), .dout(n2282));
  jnot g1641(.din(n2282), .dout(n2283));
  jnot g1642(.din(\in2[42] ), .dout(n2284));
  jand g1643(.dina(\in3[42] ), .dinb(n2284), .dout(n2285));
  jnot g1644(.din(\in2[43] ), .dout(n2286));
  jand g1645(.dina(\in3[43] ), .dinb(n2286), .dout(n2287));
  jor  g1646(.dina(n2287), .dinb(n2285), .dout(n2288));
  jor  g1647(.dina(n2288), .dinb(n2003), .dout(n2289));
  jnot g1648(.din(n2289), .dout(n2290));
  jand g1649(.dina(n2290), .dinb(n2283), .dout(n2291));
  jand g1650(.dina(n2291), .dinb(n2280), .dout(n2292));
  jnot g1651(.din(n2292), .dout(n2293));
  jor  g1652(.dina(n2293), .dinb(n2277), .dout(n2294));
  jnot g1653(.din(\in3[41] ), .dout(n2295));
  jand g1654(.dina(n2295), .dinb(\in2[41] ), .dout(n2296));
  jnot g1655(.din(\in3[42] ), .dout(n2297));
  jand g1656(.dina(n2297), .dinb(\in2[42] ), .dout(n2298));
  jor  g1657(.dina(n2298), .dinb(n2296), .dout(n2299));
  jnot g1658(.din(\in3[40] ), .dout(n2300));
  jand g1659(.dina(n2300), .dinb(\in2[40] ), .dout(n2301));
  jand g1660(.dina(n2301), .dinb(n2283), .dout(n2302));
  jor  g1661(.dina(n2302), .dinb(n2299), .dout(n2303));
  jand g1662(.dina(n2303), .dinb(n2290), .dout(n2304));
  jnot g1663(.din(n2002), .dout(n2305));
  jnot g1664(.din(\in3[45] ), .dout(n2306));
  jand g1665(.dina(n2306), .dinb(\in2[45] ), .dout(n2307));
  jnot g1666(.din(\in3[44] ), .dout(n2308));
  jand g1667(.dina(n2308), .dinb(\in2[44] ), .dout(n2309));
  jor  g1668(.dina(n2309), .dinb(n2307), .dout(n2310));
  jand g1669(.dina(n2310), .dinb(n2305), .dout(n2311));
  jnot g1670(.din(n1996), .dout(n2312));
  jnot g1671(.din(\in3[47] ), .dout(n2313));
  jand g1672(.dina(n2313), .dinb(\in2[47] ), .dout(n2314));
  jnot g1673(.din(\in3[46] ), .dout(n2315));
  jand g1674(.dina(n2315), .dinb(\in2[46] ), .dout(n2316));
  jor  g1675(.dina(n2316), .dinb(n2314), .dout(n2317));
  jand g1676(.dina(n2317), .dinb(n2312), .dout(n2318));
  jor  g1677(.dina(n2318), .dinb(n2311), .dout(n2319));
  jor  g1678(.dina(n2319), .dinb(n2304), .dout(n2320));
  jnot g1679(.din(n2320), .dout(n2321));
  jand g1680(.dina(n2321), .dinb(n2294), .dout(n2322));
  jand g1681(.dina(n2322), .dinb(n2007), .dout(n2323));
  jnot g1682(.din(\in2[48] ), .dout(n2324));
  jand g1683(.dina(\in3[48] ), .dinb(n2324), .dout(n2325));
  jnot g1684(.din(n2325), .dout(n2326));
  jnot g1685(.din(\in2[49] ), .dout(n2327));
  jand g1686(.dina(\in3[49] ), .dinb(n2327), .dout(n2328));
  jnot g1687(.din(n2328), .dout(n2329));
  jnot g1688(.din(\in2[50] ), .dout(n2330));
  jand g1689(.dina(\in3[50] ), .dinb(n2330), .dout(n2331));
  jnot g1690(.din(\in2[51] ), .dout(n2332));
  jand g1691(.dina(\in3[51] ), .dinb(n2332), .dout(n2333));
  jor  g1692(.dina(n2333), .dinb(n2331), .dout(n2334));
  jor  g1693(.dina(n2334), .dinb(n1987), .dout(n2335));
  jnot g1694(.din(n2335), .dout(n2336));
  jand g1695(.dina(n2336), .dinb(n2329), .dout(n2337));
  jand g1696(.dina(n2337), .dinb(n2326), .dout(n2338));
  jnot g1697(.din(n2338), .dout(n2339));
  jor  g1698(.dina(n2339), .dinb(n2323), .dout(n2340));
  jnot g1699(.din(\in3[49] ), .dout(n2341));
  jand g1700(.dina(n2341), .dinb(\in2[49] ), .dout(n2342));
  jnot g1701(.din(\in3[50] ), .dout(n2343));
  jand g1702(.dina(n2343), .dinb(\in2[50] ), .dout(n2344));
  jor  g1703(.dina(n2344), .dinb(n2342), .dout(n2345));
  jnot g1704(.din(\in3[48] ), .dout(n2346));
  jand g1705(.dina(n2346), .dinb(\in2[48] ), .dout(n2347));
  jand g1706(.dina(n2347), .dinb(n2329), .dout(n2348));
  jor  g1707(.dina(n2348), .dinb(n2345), .dout(n2349));
  jand g1708(.dina(n2349), .dinb(n2336), .dout(n2350));
  jnot g1709(.din(\in3[55] ), .dout(n2351));
  jand g1710(.dina(n2351), .dinb(\in2[55] ), .dout(n2352));
  jnot g1711(.din(n1983), .dout(n2353));
  jnot g1712(.din(n1978), .dout(n2354));
  jnot g1713(.din(\in3[52] ), .dout(n2355));
  jand g1714(.dina(n2355), .dinb(\in2[52] ), .dout(n2356));
  jand g1715(.dina(n2356), .dinb(n2354), .dout(n2357));
  jnot g1716(.din(\in3[54] ), .dout(n2358));
  jand g1717(.dina(n2358), .dinb(\in2[54] ), .dout(n2359));
  jnot g1718(.din(\in3[53] ), .dout(n2360));
  jand g1719(.dina(n2360), .dinb(\in2[53] ), .dout(n2361));
  jor  g1720(.dina(n2361), .dinb(n2359), .dout(n2362));
  jor  g1721(.dina(n2362), .dinb(n2357), .dout(n2363));
  jand g1722(.dina(n2363), .dinb(n2353), .dout(n2364));
  jor  g1723(.dina(n2364), .dinb(n2352), .dout(n2365));
  jor  g1724(.dina(n2365), .dinb(n2350), .dout(n2366));
  jnot g1725(.din(n2366), .dout(n2367));
  jand g1726(.dina(n2367), .dinb(n2340), .dout(n2368));
  jand g1727(.dina(n2368), .dinb(n1991), .dout(n2369));
  jnot g1728(.din(\in2[56] ), .dout(n2370));
  jand g1729(.dina(\in3[56] ), .dinb(n2370), .dout(n2371));
  jnot g1730(.din(n2371), .dout(n2372));
  jnot g1731(.din(\in2[57] ), .dout(n2373));
  jand g1732(.dina(\in3[57] ), .dinb(n2373), .dout(n2374));
  jnot g1733(.din(n2374), .dout(n2375));
  jnot g1734(.din(\in2[58] ), .dout(n2376));
  jand g1735(.dina(\in3[58] ), .dinb(n2376), .dout(n2377));
  jnot g1736(.din(\in2[59] ), .dout(n2378));
  jand g1737(.dina(\in3[59] ), .dinb(n2378), .dout(n2379));
  jor  g1738(.dina(n2379), .dinb(n2377), .dout(n2380));
  jor  g1739(.dina(n2380), .dinb(n1971), .dout(n2381));
  jnot g1740(.din(n2381), .dout(n2382));
  jand g1741(.dina(n2382), .dinb(n2375), .dout(n2383));
  jand g1742(.dina(n2383), .dinb(n2372), .dout(n2384));
  jnot g1743(.din(n2384), .dout(n2385));
  jor  g1744(.dina(n2385), .dinb(n2369), .dout(n2386));
  jnot g1745(.din(\in3[57] ), .dout(n2387));
  jand g1746(.dina(n2387), .dinb(\in2[57] ), .dout(n2388));
  jnot g1747(.din(\in3[58] ), .dout(n2389));
  jand g1748(.dina(n2389), .dinb(\in2[58] ), .dout(n2390));
  jor  g1749(.dina(n2390), .dinb(n2388), .dout(n2391));
  jnot g1750(.din(\in3[56] ), .dout(n2392));
  jand g1751(.dina(n2392), .dinb(\in2[56] ), .dout(n2393));
  jand g1752(.dina(n2393), .dinb(n2375), .dout(n2394));
  jor  g1753(.dina(n2394), .dinb(n2391), .dout(n2395));
  jand g1754(.dina(n2395), .dinb(n2382), .dout(n2396));
  jnot g1755(.din(n1970), .dout(n2397));
  jnot g1756(.din(\in3[61] ), .dout(n2398));
  jand g1757(.dina(n2398), .dinb(\in2[61] ), .dout(n2399));
  jnot g1758(.din(\in3[60] ), .dout(n2400));
  jand g1759(.dina(n2400), .dinb(\in2[60] ), .dout(n2401));
  jor  g1760(.dina(n2401), .dinb(n2399), .dout(n2402));
  jand g1761(.dina(n2402), .dinb(n2397), .dout(n2403));
  jnot g1762(.din(n1964), .dout(n2404));
  jnot g1763(.din(\in3[63] ), .dout(n2405));
  jand g1764(.dina(n2405), .dinb(\in2[63] ), .dout(n2406));
  jnot g1765(.din(\in3[62] ), .dout(n2407));
  jand g1766(.dina(n2407), .dinb(\in2[62] ), .dout(n2408));
  jor  g1767(.dina(n2408), .dinb(n2406), .dout(n2409));
  jand g1768(.dina(n2409), .dinb(n2404), .dout(n2410));
  jor  g1769(.dina(n2410), .dinb(n2403), .dout(n2411));
  jor  g1770(.dina(n2411), .dinb(n2396), .dout(n2412));
  jnot g1771(.din(n2412), .dout(n2413));
  jand g1772(.dina(n2413), .dinb(n2386), .dout(n2414));
  jand g1773(.dina(n2414), .dinb(n1975), .dout(n2415));
  jnot g1774(.din(\in2[64] ), .dout(n2416));
  jand g1775(.dina(\in3[64] ), .dinb(n2416), .dout(n2417));
  jor  g1776(.dina(n2417), .dinb(n1948), .dout(n2418));
  jor  g1777(.dina(n2418), .dinb(n2415), .dout(n2419));
  jand g1778(.dina(n2419), .dinb(n1959), .dout(n2420));
  jnot g1779(.din(\in2[67] ), .dout(n2421));
  jand g1780(.dina(\in3[67] ), .dinb(n2421), .dout(n2422));
  jnot g1781(.din(\in2[66] ), .dout(n2423));
  jand g1782(.dina(\in3[66] ), .dinb(n2423), .dout(n2424));
  jor  g1783(.dina(n2424), .dinb(n2422), .dout(n2425));
  jor  g1784(.dina(n2425), .dinb(n2420), .dout(n2426));
  jand g1785(.dina(n2426), .dinb(n1946), .dout(n2427));
  jnot g1786(.din(\in2[68] ), .dout(n2428));
  jand g1787(.dina(\in3[68] ), .dinb(n2428), .dout(n2429));
  jor  g1788(.dina(n2429), .dinb(n1927), .dout(n2430));
  jor  g1789(.dina(n2430), .dinb(n2427), .dout(n2431));
  jand g1790(.dina(n2431), .dinb(n1943), .dout(n2432));
  jnot g1791(.din(\in2[75] ), .dout(n2433));
  jand g1792(.dina(\in3[75] ), .dinb(n2433), .dout(n2434));
  jnot g1793(.din(\in2[74] ), .dout(n2435));
  jand g1794(.dina(\in3[74] ), .dinb(n2435), .dout(n2436));
  jor  g1795(.dina(n2436), .dinb(n2434), .dout(n2437));
  jnot g1796(.din(\in2[72] ), .dout(n2438));
  jand g1797(.dina(\in3[72] ), .dinb(n2438), .dout(n2439));
  jnot g1798(.din(\in2[73] ), .dout(n2440));
  jand g1799(.dina(\in3[73] ), .dinb(n2440), .dout(n2441));
  jor  g1800(.dina(n2441), .dinb(n2439), .dout(n2442));
  jor  g1801(.dina(n2442), .dinb(n2437), .dout(n2443));
  jor  g1802(.dina(n2443), .dinb(n2432), .dout(n2444));
  jnot g1803(.din(n2437), .dout(n2445));
  jnot g1804(.din(\in3[73] ), .dout(n2446));
  jand g1805(.dina(n2446), .dinb(\in2[73] ), .dout(n2447));
  jnot g1806(.din(\in3[74] ), .dout(n2448));
  jand g1807(.dina(n2448), .dinb(\in2[74] ), .dout(n2449));
  jor  g1808(.dina(n2449), .dinb(n2447), .dout(n2450));
  jnot g1809(.din(n2441), .dout(n2451));
  jnot g1810(.din(\in3[72] ), .dout(n2452));
  jand g1811(.dina(n2452), .dinb(\in2[72] ), .dout(n2453));
  jand g1812(.dina(n2453), .dinb(n2451), .dout(n2454));
  jor  g1813(.dina(n2454), .dinb(n2450), .dout(n2455));
  jand g1814(.dina(n2455), .dinb(n2445), .dout(n2456));
  jnot g1815(.din(n2456), .dout(n2457));
  jand g1816(.dina(n2457), .dinb(n2444), .dout(n2458));
  jand g1817(.dina(n2458), .dinb(n1919), .dout(n2459));
  jnot g1818(.din(\in2[76] ), .dout(n2460));
  jand g1819(.dina(\in3[76] ), .dinb(n2460), .dout(n2461));
  jor  g1820(.dina(n2461), .dinb(n1900), .dout(n2462));
  jor  g1821(.dina(n2462), .dinb(n2459), .dout(n2463));
  jand g1822(.dina(n2463), .dinb(n1916), .dout(n2464));
  jnot g1823(.din(\in2[83] ), .dout(n2465));
  jand g1824(.dina(\in3[83] ), .dinb(n2465), .dout(n2466));
  jnot g1825(.din(\in2[82] ), .dout(n2467));
  jand g1826(.dina(\in3[82] ), .dinb(n2467), .dout(n2468));
  jor  g1827(.dina(n2468), .dinb(n2466), .dout(n2469));
  jor  g1828(.dina(n2469), .dinb(n2464), .dout(n2470));
  jor  g1829(.dina(n2470), .dinb(n1892), .dout(n2471));
  jnot g1830(.din(n2469), .dout(n2472));
  jnot g1831(.din(\in3[81] ), .dout(n2473));
  jand g1832(.dina(n2473), .dinb(\in2[81] ), .dout(n2474));
  jnot g1833(.din(\in3[82] ), .dout(n2475));
  jand g1834(.dina(n2475), .dinb(\in2[82] ), .dout(n2476));
  jor  g1835(.dina(n2476), .dinb(n2474), .dout(n2477));
  jnot g1836(.din(n1889), .dout(n2478));
  jnot g1837(.din(\in3[80] ), .dout(n2479));
  jand g1838(.dina(n2479), .dinb(\in2[80] ), .dout(n2480));
  jand g1839(.dina(n2480), .dinb(n2478), .dout(n2481));
  jor  g1840(.dina(n2481), .dinb(n2477), .dout(n2482));
  jand g1841(.dina(n2482), .dinb(n2472), .dout(n2483));
  jnot g1842(.din(n2483), .dout(n2484));
  jand g1843(.dina(n2484), .dinb(n2471), .dout(n2485));
  jand g1844(.dina(n2485), .dinb(n1887), .dout(n2486));
  jnot g1845(.din(\in2[84] ), .dout(n2487));
  jand g1846(.dina(\in3[84] ), .dinb(n2487), .dout(n2488));
  jor  g1847(.dina(n2488), .dinb(n1868), .dout(n2489));
  jor  g1848(.dina(n2489), .dinb(n2486), .dout(n2490));
  jand g1849(.dina(n2490), .dinb(n1884), .dout(n2491));
  jnot g1850(.din(\in2[91] ), .dout(n2492));
  jand g1851(.dina(\in3[91] ), .dinb(n2492), .dout(n2493));
  jnot g1852(.din(\in2[90] ), .dout(n2494));
  jand g1853(.dina(\in3[90] ), .dinb(n2494), .dout(n2495));
  jor  g1854(.dina(n2495), .dinb(n2493), .dout(n2496));
  jnot g1855(.din(\in2[88] ), .dout(n2497));
  jand g1856(.dina(\in3[88] ), .dinb(n2497), .dout(n2498));
  jnot g1857(.din(\in2[89] ), .dout(n2499));
  jand g1858(.dina(\in3[89] ), .dinb(n2499), .dout(n2500));
  jor  g1859(.dina(n2500), .dinb(n2498), .dout(n2501));
  jor  g1860(.dina(n2501), .dinb(n2496), .dout(n2502));
  jor  g1861(.dina(n2502), .dinb(n2491), .dout(n2503));
  jnot g1862(.din(n2496), .dout(n2504));
  jnot g1863(.din(\in3[89] ), .dout(n2505));
  jand g1864(.dina(n2505), .dinb(\in2[89] ), .dout(n2506));
  jnot g1865(.din(\in3[90] ), .dout(n2507));
  jand g1866(.dina(n2507), .dinb(\in2[90] ), .dout(n2508));
  jor  g1867(.dina(n2508), .dinb(n2506), .dout(n2509));
  jnot g1868(.din(n2500), .dout(n2510));
  jnot g1869(.din(\in3[88] ), .dout(n2511));
  jand g1870(.dina(n2511), .dinb(\in2[88] ), .dout(n2512));
  jand g1871(.dina(n2512), .dinb(n2510), .dout(n2513));
  jor  g1872(.dina(n2513), .dinb(n2509), .dout(n2514));
  jand g1873(.dina(n2514), .dinb(n2504), .dout(n2515));
  jnot g1874(.din(n2515), .dout(n2516));
  jand g1875(.dina(n2516), .dinb(n2503), .dout(n2517));
  jand g1876(.dina(n2517), .dinb(n1860), .dout(n2518));
  jnot g1877(.din(\in2[92] ), .dout(n2519));
  jand g1878(.dina(\in3[92] ), .dinb(n2519), .dout(n2520));
  jor  g1879(.dina(n2520), .dinb(n1841), .dout(n2521));
  jor  g1880(.dina(n2521), .dinb(n2518), .dout(n2522));
  jand g1881(.dina(n2522), .dinb(n1857), .dout(n2523));
  jnot g1882(.din(\in2[99] ), .dout(n2524));
  jand g1883(.dina(\in3[99] ), .dinb(n2524), .dout(n2525));
  jnot g1884(.din(\in2[98] ), .dout(n2526));
  jand g1885(.dina(\in3[98] ), .dinb(n2526), .dout(n2527));
  jor  g1886(.dina(n2527), .dinb(n2525), .dout(n2528));
  jor  g1887(.dina(n2528), .dinb(n2523), .dout(n2529));
  jor  g1888(.dina(n2529), .dinb(n1833), .dout(n2530));
  jnot g1889(.din(n2528), .dout(n2531));
  jnot g1890(.din(\in3[97] ), .dout(n2532));
  jand g1891(.dina(n2532), .dinb(\in2[97] ), .dout(n2533));
  jnot g1892(.din(\in3[98] ), .dout(n2534));
  jand g1893(.dina(n2534), .dinb(\in2[98] ), .dout(n2535));
  jor  g1894(.dina(n2535), .dinb(n2533), .dout(n2536));
  jnot g1895(.din(n1830), .dout(n2537));
  jnot g1896(.din(\in3[96] ), .dout(n2538));
  jand g1897(.dina(n2538), .dinb(\in2[96] ), .dout(n2539));
  jand g1898(.dina(n2539), .dinb(n2537), .dout(n2540));
  jor  g1899(.dina(n2540), .dinb(n2536), .dout(n2541));
  jand g1900(.dina(n2541), .dinb(n2531), .dout(n2542));
  jnot g1901(.din(n2542), .dout(n2543));
  jand g1902(.dina(n2543), .dinb(n2530), .dout(n2544));
  jand g1903(.dina(n2544), .dinb(n1828), .dout(n2545));
  jnot g1904(.din(\in2[100] ), .dout(n2546));
  jand g1905(.dina(\in3[100] ), .dinb(n2546), .dout(n2547));
  jor  g1906(.dina(n2547), .dinb(n1809), .dout(n2548));
  jor  g1907(.dina(n2548), .dinb(n2545), .dout(n2549));
  jand g1908(.dina(n2549), .dinb(n1825), .dout(n2550));
  jnot g1909(.din(\in2[107] ), .dout(n2551));
  jand g1910(.dina(\in3[107] ), .dinb(n2551), .dout(n2552));
  jnot g1911(.din(\in2[106] ), .dout(n2553));
  jand g1912(.dina(\in3[106] ), .dinb(n2553), .dout(n2554));
  jor  g1913(.dina(n2554), .dinb(n2552), .dout(n2555));
  jnot g1914(.din(\in2[104] ), .dout(n2556));
  jand g1915(.dina(\in3[104] ), .dinb(n2556), .dout(n2557));
  jnot g1916(.din(\in2[105] ), .dout(n2558));
  jand g1917(.dina(\in3[105] ), .dinb(n2558), .dout(n2559));
  jor  g1918(.dina(n2559), .dinb(n2557), .dout(n2560));
  jor  g1919(.dina(n2560), .dinb(n2555), .dout(n2561));
  jor  g1920(.dina(n2561), .dinb(n2550), .dout(n2562));
  jnot g1921(.din(n2555), .dout(n2563));
  jnot g1922(.din(\in3[105] ), .dout(n2564));
  jand g1923(.dina(n2564), .dinb(\in2[105] ), .dout(n2565));
  jnot g1924(.din(\in3[106] ), .dout(n2566));
  jand g1925(.dina(n2566), .dinb(\in2[106] ), .dout(n2567));
  jor  g1926(.dina(n2567), .dinb(n2565), .dout(n2568));
  jnot g1927(.din(n2559), .dout(n2569));
  jnot g1928(.din(\in3[104] ), .dout(n2570));
  jand g1929(.dina(n2570), .dinb(\in2[104] ), .dout(n2571));
  jand g1930(.dina(n2571), .dinb(n2569), .dout(n2572));
  jor  g1931(.dina(n2572), .dinb(n2568), .dout(n2573));
  jand g1932(.dina(n2573), .dinb(n2563), .dout(n2574));
  jnot g1933(.din(n2574), .dout(n2575));
  jand g1934(.dina(n2575), .dinb(n2562), .dout(n2576));
  jand g1935(.dina(n2576), .dinb(n1801), .dout(n2577));
  jnot g1936(.din(\in2[108] ), .dout(n2578));
  jand g1937(.dina(\in3[108] ), .dinb(n2578), .dout(n2579));
  jor  g1938(.dina(n2579), .dinb(n1782), .dout(n2580));
  jor  g1939(.dina(n2580), .dinb(n2577), .dout(n2581));
  jand g1940(.dina(n2581), .dinb(n1798), .dout(n2582));
  jnot g1941(.din(\in2[115] ), .dout(n2583));
  jand g1942(.dina(\in3[115] ), .dinb(n2583), .dout(n2584));
  jnot g1943(.din(\in2[114] ), .dout(n2585));
  jand g1944(.dina(\in3[114] ), .dinb(n2585), .dout(n2586));
  jor  g1945(.dina(n2586), .dinb(n2584), .dout(n2587));
  jor  g1946(.dina(n2587), .dinb(n2582), .dout(n2588));
  jor  g1947(.dina(n2588), .dinb(n1774), .dout(n2589));
  jnot g1948(.din(n2587), .dout(n2590));
  jnot g1949(.din(\in3[113] ), .dout(n2591));
  jand g1950(.dina(n2591), .dinb(\in2[113] ), .dout(n2592));
  jnot g1951(.din(\in3[114] ), .dout(n2593));
  jand g1952(.dina(n2593), .dinb(\in2[114] ), .dout(n2594));
  jor  g1953(.dina(n2594), .dinb(n2592), .dout(n2595));
  jnot g1954(.din(n1771), .dout(n2596));
  jnot g1955(.din(\in3[112] ), .dout(n2597));
  jand g1956(.dina(n2597), .dinb(\in2[112] ), .dout(n2598));
  jand g1957(.dina(n2598), .dinb(n2596), .dout(n2599));
  jor  g1958(.dina(n2599), .dinb(n2595), .dout(n2600));
  jand g1959(.dina(n2600), .dinb(n2590), .dout(n2601));
  jnot g1960(.din(n2601), .dout(n2602));
  jand g1961(.dina(n2602), .dinb(n2589), .dout(n2603));
  jand g1962(.dina(n2603), .dinb(n1769), .dout(n2604));
  jnot g1963(.din(\in2[116] ), .dout(n2605));
  jand g1964(.dina(\in3[116] ), .dinb(n2605), .dout(n2606));
  jor  g1965(.dina(n2606), .dinb(n1750), .dout(n2607));
  jor  g1966(.dina(n2607), .dinb(n2604), .dout(n2608));
  jand g1967(.dina(n2608), .dinb(n1766), .dout(n2609));
  jnot g1968(.din(\in2[123] ), .dout(n2610));
  jand g1969(.dina(\in3[123] ), .dinb(n2610), .dout(n2611));
  jnot g1970(.din(\in2[122] ), .dout(n2612));
  jand g1971(.dina(\in3[122] ), .dinb(n2612), .dout(n2613));
  jor  g1972(.dina(n2613), .dinb(n2611), .dout(n2614));
  jnot g1973(.din(\in2[120] ), .dout(n2615));
  jand g1974(.dina(\in3[120] ), .dinb(n2615), .dout(n2616));
  jnot g1975(.din(\in2[121] ), .dout(n2617));
  jand g1976(.dina(\in3[121] ), .dinb(n2617), .dout(n2618));
  jor  g1977(.dina(n2618), .dinb(n2616), .dout(n2619));
  jor  g1978(.dina(n2619), .dinb(n2614), .dout(n2620));
  jor  g1979(.dina(n2620), .dinb(n2609), .dout(n2621));
  jnot g1980(.din(n2614), .dout(n2622));
  jnot g1981(.din(\in3[121] ), .dout(n2623));
  jand g1982(.dina(n2623), .dinb(\in2[121] ), .dout(n2624));
  jnot g1983(.din(\in3[122] ), .dout(n2625));
  jand g1984(.dina(n2625), .dinb(\in2[122] ), .dout(n2626));
  jor  g1985(.dina(n2626), .dinb(n2624), .dout(n2627));
  jnot g1986(.din(n2618), .dout(n2628));
  jnot g1987(.din(\in3[120] ), .dout(n2629));
  jand g1988(.dina(n2629), .dinb(\in2[120] ), .dout(n2630));
  jand g1989(.dina(n2630), .dinb(n2628), .dout(n2631));
  jor  g1990(.dina(n2631), .dinb(n2627), .dout(n2632));
  jand g1991(.dina(n2632), .dinb(n2622), .dout(n2633));
  jnot g1992(.din(n2633), .dout(n2634));
  jand g1993(.dina(n2634), .dinb(n2621), .dout(n2635));
  jand g1994(.dina(n2635), .dinb(n1742), .dout(n2636));
  jnot g1995(.din(\in2[124] ), .dout(n2637));
  jand g1996(.dina(\in3[124] ), .dinb(n2637), .dout(n2638));
  jor  g1997(.dina(n2638), .dinb(n1728), .dout(n2639));
  jnot g1998(.din(n2639), .dout(n2640));
  jand g1999(.dina(\in3[127] ), .dinb(\in2[127] ), .dout(n2641));
  jnot g2000(.din(n2641), .dout(n2642));
  jand g2001(.dina(\in1[127] ), .dinb(\in0[127] ), .dout(n2643));
  jand g2002(.dina(n2643), .dinb(n2642), .dout(n2644));
  jand g2003(.dina(n1721), .dinb(n1534), .dout(n2645));
  jand g2004(.dina(n1562), .dinb(n1554), .dout(n2646));
  jor  g2005(.dina(n2646), .dinb(n2645), .dout(n2647));
  jnot g2006(.din(\in3[127] ), .dout(n2648));
  jand g2007(.dina(n2648), .dinb(\in2[127] ), .dout(n2649));
  jnot g2008(.din(n2649), .dout(n2650));
  jnot g2009(.din(n1774), .dout(n2651));
  jnot g2010(.din(n1833), .dout(n2652));
  jnot g2011(.din(n1892), .dout(n2653));
  jnot g2012(.din(n2041), .dout(n2654));
  jnot g2013(.din(n2046), .dout(n2655));
  jnot g2014(.din(n2051), .dout(n2656));
  jnot g2015(.din(n2056), .dout(n2657));
  jnot g2016(.din(n2061), .dout(n2658));
  jnot g2017(.din(n2063), .dout(n2659));
  jnot g2018(.din(n2068), .dout(n2660));
  jnot g2019(.din(n2073), .dout(n2661));
  jnot g2020(.din(n2078), .dout(n2662));
  jnot g2021(.din(n2083), .dout(n2663));
  jnot g2022(.din(n2085), .dout(n2664));
  jnot g2023(.din(n2090), .dout(n2665));
  jnot g2024(.din(n2095), .dout(n2666));
  jnot g2025(.din(n2100), .dout(n2667));
  jnot g2026(.din(n2105), .dout(n2668));
  jnot g2027(.din(n2107), .dout(n2669));
  jnot g2028(.din(n2109), .dout(n2670));
  jor  g2029(.dina(n2110), .dinb(\in2[1] ), .dout(n2671));
  jnot g2030(.din(\in3[0] ), .dout(n2672));
  jand g2031(.dina(n2672), .dinb(\in2[0] ), .dout(n2673));
  jand g2032(.dina(n2673), .dinb(n2671), .dout(n2674));
  jor  g2033(.dina(n2674), .dinb(n2111), .dout(n2675));
  jand g2034(.dina(n2675), .dinb(n2670), .dout(n2676));
  jor  g2035(.dina(n2124), .dinb(n2676), .dout(n2677));
  jnot g2036(.din(n2128), .dout(n2678));
  jand g2037(.dina(n2678), .dinb(n2677), .dout(n2679));
  jand g2038(.dina(n2679), .dinb(n2669), .dout(n2680));
  jor  g2039(.dina(n2135), .dinb(n2680), .dout(n2681));
  jnot g2040(.din(n2142), .dout(n2682));
  jand g2041(.dina(n2682), .dinb(n2681), .dout(n2683));
  jor  g2042(.dina(n2148), .dinb(n2683), .dout(n2684));
  jnot g2043(.din(n2152), .dout(n2685));
  jand g2044(.dina(n2685), .dinb(n2684), .dout(n2686));
  jand g2045(.dina(n2686), .dinb(n2668), .dout(n2687));
  jor  g2046(.dina(n2159), .dinb(n2687), .dout(n2688));
  jnot g2047(.din(n2166), .dout(n2689));
  jand g2048(.dina(n2689), .dinb(n2688), .dout(n2690));
  jor  g2049(.dina(n2690), .dinb(n2102), .dout(n2691));
  jand g2050(.dina(n2691), .dinb(n2667), .dout(n2692));
  jor  g2051(.dina(n2692), .dinb(n2097), .dout(n2693));
  jand g2052(.dina(n2693), .dinb(n2666), .dout(n2694));
  jor  g2053(.dina(n2694), .dinb(n2092), .dout(n2695));
  jand g2054(.dina(n2695), .dinb(n2665), .dout(n2696));
  jor  g2055(.dina(n2696), .dinb(n2087), .dout(n2697));
  jand g2056(.dina(n2697), .dinb(n2664), .dout(n2698));
  jor  g2057(.dina(n2180), .dinb(n2698), .dout(n2699));
  jnot g2058(.din(n2184), .dout(n2700));
  jand g2059(.dina(n2700), .dinb(n2699), .dout(n2701));
  jand g2060(.dina(n2701), .dinb(n2663), .dout(n2702));
  jor  g2061(.dina(n2191), .dinb(n2702), .dout(n2703));
  jnot g2062(.din(n2198), .dout(n2704));
  jand g2063(.dina(n2704), .dinb(n2703), .dout(n2705));
  jor  g2064(.dina(n2705), .dinb(n2080), .dout(n2706));
  jand g2065(.dina(n2706), .dinb(n2662), .dout(n2707));
  jor  g2066(.dina(n2707), .dinb(n2075), .dout(n2708));
  jand g2067(.dina(n2708), .dinb(n2661), .dout(n2709));
  jor  g2068(.dina(n2709), .dinb(n2070), .dout(n2710));
  jand g2069(.dina(n2710), .dinb(n2660), .dout(n2711));
  jor  g2070(.dina(n2711), .dinb(n2065), .dout(n2712));
  jand g2071(.dina(n2712), .dinb(n2659), .dout(n2713));
  jor  g2072(.dina(n2212), .dinb(n2713), .dout(n2714));
  jnot g2073(.din(n2216), .dout(n2715));
  jand g2074(.dina(n2715), .dinb(n2714), .dout(n2716));
  jand g2075(.dina(n2716), .dinb(n2658), .dout(n2717));
  jor  g2076(.dina(n2223), .dinb(n2717), .dout(n2718));
  jnot g2077(.din(n2230), .dout(n2719));
  jand g2078(.dina(n2719), .dinb(n2718), .dout(n2720));
  jor  g2079(.dina(n2720), .dinb(n2058), .dout(n2721));
  jand g2080(.dina(n2721), .dinb(n2657), .dout(n2722));
  jor  g2081(.dina(n2722), .dinb(n2053), .dout(n2723));
  jand g2082(.dina(n2723), .dinb(n2656), .dout(n2724));
  jor  g2083(.dina(n2724), .dinb(n2048), .dout(n2725));
  jand g2084(.dina(n2725), .dinb(n2655), .dout(n2726));
  jor  g2085(.dina(n2726), .dinb(n2043), .dout(n2727));
  jand g2086(.dina(n2727), .dinb(n2654), .dout(n2728));
  jor  g2087(.dina(n2244), .dinb(n2728), .dout(n2729));
  jnot g2088(.din(n2253), .dout(n2730));
  jand g2089(.dina(n2730), .dinb(n2729), .dout(n2731));
  jor  g2090(.dina(n2274), .dinb(n2731), .dout(n2732));
  jor  g2091(.dina(n2732), .dinb(n2038), .dout(n2733));
  jand g2092(.dina(n2292), .dinb(n2733), .dout(n2734));
  jor  g2093(.dina(n2320), .dinb(n2734), .dout(n2735));
  jor  g2094(.dina(n2735), .dinb(n2006), .dout(n2736));
  jand g2095(.dina(n2338), .dinb(n2736), .dout(n2737));
  jor  g2096(.dina(n2366), .dinb(n2737), .dout(n2738));
  jor  g2097(.dina(n2738), .dinb(n1990), .dout(n2739));
  jand g2098(.dina(n2384), .dinb(n2739), .dout(n2740));
  jor  g2099(.dina(n2412), .dinb(n2740), .dout(n2741));
  jor  g2100(.dina(n2741), .dinb(n1974), .dout(n2742));
  jnot g2101(.din(n2418), .dout(n2743));
  jand g2102(.dina(n2743), .dinb(n2742), .dout(n2744));
  jor  g2103(.dina(n2744), .dinb(n1958), .dout(n2745));
  jnot g2104(.din(n2425), .dout(n2746));
  jand g2105(.dina(n2746), .dinb(n2745), .dout(n2747));
  jor  g2106(.dina(n2747), .dinb(n1945), .dout(n2748));
  jnot g2107(.din(n2430), .dout(n2749));
  jand g2108(.dina(n2749), .dinb(n2748), .dout(n2750));
  jor  g2109(.dina(n2750), .dinb(n1942), .dout(n2751));
  jnot g2110(.din(n2443), .dout(n2752));
  jand g2111(.dina(n2752), .dinb(n2751), .dout(n2753));
  jor  g2112(.dina(n2456), .dinb(n2753), .dout(n2754));
  jor  g2113(.dina(n2754), .dinb(n1918), .dout(n2755));
  jnot g2114(.din(n2462), .dout(n2756));
  jand g2115(.dina(n2756), .dinb(n2755), .dout(n2757));
  jor  g2116(.dina(n2757), .dinb(n1915), .dout(n2758));
  jand g2117(.dina(n2472), .dinb(n2758), .dout(n2759));
  jand g2118(.dina(n2759), .dinb(n2653), .dout(n2760));
  jor  g2119(.dina(n2483), .dinb(n2760), .dout(n2761));
  jor  g2120(.dina(n2761), .dinb(n1886), .dout(n2762));
  jnot g2121(.din(n2489), .dout(n2763));
  jand g2122(.dina(n2763), .dinb(n2762), .dout(n2764));
  jor  g2123(.dina(n2764), .dinb(n1883), .dout(n2765));
  jnot g2124(.din(n2502), .dout(n2766));
  jand g2125(.dina(n2766), .dinb(n2765), .dout(n2767));
  jor  g2126(.dina(n2515), .dinb(n2767), .dout(n2768));
  jor  g2127(.dina(n2768), .dinb(n1859), .dout(n2769));
  jnot g2128(.din(n2521), .dout(n2770));
  jand g2129(.dina(n2770), .dinb(n2769), .dout(n2771));
  jor  g2130(.dina(n2771), .dinb(n1856), .dout(n2772));
  jand g2131(.dina(n2531), .dinb(n2772), .dout(n2773));
  jand g2132(.dina(n2773), .dinb(n2652), .dout(n2774));
  jor  g2133(.dina(n2542), .dinb(n2774), .dout(n2775));
  jor  g2134(.dina(n2775), .dinb(n1827), .dout(n2776));
  jnot g2135(.din(n2548), .dout(n2777));
  jand g2136(.dina(n2777), .dinb(n2776), .dout(n2778));
  jor  g2137(.dina(n2778), .dinb(n1824), .dout(n2779));
  jnot g2138(.din(n2561), .dout(n2780));
  jand g2139(.dina(n2780), .dinb(n2779), .dout(n2781));
  jor  g2140(.dina(n2574), .dinb(n2781), .dout(n2782));
  jor  g2141(.dina(n2782), .dinb(n1800), .dout(n2783));
  jnot g2142(.din(n2580), .dout(n2784));
  jand g2143(.dina(n2784), .dinb(n2783), .dout(n2785));
  jor  g2144(.dina(n2785), .dinb(n1797), .dout(n2786));
  jand g2145(.dina(n2590), .dinb(n2786), .dout(n2787));
  jand g2146(.dina(n2787), .dinb(n2651), .dout(n2788));
  jor  g2147(.dina(n2601), .dinb(n2788), .dout(n2789));
  jor  g2148(.dina(n2789), .dinb(n1768), .dout(n2790));
  jnot g2149(.din(n2607), .dout(n2791));
  jand g2150(.dina(n2791), .dinb(n2790), .dout(n2792));
  jor  g2151(.dina(n2792), .dinb(n1765), .dout(n2793));
  jnot g2152(.din(n2620), .dout(n2794));
  jand g2153(.dina(n2794), .dinb(n2793), .dout(n2795));
  jor  g2154(.dina(n2633), .dinb(n2795), .dout(n2796));
  jor  g2155(.dina(n2796), .dinb(n1741), .dout(n2797));
  jand g2156(.dina(n2640), .dinb(n2797), .dout(n2798));
  jor  g2157(.dina(n2798), .dinb(n1738), .dout(n2799));
  jand g2158(.dina(n2799), .dinb(n2650), .dout(n2800));
  jor  g2159(.dina(n2648), .dinb(\in2[127] ), .dout(n2801));
  jnot g2160(.din(n2801), .dout(n2802));
  jor  g2161(.dina(n2802), .dinb(n2800), .dout(n2803));
  jand g2162(.dina(n2803), .dinb(n1724), .dout(n2804));
  jor  g2163(.dina(n2639), .dinb(n2636), .dout(n2805));
  jand g2164(.dina(n2805), .dinb(n1739), .dout(n2806));
  jor  g2165(.dina(n2806), .dinb(n2649), .dout(n2807));
  jand g2166(.dina(n2801), .dinb(n2807), .dout(n2808));
  jand g2167(.dina(n2808), .dinb(n1736), .dout(n2809));
  jor  g2168(.dina(n2809), .dinb(n2804), .dout(n2810));
  jnot g2169(.din(n2810), .dout(n2811));
  jand g2170(.dina(n2811), .dinb(n2647), .dout(n2812));
  jand g2171(.dina(n1721), .dinb(n1536), .dout(n2813));
  jand g2172(.dina(n1562), .dinb(n1550), .dout(n2814));
  jor  g2173(.dina(n2814), .dinb(n2813), .dout(n2815));
  jand g2174(.dina(n2803), .dinb(n1726), .dout(n2816));
  jand g2175(.dina(n2808), .dinb(n1732), .dout(n2817));
  jor  g2176(.dina(n2817), .dinb(n2816), .dout(n2818));
  jnot g2177(.din(n2818), .dout(n2819));
  jand g2178(.dina(n2819), .dinb(n2815), .dout(n2820));
  jor  g2179(.dina(n2820), .dinb(n2812), .dout(n2821));
  jnot g2180(.din(n2821), .dout(n2822));
  jand g2181(.dina(n1721), .dinb(n1539), .dout(n2823));
  jand g2182(.dina(n1562), .dinb(n1548), .dout(n2824));
  jor  g2183(.dina(n2824), .dinb(n2823), .dout(n2825));
  jnot g2184(.din(n2825), .dout(n2826));
  jand g2185(.dina(n2803), .dinb(n2637), .dout(n2827));
  jand g2186(.dina(n2808), .dinb(n1730), .dout(n2828));
  jor  g2187(.dina(n2828), .dinb(n2827), .dout(n2829));
  jand g2188(.dina(n2829), .dinb(n2826), .dout(n2830));
  jnot g2189(.din(n2815), .dout(n2831));
  jand g2190(.dina(n2818), .dinb(n2831), .dout(n2832));
  jor  g2191(.dina(n2832), .dinb(n2830), .dout(n2833));
  jand g2192(.dina(n2833), .dinb(n2822), .dout(n2834));
  jnot g2193(.din(n2647), .dout(n2835));
  jand g2194(.dina(n2810), .dinb(n2835), .dout(n2836));
  jor  g2195(.dina(n2836), .dinb(n2834), .dout(n2837));
  jnot g2196(.din(n2837), .dout(n2838));
  jnot g2197(.din(n2829), .dout(n2839));
  jand g2198(.dina(n2839), .dinb(n2825), .dout(n2840));
  jor  g2199(.dina(n2840), .dinb(n2821), .dout(n2841));
  jand g2200(.dina(n2803), .dinb(n1743), .dout(n2842));
  jand g2201(.dina(n2808), .dinb(n1761), .dout(n2843));
  jor  g2202(.dina(n2843), .dinb(n2842), .dout(n2844));
  jnot g2203(.din(n2844), .dout(n2845));
  jand g2204(.dina(n1721), .dinb(n650), .dout(n2846));
  jand g2205(.dina(n1562), .dinb(n668), .dout(n2847));
  jor  g2206(.dina(n2847), .dinb(n2846), .dout(n2848));
  jand g2207(.dina(n2848), .dinb(n2845), .dout(n2849));
  jand g2208(.dina(n1721), .dinb(n652), .dout(n2850));
  jand g2209(.dina(n1562), .dinb(n666), .dout(n2851));
  jor  g2210(.dina(n2851), .dinb(n2850), .dout(n2852));
  jand g2211(.dina(n2803), .dinb(n1745), .dout(n2853));
  jand g2212(.dina(n2808), .dinb(n1759), .dout(n2854));
  jor  g2213(.dina(n2854), .dinb(n2853), .dout(n2855));
  jnot g2214(.din(n2855), .dout(n2856));
  jand g2215(.dina(n2856), .dinb(n2852), .dout(n2857));
  jand g2216(.dina(n1721), .dinb(n654), .dout(n2858));
  jand g2217(.dina(n1562), .dinb(n659), .dout(n2859));
  jor  g2218(.dina(n2859), .dinb(n2858), .dout(n2860));
  jand g2219(.dina(n2803), .dinb(n1747), .dout(n2861));
  jand g2220(.dina(n2808), .dinb(n1752), .dout(n2862));
  jor  g2221(.dina(n2862), .dinb(n2861), .dout(n2863));
  jnot g2222(.din(n2863), .dout(n2864));
  jand g2223(.dina(n2864), .dinb(n2860), .dout(n2865));
  jor  g2224(.dina(n2865), .dinb(n2857), .dout(n2866));
  jor  g2225(.dina(n2866), .dinb(n2849), .dout(n2867));
  jnot g2226(.din(n2867), .dout(n2868));
  jnot g2227(.din(n2860), .dout(n2869));
  jand g2228(.dina(n2863), .dinb(n2869), .dout(n2870));
  jand g2229(.dina(n1721), .dinb(n1507), .dout(n2871));
  jand g2230(.dina(n1562), .dinb(n661), .dout(n2872));
  jor  g2231(.dina(n2872), .dinb(n2871), .dout(n2873));
  jnot g2232(.din(n2873), .dout(n2874));
  jand g2233(.dina(n2803), .dinb(n2605), .dout(n2875));
  jand g2234(.dina(n2808), .dinb(n1754), .dout(n2876));
  jor  g2235(.dina(n2876), .dinb(n2875), .dout(n2877));
  jand g2236(.dina(n2877), .dinb(n2874), .dout(n2878));
  jor  g2237(.dina(n2878), .dinb(n2870), .dout(n2879));
  jand g2238(.dina(n2879), .dinb(n2868), .dout(n2880));
  jnot g2239(.din(n2857), .dout(n2881));
  jnot g2240(.din(n2852), .dout(n2882));
  jand g2241(.dina(n2855), .dinb(n2882), .dout(n2883));
  jnot g2242(.din(n2848), .dout(n2884));
  jand g2243(.dina(n2884), .dinb(n2844), .dout(n2885));
  jor  g2244(.dina(n2885), .dinb(n2883), .dout(n2886));
  jand g2245(.dina(n2886), .dinb(n2881), .dout(n2887));
  jor  g2246(.dina(n2887), .dinb(n2880), .dout(n2888));
  jnot g2247(.din(n2888), .dout(n2889));
  jand g2248(.dina(n1721), .dinb(n1485), .dout(n2890));
  jand g2249(.dina(n1562), .dinb(n674), .dout(n2891));
  jor  g2250(.dina(n2891), .dinb(n2890), .dout(n2892));
  jnot g2251(.din(n2892), .dout(n2893));
  jand g2252(.dina(n2803), .dinb(n2583), .dout(n2894));
  jand g2253(.dina(n2808), .dinb(n1767), .dout(n2895));
  jor  g2254(.dina(n2895), .dinb(n2894), .dout(n2896));
  jand g2255(.dina(n2896), .dinb(n2893), .dout(n2897));
  jnot g2256(.din(n2897), .dout(n2898));
  jand g2257(.dina(n2803), .dinb(n1775), .dout(n2899));
  jand g2258(.dina(n2808), .dinb(n1793), .dout(n2900));
  jor  g2259(.dina(n2900), .dinb(n2899), .dout(n2901));
  jnot g2260(.din(n2901), .dout(n2902));
  jand g2261(.dina(n1721), .dinb(n682), .dout(n2903));
  jand g2262(.dina(n1562), .dinb(n700), .dout(n2904));
  jor  g2263(.dina(n2904), .dinb(n2903), .dout(n2905));
  jand g2264(.dina(n2905), .dinb(n2902), .dout(n2906));
  jand g2265(.dina(n1721), .dinb(n684), .dout(n2907));
  jand g2266(.dina(n1562), .dinb(n698), .dout(n2908));
  jor  g2267(.dina(n2908), .dinb(n2907), .dout(n2909));
  jand g2268(.dina(n2803), .dinb(n1777), .dout(n2910));
  jand g2269(.dina(n2808), .dinb(n1791), .dout(n2911));
  jor  g2270(.dina(n2911), .dinb(n2910), .dout(n2912));
  jnot g2271(.din(n2912), .dout(n2913));
  jand g2272(.dina(n2913), .dinb(n2909), .dout(n2914));
  jand g2273(.dina(n1721), .dinb(n686), .dout(n2915));
  jand g2274(.dina(n1562), .dinb(n691), .dout(n2916));
  jor  g2275(.dina(n2916), .dinb(n2915), .dout(n2917));
  jand g2276(.dina(n2803), .dinb(n1779), .dout(n2918));
  jand g2277(.dina(n2808), .dinb(n1784), .dout(n2919));
  jor  g2278(.dina(n2919), .dinb(n2918), .dout(n2920));
  jnot g2279(.din(n2920), .dout(n2921));
  jand g2280(.dina(n2921), .dinb(n2917), .dout(n2922));
  jor  g2281(.dina(n2922), .dinb(n2914), .dout(n2923));
  jor  g2282(.dina(n2923), .dinb(n2906), .dout(n2924));
  jnot g2283(.din(n2924), .dout(n2925));
  jnot g2284(.din(n2917), .dout(n2926));
  jand g2285(.dina(n2920), .dinb(n2926), .dout(n2927));
  jand g2286(.dina(n1721), .dinb(n1480), .dout(n2928));
  jand g2287(.dina(n1562), .dinb(n693), .dout(n2929));
  jor  g2288(.dina(n2929), .dinb(n2928), .dout(n2930));
  jnot g2289(.din(n2930), .dout(n2931));
  jand g2290(.dina(n2803), .dinb(n2578), .dout(n2932));
  jand g2291(.dina(n2808), .dinb(n1786), .dout(n2933));
  jor  g2292(.dina(n2933), .dinb(n2932), .dout(n2934));
  jand g2293(.dina(n2934), .dinb(n2931), .dout(n2935));
  jor  g2294(.dina(n2935), .dinb(n2927), .dout(n2936));
  jand g2295(.dina(n2936), .dinb(n2925), .dout(n2937));
  jnot g2296(.din(n2937), .dout(n2938));
  jnot g2297(.din(n2934), .dout(n2939));
  jand g2298(.dina(n2939), .dinb(n2930), .dout(n2940));
  jor  g2299(.dina(n2940), .dinb(n2924), .dout(n2941));
  jand g2300(.dina(n1721), .dinb(n1458), .dout(n2942));
  jand g2301(.dina(n1562), .dinb(n706), .dout(n2943));
  jor  g2302(.dina(n2943), .dinb(n2942), .dout(n2944));
  jand g2303(.dina(n2803), .dinb(n2551), .dout(n2945));
  jand g2304(.dina(n2808), .dinb(n1799), .dout(n2946));
  jor  g2305(.dina(n2946), .dinb(n2945), .dout(n2947));
  jnot g2306(.din(n2947), .dout(n2948));
  jand g2307(.dina(n2948), .dinb(n2944), .dout(n2949));
  jand g2308(.dina(n2803), .dinb(n2553), .dout(n2950));
  jand g2309(.dina(n2808), .dinb(n2566), .dout(n2951));
  jor  g2310(.dina(n2951), .dinb(n2950), .dout(n2952));
  jnot g2311(.din(n2952), .dout(n2953));
  jand g2312(.dina(n1721), .dinb(n1460), .dout(n2954));
  jand g2313(.dina(n1562), .dinb(n1468), .dout(n2955));
  jor  g2314(.dina(n2955), .dinb(n2954), .dout(n2956));
  jand g2315(.dina(n2956), .dinb(n2953), .dout(n2957));
  jor  g2316(.dina(n2957), .dinb(n2949), .dout(n2958));
  jand g2317(.dina(n1721), .dinb(n711), .dout(n2959));
  jand g2318(.dina(n1562), .dinb(n1466), .dout(n2960));
  jor  g2319(.dina(n2960), .dinb(n2959), .dout(n2961));
  jand g2320(.dina(n2803), .dinb(n2558), .dout(n2962));
  jand g2321(.dina(n2808), .dinb(n2564), .dout(n2963));
  jor  g2322(.dina(n2963), .dinb(n2962), .dout(n2964));
  jnot g2323(.din(n2964), .dout(n2965));
  jand g2324(.dina(n2965), .dinb(n2961), .dout(n2966));
  jand g2325(.dina(n2803), .dinb(n2556), .dout(n2967));
  jand g2326(.dina(n2808), .dinb(n2570), .dout(n2968));
  jor  g2327(.dina(n2968), .dinb(n2967), .dout(n2969));
  jnot g2328(.din(n2969), .dout(n2970));
  jand g2329(.dina(n1721), .dinb(n709), .dout(n2971));
  jand g2330(.dina(n1562), .dinb(n1472), .dout(n2972));
  jor  g2331(.dina(n2972), .dinb(n2971), .dout(n2973));
  jand g2332(.dina(n2973), .dinb(n2970), .dout(n2974));
  jor  g2333(.dina(n2974), .dinb(n2966), .dout(n2975));
  jor  g2334(.dina(n2975), .dinb(n2958), .dout(n2976));
  jand g2335(.dina(n1721), .dinb(n1453), .dout(n2977));
  jand g2336(.dina(n1562), .dinb(n725), .dout(n2978));
  jor  g2337(.dina(n2978), .dinb(n2977), .dout(n2979));
  jand g2338(.dina(n2803), .dinb(n2546), .dout(n2980));
  jand g2339(.dina(n2808), .dinb(n1813), .dout(n2981));
  jor  g2340(.dina(n2981), .dinb(n2980), .dout(n2982));
  jnot g2341(.din(n2982), .dout(n2983));
  jand g2342(.dina(n2983), .dinb(n2979), .dout(n2984));
  jand g2343(.dina(n2803), .dinb(n1802), .dout(n2985));
  jand g2344(.dina(n2808), .dinb(n1820), .dout(n2986));
  jor  g2345(.dina(n2986), .dinb(n2985), .dout(n2987));
  jnot g2346(.din(n2987), .dout(n2988));
  jand g2347(.dina(n1721), .dinb(n714), .dout(n2989));
  jand g2348(.dina(n1562), .dinb(n732), .dout(n2990));
  jor  g2349(.dina(n2990), .dinb(n2989), .dout(n2991));
  jand g2350(.dina(n2991), .dinb(n2988), .dout(n2992));
  jand g2351(.dina(n1721), .dinb(n716), .dout(n2993));
  jand g2352(.dina(n1562), .dinb(n730), .dout(n2994));
  jor  g2353(.dina(n2994), .dinb(n2993), .dout(n2995));
  jand g2354(.dina(n2803), .dinb(n1804), .dout(n2996));
  jand g2355(.dina(n2808), .dinb(n1818), .dout(n2997));
  jor  g2356(.dina(n2997), .dinb(n2996), .dout(n2998));
  jnot g2357(.din(n2998), .dout(n2999));
  jand g2358(.dina(n2999), .dinb(n2995), .dout(n3000));
  jand g2359(.dina(n1721), .dinb(n718), .dout(n3001));
  jand g2360(.dina(n1562), .dinb(n723), .dout(n3002));
  jor  g2361(.dina(n3002), .dinb(n3001), .dout(n3003));
  jand g2362(.dina(n2803), .dinb(n1806), .dout(n3004));
  jand g2363(.dina(n2808), .dinb(n1811), .dout(n3005));
  jor  g2364(.dina(n3005), .dinb(n3004), .dout(n3006));
  jnot g2365(.din(n3006), .dout(n3007));
  jand g2366(.dina(n3007), .dinb(n3003), .dout(n3008));
  jor  g2367(.dina(n3008), .dinb(n3000), .dout(n3009));
  jor  g2368(.dina(n3009), .dinb(n2992), .dout(n3010));
  jor  g2369(.dina(n3010), .dinb(n2984), .dout(n3011));
  jand g2370(.dina(n1721), .dinb(n1431), .dout(n3012));
  jand g2371(.dina(n1562), .dinb(n738), .dout(n3013));
  jor  g2372(.dina(n3013), .dinb(n3012), .dout(n3014));
  jand g2373(.dina(n2803), .dinb(n2524), .dout(n3015));
  jand g2374(.dina(n2808), .dinb(n1826), .dout(n3016));
  jor  g2375(.dina(n3016), .dinb(n3015), .dout(n3017));
  jnot g2376(.din(n3017), .dout(n3018));
  jand g2377(.dina(n3018), .dinb(n3014), .dout(n3019));
  jand g2378(.dina(n2803), .dinb(n2526), .dout(n3020));
  jand g2379(.dina(n2808), .dinb(n2534), .dout(n3021));
  jor  g2380(.dina(n3021), .dinb(n3020), .dout(n3022));
  jnot g2381(.din(n3022), .dout(n3023));
  jand g2382(.dina(n1721), .dinb(n1433), .dout(n3024));
  jand g2383(.dina(n1562), .dinb(n1441), .dout(n3025));
  jor  g2384(.dina(n3025), .dinb(n3024), .dout(n3026));
  jand g2385(.dina(n3026), .dinb(n3023), .dout(n3027));
  jor  g2386(.dina(n3027), .dinb(n3019), .dout(n3028));
  jand g2387(.dina(n1721), .dinb(n741), .dout(n3029));
  jand g2388(.dina(n1562), .dinb(n1439), .dout(n3030));
  jor  g2389(.dina(n3030), .dinb(n3029), .dout(n3031));
  jand g2390(.dina(n2803), .dinb(n1829), .dout(n3032));
  jand g2391(.dina(n2808), .dinb(n2532), .dout(n3033));
  jor  g2392(.dina(n3033), .dinb(n3032), .dout(n3034));
  jnot g2393(.din(n3034), .dout(n3035));
  jand g2394(.dina(n3035), .dinb(n3031), .dout(n3036));
  jand g2395(.dina(n2803), .dinb(n1831), .dout(n3037));
  jand g2396(.dina(n2808), .dinb(n2538), .dout(n3038));
  jor  g2397(.dina(n3038), .dinb(n3037), .dout(n3039));
  jnot g2398(.din(n3039), .dout(n3040));
  jand g2399(.dina(n1721), .dinb(n743), .dout(n3041));
  jand g2400(.dina(n1562), .dinb(n1445), .dout(n3042));
  jor  g2401(.dina(n3042), .dinb(n3041), .dout(n3043));
  jand g2402(.dina(n3043), .dinb(n3040), .dout(n3044));
  jor  g2403(.dina(n3044), .dinb(n3036), .dout(n3045));
  jor  g2404(.dina(n3045), .dinb(n3028), .dout(n3046));
  jand g2405(.dina(n1721), .dinb(n1426), .dout(n3047));
  jand g2406(.dina(n1562), .dinb(n757), .dout(n3048));
  jor  g2407(.dina(n3048), .dinb(n3047), .dout(n3049));
  jand g2408(.dina(n2803), .dinb(n2519), .dout(n3050));
  jand g2409(.dina(n2808), .dinb(n1845), .dout(n3051));
  jor  g2410(.dina(n3051), .dinb(n3050), .dout(n3052));
  jnot g2411(.din(n3052), .dout(n3053));
  jand g2412(.dina(n3053), .dinb(n3049), .dout(n3054));
  jand g2413(.dina(n2803), .dinb(n1834), .dout(n3055));
  jand g2414(.dina(n2808), .dinb(n1852), .dout(n3056));
  jor  g2415(.dina(n3056), .dinb(n3055), .dout(n3057));
  jnot g2416(.din(n3057), .dout(n3058));
  jand g2417(.dina(n1721), .dinb(n746), .dout(n3059));
  jand g2418(.dina(n1562), .dinb(n764), .dout(n3060));
  jor  g2419(.dina(n3060), .dinb(n3059), .dout(n3061));
  jand g2420(.dina(n3061), .dinb(n3058), .dout(n3062));
  jand g2421(.dina(n1721), .dinb(n748), .dout(n3063));
  jand g2422(.dina(n1562), .dinb(n762), .dout(n3064));
  jor  g2423(.dina(n3064), .dinb(n3063), .dout(n3065));
  jand g2424(.dina(n2803), .dinb(n1836), .dout(n3066));
  jand g2425(.dina(n2808), .dinb(n1850), .dout(n3067));
  jor  g2426(.dina(n3067), .dinb(n3066), .dout(n3068));
  jnot g2427(.din(n3068), .dout(n3069));
  jand g2428(.dina(n3069), .dinb(n3065), .dout(n3070));
  jand g2429(.dina(n1721), .dinb(n750), .dout(n3071));
  jand g2430(.dina(n1562), .dinb(n755), .dout(n3072));
  jor  g2431(.dina(n3072), .dinb(n3071), .dout(n3073));
  jand g2432(.dina(n2803), .dinb(n1838), .dout(n3074));
  jand g2433(.dina(n2808), .dinb(n1843), .dout(n3075));
  jor  g2434(.dina(n3075), .dinb(n3074), .dout(n3076));
  jnot g2435(.din(n3076), .dout(n3077));
  jand g2436(.dina(n3077), .dinb(n3073), .dout(n3078));
  jor  g2437(.dina(n3078), .dinb(n3070), .dout(n3079));
  jor  g2438(.dina(n3079), .dinb(n3062), .dout(n3080));
  jor  g2439(.dina(n3080), .dinb(n3054), .dout(n3081));
  jand g2440(.dina(n1721), .dinb(n1399), .dout(n3082));
  jand g2441(.dina(n1562), .dinb(n770), .dout(n3083));
  jor  g2442(.dina(n3083), .dinb(n3082), .dout(n3084));
  jand g2443(.dina(n2803), .dinb(n2492), .dout(n3085));
  jand g2444(.dina(n2808), .dinb(n1858), .dout(n3086));
  jor  g2445(.dina(n3086), .dinb(n3085), .dout(n3087));
  jnot g2446(.din(n3087), .dout(n3088));
  jand g2447(.dina(n3088), .dinb(n3084), .dout(n3089));
  jand g2448(.dina(n2803), .dinb(n2494), .dout(n3090));
  jand g2449(.dina(n2808), .dinb(n2507), .dout(n3091));
  jor  g2450(.dina(n3091), .dinb(n3090), .dout(n3092));
  jnot g2451(.din(n3092), .dout(n3093));
  jand g2452(.dina(n1721), .dinb(n1401), .dout(n3094));
  jand g2453(.dina(n1562), .dinb(n1414), .dout(n3095));
  jor  g2454(.dina(n3095), .dinb(n3094), .dout(n3096));
  jand g2455(.dina(n3096), .dinb(n3093), .dout(n3097));
  jor  g2456(.dina(n3097), .dinb(n3089), .dout(n3098));
  jand g2457(.dina(n1721), .dinb(n1406), .dout(n3099));
  jand g2458(.dina(n1562), .dinb(n1412), .dout(n3100));
  jor  g2459(.dina(n3100), .dinb(n3099), .dout(n3101));
  jand g2460(.dina(n2803), .dinb(n2499), .dout(n3102));
  jand g2461(.dina(n2808), .dinb(n2505), .dout(n3103));
  jor  g2462(.dina(n3103), .dinb(n3102), .dout(n3104));
  jnot g2463(.din(n3104), .dout(n3105));
  jand g2464(.dina(n3105), .dinb(n3101), .dout(n3106));
  jand g2465(.dina(n2803), .dinb(n2497), .dout(n3107));
  jand g2466(.dina(n2808), .dinb(n2511), .dout(n3108));
  jor  g2467(.dina(n3108), .dinb(n3107), .dout(n3109));
  jnot g2468(.din(n3109), .dout(n3110));
  jand g2469(.dina(n1721), .dinb(n1404), .dout(n3111));
  jand g2470(.dina(n1562), .dinb(n1418), .dout(n3112));
  jor  g2471(.dina(n3112), .dinb(n3111), .dout(n3113));
  jand g2472(.dina(n3113), .dinb(n3110), .dout(n3114));
  jor  g2473(.dina(n3114), .dinb(n3106), .dout(n3115));
  jor  g2474(.dina(n3115), .dinb(n3098), .dout(n3116));
  jand g2475(.dina(n2803), .dinb(n1861), .dout(n3117));
  jand g2476(.dina(n2808), .dinb(n1879), .dout(n3118));
  jor  g2477(.dina(n3118), .dinb(n3117), .dout(n3119));
  jnot g2478(.din(n3119), .dout(n3120));
  jand g2479(.dina(n1721), .dinb(n773), .dout(n3121));
  jand g2480(.dina(n1562), .dinb(n791), .dout(n3122));
  jor  g2481(.dina(n3122), .dinb(n3121), .dout(n3123));
  jand g2482(.dina(n3123), .dinb(n3120), .dout(n3124));
  jand g2483(.dina(n1721), .dinb(n775), .dout(n3125));
  jand g2484(.dina(n1562), .dinb(n789), .dout(n3126));
  jor  g2485(.dina(n3126), .dinb(n3125), .dout(n3127));
  jand g2486(.dina(n2803), .dinb(n1863), .dout(n3128));
  jand g2487(.dina(n2808), .dinb(n1877), .dout(n3129));
  jor  g2488(.dina(n3129), .dinb(n3128), .dout(n3130));
  jnot g2489(.din(n3130), .dout(n3131));
  jand g2490(.dina(n3131), .dinb(n3127), .dout(n3132));
  jand g2491(.dina(n1721), .dinb(n777), .dout(n3133));
  jand g2492(.dina(n1562), .dinb(n782), .dout(n3134));
  jor  g2493(.dina(n3134), .dinb(n3133), .dout(n3135));
  jand g2494(.dina(n2803), .dinb(n1865), .dout(n3136));
  jand g2495(.dina(n2808), .dinb(n1870), .dout(n3137));
  jor  g2496(.dina(n3137), .dinb(n3136), .dout(n3138));
  jnot g2497(.din(n3138), .dout(n3139));
  jand g2498(.dina(n3139), .dinb(n3135), .dout(n3140));
  jor  g2499(.dina(n3140), .dinb(n3132), .dout(n3141));
  jor  g2500(.dina(n3141), .dinb(n3124), .dout(n3142));
  jnot g2501(.din(n3142), .dout(n3143));
  jnot g2502(.din(n3135), .dout(n3144));
  jand g2503(.dina(n3138), .dinb(n3144), .dout(n3145));
  jand g2504(.dina(n1721), .dinb(n1394), .dout(n3146));
  jand g2505(.dina(n1562), .dinb(n784), .dout(n3147));
  jor  g2506(.dina(n3147), .dinb(n3146), .dout(n3148));
  jnot g2507(.din(n3148), .dout(n3149));
  jand g2508(.dina(n2803), .dinb(n2487), .dout(n3150));
  jand g2509(.dina(n2808), .dinb(n1872), .dout(n3151));
  jor  g2510(.dina(n3151), .dinb(n3150), .dout(n3152));
  jand g2511(.dina(n3152), .dinb(n3149), .dout(n3153));
  jor  g2512(.dina(n3153), .dinb(n3145), .dout(n3154));
  jand g2513(.dina(n3154), .dinb(n3143), .dout(n3155));
  jnot g2514(.din(n3155), .dout(n3156));
  jnot g2515(.din(n3132), .dout(n3157));
  jnot g2516(.din(n3127), .dout(n3158));
  jand g2517(.dina(n3130), .dinb(n3158), .dout(n3159));
  jnot g2518(.din(n3123), .dout(n3160));
  jand g2519(.dina(n3160), .dinb(n3119), .dout(n3161));
  jor  g2520(.dina(n3161), .dinb(n3159), .dout(n3162));
  jand g2521(.dina(n3162), .dinb(n3157), .dout(n3163));
  jnot g2522(.din(n3163), .dout(n3164));
  jand g2523(.dina(n1721), .dinb(n1372), .dout(n3165));
  jand g2524(.dina(n1562), .dinb(n797), .dout(n3166));
  jor  g2525(.dina(n3166), .dinb(n3165), .dout(n3167));
  jnot g2526(.din(n3167), .dout(n3168));
  jand g2527(.dina(n2803), .dinb(n2465), .dout(n3169));
  jand g2528(.dina(n2808), .dinb(n1885), .dout(n3170));
  jor  g2529(.dina(n3170), .dinb(n3169), .dout(n3171));
  jand g2530(.dina(n3171), .dinb(n3168), .dout(n3172));
  jnot g2531(.din(n3172), .dout(n3173));
  jnot g2532(.din(n3171), .dout(n3174));
  jand g2533(.dina(n3174), .dinb(n3167), .dout(n3175));
  jand g2534(.dina(n2803), .dinb(n2467), .dout(n3176));
  jand g2535(.dina(n2808), .dinb(n2475), .dout(n3177));
  jor  g2536(.dina(n3177), .dinb(n3176), .dout(n3178));
  jnot g2537(.din(n3178), .dout(n3179));
  jand g2538(.dina(n1721), .dinb(n1374), .dout(n3180));
  jand g2539(.dina(n1562), .dinb(n1382), .dout(n3181));
  jor  g2540(.dina(n3181), .dinb(n3180), .dout(n3182));
  jand g2541(.dina(n3182), .dinb(n3179), .dout(n3183));
  jor  g2542(.dina(n3183), .dinb(n3175), .dout(n3184));
  jand g2543(.dina(n1721), .dinb(n800), .dout(n3185));
  jand g2544(.dina(n1562), .dinb(n1380), .dout(n3186));
  jor  g2545(.dina(n3186), .dinb(n3185), .dout(n3187));
  jand g2546(.dina(n2803), .dinb(n1888), .dout(n3188));
  jand g2547(.dina(n2808), .dinb(n2473), .dout(n3189));
  jor  g2548(.dina(n3189), .dinb(n3188), .dout(n3190));
  jnot g2549(.din(n3190), .dout(n3191));
  jand g2550(.dina(n3191), .dinb(n3187), .dout(n3192));
  jand g2551(.dina(n2803), .dinb(n1890), .dout(n3193));
  jand g2552(.dina(n2808), .dinb(n2479), .dout(n3194));
  jor  g2553(.dina(n3194), .dinb(n3193), .dout(n3195));
  jnot g2554(.din(n3195), .dout(n3196));
  jand g2555(.dina(n1721), .dinb(n802), .dout(n3197));
  jand g2556(.dina(n1562), .dinb(n1386), .dout(n3198));
  jor  g2557(.dina(n3198), .dinb(n3197), .dout(n3199));
  jand g2558(.dina(n3199), .dinb(n3196), .dout(n3200));
  jor  g2559(.dina(n3200), .dinb(n3192), .dout(n3201));
  jor  g2560(.dina(n3201), .dinb(n3184), .dout(n3202));
  jand g2561(.dina(n1721), .dinb(n1367), .dout(n3203));
  jand g2562(.dina(n1562), .dinb(n816), .dout(n3204));
  jor  g2563(.dina(n3204), .dinb(n3203), .dout(n3205));
  jand g2564(.dina(n2803), .dinb(n2460), .dout(n3206));
  jand g2565(.dina(n2808), .dinb(n1904), .dout(n3207));
  jor  g2566(.dina(n3207), .dinb(n3206), .dout(n3208));
  jnot g2567(.din(n3208), .dout(n3209));
  jand g2568(.dina(n3209), .dinb(n3205), .dout(n3210));
  jand g2569(.dina(n2803), .dinb(n1893), .dout(n3211));
  jand g2570(.dina(n2808), .dinb(n1911), .dout(n3212));
  jor  g2571(.dina(n3212), .dinb(n3211), .dout(n3213));
  jnot g2572(.din(n3213), .dout(n3214));
  jand g2573(.dina(n1721), .dinb(n805), .dout(n3215));
  jand g2574(.dina(n1562), .dinb(n823), .dout(n3216));
  jor  g2575(.dina(n3216), .dinb(n3215), .dout(n3217));
  jand g2576(.dina(n3217), .dinb(n3214), .dout(n3218));
  jand g2577(.dina(n1721), .dinb(n807), .dout(n3219));
  jand g2578(.dina(n1562), .dinb(n821), .dout(n3220));
  jor  g2579(.dina(n3220), .dinb(n3219), .dout(n3221));
  jand g2580(.dina(n2803), .dinb(n1895), .dout(n3222));
  jand g2581(.dina(n2808), .dinb(n1909), .dout(n3223));
  jor  g2582(.dina(n3223), .dinb(n3222), .dout(n3224));
  jnot g2583(.din(n3224), .dout(n3225));
  jand g2584(.dina(n3225), .dinb(n3221), .dout(n3226));
  jand g2585(.dina(n1721), .dinb(n809), .dout(n3227));
  jand g2586(.dina(n1562), .dinb(n814), .dout(n3228));
  jor  g2587(.dina(n3228), .dinb(n3227), .dout(n3229));
  jand g2588(.dina(n2803), .dinb(n1897), .dout(n3230));
  jand g2589(.dina(n2808), .dinb(n1902), .dout(n3231));
  jor  g2590(.dina(n3231), .dinb(n3230), .dout(n3232));
  jnot g2591(.din(n3232), .dout(n3233));
  jand g2592(.dina(n3233), .dinb(n3229), .dout(n3234));
  jor  g2593(.dina(n3234), .dinb(n3226), .dout(n3235));
  jor  g2594(.dina(n3235), .dinb(n3218), .dout(n3236));
  jor  g2595(.dina(n3236), .dinb(n3210), .dout(n3237));
  jand g2596(.dina(n2803), .dinb(n1920), .dout(n3238));
  jand g2597(.dina(n2808), .dinb(n1938), .dout(n3239));
  jor  g2598(.dina(n3239), .dinb(n3238), .dout(n3240));
  jnot g2599(.din(n3240), .dout(n3241));
  jand g2600(.dina(n1721), .dinb(n837), .dout(n3242));
  jand g2601(.dina(n1562), .dinb(n855), .dout(n3243));
  jor  g2602(.dina(n3243), .dinb(n3242), .dout(n3244));
  jand g2603(.dina(n3244), .dinb(n3241), .dout(n3245));
  jand g2604(.dina(n1721), .dinb(n839), .dout(n3246));
  jand g2605(.dina(n1562), .dinb(n853), .dout(n3247));
  jor  g2606(.dina(n3247), .dinb(n3246), .dout(n3248));
  jand g2607(.dina(n2803), .dinb(n1922), .dout(n3249));
  jand g2608(.dina(n2808), .dinb(n1936), .dout(n3250));
  jor  g2609(.dina(n3250), .dinb(n3249), .dout(n3251));
  jnot g2610(.din(n3251), .dout(n3252));
  jand g2611(.dina(n3252), .dinb(n3248), .dout(n3253));
  jand g2612(.dina(n1721), .dinb(n841), .dout(n3254));
  jand g2613(.dina(n1562), .dinb(n846), .dout(n3255));
  jor  g2614(.dina(n3255), .dinb(n3254), .dout(n3256));
  jand g2615(.dina(n2803), .dinb(n1924), .dout(n3257));
  jand g2616(.dina(n2808), .dinb(n1929), .dout(n3258));
  jor  g2617(.dina(n3258), .dinb(n3257), .dout(n3259));
  jnot g2618(.din(n3259), .dout(n3260));
  jand g2619(.dina(n3260), .dinb(n3256), .dout(n3261));
  jor  g2620(.dina(n3261), .dinb(n3253), .dout(n3262));
  jor  g2621(.dina(n3262), .dinb(n3245), .dout(n3263));
  jnot g2622(.din(n3263), .dout(n3264));
  jnot g2623(.din(n3256), .dout(n3265));
  jand g2624(.dina(n3259), .dinb(n3265), .dout(n3266));
  jand g2625(.dina(n1721), .dinb(n1340), .dout(n3267));
  jand g2626(.dina(n1562), .dinb(n848), .dout(n3268));
  jor  g2627(.dina(n3268), .dinb(n3267), .dout(n3269));
  jnot g2628(.din(n3269), .dout(n3270));
  jand g2629(.dina(n2803), .dinb(n2428), .dout(n3271));
  jand g2630(.dina(n2808), .dinb(n1931), .dout(n3272));
  jor  g2631(.dina(n3272), .dinb(n3271), .dout(n3273));
  jand g2632(.dina(n3273), .dinb(n3270), .dout(n3274));
  jor  g2633(.dina(n3274), .dinb(n3266), .dout(n3275));
  jand g2634(.dina(n3275), .dinb(n3264), .dout(n3276));
  jnot g2635(.din(n3253), .dout(n3277));
  jnot g2636(.din(n3248), .dout(n3278));
  jand g2637(.dina(n3251), .dinb(n3278), .dout(n3279));
  jnot g2638(.din(n3244), .dout(n3280));
  jand g2639(.dina(n3280), .dinb(n3240), .dout(n3281));
  jor  g2640(.dina(n3281), .dinb(n3279), .dout(n3282));
  jand g2641(.dina(n3282), .dinb(n3277), .dout(n3283));
  jor  g2642(.dina(n3283), .dinb(n3276), .dout(n3284));
  jnot g2643(.din(n3284), .dout(n3285));
  jand g2644(.dina(n1721), .dinb(n1333), .dout(n3286));
  jand g2645(.dina(n1562), .dinb(n861), .dout(n3287));
  jor  g2646(.dina(n3287), .dinb(n3286), .dout(n3288));
  jnot g2647(.din(n3288), .dout(n3289));
  jand g2648(.dina(n2803), .dinb(n2421), .dout(n3290));
  jand g2649(.dina(n2808), .dinb(n1944), .dout(n3291));
  jor  g2650(.dina(n3291), .dinb(n3290), .dout(n3292));
  jand g2651(.dina(n3292), .dinb(n3289), .dout(n3293));
  jnot g2652(.din(n3293), .dout(n3294));
  jand g2653(.dina(n2803), .dinb(n2423), .dout(n3295));
  jand g2654(.dina(n2808), .dinb(n1953), .dout(n3296));
  jor  g2655(.dina(n3296), .dinb(n3295), .dout(n3297));
  jand g2656(.dina(n1721), .dinb(n1335), .dout(n3298));
  jand g2657(.dina(n1562), .dinb(n870), .dout(n3299));
  jor  g2658(.dina(n3299), .dinb(n3298), .dout(n3300));
  jnot g2659(.din(n3300), .dout(n3301));
  jand g2660(.dina(n3301), .dinb(n3297), .dout(n3302));
  jand g2661(.dina(n1721), .dinb(n864), .dout(n3303));
  jand g2662(.dina(n1562), .dinb(n872), .dout(n3304));
  jor  g2663(.dina(n3304), .dinb(n3303), .dout(n3305));
  jnot g2664(.din(n3305), .dout(n3306));
  jand g2665(.dina(n2803), .dinb(n1947), .dout(n3307));
  jand g2666(.dina(n2808), .dinb(n1955), .dout(n3308));
  jor  g2667(.dina(n3308), .dinb(n3307), .dout(n3309));
  jand g2668(.dina(n3309), .dinb(n3306), .dout(n3310));
  jnot g2669(.din(n3309), .dout(n3311));
  jand g2670(.dina(n3311), .dinb(n3305), .dout(n3312));
  jnot g2671(.din(n3312), .dout(n3313));
  jand g2672(.dina(n2803), .dinb(n2416), .dout(n3314));
  jand g2673(.dina(n2808), .dinb(n1950), .dout(n3315));
  jor  g2674(.dina(n3315), .dinb(n3314), .dout(n3316));
  jand g2675(.dina(n1721), .dinb(n1328), .dout(n3317));
  jand g2676(.dina(n1562), .dinb(n867), .dout(n3318));
  jor  g2677(.dina(n3318), .dinb(n3317), .dout(n3319));
  jnot g2678(.din(n3319), .dout(n3320));
  jand g2679(.dina(n3320), .dinb(n3316), .dout(n3321));
  jand g2680(.dina(n3321), .dinb(n3313), .dout(n3322));
  jor  g2681(.dina(n3322), .dinb(n3310), .dout(n3323));
  jor  g2682(.dina(n3323), .dinb(n3302), .dout(n3324));
  jnot g2683(.din(n3324), .dout(n3325));
  jand g2684(.dina(n1721), .dinb(n878), .dout(n3326));
  jand g2685(.dina(n1562), .dinb(n1312), .dout(n3327));
  jor  g2686(.dina(n3327), .dinb(n3326), .dout(n3328));
  jand g2687(.dina(n2803), .dinb(n1961), .dout(n3329));
  jand g2688(.dina(n2808), .dinb(n2400), .dout(n3330));
  jor  g2689(.dina(n3330), .dinb(n3329), .dout(n3331));
  jnot g2690(.din(n3331), .dout(n3332));
  jand g2691(.dina(n3332), .dinb(n3328), .dout(n3333));
  jand g2692(.dina(n2803), .dinb(n1967), .dout(n3334));
  jand g2693(.dina(n2808), .dinb(n2407), .dout(n3335));
  jor  g2694(.dina(n3335), .dinb(n3334), .dout(n3336));
  jnot g2695(.din(n3336), .dout(n3337));
  jand g2696(.dina(n1721), .dinb(n884), .dout(n3338));
  jand g2697(.dina(n1562), .dinb(n1319), .dout(n3339));
  jor  g2698(.dina(n3339), .dinb(n3338), .dout(n3340));
  jand g2699(.dina(n3340), .dinb(n3337), .dout(n3341));
  jand g2700(.dina(n1721), .dinb(n880), .dout(n3342));
  jand g2701(.dina(n1562), .dinb(n1317), .dout(n3343));
  jor  g2702(.dina(n3343), .dinb(n3342), .dout(n3344));
  jand g2703(.dina(n2803), .dinb(n1963), .dout(n3345));
  jand g2704(.dina(n2808), .dinb(n2405), .dout(n3346));
  jor  g2705(.dina(n3346), .dinb(n3345), .dout(n3347));
  jnot g2706(.din(n3347), .dout(n3348));
  jand g2707(.dina(n3348), .dinb(n3344), .dout(n3349));
  jand g2708(.dina(n1721), .dinb(n882), .dout(n3350));
  jand g2709(.dina(n1562), .dinb(n1310), .dout(n3351));
  jor  g2710(.dina(n3351), .dinb(n3350), .dout(n3352));
  jand g2711(.dina(n2803), .dinb(n1965), .dout(n3353));
  jand g2712(.dina(n2808), .dinb(n2398), .dout(n3354));
  jor  g2713(.dina(n3354), .dinb(n3353), .dout(n3355));
  jnot g2714(.din(n3355), .dout(n3356));
  jand g2715(.dina(n3356), .dinb(n3352), .dout(n3357));
  jor  g2716(.dina(n3357), .dinb(n3349), .dout(n3358));
  jor  g2717(.dina(n3358), .dinb(n3341), .dout(n3359));
  jor  g2718(.dina(n3359), .dinb(n3333), .dout(n3360));
  jnot g2719(.din(n3360), .dout(n3361));
  jand g2720(.dina(n1721), .dinb(n1290), .dout(n3362));
  jand g2721(.dina(n1562), .dinb(n877), .dout(n3363));
  jor  g2722(.dina(n3363), .dinb(n3362), .dout(n3364));
  jnot g2723(.din(n3364), .dout(n3365));
  jand g2724(.dina(n2803), .dinb(n2378), .dout(n3366));
  jand g2725(.dina(n2808), .dinb(n1960), .dout(n3367));
  jor  g2726(.dina(n3367), .dinb(n3366), .dout(n3368));
  jand g2727(.dina(n3368), .dinb(n3365), .dout(n3369));
  jnot g2728(.din(n3368), .dout(n3370));
  jand g2729(.dina(n3370), .dinb(n3364), .dout(n3371));
  jand g2730(.dina(n1721), .dinb(n1288), .dout(n3372));
  jand g2731(.dina(n1562), .dinb(n1301), .dout(n3373));
  jor  g2732(.dina(n3373), .dinb(n3372), .dout(n3374));
  jand g2733(.dina(n2803), .dinb(n2376), .dout(n3375));
  jand g2734(.dina(n2808), .dinb(n2389), .dout(n3376));
  jor  g2735(.dina(n3376), .dinb(n3375), .dout(n3377));
  jnot g2736(.din(n3377), .dout(n3378));
  jand g2737(.dina(n3378), .dinb(n3374), .dout(n3379));
  jor  g2738(.dina(n3379), .dinb(n3371), .dout(n3380));
  jnot g2739(.din(n3380), .dout(n3381));
  jnot g2740(.din(n3374), .dout(n3382));
  jand g2741(.dina(n3377), .dinb(n3382), .dout(n3383));
  jand g2742(.dina(n1721), .dinb(n1285), .dout(n3384));
  jand g2743(.dina(n1562), .dinb(n1299), .dout(n3385));
  jor  g2744(.dina(n3385), .dinb(n3384), .dout(n3386));
  jand g2745(.dina(n2803), .dinb(n2373), .dout(n3387));
  jand g2746(.dina(n2808), .dinb(n2387), .dout(n3388));
  jor  g2747(.dina(n3388), .dinb(n3387), .dout(n3389));
  jnot g2748(.din(n3389), .dout(n3390));
  jand g2749(.dina(n3390), .dinb(n3386), .dout(n3391));
  jnot g2750(.din(n3391), .dout(n3392));
  jand g2751(.dina(n1721), .dinb(n1282), .dout(n3393));
  jand g2752(.dina(n1562), .dinb(n1304), .dout(n3394));
  jor  g2753(.dina(n3394), .dinb(n3393), .dout(n3395));
  jnot g2754(.din(n3395), .dout(n3396));
  jand g2755(.dina(n2803), .dinb(n2370), .dout(n3397));
  jand g2756(.dina(n2808), .dinb(n2392), .dout(n3398));
  jor  g2757(.dina(n3398), .dinb(n3397), .dout(n3399));
  jand g2758(.dina(n3399), .dinb(n3396), .dout(n3400));
  jand g2759(.dina(n3400), .dinb(n3392), .dout(n3401));
  jnot g2760(.din(n3386), .dout(n3402));
  jand g2761(.dina(n3389), .dinb(n3402), .dout(n3403));
  jor  g2762(.dina(n3403), .dinb(n3401), .dout(n3404));
  jor  g2763(.dina(n3404), .dinb(n3383), .dout(n3405));
  jand g2764(.dina(n3405), .dinb(n3381), .dout(n3406));
  jor  g2765(.dina(n3406), .dinb(n3369), .dout(n3407));
  jand g2766(.dina(n3407), .dinb(n3361), .dout(n3408));
  jnot g2767(.din(n3408), .dout(n3409));
  jand g2768(.dina(n1721), .dinb(n896), .dout(n3410));
  jand g2769(.dina(n1562), .dinb(n1263), .dout(n3411));
  jor  g2770(.dina(n3411), .dinb(n3410), .dout(n3412));
  jnot g2771(.din(n3412), .dout(n3413));
  jand g2772(.dina(n2803), .dinb(n1979), .dout(n3414));
  jand g2773(.dina(n2808), .dinb(n2351), .dout(n3415));
  jor  g2774(.dina(n3415), .dinb(n3414), .dout(n3416));
  jand g2775(.dina(n3416), .dinb(n3413), .dout(n3417));
  jnot g2776(.din(n3417), .dout(n3418));
  jand g2777(.dina(n2803), .dinb(n2286), .dout(n3419));
  jand g2778(.dina(n2808), .dinb(n1992), .dout(n3420));
  jor  g2779(.dina(n3420), .dinb(n3419), .dout(n3421));
  jand g2780(.dina(n1721), .dinb(n909), .dout(n3422));
  jand g2781(.dina(n1562), .dinb(n1218), .dout(n3423));
  jor  g2782(.dina(n3423), .dinb(n3422), .dout(n3424));
  jand g2783(.dina(n2803), .dinb(n1993), .dout(n3425));
  jand g2784(.dina(n2808), .dinb(n2308), .dout(n3426));
  jor  g2785(.dina(n3426), .dinb(n3425), .dout(n3427));
  jnot g2786(.din(n3427), .dout(n3428));
  jand g2787(.dina(n3428), .dinb(n3424), .dout(n3429));
  jnot g2788(.din(n3429), .dout(n3430));
  jand g2789(.dina(n1721), .dinb(n911), .dout(n3431));
  jand g2790(.dina(n1562), .dinb(n1223), .dout(n3432));
  jor  g2791(.dina(n3432), .dinb(n3431), .dout(n3433));
  jand g2792(.dina(n2803), .dinb(n1995), .dout(n3434));
  jand g2793(.dina(n2808), .dinb(n2313), .dout(n3435));
  jor  g2794(.dina(n3435), .dinb(n3434), .dout(n3436));
  jnot g2795(.din(n3436), .dout(n3437));
  jand g2796(.dina(n3437), .dinb(n3433), .dout(n3438));
  jand g2797(.dina(n2803), .dinb(n1999), .dout(n3439));
  jand g2798(.dina(n2808), .dinb(n2315), .dout(n3440));
  jor  g2799(.dina(n3440), .dinb(n3439), .dout(n3441));
  jnot g2800(.din(n3441), .dout(n3442));
  jand g2801(.dina(n1721), .dinb(n915), .dout(n3443));
  jand g2802(.dina(n1562), .dinb(n1225), .dout(n3444));
  jor  g2803(.dina(n3444), .dinb(n3443), .dout(n3445));
  jand g2804(.dina(n3445), .dinb(n3442), .dout(n3446));
  jor  g2805(.dina(n3446), .dinb(n3438), .dout(n3447));
  jnot g2806(.din(n3447), .dout(n3448));
  jand g2807(.dina(n1721), .dinb(n913), .dout(n3449));
  jand g2808(.dina(n1562), .dinb(n1216), .dout(n3450));
  jor  g2809(.dina(n3450), .dinb(n3449), .dout(n3451));
  jand g2810(.dina(n2803), .dinb(n1997), .dout(n3452));
  jand g2811(.dina(n2808), .dinb(n2306), .dout(n3453));
  jor  g2812(.dina(n3453), .dinb(n3452), .dout(n3454));
  jnot g2813(.din(n3454), .dout(n3455));
  jand g2814(.dina(n3455), .dinb(n3451), .dout(n3456));
  jnot g2815(.din(n3456), .dout(n3457));
  jand g2816(.dina(n3457), .dinb(n3448), .dout(n3458));
  jand g2817(.dina(n3458), .dinb(n3430), .dout(n3459));
  jand g2818(.dina(n1721), .dinb(n922), .dout(n3460));
  jnot g2819(.din(n3460), .dout(n3461));
  jor  g2820(.dina(n1721), .dinb(\in1[43] ), .dout(n3462));
  jand g2821(.dina(n3462), .dinb(n3461), .dout(n3463));
  jand g2822(.dina(n3463), .dinb(n3459), .dout(n3464));
  jand g2823(.dina(n3464), .dinb(n3421), .dout(n3465));
  jnot g2824(.din(n3465), .dout(n3466));
  jand g2825(.dina(n1721), .dinb(n962), .dout(n3467));
  jand g2826(.dina(n1562), .dinb(n1198), .dout(n3468));
  jor  g2827(.dina(n3468), .dinb(n3467), .dout(n3469));
  jand g2828(.dina(n2803), .dinb(n2029), .dout(n3470));
  jand g2829(.dina(n2808), .dinb(n2266), .dout(n3471));
  jor  g2830(.dina(n3471), .dinb(n3470), .dout(n3472));
  jnot g2831(.din(n3472), .dout(n3473));
  jand g2832(.dina(n3473), .dinb(n3469), .dout(n3474));
  jnot g2833(.din(n3474), .dout(n3475));
  jand g2834(.dina(n2803), .dinb(n2027), .dout(n3476));
  jand g2835(.dina(n2808), .dinb(n2269), .dout(n3477));
  jor  g2836(.dina(n3477), .dinb(n3476), .dout(n3478));
  jnot g2837(.din(n3478), .dout(n3479));
  jand g2838(.dina(n1721), .dinb(n960), .dout(n3480));
  jand g2839(.dina(n1562), .dinb(n1201), .dout(n3481));
  jor  g2840(.dina(n3481), .dinb(n3480), .dout(n3482));
  jand g2841(.dina(n3482), .dinb(n3479), .dout(n3483));
  jand g2842(.dina(n1721), .dinb(n964), .dout(n3484));
  jand g2843(.dina(n1562), .dinb(n1188), .dout(n3485));
  jor  g2844(.dina(n3485), .dinb(n3484), .dout(n3486));
  jand g2845(.dina(n2803), .dinb(n2031), .dout(n3487));
  jand g2846(.dina(n2808), .dinb(n2256), .dout(n3488));
  jor  g2847(.dina(n3488), .dinb(n3487), .dout(n3489));
  jnot g2848(.din(n3489), .dout(n3490));
  jand g2849(.dina(n3490), .dinb(n3486), .dout(n3491));
  jor  g2850(.dina(n3491), .dinb(n3483), .dout(n3492));
  jnot g2851(.din(n3492), .dout(n3493));
  jnot g2852(.din(n3486), .dout(n3494));
  jand g2853(.dina(n3489), .dinb(n3494), .dout(n3495));
  jand g2854(.dina(n1721), .dinb(n958), .dout(n3496));
  jand g2855(.dina(n1562), .dinb(n1190), .dout(n3497));
  jor  g2856(.dina(n3497), .dinb(n3496), .dout(n3498));
  jnot g2857(.din(n3498), .dout(n3499));
  jand g2858(.dina(n2803), .dinb(n2025), .dout(n3500));
  jand g2859(.dina(n2808), .dinb(n2258), .dout(n3501));
  jor  g2860(.dina(n3501), .dinb(n3500), .dout(n3502));
  jand g2861(.dina(n3502), .dinb(n3499), .dout(n3503));
  jor  g2862(.dina(n3503), .dinb(n3495), .dout(n3504));
  jnot g2863(.din(n3502), .dout(n3505));
  jand g2864(.dina(n3505), .dinb(n3498), .dout(n3506));
  jnot g2865(.din(n3506), .dout(n3507));
  jand g2866(.dina(n1721), .dinb(n953), .dout(n3508));
  jand g2867(.dina(n1562), .dinb(n1195), .dout(n3509));
  jor  g2868(.dina(n3509), .dinb(n3508), .dout(n3510));
  jand g2869(.dina(n2803), .dinb(n2020), .dout(n3511));
  jand g2870(.dina(n2808), .dinb(n2263), .dout(n3512));
  jor  g2871(.dina(n3512), .dinb(n3511), .dout(n3513));
  jnot g2872(.din(n3513), .dout(n3514));
  jand g2873(.dina(n3514), .dinb(n3510), .dout(n3515));
  jnot g2874(.din(n3515), .dout(n3516));
  jand g2875(.dina(n1721), .dinb(n946), .dout(n3517));
  jand g2876(.dina(n1562), .dinb(n941), .dout(n3518));
  jor  g2877(.dina(n3518), .dinb(n3517), .dout(n3519));
  jand g2878(.dina(n2803), .dinb(n2013), .dout(n3520));
  jand g2879(.dina(n2808), .dinb(n2008), .dout(n3521));
  jor  g2880(.dina(n3521), .dinb(n3520), .dout(n3522));
  jnot g2881(.din(n3522), .dout(n3523));
  jand g2882(.dina(n3523), .dinb(n3519), .dout(n3524));
  jand g2883(.dina(n2803), .dinb(n2022), .dout(n3525));
  jand g2884(.dina(n2808), .dinb(n2010), .dout(n3526));
  jor  g2885(.dina(n3526), .dinb(n3525), .dout(n3527));
  jnot g2886(.din(n3527), .dout(n3528));
  jand g2887(.dina(n1721), .dinb(n955), .dout(n3529));
  jand g2888(.dina(n1562), .dinb(n943), .dout(n3530));
  jor  g2889(.dina(n3530), .dinb(n3529), .dout(n3531));
  jand g2890(.dina(n3531), .dinb(n3528), .dout(n3532));
  jor  g2891(.dina(n3532), .dinb(n3524), .dout(n3533));
  jnot g2892(.din(n3533), .dout(n3534));
  jand g2893(.dina(n2803), .dinb(n2249), .dout(n3535));
  jand g2894(.dina(n2808), .dinb(n2016), .dout(n3536));
  jor  g2895(.dina(n3536), .dinb(n3535), .dout(n3537));
  jand g2896(.dina(n1721), .dinb(n1181), .dout(n3538));
  jand g2897(.dina(n1562), .dinb(n949), .dout(n3539));
  jor  g2898(.dina(n3539), .dinb(n3538), .dout(n3540));
  jnot g2899(.din(n3540), .dout(n3541));
  jand g2900(.dina(n3541), .dinb(n3537), .dout(n3542));
  jnot g2901(.din(n3519), .dout(n3543));
  jand g2902(.dina(n3522), .dinb(n3543), .dout(n3544));
  jor  g2903(.dina(n3544), .dinb(n3542), .dout(n3545));
  jand g2904(.dina(n3545), .dinb(n3534), .dout(n3546));
  jnot g2905(.din(n3510), .dout(n3547));
  jand g2906(.dina(n3513), .dinb(n3547), .dout(n3548));
  jnot g2907(.din(n3531), .dout(n3549));
  jand g2908(.dina(n3549), .dinb(n3527), .dout(n3550));
  jor  g2909(.dina(n3550), .dinb(n3548), .dout(n3551));
  jor  g2910(.dina(n3551), .dinb(n3546), .dout(n3552));
  jand g2911(.dina(n3552), .dinb(n3516), .dout(n3553));
  jand g2912(.dina(n3553), .dinb(n3507), .dout(n3554));
  jor  g2913(.dina(n3554), .dinb(n3504), .dout(n3555));
  jand g2914(.dina(n3555), .dinb(n3493), .dout(n3556));
  jnot g2915(.din(n3469), .dout(n3557));
  jand g2916(.dina(n3472), .dinb(n3557), .dout(n3558));
  jnot g2917(.din(n3482), .dout(n3559));
  jand g2918(.dina(n3559), .dinb(n3478), .dout(n3560));
  jor  g2919(.dina(n3560), .dinb(n3558), .dout(n3561));
  jor  g2920(.dina(n3561), .dinb(n3556), .dout(n3562));
  jand g2921(.dina(n3562), .dinb(n3475), .dout(n3563));
  jnot g2922(.din(n3563), .dout(n3564));
  jand g2923(.dina(n1721), .dinb(n1179), .dout(n3565));
  jand g2924(.dina(n1562), .dinb(n1172), .dout(n3566));
  jor  g2925(.dina(n3566), .dinb(n3565), .dout(n3567));
  jnot g2926(.din(n3567), .dout(n3568));
  jand g2927(.dina(n2803), .dinb(n2247), .dout(n3569));
  jand g2928(.dina(n2808), .dinb(n2240), .dout(n3570));
  jor  g2929(.dina(n3570), .dinb(n3569), .dout(n3571));
  jand g2930(.dina(n3571), .dinb(n3568), .dout(n3572));
  jnot g2931(.din(n3572), .dout(n3573));
  jand g2932(.dina(n1721), .dinb(n978), .dout(n3574));
  jand g2933(.dina(n1562), .dinb(n975), .dout(n3575));
  jor  g2934(.dina(n3575), .dinb(n3574), .dout(n3576));
  jand g2935(.dina(n2803), .dinb(n2045), .dout(n3577));
  jand g2936(.dina(n2808), .dinb(n2042), .dout(n3578));
  jor  g2937(.dina(n3578), .dinb(n3577), .dout(n3579));
  jnot g2938(.din(n3579), .dout(n3580));
  jand g2939(.dina(n3580), .dinb(n3576), .dout(n3581));
  jand g2940(.dina(n1721), .dinb(n983), .dout(n3582));
  jand g2941(.dina(n1562), .dinb(n980), .dout(n3583));
  jor  g2942(.dina(n3583), .dinb(n3582), .dout(n3584));
  jnot g2943(.din(n3584), .dout(n3585));
  jand g2944(.dina(n2803), .dinb(n2050), .dout(n3586));
  jand g2945(.dina(n2808), .dinb(n2047), .dout(n3587));
  jor  g2946(.dina(n3587), .dinb(n3586), .dout(n3588));
  jand g2947(.dina(n3588), .dinb(n3585), .dout(n3589));
  jnot g2948(.din(n3589), .dout(n3590));
  jand g2949(.dina(n1721), .dinb(n1158), .dout(n3591));
  jand g2950(.dina(n1562), .dinb(n990), .dout(n3592));
  jor  g2951(.dina(n3592), .dinb(n3591), .dout(n3593));
  jand g2952(.dina(n2803), .dinb(n2226), .dout(n3594));
  jand g2953(.dina(n2808), .dinb(n2057), .dout(n3595));
  jor  g2954(.dina(n3595), .dinb(n3594), .dout(n3596));
  jnot g2955(.din(n3596), .dout(n3597));
  jand g2956(.dina(n3597), .dinb(n3593), .dout(n3598));
  jand g2957(.dina(n2803), .dinb(n2215), .dout(n3599));
  jand g2958(.dina(n2808), .dinb(n2219), .dout(n3600));
  jor  g2959(.dina(n3600), .dinb(n3599), .dout(n3601));
  jand g2960(.dina(n1721), .dinb(n1147), .dout(n3602));
  jand g2961(.dina(n1562), .dinb(n1151), .dout(n3603));
  jor  g2962(.dina(n3603), .dinb(n3602), .dout(n3604));
  jnot g2963(.din(n3604), .dout(n3605));
  jand g2964(.dina(n3605), .dinb(n3601), .dout(n3606));
  jand g2965(.dina(n2803), .dinb(n2228), .dout(n3607));
  jand g2966(.dina(n2808), .dinb(n2221), .dout(n3608));
  jor  g2967(.dina(n3608), .dinb(n3607), .dout(n3609));
  jand g2968(.dina(n1721), .dinb(n1160), .dout(n3610));
  jand g2969(.dina(n1562), .dinb(n1153), .dout(n3611));
  jor  g2970(.dina(n3611), .dinb(n3610), .dout(n3612));
  jnot g2971(.din(n3612), .dout(n3613));
  jand g2972(.dina(n3613), .dinb(n3609), .dout(n3614));
  jor  g2973(.dina(n3614), .dinb(n3606), .dout(n3615));
  jnot g2974(.din(n3615), .dout(n3616));
  jand g2975(.dina(n1721), .dinb(n993), .dout(n3617));
  jand g2976(.dina(n1562), .dinb(n1140), .dout(n3618));
  jor  g2977(.dina(n3618), .dinb(n3617), .dout(n3619));
  jnot g2978(.din(n3619), .dout(n3620));
  jand g2979(.dina(n2803), .dinb(n2060), .dout(n3621));
  jand g2980(.dina(n2808), .dinb(n2208), .dout(n3622));
  jor  g2981(.dina(n3622), .dinb(n3621), .dout(n3623));
  jand g2982(.dina(n3623), .dinb(n3620), .dout(n3624));
  jnot g2983(.din(n3624), .dout(n3625));
  jand g2984(.dina(n1721), .dinb(n995), .dout(n3626));
  jand g2985(.dina(n1562), .dinb(n1142), .dout(n3627));
  jor  g2986(.dina(n3627), .dinb(n3626), .dout(n3628));
  jand g2987(.dina(n2803), .dinb(n2062), .dout(n3629));
  jand g2988(.dina(n2808), .dinb(n2210), .dout(n3630));
  jor  g2989(.dina(n3630), .dinb(n3629), .dout(n3631));
  jnot g2990(.din(n3631), .dout(n3632));
  jand g2991(.dina(n3632), .dinb(n3628), .dout(n3633));
  jand g2992(.dina(n1721), .dinb(n1005), .dout(n3634));
  jand g2993(.dina(n1562), .dinb(n1002), .dout(n3635));
  jor  g2994(.dina(n3635), .dinb(n3634), .dout(n3636));
  jand g2995(.dina(n2803), .dinb(n2072), .dout(n3637));
  jand g2996(.dina(n2808), .dinb(n2069), .dout(n3638));
  jor  g2997(.dina(n3638), .dinb(n3637), .dout(n3639));
  jnot g2998(.din(n3639), .dout(n3640));
  jand g2999(.dina(n3640), .dinb(n3636), .dout(n3641));
  jnot g3000(.din(n3636), .dout(n3642));
  jand g3001(.dina(n3639), .dinb(n3642), .dout(n3643));
  jnot g3002(.din(n3643), .dout(n3644));
  jand g3003(.dina(n1721), .dinb(n1010), .dout(n3645));
  jand g3004(.dina(n1562), .dinb(n1007), .dout(n3646));
  jor  g3005(.dina(n3646), .dinb(n3645), .dout(n3647));
  jand g3006(.dina(n2803), .dinb(n2077), .dout(n3648));
  jand g3007(.dina(n2808), .dinb(n2074), .dout(n3649));
  jor  g3008(.dina(n3649), .dinb(n3648), .dout(n3650));
  jnot g3009(.din(n3650), .dout(n3651));
  jand g3010(.dina(n3651), .dinb(n3647), .dout(n3652));
  jand g3011(.dina(n1721), .dinb(n1126), .dout(n3653));
  jand g3012(.dina(n1562), .dinb(n1012), .dout(n3654));
  jor  g3013(.dina(n3654), .dinb(n3653), .dout(n3655));
  jand g3014(.dina(n2803), .dinb(n2194), .dout(n3656));
  jand g3015(.dina(n2808), .dinb(n2079), .dout(n3657));
  jor  g3016(.dina(n3657), .dinb(n3656), .dout(n3658));
  jnot g3017(.din(n3658), .dout(n3659));
  jand g3018(.dina(n3659), .dinb(n3655), .dout(n3660));
  jand g3019(.dina(n2803), .dinb(n2183), .dout(n3661));
  jand g3020(.dina(n2808), .dinb(n2187), .dout(n3662));
  jor  g3021(.dina(n3662), .dinb(n3661), .dout(n3663));
  jand g3022(.dina(n1721), .dinb(n1115), .dout(n3664));
  jand g3023(.dina(n1562), .dinb(n1119), .dout(n3665));
  jor  g3024(.dina(n3665), .dinb(n3664), .dout(n3666));
  jnot g3025(.din(n3666), .dout(n3667));
  jand g3026(.dina(n3667), .dinb(n3663), .dout(n3668));
  jnot g3027(.din(n3668), .dout(n3669));
  jand g3028(.dina(n1721), .dinb(n1015), .dout(n3670));
  jand g3029(.dina(n1562), .dinb(n1108), .dout(n3671));
  jor  g3030(.dina(n3671), .dinb(n3670), .dout(n3672));
  jand g3031(.dina(n2803), .dinb(n2082), .dout(n3673));
  jand g3032(.dina(n2808), .dinb(n2176), .dout(n3674));
  jor  g3033(.dina(n3674), .dinb(n3673), .dout(n3675));
  jnot g3034(.din(n3675), .dout(n3676));
  jand g3035(.dina(n3676), .dinb(n3672), .dout(n3677));
  jand g3036(.dina(n1721), .dinb(n1017), .dout(n3678));
  jand g3037(.dina(n1562), .dinb(n1110), .dout(n3679));
  jor  g3038(.dina(n3679), .dinb(n3678), .dout(n3680));
  jand g3039(.dina(n2803), .dinb(n2084), .dout(n3681));
  jand g3040(.dina(n2808), .dinb(n2178), .dout(n3682));
  jor  g3041(.dina(n3682), .dinb(n3681), .dout(n3683));
  jnot g3042(.din(n3683), .dout(n3684));
  jand g3043(.dina(n3684), .dinb(n3680), .dout(n3685));
  jand g3044(.dina(n1721), .dinb(n1022), .dout(n3686));
  jand g3045(.dina(n1562), .dinb(n1019), .dout(n3687));
  jor  g3046(.dina(n3687), .dinb(n3686), .dout(n3688));
  jnot g3047(.din(n3688), .dout(n3689));
  jand g3048(.dina(n2803), .dinb(n2089), .dout(n3690));
  jand g3049(.dina(n2808), .dinb(n2086), .dout(n3691));
  jor  g3050(.dina(n3691), .dinb(n3690), .dout(n3692));
  jand g3051(.dina(n3692), .dinb(n3689), .dout(n3693));
  jnot g3052(.din(n3693), .dout(n3694));
  jnot g3053(.din(n3692), .dout(n3695));
  jand g3054(.dina(n3695), .dinb(n3688), .dout(n3696));
  jand g3055(.dina(n1721), .dinb(n1027), .dout(n3697));
  jand g3056(.dina(n1562), .dinb(n1024), .dout(n3698));
  jor  g3057(.dina(n3698), .dinb(n3697), .dout(n3699));
  jnot g3058(.din(n3699), .dout(n3700));
  jand g3059(.dina(n2803), .dinb(n2094), .dout(n3701));
  jand g3060(.dina(n2808), .dinb(n2091), .dout(n3702));
  jor  g3061(.dina(n3702), .dinb(n3701), .dout(n3703));
  jand g3062(.dina(n3703), .dinb(n3700), .dout(n3704));
  jnot g3063(.din(n3704), .dout(n3705));
  jand g3064(.dina(n1721), .dinb(n1094), .dout(n3706));
  jand g3065(.dina(n1562), .dinb(n1034), .dout(n3707));
  jor  g3066(.dina(n3707), .dinb(n3706), .dout(n3708));
  jand g3067(.dina(n2803), .dinb(n2162), .dout(n3709));
  jand g3068(.dina(n2808), .dinb(n2101), .dout(n3710));
  jor  g3069(.dina(n3710), .dinb(n3709), .dout(n3711));
  jnot g3070(.din(n3711), .dout(n3712));
  jand g3071(.dina(n3712), .dinb(n3708), .dout(n3713));
  jand g3072(.dina(n2803), .dinb(n2151), .dout(n3714));
  jand g3073(.dina(n2808), .dinb(n2155), .dout(n3715));
  jor  g3074(.dina(n3715), .dinb(n3714), .dout(n3716));
  jand g3075(.dina(n1721), .dinb(n1083), .dout(n3717));
  jand g3076(.dina(n1562), .dinb(n1087), .dout(n3718));
  jor  g3077(.dina(n3718), .dinb(n3717), .dout(n3719));
  jnot g3078(.din(n3719), .dout(n3720));
  jand g3079(.dina(n3720), .dinb(n3716), .dout(n3721));
  jnot g3080(.din(n3721), .dout(n3722));
  jand g3081(.dina(n1721), .dinb(n1037), .dout(n3723));
  jand g3082(.dina(n1562), .dinb(n1076), .dout(n3724));
  jor  g3083(.dina(n3724), .dinb(n3723), .dout(n3725));
  jand g3084(.dina(n2803), .dinb(n2104), .dout(n3726));
  jand g3085(.dina(n2808), .dinb(n2144), .dout(n3727));
  jor  g3086(.dina(n3727), .dinb(n3726), .dout(n3728));
  jnot g3087(.din(n3728), .dout(n3729));
  jand g3088(.dina(n3729), .dinb(n3725), .dout(n3730));
  jand g3089(.dina(n2803), .dinb(n2138), .dout(n3731));
  jand g3090(.dina(n2808), .dinb(n2146), .dout(n3732));
  jor  g3091(.dina(n3732), .dinb(n3731), .dout(n3733));
  jnot g3092(.din(n3733), .dout(n3734));
  jand g3093(.dina(n1721), .dinb(n1070), .dout(n3735));
  jand g3094(.dina(n1562), .dinb(n1078), .dout(n3736));
  jor  g3095(.dina(n3736), .dinb(n3735), .dout(n3737));
  jand g3096(.dina(n3737), .dinb(n3734), .dout(n3738));
  jand g3097(.dina(n2803), .dinb(n2140), .dout(n3739));
  jand g3098(.dina(n2808), .dinb(n2133), .dout(n3740));
  jor  g3099(.dina(n3740), .dinb(n3739), .dout(n3741));
  jand g3100(.dina(n1721), .dinb(n1072), .dout(n3742));
  jand g3101(.dina(n1562), .dinb(n1065), .dout(n3743));
  jor  g3102(.dina(n3743), .dinb(n3742), .dout(n3744));
  jnot g3103(.din(n3744), .dout(n3745));
  jand g3104(.dina(n3745), .dinb(n3741), .dout(n3746));
  jnot g3105(.din(n3746), .dout(n3747));
  jnot g3106(.din(n3741), .dout(n3748));
  jand g3107(.dina(n3744), .dinb(n3748), .dout(n3749));
  jand g3108(.dina(n2803), .dinb(n2127), .dout(n3750));
  jand g3109(.dina(n2808), .dinb(n2131), .dout(n3751));
  jor  g3110(.dina(n3751), .dinb(n3750), .dout(n3752));
  jand g3111(.dina(n1721), .dinb(n1059), .dout(n3753));
  jand g3112(.dina(n1562), .dinb(n1063), .dout(n3754));
  jor  g3113(.dina(n3754), .dinb(n3753), .dout(n3755));
  jnot g3114(.din(n3755), .dout(n3756));
  jand g3115(.dina(n3756), .dinb(n3752), .dout(n3757));
  jnot g3116(.din(n3757), .dout(n3758));
  jor  g3117(.dina(n2808), .dinb(\in2[1] ), .dout(n3759));
  jor  g3118(.dina(n2803), .dinb(\in3[1] ), .dout(n3760));
  jand g3119(.dina(n3760), .dinb(n3759), .dout(n3761));
  jand g3120(.dina(n1721), .dinb(n1044), .dout(n3762));
  jand g3121(.dina(n1562), .dinb(n1586), .dout(n3763));
  jor  g3122(.dina(n3763), .dinb(n3762), .dout(n3764));
  jor  g3123(.dina(n3764), .dinb(n3761), .dout(n3765));
  jand g3124(.dina(n1721), .dinb(n1046), .dout(n3766));
  jand g3125(.dina(n1562), .dinb(n1588), .dout(n3767));
  jor  g3126(.dina(n3767), .dinb(n3766), .dout(n3768));
  jor  g3127(.dina(n2808), .dinb(\in2[0] ), .dout(n3769));
  jor  g3128(.dina(n2803), .dinb(\in3[0] ), .dout(n3770));
  jand g3129(.dina(n3770), .dinb(n3769), .dout(n3771));
  jor  g3130(.dina(n3771), .dinb(n3768), .dout(n3772));
  jand g3131(.dina(n3772), .dinb(n3765), .dout(n3773));
  jand g3132(.dina(n1721), .dinb(n1049), .dout(n3774));
  jand g3133(.dina(n1562), .dinb(n1041), .dout(n3775));
  jor  g3134(.dina(n3775), .dinb(n3774), .dout(n3776));
  jor  g3135(.dina(n2808), .dinb(\in2[2] ), .dout(n3777));
  jor  g3136(.dina(n2803), .dinb(\in3[2] ), .dout(n3778));
  jand g3137(.dina(n3778), .dinb(n3777), .dout(n3779));
  jand g3138(.dina(n3779), .dinb(n3776), .dout(n3780));
  jand g3139(.dina(n3764), .dinb(n3761), .dout(n3781));
  jor  g3140(.dina(n3781), .dinb(n3780), .dout(n3782));
  jor  g3141(.dina(n3782), .dinb(n3773), .dout(n3783));
  jor  g3142(.dina(n3779), .dinb(n3776), .dout(n3784));
  jand g3143(.dina(n1721), .dinb(n1039), .dout(n3785));
  jand g3144(.dina(n1562), .dinb(n1054), .dout(n3786));
  jor  g3145(.dina(n3786), .dinb(n3785), .dout(n3787));
  jand g3146(.dina(n2803), .dinb(n2106), .dout(n3788));
  jand g3147(.dina(n2808), .dinb(n2120), .dout(n3789));
  jor  g3148(.dina(n3789), .dinb(n3788), .dout(n3790));
  jnot g3149(.din(n3790), .dout(n3791));
  jor  g3150(.dina(n3791), .dinb(n3787), .dout(n3792));
  jand g3151(.dina(n3792), .dinb(n3784), .dout(n3793));
  jand g3152(.dina(n3793), .dinb(n3783), .dout(n3794));
  jnot g3153(.din(n3752), .dout(n3795));
  jand g3154(.dina(n3755), .dinb(n3795), .dout(n3796));
  jand g3155(.dina(n3791), .dinb(n3787), .dout(n3797));
  jor  g3156(.dina(n3797), .dinb(n3796), .dout(n3798));
  jor  g3157(.dina(n3798), .dinb(n3794), .dout(n3799));
  jand g3158(.dina(n3799), .dinb(n3758), .dout(n3800));
  jor  g3159(.dina(n3800), .dinb(n3749), .dout(n3801));
  jand g3160(.dina(n3801), .dinb(n3747), .dout(n3802));
  jor  g3161(.dina(n3802), .dinb(n3738), .dout(n3803));
  jnot g3162(.din(n3725), .dout(n3804));
  jand g3163(.dina(n3728), .dinb(n3804), .dout(n3805));
  jnot g3164(.din(n3737), .dout(n3806));
  jand g3165(.dina(n3806), .dinb(n3733), .dout(n3807));
  jor  g3166(.dina(n3807), .dinb(n3805), .dout(n3808));
  jnot g3167(.din(n3808), .dout(n3809));
  jand g3168(.dina(n3809), .dinb(n3803), .dout(n3810));
  jnot g3169(.din(n3716), .dout(n3811));
  jand g3170(.dina(n3719), .dinb(n3811), .dout(n3812));
  jor  g3171(.dina(n3812), .dinb(n3810), .dout(n3813));
  jor  g3172(.dina(n3813), .dinb(n3730), .dout(n3814));
  jand g3173(.dina(n2803), .dinb(n2164), .dout(n3815));
  jand g3174(.dina(n2808), .dinb(n2157), .dout(n3816));
  jor  g3175(.dina(n3816), .dinb(n3815), .dout(n3817));
  jand g3176(.dina(n1721), .dinb(n1096), .dout(n3818));
  jand g3177(.dina(n1562), .dinb(n1089), .dout(n3819));
  jor  g3178(.dina(n3819), .dinb(n3818), .dout(n3820));
  jnot g3179(.din(n3820), .dout(n3821));
  jand g3180(.dina(n3821), .dinb(n3817), .dout(n3822));
  jnot g3181(.din(n3822), .dout(n3823));
  jand g3182(.dina(n3823), .dinb(n3814), .dout(n3824));
  jand g3183(.dina(n3824), .dinb(n3722), .dout(n3825));
  jnot g3184(.din(n3817), .dout(n3826));
  jand g3185(.dina(n3820), .dinb(n3826), .dout(n3827));
  jor  g3186(.dina(n3827), .dinb(n3825), .dout(n3828));
  jor  g3187(.dina(n3828), .dinb(n3713), .dout(n3829));
  jnot g3188(.din(n3708), .dout(n3830));
  jand g3189(.dina(n3711), .dinb(n3830), .dout(n3831));
  jand g3190(.dina(n1721), .dinb(n1032), .dout(n3832));
  jand g3191(.dina(n1562), .dinb(n1029), .dout(n3833));
  jor  g3192(.dina(n3833), .dinb(n3832), .dout(n3834));
  jnot g3193(.din(n3834), .dout(n3835));
  jand g3194(.dina(n2803), .dinb(n2099), .dout(n3836));
  jand g3195(.dina(n2808), .dinb(n2096), .dout(n3837));
  jor  g3196(.dina(n3837), .dinb(n3836), .dout(n3838));
  jand g3197(.dina(n3838), .dinb(n3835), .dout(n3839));
  jor  g3198(.dina(n3839), .dinb(n3831), .dout(n3840));
  jnot g3199(.din(n3840), .dout(n3841));
  jand g3200(.dina(n3841), .dinb(n3829), .dout(n3842));
  jnot g3201(.din(n3703), .dout(n3843));
  jand g3202(.dina(n3843), .dinb(n3699), .dout(n3844));
  jnot g3203(.din(n3838), .dout(n3845));
  jand g3204(.dina(n3845), .dinb(n3834), .dout(n3846));
  jor  g3205(.dina(n3846), .dinb(n3844), .dout(n3847));
  jor  g3206(.dina(n3847), .dinb(n3842), .dout(n3848));
  jand g3207(.dina(n3848), .dinb(n3705), .dout(n3849));
  jor  g3208(.dina(n3849), .dinb(n3696), .dout(n3850));
  jand g3209(.dina(n3850), .dinb(n3694), .dout(n3851));
  jor  g3210(.dina(n3851), .dinb(n3685), .dout(n3852));
  jnot g3211(.din(n3672), .dout(n3853));
  jand g3212(.dina(n3675), .dinb(n3853), .dout(n3854));
  jnot g3213(.din(n3680), .dout(n3855));
  jand g3214(.dina(n3683), .dinb(n3855), .dout(n3856));
  jor  g3215(.dina(n3856), .dinb(n3854), .dout(n3857));
  jnot g3216(.din(n3857), .dout(n3858));
  jand g3217(.dina(n3858), .dinb(n3852), .dout(n3859));
  jnot g3218(.din(n3663), .dout(n3860));
  jand g3219(.dina(n3666), .dinb(n3860), .dout(n3861));
  jor  g3220(.dina(n3861), .dinb(n3859), .dout(n3862));
  jor  g3221(.dina(n3862), .dinb(n3677), .dout(n3863));
  jand g3222(.dina(n2803), .dinb(n2196), .dout(n3864));
  jand g3223(.dina(n2808), .dinb(n2189), .dout(n3865));
  jor  g3224(.dina(n3865), .dinb(n3864), .dout(n3866));
  jand g3225(.dina(n1721), .dinb(n1128), .dout(n3867));
  jand g3226(.dina(n1562), .dinb(n1121), .dout(n3868));
  jor  g3227(.dina(n3868), .dinb(n3867), .dout(n3869));
  jnot g3228(.din(n3869), .dout(n3870));
  jand g3229(.dina(n3870), .dinb(n3866), .dout(n3871));
  jnot g3230(.din(n3871), .dout(n3872));
  jand g3231(.dina(n3872), .dinb(n3863), .dout(n3873));
  jand g3232(.dina(n3873), .dinb(n3669), .dout(n3874));
  jnot g3233(.din(n3866), .dout(n3875));
  jand g3234(.dina(n3869), .dinb(n3875), .dout(n3876));
  jor  g3235(.dina(n3876), .dinb(n3874), .dout(n3877));
  jor  g3236(.dina(n3877), .dinb(n3660), .dout(n3878));
  jnot g3237(.din(n3655), .dout(n3879));
  jand g3238(.dina(n3658), .dinb(n3879), .dout(n3880));
  jnot g3239(.din(n3647), .dout(n3881));
  jand g3240(.dina(n3650), .dinb(n3881), .dout(n3882));
  jor  g3241(.dina(n3882), .dinb(n3880), .dout(n3883));
  jnot g3242(.din(n3883), .dout(n3884));
  jand g3243(.dina(n3884), .dinb(n3878), .dout(n3885));
  jor  g3244(.dina(n3885), .dinb(n3652), .dout(n3886));
  jand g3245(.dina(n3886), .dinb(n3644), .dout(n3887));
  jand g3246(.dina(n1721), .dinb(n1000), .dout(n3888));
  jand g3247(.dina(n1562), .dinb(n997), .dout(n3889));
  jor  g3248(.dina(n3889), .dinb(n3888), .dout(n3890));
  jand g3249(.dina(n2803), .dinb(n2067), .dout(n3891));
  jand g3250(.dina(n2808), .dinb(n2064), .dout(n3892));
  jor  g3251(.dina(n3892), .dinb(n3891), .dout(n3893));
  jnot g3252(.din(n3893), .dout(n3894));
  jand g3253(.dina(n3894), .dinb(n3890), .dout(n3895));
  jor  g3254(.dina(n3895), .dinb(n3887), .dout(n3896));
  jor  g3255(.dina(n3896), .dinb(n3641), .dout(n3897));
  jnot g3256(.din(n3890), .dout(n3898));
  jand g3257(.dina(n3893), .dinb(n3898), .dout(n3899));
  jnot g3258(.din(n3628), .dout(n3900));
  jand g3259(.dina(n3631), .dinb(n3900), .dout(n3901));
  jor  g3260(.dina(n3901), .dinb(n3899), .dout(n3902));
  jnot g3261(.din(n3902), .dout(n3903));
  jand g3262(.dina(n3903), .dinb(n3897), .dout(n3904));
  jor  g3263(.dina(n3904), .dinb(n3633), .dout(n3905));
  jand g3264(.dina(n3905), .dinb(n3625), .dout(n3906));
  jnot g3265(.din(n3623), .dout(n3907));
  jand g3266(.dina(n3907), .dinb(n3619), .dout(n3908));
  jnot g3267(.din(n3601), .dout(n3909));
  jand g3268(.dina(n3604), .dinb(n3909), .dout(n3910));
  jor  g3269(.dina(n3910), .dinb(n3908), .dout(n3911));
  jor  g3270(.dina(n3911), .dinb(n3906), .dout(n3912));
  jand g3271(.dina(n3912), .dinb(n3616), .dout(n3913));
  jnot g3272(.din(n3609), .dout(n3914));
  jand g3273(.dina(n3612), .dinb(n3914), .dout(n3915));
  jor  g3274(.dina(n3915), .dinb(n3913), .dout(n3916));
  jor  g3275(.dina(n3916), .dinb(n3598), .dout(n3917));
  jnot g3276(.din(n3593), .dout(n3918));
  jand g3277(.dina(n3596), .dinb(n3918), .dout(n3919));
  jand g3278(.dina(n1721), .dinb(n988), .dout(n3920));
  jand g3279(.dina(n1562), .dinb(n985), .dout(n3921));
  jor  g3280(.dina(n3921), .dinb(n3920), .dout(n3922));
  jnot g3281(.din(n3922), .dout(n3923));
  jand g3282(.dina(n2803), .dinb(n2055), .dout(n3924));
  jand g3283(.dina(n2808), .dinb(n2052), .dout(n3925));
  jor  g3284(.dina(n3925), .dinb(n3924), .dout(n3926));
  jand g3285(.dina(n3926), .dinb(n3923), .dout(n3927));
  jor  g3286(.dina(n3927), .dinb(n3919), .dout(n3928));
  jnot g3287(.din(n3928), .dout(n3929));
  jand g3288(.dina(n3929), .dinb(n3917), .dout(n3930));
  jnot g3289(.din(n3588), .dout(n3931));
  jand g3290(.dina(n3931), .dinb(n3584), .dout(n3932));
  jnot g3291(.din(n3926), .dout(n3933));
  jand g3292(.dina(n3933), .dinb(n3922), .dout(n3934));
  jor  g3293(.dina(n3934), .dinb(n3932), .dout(n3935));
  jor  g3294(.dina(n3935), .dinb(n3930), .dout(n3936));
  jand g3295(.dina(n3936), .dinb(n3590), .dout(n3937));
  jor  g3296(.dina(n3937), .dinb(n3581), .dout(n3938));
  jand g3297(.dina(n1721), .dinb(n973), .dout(n3939));
  jand g3298(.dina(n1562), .dinb(n1174), .dout(n3940));
  jor  g3299(.dina(n3940), .dinb(n3939), .dout(n3941));
  jnot g3300(.din(n3941), .dout(n3942));
  jand g3301(.dina(n2803), .dinb(n2040), .dout(n3943));
  jand g3302(.dina(n2808), .dinb(n2242), .dout(n3944));
  jor  g3303(.dina(n3944), .dinb(n3943), .dout(n3945));
  jand g3304(.dina(n3945), .dinb(n3942), .dout(n3946));
  jnot g3305(.din(n3576), .dout(n3947));
  jand g3306(.dina(n3579), .dinb(n3947), .dout(n3948));
  jor  g3307(.dina(n3948), .dinb(n3946), .dout(n3949));
  jnot g3308(.din(n3949), .dout(n3950));
  jand g3309(.dina(n3950), .dinb(n3938), .dout(n3951));
  jnot g3310(.din(n3571), .dout(n3952));
  jand g3311(.dina(n3952), .dinb(n3567), .dout(n3953));
  jnot g3312(.din(n3945), .dout(n3954));
  jand g3313(.dina(n3954), .dinb(n3941), .dout(n3955));
  jor  g3314(.dina(n3955), .dinb(n3953), .dout(n3956));
  jor  g3315(.dina(n3956), .dinb(n3951), .dout(n3957));
  jand g3316(.dina(n3957), .dinb(n3573), .dout(n3958));
  jand g3317(.dina(n3507), .dinb(n3475), .dout(n3959));
  jnot g3318(.din(n3537), .dout(n3960));
  jand g3319(.dina(n3540), .dinb(n3960), .dout(n3961));
  jor  g3320(.dina(n3961), .dinb(n3515), .dout(n3962));
  jnot g3321(.din(n3962), .dout(n3963));
  jand g3322(.dina(n3963), .dinb(n3959), .dout(n3964));
  jand g3323(.dina(n3964), .dinb(n3493), .dout(n3965));
  jnot g3324(.din(n3965), .dout(n3966));
  jor  g3325(.dina(n3966), .dinb(n3958), .dout(n3967));
  jor  g3326(.dina(n3967), .dinb(n3533), .dout(n3968));
  jand g3327(.dina(n3968), .dinb(n3564), .dout(n3969));
  jand g3328(.dina(n1721), .dinb(n931), .dout(n3970));
  jand g3329(.dina(n1562), .dinb(n929), .dout(n3971));
  jor  g3330(.dina(n3971), .dinb(n3970), .dout(n3972));
  jand g3331(.dina(n2803), .dinb(n2281), .dout(n3973));
  jand g3332(.dina(n2808), .dinb(n2295), .dout(n3974));
  jor  g3333(.dina(n3974), .dinb(n3973), .dout(n3975));
  jnot g3334(.din(n3975), .dout(n3976));
  jand g3335(.dina(n3976), .dinb(n3972), .dout(n3977));
  jand g3336(.dina(n1721), .dinb(n1210), .dout(n3978));
  jand g3337(.dina(n1562), .dinb(n934), .dout(n3979));
  jor  g3338(.dina(n3979), .dinb(n3978), .dout(n3980));
  jand g3339(.dina(n2803), .dinb(n2278), .dout(n3981));
  jand g3340(.dina(n2808), .dinb(n2300), .dout(n3982));
  jor  g3341(.dina(n3982), .dinb(n3981), .dout(n3983));
  jnot g3342(.din(n3983), .dout(n3984));
  jand g3343(.dina(n3984), .dinb(n3980), .dout(n3985));
  jand g3344(.dina(n1721), .dinb(n920), .dout(n3986));
  jand g3345(.dina(n1562), .dinb(n927), .dout(n3987));
  jor  g3346(.dina(n3987), .dinb(n3986), .dout(n3988));
  jand g3347(.dina(n2803), .dinb(n2284), .dout(n3989));
  jand g3348(.dina(n2808), .dinb(n2297), .dout(n3990));
  jor  g3349(.dina(n3990), .dinb(n3989), .dout(n3991));
  jnot g3350(.din(n3991), .dout(n3992));
  jand g3351(.dina(n3992), .dinb(n3988), .dout(n3993));
  jnot g3352(.din(n3993), .dout(n3994));
  jor  g3353(.dina(n3463), .dinb(n3421), .dout(n3995));
  jand g3354(.dina(n3995), .dinb(n3994), .dout(n3996));
  jand g3355(.dina(n3996), .dinb(n3459), .dout(n3997));
  jnot g3356(.din(n3997), .dout(n3998));
  jor  g3357(.dina(n3998), .dinb(n3985), .dout(n3999));
  jor  g3358(.dina(n3999), .dinb(n3977), .dout(n4000));
  jor  g3359(.dina(n4000), .dinb(n3969), .dout(n4001));
  jnot g3360(.din(n3988), .dout(n4002));
  jand g3361(.dina(n3991), .dinb(n4002), .dout(n4003));
  jnot g3362(.din(n3977), .dout(n4004));
  jnot g3363(.din(n3980), .dout(n4005));
  jand g3364(.dina(n3983), .dinb(n4005), .dout(n4006));
  jand g3365(.dina(n4006), .dinb(n4004), .dout(n4007));
  jnot g3366(.din(n3972), .dout(n4008));
  jand g3367(.dina(n3975), .dinb(n4008), .dout(n4009));
  jor  g3368(.dina(n4009), .dinb(n4007), .dout(n4010));
  jor  g3369(.dina(n4010), .dinb(n4003), .dout(n4011));
  jand g3370(.dina(n4011), .dinb(n3997), .dout(n4012));
  jnot g3371(.din(n3451), .dout(n4013));
  jand g3372(.dina(n3454), .dinb(n4013), .dout(n4014));
  jnot g3373(.din(n3424), .dout(n4015));
  jand g3374(.dina(n3427), .dinb(n4015), .dout(n4016));
  jor  g3375(.dina(n4016), .dinb(n4014), .dout(n4017));
  jand g3376(.dina(n4017), .dinb(n3457), .dout(n4018));
  jand g3377(.dina(n4018), .dinb(n3448), .dout(n4019));
  jnot g3378(.din(n3438), .dout(n4020));
  jnot g3379(.din(n3433), .dout(n4021));
  jand g3380(.dina(n3436), .dinb(n4021), .dout(n4022));
  jnot g3381(.din(n3445), .dout(n4023));
  jand g3382(.dina(n4023), .dinb(n3441), .dout(n4024));
  jor  g3383(.dina(n4024), .dinb(n4022), .dout(n4025));
  jand g3384(.dina(n4025), .dinb(n4020), .dout(n4026));
  jor  g3385(.dina(n4026), .dinb(n4019), .dout(n4027));
  jor  g3386(.dina(n4027), .dinb(n4012), .dout(n4028));
  jnot g3387(.din(n4028), .dout(n4029));
  jand g3388(.dina(n4029), .dinb(n4001), .dout(n4030));
  jand g3389(.dina(n4030), .dinb(n3466), .dout(n4031));
  jand g3390(.dina(n1721), .dinb(n1239), .dout(n4032));
  jand g3391(.dina(n1562), .dinb(n1253), .dout(n4033));
  jor  g3392(.dina(n4033), .dinb(n4032), .dout(n4034));
  jand g3393(.dina(n2803), .dinb(n2327), .dout(n4035));
  jand g3394(.dina(n2808), .dinb(n2341), .dout(n4036));
  jor  g3395(.dina(n4036), .dinb(n4035), .dout(n4037));
  jnot g3396(.din(n4037), .dout(n4038));
  jand g3397(.dina(n4038), .dinb(n4034), .dout(n4039));
  jand g3398(.dina(n2803), .dinb(n2330), .dout(n4040));
  jand g3399(.dina(n2808), .dinb(n2343), .dout(n4041));
  jor  g3400(.dina(n4041), .dinb(n4040), .dout(n4042));
  jnot g3401(.din(n4042), .dout(n4043));
  jand g3402(.dina(n1721), .dinb(n1242), .dout(n4044));
  jand g3403(.dina(n1562), .dinb(n1255), .dout(n4045));
  jor  g3404(.dina(n4045), .dinb(n4044), .dout(n4046));
  jand g3405(.dina(n4046), .dinb(n4043), .dout(n4047));
  jor  g3406(.dina(n4047), .dinb(n4039), .dout(n4048));
  jand g3407(.dina(n2803), .dinb(n1984), .dout(n4049));
  jand g3408(.dina(n2808), .dinb(n2355), .dout(n4050));
  jor  g3409(.dina(n4050), .dinb(n4049), .dout(n4051));
  jnot g3410(.din(n4051), .dout(n4052));
  jand g3411(.dina(n1721), .dinb(n901), .dout(n4053));
  jand g3412(.dina(n1562), .dinb(n1267), .dout(n4054));
  jor  g3413(.dina(n4054), .dinb(n4053), .dout(n4055));
  jand g3414(.dina(n4055), .dinb(n4052), .dout(n4056));
  jand g3415(.dina(n1721), .dinb(n894), .dout(n4057));
  jand g3416(.dina(n1562), .dinb(n1272), .dout(n4058));
  jor  g3417(.dina(n4058), .dinb(n4057), .dout(n4059));
  jand g3418(.dina(n2803), .dinb(n1977), .dout(n4060));
  jand g3419(.dina(n2808), .dinb(n2360), .dout(n4061));
  jor  g3420(.dina(n4061), .dinb(n4060), .dout(n4062));
  jnot g3421(.din(n4062), .dout(n4063));
  jand g3422(.dina(n4063), .dinb(n4059), .dout(n4064));
  jor  g3423(.dina(n4064), .dinb(n4056), .dout(n4065));
  jnot g3424(.din(n3416), .dout(n4066));
  jand g3425(.dina(n4066), .dinb(n3412), .dout(n4067));
  jand g3426(.dina(n2803), .dinb(n1981), .dout(n4068));
  jand g3427(.dina(n2808), .dinb(n2358), .dout(n4069));
  jor  g3428(.dina(n4069), .dinb(n4068), .dout(n4070));
  jnot g3429(.din(n4070), .dout(n4071));
  jand g3430(.dina(n1721), .dinb(n898), .dout(n4072));
  jand g3431(.dina(n1562), .dinb(n1270), .dout(n4073));
  jor  g3432(.dina(n4073), .dinb(n4072), .dout(n4074));
  jand g3433(.dina(n4074), .dinb(n4071), .dout(n4075));
  jor  g3434(.dina(n4075), .dinb(n4067), .dout(n4076));
  jand g3435(.dina(n2803), .dinb(n2324), .dout(n4077));
  jand g3436(.dina(n2808), .dinb(n2346), .dout(n4078));
  jor  g3437(.dina(n4078), .dinb(n4077), .dout(n4079));
  jnot g3438(.din(n4079), .dout(n4080));
  jand g3439(.dina(n1721), .dinb(n1236), .dout(n4081));
  jand g3440(.dina(n1562), .dinb(n1258), .dout(n4082));
  jor  g3441(.dina(n4082), .dinb(n4081), .dout(n4083));
  jand g3442(.dina(n4083), .dinb(n4080), .dout(n4084));
  jand g3443(.dina(n1721), .dinb(n1244), .dout(n4085));
  jand g3444(.dina(n1562), .dinb(n893), .dout(n4086));
  jor  g3445(.dina(n4086), .dinb(n4085), .dout(n4087));
  jand g3446(.dina(n2803), .dinb(n2332), .dout(n4088));
  jand g3447(.dina(n2808), .dinb(n1976), .dout(n4089));
  jor  g3448(.dina(n4089), .dinb(n4088), .dout(n4090));
  jnot g3449(.din(n4090), .dout(n4091));
  jand g3450(.dina(n4091), .dinb(n4087), .dout(n4092));
  jor  g3451(.dina(n4092), .dinb(n4084), .dout(n4093));
  jor  g3452(.dina(n4093), .dinb(n4076), .dout(n4094));
  jor  g3453(.dina(n4094), .dinb(n4065), .dout(n4095));
  jor  g3454(.dina(n4095), .dinb(n4048), .dout(n4096));
  jor  g3455(.dina(n4096), .dinb(n4031), .dout(n4097));
  jnot g3456(.din(n4076), .dout(n4098));
  jnot g3457(.din(n4059), .dout(n4099));
  jand g3458(.dina(n4062), .dinb(n4099), .dout(n4100));
  jnot g3459(.din(n4074), .dout(n4101));
  jand g3460(.dina(n4101), .dinb(n4070), .dout(n4102));
  jnot g3461(.din(n4065), .dout(n4103));
  jnot g3462(.din(n4055), .dout(n4104));
  jand g3463(.dina(n4104), .dinb(n4051), .dout(n4105));
  jnot g3464(.din(n4092), .dout(n4106));
  jnot g3465(.din(n4048), .dout(n4107));
  jnot g3466(.din(n4083), .dout(n4108));
  jand g3467(.dina(n4108), .dinb(n4079), .dout(n4109));
  jnot g3468(.din(n4034), .dout(n4110));
  jand g3469(.dina(n4037), .dinb(n4110), .dout(n4111));
  jor  g3470(.dina(n4111), .dinb(n4109), .dout(n4112));
  jand g3471(.dina(n4112), .dinb(n4107), .dout(n4113));
  jnot g3472(.din(n4087), .dout(n4114));
  jand g3473(.dina(n4090), .dinb(n4114), .dout(n4115));
  jnot g3474(.din(n4046), .dout(n4116));
  jand g3475(.dina(n4116), .dinb(n4042), .dout(n4117));
  jor  g3476(.dina(n4117), .dinb(n4115), .dout(n4118));
  jor  g3477(.dina(n4118), .dinb(n4113), .dout(n4119));
  jand g3478(.dina(n4119), .dinb(n4106), .dout(n4120));
  jor  g3479(.dina(n4120), .dinb(n4105), .dout(n4121));
  jand g3480(.dina(n4121), .dinb(n4103), .dout(n4122));
  jor  g3481(.dina(n4122), .dinb(n4102), .dout(n4123));
  jor  g3482(.dina(n4123), .dinb(n4100), .dout(n4124));
  jand g3483(.dina(n4124), .dinb(n4098), .dout(n4125));
  jnot g3484(.din(n4125), .dout(n4126));
  jand g3485(.dina(n4126), .dinb(n4097), .dout(n4127));
  jand g3486(.dina(n4127), .dinb(n3418), .dout(n4128));
  jnot g3487(.din(n3399), .dout(n4129));
  jand g3488(.dina(n4129), .dinb(n3395), .dout(n4130));
  jor  g3489(.dina(n4130), .dinb(n3391), .dout(n4131));
  jor  g3490(.dina(n4131), .dinb(n3380), .dout(n4132));
  jor  g3491(.dina(n4132), .dinb(n3360), .dout(n4133));
  jor  g3492(.dina(n4133), .dinb(n4128), .dout(n4134));
  jnot g3493(.din(n3359), .dout(n4135));
  jnot g3494(.din(n3352), .dout(n4136));
  jand g3495(.dina(n3355), .dinb(n4136), .dout(n4137));
  jnot g3496(.din(n3328), .dout(n4138));
  jand g3497(.dina(n3331), .dinb(n4138), .dout(n4139));
  jor  g3498(.dina(n4139), .dinb(n4137), .dout(n4140));
  jand g3499(.dina(n4140), .dinb(n4135), .dout(n4141));
  jnot g3500(.din(n3349), .dout(n4142));
  jnot g3501(.din(n3344), .dout(n4143));
  jand g3502(.dina(n3347), .dinb(n4143), .dout(n4144));
  jnot g3503(.din(n3340), .dout(n4145));
  jand g3504(.dina(n4145), .dinb(n3336), .dout(n4146));
  jor  g3505(.dina(n4146), .dinb(n4144), .dout(n4147));
  jand g3506(.dina(n4147), .dinb(n4142), .dout(n4148));
  jor  g3507(.dina(n4148), .dinb(n4141), .dout(n4149));
  jnot g3508(.din(n4149), .dout(n4150));
  jand g3509(.dina(n4150), .dinb(n4134), .dout(n4151));
  jand g3510(.dina(n4151), .dinb(n3409), .dout(n4152));
  jnot g3511(.din(n3316), .dout(n4153));
  jand g3512(.dina(n3319), .dinb(n4153), .dout(n4154));
  jor  g3513(.dina(n4154), .dinb(n3312), .dout(n4155));
  jor  g3514(.dina(n4155), .dinb(n4152), .dout(n4156));
  jand g3515(.dina(n4156), .dinb(n3325), .dout(n4157));
  jnot g3516(.din(n3292), .dout(n4158));
  jand g3517(.dina(n4158), .dinb(n3288), .dout(n4159));
  jnot g3518(.din(n3297), .dout(n4160));
  jand g3519(.dina(n3300), .dinb(n4160), .dout(n4161));
  jor  g3520(.dina(n4161), .dinb(n4159), .dout(n4162));
  jor  g3521(.dina(n4162), .dinb(n4157), .dout(n4163));
  jand g3522(.dina(n4163), .dinb(n3294), .dout(n4164));
  jnot g3523(.din(n3273), .dout(n4165));
  jand g3524(.dina(n4165), .dinb(n3269), .dout(n4166));
  jor  g3525(.dina(n4166), .dinb(n3263), .dout(n4167));
  jor  g3526(.dina(n4167), .dinb(n4164), .dout(n4168));
  jand g3527(.dina(n4168), .dinb(n3285), .dout(n4169));
  jand g3528(.dina(n2803), .dinb(n2438), .dout(n4170));
  jand g3529(.dina(n2808), .dinb(n2452), .dout(n4171));
  jor  g3530(.dina(n4171), .dinb(n4170), .dout(n4172));
  jnot g3531(.din(n4172), .dout(n4173));
  jand g3532(.dina(n1721), .dinb(n832), .dout(n4174));
  jand g3533(.dina(n1562), .dinb(n1359), .dout(n4175));
  jor  g3534(.dina(n4175), .dinb(n4174), .dout(n4176));
  jand g3535(.dina(n4176), .dinb(n4173), .dout(n4177));
  jnot g3536(.din(n4177), .dout(n4178));
  jand g3537(.dina(n1721), .dinb(n1345), .dout(n4179));
  jand g3538(.dina(n1562), .dinb(n829), .dout(n4180));
  jor  g3539(.dina(n4180), .dinb(n4179), .dout(n4181));
  jand g3540(.dina(n2803), .dinb(n2433), .dout(n4182));
  jand g3541(.dina(n2808), .dinb(n1917), .dout(n4183));
  jor  g3542(.dina(n4183), .dinb(n4182), .dout(n4184));
  jnot g3543(.din(n4184), .dout(n4185));
  jand g3544(.dina(n4185), .dinb(n4181), .dout(n4186));
  jand g3545(.dina(n2803), .dinb(n2435), .dout(n4187));
  jand g3546(.dina(n2808), .dinb(n2448), .dout(n4188));
  jor  g3547(.dina(n4188), .dinb(n4187), .dout(n4189));
  jnot g3548(.din(n4189), .dout(n4190));
  jand g3549(.dina(n1721), .dinb(n1347), .dout(n4191));
  jand g3550(.dina(n1562), .dinb(n1355), .dout(n4192));
  jor  g3551(.dina(n4192), .dinb(n4191), .dout(n4193));
  jand g3552(.dina(n4193), .dinb(n4190), .dout(n4194));
  jor  g3553(.dina(n4194), .dinb(n4186), .dout(n4195));
  jnot g3554(.din(n4195), .dout(n4196));
  jand g3555(.dina(n1721), .dinb(n834), .dout(n4197));
  jand g3556(.dina(n1562), .dinb(n1353), .dout(n4198));
  jor  g3557(.dina(n4198), .dinb(n4197), .dout(n4199));
  jand g3558(.dina(n2803), .dinb(n2440), .dout(n4200));
  jand g3559(.dina(n2808), .dinb(n2446), .dout(n4201));
  jor  g3560(.dina(n4201), .dinb(n4200), .dout(n4202));
  jnot g3561(.din(n4202), .dout(n4203));
  jand g3562(.dina(n4203), .dinb(n4199), .dout(n4204));
  jnot g3563(.din(n4204), .dout(n4205));
  jand g3564(.dina(n4205), .dinb(n4196), .dout(n4206));
  jand g3565(.dina(n4206), .dinb(n4178), .dout(n4207));
  jnot g3566(.din(n4207), .dout(n4208));
  jor  g3567(.dina(n4208), .dinb(n4169), .dout(n4209));
  jnot g3568(.din(n4181), .dout(n4210));
  jand g3569(.dina(n4184), .dinb(n4210), .dout(n4211));
  jnot g3570(.din(n4193), .dout(n4212));
  jand g3571(.dina(n4212), .dinb(n4189), .dout(n4213));
  jnot g3572(.din(n4176), .dout(n4214));
  jand g3573(.dina(n4214), .dinb(n4172), .dout(n4215));
  jand g3574(.dina(n4215), .dinb(n4205), .dout(n4216));
  jnot g3575(.din(n4199), .dout(n4217));
  jand g3576(.dina(n4202), .dinb(n4217), .dout(n4218));
  jor  g3577(.dina(n4218), .dinb(n4216), .dout(n4219));
  jor  g3578(.dina(n4219), .dinb(n4213), .dout(n4220));
  jand g3579(.dina(n4220), .dinb(n4196), .dout(n4221));
  jor  g3580(.dina(n4221), .dinb(n4211), .dout(n4222));
  jnot g3581(.din(n4222), .dout(n4223));
  jand g3582(.dina(n4223), .dinb(n4209), .dout(n4224));
  jor  g3583(.dina(n4224), .dinb(n3237), .dout(n4225));
  jnot g3584(.din(n3236), .dout(n4226));
  jnot g3585(.din(n3229), .dout(n4227));
  jand g3586(.dina(n3232), .dinb(n4227), .dout(n4228));
  jnot g3587(.din(n3205), .dout(n4229));
  jand g3588(.dina(n3208), .dinb(n4229), .dout(n4230));
  jor  g3589(.dina(n4230), .dinb(n4228), .dout(n4231));
  jand g3590(.dina(n4231), .dinb(n4226), .dout(n4232));
  jnot g3591(.din(n3226), .dout(n4233));
  jnot g3592(.din(n3221), .dout(n4234));
  jand g3593(.dina(n3224), .dinb(n4234), .dout(n4235));
  jnot g3594(.din(n3217), .dout(n4236));
  jand g3595(.dina(n4236), .dinb(n3213), .dout(n4237));
  jor  g3596(.dina(n4237), .dinb(n4235), .dout(n4238));
  jand g3597(.dina(n4238), .dinb(n4233), .dout(n4239));
  jor  g3598(.dina(n4239), .dinb(n4232), .dout(n4240));
  jnot g3599(.din(n4240), .dout(n4241));
  jand g3600(.dina(n4241), .dinb(n4225), .dout(n4242));
  jor  g3601(.dina(n4242), .dinb(n3202), .dout(n4243));
  jnot g3602(.din(n3184), .dout(n4244));
  jnot g3603(.din(n3182), .dout(n4245));
  jand g3604(.dina(n4245), .dinb(n3178), .dout(n4246));
  jnot g3605(.din(n3192), .dout(n4247));
  jnot g3606(.din(n3199), .dout(n4248));
  jand g3607(.dina(n4248), .dinb(n3195), .dout(n4249));
  jand g3608(.dina(n4249), .dinb(n4247), .dout(n4250));
  jnot g3609(.din(n3187), .dout(n4251));
  jand g3610(.dina(n3190), .dinb(n4251), .dout(n4252));
  jor  g3611(.dina(n4252), .dinb(n4250), .dout(n4253));
  jor  g3612(.dina(n4253), .dinb(n4246), .dout(n4254));
  jand g3613(.dina(n4254), .dinb(n4244), .dout(n4255));
  jnot g3614(.din(n4255), .dout(n4256));
  jand g3615(.dina(n4256), .dinb(n4243), .dout(n4257));
  jand g3616(.dina(n4257), .dinb(n3173), .dout(n4258));
  jnot g3617(.din(n3152), .dout(n4259));
  jand g3618(.dina(n4259), .dinb(n3148), .dout(n4260));
  jor  g3619(.dina(n4260), .dinb(n3142), .dout(n4261));
  jor  g3620(.dina(n4261), .dinb(n4258), .dout(n4262));
  jand g3621(.dina(n4262), .dinb(n3164), .dout(n4263));
  jand g3622(.dina(n4263), .dinb(n3156), .dout(n4264));
  jor  g3623(.dina(n4264), .dinb(n3116), .dout(n4265));
  jnot g3624(.din(n3084), .dout(n4266));
  jand g3625(.dina(n3087), .dinb(n4266), .dout(n4267));
  jnot g3626(.din(n3098), .dout(n4268));
  jnot g3627(.din(n3096), .dout(n4269));
  jand g3628(.dina(n4269), .dinb(n3092), .dout(n4270));
  jnot g3629(.din(n3106), .dout(n4271));
  jnot g3630(.din(n3113), .dout(n4272));
  jand g3631(.dina(n4272), .dinb(n3109), .dout(n4273));
  jand g3632(.dina(n4273), .dinb(n4271), .dout(n4274));
  jnot g3633(.din(n3101), .dout(n4275));
  jand g3634(.dina(n3104), .dinb(n4275), .dout(n4276));
  jor  g3635(.dina(n4276), .dinb(n4274), .dout(n4277));
  jor  g3636(.dina(n4277), .dinb(n4270), .dout(n4278));
  jand g3637(.dina(n4278), .dinb(n4268), .dout(n4279));
  jor  g3638(.dina(n4279), .dinb(n4267), .dout(n4280));
  jnot g3639(.din(n4280), .dout(n4281));
  jand g3640(.dina(n4281), .dinb(n4265), .dout(n4282));
  jor  g3641(.dina(n4282), .dinb(n3081), .dout(n4283));
  jnot g3642(.din(n3080), .dout(n4284));
  jnot g3643(.din(n3073), .dout(n4285));
  jand g3644(.dina(n3076), .dinb(n4285), .dout(n4286));
  jnot g3645(.din(n3049), .dout(n4287));
  jand g3646(.dina(n3052), .dinb(n4287), .dout(n4288));
  jor  g3647(.dina(n4288), .dinb(n4286), .dout(n4289));
  jand g3648(.dina(n4289), .dinb(n4284), .dout(n4290));
  jnot g3649(.din(n3070), .dout(n4291));
  jnot g3650(.din(n3065), .dout(n4292));
  jand g3651(.dina(n3068), .dinb(n4292), .dout(n4293));
  jnot g3652(.din(n3061), .dout(n4294));
  jand g3653(.dina(n4294), .dinb(n3057), .dout(n4295));
  jor  g3654(.dina(n4295), .dinb(n4293), .dout(n4296));
  jand g3655(.dina(n4296), .dinb(n4291), .dout(n4297));
  jor  g3656(.dina(n4297), .dinb(n4290), .dout(n4298));
  jnot g3657(.din(n4298), .dout(n4299));
  jand g3658(.dina(n4299), .dinb(n4283), .dout(n4300));
  jor  g3659(.dina(n4300), .dinb(n3046), .dout(n4301));
  jnot g3660(.din(n3014), .dout(n4302));
  jand g3661(.dina(n3017), .dinb(n4302), .dout(n4303));
  jnot g3662(.din(n3028), .dout(n4304));
  jnot g3663(.din(n3026), .dout(n4305));
  jand g3664(.dina(n4305), .dinb(n3022), .dout(n4306));
  jnot g3665(.din(n3036), .dout(n4307));
  jnot g3666(.din(n3043), .dout(n4308));
  jand g3667(.dina(n4308), .dinb(n3039), .dout(n4309));
  jand g3668(.dina(n4309), .dinb(n4307), .dout(n4310));
  jnot g3669(.din(n3031), .dout(n4311));
  jand g3670(.dina(n3034), .dinb(n4311), .dout(n4312));
  jor  g3671(.dina(n4312), .dinb(n4310), .dout(n4313));
  jor  g3672(.dina(n4313), .dinb(n4306), .dout(n4314));
  jand g3673(.dina(n4314), .dinb(n4304), .dout(n4315));
  jor  g3674(.dina(n4315), .dinb(n4303), .dout(n4316));
  jnot g3675(.din(n4316), .dout(n4317));
  jand g3676(.dina(n4317), .dinb(n4301), .dout(n4318));
  jor  g3677(.dina(n4318), .dinb(n3011), .dout(n4319));
  jnot g3678(.din(n3010), .dout(n4320));
  jnot g3679(.din(n3003), .dout(n4321));
  jand g3680(.dina(n3006), .dinb(n4321), .dout(n4322));
  jnot g3681(.din(n2979), .dout(n4323));
  jand g3682(.dina(n2982), .dinb(n4323), .dout(n4324));
  jor  g3683(.dina(n4324), .dinb(n4322), .dout(n4325));
  jand g3684(.dina(n4325), .dinb(n4320), .dout(n4326));
  jnot g3685(.din(n3000), .dout(n4327));
  jnot g3686(.din(n2995), .dout(n4328));
  jand g3687(.dina(n2998), .dinb(n4328), .dout(n4329));
  jnot g3688(.din(n2991), .dout(n4330));
  jand g3689(.dina(n4330), .dinb(n2987), .dout(n4331));
  jor  g3690(.dina(n4331), .dinb(n4329), .dout(n4332));
  jand g3691(.dina(n4332), .dinb(n4327), .dout(n4333));
  jor  g3692(.dina(n4333), .dinb(n4326), .dout(n4334));
  jnot g3693(.din(n4334), .dout(n4335));
  jand g3694(.dina(n4335), .dinb(n4319), .dout(n4336));
  jor  g3695(.dina(n4336), .dinb(n2976), .dout(n4337));
  jnot g3696(.din(n2944), .dout(n4338));
  jand g3697(.dina(n2947), .dinb(n4338), .dout(n4339));
  jnot g3698(.din(n2958), .dout(n4340));
  jnot g3699(.din(n2956), .dout(n4341));
  jand g3700(.dina(n4341), .dinb(n2952), .dout(n4342));
  jnot g3701(.din(n2966), .dout(n4343));
  jnot g3702(.din(n2973), .dout(n4344));
  jand g3703(.dina(n4344), .dinb(n2969), .dout(n4345));
  jand g3704(.dina(n4345), .dinb(n4343), .dout(n4346));
  jnot g3705(.din(n2961), .dout(n4347));
  jand g3706(.dina(n2964), .dinb(n4347), .dout(n4348));
  jor  g3707(.dina(n4348), .dinb(n4346), .dout(n4349));
  jor  g3708(.dina(n4349), .dinb(n4342), .dout(n4350));
  jand g3709(.dina(n4350), .dinb(n4340), .dout(n4351));
  jor  g3710(.dina(n4351), .dinb(n4339), .dout(n4352));
  jnot g3711(.din(n4352), .dout(n4353));
  jand g3712(.dina(n4353), .dinb(n4337), .dout(n4354));
  jor  g3713(.dina(n4354), .dinb(n2941), .dout(n4355));
  jnot g3714(.din(n2914), .dout(n4356));
  jnot g3715(.din(n2909), .dout(n4357));
  jand g3716(.dina(n2912), .dinb(n4357), .dout(n4358));
  jnot g3717(.din(n2905), .dout(n4359));
  jand g3718(.dina(n4359), .dinb(n2901), .dout(n4360));
  jor  g3719(.dina(n4360), .dinb(n4358), .dout(n4361));
  jand g3720(.dina(n4361), .dinb(n4356), .dout(n4362));
  jnot g3721(.din(n4362), .dout(n4363));
  jand g3722(.dina(n4363), .dinb(n4355), .dout(n4364));
  jand g3723(.dina(n4364), .dinb(n2938), .dout(n4365));
  jand g3724(.dina(n1721), .dinb(n677), .dout(n4366));
  jand g3725(.dina(n1562), .dinb(n1493), .dout(n4367));
  jor  g3726(.dina(n4367), .dinb(n4366), .dout(n4368));
  jand g3727(.dina(n2803), .dinb(n1770), .dout(n4369));
  jand g3728(.dina(n2808), .dinb(n2591), .dout(n4370));
  jor  g3729(.dina(n4370), .dinb(n4369), .dout(n4371));
  jnot g3730(.din(n4371), .dout(n4372));
  jand g3731(.dina(n4372), .dinb(n4368), .dout(n4373));
  jnot g3732(.din(n2896), .dout(n4374));
  jand g3733(.dina(n4374), .dinb(n2892), .dout(n4375));
  jand g3734(.dina(n2803), .dinb(n2585), .dout(n4376));
  jand g3735(.dina(n2808), .dinb(n2593), .dout(n4377));
  jor  g3736(.dina(n4377), .dinb(n4376), .dout(n4378));
  jnot g3737(.din(n4378), .dout(n4379));
  jand g3738(.dina(n1721), .dinb(n1487), .dout(n4380));
  jand g3739(.dina(n1562), .dinb(n1495), .dout(n4381));
  jor  g3740(.dina(n4381), .dinb(n4380), .dout(n4382));
  jand g3741(.dina(n4382), .dinb(n4379), .dout(n4383));
  jor  g3742(.dina(n4383), .dinb(n4375), .dout(n4384));
  jand g3743(.dina(n2803), .dinb(n1772), .dout(n4385));
  jand g3744(.dina(n2808), .dinb(n2597), .dout(n4386));
  jor  g3745(.dina(n4386), .dinb(n4385), .dout(n4387));
  jnot g3746(.din(n4387), .dout(n4388));
  jand g3747(.dina(n1721), .dinb(n679), .dout(n4389));
  jand g3748(.dina(n1562), .dinb(n1499), .dout(n4390));
  jor  g3749(.dina(n4390), .dinb(n4389), .dout(n4391));
  jand g3750(.dina(n4391), .dinb(n4388), .dout(n4392));
  jor  g3751(.dina(n4392), .dinb(n4384), .dout(n4393));
  jor  g3752(.dina(n4393), .dinb(n4373), .dout(n4394));
  jor  g3753(.dina(n4394), .dinb(n4365), .dout(n4395));
  jnot g3754(.din(n4384), .dout(n4396));
  jnot g3755(.din(n4382), .dout(n4397));
  jand g3756(.dina(n4397), .dinb(n4378), .dout(n4398));
  jnot g3757(.din(n4373), .dout(n4399));
  jnot g3758(.din(n4391), .dout(n4400));
  jand g3759(.dina(n4400), .dinb(n4387), .dout(n4401));
  jand g3760(.dina(n4401), .dinb(n4399), .dout(n4402));
  jnot g3761(.din(n4368), .dout(n4403));
  jand g3762(.dina(n4371), .dinb(n4403), .dout(n4404));
  jor  g3763(.dina(n4404), .dinb(n4402), .dout(n4405));
  jor  g3764(.dina(n4405), .dinb(n4398), .dout(n4406));
  jand g3765(.dina(n4406), .dinb(n4396), .dout(n4407));
  jnot g3766(.din(n4407), .dout(n4408));
  jand g3767(.dina(n4408), .dinb(n4395), .dout(n4409));
  jand g3768(.dina(n4409), .dinb(n2898), .dout(n4410));
  jnot g3769(.din(n2877), .dout(n4411));
  jand g3770(.dina(n4411), .dinb(n2873), .dout(n4412));
  jor  g3771(.dina(n4412), .dinb(n2867), .dout(n4413));
  jor  g3772(.dina(n4413), .dinb(n4410), .dout(n4414));
  jand g3773(.dina(n4414), .dinb(n2889), .dout(n4415));
  jand g3774(.dina(n2803), .dinb(n2615), .dout(n4416));
  jand g3775(.dina(n2808), .dinb(n2629), .dout(n4417));
  jor  g3776(.dina(n4417), .dinb(n4416), .dout(n4418));
  jnot g3777(.din(n4418), .dout(n4419));
  jand g3778(.dina(n1721), .dinb(n645), .dout(n4420));
  jand g3779(.dina(n1562), .dinb(n1526), .dout(n4421));
  jor  g3780(.dina(n4421), .dinb(n4420), .dout(n4422));
  jand g3781(.dina(n4422), .dinb(n4419), .dout(n4423));
  jnot g3782(.din(n4423), .dout(n4424));
  jand g3783(.dina(n1721), .dinb(n1512), .dout(n4425));
  jand g3784(.dina(n1562), .dinb(n642), .dout(n4426));
  jor  g3785(.dina(n4426), .dinb(n4425), .dout(n4427));
  jand g3786(.dina(n2803), .dinb(n2610), .dout(n4428));
  jand g3787(.dina(n2808), .dinb(n1740), .dout(n4429));
  jor  g3788(.dina(n4429), .dinb(n4428), .dout(n4430));
  jnot g3789(.din(n4430), .dout(n4431));
  jand g3790(.dina(n4431), .dinb(n4427), .dout(n4432));
  jand g3791(.dina(n2803), .dinb(n2612), .dout(n4433));
  jand g3792(.dina(n2808), .dinb(n2625), .dout(n4434));
  jor  g3793(.dina(n4434), .dinb(n4433), .dout(n4435));
  jnot g3794(.din(n4435), .dout(n4436));
  jand g3795(.dina(n1721), .dinb(n1514), .dout(n4437));
  jand g3796(.dina(n1562), .dinb(n1522), .dout(n4438));
  jor  g3797(.dina(n4438), .dinb(n4437), .dout(n4439));
  jand g3798(.dina(n4439), .dinb(n4436), .dout(n4440));
  jor  g3799(.dina(n4440), .dinb(n4432), .dout(n4441));
  jnot g3800(.din(n4441), .dout(n4442));
  jand g3801(.dina(n1721), .dinb(n647), .dout(n4443));
  jand g3802(.dina(n1562), .dinb(n1520), .dout(n4444));
  jor  g3803(.dina(n4444), .dinb(n4443), .dout(n4445));
  jand g3804(.dina(n2803), .dinb(n2617), .dout(n4446));
  jand g3805(.dina(n2808), .dinb(n2623), .dout(n4447));
  jor  g3806(.dina(n4447), .dinb(n4446), .dout(n4448));
  jnot g3807(.din(n4448), .dout(n4449));
  jand g3808(.dina(n4449), .dinb(n4445), .dout(n4450));
  jnot g3809(.din(n4450), .dout(n4451));
  jand g3810(.dina(n4451), .dinb(n4442), .dout(n4452));
  jand g3811(.dina(n4452), .dinb(n4424), .dout(n4453));
  jnot g3812(.din(n4453), .dout(n4454));
  jor  g3813(.dina(n4454), .dinb(n4415), .dout(n4455));
  jnot g3814(.din(n4427), .dout(n4456));
  jand g3815(.dina(n4430), .dinb(n4456), .dout(n4457));
  jnot g3816(.din(n4439), .dout(n4458));
  jand g3817(.dina(n4458), .dinb(n4435), .dout(n4459));
  jnot g3818(.din(n4422), .dout(n4460));
  jand g3819(.dina(n4460), .dinb(n4418), .dout(n4461));
  jand g3820(.dina(n4461), .dinb(n4451), .dout(n4462));
  jnot g3821(.din(n4445), .dout(n4463));
  jand g3822(.dina(n4448), .dinb(n4463), .dout(n4464));
  jor  g3823(.dina(n4464), .dinb(n4462), .dout(n4465));
  jor  g3824(.dina(n4465), .dinb(n4459), .dout(n4466));
  jand g3825(.dina(n4466), .dinb(n4442), .dout(n4467));
  jor  g3826(.dina(n4467), .dinb(n4457), .dout(n4468));
  jnot g3827(.din(n4468), .dout(n4469));
  jand g3828(.dina(n4469), .dinb(n4455), .dout(n4470));
  jor  g3829(.dina(n4470), .dinb(n2841), .dout(n4471));
  jand g3830(.dina(n4471), .dinb(n2838), .dout(n4472));
  jor  g3831(.dina(n4472), .dinb(n2644), .dout(n4473));
  jand g3832(.dina(n4473), .dinb(n2642), .dout(n4474));
  jand g3833(.dina(n4473), .dinb(n2643), .dout(n4475));
  jor  g3834(.dina(n4475), .dinb(n4474), .dout(\address[1] ));
  jor  g3835(.dina(\address[1] ), .dinb(n1723), .dout(n4477));
  jnot g3836(.din(n2644), .dout(n4478));
  jnot g3837(.din(n2841), .dout(n4479));
  jnot g3838(.din(n2941), .dout(n4480));
  jnot g3839(.din(n2976), .dout(n4481));
  jnot g3840(.din(n3011), .dout(n4482));
  jnot g3841(.din(n3046), .dout(n4483));
  jnot g3842(.din(n3081), .dout(n4484));
  jnot g3843(.din(n3116), .dout(n4485));
  jnot g3844(.din(n3202), .dout(n4486));
  jnot g3845(.din(n3237), .dout(n4487));
  jnot g3846(.din(n3581), .dout(n4488));
  jnot g3847(.din(n3598), .dout(n4489));
  jnot g3848(.din(n3633), .dout(n4490));
  jnot g3849(.din(n3641), .dout(n4491));
  jnot g3850(.din(n3652), .dout(n4492));
  jnot g3851(.din(n3660), .dout(n4493));
  jnot g3852(.din(n3677), .dout(n4494));
  jnot g3853(.din(n3685), .dout(n4495));
  jnot g3854(.din(n3696), .dout(n4496));
  jnot g3855(.din(n3713), .dout(n4497));
  jnot g3856(.din(n3730), .dout(n4498));
  jnot g3857(.din(n3738), .dout(n4499));
  jnot g3858(.din(n3749), .dout(n4500));
  jand g3859(.dina(n2803), .dinb(n2113), .dout(n4501));
  jand g3860(.dina(n2808), .dinb(n2110), .dout(n4502));
  jor  g3861(.dina(n4502), .dinb(n4501), .dout(n4503));
  jor  g3862(.dina(n1562), .dinb(\in0[1] ), .dout(n4504));
  jor  g3863(.dina(n1721), .dinb(\in1[1] ), .dout(n4505));
  jand g3864(.dina(n4505), .dinb(n4504), .dout(n4506));
  jand g3865(.dina(n4506), .dinb(n4503), .dout(n4507));
  jand g3866(.dina(n2803), .dinb(n2115), .dout(n4508));
  jand g3867(.dina(n2808), .dinb(n2672), .dout(n4509));
  jor  g3868(.dina(n4509), .dinb(n4508), .dout(n4510));
  jand g3869(.dina(n4510), .dinb(n1723), .dout(n4511));
  jor  g3870(.dina(n4511), .dinb(n4507), .dout(n4512));
  jor  g3871(.dina(n1562), .dinb(\in0[2] ), .dout(n4513));
  jor  g3872(.dina(n1721), .dinb(\in1[2] ), .dout(n4514));
  jand g3873(.dina(n4514), .dinb(n4513), .dout(n4515));
  jand g3874(.dina(n2803), .dinb(n2108), .dout(n4516));
  jand g3875(.dina(n2808), .dinb(n2122), .dout(n4517));
  jor  g3876(.dina(n4517), .dinb(n4516), .dout(n4518));
  jor  g3877(.dina(n4518), .dinb(n4515), .dout(n4519));
  jor  g3878(.dina(n4506), .dinb(n4503), .dout(n4520));
  jand g3879(.dina(n4520), .dinb(n4519), .dout(n4521));
  jand g3880(.dina(n4521), .dinb(n4512), .dout(n4522));
  jand g3881(.dina(n4518), .dinb(n4515), .dout(n4523));
  jor  g3882(.dina(n1562), .dinb(\in0[3] ), .dout(n4524));
  jor  g3883(.dina(n1721), .dinb(\in1[3] ), .dout(n4525));
  jand g3884(.dina(n4525), .dinb(n4524), .dout(n4526));
  jand g3885(.dina(n3790), .dinb(n4526), .dout(n4527));
  jor  g3886(.dina(n4527), .dinb(n4523), .dout(n4528));
  jor  g3887(.dina(n4528), .dinb(n4522), .dout(n4529));
  jnot g3888(.din(n3798), .dout(n4530));
  jand g3889(.dina(n4530), .dinb(n4529), .dout(n4531));
  jor  g3890(.dina(n4531), .dinb(n3757), .dout(n4532));
  jand g3891(.dina(n4532), .dinb(n4500), .dout(n4533));
  jor  g3892(.dina(n4533), .dinb(n3746), .dout(n4534));
  jand g3893(.dina(n4534), .dinb(n4499), .dout(n4535));
  jor  g3894(.dina(n3808), .dinb(n4535), .dout(n4536));
  jnot g3895(.din(n3812), .dout(n4537));
  jand g3896(.dina(n4537), .dinb(n4536), .dout(n4538));
  jand g3897(.dina(n4538), .dinb(n4498), .dout(n4539));
  jor  g3898(.dina(n3822), .dinb(n4539), .dout(n4540));
  jor  g3899(.dina(n4540), .dinb(n3721), .dout(n4541));
  jnot g3900(.din(n3827), .dout(n4542));
  jand g3901(.dina(n4542), .dinb(n4541), .dout(n4543));
  jand g3902(.dina(n4543), .dinb(n4497), .dout(n4544));
  jor  g3903(.dina(n3840), .dinb(n4544), .dout(n4545));
  jnot g3904(.din(n3847), .dout(n4546));
  jand g3905(.dina(n4546), .dinb(n4545), .dout(n4547));
  jor  g3906(.dina(n4547), .dinb(n3704), .dout(n4548));
  jand g3907(.dina(n4548), .dinb(n4496), .dout(n4549));
  jor  g3908(.dina(n4549), .dinb(n3693), .dout(n4550));
  jand g3909(.dina(n4550), .dinb(n4495), .dout(n4551));
  jor  g3910(.dina(n3857), .dinb(n4551), .dout(n4552));
  jnot g3911(.din(n3861), .dout(n4553));
  jand g3912(.dina(n4553), .dinb(n4552), .dout(n4554));
  jand g3913(.dina(n4554), .dinb(n4494), .dout(n4555));
  jor  g3914(.dina(n3871), .dinb(n4555), .dout(n4556));
  jor  g3915(.dina(n4556), .dinb(n3668), .dout(n4557));
  jnot g3916(.din(n3876), .dout(n4558));
  jand g3917(.dina(n4558), .dinb(n4557), .dout(n4559));
  jand g3918(.dina(n4559), .dinb(n4493), .dout(n4560));
  jor  g3919(.dina(n3883), .dinb(n4560), .dout(n4561));
  jand g3920(.dina(n4561), .dinb(n4492), .dout(n4562));
  jor  g3921(.dina(n4562), .dinb(n3643), .dout(n4563));
  jnot g3922(.din(n3895), .dout(n4564));
  jand g3923(.dina(n4564), .dinb(n4563), .dout(n4565));
  jand g3924(.dina(n4565), .dinb(n4491), .dout(n4566));
  jor  g3925(.dina(n3902), .dinb(n4566), .dout(n4567));
  jand g3926(.dina(n4567), .dinb(n4490), .dout(n4568));
  jor  g3927(.dina(n4568), .dinb(n3624), .dout(n4569));
  jnot g3928(.din(n3911), .dout(n4570));
  jand g3929(.dina(n4570), .dinb(n4569), .dout(n4571));
  jor  g3930(.dina(n4571), .dinb(n3615), .dout(n4572));
  jnot g3931(.din(n3915), .dout(n4573));
  jand g3932(.dina(n4573), .dinb(n4572), .dout(n4574));
  jand g3933(.dina(n4574), .dinb(n4489), .dout(n4575));
  jor  g3934(.dina(n3928), .dinb(n4575), .dout(n4576));
  jnot g3935(.din(n3935), .dout(n4577));
  jand g3936(.dina(n4577), .dinb(n4576), .dout(n4578));
  jor  g3937(.dina(n4578), .dinb(n3589), .dout(n4579));
  jand g3938(.dina(n4579), .dinb(n4488), .dout(n4580));
  jor  g3939(.dina(n3949), .dinb(n4580), .dout(n4581));
  jnot g3940(.din(n3956), .dout(n4582));
  jand g3941(.dina(n4582), .dinb(n4581), .dout(n4583));
  jor  g3942(.dina(n4583), .dinb(n3572), .dout(n4584));
  jand g3943(.dina(n3965), .dinb(n4584), .dout(n4585));
  jand g3944(.dina(n4585), .dinb(n3534), .dout(n4586));
  jor  g3945(.dina(n4586), .dinb(n3563), .dout(n4587));
  jnot g3946(.din(n4000), .dout(n4588));
  jand g3947(.dina(n4588), .dinb(n4587), .dout(n4589));
  jor  g3948(.dina(n4028), .dinb(n4589), .dout(n4590));
  jor  g3949(.dina(n4590), .dinb(n3465), .dout(n4591));
  jnot g3950(.din(n4096), .dout(n4592));
  jand g3951(.dina(n4592), .dinb(n4591), .dout(n4593));
  jor  g3952(.dina(n4125), .dinb(n4593), .dout(n4594));
  jor  g3953(.dina(n4594), .dinb(n3417), .dout(n4595));
  jnot g3954(.din(n4133), .dout(n4596));
  jand g3955(.dina(n4596), .dinb(n4595), .dout(n4597));
  jor  g3956(.dina(n4149), .dinb(n4597), .dout(n4598));
  jor  g3957(.dina(n4598), .dinb(n3408), .dout(n4599));
  jnot g3958(.din(n4155), .dout(n4600));
  jand g3959(.dina(n4600), .dinb(n4599), .dout(n4601));
  jor  g3960(.dina(n4601), .dinb(n3324), .dout(n4602));
  jnot g3961(.din(n4162), .dout(n4603));
  jand g3962(.dina(n4603), .dinb(n4602), .dout(n4604));
  jor  g3963(.dina(n4604), .dinb(n3293), .dout(n4605));
  jnot g3964(.din(n4167), .dout(n4606));
  jand g3965(.dina(n4606), .dinb(n4605), .dout(n4607));
  jor  g3966(.dina(n4607), .dinb(n3284), .dout(n4608));
  jand g3967(.dina(n4207), .dinb(n4608), .dout(n4609));
  jor  g3968(.dina(n4222), .dinb(n4609), .dout(n4610));
  jand g3969(.dina(n4610), .dinb(n4487), .dout(n4611));
  jor  g3970(.dina(n4240), .dinb(n4611), .dout(n4612));
  jand g3971(.dina(n4612), .dinb(n4486), .dout(n4613));
  jor  g3972(.dina(n4255), .dinb(n4613), .dout(n4614));
  jor  g3973(.dina(n4614), .dinb(n3172), .dout(n4615));
  jnot g3974(.din(n4261), .dout(n4616));
  jand g3975(.dina(n4616), .dinb(n4615), .dout(n4617));
  jor  g3976(.dina(n4617), .dinb(n3163), .dout(n4618));
  jor  g3977(.dina(n4618), .dinb(n3155), .dout(n4619));
  jand g3978(.dina(n4619), .dinb(n4485), .dout(n4620));
  jor  g3979(.dina(n4280), .dinb(n4620), .dout(n4621));
  jand g3980(.dina(n4621), .dinb(n4484), .dout(n4622));
  jor  g3981(.dina(n4298), .dinb(n4622), .dout(n4623));
  jand g3982(.dina(n4623), .dinb(n4483), .dout(n4624));
  jor  g3983(.dina(n4316), .dinb(n4624), .dout(n4625));
  jand g3984(.dina(n4625), .dinb(n4482), .dout(n4626));
  jor  g3985(.dina(n4334), .dinb(n4626), .dout(n4627));
  jand g3986(.dina(n4627), .dinb(n4481), .dout(n4628));
  jor  g3987(.dina(n4352), .dinb(n4628), .dout(n4629));
  jand g3988(.dina(n4629), .dinb(n4480), .dout(n4630));
  jor  g3989(.dina(n4362), .dinb(n4630), .dout(n4631));
  jor  g3990(.dina(n4631), .dinb(n2937), .dout(n4632));
  jnot g3991(.din(n4394), .dout(n4633));
  jand g3992(.dina(n4633), .dinb(n4632), .dout(n4634));
  jor  g3993(.dina(n4407), .dinb(n4634), .dout(n4635));
  jor  g3994(.dina(n4635), .dinb(n2897), .dout(n4636));
  jnot g3995(.din(n4413), .dout(n4637));
  jand g3996(.dina(n4637), .dinb(n4636), .dout(n4638));
  jor  g3997(.dina(n4638), .dinb(n2888), .dout(n4639));
  jand g3998(.dina(n4453), .dinb(n4639), .dout(n4640));
  jor  g3999(.dina(n4468), .dinb(n4640), .dout(n4641));
  jand g4000(.dina(n4641), .dinb(n4479), .dout(n4642));
  jor  g4001(.dina(n4642), .dinb(n2837), .dout(n4643));
  jand g4002(.dina(n4643), .dinb(n4478), .dout(n4644));
  jor  g4003(.dina(n4644), .dinb(n2641), .dout(n4645));
  jnot g4004(.din(n2643), .dout(n4646));
  jor  g4005(.dina(n4644), .dinb(n4646), .dout(n4647));
  jand g4006(.dina(n4647), .dinb(n4645), .dout(n4648));
  jor  g4007(.dina(n4648), .dinb(n3771), .dout(n4649));
  jand g4008(.dina(n4649), .dinb(n4477), .dout(\result[0] ));
  jor  g4009(.dina(\address[1] ), .dinb(n4506), .dout(n4651));
  jor  g4010(.dina(n4648), .dinb(n3761), .dout(n4652));
  jand g4011(.dina(n4652), .dinb(n4651), .dout(\result[1] ));
  jor  g4012(.dina(\address[1] ), .dinb(n4515), .dout(n4654));
  jor  g4013(.dina(n4648), .dinb(n3779), .dout(n4655));
  jand g4014(.dina(n4655), .dinb(n4654), .dout(\result[2] ));
  jor  g4015(.dina(\address[1] ), .dinb(n4526), .dout(n4657));
  jor  g4016(.dina(n4648), .dinb(n3791), .dout(n4658));
  jand g4017(.dina(n4658), .dinb(n4657), .dout(\result[3] ));
  jor  g4018(.dina(\address[1] ), .dinb(n3756), .dout(n4660));
  jor  g4019(.dina(n4648), .dinb(n3795), .dout(n4661));
  jand g4020(.dina(n4661), .dinb(n4660), .dout(\result[4] ));
  jor  g4021(.dina(\address[1] ), .dinb(n3745), .dout(n4663));
  jor  g4022(.dina(n4648), .dinb(n3748), .dout(n4664));
  jand g4023(.dina(n4664), .dinb(n4663), .dout(\result[5] ));
  jor  g4024(.dina(\address[1] ), .dinb(n3806), .dout(n4666));
  jor  g4025(.dina(n4648), .dinb(n3734), .dout(n4667));
  jand g4026(.dina(n4667), .dinb(n4666), .dout(\result[6] ));
  jor  g4027(.dina(\address[1] ), .dinb(n3804), .dout(n4669));
  jor  g4028(.dina(n4648), .dinb(n3729), .dout(n4670));
  jand g4029(.dina(n4670), .dinb(n4669), .dout(\result[7] ));
  jor  g4030(.dina(\address[1] ), .dinb(n3720), .dout(n4672));
  jor  g4031(.dina(n4648), .dinb(n3811), .dout(n4673));
  jand g4032(.dina(n4673), .dinb(n4672), .dout(\result[8] ));
  jor  g4033(.dina(\address[1] ), .dinb(n3821), .dout(n4675));
  jor  g4034(.dina(n4648), .dinb(n3826), .dout(n4676));
  jand g4035(.dina(n4676), .dinb(n4675), .dout(\result[9] ));
  jor  g4036(.dina(\address[1] ), .dinb(n3830), .dout(n4678));
  jor  g4037(.dina(n4648), .dinb(n3712), .dout(n4679));
  jand g4038(.dina(n4679), .dinb(n4678), .dout(\result[10] ));
  jor  g4039(.dina(\address[1] ), .dinb(n3835), .dout(n4681));
  jor  g4040(.dina(n4648), .dinb(n3845), .dout(n4682));
  jand g4041(.dina(n4682), .dinb(n4681), .dout(\result[11] ));
  jor  g4042(.dina(\address[1] ), .dinb(n3700), .dout(n4684));
  jor  g4043(.dina(n4648), .dinb(n3843), .dout(n4685));
  jand g4044(.dina(n4685), .dinb(n4684), .dout(\result[12] ));
  jor  g4045(.dina(\address[1] ), .dinb(n3689), .dout(n4687));
  jor  g4046(.dina(n4648), .dinb(n3695), .dout(n4688));
  jand g4047(.dina(n4688), .dinb(n4687), .dout(\result[13] ));
  jor  g4048(.dina(\address[1] ), .dinb(n3855), .dout(n4690));
  jor  g4049(.dina(n4648), .dinb(n3684), .dout(n4691));
  jand g4050(.dina(n4691), .dinb(n4690), .dout(\result[14] ));
  jor  g4051(.dina(\address[1] ), .dinb(n3853), .dout(n4693));
  jor  g4052(.dina(n4648), .dinb(n3676), .dout(n4694));
  jand g4053(.dina(n4694), .dinb(n4693), .dout(\result[15] ));
  jor  g4054(.dina(\address[1] ), .dinb(n3667), .dout(n4696));
  jor  g4055(.dina(n4648), .dinb(n3860), .dout(n4697));
  jand g4056(.dina(n4697), .dinb(n4696), .dout(\result[16] ));
  jor  g4057(.dina(\address[1] ), .dinb(n3870), .dout(n4699));
  jor  g4058(.dina(n4648), .dinb(n3875), .dout(n4700));
  jand g4059(.dina(n4700), .dinb(n4699), .dout(\result[17] ));
  jor  g4060(.dina(\address[1] ), .dinb(n3879), .dout(n4702));
  jor  g4061(.dina(n4648), .dinb(n3659), .dout(n4703));
  jand g4062(.dina(n4703), .dinb(n4702), .dout(\result[18] ));
  jor  g4063(.dina(\address[1] ), .dinb(n3881), .dout(n4705));
  jor  g4064(.dina(n4648), .dinb(n3651), .dout(n4706));
  jand g4065(.dina(n4706), .dinb(n4705), .dout(\result[19] ));
  jor  g4066(.dina(\address[1] ), .dinb(n3642), .dout(n4708));
  jor  g4067(.dina(n4648), .dinb(n3640), .dout(n4709));
  jand g4068(.dina(n4709), .dinb(n4708), .dout(\result[20] ));
  jor  g4069(.dina(\address[1] ), .dinb(n3898), .dout(n4711));
  jor  g4070(.dina(n4648), .dinb(n3894), .dout(n4712));
  jand g4071(.dina(n4712), .dinb(n4711), .dout(\result[21] ));
  jor  g4072(.dina(\address[1] ), .dinb(n3900), .dout(n4714));
  jor  g4073(.dina(n4648), .dinb(n3632), .dout(n4715));
  jand g4074(.dina(n4715), .dinb(n4714), .dout(\result[22] ));
  jor  g4075(.dina(\address[1] ), .dinb(n3620), .dout(n4717));
  jor  g4076(.dina(n4648), .dinb(n3907), .dout(n4718));
  jand g4077(.dina(n4718), .dinb(n4717), .dout(\result[23] ));
  jor  g4078(.dina(\address[1] ), .dinb(n3605), .dout(n4720));
  jor  g4079(.dina(n4648), .dinb(n3909), .dout(n4721));
  jand g4080(.dina(n4721), .dinb(n4720), .dout(\result[24] ));
  jor  g4081(.dina(\address[1] ), .dinb(n3613), .dout(n4723));
  jor  g4082(.dina(n4648), .dinb(n3914), .dout(n4724));
  jand g4083(.dina(n4724), .dinb(n4723), .dout(\result[25] ));
  jor  g4084(.dina(\address[1] ), .dinb(n3918), .dout(n4726));
  jor  g4085(.dina(n4648), .dinb(n3597), .dout(n4727));
  jand g4086(.dina(n4727), .dinb(n4726), .dout(\result[26] ));
  jor  g4087(.dina(\address[1] ), .dinb(n3923), .dout(n4729));
  jor  g4088(.dina(n4648), .dinb(n3933), .dout(n4730));
  jand g4089(.dina(n4730), .dinb(n4729), .dout(\result[27] ));
  jor  g4090(.dina(\address[1] ), .dinb(n3585), .dout(n4732));
  jor  g4091(.dina(n4648), .dinb(n3931), .dout(n4733));
  jand g4092(.dina(n4733), .dinb(n4732), .dout(\result[28] ));
  jor  g4093(.dina(\address[1] ), .dinb(n3947), .dout(n4735));
  jor  g4094(.dina(n4648), .dinb(n3580), .dout(n4736));
  jand g4095(.dina(n4736), .dinb(n4735), .dout(\result[29] ));
  jor  g4096(.dina(\address[1] ), .dinb(n3942), .dout(n4738));
  jor  g4097(.dina(n4648), .dinb(n3954), .dout(n4739));
  jand g4098(.dina(n4739), .dinb(n4738), .dout(\result[30] ));
  jor  g4099(.dina(\address[1] ), .dinb(n3568), .dout(n4741));
  jor  g4100(.dina(n4648), .dinb(n3952), .dout(n4742));
  jand g4101(.dina(n4742), .dinb(n4741), .dout(\result[31] ));
  jor  g4102(.dina(\address[1] ), .dinb(n3541), .dout(n4744));
  jor  g4103(.dina(n4648), .dinb(n3960), .dout(n4745));
  jand g4104(.dina(n4745), .dinb(n4744), .dout(\result[32] ));
  jor  g4105(.dina(\address[1] ), .dinb(n3543), .dout(n4747));
  jor  g4106(.dina(n4648), .dinb(n3523), .dout(n4748));
  jand g4107(.dina(n4748), .dinb(n4747), .dout(\result[33] ));
  jor  g4108(.dina(\address[1] ), .dinb(n3549), .dout(n4750));
  jor  g4109(.dina(n4648), .dinb(n3528), .dout(n4751));
  jand g4110(.dina(n4751), .dinb(n4750), .dout(\result[34] ));
  jor  g4111(.dina(\address[1] ), .dinb(n3547), .dout(n4753));
  jor  g4112(.dina(n4648), .dinb(n3514), .dout(n4754));
  jand g4113(.dina(n4754), .dinb(n4753), .dout(\result[35] ));
  jor  g4114(.dina(\address[1] ), .dinb(n3499), .dout(n4756));
  jor  g4115(.dina(n4648), .dinb(n3505), .dout(n4757));
  jand g4116(.dina(n4757), .dinb(n4756), .dout(\result[36] ));
  jor  g4117(.dina(\address[1] ), .dinb(n3494), .dout(n4759));
  jor  g4118(.dina(n4648), .dinb(n3490), .dout(n4760));
  jand g4119(.dina(n4760), .dinb(n4759), .dout(\result[37] ));
  jor  g4120(.dina(\address[1] ), .dinb(n3559), .dout(n4762));
  jor  g4121(.dina(n4648), .dinb(n3479), .dout(n4763));
  jand g4122(.dina(n4763), .dinb(n4762), .dout(\result[38] ));
  jor  g4123(.dina(\address[1] ), .dinb(n3557), .dout(n4765));
  jor  g4124(.dina(n4648), .dinb(n3473), .dout(n4766));
  jand g4125(.dina(n4766), .dinb(n4765), .dout(\result[39] ));
  jor  g4126(.dina(\address[1] ), .dinb(n4005), .dout(n4768));
  jor  g4127(.dina(n4648), .dinb(n3984), .dout(n4769));
  jand g4128(.dina(n4769), .dinb(n4768), .dout(\result[40] ));
  jor  g4129(.dina(\address[1] ), .dinb(n4008), .dout(n4771));
  jor  g4130(.dina(n4648), .dinb(n3976), .dout(n4772));
  jand g4131(.dina(n4772), .dinb(n4771), .dout(\result[41] ));
  jor  g4132(.dina(\address[1] ), .dinb(n4002), .dout(n4774));
  jor  g4133(.dina(n4648), .dinb(n3992), .dout(n4775));
  jand g4134(.dina(n4775), .dinb(n4774), .dout(\result[42] ));
  jor  g4135(.dina(\address[1] ), .dinb(n3463), .dout(n4777));
  jnot g4136(.din(n3421), .dout(n4778));
  jor  g4137(.dina(n4648), .dinb(n4778), .dout(n4779));
  jand g4138(.dina(n4779), .dinb(n4777), .dout(\result[43] ));
  jor  g4139(.dina(\address[1] ), .dinb(n4015), .dout(n4781));
  jor  g4140(.dina(n4648), .dinb(n3428), .dout(n4782));
  jand g4141(.dina(n4782), .dinb(n4781), .dout(\result[44] ));
  jor  g4142(.dina(\address[1] ), .dinb(n4013), .dout(n4784));
  jor  g4143(.dina(n4648), .dinb(n3455), .dout(n4785));
  jand g4144(.dina(n4785), .dinb(n4784), .dout(\result[45] ));
  jor  g4145(.dina(\address[1] ), .dinb(n4023), .dout(n4787));
  jor  g4146(.dina(n4648), .dinb(n3442), .dout(n4788));
  jand g4147(.dina(n4788), .dinb(n4787), .dout(\result[46] ));
  jor  g4148(.dina(\address[1] ), .dinb(n4021), .dout(n4790));
  jor  g4149(.dina(n4648), .dinb(n3437), .dout(n4791));
  jand g4150(.dina(n4791), .dinb(n4790), .dout(\result[47] ));
  jor  g4151(.dina(\address[1] ), .dinb(n4108), .dout(n4793));
  jor  g4152(.dina(n4648), .dinb(n4080), .dout(n4794));
  jand g4153(.dina(n4794), .dinb(n4793), .dout(\result[48] ));
  jor  g4154(.dina(\address[1] ), .dinb(n4110), .dout(n4796));
  jor  g4155(.dina(n4648), .dinb(n4038), .dout(n4797));
  jand g4156(.dina(n4797), .dinb(n4796), .dout(\result[49] ));
  jor  g4157(.dina(\address[1] ), .dinb(n4116), .dout(n4799));
  jor  g4158(.dina(n4648), .dinb(n4043), .dout(n4800));
  jand g4159(.dina(n4800), .dinb(n4799), .dout(\result[50] ));
  jor  g4160(.dina(\address[1] ), .dinb(n4114), .dout(n4802));
  jor  g4161(.dina(n4648), .dinb(n4091), .dout(n4803));
  jand g4162(.dina(n4803), .dinb(n4802), .dout(\result[51] ));
  jor  g4163(.dina(\address[1] ), .dinb(n4104), .dout(n4805));
  jor  g4164(.dina(n4648), .dinb(n4052), .dout(n4806));
  jand g4165(.dina(n4806), .dinb(n4805), .dout(\result[52] ));
  jor  g4166(.dina(\address[1] ), .dinb(n4099), .dout(n4808));
  jor  g4167(.dina(n4648), .dinb(n4063), .dout(n4809));
  jand g4168(.dina(n4809), .dinb(n4808), .dout(\result[53] ));
  jor  g4169(.dina(\address[1] ), .dinb(n4101), .dout(n4811));
  jor  g4170(.dina(n4648), .dinb(n4071), .dout(n4812));
  jand g4171(.dina(n4812), .dinb(n4811), .dout(\result[54] ));
  jor  g4172(.dina(\address[1] ), .dinb(n3413), .dout(n4814));
  jor  g4173(.dina(n4648), .dinb(n4066), .dout(n4815));
  jand g4174(.dina(n4815), .dinb(n4814), .dout(\result[55] ));
  jor  g4175(.dina(\address[1] ), .dinb(n3396), .dout(n4817));
  jor  g4176(.dina(n4648), .dinb(n4129), .dout(n4818));
  jand g4177(.dina(n4818), .dinb(n4817), .dout(\result[56] ));
  jor  g4178(.dina(\address[1] ), .dinb(n3402), .dout(n4820));
  jor  g4179(.dina(n4648), .dinb(n3390), .dout(n4821));
  jand g4180(.dina(n4821), .dinb(n4820), .dout(\result[57] ));
  jor  g4181(.dina(\address[1] ), .dinb(n3382), .dout(n4823));
  jor  g4182(.dina(n4648), .dinb(n3378), .dout(n4824));
  jand g4183(.dina(n4824), .dinb(n4823), .dout(\result[58] ));
  jor  g4184(.dina(\address[1] ), .dinb(n3365), .dout(n4826));
  jor  g4185(.dina(n4648), .dinb(n3370), .dout(n4827));
  jand g4186(.dina(n4827), .dinb(n4826), .dout(\result[59] ));
  jor  g4187(.dina(\address[1] ), .dinb(n4138), .dout(n4829));
  jor  g4188(.dina(n4648), .dinb(n3332), .dout(n4830));
  jand g4189(.dina(n4830), .dinb(n4829), .dout(\result[60] ));
  jor  g4190(.dina(\address[1] ), .dinb(n4136), .dout(n4832));
  jor  g4191(.dina(n4648), .dinb(n3356), .dout(n4833));
  jand g4192(.dina(n4833), .dinb(n4832), .dout(\result[61] ));
  jor  g4193(.dina(\address[1] ), .dinb(n4145), .dout(n4835));
  jor  g4194(.dina(n4648), .dinb(n3337), .dout(n4836));
  jand g4195(.dina(n4836), .dinb(n4835), .dout(\result[62] ));
  jor  g4196(.dina(\address[1] ), .dinb(n4143), .dout(n4838));
  jor  g4197(.dina(n4648), .dinb(n3348), .dout(n4839));
  jand g4198(.dina(n4839), .dinb(n4838), .dout(\result[63] ));
  jor  g4199(.dina(\address[1] ), .dinb(n3320), .dout(n4841));
  jor  g4200(.dina(n4648), .dinb(n4153), .dout(n4842));
  jand g4201(.dina(n4842), .dinb(n4841), .dout(\result[64] ));
  jor  g4202(.dina(\address[1] ), .dinb(n3306), .dout(n4844));
  jor  g4203(.dina(n4648), .dinb(n3311), .dout(n4845));
  jand g4204(.dina(n4845), .dinb(n4844), .dout(\result[65] ));
  jor  g4205(.dina(\address[1] ), .dinb(n3301), .dout(n4847));
  jor  g4206(.dina(n4648), .dinb(n4160), .dout(n4848));
  jand g4207(.dina(n4848), .dinb(n4847), .dout(\result[66] ));
  jor  g4208(.dina(\address[1] ), .dinb(n3289), .dout(n4850));
  jor  g4209(.dina(n4648), .dinb(n4158), .dout(n4851));
  jand g4210(.dina(n4851), .dinb(n4850), .dout(\result[67] ));
  jor  g4211(.dina(\address[1] ), .dinb(n3270), .dout(n4853));
  jor  g4212(.dina(n4648), .dinb(n4165), .dout(n4854));
  jand g4213(.dina(n4854), .dinb(n4853), .dout(\result[68] ));
  jor  g4214(.dina(\address[1] ), .dinb(n3265), .dout(n4856));
  jor  g4215(.dina(n4648), .dinb(n3260), .dout(n4857));
  jand g4216(.dina(n4857), .dinb(n4856), .dout(\result[69] ));
  jor  g4217(.dina(\address[1] ), .dinb(n3280), .dout(n4859));
  jor  g4218(.dina(n4648), .dinb(n3241), .dout(n4860));
  jand g4219(.dina(n4860), .dinb(n4859), .dout(\result[70] ));
  jor  g4220(.dina(\address[1] ), .dinb(n3278), .dout(n4862));
  jor  g4221(.dina(n4648), .dinb(n3252), .dout(n4863));
  jand g4222(.dina(n4863), .dinb(n4862), .dout(\result[71] ));
  jor  g4223(.dina(\address[1] ), .dinb(n4214), .dout(n4865));
  jor  g4224(.dina(n4648), .dinb(n4173), .dout(n4866));
  jand g4225(.dina(n4866), .dinb(n4865), .dout(\result[72] ));
  jor  g4226(.dina(\address[1] ), .dinb(n4217), .dout(n4868));
  jor  g4227(.dina(n4648), .dinb(n4203), .dout(n4869));
  jand g4228(.dina(n4869), .dinb(n4868), .dout(\result[73] ));
  jor  g4229(.dina(\address[1] ), .dinb(n4212), .dout(n4871));
  jor  g4230(.dina(n4648), .dinb(n4190), .dout(n4872));
  jand g4231(.dina(n4872), .dinb(n4871), .dout(\result[74] ));
  jor  g4232(.dina(\address[1] ), .dinb(n4210), .dout(n4874));
  jor  g4233(.dina(n4648), .dinb(n4185), .dout(n4875));
  jand g4234(.dina(n4875), .dinb(n4874), .dout(\result[75] ));
  jor  g4235(.dina(\address[1] ), .dinb(n4229), .dout(n4877));
  jor  g4236(.dina(n4648), .dinb(n3209), .dout(n4878));
  jand g4237(.dina(n4878), .dinb(n4877), .dout(\result[76] ));
  jor  g4238(.dina(\address[1] ), .dinb(n4227), .dout(n4880));
  jor  g4239(.dina(n4648), .dinb(n3233), .dout(n4881));
  jand g4240(.dina(n4881), .dinb(n4880), .dout(\result[77] ));
  jor  g4241(.dina(\address[1] ), .dinb(n4236), .dout(n4883));
  jor  g4242(.dina(n4648), .dinb(n3214), .dout(n4884));
  jand g4243(.dina(n4884), .dinb(n4883), .dout(\result[78] ));
  jor  g4244(.dina(\address[1] ), .dinb(n4234), .dout(n4886));
  jor  g4245(.dina(n4648), .dinb(n3225), .dout(n4887));
  jand g4246(.dina(n4887), .dinb(n4886), .dout(\result[79] ));
  jor  g4247(.dina(\address[1] ), .dinb(n4248), .dout(n4889));
  jor  g4248(.dina(n4648), .dinb(n3196), .dout(n4890));
  jand g4249(.dina(n4890), .dinb(n4889), .dout(\result[80] ));
  jor  g4250(.dina(\address[1] ), .dinb(n4251), .dout(n4892));
  jor  g4251(.dina(n4648), .dinb(n3191), .dout(n4893));
  jand g4252(.dina(n4893), .dinb(n4892), .dout(\result[81] ));
  jor  g4253(.dina(\address[1] ), .dinb(n4245), .dout(n4895));
  jor  g4254(.dina(n4648), .dinb(n3179), .dout(n4896));
  jand g4255(.dina(n4896), .dinb(n4895), .dout(\result[82] ));
  jor  g4256(.dina(\address[1] ), .dinb(n3168), .dout(n4898));
  jor  g4257(.dina(n4648), .dinb(n3174), .dout(n4899));
  jand g4258(.dina(n4899), .dinb(n4898), .dout(\result[83] ));
  jor  g4259(.dina(\address[1] ), .dinb(n3149), .dout(n4901));
  jor  g4260(.dina(n4648), .dinb(n4259), .dout(n4902));
  jand g4261(.dina(n4902), .dinb(n4901), .dout(\result[84] ));
  jor  g4262(.dina(\address[1] ), .dinb(n3144), .dout(n4904));
  jor  g4263(.dina(n4648), .dinb(n3139), .dout(n4905));
  jand g4264(.dina(n4905), .dinb(n4904), .dout(\result[85] ));
  jor  g4265(.dina(\address[1] ), .dinb(n3160), .dout(n4907));
  jor  g4266(.dina(n4648), .dinb(n3120), .dout(n4908));
  jand g4267(.dina(n4908), .dinb(n4907), .dout(\result[86] ));
  jor  g4268(.dina(\address[1] ), .dinb(n3158), .dout(n4910));
  jor  g4269(.dina(n4648), .dinb(n3131), .dout(n4911));
  jand g4270(.dina(n4911), .dinb(n4910), .dout(\result[87] ));
  jor  g4271(.dina(\address[1] ), .dinb(n4272), .dout(n4913));
  jor  g4272(.dina(n4648), .dinb(n3110), .dout(n4914));
  jand g4273(.dina(n4914), .dinb(n4913), .dout(\result[88] ));
  jor  g4274(.dina(\address[1] ), .dinb(n4275), .dout(n4916));
  jor  g4275(.dina(n4648), .dinb(n3105), .dout(n4917));
  jand g4276(.dina(n4917), .dinb(n4916), .dout(\result[89] ));
  jor  g4277(.dina(\address[1] ), .dinb(n4269), .dout(n4919));
  jor  g4278(.dina(n4648), .dinb(n3093), .dout(n4920));
  jand g4279(.dina(n4920), .dinb(n4919), .dout(\result[90] ));
  jor  g4280(.dina(\address[1] ), .dinb(n4266), .dout(n4922));
  jor  g4281(.dina(n4648), .dinb(n3088), .dout(n4923));
  jand g4282(.dina(n4923), .dinb(n4922), .dout(\result[91] ));
  jor  g4283(.dina(\address[1] ), .dinb(n4287), .dout(n4925));
  jor  g4284(.dina(n4648), .dinb(n3053), .dout(n4926));
  jand g4285(.dina(n4926), .dinb(n4925), .dout(\result[92] ));
  jor  g4286(.dina(\address[1] ), .dinb(n4285), .dout(n4928));
  jor  g4287(.dina(n4648), .dinb(n3077), .dout(n4929));
  jand g4288(.dina(n4929), .dinb(n4928), .dout(\result[93] ));
  jor  g4289(.dina(\address[1] ), .dinb(n4294), .dout(n4931));
  jor  g4290(.dina(n4648), .dinb(n3058), .dout(n4932));
  jand g4291(.dina(n4932), .dinb(n4931), .dout(\result[94] ));
  jor  g4292(.dina(\address[1] ), .dinb(n4292), .dout(n4934));
  jor  g4293(.dina(n4648), .dinb(n3069), .dout(n4935));
  jand g4294(.dina(n4935), .dinb(n4934), .dout(\result[95] ));
  jor  g4295(.dina(\address[1] ), .dinb(n4308), .dout(n4937));
  jor  g4296(.dina(n4648), .dinb(n3040), .dout(n4938));
  jand g4297(.dina(n4938), .dinb(n4937), .dout(\result[96] ));
  jor  g4298(.dina(\address[1] ), .dinb(n4311), .dout(n4940));
  jor  g4299(.dina(n4648), .dinb(n3035), .dout(n4941));
  jand g4300(.dina(n4941), .dinb(n4940), .dout(\result[97] ));
  jor  g4301(.dina(\address[1] ), .dinb(n4305), .dout(n4943));
  jor  g4302(.dina(n4648), .dinb(n3023), .dout(n4944));
  jand g4303(.dina(n4944), .dinb(n4943), .dout(\result[98] ));
  jor  g4304(.dina(\address[1] ), .dinb(n4302), .dout(n4946));
  jor  g4305(.dina(n4648), .dinb(n3018), .dout(n4947));
  jand g4306(.dina(n4947), .dinb(n4946), .dout(\result[99] ));
  jor  g4307(.dina(\address[1] ), .dinb(n4323), .dout(n4949));
  jor  g4308(.dina(n4648), .dinb(n2983), .dout(n4950));
  jand g4309(.dina(n4950), .dinb(n4949), .dout(\result[100] ));
  jor  g4310(.dina(\address[1] ), .dinb(n4321), .dout(n4952));
  jor  g4311(.dina(n4648), .dinb(n3007), .dout(n4953));
  jand g4312(.dina(n4953), .dinb(n4952), .dout(\result[101] ));
  jor  g4313(.dina(\address[1] ), .dinb(n4330), .dout(n4955));
  jor  g4314(.dina(n4648), .dinb(n2988), .dout(n4956));
  jand g4315(.dina(n4956), .dinb(n4955), .dout(\result[102] ));
  jor  g4316(.dina(\address[1] ), .dinb(n4328), .dout(n4958));
  jor  g4317(.dina(n4648), .dinb(n2999), .dout(n4959));
  jand g4318(.dina(n4959), .dinb(n4958), .dout(\result[103] ));
  jor  g4319(.dina(\address[1] ), .dinb(n4344), .dout(n4961));
  jor  g4320(.dina(n4648), .dinb(n2970), .dout(n4962));
  jand g4321(.dina(n4962), .dinb(n4961), .dout(\result[104] ));
  jor  g4322(.dina(\address[1] ), .dinb(n4347), .dout(n4964));
  jor  g4323(.dina(n4648), .dinb(n2965), .dout(n4965));
  jand g4324(.dina(n4965), .dinb(n4964), .dout(\result[105] ));
  jor  g4325(.dina(\address[1] ), .dinb(n4341), .dout(n4967));
  jor  g4326(.dina(n4648), .dinb(n2953), .dout(n4968));
  jand g4327(.dina(n4968), .dinb(n4967), .dout(\result[106] ));
  jor  g4328(.dina(\address[1] ), .dinb(n4338), .dout(n4970));
  jor  g4329(.dina(n4648), .dinb(n2948), .dout(n4971));
  jand g4330(.dina(n4971), .dinb(n4970), .dout(\result[107] ));
  jor  g4331(.dina(\address[1] ), .dinb(n2931), .dout(n4973));
  jor  g4332(.dina(n4648), .dinb(n2939), .dout(n4974));
  jand g4333(.dina(n4974), .dinb(n4973), .dout(\result[108] ));
  jor  g4334(.dina(\address[1] ), .dinb(n2926), .dout(n4976));
  jor  g4335(.dina(n4648), .dinb(n2921), .dout(n4977));
  jand g4336(.dina(n4977), .dinb(n4976), .dout(\result[109] ));
  jor  g4337(.dina(\address[1] ), .dinb(n4359), .dout(n4979));
  jor  g4338(.dina(n4648), .dinb(n2902), .dout(n4980));
  jand g4339(.dina(n4980), .dinb(n4979), .dout(\result[110] ));
  jor  g4340(.dina(\address[1] ), .dinb(n4357), .dout(n4982));
  jor  g4341(.dina(n4648), .dinb(n2913), .dout(n4983));
  jand g4342(.dina(n4983), .dinb(n4982), .dout(\result[111] ));
  jor  g4343(.dina(\address[1] ), .dinb(n4400), .dout(n4985));
  jor  g4344(.dina(n4648), .dinb(n4388), .dout(n4986));
  jand g4345(.dina(n4986), .dinb(n4985), .dout(\result[112] ));
  jor  g4346(.dina(\address[1] ), .dinb(n4403), .dout(n4988));
  jor  g4347(.dina(n4648), .dinb(n4372), .dout(n4989));
  jand g4348(.dina(n4989), .dinb(n4988), .dout(\result[113] ));
  jor  g4349(.dina(\address[1] ), .dinb(n4397), .dout(n4991));
  jor  g4350(.dina(n4648), .dinb(n4379), .dout(n4992));
  jand g4351(.dina(n4992), .dinb(n4991), .dout(\result[114] ));
  jor  g4352(.dina(\address[1] ), .dinb(n2893), .dout(n4994));
  jor  g4353(.dina(n4648), .dinb(n4374), .dout(n4995));
  jand g4354(.dina(n4995), .dinb(n4994), .dout(\result[115] ));
  jor  g4355(.dina(\address[1] ), .dinb(n2874), .dout(n4997));
  jor  g4356(.dina(n4648), .dinb(n4411), .dout(n4998));
  jand g4357(.dina(n4998), .dinb(n4997), .dout(\result[116] ));
  jor  g4358(.dina(\address[1] ), .dinb(n2869), .dout(n5000));
  jor  g4359(.dina(n4648), .dinb(n2864), .dout(n5001));
  jand g4360(.dina(n5001), .dinb(n5000), .dout(\result[117] ));
  jor  g4361(.dina(\address[1] ), .dinb(n2884), .dout(n5003));
  jor  g4362(.dina(n4648), .dinb(n2845), .dout(n5004));
  jand g4363(.dina(n5004), .dinb(n5003), .dout(\result[118] ));
  jor  g4364(.dina(\address[1] ), .dinb(n2882), .dout(n5006));
  jor  g4365(.dina(n4648), .dinb(n2856), .dout(n5007));
  jand g4366(.dina(n5007), .dinb(n5006), .dout(\result[119] ));
  jor  g4367(.dina(\address[1] ), .dinb(n4460), .dout(n5009));
  jor  g4368(.dina(n4648), .dinb(n4419), .dout(n5010));
  jand g4369(.dina(n5010), .dinb(n5009), .dout(\result[120] ));
  jor  g4370(.dina(\address[1] ), .dinb(n4463), .dout(n5012));
  jor  g4371(.dina(n4648), .dinb(n4449), .dout(n5013));
  jand g4372(.dina(n5013), .dinb(n5012), .dout(\result[121] ));
  jor  g4373(.dina(\address[1] ), .dinb(n4458), .dout(n5015));
  jor  g4374(.dina(n4648), .dinb(n4436), .dout(n5016));
  jand g4375(.dina(n5016), .dinb(n5015), .dout(\result[122] ));
  jor  g4376(.dina(\address[1] ), .dinb(n4456), .dout(n5018));
  jor  g4377(.dina(n4648), .dinb(n4431), .dout(n5019));
  jand g4378(.dina(n5019), .dinb(n5018), .dout(\result[123] ));
  jor  g4379(.dina(\address[1] ), .dinb(n2826), .dout(n5021));
  jor  g4380(.dina(n4648), .dinb(n2839), .dout(n5022));
  jand g4381(.dina(n5022), .dinb(n5021), .dout(\result[124] ));
  jor  g4382(.dina(\address[1] ), .dinb(n2831), .dout(n5024));
  jor  g4383(.dina(n4648), .dinb(n2819), .dout(n5025));
  jand g4384(.dina(n5025), .dinb(n5024), .dout(\result[125] ));
  jor  g4385(.dina(\address[1] ), .dinb(n2835), .dout(n5027));
  jor  g4386(.dina(n4648), .dinb(n2811), .dout(n5028));
  jand g4387(.dina(n5028), .dinb(n5027), .dout(\result[126] ));
  jand g4388(.dina(n2643), .dinb(n2641), .dout(\result[127] ));
  jor  g4389(.dina(\address[1] ), .dinb(n1562), .dout(n5031));
  jor  g4390(.dina(n4648), .dinb(n2808), .dout(n5032));
  jand g4391(.dina(n5032), .dinb(n5031), .dout(\address[0] ));
endmodule


