module rf_c432(G115gat, G108gat, G102gat, G99gat, G112gat, G95gat, G92gat, G105gat, G37gat, G4gat, G69gat, G17gat, G34gat, G1gat, G79gat, G30gat, G14gat, G21gat, G53gat, G60gat, G8gat, G63gat, G11gat, G24gat, G40gat, G43gat, G82gat, G47gat, G50gat, G56gat, G66gat, G73gat, G89gat, G76gat, G27gat, G86gat, G432gat, G430gat, G421gat, G431gat, G370gat, G329gat, G223gat);
    input G115gat, G108gat, G102gat, G99gat, G112gat, G95gat, G92gat, G105gat, G37gat, G4gat, G69gat, G17gat, G34gat, G1gat, G79gat, G30gat, G14gat, G21gat, G53gat, G60gat, G8gat, G63gat, G11gat, G24gat, G40gat, G43gat, G82gat, G47gat, G50gat, G56gat, G66gat, G73gat, G89gat, G76gat, G27gat, G86gat;
    output G432gat, G430gat, G421gat, G431gat, G370gat, G329gat, G223gat;
    wire n45;
    wire n49;
    wire n52;
    wire n56;
    wire n59;
    wire n63;
    wire n67;
    wire n71;
    wire n74;
    wire n78;
    wire n81;
    wire n85;
    wire n89;
    wire n92;
    wire n96;
    wire n99;
    wire n103;
    wire n107;
    wire n110;
    wire n114;
    wire n117;
    wire n121;
    wire n125;
    wire n129;
    wire n133;
    wire n137;
    wire n140;
    wire n143;
    wire n146;
    wire n150;
    wire n153;
    wire n157;
    wire n161;
    wire n165;
    wire n168;
    wire n172;
    wire n175;
    wire n179;
    wire n183;
    wire n186;
    wire n190;
    wire n193;
    wire n197;
    wire n201;
    wire n204;
    wire n208;
    wire n211;
    wire n215;
    wire n219;
    wire n223;
    wire n227;
    wire n231;
    wire n235;
    wire n239;
    wire n243;
    wire n246;
    wire n250;
    wire n254;
    wire n258;
    wire n262;
    wire n265;
    wire n269;
    wire n273;
    wire n277;
    wire n280;
    wire n284;
    wire n288;
    wire n292;
    wire n296;
    wire n300;
    wire n304;
    wire n308;
    wire n312;
    wire n315;
    wire n318;
    wire n322;
    wire n326;
    wire n330;
    wire n334;
    wire n337;
    wire n341;
    wire n345;
    wire n349;
    wire n352;
    wire n356;
    wire n360;
    wire n364;
    wire n367;
    wire n371;
    wire n375;
    wire n379;
    wire n383;
    wire n387;
    wire n391;
    wire n395;
    wire n399;
    wire n403;
    wire n407;
    wire n411;
    wire n415;
    wire n418;
    wire n422;
    wire n426;
    wire n430;
    wire n434;
    wire n437;
    wire n440;
    wire n444;
    wire n448;
    wire n451;
    wire n455;
    wire n459;
    wire n463;
    wire n467;
    wire n471;
    wire n475;
    wire n479;
    wire n483;
    wire n487;
    wire n491;
    wire n495;
    wire n499;
    wire n503;
    wire n507;
    wire n510;
    wire n514;
    wire n518;
    wire n521;
    wire n525;
    wire n529;
    wire n533;
    wire n537;
    wire n541;
    wire n545;
    wire n549;
    wire n553;
    wire n557;
    wire n561;
    wire n565;
    wire n569;
    wire n573;
    wire n577;
    wire n581;
    wire n585;
    wire n588;
    wire n591;
    wire n595;
    wire n599;
    wire n603;
    wire n607;
    wire n611;
    wire n614;
    wire n618;
    wire n622;
    wire n626;
    wire n630;
    wire n634;
    wire n638;
    wire n641;
    wire n645;
    wire n649;
    wire n653;
    wire n656;
    wire n660;
    wire n664;
    wire n668;
    wire n672;
    wire n675;
    wire n679;
    wire n682;
    wire n685;
    wire n689;
    wire n693;
    wire n696;
    wire n700;
    wire n704;
    wire n708;
    wire n712;
    wire n716;
    wire n720;
    wire n724;
    wire n728;
    wire n732;
    wire n736;
    wire n740;
    wire n743;
    wire n747;
    wire n751;
    wire n755;
    wire n759;
    wire n763;
    wire n767;
    wire n770;
    wire n774;
    wire n778;
    wire n782;
    wire n786;
    wire n790;
    wire n794;
    wire n798;
    wire n802;
    wire n806;
    wire n810;
    wire n814;
    wire n818;
    wire n822;
    wire n826;
    wire n830;
    wire n833;
    wire n837;
    wire n841;
    wire n845;
    wire n849;
    wire n853;
    wire n857;
    wire n861;
    wire n865;
    wire n869;
    wire n873;
    wire n877;
    wire n880;
    wire n884;
    wire n888;
    wire n892;
    wire n896;
    wire n900;
    wire n904;
    wire n907;
    wire n911;
    wire n915;
    wire n919;
    wire n923;
    wire n927;
    wire n931;
    wire n934;
    wire n938;
    wire n942;
    wire n946;
    wire n950;
    wire n954;
    wire n958;
    wire n962;
    wire n966;
    wire n969;
    wire n972;
    wire n976;
    wire n980;
    wire n984;
    wire n988;
    wire n992;
    wire n996;
    wire n1000;
    wire n1008;
    wire n1012;
    wire n1016;
    wire n1020;
    wire n1024;
    wire n1028;
    wire n1032;
    wire n1036;
    wire n1040;
    wire n1044;
    wire n1048;
    wire n1056;
    wire n1060;
    wire n1064;
    wire n1068;
    wire n1072;
    wire n1076;
    wire n1080;
    wire n1084;
    wire n1574;
    wire n1577;
    wire n1580;
    wire n1583;
    wire n1586;
    wire n1589;
    wire n1592;
    wire n1595;
    wire n1598;
    wire n1600;
    wire n1604;
    wire n1607;
    wire n1610;
    wire n1613;
    wire n1616;
    wire n1618;
    wire n1622;
    wire n1625;
    wire n1628;
    wire n1631;
    wire n1634;
    wire n1637;
    wire n1639;
    wire n1642;
    wire n1645;
    wire n1648;
    wire n1651;
    wire n1654;
    wire n1657;
    wire n1661;
    wire n1664;
    wire n1667;
    wire n1670;
    wire n1673;
    wire n1676;
    wire n1679;
    wire n1682;
    wire n1685;
    wire n1688;
    wire n1691;
    wire n1694;
    wire n1697;
    wire n1700;
    wire n1703;
    wire n1706;
    wire n1709;
    wire n1712;
    wire n1715;
    wire n1718;
    wire n1721;
    wire n1724;
    wire n1727;
    wire n1730;
    wire n1733;
    wire n1736;
    wire n1739;
    wire n1742;
    wire n1745;
    wire n1748;
    wire n1750;
    wire n1753;
    wire n1756;
    wire n1759;
    wire n1762;
    wire n1765;
    wire n1769;
    wire n1772;
    wire n1775;
    wire n1778;
    wire n1781;
    wire n1784;
    wire n1787;
    wire n1790;
    wire n1793;
    wire n1796;
    wire n1799;
    wire n1801;
    wire n1804;
    wire n1807;
    wire n1810;
    wire n1813;
    wire n1816;
    wire n1819;
    wire n1822;
    wire n1825;
    wire n1828;
    wire n1831;
    wire n1834;
    wire n1837;
    wire n1840;
    wire n1843;
    wire n1846;
    wire n1849;
    wire n1852;
    wire n1856;
    wire n1859;
    wire n1862;
    wire n1865;
    wire n1868;
    wire n1871;
    wire n1874;
    wire n1877;
    wire n1880;
    wire n1882;
    wire n1885;
    wire n1888;
    wire n1891;
    wire n1894;
    wire n1897;
    wire n1900;
    wire n1903;
    wire n1906;
    wire n1909;
    wire n1912;
    wire n1916;
    wire n1919;
    wire n1922;
    wire n1925;
    wire n1928;
    wire n1931;
    wire n1934;
    wire n1937;
    wire n1940;
    wire n1943;
    wire n1946;
    wire n1949;
    wire n1952;
    wire n1955;
    wire n1957;
    wire n1960;
    wire n1963;
    wire n1966;
    wire n1969;
    wire n1972;
    wire n1975;
    wire n1978;
    wire n1981;
    wire n1984;
    wire n1987;
    wire n1990;
    wire n1993;
    wire n1996;
    wire n1999;
    wire n2002;
    wire n2005;
    wire n2008;
    wire n2011;
    wire n2014;
    wire n2017;
    wire n2020;
    wire n2023;
    wire n2026;
    wire n2029;
    wire n2032;
    wire n2035;
    wire n2038;
    wire n2041;
    wire n2044;
    wire n2048;
    wire n2051;
    wire n2054;
    wire n2057;
    wire n2060;
    wire n2063;
    wire n2066;
    wire n2069;
    wire n2071;
    wire n2074;
    wire n2077;
    wire n2080;
    wire n2083;
    wire n2086;
    wire n2089;
    wire n2092;
    wire n2095;
    wire n2098;
    wire n2101;
    wire n2104;
    wire n2107;
    wire n2110;
    wire n2113;
    wire n2116;
    wire n2119;
    wire n2122;
    wire n2125;
    wire n2128;
    wire n2132;
    wire n2135;
    wire n2138;
    wire n2141;
    wire n2144;
    wire n2147;
    wire n2150;
    wire n2153;
    wire n2156;
    wire n2159;
    wire n2162;
    wire n2165;
    wire n2168;
    wire n2171;
    wire n2174;
    wire n2177;
    wire n2180;
    wire n2183;
    wire n2186;
    wire n2189;
    wire n2192;
    wire n2195;
    wire n2198;
    wire n2201;
    wire n2204;
    wire n2207;
    wire n2209;
    wire n2212;
    wire n2215;
    wire n2218;
    wire n2221;
    wire n2224;
    wire n2227;
    wire n2230;
    wire n2233;
    wire n2236;
    wire n2239;
    wire n2242;
    wire n2245;
    wire n2248;
    wire n2251;
    wire n2254;
    wire n2257;
    wire n2260;
    wire n2263;
    wire n2266;
    wire n2269;
    wire n2272;
    wire n2275;
    wire n2278;
    wire n2281;
    wire n2284;
    wire n2287;
    wire n2290;
    wire n2293;
    wire n2296;
    wire n2299;
    wire n2302;
    wire n2305;
    wire n2308;
    wire n2311;
    wire n2314;
    wire n2317;
    wire n2320;
    wire n2323;
    wire n2326;
    wire n2329;
    wire n2333;
    wire n2336;
    wire n2339;
    wire n2342;
    wire n2345;
    wire n2348;
    wire n2351;
    wire n2354;
    wire n2357;
    wire n2360;
    wire n2363;
    wire n2366;
    wire n2369;
    wire n2371;
    wire n2374;
    wire n2377;
    wire n2380;
    wire n2383;
    wire n2386;
    wire n2389;
    wire n2392;
    wire n2395;
    wire n2398;
    wire n2401;
    wire n2404;
    wire n2407;
    wire n2410;
    wire n2413;
    wire n2416;
    wire n2419;
    wire n2422;
    wire n2425;
    wire n2428;
    wire n2431;
    wire n2434;
    wire n2437;
    wire n2440;
    wire n2443;
    wire n2446;
    wire n2449;
    wire n2452;
    wire n2455;
    wire n2458;
    wire n2461;
    wire n2464;
    wire n2467;
    wire n2470;
    wire n2473;
    wire n2476;
    wire n2479;
    wire n2482;
    wire n2485;
    wire n2488;
    wire n2491;
    wire n2494;
    wire n2497;
    wire n2500;
    wire n2503;
    wire n2506;
    wire n2510;
    wire n2513;
    wire n2516;
    wire n2519;
    wire n2522;
    wire n2525;
    wire n2528;
    wire n2531;
    wire n2534;
    wire n2537;
    wire n2540;
    wire n2543;
    wire n2546;
    wire n2548;
    wire n2551;
    wire n2554;
    wire n2557;
    wire n2560;
    wire n2563;
    wire n2566;
    wire n2569;
    wire n2572;
    wire n2575;
    wire n2578;
    wire n2581;
    wire n2584;
    wire n2587;
    wire n2590;
    wire n2593;
    wire n2596;
    wire n2599;
    wire n2602;
    wire n2605;
    wire n2608;
    wire n2611;
    wire n2614;
    wire n2617;
    wire n2620;
    wire n2623;
    wire n2626;
    wire n2630;
    wire n2633;
    wire n2636;
    wire n2639;
    wire n2642;
    wire n2644;
    wire n2647;
    wire n2650;
    wire n2653;
    wire n2656;
    wire n2659;
    wire n2662;
    wire n2665;
    wire n2668;
    wire n2671;
    wire n2674;
    wire n2677;
    wire n2680;
    wire n2683;
    wire n2686;
    wire n2689;
    wire n2692;
    wire n2695;
    wire n2698;
    wire n2701;
    wire n2704;
    wire n2707;
    wire n2710;
    wire n2713;
    wire n2716;
    wire n2719;
    wire n2722;
    wire n2725;
    wire n2728;
    wire n2731;
    wire n2734;
    wire n2737;
    wire n2740;
    wire n2743;
    wire n2746;
    wire n2749;
    wire n2752;
    wire n2755;
    wire n2758;
    wire n2761;
    wire n2764;
    wire n2767;
    wire n2770;
    wire n2773;
    wire n2776;
    wire n2780;
    wire n2782;
    wire n2785;
    wire n2788;
    wire n2791;
    wire n2794;
    wire n2797;
    wire n2800;
    wire n2803;
    wire n2806;
    wire n2809;
    wire n2812;
    wire n2815;
    wire n2819;
    wire n2822;
    wire n2825;
    wire n2828;
    wire n2831;
    wire n2834;
    wire n2836;
    wire n2839;
    wire n2842;
    wire n2845;
    wire n2849;
    wire n2852;
    wire n2855;
    wire n2858;
    wire n2861;
    wire n2863;
    wire n2866;
    wire n2869;
    wire n2872;
    wire n2875;
    wire n2878;
    wire n2881;
    wire n2884;
    wire n2887;
    wire n2890;
    wire n2893;
    wire n2896;
    wire n2899;
    wire n2902;
    wire n2905;
    wire n2908;
    wire n2911;
    wire n2914;
    wire n2917;
    wire n2920;
    wire n2923;
    wire n2926;
    wire n2929;
    wire n2933;
    wire n2936;
    wire n2939;
    wire n2942;
    wire n2945;
    wire n2948;
    wire n2951;
    wire n2954;
    wire n2957;
    wire n2960;
    wire n2963;
    wire n2966;
    wire n2969;
    wire n2972;
    wire n2974;
    wire n2977;
    wire n2980;
    wire n2983;
    wire n2986;
    wire n2989;
    wire n2992;
    wire n2995;
    wire n2998;
    wire n3001;
    wire n3004;
    wire n3007;
    wire n3010;
    wire n3013;
    wire n3016;
    wire n3019;
    wire n3022;
    wire n3025;
    wire n3028;
    wire n3031;
    wire n3034;
    wire n3037;
    wire n3040;
    wire n3043;
    wire n3046;
    wire n3049;
    wire n3052;
    wire n3055;
    wire n3058;
    wire n3061;
    wire n3064;
    wire n3067;
    wire n3070;
    wire n3074;
    wire n3077;
    wire n3080;
    wire n3083;
    wire n3086;
    wire n3089;
    wire n3092;
    wire n3094;
    wire n3097;
    wire n3100;
    wire n3103;
    wire n3106;
    wire n3109;
    wire n3112;
    wire n3115;
    wire n3118;
    wire n3121;
    wire n3124;
    wire n3127;
    wire n3130;
    wire n3133;
    wire n3136;
    wire n3139;
    wire n3142;
    wire n3145;
    wire n3148;
    wire n3151;
    wire n3154;
    wire n3157;
    wire n3160;
    wire n3163;
    wire n3166;
    wire n3169;
    wire n3172;
    wire n3175;
    wire n3178;
    wire n3181;
    wire n3184;
    wire n3188;
    wire n3191;
    wire n3193;
    wire n3196;
    wire n3199;
    wire n3202;
    wire n3205;
    wire n3208;
    wire n3211;
    wire n3214;
    wire n3217;
    wire n3220;
    wire n3223;
    wire n3226;
    wire n3229;
    wire n3232;
    wire n3235;
    wire n3238;
    wire n3242;
    wire n3245;
    wire n3248;
    wire n3251;
    wire n3254;
    wire n3257;
    wire n3260;
    wire n3262;
    wire n3265;
    wire n3268;
    wire n3271;
    wire n3274;
    wire n3277;
    wire n3280;
    wire n3283;
    wire n3286;
    wire n3289;
    wire n3292;
    wire n3295;
    wire n3298;
    wire n3301;
    wire n3304;
    wire n3307;
    wire n3310;
    wire n3313;
    wire n3316;
    wire n3319;
    wire n3322;
    wire n3325;
    wire n3328;
    wire n3331;
    wire n3334;
    wire n3337;
    wire n3340;
    wire n3343;
    wire n3346;
    wire n3349;
    wire n3352;
    wire n3355;
    wire n3358;
    wire n3361;
    wire n3364;
    wire n3367;
    wire n3370;
    wire n3373;
    wire n3376;
    wire n3379;
    wire n3382;
    wire n3385;
    wire n3388;
    wire n3391;
    wire n3394;
    wire n3397;
    wire n3400;
    wire n3403;
    wire n3406;
    wire n3409;
    wire n3413;
    wire n3416;
    wire n3419;
    wire n3422;
    wire n3425;
    wire n3428;
    wire n3431;
    wire n3433;
    wire n3436;
    wire n3439;
    wire n3442;
    wire n3445;
    wire n3448;
    wire n3451;
    wire n3454;
    wire n3457;
    wire n3460;
    wire n3463;
    wire n3466;
    wire n3469;
    wire n3472;
    wire n3475;
    wire n3478;
    wire n3481;
    wire n3484;
    wire n3487;
    wire n3490;
    wire n3493;
    wire n3496;
    wire n3499;
    wire n3502;
    wire n3505;
    wire n3508;
    wire n3511;
    wire n3514;
    wire n3517;
    wire n3520;
    wire n3523;
    wire n3526;
    wire n3529;
    wire n3532;
    wire n3536;
    wire n3538;
    wire n3541;
    wire n3544;
    wire n3547;
    wire n3550;
    wire n3553;
    wire n3556;
    wire n3559;
    wire n3562;
    wire n3565;
    wire n3568;
    wire n3571;
    wire n3574;
    wire n3577;
    wire n3580;
    wire n3583;
    wire n3586;
    wire n3589;
    wire n3593;
    wire n3596;
    wire n3599;
    wire n3602;
    wire n3605;
    wire n3608;
    wire n3611;
    wire n3613;
    wire n3616;
    wire n3619;
    wire n3622;
    wire n3625;
    wire n3628;
    wire n3631;
    wire n3634;
    wire n3637;
    wire n3640;
    wire n3643;
    wire n3646;
    wire n3649;
    wire n3652;
    wire n3655;
    wire n3658;
    wire n3661;
    wire n3664;
    wire n3667;
    wire n3670;
    wire n3673;
    wire n3676;
    wire n3679;
    wire n3682;
    wire n3685;
    wire n3688;
    wire n3691;
    wire n3694;
    wire n3697;
    wire n3700;
    wire n3703;
    wire n3706;
    wire n3709;
    wire n3712;
    wire n3715;
    wire n3718;
    wire n3721;
    wire n3724;
    wire n3727;
    wire n3730;
    wire n3733;
    wire n3736;
    wire n3739;
    wire n3742;
    wire n3745;
    wire n3748;
    wire n3751;
    wire n3754;
    wire n3757;
    wire n3760;
    wire n3763;
    wire n3766;
    wire n3769;
    wire n3772;
    wire n3775;
    wire n3778;
    wire n3781;
    wire n3784;
    wire n3787;
    wire n3790;
    wire n3793;
    wire n3797;
    wire n3800;
    wire n3803;
    wire n3806;
    wire n3809;
    wire n3812;
    wire n3815;
    wire n3817;
    wire n3820;
    wire n3823;
    wire n3826;
    wire n3829;
    wire n3832;
    wire n3835;
    wire n3838;
    wire n3841;
    wire n3844;
    wire n3847;
    wire n3850;
    wire n3853;
    wire n3856;
    wire n3859;
    wire n3862;
    wire n3865;
    wire n3868;
    wire n3871;
    wire n3874;
    wire n3877;
    wire n3881;
    wire n3884;
    wire n3887;
    wire n3890;
    wire n3893;
    wire n3896;
    wire n3899;
    wire n3901;
    wire n3904;
    wire n3907;
    wire n3910;
    wire n3913;
    wire n3916;
    wire n3919;
    wire n3922;
    wire n3925;
    wire n3928;
    wire n3931;
    wire n3934;
    wire n3937;
    wire n3940;
    wire n3943;
    wire n3946;
    wire n3949;
    wire n3952;
    wire n3955;
    wire n3958;
    wire n3961;
    wire n3964;
    wire n3967;
    wire n3970;
    wire n3973;
    wire n3976;
    wire n3979;
    wire n3982;
    wire n3985;
    wire n3988;
    wire n3991;
    wire n3994;
    wire n3998;
    wire n4001;
    wire n4004;
    wire n4007;
    wire n4010;
    wire n4013;
    wire n4016;
    wire n4018;
    wire n4021;
    wire n4024;
    wire n4027;
    wire n4030;
    wire n4033;
    wire n4036;
    wire n4039;
    wire n4042;
    wire n4045;
    wire n4048;
    wire n4051;
    wire n4054;
    wire n4057;
    wire n4060;
    wire n4063;
    wire n4066;
    wire n4069;
    wire n4072;
    wire n4075;
    wire n4078;
    wire n4081;
    wire n4084;
    wire n4087;
    wire n4090;
    wire n4093;
    wire n4096;
    wire n4100;
    wire n4103;
    wire n4105;
    wire n4108;
    wire n4111;
    wire n4114;
    wire n4117;
    wire n4120;
    wire n4123;
    wire n4126;
    wire n4129;
    wire n4132;
    wire n4135;
    wire n4138;
    wire n4141;
    wire n4144;
    wire n4147;
    wire n4150;
    wire n4153;
    wire n4156;
    wire n4159;
    wire n4162;
    wire n4165;
    wire n4168;
    wire n4171;
    wire n4174;
    wire n4177;
    wire n4180;
    wire n4183;
    wire n4186;
    wire n4189;
    wire n4192;
    wire n4195;
    wire n4198;
    wire n4201;
    wire n4204;
    wire n4207;
    wire n4210;
    wire n4213;
    wire n4216;
    wire n4219;
    wire n4222;
    wire n4225;
    wire n4228;
    wire n4231;
    wire n4234;
    wire n4237;
    wire n4240;
    wire n4243;
    wire n4246;
    wire n4249;
    wire n4252;
    wire n4255;
    wire n4258;
    wire n4261;
    wire n4264;
    wire n4267;
    wire n4271;
    wire n4274;
    wire n4277;
    wire n4280;
    wire n4283;
    wire n4286;
    wire n4289;
    wire n4291;
    wire n4294;
    wire n4297;
    wire n4300;
    wire n4303;
    wire n4306;
    wire n4309;
    wire n4312;
    wire n4315;
    wire n4318;
    wire n4321;
    wire n4324;
    wire n4327;
    wire n4330;
    wire n4333;
    wire n4336;
    wire n4339;
    wire n4342;
    wire n4345;
    wire n4348;
    wire n4351;
    wire n4354;
    wire n4357;
    wire n4360;
    wire n4363;
    wire n4366;
    wire n4369;
    wire n4373;
    wire n4376;
    wire n4378;
    wire n4381;
    wire n4384;
    wire n4387;
    wire n4390;
    wire n4393;
    wire n4396;
    wire n4399;
    wire n4402;
    wire n4405;
    wire n4408;
    wire n4411;
    wire n4414;
    wire n4417;
    wire n4420;
    wire n4423;
    wire n4426;
    wire n4429;
    wire n4432;
    wire n4435;
    wire n4438;
    wire n4441;
    wire n4444;
    wire n4447;
    wire n4450;
    wire n4453;
    wire n4456;
    wire n4459;
    wire n4462;
    wire n4465;
    wire n4468;
    wire n4471;
    wire n4474;
    wire n4477;
    wire n4480;
    wire n4483;
    wire n4486;
    wire n4489;
    wire n4492;
    wire n4495;
    wire n4498;
    wire n4501;
    wire n4504;
    wire n4507;
    wire n4510;
    wire n4513;
    wire n4516;
    wire n4519;
    wire n4522;
    wire n4525;
    wire n4528;
    wire n4531;
    wire n4534;
    wire n4537;
    wire n4540;
    wire n4543;
    wire n4546;
    wire n4549;
    wire n4552;
    wire n4555;
    wire n4558;
    wire n4561;
    wire n4564;
    wire n4567;
    wire n4570;
    wire n4573;
    wire n4576;
    wire n4579;
    wire n4582;
    wire n4585;
    wire n4588;
    wire n4591;
    wire n4594;
    wire n4597;
    wire n4600;
    wire n4603;
    wire n4606;
    wire n4609;
    wire n4612;
    wire n4615;
    wire n4618;
    wire n4621;
    wire n4624;
    wire n4627;
    wire n4630;
    wire n4633;
    wire n4636;
    wire n4639;
    wire n4642;
    wire n4645;
    wire n4648;
    wire n4651;
    wire n4654;
    wire n4657;
    wire n4660;
    wire n4663;
    wire n4666;
    wire n4669;
    wire n4672;
    wire n4675;
    wire n4678;
    wire n4681;
    wire n4684;
    wire n4687;
    wire n4690;
    wire n4693;
    wire n4696;
    wire n4699;
    wire n4702;
    wire n4705;
    wire n4708;
    wire n4711;
    wire n4714;
    wire n4717;
    wire n4720;
    wire n4723;
    wire n4726;
    wire n4729;
    wire n4732;
    wire n4735;
    wire n4738;
    wire n4741;
    wire n4744;
    wire n4747;
    wire n4750;
    wire n4753;
    wire n4756;
    wire n4759;
    wire n4762;
    wire n4765;
    wire n4768;
    wire n4771;
    wire n4774;
    wire n4777;
    wire n4780;
    wire n4783;
    wire n4786;
    wire n4789;
    wire n4792;
    wire n4795;
    wire n4798;
    wire n4801;
    wire n4804;
    wire n4807;
    wire n4810;
    wire n4813;
    wire n4816;
    wire n4819;
    wire n4822;
    wire n4825;
    wire n4828;
    wire n4831;
    wire n4834;
    wire n4837;
    wire n4840;
    wire n4843;
    wire n4846;
    wire n4849;
    wire n4852;
    wire n4855;
    wire n4858;
    wire n4861;
    wire n4864;
    wire n4867;
    wire n4870;
    wire n4873;
    wire n4876;
    wire n4879;
    wire n4882;
    wire n4885;
    wire n4888;
    wire n4891;
    wire n4894;
    wire n4897;
    wire n4900;
    wire n4903;
    wire n4906;
    wire n4909;
    wire n4912;
    wire n4915;
    wire n4918;
    wire n4921;
    wire n4924;
    wire n4927;
    wire n4930;
    wire n4933;
    wire n4936;
    wire n4939;
    wire n4942;
    wire n4945;
    wire n4948;
    wire n4951;
    wire n4954;
    wire n4957;
    wire n4960;
    wire n4963;
    wire n4969;
    wire n4972;
    wire n4975;
    wire n4978;
    wire n4981;
    wire n4984;
    wire n4987;
    wire n4990;
    wire n4993;
    wire n4996;
    wire n4999;
    wire n5002;
    wire n5008;
    wire n5011;
    wire n5014;
    wire n5017;
    wire n5020;
    wire n5026;
    jnot g000(.din(G76gat), .dout(n45));
    jand g001(.dinb(n45), .dina(n4786), .dout(n49));
    jnot g002(.din(G24gat), .dout(n52));
    jand g003(.dinb(n52), .dina(n4756), .dout(n56));
    jnot g004(.din(G11gat), .dout(n59));
    jand g005(.dinb(n59), .dina(n4717), .dout(n63));
    jor g006(.dinb(n56), .dina(n63), .dout(n67));
    jor g007(.dinb(n4762), .dina(n67), .dout(n71));
    jnot g008(.din(G37gat), .dout(n74));
    jand g009(.dinb(n74), .dina(n4666), .dout(n78));
    jnot g010(.din(G63gat), .dout(n81));
    jand g011(.dinb(n81), .dina(n4615), .dout(n85));
    jor g012(.dinb(n78), .dina(n85), .dout(n89));
    jnot g013(.din(G102gat), .dout(n92));
    jand g014(.dinb(n92), .dina(n4555), .dout(n96));
    jnot g015(.din(G50gat), .dout(n99));
    jand g016(.dinb(n99), .dina(n4495), .dout(n103));
    jor g017(.dinb(n96), .dina(n103), .dout(n107));
    jnot g018(.din(G89gat), .dout(n110));
    jand g019(.dinb(n110), .dina(n4861), .dout(n114));
    jnot g020(.din(G1gat), .dout(n117));
    jand g021(.dinb(n117), .dina(n4399), .dout(n121));
    jor g022(.dinb(n114), .dina(n121), .dout(n125));
    jor g023(.dinb(n107), .dina(n125), .dout(n129));
    jor g024(.dinb(n4376), .dina(n129), .dout(n133));
    jor g025(.dinb(n4373), .dina(n133), .dout(n137));
    jnot g026(.din(G112gat), .dout(n140));
    jnot g027(.din(n49), .dout(n143));
    jnot g028(.din(G30gat), .dout(n146));
    jor g029(.dinb(n4759), .dina(n146), .dout(n150));
    jnot g030(.din(G17gat), .dout(n153));
    jor g031(.dinb(n4753), .dina(n153), .dout(n157));
    jand g032(.dinb(n150), .dina(n157), .dout(n161));
    jand g033(.dinb(n143), .dina(n161), .dout(n165));
    jnot g034(.din(G43gat), .dout(n168));
    jor g035(.dinb(n4693), .dina(n168), .dout(n172));
    jnot g036(.din(G69gat), .dout(n175));
    jor g037(.dinb(n4651), .dina(n175), .dout(n179));
    jand g038(.dinb(n172), .dina(n179), .dout(n183));
    jnot g039(.din(G108gat), .dout(n186));
    jor g040(.dinb(n4591), .dina(n186), .dout(n190));
    jnot g041(.din(G56gat), .dout(n193));
    jor g042(.dinb(n4531), .dina(n193), .dout(n197));
    jand g043(.dinb(n190), .dina(n197), .dout(n201));
    jnot g044(.din(G95gat), .dout(n204));
    jor g045(.dinb(n4471), .dina(n204), .dout(n208));
    jnot g046(.din(G4gat), .dout(n211));
    jor g047(.dinb(n4435), .dina(n211), .dout(n215));
    jand g048(.dinb(n208), .dina(n215), .dout(n219));
    jand g049(.dinb(n201), .dina(n219), .dout(n223));
    jand g050(.dinb(n4103), .dina(n223), .dout(n227));
    jand g051(.dinb(n4100), .dina(n227), .dout(n231));
    jor g052(.dinb(n4558), .dina(n231), .dout(n235));
    jand g053(.dinb(n4534), .dina(n235), .dout(n239));
    jand g054(.dinb(n4289), .dina(n239), .dout(n243));
    jnot g055(.din(G8gat), .dout(n246));
    jor g056(.dinb(n4402), .dina(n231), .dout(n250));
    jand g057(.dinb(n4378), .dina(n250), .dout(n254));
    jand g058(.dinb(n4016), .dina(n254), .dout(n258));
    jor g059(.dinb(n243), .dina(n258), .dout(n262));
    jnot g060(.din(G99gat), .dout(n265));
    jor g061(.dinb(n4438), .dina(n231), .dout(n269));
    jand g062(.dinb(n4840), .dina(n269), .dout(n273));
    jand g063(.dinb(n3899), .dina(n273), .dout(n277));
    jnot g064(.din(G73gat), .dout(n280));
    jor g065(.dinb(n4618), .dina(n231), .dout(n284));
    jand g066(.dinb(n4594), .dina(n284), .dout(n288));
    jand g067(.dinb(n3815), .dina(n288), .dout(n292));
    jor g068(.dinb(n277), .dina(n292), .dout(n296));
    jor g069(.dinb(n262), .dina(n296), .dout(n300));
    jxor g070(.dinb(n4225), .dina(n231), .dout(n304));
    jor g071(.dinb(n4237), .dina(n304), .dout(n308));
    jor g072(.dinb(n3739), .dina(n308), .dout(n312));
    jnot g073(.din(n312), .dout(n315));
    jnot g074(.din(G60gat), .dout(n318));
    jor g075(.dinb(n4498), .dina(n231), .dout(n322));
    jand g076(.dinb(n4474), .dina(n322), .dout(n326));
    jand g077(.dinb(n3611), .dina(n326), .dout(n330));
    jxor g078(.dinb(n4654), .dina(n231), .dout(n334));
    jnot g079(.din(G47gat), .dout(n337));
    jand g080(.dinb(n4672), .dina(n337), .dout(n341));
    jand g081(.dinb(n334), .dina(n3538), .dout(n345));
    jor g082(.dinb(n330), .dina(n3536), .dout(n349));
    jnot g083(.din(G86gat), .dout(n352));
    jor g084(.dinb(n4789), .dina(n231), .dout(n356));
    jand g085(.dinb(n4765), .dina(n356), .dout(n360));
    jand g086(.dinb(n3431), .dina(n360), .dout(n364));
    jnot g087(.din(G21gat), .dout(n367));
    jor g088(.dinb(n4720), .dina(n231), .dout(n371));
    jand g089(.dinb(n4696), .dina(n371), .dout(n375));
    jand g090(.dinb(n3260), .dina(n375), .dout(n379));
    jor g091(.dinb(n364), .dina(n379), .dout(n383));
    jor g092(.dinb(n349), .dina(n383), .dout(n387));
    jor g093(.dinb(n3191), .dina(n387), .dout(n391));
    jor g094(.dinb(n3188), .dina(n391), .dout(n395));
    jand g095(.dinb(n4453), .dina(n137), .dout(n399));
    jor g096(.dinb(n4822), .dina(n399), .dout(n403));
    jand g097(.dinb(n3925), .dina(n395), .dout(n407));
    jor g098(.dinb(n4354), .dina(n407), .dout(n411));
    jor g099(.dinb(n4864), .dina(n411), .dout(n415));
    jnot g100(.din(n415), .dout(n418));
    jand g101(.dinb(n4513), .dina(n137), .dout(n422));
    jor g102(.dinb(n4123), .dina(n422), .dout(n426));
    jor g103(.dinb(n3652), .dina(n426), .dout(n430));
    jand g104(.dinb(n3154), .dina(n395), .dout(n434));
    jnot g105(.din(n434), .dout(n437));
    jnot g106(.din(G66gat), .dout(n440));
    jand g107(.dinb(n3092), .dina(n326), .dout(n444));
    jand g108(.dinb(n437), .dina(n3019), .dout(n448));
    jnot g109(.din(G79gat), .dout(n451));
    jand g110(.dinb(n4573), .dina(n137), .dout(n455));
    jor g111(.dinb(n4141), .dina(n455), .dout(n459));
    jor g112(.dinb(n4330), .dina(n459), .dout(n463));
    jand g113(.dinb(n4417), .dina(n137), .dout(n467));
    jor g114(.dinb(n4105), .dina(n467), .dout(n471));
    jor g115(.dinb(n4057), .dina(n471), .dout(n475));
    jand g116(.dinb(n463), .dina(n475), .dout(n479));
    jor g117(.dinb(n3901), .dina(n403), .dout(n483));
    jand g118(.dinb(n4633), .dina(n137), .dout(n487));
    jor g119(.dinb(n4159), .dina(n487), .dout(n491));
    jor g120(.dinb(n3856), .dina(n491), .dout(n495));
    jand g121(.dinb(n483), .dina(n495), .dout(n499));
    jand g122(.dinb(n479), .dina(n499), .dout(n503));
    jxor g123(.dinb(n4177), .dina(n231), .dout(n507));
    jnot g124(.din(n341), .dout(n510));
    jor g125(.dinb(n507), .dina(n2861), .dout(n514));
    jand g126(.dinb(n430), .dina(n2849), .dout(n518));
    jnot g127(.din(G82gat), .dout(n521));
    jand g128(.dinb(n4804), .dina(n137), .dout(n525));
    jor g129(.dinb(n2834), .dina(n525), .dout(n529));
    jor g130(.dinb(n3433), .dina(n529), .dout(n533));
    jand g131(.dinb(n4735), .dina(n137), .dout(n537));
    jor g132(.dinb(n4207), .dina(n537), .dout(n541));
    jor g133(.dinb(n3262), .dina(n541), .dout(n545));
    jand g134(.dinb(n533), .dina(n545), .dout(n549));
    jand g135(.dinb(n518), .dina(n549), .dout(n553));
    jand g136(.dinb(n3676), .dina(n553), .dout(n557));
    jand g137(.dinb(n2780), .dina(n557), .dout(n561));
    jor g138(.dinb(n3781), .dina(n561), .dout(n565));
    jand g139(.dinb(n3763), .dina(n565), .dout(n569));
    jand g140(.dinb(n2972), .dina(n569), .dout(n573));
    jor g141(.dinb(n448), .dina(n573), .dout(n577));
    jor g142(.dinb(n418), .dina(n577), .dout(n581));
    jand g143(.dinb(n2836), .dina(n395), .dout(n585));
    jnot g144(.din(n585), .dout(n588));
    jnot g145(.din(G53gat), .dout(n591));
    jand g146(.dinb(n4669), .dina(n591), .dout(n595));
    jand g147(.dinb(n334), .dina(n2642), .dout(n599));
    jand g148(.dinb(n588), .dina(n2608), .dout(n603));
    jor g149(.dinb(n3226), .dina(n561), .dout(n607));
    jand g150(.dinb(n3193), .dina(n607), .dout(n611));
    jnot g151(.din(G27gat), .dout(n614));
    jor g152(.dinb(n3325), .dina(n395), .dout(n618));
    jand g153(.dinb(n2546), .dina(n618), .dout(n622));
    jand g154(.dinb(n611), .dina(n622), .dout(n626));
    jor g155(.dinb(n603), .dina(n626), .dout(n630));
    jor g156(.dinb(n3397), .dina(n561), .dout(n634));
    jand g157(.dinb(n3364), .dina(n634), .dout(n638));
    jnot g158(.din(G92gat), .dout(n641));
    jor g159(.dinb(n3496), .dina(n395), .dout(n645));
    jand g160(.dinb(n2369), .dina(n645), .dout(n649));
    jand g161(.dinb(n638), .dina(n649), .dout(n653));
    jnot g162(.din(G14gat), .dout(n656));
    jor g163(.dinb(n3982), .dina(n561), .dout(n660));
    jand g164(.dinb(n3964), .dina(n660), .dout(n664));
    jand g165(.dinb(n2207), .dina(n664), .dout(n668));
    jor g166(.dinb(n653), .dina(n668), .dout(n672));
    jnot g167(.din(G34gat), .dout(n675));
    jor g168(.dinb(n2165), .dina(n561), .dout(n679));
    jnot g169(.din(G40gat), .dout(n682));
    jnot g170(.din(n308), .dout(n685));
    jand g171(.dinb(n2069), .dina(n685), .dout(n689));
    jand g172(.dinb(n679), .dina(n2002), .dout(n693));
    jnot g173(.din(G115gat), .dout(n696));
    jor g174(.dinb(n4255), .dina(n561), .dout(n700));
    jand g175(.dinb(n4081), .dina(n700), .dout(n704));
    jand g176(.dinb(n1955), .dina(n704), .dout(n708));
    jor g177(.dinb(n1880), .dina(n708), .dout(n712));
    jor g178(.dinb(n672), .dina(n712), .dout(n716));
    jor g179(.dinb(n1877), .dina(n716), .dout(n720));
    jor g180(.dinb(n1874), .dina(n720), .dout(n724));
    jand g181(.dinb(n4018), .dina(n395), .dout(n728));
    jor g182(.dinb(n2881), .dina(n728), .dout(n732));
    jand g183(.dinb(n2254), .dina(n724), .dout(n736));
    jor g184(.dinb(n1750), .dina(n736), .dout(n740));
    jnot g185(.din(n444), .dout(n743));
    jor g186(.dinb(n434), .dina(n1799), .dout(n747));
    jand g187(.dinb(n3817), .dina(n395), .dout(n751));
    jor g188(.dinb(n2863), .dina(n751), .dout(n755));
    jor g189(.dinb(n2974), .dina(n755), .dout(n759));
    jand g190(.dinb(n1787), .dina(n759), .dout(n763));
    jand g191(.dinb(n3184), .dina(n763), .dout(n767));
    jnot g192(.din(n599), .dout(n770));
    jor g193(.dinb(n585), .dina(n1784), .dout(n774));
    jand g194(.dinb(n3286), .dina(n395), .dout(n778));
    jor g195(.dinb(n2782), .dina(n778), .dout(n782));
    jand g196(.dinb(n3211), .dina(n561), .dout(n786));
    jor g197(.dinb(n2548), .dina(n786), .dout(n790));
    jor g198(.dinb(n782), .dina(n790), .dout(n794));
    jand g199(.dinb(n1769), .dina(n794), .dout(n798));
    jand g200(.dinb(n3457), .dina(n395), .dout(n802));
    jor g201(.dinb(n2800), .dina(n802), .dout(n806));
    jand g202(.dinb(n3382), .dina(n561), .dout(n810));
    jor g203(.dinb(n2431), .dina(n810), .dout(n814));
    jor g204(.dinb(n806), .dina(n814), .dout(n818));
    jor g205(.dinb(n2209), .dina(n732), .dout(n822));
    jand g206(.dinb(n818), .dina(n822), .dout(n826));
    jand g207(.dinb(n3700), .dina(n395), .dout(n830));
    jnot g208(.din(n689), .dout(n833));
    jor g209(.dinb(n830), .dina(n1748), .dout(n837));
    jand g210(.dinb(n4291), .dina(n395), .dout(n841));
    jor g211(.dinb(n2899), .dina(n841), .dout(n845));
    jor g212(.dinb(n1957), .dina(n845), .dout(n849));
    jand g213(.dinb(n1739), .dina(n849), .dout(n853));
    jand g214(.dinb(n826), .dina(n853), .dout(n857));
    jand g215(.dinb(n1736), .dina(n857), .dout(n861));
    jand g216(.dinb(n1733), .dina(n861), .dout(n865));
    jor g217(.dinb(n3037), .dina(n865), .dout(n869));
    jand g218(.dinb(n3613), .dina(n395), .dout(n873));
    jor g219(.dinb(n3166), .dina(n873), .dout(n877));
    jnot g220(.din(n877), .dout(n880));
    jand g221(.dinb(n869), .dina(n1595), .dout(n884));
    jor g222(.dinb(n2644), .dina(n865), .dout(n888));
    jand g223(.dinb(n3553), .dina(n395), .dout(n892));
    jand g224(.dinb(n4675), .dina(n137), .dout(n896));
    jor g225(.dinb(n4189), .dina(n896), .dout(n900));
    jor g226(.dinb(n892), .dina(n1871), .dout(n904));
    jnot g227(.din(n904), .dout(n907));
    jand g228(.dinb(n888), .dina(n1637), .dout(n911));
    jor g229(.dinb(n884), .dina(n911), .dout(n915));
    jor g230(.dinb(n2491), .dina(n865), .dout(n919));
    jand g231(.dinb(n2590), .dina(n919), .dout(n923));
    jor g232(.dinb(n2014), .dina(n865), .dout(n927));
    jor g233(.dinb(n830), .dina(n3682), .dout(n931));
    jnot g234(.din(n931), .dout(n934));
    jand g235(.dinb(n927), .dina(n1616), .dout(n938));
    jor g236(.dinb(n923), .dina(n938), .dout(n942));
    jor g237(.dinb(n915), .dina(n942), .dout(n946));
    jor g238(.dinb(n2314), .dina(n865), .dout(n950));
    jand g239(.dinb(n2473), .dina(n950), .dout(n954));
    jor g240(.dinb(n1900), .dina(n865), .dout(n958));
    jand g241(.dinb(n1882), .dina(n958), .dout(n962));
    jor g242(.dinb(n954), .dina(n962), .dout(n966));
    jnot g243(.din(n411), .dout(n969));
    jnot g244(.din(G105gat), .dout(n972));
    jor g245(.dinb(n1730), .dina(n865), .dout(n976));
    jand g246(.dinb(n1673), .dina(n976), .dout(n980));
    jor g247(.dinb(n2917), .dina(n865), .dout(n984));
    jand g248(.dinb(n2761), .dina(n984), .dout(n988));
    jor g249(.dinb(n980), .dina(n988), .dout(n992));
    jor g250(.dinb(n966), .dina(n992), .dout(n996));
    jor g251(.dinb(n946), .dina(n996), .dout(n1000));
    jand g252(.dinb(n1580), .dina(n1000), .dout(G421gat));
    jand g253(.dinb(n3094), .dina(n724), .dout(n1008));
    jor g254(.dinb(n1008), .dina(n1642), .dout(n1012));
    jand g255(.dinb(n2701), .dina(n724), .dout(n1016));
    jor g256(.dinb(n1016), .dina(n1837), .dout(n1020));
    jand g257(.dinb(n1012), .dina(n1020), .dout(n1024));
    jand g258(.dinb(n1024), .dina(n1618), .dout(n1028));
    jand g259(.dinb(n2071), .dina(n724), .dout(n1032));
    jor g260(.dinb(n1032), .dina(n1801), .dout(n1036));
    jand g261(.dinb(n1036), .dina(n988), .dout(n1040));
    jand g262(.dinb(n1024), .dina(n1040), .dout(n1044));
    jor g263(.dinb(n1600), .dina(n1044), .dout(n1048));
    jor g264(.dinb(n1598), .dina(n1048), .dout(G431gat));
    jand g265(.dinb(n2371), .dina(n724), .dout(n1056));
    jor g266(.dinb(n1819), .dina(n1056), .dout(n1060));
    jand g267(.dinb(n1020), .dina(n1060), .dout(n1064));
    jand g268(.dinb(n1036), .dina(n980), .dout(n1068));
    jand g269(.dinb(n1064), .dina(n1068), .dout(n1072));
    jand g270(.dinb(n911), .dina(n1036), .dout(n1076));
    jor g271(.dinb(n1639), .dina(n1076), .dout(n1080));
    jor g272(.dinb(n1044), .dina(n1080), .dout(n1084));
    jor g273(.dinb(n1622), .dina(n1084), .dout(G432gat));
    jdff dff_A_9J82KA3Q7_0(.din(n5026), .dout(G430gat));
    jdff dff_A_RCUy6P1j0_1(.din(n946), .dout(n5026));
    jdff dff_A_vrpEtuVb5_0(.din(n5020), .dout(G370gat));
    jdff dff_A_ZswGhIHK6_0(.din(n5017), .dout(n5020));
    jdff dff_A_wAmORMbX5_0(.din(n5014), .dout(n5017));
    jdff dff_A_FiOshWDZ9_0(.din(n5011), .dout(n5014));
    jdff dff_A_KJlCgD6r5_0(.din(n5008), .dout(n5011));
    jdff dff_A_cgYnHa567_1(.din(n724), .dout(n5008));
    jdff dff_A_zl0zYyGv5_0(.din(n5002), .dout(G329gat));
    jdff dff_A_ALrhgiIh9_0(.din(n4999), .dout(n5002));
    jdff dff_A_4ZYY7OJs4_0(.din(n4996), .dout(n4999));
    jdff dff_A_CfF1bmPV9_0(.din(n4993), .dout(n4996));
    jdff dff_A_FJfEB19U4_0(.din(n4990), .dout(n4993));
    jdff dff_A_QsnA1HsA9_0(.din(n4987), .dout(n4990));
    jdff dff_A_0k8GlC1P6_0(.din(n4984), .dout(n4987));
    jdff dff_A_w4Gaq2Dg0_0(.din(n4981), .dout(n4984));
    jdff dff_A_BWbWi0ka0_0(.din(n4978), .dout(n4981));
    jdff dff_A_qQXOIv9C2_0(.din(n4975), .dout(n4978));
    jdff dff_A_4ifcTakD8_0(.din(n4972), .dout(n4975));
    jdff dff_A_Gw6NYGQ52_0(.din(n4969), .dout(n4972));
    jdff dff_A_R3l9X8Gn8_1(.din(n395), .dout(n4969));
    jdff dff_A_GlggAXEA0_0(.din(n4963), .dout(G223gat));
    jdff dff_A_cjO7Z7sD3_0(.din(n4960), .dout(n4963));
    jdff dff_A_B9DHgZ8K7_0(.din(n4957), .dout(n4960));
    jdff dff_A_okGHrDh63_0(.din(n4954), .dout(n4957));
    jdff dff_A_sgcmtF7V4_0(.din(n4951), .dout(n4954));
    jdff dff_A_CKJaqjPo3_0(.din(n4948), .dout(n4951));
    jdff dff_A_51UUfiLp3_0(.din(n4945), .dout(n4948));
    jdff dff_A_VWaVx4QM1_0(.din(n4942), .dout(n4945));
    jdff dff_A_7RCADPY52_0(.din(n4939), .dout(n4942));
    jdff dff_A_h0b9DVmg1_0(.din(n4936), .dout(n4939));
    jdff dff_A_iTGutd682_0(.din(n4933), .dout(n4936));
    jdff dff_A_Z928laBU1_0(.din(n4930), .dout(n4933));
    jdff dff_A_auaaU9JO5_0(.din(n4927), .dout(n4930));
    jdff dff_A_G2P8yfdL6_0(.din(n4924), .dout(n4927));
    jdff dff_A_NAzGTNyg9_0(.din(n4921), .dout(n4924));
    jdff dff_A_uL6REXsy7_0(.din(n4918), .dout(n4921));
    jdff dff_A_QWADezyW3_0(.din(n4915), .dout(n4918));
    jdff dff_A_RxCxpIGD6_0(.din(n4912), .dout(n4915));
    jdff dff_A_4a1iUSTY4_0(.din(n4909), .dout(n4912));
    jdff dff_A_MaxiYCp89_2(.din(n137), .dout(n4909));
    jdff dff_A_PYJI8UMC6_1(.din(G105gat), .dout(n4906));
    jdff dff_A_wxwzoTvF1_1(.din(n4906), .dout(n4903));
    jdff dff_A_2gHoIhD52_1(.din(n4903), .dout(n4900));
    jdff dff_A_0Re8soi95_1(.din(n4900), .dout(n4897));
    jdff dff_A_KdNP7kkJ2_1(.din(n4897), .dout(n4894));
    jdff dff_A_lxZPLhBu6_1(.din(n4894), .dout(n4891));
    jdff dff_A_R2AnmVBV4_1(.din(n4891), .dout(n4888));
    jdff dff_A_y6qefsw96_1(.din(n4888), .dout(n4885));
    jdff dff_A_fDZDKLkV4_1(.din(n4885), .dout(n4882));
    jdff dff_A_5HP8BIJ01_1(.din(n4882), .dout(n4879));
    jdff dff_A_B6clcUBo2_1(.din(n4879), .dout(n4876));
    jdff dff_A_rIMszMo84_1(.din(n4876), .dout(n4873));
    jdff dff_A_HMT7AyUD1_1(.din(n4873), .dout(n4870));
    jdff dff_A_YC0wFypt7_1(.din(n4870), .dout(n4867));
    jdff dff_A_tkBIfQCV9_1(.din(n4867), .dout(n4864));
    jdff dff_A_AcISA6RU7_2(.din(G95gat), .dout(n4861));
    jdff dff_A_F2J5LdON6_0(.din(G95gat), .dout(n4858));
    jdff dff_A_nGIOe9D07_0(.din(n4858), .dout(n4855));
    jdff dff_A_j00AEJWg8_0(.din(n4855), .dout(n4852));
    jdff dff_A_I6MPMl0M1_0(.din(n4852), .dout(n4849));
    jdff dff_A_pN3ggmc15_0(.din(n4849), .dout(n4846));
    jdff dff_A_retoFnjf2_0(.din(n4846), .dout(n4843));
    jdff dff_A_gp6QfW5O2_0(.din(n4843), .dout(n4840));
    jdff dff_A_st7JVpjz6_0(.din(n204), .dout(n4837));
    jdff dff_A_g0XFfzZl5_0(.din(n4837), .dout(n4834));
    jdff dff_A_E9ik2gEm3_0(.din(n4834), .dout(n4831));
    jdff dff_A_jdyjcmOa7_0(.din(n4831), .dout(n4828));
    jdff dff_A_Vr9TnkqD2_0(.din(n4828), .dout(n4825));
    jdff dff_A_PUZJsGRG5_0(.din(n4825), .dout(n4822));
    jdff dff_A_Z8LXqTPZ1_0(.din(G76gat), .dout(n4819));
    jdff dff_A_3N6aZG4V1_0(.din(n4819), .dout(n4816));
    jdff dff_A_RgKDmBCP5_0(.din(n4816), .dout(n4813));
    jdff dff_A_JODcJSlN7_0(.din(n4813), .dout(n4810));
    jdff dff_A_WsAkDPUO5_0(.din(n4810), .dout(n4807));
    jdff dff_A_kmbyvGTf0_0(.din(n4807), .dout(n4804));
    jdff dff_A_1S6iYLtK3_0(.din(n45), .dout(n4801));
    jdff dff_A_58tyhiZ74_0(.din(n4801), .dout(n4798));
    jdff dff_A_9aYZ00BV6_0(.din(n4798), .dout(n4795));
    jdff dff_A_lmUF8aNa7_0(.din(n4795), .dout(n4792));
    jdff dff_A_a5LUy0Jh0_0(.din(n4792), .dout(n4789));
    jdff dff_A_iYOw4pOk9_2(.din(G82gat), .dout(n4786));
    jdff dff_A_7hgsGo9G1_1(.din(G82gat), .dout(n4783));
    jdff dff_A_YrRtR3Ve0_1(.din(n4783), .dout(n4780));
    jdff dff_A_rZNTymzR4_1(.din(n4780), .dout(n4777));
    jdff dff_A_RTUJgqj54_1(.din(n4777), .dout(n4774));
    jdff dff_A_y1wdbJ7V5_1(.din(n4774), .dout(n4771));
    jdff dff_A_JHlZvLiu2_1(.din(n4771), .dout(n4768));
    jdff dff_A_G8whc0Pr5_1(.din(n4768), .dout(n4765));
    jdff dff_A_DMrYvpqC1_1(.din(n49), .dout(n4762));
    jdff dff_A_8fNpvyNO4_0(.din(G24gat), .dout(n4759));
    jdff dff_A_vq767C681_1(.din(G30gat), .dout(n4756));
    jdff dff_A_scHdCel47_1(.din(G11gat), .dout(n4753));
    jdff dff_A_MQd5T3JC6_0(.din(G11gat), .dout(n4750));
    jdff dff_A_mtSJ8G1E7_0(.din(n4750), .dout(n4747));
    jdff dff_A_ZFI4vkSL7_0(.din(n4747), .dout(n4744));
    jdff dff_A_s83XpgJt9_0(.din(n4744), .dout(n4741));
    jdff dff_A_YqfOQ8zT2_0(.din(n4741), .dout(n4738));
    jdff dff_A_n9yPRBbA0_0(.din(n4738), .dout(n4735));
    jdff dff_A_jrm4zwtG2_0(.din(n59), .dout(n4732));
    jdff dff_A_PSEeBRYd0_0(.din(n4732), .dout(n4729));
    jdff dff_A_thtnU7wY1_0(.din(n4729), .dout(n4726));
    jdff dff_A_KRiWLSeP7_0(.din(n4726), .dout(n4723));
    jdff dff_A_cjWThgh89_0(.din(n4723), .dout(n4720));
    jdff dff_A_eny0RcZF5_2(.din(G17gat), .dout(n4717));
    jdff dff_A_xXeOIwou4_0(.din(G17gat), .dout(n4714));
    jdff dff_A_IAVnKPJE6_0(.din(n4714), .dout(n4711));
    jdff dff_A_nAqjQpYU9_0(.din(n4711), .dout(n4708));
    jdff dff_A_yjFjDUBe5_0(.din(n4708), .dout(n4705));
    jdff dff_A_RUCOTxEn2_0(.din(n4705), .dout(n4702));
    jdff dff_A_KSeK94Xh3_0(.din(n4702), .dout(n4699));
    jdff dff_A_DbMQvbvi3_0(.din(n4699), .dout(n4696));
    jdff dff_A_iK9sgUV75_1(.din(G37gat), .dout(n4693));
    jdff dff_A_N4JjRjiX8_0(.din(G37gat), .dout(n4690));
    jdff dff_A_baAoJW3O6_0(.din(n4690), .dout(n4687));
    jdff dff_A_9KzMed2U8_0(.din(n4687), .dout(n4684));
    jdff dff_A_msD5FqKo8_0(.din(n4684), .dout(n4681));
    jdff dff_A_vKMgwbGJ8_0(.din(n4681), .dout(n4678));
    jdff dff_A_rMRatPpU3_0(.din(n4678), .dout(n4675));
    jdff dff_A_Pjmk4a686_2(.din(G43gat), .dout(n4672));
    jdff dff_A_xghP78uJ2_1(.din(G43gat), .dout(n4669));
    jdff dff_A_wAnMmerE8_1(.din(G43gat), .dout(n4666));
    jdff dff_A_3ykacEbC4_0(.din(n78), .dout(n4663));
    jdff dff_A_9EIHA2mN8_0(.din(n4663), .dout(n4660));
    jdff dff_A_kxm4TQ1o1_0(.din(n4660), .dout(n4657));
    jdff dff_A_9XmdiHfa7_0(.din(n4657), .dout(n4654));
    jdff dff_A_U0O983TN1_1(.din(G63gat), .dout(n4651));
    jdff dff_A_HZbKt9s03_0(.din(G63gat), .dout(n4648));
    jdff dff_A_IO7KywT24_0(.din(n4648), .dout(n4645));
    jdff dff_A_VMN1DwnB5_0(.din(n4645), .dout(n4642));
    jdff dff_A_zy3GkgzL0_0(.din(n4642), .dout(n4639));
    jdff dff_A_38LifaDN7_0(.din(n4639), .dout(n4636));
    jdff dff_A_cOVi5QN32_0(.din(n4636), .dout(n4633));
    jdff dff_A_QQxypFdR7_0(.din(n81), .dout(n4630));
    jdff dff_A_8un81v9g3_0(.din(n4630), .dout(n4627));
    jdff dff_A_7HGOLgLQ0_0(.din(n4627), .dout(n4624));
    jdff dff_A_iqYffsIx4_0(.din(n4624), .dout(n4621));
    jdff dff_A_BWUVzlYy0_0(.din(n4621), .dout(n4618));
    jdff dff_A_4g578riZ3_2(.din(G69gat), .dout(n4615));
    jdff dff_A_Ge8B9hJt4_0(.din(G69gat), .dout(n4612));
    jdff dff_A_dvRx08Gc4_0(.din(n4612), .dout(n4609));
    jdff dff_A_isRDBUU88_0(.din(n4609), .dout(n4606));
    jdff dff_A_zK5BxrtN3_0(.din(n4606), .dout(n4603));
    jdff dff_A_5EXQ7Kn36_0(.din(n4603), .dout(n4600));
    jdff dff_B_95uf8pzk0_1(.din(n740), .dout(n1574));
    jdff dff_B_letGXm1p6_1(.din(n1574), .dout(n1577));
    jdff dff_B_TBCYFE2o0_1(.din(n1577), .dout(n1580));
    jdff dff_B_pTm7TwKv4_0(.din(n880), .dout(n1583));
    jdff dff_B_ZFViDVo62_0(.din(n1583), .dout(n1586));
    jdff dff_B_M4uKZ33d6_0(.din(n1586), .dout(n1589));
    jdff dff_B_BzQbd4wn1_0(.din(n1589), .dout(n1592));
    jdff dff_B_2aQgTpKd8_0(.din(n1592), .dout(n1595));
    jdff dff_B_zqiK0Xpw6_1(.din(n1028), .dout(n1598));
    jdff dff_A_ap4p4pgH8_0(.din(n942), .dout(n1600));
    jdff dff_B_Zb5l6RDP0_0(.din(n934), .dout(n1604));
    jdff dff_B_XihP7rBk7_0(.din(n1604), .dout(n1607));
    jdff dff_B_tm2ksOGf1_0(.din(n1607), .dout(n1610));
    jdff dff_B_mKHebEnU9_0(.din(n1610), .dout(n1613));
    jdff dff_B_TNL17A3L5_0(.din(n1613), .dout(n1616));
    jdff dff_A_bhTq7Q2L7_0(.din(n954), .dout(n1618));
    jdff dff_B_RIYvRidS5_1(.din(n1072), .dout(n1622));
    jdff dff_B_LSjvtylg8_0(.din(n907), .dout(n1625));
    jdff dff_B_MqE7YZoz4_0(.din(n1625), .dout(n1628));
    jdff dff_B_ZTCuf4J51_0(.din(n1628), .dout(n1631));
    jdff dff_B_KlpllYaD6_0(.din(n1631), .dout(n1634));
    jdff dff_B_DkoggYqW3_0(.din(n1634), .dout(n1637));
    jdff dff_A_lUbJeBKw1_0(.din(n923), .dout(n1639));
    jdff dff_A_Ht0QTSse1_0(.din(n1645), .dout(n1642));
    jdff dff_A_qS4YkDag0_0(.din(n1648), .dout(n1645));
    jdff dff_A_DxhtPWx42_0(.din(n1651), .dout(n1648));
    jdff dff_A_Y6V6tujw5_0(.din(n1654), .dout(n1651));
    jdff dff_A_YbFHvBUL5_0(.din(n1657), .dout(n1654));
    jdff dff_A_ww5EVM0P1_0(.din(n877), .dout(n1657));
    jdff dff_B_61851nHU8_1(.din(n969), .dout(n1661));
    jdff dff_B_Vy3M2GSb4_1(.din(n1661), .dout(n1664));
    jdff dff_B_lsmVxR8I6_1(.din(n1664), .dout(n1667));
    jdff dff_B_OGRnpnlf3_1(.din(n1667), .dout(n1670));
    jdff dff_B_IOwF4Glq7_1(.din(n1670), .dout(n1673));
    jdff dff_B_63lnhOn55_1(.din(n972), .dout(n1676));
    jdff dff_B_sMrOjCU75_1(.din(n1676), .dout(n1679));
    jdff dff_B_sFDJB6s57_1(.din(n1679), .dout(n1682));
    jdff dff_B_ZAn4Sgqp9_1(.din(n1682), .dout(n1685));
    jdff dff_B_P06ILHvw6_1(.din(n1685), .dout(n1688));
    jdff dff_B_zZX3Faph4_1(.din(n1688), .dout(n1691));
    jdff dff_B_XaagROtF9_1(.din(n1691), .dout(n1694));
    jdff dff_B_QEnaAqci1_1(.din(n1694), .dout(n1697));
    jdff dff_B_EYcpcktT1_1(.din(n1697), .dout(n1700));
    jdff dff_B_s5oZxAZy6_1(.din(n1700), .dout(n1703));
    jdff dff_B_Y3tVv5mi2_1(.din(n1703), .dout(n1706));
    jdff dff_B_4EwAZuwG0_1(.din(n1706), .dout(n1709));
    jdff dff_B_bPVohXzw7_1(.din(n1709), .dout(n1712));
    jdff dff_B_XMUnQGRf5_1(.din(n1712), .dout(n1715));
    jdff dff_B_XvNhl9Hs3_1(.din(n1715), .dout(n1718));
    jdff dff_B_87glUefm9_1(.din(n1718), .dout(n1721));
    jdff dff_B_l5MATZEJ2_1(.din(n1721), .dout(n1724));
    jdff dff_B_vCzdesii0_1(.din(n1724), .dout(n1727));
    jdff dff_B_jfxZeJNT7_1(.din(n1727), .dout(n1730));
    jdff dff_B_erZJyVKo4_1(.din(n767), .dout(n1733));
    jdff dff_B_RwErxWos9_1(.din(n798), .dout(n1736));
    jdff dff_B_eADzKhT00_1(.din(n837), .dout(n1739));
    jdff dff_B_zDm1Bszp8_0(.din(n833), .dout(n1742));
    jdff dff_B_yx1vB4yl4_0(.din(n1742), .dout(n1745));
    jdff dff_B_Gh5mMvPZ6_0(.din(n1745), .dout(n1748));
    jdff dff_A_YvsfF6k72_1(.din(n1753), .dout(n1750));
    jdff dff_A_yqcP8mIO8_1(.din(n1756), .dout(n1753));
    jdff dff_A_p4YkqInR2_1(.din(n1759), .dout(n1756));
    jdff dff_A_wfABZNCu4_1(.din(n1762), .dout(n1759));
    jdff dff_A_nu4IWkEs7_1(.din(n1765), .dout(n1762));
    jdff dff_A_ZkBAqm027_1(.din(n732), .dout(n1765));
    jdff dff_B_Vhe6vJ0b1_1(.din(n774), .dout(n1769));
    jdff dff_B_tXGSSCjs9_0(.din(n770), .dout(n1772));
    jdff dff_B_V4QtIwkQ2_0(.din(n1772), .dout(n1775));
    jdff dff_B_rnzU1YTc2_0(.din(n1775), .dout(n1778));
    jdff dff_B_wszG0AMj8_0(.din(n1778), .dout(n1781));
    jdff dff_B_sJNE8zIO8_0(.din(n1781), .dout(n1784));
    jdff dff_B_a1rqcxTg0_1(.din(n747), .dout(n1787));
    jdff dff_B_qUUUr8lb5_0(.din(n743), .dout(n1790));
    jdff dff_B_maInDkaC0_0(.din(n1790), .dout(n1793));
    jdff dff_B_39ayU2Sl8_0(.din(n1793), .dout(n1796));
    jdff dff_B_iR4wkDcl9_0(.din(n1796), .dout(n1799));
    jdff dff_A_3WSsRxUf9_0(.din(n1804), .dout(n1801));
    jdff dff_A_se6up4Ss9_0(.din(n1807), .dout(n1804));
    jdff dff_A_cHk6rDJq0_0(.din(n1810), .dout(n1807));
    jdff dff_A_jCNboXfa1_0(.din(n1813), .dout(n1810));
    jdff dff_A_IMLsThk60_0(.din(n1816), .dout(n1813));
    jdff dff_A_GzvYsrTd6_0(.din(n931), .dout(n1816));
    jdff dff_A_SKKqbJ652_0(.din(n1822), .dout(n1819));
    jdff dff_A_8zBGWutK1_0(.din(n1825), .dout(n1822));
    jdff dff_A_jT2p71gI7_0(.din(n1828), .dout(n1825));
    jdff dff_A_SXoqwkCD7_0(.din(n1831), .dout(n1828));
    jdff dff_A_k33Srw5y6_0(.din(n1834), .dout(n1831));
    jdff dff_A_kM1VUIek2_0(.din(n806), .dout(n1834));
    jdff dff_A_eb3iF4Np2_0(.din(n1840), .dout(n1837));
    jdff dff_A_nC1hyU7V1_0(.din(n1843), .dout(n1840));
    jdff dff_A_Ux3zMEJf2_0(.din(n1846), .dout(n1843));
    jdff dff_A_BJy6mq5s7_0(.din(n1849), .dout(n1846));
    jdff dff_A_q8Bkd44h3_0(.din(n1852), .dout(n1849));
    jdff dff_A_tVDtwLTa1_0(.din(n904), .dout(n1852));
    jdff dff_B_akSLQiSm2_0(.din(n900), .dout(n1856));
    jdff dff_B_LBaWGVAn0_0(.din(n1856), .dout(n1859));
    jdff dff_B_5AGmBoIP4_0(.din(n1859), .dout(n1862));
    jdff dff_B_kauUpNH26_0(.din(n1862), .dout(n1865));
    jdff dff_B_Cje7cwRF8_0(.din(n1865), .dout(n1868));
    jdff dff_B_uXF6yqlK1_0(.din(n1868), .dout(n1871));
    jdff dff_B_moVH5SBR5_1(.din(n581), .dout(n1874));
    jdff dff_B_0pCmD9204_1(.din(n630), .dout(n1877));
    jdff dff_B_WWvHWYd57_1(.din(n693), .dout(n1880));
    jdff dff_A_ux7bgzkJ7_0(.din(n1885), .dout(n1882));
    jdff dff_A_IPNqJfBU6_0(.din(n1888), .dout(n1885));
    jdff dff_A_KxMR96IR3_0(.din(n1891), .dout(n1888));
    jdff dff_A_cNOtW5Mx9_0(.din(n1894), .dout(n1891));
    jdff dff_A_qOv4CHeU1_0(.din(n1897), .dout(n1894));
    jdff dff_A_6c6mhX8v0_0(.din(n704), .dout(n1897));
    jdff dff_A_fDii76br6_0(.din(n1903), .dout(n1900));
    jdff dff_A_zpHB0f9z4_0(.din(n1906), .dout(n1903));
    jdff dff_A_llTFJ1Qm0_0(.din(n1909), .dout(n1906));
    jdff dff_A_ybiPwF451_0(.din(n1912), .dout(n1909));
    jdff dff_A_UrpyTP039_0(.din(n1955), .dout(n1912));
    jdff dff_B_T3Is5w2W2_2(.din(n696), .dout(n1916));
    jdff dff_B_pKTwd5Z91_2(.din(n1916), .dout(n1919));
    jdff dff_B_CqtvmWDt2_2(.din(n1919), .dout(n1922));
    jdff dff_B_08764Txh0_2(.din(n1922), .dout(n1925));
    jdff dff_B_pXtP3Vtx6_2(.din(n1925), .dout(n1928));
    jdff dff_B_eKkeObvC3_2(.din(n1928), .dout(n1931));
    jdff dff_B_OJgdGmN87_2(.din(n1931), .dout(n1934));
    jdff dff_B_pSVPQ7HT1_2(.din(n1934), .dout(n1937));
    jdff dff_B_t92uup1W4_2(.din(n1937), .dout(n1940));
    jdff dff_B_vlqbdS308_2(.din(n1940), .dout(n1943));
    jdff dff_B_jnVQKEtB0_2(.din(n1943), .dout(n1946));
    jdff dff_B_6aDjtOHo2_2(.din(n1946), .dout(n1949));
    jdff dff_B_12btdkct8_2(.din(n1949), .dout(n1952));
    jdff dff_B_gbWZni8G5_2(.din(n1952), .dout(n1955));
    jdff dff_A_Grp4gKbN7_0(.din(n1960), .dout(n1957));
    jdff dff_A_ITG7dhPe3_0(.din(n1963), .dout(n1960));
    jdff dff_A_rOAgBkxG5_0(.din(n1966), .dout(n1963));
    jdff dff_A_e8bdT4yK3_0(.din(n1969), .dout(n1966));
    jdff dff_A_SDe99cyn0_0(.din(n1972), .dout(n1969));
    jdff dff_A_e8PApaLy4_0(.din(n1975), .dout(n1972));
    jdff dff_A_KHl453nB9_0(.din(n1978), .dout(n1975));
    jdff dff_A_Jz1BAu5o4_0(.din(n1981), .dout(n1978));
    jdff dff_A_W99BY7sm6_0(.din(n1984), .dout(n1981));
    jdff dff_A_8UNSU2Zm8_0(.din(n1987), .dout(n1984));
    jdff dff_A_vo7ecOzY8_0(.din(n1990), .dout(n1987));
    jdff dff_A_cNYE0Rxi5_0(.din(n1993), .dout(n1990));
    jdff dff_A_oM79tBM66_0(.din(n1996), .dout(n1993));
    jdff dff_A_JO4lQiNv4_0(.din(n1999), .dout(n1996));
    jdff dff_A_AvwkGZtH5_0(.din(G115gat), .dout(n1999));
    jdff dff_A_9KkDxQ5a3_1(.din(n2005), .dout(n2002));
    jdff dff_A_d8smjoO24_1(.din(n2008), .dout(n2005));
    jdff dff_A_iYCqwx7Q1_1(.din(n2011), .dout(n2008));
    jdff dff_A_LmDCxI092_1(.din(n689), .dout(n2011));
    jdff dff_A_RzoDSxuh6_0(.din(n2017), .dout(n2014));
    jdff dff_A_87mnJcZt7_0(.din(n2020), .dout(n2017));
    jdff dff_A_Cn4HUcMZ8_0(.din(n2023), .dout(n2020));
    jdff dff_A_4WHONs2a7_0(.din(n2026), .dout(n2023));
    jdff dff_A_tf2Eq1HF3_0(.din(n2029), .dout(n2026));
    jdff dff_A_5dQwUhWN5_0(.din(n2032), .dout(n2029));
    jdff dff_A_XVPZIjSM2_0(.din(n2035), .dout(n2032));
    jdff dff_A_bKBSNtxC2_0(.din(n2038), .dout(n2035));
    jdff dff_A_hQecb5Yc4_0(.din(n2041), .dout(n2038));
    jdff dff_A_GYxAzLjh8_0(.din(n2044), .dout(n2041));
    jdff dff_A_zSHVQ4E95_0(.din(n2069), .dout(n2044));
    jdff dff_B_nMRYpbD35_2(.din(n682), .dout(n2048));
    jdff dff_B_vCdUxLIY4_2(.din(n2048), .dout(n2051));
    jdff dff_B_ZIWcIQdJ4_2(.din(n2051), .dout(n2054));
    jdff dff_B_JyJZ34XK2_2(.din(n2054), .dout(n2057));
    jdff dff_B_zRU6HOQA3_2(.din(n2057), .dout(n2060));
    jdff dff_B_qAJHj5iF4_2(.din(n2060), .dout(n2063));
    jdff dff_B_Z2zh11bp5_2(.din(n2063), .dout(n2066));
    jdff dff_B_fgU23e0C8_2(.din(n2066), .dout(n2069));
    jdff dff_A_8xMlCICc9_0(.din(n2074), .dout(n2071));
    jdff dff_A_n85eMn4U7_0(.din(n2077), .dout(n2074));
    jdff dff_A_hP8Jo5fs6_0(.din(n2080), .dout(n2077));
    jdff dff_A_3GJcADem5_0(.din(n2083), .dout(n2080));
    jdff dff_A_ayoFeQod0_0(.din(n2086), .dout(n2083));
    jdff dff_A_qpPAXIMO3_0(.din(n2089), .dout(n2086));
    jdff dff_A_wXmZkkXC5_0(.din(n2092), .dout(n2089));
    jdff dff_A_Ztxnv9k10_0(.din(n2095), .dout(n2092));
    jdff dff_A_hzillUTC0_0(.din(n2098), .dout(n2095));
    jdff dff_A_OybFytYO1_0(.din(n2101), .dout(n2098));
    jdff dff_A_kwAPfovI5_0(.din(n2104), .dout(n2101));
    jdff dff_A_T4MwwXy39_0(.din(n2107), .dout(n2104));
    jdff dff_A_0iTrAXob9_0(.din(n2110), .dout(n2107));
    jdff dff_A_piB35lYS0_0(.din(n2113), .dout(n2110));
    jdff dff_A_kYFkFj4w9_0(.din(n2116), .dout(n2113));
    jdff dff_A_pXpSgiNB9_0(.din(n2119), .dout(n2116));
    jdff dff_A_y6Ii1q5d4_0(.din(n2122), .dout(n2119));
    jdff dff_A_KA6riDI94_0(.din(n2125), .dout(n2122));
    jdff dff_A_flqTqVj67_0(.din(n2128), .dout(n2125));
    jdff dff_A_diYIX76x0_0(.din(G40gat), .dout(n2128));
    jdff dff_B_lnn5Uzfq6_1(.din(n675), .dout(n2132));
    jdff dff_B_U98fcXty5_1(.din(n2132), .dout(n2135));
    jdff dff_B_xlcXHhRu7_1(.din(n2135), .dout(n2138));
    jdff dff_B_efK2R0bh5_1(.din(n2138), .dout(n2141));
    jdff dff_B_X67VoH9R1_1(.din(n2141), .dout(n2144));
    jdff dff_B_TGwtTXDD7_1(.din(n2144), .dout(n2147));
    jdff dff_B_00zlxIno6_1(.din(n2147), .dout(n2150));
    jdff dff_B_6KJG3Flh1_1(.din(n2150), .dout(n2153));
    jdff dff_B_fALiyNYM4_1(.din(n2153), .dout(n2156));
    jdff dff_B_z1LzTmC00_1(.din(n2156), .dout(n2159));
    jdff dff_B_B01hDh9Y3_1(.din(n2159), .dout(n2162));
    jdff dff_B_o98iBe3S6_1(.din(n2162), .dout(n2165));
    jdff dff_B_xElPkw5s0_1(.din(n656), .dout(n2168));
    jdff dff_B_W5Y98niU1_1(.din(n2168), .dout(n2171));
    jdff dff_B_1hD0ELZz5_1(.din(n2171), .dout(n2174));
    jdff dff_B_L28FJEj32_1(.din(n2174), .dout(n2177));
    jdff dff_B_bUzvdw0K2_1(.din(n2177), .dout(n2180));
    jdff dff_B_AXbgqMsT7_1(.din(n2180), .dout(n2183));
    jdff dff_B_EGEo9Tis2_1(.din(n2183), .dout(n2186));
    jdff dff_B_krtebK9K0_1(.din(n2186), .dout(n2189));
    jdff dff_B_qitdhjvU1_1(.din(n2189), .dout(n2192));
    jdff dff_B_YrtmM10h8_1(.din(n2192), .dout(n2195));
    jdff dff_B_HmraLxQV5_1(.din(n2195), .dout(n2198));
    jdff dff_B_A6mZnrIx9_1(.din(n2198), .dout(n2201));
    jdff dff_B_IRfLmUY64_1(.din(n2201), .dout(n2204));
    jdff dff_B_dpOwkNU81_1(.din(n2204), .dout(n2207));
    jdff dff_A_TpSj3xwa4_0(.din(n2212), .dout(n2209));
    jdff dff_A_cnwC30Rj0_0(.din(n2215), .dout(n2212));
    jdff dff_A_YUca2dnA6_0(.din(n2218), .dout(n2215));
    jdff dff_A_nyA0KeG70_0(.din(n2221), .dout(n2218));
    jdff dff_A_87Dcb33u9_0(.din(n2224), .dout(n2221));
    jdff dff_A_QRl0R2Rj7_0(.din(n2227), .dout(n2224));
    jdff dff_A_hNQMmCzg6_0(.din(n2230), .dout(n2227));
    jdff dff_A_LLwNLMZU3_0(.din(n2233), .dout(n2230));
    jdff dff_A_zSyOxV917_0(.din(n2236), .dout(n2233));
    jdff dff_A_I6lDnbCy9_0(.din(n2239), .dout(n2236));
    jdff dff_A_aSyy6zo64_0(.din(n2242), .dout(n2239));
    jdff dff_A_aNyeiOYG6_0(.din(n2245), .dout(n2242));
    jdff dff_A_Srj0DVv62_0(.din(n2248), .dout(n2245));
    jdff dff_A_7g9FVgZL0_0(.din(n2251), .dout(n2248));
    jdff dff_A_X0N0VDcb5_0(.din(G14gat), .dout(n2251));
    jdff dff_A_ZqZMyaQl6_1(.din(n2257), .dout(n2254));
    jdff dff_A_aTIWMwVj2_1(.din(n2260), .dout(n2257));
    jdff dff_A_le4NPD2O9_1(.din(n2263), .dout(n2260));
    jdff dff_A_ybQYTo8r8_1(.din(n2266), .dout(n2263));
    jdff dff_A_pLdptZsi5_1(.din(n2269), .dout(n2266));
    jdff dff_A_QL7Q4aix8_1(.din(n2272), .dout(n2269));
    jdff dff_A_vkziZMf91_1(.din(n2275), .dout(n2272));
    jdff dff_A_8zERPKfg0_1(.din(n2278), .dout(n2275));
    jdff dff_A_WxUBDYyB5_1(.din(n2281), .dout(n2278));
    jdff dff_A_GCO729jO1_1(.din(n2284), .dout(n2281));
    jdff dff_A_Sg2vU5sp9_1(.din(n2287), .dout(n2284));
    jdff dff_A_n2X8c3xd3_1(.din(n2290), .dout(n2287));
    jdff dff_A_bQX8fFmd2_1(.din(n2293), .dout(n2290));
    jdff dff_A_FukfDVB72_1(.din(n2296), .dout(n2293));
    jdff dff_A_IVEt6Yi41_1(.din(n2299), .dout(n2296));
    jdff dff_A_rnL2bv6w1_1(.din(n2302), .dout(n2299));
    jdff dff_A_9zWOeDKj4_1(.din(n2305), .dout(n2302));
    jdff dff_A_PX4wzWm83_1(.din(n2308), .dout(n2305));
    jdff dff_A_F43mayrn8_1(.din(n2311), .dout(n2308));
    jdff dff_A_reYrKxhI4_1(.din(G14gat), .dout(n2311));
    jdff dff_A_5O11Kk6m7_0(.din(n2317), .dout(n2314));
    jdff dff_A_jHfTwugk2_0(.din(n2320), .dout(n2317));
    jdff dff_A_Z39AWxCp2_0(.din(n2323), .dout(n2320));
    jdff dff_A_QncNGc8c7_0(.din(n2326), .dout(n2323));
    jdff dff_A_OnOWwz199_0(.din(n2329), .dout(n2326));
    jdff dff_A_mutchN9n9_0(.din(n2369), .dout(n2329));
    jdff dff_B_5na9E6hu8_2(.din(n641), .dout(n2333));
    jdff dff_B_lldkz9KD6_2(.din(n2333), .dout(n2336));
    jdff dff_B_eXp3ymoj3_2(.din(n2336), .dout(n2339));
    jdff dff_B_w50sHWmX1_2(.din(n2339), .dout(n2342));
    jdff dff_B_momk3OCZ7_2(.din(n2342), .dout(n2345));
    jdff dff_B_VPnhVvQf6_2(.din(n2345), .dout(n2348));
    jdff dff_B_i7T2ylon8_2(.din(n2348), .dout(n2351));
    jdff dff_B_Hg1wGNpr9_2(.din(n2351), .dout(n2354));
    jdff dff_B_XQEDxvVJ3_2(.din(n2354), .dout(n2357));
    jdff dff_B_8WWWUYmp0_2(.din(n2357), .dout(n2360));
    jdff dff_B_pPgTgPVb9_2(.din(n2360), .dout(n2363));
    jdff dff_B_b3BVX2oY0_2(.din(n2363), .dout(n2366));
    jdff dff_B_uUvTNaPX9_2(.din(n2366), .dout(n2369));
    jdff dff_A_2VNDQKNF4_0(.din(n2374), .dout(n2371));
    jdff dff_A_VRPZQ8vi8_0(.din(n2377), .dout(n2374));
    jdff dff_A_K0v8OTU29_0(.din(n2380), .dout(n2377));
    jdff dff_A_6O5rJf7T4_0(.din(n2383), .dout(n2380));
    jdff dff_A_6cl3ISZv3_0(.din(n2386), .dout(n2383));
    jdff dff_A_dLTShI6e4_0(.din(n2389), .dout(n2386));
    jdff dff_A_lEY5TJhc5_0(.din(n2392), .dout(n2389));
    jdff dff_A_YSebzq7q0_0(.din(n2395), .dout(n2392));
    jdff dff_A_EPWGFcJD8_0(.din(n2398), .dout(n2395));
    jdff dff_A_IVYwyVLb4_0(.din(n2401), .dout(n2398));
    jdff dff_A_TNf5Xzci9_0(.din(n2404), .dout(n2401));
    jdff dff_A_SRzfEq2P7_0(.din(n2407), .dout(n2404));
    jdff dff_A_Sa2BPSPj2_0(.din(n2410), .dout(n2407));
    jdff dff_A_ZNR42zaU9_0(.din(n2413), .dout(n2410));
    jdff dff_A_RlohIgWY0_0(.din(n2416), .dout(n2413));
    jdff dff_A_8YKBPe6X5_0(.din(n2419), .dout(n2416));
    jdff dff_A_Xs0xBlaI4_0(.din(n2422), .dout(n2419));
    jdff dff_A_xMwM09Dw7_0(.din(n2425), .dout(n2422));
    jdff dff_A_ec6FnCUB3_0(.din(n2428), .dout(n2425));
    jdff dff_A_hTvL5vzG1_0(.din(G92gat), .dout(n2428));
    jdff dff_A_83dePEjo1_1(.din(n2434), .dout(n2431));
    jdff dff_A_2kmHN2nr2_1(.din(n2437), .dout(n2434));
    jdff dff_A_bICRxTcp6_1(.din(n2440), .dout(n2437));
    jdff dff_A_A6pcBdQW9_1(.din(n2443), .dout(n2440));
    jdff dff_A_dqA1iTsp5_1(.din(n2446), .dout(n2443));
    jdff dff_A_2p6TzBdR0_1(.din(n2449), .dout(n2446));
    jdff dff_A_nOdvEM2O8_1(.din(n2452), .dout(n2449));
    jdff dff_A_lem8xaPx7_1(.din(n2455), .dout(n2452));
    jdff dff_A_w29xGCwv0_1(.din(n2458), .dout(n2455));
    jdff dff_A_EyvGYo8f4_1(.din(n2461), .dout(n2458));
    jdff dff_A_rNyqQz2R0_1(.din(n2464), .dout(n2461));
    jdff dff_A_ZkEt66zK0_1(.din(n2467), .dout(n2464));
    jdff dff_A_b8m4tGwy5_1(.din(n2470), .dout(n2467));
    jdff dff_A_Cja6zkSj7_1(.din(G92gat), .dout(n2470));
    jdff dff_A_lzEL013z8_0(.din(n2476), .dout(n2473));
    jdff dff_A_HitMEIcW0_0(.din(n2479), .dout(n2476));
    jdff dff_A_Z1SZBG4I3_0(.din(n2482), .dout(n2479));
    jdff dff_A_vgxR4BZu9_0(.din(n2485), .dout(n2482));
    jdff dff_A_OcK3Z1p87_0(.din(n2488), .dout(n2485));
    jdff dff_A_kJY4IHWD0_0(.din(n638), .dout(n2488));
    jdff dff_A_VlCqvEiy4_0(.din(n2494), .dout(n2491));
    jdff dff_A_3UtBEZuj6_0(.din(n2497), .dout(n2494));
    jdff dff_A_fHwwK6F40_0(.din(n2500), .dout(n2497));
    jdff dff_A_UKVnAVN40_0(.din(n2503), .dout(n2500));
    jdff dff_A_gGr99vMR6_0(.din(n2506), .dout(n2503));
    jdff dff_A_0CyklLM18_0(.din(n2546), .dout(n2506));
    jdff dff_B_qUqSm9GJ4_2(.din(n614), .dout(n2510));
    jdff dff_B_7fuvmvCx4_2(.din(n2510), .dout(n2513));
    jdff dff_B_az7TCeYd7_2(.din(n2513), .dout(n2516));
    jdff dff_B_7RL1TIQc5_2(.din(n2516), .dout(n2519));
    jdff dff_B_SVdhd0Dc8_2(.din(n2519), .dout(n2522));
    jdff dff_B_0MyRwGPc8_2(.din(n2522), .dout(n2525));
    jdff dff_B_D9yHKpXV5_2(.din(n2525), .dout(n2528));
    jdff dff_B_np3gfNno3_2(.din(n2528), .dout(n2531));
    jdff dff_B_XoQwXwxj0_2(.din(n2531), .dout(n2534));
    jdff dff_B_BAQRRF1l2_2(.din(n2534), .dout(n2537));
    jdff dff_B_5VtNxWne5_2(.din(n2537), .dout(n2540));
    jdff dff_B_XBhqH1475_2(.din(n2540), .dout(n2543));
    jdff dff_B_fyrZXCvG0_2(.din(n2543), .dout(n2546));
    jdff dff_A_P4E9OfrU2_0(.din(n2551), .dout(n2548));
    jdff dff_A_NfnO9f7r4_0(.din(n2554), .dout(n2551));
    jdff dff_A_oF9666GH5_0(.din(n2557), .dout(n2554));
    jdff dff_A_TMJ6cU6F7_0(.din(n2560), .dout(n2557));
    jdff dff_A_q40O1sGG4_0(.din(n2563), .dout(n2560));
    jdff dff_A_KdSzsY7L4_0(.din(n2566), .dout(n2563));
    jdff dff_A_TDSvuKZa7_0(.din(n2569), .dout(n2566));
    jdff dff_A_Z0zALdGJ2_0(.din(n2572), .dout(n2569));
    jdff dff_A_14tCVaq02_0(.din(n2575), .dout(n2572));
    jdff dff_A_9ASsQCif4_0(.din(n2578), .dout(n2575));
    jdff dff_A_Yb4EtMYG4_0(.din(n2581), .dout(n2578));
    jdff dff_A_AOjEDhQx8_0(.din(n2584), .dout(n2581));
    jdff dff_A_NeiQxvBq5_0(.din(n2587), .dout(n2584));
    jdff dff_A_O0PhjXJJ1_0(.din(G27gat), .dout(n2587));
    jdff dff_A_3DkbUKqV4_0(.din(n2593), .dout(n2590));
    jdff dff_A_q4PeoTyl5_0(.din(n2596), .dout(n2593));
    jdff dff_A_32hI6N2n9_0(.din(n2599), .dout(n2596));
    jdff dff_A_IYUO0ecr1_0(.din(n2602), .dout(n2599));
    jdff dff_A_11nRX98N3_0(.din(n2605), .dout(n2602));
    jdff dff_A_T30xqLpp4_0(.din(n611), .dout(n2605));
    jdff dff_A_2gpDt1rw1_1(.din(n2611), .dout(n2608));
    jdff dff_A_z4WWpocZ0_1(.din(n2614), .dout(n2611));
    jdff dff_A_BiEMJDwr2_1(.din(n2617), .dout(n2614));
    jdff dff_A_x3s1wrdr0_1(.din(n2620), .dout(n2617));
    jdff dff_A_CUXDsklJ4_1(.din(n2623), .dout(n2620));
    jdff dff_A_9Jbz5w6N9_1(.din(n2626), .dout(n2623));
    jdff dff_A_s6t7iNYI6_1(.din(n599), .dout(n2626));
    jdff dff_B_4QZ46xG08_0(.din(n595), .dout(n2630));
    jdff dff_B_b6nSR68a2_0(.din(n2630), .dout(n2633));
    jdff dff_B_NJHj4LJQ3_0(.din(n2633), .dout(n2636));
    jdff dff_B_cylbLnVE1_0(.din(n2636), .dout(n2639));
    jdff dff_B_0xlbnkxf7_0(.din(n2639), .dout(n2642));
    jdff dff_A_kkuwY2iN0_0(.din(n2647), .dout(n2644));
    jdff dff_A_xEo5DSXc0_0(.din(n2650), .dout(n2647));
    jdff dff_A_JxBinVoZ4_0(.din(n2653), .dout(n2650));
    jdff dff_A_nUTgCvt80_0(.din(n2656), .dout(n2653));
    jdff dff_A_r7iu4eT31_0(.din(n2659), .dout(n2656));
    jdff dff_A_PZtx4D5a9_0(.din(n2662), .dout(n2659));
    jdff dff_A_D1zSyuGG8_0(.din(n2665), .dout(n2662));
    jdff dff_A_4WhcggbI7_0(.din(n2668), .dout(n2665));
    jdff dff_A_6VDJmKIe8_0(.din(n2671), .dout(n2668));
    jdff dff_A_AGZU92X91_0(.din(n2674), .dout(n2671));
    jdff dff_A_7EfEMMAw2_0(.din(n2677), .dout(n2674));
    jdff dff_A_gn9Dwxgk1_0(.din(n2680), .dout(n2677));
    jdff dff_A_nbLpy6kM5_0(.din(n2683), .dout(n2680));
    jdff dff_A_JYv7xi7H3_0(.din(n2686), .dout(n2683));
    jdff dff_A_Y4jSUqGe3_0(.din(n2689), .dout(n2686));
    jdff dff_A_1xfANVUj8_0(.din(n2692), .dout(n2689));
    jdff dff_A_wYFRCQu26_0(.din(n2695), .dout(n2692));
    jdff dff_A_CHVy6Qct6_0(.din(n2698), .dout(n2695));
    jdff dff_A_NztlICNx4_0(.din(n591), .dout(n2698));
    jdff dff_A_K70pXfwm2_0(.din(n2704), .dout(n2701));
    jdff dff_A_rhgUzpww6_0(.din(n2707), .dout(n2704));
    jdff dff_A_lPudnZzQ4_0(.din(n2710), .dout(n2707));
    jdff dff_A_Tqzg5ZiU4_0(.din(n2713), .dout(n2710));
    jdff dff_A_is7xcMgr9_0(.din(n2716), .dout(n2713));
    jdff dff_A_ZSidA31H8_0(.din(n2719), .dout(n2716));
    jdff dff_A_AdleOg1T4_0(.din(n2722), .dout(n2719));
    jdff dff_A_2kr83mvm7_0(.din(n2725), .dout(n2722));
    jdff dff_A_7YB8gEZS0_0(.din(n2728), .dout(n2725));
    jdff dff_A_72YPSi479_0(.din(n2731), .dout(n2728));
    jdff dff_A_g7Y78fgg7_0(.din(n2734), .dout(n2731));
    jdff dff_A_ijzhXmIl2_0(.din(n2737), .dout(n2734));
    jdff dff_A_5mq645bi0_0(.din(n2740), .dout(n2737));
    jdff dff_A_vOdb2YxJ8_0(.din(n2743), .dout(n2740));
    jdff dff_A_Rp8YjN2A0_0(.din(n2746), .dout(n2743));
    jdff dff_A_wXz8MI1r6_0(.din(n2749), .dout(n2746));
    jdff dff_A_iPjsRmrz4_0(.din(n2752), .dout(n2749));
    jdff dff_A_Qiowc9UD7_0(.din(n2755), .dout(n2752));
    jdff dff_A_eS2VW7jv4_0(.din(n2758), .dout(n2755));
    jdff dff_A_OYC4wMHD3_0(.din(G53gat), .dout(n2758));
    jdff dff_A_rvv8PztO5_0(.din(n2764), .dout(n2761));
    jdff dff_A_39boRS979_0(.din(n2767), .dout(n2764));
    jdff dff_A_NvpKZUwL4_0(.din(n2770), .dout(n2767));
    jdff dff_A_ySeg3elV5_0(.din(n2773), .dout(n2770));
    jdff dff_A_CfgtonVu2_0(.din(n2776), .dout(n2773));
    jdff dff_A_ajlO7iq04_0(.din(n569), .dout(n2776));
    jdff dff_B_TULCKkIv7_1(.din(n503), .dout(n2780));
    jdff dff_A_lOfZMnf54_0(.din(n2785), .dout(n2782));
    jdff dff_A_n6hXZ9SH3_0(.din(n2788), .dout(n2785));
    jdff dff_A_jUYZU3kF9_0(.din(n2791), .dout(n2788));
    jdff dff_A_gevSWNzF0_0(.din(n2794), .dout(n2791));
    jdff dff_A_6BGROkuE9_0(.din(n2797), .dout(n2794));
    jdff dff_A_eV97XeUj9_0(.din(n541), .dout(n2797));
    jdff dff_A_Kf3ddpAR8_0(.din(n2803), .dout(n2800));
    jdff dff_A_AC3V1HOO4_0(.din(n2806), .dout(n2803));
    jdff dff_A_WE7qvhvl3_0(.din(n2809), .dout(n2806));
    jdff dff_A_VMbfIxYJ9_0(.din(n2812), .dout(n2809));
    jdff dff_A_Iyn24Ir93_0(.din(n2815), .dout(n2812));
    jdff dff_A_1NHobVf29_0(.din(n529), .dout(n2815));
    jdff dff_B_OOZQruHx0_1(.din(n521), .dout(n2819));
    jdff dff_B_c5c18Uis1_1(.din(n2819), .dout(n2822));
    jdff dff_B_PVqFOUhM9_1(.din(n2822), .dout(n2825));
    jdff dff_B_sgkt7iPm9_1(.din(n2825), .dout(n2828));
    jdff dff_B_5SkpzC2A4_1(.din(n2828), .dout(n2831));
    jdff dff_B_vuzsV2FC6_1(.din(n2831), .dout(n2834));
    jdff dff_A_nC9RLLDY4_0(.din(n2839), .dout(n2836));
    jdff dff_A_fSU0j8Yn2_0(.din(n2842), .dout(n2839));
    jdff dff_A_5UjwFNuN8_0(.din(n2845), .dout(n2842));
    jdff dff_A_I0B4DkU05_0(.din(n2849), .dout(n2845));
    jdff dff_B_DacFIcBk5_2(.din(n514), .dout(n2849));
    jdff dff_B_i2Sflq2H1_0(.din(n510), .dout(n2852));
    jdff dff_B_SlHUmUsE1_0(.din(n2852), .dout(n2855));
    jdff dff_B_nQ6YaW0S4_0(.din(n2855), .dout(n2858));
    jdff dff_B_i8ozyrsk5_0(.din(n2858), .dout(n2861));
    jdff dff_A_mIghtVWN7_0(.din(n2866), .dout(n2863));
    jdff dff_A_U6hHS9oy6_0(.din(n2869), .dout(n2866));
    jdff dff_A_3A1so0WA4_0(.din(n2872), .dout(n2869));
    jdff dff_A_M2mwOCZz0_0(.din(n2875), .dout(n2872));
    jdff dff_A_2TjCq7Hh6_0(.din(n2878), .dout(n2875));
    jdff dff_A_P8mWUwpS3_0(.din(n491), .dout(n2878));
    jdff dff_A_X4qN0ZtE2_0(.din(n2884), .dout(n2881));
    jdff dff_A_ZnHftyNV4_0(.din(n2887), .dout(n2884));
    jdff dff_A_9cQavNd13_0(.din(n2890), .dout(n2887));
    jdff dff_A_pbaOLV8f9_0(.din(n2893), .dout(n2890));
    jdff dff_A_Ar5obENu8_0(.din(n2896), .dout(n2893));
    jdff dff_A_3fWF9Vay3_0(.din(n471), .dout(n2896));
    jdff dff_A_X9fM55LS2_0(.din(n2902), .dout(n2899));
    jdff dff_A_5Q738wrw6_0(.din(n2905), .dout(n2902));
    jdff dff_A_DATfAEHS4_0(.din(n2908), .dout(n2905));
    jdff dff_A_gVjaJtsn2_0(.din(n2911), .dout(n2908));
    jdff dff_A_bRsrjABE0_0(.din(n2914), .dout(n2911));
    jdff dff_A_ZOGdPGs42_0(.din(n459), .dout(n2914));
    jdff dff_A_upZOs5PZ5_0(.din(n2920), .dout(n2917));
    jdff dff_A_BdUgGSAh2_0(.din(n2923), .dout(n2920));
    jdff dff_A_Nc2x7Jwl2_0(.din(n2926), .dout(n2923));
    jdff dff_A_1mU1ZLEm8_0(.din(n2929), .dout(n2926));
    jdff dff_A_nl7IyFXG9_0(.din(n2972), .dout(n2929));
    jdff dff_B_ih3E6Wpi6_2(.din(n451), .dout(n2933));
    jdff dff_B_D617FD3g6_2(.din(n2933), .dout(n2936));
    jdff dff_B_TAsBmQD71_2(.din(n2936), .dout(n2939));
    jdff dff_B_m9OscV3G6_2(.din(n2939), .dout(n2942));
    jdff dff_B_0C65iaNx5_2(.din(n2942), .dout(n2945));
    jdff dff_B_f4x8NmUE9_2(.din(n2945), .dout(n2948));
    jdff dff_B_6g7kN7jm8_2(.din(n2948), .dout(n2951));
    jdff dff_B_MybpwxhO4_2(.din(n2951), .dout(n2954));
    jdff dff_B_Rv3whGh50_2(.din(n2954), .dout(n2957));
    jdff dff_B_ujhZzmE93_2(.din(n2957), .dout(n2960));
    jdff dff_B_p9htagI23_2(.din(n2960), .dout(n2963));
    jdff dff_B_7tnf8wmb0_2(.din(n2963), .dout(n2966));
    jdff dff_B_IR8Bvya77_2(.din(n2966), .dout(n2969));
    jdff dff_B_ynVHqGdP0_2(.din(n2969), .dout(n2972));
    jdff dff_A_3OPq8lC90_0(.din(n2977), .dout(n2974));
    jdff dff_A_qLM8c9x33_0(.din(n2980), .dout(n2977));
    jdff dff_A_K8uVWCHg2_0(.din(n2983), .dout(n2980));
    jdff dff_A_wQUjB8Sy9_0(.din(n2986), .dout(n2983));
    jdff dff_A_dLf5Wvxq3_0(.din(n2989), .dout(n2986));
    jdff dff_A_3QiR7ewA2_0(.din(n2992), .dout(n2989));
    jdff dff_A_iWa6xviI8_0(.din(n2995), .dout(n2992));
    jdff dff_A_eklnG9MQ6_0(.din(n2998), .dout(n2995));
    jdff dff_A_GBFYKOkz5_0(.din(n3001), .dout(n2998));
    jdff dff_A_c63E0tea8_0(.din(n3004), .dout(n3001));
    jdff dff_A_qMmAYXyr9_0(.din(n3007), .dout(n3004));
    jdff dff_A_qahQb5Qc7_0(.din(n3010), .dout(n3007));
    jdff dff_A_FT22x3K41_0(.din(n3013), .dout(n3010));
    jdff dff_A_FjkyvDqN9_0(.din(n3016), .dout(n3013));
    jdff dff_A_IcPR62ao3_0(.din(G79gat), .dout(n3016));
    jdff dff_A_dMFpHtVm4_1(.din(n3022), .dout(n3019));
    jdff dff_A_7bWL3VEH3_1(.din(n3025), .dout(n3022));
    jdff dff_A_3vDhBz6t5_1(.din(n3028), .dout(n3025));
    jdff dff_A_d05E4w361_1(.din(n3031), .dout(n3028));
    jdff dff_A_2wwBRVl54_1(.din(n3034), .dout(n3031));
    jdff dff_A_iswuUbvY4_1(.din(n444), .dout(n3034));
    jdff dff_A_wSS7Uavd7_0(.din(n3040), .dout(n3037));
    jdff dff_A_ahDzLQV77_0(.din(n3043), .dout(n3040));
    jdff dff_A_tyBqzzah5_0(.din(n3046), .dout(n3043));
    jdff dff_A_lkFuCNfX4_0(.din(n3049), .dout(n3046));
    jdff dff_A_YbFSinoe7_0(.din(n3052), .dout(n3049));
    jdff dff_A_t3Hryi672_0(.din(n3055), .dout(n3052));
    jdff dff_A_yj0eJcbk9_0(.din(n3058), .dout(n3055));
    jdff dff_A_iS7P584Y7_0(.din(n3061), .dout(n3058));
    jdff dff_A_R5mgsJEh5_0(.din(n3064), .dout(n3061));
    jdff dff_A_KNtmxcGp2_0(.din(n3067), .dout(n3064));
    jdff dff_A_FP4D0iMU9_0(.din(n3070), .dout(n3067));
    jdff dff_A_b787DLJQ7_0(.din(n3092), .dout(n3070));
    jdff dff_B_3suSYngp4_2(.din(n440), .dout(n3074));
    jdff dff_B_ryLnhs7O7_2(.din(n3074), .dout(n3077));
    jdff dff_B_nck2wWvV9_2(.din(n3077), .dout(n3080));
    jdff dff_B_SgbJxtLR8_2(.din(n3080), .dout(n3083));
    jdff dff_B_1bgoMqsc2_2(.din(n3083), .dout(n3086));
    jdff dff_B_4737DIKd2_2(.din(n3086), .dout(n3089));
    jdff dff_B_oJ0khUTh6_2(.din(n3089), .dout(n3092));
    jdff dff_A_CBhlU5Vi0_0(.din(n3097), .dout(n3094));
    jdff dff_A_Rhp8TIeZ8_0(.din(n3100), .dout(n3097));
    jdff dff_A_hqIttyzW7_0(.din(n3103), .dout(n3100));
    jdff dff_A_ggH5p7q20_0(.din(n3106), .dout(n3103));
    jdff dff_A_4LvNKKTI7_0(.din(n3109), .dout(n3106));
    jdff dff_A_2Aj9k8949_0(.din(n3112), .dout(n3109));
    jdff dff_A_WvQViioJ4_0(.din(n3115), .dout(n3112));
    jdff dff_A_36KIvm9k9_0(.din(n3118), .dout(n3115));
    jdff dff_A_rrQ8oGqq8_0(.din(n3121), .dout(n3118));
    jdff dff_A_grHjRU1c6_0(.din(n3124), .dout(n3121));
    jdff dff_A_38u79YLn2_0(.din(n3127), .dout(n3124));
    jdff dff_A_Ip7mFw6K8_0(.din(n3130), .dout(n3127));
    jdff dff_A_ylJ6p2Hj3_0(.din(n3133), .dout(n3130));
    jdff dff_A_lpLg8iFg3_0(.din(n3136), .dout(n3133));
    jdff dff_A_tbpptluP1_0(.din(n3139), .dout(n3136));
    jdff dff_A_MxJo78O71_0(.din(n3142), .dout(n3139));
    jdff dff_A_LPShTF3E9_0(.din(n3145), .dout(n3142));
    jdff dff_A_YLc1MDH15_0(.din(n3148), .dout(n3145));
    jdff dff_A_TfSFkQUk7_0(.din(n3151), .dout(n3148));
    jdff dff_A_4L7SPVuI9_0(.din(G66gat), .dout(n3151));
    jdff dff_A_qKQ1EjVd3_1(.din(n3157), .dout(n3154));
    jdff dff_A_CWr6yg7X2_1(.din(n3160), .dout(n3157));
    jdff dff_A_OPhQx6q53_1(.din(n3163), .dout(n3160));
    jdff dff_A_YDMdgSf06_1(.din(n430), .dout(n3163));
    jdff dff_A_NHH8y1P76_0(.din(n3169), .dout(n3166));
    jdff dff_A_dy9ywEpf3_0(.din(n3172), .dout(n3169));
    jdff dff_A_4Yn67P8E2_0(.din(n3175), .dout(n3172));
    jdff dff_A_36qhM1LE6_0(.din(n3178), .dout(n3175));
    jdff dff_A_rqGOiAIo8_0(.din(n3181), .dout(n3178));
    jdff dff_A_jggaCk2R5_0(.din(n426), .dout(n3181));
    jdff dff_A_TH3VM6Wq8_0(.din(n415), .dout(n3184));
    jdff dff_B_L8xAIm631_1(.din(n300), .dout(n3188));
    jdff dff_B_5HVIxTto7_1(.din(n315), .dout(n3191));
    jdff dff_A_KvN69eRv0_0(.din(n3196), .dout(n3193));
    jdff dff_A_8qC8Bxil9_0(.din(n3199), .dout(n3196));
    jdff dff_A_Ahft7AOV4_0(.din(n3202), .dout(n3199));
    jdff dff_A_EvMmlDyf5_0(.din(n3205), .dout(n3202));
    jdff dff_A_0KBaRO998_0(.din(n3208), .dout(n3205));
    jdff dff_A_HxjKhfpm3_0(.din(n375), .dout(n3208));
    jdff dff_A_FYfj79HQ6_0(.din(n3214), .dout(n3211));
    jdff dff_A_nqUp2RTk9_0(.din(n3217), .dout(n3214));
    jdff dff_A_5TRk2knt2_0(.din(n3220), .dout(n3217));
    jdff dff_A_55IHtMGb3_0(.din(n3223), .dout(n3220));
    jdff dff_A_ikW0gD047_0(.din(n3260), .dout(n3223));
    jdff dff_A_rvw2qnGv6_1(.din(n3229), .dout(n3226));
    jdff dff_A_LzYGizPC2_1(.din(n3232), .dout(n3229));
    jdff dff_A_SrzJZZRR9_1(.din(n3235), .dout(n3232));
    jdff dff_A_8EMDDm7r3_1(.din(n3238), .dout(n3235));
    jdff dff_A_Ss3t7B913_1(.din(n3260), .dout(n3238));
    jdff dff_B_esKR7kkk1_3(.din(n367), .dout(n3242));
    jdff dff_B_yQY2moTH4_3(.din(n3242), .dout(n3245));
    jdff dff_B_oeXp4PmU3_3(.din(n3245), .dout(n3248));
    jdff dff_B_ttlJSbP61_3(.din(n3248), .dout(n3251));
    jdff dff_B_Qfl55UKq8_3(.din(n3251), .dout(n3254));
    jdff dff_B_mKkf82ms6_3(.din(n3254), .dout(n3257));
    jdff dff_B_duBsfNaE5_3(.din(n3257), .dout(n3260));
    jdff dff_A_hnpq7YPZ0_0(.din(n3265), .dout(n3262));
    jdff dff_A_6ZzR6NVO8_0(.din(n3268), .dout(n3265));
    jdff dff_A_IhUCNGIH8_0(.din(n3271), .dout(n3268));
    jdff dff_A_yaCqGn8t2_0(.din(n3274), .dout(n3271));
    jdff dff_A_unDrCpin6_0(.din(n3277), .dout(n3274));
    jdff dff_A_alPvvsFh2_0(.din(n3280), .dout(n3277));
    jdff dff_A_Mr5eIYlc5_0(.din(n3283), .dout(n3280));
    jdff dff_A_6wYury1T2_0(.din(G21gat), .dout(n3283));
    jdff dff_A_vz536jsF4_1(.din(n3289), .dout(n3286));
    jdff dff_A_zOFjjEo51_1(.din(n3292), .dout(n3289));
    jdff dff_A_OjvD6dLG8_1(.din(n3295), .dout(n3292));
    jdff dff_A_JjBEHFzh0_1(.din(n3298), .dout(n3295));
    jdff dff_A_GIjglU9u6_1(.din(n3301), .dout(n3298));
    jdff dff_A_elrsTPmC6_1(.din(n3304), .dout(n3301));
    jdff dff_A_gzX4iWzT6_1(.din(n3307), .dout(n3304));
    jdff dff_A_wf3DvDfL8_1(.din(n3310), .dout(n3307));
    jdff dff_A_WHh6n79A7_1(.din(n3313), .dout(n3310));
    jdff dff_A_LSGuI2nP5_1(.din(n3316), .dout(n3313));
    jdff dff_A_MIwgaU5U1_1(.din(n3319), .dout(n3316));
    jdff dff_A_BmWdvScP5_1(.din(n3322), .dout(n3319));
    jdff dff_A_ylkeI8A80_1(.din(G21gat), .dout(n3322));
    jdff dff_A_P90YzDTl9_2(.din(n3328), .dout(n3325));
    jdff dff_A_kkPlUJ2S0_2(.din(n3331), .dout(n3328));
    jdff dff_A_boGCpCYk7_2(.din(n3334), .dout(n3331));
    jdff dff_A_r0km9SAv1_2(.din(n3337), .dout(n3334));
    jdff dff_A_cbe27X4j3_2(.din(n3340), .dout(n3337));
    jdff dff_A_FtHp9jB85_2(.din(n3343), .dout(n3340));
    jdff dff_A_1cc9wIDL4_2(.din(n3346), .dout(n3343));
    jdff dff_A_2S56qNHh7_2(.din(n3349), .dout(n3346));
    jdff dff_A_ngVAlWUj2_2(.din(n3352), .dout(n3349));
    jdff dff_A_1LyjpzAE0_2(.din(n3355), .dout(n3352));
    jdff dff_A_8bhxMlF20_2(.din(n3358), .dout(n3355));
    jdff dff_A_CgRXMc1o9_2(.din(n3361), .dout(n3358));
    jdff dff_A_8CzVoGhG7_2(.din(G21gat), .dout(n3361));
    jdff dff_A_pCSGokb38_0(.din(n3367), .dout(n3364));
    jdff dff_A_IWZY9deA1_0(.din(n3370), .dout(n3367));
    jdff dff_A_Qx3ogJgN7_0(.din(n3373), .dout(n3370));
    jdff dff_A_xCyHPCLS3_0(.din(n3376), .dout(n3373));
    jdff dff_A_dRSkMPP55_0(.din(n3379), .dout(n3376));
    jdff dff_A_nFqf8QzF1_0(.din(n360), .dout(n3379));
    jdff dff_A_2zuZ6jFB0_0(.din(n3385), .dout(n3382));
    jdff dff_A_D64y7Lok3_0(.din(n3388), .dout(n3385));
    jdff dff_A_nfY9ctfx9_0(.din(n3391), .dout(n3388));
    jdff dff_A_6DMYWMBQ7_0(.din(n3394), .dout(n3391));
    jdff dff_A_QLBicpOR7_0(.din(n3431), .dout(n3394));
    jdff dff_A_C7ESVwgH7_1(.din(n3400), .dout(n3397));
    jdff dff_A_SNot2wgA3_1(.din(n3403), .dout(n3400));
    jdff dff_A_p5ML6ha55_1(.din(n3406), .dout(n3403));
    jdff dff_A_sgt5feMI3_1(.din(n3409), .dout(n3406));
    jdff dff_A_u7RDWOiz3_1(.din(n3431), .dout(n3409));
    jdff dff_B_7iFtbWKM7_3(.din(n352), .dout(n3413));
    jdff dff_B_uckc6IQQ9_3(.din(n3413), .dout(n3416));
    jdff dff_B_GtsIZzQw2_3(.din(n3416), .dout(n3419));
    jdff dff_B_QL9zLZh95_3(.din(n3419), .dout(n3422));
    jdff dff_B_C9hIiv3k6_3(.din(n3422), .dout(n3425));
    jdff dff_B_DnfFyvX56_3(.din(n3425), .dout(n3428));
    jdff dff_B_SWO0A4BS1_3(.din(n3428), .dout(n3431));
    jdff dff_A_kcobK8Is2_0(.din(n3436), .dout(n3433));
    jdff dff_A_CQM9eZFe7_0(.din(n3439), .dout(n3436));
    jdff dff_A_slPQWZ2C3_0(.din(n3442), .dout(n3439));
    jdff dff_A_TFALbzua9_0(.din(n3445), .dout(n3442));
    jdff dff_A_9EKSZZo06_0(.din(n3448), .dout(n3445));
    jdff dff_A_cjXAEE6s3_0(.din(n3451), .dout(n3448));
    jdff dff_A_BtYnkijl0_0(.din(n3454), .dout(n3451));
    jdff dff_A_zpvm1eo74_0(.din(G86gat), .dout(n3454));
    jdff dff_A_yvnGjsRs8_1(.din(n3460), .dout(n3457));
    jdff dff_A_rw8qT8P43_1(.din(n3463), .dout(n3460));
    jdff dff_A_jlDVpJ7x8_1(.din(n3466), .dout(n3463));
    jdff dff_A_bOKXQDzp5_1(.din(n3469), .dout(n3466));
    jdff dff_A_ve1rEFdc6_1(.din(n3472), .dout(n3469));
    jdff dff_A_sVMokOZU3_1(.din(n3475), .dout(n3472));
    jdff dff_A_KFc4OUjj6_1(.din(n3478), .dout(n3475));
    jdff dff_A_GPzwGosk0_1(.din(n3481), .dout(n3478));
    jdff dff_A_lRCmjHhC6_1(.din(n3484), .dout(n3481));
    jdff dff_A_0xwpSxdc4_1(.din(n3487), .dout(n3484));
    jdff dff_A_4OjroygO6_1(.din(n3490), .dout(n3487));
    jdff dff_A_xsWauW9u4_1(.din(n3493), .dout(n3490));
    jdff dff_A_3RY14p7Q2_1(.din(G86gat), .dout(n3493));
    jdff dff_A_ABVZFhL37_2(.din(n3499), .dout(n3496));
    jdff dff_A_zuVWxMWC9_2(.din(n3502), .dout(n3499));
    jdff dff_A_WNcFqDLe9_2(.din(n3505), .dout(n3502));
    jdff dff_A_fzOGFt1a7_2(.din(n3508), .dout(n3505));
    jdff dff_A_ubA3NRgw2_2(.din(n3511), .dout(n3508));
    jdff dff_A_OOhARacv6_2(.din(n3514), .dout(n3511));
    jdff dff_A_hE7n0a4I7_2(.din(n3517), .dout(n3514));
    jdff dff_A_UoDmrJph5_2(.din(n3520), .dout(n3517));
    jdff dff_A_zIohYmyg3_2(.din(n3523), .dout(n3520));
    jdff dff_A_Bq1laqnH5_2(.din(n3526), .dout(n3523));
    jdff dff_A_RsgW4ij96_2(.din(n3529), .dout(n3526));
    jdff dff_A_ktF3Za192_2(.din(n3532), .dout(n3529));
    jdff dff_A_kTePh0YY1_2(.din(G86gat), .dout(n3532));
    jdff dff_B_rsRN4gi21_0(.din(n345), .dout(n3536));
    jdff dff_A_DD2EwS6E1_1(.din(n3541), .dout(n3538));
    jdff dff_A_3mO9yJA19_1(.din(n3544), .dout(n3541));
    jdff dff_A_GqZtSLYu0_1(.din(n3547), .dout(n3544));
    jdff dff_A_LNLRBGh42_1(.din(n3550), .dout(n3547));
    jdff dff_A_0GVK19w73_1(.din(n341), .dout(n3550));
    jdff dff_A_EUSJa4NQ3_0(.din(n3556), .dout(n3553));
    jdff dff_A_UzJrRbZe3_0(.din(n3559), .dout(n3556));
    jdff dff_A_vFgpuMpX8_0(.din(n3562), .dout(n3559));
    jdff dff_A_jJt15PHk3_0(.din(n3565), .dout(n3562));
    jdff dff_A_gObTqNUE4_0(.din(n3568), .dout(n3565));
    jdff dff_A_jE8scXq03_0(.din(n3571), .dout(n3568));
    jdff dff_A_qyEOFRol2_0(.din(n3574), .dout(n3571));
    jdff dff_A_RezMjxAs2_0(.din(n3577), .dout(n3574));
    jdff dff_A_s2sk7ri67_0(.din(n3580), .dout(n3577));
    jdff dff_A_0Hp699qs0_0(.din(n3583), .dout(n3580));
    jdff dff_A_4bkjgAZJ1_0(.din(n3586), .dout(n3583));
    jdff dff_A_cENlmcPz9_0(.din(n3589), .dout(n3586));
    jdff dff_A_7wffRQjy9_0(.din(G47gat), .dout(n3589));
    jdff dff_B_Fv6m2CzD8_1(.din(n318), .dout(n3593));
    jdff dff_B_TmclbHEC8_1(.din(n3593), .dout(n3596));
    jdff dff_B_KBCDqDzO1_1(.din(n3596), .dout(n3599));
    jdff dff_B_YhorwD8j4_1(.din(n3599), .dout(n3602));
    jdff dff_B_wKH6W4uK7_1(.din(n3602), .dout(n3605));
    jdff dff_B_aokus66T8_1(.din(n3605), .dout(n3608));
    jdff dff_B_u6r39nYs8_1(.din(n3608), .dout(n3611));
    jdff dff_A_it2qwHqH0_0(.din(n3616), .dout(n3613));
    jdff dff_A_qwn3zPLH3_0(.din(n3619), .dout(n3616));
    jdff dff_A_cyDwvHrD6_0(.din(n3622), .dout(n3619));
    jdff dff_A_wHUrBUHx2_0(.din(n3625), .dout(n3622));
    jdff dff_A_tm1iovNG2_0(.din(n3628), .dout(n3625));
    jdff dff_A_fOcwSh3o6_0(.din(n3631), .dout(n3628));
    jdff dff_A_ECDtJwif4_0(.din(n3634), .dout(n3631));
    jdff dff_A_2GhpTHQo1_0(.din(n3637), .dout(n3634));
    jdff dff_A_2S4R9faL7_0(.din(n3640), .dout(n3637));
    jdff dff_A_ODmWjlRV5_0(.din(n3643), .dout(n3640));
    jdff dff_A_rd3Fba8s6_0(.din(n3646), .dout(n3643));
    jdff dff_A_tko4XCxQ2_0(.din(n3649), .dout(n3646));
    jdff dff_A_tKksQxqR6_0(.din(G60gat), .dout(n3649));
    jdff dff_A_KEyb8s4Y9_1(.din(n3655), .dout(n3652));
    jdff dff_A_U5B2XVT57_1(.din(n3658), .dout(n3655));
    jdff dff_A_tgiBVSHu4_1(.din(n3661), .dout(n3658));
    jdff dff_A_eucTybFG0_1(.din(n3664), .dout(n3661));
    jdff dff_A_dyrbwCaQ3_1(.din(n3667), .dout(n3664));
    jdff dff_A_zPHajorB1_1(.din(n3670), .dout(n3667));
    jdff dff_A_0r1rFZJN2_1(.din(n3673), .dout(n3670));
    jdff dff_A_gtyfAx5u2_1(.din(G60gat), .dout(n3673));
    jdff dff_A_lyQsZuTS8_0(.din(n3679), .dout(n3676));
    jdff dff_A_8PsZVu7s4_0(.din(n312), .dout(n3679));
    jdff dff_A_4x2ufxxD8_0(.din(n3685), .dout(n3682));
    jdff dff_A_5P6RYtYA6_0(.din(n3688), .dout(n3685));
    jdff dff_A_z7doHYr38_0(.din(n3691), .dout(n3688));
    jdff dff_A_bU20rqy65_0(.din(n3694), .dout(n3691));
    jdff dff_A_O709u4Bz7_0(.din(n3697), .dout(n3694));
    jdff dff_A_2iAQPlyp8_0(.din(n308), .dout(n3697));
    jdff dff_A_hiYXJa653_0(.din(n3703), .dout(n3700));
    jdff dff_A_ZkJX8wsO7_0(.din(n3706), .dout(n3703));
    jdff dff_A_O1gGKJgq3_0(.din(n3709), .dout(n3706));
    jdff dff_A_w1nJKGU09_0(.din(n3712), .dout(n3709));
    jdff dff_A_GsPdezS24_0(.din(n3715), .dout(n3712));
    jdff dff_A_EZTCzFBR7_0(.din(n3718), .dout(n3715));
    jdff dff_A_hAAFYBmp5_0(.din(n3721), .dout(n3718));
    jdff dff_A_kAASZgl22_0(.din(n3724), .dout(n3721));
    jdff dff_A_XCqU0mN41_0(.din(n3727), .dout(n3724));
    jdff dff_A_ay6l1FQL0_0(.din(n3730), .dout(n3727));
    jdff dff_A_doOqM7bH5_0(.din(n3733), .dout(n3730));
    jdff dff_A_Ctzd03QN7_0(.din(n3736), .dout(n3733));
    jdff dff_A_kTjO4ryG8_0(.din(G34gat), .dout(n3736));
    jdff dff_A_2Esfz2Cc2_2(.din(n3742), .dout(n3739));
    jdff dff_A_kA7UKfZ70_2(.din(n3745), .dout(n3742));
    jdff dff_A_FNMcSjCE6_2(.din(n3748), .dout(n3745));
    jdff dff_A_Sf7DTXvw4_2(.din(n3751), .dout(n3748));
    jdff dff_A_IodsmCM40_2(.din(n3754), .dout(n3751));
    jdff dff_A_OGXhtmPX5_2(.din(n3757), .dout(n3754));
    jdff dff_A_PJ5ac82i5_2(.din(n3760), .dout(n3757));
    jdff dff_A_HLRxu9hC8_2(.din(G34gat), .dout(n3760));
    jdff dff_A_pdZLw88M9_0(.din(n3766), .dout(n3763));
    jdff dff_A_3T5QZSFe4_0(.din(n3769), .dout(n3766));
    jdff dff_A_Ix1wpVIR0_0(.din(n3772), .dout(n3769));
    jdff dff_A_QAVbQ8KG3_0(.din(n3775), .dout(n3772));
    jdff dff_A_ousPHLrB5_0(.din(n3778), .dout(n3775));
    jdff dff_A_riHUICMo6_0(.din(n288), .dout(n3778));
    jdff dff_A_1BCrSjlV2_0(.din(n3784), .dout(n3781));
    jdff dff_A_ad8fcmtR1_0(.din(n3787), .dout(n3784));
    jdff dff_A_XH5Xx23o7_0(.din(n3790), .dout(n3787));
    jdff dff_A_MJcv7u0l3_0(.din(n3793), .dout(n3790));
    jdff dff_A_Klo8Z9nq0_0(.din(n3815), .dout(n3793));
    jdff dff_B_vbNPuuRj4_2(.din(n280), .dout(n3797));
    jdff dff_B_wXu0phGn4_2(.din(n3797), .dout(n3800));
    jdff dff_B_TC71sZVX0_2(.din(n3800), .dout(n3803));
    jdff dff_B_riSjZN5b5_2(.din(n3803), .dout(n3806));
    jdff dff_B_yXinODag7_2(.din(n3806), .dout(n3809));
    jdff dff_B_Qo2yRTwU3_2(.din(n3809), .dout(n3812));
    jdff dff_B_Qpnbjv8i6_2(.din(n3812), .dout(n3815));
    jdff dff_A_1jLi4RYx1_0(.din(n3820), .dout(n3817));
    jdff dff_A_hdwRdQAI2_0(.din(n3823), .dout(n3820));
    jdff dff_A_I0FAqYFk4_0(.din(n3826), .dout(n3823));
    jdff dff_A_RPQm22uG9_0(.din(n3829), .dout(n3826));
    jdff dff_A_ToZX8LuQ5_0(.din(n3832), .dout(n3829));
    jdff dff_A_Eqvtuz0k7_0(.din(n3835), .dout(n3832));
    jdff dff_A_9Iq4itu71_0(.din(n3838), .dout(n3835));
    jdff dff_A_hgpJNaHG9_0(.din(n3841), .dout(n3838));
    jdff dff_A_GEyPZXY59_0(.din(n3844), .dout(n3841));
    jdff dff_A_85mXJdqJ6_0(.din(n3847), .dout(n3844));
    jdff dff_A_XiE6s5Pe4_0(.din(n3850), .dout(n3847));
    jdff dff_A_OxhLI8F16_0(.din(n3853), .dout(n3850));
    jdff dff_A_Uf4wyVZi1_0(.din(G73gat), .dout(n3853));
    jdff dff_A_bmHSz2Tj0_1(.din(n3859), .dout(n3856));
    jdff dff_A_qlobzmpw6_1(.din(n3862), .dout(n3859));
    jdff dff_A_R441xY9b2_1(.din(n3865), .dout(n3862));
    jdff dff_A_V0yOCIhw4_1(.din(n3868), .dout(n3865));
    jdff dff_A_gGJtaM9k0_1(.din(n3871), .dout(n3868));
    jdff dff_A_bRpoo7C77_1(.din(n3874), .dout(n3871));
    jdff dff_A_0C47CxO73_1(.din(n3877), .dout(n3874));
    jdff dff_A_LFlt7WTf2_1(.din(G73gat), .dout(n3877));
    jdff dff_B_FIU4XNhX5_1(.din(n265), .dout(n3881));
    jdff dff_B_E79sbgNT4_1(.din(n3881), .dout(n3884));
    jdff dff_B_sox4Yx8h2_1(.din(n3884), .dout(n3887));
    jdff dff_B_BH8cCgRW1_1(.din(n3887), .dout(n3890));
    jdff dff_B_1PvCAizf9_1(.din(n3890), .dout(n3893));
    jdff dff_B_IY29OhhM2_1(.din(n3893), .dout(n3896));
    jdff dff_B_4aXRGgFB2_1(.din(n3896), .dout(n3899));
    jdff dff_A_Bl0vePuy3_0(.din(n3904), .dout(n3901));
    jdff dff_A_WPByknKX0_0(.din(n3907), .dout(n3904));
    jdff dff_A_psbqyxzE7_0(.din(n3910), .dout(n3907));
    jdff dff_A_vAiuKXTl7_0(.din(n3913), .dout(n3910));
    jdff dff_A_YDBVrOPt0_0(.din(n3916), .dout(n3913));
    jdff dff_A_KHOofYdl2_0(.din(n3919), .dout(n3916));
    jdff dff_A_BlT9XUv15_0(.din(n3922), .dout(n3919));
    jdff dff_A_4MmouBb57_0(.din(G99gat), .dout(n3922));
    jdff dff_A_ryZQ9wY16_1(.din(n3928), .dout(n3925));
    jdff dff_A_NzIrbV8u5_1(.din(n3931), .dout(n3928));
    jdff dff_A_NumHLs2G7_1(.din(n3934), .dout(n3931));
    jdff dff_A_mZHBZK701_1(.din(n3937), .dout(n3934));
    jdff dff_A_70pygJTa6_1(.din(n3940), .dout(n3937));
    jdff dff_A_PNlwz2hy0_1(.din(n3943), .dout(n3940));
    jdff dff_A_5DxUnceN5_1(.din(n3946), .dout(n3943));
    jdff dff_A_u0Reuen91_1(.din(n3949), .dout(n3946));
    jdff dff_A_3S0Noii19_1(.din(n3952), .dout(n3949));
    jdff dff_A_HOdmcer34_1(.din(n3955), .dout(n3952));
    jdff dff_A_Js6aPtXj6_1(.din(n3958), .dout(n3955));
    jdff dff_A_ixIbOInX5_1(.din(n3961), .dout(n3958));
    jdff dff_A_3q3Udb6f2_1(.din(G99gat), .dout(n3961));
    jdff dff_A_3WhSAtBC6_0(.din(n3967), .dout(n3964));
    jdff dff_A_C4yHK1bg7_0(.din(n3970), .dout(n3967));
    jdff dff_A_OHNi3BtC2_0(.din(n3973), .dout(n3970));
    jdff dff_A_tmvUf1fZ7_0(.din(n3976), .dout(n3973));
    jdff dff_A_vry5MGvC5_0(.din(n3979), .dout(n3976));
    jdff dff_A_FycskBfx6_0(.din(n254), .dout(n3979));
    jdff dff_A_WYcYWevu1_0(.din(n3985), .dout(n3982));
    jdff dff_A_bNclPy5R3_0(.din(n3988), .dout(n3985));
    jdff dff_A_SBDThDsY3_0(.din(n3991), .dout(n3988));
    jdff dff_A_buxUTz049_0(.din(n3994), .dout(n3991));
    jdff dff_A_QQALszhd2_0(.din(n4016), .dout(n3994));
    jdff dff_B_3SWlJP7U6_2(.din(n246), .dout(n3998));
    jdff dff_B_H7EoF3O72_2(.din(n3998), .dout(n4001));
    jdff dff_B_f6U0AA6u9_2(.din(n4001), .dout(n4004));
    jdff dff_B_jiu8K6Mv4_2(.din(n4004), .dout(n4007));
    jdff dff_B_h5wiugK65_2(.din(n4007), .dout(n4010));
    jdff dff_B_0L1AhYIW6_2(.din(n4010), .dout(n4013));
    jdff dff_B_zzOnSQo75_2(.din(n4013), .dout(n4016));
    jdff dff_A_pKoZdVtq3_0(.din(n4021), .dout(n4018));
    jdff dff_A_LBmYrF4v2_0(.din(n4024), .dout(n4021));
    jdff dff_A_vkLkEUDb0_0(.din(n4027), .dout(n4024));
    jdff dff_A_8nGOXfmL3_0(.din(n4030), .dout(n4027));
    jdff dff_A_tckeineN2_0(.din(n4033), .dout(n4030));
    jdff dff_A_V0OZ0ex87_0(.din(n4036), .dout(n4033));
    jdff dff_A_RAQ7soBi6_0(.din(n4039), .dout(n4036));
    jdff dff_A_3gY0AY0h1_0(.din(n4042), .dout(n4039));
    jdff dff_A_stDXda203_0(.din(n4045), .dout(n4042));
    jdff dff_A_4wrPObSd0_0(.din(n4048), .dout(n4045));
    jdff dff_A_inT0k7Z87_0(.din(n4051), .dout(n4048));
    jdff dff_A_5z3gmTeW9_0(.din(n4054), .dout(n4051));
    jdff dff_A_BF8gCdAp4_0(.din(G8gat), .dout(n4054));
    jdff dff_A_MGDYFj995_1(.din(n4060), .dout(n4057));
    jdff dff_A_2T4XnEqm3_1(.din(n4063), .dout(n4060));
    jdff dff_A_Gm0vMFkY0_1(.din(n4066), .dout(n4063));
    jdff dff_A_n64ETrL61_1(.din(n4069), .dout(n4066));
    jdff dff_A_s1VW2A2j8_1(.din(n4072), .dout(n4069));
    jdff dff_A_mPsWAnai9_1(.din(n4075), .dout(n4072));
    jdff dff_A_iXdroaPO2_1(.din(n4078), .dout(n4075));
    jdff dff_A_6l4mxBtJ8_1(.din(G8gat), .dout(n4078));
    jdff dff_A_ZAq4GogY7_0(.din(n4084), .dout(n4081));
    jdff dff_A_Zjd3FBVm9_0(.din(n4087), .dout(n4084));
    jdff dff_A_hP8e5VEY4_0(.din(n4090), .dout(n4087));
    jdff dff_A_E5jsua8o5_0(.din(n4093), .dout(n4090));
    jdff dff_A_x77Iu3pY1_0(.din(n4096), .dout(n4093));
    jdff dff_A_F1VAy6oj4_0(.din(n239), .dout(n4096));
    jdff dff_B_1g27YgFr7_1(.din(n165), .dout(n4100));
    jdff dff_B_7jHgBMXL3_1(.din(n183), .dout(n4103));
    jdff dff_A_YS5WvG4O8_0(.din(n4108), .dout(n4105));
    jdff dff_A_RdscfmSd6_0(.din(n4111), .dout(n4108));
    jdff dff_A_vs4Yte5a6_0(.din(n4114), .dout(n4111));
    jdff dff_A_McmLrzke5_0(.din(n4117), .dout(n4114));
    jdff dff_A_TTdqR00b8_0(.din(n4120), .dout(n4117));
    jdff dff_A_vcoSxdJH7_0(.din(n211), .dout(n4120));
    jdff dff_A_FNBBFI7k1_0(.din(n4126), .dout(n4123));
    jdff dff_A_egyvezmP1_0(.din(n4129), .dout(n4126));
    jdff dff_A_KAqRUqc41_0(.din(n4132), .dout(n4129));
    jdff dff_A_tNomMc159_0(.din(n4135), .dout(n4132));
    jdff dff_A_xxDRcru73_0(.din(n4138), .dout(n4135));
    jdff dff_A_t6pyZeN27_0(.din(n193), .dout(n4138));
    jdff dff_A_0tDbL01y9_0(.din(n4144), .dout(n4141));
    jdff dff_A_QgsUMgbR2_0(.din(n4147), .dout(n4144));
    jdff dff_A_zSvERz9r7_0(.din(n4150), .dout(n4147));
    jdff dff_A_D8HQEZDm7_0(.din(n4153), .dout(n4150));
    jdff dff_A_VUMppq5o2_0(.din(n4156), .dout(n4153));
    jdff dff_A_PftCV0974_0(.din(n186), .dout(n4156));
    jdff dff_A_H77QyUzX6_0(.din(n4162), .dout(n4159));
    jdff dff_A_ikqDVpKe9_0(.din(n4165), .dout(n4162));
    jdff dff_A_6IvXc7H93_0(.din(n4168), .dout(n4165));
    jdff dff_A_IEeZPfcm7_0(.din(n4171), .dout(n4168));
    jdff dff_A_E3m0gHHM1_0(.din(n4174), .dout(n4171));
    jdff dff_A_0iX5VOvF3_0(.din(n175), .dout(n4174));
    jdff dff_A_0KSjwQtd3_0(.din(n4180), .dout(n4177));
    jdff dff_A_tJBtmbww6_0(.din(n4183), .dout(n4180));
    jdff dff_A_KIGRHkPL2_0(.din(n4186), .dout(n4183));
    jdff dff_A_3oa89vUu6_0(.din(n172), .dout(n4186));
    jdff dff_A_CAjglNfV7_0(.din(n4192), .dout(n4189));
    jdff dff_A_OU2Z0wSZ9_0(.din(n4195), .dout(n4192));
    jdff dff_A_LbP9gmM75_0(.din(n4198), .dout(n4195));
    jdff dff_A_qKygx8oj3_0(.din(n4201), .dout(n4198));
    jdff dff_A_H49QXB351_0(.din(n4204), .dout(n4201));
    jdff dff_A_DQdR1sTx9_0(.din(n168), .dout(n4204));
    jdff dff_A_0WKc5XU48_0(.din(n4210), .dout(n4207));
    jdff dff_A_1eDK6lYR9_0(.din(n4213), .dout(n4210));
    jdff dff_A_b8Ik8HGI4_0(.din(n4216), .dout(n4213));
    jdff dff_A_d4CkhFFo4_0(.din(n4219), .dout(n4216));
    jdff dff_A_Km5hpih89_0(.din(n4222), .dout(n4219));
    jdff dff_A_p5hPemGS8_0(.din(n153), .dout(n4222));
    jdff dff_A_wgydJpYc2_0(.din(n4228), .dout(n4225));
    jdff dff_A_Fevppzgi7_0(.din(n4231), .dout(n4228));
    jdff dff_A_4rThsRKZ8_0(.din(n4234), .dout(n4231));
    jdff dff_A_mjNe2c9q6_0(.din(n150), .dout(n4234));
    jdff dff_A_UN8sB5N10_0(.din(n4240), .dout(n4237));
    jdff dff_A_cQUYckR48_0(.din(n4243), .dout(n4240));
    jdff dff_A_vyhN0RL21_0(.din(n4246), .dout(n4243));
    jdff dff_A_XmSAc9Y30_0(.din(n4249), .dout(n4246));
    jdff dff_A_nPf3tF7K5_0(.din(n4252), .dout(n4249));
    jdff dff_A_im35mc7u0_0(.din(n146), .dout(n4252));
    jdff dff_A_ibEiz88q1_0(.din(n4258), .dout(n4255));
    jdff dff_A_NQDn57kM7_0(.din(n4261), .dout(n4258));
    jdff dff_A_k8AqYqB49_0(.din(n4264), .dout(n4261));
    jdff dff_A_UEpzuz7S1_0(.din(n4267), .dout(n4264));
    jdff dff_A_9tiFhrMz9_0(.din(n4289), .dout(n4267));
    jdff dff_B_N7AGX4IP8_2(.din(n140), .dout(n4271));
    jdff dff_B_6G06KosA9_2(.din(n4271), .dout(n4274));
    jdff dff_B_KOAIJrsW4_2(.din(n4274), .dout(n4277));
    jdff dff_B_B4a7me5l3_2(.din(n4277), .dout(n4280));
    jdff dff_B_fHVpo0DQ5_2(.din(n4280), .dout(n4283));
    jdff dff_B_YCdv7NHY3_2(.din(n4283), .dout(n4286));
    jdff dff_B_R69DaiPJ4_2(.din(n4286), .dout(n4289));
    jdff dff_A_68eKiuOq4_0(.din(n4294), .dout(n4291));
    jdff dff_A_7s7x76Wm0_0(.din(n4297), .dout(n4294));
    jdff dff_A_5VbRwkNE8_0(.din(n4300), .dout(n4297));
    jdff dff_A_DyW161X97_0(.din(n4303), .dout(n4300));
    jdff dff_A_W2PdFSHR5_0(.din(n4306), .dout(n4303));
    jdff dff_A_D6w4JkDp7_0(.din(n4309), .dout(n4306));
    jdff dff_A_8JH5ryuG1_0(.din(n4312), .dout(n4309));
    jdff dff_A_bNWg9gOY3_0(.din(n4315), .dout(n4312));
    jdff dff_A_5LwtncGv2_0(.din(n4318), .dout(n4315));
    jdff dff_A_SY7nT9p57_0(.din(n4321), .dout(n4318));
    jdff dff_A_qDDjToK53_0(.din(n4324), .dout(n4321));
    jdff dff_A_MEWjSqDL2_0(.din(n4327), .dout(n4324));
    jdff dff_A_y0ynk3B09_0(.din(G112gat), .dout(n4327));
    jdff dff_A_aPcuxAQt9_1(.din(n4333), .dout(n4330));
    jdff dff_A_j4NiqdiA4_1(.din(n4336), .dout(n4333));
    jdff dff_A_ggz7T9v59_1(.din(n4339), .dout(n4336));
    jdff dff_A_QceUSftn8_1(.din(n4342), .dout(n4339));
    jdff dff_A_q5xRitIL5_1(.din(n4345), .dout(n4342));
    jdff dff_A_tXyKoq2u0_1(.din(n4348), .dout(n4345));
    jdff dff_A_PidPrwjK1_1(.din(n4351), .dout(n4348));
    jdff dff_A_nAPqZLqT6_1(.din(G112gat), .dout(n4351));
    jdff dff_A_gJ6hF6OQ1_1(.din(n4357), .dout(n4354));
    jdff dff_A_SqMnunAP0_1(.din(n4360), .dout(n4357));
    jdff dff_A_x8GueNsS5_1(.din(n4363), .dout(n4360));
    jdff dff_A_69bqsicp0_1(.din(n4366), .dout(n4363));
    jdff dff_A_VEwuRhUd5_1(.din(n4369), .dout(n4366));
    jdff dff_A_8uzRIjdi1_1(.din(n403), .dout(n4369));
    jdff dff_B_psk07u3V0_1(.din(n71), .dout(n4373));
    jdff dff_B_oqycvCM21_1(.din(n89), .dout(n4376));
    jdff dff_A_MMSOLrkf9_0(.din(n4381), .dout(n4378));
    jdff dff_A_EmbrQ3OK4_0(.din(n4384), .dout(n4381));
    jdff dff_A_5EwA2DpY9_0(.din(n4387), .dout(n4384));
    jdff dff_A_sSsn89L83_0(.din(n4390), .dout(n4387));
    jdff dff_A_5ABIk3ha6_0(.din(n4393), .dout(n4390));
    jdff dff_A_Rd3Iqsut7_0(.din(n4396), .dout(n4393));
    jdff dff_A_B0KcFS5N3_0(.din(G4gat), .dout(n4396));
    jdff dff_A_OXR4KdRt3_2(.din(G4gat), .dout(n4399));
    jdff dff_A_HGZVjoyq2_0(.din(n4405), .dout(n4402));
    jdff dff_A_y3JgxNnQ8_0(.din(n4408), .dout(n4405));
    jdff dff_A_xSbHDy8M1_0(.din(n4411), .dout(n4408));
    jdff dff_A_Zh6Zzmpx9_0(.din(n4414), .dout(n4411));
    jdff dff_A_GHmMaPQz1_0(.din(n117), .dout(n4414));
    jdff dff_A_zxg6pJ4q5_0(.din(n4420), .dout(n4417));
    jdff dff_A_KlkLvP1s6_0(.din(n4423), .dout(n4420));
    jdff dff_A_l6Ex0cdx4_0(.din(n4426), .dout(n4423));
    jdff dff_A_wQCdnG0t0_0(.din(n4429), .dout(n4426));
    jdff dff_A_unlN3uPJ9_0(.din(n4432), .dout(n4429));
    jdff dff_A_qMJdKDQo4_0(.din(G1gat), .dout(n4432));
    jdff dff_A_A24A1gXq5_1(.din(G1gat), .dout(n4435));
    jdff dff_A_poMtGWKM2_0(.din(n4441), .dout(n4438));
    jdff dff_A_BGrAfOEQ2_0(.din(n4444), .dout(n4441));
    jdff dff_A_KOnpoR7X3_0(.din(n4447), .dout(n4444));
    jdff dff_A_xyIwAmPi0_0(.din(n4450), .dout(n4447));
    jdff dff_A_0ee1nJSj0_0(.din(n110), .dout(n4450));
    jdff dff_A_mXeuhKAh9_0(.din(n4456), .dout(n4453));
    jdff dff_A_WiEggLot0_0(.din(n4459), .dout(n4456));
    jdff dff_A_k2SMsEB40_0(.din(n4462), .dout(n4459));
    jdff dff_A_Pdt8fVrR5_0(.din(n4465), .dout(n4462));
    jdff dff_A_Xslwsn9A7_0(.din(n4468), .dout(n4465));
    jdff dff_A_VTHH7CAn5_0(.din(G89gat), .dout(n4468));
    jdff dff_A_wx4vqfXc1_1(.din(G89gat), .dout(n4471));
    jdff dff_A_OtuWHIYh9_0(.din(n4477), .dout(n4474));
    jdff dff_A_CQZXVABP2_0(.din(n4480), .dout(n4477));
    jdff dff_A_t8svVLG17_0(.din(n4483), .dout(n4480));
    jdff dff_A_4DJWQcyM2_0(.din(n4486), .dout(n4483));
    jdff dff_A_Gj9lJwna2_0(.din(n4489), .dout(n4486));
    jdff dff_A_fsi7MOdP6_0(.din(n4492), .dout(n4489));
    jdff dff_A_MpS27uXT9_0(.din(G56gat), .dout(n4492));
    jdff dff_A_LTw6E6Ql5_2(.din(G56gat), .dout(n4495));
    jdff dff_A_b7HwALh75_0(.din(n4501), .dout(n4498));
    jdff dff_A_tUTfemSi8_0(.din(n4504), .dout(n4501));
    jdff dff_A_1qWtbnpy2_0(.din(n4507), .dout(n4504));
    jdff dff_A_ZnTlYI2p8_0(.din(n4510), .dout(n4507));
    jdff dff_A_bmwWrFaJ6_0(.din(n99), .dout(n4510));
    jdff dff_A_SbywBC6r8_0(.din(n4516), .dout(n4513));
    jdff dff_A_2oG41Q1J2_0(.din(n4519), .dout(n4516));
    jdff dff_A_368eFpuS7_0(.din(n4522), .dout(n4519));
    jdff dff_A_EeKppYKU2_0(.din(n4525), .dout(n4522));
    jdff dff_A_e8Vraddr0_0(.din(n4528), .dout(n4525));
    jdff dff_A_XquBIlvv5_0(.din(G50gat), .dout(n4528));
    jdff dff_A_o0bLKkPz9_1(.din(G50gat), .dout(n4531));
    jdff dff_A_sxEaZZfL4_0(.din(n4537), .dout(n4534));
    jdff dff_A_3uv68hd12_0(.din(n4540), .dout(n4537));
    jdff dff_A_tMi8ojkN1_0(.din(n4543), .dout(n4540));
    jdff dff_A_gOAH3kGN4_0(.din(n4546), .dout(n4543));
    jdff dff_A_1NtzMFup5_0(.din(n4549), .dout(n4546));
    jdff dff_A_saW5UnnJ7_0(.din(n4552), .dout(n4549));
    jdff dff_A_Z5ttAmgn2_0(.din(G108gat), .dout(n4552));
    jdff dff_A_WgCxUncS6_2(.din(G108gat), .dout(n4555));
    jdff dff_A_zpHSg7Vy4_0(.din(n4561), .dout(n4558));
    jdff dff_A_LL1rQsT87_0(.din(n4564), .dout(n4561));
    jdff dff_A_KVTmalWt2_0(.din(n4567), .dout(n4564));
    jdff dff_A_5OMAOq8G4_0(.din(n4570), .dout(n4567));
    jdff dff_A_UoMNT9Qa5_0(.din(n92), .dout(n4570));
    jdff dff_A_C4ohPfNl4_0(.din(n4576), .dout(n4573));
    jdff dff_A_iUHYDX1B0_0(.din(n4579), .dout(n4576));
    jdff dff_A_PWJzbRI75_0(.din(n4582), .dout(n4579));
    jdff dff_A_2ulqc1dc6_0(.din(n4585), .dout(n4582));
    jdff dff_A_KjHMfl831_0(.din(n4588), .dout(n4585));
    jdff dff_A_VjTQ0GMX3_0(.din(G102gat), .dout(n4588));
    jdff dff_A_uTzSJXu04_1(.din(G102gat), .dout(n4591));
    jdff dff_A_fBEA9jxP0_0(.din(n4597), .dout(n4594));
    jdff dff_A_OLfa3rfG0_0(.din(n4600), .dout(n4597));
endmodule

