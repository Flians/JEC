/*

c6288:
	jxor: 446
	jspl: 940
	jspl3: 260
	jnot: 330
	jdff: 8448
	jand: 683
	jor: 331

Summary:
	jxor: 446
	jspl: 940
	jspl3: 260
	jnot: 330
	jdff: 8448
	jand: 683
	jor: 331
*/

module c6288(gclk, G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat, G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat, G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat, G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat, G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat, G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat, G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat, G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat, G6270gat, G6280gat, G6287gat, G6288gat);
	input gclk;
	input G1gat;
	input G18gat;
	input G35gat;
	input G52gat;
	input G69gat;
	input G86gat;
	input G103gat;
	input G120gat;
	input G137gat;
	input G154gat;
	input G171gat;
	input G188gat;
	input G205gat;
	input G222gat;
	input G239gat;
	input G256gat;
	input G273gat;
	input G290gat;
	input G307gat;
	input G324gat;
	input G341gat;
	input G358gat;
	input G375gat;
	input G392gat;
	input G409gat;
	input G426gat;
	input G443gat;
	input G460gat;
	input G477gat;
	input G494gat;
	input G511gat;
	input G528gat;
	output G545gat;
	output G1581gat;
	output G1901gat;
	output G2223gat;
	output G2548gat;
	output G2877gat;
	output G3211gat;
	output G3552gat;
	output G3895gat;
	output G4241gat;
	output G4591gat;
	output G4946gat;
	output G5308gat;
	output G5672gat;
	output G5971gat;
	output G6123gat;
	output G6150gat;
	output G6160gat;
	output G6170gat;
	output G6180gat;
	output G6190gat;
	output G6200gat;
	output G6210gat;
	output G6220gat;
	output G6230gat;
	output G6240gat;
	output G6250gat;
	output G6260gat;
	output G6270gat;
	output G6280gat;
	output G6287gat;
	output G6288gat;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n70;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1667;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1684;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1690;
	wire n1691;
	wire n1692;
	wire n1693;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1707;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire n1718;
	wire n1719;
	wire n1720;
	wire n1722;
	wire n1723;
	wire n1724;
	wire n1725;
	wire n1726;
	wire n1727;
	wire n1728;
	wire n1729;
	wire n1730;
	wire n1731;
	wire n1732;
	wire n1733;
	wire n1734;
	wire n1735;
	wire n1736;
	wire n1737;
	wire n1738;
	wire n1739;
	wire n1740;
	wire n1741;
	wire n1742;
	wire n1743;
	wire n1744;
	wire n1745;
	wire n1746;
	wire n1747;
	wire n1748;
	wire n1749;
	wire n1750;
	wire n1751;
	wire n1752;
	wire n1753;
	wire n1754;
	wire n1755;
	wire n1756;
	wire n1757;
	wire n1758;
	wire n1760;
	wire n1761;
	wire n1762;
	wire n1763;
	wire n1764;
	wire n1765;
	wire n1766;
	wire n1767;
	wire n1768;
	wire n1769;
	wire n1770;
	wire n1771;
	wire n1772;
	wire n1773;
	wire n1774;
	wire n1775;
	wire n1776;
	wire n1777;
	wire n1778;
	wire n1779;
	wire n1780;
	wire n1781;
	wire n1782;
	wire n1783;
	wire n1784;
	wire n1785;
	wire n1786;
	wire n1787;
	wire n1788;
	wire n1789;
	wire n1790;
	wire n1791;
	wire n1793;
	wire n1794;
	wire n1795;
	wire n1796;
	wire n1797;
	wire n1798;
	wire n1799;
	wire n1800;
	wire n1801;
	wire n1802;
	wire n1803;
	wire n1804;
	wire n1805;
	wire n1806;
	wire n1807;
	wire n1808;
	wire n1809;
	wire n1810;
	wire n1811;
	wire n1812;
	wire n1813;
	wire n1814;
	wire n1815;
	wire n1816;
	wire n1817;
	wire n1819;
	wire n1820;
	wire n1821;
	wire n1822;
	wire n1823;
	wire n1824;
	wire n1825;
	wire n1826;
	wire n1827;
	wire n1828;
	wire n1829;
	wire n1830;
	wire n1831;
	wire n1832;
	wire n1833;
	wire n1834;
	wire n1835;
	wire n1836;
	wire n1838;
	wire n1839;
	wire n1840;
	wire n1841;
	wire n1842;
	wire n1843;
	wire n1844;
	wire n1845;
	wire n1846;
	wire n1847;
	wire n1848;
	wire n1849;
	wire n1850;
	wire n1851;
	wire[2:0] w_G1gat_0;
	wire[2:0] w_G1gat_1;
	wire[2:0] w_G1gat_2;
	wire[2:0] w_G1gat_3;
	wire[2:0] w_G1gat_4;
	wire[2:0] w_G1gat_5;
	wire[2:0] w_G1gat_6;
	wire[1:0] w_G1gat_7;
	wire[2:0] w_G18gat_0;
	wire[2:0] w_G18gat_1;
	wire[2:0] w_G18gat_2;
	wire[2:0] w_G18gat_3;
	wire[2:0] w_G18gat_4;
	wire[2:0] w_G18gat_5;
	wire[2:0] w_G18gat_6;
	wire[2:0] w_G18gat_7;
	wire[2:0] w_G35gat_0;
	wire[2:0] w_G35gat_1;
	wire[2:0] w_G35gat_2;
	wire[2:0] w_G35gat_3;
	wire[2:0] w_G35gat_4;
	wire[2:0] w_G35gat_5;
	wire[2:0] w_G35gat_6;
	wire[2:0] w_G35gat_7;
	wire[2:0] w_G52gat_0;
	wire[2:0] w_G52gat_1;
	wire[2:0] w_G52gat_2;
	wire[2:0] w_G52gat_3;
	wire[2:0] w_G52gat_4;
	wire[2:0] w_G52gat_5;
	wire[2:0] w_G52gat_6;
	wire[2:0] w_G52gat_7;
	wire[2:0] w_G69gat_0;
	wire[2:0] w_G69gat_1;
	wire[2:0] w_G69gat_2;
	wire[2:0] w_G69gat_3;
	wire[2:0] w_G69gat_4;
	wire[2:0] w_G69gat_5;
	wire[2:0] w_G69gat_6;
	wire[1:0] w_G69gat_7;
	wire[2:0] w_G86gat_0;
	wire[2:0] w_G86gat_1;
	wire[2:0] w_G86gat_2;
	wire[2:0] w_G86gat_3;
	wire[2:0] w_G86gat_4;
	wire[2:0] w_G86gat_5;
	wire[2:0] w_G86gat_6;
	wire[1:0] w_G86gat_7;
	wire[2:0] w_G103gat_0;
	wire[2:0] w_G103gat_1;
	wire[2:0] w_G103gat_2;
	wire[2:0] w_G103gat_3;
	wire[2:0] w_G103gat_4;
	wire[2:0] w_G103gat_5;
	wire[2:0] w_G103gat_6;
	wire[1:0] w_G103gat_7;
	wire[2:0] w_G120gat_0;
	wire[2:0] w_G120gat_1;
	wire[2:0] w_G120gat_2;
	wire[2:0] w_G120gat_3;
	wire[2:0] w_G120gat_4;
	wire[2:0] w_G120gat_5;
	wire[2:0] w_G120gat_6;
	wire[1:0] w_G120gat_7;
	wire[2:0] w_G137gat_0;
	wire[2:0] w_G137gat_1;
	wire[2:0] w_G137gat_2;
	wire[2:0] w_G137gat_3;
	wire[2:0] w_G137gat_4;
	wire[2:0] w_G137gat_5;
	wire[2:0] w_G137gat_6;
	wire[1:0] w_G137gat_7;
	wire[2:0] w_G154gat_0;
	wire[2:0] w_G154gat_1;
	wire[2:0] w_G154gat_2;
	wire[2:0] w_G154gat_3;
	wire[2:0] w_G154gat_4;
	wire[2:0] w_G154gat_5;
	wire[2:0] w_G154gat_6;
	wire[1:0] w_G154gat_7;
	wire[2:0] w_G171gat_0;
	wire[2:0] w_G171gat_1;
	wire[2:0] w_G171gat_2;
	wire[2:0] w_G171gat_3;
	wire[2:0] w_G171gat_4;
	wire[2:0] w_G171gat_5;
	wire[2:0] w_G171gat_6;
	wire[1:0] w_G171gat_7;
	wire[2:0] w_G188gat_0;
	wire[2:0] w_G188gat_1;
	wire[2:0] w_G188gat_2;
	wire[2:0] w_G188gat_3;
	wire[2:0] w_G188gat_4;
	wire[2:0] w_G188gat_5;
	wire[2:0] w_G188gat_6;
	wire[1:0] w_G188gat_7;
	wire[2:0] w_G205gat_0;
	wire[2:0] w_G205gat_1;
	wire[2:0] w_G205gat_2;
	wire[2:0] w_G205gat_3;
	wire[2:0] w_G205gat_4;
	wire[2:0] w_G205gat_5;
	wire[2:0] w_G205gat_6;
	wire[1:0] w_G205gat_7;
	wire[2:0] w_G222gat_0;
	wire[2:0] w_G222gat_1;
	wire[2:0] w_G222gat_2;
	wire[2:0] w_G222gat_3;
	wire[2:0] w_G222gat_4;
	wire[2:0] w_G222gat_5;
	wire[2:0] w_G222gat_6;
	wire[1:0] w_G222gat_7;
	wire[2:0] w_G239gat_0;
	wire[2:0] w_G239gat_1;
	wire[2:0] w_G239gat_2;
	wire[2:0] w_G239gat_3;
	wire[2:0] w_G239gat_4;
	wire[2:0] w_G239gat_5;
	wire[2:0] w_G239gat_6;
	wire[1:0] w_G239gat_7;
	wire[2:0] w_G256gat_0;
	wire[2:0] w_G256gat_1;
	wire[2:0] w_G256gat_2;
	wire[2:0] w_G256gat_3;
	wire[2:0] w_G256gat_4;
	wire[2:0] w_G256gat_5;
	wire[2:0] w_G256gat_6;
	wire[1:0] w_G256gat_7;
	wire[2:0] w_G273gat_0;
	wire[2:0] w_G273gat_1;
	wire[2:0] w_G273gat_2;
	wire[2:0] w_G273gat_3;
	wire[2:0] w_G273gat_4;
	wire[2:0] w_G273gat_5;
	wire[2:0] w_G273gat_6;
	wire[2:0] w_G273gat_7;
	wire[2:0] w_G290gat_0;
	wire[2:0] w_G290gat_1;
	wire[2:0] w_G290gat_2;
	wire[2:0] w_G290gat_3;
	wire[2:0] w_G290gat_4;
	wire[2:0] w_G290gat_5;
	wire[2:0] w_G290gat_6;
	wire[2:0] w_G290gat_7;
	wire[2:0] w_G307gat_0;
	wire[2:0] w_G307gat_1;
	wire[2:0] w_G307gat_2;
	wire[2:0] w_G307gat_3;
	wire[2:0] w_G307gat_4;
	wire[2:0] w_G307gat_5;
	wire[2:0] w_G307gat_6;
	wire[2:0] w_G307gat_7;
	wire[2:0] w_G324gat_0;
	wire[2:0] w_G324gat_1;
	wire[2:0] w_G324gat_2;
	wire[2:0] w_G324gat_3;
	wire[2:0] w_G324gat_4;
	wire[2:0] w_G324gat_5;
	wire[2:0] w_G324gat_6;
	wire[1:0] w_G324gat_7;
	wire[2:0] w_G341gat_0;
	wire[2:0] w_G341gat_1;
	wire[2:0] w_G341gat_2;
	wire[2:0] w_G341gat_3;
	wire[2:0] w_G341gat_4;
	wire[2:0] w_G341gat_5;
	wire[2:0] w_G341gat_6;
	wire[1:0] w_G341gat_7;
	wire[2:0] w_G358gat_0;
	wire[2:0] w_G358gat_1;
	wire[2:0] w_G358gat_2;
	wire[2:0] w_G358gat_3;
	wire[2:0] w_G358gat_4;
	wire[2:0] w_G358gat_5;
	wire[2:0] w_G358gat_6;
	wire[1:0] w_G358gat_7;
	wire[2:0] w_G375gat_0;
	wire[2:0] w_G375gat_1;
	wire[2:0] w_G375gat_2;
	wire[2:0] w_G375gat_3;
	wire[2:0] w_G375gat_4;
	wire[2:0] w_G375gat_5;
	wire[2:0] w_G375gat_6;
	wire[1:0] w_G375gat_7;
	wire[2:0] w_G392gat_0;
	wire[2:0] w_G392gat_1;
	wire[2:0] w_G392gat_2;
	wire[2:0] w_G392gat_3;
	wire[2:0] w_G392gat_4;
	wire[2:0] w_G392gat_5;
	wire[2:0] w_G392gat_6;
	wire[1:0] w_G392gat_7;
	wire[2:0] w_G409gat_0;
	wire[2:0] w_G409gat_1;
	wire[2:0] w_G409gat_2;
	wire[2:0] w_G409gat_3;
	wire[2:0] w_G409gat_4;
	wire[2:0] w_G409gat_5;
	wire[2:0] w_G409gat_6;
	wire[1:0] w_G409gat_7;
	wire[2:0] w_G426gat_0;
	wire[2:0] w_G426gat_1;
	wire[2:0] w_G426gat_2;
	wire[2:0] w_G426gat_3;
	wire[2:0] w_G426gat_4;
	wire[2:0] w_G426gat_5;
	wire[2:0] w_G426gat_6;
	wire[1:0] w_G426gat_7;
	wire[2:0] w_G443gat_0;
	wire[2:0] w_G443gat_1;
	wire[2:0] w_G443gat_2;
	wire[2:0] w_G443gat_3;
	wire[2:0] w_G443gat_4;
	wire[2:0] w_G443gat_5;
	wire[2:0] w_G443gat_6;
	wire[1:0] w_G443gat_7;
	wire[2:0] w_G460gat_0;
	wire[2:0] w_G460gat_1;
	wire[2:0] w_G460gat_2;
	wire[2:0] w_G460gat_3;
	wire[2:0] w_G460gat_4;
	wire[2:0] w_G460gat_5;
	wire[2:0] w_G460gat_6;
	wire[1:0] w_G460gat_7;
	wire[2:0] w_G477gat_0;
	wire[2:0] w_G477gat_1;
	wire[2:0] w_G477gat_2;
	wire[2:0] w_G477gat_3;
	wire[2:0] w_G477gat_4;
	wire[2:0] w_G477gat_5;
	wire[2:0] w_G477gat_6;
	wire[1:0] w_G477gat_7;
	wire[2:0] w_G494gat_0;
	wire[2:0] w_G494gat_1;
	wire[2:0] w_G494gat_2;
	wire[2:0] w_G494gat_3;
	wire[2:0] w_G494gat_4;
	wire[2:0] w_G494gat_5;
	wire[2:0] w_G494gat_6;
	wire[1:0] w_G494gat_7;
	wire[2:0] w_G511gat_0;
	wire[2:0] w_G511gat_1;
	wire[2:0] w_G511gat_2;
	wire[2:0] w_G511gat_3;
	wire[2:0] w_G511gat_4;
	wire[2:0] w_G511gat_5;
	wire[2:0] w_G511gat_6;
	wire[1:0] w_G511gat_7;
	wire[2:0] w_G528gat_0;
	wire[2:0] w_G528gat_1;
	wire[2:0] w_G528gat_2;
	wire[2:0] w_G528gat_3;
	wire[2:0] w_G528gat_4;
	wire[2:0] w_G528gat_5;
	wire[2:0] w_G528gat_6;
	wire[1:0] w_G528gat_7;
	wire w_G545gat_0;
	wire G545gat_fa_;
	wire[1:0] w_n65_0;
	wire[1:0] w_n69_0;
	wire[1:0] w_n70_0;
	wire[1:0] w_n72_0;
	wire[1:0] w_n75_0;
	wire[1:0] w_n77_0;
	wire[1:0] w_n78_0;
	wire[1:0] w_n81_0;
	wire[2:0] w_n82_0;
	wire[1:0] w_n82_1;
	wire[1:0] w_n84_0;
	wire[1:0] w_n85_0;
	wire[1:0] w_n87_0;
	wire[1:0] w_n89_0;
	wire[1:0] w_n93_0;
	wire[1:0] w_n94_0;
	wire[1:0] w_n96_0;
	wire[1:0] w_n99_0;
	wire[2:0] w_n100_0;
	wire[1:0] w_n100_1;
	wire[2:0] w_n101_0;
	wire[1:0] w_n103_0;
	wire[1:0] w_n104_0;
	wire[1:0] w_n107_0;
	wire[1:0] w_n108_0;
	wire[1:0] w_n110_0;
	wire[1:0] w_n115_0;
	wire[1:0] w_n116_0;
	wire[2:0] w_n126_0;
	wire[1:0] w_n128_0;
	wire[1:0] w_n129_0;
	wire[1:0] w_n130_0;
	wire[1:0] w_n131_0;
	wire[2:0] w_n132_0;
	wire[2:0] w_n133_0;
	wire[1:0] w_n138_0;
	wire[1:0] w_n139_0;
	wire[1:0] w_n140_0;
	wire[1:0] w_n142_0;
	wire[1:0] w_n143_0;
	wire[1:0] w_n145_0;
	wire[1:0] w_n150_0;
	wire[1:0] w_n151_0;
	wire[2:0] w_n156_0;
	wire[1:0] w_n158_0;
	wire[1:0] w_n163_0;
	wire[1:0] w_n165_0;
	wire[1:0] w_n166_0;
	wire[1:0] w_n168_0;
	wire[2:0] w_n169_0;
	wire[1:0] w_n170_0;
	wire[1:0] w_n172_0;
	wire[1:0] w_n174_0;
	wire[1:0] w_n175_0;
	wire[1:0] w_n176_0;
	wire[1:0] w_n177_0;
	wire[1:0] w_n178_0;
	wire[1:0] w_n180_0;
	wire[1:0] w_n181_0;
	wire[1:0] w_n183_0;
	wire[1:0] w_n188_0;
	wire[1:0] w_n189_0;
	wire[2:0] w_n194_0;
	wire[1:0] w_n196_0;
	wire[1:0] w_n199_0;
	wire[1:0] w_n201_0;
	wire[1:0] w_n204_0;
	wire[1:0] w_n206_0;
	wire[1:0] w_n207_0;
	wire[1:0] w_n209_0;
	wire[2:0] w_n210_0;
	wire[1:0] w_n210_1;
	wire[1:0] w_n213_0;
	wire[1:0] w_n215_0;
	wire[1:0] w_n216_0;
	wire[1:0] w_n217_0;
	wire[1:0] w_n218_0;
	wire[1:0] w_n219_0;
	wire[1:0] w_n220_0;
	wire[1:0] w_n221_0;
	wire[1:0] w_n223_0;
	wire[1:0] w_n224_0;
	wire[1:0] w_n226_0;
	wire[1:0] w_n231_0;
	wire[1:0] w_n232_0;
	wire[2:0] w_n237_0;
	wire[1:0] w_n239_0;
	wire[1:0] w_n242_0;
	wire[1:0] w_n244_0;
	wire[1:0] w_n247_0;
	wire[1:0] w_n249_0;
	wire[1:0] w_n252_0;
	wire[1:0] w_n254_0;
	wire[1:0] w_n255_0;
	wire[1:0] w_n257_0;
	wire[2:0] w_n258_0;
	wire[1:0] w_n259_0;
	wire[1:0] w_n261_0;
	wire[1:0] w_n264_0;
	wire[1:0] w_n265_0;
	wire[1:0] w_n266_0;
	wire[1:0] w_n267_0;
	wire[1:0] w_n268_0;
	wire[1:0] w_n269_0;
	wire[1:0] w_n270_0;
	wire[1:0] w_n271_0;
	wire[1:0] w_n272_0;
	wire[1:0] w_n274_0;
	wire[1:0] w_n275_0;
	wire[1:0] w_n277_0;
	wire[1:0] w_n282_0;
	wire[1:0] w_n283_0;
	wire[2:0] w_n288_0;
	wire[1:0] w_n290_0;
	wire[1:0] w_n293_0;
	wire[1:0] w_n295_0;
	wire[1:0] w_n298_0;
	wire[1:0] w_n300_0;
	wire[1:0] w_n303_0;
	wire[1:0] w_n305_0;
	wire[1:0] w_n308_0;
	wire[1:0] w_n310_0;
	wire[1:0] w_n311_0;
	wire[1:0] w_n313_0;
	wire[2:0] w_n314_0;
	wire[1:0] w_n315_0;
	wire[1:0] w_n317_0;
	wire[1:0] w_n320_0;
	wire[1:0] w_n321_0;
	wire[1:0] w_n322_0;
	wire[1:0] w_n323_0;
	wire[1:0] w_n324_0;
	wire[1:0] w_n325_0;
	wire[1:0] w_n326_0;
	wire[1:0] w_n327_0;
	wire[1:0] w_n328_0;
	wire[1:0] w_n329_0;
	wire[1:0] w_n330_0;
	wire[1:0] w_n332_0;
	wire[1:0] w_n333_0;
	wire[1:0] w_n335_0;
	wire[1:0] w_n340_0;
	wire[1:0] w_n341_0;
	wire[2:0] w_n346_0;
	wire[1:0] w_n348_0;
	wire[1:0] w_n351_0;
	wire[1:0] w_n353_0;
	wire[1:0] w_n356_0;
	wire[1:0] w_n358_0;
	wire[1:0] w_n361_0;
	wire[1:0] w_n363_0;
	wire[1:0] w_n366_0;
	wire[1:0] w_n368_0;
	wire[1:0] w_n371_0;
	wire[1:0] w_n372_0;
	wire[1:0] w_n373_0;
	wire[1:0] w_n375_0;
	wire[2:0] w_n376_0;
	wire[1:0] w_n377_0;
	wire[1:0] w_n380_0;
	wire[1:0] w_n382_0;
	wire[1:0] w_n383_0;
	wire[1:0] w_n384_0;
	wire[1:0] w_n385_0;
	wire[1:0] w_n386_0;
	wire[1:0] w_n387_0;
	wire[1:0] w_n388_0;
	wire[1:0] w_n389_0;
	wire[1:0] w_n390_0;
	wire[1:0] w_n391_0;
	wire[1:0] w_n392_0;
	wire[1:0] w_n393_0;
	wire[1:0] w_n394_0;
	wire[1:0] w_n396_0;
	wire[1:0] w_n397_0;
	wire[1:0] w_n399_0;
	wire[1:0] w_n404_0;
	wire[1:0] w_n405_0;
	wire[2:0] w_n410_0;
	wire[1:0] w_n412_0;
	wire[1:0] w_n415_0;
	wire[1:0] w_n417_0;
	wire[1:0] w_n420_0;
	wire[1:0] w_n422_0;
	wire[1:0] w_n425_0;
	wire[1:0] w_n427_0;
	wire[1:0] w_n430_0;
	wire[1:0] w_n432_0;
	wire[1:0] w_n435_0;
	wire[1:0] w_n437_0;
	wire[1:0] w_n441_0;
	wire[1:0] w_n442_0;
	wire[1:0] w_n443_0;
	wire[1:0] w_n445_0;
	wire[2:0] w_n446_0;
	wire[1:0] w_n447_0;
	wire[1:0] w_n450_0;
	wire[1:0] w_n452_0;
	wire[1:0] w_n453_0;
	wire[1:0] w_n454_0;
	wire[1:0] w_n455_0;
	wire[1:0] w_n456_0;
	wire[1:0] w_n457_0;
	wire[1:0] w_n458_0;
	wire[1:0] w_n459_0;
	wire[1:0] w_n460_0;
	wire[1:0] w_n461_0;
	wire[1:0] w_n462_0;
	wire[1:0] w_n463_0;
	wire[1:0] w_n464_0;
	wire[1:0] w_n465_0;
	wire[1:0] w_n466_0;
	wire[1:0] w_n468_0;
	wire[1:0] w_n469_0;
	wire[1:0] w_n471_0;
	wire[1:0] w_n476_0;
	wire[1:0] w_n477_0;
	wire[2:0] w_n482_0;
	wire[1:0] w_n484_0;
	wire[1:0] w_n487_0;
	wire[1:0] w_n489_0;
	wire[1:0] w_n492_0;
	wire[1:0] w_n494_0;
	wire[1:0] w_n497_0;
	wire[1:0] w_n499_0;
	wire[1:0] w_n502_0;
	wire[1:0] w_n504_0;
	wire[1:0] w_n507_0;
	wire[1:0] w_n509_0;
	wire[1:0] w_n512_0;
	wire[1:0] w_n514_0;
	wire[1:0] w_n518_0;
	wire[1:0] w_n519_0;
	wire[1:0] w_n520_0;
	wire[1:0] w_n522_0;
	wire[2:0] w_n523_0;
	wire[1:0] w_n524_0;
	wire[1:0] w_n527_0;
	wire[1:0] w_n529_0;
	wire[1:0] w_n530_0;
	wire[1:0] w_n531_0;
	wire[1:0] w_n532_0;
	wire[1:0] w_n533_0;
	wire[1:0] w_n534_0;
	wire[1:0] w_n535_0;
	wire[1:0] w_n536_0;
	wire[1:0] w_n537_0;
	wire[1:0] w_n538_0;
	wire[1:0] w_n539_0;
	wire[1:0] w_n540_0;
	wire[1:0] w_n541_0;
	wire[1:0] w_n542_0;
	wire[1:0] w_n543_0;
	wire[1:0] w_n544_0;
	wire[1:0] w_n545_0;
	wire[1:0] w_n547_0;
	wire[1:0] w_n548_0;
	wire[1:0] w_n550_0;
	wire[1:0] w_n555_0;
	wire[1:0] w_n556_0;
	wire[2:0] w_n561_0;
	wire[1:0] w_n563_0;
	wire[1:0] w_n566_0;
	wire[1:0] w_n568_0;
	wire[1:0] w_n571_0;
	wire[1:0] w_n573_0;
	wire[1:0] w_n576_0;
	wire[1:0] w_n578_0;
	wire[1:0] w_n581_0;
	wire[1:0] w_n583_0;
	wire[1:0] w_n586_0;
	wire[1:0] w_n588_0;
	wire[1:0] w_n591_0;
	wire[1:0] w_n593_0;
	wire[1:0] w_n596_0;
	wire[1:0] w_n598_0;
	wire[1:0] w_n602_0;
	wire[1:0] w_n603_0;
	wire[1:0] w_n604_0;
	wire[1:0] w_n606_0;
	wire[2:0] w_n607_0;
	wire[1:0] w_n608_0;
	wire[1:0] w_n611_0;
	wire[1:0] w_n613_0;
	wire[1:0] w_n614_0;
	wire[1:0] w_n615_0;
	wire[1:0] w_n616_0;
	wire[1:0] w_n617_0;
	wire[1:0] w_n618_0;
	wire[1:0] w_n619_0;
	wire[1:0] w_n620_0;
	wire[1:0] w_n621_0;
	wire[1:0] w_n622_0;
	wire[1:0] w_n623_0;
	wire[1:0] w_n624_0;
	wire[1:0] w_n625_0;
	wire[1:0] w_n626_0;
	wire[1:0] w_n627_0;
	wire[1:0] w_n628_0;
	wire[1:0] w_n629_0;
	wire[1:0] w_n630_0;
	wire[1:0] w_n631_0;
	wire[1:0] w_n633_0;
	wire[1:0] w_n634_0;
	wire[1:0] w_n636_0;
	wire[1:0] w_n641_0;
	wire[1:0] w_n642_0;
	wire[2:0] w_n647_0;
	wire[1:0] w_n649_0;
	wire[1:0] w_n652_0;
	wire[1:0] w_n654_0;
	wire[1:0] w_n657_0;
	wire[1:0] w_n659_0;
	wire[1:0] w_n662_0;
	wire[1:0] w_n664_0;
	wire[1:0] w_n667_0;
	wire[1:0] w_n669_0;
	wire[1:0] w_n672_0;
	wire[1:0] w_n674_0;
	wire[1:0] w_n677_0;
	wire[1:0] w_n679_0;
	wire[1:0] w_n682_0;
	wire[1:0] w_n684_0;
	wire[1:0] w_n687_0;
	wire[1:0] w_n689_0;
	wire[1:0] w_n693_0;
	wire[1:0] w_n694_0;
	wire[2:0] w_n695_0;
	wire[1:0] w_n697_0;
	wire[2:0] w_n698_0;
	wire[1:0] w_n699_0;
	wire[1:0] w_n702_0;
	wire[1:0] w_n704_0;
	wire[1:0] w_n705_0;
	wire[1:0] w_n706_0;
	wire[1:0] w_n707_0;
	wire[1:0] w_n708_0;
	wire[1:0] w_n709_0;
	wire[1:0] w_n710_0;
	wire[1:0] w_n711_0;
	wire[1:0] w_n712_0;
	wire[1:0] w_n713_0;
	wire[1:0] w_n714_0;
	wire[1:0] w_n715_0;
	wire[1:0] w_n716_0;
	wire[1:0] w_n717_0;
	wire[1:0] w_n718_0;
	wire[1:0] w_n719_0;
	wire[1:0] w_n720_0;
	wire[1:0] w_n721_0;
	wire[1:0] w_n722_0;
	wire[1:0] w_n723_0;
	wire[1:0] w_n724_0;
	wire[1:0] w_n726_0;
	wire[1:0] w_n727_0;
	wire[1:0] w_n729_0;
	wire[1:0] w_n734_0;
	wire[1:0] w_n735_0;
	wire[2:0] w_n740_0;
	wire[1:0] w_n742_0;
	wire[1:0] w_n745_0;
	wire[1:0] w_n747_0;
	wire[1:0] w_n750_0;
	wire[1:0] w_n752_0;
	wire[1:0] w_n755_0;
	wire[1:0] w_n757_0;
	wire[1:0] w_n760_0;
	wire[1:0] w_n762_0;
	wire[1:0] w_n765_0;
	wire[1:0] w_n767_0;
	wire[1:0] w_n770_0;
	wire[1:0] w_n772_0;
	wire[1:0] w_n775_0;
	wire[1:0] w_n777_0;
	wire[1:0] w_n780_0;
	wire[1:0] w_n782_0;
	wire[1:0] w_n785_0;
	wire[1:0] w_n787_0;
	wire[1:0] w_n791_0;
	wire[1:0] w_n792_0;
	wire[1:0] w_n793_0;
	wire[1:0] w_n795_0;
	wire[2:0] w_n797_0;
	wire[1:0] w_n800_0;
	wire[1:0] w_n802_0;
	wire[1:0] w_n803_0;
	wire[1:0] w_n804_0;
	wire[1:0] w_n805_0;
	wire[1:0] w_n806_0;
	wire[1:0] w_n807_0;
	wire[1:0] w_n808_0;
	wire[1:0] w_n809_0;
	wire[1:0] w_n810_0;
	wire[1:0] w_n811_0;
	wire[1:0] w_n812_0;
	wire[1:0] w_n813_0;
	wire[1:0] w_n814_0;
	wire[1:0] w_n815_0;
	wire[1:0] w_n816_0;
	wire[1:0] w_n817_0;
	wire[1:0] w_n818_0;
	wire[1:0] w_n819_0;
	wire[1:0] w_n820_0;
	wire[1:0] w_n821_0;
	wire[1:0] w_n822_0;
	wire[1:0] w_n823_0;
	wire[1:0] w_n824_0;
	wire[1:0] w_n826_0;
	wire[1:0] w_n827_0;
	wire[1:0] w_n829_0;
	wire[1:0] w_n834_0;
	wire[1:0] w_n835_0;
	wire[1:0] w_n839_0;
	wire[1:0] w_n840_0;
	wire[2:0] w_n844_0;
	wire[1:0] w_n846_0;
	wire[1:0] w_n849_0;
	wire[1:0] w_n851_0;
	wire[1:0] w_n854_0;
	wire[1:0] w_n856_0;
	wire[1:0] w_n859_0;
	wire[1:0] w_n861_0;
	wire[1:0] w_n864_0;
	wire[1:0] w_n866_0;
	wire[1:0] w_n869_0;
	wire[1:0] w_n871_0;
	wire[1:0] w_n874_0;
	wire[1:0] w_n876_0;
	wire[1:0] w_n879_0;
	wire[1:0] w_n881_0;
	wire[1:0] w_n884_0;
	wire[1:0] w_n886_0;
	wire[1:0] w_n889_0;
	wire[1:0] w_n891_0;
	wire[1:0] w_n895_0;
	wire[1:0] w_n896_0;
	wire[1:0] w_n897_0;
	wire[1:0] w_n898_0;
	wire[1:0] w_n901_0;
	wire[1:0] w_n903_0;
	wire[1:0] w_n906_0;
	wire[1:0] w_n907_0;
	wire[1:0] w_n908_0;
	wire[1:0] w_n909_0;
	wire[1:0] w_n910_0;
	wire[1:0] w_n911_0;
	wire[1:0] w_n912_0;
	wire[1:0] w_n913_0;
	wire[1:0] w_n914_0;
	wire[1:0] w_n915_0;
	wire[1:0] w_n916_0;
	wire[1:0] w_n917_0;
	wire[1:0] w_n918_0;
	wire[1:0] w_n919_0;
	wire[1:0] w_n920_0;
	wire[1:0] w_n921_0;
	wire[1:0] w_n922_0;
	wire[1:0] w_n923_0;
	wire[1:0] w_n924_0;
	wire[1:0] w_n925_0;
	wire[1:0] w_n926_0;
	wire[2:0] w_n927_0;
	wire[1:0] w_n929_0;
	wire[1:0] w_n930_0;
	wire[1:0] w_n931_0;
	wire[1:0] w_n932_0;
	wire[1:0] w_n937_0;
	wire[1:0] w_n938_0;
	wire[2:0] w_n942_0;
	wire[1:0] w_n943_0;
	wire[1:0] w_n949_0;
	wire[1:0] w_n951_0;
	wire[1:0] w_n954_0;
	wire[1:0] w_n956_0;
	wire[1:0] w_n959_0;
	wire[1:0] w_n961_0;
	wire[1:0] w_n964_0;
	wire[1:0] w_n966_0;
	wire[1:0] w_n969_0;
	wire[1:0] w_n971_0;
	wire[1:0] w_n974_0;
	wire[1:0] w_n976_0;
	wire[1:0] w_n979_0;
	wire[1:0] w_n981_0;
	wire[1:0] w_n984_0;
	wire[1:0] w_n986_0;
	wire[1:0] w_n989_0;
	wire[1:0] w_n991_0;
	wire[1:0] w_n994_0;
	wire[1:0] w_n996_0;
	wire[1:0] w_n999_0;
	wire[1:0] w_n1001_0;
	wire[1:0] w_n1005_0;
	wire[1:0] w_n1006_0;
	wire[1:0] w_n1008_0;
	wire[1:0] w_n1009_0;
	wire[1:0] w_n1010_0;
	wire[1:0] w_n1011_0;
	wire[1:0] w_n1012_0;
	wire[1:0] w_n1013_0;
	wire[1:0] w_n1014_0;
	wire[1:0] w_n1015_0;
	wire[1:0] w_n1016_0;
	wire[1:0] w_n1017_0;
	wire[1:0] w_n1018_0;
	wire[1:0] w_n1019_0;
	wire[1:0] w_n1020_0;
	wire[1:0] w_n1021_0;
	wire[1:0] w_n1022_0;
	wire[1:0] w_n1023_0;
	wire[1:0] w_n1024_0;
	wire[1:0] w_n1025_0;
	wire[1:0] w_n1026_0;
	wire[1:0] w_n1027_0;
	wire[1:0] w_n1028_0;
	wire[1:0] w_n1029_0;
	wire[1:0] w_n1030_0;
	wire[1:0] w_n1031_0;
	wire[1:0] w_n1032_0;
	wire[1:0] w_n1033_0;
	wire[1:0] w_n1034_0;
	wire[1:0] w_n1035_0;
	wire[1:0] w_n1037_0;
	wire[1:0] w_n1039_0;
	wire[1:0] w_n1043_0;
	wire[1:0] w_n1044_0;
	wire[1:0] w_n1048_0;
	wire[1:0] w_n1049_0;
	wire[1:0] w_n1052_0;
	wire[1:0] w_n1054_0;
	wire[1:0] w_n1057_0;
	wire[1:0] w_n1059_0;
	wire[1:0] w_n1062_0;
	wire[1:0] w_n1064_0;
	wire[1:0] w_n1067_0;
	wire[1:0] w_n1069_0;
	wire[1:0] w_n1072_0;
	wire[1:0] w_n1074_0;
	wire[1:0] w_n1077_0;
	wire[1:0] w_n1079_0;
	wire[1:0] w_n1082_0;
	wire[1:0] w_n1084_0;
	wire[1:0] w_n1087_0;
	wire[1:0] w_n1089_0;
	wire[1:0] w_n1092_0;
	wire[1:0] w_n1094_0;
	wire[1:0] w_n1097_0;
	wire[1:0] w_n1099_0;
	wire[1:0] w_n1102_0;
	wire[1:0] w_n1103_0;
	wire[1:0] w_n1109_0;
	wire[1:0] w_n1110_0;
	wire[1:0] w_n1114_0;
	wire[1:0] w_n1115_0;
	wire[1:0] w_n1116_0;
	wire[1:0] w_n1117_0;
	wire[1:0] w_n1118_0;
	wire[1:0] w_n1119_0;
	wire[1:0] w_n1120_0;
	wire[1:0] w_n1121_0;
	wire[1:0] w_n1122_0;
	wire[1:0] w_n1123_0;
	wire[1:0] w_n1124_0;
	wire[1:0] w_n1125_0;
	wire[1:0] w_n1126_0;
	wire[1:0] w_n1127_0;
	wire[1:0] w_n1128_0;
	wire[1:0] w_n1129_0;
	wire[1:0] w_n1130_0;
	wire[1:0] w_n1131_0;
	wire[1:0] w_n1132_0;
	wire[1:0] w_n1133_0;
	wire[1:0] w_n1134_0;
	wire[1:0] w_n1135_0;
	wire[1:0] w_n1137_0;
	wire[1:0] w_n1138_0;
	wire[1:0] w_n1139_0;
	wire[1:0] w_n1140_0;
	wire[1:0] w_n1141_0;
	wire[1:0] w_n1147_0;
	wire[1:0] w_n1151_0;
	wire[1:0] w_n1152_0;
	wire[1:0] w_n1156_0;
	wire[1:0] w_n1158_0;
	wire[1:0] w_n1161_0;
	wire[1:0] w_n1163_0;
	wire[1:0] w_n1166_0;
	wire[1:0] w_n1168_0;
	wire[1:0] w_n1171_0;
	wire[1:0] w_n1173_0;
	wire[1:0] w_n1176_0;
	wire[1:0] w_n1178_0;
	wire[1:0] w_n1181_0;
	wire[1:0] w_n1183_0;
	wire[1:0] w_n1186_0;
	wire[1:0] w_n1188_0;
	wire[1:0] w_n1191_0;
	wire[1:0] w_n1193_0;
	wire[1:0] w_n1196_0;
	wire[1:0] w_n1198_0;
	wire[1:0] w_n1201_0;
	wire[1:0] w_n1203_0;
	wire[1:0] w_n1206_0;
	wire[1:0] w_n1207_0;
	wire[1:0] w_n1208_0;
	wire[1:0] w_n1210_0;
	wire[1:0] w_n1212_0;
	wire[1:0] w_n1213_0;
	wire[1:0] w_n1214_0;
	wire[1:0] w_n1215_0;
	wire[1:0] w_n1216_0;
	wire[1:0] w_n1217_0;
	wire[1:0] w_n1218_0;
	wire[1:0] w_n1219_0;
	wire[1:0] w_n1220_0;
	wire[1:0] w_n1221_0;
	wire[1:0] w_n1222_0;
	wire[1:0] w_n1223_0;
	wire[1:0] w_n1224_0;
	wire[1:0] w_n1225_0;
	wire[1:0] w_n1226_0;
	wire[1:0] w_n1227_0;
	wire[1:0] w_n1228_0;
	wire[1:0] w_n1229_0;
	wire[1:0] w_n1230_0;
	wire[1:0] w_n1231_0;
	wire[1:0] w_n1232_0;
	wire[1:0] w_n1234_0;
	wire[1:0] w_n1236_0;
	wire[1:0] w_n1237_0;
	wire[1:0] w_n1238_0;
	wire[1:0] w_n1244_0;
	wire[1:0] w_n1247_0;
	wire[1:0] w_n1248_0;
	wire[1:0] w_n1251_0;
	wire[1:0] w_n1253_0;
	wire[1:0] w_n1256_0;
	wire[1:0] w_n1258_0;
	wire[1:0] w_n1261_0;
	wire[1:0] w_n1263_0;
	wire[1:0] w_n1266_0;
	wire[1:0] w_n1268_0;
	wire[1:0] w_n1271_0;
	wire[1:0] w_n1273_0;
	wire[1:0] w_n1276_0;
	wire[1:0] w_n1278_0;
	wire[1:0] w_n1281_0;
	wire[1:0] w_n1283_0;
	wire[1:0] w_n1286_0;
	wire[1:0] w_n1288_0;
	wire[1:0] w_n1291_0;
	wire[1:0] w_n1293_0;
	wire[1:0] w_n1296_0;
	wire[1:0] w_n1297_0;
	wire[1:0] w_n1298_0;
	wire[1:0] w_n1301_0;
	wire[1:0] w_n1303_0;
	wire[1:0] w_n1304_0;
	wire[1:0] w_n1305_0;
	wire[1:0] w_n1306_0;
	wire[1:0] w_n1307_0;
	wire[1:0] w_n1308_0;
	wire[1:0] w_n1309_0;
	wire[1:0] w_n1310_0;
	wire[1:0] w_n1311_0;
	wire[1:0] w_n1312_0;
	wire[1:0] w_n1313_0;
	wire[1:0] w_n1314_0;
	wire[1:0] w_n1315_0;
	wire[1:0] w_n1316_0;
	wire[1:0] w_n1317_0;
	wire[1:0] w_n1318_0;
	wire[1:0] w_n1319_0;
	wire[1:0] w_n1320_0;
	wire[1:0] w_n1321_0;
	wire[1:0] w_n1322_0;
	wire[1:0] w_n1324_0;
	wire[1:0] w_n1325_0;
	wire[1:0] w_n1326_0;
	wire[1:0] w_n1332_0;
	wire[1:0] w_n1337_0;
	wire[1:0] w_n1338_0;
	wire[1:0] w_n1341_0;
	wire[1:0] w_n1343_0;
	wire[1:0] w_n1346_0;
	wire[1:0] w_n1348_0;
	wire[1:0] w_n1351_0;
	wire[1:0] w_n1353_0;
	wire[1:0] w_n1356_0;
	wire[1:0] w_n1358_0;
	wire[1:0] w_n1361_0;
	wire[1:0] w_n1363_0;
	wire[1:0] w_n1366_0;
	wire[1:0] w_n1368_0;
	wire[1:0] w_n1371_0;
	wire[1:0] w_n1373_0;
	wire[1:0] w_n1376_0;
	wire[1:0] w_n1378_0;
	wire[1:0] w_n1381_0;
	wire[1:0] w_n1382_0;
	wire[1:0] w_n1383_0;
	wire[1:0] w_n1386_0;
	wire[1:0] w_n1388_0;
	wire[1:0] w_n1389_0;
	wire[1:0] w_n1390_0;
	wire[1:0] w_n1391_0;
	wire[1:0] w_n1392_0;
	wire[1:0] w_n1393_0;
	wire[1:0] w_n1394_0;
	wire[1:0] w_n1395_0;
	wire[1:0] w_n1396_0;
	wire[1:0] w_n1397_0;
	wire[1:0] w_n1398_0;
	wire[1:0] w_n1399_0;
	wire[1:0] w_n1400_0;
	wire[1:0] w_n1401_0;
	wire[1:0] w_n1402_0;
	wire[1:0] w_n1403_0;
	wire[1:0] w_n1404_0;
	wire[1:0] w_n1405_0;
	wire[1:0] w_n1407_0;
	wire[1:0] w_n1409_0;
	wire[1:0] w_n1410_0;
	wire[1:0] w_n1415_0;
	wire[1:0] w_n1420_0;
	wire[1:0] w_n1421_0;
	wire[1:0] w_n1424_0;
	wire[1:0] w_n1426_0;
	wire[1:0] w_n1429_0;
	wire[1:0] w_n1431_0;
	wire[1:0] w_n1434_0;
	wire[1:0] w_n1436_0;
	wire[1:0] w_n1439_0;
	wire[1:0] w_n1441_0;
	wire[1:0] w_n1444_0;
	wire[1:0] w_n1446_0;
	wire[1:0] w_n1449_0;
	wire[1:0] w_n1451_0;
	wire[1:0] w_n1454_0;
	wire[1:0] w_n1456_0;
	wire[1:0] w_n1459_0;
	wire[1:0] w_n1460_0;
	wire[1:0] w_n1461_0;
	wire[1:0] w_n1464_0;
	wire[1:0] w_n1466_0;
	wire[1:0] w_n1467_0;
	wire[1:0] w_n1468_0;
	wire[1:0] w_n1469_0;
	wire[1:0] w_n1470_0;
	wire[1:0] w_n1471_0;
	wire[1:0] w_n1472_0;
	wire[1:0] w_n1473_0;
	wire[1:0] w_n1474_0;
	wire[1:0] w_n1475_0;
	wire[1:0] w_n1476_0;
	wire[1:0] w_n1477_0;
	wire[1:0] w_n1478_0;
	wire[1:0] w_n1479_0;
	wire[1:0] w_n1480_0;
	wire[1:0] w_n1481_0;
	wire[1:0] w_n1483_0;
	wire[1:0] w_n1485_0;
	wire[1:0] w_n1486_0;
	wire[1:0] w_n1491_0;
	wire[1:0] w_n1496_0;
	wire[1:0] w_n1497_0;
	wire[1:0] w_n1500_0;
	wire[1:0] w_n1502_0;
	wire[1:0] w_n1505_0;
	wire[1:0] w_n1507_0;
	wire[1:0] w_n1510_0;
	wire[1:0] w_n1512_0;
	wire[1:0] w_n1515_0;
	wire[1:0] w_n1517_0;
	wire[1:0] w_n1520_0;
	wire[1:0] w_n1522_0;
	wire[1:0] w_n1525_0;
	wire[1:0] w_n1527_0;
	wire[1:0] w_n1530_0;
	wire[1:0] w_n1531_0;
	wire[1:0] w_n1532_0;
	wire[1:0] w_n1535_0;
	wire[1:0] w_n1537_0;
	wire[1:0] w_n1538_0;
	wire[1:0] w_n1539_0;
	wire[1:0] w_n1540_0;
	wire[1:0] w_n1541_0;
	wire[1:0] w_n1542_0;
	wire[1:0] w_n1543_0;
	wire[1:0] w_n1544_0;
	wire[1:0] w_n1545_0;
	wire[1:0] w_n1546_0;
	wire[1:0] w_n1547_0;
	wire[1:0] w_n1548_0;
	wire[1:0] w_n1549_0;
	wire[1:0] w_n1550_0;
	wire[1:0] w_n1552_0;
	wire[1:0] w_n1554_0;
	wire[1:0] w_n1555_0;
	wire[1:0] w_n1560_0;
	wire[1:0] w_n1565_0;
	wire[1:0] w_n1566_0;
	wire[1:0] w_n1569_0;
	wire[1:0] w_n1571_0;
	wire[1:0] w_n1574_0;
	wire[1:0] w_n1576_0;
	wire[1:0] w_n1579_0;
	wire[1:0] w_n1581_0;
	wire[1:0] w_n1584_0;
	wire[1:0] w_n1586_0;
	wire[1:0] w_n1589_0;
	wire[1:0] w_n1591_0;
	wire[1:0] w_n1594_0;
	wire[1:0] w_n1595_0;
	wire[1:0] w_n1596_0;
	wire[1:0] w_n1599_0;
	wire[1:0] w_n1601_0;
	wire[1:0] w_n1602_0;
	wire[1:0] w_n1603_0;
	wire[1:0] w_n1604_0;
	wire[1:0] w_n1605_0;
	wire[1:0] w_n1606_0;
	wire[1:0] w_n1607_0;
	wire[1:0] w_n1608_0;
	wire[1:0] w_n1609_0;
	wire[1:0] w_n1610_0;
	wire[1:0] w_n1611_0;
	wire[1:0] w_n1612_0;
	wire[1:0] w_n1614_0;
	wire[1:0] w_n1616_0;
	wire[1:0] w_n1617_0;
	wire[1:0] w_n1622_0;
	wire[1:0] w_n1627_0;
	wire[1:0] w_n1628_0;
	wire[1:0] w_n1631_0;
	wire[1:0] w_n1633_0;
	wire[1:0] w_n1636_0;
	wire[1:0] w_n1638_0;
	wire[1:0] w_n1641_0;
	wire[1:0] w_n1643_0;
	wire[1:0] w_n1646_0;
	wire[1:0] w_n1648_0;
	wire[1:0] w_n1651_0;
	wire[1:0] w_n1652_0;
	wire[1:0] w_n1653_0;
	wire[1:0] w_n1656_0;
	wire[1:0] w_n1658_0;
	wire[1:0] w_n1659_0;
	wire[1:0] w_n1660_0;
	wire[1:0] w_n1661_0;
	wire[1:0] w_n1662_0;
	wire[1:0] w_n1663_0;
	wire[1:0] w_n1664_0;
	wire[1:0] w_n1665_0;
	wire[1:0] w_n1666_0;
	wire[1:0] w_n1667_0;
	wire[1:0] w_n1669_0;
	wire[1:0] w_n1671_0;
	wire[1:0] w_n1672_0;
	wire[1:0] w_n1677_0;
	wire[1:0] w_n1682_0;
	wire[1:0] w_n1684_0;
	wire[1:0] w_n1687_0;
	wire[1:0] w_n1689_0;
	wire[1:0] w_n1692_0;
	wire[1:0] w_n1694_0;
	wire[1:0] w_n1697_0;
	wire[1:0] w_n1699_0;
	wire[1:0] w_n1702_0;
	wire[1:0] w_n1703_0;
	wire[1:0] w_n1704_0;
	wire[1:0] w_n1707_0;
	wire[1:0] w_n1709_0;
	wire[1:0] w_n1710_0;
	wire[1:0] w_n1711_0;
	wire[1:0] w_n1712_0;
	wire[1:0] w_n1713_0;
	wire[1:0] w_n1714_0;
	wire[1:0] w_n1715_0;
	wire[1:0] w_n1716_0;
	wire[1:0] w_n1717_0;
	wire[1:0] w_n1719_0;
	wire[1:0] w_n1720_0;
	wire[1:0] w_n1725_0;
	wire[1:0] w_n1728_0;
	wire[1:0] w_n1730_0;
	wire[1:0] w_n1733_0;
	wire[1:0] w_n1735_0;
	wire[1:0] w_n1738_0;
	wire[1:0] w_n1740_0;
	wire[1:0] w_n1743_0;
	wire[1:0] w_n1744_0;
	wire[1:0] w_n1745_0;
	wire[1:0] w_n1748_0;
	wire[1:0] w_n1750_0;
	wire[1:0] w_n1751_0;
	wire[1:0] w_n1752_0;
	wire[1:0] w_n1753_0;
	wire[1:0] w_n1754_0;
	wire[1:0] w_n1755_0;
	wire[1:0] w_n1756_0;
	wire[1:0] w_n1757_0;
	wire[1:0] w_n1758_0;
	wire[1:0] w_n1765_0;
	wire[1:0] w_n1768_0;
	wire[1:0] w_n1770_0;
	wire[1:0] w_n1773_0;
	wire[1:0] w_n1775_0;
	wire[1:0] w_n1778_0;
	wire[1:0] w_n1779_0;
	wire[1:0] w_n1780_0;
	wire[1:0] w_n1783_0;
	wire[1:0] w_n1785_0;
	wire[1:0] w_n1786_0;
	wire[1:0] w_n1787_0;
	wire[1:0] w_n1788_0;
	wire[1:0] w_n1789_0;
	wire[1:0] w_n1790_0;
	wire[1:0] w_n1791_0;
	wire[1:0] w_n1798_0;
	wire[1:0] w_n1801_0;
	wire[1:0] w_n1803_0;
	wire[1:0] w_n1806_0;
	wire[1:0] w_n1807_0;
	wire[1:0] w_n1808_0;
	wire[1:0] w_n1811_0;
	wire[1:0] w_n1813_0;
	wire[1:0] w_n1814_0;
	wire[1:0] w_n1815_0;
	wire[1:0] w_n1816_0;
	wire[1:0] w_n1817_0;
	wire[1:0] w_n1824_0;
	wire[1:0] w_n1827_0;
	wire[1:0] w_n1828_0;
	wire[1:0] w_n1829_0;
	wire[1:0] w_n1832_0;
	wire[1:0] w_n1834_0;
	wire[1:0] w_n1835_0;
	wire[1:0] w_n1836_0;
	wire[1:0] w_n1838_0;
	wire[1:0] w_n1841_0;
	wire[1:0] w_n1848_0;
	wire[1:0] w_n1849_0;
	wire w_dff_B_3FRV3OSY1_1;
	wire w_dff_B_tzS6DnrW4_1;
	wire w_dff_B_VxIDHxam6_1;
	wire w_dff_B_ha9tIQWA4_1;
	wire w_dff_B_jMMSq32A1_1;
	wire w_dff_B_ZlFNlmzc9_1;
	wire w_dff_B_6XD066jy3_1;
	wire w_dff_B_9OzVm5of4_1;
	wire w_dff_B_veTJQclE4_1;
	wire w_dff_B_x5apiaGv1_1;
	wire w_dff_B_1mlkccCS3_1;
	wire w_dff_B_cSsKQ9UH7_1;
	wire w_dff_B_TqF3Kyx21_1;
	wire w_dff_B_YjBbOTB80_1;
	wire w_dff_B_BOxqgtoR5_1;
	wire w_dff_B_Xxmuud8I0_1;
	wire w_dff_B_b1tBh9bS4_1;
	wire w_dff_B_UsYlwApm6_1;
	wire w_dff_B_DsS1jNqW1_1;
	wire w_dff_B_8wetMZx70_1;
	wire w_dff_B_l6ggz8262_1;
	wire w_dff_B_8JplcJiB0_1;
	wire w_dff_B_XbHPK9DO3_1;
	wire w_dff_B_e6cgpSpf1_1;
	wire w_dff_B_2KBjygSb8_1;
	wire w_dff_B_8yoM9yav3_1;
	wire w_dff_B_tlcf4OLo2_1;
	wire w_dff_B_4imTgWz93_1;
	wire w_dff_B_jb3PVe8J8_1;
	wire w_dff_B_3BUodJPE9_1;
	wire w_dff_B_0574HHts2_1;
	wire w_dff_B_1mRT852b6_1;
	wire w_dff_B_r5OIKcNp3_1;
	wire w_dff_B_ywNGUkGh3_1;
	wire w_dff_B_QcEJJi5q5_1;
	wire w_dff_B_2sZeV0CD3_1;
	wire w_dff_B_ghT6ytBR1_1;
	wire w_dff_B_ysQBawSr4_1;
	wire w_dff_B_pveCeIwn2_1;
	wire w_dff_B_VObvQZJ06_1;
	wire w_dff_B_ExXvj7BS1_1;
	wire w_dff_B_j1cevLAF1_1;
	wire w_dff_B_GxfvPRXo7_1;
	wire w_dff_B_HhQvWPrz0_1;
	wire w_dff_B_mnqfQLlW2_1;
	wire w_dff_B_z9VEiMmP8_1;
	wire w_dff_B_xMn0ITae1_1;
	wire w_dff_B_ewCwHZCZ0_1;
	wire w_dff_B_QoLFz0zf3_1;
	wire w_dff_B_l86IBcNm1_1;
	wire w_dff_B_kiwggGnl5_1;
	wire w_dff_B_abxSj8tI2_1;
	wire w_dff_B_fmM58jD45_1;
	wire w_dff_B_SVDUn8oa2_1;
	wire w_dff_B_j3ONxwAh5_1;
	wire w_dff_B_aw7WoDnN4_1;
	wire w_dff_B_7GY3ZO541_1;
	wire w_dff_B_lOjagvgO9_1;
	wire w_dff_B_vYASkG8n9_1;
	wire w_dff_B_U1Pd7OVs7_1;
	wire w_dff_B_5zUAPdQo9_1;
	wire w_dff_B_GsaYMcr60_1;
	wire w_dff_B_cknEWKCP9_1;
	wire w_dff_B_RTzxDbo07_1;
	wire w_dff_B_tfuvyd3x2_1;
	wire w_dff_B_AF5hPx0J7_1;
	wire w_dff_B_uXxDI9bO5_1;
	wire w_dff_B_rjvlO9LX2_1;
	wire w_dff_B_LDGGGVfw2_1;
	wire w_dff_B_TAGRaUJf0_1;
	wire w_dff_B_m3IXWPoE5_1;
	wire w_dff_B_fq4LRnHV2_1;
	wire w_dff_B_P0aUQM8E8_1;
	wire w_dff_B_RyggImi25_1;
	wire w_dff_B_s5qXbtjj8_1;
	wire w_dff_B_yarOBbtK5_1;
	wire w_dff_B_4iVZKolt8_1;
	wire w_dff_B_i7QAnRf78_1;
	wire w_dff_B_L4G8jCl37_1;
	wire w_dff_B_eGvjOvZb0_1;
	wire w_dff_B_OEpOfUij9_1;
	wire w_dff_B_LpCIXDfk1_1;
	wire w_dff_B_f7FUm4Yq4_1;
	wire w_dff_B_LgnLW0fG9_1;
	wire w_dff_B_OdqFMnh06_1;
	wire w_dff_B_nB35EGLw1_1;
	wire w_dff_B_IUKdWtAb3_1;
	wire w_dff_B_0GZO3Pon4_1;
	wire w_dff_B_MCKfq1186_1;
	wire w_dff_B_VND7Ereb9_1;
	wire w_dff_B_WDv7auJn1_1;
	wire w_dff_B_NtzpAMMQ5_1;
	wire w_dff_B_tM6B2SdG8_1;
	wire w_dff_B_hxb9EYi46_1;
	wire w_dff_B_HAvgtCbm0_1;
	wire w_dff_B_xlDvBJx33_1;
	wire w_dff_B_I3fXIWZ77_1;
	wire w_dff_B_mnw3fniH1_1;
	wire w_dff_B_zvg1jZKl6_1;
	wire w_dff_B_dluCOjUp9_1;
	wire w_dff_B_U0UsSENG4_1;
	wire w_dff_B_NyKtFR510_1;
	wire w_dff_B_jj6fPb5s9_1;
	wire w_dff_B_emUqo5MA2_1;
	wire w_dff_B_09jwJg3T4_1;
	wire w_dff_B_QI2QzpDT6_1;
	wire w_dff_B_AJT4CnW13_1;
	wire w_dff_B_emjodvUZ5_1;
	wire w_dff_B_LVmnjLSK7_1;
	wire w_dff_B_HMddPGFz1_1;
	wire w_dff_B_xCTg7QvE2_1;
	wire w_dff_B_d8mlmS3d1_1;
	wire w_dff_B_6rj66GPP9_1;
	wire w_dff_B_BegVnqY61_1;
	wire w_dff_B_nlzDf3JQ8_1;
	wire w_dff_B_p5ZFmHRw7_1;
	wire w_dff_B_7PYVdMoG0_1;
	wire w_dff_B_f7ERvtf70_1;
	wire w_dff_B_wiUZgfzF6_1;
	wire w_dff_B_HhkEzole3_1;
	wire w_dff_B_ClOxpV8b1_1;
	wire w_dff_B_fAWMF5Wi6_1;
	wire w_dff_B_j4ubxkx71_1;
	wire w_dff_B_g0qfZzsD4_1;
	wire w_dff_B_7qAExO8r4_1;
	wire w_dff_B_2qeprMuU1_1;
	wire w_dff_B_YTgH9Afm7_1;
	wire w_dff_B_zcqFA8Wl0_1;
	wire w_dff_B_zOMgdbVA7_1;
	wire w_dff_B_lVWfBE479_1;
	wire w_dff_B_rWv6YpuE1_1;
	wire w_dff_B_slmxmLJT8_1;
	wire w_dff_B_JoeVYMHM5_1;
	wire w_dff_B_zSendvSt1_1;
	wire w_dff_B_S15Yp8XT0_1;
	wire w_dff_B_ot8aqExn0_1;
	wire w_dff_B_CFn3SMXg3_1;
	wire w_dff_B_mn1cQTSZ7_1;
	wire w_dff_B_fb82xcaX4_1;
	wire w_dff_B_oU3W5YhB5_1;
	wire w_dff_B_mBXNtslG7_1;
	wire w_dff_B_f2vFp1tY3_1;
	wire w_dff_B_0TqlkH5f5_1;
	wire w_dff_B_KpMIxvXc7_1;
	wire w_dff_B_N82dfrYa9_1;
	wire w_dff_B_vV4gSXGs0_1;
	wire w_dff_B_o8lrPJoM1_1;
	wire w_dff_B_r0o7HmVf9_1;
	wire w_dff_B_bjGuhllO6_1;
	wire w_dff_B_T1AUH2Ff3_1;
	wire w_dff_B_5aQGEkCr3_1;
	wire w_dff_B_atN5qAza3_1;
	wire w_dff_B_x6V5G3zo2_1;
	wire w_dff_B_6mRlSyiG1_1;
	wire w_dff_B_2HrLUCD95_1;
	wire w_dff_B_SAwXU5909_1;
	wire w_dff_B_alzmbQ5D8_1;
	wire w_dff_B_uos9j3hj8_1;
	wire w_dff_B_p6s9f53C7_1;
	wire w_dff_B_23sqyV4G0_1;
	wire w_dff_B_tmRTLLGG7_1;
	wire w_dff_B_LdNvkQAU9_1;
	wire w_dff_B_ksqaA3H48_1;
	wire w_dff_B_n4wnCgRt3_1;
	wire w_dff_B_tHAqzUIO9_1;
	wire w_dff_B_LiPwz7S20_1;
	wire w_dff_B_fS7HDFdk1_1;
	wire w_dff_B_vd6OvMni6_1;
	wire w_dff_B_X402efUH3_1;
	wire w_dff_B_YBmjWnM61_1;
	wire w_dff_B_wttfy1U82_1;
	wire w_dff_B_DBNqSZ240_1;
	wire w_dff_B_d8wE2Uer4_1;
	wire w_dff_B_QZdtZDCn1_1;
	wire w_dff_B_Yr1vIQ269_1;
	wire w_dff_B_rp1raYfx8_1;
	wire w_dff_B_kCXG7ccs1_1;
	wire w_dff_B_tfPxnPeR4_1;
	wire w_dff_B_KyjXoe9I9_1;
	wire w_dff_B_WXo3Jx9S1_1;
	wire w_dff_B_CQWxuADi2_1;
	wire w_dff_B_ewuybWPi6_1;
	wire w_dff_B_nFucVkYg9_1;
	wire w_dff_B_OEPrANys4_1;
	wire w_dff_B_3FMTbEV32_1;
	wire w_dff_B_cVsX0Vlq1_1;
	wire w_dff_B_7yipnxMK4_1;
	wire w_dff_B_mZLm2enn4_1;
	wire w_dff_B_Mld6iIyQ6_1;
	wire w_dff_B_alg5Gp4J8_1;
	wire w_dff_B_M7md7Umi8_1;
	wire w_dff_B_4VdDZshB9_1;
	wire w_dff_B_kqR09lbr4_1;
	wire w_dff_B_QPegivjI8_1;
	wire w_dff_B_SDOqiyuU7_1;
	wire w_dff_B_oBlrIWPA2_1;
	wire w_dff_B_B5qQ1p6k5_1;
	wire w_dff_B_GYsVnjmm1_1;
	wire w_dff_B_be6zHySW2_1;
	wire w_dff_B_SWoxspAq3_1;
	wire w_dff_B_6m5zXTgz9_1;
	wire w_dff_B_DAUafqyZ5_1;
	wire w_dff_B_hZnynIeh0_1;
	wire w_dff_B_ifkqVlaJ3_1;
	wire w_dff_B_29WaMTkW6_1;
	wire w_dff_B_QUYCBp1w1_1;
	wire w_dff_B_MYLIJuEe3_1;
	wire w_dff_B_pAA7W6Lg1_1;
	wire w_dff_B_gL4nA4Lz8_1;
	wire w_dff_B_3CG9xstA3_1;
	wire w_dff_B_1Qz7w2UC3_1;
	wire w_dff_B_8vGu5hgd2_1;
	wire w_dff_B_rOZ0ysnI4_1;
	wire w_dff_B_8NtzV6A68_1;
	wire w_dff_B_Yb6stWZa1_1;
	wire w_dff_B_Uv0qjueR9_1;
	wire w_dff_B_evmr8apB2_1;
	wire w_dff_B_Q0tinFuv6_1;
	wire w_dff_B_PmDzMrum9_1;
	wire w_dff_B_gE6BLSiU0_1;
	wire w_dff_B_ZYRBFtCg1_1;
	wire w_dff_B_6M1Gccuy5_1;
	wire w_dff_B_c4FUp6yr5_1;
	wire w_dff_B_9uueaT3B7_1;
	wire w_dff_B_n74dByiy5_1;
	wire w_dff_B_i5xs0pLM2_1;
	wire w_dff_B_D8QHiqNG5_1;
	wire w_dff_B_WEtqzBk58_1;
	wire w_dff_B_XxrgRmDw6_1;
	wire w_dff_B_ux8VR4h52_1;
	wire w_dff_B_0FWt9EOj8_1;
	wire w_dff_B_OeLgFibZ7_1;
	wire w_dff_B_8gitHIJ50_1;
	wire w_dff_B_3WcVn7vX6_1;
	wire w_dff_B_rEOHq21o6_1;
	wire w_dff_B_6NhvmuVH1_1;
	wire w_dff_B_RWn2bz0N6_1;
	wire w_dff_B_EWMTpNai1_1;
	wire w_dff_B_MerO0PB70_1;
	wire w_dff_B_kFLXeI0q6_1;
	wire w_dff_B_cyMf9eUe5_1;
	wire w_dff_B_1ZEggp9p7_1;
	wire w_dff_B_xLb88RAj3_1;
	wire w_dff_B_mtv59oc30_1;
	wire w_dff_B_Isi4F8E74_1;
	wire w_dff_B_Qcd02HFj4_1;
	wire w_dff_B_tPTGsLaV0_1;
	wire w_dff_B_sFUxrmKn2_1;
	wire w_dff_B_a9lb9UVr0_1;
	wire w_dff_B_hCoDeQjV6_1;
	wire w_dff_B_gzVFP90e4_1;
	wire w_dff_B_0WQxg2FI6_1;
	wire w_dff_B_7NcIjERV3_1;
	wire w_dff_B_nKF7123N6_1;
	wire w_dff_B_Ll9sTDLV6_1;
	wire w_dff_B_UiPn8pnG6_1;
	wire w_dff_B_B3QeUWtN6_1;
	wire w_dff_B_jjvuWWT53_1;
	wire w_dff_B_Cy24TzKo4_1;
	wire w_dff_B_AvrJc9Fh3_1;
	wire w_dff_B_7P7v1f2R5_1;
	wire w_dff_B_Ftur8imG0_1;
	wire w_dff_B_EuNF3oqt9_1;
	wire w_dff_B_ROre4ehw0_1;
	wire w_dff_B_Icv5Cas06_1;
	wire w_dff_B_6C3O9f618_1;
	wire w_dff_B_rtFAHHBq0_1;
	wire w_dff_B_SUPdgmT26_1;
	wire w_dff_B_HWA83ljg1_1;
	wire w_dff_B_3tb95YT87_1;
	wire w_dff_B_QlWV5ZWu3_1;
	wire w_dff_B_QYVvlqZl4_1;
	wire w_dff_B_tPk13MuO0_1;
	wire w_dff_B_NoJYw5590_1;
	wire w_dff_B_NfP8PkSF3_1;
	wire w_dff_B_tQwdKdFd9_1;
	wire w_dff_B_t68SnBns4_1;
	wire w_dff_B_5eOFGvez3_1;
	wire w_dff_B_EiwBf9Ie5_1;
	wire w_dff_B_cp3TvIVf9_1;
	wire w_dff_B_YUC97WWG0_1;
	wire w_dff_B_PXBcDd5b3_1;
	wire w_dff_B_hsZqMFhJ3_1;
	wire w_dff_B_bqNHNd9T7_1;
	wire w_dff_B_R6d7TecP0_1;
	wire w_dff_B_IFujLWY08_1;
	wire w_dff_B_xMYa2SRa8_1;
	wire w_dff_B_oCldZxq23_1;
	wire w_dff_B_IGGrZXnp3_1;
	wire w_dff_B_CTGbThQI0_1;
	wire w_dff_B_s79fFjKv1_1;
	wire w_dff_B_REH0IWYZ2_1;
	wire w_dff_B_083CD5wE9_1;
	wire w_dff_B_VSl1wgOi2_1;
	wire w_dff_B_aIONJ2mi4_1;
	wire w_dff_B_abvVIJ2j0_1;
	wire w_dff_B_0Y8Nd7JK9_1;
	wire w_dff_B_vwbuSnOT1_1;
	wire w_dff_B_7le6HbYy0_1;
	wire w_dff_B_UMLSg4MG9_1;
	wire w_dff_B_Js5upuCB5_1;
	wire w_dff_B_xsZlMiFw6_1;
	wire w_dff_B_tCrQe8HZ1_1;
	wire w_dff_B_JboN2GVL0_1;
	wire w_dff_B_VyhYR3BZ3_1;
	wire w_dff_B_aHGbkyCo1_1;
	wire w_dff_B_3QxYAQfJ2_1;
	wire w_dff_B_zLHK66928_1;
	wire w_dff_B_3BYEE1pX4_1;
	wire w_dff_B_9BFhlPnb4_1;
	wire w_dff_B_AP6uzT607_1;
	wire w_dff_B_DnPi3aFF2_1;
	wire w_dff_B_jUOIzjKU2_1;
	wire w_dff_B_EUCmrPbZ2_1;
	wire w_dff_B_RdmUctx22_1;
	wire w_dff_B_oZkFp8qa8_1;
	wire w_dff_B_pWo908Su2_1;
	wire w_dff_B_hTbA170c1_1;
	wire w_dff_B_4aWxsDc90_1;
	wire w_dff_B_91vhNdIB6_1;
	wire w_dff_B_94Tj5YPh4_1;
	wire w_dff_B_UQjdE8xZ5_1;
	wire w_dff_B_VnsM0W395_1;
	wire w_dff_B_wdDfIAoD4_1;
	wire w_dff_B_Ni3DAazg6_1;
	wire w_dff_B_AcOt0G3U1_1;
	wire w_dff_B_Njn7T5vJ0_1;
	wire w_dff_B_FDPn5Wpe1_1;
	wire w_dff_B_DFYNvs9J6_1;
	wire w_dff_B_eG6R2dfb6_1;
	wire w_dff_B_nYPmOVXp3_0;
	wire w_dff_B_h2NQdNi83_1;
	wire w_dff_B_w6xAud9Y6_1;
	wire w_dff_B_j1HUws5y5_1;
	wire w_dff_B_weuFHwps7_1;
	wire w_dff_B_K4gMSjdJ2_1;
	wire w_dff_B_UK1pMBul3_1;
	wire w_dff_B_dpAYw9U66_1;
	wire w_dff_B_3FPqNqRg6_1;
	wire w_dff_B_RMgXq30i1_1;
	wire w_dff_B_GuIkOsrU9_1;
	wire w_dff_B_eOPWVIyh9_1;
	wire w_dff_B_98YfWaMd6_1;
	wire w_dff_B_AJQXN7UJ4_1;
	wire w_dff_B_39OHMP0W1_0;
	wire w_dff_B_OUfenZMD6_0;
	wire w_dff_B_L6Be0ODT9_0;
	wire w_dff_B_Zy4gqZv55_0;
	wire w_dff_B_15S0DRQx3_0;
	wire w_dff_B_NGHghf4S2_0;
	wire w_dff_B_yATPcVva5_0;
	wire w_dff_B_P11wpji41_0;
	wire w_dff_B_xYQC0U1N6_0;
	wire w_dff_B_r8nRu9jp0_0;
	wire w_dff_B_6I7wTHAp0_0;
	wire w_dff_A_ut6G07172_0;
	wire w_dff_A_j8oWk5Pk2_0;
	wire w_dff_A_4eV7sBfX8_0;
	wire w_dff_A_2MoJfxAt0_0;
	wire w_dff_A_VCXPxjPL6_0;
	wire w_dff_A_EwPuKEHs2_0;
	wire w_dff_A_zj2c6nf41_0;
	wire w_dff_A_ZhxcM4KJ4_0;
	wire w_dff_A_lugix02b7_0;
	wire w_dff_A_IPF9IkbT3_0;
	wire w_dff_A_284Si4af7_0;
	wire w_dff_A_QBk0R33Z3_0;
	wire w_dff_B_xVnw1T4P0_1;
	wire w_dff_B_WeG7aV7r0_1;
	wire w_dff_B_ge5YKwtn3_2;
	wire w_dff_B_uOnjh6FF0_2;
	wire w_dff_B_7dltARmO9_2;
	wire w_dff_B_dYqFSJCv4_2;
	wire w_dff_B_hDWLPYSj5_2;
	wire w_dff_B_ktoieRTt7_2;
	wire w_dff_B_eGcA9lNu1_2;
	wire w_dff_B_GLCtRJhO2_2;
	wire w_dff_B_UhUHDKJs4_2;
	wire w_dff_B_v8rodcin4_2;
	wire w_dff_B_9D2a0kP39_2;
	wire w_dff_B_IRruBjsc7_2;
	wire w_dff_B_9SBKtdGh8_2;
	wire w_dff_B_MCcCQBYY6_2;
	wire w_dff_B_HZ0SNEbB3_2;
	wire w_dff_B_xsA2ur2w2_2;
	wire w_dff_B_ZfUXriGL6_2;
	wire w_dff_B_ZyGa1XKK1_2;
	wire w_dff_B_noLV7L8v9_2;
	wire w_dff_B_pwctVWsi5_2;
	wire w_dff_B_ALlT3D7p5_2;
	wire w_dff_B_9zlQwrjG4_2;
	wire w_dff_B_5Hh2I43g5_2;
	wire w_dff_B_3Z2Abyrm9_2;
	wire w_dff_B_QVE63Xpr3_2;
	wire w_dff_B_gMekOidd8_2;
	wire w_dff_B_WlBOIRCB2_2;
	wire w_dff_B_bi5BQzpe5_2;
	wire w_dff_B_P91ieAHo2_2;
	wire w_dff_B_wilyBuqr6_2;
	wire w_dff_B_ERYonw4I7_2;
	wire w_dff_B_Lr5wXo5p7_2;
	wire w_dff_B_P9xRXVrX5_2;
	wire w_dff_B_ilDlmYak6_2;
	wire w_dff_B_WwsrPN2o0_2;
	wire w_dff_B_13jMJ3xx1_2;
	wire w_dff_B_JRJiaY1R1_2;
	wire w_dff_B_yH53UUPr2_2;
	wire w_dff_B_2m82q0HC0_2;
	wire w_dff_B_uQcGInwi9_2;
	wire w_dff_B_nZrOZltL0_2;
	wire w_dff_B_etKkFuI77_2;
	wire w_dff_B_1fFlJiSp1_2;
	wire w_dff_B_Ttqu1gge7_2;
	wire w_dff_B_P0vgnwCv1_2;
	wire w_dff_B_voaJivia8_2;
	wire w_dff_B_Kk9wTNeM2_2;
	wire w_dff_B_18GxfdaB7_2;
	wire w_dff_B_LyHkaUR49_2;
	wire w_dff_B_oIOR0dmo3_2;
	wire w_dff_B_Iz8tKzEp8_2;
	wire w_dff_B_shPZTjE78_2;
	wire w_dff_B_A68aUUPC3_2;
	wire w_dff_B_jhc8pLKm4_2;
	wire w_dff_B_U9JniUaH8_2;
	wire w_dff_B_oJdtqV5z9_2;
	wire w_dff_B_aYCWcGSM8_2;
	wire w_dff_B_COra2qfM4_2;
	wire w_dff_B_7UCxlYQc8_2;
	wire w_dff_B_Z1zRk0uY1_2;
	wire w_dff_B_o9ACfJgY0_1;
	wire w_dff_B_cPOEvITt8_1;
	wire w_dff_B_XGwvc5G29_1;
	wire w_dff_B_o8h1KEpz0_1;
	wire w_dff_B_FhFui9Xf6_1;
	wire w_dff_B_3RwaW1OU2_1;
	wire w_dff_B_qiqCAw8V7_1;
	wire w_dff_B_KkPLgnen0_1;
	wire w_dff_B_Z9C3wXrT3_1;
	wire w_dff_B_cQs5ZD5z6_1;
	wire w_dff_B_axl2M9jY6_1;
	wire w_dff_B_d8alS8uA0_0;
	wire w_dff_B_5sHni9tO0_0;
	wire w_dff_B_1SUwnsbX8_0;
	wire w_dff_B_mLEFg69p4_0;
	wire w_dff_B_j4DcIPp68_0;
	wire w_dff_B_R1K5cPig8_0;
	wire w_dff_B_so0dxkMW6_0;
	wire w_dff_B_iEzwuLDR8_0;
	wire w_dff_B_3jds2xVB2_0;
	wire w_dff_B_SRiaM2L53_0;
	wire w_dff_A_7VKAsHle8_1;
	wire w_dff_A_UZY1CrhJ1_1;
	wire w_dff_A_ViV3GljL8_1;
	wire w_dff_A_bcsj0KjH5_1;
	wire w_dff_A_ijZFIdMx3_1;
	wire w_dff_A_0YRQSRgp9_1;
	wire w_dff_A_guFOqtuK1_1;
	wire w_dff_A_87hGvDmh0_1;
	wire w_dff_A_Y9aOEV3y0_1;
	wire w_dff_A_YWfTYHQ56_1;
	wire w_dff_A_0qrSNxvr5_1;
	wire w_dff_B_YEAzskLF4_1;
	wire w_dff_B_rMusndVY0_1;
	wire w_dff_B_5gi6yClv4_1;
	wire w_dff_B_ZmqVvHfH9_1;
	wire w_dff_B_V4WhLO7C5_1;
	wire w_dff_B_BQPEx8m24_1;
	wire w_dff_B_3kphcJ8Y9_1;
	wire w_dff_B_LZt5y3kR9_1;
	wire w_dff_B_YEMg0A4Q4_1;
	wire w_dff_B_6Hr1ygcP3_1;
	wire w_dff_B_bXC1YG0R2_1;
	wire w_dff_B_ianbkAXR0_0;
	wire w_dff_B_BwzHQZTA6_0;
	wire w_dff_B_0fFYEaoK5_0;
	wire w_dff_B_pdEzTE1M5_0;
	wire w_dff_B_EvVAsKtu6_0;
	wire w_dff_B_7A4DT3zN2_0;
	wire w_dff_B_qB0lheFZ7_0;
	wire w_dff_B_SoNZnL051_0;
	wire w_dff_B_67VTckUz2_0;
	wire w_dff_B_E29MaRkv1_0;
	wire w_dff_A_Mj40EOBe6_1;
	wire w_dff_A_bsSvo46Y5_1;
	wire w_dff_A_HkR7Ylcm6_1;
	wire w_dff_A_F3AxsMFG9_1;
	wire w_dff_A_U20mPH2w6_1;
	wire w_dff_A_H8pWA1CF4_1;
	wire w_dff_A_yAmQbFP07_1;
	wire w_dff_A_sKtmNH8T0_1;
	wire w_dff_A_xDVMtuT66_1;
	wire w_dff_A_ScOg4b7Q9_1;
	wire w_dff_A_eIaV6tH83_1;
	wire w_dff_B_5YvjGBAs8_1;
	wire w_dff_B_8UiDUOn22_1;
	wire w_dff_B_bZ1rNLCr2_1;
	wire w_dff_B_ONt2Z9LH7_1;
	wire w_dff_B_t39CgGCb0_1;
	wire w_dff_B_zL86rSCx0_1;
	wire w_dff_B_q5XuGfCR8_1;
	wire w_dff_B_G55bmCv26_1;
	wire w_dff_B_Eh9dYSzZ7_1;
	wire w_dff_B_d9jDqZ8E4_1;
	wire w_dff_B_7um8b3989_1;
	wire w_dff_B_749dpsfz8_0;
	wire w_dff_B_skbY2O4v8_0;
	wire w_dff_B_DMlJozVD5_0;
	wire w_dff_B_fhmqYWYx6_0;
	wire w_dff_B_GzG1hbKr7_0;
	wire w_dff_B_UidKZxkQ4_0;
	wire w_dff_B_1dzjzpZw2_0;
	wire w_dff_B_e3bYoBsL9_0;
	wire w_dff_B_MMAW9hxB9_0;
	wire w_dff_B_sqeRZOro5_0;
	wire w_dff_A_mswBxS1X9_1;
	wire w_dff_A_UeLFYQ4b1_1;
	wire w_dff_A_TYKipJmp5_1;
	wire w_dff_A_YL9q3rcN2_1;
	wire w_dff_A_b5X0aJG49_1;
	wire w_dff_A_Ok1SW55K5_1;
	wire w_dff_A_t08ZGmFO9_1;
	wire w_dff_A_xhE2jIkx8_1;
	wire w_dff_A_xAT2xVsN4_1;
	wire w_dff_A_drFri1Aq6_1;
	wire w_dff_A_IoAnXfgU6_1;
	wire w_dff_B_arrQLrjA0_1;
	wire w_dff_B_wdj2zzep9_1;
	wire w_dff_B_cv8hbwiA3_1;
	wire w_dff_B_mBMwSrKI0_1;
	wire w_dff_B_ZNrIb3Ob7_1;
	wire w_dff_B_62OmB0kE6_1;
	wire w_dff_B_TC6QIwv07_1;
	wire w_dff_B_yQECvr7t1_1;
	wire w_dff_B_DYxvsUTe6_1;
	wire w_dff_B_bg5QWs855_1;
	wire w_dff_B_yshrl5Ud5_1;
	wire w_dff_B_2rU6hWhb0_0;
	wire w_dff_B_gCDpAbbi9_0;
	wire w_dff_B_4h9QGvdW3_0;
	wire w_dff_B_syhtqtz50_0;
	wire w_dff_B_DhS074Qe9_0;
	wire w_dff_B_rfxAJ5Yw9_0;
	wire w_dff_B_OkSZCMOR4_0;
	wire w_dff_B_OCfgNTLu2_0;
	wire w_dff_B_61oQJSTp8_0;
	wire w_dff_B_W6zUBB6O9_0;
	wire w_dff_A_mxwr8UYm7_1;
	wire w_dff_A_IFCPKTSb9_1;
	wire w_dff_A_t0TQDQ423_1;
	wire w_dff_A_Btn4SYhf5_1;
	wire w_dff_A_4uPoGXNf8_1;
	wire w_dff_A_kps6M7715_1;
	wire w_dff_A_tqWCwPQ50_1;
	wire w_dff_A_aFTLbqF16_1;
	wire w_dff_A_B98nMDlS7_1;
	wire w_dff_A_cOOiRZiJ6_1;
	wire w_dff_A_3bR1yH9e9_1;
	wire w_dff_B_WnJUfAew8_1;
	wire w_dff_B_Kj1H0aPJ0_1;
	wire w_dff_B_L7PzYaCk1_1;
	wire w_dff_B_TYZClh2K1_1;
	wire w_dff_B_0u6ciJRm1_1;
	wire w_dff_B_2lCvsLXn6_1;
	wire w_dff_B_DjyO0dHN9_1;
	wire w_dff_B_UJGNFLuM7_1;
	wire w_dff_B_fWiL7Xtt8_1;
	wire w_dff_B_q2RjPvxV1_1;
	wire w_dff_B_XjLyrqrv9_1;
	wire w_dff_B_dC54bDG36_0;
	wire w_dff_B_YhLA8U5Y5_0;
	wire w_dff_B_EOwbEmdX9_0;
	wire w_dff_B_XE0L8f0U6_0;
	wire w_dff_B_5gv2pbhi4_0;
	wire w_dff_B_cekxpdly7_0;
	wire w_dff_B_pL8ykWlX0_0;
	wire w_dff_B_46e03LDC6_0;
	wire w_dff_B_5CmIey8H7_0;
	wire w_dff_A_u380fZG16_1;
	wire w_dff_A_dayGIxwK3_1;
	wire w_dff_A_nnaOHHwf3_1;
	wire w_dff_A_RLPkLiQf4_1;
	wire w_dff_A_mF3z3wDM0_1;
	wire w_dff_A_gtl5zLcf6_1;
	wire w_dff_A_rEqRhFPT8_1;
	wire w_dff_A_KnR9i2lp7_1;
	wire w_dff_A_FDqqWS4F2_1;
	wire w_dff_A_4SVq3Cyq9_1;
	wire w_dff_B_MsVoWa3L2_1;
	wire w_dff_B_60a7kRpr4_1;
	wire w_dff_B_Np9BxNl36_1;
	wire w_dff_B_XlZxtOUp8_1;
	wire w_dff_B_aAK0I0uV1_1;
	wire w_dff_B_YioF7NQx9_1;
	wire w_dff_B_0Px2zpau2_1;
	wire w_dff_B_vY0YaZ6a4_1;
	wire w_dff_B_4qelXxch3_1;
	wire w_dff_B_mtlvViN33_1;
	wire w_dff_B_liyKuP360_0;
	wire w_dff_B_szUbbBuD2_0;
	wire w_dff_B_sQKoR2ul9_0;
	wire w_dff_B_jsPi28bt0_0;
	wire w_dff_B_n3mW5Eo46_0;
	wire w_dff_B_BlcJPBFe0_0;
	wire w_dff_B_6UsnmYeN3_0;
	wire w_dff_B_Tze7IZDs2_0;
	wire w_dff_A_hkeAjjSB2_1;
	wire w_dff_A_8YjD7zZi1_1;
	wire w_dff_A_5lkyAW9x8_1;
	wire w_dff_A_xBHAMgpt6_1;
	wire w_dff_A_HDJofp8d4_1;
	wire w_dff_A_KwCiN0Sy0_1;
	wire w_dff_A_Hhxneuyj6_1;
	wire w_dff_A_hzYJS89d0_1;
	wire w_dff_A_PseeWV7o8_1;
	wire w_dff_B_a7YIOk8M8_1;
	wire w_dff_B_dZbbqaue6_1;
	wire w_dff_B_o19TEuSk0_1;
	wire w_dff_B_LU2YWc9d6_1;
	wire w_dff_B_SAjuZs1F7_1;
	wire w_dff_B_kAZFaCcr0_1;
	wire w_dff_B_dhgKUgDp9_1;
	wire w_dff_B_vZYIiGeW8_1;
	wire w_dff_B_osgi03YI5_1;
	wire w_dff_B_ARhsUsw33_1;
	wire w_dff_B_eqChqEf42_0;
	wire w_dff_B_9xaitLE90_0;
	wire w_dff_B_5vca0cLj1_0;
	wire w_dff_B_hxYnyNWb0_0;
	wire w_dff_B_inrFCRUM7_0;
	wire w_dff_B_eOcvstmW6_0;
	wire w_dff_B_32WcYKRw9_0;
	wire w_dff_B_6YQoVxFh5_0;
	wire w_dff_A_mA5lx3FM3_1;
	wire w_dff_A_taLSbNYm3_1;
	wire w_dff_A_DRq3fT7G6_1;
	wire w_dff_A_dofAhVII2_1;
	wire w_dff_A_hfR7aPfM0_1;
	wire w_dff_A_SkuTR7Ef7_1;
	wire w_dff_A_FJjl9Pkl0_1;
	wire w_dff_A_uRC3vwxj8_1;
	wire w_dff_A_9NTLJcnU8_1;
	wire w_dff_B_H92v0Rrm3_1;
	wire w_dff_B_8B6yT9DT0_1;
	wire w_dff_B_kG9W971c6_1;
	wire w_dff_B_ezsMz3ps2_1;
	wire w_dff_B_bQtBB8yb6_1;
	wire w_dff_B_N1gPcbpr7_1;
	wire w_dff_B_Xd7nkYJJ5_1;
	wire w_dff_B_EAv8BngY7_1;
	wire w_dff_B_hhXVJfRN7_0;
	wire w_dff_B_jOg8jmyr1_0;
	wire w_dff_B_ASlbXrhA5_0;
	wire w_dff_B_XW7fl4cO5_0;
	wire w_dff_B_htQ0YOcZ4_0;
	wire w_dff_B_m0hmfefD1_0;
	wire w_dff_A_GarCRriD1_1;
	wire w_dff_A_TA1hEKgS4_1;
	wire w_dff_A_Qn41WNQI1_1;
	wire w_dff_A_IsTiWrYf3_1;
	wire w_dff_A_daiH8hST4_1;
	wire w_dff_A_OWyDLyKj7_1;
	wire w_dff_A_xmslFCKQ7_1;
	wire w_dff_B_atpQrkQn9_1;
	wire w_dff_B_s36uqheW1_1;
	wire w_dff_B_JFKjl0bP0_1;
	wire w_dff_B_mcZUAll60_1;
	wire w_dff_B_FnujWyla8_1;
	wire w_dff_B_D2ZhCCaW9_1;
	wire w_dff_B_KasjwAkM9_1;
	wire w_dff_B_6kN2imgs3_0;
	wire w_dff_B_EiultIJq1_0;
	wire w_dff_B_aE74eXWs0_0;
	wire w_dff_B_23oOUYVq6_0;
	wire w_dff_B_cotjRpX83_0;
	wire w_dff_A_rMpQbARe6_1;
	wire w_dff_A_HBMx0F6Y6_1;
	wire w_dff_A_acFAoB715_1;
	wire w_dff_A_gELSl4NY6_1;
	wire w_dff_A_pc60ZrUb1_1;
	wire w_dff_A_njEHyu7l3_1;
	wire w_dff_B_q05ACBSj4_1;
	wire w_dff_B_xZx0QW7B2_1;
	wire w_dff_B_fWrkI66s4_1;
	wire w_dff_B_GlgzqquN0_1;
	wire w_dff_B_w0BcUHRx3_1;
	wire w_dff_B_0wQXfKuk2_1;
	wire w_dff_B_d1g90P6Y5_0;
	wire w_dff_B_CpLBWBme5_0;
	wire w_dff_B_YpiA6JQf3_0;
	wire w_dff_B_w6qGUp2q7_0;
	wire w_dff_A_qRWrLJHO5_1;
	wire w_dff_A_rLQ3MIbx8_1;
	wire w_dff_A_wshycQhA0_1;
	wire w_dff_A_PZSan8Hh2_1;
	wire w_dff_A_vT4dEFkO3_1;
	wire w_dff_B_TneMuxcJ0_1;
	wire w_dff_B_R5r31NiQ5_1;
	wire w_dff_B_W6JW4JY46_1;
	wire w_dff_A_hPDweS9h2_0;
	wire w_dff_A_GY0tRlvX7_0;
	wire w_dff_B_BBetNlil1_1;
	wire w_dff_A_3F2qeiCQ3_0;
	wire w_dff_B_OmGa2UCE3_1;
	wire w_dff_A_hrBreWcA4_1;
	wire w_dff_B_k77NgaMe2_2;
	wire w_dff_B_2Jd0iHVW5_1;
	wire w_dff_A_XztLsaWI3_0;
	wire w_dff_A_xnlAbdHd7_0;
	wire w_dff_A_IZBE0o1x6_0;
	wire w_dff_A_WYzqc2nb3_0;
	wire w_dff_A_rMekzOQB9_0;
	wire w_dff_A_2uvANXjR1_0;
	wire w_dff_A_GKRicQKM4_0;
	wire w_dff_A_iK5LrSOU7_0;
	wire w_dff_A_HtoL1htq2_0;
	wire w_dff_A_giro5rPs9_0;
	wire w_dff_A_TNBabMUo3_0;
	wire w_dff_A_UQiFp3kU6_0;
	wire w_dff_A_YxTF7zei4_0;
	wire w_dff_A_uQYrV3Kw3_0;
	wire w_dff_A_dzzTosjp0_0;
	wire w_dff_A_lJw1AJoj7_0;
	wire w_dff_A_uCWYDUEs9_0;
	wire w_dff_A_UrefqLHB0_0;
	wire w_dff_A_QqBQw9H95_0;
	wire w_dff_A_iUYgljVi1_0;
	wire w_dff_A_tQvnKtQ70_0;
	wire w_dff_A_oPVbxvsv2_0;
	wire w_dff_A_itqnddGD8_0;
	wire w_dff_A_3JlSNcIc5_0;
	wire w_dff_A_raRNB5ki5_0;
	wire w_dff_A_5WqZGXYg5_0;
	wire w_dff_A_dewhXr0h6_0;
	wire w_dff_A_QSqF0f3R4_0;
	wire w_dff_A_cXIP6Qxb4_0;
	wire w_dff_A_veMi3zVL4_0;
	wire w_dff_A_W5I2SHU40_0;
	wire w_dff_A_W8t6BoxU0_0;
	wire w_dff_A_1fyNjCk01_0;
	wire w_dff_A_9PvjUJ8f1_0;
	wire w_dff_A_qYzi9ijr9_0;
	wire w_dff_A_M1TmlG254_0;
	wire w_dff_A_5G5kckfl5_0;
	wire w_dff_A_mPZQ5b8e5_0;
	wire w_dff_A_MqVzcWX48_0;
	wire w_dff_A_Iu5dIaPF2_0;
	wire w_dff_A_bqv7GY0M5_0;
	wire w_dff_A_S72Wv5Nx9_0;
	wire w_dff_A_z6gwAQrs2_0;
	wire w_dff_A_UeowzV526_0;
	wire w_dff_A_hQoEVyXq2_1;
	wire w_dff_B_WgXmBxuA8_1;
	wire w_dff_A_PiiIzt3R8_0;
	wire w_dff_A_I6e6MBN94_0;
	wire w_dff_A_DI0hUnOy4_0;
	wire w_dff_A_j2gyYtOg8_0;
	wire w_dff_A_FUuFRAB05_0;
	wire w_dff_A_PC4p1H1m1_0;
	wire w_dff_A_ff5HL2R95_0;
	wire w_dff_A_Ed77mGnc4_0;
	wire w_dff_A_BJEJ6zXE4_0;
	wire w_dff_A_Rw5MsoPp1_0;
	wire w_dff_A_vt7VItj09_0;
	wire w_dff_A_2ikhUUUE6_0;
	wire w_dff_A_9vdDxUv13_0;
	wire w_dff_A_B3Q9oF6k0_0;
	wire w_dff_A_bKwww85G7_0;
	wire w_dff_A_2b9e82EN5_0;
	wire w_dff_A_P19Sqdo77_0;
	wire w_dff_A_SZzxIYQ15_0;
	wire w_dff_A_cB4yQMR73_0;
	wire w_dff_A_c0vytwfD9_0;
	wire w_dff_A_c8KSx1ND0_0;
	wire w_dff_A_JiHQIVAM4_0;
	wire w_dff_A_kYty4V296_0;
	wire w_dff_A_RojqhZIA9_0;
	wire w_dff_A_wP5F6fzZ2_0;
	wire w_dff_A_QZY8CUOS1_0;
	wire w_dff_A_jGHnAh5L7_0;
	wire w_dff_A_nXyRtF1i2_0;
	wire w_dff_A_XwPGBhfq3_0;
	wire w_dff_A_222ylpW08_0;
	wire w_dff_A_NuBlYdaU7_0;
	wire w_dff_A_iqjfqWP06_0;
	wire w_dff_A_6NZ3krYe9_0;
	wire w_dff_A_3pOUc97J3_0;
	wire w_dff_A_dp2Y069B6_0;
	wire w_dff_A_t8XThZsf8_0;
	wire w_dff_A_oz8NCmJL2_0;
	wire w_dff_A_9CdNR69I7_0;
	wire w_dff_A_L1XzuGHU3_0;
	wire w_dff_A_WhIZKAjF7_0;
	wire w_dff_A_v4PrTfen7_0;
	wire w_dff_A_ls7XPJqC5_1;
	wire w_dff_B_8VzzC10B8_1;
	wire w_dff_B_lW2Bhz3d1_1;
	wire w_dff_B_GszznvkK5_1;
	wire w_dff_B_dIqA0EZB7_1;
	wire w_dff_B_IjjNUSPc6_1;
	wire w_dff_B_kNGsYjop5_1;
	wire w_dff_B_B1YHmoVt1_1;
	wire w_dff_B_Bblgcefy8_1;
	wire w_dff_B_5op6F0yd7_1;
	wire w_dff_B_m0G09LZF4_1;
	wire w_dff_B_Qi8aYOEC6_1;
	wire w_dff_B_kCqh92Sm3_1;
	wire w_dff_B_qPkrqY9x8_1;
	wire w_dff_B_Df7brTSZ1_1;
	wire w_dff_B_dsPxwSMv0_1;
	wire w_dff_B_1aRYIuQ52_1;
	wire w_dff_B_A610nrWP2_1;
	wire w_dff_B_gGKQdiBh5_1;
	wire w_dff_B_qEuix4A42_1;
	wire w_dff_B_d1zF20rF8_1;
	wire w_dff_B_gf3e94Nk0_1;
	wire w_dff_B_e084yyqQ9_1;
	wire w_dff_B_pKqFTqWp9_1;
	wire w_dff_B_9pu5oilm6_1;
	wire w_dff_B_7q7EsWDB4_1;
	wire w_dff_B_idov8ouX8_1;
	wire w_dff_B_anLHWe976_1;
	wire w_dff_B_XJxIqut58_1;
	wire w_dff_B_0oEBqDHD6_1;
	wire w_dff_B_5uNkM3F92_1;
	wire w_dff_B_Y3RneUl01_1;
	wire w_dff_B_z0sf1KzW4_1;
	wire w_dff_B_uHKisNI68_1;
	wire w_dff_B_YMFs8YlH7_1;
	wire w_dff_B_hkwLdqAe5_1;
	wire w_dff_B_sig7arG82_1;
	wire w_dff_B_xjv428pr0_1;
	wire w_dff_B_DpzuuPns0_1;
	wire w_dff_A_nA9jw31B6_0;
	wire w_dff_A_23tyB7qe4_0;
	wire w_dff_A_XwaEOSLh7_0;
	wire w_dff_A_vE5fslys9_0;
	wire w_dff_A_6YvIlmwi6_0;
	wire w_dff_A_YYyqgfnK7_0;
	wire w_dff_A_2EN1hU2K0_0;
	wire w_dff_A_hzwtpl9Z3_0;
	wire w_dff_A_90gH4jFa1_0;
	wire w_dff_A_FgzVbrpY4_0;
	wire w_dff_A_1XcERHTm8_0;
	wire w_dff_A_wBvetjQi4_0;
	wire w_dff_A_ZgbRKsPe0_0;
	wire w_dff_A_fjrB3MRu2_0;
	wire w_dff_A_4viJ7sGW2_0;
	wire w_dff_A_ZWMKS3Hy3_0;
	wire w_dff_A_mjQvio0T8_0;
	wire w_dff_A_kLFRzyFN5_0;
	wire w_dff_A_mWy1c4T31_0;
	wire w_dff_A_HCg9oAAy7_0;
	wire w_dff_A_djxzIVmo4_0;
	wire w_dff_A_R5abQt844_0;
	wire w_dff_A_CmWCl49J9_0;
	wire w_dff_A_z0bjo0uP4_0;
	wire w_dff_A_JXVj8edD7_0;
	wire w_dff_A_fyaOQ5gL1_0;
	wire w_dff_A_i7Zvo5oI9_0;
	wire w_dff_A_1t8sO5HL6_0;
	wire w_dff_A_q8C2996N9_0;
	wire w_dff_A_WzsIyWS02_0;
	wire w_dff_A_UKKkdDDR4_0;
	wire w_dff_A_LVFMzPm42_0;
	wire w_dff_A_5IrwuyqO3_0;
	wire w_dff_A_LXmC66Bo0_0;
	wire w_dff_A_WusR1u5e7_0;
	wire w_dff_A_gSX6UWhN7_0;
	wire w_dff_A_Jb2z1ag75_0;
	wire w_dff_A_evevrTmx4_0;
	wire w_dff_A_90iIDhbQ1_1;
	wire w_dff_B_8GwMWOwi5_1;
	wire w_dff_B_wjSGixRt4_1;
	wire w_dff_B_PfTadJ1a7_1;
	wire w_dff_B_xbIpS5bo9_1;
	wire w_dff_B_rjAWUfle1_1;
	wire w_dff_B_3hSQSrmw5_1;
	wire w_dff_B_IGCzFkC48_1;
	wire w_dff_B_TTqoxdy02_1;
	wire w_dff_B_EbOVk6836_1;
	wire w_dff_B_Nd3oec7e5_1;
	wire w_dff_B_aK7nwTNr0_1;
	wire w_dff_B_mBYciLTO1_1;
	wire w_dff_B_LZfPGB4O3_1;
	wire w_dff_B_PkFReVkE7_1;
	wire w_dff_B_8E8txXkl3_1;
	wire w_dff_B_rk4MerAO0_1;
	wire w_dff_B_1B0G0wJu3_1;
	wire w_dff_B_Ypa3paFi0_1;
	wire w_dff_B_BepEl4gS3_1;
	wire w_dff_B_zw0CxJy35_1;
	wire w_dff_B_XCArx3YC5_1;
	wire w_dff_B_Tfpplh7L3_1;
	wire w_dff_B_npfMN3jQ8_1;
	wire w_dff_B_zcm2AJ8X1_1;
	wire w_dff_B_TJysLcki0_1;
	wire w_dff_B_ATal7wO17_1;
	wire w_dff_B_V5qXykAA4_1;
	wire w_dff_B_AwxioecJ7_1;
	wire w_dff_B_m0V5luZO3_1;
	wire w_dff_B_G3AF7vZ51_1;
	wire w_dff_B_FhKe6taQ1_1;
	wire w_dff_B_FxSvqxgM2_1;
	wire w_dff_B_0FnM0RF66_1;
	wire w_dff_B_ecnqGgPb9_1;
	wire w_dff_B_y1OoywVh9_1;
	wire w_dff_A_wjHhreBH5_0;
	wire w_dff_A_kHIIfzcz3_0;
	wire w_dff_A_pNw3Vfkk7_0;
	wire w_dff_A_CuI1nMiy9_0;
	wire w_dff_A_WjdbFQ856_0;
	wire w_dff_A_8FPxcX2V4_0;
	wire w_dff_A_6V0mvtf37_0;
	wire w_dff_A_eCAGxrrg2_0;
	wire w_dff_A_ltU7wmsA2_0;
	wire w_dff_A_2xJ5iN1W9_0;
	wire w_dff_A_sSc3NPIN9_0;
	wire w_dff_A_vbGXJaMS9_0;
	wire w_dff_A_CMML3V2z0_0;
	wire w_dff_A_ka4veQaB0_0;
	wire w_dff_A_uBByO3HM8_0;
	wire w_dff_A_pWQUe7gN1_0;
	wire w_dff_A_rw4GaEQf6_0;
	wire w_dff_A_asnyFLVr1_0;
	wire w_dff_A_Iwagun5z0_0;
	wire w_dff_A_QjD8yeB65_0;
	wire w_dff_A_i8nJWRvf8_0;
	wire w_dff_A_XOYjXaGu2_0;
	wire w_dff_A_Efev6IZb6_0;
	wire w_dff_A_oRSD7Bg98_0;
	wire w_dff_A_4Ew5CFO26_0;
	wire w_dff_A_s9G4wvIg4_0;
	wire w_dff_A_rfCgWFzs2_0;
	wire w_dff_A_GCa1fvs20_0;
	wire w_dff_A_6ZEIhEwW2_0;
	wire w_dff_A_H1nUe7rP0_0;
	wire w_dff_A_jSl38lnw2_0;
	wire w_dff_A_SP3GChog1_0;
	wire w_dff_A_S0GLViYs8_0;
	wire w_dff_A_hrtsktC32_0;
	wire w_dff_A_aYONlrSn6_0;
	wire w_dff_A_XitmDLyL7_1;
	wire w_dff_B_bQKhF1F47_1;
	wire w_dff_B_vjuSIyUB2_1;
	wire w_dff_B_PcHPSCLQ2_1;
	wire w_dff_B_QdtqTTb28_1;
	wire w_dff_B_qXnzfyTX4_1;
	wire w_dff_B_qIzEorvX0_1;
	wire w_dff_B_nL0F2n6x6_1;
	wire w_dff_B_yvW3kLcj1_1;
	wire w_dff_B_fFf8iiWK8_1;
	wire w_dff_B_RLagDZks1_1;
	wire w_dff_B_Ut3jzycM5_1;
	wire w_dff_B_doUVHaHM0_1;
	wire w_dff_B_p50seZT68_1;
	wire w_dff_B_U9Ml2wZm5_1;
	wire w_dff_B_MREcElIB3_1;
	wire w_dff_B_YW9BFBrY3_1;
	wire w_dff_B_mHPEN9Xj0_1;
	wire w_dff_B_5br7u1YE9_1;
	wire w_dff_B_rW3gkcug8_1;
	wire w_dff_B_VpOX9ND18_1;
	wire w_dff_B_RnKFdvZv0_1;
	wire w_dff_B_4BS9jKbC4_1;
	wire w_dff_B_tOPjf5nt5_1;
	wire w_dff_B_hblLleH77_1;
	wire w_dff_B_6OcBKw6m0_1;
	wire w_dff_B_buaxEEK13_1;
	wire w_dff_B_rFvh3htF3_1;
	wire w_dff_B_9Yvcven91_1;
	wire w_dff_B_8cNmkGp30_1;
	wire w_dff_B_M7jHNoC75_1;
	wire w_dff_B_Ga7CVoxM6_1;
	wire w_dff_B_XVNnUZs48_1;
	wire w_dff_A_cup175MQ3_0;
	wire w_dff_A_VGGhTwsL0_0;
	wire w_dff_A_8JxtuMRC3_0;
	wire w_dff_A_p7tuihX95_0;
	wire w_dff_A_PbganX0l8_0;
	wire w_dff_A_WDaqGhkC0_0;
	wire w_dff_A_f0j3Hkkh9_0;
	wire w_dff_A_9hW3Rs4c1_0;
	wire w_dff_A_pAF6pTS79_0;
	wire w_dff_A_SJTcTBc30_0;
	wire w_dff_A_68QkYdto2_0;
	wire w_dff_A_ILiET0zh3_0;
	wire w_dff_A_ZO5bSGG75_0;
	wire w_dff_A_3u8TvXnr2_0;
	wire w_dff_A_H2nB6pCw4_0;
	wire w_dff_A_RZTEJqO27_0;
	wire w_dff_A_JoNuCgjT2_0;
	wire w_dff_A_qL8ypbtA8_0;
	wire w_dff_A_2aoblbmy5_0;
	wire w_dff_A_OhyDLvdh6_0;
	wire w_dff_A_iSskpdNs3_0;
	wire w_dff_A_hQfPfrTh2_0;
	wire w_dff_A_u0aQlJdh3_0;
	wire w_dff_A_DOmuxUPB5_0;
	wire w_dff_A_GuuIyRFy5_0;
	wire w_dff_A_1DyrCIQR3_0;
	wire w_dff_A_Sz2mTKNr3_0;
	wire w_dff_A_7RPHRJMB6_0;
	wire w_dff_A_Yngj7ojn7_0;
	wire w_dff_A_VegrjOOJ0_0;
	wire w_dff_A_GpCWbGKG9_0;
	wire w_dff_A_YKx6JKpo5_0;
	wire w_dff_A_J8sheeoS5_1;
	wire w_dff_B_jrF5iNMt4_1;
	wire w_dff_B_hMXa6umq4_1;
	wire w_dff_B_33VFdYq93_1;
	wire w_dff_B_CqaD6UHH1_1;
	wire w_dff_B_UfUEr0xq4_1;
	wire w_dff_B_pQzfiOQg9_1;
	wire w_dff_B_D8CY7Prf3_1;
	wire w_dff_B_iQni8Os93_1;
	wire w_dff_B_4JPkIfmu0_1;
	wire w_dff_B_gPMIkARU2_1;
	wire w_dff_B_jv1RGV173_1;
	wire w_dff_B_uskEw4QF4_1;
	wire w_dff_B_NIyWbGYb4_1;
	wire w_dff_B_mpsZPCTS8_1;
	wire w_dff_B_66iPT5vT4_1;
	wire w_dff_B_m0XG0Q223_1;
	wire w_dff_B_1TFWPF3C5_1;
	wire w_dff_B_a6UUGYvC2_1;
	wire w_dff_B_zTNQmmtu5_1;
	wire w_dff_B_TfPXk9OU3_1;
	wire w_dff_B_wkDuxIzr9_1;
	wire w_dff_B_ds9l8EH26_1;
	wire w_dff_B_nbv2E0wK9_1;
	wire w_dff_B_7sfGItpL4_1;
	wire w_dff_B_lkAEWT7l6_1;
	wire w_dff_B_9MUXxqf55_1;
	wire w_dff_B_IwBOIOfu2_1;
	wire w_dff_B_i7Y5QUbp9_1;
	wire w_dff_B_Sas486Fy7_1;
	wire w_dff_A_clNM4O544_0;
	wire w_dff_A_FRDKW83e5_0;
	wire w_dff_A_2pubCDBU9_0;
	wire w_dff_A_u6cC8iEo2_0;
	wire w_dff_A_bihMRFSc1_0;
	wire w_dff_A_Tp5ukWrU6_0;
	wire w_dff_A_PQHBQeQ88_0;
	wire w_dff_A_6hKGXp2n6_0;
	wire w_dff_A_2hLXjuSt9_0;
	wire w_dff_A_VT9uk01s8_0;
	wire w_dff_A_ba218ma79_0;
	wire w_dff_A_LH6i8iDf7_0;
	wire w_dff_A_k0fnviVx3_0;
	wire w_dff_A_pcNzs3g52_0;
	wire w_dff_A_SKeRgjCD9_0;
	wire w_dff_A_DlXmu2b54_0;
	wire w_dff_A_IcQ1nQXP5_0;
	wire w_dff_A_9j7mjvKU0_0;
	wire w_dff_A_isWUtwEk6_0;
	wire w_dff_A_c2KFI1wt8_0;
	wire w_dff_A_zUYihYQ72_0;
	wire w_dff_A_S80ML2T33_0;
	wire w_dff_A_2kzZNoJ95_0;
	wire w_dff_A_uwNEA9JR7_0;
	wire w_dff_A_zMfLwwtg2_0;
	wire w_dff_A_MKBp2C5v8_0;
	wire w_dff_A_nLBL5pzN6_0;
	wire w_dff_A_YLBwudag3_0;
	wire w_dff_A_R4ZeTc807_0;
	wire w_dff_A_q8tDLDGG5_1;
	wire w_dff_B_ZL5VaW9n3_1;
	wire w_dff_B_JsJNkWNH7_1;
	wire w_dff_B_dEhn0jED6_1;
	wire w_dff_B_7dYbH2lr6_1;
	wire w_dff_B_WAvn0rNU6_1;
	wire w_dff_B_2qcrzXlP2_1;
	wire w_dff_B_qqCwWwgw5_1;
	wire w_dff_B_D7WDdV4b2_1;
	wire w_dff_B_Vfe8ybqM6_1;
	wire w_dff_B_Vm90iu193_1;
	wire w_dff_B_gplyiiRe7_1;
	wire w_dff_B_tPqXlddp7_1;
	wire w_dff_B_KIn84tUX8_1;
	wire w_dff_B_gdAerqbx6_1;
	wire w_dff_B_X6cvKOX49_1;
	wire w_dff_B_QauYEzdS0_1;
	wire w_dff_B_dftS0TZo7_1;
	wire w_dff_B_1q90oM0k9_1;
	wire w_dff_B_AoFvBdpB5_1;
	wire w_dff_B_KFqcFrUX6_1;
	wire w_dff_B_RRU6Zs145_1;
	wire w_dff_B_WPcY44fS0_1;
	wire w_dff_B_UlbgQ8MC5_1;
	wire w_dff_B_gzwSsxYP3_1;
	wire w_dff_B_vfMFIONK9_1;
	wire w_dff_B_r79Ag4N17_1;
	wire w_dff_A_07XvEf3d4_0;
	wire w_dff_A_S71DeJ4S7_0;
	wire w_dff_A_AyP7AboR5_0;
	wire w_dff_A_1RfPkj7S2_0;
	wire w_dff_A_3JrGAypj5_0;
	wire w_dff_A_SGAlmRUy8_0;
	wire w_dff_A_vRWkMEVA7_0;
	wire w_dff_A_eYZc56bQ0_0;
	wire w_dff_A_AL1Jq1aZ1_0;
	wire w_dff_A_tiCsG0FA5_0;
	wire w_dff_A_ZM8KHHC41_0;
	wire w_dff_A_yG9RquUF1_0;
	wire w_dff_A_BQAGjrTr2_0;
	wire w_dff_A_VKyZLDAL4_0;
	wire w_dff_A_sXRZKFtq1_0;
	wire w_dff_A_WcV7LFru5_0;
	wire w_dff_A_KyVO6UQE1_0;
	wire w_dff_A_bADsdaOd3_0;
	wire w_dff_A_VaKaZm7P5_0;
	wire w_dff_A_iQtCWTZW2_0;
	wire w_dff_A_9rJU7ldF3_0;
	wire w_dff_A_BOGCJ2fr5_0;
	wire w_dff_A_3yB3pTCZ0_0;
	wire w_dff_A_pedVWmIY0_0;
	wire w_dff_A_rxJ6Gxda0_0;
	wire w_dff_A_KQ2O2otq9_0;
	wire w_dff_A_pdtZY1cb0_1;
	wire w_dff_B_uaji9XrL9_1;
	wire w_dff_B_V2XGEC8k2_1;
	wire w_dff_B_8ddoDOuH7_1;
	wire w_dff_B_MzbcbGUO3_1;
	wire w_dff_B_3nXnYQNm5_1;
	wire w_dff_B_3DZjDbuJ3_1;
	wire w_dff_B_zEBeWXrs6_1;
	wire w_dff_B_7u9uNGiF4_1;
	wire w_dff_B_iC2ahARG7_1;
	wire w_dff_B_B77UuNaF2_1;
	wire w_dff_B_7NcS5zV68_1;
	wire w_dff_B_6n4SH0qe0_1;
	wire w_dff_B_z1Jwm19L5_1;
	wire w_dff_B_DNVYFIAU3_1;
	wire w_dff_B_T3LTlcff9_1;
	wire w_dff_B_LHX2JYat5_1;
	wire w_dff_B_48TZ66Tv1_1;
	wire w_dff_B_RnpQ5oW77_1;
	wire w_dff_B_KQtljAQK4_1;
	wire w_dff_B_0kHpSL6g5_1;
	wire w_dff_B_cwlt9MPQ2_1;
	wire w_dff_B_9zhxnigc6_1;
	wire w_dff_B_G2a9mku59_1;
	wire w_dff_A_WNAubkdK7_0;
	wire w_dff_A_Gko9mBMh7_0;
	wire w_dff_A_PnNbR9Vs1_0;
	wire w_dff_A_4tqugQMX6_0;
	wire w_dff_A_VOBEbYy45_0;
	wire w_dff_A_PKufTHoC4_0;
	wire w_dff_A_pOyXgVy32_0;
	wire w_dff_A_EiDPqxd47_0;
	wire w_dff_A_onxi8iqR4_0;
	wire w_dff_A_36dRa3KG5_0;
	wire w_dff_A_HQNQH4wm9_0;
	wire w_dff_A_1utdlHDO5_0;
	wire w_dff_A_TOHpIvxF1_0;
	wire w_dff_A_Kujq2QhY2_0;
	wire w_dff_A_kKiCe1CS3_0;
	wire w_dff_A_AyFQGTNA1_0;
	wire w_dff_A_gIufiRDE7_0;
	wire w_dff_A_YDtrAI5W8_0;
	wire w_dff_A_yoD1KkwS9_0;
	wire w_dff_A_61wkXLfz2_0;
	wire w_dff_A_M9Vj75ie0_0;
	wire w_dff_A_Yi0R7pV94_0;
	wire w_dff_A_NzASmWdC1_0;
	wire w_dff_A_ZBNkQBen1_1;
	wire w_dff_B_sQHggNVV2_1;
	wire w_dff_B_0a2EIjzn2_1;
	wire w_dff_B_g74iP5qI6_1;
	wire w_dff_B_mgLSvAeH6_1;
	wire w_dff_B_TpEiFXiZ6_1;
	wire w_dff_B_tDN3qfWj5_1;
	wire w_dff_B_3JPPXOvh9_1;
	wire w_dff_B_UtoxWck83_1;
	wire w_dff_B_2yGWQ7121_1;
	wire w_dff_B_jB9nM9qL7_1;
	wire w_dff_B_FARCtiGb1_1;
	wire w_dff_B_giBP00WZ2_1;
	wire w_dff_B_VwapzuL72_1;
	wire w_dff_B_HmBmlcBA0_1;
	wire w_dff_B_mrciLR6N7_1;
	wire w_dff_B_GSMkC0mH3_1;
	wire w_dff_B_guxh1W8Y9_1;
	wire w_dff_B_RVtFTpM18_1;
	wire w_dff_B_1NeGTeA62_1;
	wire w_dff_B_EtRKUMoM0_1;
	wire w_dff_A_yd2wSgOJ3_0;
	wire w_dff_A_dTud4PkE8_0;
	wire w_dff_A_16Otk0LG3_0;
	wire w_dff_A_VrZ2eqAD3_0;
	wire w_dff_A_394mG6D45_0;
	wire w_dff_A_CcPw8DQa1_0;
	wire w_dff_A_8zxqr1RF4_0;
	wire w_dff_A_8INlV0gl9_0;
	wire w_dff_A_B8Ldhac90_0;
	wire w_dff_A_KQZqEpd62_0;
	wire w_dff_A_PSu4PeRC0_0;
	wire w_dff_A_MxZaryhj4_0;
	wire w_dff_A_PaFBBoOj8_0;
	wire w_dff_A_2Vf80ylI8_0;
	wire w_dff_A_gFaHzqXF3_0;
	wire w_dff_A_rsFsgka31_0;
	wire w_dff_A_47xJSKVp3_0;
	wire w_dff_A_EbhXl6AE0_0;
	wire w_dff_A_mADN9N8V2_0;
	wire w_dff_A_JPXdPWUu5_0;
	wire w_dff_A_dd2KuOew4_1;
	wire w_dff_B_F1mXoP8m7_1;
	wire w_dff_B_cnK0nCHN4_1;
	wire w_dff_B_mtYEvDP34_1;
	wire w_dff_B_qzSAt64H2_1;
	wire w_dff_B_InDJSpJP6_1;
	wire w_dff_B_e9LzUf0S0_1;
	wire w_dff_B_yttmxCRk8_1;
	wire w_dff_B_3JdfAORd1_1;
	wire w_dff_B_fpJaDYb26_1;
	wire w_dff_B_RU9jkWQh0_1;
	wire w_dff_B_9u5QYrI36_1;
	wire w_dff_B_A51qYh7k0_1;
	wire w_dff_B_5wXpyIlb9_1;
	wire w_dff_B_n6hjHG9P8_1;
	wire w_dff_B_ghI2TLLK7_1;
	wire w_dff_B_2sGGj5117_1;
	wire w_dff_B_MLjx4sMy3_1;
	wire w_dff_A_jIPo6DQn7_0;
	wire w_dff_A_BEoNHnEm8_0;
	wire w_dff_A_UoeXRQNw2_0;
	wire w_dff_A_jgtar52N4_0;
	wire w_dff_A_qSSw6ntj5_0;
	wire w_dff_A_T7JiqPbL0_0;
	wire w_dff_A_tgdsUr972_0;
	wire w_dff_A_MYKZjBnC5_0;
	wire w_dff_A_X2TWBBO39_0;
	wire w_dff_A_tdEjQUA01_0;
	wire w_dff_A_rkvro7cG4_0;
	wire w_dff_A_ckoPgMau3_0;
	wire w_dff_A_FghHqTZj2_0;
	wire w_dff_A_J97Nnlbp0_0;
	wire w_dff_A_JJYQDiXV5_0;
	wire w_dff_A_6zj07BYk5_0;
	wire w_dff_A_wIZmNCxX4_0;
	wire w_dff_A_G11zUqc14_1;
	wire w_dff_B_msPiOmBT6_1;
	wire w_dff_B_9K8Fc5g41_1;
	wire w_dff_B_7Y8ID8hz4_1;
	wire w_dff_B_m7TJb8T42_1;
	wire w_dff_B_KjcKKkyc3_1;
	wire w_dff_B_XOmIvBiT7_1;
	wire w_dff_B_b4BIqd5J5_1;
	wire w_dff_B_QlSxxFjz7_1;
	wire w_dff_B_uMAiGIYJ8_1;
	wire w_dff_B_FUD1bpmc2_1;
	wire w_dff_B_whOG2x2d8_1;
	wire w_dff_B_5vO4kvi22_1;
	wire w_dff_B_TzMqASIS7_1;
	wire w_dff_B_pbsMynBF6_1;
	wire w_dff_A_1zRpXd2X4_0;
	wire w_dff_A_rMclxszd8_0;
	wire w_dff_A_X7OvdmMJ0_0;
	wire w_dff_A_pOInmols4_0;
	wire w_dff_A_LydU78NP4_0;
	wire w_dff_A_fgn7zzmi1_0;
	wire w_dff_A_3UFqp5xG1_0;
	wire w_dff_A_rbqVl4It0_0;
	wire w_dff_A_Ve2xpuXI7_0;
	wire w_dff_A_bIJGbnrZ6_0;
	wire w_dff_A_R8xzFM1X6_0;
	wire w_dff_A_WbyxWmyk1_0;
	wire w_dff_A_c8emaS972_0;
	wire w_dff_A_vuvYPKsd0_0;
	wire w_dff_A_abjFZba61_1;
	wire w_dff_B_znPVCf3g9_1;
	wire w_dff_B_uTY9VtKv1_1;
	wire w_dff_B_QvttyXg92_1;
	wire w_dff_B_ow2AcIkY8_1;
	wire w_dff_B_VsT4Cj7R0_1;
	wire w_dff_B_kPhGAsQz8_1;
	wire w_dff_B_sephocXF6_1;
	wire w_dff_B_7IqEQ2Rw3_1;
	wire w_dff_B_R7Ngk5aT2_1;
	wire w_dff_B_Y8lCDkCI6_1;
	wire w_dff_B_3eb8cAjZ3_1;
	wire w_dff_A_1yPGyo8y2_0;
	wire w_dff_A_EjRqAhi79_0;
	wire w_dff_A_JIpqIlhj3_0;
	wire w_dff_A_tzommCdL5_0;
	wire w_dff_A_LIEnoCqY8_0;
	wire w_dff_A_gHrsytin8_0;
	wire w_dff_A_fT46BE4Z8_0;
	wire w_dff_A_aFpAwGkv1_0;
	wire w_dff_A_K3J3VhNi6_0;
	wire w_dff_A_jdGnuqf83_0;
	wire w_dff_A_EVKqHyce1_0;
	wire w_dff_A_Bw9625kf4_1;
	wire w_dff_B_5lTOWi381_1;
	wire w_dff_B_nKOywrTp7_1;
	wire w_dff_B_ivFGV6Zl1_1;
	wire w_dff_B_Oeuj6ZRK6_1;
	wire w_dff_B_YknQjzgM1_1;
	wire w_dff_B_4ez6oAxy9_1;
	wire w_dff_B_z5yrB3Ls7_1;
	wire w_dff_B_xBBblVJN9_1;
	wire w_dff_A_O17b2fkp1_0;
	wire w_dff_A_Y4F5XlY71_0;
	wire w_dff_A_fUs8N7ld7_0;
	wire w_dff_A_MMsPaLNi4_0;
	wire w_dff_A_OVUgk53k2_0;
	wire w_dff_A_R6l0TgAt6_0;
	wire w_dff_A_VzizVc8V0_0;
	wire w_dff_A_kiy2BO7f5_0;
	wire w_dff_A_4iAploSe2_1;
	wire w_dff_B_xhEpL6TF3_1;
	wire w_dff_B_G4j0ydwA7_1;
	wire w_dff_B_KJVIe0q63_1;
	wire w_dff_B_Mc0qdUx74_1;
	wire w_dff_B_s2BIrOrl5_1;
	wire w_dff_B_PSo8MNph8_0;
	wire w_dff_A_TcIp6Mog2_0;
	wire w_dff_A_sRvmt9jy6_0;
	wire w_dff_A_butF18JX5_0;
	wire w_dff_A_1Eby9pJV6_0;
	wire w_dff_A_OX7nFsGl7_0;
	wire w_dff_A_x31Ir6Po7_0;
	wire w_dff_A_YDMEMreQ6_0;
	wire w_dff_A_ZxkjIyrc9_1;
	wire w_dff_B_RiwhK7vq5_1;
	wire w_dff_B_wlm8K5mf0_2;
	wire w_dff_B_9DyEIpxU0_2;
	wire w_dff_B_QOBEJ13A7_2;
	wire w_dff_B_eKOMNCZY4_2;
	wire w_dff_B_IHNDThLe2_2;
	wire w_dff_B_DO2laoWd9_2;
	wire w_dff_B_3ILXNG2K0_2;
	wire w_dff_B_XwxPcHRt9_2;
	wire w_dff_B_cWQYjVO54_2;
	wire w_dff_B_u4zv1JeY5_2;
	wire w_dff_B_Mfvhq5wL2_2;
	wire w_dff_B_7k9eOmYL7_2;
	wire w_dff_B_zqDm2X7C0_2;
	wire w_dff_B_bsSSdUYK4_2;
	wire w_dff_B_fAI1qAow0_2;
	wire w_dff_B_pDPQ9iTi9_2;
	wire w_dff_B_JjtxkxWH7_2;
	wire w_dff_B_TrlfOvVw6_2;
	wire w_dff_B_mxlSVfqZ6_2;
	wire w_dff_B_p0eQka6R1_2;
	wire w_dff_B_nuCChVu33_2;
	wire w_dff_B_M68hpCGC0_2;
	wire w_dff_B_3EgGeu4s0_2;
	wire w_dff_B_TBLieZRy2_2;
	wire w_dff_B_u2iHJdBs5_2;
	wire w_dff_B_BMsMvpkg9_2;
	wire w_dff_B_LvuS2iwE2_2;
	wire w_dff_B_2I2ldc0Q1_2;
	wire w_dff_B_ZT3XjHeo4_2;
	wire w_dff_B_bvi7awdg8_2;
	wire w_dff_B_rocixNWt1_2;
	wire w_dff_B_Su9B3HDt0_2;
	wire w_dff_B_RJTu95gr9_2;
	wire w_dff_B_vuVW65hV3_2;
	wire w_dff_B_GpdtCDhE0_2;
	wire w_dff_B_EtbdMEIt7_2;
	wire w_dff_B_gL9dlKkl5_2;
	wire w_dff_B_wbzRpzcA5_2;
	wire w_dff_B_iVbP97Cc2_2;
	wire w_dff_B_NNZxI4Y85_2;
	wire w_dff_B_zO54pNgP7_2;
	wire w_dff_B_zxiSrnG13_2;
	wire w_dff_B_Vlr8Yz1X6_2;
	wire w_dff_B_wKqaqs3V7_2;
	wire w_dff_A_oCU1WYQG2_0;
	wire w_dff_B_sU9bcwMw6_1;
	wire w_dff_B_VJypzdYV9_2;
	wire w_dff_B_Y2k4OLYn9_2;
	wire w_dff_B_BjMOCRay1_2;
	wire w_dff_B_imY2ErmR9_2;
	wire w_dff_B_TY4unhCk6_2;
	wire w_dff_B_7gY5SbKn7_2;
	wire w_dff_B_7WMmc1Q55_2;
	wire w_dff_B_Z7pnereq8_2;
	wire w_dff_B_uky2RO3m1_2;
	wire w_dff_B_WCkNCACs6_2;
	wire w_dff_B_skYH6HWA4_2;
	wire w_dff_B_DDRNHVOi9_2;
	wire w_dff_B_IfW36s7h2_2;
	wire w_dff_B_wZmO0LWb3_2;
	wire w_dff_B_CfzwRqWY3_2;
	wire w_dff_B_tqabiXk82_2;
	wire w_dff_B_Y9CPakYO9_2;
	wire w_dff_B_v9p8bOxX9_2;
	wire w_dff_B_haKXbpP99_2;
	wire w_dff_B_udy1DNGD2_2;
	wire w_dff_B_WKiDCyR22_2;
	wire w_dff_B_WlRhaTgl7_2;
	wire w_dff_B_t5Hj2OAO4_2;
	wire w_dff_B_4NhvaBxW3_2;
	wire w_dff_B_UbmjPo4v2_2;
	wire w_dff_B_VczT7VEE2_2;
	wire w_dff_B_cB3JZs4O7_2;
	wire w_dff_B_2xd6d1XP0_2;
	wire w_dff_B_tOKVNuNH8_2;
	wire w_dff_B_LYhKJWIc2_2;
	wire w_dff_B_nBqCEzFN0_2;
	wire w_dff_B_84Bzju1Y5_2;
	wire w_dff_B_ynuEwP5C3_2;
	wire w_dff_B_k8s1KtEa8_2;
	wire w_dff_B_ayWRMvj83_2;
	wire w_dff_B_sLv6jA1Q2_2;
	wire w_dff_B_p0TIb4wo2_2;
	wire w_dff_B_PKqJBaaX4_2;
	wire w_dff_B_PuUXjBx90_2;
	wire w_dff_B_ihQYhirz0_2;
	wire w_dff_B_AQetBEn90_2;
	wire w_dff_A_cONBtyJ46_1;
	wire w_dff_B_AvjPNMHL6_1;
	wire w_dff_B_mqiQvk0p7_1;
	wire w_dff_B_acdaogRU1_1;
	wire w_dff_B_qgxLf77o2_1;
	wire w_dff_B_fFsmRr6I2_1;
	wire w_dff_B_jcUMisnA9_1;
	wire w_dff_B_2eOApgTo6_1;
	wire w_dff_B_6scP1DdX7_1;
	wire w_dff_B_TSPbQ89E1_1;
	wire w_dff_B_fGWUI9Tp2_1;
	wire w_dff_B_M3u0kNba0_1;
	wire w_dff_B_VIQCteMv2_1;
	wire w_dff_B_SRQYIHw39_1;
	wire w_dff_B_MmkCkwgi4_1;
	wire w_dff_B_lxBhCIgM5_1;
	wire w_dff_B_6ED25RvQ3_1;
	wire w_dff_B_WBldEzQT6_1;
	wire w_dff_B_CPlagn032_1;
	wire w_dff_B_2DjvS6QV6_1;
	wire w_dff_B_jmOwVMch1_1;
	wire w_dff_B_MLvqnb6r0_1;
	wire w_dff_B_xZtk7he16_1;
	wire w_dff_B_D1HSzlMy5_1;
	wire w_dff_B_USsH6uLG6_1;
	wire w_dff_B_63BIwxNr4_1;
	wire w_dff_B_MkaGDmVJ4_1;
	wire w_dff_B_fzUX9pqF2_1;
	wire w_dff_B_ZEqeuxXy8_1;
	wire w_dff_B_YH8ylwvq8_1;
	wire w_dff_B_bOLYBQKJ0_1;
	wire w_dff_B_adV0flcJ0_1;
	wire w_dff_B_DPKHiAnn9_1;
	wire w_dff_B_9NcFDRM84_1;
	wire w_dff_B_n67DSODH3_1;
	wire w_dff_B_7l2d7zuR9_1;
	wire w_dff_B_6DCynWGq4_1;
	wire w_dff_B_7RVIsGbA0_1;
	wire w_dff_B_ovdRJMmp2_1;
	wire w_dff_A_UVdQvCkA8_0;
	wire w_dff_A_04aJCo1j7_0;
	wire w_dff_A_UxLiuMz43_0;
	wire w_dff_A_KhvWNSVw3_0;
	wire w_dff_A_ms6nHWDr4_0;
	wire w_dff_A_CIWGLgWw2_0;
	wire w_dff_A_xkzRNhBk4_0;
	wire w_dff_A_xTzD6xi55_0;
	wire w_dff_A_lszBqshw8_0;
	wire w_dff_A_BQj4aOpR2_0;
	wire w_dff_A_0xU5GpCO3_0;
	wire w_dff_A_Qv7ZXBIv3_0;
	wire w_dff_A_k7Df8nbQ4_0;
	wire w_dff_A_QQiiX0Vu0_0;
	wire w_dff_A_9piMC1ul0_0;
	wire w_dff_A_6AQH89uj8_0;
	wire w_dff_A_4xNyVkIb0_0;
	wire w_dff_A_6WqT3W6u4_0;
	wire w_dff_A_kiUOKrWm1_0;
	wire w_dff_A_AeuFT1PZ5_0;
	wire w_dff_A_oa8WIHar6_0;
	wire w_dff_A_Fd0sMzLa5_0;
	wire w_dff_A_vOuxIzFn3_0;
	wire w_dff_A_VdoUm5ic5_0;
	wire w_dff_A_WTkvgKrv1_0;
	wire w_dff_A_bp7H5e9c0_0;
	wire w_dff_A_u6MW3VeA7_0;
	wire w_dff_A_wMp9Fyq01_0;
	wire w_dff_A_qyK09UQA0_0;
	wire w_dff_A_Vvrmtr2d3_0;
	wire w_dff_A_phSzcfPN8_0;
	wire w_dff_A_tDjoEEd31_0;
	wire w_dff_A_W39d1HSr2_0;
	wire w_dff_A_Amm4FCpX8_0;
	wire w_dff_A_vqcRHNxM6_0;
	wire w_dff_A_r8hunF2l9_0;
	wire w_dff_A_Mz91aW7g2_0;
	wire w_dff_A_gv2XXJR31_0;
	wire w_dff_A_pNJ353jV9_0;
	wire w_dff_B_EyD3ZNz90_1;
	wire w_dff_A_HuXg3usU8_0;
	wire w_dff_A_VhUgFByC0_0;
	wire w_dff_A_T8OBfhSl4_0;
	wire w_dff_A_ZTw5wOAj9_0;
	wire w_dff_A_Iq7nWvCZ3_0;
	wire w_dff_A_yAVt7SLb7_0;
	wire w_dff_A_3T4qwT0d2_0;
	wire w_dff_A_tloxYKW44_0;
	wire w_dff_A_ICBfhIee0_0;
	wire w_dff_A_6pWsmhI01_0;
	wire w_dff_A_OMfI1VVd3_0;
	wire w_dff_A_31gBrAmU9_0;
	wire w_dff_A_KYey5Sve1_0;
	wire w_dff_A_HVEucIQN2_0;
	wire w_dff_A_rkunZU9h1_0;
	wire w_dff_A_j1oYindC5_0;
	wire w_dff_A_VYrKM87F3_0;
	wire w_dff_A_EKz6TQDI9_0;
	wire w_dff_A_f2mVVxbV6_0;
	wire w_dff_A_jLXU7hEw3_0;
	wire w_dff_A_Dh7TuOOs1_0;
	wire w_dff_A_gee1VQJY0_0;
	wire w_dff_A_UiBaxkEB2_0;
	wire w_dff_A_gF0DgSDn7_0;
	wire w_dff_A_5nJP6kj45_0;
	wire w_dff_A_5YlSKAyw2_0;
	wire w_dff_A_9UrDpWcG8_0;
	wire w_dff_A_0xb8Nnld4_0;
	wire w_dff_A_b0OUSrwL9_0;
	wire w_dff_A_tKVgjKau1_0;
	wire w_dff_A_NhYBq0aE6_0;
	wire w_dff_A_294attYK5_0;
	wire w_dff_A_tGA5ayuD0_0;
	wire w_dff_A_1U8j3zsV2_0;
	wire w_dff_A_KkeADDaJ8_0;
	wire w_dff_A_TUptm82n2_0;
	wire w_dff_B_BZtiQIGW5_1;
	wire w_dff_A_YmDAWMXy9_0;
	wire w_dff_A_3sjevCOi3_0;
	wire w_dff_A_LuA94Ww84_0;
	wire w_dff_A_ZEFFbOkh0_0;
	wire w_dff_A_36Ksepbw6_0;
	wire w_dff_A_BqwJaW1i7_0;
	wire w_dff_A_WV7QDBiF0_0;
	wire w_dff_A_Q9VywNaz5_0;
	wire w_dff_A_dRGyk5DL1_0;
	wire w_dff_A_a6JJmDOB4_0;
	wire w_dff_A_8sF6Pv531_0;
	wire w_dff_A_PVGlaclK5_0;
	wire w_dff_A_AVHr9Sag9_0;
	wire w_dff_A_9yEu5N526_0;
	wire w_dff_A_FFbwqjPf7_0;
	wire w_dff_A_BN9ZPw1b9_0;
	wire w_dff_A_d622n9di5_0;
	wire w_dff_A_xxYF6zzz1_0;
	wire w_dff_A_LwGpTb137_0;
	wire w_dff_A_B31UjaJ41_0;
	wire w_dff_A_umLnOgFL4_0;
	wire w_dff_A_sjVppoKo5_0;
	wire w_dff_A_oGxl3qyH6_0;
	wire w_dff_A_uK2dd1MW6_0;
	wire w_dff_A_og1RfghJ3_0;
	wire w_dff_A_NBSdpVgE9_0;
	wire w_dff_A_X2au5xLe7_0;
	wire w_dff_A_faA1aRbu0_0;
	wire w_dff_A_uorRZza72_0;
	wire w_dff_A_sOpgKyRl1_0;
	wire w_dff_A_HnJjiojV1_0;
	wire w_dff_A_Jpe6BBw50_0;
	wire w_dff_A_XG0hYoUi2_0;
	wire w_dff_B_wMbzty9e4_1;
	wire w_dff_A_KaHITHHw3_0;
	wire w_dff_A_YHcdlSYS8_0;
	wire w_dff_A_71bnE8T27_0;
	wire w_dff_A_IcYZhxDj6_0;
	wire w_dff_A_MeUppa0m2_0;
	wire w_dff_A_vDoUtolz6_0;
	wire w_dff_A_FtzTPT0R4_0;
	wire w_dff_A_qkDOJSN16_0;
	wire w_dff_A_Exg6Qtis6_0;
	wire w_dff_A_w2w9PQBI8_0;
	wire w_dff_A_J2LgcBq67_0;
	wire w_dff_A_DeMBVa2p6_0;
	wire w_dff_A_dzqe0GZw0_0;
	wire w_dff_A_IcvYiBy34_0;
	wire w_dff_A_t5ToewZA2_0;
	wire w_dff_A_5CZrI5LA4_0;
	wire w_dff_A_AxmcDDgY1_0;
	wire w_dff_A_K7y1rP592_0;
	wire w_dff_A_MVOJowLq9_0;
	wire w_dff_A_IAsHkHwr8_0;
	wire w_dff_A_6Z8LPAIr1_0;
	wire w_dff_A_rT5Ohd2b5_0;
	wire w_dff_A_zfIy0Op68_0;
	wire w_dff_A_z2sX11c36_0;
	wire w_dff_A_XVEZyGxX8_0;
	wire w_dff_A_6oUrGpVr9_0;
	wire w_dff_A_vozhl1db5_0;
	wire w_dff_A_AX55zDq92_0;
	wire w_dff_A_VqxSOFmS0_0;
	wire w_dff_A_2N5I4kY78_0;
	wire w_dff_B_FEoRVAiC6_1;
	wire w_dff_A_rSSfFkGL7_0;
	wire w_dff_A_2P6IX7Vy4_0;
	wire w_dff_A_jZ0Pp9hB4_0;
	wire w_dff_A_FuL9DUHR5_0;
	wire w_dff_A_nFAIsQCq7_0;
	wire w_dff_A_gcJcQK3r4_0;
	wire w_dff_A_eUkOJ6RB7_0;
	wire w_dff_A_Bzw9U4m02_0;
	wire w_dff_A_mf73h0d85_0;
	wire w_dff_A_OhHNfjlm2_0;
	wire w_dff_A_B2Fb4YMo2_0;
	wire w_dff_A_u6twTcmm9_0;
	wire w_dff_A_wAzQ8J249_0;
	wire w_dff_A_apdojfAh8_0;
	wire w_dff_A_VGhAByjY6_0;
	wire w_dff_A_VM7tfSf83_0;
	wire w_dff_A_J7xDq3NS9_0;
	wire w_dff_A_GMkWIvKo6_0;
	wire w_dff_A_plhgGVHr5_0;
	wire w_dff_A_PXn4uhnT1_0;
	wire w_dff_A_tBZUMiHN1_0;
	wire w_dff_A_16NOPfRQ9_0;
	wire w_dff_A_zmfxMyyQ8_0;
	wire w_dff_A_CNh7Nu3u2_0;
	wire w_dff_A_gtpigkUz9_0;
	wire w_dff_A_ymql107S1_0;
	wire w_dff_A_14eYYD6s0_0;
	wire w_dff_B_kPMvTxiM2_1;
	wire w_dff_A_YeJVYQXg0_0;
	wire w_dff_A_R38Uz8Qr5_0;
	wire w_dff_A_YeDyhrtn7_0;
	wire w_dff_A_JRTqZJJi4_0;
	wire w_dff_A_GppyQCC35_0;
	wire w_dff_A_ZVfjUG6W6_0;
	wire w_dff_A_HUEjaspn9_0;
	wire w_dff_A_Eycn70NM7_0;
	wire w_dff_A_1dG69cYp3_0;
	wire w_dff_A_LEBvhOVo8_0;
	wire w_dff_A_um5d6ucm7_0;
	wire w_dff_A_yDEYgugP7_0;
	wire w_dff_A_fFN5noq34_0;
	wire w_dff_A_th0X1hPA4_0;
	wire w_dff_A_xENboy8f2_0;
	wire w_dff_A_uP4UVEoX6_0;
	wire w_dff_A_SdN53j033_0;
	wire w_dff_A_uud2UxEa9_0;
	wire w_dff_A_6rdpdBqO0_0;
	wire w_dff_A_AFdo8ZFi4_0;
	wire w_dff_A_arRcaiPL9_0;
	wire w_dff_A_wNODA5kc9_0;
	wire w_dff_A_4O2bYNf23_0;
	wire w_dff_A_f6dTGFVx1_0;
	wire w_dff_B_fe1ABSNx2_1;
	wire w_dff_A_v4h6FCT37_0;
	wire w_dff_A_xurBvHRF2_0;
	wire w_dff_A_thaJ0oX79_0;
	wire w_dff_A_3J2MmRBC0_0;
	wire w_dff_A_EoRG3Vju7_0;
	wire w_dff_A_fPKf6J8R7_0;
	wire w_dff_A_HfWU2cp27_0;
	wire w_dff_A_S3sF77xW4_0;
	wire w_dff_A_qnzCvVW00_0;
	wire w_dff_A_Oo8rQiay1_0;
	wire w_dff_A_aZ8uug2N0_0;
	wire w_dff_A_O9TNbANi8_0;
	wire w_dff_A_UsrYieBD6_0;
	wire w_dff_A_LxWqcRCL8_0;
	wire w_dff_A_LhjZQx3V7_0;
	wire w_dff_A_xp19xgGk1_0;
	wire w_dff_A_6wr8L5QS8_0;
	wire w_dff_A_Il3ZipLs2_0;
	wire w_dff_A_W4SPQo6p9_0;
	wire w_dff_A_fWFkXRlH4_0;
	wire w_dff_A_QRKEAwBf9_0;
	wire w_dff_B_O8JHUWz01_1;
	wire w_dff_A_9POCDiGY1_0;
	wire w_dff_A_ZCHKqSSI1_0;
	wire w_dff_A_0S0TpdwX1_0;
	wire w_dff_A_Mdz7uxmj4_0;
	wire w_dff_A_I4W6y1b86_0;
	wire w_dff_A_w9YcuNlA4_0;
	wire w_dff_A_4Yyi2UMC7_0;
	wire w_dff_A_m6OJCe4J6_0;
	wire w_dff_A_T10kneES8_0;
	wire w_dff_A_LY7tWZne4_0;
	wire w_dff_A_ixXQUpog3_0;
	wire w_dff_A_JesL3Qq71_0;
	wire w_dff_A_RwR5CIS09_0;
	wire w_dff_A_awMZdQbR4_0;
	wire w_dff_A_wdugtVvB2_0;
	wire w_dff_A_4J1mDx4A8_0;
	wire w_dff_A_9rl5Eyhd7_0;
	wire w_dff_A_MysAQcee9_0;
	wire w_dff_B_cbtQ91dg3_1;
	wire w_dff_A_4IDSjOmg1_0;
	wire w_dff_A_yeXiaizK6_0;
	wire w_dff_A_BRa5oHz15_0;
	wire w_dff_A_8A3KkQU06_0;
	wire w_dff_A_dKFWCrB36_0;
	wire w_dff_A_GbwxdbAl8_0;
	wire w_dff_A_wxEnhyk05_0;
	wire w_dff_A_SxUNq4le0_0;
	wire w_dff_A_vx89NLt18_0;
	wire w_dff_A_TS2dk8aB6_0;
	wire w_dff_A_Ft1061mu7_0;
	wire w_dff_A_CO63azFW2_0;
	wire w_dff_A_sbQXxpaQ1_0;
	wire w_dff_A_4hwEkcxO6_0;
	wire w_dff_A_UvMWN99Q9_0;
	wire w_dff_B_eeFZZLUH4_1;
	wire w_dff_A_dkxWOv9F3_0;
	wire w_dff_A_2T6ae3xM2_0;
	wire w_dff_A_ma8HyiPD1_0;
	wire w_dff_A_U2wuna6b7_0;
	wire w_dff_A_UpQ6p02F9_0;
	wire w_dff_A_deECsCTN8_0;
	wire w_dff_A_SK85NqZm4_0;
	wire w_dff_A_yIvN9eRV9_0;
	wire w_dff_A_ibvQb0Gk5_0;
	wire w_dff_A_LjPZjcXj8_0;
	wire w_dff_A_HWEN1MZi5_0;
	wire w_dff_A_AQPO0Rr33_0;
	wire w_dff_B_1ANJNn590_1;
	wire w_dff_A_zrNSo0n93_0;
	wire w_dff_A_lOpvbmHH4_0;
	wire w_dff_A_AntLwJ2t4_0;
	wire w_dff_A_gk6giD027_0;
	wire w_dff_A_sCloH9aA0_0;
	wire w_dff_A_IBKEFPBT2_0;
	wire w_dff_A_7Xa03SXm3_0;
	wire w_dff_A_NiDcVqga0_0;
	wire w_dff_A_SwFztyXO9_0;
	wire w_dff_A_tW1bCqem0_0;
	wire w_dff_A_MmWWRJ4h6_0;
	wire w_dff_A_latRsa6l4_1;
	wire w_dff_A_tARccCuP3_0;
	wire w_dff_A_2FdPF67W0_0;
	wire w_dff_A_4pnYCnEO6_0;
	wire w_dff_A_kb4H3JFE0_0;
	wire w_dff_A_GfrnQwgt6_0;
	wire w_dff_A_dAinsZSM4_0;
	wire w_dff_A_nDVYqqP91_0;
	wire w_dff_B_OcM2U1nk7_1;
	wire w_dff_A_balw0lKA6_1;
	wire w_dff_A_z69XGoAz2_2;
	wire w_dff_A_jO2YVfKU2_2;
	wire w_dff_A_NPQRlaQD6_0;
	wire w_dff_B_QGHX3ctl8_2;
	wire w_dff_B_MHoeFrk23_2;
	wire w_dff_B_gws117dq8_2;
	wire w_dff_B_tifPlCMi5_2;
	wire w_dff_B_Rj64qouw7_2;
	wire w_dff_B_kQlaz3Tw8_2;
	wire w_dff_B_rRtv8xqQ1_2;
	wire w_dff_B_ey2UuyBs2_2;
	wire w_dff_B_F0p8rIpF7_2;
	wire w_dff_B_Br6ydx2a0_2;
	wire w_dff_B_2zzmWZYw0_2;
	wire w_dff_B_vp6DkEgp1_2;
	wire w_dff_B_MDnTEYkg5_2;
	wire w_dff_B_F3di0N1X6_2;
	wire w_dff_B_GAOlDm706_2;
	wire w_dff_B_7jCxRxhH3_2;
	wire w_dff_B_ifmk5Njb2_2;
	wire w_dff_B_aIOg3fAo8_2;
	wire w_dff_B_0ATg7qQP5_2;
	wire w_dff_B_7H3zKe8G2_2;
	wire w_dff_B_k910qDAn8_2;
	wire w_dff_B_Xxr9HxW06_2;
	wire w_dff_B_wOXhzEnW7_2;
	wire w_dff_B_d1jkG5A91_2;
	wire w_dff_B_Zvy5EmfT8_2;
	wire w_dff_B_M7Dc5XBP8_2;
	wire w_dff_B_18qI0mSA0_2;
	wire w_dff_B_uUHLfI278_2;
	wire w_dff_B_idxkNm928_2;
	wire w_dff_B_icSfbRwi4_2;
	wire w_dff_B_LcGvbYJG9_2;
	wire w_dff_B_RupLQkck6_2;
	wire w_dff_B_SqA6HFO79_2;
	wire w_dff_B_8ZUQ4tkS4_2;
	wire w_dff_B_ag5IAlUv0_2;
	wire w_dff_B_PNcUOeWy6_2;
	wire w_dff_B_FY9qpg459_2;
	wire w_dff_B_OeklvmLV9_2;
	wire w_dff_B_XWAljari1_2;
	wire w_dff_B_iJHGWhC59_2;
	wire w_dff_B_Qrjc45HK0_2;
	wire w_dff_B_RrNwMvPl4_2;
	wire w_dff_B_ObwdBbpI9_2;
	wire w_dff_B_V7ssezCX9_2;
	wire w_dff_B_RMjRo5a85_2;
	wire w_dff_A_Gr7HxICE1_0;
	wire w_dff_B_C5C6vHsw0_1;
	wire w_dff_B_iaZRAhFW6_2;
	wire w_dff_B_2TDY65Zz8_2;
	wire w_dff_B_0fhOpMHw5_2;
	wire w_dff_B_vvzU0n9K2_2;
	wire w_dff_B_10vFc8aT8_2;
	wire w_dff_B_SMvp4JlQ5_2;
	wire w_dff_B_tP7UwAxs3_2;
	wire w_dff_B_JfNg4S6k6_2;
	wire w_dff_B_bYrUj9De7_2;
	wire w_dff_B_Cgosjsxv6_2;
	wire w_dff_B_Aml9V9434_2;
	wire w_dff_B_a7R85p2m3_2;
	wire w_dff_B_5xuTbzze6_2;
	wire w_dff_B_V0r0Cty86_2;
	wire w_dff_B_wbkapKat3_2;
	wire w_dff_B_X0QoIk4I0_2;
	wire w_dff_B_ika6nGXW6_2;
	wire w_dff_B_wyaMoXPG7_2;
	wire w_dff_B_JNFVLx476_2;
	wire w_dff_B_x6WgiwO93_2;
	wire w_dff_B_JMVRf94X0_2;
	wire w_dff_B_BoPQ9V3g4_2;
	wire w_dff_B_ZYOlnaYm7_2;
	wire w_dff_B_4jhnZ5ka0_2;
	wire w_dff_B_eIRitcNo3_2;
	wire w_dff_B_TvqE9uf95_2;
	wire w_dff_B_3bKDlMsj1_2;
	wire w_dff_B_DcS1Cs1W5_2;
	wire w_dff_B_fonBbvhv6_2;
	wire w_dff_B_y1KNow2p2_2;
	wire w_dff_B_BIs2VB3x1_2;
	wire w_dff_B_Czt5w7if6_2;
	wire w_dff_B_9GKbfECR6_2;
	wire w_dff_B_0VfGIVGN6_2;
	wire w_dff_B_0bHdgDPC4_2;
	wire w_dff_B_spyQcbM83_2;
	wire w_dff_B_QJYOa0LS2_2;
	wire w_dff_B_CF9HbN4S9_2;
	wire w_dff_B_cPZGtjOu4_2;
	wire w_dff_B_IJd8LxC51_2;
	wire w_dff_B_YoBgo9Qz8_2;
	wire w_dff_A_Voa2nWZi3_1;
	wire w_dff_A_wffRyLGQ2_0;
	wire w_dff_A_Jiev30sR6_0;
	wire w_dff_A_yRzzr99x9_0;
	wire w_dff_A_okwQI6dM4_0;
	wire w_dff_A_WlfA4e3J1_0;
	wire w_dff_A_9izv6p7Q0_0;
	wire w_dff_A_oG2l49pI2_0;
	wire w_dff_A_JrvRMgIl1_0;
	wire w_dff_A_o6Cj6fUe2_0;
	wire w_dff_A_AZb03TZg5_0;
	wire w_dff_A_AYp5yxnn5_0;
	wire w_dff_A_M83VFdcT0_0;
	wire w_dff_A_vgfgNsFQ8_0;
	wire w_dff_A_AbLuLFGa1_0;
	wire w_dff_A_0enXMpnx4_0;
	wire w_dff_A_2SNGlnfv3_0;
	wire w_dff_A_DuIUZFrL8_0;
	wire w_dff_A_8fEtIe8F0_0;
	wire w_dff_A_NIK03Wgq9_0;
	wire w_dff_A_QjXnEzaT1_0;
	wire w_dff_A_bzEBMzYu8_0;
	wire w_dff_A_oa3qovs33_0;
	wire w_dff_A_j22LvmOX9_0;
	wire w_dff_A_WO8fjwTM6_0;
	wire w_dff_A_k4v5EosN3_0;
	wire w_dff_A_bvLb5Hwb9_0;
	wire w_dff_A_gl2Xkir28_0;
	wire w_dff_A_cKB4c44g8_0;
	wire w_dff_A_fIXzMqHS5_0;
	wire w_dff_A_DtHx8EY68_0;
	wire w_dff_A_8PxlBvTy6_0;
	wire w_dff_A_yC00dDdR2_0;
	wire w_dff_A_DkrMaw6R4_0;
	wire w_dff_A_PddTMFSd3_0;
	wire w_dff_A_X1EWdI6e8_0;
	wire w_dff_A_gEHaypot5_0;
	wire w_dff_A_aGBweFga6_0;
	wire w_dff_A_rddEyTe76_0;
	wire w_dff_A_wALpsxUl8_1;
	wire w_dff_A_9OrlJGK70_2;
	wire w_dff_B_fW2vjjGI2_1;
	wire w_dff_B_IJ5OlnYO2_2;
	wire w_dff_B_8IgOr1vF2_2;
	wire w_dff_B_rl6nwMBb7_2;
	wire w_dff_B_TStHV4gC1_2;
	wire w_dff_B_VS3KmYDs1_2;
	wire w_dff_B_RDOWJLpY9_2;
	wire w_dff_B_F4WPU77a4_2;
	wire w_dff_B_MsPTZtWX0_2;
	wire w_dff_B_N7hLyVMd8_2;
	wire w_dff_B_UaRHLEQh0_2;
	wire w_dff_B_KKTM7mhX0_2;
	wire w_dff_B_eFNfMcul8_2;
	wire w_dff_B_CGWKM9Es8_2;
	wire w_dff_B_SKRDRi1s4_2;
	wire w_dff_B_gSelskiQ9_2;
	wire w_dff_B_O39CEEfe2_2;
	wire w_dff_B_Hn0InsQg1_2;
	wire w_dff_B_CE985Xd50_2;
	wire w_dff_B_GtU9kTDA0_2;
	wire w_dff_B_OB8Bx5xK2_2;
	wire w_dff_B_GLYUIhhM4_2;
	wire w_dff_B_kYmFj8NL4_2;
	wire w_dff_B_LatTYkkC1_2;
	wire w_dff_B_dQMelPoN9_2;
	wire w_dff_B_RGqQmZMC8_2;
	wire w_dff_B_oOjENsPs8_2;
	wire w_dff_B_rkcCQZ1A9_2;
	wire w_dff_B_QOlkaEfQ8_2;
	wire w_dff_B_1IeHQctC1_2;
	wire w_dff_B_HeUSRud13_2;
	wire w_dff_B_SaltxAMU0_2;
	wire w_dff_B_9V9GPrAc5_2;
	wire w_dff_B_YFh1Hbc80_2;
	wire w_dff_B_XHgoh4ZN7_2;
	wire w_dff_B_xlzt7Jp13_2;
	wire w_dff_B_oSL6BcdO5_1;
	wire w_dff_B_iMdscc0W2_2;
	wire w_dff_B_jFQW4TTe5_2;
	wire w_dff_B_tGPVsApc9_2;
	wire w_dff_B_pGsXkn8C9_2;
	wire w_dff_B_057dNnmj0_2;
	wire w_dff_B_OY10Ofyj4_2;
	wire w_dff_B_rbpXlvB25_2;
	wire w_dff_B_Bqq1RtNr1_2;
	wire w_dff_B_liNTPTn07_2;
	wire w_dff_B_ZgOedF5v2_2;
	wire w_dff_B_UTHrbvr56_2;
	wire w_dff_B_Z1kbUkjJ4_2;
	wire w_dff_B_r2aTpHtA9_2;
	wire w_dff_B_TQBDAibS2_2;
	wire w_dff_B_UFo8eQQv2_2;
	wire w_dff_B_Zmc2OscO3_2;
	wire w_dff_B_QroViJCe0_2;
	wire w_dff_B_5vHej5g29_2;
	wire w_dff_B_balQTqqz3_2;
	wire w_dff_B_3sTWP1yL3_2;
	wire w_dff_B_YT72ouv26_2;
	wire w_dff_B_5ODYHuU70_2;
	wire w_dff_B_BigxqMvF8_2;
	wire w_dff_B_AVo9YrBg9_2;
	wire w_dff_B_GcNonWx66_2;
	wire w_dff_B_UKi28Gol0_2;
	wire w_dff_B_zOMFcPxr4_2;
	wire w_dff_B_bZJxbUq97_2;
	wire w_dff_B_CVPIZxQW3_2;
	wire w_dff_B_mWtJKION0_2;
	wire w_dff_B_53epCT4a7_2;
	wire w_dff_B_ZBEN2qtH8_2;
	wire w_dff_B_mEGkhFkZ1_1;
	wire w_dff_B_QNY9H9gw2_2;
	wire w_dff_B_qMXoEl3D7_2;
	wire w_dff_B_FInI1Q5Q0_2;
	wire w_dff_B_Hj0o3xIa6_2;
	wire w_dff_B_PpNK2lKF5_2;
	wire w_dff_B_6ruxRVpm7_2;
	wire w_dff_B_l1sk7anW1_2;
	wire w_dff_B_0LpA89Jc7_2;
	wire w_dff_B_1XyAd6jb9_2;
	wire w_dff_B_roRoidhf6_2;
	wire w_dff_B_Vh5jt5Ez2_2;
	wire w_dff_B_hZMrdm1s0_2;
	wire w_dff_B_bt2OBplg4_2;
	wire w_dff_B_2CCavDMt0_2;
	wire w_dff_B_pAgxNNHr2_2;
	wire w_dff_B_uTiVbRAA8_2;
	wire w_dff_B_Zbqh0ZSs0_2;
	wire w_dff_B_w5XslQ6o1_2;
	wire w_dff_B_5DNGVSKm0_2;
	wire w_dff_B_EewqZM6m7_2;
	wire w_dff_B_KnMiODfg2_2;
	wire w_dff_B_ptY0swbn7_2;
	wire w_dff_B_kjBbuBWi9_2;
	wire w_dff_B_D96xFsyD7_2;
	wire w_dff_B_LoGBgwd11_2;
	wire w_dff_B_XYasrhLl9_2;
	wire w_dff_B_xk4ibRrF9_2;
	wire w_dff_B_S0rXoPdI4_2;
	wire w_dff_B_9FCmbrcm4_2;
	wire w_dff_B_qm7W71SE7_1;
	wire w_dff_B_UJCveD5s6_2;
	wire w_dff_B_XhEtsp7o1_2;
	wire w_dff_B_7TDTOO5L2_2;
	wire w_dff_B_j6oRqiWS4_2;
	wire w_dff_B_2GhB4nT59_2;
	wire w_dff_B_ccEB6Pcf4_2;
	wire w_dff_B_oBomMU8s7_2;
	wire w_dff_B_KNKsVjQm0_2;
	wire w_dff_B_nt40BZEQ4_2;
	wire w_dff_B_Rwy0X4qp1_2;
	wire w_dff_B_k9NhsHdL9_2;
	wire w_dff_B_OgDnLGtX7_2;
	wire w_dff_B_pPJF5NhR9_2;
	wire w_dff_B_kc4KIVQx5_2;
	wire w_dff_B_IC22vasF6_2;
	wire w_dff_B_f1wTeq276_2;
	wire w_dff_B_vBVb1UCN5_2;
	wire w_dff_B_BhBeVO2I9_2;
	wire w_dff_B_FSxNYMdQ9_2;
	wire w_dff_B_N8DuCpGu2_2;
	wire w_dff_B_kiSpnneP1_2;
	wire w_dff_B_YPdz383g3_2;
	wire w_dff_B_GgPbChkp9_2;
	wire w_dff_B_I8e2cYpL6_2;
	wire w_dff_B_CCND9ubK0_2;
	wire w_dff_B_WcIQi2vz7_2;
	wire w_dff_B_Voqlg2Yh1_1;
	wire w_dff_B_sdAh0Vr59_2;
	wire w_dff_B_HWYeEN6q5_2;
	wire w_dff_B_EbCUtrqW3_2;
	wire w_dff_B_pybQll3U4_2;
	wire w_dff_B_F7jBQweO7_2;
	wire w_dff_B_2vXrbfAh1_2;
	wire w_dff_B_0YqPQxRO0_2;
	wire w_dff_B_o4abx7OD4_2;
	wire w_dff_B_BbHWM7GS3_2;
	wire w_dff_B_O3NBLQHP3_2;
	wire w_dff_B_HfLyjiRQ8_2;
	wire w_dff_B_GlUM8oqM5_2;
	wire w_dff_B_6HUbN8uF2_2;
	wire w_dff_B_nkT76NXQ8_2;
	wire w_dff_B_fX5wZIZn9_2;
	wire w_dff_B_rvPz3zkP7_2;
	wire w_dff_B_ljo04jbn2_2;
	wire w_dff_B_V1ZSVRvV4_2;
	wire w_dff_B_YvxezPYK2_2;
	wire w_dff_B_M3KLAOSb8_2;
	wire w_dff_B_QdKVDZSg5_2;
	wire w_dff_B_m3egyPwj4_2;
	wire w_dff_B_A822Pj3E2_2;
	wire w_dff_B_NdpLZSRB4_1;
	wire w_dff_B_XUqUdk527_2;
	wire w_dff_B_mfiIfL1c9_2;
	wire w_dff_B_CaB7WW3i5_2;
	wire w_dff_B_a7SQIuAl9_2;
	wire w_dff_B_i1YtFsae0_2;
	wire w_dff_B_LgQKcvdf3_2;
	wire w_dff_B_iHry2Aq55_2;
	wire w_dff_B_mMgSrYur5_2;
	wire w_dff_B_eNYHndts9_2;
	wire w_dff_B_L2PolUdN0_2;
	wire w_dff_B_ajjNMWC26_2;
	wire w_dff_B_zfI7wkQw6_2;
	wire w_dff_B_qCWSYLrs6_2;
	wire w_dff_B_1wvC4odU9_2;
	wire w_dff_B_PUpj6HfG9_2;
	wire w_dff_B_LMGXKl6t7_2;
	wire w_dff_B_5BpYIurk2_2;
	wire w_dff_B_ag9VBo1Y6_2;
	wire w_dff_B_o72n8RB88_2;
	wire w_dff_B_ce9XI3zW7_2;
	wire w_dff_B_jDbqou9V2_1;
	wire w_dff_B_7GHg35vR0_2;
	wire w_dff_B_oCDg3lK08_2;
	wire w_dff_B_TcUJFPef2_2;
	wire w_dff_B_HzEkmRhg0_2;
	wire w_dff_B_LWuWehQz4_2;
	wire w_dff_B_5P0B3daq3_2;
	wire w_dff_B_QLyzIFN62_2;
	wire w_dff_B_QWjgs8c67_2;
	wire w_dff_B_snrHGHww9_2;
	wire w_dff_B_NXZQbBGI2_2;
	wire w_dff_B_uvL3rfcW6_2;
	wire w_dff_B_m7NKtxLp4_2;
	wire w_dff_B_EYmoJy0P8_2;
	wire w_dff_B_oXEPrpvp0_2;
	wire w_dff_B_B8d0Foqb2_2;
	wire w_dff_B_9vo0u5m23_2;
	wire w_dff_B_3RE2EL7P0_2;
	wire w_dff_B_al8aNhS70_1;
	wire w_dff_B_k6V0TNG19_2;
	wire w_dff_B_MXawkFPT4_2;
	wire w_dff_B_1othvyRy4_2;
	wire w_dff_B_r2xHZHD81_2;
	wire w_dff_B_mO3HnqJG0_2;
	wire w_dff_B_D7ZVLqB92_2;
	wire w_dff_B_N433o7ZI4_2;
	wire w_dff_B_BdcSgprP4_2;
	wire w_dff_B_qRGWIEP82_2;
	wire w_dff_B_22AIujaK0_2;
	wire w_dff_B_03nXaE3f7_2;
	wire w_dff_B_UjOpp8Dk8_2;
	wire w_dff_B_psODmytO6_2;
	wire w_dff_B_DveKxQYH6_2;
	wire w_dff_B_2fcWdJM90_1;
	wire w_dff_B_v1Z9jLdn7_2;
	wire w_dff_B_OGDdeCCB7_2;
	wire w_dff_B_G8xzG6C29_2;
	wire w_dff_B_UERly8ar0_2;
	wire w_dff_B_2xCgGoC53_2;
	wire w_dff_B_Yrxj0Kgk9_2;
	wire w_dff_B_4WYVfu2E8_2;
	wire w_dff_B_vMZ5OOKg0_2;
	wire w_dff_B_d8kcAuRM0_2;
	wire w_dff_B_tViMIGoP6_2;
	wire w_dff_B_LYxRxdqy1_2;
	wire w_dff_B_5TW31LH74_1;
	wire w_dff_B_pklqfeAD2_2;
	wire w_dff_B_VIApfomQ3_2;
	wire w_dff_B_znQYor7B9_2;
	wire w_dff_B_kDZqI6jJ4_2;
	wire w_dff_B_q4MDs3Rk9_2;
	wire w_dff_B_dCnCZZZE5_2;
	wire w_dff_B_p6mphz8N5_2;
	wire w_dff_B_JHKovzKr2_2;
	wire w_dff_B_Lo1si02i0_1;
	wire w_dff_B_xBFu5Phx7_1;
	wire w_dff_B_98WjUXC83_2;
	wire w_dff_B_cZeyvtrC4_2;
	wire w_dff_B_fODRA8fO1_2;
	wire w_dff_B_s8Xsddgu1_2;
	wire w_dff_A_R32qMOHF2_1;
	wire w_dff_A_D2IVofeZ1_0;
	wire w_dff_A_9S0is7Qi5_0;
	wire w_dff_A_8BlzFoWF9_1;
	wire w_dff_A_NwSCs7bj4_2;
	wire w_dff_A_ZXYPmR2t3_2;
	wire w_dff_B_yOr46Oam9_0;
	wire w_dff_A_U692QmXf8_1;
	wire w_dff_A_IPnXeFHN0_1;
	wire w_dff_B_i5Q5GgX24_1;
	wire w_dff_B_JNPv3mIo9_1;
	wire w_dff_B_jAaslnVt5_2;
	wire w_dff_B_WDRKdxAH1_2;
	wire w_dff_B_f9uoqLHw5_2;
	wire w_dff_B_AMSHqjDG7_2;
	wire w_dff_B_o9VwloPg3_2;
	wire w_dff_B_ay0dwz2M9_2;
	wire w_dff_B_rkuvduRC8_2;
	wire w_dff_B_SxoeFFU92_2;
	wire w_dff_B_nrRDnhYj9_2;
	wire w_dff_B_P9wYd6x00_2;
	wire w_dff_B_u1Gkuo0E9_2;
	wire w_dff_B_TiZHioho0_2;
	wire w_dff_B_xicjWSWt0_2;
	wire w_dff_B_Z9PyoSK47_2;
	wire w_dff_B_2ifOi42V8_2;
	wire w_dff_B_XhAMf2eX6_2;
	wire w_dff_B_eaDWm4203_2;
	wire w_dff_B_6vWy6wCL8_2;
	wire w_dff_B_qxi5hrBP4_2;
	wire w_dff_B_VyECjBLD2_2;
	wire w_dff_B_e6XjtRon2_2;
	wire w_dff_B_CrYiwVtH3_2;
	wire w_dff_B_kCnhktvL1_2;
	wire w_dff_B_fqGu5zJg1_2;
	wire w_dff_B_scwyyet63_2;
	wire w_dff_B_0guQVbUe6_2;
	wire w_dff_B_h1VlblDI5_2;
	wire w_dff_B_EA0GKumX9_2;
	wire w_dff_B_uP1G5RxD5_2;
	wire w_dff_B_WVF5oxW86_2;
	wire w_dff_B_RU3lt3cc7_2;
	wire w_dff_B_u0KFp77y1_2;
	wire w_dff_B_S09I4NAK0_2;
	wire w_dff_B_1iXi2EKq2_2;
	wire w_dff_B_We1EybXJ2_2;
	wire w_dff_B_wAilYS1r5_2;
	wire w_dff_B_ChOaTK1q7_2;
	wire w_dff_B_seCLvjU91_2;
	wire w_dff_B_zhzxnqSk0_2;
	wire w_dff_B_Od0HTU9o4_2;
	wire w_dff_B_BITHYmtq6_2;
	wire w_dff_B_efLQbOd50_2;
	wire w_dff_B_u5obT7YS6_2;
	wire w_dff_B_K0dT0OMv0_2;
	wire w_dff_B_OtPzkkDJ3_2;
	wire w_dff_B_Ycu9g66M0_2;
	wire w_dff_B_DxnsUaBS1_2;
	wire w_dff_B_DOH2dNe61_1;
	wire w_dff_B_Dm35Epxf3_2;
	wire w_dff_B_spdaXV6m5_2;
	wire w_dff_B_6FcRjeyT7_2;
	wire w_dff_B_Eab1VxWV3_2;
	wire w_dff_B_XEXLONgk2_2;
	wire w_dff_B_y8ZMA8v00_2;
	wire w_dff_B_WHEhknZP7_2;
	wire w_dff_B_PwaeNsOc6_2;
	wire w_dff_B_PKsSXaIl1_2;
	wire w_dff_B_M81eb61a7_2;
	wire w_dff_B_scetwMPr7_2;
	wire w_dff_B_X7d9ZqKg6_2;
	wire w_dff_B_B5jRDPeS3_2;
	wire w_dff_B_dCPPhaFI7_2;
	wire w_dff_B_J3QBwTyD9_2;
	wire w_dff_B_KtSpz4A72_2;
	wire w_dff_B_X7xx28KV1_2;
	wire w_dff_B_20jGAzNF7_2;
	wire w_dff_B_dH5f8ZMy5_2;
	wire w_dff_B_92asM1Ah7_2;
	wire w_dff_B_nRLOAZKs0_2;
	wire w_dff_B_2Mjul4hS6_2;
	wire w_dff_B_OUHK7XmR8_2;
	wire w_dff_B_QLKb3DCw2_2;
	wire w_dff_B_kbi6UYoJ0_2;
	wire w_dff_B_W9BWA3aT2_2;
	wire w_dff_B_p8H4l33e3_2;
	wire w_dff_B_DhC8iWBV8_2;
	wire w_dff_B_MHEttRoN0_2;
	wire w_dff_B_YjRiMxhe4_2;
	wire w_dff_B_kpnditTe6_2;
	wire w_dff_B_eN0tyKXH9_2;
	wire w_dff_B_p2tJ8tsJ5_2;
	wire w_dff_B_5AH076gK6_2;
	wire w_dff_B_Bf1i3PuS7_2;
	wire w_dff_B_6y5Is34i5_2;
	wire w_dff_B_2NieMKZc8_2;
	wire w_dff_B_VUAU0JZs5_2;
	wire w_dff_B_NBxWaCyk3_2;
	wire w_dff_B_fsZIy8ab7_2;
	wire w_dff_B_Lk7lfpJo0_2;
	wire w_dff_B_9Ia7o4WF4_2;
	wire w_dff_B_xK3sLJvh1_2;
	wire w_dff_B_ReanFiuq9_1;
	wire w_dff_B_kd5W7eq48_2;
	wire w_dff_B_bSqiJIAL2_2;
	wire w_dff_B_s9AVR4QJ7_2;
	wire w_dff_B_uOvxAZgz8_2;
	wire w_dff_B_yCNIsvPl7_2;
	wire w_dff_B_4gRAYFMp6_2;
	wire w_dff_B_1HFBDYUU6_2;
	wire w_dff_B_p5h5Y9lv0_2;
	wire w_dff_B_n8BAi0lj0_2;
	wire w_dff_B_IZZl6UlQ7_2;
	wire w_dff_B_TtO1xaW49_2;
	wire w_dff_B_L92VncoI1_2;
	wire w_dff_B_knM46jCd4_2;
	wire w_dff_B_k9r9QfiP1_2;
	wire w_dff_B_i9B2Xl7L9_2;
	wire w_dff_B_077RMbcc9_2;
	wire w_dff_B_z9sBgvdy8_2;
	wire w_dff_B_jVRchJe06_2;
	wire w_dff_B_ZMeHh2362_2;
	wire w_dff_B_0vpAugcX0_2;
	wire w_dff_B_RlEOiPQl5_2;
	wire w_dff_B_JJxAOLQ72_2;
	wire w_dff_B_VflyZQf91_2;
	wire w_dff_B_3GwdQ9y38_2;
	wire w_dff_B_NYtYSTII0_2;
	wire w_dff_B_A2GR43w15_2;
	wire w_dff_B_bh7xWzCl8_2;
	wire w_dff_B_rV1Cd45P9_2;
	wire w_dff_B_FPPMKExE6_2;
	wire w_dff_B_M8ZdatmK8_2;
	wire w_dff_B_FqWQonU96_2;
	wire w_dff_B_PakFZR2O0_2;
	wire w_dff_B_mkgt8N1q3_2;
	wire w_dff_B_tJknHRp68_2;
	wire w_dff_B_yzHuByxt2_2;
	wire w_dff_B_7ojqKWlw1_2;
	wire w_dff_B_NQ7tOS5e6_2;
	wire w_dff_B_7fn1wqLK1_2;
	wire w_dff_B_veTUZf680_1;
	wire w_dff_B_1MFlNQlG1_2;
	wire w_dff_B_0eN4ZT366_2;
	wire w_dff_B_4ojSBjCe6_2;
	wire w_dff_B_zo6D3ETH3_2;
	wire w_dff_B_KruONTMx9_2;
	wire w_dff_B_o0qIjMcI0_2;
	wire w_dff_B_WiooH75D1_2;
	wire w_dff_B_J5bK2PNU9_2;
	wire w_dff_B_8mZNg4Bt8_2;
	wire w_dff_B_sPXgLBGy4_2;
	wire w_dff_B_RljsrN7P1_2;
	wire w_dff_B_4kslgDHs2_2;
	wire w_dff_B_iL4uqpSt0_2;
	wire w_dff_B_lSTVk3zs6_2;
	wire w_dff_B_bndFLteT9_2;
	wire w_dff_B_XFXya9ej0_2;
	wire w_dff_B_7UGjaJmc3_2;
	wire w_dff_B_NyH3w9a65_2;
	wire w_dff_B_Cfij2J5D3_2;
	wire w_dff_B_hxt3pRNb1_2;
	wire w_dff_B_iZ9qV8Xy0_2;
	wire w_dff_B_lRQXa5jr7_2;
	wire w_dff_B_Mp2o1zNl5_2;
	wire w_dff_B_oRPwrnrs1_2;
	wire w_dff_B_SNSed7v20_2;
	wire w_dff_B_ilCQwkt75_2;
	wire w_dff_B_rdJAEZub9_2;
	wire w_dff_B_SOy1ZkQG2_2;
	wire w_dff_B_Ucw9Lnho8_2;
	wire w_dff_B_xpm8tpan2_2;
	wire w_dff_B_bbJOOXCc6_2;
	wire w_dff_B_qHtDA7VN9_2;
	wire w_dff_B_j4Sgkr0I9_2;
	wire w_dff_B_oW3OI4Cm9_2;
	wire w_dff_B_k1sYNB9t6_2;
	wire w_dff_B_zMMYx8m05_1;
	wire w_dff_B_hLjqSoFN7_2;
	wire w_dff_B_APoPfVjO3_2;
	wire w_dff_B_Bra40SYJ4_2;
	wire w_dff_B_uHVFLnpZ9_2;
	wire w_dff_B_JYAUm4iW2_2;
	wire w_dff_B_LCVNXzDv4_2;
	wire w_dff_B_kjKg7emo8_2;
	wire w_dff_B_51pMvQNO7_2;
	wire w_dff_B_jd3hHe7a2_2;
	wire w_dff_B_ggBOShHj9_2;
	wire w_dff_B_HwbKrmSb1_2;
	wire w_dff_B_EET26NwP6_2;
	wire w_dff_B_bgYwDUoa3_2;
	wire w_dff_B_ELpMcuE14_2;
	wire w_dff_B_KcuxWioZ5_2;
	wire w_dff_B_0dGhzTqP6_2;
	wire w_dff_B_7ghHuPuN3_2;
	wire w_dff_B_ebQO4LoM7_2;
	wire w_dff_B_o0GDCZ3h2_2;
	wire w_dff_B_xDjETYky4_2;
	wire w_dff_B_AsUrr5bl6_2;
	wire w_dff_B_NqiSNVvD0_2;
	wire w_dff_B_9x5qZPpR0_2;
	wire w_dff_B_Pu9DKG484_2;
	wire w_dff_B_8LSz4q5N1_2;
	wire w_dff_B_uHWOdmql1_2;
	wire w_dff_B_mlwlzIqc9_2;
	wire w_dff_B_w0kTrk9X0_2;
	wire w_dff_B_GtifgqIH0_2;
	wire w_dff_B_9lXJlrPk0_2;
	wire w_dff_B_MZeffkU02_2;
	wire w_dff_B_NrvwmNJd9_2;
	wire w_dff_B_HCj8WZ5M8_1;
	wire w_dff_B_1nUfeMI19_2;
	wire w_dff_B_r4TgFsLg4_2;
	wire w_dff_B_U7eK7ras0_2;
	wire w_dff_B_zrvC81M98_2;
	wire w_dff_B_27TquYjo6_2;
	wire w_dff_B_TRzeehci4_2;
	wire w_dff_B_FADVWIPW6_2;
	wire w_dff_B_owwTMn0U6_2;
	wire w_dff_B_6k6UJhV44_2;
	wire w_dff_B_wf9KYBtm9_2;
	wire w_dff_B_dpSXt6cN0_2;
	wire w_dff_B_WmjDN2X53_2;
	wire w_dff_B_9rOUK7gv4_2;
	wire w_dff_B_0ntmxdeh9_2;
	wire w_dff_B_IYb19NAp3_2;
	wire w_dff_B_BNwk8ty04_2;
	wire w_dff_B_SVIbwp204_2;
	wire w_dff_B_7TVy182l6_2;
	wire w_dff_B_BdpKSbg85_2;
	wire w_dff_B_3E69npys3_2;
	wire w_dff_B_gUBw3JOx5_2;
	wire w_dff_B_pQ6i6UA62_2;
	wire w_dff_B_OcfXnWdd8_2;
	wire w_dff_B_VJgSELb14_2;
	wire w_dff_B_67gh5KcN0_2;
	wire w_dff_B_NrHTQXjL7_2;
	wire w_dff_B_UzLe5UKv6_2;
	wire w_dff_B_za3ROloz1_2;
	wire w_dff_B_fkjO06sJ2_2;
	wire w_dff_B_oNQaC9jL0_1;
	wire w_dff_B_JhXoKu6z7_2;
	wire w_dff_B_Cch5dsic8_2;
	wire w_dff_B_LFIHne1m0_2;
	wire w_dff_B_u9d8O3ND9_2;
	wire w_dff_B_Ov5TIUFx9_2;
	wire w_dff_B_RqyCoBIX2_2;
	wire w_dff_B_OFcUnF6F3_2;
	wire w_dff_B_0zouLgnG1_2;
	wire w_dff_B_toc16hBi5_2;
	wire w_dff_B_TXI1F9mV5_2;
	wire w_dff_B_btvoys767_2;
	wire w_dff_B_ubAH73YH1_2;
	wire w_dff_B_WKnDMv1C8_2;
	wire w_dff_B_WbdYm6aS0_2;
	wire w_dff_B_CPeD9D6j4_2;
	wire w_dff_B_OkSrRGy12_2;
	wire w_dff_B_RUrXO1uE5_2;
	wire w_dff_B_OpurLFzk8_2;
	wire w_dff_B_6k1b1P5b2_2;
	wire w_dff_B_qcQUQ9rg3_2;
	wire w_dff_B_4Cjcde9o2_2;
	wire w_dff_B_OyySodQ52_2;
	wire w_dff_B_Ni0jIFDv4_2;
	wire w_dff_B_jtDwDZT59_2;
	wire w_dff_B_w04eOjon8_2;
	wire w_dff_B_TPz8dDkP1_2;
	wire w_dff_B_T5RspWwv6_1;
	wire w_dff_B_fSNe4Gi35_2;
	wire w_dff_B_MGVDY3nQ9_2;
	wire w_dff_B_LKhWCFMS9_2;
	wire w_dff_B_JvBHsJIQ3_2;
	wire w_dff_B_os76MLwk6_2;
	wire w_dff_B_tUa7eqWR4_2;
	wire w_dff_B_R9yK3csS1_2;
	wire w_dff_B_eqDiBzSp9_2;
	wire w_dff_B_XwtrnRCF6_2;
	wire w_dff_B_hsqfgo138_2;
	wire w_dff_B_lkSsZcwb9_2;
	wire w_dff_B_fYJXpoVy8_2;
	wire w_dff_B_8kgu35s13_2;
	wire w_dff_B_AWLHZFl22_2;
	wire w_dff_B_NNc4Skoq2_2;
	wire w_dff_B_UnMGkXVj1_2;
	wire w_dff_B_Oa8tzeVT3_2;
	wire w_dff_B_y4oUdMDz2_2;
	wire w_dff_B_j68deaQ98_2;
	wire w_dff_B_mBouTcgA7_2;
	wire w_dff_B_HU2a7Mqb4_2;
	wire w_dff_B_lXtCB2Gg5_2;
	wire w_dff_B_y0jHMrmq7_2;
	wire w_dff_B_o0IytErQ1_1;
	wire w_dff_B_ucXkrZDx5_2;
	wire w_dff_B_ydJOXd4d9_2;
	wire w_dff_B_LWpnIXHO7_2;
	wire w_dff_B_Bcbw6A0V4_2;
	wire w_dff_B_qoT6i7rj0_2;
	wire w_dff_B_LDqagPD31_2;
	wire w_dff_B_WAjYjVyj0_2;
	wire w_dff_B_C9xGoUl13_2;
	wire w_dff_B_qmBgromb0_2;
	wire w_dff_B_PYnyeRYe8_2;
	wire w_dff_B_F3Z9RT8L7_2;
	wire w_dff_B_9LT574Eg5_2;
	wire w_dff_B_y8MtH8ep3_2;
	wire w_dff_B_7NlvxpPL2_2;
	wire w_dff_B_XPNeS3VR2_2;
	wire w_dff_B_wEMM3LnP6_2;
	wire w_dff_B_YWnGqG0v9_2;
	wire w_dff_B_w8wLh6XU3_2;
	wire w_dff_B_NH7vxheQ8_2;
	wire w_dff_B_PUBqbE3j7_2;
	wire w_dff_B_6lk4vICq9_1;
	wire w_dff_B_u2ild03L2_2;
	wire w_dff_B_ZeVZeRrl4_2;
	wire w_dff_B_W4FDz4uA4_2;
	wire w_dff_B_STI5qzlE4_2;
	wire w_dff_B_HPYReZu66_2;
	wire w_dff_B_jdO8fL5H8_2;
	wire w_dff_B_fKNculjk0_2;
	wire w_dff_B_J7DP4vnD7_2;
	wire w_dff_B_oUbEnMrs0_2;
	wire w_dff_B_x8DoXHst6_2;
	wire w_dff_B_7PvO9cLP0_2;
	wire w_dff_B_RPRND2GF9_2;
	wire w_dff_B_JI98W9DV0_2;
	wire w_dff_B_wWwjP0kI7_2;
	wire w_dff_B_g8Jwdm8a4_2;
	wire w_dff_B_odjSL4HC4_2;
	wire w_dff_B_CqLjs5BL4_2;
	wire w_dff_B_xT0WLZwq2_1;
	wire w_dff_B_RKKdMgNN3_2;
	wire w_dff_B_0DpLjLmY6_2;
	wire w_dff_B_v29ksKNL0_2;
	wire w_dff_B_G98R3u7e8_2;
	wire w_dff_B_gXyykDV45_2;
	wire w_dff_B_oCySopo13_2;
	wire w_dff_B_BdqtUJ2l9_2;
	wire w_dff_B_tT89ZdvF9_2;
	wire w_dff_B_3oAWeIJS4_2;
	wire w_dff_B_AQuR4vss1_2;
	wire w_dff_B_hBQ9ltan8_2;
	wire w_dff_B_vYU6pmby5_2;
	wire w_dff_B_zfj2YvDS8_2;
	wire w_dff_B_nj6Se62c5_2;
	wire w_dff_B_TaolNwSg5_1;
	wire w_dff_B_XOMwYQ1g5_2;
	wire w_dff_B_RjhhO5uD1_2;
	wire w_dff_B_aOsYWP852_2;
	wire w_dff_B_faJLiB5J2_2;
	wire w_dff_B_GLqZUqOV1_2;
	wire w_dff_B_XGMTY2iG4_2;
	wire w_dff_B_cT7NVXqe5_2;
	wire w_dff_B_5TKpctYA4_2;
	wire w_dff_B_VsouEbG68_2;
	wire w_dff_B_kXxIFRYn3_2;
	wire w_dff_B_LhM19GdE6_2;
	wire w_dff_B_63xYh7mI9_1;
	wire w_dff_B_lUvToWTD5_2;
	wire w_dff_B_nT9XyHk90_2;
	wire w_dff_B_fAvqAzWA9_2;
	wire w_dff_B_ziFl5Luj2_2;
	wire w_dff_B_0jAIa8Ra8_2;
	wire w_dff_B_nOvOlYwI9_2;
	wire w_dff_B_8cqyc2hd9_2;
	wire w_dff_B_NuTfgCbl3_2;
	wire w_dff_B_840c3GDk4_1;
	wire w_dff_B_y5d7qXEA7_0;
	wire w_dff_B_MvKZ4hK44_2;
	wire w_dff_B_i0AiXt3t0_2;
	wire w_dff_B_bLePfPt96_2;
	wire w_dff_B_MwjjekUY8_2;
	wire w_dff_B_KKHmuLIX0_1;
	wire w_dff_A_8E5w6H2V9_0;
	wire w_dff_A_kW5i3c4R9_0;
	wire w_dff_A_fhzCCFL74_1;
	wire w_dff_B_FYr4FdfB3_1;
	wire w_dff_B_97dahFt13_2;
	wire w_dff_B_kM2w0pJj4_2;
	wire w_dff_B_sdvDUFMH0_2;
	wire w_dff_B_ye70Y0S27_2;
	wire w_dff_B_tOA5M8gj2_2;
	wire w_dff_B_canzLa4y0_2;
	wire w_dff_B_z2WiqUud6_2;
	wire w_dff_B_wb7ixjfM7_2;
	wire w_dff_B_KOEcrsUM2_2;
	wire w_dff_B_eZqMxb2o3_2;
	wire w_dff_B_lxWqMd960_2;
	wire w_dff_B_Vzi2AMkV3_2;
	wire w_dff_B_yjBAKb3p0_2;
	wire w_dff_B_1QmP0zAE6_2;
	wire w_dff_B_Clfefpkr0_2;
	wire w_dff_B_wvS48xXe8_2;
	wire w_dff_B_FMFdajSE8_2;
	wire w_dff_B_F0U9BQuG0_2;
	wire w_dff_B_jp4O6DnO3_2;
	wire w_dff_B_NpJKpymw5_2;
	wire w_dff_B_NWlGvxaR1_2;
	wire w_dff_B_BRLxfiIB6_2;
	wire w_dff_B_Xnznz3Hc7_2;
	wire w_dff_B_IkTFQmgJ4_2;
	wire w_dff_B_xfdBIZhg2_2;
	wire w_dff_B_zHvjn4iN1_2;
	wire w_dff_B_Vsu5ghWg6_2;
	wire w_dff_B_daI5tDWJ4_2;
	wire w_dff_B_tqj6Turq9_2;
	wire w_dff_B_yWe4buxL1_2;
	wire w_dff_B_ojg5zu0o8_2;
	wire w_dff_B_tvYn0OcY7_2;
	wire w_dff_B_pfHaJ1on5_2;
	wire w_dff_B_eFlPGGgw9_2;
	wire w_dff_B_wTqoOGBS9_2;
	wire w_dff_B_1w1TVNSQ3_2;
	wire w_dff_B_SN7CToZX4_2;
	wire w_dff_B_2azUBcUx4_2;
	wire w_dff_B_Uh8vgPYg3_2;
	wire w_dff_B_UjghNXSM2_2;
	wire w_dff_B_Vl97vaTn6_2;
	wire w_dff_B_P26eiy1G5_2;
	wire w_dff_B_NO15k2Oc6_2;
	wire w_dff_B_QNpmEh2r7_2;
	wire w_dff_B_TkXN03tm1_2;
	wire w_dff_B_ErSGtDO89_0;
	wire w_dff_A_kYtAJoyj3_1;
	wire w_dff_B_PO12R7st0_1;
	wire w_dff_B_G1maRCRW3_2;
	wire w_dff_B_Q64g7U0e7_2;
	wire w_dff_B_UbQ2xhCw9_2;
	wire w_dff_B_GchuL2Ck6_2;
	wire w_dff_B_Y2h6OELG8_2;
	wire w_dff_B_SmnIKM9c9_2;
	wire w_dff_B_T6OUy6Wr5_2;
	wire w_dff_B_MAVHHYY07_2;
	wire w_dff_B_nI5hRsFM4_2;
	wire w_dff_B_VPiU3bUU2_2;
	wire w_dff_B_VO0rdYS86_2;
	wire w_dff_B_xnIqzth18_2;
	wire w_dff_B_PHhCAjey3_2;
	wire w_dff_B_gYLMXeYr0_2;
	wire w_dff_B_sfVftEcX5_2;
	wire w_dff_B_iHWmKDPY2_2;
	wire w_dff_B_lWA7B3iK7_2;
	wire w_dff_B_G23HMgzn4_2;
	wire w_dff_B_ucLvddoU5_2;
	wire w_dff_B_nvPwtDLH3_2;
	wire w_dff_B_XMI1GGMD8_2;
	wire w_dff_B_dj8YkQ9B8_2;
	wire w_dff_B_neCjZH8g0_2;
	wire w_dff_B_mwiq29ZP1_2;
	wire w_dff_B_oWVLYtYp5_2;
	wire w_dff_B_2ph7WAf20_2;
	wire w_dff_B_To9WhxcV1_2;
	wire w_dff_B_xPwgAhsL9_2;
	wire w_dff_B_uXZKAVL43_2;
	wire w_dff_B_nfefX84y6_2;
	wire w_dff_B_bLHxjmhz6_2;
	wire w_dff_B_yBHXCI0G8_2;
	wire w_dff_B_6Xd9MZD60_2;
	wire w_dff_B_xHJA97rU7_2;
	wire w_dff_B_O3NERh0V7_2;
	wire w_dff_B_VeJfhk6p7_2;
	wire w_dff_B_w5VGHhFp4_2;
	wire w_dff_B_hcXKlHQ22_2;
	wire w_dff_B_x3gphihD4_2;
	wire w_dff_B_C1CopPj13_2;
	wire w_dff_B_yl0l0a1u5_2;
	wire w_dff_B_1FdTulTQ5_1;
	wire w_dff_B_WDUMuBKs2_2;
	wire w_dff_B_tHPoC6bH8_2;
	wire w_dff_B_iuPXHBei1_2;
	wire w_dff_B_wOLEZ0023_2;
	wire w_dff_B_3CbNm7mZ3_2;
	wire w_dff_B_33K1CaVa9_2;
	wire w_dff_B_NuYLS1BX4_2;
	wire w_dff_B_NG9JutYO9_2;
	wire w_dff_B_tMct18bU3_2;
	wire w_dff_B_6ytrvTXf3_2;
	wire w_dff_B_J0a2xsRx4_2;
	wire w_dff_B_qOZOIK6A6_2;
	wire w_dff_B_FrL6L2WZ9_2;
	wire w_dff_B_1Hhp8gWr8_2;
	wire w_dff_B_wybK3zaP9_2;
	wire w_dff_B_e4Ywqcf42_2;
	wire w_dff_B_T4vBLDra3_2;
	wire w_dff_B_vVwrYBw38_2;
	wire w_dff_B_Bb3YooaZ9_2;
	wire w_dff_B_J64LuYsM8_2;
	wire w_dff_B_pcviOWKM5_2;
	wire w_dff_B_YSQZGqYA8_2;
	wire w_dff_B_LTyKT05K8_2;
	wire w_dff_B_ZbNZszgQ1_2;
	wire w_dff_B_xCevtBru7_2;
	wire w_dff_B_Z1Yh5kcX9_2;
	wire w_dff_B_zYtxJ5f01_2;
	wire w_dff_B_pSBAOqev4_2;
	wire w_dff_B_qjoQU56g2_2;
	wire w_dff_B_doZPJe446_2;
	wire w_dff_B_fBFLnPRJ9_2;
	wire w_dff_B_R8Mu0ulb9_2;
	wire w_dff_B_xcIS3Db01_2;
	wire w_dff_B_LDj1WWAe8_2;
	wire w_dff_B_eQ3WmxFV6_2;
	wire w_dff_B_50d97sJh9_2;
	wire w_dff_B_SPEl12Do8_2;
	wire w_dff_B_dwHvenCd1_2;
	wire w_dff_B_e7fGPhgE3_1;
	wire w_dff_B_LmsiQImZ3_2;
	wire w_dff_B_8CLIK6zu7_2;
	wire w_dff_B_4bWhRPM23_2;
	wire w_dff_B_6YuIOJ1G8_2;
	wire w_dff_B_OuAbxXVj7_2;
	wire w_dff_B_rTGNjhvs5_2;
	wire w_dff_B_IzYZFxIU4_2;
	wire w_dff_B_1h37I6P49_2;
	wire w_dff_B_b7RuuJtX6_2;
	wire w_dff_B_rq5qyBfF8_2;
	wire w_dff_B_WNWLDnI84_2;
	wire w_dff_B_cO8QrZAa1_2;
	wire w_dff_B_msLjvfIU6_2;
	wire w_dff_B_MGLBF5eC1_2;
	wire w_dff_B_lDkGGy7K7_2;
	wire w_dff_B_TeVGVNDj4_2;
	wire w_dff_B_cwoCL9eg1_2;
	wire w_dff_B_GQukG6X37_2;
	wire w_dff_B_J239FyPX1_2;
	wire w_dff_B_sA8k7kSF3_2;
	wire w_dff_B_RDMpURB99_2;
	wire w_dff_B_5iE0CbGz1_2;
	wire w_dff_B_PX3zf5Gz8_2;
	wire w_dff_B_IhNFsn7B3_2;
	wire w_dff_B_pORJCIuw4_2;
	wire w_dff_B_wGuVFKaH5_2;
	wire w_dff_B_3uCZmPoo8_2;
	wire w_dff_B_gPlS9qr43_2;
	wire w_dff_B_ktyEjLTY7_2;
	wire w_dff_B_9CtZTChJ3_2;
	wire w_dff_B_Fhb1x64I8_2;
	wire w_dff_B_5hKuInnK9_2;
	wire w_dff_B_hws0KtPy6_2;
	wire w_dff_B_65svk5wf5_2;
	wire w_dff_B_j5PCsBuH8_2;
	wire w_dff_B_pBI9Lvgg8_1;
	wire w_dff_B_wzDJ8GCf6_2;
	wire w_dff_B_OpDI0DFm5_2;
	wire w_dff_B_IvLQERmA4_2;
	wire w_dff_B_TOp3wvWf0_2;
	wire w_dff_B_A3nHQHCi0_2;
	wire w_dff_B_B3ko1R7p6_2;
	wire w_dff_B_fNYjTCIu3_2;
	wire w_dff_B_SOwTlDjF2_2;
	wire w_dff_B_TCvgAghv5_2;
	wire w_dff_B_iyMBxWQQ9_2;
	wire w_dff_B_D5ACEWdk6_2;
	wire w_dff_B_IHkhM8kn8_2;
	wire w_dff_B_ZhaEjqcn4_2;
	wire w_dff_B_8eldP4aa5_2;
	wire w_dff_B_UAtNCGJR1_2;
	wire w_dff_B_Pb1SEEpV5_2;
	wire w_dff_B_VZjmkF8E2_2;
	wire w_dff_B_SQ1korkG5_2;
	wire w_dff_B_rKvf5muT9_2;
	wire w_dff_B_Zjp6PeYn3_2;
	wire w_dff_B_8iRFxlKX4_2;
	wire w_dff_B_bPyhQSOP4_2;
	wire w_dff_B_Wtx5tA226_2;
	wire w_dff_B_Vh4MYR6s0_2;
	wire w_dff_B_UBhSE7YF7_2;
	wire w_dff_B_Q9jpslpw3_2;
	wire w_dff_B_L2o0Hqbn7_2;
	wire w_dff_B_8bwieWx31_2;
	wire w_dff_B_lL1GPZWx1_2;
	wire w_dff_B_d5zoKY9j2_2;
	wire w_dff_B_FvJ5VlAH2_2;
	wire w_dff_B_r0eWN7pX6_2;
	wire w_dff_B_ts1N6ri07_1;
	wire w_dff_B_YqdZnYp53_2;
	wire w_dff_B_kmMz4Gf42_2;
	wire w_dff_B_43mAdFk75_2;
	wire w_dff_B_6i7Y3gjJ6_2;
	wire w_dff_B_TPqjHbOt1_2;
	wire w_dff_B_gPv13XMD8_2;
	wire w_dff_B_JDbgwmlQ8_2;
	wire w_dff_B_nxTYpnUK8_2;
	wire w_dff_B_bRG6w92b1_2;
	wire w_dff_B_uullTJNc3_2;
	wire w_dff_B_Vchd5S709_2;
	wire w_dff_B_lYzj0mSx3_2;
	wire w_dff_B_OTVnSV1y4_2;
	wire w_dff_B_X9qIEM6a7_2;
	wire w_dff_B_jyz3z9Kz0_2;
	wire w_dff_B_Zq7N5mJb5_2;
	wire w_dff_B_VCjJqEBn3_2;
	wire w_dff_B_yenbJd053_2;
	wire w_dff_B_xulcjw5X0_2;
	wire w_dff_B_evc9jos05_2;
	wire w_dff_B_5SfTaJ0x0_2;
	wire w_dff_B_QUB7MmDY1_2;
	wire w_dff_B_aOnfFLsY0_2;
	wire w_dff_B_WLQ1ZuIR2_2;
	wire w_dff_B_jAPbVsbm7_2;
	wire w_dff_B_E0p2adVD9_2;
	wire w_dff_B_ZNy59xiD0_2;
	wire w_dff_B_vREFlxaq6_2;
	wire w_dff_B_6ugO9nhT4_2;
	wire w_dff_B_ScF5DwwC9_1;
	wire w_dff_B_PvOC5jrK0_2;
	wire w_dff_B_4tPRFRgg6_2;
	wire w_dff_B_kudyrlO27_2;
	wire w_dff_B_qfalpslK9_2;
	wire w_dff_B_V3HQj16c1_2;
	wire w_dff_B_QDyQD9Zb0_2;
	wire w_dff_B_DaCLurpc9_2;
	wire w_dff_B_6QTSgAb25_2;
	wire w_dff_B_2euEQrjF8_2;
	wire w_dff_B_paSe0hMp1_2;
	wire w_dff_B_n5Tgybgr7_2;
	wire w_dff_B_xsJ9fH2c7_2;
	wire w_dff_B_oXKF7KbU7_2;
	wire w_dff_B_uEedBUuE2_2;
	wire w_dff_B_iKwcjPnB7_2;
	wire w_dff_B_ou0gdfKh1_2;
	wire w_dff_B_myqiBtY24_2;
	wire w_dff_B_SKuD2mDk0_2;
	wire w_dff_B_oDNeadf12_2;
	wire w_dff_B_IPPejWRp4_2;
	wire w_dff_B_3TBBLLiv7_2;
	wire w_dff_B_KRrt0mCn7_2;
	wire w_dff_B_v7HP5egH3_2;
	wire w_dff_B_l2K1yHub2_2;
	wire w_dff_B_2n9qfHGe5_2;
	wire w_dff_B_Jf9q3FuV5_2;
	wire w_dff_B_ambeZDru3_1;
	wire w_dff_B_pT211enw6_2;
	wire w_dff_B_5RbJpCSr5_2;
	wire w_dff_B_BnSh8e9n1_2;
	wire w_dff_B_Oa3AfMKN1_2;
	wire w_dff_B_FUq7BMzz2_2;
	wire w_dff_B_69ytwXJt8_2;
	wire w_dff_B_kAl9rvsN4_2;
	wire w_dff_B_4ccqOJDd4_2;
	wire w_dff_B_Shtvuj1w8_2;
	wire w_dff_B_4irAzCcn9_2;
	wire w_dff_B_cc4iG2Le1_2;
	wire w_dff_B_Acxl081n6_2;
	wire w_dff_B_fWheg23y9_2;
	wire w_dff_B_NKNkC2Cm6_2;
	wire w_dff_B_GS2PR2bm7_2;
	wire w_dff_B_rV9VqsnX6_2;
	wire w_dff_B_WGkWsx5q0_2;
	wire w_dff_B_u1wLJopG9_2;
	wire w_dff_B_MwQPq3qX3_2;
	wire w_dff_B_F2UjT6mZ9_2;
	wire w_dff_B_j4WSWt6l8_2;
	wire w_dff_B_YtxsDGOU2_2;
	wire w_dff_B_smBEFrpg5_2;
	wire w_dff_B_7S1vnxda9_1;
	wire w_dff_B_uWHYvu380_2;
	wire w_dff_B_LJhkuRgl3_2;
	wire w_dff_B_mvKh69Z53_2;
	wire w_dff_B_F6qK8rmi9_2;
	wire w_dff_B_cwclJGCG1_2;
	wire w_dff_B_izOQKGti7_2;
	wire w_dff_B_FS2E4zBV6_2;
	wire w_dff_B_9SNvCuRv9_2;
	wire w_dff_B_xQyJCR9W3_2;
	wire w_dff_B_RgON4shO5_2;
	wire w_dff_B_XmO9pUmN1_2;
	wire w_dff_B_rIKw22Tb8_2;
	wire w_dff_B_zCITm22H5_2;
	wire w_dff_B_u899r1GP3_2;
	wire w_dff_B_UVKIPfSg1_2;
	wire w_dff_B_uhNwhAlK3_2;
	wire w_dff_B_zq1Xb35I2_2;
	wire w_dff_B_TryxKBJx8_2;
	wire w_dff_B_6D0AnOxI9_2;
	wire w_dff_B_60jCzz1X6_2;
	wire w_dff_B_0ub2UGTJ6_1;
	wire w_dff_B_hZP5Pcea3_2;
	wire w_dff_B_xaF7K1LR1_2;
	wire w_dff_B_6NBxfdrw1_2;
	wire w_dff_B_DzFcIKYo9_2;
	wire w_dff_B_cIXviL1N7_2;
	wire w_dff_B_GKUwsO8n9_2;
	wire w_dff_B_zQ5YPaKt5_2;
	wire w_dff_B_A8lGErrZ9_2;
	wire w_dff_B_7PCCRPQf4_2;
	wire w_dff_B_XFS9fUwq4_2;
	wire w_dff_B_04UenHlJ6_2;
	wire w_dff_B_VJuDTfFt3_2;
	wire w_dff_B_Lh6ghqtr8_2;
	wire w_dff_B_BkLOlcoO5_2;
	wire w_dff_B_GoYdnHUq3_2;
	wire w_dff_B_DMYriVf68_2;
	wire w_dff_B_99G06CEw4_2;
	wire w_dff_B_VavVFlVG0_1;
	wire w_dff_B_l6lJxTBy4_2;
	wire w_dff_B_Zu9RzIMr3_2;
	wire w_dff_B_meauC6jk3_2;
	wire w_dff_B_F4RgRU7D9_2;
	wire w_dff_B_XRQJSKkf0_2;
	wire w_dff_B_bzJFWsZ66_2;
	wire w_dff_B_2Rga0I6R9_2;
	wire w_dff_B_Q8fkGh5e6_2;
	wire w_dff_B_y92OjV0m5_2;
	wire w_dff_B_Z2uRmlb57_2;
	wire w_dff_B_ENARae1N1_2;
	wire w_dff_B_BW0Xlbkn2_2;
	wire w_dff_B_z3z38aMv1_2;
	wire w_dff_B_mh08k7Jk4_2;
	wire w_dff_B_wBflJaNu9_1;
	wire w_dff_B_Hg4HGYb48_2;
	wire w_dff_B_EGYQy1GI8_2;
	wire w_dff_B_wtoysNb52_2;
	wire w_dff_B_nnmYLzoN4_2;
	wire w_dff_B_BgbXiQmy6_2;
	wire w_dff_B_5DaD8okL6_2;
	wire w_dff_B_1qb0wsjc3_2;
	wire w_dff_B_2OvjnneS9_2;
	wire w_dff_B_MOR0XDjc2_2;
	wire w_dff_B_Fh9L8oXW3_2;
	wire w_dff_B_3l4SKcDE9_2;
	wire w_dff_B_4pUskhmR3_1;
	wire w_dff_B_Zffz6OVe5_2;
	wire w_dff_B_mqFqbXDs5_2;
	wire w_dff_B_eDp7MZDI5_2;
	wire w_dff_B_90Go2Bhy0_2;
	wire w_dff_B_8ojogRrX5_2;
	wire w_dff_B_i3BNk4I12_2;
	wire w_dff_B_NzaK6og78_2;
	wire w_dff_B_2ZFijG8y4_2;
	wire w_dff_B_KmYDFXAP3_1;
	wire w_dff_B_K5WYOovD9_0;
	wire w_dff_B_NYY6r2fA2_2;
	wire w_dff_B_e0vTI1iP1_2;
	wire w_dff_B_tnEQxkZm4_2;
	wire w_dff_B_sgCcalFI4_2;
	wire w_dff_B_4EFGqvCf7_1;
	wire w_dff_A_1dikcfgM7_0;
	wire w_dff_A_vdeHAEpJ2_0;
	wire w_dff_A_S5jpLcNQ9_0;
	wire w_dff_A_0436c07I2_1;
	wire w_dff_B_16GkUzZv0_2;
	wire w_dff_B_LlyAvuTl5_1;
	wire w_dff_B_oEuP862p2_2;
	wire w_dff_B_2FCJ6bpK1_2;
	wire w_dff_B_qXX7wsY90_2;
	wire w_dff_B_MnL8R5MZ8_2;
	wire w_dff_B_rmY4Ptp70_2;
	wire w_dff_B_8ctsjS5W8_2;
	wire w_dff_B_BoSfgg6J1_2;
	wire w_dff_B_QdedzU871_2;
	wire w_dff_B_0UnuHLDC7_2;
	wire w_dff_B_eNHY3aZ41_2;
	wire w_dff_B_OYthKwP47_2;
	wire w_dff_B_N22Abqi71_2;
	wire w_dff_B_nS1bcpwc5_2;
	wire w_dff_B_zVmWG6I28_2;
	wire w_dff_B_aWVtrNGj7_2;
	wire w_dff_B_zyJ1kUiO0_2;
	wire w_dff_B_j02usAVa0_2;
	wire w_dff_B_4SqEQTPA9_2;
	wire w_dff_B_Ur1Yvhqh7_2;
	wire w_dff_B_ttgQNeSP6_2;
	wire w_dff_B_RTUYvkxv7_2;
	wire w_dff_B_VChcbkYF1_2;
	wire w_dff_B_Mymb4dbm0_2;
	wire w_dff_B_MRo1fH5Q9_2;
	wire w_dff_B_Cad5qNF82_2;
	wire w_dff_B_b1nxdM0V6_2;
	wire w_dff_B_NwW9LOgV5_2;
	wire w_dff_B_BunGjR6r7_2;
	wire w_dff_B_FsOwk66u3_2;
	wire w_dff_B_uNqCDQEp1_2;
	wire w_dff_B_uhVxvnRV0_2;
	wire w_dff_B_8jOKIvXi1_2;
	wire w_dff_B_7N7nnwl53_2;
	wire w_dff_B_DVINhr4B0_2;
	wire w_dff_B_4hZRj11s0_2;
	wire w_dff_B_eFxfwSUJ7_2;
	wire w_dff_B_aiTdjmL76_2;
	wire w_dff_B_K0232ANi8_2;
	wire w_dff_B_te5GG3Dy5_2;
	wire w_dff_B_F2cji9dj0_2;
	wire w_dff_B_1AcWBykD1_2;
	wire w_dff_B_3WeEeyUq7_2;
	wire w_dff_B_nP6Q6lid7_2;
	wire w_dff_B_HBO5oRPH1_2;
	wire w_dff_B_CAjFbE2G4_2;
	wire w_dff_B_pdJuQq7B8_1;
	wire w_dff_B_chTdOyU17_2;
	wire w_dff_B_Z2Q8o9qI7_2;
	wire w_dff_B_N4xaF1I83_2;
	wire w_dff_B_fnokAywJ5_2;
	wire w_dff_B_NM8bVZpu9_2;
	wire w_dff_B_2liClNdT1_2;
	wire w_dff_B_6NSKfvJq5_2;
	wire w_dff_B_Gvfcs4qJ3_2;
	wire w_dff_B_aB3ZMS1L8_2;
	wire w_dff_B_u9npDKRN6_2;
	wire w_dff_B_B9aHE3oi2_2;
	wire w_dff_B_Ei6sL0dE9_2;
	wire w_dff_B_oo9UdODz6_2;
	wire w_dff_B_tBI6EE1Q0_2;
	wire w_dff_B_tZzyRcw01_2;
	wire w_dff_B_A5maOp4O6_2;
	wire w_dff_B_j1UCzGsH7_2;
	wire w_dff_B_iSYxG9pj5_2;
	wire w_dff_B_UMJ4k9Yu1_2;
	wire w_dff_B_ZDpuUfWg8_2;
	wire w_dff_B_BRKGf0Ev2_2;
	wire w_dff_B_7l7sEoCG9_2;
	wire w_dff_B_nOgqgypv4_2;
	wire w_dff_B_YclXjoTc9_2;
	wire w_dff_B_xatqhX4U5_2;
	wire w_dff_B_M7p0NrRz6_2;
	wire w_dff_B_0TSKVTvp0_2;
	wire w_dff_B_SCIfQhJ49_2;
	wire w_dff_B_gq05zGsY8_2;
	wire w_dff_B_LtheA07r3_2;
	wire w_dff_B_ojVqX1w55_2;
	wire w_dff_B_wSZW6EuG9_2;
	wire w_dff_B_At1IcBmn8_2;
	wire w_dff_B_iGi0t4qg6_2;
	wire w_dff_B_lkkK2CV79_2;
	wire w_dff_B_6ObnPa4j5_2;
	wire w_dff_B_hn6oqsic3_2;
	wire w_dff_B_pzi2CGvT6_2;
	wire w_dff_B_PnKzv59X5_2;
	wire w_dff_B_ohmRqlak2_2;
	wire w_dff_B_lpCrGuqL4_1;
	wire w_dff_B_xMSg6Pv57_2;
	wire w_dff_B_E9U3GXRQ5_2;
	wire w_dff_B_CP7JYHcq8_2;
	wire w_dff_B_L9GOE1g96_2;
	wire w_dff_B_NoW9bIoI4_2;
	wire w_dff_B_YFVVYW8j0_2;
	wire w_dff_B_a0Rvi3PB2_2;
	wire w_dff_B_LBrZgVoU5_2;
	wire w_dff_B_tk3aPc7C7_2;
	wire w_dff_B_u9ssFZvA8_2;
	wire w_dff_B_Fl0OUili8_2;
	wire w_dff_B_hYDrS2Ux9_2;
	wire w_dff_B_DfHYd1zE0_2;
	wire w_dff_B_jqxNP8hZ4_2;
	wire w_dff_B_kuYCNlZG7_2;
	wire w_dff_B_Px6qQJVb1_2;
	wire w_dff_B_VV58nyGG9_2;
	wire w_dff_B_8eEwJLS32_2;
	wire w_dff_B_z2gX4LoL0_2;
	wire w_dff_B_tZ7WiEt35_2;
	wire w_dff_B_kTUwXg5W8_2;
	wire w_dff_B_tTmRNDrj0_2;
	wire w_dff_B_LKiUVsHw3_2;
	wire w_dff_B_LnJBXjGF4_2;
	wire w_dff_B_8ymCK2S00_2;
	wire w_dff_B_l0TVVT9J5_2;
	wire w_dff_B_lnSV6onm5_2;
	wire w_dff_B_oIsHcuvu5_2;
	wire w_dff_B_TD1EOJbO4_2;
	wire w_dff_B_GTscYVNi9_2;
	wire w_dff_B_0Pyrvwmj5_2;
	wire w_dff_B_ReYYuzyW9_2;
	wire w_dff_B_QzHvZwvc8_2;
	wire w_dff_B_nBE31lqW3_2;
	wire w_dff_B_M6j72Ivz5_2;
	wire w_dff_B_tsGImOhK0_2;
	wire w_dff_B_8aqOsc927_2;
	wire w_dff_B_adC3VRFf2_1;
	wire w_dff_B_nZwFZUuS8_2;
	wire w_dff_B_fghC81nT8_2;
	wire w_dff_B_W84BEZuG4_2;
	wire w_dff_B_Q9Kvb8bM8_2;
	wire w_dff_B_n8tv2Y4G5_2;
	wire w_dff_B_MQ79rhWR4_2;
	wire w_dff_B_CLBbNLD51_2;
	wire w_dff_B_HeqE217R7_2;
	wire w_dff_B_vID76VdG3_2;
	wire w_dff_B_ND2md9je1_2;
	wire w_dff_B_a5u4UEfa0_2;
	wire w_dff_B_gb6uSkQw7_2;
	wire w_dff_B_PIyZ6Yf77_2;
	wire w_dff_B_Q9uXNTZf7_2;
	wire w_dff_B_eEQSogE30_2;
	wire w_dff_B_rCIWTCVw9_2;
	wire w_dff_B_C3Y2j74P1_2;
	wire w_dff_B_hNCZ22lm5_2;
	wire w_dff_B_r7At73XZ7_2;
	wire w_dff_B_at497RtK3_2;
	wire w_dff_B_oIaN6k833_2;
	wire w_dff_B_z4ZJdOQc2_2;
	wire w_dff_B_Z3NA1rv65_2;
	wire w_dff_B_O8QjDOkw8_2;
	wire w_dff_B_JSWpm2pQ9_2;
	wire w_dff_B_P6ywCwKw3_2;
	wire w_dff_B_tgNWZzZ02_2;
	wire w_dff_B_NB4urrU51_2;
	wire w_dff_B_5GDDgcpi7_2;
	wire w_dff_B_IxXY4A5c0_2;
	wire w_dff_B_b8TbJFpE6_2;
	wire w_dff_B_7E5RzLfs3_2;
	wire w_dff_B_Gx4FnGt11_2;
	wire w_dff_B_hezCouQL0_2;
	wire w_dff_B_5UvB3LGI1_1;
	wire w_dff_B_mCXEI6MU7_2;
	wire w_dff_B_O0VDQWk33_2;
	wire w_dff_B_CzGRzmdV8_2;
	wire w_dff_B_Zy6iEuIS8_2;
	wire w_dff_B_Rzq0WHkh1_2;
	wire w_dff_B_3jIJbPnN8_2;
	wire w_dff_B_vSRM9jtN1_2;
	wire w_dff_B_C064Ldx37_2;
	wire w_dff_B_UqCfUbbl0_2;
	wire w_dff_B_4gNqZQ6U3_2;
	wire w_dff_B_a3Pynn9J5_2;
	wire w_dff_B_c7KDfeEO5_2;
	wire w_dff_B_gBzgjfyH6_2;
	wire w_dff_B_5SEIbU7t3_2;
	wire w_dff_B_415qIkVG1_2;
	wire w_dff_B_v3rUocvQ8_2;
	wire w_dff_B_3haXmg0g8_2;
	wire w_dff_B_KNCiGKZ97_2;
	wire w_dff_B_rf24kMxm6_2;
	wire w_dff_B_lNUudiTQ0_2;
	wire w_dff_B_2UpIYckQ7_2;
	wire w_dff_B_QQtLohz15_2;
	wire w_dff_B_aYNdfhs14_2;
	wire w_dff_B_L1fuHQAh4_2;
	wire w_dff_B_MTCZ4dim3_2;
	wire w_dff_B_qt7G1FVR1_2;
	wire w_dff_B_NP9hEVwk7_2;
	wire w_dff_B_U4zjTHIe6_2;
	wire w_dff_B_dYxUp4ZZ2_2;
	wire w_dff_B_ftWiGBnT3_2;
	wire w_dff_B_9hb6a1Uh9_2;
	wire w_dff_B_hgj8ijXl0_1;
	wire w_dff_B_SVC12NAg3_2;
	wire w_dff_B_T8Zumf2g3_2;
	wire w_dff_B_6qLkuQYL8_2;
	wire w_dff_B_fqbulSk57_2;
	wire w_dff_B_iDJaM1gZ3_2;
	wire w_dff_B_KGVodRJG6_2;
	wire w_dff_B_Ranb23lH1_2;
	wire w_dff_B_T7WTgaHo4_2;
	wire w_dff_B_NuDEaQ5W8_2;
	wire w_dff_B_USGlNJi82_2;
	wire w_dff_B_r1SfLcPh4_2;
	wire w_dff_B_rlHly6nH8_2;
	wire w_dff_B_E0ZwuUQ76_2;
	wire w_dff_B_Wd3YRfVH6_2;
	wire w_dff_B_USoAhaje4_2;
	wire w_dff_B_1A3IAvez5_2;
	wire w_dff_B_uwKaJnVk3_2;
	wire w_dff_B_52vhSuAy0_2;
	wire w_dff_B_MzU2Z5P66_2;
	wire w_dff_B_rFlLrsM89_2;
	wire w_dff_B_FoivV4FK2_2;
	wire w_dff_B_1lSY83kJ5_2;
	wire w_dff_B_U6pn8MCV0_2;
	wire w_dff_B_FRwaVpTt6_2;
	wire w_dff_B_YbsbpVBo5_2;
	wire w_dff_B_DogKVEKI8_2;
	wire w_dff_B_EvPQsQTx9_2;
	wire w_dff_B_lyf6aRnj3_2;
	wire w_dff_B_ejihLi905_1;
	wire w_dff_B_8tmlnGSw0_2;
	wire w_dff_B_jYs3cOUC2_2;
	wire w_dff_B_rnlV4XhB4_2;
	wire w_dff_B_5bgru6wk6_2;
	wire w_dff_B_5FJUSTER4_2;
	wire w_dff_B_TgHwNfGx5_2;
	wire w_dff_B_BIfroLRr4_2;
	wire w_dff_B_KLTNwEvz7_2;
	wire w_dff_B_A9JB9CBx1_2;
	wire w_dff_B_B79SkSOP5_2;
	wire w_dff_B_kVzTENRN5_2;
	wire w_dff_B_HOolG97J3_2;
	wire w_dff_B_ub6LlqDt7_2;
	wire w_dff_B_rXfaiVXV7_2;
	wire w_dff_B_OmLrzGUh4_2;
	wire w_dff_B_rVcu2sb88_2;
	wire w_dff_B_tiC8XncD4_2;
	wire w_dff_B_NFzBo2b02_2;
	wire w_dff_B_4oNoGlTu0_2;
	wire w_dff_B_zkskbeVv0_2;
	wire w_dff_B_DBALOCue2_2;
	wire w_dff_B_exPGFf5H8_2;
	wire w_dff_B_X27X6G9E4_2;
	wire w_dff_B_rVdzUtEe9_2;
	wire w_dff_B_kRNE0XN38_2;
	wire w_dff_B_bcO87PmO5_1;
	wire w_dff_B_15o0CNIv7_2;
	wire w_dff_B_xDZqN6vV3_2;
	wire w_dff_B_WxaKVyv42_2;
	wire w_dff_B_1oUppQOW7_2;
	wire w_dff_B_RTD3wpxT4_2;
	wire w_dff_B_O6tY3K6D3_2;
	wire w_dff_B_VIM8IrZv5_2;
	wire w_dff_B_zZP8cuCn5_2;
	wire w_dff_B_SggYFhFN6_2;
	wire w_dff_B_w3hIOeJM8_2;
	wire w_dff_B_bgnhEpoc2_2;
	wire w_dff_B_9aT2FqOb2_2;
	wire w_dff_B_XF7sNaeb1_2;
	wire w_dff_B_g8ZFeTXx7_2;
	wire w_dff_B_juyLj4hL1_2;
	wire w_dff_B_VoESLRuS1_2;
	wire w_dff_B_AqrnZTjL2_2;
	wire w_dff_B_RZYSF6Ie9_2;
	wire w_dff_B_zu2LB1KE1_2;
	wire w_dff_B_bwquSfY57_2;
	wire w_dff_B_sOd524Ka7_2;
	wire w_dff_B_aetrGM480_2;
	wire w_dff_B_URPxwRpp9_1;
	wire w_dff_B_JX1JPsH39_2;
	wire w_dff_B_LzIMJpeT5_2;
	wire w_dff_B_RHRCl1m07_2;
	wire w_dff_B_kVRLkMIe7_2;
	wire w_dff_B_JrghY2dp3_2;
	wire w_dff_B_VIqPRXn84_2;
	wire w_dff_B_86Mvjovt1_2;
	wire w_dff_B_tJqfScUJ3_2;
	wire w_dff_B_pHeX8w844_2;
	wire w_dff_B_gxYV5lXF4_2;
	wire w_dff_B_j4FeBo5q3_2;
	wire w_dff_B_A4h8XyKt2_2;
	wire w_dff_B_fxIZkuyq5_2;
	wire w_dff_B_OVMCcV4M9_2;
	wire w_dff_B_d4lPeMhm0_2;
	wire w_dff_B_gxhFJIEX7_2;
	wire w_dff_B_PfbytpzH3_2;
	wire w_dff_B_9p9WPMGU1_2;
	wire w_dff_B_36Zt8hAt2_2;
	wire w_dff_B_mt15VX7D5_1;
	wire w_dff_B_QDVq3hhf5_2;
	wire w_dff_B_laVjKb8a7_2;
	wire w_dff_B_13uV7ovM8_2;
	wire w_dff_B_TWvCCRVY6_2;
	wire w_dff_B_SV5xxY753_2;
	wire w_dff_B_5Vk9CDUZ0_2;
	wire w_dff_B_sqsRiXlB5_2;
	wire w_dff_B_HsnvKVp48_2;
	wire w_dff_B_m50m7EFJ1_2;
	wire w_dff_B_CLPglvEP6_2;
	wire w_dff_B_41jZgiFH2_2;
	wire w_dff_B_iWxlPfgi3_2;
	wire w_dff_B_VzJY0HY34_2;
	wire w_dff_B_BtmYRip35_2;
	wire w_dff_B_NiKik2ow3_2;
	wire w_dff_B_En3EkI4x6_2;
	wire w_dff_B_6mIyvaqr8_1;
	wire w_dff_B_ZkG2sCKQ3_2;
	wire w_dff_B_yz6FXYRl2_2;
	wire w_dff_B_PvE48pp64_2;
	wire w_dff_B_RzRloISO6_2;
	wire w_dff_B_DpzYwDeu2_2;
	wire w_dff_B_auSHm8h75_2;
	wire w_dff_B_UTZuA6aA1_2;
	wire w_dff_B_aLw4IxKS5_2;
	wire w_dff_B_a5EYDvMD5_2;
	wire w_dff_B_jCqgFF7T6_2;
	wire w_dff_B_bbkjXoID6_2;
	wire w_dff_B_B72SyqhR8_2;
	wire w_dff_B_7NIX7gzS4_2;
	wire w_dff_B_WEau1fSs0_1;
	wire w_dff_B_o8LENZfH4_2;
	wire w_dff_B_mYcDDcaN1_2;
	wire w_dff_B_3xPx2mjP2_2;
	wire w_dff_B_EU0XWfQ37_2;
	wire w_dff_B_1WI1LxuM9_2;
	wire w_dff_B_Mq67UBh45_2;
	wire w_dff_B_GkKC40wH3_2;
	wire w_dff_B_Vd9qOpJS2_2;
	wire w_dff_B_1I7m3Dei3_2;
	wire w_dff_B_21WflzzA2_2;
	wire w_dff_B_hGv4qMwx9_2;
	wire w_dff_B_BRvDgPUz5_1;
	wire w_dff_B_gkTAIXDB4_2;
	wire w_dff_B_5AEfshf03_2;
	wire w_dff_B_sn5xgl242_2;
	wire w_dff_B_StLJC8py1_2;
	wire w_dff_B_3aGprczc4_2;
	wire w_dff_B_BuSQx6z12_2;
	wire w_dff_B_6rTgYPtY9_2;
	wire w_dff_B_VPsceqs67_2;
	wire w_dff_B_zXRprNEB1_1;
	wire w_dff_B_pfL42Ayq3_2;
	wire w_dff_B_qx0OKX9I8_2;
	wire w_dff_B_DPBQgWQQ8_2;
	wire w_dff_B_u3Vi490M7_2;
	wire w_dff_B_9hPIJqTT8_1;
	wire w_dff_A_mTvMtSiG7_1;
	wire w_dff_A_9AFadnxN6_2;
	wire w_dff_A_Y3Yw9DWj9_2;
	wire w_dff_B_af4nwA5n9_2;
	wire w_dff_B_lyPa9dUU4_1;
	wire w_dff_B_b91cSgik3_2;
	wire w_dff_B_oSg7x4ko5_2;
	wire w_dff_B_qjZqg0KE8_2;
	wire w_dff_B_u7AMRP7r4_2;
	wire w_dff_B_FCrRxCp12_2;
	wire w_dff_B_e9lWhaMh6_2;
	wire w_dff_B_2Jin6f3F3_2;
	wire w_dff_B_8JFB5qkn8_2;
	wire w_dff_B_0EMXC8208_2;
	wire w_dff_B_NuzJ0KOO9_2;
	wire w_dff_B_u46PCaA40_2;
	wire w_dff_B_0ErCbtZ50_2;
	wire w_dff_B_uM9twtl81_2;
	wire w_dff_B_3LU7KrCG1_2;
	wire w_dff_B_Ql0WrQ9X9_2;
	wire w_dff_B_RkAULWx05_2;
	wire w_dff_B_6vocVvua1_2;
	wire w_dff_B_tW9KBL286_2;
	wire w_dff_B_ZyUpNRHt8_2;
	wire w_dff_B_biC251xL4_2;
	wire w_dff_B_e92ZTNfs3_2;
	wire w_dff_B_bNC18lju6_2;
	wire w_dff_B_cRmE4bC50_2;
	wire w_dff_B_lfOlE06q1_2;
	wire w_dff_B_eoX6Bakl1_2;
	wire w_dff_B_9TVjwXdf9_2;
	wire w_dff_B_YTqThHKS5_2;
	wire w_dff_B_xlThTkhQ4_2;
	wire w_dff_B_Nx0zpbCt3_2;
	wire w_dff_B_bij20Ba39_2;
	wire w_dff_B_C8CaNbL76_2;
	wire w_dff_B_N5WoFur92_2;
	wire w_dff_B_mZ5Xmqrh6_2;
	wire w_dff_B_0Ag6xAvX4_2;
	wire w_dff_B_U0zwXmFV7_2;
	wire w_dff_B_CuCPYtPz5_2;
	wire w_dff_B_pxy1iGAq9_2;
	wire w_dff_B_jR0iFg8K1_2;
	wire w_dff_B_1J0Cuqgg8_2;
	wire w_dff_B_apvSUipR6_2;
	wire w_dff_B_q7suo3Om0_2;
	wire w_dff_B_So1lJT9J4_2;
	wire w_dff_B_UMZT43dn0_2;
	wire w_dff_B_KtAuF9hr8_2;
	wire w_dff_B_yHuuOPrg8_2;
	wire w_dff_B_mHXheFJ27_2;
	wire w_dff_B_0sLmQqVT3_1;
	wire w_dff_B_5tJmI57P5_2;
	wire w_dff_B_9QME0q2B4_2;
	wire w_dff_B_7xhXWA223_2;
	wire w_dff_B_dJOUgNBE3_2;
	wire w_dff_B_TwqBUNJx6_2;
	wire w_dff_B_OT7Snrp47_2;
	wire w_dff_B_pDi4Wbia3_2;
	wire w_dff_B_AUAjYsRO8_2;
	wire w_dff_B_2HlyQ3Bq3_2;
	wire w_dff_B_QDoAMHQW1_2;
	wire w_dff_B_kNc6j2k42_2;
	wire w_dff_B_S9UkJYeo5_2;
	wire w_dff_B_ullc4rfi4_2;
	wire w_dff_B_IQtjO9Gk3_2;
	wire w_dff_B_wMJgVePA9_2;
	wire w_dff_B_z3dhxdxZ4_2;
	wire w_dff_B_h61JaaDv8_2;
	wire w_dff_B_2UEESRfr9_2;
	wire w_dff_B_tyLtbAUh7_2;
	wire w_dff_B_ign3mPvn2_2;
	wire w_dff_B_BKmplsR23_2;
	wire w_dff_B_ACE7mfZj3_2;
	wire w_dff_B_7ilA3YS45_2;
	wire w_dff_B_w5rh1REM0_2;
	wire w_dff_B_k3j7mOcY8_2;
	wire w_dff_B_z5EWQJTw5_2;
	wire w_dff_B_FXUl9Wqj3_2;
	wire w_dff_B_lt5yDCXU4_2;
	wire w_dff_B_VAv23shb7_2;
	wire w_dff_B_iHuUAZne0_2;
	wire w_dff_B_gHdQwUYq2_2;
	wire w_dff_B_nQBWvc5R7_2;
	wire w_dff_B_10SL5MYS1_2;
	wire w_dff_B_LWPKLSUN0_2;
	wire w_dff_B_OOad25P37_2;
	wire w_dff_B_RZEtVhtQ4_2;
	wire w_dff_B_Ayb7RcQF5_2;
	wire w_dff_B_GiRCWBgL6_2;
	wire w_dff_B_GFOoJ2eq1_2;
	wire w_dff_B_8QCyBW503_2;
	wire w_dff_B_y92mo1M43_2;
	wire w_dff_B_bDocydhb6_1;
	wire w_dff_B_Ail7x0LW9_2;
	wire w_dff_B_xavbA5MR9_2;
	wire w_dff_B_vHrddRzb8_2;
	wire w_dff_B_NJui82fM2_2;
	wire w_dff_B_RskdySKq1_2;
	wire w_dff_B_hw3E776r6_2;
	wire w_dff_B_XIN9RZpx1_2;
	wire w_dff_B_d4Zgy1eJ0_2;
	wire w_dff_B_0NtEvgCP8_2;
	wire w_dff_B_RlnOtElS8_2;
	wire w_dff_B_IfUQm2lL0_2;
	wire w_dff_B_i5zHiUAi2_2;
	wire w_dff_B_KkSADCCF8_2;
	wire w_dff_B_8g0Ewo7V6_2;
	wire w_dff_B_HSIJxpFC1_2;
	wire w_dff_B_DAgV7bOd7_2;
	wire w_dff_B_dsajmSpj9_2;
	wire w_dff_B_Pk4fXni59_2;
	wire w_dff_B_OVThfzDU0_2;
	wire w_dff_B_zWenA68s5_2;
	wire w_dff_B_Eu3jSEHU6_2;
	wire w_dff_B_RVVbgxur4_2;
	wire w_dff_B_DuuBdalP3_2;
	wire w_dff_B_REGAyUM73_2;
	wire w_dff_B_a2ns7YfN0_2;
	wire w_dff_B_3fS8brj32_2;
	wire w_dff_B_Hgfq9Fns9_2;
	wire w_dff_B_IOp36Eyd7_2;
	wire w_dff_B_McR7QJ8w7_2;
	wire w_dff_B_xciPzj6d2_2;
	wire w_dff_B_HCGnocdg4_2;
	wire w_dff_B_85Xw2VgO6_2;
	wire w_dff_B_5voB3PvG2_2;
	wire w_dff_B_mWk1ScFL8_2;
	wire w_dff_B_Pg428fCG4_2;
	wire w_dff_B_shBRayP63_2;
	wire w_dff_B_OTJVvwQm7_2;
	wire w_dff_B_jqkbv9TZ6_2;
	wire w_dff_B_zK7yrA7e2_1;
	wire w_dff_B_7uyajVL02_2;
	wire w_dff_B_aJI8Ek0i5_2;
	wire w_dff_B_mlSvc89j3_2;
	wire w_dff_B_casXwag60_2;
	wire w_dff_B_gtm8WN0E9_2;
	wire w_dff_B_8MCiHWbo3_2;
	wire w_dff_B_cYymuwiC9_2;
	wire w_dff_B_9iBaMvuu7_2;
	wire w_dff_B_PFTMqEUl0_2;
	wire w_dff_B_M8nr22Pk2_2;
	wire w_dff_B_D8TWBapD3_2;
	wire w_dff_B_pbZqulTo2_2;
	wire w_dff_B_wMTcAZ8Y7_2;
	wire w_dff_B_4tgce4Oe3_2;
	wire w_dff_B_B0kY7cIH1_2;
	wire w_dff_B_c076dEod8_2;
	wire w_dff_B_5AyQ7Kps5_2;
	wire w_dff_B_zCdsglMz7_2;
	wire w_dff_B_7sk5J8Lk6_2;
	wire w_dff_B_3QNWTExY5_2;
	wire w_dff_B_CfXARsHa5_2;
	wire w_dff_B_UQzIMyu93_2;
	wire w_dff_B_I1spHyv23_2;
	wire w_dff_B_iWjL12xB1_2;
	wire w_dff_B_neoiNxse3_2;
	wire w_dff_B_8FspEcO81_2;
	wire w_dff_B_8f7XQWKB3_2;
	wire w_dff_B_lALwfbKI4_2;
	wire w_dff_B_m9RP6cwh6_2;
	wire w_dff_B_SSSYWT8j9_2;
	wire w_dff_B_7VQRIbGZ3_2;
	wire w_dff_B_V6QtCvTC6_2;
	wire w_dff_B_WtOJPJKQ0_2;
	wire w_dff_B_EDZ0dM3p1_2;
	wire w_dff_B_E2OoLQUy0_2;
	wire w_dff_B_XCy6AqqE0_1;
	wire w_dff_B_mOhtwAco6_2;
	wire w_dff_B_x0ipWgB22_2;
	wire w_dff_B_zf7ubohQ5_2;
	wire w_dff_B_PeLc1mhz9_2;
	wire w_dff_B_whT14DNR7_2;
	wire w_dff_B_HWEOoNUW5_2;
	wire w_dff_B_VvaK21gh7_2;
	wire w_dff_B_f7Ewsdfj0_2;
	wire w_dff_B_Uw2GXW670_2;
	wire w_dff_B_JoyZDAp41_2;
	wire w_dff_B_OKEVUuN66_2;
	wire w_dff_B_s2pdcjXa7_2;
	wire w_dff_B_jPZTSIGX5_2;
	wire w_dff_B_sKgUjKXE1_2;
	wire w_dff_B_9PaQxmQP1_2;
	wire w_dff_B_ywhxro8M9_2;
	wire w_dff_B_LptVu05a3_2;
	wire w_dff_B_IuiQWMej4_2;
	wire w_dff_B_fNhIjUJw6_2;
	wire w_dff_B_OSaYeidp7_2;
	wire w_dff_B_6Jqctgxu6_2;
	wire w_dff_B_6vbSIVrz5_2;
	wire w_dff_B_hc25mcsi0_2;
	wire w_dff_B_BHvM9pOO0_2;
	wire w_dff_B_vZjccCfE4_2;
	wire w_dff_B_KO3LgFCP8_2;
	wire w_dff_B_K2se7K8b0_2;
	wire w_dff_B_33bsCwZD8_2;
	wire w_dff_B_LPZAWkT82_2;
	wire w_dff_B_rdNKtdbr7_2;
	wire w_dff_B_bzUD0DS71_2;
	wire w_dff_B_NrD0JuhJ0_2;
	wire w_dff_B_oBxkf0G21_1;
	wire w_dff_B_nyQzncQx5_2;
	wire w_dff_B_hENfEriK5_2;
	wire w_dff_B_uC9fZBbf0_2;
	wire w_dff_B_95qiEZUQ9_2;
	wire w_dff_B_Q0983WCM7_2;
	wire w_dff_B_t5DBuE1C2_2;
	wire w_dff_B_xPq4QyHT7_2;
	wire w_dff_B_QnUdnQ4N2_2;
	wire w_dff_B_DeNrO5LU5_2;
	wire w_dff_B_lzcae39c3_2;
	wire w_dff_B_jjAg2ibS9_2;
	wire w_dff_B_HfQroRc54_2;
	wire w_dff_B_UnysazIq1_2;
	wire w_dff_B_B2BlSJOF6_2;
	wire w_dff_B_2ifCDld99_2;
	wire w_dff_B_KbyW8fFN2_2;
	wire w_dff_B_MPuTgbVK7_2;
	wire w_dff_B_tWotBzHZ0_2;
	wire w_dff_B_KeyjJanE4_2;
	wire w_dff_B_zWDtDGxn6_2;
	wire w_dff_B_DS3KBvOr0_2;
	wire w_dff_B_CG1L7VNh1_2;
	wire w_dff_B_zhuitS4c0_2;
	wire w_dff_B_V8xvLMEC0_2;
	wire w_dff_B_1mwnz31j4_2;
	wire w_dff_B_o8JfBlew1_2;
	wire w_dff_B_NnywUvYP6_2;
	wire w_dff_B_AJzwcfb63_2;
	wire w_dff_B_JKhRRn0h9_2;
	wire w_dff_B_E28e5hOE1_1;
	wire w_dff_B_XOMImEQL4_2;
	wire w_dff_B_qGKIcVa97_2;
	wire w_dff_B_HqFOYD4u0_2;
	wire w_dff_B_lcSgrEP82_2;
	wire w_dff_B_AljT9tO11_2;
	wire w_dff_B_FruXNmDq8_2;
	wire w_dff_B_3603w8rk5_2;
	wire w_dff_B_OFuueyCD7_2;
	wire w_dff_B_Oi6COfNE5_2;
	wire w_dff_B_Ku37XT687_2;
	wire w_dff_B_5IOc2Odm5_2;
	wire w_dff_B_KSCjAnzz0_2;
	wire w_dff_B_k0txzxyL3_2;
	wire w_dff_B_P8ezx6NU1_2;
	wire w_dff_B_SaaKk0rA0_2;
	wire w_dff_B_B717Sm6c3_2;
	wire w_dff_B_m7ZYFU6e0_2;
	wire w_dff_B_uAifJrff4_2;
	wire w_dff_B_SGZ4B0SC9_2;
	wire w_dff_B_Yl81yMHH5_2;
	wire w_dff_B_pB7p2nKL1_2;
	wire w_dff_B_KtKs2P754_2;
	wire w_dff_B_Bdt25Oma6_2;
	wire w_dff_B_liaGK4Oh9_2;
	wire w_dff_B_753rPRre9_2;
	wire w_dff_B_OIsxnejw5_2;
	wire w_dff_B_BjPK4aKx5_1;
	wire w_dff_B_DMqxYSwQ6_2;
	wire w_dff_B_Z2s64YQC9_2;
	wire w_dff_B_cuSyWlnS8_2;
	wire w_dff_B_Nbzw6ON34_2;
	wire w_dff_B_HH89iHAK3_2;
	wire w_dff_B_C6LyLxPP1_2;
	wire w_dff_B_hcv6tpdE9_2;
	wire w_dff_B_0szlR8g17_2;
	wire w_dff_B_ArXzfoTA0_2;
	wire w_dff_B_1B7dMboQ7_2;
	wire w_dff_B_a5FZGSEl5_2;
	wire w_dff_B_0Yhipu7D7_2;
	wire w_dff_B_1NUpT4y28_2;
	wire w_dff_B_8xQEpUDT5_2;
	wire w_dff_B_P6n3vYq81_2;
	wire w_dff_B_p5tsQIBi6_2;
	wire w_dff_B_LuONwujo3_2;
	wire w_dff_B_kvuIYBN82_2;
	wire w_dff_B_B1AggMv63_2;
	wire w_dff_B_6AdCB4FG6_2;
	wire w_dff_B_LLHzkkIu4_2;
	wire w_dff_B_xGKzri6L1_2;
	wire w_dff_B_ZHXhiKye4_2;
	wire w_dff_B_OItvkCtj8_1;
	wire w_dff_B_9iip8WQh6_2;
	wire w_dff_B_UZ6QsmhZ9_2;
	wire w_dff_B_CN2r3IKi5_2;
	wire w_dff_B_55AyiywL1_2;
	wire w_dff_B_sR5FerlT7_2;
	wire w_dff_B_8geRG4Xy3_2;
	wire w_dff_B_DePmAgkt6_2;
	wire w_dff_B_iU6G1aGu4_2;
	wire w_dff_B_FqTiiNcf0_2;
	wire w_dff_B_QEpK86Ut0_2;
	wire w_dff_B_T56r6L5y9_2;
	wire w_dff_B_P48ZY4Fs4_2;
	wire w_dff_B_Bjh8NZoH4_2;
	wire w_dff_B_BUMgbZW81_2;
	wire w_dff_B_Czt1wo8U3_2;
	wire w_dff_B_YvoKr5Zw3_2;
	wire w_dff_B_LcymxrAF2_2;
	wire w_dff_B_jrHV2jSQ8_2;
	wire w_dff_B_CPoqtNDM3_2;
	wire w_dff_B_gvaO9FrA4_2;
	wire w_dff_B_wUqJfUUX3_1;
	wire w_dff_B_kFLC2GR77_2;
	wire w_dff_B_TIqJxy468_2;
	wire w_dff_B_68EIUyMI6_2;
	wire w_dff_B_d73FkaNb1_2;
	wire w_dff_B_rswHVzdp1_2;
	wire w_dff_B_yGhtyHuM2_2;
	wire w_dff_B_H36rjuGp4_2;
	wire w_dff_B_NPyD8V6Q4_2;
	wire w_dff_B_kkvFLeXN6_2;
	wire w_dff_B_MOs6bbNg7_2;
	wire w_dff_B_XgJLOM088_2;
	wire w_dff_B_Jqb2q0UQ9_2;
	wire w_dff_B_23u9yKB51_2;
	wire w_dff_B_vFV6DZay9_2;
	wire w_dff_B_ljWA7UnI5_2;
	wire w_dff_B_oIEOGCbR3_2;
	wire w_dff_B_FnvGQ8Bn4_2;
	wire w_dff_B_fglGzeOF8_1;
	wire w_dff_B_GmEdFwzt9_2;
	wire w_dff_B_Wet41jYg8_2;
	wire w_dff_B_0IM08Xhr6_2;
	wire w_dff_B_Nm7ohPpE8_2;
	wire w_dff_B_799TdZwW8_2;
	wire w_dff_B_RCFvNIZR1_2;
	wire w_dff_B_FSi5VrUN6_2;
	wire w_dff_B_QZz8XZda1_2;
	wire w_dff_B_WZuxoPR85_2;
	wire w_dff_B_PXzCCsIk5_2;
	wire w_dff_B_IaG5tIM03_2;
	wire w_dff_B_EZJV2KLH4_2;
	wire w_dff_B_g1cfKTTf9_2;
	wire w_dff_B_teV2fcSQ9_2;
	wire w_dff_B_Vf2dWUQs7_1;
	wire w_dff_B_cMyEysnW7_2;
	wire w_dff_B_ZS1GBwxJ1_2;
	wire w_dff_B_z8q1Xxtq9_2;
	wire w_dff_B_88FlmuEy4_2;
	wire w_dff_B_C0jFK4sV5_2;
	wire w_dff_B_A58XZpTV7_2;
	wire w_dff_B_kPCrZGqh9_2;
	wire w_dff_B_9eO8g0EC0_2;
	wire w_dff_B_Bb2lQgUJ4_2;
	wire w_dff_B_xj0jtopr1_2;
	wire w_dff_B_mcltNOjw8_2;
	wire w_dff_B_qWfI2QVG8_2;
	wire w_dff_B_Q5Fcfau46_1;
	wire w_dff_B_U2vHbwWV2_2;
	wire w_dff_B_4MUSLB1k8_2;
	wire w_dff_B_cJrien2v6_2;
	wire w_dff_B_yGpplbgN8_2;
	wire w_dff_B_oeqtDQfZ4_2;
	wire w_dff_B_P2HwkiEj0_2;
	wire w_dff_B_BeecgaRi2_2;
	wire w_dff_B_frfc0sZl2_1;
	wire w_dff_B_kEXGgwSC7_2;
	wire w_dff_B_u817jq6I1_2;
	wire w_dff_B_hT7sTadY8_2;
	wire w_dff_B_Vr0RTiuP0_2;
	wire w_dff_B_oBTVm2AH7_1;
	wire w_dff_A_AvuFHgdL3_0;
	wire w_dff_A_7C2puQDr9_1;
	wire w_dff_A_jWxdfK7Z8_1;
	wire w_dff_B_a7Ek4TkY8_1;
	wire w_dff_B_6OiQ7KOP5_2;
	wire w_dff_B_VAkpoyWb1_2;
	wire w_dff_B_JxIrZkrD4_2;
	wire w_dff_B_iQLfoj5c4_2;
	wire w_dff_B_YxIZrGR83_2;
	wire w_dff_B_o6gtRhGj2_2;
	wire w_dff_B_TW9KYJLO6_2;
	wire w_dff_B_k6VH2Q193_2;
	wire w_dff_B_25UzyUww6_2;
	wire w_dff_B_6km1JTS97_2;
	wire w_dff_B_VKnZfUOf9_2;
	wire w_dff_B_38KD7hC70_2;
	wire w_dff_B_b8etlaOw9_2;
	wire w_dff_B_hjrHoEkS4_2;
	wire w_dff_B_kEykrjUL0_2;
	wire w_dff_B_vq3QEiX60_2;
	wire w_dff_B_EnuqSSC76_2;
	wire w_dff_B_RyGsuda15_2;
	wire w_dff_B_gXBYITOv9_2;
	wire w_dff_B_s8ONbQNv6_2;
	wire w_dff_B_wGlfMzgV9_2;
	wire w_dff_B_zYRG2Gs04_2;
	wire w_dff_B_c91Sn8wm0_2;
	wire w_dff_B_eus8bNGi7_2;
	wire w_dff_B_w9D4qMMB1_2;
	wire w_dff_B_AxNKrLfK5_2;
	wire w_dff_B_j7ItMyId4_2;
	wire w_dff_B_fiq6Y3Uz5_2;
	wire w_dff_B_Ehj2jM1H8_2;
	wire w_dff_B_XxuADOnt9_2;
	wire w_dff_B_suFlq2yO6_2;
	wire w_dff_B_9XRI0iW76_2;
	wire w_dff_B_DYWbz1V77_2;
	wire w_dff_B_t2OAjFSP9_2;
	wire w_dff_B_rQhOI8dt1_2;
	wire w_dff_B_aXoHWW1L3_2;
	wire w_dff_B_bb8YBTnX9_2;
	wire w_dff_B_V0we07Ct8_2;
	wire w_dff_B_4J5hfqI36_2;
	wire w_dff_B_gjALG9Sg6_2;
	wire w_dff_B_vcd18Xy44_2;
	wire w_dff_B_MaBGK2ZJ6_2;
	wire w_dff_B_rdBsrFSB6_2;
	wire w_dff_B_fOTeTZGn3_2;
	wire w_dff_B_CglMBADb8_2;
	wire w_dff_B_tJOgbhkn2_2;
	wire w_dff_B_tUghYg4N8_2;
	wire w_dff_B_s9pv34mm5_0;
	wire w_dff_A_F5DGNIku5_1;
	wire w_dff_B_e2bwT7h06_1;
	wire w_dff_B_CRk1sifL2_2;
	wire w_dff_B_Ju8zlzNq1_2;
	wire w_dff_B_BY1FXfIO0_2;
	wire w_dff_B_WfLnq02U3_2;
	wire w_dff_B_ksq5eyME8_2;
	wire w_dff_B_l6MKBJQM9_2;
	wire w_dff_B_930jjDuG8_2;
	wire w_dff_B_EsZfHCgp1_2;
	wire w_dff_B_JnaD8V9o0_2;
	wire w_dff_B_BjsTLkAz3_2;
	wire w_dff_B_RL6P5p603_2;
	wire w_dff_B_hIKrwDcf8_2;
	wire w_dff_B_ogz0763N5_2;
	wire w_dff_B_PfZnDpBT2_2;
	wire w_dff_B_tnuc2eg79_2;
	wire w_dff_B_7k1bm7ej2_2;
	wire w_dff_B_zvaQSFfi3_2;
	wire w_dff_B_cLNwiovw4_2;
	wire w_dff_B_8wOJKZMX3_2;
	wire w_dff_B_SLA6GgvG4_2;
	wire w_dff_B_amgcxnxY8_2;
	wire w_dff_B_v4Dq6eWx9_2;
	wire w_dff_B_yNxQI4gv3_2;
	wire w_dff_B_FGIvQC5V9_2;
	wire w_dff_B_FndKnCOF7_2;
	wire w_dff_B_wIsyC8f90_2;
	wire w_dff_B_OuhIXG5k1_2;
	wire w_dff_B_fM5tUCeI0_2;
	wire w_dff_B_cwCqhBH69_2;
	wire w_dff_B_Pw1ZbvxO1_2;
	wire w_dff_B_JyhtQZQO0_2;
	wire w_dff_B_5Dh4twdb5_2;
	wire w_dff_B_UfOpPLRJ1_2;
	wire w_dff_B_g28XbUXD3_2;
	wire w_dff_B_zYdXWDBQ3_2;
	wire w_dff_B_uSFFYiaJ4_2;
	wire w_dff_B_j8gS4rYn5_2;
	wire w_dff_B_cpus0BYS8_2;
	wire w_dff_B_DnWkXHHD1_2;
	wire w_dff_B_0UOEMpfM8_2;
	wire w_dff_B_HVbczsyo8_2;
	wire w_dff_B_EZtOMoZi1_2;
	wire w_dff_B_tAhCEUVg1_2;
	wire w_dff_B_ZSPAhZlk1_1;
	wire w_dff_B_BBihBqEI5_2;
	wire w_dff_B_jDDh1dZe2_2;
	wire w_dff_B_GgoR3HXw2_2;
	wire w_dff_B_HiHWYSxc4_2;
	wire w_dff_B_v3TXDpmH7_2;
	wire w_dff_B_9oJoUrMx1_2;
	wire w_dff_B_ISiofFKw6_2;
	wire w_dff_B_xRZfEihv5_2;
	wire w_dff_B_hIyYMjOF2_2;
	wire w_dff_B_X6nD6tSp8_2;
	wire w_dff_B_WKhHgbCe4_2;
	wire w_dff_B_kQ7EQnuO3_2;
	wire w_dff_B_5zgnJw3n2_2;
	wire w_dff_B_wHnUWgf08_2;
	wire w_dff_B_VekJkxUo3_2;
	wire w_dff_B_DBhouzLf2_2;
	wire w_dff_B_Zfm53BT94_2;
	wire w_dff_B_IBqI79TY6_2;
	wire w_dff_B_68jk4Xgo4_2;
	wire w_dff_B_sTWsASjY0_2;
	wire w_dff_B_aGyb8gCw7_2;
	wire w_dff_B_QVHn0I109_2;
	wire w_dff_B_79NxnVDp1_2;
	wire w_dff_B_s7opvF8h8_2;
	wire w_dff_B_t78o9VrW6_2;
	wire w_dff_B_YrlfMDkA7_2;
	wire w_dff_B_3PDqQoUz8_2;
	wire w_dff_B_6rpQnCHN7_2;
	wire w_dff_B_2JdcIaBd0_2;
	wire w_dff_B_eKtQYpni8_2;
	wire w_dff_B_cIpnUKxG6_2;
	wire w_dff_B_2EQaBGhu3_2;
	wire w_dff_B_TG6jqPYo9_2;
	wire w_dff_B_JIKEOoQC7_2;
	wire w_dff_B_dGFEP0HU9_2;
	wire w_dff_B_moFxXqUc3_2;
	wire w_dff_B_zrGK7h9Q9_2;
	wire w_dff_B_yajQF2IL8_2;
	wire w_dff_B_1mUiIhGD0_2;
	wire w_dff_B_h43tcy7G1_2;
	wire w_dff_B_wy76JoGg3_1;
	wire w_dff_B_NeX1hRvQ1_2;
	wire w_dff_B_RWBEAAdS1_2;
	wire w_dff_B_RVTA9aVm7_2;
	wire w_dff_B_zf0beyWt6_2;
	wire w_dff_B_ACwv2XYC1_2;
	wire w_dff_B_ueVYOmkw0_2;
	wire w_dff_B_LgATYXHV8_2;
	wire w_dff_B_uwK8qIgI7_2;
	wire w_dff_B_u0jfZRod8_2;
	wire w_dff_B_EHBcFeNq6_2;
	wire w_dff_B_OJxLDOx33_2;
	wire w_dff_B_rewFnKMG4_2;
	wire w_dff_B_4lNU28JW5_2;
	wire w_dff_B_8mQQWD5G9_2;
	wire w_dff_B_ShnYhHWD6_2;
	wire w_dff_B_xlD0g9lO1_2;
	wire w_dff_B_fF2yctoZ7_2;
	wire w_dff_B_Y1wkKzun8_2;
	wire w_dff_B_dNSLuPXO6_2;
	wire w_dff_B_G8qqZ5KO9_2;
	wire w_dff_B_OERPKPWq2_2;
	wire w_dff_B_Dueiev5m7_2;
	wire w_dff_B_G9m2nPnM6_2;
	wire w_dff_B_P8kuslus2_2;
	wire w_dff_B_Lj7OmQTa2_2;
	wire w_dff_B_DZv6EsN07_2;
	wire w_dff_B_08JtWV9c9_2;
	wire w_dff_B_4FmvezaM7_2;
	wire w_dff_B_ttAipD6f0_2;
	wire w_dff_B_c6VXBlo29_2;
	wire w_dff_B_sSyisVPl4_2;
	wire w_dff_B_XZx3L21p3_2;
	wire w_dff_B_BirgbWRu8_2;
	wire w_dff_B_HGNURKlE3_2;
	wire w_dff_B_7HTfMSpd3_2;
	wire w_dff_B_xJ4lo3gy1_2;
	wire w_dff_B_j4ccORpw4_2;
	wire w_dff_B_pso4BWIG7_1;
	wire w_dff_B_1358zHiR8_2;
	wire w_dff_B_CYXUL9BU8_2;
	wire w_dff_B_ZSNxD25b5_2;
	wire w_dff_B_AYe82MC54_2;
	wire w_dff_B_UQRwkBIb4_2;
	wire w_dff_B_AdAe421E2_2;
	wire w_dff_B_6asGMBeO7_2;
	wire w_dff_B_nKGYjs7M3_2;
	wire w_dff_B_uPiQvcUB2_2;
	wire w_dff_B_MWdC6FJw8_2;
	wire w_dff_B_4OLM8gYH6_2;
	wire w_dff_B_YGzHT0Ke1_2;
	wire w_dff_B_vcWwLAXK1_2;
	wire w_dff_B_fzaBfLtr1_2;
	wire w_dff_B_MfQrkHRc2_2;
	wire w_dff_B_silPUtMO9_2;
	wire w_dff_B_S0Z2uyZL2_2;
	wire w_dff_B_8yEk5SvW4_2;
	wire w_dff_B_pEDkgknt9_2;
	wire w_dff_B_OTlGUdHG2_2;
	wire w_dff_B_uofPgif12_2;
	wire w_dff_B_ChPGCqtO6_2;
	wire w_dff_B_zcb7UaWP0_2;
	wire w_dff_B_GYbfLOCB6_2;
	wire w_dff_B_mqJNDizi8_2;
	wire w_dff_B_YGE03wAb8_2;
	wire w_dff_B_Q292y9IC7_2;
	wire w_dff_B_WCye4B1L3_2;
	wire w_dff_B_B58ROhoa7_2;
	wire w_dff_B_MAo13koB8_2;
	wire w_dff_B_Vcwkr3mJ5_2;
	wire w_dff_B_jX9rnMVy8_2;
	wire w_dff_B_j1oyz5BA5_2;
	wire w_dff_B_9lJINcr55_2;
	wire w_dff_B_G4BLumyx3_1;
	wire w_dff_B_Q3jPNhJv6_2;
	wire w_dff_B_wbRrDhLM7_2;
	wire w_dff_B_ZUZcUyXr0_2;
	wire w_dff_B_gIIwQgTX3_2;
	wire w_dff_B_xuS6p7uN6_2;
	wire w_dff_B_0iImqIBf5_2;
	wire w_dff_B_vbz6hfqB8_2;
	wire w_dff_B_qnixko3u2_2;
	wire w_dff_B_FTMFh1rF0_2;
	wire w_dff_B_AU68H9Ma6_2;
	wire w_dff_B_PXvKcBjt5_2;
	wire w_dff_B_KAXABrBD4_2;
	wire w_dff_B_gdYoejx88_2;
	wire w_dff_B_sVMqajT57_2;
	wire w_dff_B_wsJfr5GO5_2;
	wire w_dff_B_9QDL4fAG9_2;
	wire w_dff_B_kl0hNwtY1_2;
	wire w_dff_B_Moe8oQkM1_2;
	wire w_dff_B_Z0tkFoNr0_2;
	wire w_dff_B_VGf10PbV4_2;
	wire w_dff_B_rQQEUbGa5_2;
	wire w_dff_B_i4zFlsOZ1_2;
	wire w_dff_B_UnitFUWO0_2;
	wire w_dff_B_xkZ4nLUA8_2;
	wire w_dff_B_Lgee2QSR6_2;
	wire w_dff_B_yO2qVK7s6_2;
	wire w_dff_B_2NTOnvvt3_2;
	wire w_dff_B_doNzjmTP1_2;
	wire w_dff_B_Dgg0nkJt3_2;
	wire w_dff_B_GJjsYhnp3_2;
	wire w_dff_B_kDDcdUhh8_2;
	wire w_dff_B_Te2DMkeV2_1;
	wire w_dff_B_Jsa86ADT8_2;
	wire w_dff_B_WL9chbz29_2;
	wire w_dff_B_ULj5iaHx7_2;
	wire w_dff_B_DHBfNhz54_2;
	wire w_dff_B_2qGWFMQl2_2;
	wire w_dff_B_aQGaA4Za0_2;
	wire w_dff_B_mjHKD8rN8_2;
	wire w_dff_B_oBXeoxYE2_2;
	wire w_dff_B_UlvHVh8l3_2;
	wire w_dff_B_yrL2DVxN3_2;
	wire w_dff_B_NkKw86oq4_2;
	wire w_dff_B_14l0rrfd8_2;
	wire w_dff_B_kXV8kFB23_2;
	wire w_dff_B_kSCqlgoC6_2;
	wire w_dff_B_3iU9ar9N8_2;
	wire w_dff_B_Gw5pAFzS1_2;
	wire w_dff_B_rVHpWqyr2_2;
	wire w_dff_B_qrzvK4L54_2;
	wire w_dff_B_kM7teKYt7_2;
	wire w_dff_B_ES7MMwfb4_2;
	wire w_dff_B_yhxDzAL87_2;
	wire w_dff_B_6vJfkKJo8_2;
	wire w_dff_B_coBziEtT1_2;
	wire w_dff_B_9Hzk6QpC5_2;
	wire w_dff_B_owkWELKf1_2;
	wire w_dff_B_WJPbcDJ61_2;
	wire w_dff_B_0GgBGg4k2_2;
	wire w_dff_B_zSTRPc7K1_2;
	wire w_dff_B_EmgwCGB41_1;
	wire w_dff_B_3nxafNs61_2;
	wire w_dff_B_UVOgzU6u1_2;
	wire w_dff_B_GUrKVJXz2_2;
	wire w_dff_B_NJZcMozq2_2;
	wire w_dff_B_NDV9Pm8I8_2;
	wire w_dff_B_o2j6B1N85_2;
	wire w_dff_B_vH3utIIh2_2;
	wire w_dff_B_wCKZoReK9_2;
	wire w_dff_B_UCXrvMmd6_2;
	wire w_dff_B_ohqaDXTR8_2;
	wire w_dff_B_LdsytaWj7_2;
	wire w_dff_B_0fx8rzbe7_2;
	wire w_dff_B_6b4szKvX3_2;
	wire w_dff_B_rUdwhUp44_2;
	wire w_dff_B_W7VYc7rs4_2;
	wire w_dff_B_HGTTSMio6_2;
	wire w_dff_B_aeVR1pgf9_2;
	wire w_dff_B_GcMdokl36_2;
	wire w_dff_B_4LTIuvhI7_2;
	wire w_dff_B_bk8ANp4Q0_2;
	wire w_dff_B_VkVesc1V1_2;
	wire w_dff_B_CCcb015G0_2;
	wire w_dff_B_gPYa9o3J8_2;
	wire w_dff_B_krEo57156_2;
	wire w_dff_B_KJRKARdL5_2;
	wire w_dff_B_PslMiuzK5_1;
	wire w_dff_B_3wzpqXid2_2;
	wire w_dff_B_ozkBiLVY8_2;
	wire w_dff_B_eA6gvZl36_2;
	wire w_dff_B_hsfvYqfn4_2;
	wire w_dff_B_7IV9eM1K8_2;
	wire w_dff_B_3IQy30G14_2;
	wire w_dff_B_QF05wyeV8_2;
	wire w_dff_B_6gY4hOPR1_2;
	wire w_dff_B_hYDsCOy90_2;
	wire w_dff_B_Iq8m2WdW3_2;
	wire w_dff_B_Fo6RKRtK0_2;
	wire w_dff_B_PPbiLaxP4_2;
	wire w_dff_B_qfUqshtS3_2;
	wire w_dff_B_HAn7BQya3_2;
	wire w_dff_B_o6nKKGqA4_2;
	wire w_dff_B_W3KqP1vG5_2;
	wire w_dff_B_7HT5c9Ez2_2;
	wire w_dff_B_P5rom5oU2_2;
	wire w_dff_B_aIRjaaT32_2;
	wire w_dff_B_qhDAxbfJ7_2;
	wire w_dff_B_AjlORad90_2;
	wire w_dff_B_wXnEFDJP0_2;
	wire w_dff_B_akapbC7f5_1;
	wire w_dff_B_Cdhe2alZ3_2;
	wire w_dff_B_Xc8s8caI0_2;
	wire w_dff_B_3urXrUrZ3_2;
	wire w_dff_B_56jTcQuB8_2;
	wire w_dff_B_YA83Q8Oi2_2;
	wire w_dff_B_Ddzte2yZ6_2;
	wire w_dff_B_kcdaRHzb4_2;
	wire w_dff_B_LDt8Pycl5_2;
	wire w_dff_B_8RBtMjv79_2;
	wire w_dff_B_pZRsApnk2_2;
	wire w_dff_B_2j6luKJ57_2;
	wire w_dff_B_nCotYWDx6_2;
	wire w_dff_B_HBBJkLbV5_2;
	wire w_dff_B_Zk2TiZMg6_2;
	wire w_dff_B_Scitgxlo9_2;
	wire w_dff_B_zVYTE8Q64_2;
	wire w_dff_B_htiST99C0_2;
	wire w_dff_B_CsMAmuPH7_2;
	wire w_dff_B_TlpexhRO4_2;
	wire w_dff_B_50KEP5WD7_1;
	wire w_dff_B_Z1TeaOf85_2;
	wire w_dff_B_fccJNTth2_2;
	wire w_dff_B_muVYIs6Z0_2;
	wire w_dff_B_2QHyCNqZ1_2;
	wire w_dff_B_eEE9d9w62_2;
	wire w_dff_B_piToqil80_2;
	wire w_dff_B_oQCZKjdf1_2;
	wire w_dff_B_xLwPjdD22_2;
	wire w_dff_B_1LUUEQ075_2;
	wire w_dff_B_RAJxfbuE4_2;
	wire w_dff_B_6uxPmr7A3_2;
	wire w_dff_B_92CiVAVv7_2;
	wire w_dff_B_Zu1tM6Io1_2;
	wire w_dff_B_SucoWBa65_2;
	wire w_dff_B_8pJGz1xv6_2;
	wire w_dff_B_hOcmHsaa3_2;
	wire w_dff_B_TXZvMaLp9_1;
	wire w_dff_B_hvmf0dpK5_2;
	wire w_dff_B_vc5hhF7P3_2;
	wire w_dff_B_vAboxJed7_2;
	wire w_dff_B_GDaAzkyS8_2;
	wire w_dff_B_gDNdf3p49_2;
	wire w_dff_B_FxfT3svE7_2;
	wire w_dff_B_guMEdJmj5_2;
	wire w_dff_B_CtvSUjyT0_2;
	wire w_dff_B_oO173jvh5_2;
	wire w_dff_B_gPYgbGhE7_2;
	wire w_dff_B_iZulZs0t8_2;
	wire w_dff_B_FoTdDfnG1_2;
	wire w_dff_B_HiolJOlV9_2;
	wire w_dff_B_NrstpOeQ0_1;
	wire w_dff_B_GQeXlzud5_2;
	wire w_dff_B_0beilgAt0_2;
	wire w_dff_B_3ss2RhTb5_2;
	wire w_dff_B_Q3DYyzPh2_2;
	wire w_dff_B_719WvJAH0_2;
	wire w_dff_B_LQSDncny9_2;
	wire w_dff_B_7rBiztZi3_2;
	wire w_dff_B_60wxpPpz4_2;
	wire w_dff_B_45LVaV9I9_2;
	wire w_dff_B_8C6irrye9_2;
	wire w_dff_B_lYkQHvFO0_2;
	wire w_dff_B_BsPgbHp52_1;
	wire w_dff_B_ueJL4jap8_1;
	wire w_dff_B_QnoYSYpE9_1;
	wire w_dff_B_O29eXEyM1_1;
	wire w_dff_B_B5BTH9ym8_1;
	wire w_dff_B_aSZoaJ0K5_1;
	wire w_dff_B_rcbFvTAZ5_0;
	wire w_dff_B_KMrHkR3x1_0;
	wire w_dff_A_rRBiOC0i3_0;
	wire w_dff_A_y1T94mrB0_0;
	wire w_dff_A_wYtxhkNR9_0;
	wire w_dff_B_wP9WFB291_1;
	wire w_dff_A_ahOAYgm48_0;
	wire w_dff_A_j98TKgFe4_1;
	wire w_dff_A_N92C5aQQ8_1;
	wire w_dff_A_HgPoA1yu6_1;
	wire w_dff_A_dolF8lSb0_1;
	wire w_dff_A_0eUDpDWO3_1;
	wire w_dff_A_YOjFMLg99_1;
	wire w_dff_A_gnSkQPUF5_1;
	wire w_dff_A_evwGOEkL4_1;
	wire w_dff_B_6I2knGDc5_2;
	wire w_dff_B_DlNTa9EC7_2;
	wire w_dff_B_EkZtMXUx2_1;
	wire w_dff_B_ubP4Wdas1_2;
	wire w_dff_B_dS7lo7wE7_2;
	wire w_dff_B_3lAGRwe02_2;
	wire w_dff_B_DF2O6JJH6_2;
	wire w_dff_B_z6aCkRW00_2;
	wire w_dff_B_2etEtMpm6_2;
	wire w_dff_B_dM4QFiMw2_2;
	wire w_dff_B_2yQ2y7g95_2;
	wire w_dff_B_wKWoGesb3_2;
	wire w_dff_B_84NLMqOb9_2;
	wire w_dff_B_uf1EqLnv8_2;
	wire w_dff_B_3QbwMOam5_2;
	wire w_dff_B_SO8TDBDr4_2;
	wire w_dff_B_4tgEq3PU0_2;
	wire w_dff_B_Spu0gkCn5_2;
	wire w_dff_B_NJAlfSUW4_2;
	wire w_dff_B_x5OsXYSJ8_2;
	wire w_dff_B_KdhXDiYh3_2;
	wire w_dff_B_CKwbgnXW0_2;
	wire w_dff_B_kcByU88V1_2;
	wire w_dff_B_heUYiaTb6_2;
	wire w_dff_B_CWZPdP6U1_2;
	wire w_dff_B_DUHs937k4_2;
	wire w_dff_B_IioNZuZc3_2;
	wire w_dff_B_B9vIPMFR2_2;
	wire w_dff_B_N80iKUl86_2;
	wire w_dff_B_ttFVcsjR6_2;
	wire w_dff_B_THKSeorq9_2;
	wire w_dff_B_w0GMMlyp1_2;
	wire w_dff_B_Yxrf35pC7_2;
	wire w_dff_B_4Il2zcGd3_2;
	wire w_dff_B_hS6HtJUS4_2;
	wire w_dff_B_OYsJtcii9_2;
	wire w_dff_B_teUgY3HQ3_2;
	wire w_dff_B_u5c6ACBd6_2;
	wire w_dff_B_3VTx7P0T4_2;
	wire w_dff_B_g0Tf01TQ6_2;
	wire w_dff_B_WklhyrFh5_2;
	wire w_dff_B_31PN68Rk6_2;
	wire w_dff_B_TVlstJ6z2_2;
	wire w_dff_B_AjfAb4Rw8_2;
	wire w_dff_B_gBeuXSrg7_2;
	wire w_dff_B_5W3R03Kh1_2;
	wire w_dff_B_1aagcxQJ3_2;
	wire w_dff_B_610dQHof7_2;
	wire w_dff_B_ue8UUm0w1_2;
	wire w_dff_B_EVsqjVM83_2;
	wire w_dff_B_CdmtuydS5_1;
	wire w_dff_B_sxuDsbth0_2;
	wire w_dff_B_HzuHDBeP6_2;
	wire w_dff_B_T7oGcoNR3_2;
	wire w_dff_B_VQjfX0IM0_2;
	wire w_dff_B_h9BWaBXz0_2;
	wire w_dff_B_bTqfafHR7_2;
	wire w_dff_B_VMReU0S91_2;
	wire w_dff_B_P0hUCw0P0_2;
	wire w_dff_B_1HrcFrfi5_2;
	wire w_dff_B_uesnWeIG6_2;
	wire w_dff_B_vy6soyIt7_2;
	wire w_dff_B_2MKAJuKf8_2;
	wire w_dff_B_kZu3kG5s9_2;
	wire w_dff_B_IXH8WcCY9_2;
	wire w_dff_B_WjKF1KD99_2;
	wire w_dff_B_Dplf3ms51_2;
	wire w_dff_B_toTQhYKo8_2;
	wire w_dff_B_ibv82bX53_2;
	wire w_dff_B_jfiRjN7D4_2;
	wire w_dff_B_u8pQr0sd9_2;
	wire w_dff_B_WzRyQTej3_2;
	wire w_dff_B_ZqudcncV3_2;
	wire w_dff_B_Mv27uzwL3_2;
	wire w_dff_B_9duGwFgx7_2;
	wire w_dff_B_rVOXfMG23_2;
	wire w_dff_B_9zZnf4xZ4_2;
	wire w_dff_B_pICOT8mK6_2;
	wire w_dff_B_mZ2Pe8Zs1_2;
	wire w_dff_B_5VafzWNx4_2;
	wire w_dff_B_T20zpEtB5_2;
	wire w_dff_B_naGH2sfc0_2;
	wire w_dff_B_SmYMYUcR2_2;
	wire w_dff_B_dfywWW1T7_2;
	wire w_dff_B_FSTInDsE4_2;
	wire w_dff_B_oU7SjGEV6_2;
	wire w_dff_B_DhItVa4b0_2;
	wire w_dff_B_DM4qzMub8_2;
	wire w_dff_B_jr1AaHBJ1_2;
	wire w_dff_B_OBes7WtX2_2;
	wire w_dff_B_iJMIQNGM2_2;
	wire w_dff_B_OgRPnqI63_2;
	wire w_dff_B_TLbaPM3u0_2;
	wire w_dff_B_OzTc8R7Z8_2;
	wire w_dff_B_aRK956Io7_1;
	wire w_dff_B_7OEaWOFM5_2;
	wire w_dff_B_vbdHOdD61_2;
	wire w_dff_B_MgOg3O739_2;
	wire w_dff_B_r3VCoTHa5_2;
	wire w_dff_B_4L3JdPvB6_2;
	wire w_dff_B_slHNYECG7_2;
	wire w_dff_B_xEOONrcV2_2;
	wire w_dff_B_bwZdFMpz3_2;
	wire w_dff_B_zrS0wVTp4_2;
	wire w_dff_B_BgugZ0gV1_2;
	wire w_dff_B_39Q4ytw93_2;
	wire w_dff_B_Ir3EyOh10_2;
	wire w_dff_B_x6LYUNE72_2;
	wire w_dff_B_lNsOoBoq9_2;
	wire w_dff_B_MK4LfCtl3_2;
	wire w_dff_B_nNNIllSw4_2;
	wire w_dff_B_ORf6ql5j2_2;
	wire w_dff_B_VpXoKOYz5_2;
	wire w_dff_B_praYt60y0_2;
	wire w_dff_B_uUTCZeEs8_2;
	wire w_dff_B_aAIaCyAP8_2;
	wire w_dff_B_l5uhyDoT0_2;
	wire w_dff_B_gUGeMuOa0_2;
	wire w_dff_B_0vH9r3UA2_2;
	wire w_dff_B_QPujcOcK3_2;
	wire w_dff_B_uXk0qGrU1_2;
	wire w_dff_B_Cd5vAkuo7_2;
	wire w_dff_B_HrNndOAC0_2;
	wire w_dff_B_ZjZLhMMJ0_2;
	wire w_dff_B_NA0zjnQs9_2;
	wire w_dff_B_bKvuNu7H1_2;
	wire w_dff_B_anbhfeed7_2;
	wire w_dff_B_TyEoFMTR6_2;
	wire w_dff_B_brb85nqy7_2;
	wire w_dff_B_t1hNhFKR7_2;
	wire w_dff_B_A552WBmt3_2;
	wire w_dff_B_0G3AblGa3_2;
	wire w_dff_B_Lrp9Mhk18_2;
	wire w_dff_B_xqaVoTr96_2;
	wire w_dff_B_gCURn5tp9_2;
	wire w_dff_B_BlR6EJkB2_1;
	wire w_dff_B_AZN01NqR1_2;
	wire w_dff_B_HarpwzLK1_2;
	wire w_dff_B_RRrPOGVW4_2;
	wire w_dff_B_uXVhy4AP5_2;
	wire w_dff_B_CqD4oQ3g5_2;
	wire w_dff_B_7EUXIAYI3_2;
	wire w_dff_B_o1Nf8nId1_2;
	wire w_dff_B_XCXBjBFW6_2;
	wire w_dff_B_kmLVOZc66_2;
	wire w_dff_B_aUlj0tMX7_2;
	wire w_dff_B_VjgxiZoj7_2;
	wire w_dff_B_4AaBljX49_2;
	wire w_dff_B_FHdesKAm3_2;
	wire w_dff_B_dkpHPHTX8_2;
	wire w_dff_B_NSvE7o3u9_2;
	wire w_dff_B_Kvrrxyx49_2;
	wire w_dff_B_t3NzRcBg1_2;
	wire w_dff_B_5gohuiQp0_2;
	wire w_dff_B_eCKb4z697_2;
	wire w_dff_B_4T2rRRjW8_2;
	wire w_dff_B_v8jP46p51_2;
	wire w_dff_B_mQDVsplr8_2;
	wire w_dff_B_XRcFEKP07_2;
	wire w_dff_B_miN0aHYX5_2;
	wire w_dff_B_f8tEK2dq2_2;
	wire w_dff_B_KUJuGNsV2_2;
	wire w_dff_B_pHDRcmR51_2;
	wire w_dff_B_YHtoN35Y2_2;
	wire w_dff_B_nisqSuFC3_2;
	wire w_dff_B_Vcs2YyyL3_2;
	wire w_dff_B_YRJXmm4d1_2;
	wire w_dff_B_avE36V7U8_2;
	wire w_dff_B_gupLnxqX3_2;
	wire w_dff_B_enY74l0d2_2;
	wire w_dff_B_xEAcDscs6_2;
	wire w_dff_B_Patk0o6B2_2;
	wire w_dff_B_PpKZCrKf2_2;
	wire w_dff_B_FzF9b9Ge7_1;
	wire w_dff_B_lPFQZYYF1_2;
	wire w_dff_B_iJQN5Sud1_2;
	wire w_dff_B_zSCAmNSA4_2;
	wire w_dff_B_TbaZtBKf4_2;
	wire w_dff_B_pgY9WjaR5_2;
	wire w_dff_B_i2miKn7D5_2;
	wire w_dff_B_dwGCvwxX2_2;
	wire w_dff_B_nCRjsMjQ9_2;
	wire w_dff_B_tVoIQ5wF4_2;
	wire w_dff_B_I9YAnaHK0_2;
	wire w_dff_B_FbkEBOwC4_2;
	wire w_dff_B_vaBNNtNn3_2;
	wire w_dff_B_LbtjHO9Z6_2;
	wire w_dff_B_UHx5HpJW3_2;
	wire w_dff_B_oMYBigI99_2;
	wire w_dff_B_0VTcO1vk3_2;
	wire w_dff_B_s0tQSQD75_2;
	wire w_dff_B_cxYAnOAR4_2;
	wire w_dff_B_Jc4RGxH64_2;
	wire w_dff_B_XfhYZyNu6_2;
	wire w_dff_B_YH5mPmX65_2;
	wire w_dff_B_bZMqbk7c3_2;
	wire w_dff_B_PKKC6atd7_2;
	wire w_dff_B_wAHjK5OM4_2;
	wire w_dff_B_Iw5ueGsH7_2;
	wire w_dff_B_BOUJUf7R6_2;
	wire w_dff_B_YeExXbwh8_2;
	wire w_dff_B_lAYEKKoZ4_2;
	wire w_dff_B_mLTDj1ur8_2;
	wire w_dff_B_8oYXsYGA1_2;
	wire w_dff_B_VggqWUL69_2;
	wire w_dff_B_swd6VmrS0_2;
	wire w_dff_B_20xgkSPY9_2;
	wire w_dff_B_xSk7omfA1_2;
	wire w_dff_B_ScPyrVF34_1;
	wire w_dff_B_sFiR5tEY5_2;
	wire w_dff_B_UnPw4Kie4_2;
	wire w_dff_B_ohWgRbZY0_2;
	wire w_dff_B_ZLwjlKpF3_2;
	wire w_dff_B_6F7TUjP04_2;
	wire w_dff_B_HZv5SsZW7_2;
	wire w_dff_B_1XqV9wbH1_2;
	wire w_dff_B_f92aTyxH2_2;
	wire w_dff_B_3OWiSrvp2_2;
	wire w_dff_B_DK6jW7Me2_2;
	wire w_dff_B_F2LSVmmD7_2;
	wire w_dff_B_3eVzFBCr0_2;
	wire w_dff_B_DdwjIYGD6_2;
	wire w_dff_B_h9UXEoPm3_2;
	wire w_dff_B_rs5s9YpB4_2;
	wire w_dff_B_SZ1YAXcV1_2;
	wire w_dff_B_rDpriOgC5_2;
	wire w_dff_B_uqTahcw47_2;
	wire w_dff_B_bsdKYveB5_2;
	wire w_dff_B_ga8Y9ufL9_2;
	wire w_dff_B_IdXGlFdY1_2;
	wire w_dff_B_jxx4Skw51_2;
	wire w_dff_B_KDyzA9ow3_2;
	wire w_dff_B_EApnyhfk6_2;
	wire w_dff_B_I2hBWnyA5_2;
	wire w_dff_B_7uvoe9dF3_2;
	wire w_dff_B_kwO31D1A2_2;
	wire w_dff_B_g3DsQ5Nu8_2;
	wire w_dff_B_Lnnx9r0k6_2;
	wire w_dff_B_2l75t1df1_2;
	wire w_dff_B_06mQNvWb6_2;
	wire w_dff_B_buQPiXvj6_1;
	wire w_dff_B_lKOzpYjF5_2;
	wire w_dff_B_QtOqGyEj6_2;
	wire w_dff_B_vXbR900i4_2;
	wire w_dff_B_PJZ4Sj7W5_2;
	wire w_dff_B_5zxKD1uS1_2;
	wire w_dff_B_u5umJbrT3_2;
	wire w_dff_B_4DbieKDR6_2;
	wire w_dff_B_8Xc0qH8Q7_2;
	wire w_dff_B_3IwaWNBe9_2;
	wire w_dff_B_lstUPp760_2;
	wire w_dff_B_ObUwMK1Z5_2;
	wire w_dff_B_SEy8Udo97_2;
	wire w_dff_B_E2Sd5Uo40_2;
	wire w_dff_B_hVoxkf8Y0_2;
	wire w_dff_B_uly6CBGn7_2;
	wire w_dff_B_VNy9mvCG3_2;
	wire w_dff_B_osQLCnzQ4_2;
	wire w_dff_B_zV4r5tJg0_2;
	wire w_dff_B_V8ecpqJ66_2;
	wire w_dff_B_97GtppLO6_2;
	wire w_dff_B_cCGH2UfC9_2;
	wire w_dff_B_LegMgFmk3_2;
	wire w_dff_B_ugYc6VgR7_2;
	wire w_dff_B_IQpYjBsH7_2;
	wire w_dff_B_HSFqCjXr2_2;
	wire w_dff_B_vURq43Iq4_2;
	wire w_dff_B_2OVZiyHD6_2;
	wire w_dff_B_o0s09aK91_2;
	wire w_dff_B_EkaceZ4V3_1;
	wire w_dff_B_WZraOng41_2;
	wire w_dff_B_tuXRDdq15_2;
	wire w_dff_B_aV6kqfA96_2;
	wire w_dff_B_kbbTU9Lb3_2;
	wire w_dff_B_rBBeuNnG8_2;
	wire w_dff_B_4g6d9G5j8_2;
	wire w_dff_B_5f7ZHxoN4_2;
	wire w_dff_B_2X1I82Bi2_2;
	wire w_dff_B_O2ugICkc3_2;
	wire w_dff_B_9aP4QBAP7_2;
	wire w_dff_B_EqxxATn63_2;
	wire w_dff_B_aGWVTnKh6_2;
	wire w_dff_B_emYZGCaH5_2;
	wire w_dff_B_QDRa7PTO6_2;
	wire w_dff_B_AZXS3gTZ3_2;
	wire w_dff_B_cXO8BBRn6_2;
	wire w_dff_B_vmkl23lR7_2;
	wire w_dff_B_cLXB7JSd8_2;
	wire w_dff_B_e9xHyCbH4_2;
	wire w_dff_B_QXk2LXtD6_2;
	wire w_dff_B_sJ9jJqfW3_2;
	wire w_dff_B_XsdUtOc81_2;
	wire w_dff_B_NIfLEVKF7_2;
	wire w_dff_B_5gsdl4R01_2;
	wire w_dff_B_CuRktE837_2;
	wire w_dff_B_nncCmUwm5_1;
	wire w_dff_B_Wydq4k9Q5_2;
	wire w_dff_B_QTUOfhUV6_2;
	wire w_dff_B_ItN14GvT0_2;
	wire w_dff_B_lJoiSbgk9_2;
	wire w_dff_B_m18D4wSX1_2;
	wire w_dff_B_zbnIlKzT9_2;
	wire w_dff_B_3naIsnxH6_2;
	wire w_dff_B_1CPGJZLE6_2;
	wire w_dff_B_86oTyfjN9_2;
	wire w_dff_B_xPyKY8817_2;
	wire w_dff_B_9kAEL1bO5_2;
	wire w_dff_B_9b3RdcXm4_2;
	wire w_dff_B_3hpc6nPF2_2;
	wire w_dff_B_uMtkItIw9_2;
	wire w_dff_B_MKmObVUb1_2;
	wire w_dff_B_VuzFrZNL5_2;
	wire w_dff_B_pbb5q2Zf8_2;
	wire w_dff_B_wkoLnsZ62_2;
	wire w_dff_B_bi7cHT8i5_2;
	wire w_dff_B_4Kydrbx06_2;
	wire w_dff_B_6nbRevOp8_2;
	wire w_dff_B_4QWmYAAQ7_2;
	wire w_dff_B_jyFNJZ921_1;
	wire w_dff_B_lcdzaeZM2_2;
	wire w_dff_B_qaTI2bvq7_2;
	wire w_dff_B_96YTQVBa9_2;
	wire w_dff_B_TRZdrml47_2;
	wire w_dff_B_6AYmfj6H6_2;
	wire w_dff_B_XuBtdsvm0_2;
	wire w_dff_B_R5pZwYaa1_2;
	wire w_dff_B_hBEez6Zn9_2;
	wire w_dff_B_FNz6hEYy3_2;
	wire w_dff_B_MuE07MkQ4_2;
	wire w_dff_B_Yc33j1h25_2;
	wire w_dff_B_xjQuS2G13_2;
	wire w_dff_B_Mgmt5gov8_2;
	wire w_dff_B_b5oeM0lI5_2;
	wire w_dff_B_qgLEczf59_2;
	wire w_dff_B_fT5eBe3o3_2;
	wire w_dff_B_BaqnRUWR7_2;
	wire w_dff_B_IgHq9uxs3_2;
	wire w_dff_B_Z9zB7At31_2;
	wire w_dff_B_X2359Wtm1_1;
	wire w_dff_B_wHreRi5L3_2;
	wire w_dff_B_aF6BvOZO9_2;
	wire w_dff_B_mY8Jb0KE5_2;
	wire w_dff_B_6Q0BL26h6_2;
	wire w_dff_B_KwP8AI9b1_2;
	wire w_dff_B_gXZ7ufps6_2;
	wire w_dff_B_SFGv87qC9_2;
	wire w_dff_B_3SEij5VD0_2;
	wire w_dff_B_sME06cnY8_2;
	wire w_dff_B_OD1yKOzs3_2;
	wire w_dff_B_TvCgD8ks9_2;
	wire w_dff_B_dmQnRqLb9_2;
	wire w_dff_B_rztMr0lF8_2;
	wire w_dff_B_fzIesVWp9_2;
	wire w_dff_B_RJPkQgDR3_2;
	wire w_dff_B_hrRlyOSk0_2;
	wire w_dff_B_ylrELTML5_1;
	wire w_dff_B_5WgVRk198_2;
	wire w_dff_B_9En3TXtx4_2;
	wire w_dff_B_RC63I0fB5_2;
	wire w_dff_B_odALINGx2_2;
	wire w_dff_B_D1GKbF0c6_2;
	wire w_dff_B_7sCYzbVI1_2;
	wire w_dff_B_si04EEu89_2;
	wire w_dff_B_AiT3i1To3_2;
	wire w_dff_B_vMDhyFHi7_2;
	wire w_dff_B_JU5pyfFM9_2;
	wire w_dff_B_ekup89cH3_2;
	wire w_dff_B_T57MD6st6_2;
	wire w_dff_B_HPEZ81tM1_2;
	wire w_dff_B_0hhdmz5A7_1;
	wire w_dff_B_GJ0sQQWE4_2;
	wire w_dff_B_BMAXM5ca2_2;
	wire w_dff_B_rgAEmIhb9_2;
	wire w_dff_B_z9jxILgS7_2;
	wire w_dff_B_Yn1lVPN73_2;
	wire w_dff_B_xELfyWBf3_2;
	wire w_dff_B_7FJmKZb81_2;
	wire w_dff_B_PamvgK1M7_2;
	wire w_dff_B_aESPuByd0_2;
	wire w_dff_B_dk64gEpf4_2;
	wire w_dff_B_0jqNEiRK1_2;
	wire w_dff_B_0cZVaPms4_1;
	wire w_dff_B_J9N6v84s1_1;
	wire w_dff_B_ATxOrPEq5_1;
	wire w_dff_B_Gp0urcmt4_1;
	wire w_dff_B_fKbhMkZJ9_1;
	wire w_dff_B_7b9zcMbq5_1;
	wire w_dff_B_qt3Ns1xz6_0;
	wire w_dff_B_UK5oVL1A8_0;
	wire w_dff_A_4mbiZx7q8_0;
	wire w_dff_A_c7F6NGBy7_0;
	wire w_dff_A_PLejDV5i4_0;
	wire w_dff_B_B7uYD8kd4_1;
	wire w_dff_A_xQ8IgenW8_0;
	wire w_dff_A_gZ3zpvUA2_1;
	wire w_dff_A_xriyLzyx7_1;
	wire w_dff_A_oBtVO8qU7_1;
	wire w_dff_A_wFrnZpCI9_1;
	wire w_dff_A_FU0O2HPX9_1;
	wire w_dff_A_PF47EiG56_1;
	wire w_dff_A_7OB2ckyA4_1;
	wire w_dff_A_BbMEquCd0_1;
	wire w_dff_B_HeUhQdQa6_2;
	wire w_dff_B_lVy3GB6O5_1;
	wire w_dff_B_dQ3WJGGw7_2;
	wire w_dff_B_ldTcfqoU8_2;
	wire w_dff_B_yZ6BmJrI4_2;
	wire w_dff_B_xNLBdxsk3_2;
	wire w_dff_B_qNahotcy8_2;
	wire w_dff_B_mOawhLJI5_2;
	wire w_dff_B_TZUyEKTw9_2;
	wire w_dff_B_wsvjI5u81_2;
	wire w_dff_B_E6fgUefI1_2;
	wire w_dff_B_ktuDovzW2_2;
	wire w_dff_B_o1Wt4ZNl8_2;
	wire w_dff_B_JehvfdXY1_2;
	wire w_dff_B_pCYdOBkA6_2;
	wire w_dff_B_aZ9m9OjY1_2;
	wire w_dff_B_6GX5ZKiK9_2;
	wire w_dff_B_YS5Xjf8n2_2;
	wire w_dff_B_z459SVYz5_2;
	wire w_dff_B_vZsySrL29_2;
	wire w_dff_B_Tp1rGKHW1_2;
	wire w_dff_B_xxkAWJ7F4_2;
	wire w_dff_B_xHCqNPXw2_2;
	wire w_dff_B_UE3jvtuC3_2;
	wire w_dff_B_EkKxvFEV9_2;
	wire w_dff_B_wIkZEgwB4_2;
	wire w_dff_B_cwMFckBl9_2;
	wire w_dff_B_Lp9EeNir3_2;
	wire w_dff_B_BddIGRgw3_2;
	wire w_dff_B_JRcY3adb9_2;
	wire w_dff_B_Nmfldyfe3_2;
	wire w_dff_B_4r3f1oaR5_2;
	wire w_dff_B_M1cAbZWF5_2;
	wire w_dff_B_bSafRusd4_2;
	wire w_dff_B_NTkWFEcR1_2;
	wire w_dff_B_mtWm4W9N8_2;
	wire w_dff_B_OBp95y760_2;
	wire w_dff_B_yhdYSiQ66_2;
	wire w_dff_B_zkNt7NFy7_2;
	wire w_dff_B_GxcqJDat1_2;
	wire w_dff_B_ulZu1MnZ8_2;
	wire w_dff_B_GofV90ru9_2;
	wire w_dff_B_Hk0erdO04_2;
	wire w_dff_B_WQuHzJOg2_2;
	wire w_dff_B_iLUMRCel7_2;
	wire w_dff_B_Hp2dnVpw2_2;
	wire w_dff_B_6PCJZvOy1_2;
	wire w_dff_B_vKAYiyDw8_2;
	wire w_dff_B_rkJpFx9l6_2;
	wire w_dff_B_FkJQaaKQ6_2;
	wire w_dff_B_Zcxv3EB42_2;
	wire w_dff_B_1uK7f00G7_1;
	wire w_dff_A_zzjBz9dq1_1;
	wire w_dff_B_8piwo4me2_1;
	wire w_dff_B_GNtZnVvZ6_2;
	wire w_dff_B_BC58j5F35_2;
	wire w_dff_B_tBUC1MJV0_2;
	wire w_dff_B_W3BlvzBt7_2;
	wire w_dff_B_fkrU0qgZ0_2;
	wire w_dff_B_0IJ2MFpn8_2;
	wire w_dff_B_NtEEfmxq6_2;
	wire w_dff_B_oDfhuqqw5_2;
	wire w_dff_B_O1v0LXH27_2;
	wire w_dff_B_6hsAkfUT4_2;
	wire w_dff_B_uKeW7jMU2_2;
	wire w_dff_B_telpEeq35_2;
	wire w_dff_B_WjQ3XbRQ8_2;
	wire w_dff_B_ljMxDcrC3_2;
	wire w_dff_B_LYdDuLik0_2;
	wire w_dff_B_3bvJ530v8_2;
	wire w_dff_B_85rzEYy74_2;
	wire w_dff_B_6bfBNvak7_2;
	wire w_dff_B_nKxXDu9m9_2;
	wire w_dff_B_ZK55cj8A1_2;
	wire w_dff_B_v7Jz1dQl8_2;
	wire w_dff_B_GSQbuvq19_2;
	wire w_dff_B_BHwTPlm92_2;
	wire w_dff_B_0O5ul9Ub9_2;
	wire w_dff_B_T7aQKPFW2_2;
	wire w_dff_B_pn3FhFV56_2;
	wire w_dff_B_mWeyXP3g8_2;
	wire w_dff_B_wuBXv44K0_2;
	wire w_dff_B_RyPlMtWv9_2;
	wire w_dff_B_euzJQrrl4_2;
	wire w_dff_B_97zkkpKf2_2;
	wire w_dff_B_gA1ogjDf1_2;
	wire w_dff_B_ZN5G2luJ2_2;
	wire w_dff_B_sa8PHzss0_2;
	wire w_dff_B_1OPCSsHP9_2;
	wire w_dff_B_HAPxhBxl3_2;
	wire w_dff_B_DKbrqyWa3_2;
	wire w_dff_B_9qOsFu9L6_2;
	wire w_dff_B_SKOBbt7E1_2;
	wire w_dff_B_Ylbd4SZn3_2;
	wire w_dff_B_XCDLpu8W2_2;
	wire w_dff_B_yCq2Ccq29_2;
	wire w_dff_B_wG1Npweu9_2;
	wire w_dff_B_Noqgof8s2_2;
	wire w_dff_B_tX56hz7o5_1;
	wire w_dff_B_9FCnLDfC0_2;
	wire w_dff_B_QILD84OU0_2;
	wire w_dff_B_SlzcR0VO9_2;
	wire w_dff_B_UBgjGxke7_2;
	wire w_dff_B_0cXQYiqv7_2;
	wire w_dff_B_DRzKXMe08_2;
	wire w_dff_B_txBI72Yv5_2;
	wire w_dff_B_GtA5nQ8y6_2;
	wire w_dff_B_21a9CdXg4_2;
	wire w_dff_B_b3WqfLXW9_2;
	wire w_dff_B_0R5jye7Y0_2;
	wire w_dff_B_qxEdKKvB9_2;
	wire w_dff_B_8FHL79Kr7_2;
	wire w_dff_B_lKwL8on02_2;
	wire w_dff_B_T6cuERnm2_2;
	wire w_dff_B_hbNV5vVv1_2;
	wire w_dff_B_V1usOsl04_2;
	wire w_dff_B_YNtdHl5H2_2;
	wire w_dff_B_41oDOv7S4_2;
	wire w_dff_B_Av24EUB60_2;
	wire w_dff_B_etygBPsg4_2;
	wire w_dff_B_37pUb7NC7_2;
	wire w_dff_B_O76lKCOF6_2;
	wire w_dff_B_nORxJQ7s2_2;
	wire w_dff_B_VzZVCbWW8_2;
	wire w_dff_B_mZa67PnZ2_2;
	wire w_dff_B_X6RWB88F6_2;
	wire w_dff_B_CwGiKdgi9_2;
	wire w_dff_B_4itIrE3x9_2;
	wire w_dff_B_dTG4LYCM5_2;
	wire w_dff_B_CuIpjjBq1_2;
	wire w_dff_B_jy9S97pJ4_2;
	wire w_dff_B_OuLfGXr64_2;
	wire w_dff_B_vnVYfSRN1_2;
	wire w_dff_B_0nkKLhek2_2;
	wire w_dff_B_JKtBWnzS4_2;
	wire w_dff_B_fkcq9az63_2;
	wire w_dff_B_kDxvW6Z86_2;
	wire w_dff_B_k7ju0uw85_2;
	wire w_dff_B_6NaOW2oA3_1;
	wire w_dff_B_nF1gvEjr2_2;
	wire w_dff_B_CsWCo8Xl3_2;
	wire w_dff_B_aR9Py4x91_2;
	wire w_dff_B_ZkldLel05_2;
	wire w_dff_B_WmGppmAH4_2;
	wire w_dff_B_83D1O2ez9_2;
	wire w_dff_B_V0QG3D9p3_2;
	wire w_dff_B_d2eu5nKd1_2;
	wire w_dff_B_veuu8M036_2;
	wire w_dff_B_yRRLMSK59_2;
	wire w_dff_B_8fR9fykw8_2;
	wire w_dff_B_epPw27jC9_2;
	wire w_dff_B_l0jY552I6_2;
	wire w_dff_B_ulOYps4L6_2;
	wire w_dff_B_RKaAF2Bz0_2;
	wire w_dff_B_hixJMzbZ9_2;
	wire w_dff_B_SqpKesEp6_2;
	wire w_dff_B_eVOb76Xz6_2;
	wire w_dff_B_XCkHZtnd5_2;
	wire w_dff_B_TdGdLDEh4_2;
	wire w_dff_B_wyMWoNYX2_2;
	wire w_dff_B_mGxCDdZ50_2;
	wire w_dff_B_YEuEAVZI6_2;
	wire w_dff_B_WFzf4FDq0_2;
	wire w_dff_B_iRgy355T2_2;
	wire w_dff_B_dtcmYRqc6_2;
	wire w_dff_B_MOJ18p1E3_2;
	wire w_dff_B_KOtE8ltQ8_2;
	wire w_dff_B_ghuSZZYC5_2;
	wire w_dff_B_npqSoASv5_2;
	wire w_dff_B_jBDlSCiV5_2;
	wire w_dff_B_A3VBZ0HC6_2;
	wire w_dff_B_t3u4FL7p9_2;
	wire w_dff_B_TQfQi3H54_2;
	wire w_dff_B_CFl6tAIv5_2;
	wire w_dff_B_apora1Ov2_2;
	wire w_dff_B_Jmxx0iWk6_2;
	wire w_dff_B_0zbkiSiI3_1;
	wire w_dff_B_ULwV9H8K6_2;
	wire w_dff_B_xLGopkgf0_2;
	wire w_dff_B_kNmXhQ9E1_2;
	wire w_dff_B_x645mFm42_2;
	wire w_dff_B_X4QKCLC96_2;
	wire w_dff_B_fz3qGhTS1_2;
	wire w_dff_B_8zP02RlI7_2;
	wire w_dff_B_logvZ88f8_2;
	wire w_dff_B_Z2Id0T8t7_2;
	wire w_dff_B_4V1y7eKD5_2;
	wire w_dff_B_Ml2hwIKz8_2;
	wire w_dff_B_zCSbThxH9_2;
	wire w_dff_B_jGWAjlyS7_2;
	wire w_dff_B_zFz9ZT6K1_2;
	wire w_dff_B_yuzxBeyp6_2;
	wire w_dff_B_FawMs8CI6_2;
	wire w_dff_B_4nMrm7rk6_2;
	wire w_dff_B_O4o09TlU8_2;
	wire w_dff_B_L130e9Lv0_2;
	wire w_dff_B_AgqRvNee2_2;
	wire w_dff_B_9gYvM1Gb5_2;
	wire w_dff_B_Gz9EnSyV9_2;
	wire w_dff_B_F2YcDJsJ5_2;
	wire w_dff_B_6Ous1wom8_2;
	wire w_dff_B_QMsrHuJN5_2;
	wire w_dff_B_QXh3l63O4_2;
	wire w_dff_B_V5mVErpJ3_2;
	wire w_dff_B_Q9VBhwBD2_2;
	wire w_dff_B_uXcl4qyC6_2;
	wire w_dff_B_iGM9JZXL6_2;
	wire w_dff_B_NfLRQCCH1_2;
	wire w_dff_B_K4Osp7Zy8_2;
	wire w_dff_B_ZKhslv1z7_2;
	wire w_dff_B_wETVknfo3_2;
	wire w_dff_B_CE7lS43i5_1;
	wire w_dff_B_oSkge1wz6_2;
	wire w_dff_B_OZNWplzX5_2;
	wire w_dff_B_i2w7qUCi6_2;
	wire w_dff_B_WBafffGL1_2;
	wire w_dff_B_U9IasaPX0_2;
	wire w_dff_B_7oxxEOqn1_2;
	wire w_dff_B_hOVdS20Q4_2;
	wire w_dff_B_jzhZiZJb8_2;
	wire w_dff_B_jTONLOKF2_2;
	wire w_dff_B_eAELwhp47_2;
	wire w_dff_B_FB2ZC8Lh0_2;
	wire w_dff_B_hYGyFPaf4_2;
	wire w_dff_B_Ud8xlKNQ2_2;
	wire w_dff_B_ILOug0Gv0_2;
	wire w_dff_B_o7fHHtYa3_2;
	wire w_dff_B_e3JSNZto0_2;
	wire w_dff_B_XkPs0ArA9_2;
	wire w_dff_B_HZ29W4hh4_2;
	wire w_dff_B_ohXKGGyO3_2;
	wire w_dff_B_kHmhPEwo2_2;
	wire w_dff_B_P6WKDGfg9_2;
	wire w_dff_B_j2uuOPfn3_2;
	wire w_dff_B_MdQBCLTg5_2;
	wire w_dff_B_zthjBxNu4_2;
	wire w_dff_B_nWdVCvXM9_2;
	wire w_dff_B_2teXDn471_2;
	wire w_dff_B_YVTNBWn52_2;
	wire w_dff_B_FOsclKzN3_2;
	wire w_dff_B_YSkeVL2d6_2;
	wire w_dff_B_w0rM8Gjh0_2;
	wire w_dff_B_rTBOuZFw4_2;
	wire w_dff_B_2pzKa2wU6_1;
	wire w_dff_B_ZUlZ66mh1_2;
	wire w_dff_B_X2hyDXX12_2;
	wire w_dff_B_lP4BmWsy2_2;
	wire w_dff_B_gDpP7nfq6_2;
	wire w_dff_B_J5CRVO5y2_2;
	wire w_dff_B_glqvyk642_2;
	wire w_dff_B_SxCFBQLJ0_2;
	wire w_dff_B_Yy3lo1wa7_2;
	wire w_dff_B_yV4xYn2e2_2;
	wire w_dff_B_n3kDKDkW6_2;
	wire w_dff_B_OugAvdJv6_2;
	wire w_dff_B_WwZaeYDE7_2;
	wire w_dff_B_sSENcVUd2_2;
	wire w_dff_B_drzbCvJF2_2;
	wire w_dff_B_6pnHQkNz0_2;
	wire w_dff_B_GHGRV3z03_2;
	wire w_dff_B_kx2W5BoE2_2;
	wire w_dff_B_fCBQU8gt7_2;
	wire w_dff_B_Kwpo1Oyz0_2;
	wire w_dff_B_voDm8Txc9_2;
	wire w_dff_B_GhN36jN26_2;
	wire w_dff_B_jxzTPCt39_2;
	wire w_dff_B_WX55OYxl8_2;
	wire w_dff_B_jQb6Iy5f1_2;
	wire w_dff_B_MUmWnAOJ1_2;
	wire w_dff_B_aLcJ985A1_2;
	wire w_dff_B_UAI8SVqq1_2;
	wire w_dff_B_Z0a9KuK07_2;
	wire w_dff_B_fvxKhTZJ1_1;
	wire w_dff_B_veLj3kF07_2;
	wire w_dff_B_O7PMupaH6_2;
	wire w_dff_B_YOWYBIXb8_2;
	wire w_dff_B_DQTMxhKZ0_2;
	wire w_dff_B_AMbMvFhE4_2;
	wire w_dff_B_IbYMGAOT7_2;
	wire w_dff_B_yAzojypG2_2;
	wire w_dff_B_GDrmqKIT8_2;
	wire w_dff_B_z0gKijmK6_2;
	wire w_dff_B_aQoWeWUe4_2;
	wire w_dff_B_D00xBbtZ1_2;
	wire w_dff_B_AMRwQ9s03_2;
	wire w_dff_B_WYyPk8ze3_2;
	wire w_dff_B_6jHS5wNb1_2;
	wire w_dff_B_5aKXzY7B5_2;
	wire w_dff_B_O84dZUmr6_2;
	wire w_dff_B_2CR7ZkHZ7_2;
	wire w_dff_B_BjioOdj92_2;
	wire w_dff_B_iCCPp6X70_2;
	wire w_dff_B_3f60c6z12_2;
	wire w_dff_B_6XKfNODF8_2;
	wire w_dff_B_QT9H3YyO9_2;
	wire w_dff_B_WpwaJj4C1_2;
	wire w_dff_B_RiuwrtiS3_2;
	wire w_dff_B_CcpcWgtq1_2;
	wire w_dff_B_RJaWybtq6_1;
	wire w_dff_B_gZBphBBI3_2;
	wire w_dff_B_SR17P8wr8_2;
	wire w_dff_B_FxIyvZ0Q3_2;
	wire w_dff_B_Rjvzmweo7_2;
	wire w_dff_B_dQXVGhtG9_2;
	wire w_dff_B_d6NWEL8l7_2;
	wire w_dff_B_qtRC3AJQ5_2;
	wire w_dff_B_xPABRAl62_2;
	wire w_dff_B_004D1zQR1_2;
	wire w_dff_B_sZxMmARE0_2;
	wire w_dff_B_mDvlIhhp8_2;
	wire w_dff_B_NItKVYYn2_2;
	wire w_dff_B_rj8huoSf4_2;
	wire w_dff_B_blTyxex25_2;
	wire w_dff_B_yCObGZKb5_2;
	wire w_dff_B_mWNBCjqY6_2;
	wire w_dff_B_XqvcoNFE0_2;
	wire w_dff_B_s3P77hdo3_2;
	wire w_dff_B_hW4utQGO1_2;
	wire w_dff_B_7I4Blpxa0_2;
	wire w_dff_B_L1lMMz1t6_2;
	wire w_dff_B_TUzQBg6C0_2;
	wire w_dff_B_og15hhse0_1;
	wire w_dff_B_NTBdzeu70_2;
	wire w_dff_B_o8lAKN3h5_2;
	wire w_dff_B_0JO8cvJI1_2;
	wire w_dff_B_apTJhYpV8_2;
	wire w_dff_B_rgKonn0v0_2;
	wire w_dff_B_fApqZ5Nf5_2;
	wire w_dff_B_qOp703cz8_2;
	wire w_dff_B_ylc0NLGw3_2;
	wire w_dff_B_IIPZQFjA2_2;
	wire w_dff_B_I3Y7cDo83_2;
	wire w_dff_B_JEheRk3y4_2;
	wire w_dff_B_MNdHRZgK1_2;
	wire w_dff_B_HuO5DTko5_2;
	wire w_dff_B_5byUhrvB8_2;
	wire w_dff_B_TGNBIzIj4_2;
	wire w_dff_B_iNOV77LL4_2;
	wire w_dff_B_8OHwCIHs5_2;
	wire w_dff_B_TXHiw2xj9_2;
	wire w_dff_B_C2tPhRZm2_2;
	wire w_dff_B_I2zCEZrO8_1;
	wire w_dff_B_3GSWQHF03_2;
	wire w_dff_B_WzhtIyi69_2;
	wire w_dff_B_KNNWknm91_2;
	wire w_dff_B_zXi14C1v5_2;
	wire w_dff_B_u93RiUpC9_2;
	wire w_dff_B_DYSMGqam8_2;
	wire w_dff_B_pYaZClYR5_2;
	wire w_dff_B_lmerLkGA4_2;
	wire w_dff_B_hsQramjb0_2;
	wire w_dff_B_ehVgmDyt9_2;
	wire w_dff_B_GvKI84w06_2;
	wire w_dff_B_33xAjp1R9_2;
	wire w_dff_B_EQnXRH0y8_2;
	wire w_dff_B_I8zPB7qr6_2;
	wire w_dff_B_e9sc4Qcq2_2;
	wire w_dff_B_3AHQoFUj2_2;
	wire w_dff_B_AAYbOxiG6_1;
	wire w_dff_B_9BcOlL2r4_2;
	wire w_dff_B_G7qarGdR7_2;
	wire w_dff_B_EIgsg5sb1_2;
	wire w_dff_B_eouyq3bX3_2;
	wire w_dff_B_BmKJk8Qk9_2;
	wire w_dff_B_16jA1Ug15_2;
	wire w_dff_B_wTA4GIow3_2;
	wire w_dff_B_VycL0m8f3_2;
	wire w_dff_B_hmV5wMXC0_2;
	wire w_dff_B_SiwSrSmM3_2;
	wire w_dff_B_gxMSgUNz3_2;
	wire w_dff_B_1XoMUMZI6_2;
	wire w_dff_B_3ZxVpABO3_2;
	wire w_dff_B_Lv9VvjLv5_1;
	wire w_dff_B_cUdok9yr9_2;
	wire w_dff_B_sxjP9MWd4_2;
	wire w_dff_B_e4GuuxXM5_2;
	wire w_dff_B_hcW5uvqd2_2;
	wire w_dff_B_nxG1Sv2Z9_2;
	wire w_dff_B_Lx6rwnjp9_2;
	wire w_dff_B_uImVwb7e6_2;
	wire w_dff_B_mD5yxOv23_2;
	wire w_dff_B_aiLqEprQ5_2;
	wire w_dff_B_k4hePdx60_2;
	wire w_dff_B_2FQMyY2l4_2;
	wire w_dff_B_kqE9i7Nb1_1;
	wire w_dff_B_e5UcNpW79_1;
	wire w_dff_B_uhZNfmV57_1;
	wire w_dff_B_yUGuLAXp2_1;
	wire w_dff_B_jAyon4UW6_1;
	wire w_dff_B_bUtnm8xz7_1;
	wire w_dff_B_jTeyabpQ6_0;
	wire w_dff_B_BR1rDjUz4_0;
	wire w_dff_A_v4WlWYID6_0;
	wire w_dff_A_j08K9JPj0_0;
	wire w_dff_A_FLv3uGPk2_0;
	wire w_dff_B_O5bHpvuc3_1;
	wire w_dff_A_B9LfuwoA9_0;
	wire w_dff_A_8Or30avU8_1;
	wire w_dff_A_KPFWeGym0_1;
	wire w_dff_A_nWoJEuQb5_1;
	wire w_dff_A_fmU5U7Rz6_1;
	wire w_dff_A_7n3N5W964_1;
	wire w_dff_A_tLR7lvQq3_1;
	wire w_dff_A_YQ3K9KNn2_1;
	wire w_dff_A_fhhOmcMR1_1;
	wire w_dff_B_e7rQmgAM9_1;
	wire w_dff_A_KDTpLwao3_1;
	wire w_dff_B_2R8ssFfu8_1;
	wire w_dff_B_4iEGNX4k6_2;
	wire w_dff_B_bkqm7Fyg4_2;
	wire w_dff_B_Asz62aTZ5_2;
	wire w_dff_B_KWL87JfM9_2;
	wire w_dff_B_g0ZBFLtY1_2;
	wire w_dff_B_oP6nXBda2_2;
	wire w_dff_B_hch7V9117_2;
	wire w_dff_B_nZY7GlY08_2;
	wire w_dff_B_VwdoIWdU2_2;
	wire w_dff_B_yz6C6NLB2_2;
	wire w_dff_B_XoeOYaGt0_2;
	wire w_dff_B_e87aAuAG6_2;
	wire w_dff_B_WbPBm8bm5_2;
	wire w_dff_B_9mvFTDlZ6_2;
	wire w_dff_B_TnF7dwqv5_2;
	wire w_dff_B_9vMO3mb44_2;
	wire w_dff_B_xfAlWrTt6_2;
	wire w_dff_B_iKcIK2D28_2;
	wire w_dff_B_EtPQ2LJz7_2;
	wire w_dff_B_iedRFMJC1_2;
	wire w_dff_B_fhj2ej8M5_2;
	wire w_dff_B_UNn6pOEv9_2;
	wire w_dff_B_nJQaEDV28_2;
	wire w_dff_B_iL0B8Hav0_2;
	wire w_dff_B_bbmwxhks0_2;
	wire w_dff_B_1Yc9nh9s0_2;
	wire w_dff_B_8cqLZpNH1_2;
	wire w_dff_B_cI5Fv32S6_2;
	wire w_dff_B_GoHKKvWu2_2;
	wire w_dff_B_tBnbRVxq3_2;
	wire w_dff_B_jYejXZNb8_2;
	wire w_dff_B_WYnXZsUE5_2;
	wire w_dff_B_KfJcRmMU6_2;
	wire w_dff_B_Q6oF7kVo0_2;
	wire w_dff_B_6i1qVTkJ0_2;
	wire w_dff_B_lEKhbbch0_2;
	wire w_dff_B_9CUcbquI8_2;
	wire w_dff_B_76qYG72q0_2;
	wire w_dff_B_8LbPNQOY7_2;
	wire w_dff_B_phyzLvqW6_2;
	wire w_dff_B_AXkeI9wH9_2;
	wire w_dff_B_wWFUPvyS6_2;
	wire w_dff_B_al3nY6R34_2;
	wire w_dff_B_d02Ejx0N3_2;
	wire w_dff_B_JqS5l66B8_2;
	wire w_dff_B_MJeIncJl2_2;
	wire w_dff_B_3RPeXNwE6_2;
	wire w_dff_B_BKXFm4qV6_2;
	wire w_dff_B_eRWRvYFs0_2;
	wire w_dff_B_vidOmM8E0_2;
	wire w_dff_B_6E1WzGAH5_1;
	wire w_dff_B_GMXVFmo87_2;
	wire w_dff_B_VhYiU9p90_2;
	wire w_dff_B_7VmPgVOa7_2;
	wire w_dff_B_UBk9Vfuf4_2;
	wire w_dff_B_z95ndv0s8_2;
	wire w_dff_B_Gj9vx9kH3_2;
	wire w_dff_B_HHglZIgO7_2;
	wire w_dff_B_WmX87N4j8_2;
	wire w_dff_B_aCjEWD9j5_2;
	wire w_dff_B_M0JZtGP57_2;
	wire w_dff_B_ID2B8IpB5_2;
	wire w_dff_B_X9mdq5Y74_2;
	wire w_dff_B_rVSyZLor2_2;
	wire w_dff_B_WPn96d4Q4_2;
	wire w_dff_B_Z71cg9912_2;
	wire w_dff_B_ggK1QwuK4_2;
	wire w_dff_B_q9RypAz71_2;
	wire w_dff_B_D8UPfHhv9_2;
	wire w_dff_B_f6zRBvxY1_2;
	wire w_dff_B_V8j1UlyI1_2;
	wire w_dff_B_2C6bwF0m4_2;
	wire w_dff_B_nmDxdhXZ6_2;
	wire w_dff_B_n5eS17F55_2;
	wire w_dff_B_LVAZMxIP2_2;
	wire w_dff_B_LXhgr5xo7_2;
	wire w_dff_B_kWigknG92_2;
	wire w_dff_B_7gnDFMqR8_2;
	wire w_dff_B_Yw4uZofs5_2;
	wire w_dff_B_qQ3UMM6B4_2;
	wire w_dff_B_lpDWz5xn2_2;
	wire w_dff_B_A2nZeAre6_2;
	wire w_dff_B_PKbWz6PF5_2;
	wire w_dff_B_DHZPbG821_2;
	wire w_dff_B_KSbdqQjN2_2;
	wire w_dff_B_beORuMVy1_2;
	wire w_dff_B_R7JfVrcH7_2;
	wire w_dff_B_GI5B6ONl5_2;
	wire w_dff_B_ntopK4Fq5_2;
	wire w_dff_B_lNBBb5Mf1_2;
	wire w_dff_B_tkZPKKnO0_2;
	wire w_dff_B_AGe4Ytyv9_2;
	wire w_dff_B_7gf4WLNu5_2;
	wire w_dff_B_N4mBQkgr0_2;
	wire w_dff_B_CzETjaGO4_2;
	wire w_dff_B_oltETmjT9_2;
	wire w_dff_B_dpZfKvVX0_2;
	wire w_dff_B_QKibgKDa8_1;
	wire w_dff_B_1s5tCjko0_2;
	wire w_dff_B_0cI17qcD8_2;
	wire w_dff_B_58pf3EQF6_2;
	wire w_dff_B_8IaurN1Q8_2;
	wire w_dff_B_km3FnPFm5_2;
	wire w_dff_B_y6yZ3j9W2_2;
	wire w_dff_B_gocjZram1_2;
	wire w_dff_B_1IGagMmn9_2;
	wire w_dff_B_BoHTvwfo6_2;
	wire w_dff_B_uqe3gkPo4_2;
	wire w_dff_B_wyfTh3fA1_2;
	wire w_dff_B_ItWn1yZr3_2;
	wire w_dff_B_rGeIIq0s7_2;
	wire w_dff_B_liAHa5p55_2;
	wire w_dff_B_1DOurXRH0_2;
	wire w_dff_B_tuA5QtV19_2;
	wire w_dff_B_NpocvfLw3_2;
	wire w_dff_B_TmzCbW5E0_2;
	wire w_dff_B_voIYm9O80_2;
	wire w_dff_B_9RW5tuQa4_2;
	wire w_dff_B_2qZB7d1W7_2;
	wire w_dff_B_oFQGmyHB9_2;
	wire w_dff_B_MleDO6jT0_2;
	wire w_dff_B_TjcQ3fL30_2;
	wire w_dff_B_iZRbspGT7_2;
	wire w_dff_B_d0tsRWLF2_2;
	wire w_dff_B_jUZ15Anr9_2;
	wire w_dff_B_pyT6AlUX6_2;
	wire w_dff_B_mNHUaxJS4_2;
	wire w_dff_B_NSULHQX49_2;
	wire w_dff_B_OJuYZUPj1_2;
	wire w_dff_B_2CPpwImG4_2;
	wire w_dff_B_R4gpfeSf6_2;
	wire w_dff_B_OE06QjU20_2;
	wire w_dff_B_GJgtE1tx4_2;
	wire w_dff_B_EQnZijLD5_2;
	wire w_dff_B_grvRkOlY1_2;
	wire w_dff_B_FOsTG4KS8_2;
	wire w_dff_B_Uu4Xc0fB8_2;
	wire w_dff_B_bVmSKT6a5_2;
	wire w_dff_B_gEEO3E7I5_2;
	wire w_dff_B_cPxo96Ll1_2;
	wire w_dff_B_T6U1i5sD6_1;
	wire w_dff_B_97QZtcbo8_2;
	wire w_dff_B_c8yOQlVH8_2;
	wire w_dff_B_jX9lxqyI9_2;
	wire w_dff_B_r0VF3OLf9_2;
	wire w_dff_B_tFA5BSjr3_2;
	wire w_dff_B_uA5NaYnK9_2;
	wire w_dff_B_Jk9CC1OT6_2;
	wire w_dff_B_F7eTZm5u2_2;
	wire w_dff_B_ic8D8o6W3_2;
	wire w_dff_B_GSgUbhqP6_2;
	wire w_dff_B_BoKDD3bt7_2;
	wire w_dff_B_LWAtVUJ64_2;
	wire w_dff_B_RR532V0c8_2;
	wire w_dff_B_tXPXIhhT1_2;
	wire w_dff_B_QWD7vBpy0_2;
	wire w_dff_B_AyJpJwkY8_2;
	wire w_dff_B_Iv6ujFZS5_2;
	wire w_dff_B_bRWMaYzq4_2;
	wire w_dff_B_8HPVWGUP1_2;
	wire w_dff_B_3Horefdt7_2;
	wire w_dff_B_AOXHcnsf1_2;
	wire w_dff_B_Us2NEt0j0_2;
	wire w_dff_B_IKAzVBRv4_2;
	wire w_dff_B_HwS2VOr40_2;
	wire w_dff_B_WSNp20hW8_2;
	wire w_dff_B_bYZ5SP0d3_2;
	wire w_dff_B_vLE5msUt3_2;
	wire w_dff_B_nhQYtNyl6_2;
	wire w_dff_B_1W8p3sVY5_2;
	wire w_dff_B_cvQ4GP5F6_2;
	wire w_dff_B_4I6nkLkQ3_2;
	wire w_dff_B_Jej9mtvo4_2;
	wire w_dff_B_41G6egtG0_2;
	wire w_dff_B_b7RFWKmF2_2;
	wire w_dff_B_NtiGoyX29_2;
	wire w_dff_B_mJ5yHz6i7_2;
	wire w_dff_B_64mFQgHf1_2;
	wire w_dff_B_a5IKWAgM2_2;
	wire w_dff_B_yhcxjPXC0_1;
	wire w_dff_B_pFIWHQes1_2;
	wire w_dff_B_GotnhCGT2_2;
	wire w_dff_B_LTlYs43I3_2;
	wire w_dff_B_RHS81jZB5_2;
	wire w_dff_B_S3RJH4Ws2_2;
	wire w_dff_B_Tm3D5mPt7_2;
	wire w_dff_B_WE3qqVPP9_2;
	wire w_dff_B_uxT1D6338_2;
	wire w_dff_B_jMx5779a0_2;
	wire w_dff_B_v2xwKHeb4_2;
	wire w_dff_B_9jKtpsFI6_2;
	wire w_dff_B_htM14mEC7_2;
	wire w_dff_B_n9F98El57_2;
	wire w_dff_B_xoMEQcR57_2;
	wire w_dff_B_WNos43pr2_2;
	wire w_dff_B_Mh1PnJ7f7_2;
	wire w_dff_B_RpQVY65J4_2;
	wire w_dff_B_93VvMLb58_2;
	wire w_dff_B_ZQYaCXxO8_2;
	wire w_dff_B_t3EzFkF37_2;
	wire w_dff_B_K25tA2PS5_2;
	wire w_dff_B_zWRsC3bq5_2;
	wire w_dff_B_7cyJ4ttE1_2;
	wire w_dff_B_d0ojW1mo2_2;
	wire w_dff_B_w4yjCdvI7_2;
	wire w_dff_B_6c103qEE8_2;
	wire w_dff_B_Hmw166ZA9_2;
	wire w_dff_B_Q768gosW6_2;
	wire w_dff_B_bxhmf6Jn1_2;
	wire w_dff_B_mR8i586u6_2;
	wire w_dff_B_hbex8qap6_2;
	wire w_dff_B_4AVorcFG1_2;
	wire w_dff_B_eriIFOdA8_2;
	wire w_dff_B_ZYR8bUcq9_1;
	wire w_dff_B_4ssvc3ki2_2;
	wire w_dff_B_kDp4w20w5_2;
	wire w_dff_B_rbm0nJuE1_2;
	wire w_dff_B_CRhPGjLx1_2;
	wire w_dff_B_VR0TY0En9_2;
	wire w_dff_B_w7067A6k8_2;
	wire w_dff_B_ublLwUk06_2;
	wire w_dff_B_ONZshlIA3_2;
	wire w_dff_B_vS4z9xBE7_2;
	wire w_dff_B_RZGrnvTw7_2;
	wire w_dff_B_4LIAl3iU5_2;
	wire w_dff_B_iVirvHAg5_2;
	wire w_dff_B_tZsvH4Io2_2;
	wire w_dff_B_9ucynOSd9_2;
	wire w_dff_B_N5DiDxSP7_2;
	wire w_dff_B_5BWeoAYm9_2;
	wire w_dff_B_ZHtrGXRZ0_2;
	wire w_dff_B_hIsLXNHo6_2;
	wire w_dff_B_Vh3Zg9Df7_2;
	wire w_dff_B_CLMI8uF79_2;
	wire w_dff_B_L1Qd1uLb3_2;
	wire w_dff_B_IQcUPQV88_2;
	wire w_dff_B_bpggpXnK0_2;
	wire w_dff_B_yfeROOuA0_2;
	wire w_dff_B_gn6fMtlZ4_2;
	wire w_dff_B_KvxMmyCb4_2;
	wire w_dff_B_sOps9xw27_2;
	wire w_dff_B_q8M89MVA6_2;
	wire w_dff_B_9btL855A4_2;
	wire w_dff_B_7yT6s86O9_2;
	wire w_dff_B_N7HFNmL51_2;
	wire w_dff_B_3PqYq3sP3_1;
	wire w_dff_B_OtXlyWkF9_2;
	wire w_dff_B_MZJd5AlY4_2;
	wire w_dff_B_qM1O2MMg5_2;
	wire w_dff_B_XL6K4SKI0_2;
	wire w_dff_B_nPak7Bnr0_2;
	wire w_dff_B_6CFPvWJB5_2;
	wire w_dff_B_iVhXdDKL5_2;
	wire w_dff_B_K7NKydnj0_2;
	wire w_dff_B_AGFIL2cr7_2;
	wire w_dff_B_WUVTxoag8_2;
	wire w_dff_B_Qmh1s1rS4_2;
	wire w_dff_B_hhUp20oT9_2;
	wire w_dff_B_SjsIbhE67_2;
	wire w_dff_B_0RFOmsFX8_2;
	wire w_dff_B_vYHVJ21a4_2;
	wire w_dff_B_iWxfl3AW9_2;
	wire w_dff_B_noptbPDu7_2;
	wire w_dff_B_lAevw6P08_2;
	wire w_dff_B_ERzJiIhE7_2;
	wire w_dff_B_b1fEkFM42_2;
	wire w_dff_B_jqWeuXVU8_2;
	wire w_dff_B_xNkw5Xi87_2;
	wire w_dff_B_aZQysVSF8_2;
	wire w_dff_B_N9BdXA5F1_2;
	wire w_dff_B_cIzcRSxX1_2;
	wire w_dff_B_qAVhMp1z9_2;
	wire w_dff_B_rCZSACc71_2;
	wire w_dff_B_JzaWxUPK5_2;
	wire w_dff_B_GEWdfR901_1;
	wire w_dff_B_NjmbRh5y1_2;
	wire w_dff_B_3TUKA2cL3_2;
	wire w_dff_B_tQRABHbm6_2;
	wire w_dff_B_TWULv2pj6_2;
	wire w_dff_B_Zlz2yOhk7_2;
	wire w_dff_B_v6HjMCBG8_2;
	wire w_dff_B_AgvHnm2u6_2;
	wire w_dff_B_K0LGHv5S3_2;
	wire w_dff_B_tfnngBfj8_2;
	wire w_dff_B_FZfGiIqE5_2;
	wire w_dff_B_H9JVhHAc0_2;
	wire w_dff_B_MHKDtimG9_2;
	wire w_dff_B_59xidWHp8_2;
	wire w_dff_B_zIisVie89_2;
	wire w_dff_B_WmJUN1np3_2;
	wire w_dff_B_WgULM6H93_2;
	wire w_dff_B_fedn4pvG9_2;
	wire w_dff_B_BOXrLKuW2_2;
	wire w_dff_B_uvlFfCrR9_2;
	wire w_dff_B_gSqHp4Qn3_2;
	wire w_dff_B_9tzzqx2D9_2;
	wire w_dff_B_PfRVapns3_2;
	wire w_dff_B_QBrN1hbE8_2;
	wire w_dff_B_OX7pxmD05_2;
	wire w_dff_B_D9ufeY0w9_2;
	wire w_dff_B_OGayP6UF0_1;
	wire w_dff_B_pPoq0s3E5_2;
	wire w_dff_B_7YDyOhI02_2;
	wire w_dff_B_Mgyzczwn7_2;
	wire w_dff_B_WptxvJo90_2;
	wire w_dff_B_Z5oEdZZJ9_2;
	wire w_dff_B_CiRB4mgs6_2;
	wire w_dff_B_UyNeCXGl9_2;
	wire w_dff_B_LQ7cMm0f9_2;
	wire w_dff_B_CGHJPGSj3_2;
	wire w_dff_B_mhRCrGfW5_2;
	wire w_dff_B_3nlWnsGa8_2;
	wire w_dff_B_Pkf2jpEu2_2;
	wire w_dff_B_Y4zq1sGt3_2;
	wire w_dff_B_Yw5WNjbN2_2;
	wire w_dff_B_TtLTdCew5_2;
	wire w_dff_B_2I0LAd8o8_2;
	wire w_dff_B_5wyvDAza6_2;
	wire w_dff_B_CASYQ0eH7_2;
	wire w_dff_B_5WBTIYFa4_2;
	wire w_dff_B_BxoRNNht1_2;
	wire w_dff_B_7bZcCXZS1_2;
	wire w_dff_B_GbmpGLAX9_2;
	wire w_dff_B_gCRseKSX3_1;
	wire w_dff_B_mlDj4PGA0_2;
	wire w_dff_B_60JDDtxq8_2;
	wire w_dff_B_dXKPNGaB6_2;
	wire w_dff_B_BcmT4in45_2;
	wire w_dff_B_nXsgOr2e6_2;
	wire w_dff_B_b3xcDoic3_2;
	wire w_dff_B_85kXD39g6_2;
	wire w_dff_B_TDjDuefu0_2;
	wire w_dff_B_GkPCBVRA0_2;
	wire w_dff_B_k7XBf9yh1_2;
	wire w_dff_B_KLP56cjr7_2;
	wire w_dff_B_QoIdJcCd5_2;
	wire w_dff_B_d6bmIbUv2_2;
	wire w_dff_B_mqnz2Oec4_2;
	wire w_dff_B_NczUmfie4_2;
	wire w_dff_B_ScNqzfOL9_2;
	wire w_dff_B_4mkaHuoa0_2;
	wire w_dff_B_SYNboMum6_2;
	wire w_dff_B_xixEthtw6_2;
	wire w_dff_B_qeu9lj3P5_1;
	wire w_dff_B_HmnumnpZ7_2;
	wire w_dff_B_sOrVGgvY5_2;
	wire w_dff_B_iEXFjpRo6_2;
	wire w_dff_B_2GYSVV2G5_2;
	wire w_dff_B_eojb1KFr7_2;
	wire w_dff_B_w2CaxaxL6_2;
	wire w_dff_B_fvZqbBQc7_2;
	wire w_dff_B_4pObe9bz1_2;
	wire w_dff_B_yyPU1AZ42_2;
	wire w_dff_B_rDT0YzAj1_2;
	wire w_dff_B_3nyNm6ik4_2;
	wire w_dff_B_4VG4T8j56_2;
	wire w_dff_B_oDQCTvP72_2;
	wire w_dff_B_jN30JHwD0_2;
	wire w_dff_B_hZonOQGc3_2;
	wire w_dff_B_VPqAJya48_2;
	wire w_dff_B_mzUSu3Sl6_1;
	wire w_dff_B_U2zLMTSV7_2;
	wire w_dff_B_FKFziUga8_2;
	wire w_dff_B_VB0madkY1_2;
	wire w_dff_B_ndr0xpYE1_2;
	wire w_dff_B_esdRrUru9_2;
	wire w_dff_B_LaW8pPi32_2;
	wire w_dff_B_R5w4YP2I5_2;
	wire w_dff_B_cbGvOLHq5_2;
	wire w_dff_B_NcjOMpo80_2;
	wire w_dff_B_rJhexsno1_2;
	wire w_dff_B_lFlZ85i59_2;
	wire w_dff_B_qZbZfeDP3_2;
	wire w_dff_B_fwDr6czM6_2;
	wire w_dff_B_5vWzdcRT7_1;
	wire w_dff_B_8LTdD9Av0_2;
	wire w_dff_B_az2n5Dvx8_2;
	wire w_dff_B_hLCyo4IY1_2;
	wire w_dff_B_KTHieP3o9_2;
	wire w_dff_B_QJRV6pjR8_2;
	wire w_dff_B_vYcwUBYG0_2;
	wire w_dff_B_zp5mS1ME4_2;
	wire w_dff_B_dVTQh3y36_2;
	wire w_dff_B_kW0xO70A7_2;
	wire w_dff_B_Yft6KHAR0_2;
	wire w_dff_B_Q9usjkEE9_2;
	wire w_dff_B_uDBHMAkV3_1;
	wire w_dff_B_hw5kRXTC8_1;
	wire w_dff_B_xZ9luDGZ0_1;
	wire w_dff_B_p6Xw8KO09_1;
	wire w_dff_B_iU6lThHJ5_1;
	wire w_dff_B_zSBRfi7M7_1;
	wire w_dff_B_HDVF1MKI9_0;
	wire w_dff_B_EekNaYkb0_0;
	wire w_dff_A_N1glNa8a6_0;
	wire w_dff_A_XdFrbmsi7_0;
	wire w_dff_A_uWveNDfc0_0;
	wire w_dff_B_8Jm3I2aR8_1;
	wire w_dff_A_dGQ0nULC2_0;
	wire w_dff_A_KSL9U9ae5_1;
	wire w_dff_A_KSo3umKP5_1;
	wire w_dff_A_Kw2ZnM0o7_1;
	wire w_dff_A_dpJ3ydDa4_1;
	wire w_dff_A_u14aLw1x1_1;
	wire w_dff_A_8HGtWYyN0_1;
	wire w_dff_A_XiL1B0KF5_1;
	wire w_dff_A_zum0rnsQ5_1;
	wire w_dff_B_r5DeWLnr2_1;
	wire w_dff_A_NXdfcoJP4_1;
	wire w_dff_B_GY0AmhZ59_1;
	wire w_dff_B_ePK80bvI7_2;
	wire w_dff_B_cCfugXea4_2;
	wire w_dff_B_HNzP4zuC9_2;
	wire w_dff_B_xLjwrGpg1_2;
	wire w_dff_B_nlfY0wlw1_2;
	wire w_dff_B_Pzt54vDd6_2;
	wire w_dff_B_x1sVaed98_2;
	wire w_dff_B_Ke4Ut6Fp8_2;
	wire w_dff_B_qfNMeWtP7_2;
	wire w_dff_B_fqWe8lct2_2;
	wire w_dff_B_CuW57XJU7_2;
	wire w_dff_B_o0dZ6yOj0_2;
	wire w_dff_B_Nay2pum26_2;
	wire w_dff_B_ANHQpEA33_2;
	wire w_dff_B_IbVan7kt7_2;
	wire w_dff_B_HDABYoca9_2;
	wire w_dff_B_I2vE2NPk8_2;
	wire w_dff_B_fZjbahRI0_2;
	wire w_dff_B_6EEMmO5J1_2;
	wire w_dff_B_NqDLBXqy3_2;
	wire w_dff_B_5iYD0Zbd8_2;
	wire w_dff_B_u0fiProG1_2;
	wire w_dff_B_i1p3lPvA3_2;
	wire w_dff_B_JxbbM03X2_2;
	wire w_dff_B_jjbOOJty0_2;
	wire w_dff_B_LLxWuUlF7_2;
	wire w_dff_B_DwzoH0JF1_2;
	wire w_dff_B_Ca5xTHUO0_2;
	wire w_dff_B_m5J8wfJ60_2;
	wire w_dff_B_iZnl4Rt58_2;
	wire w_dff_B_DGDq6EMk9_2;
	wire w_dff_B_hNRTvzt02_2;
	wire w_dff_B_31xG7Nmt6_2;
	wire w_dff_B_TQKvFGPy5_2;
	wire w_dff_B_KdSJ1KoX0_2;
	wire w_dff_B_PzXFJFzi7_2;
	wire w_dff_B_aGujVf8T0_2;
	wire w_dff_B_VoPYT5206_2;
	wire w_dff_B_ILRjO57R8_2;
	wire w_dff_B_pw6AlegW4_2;
	wire w_dff_B_tbcR3mhi0_2;
	wire w_dff_B_ocZ4SEGP9_2;
	wire w_dff_B_TKwQSZXY8_2;
	wire w_dff_B_MU1aIrer5_2;
	wire w_dff_B_d2o0mNql3_2;
	wire w_dff_B_NOHnhdVs3_2;
	wire w_dff_B_8q2A1Z6i4_2;
	wire w_dff_B_4ZrVkaSV6_2;
	wire w_dff_B_lJgWZslt3_2;
	wire w_dff_B_DUsgVNnI2_2;
	wire w_dff_B_9RcW6zgb1_2;
	wire w_dff_B_xqDSkUBz5_2;
	wire w_dff_B_gNgsEzPQ0_1;
	wire w_dff_B_UeJy3oBG9_2;
	wire w_dff_B_7S71IYYJ9_2;
	wire w_dff_B_RXNEyLjz0_2;
	wire w_dff_B_dvGNkrd43_2;
	wire w_dff_B_dIE8lYaJ6_2;
	wire w_dff_B_7zSgs2rL9_2;
	wire w_dff_B_AOYRtnH48_2;
	wire w_dff_B_xVlfDaRu6_2;
	wire w_dff_B_Q5Q2WDhV2_2;
	wire w_dff_B_IB18Sr8k6_2;
	wire w_dff_B_RofjhBv10_2;
	wire w_dff_B_Ejvc9xEw2_2;
	wire w_dff_B_mWE9sFZR3_2;
	wire w_dff_B_cYLcsKcj5_2;
	wire w_dff_B_6s16I7Nh2_2;
	wire w_dff_B_wLve7vrG2_2;
	wire w_dff_B_QpVrswoV0_2;
	wire w_dff_B_FvWZoqPa6_2;
	wire w_dff_B_PTLvPhbQ4_2;
	wire w_dff_B_6h3tks1C3_2;
	wire w_dff_B_6MDofNqx3_2;
	wire w_dff_B_lvbNRr7F0_2;
	wire w_dff_B_KhifAR572_2;
	wire w_dff_B_pKmY9tj21_2;
	wire w_dff_B_HDS0TLWb8_2;
	wire w_dff_B_SGCr3OSu3_2;
	wire w_dff_B_kZSg5kYB2_2;
	wire w_dff_B_bDech5iz6_2;
	wire w_dff_B_flcFECST9_2;
	wire w_dff_B_F7zz0rJa6_2;
	wire w_dff_B_oHMzqdI25_2;
	wire w_dff_B_zEyIqyRd9_2;
	wire w_dff_B_1LFhMdCH5_2;
	wire w_dff_B_udmTubbg5_2;
	wire w_dff_B_YLrErCGP1_2;
	wire w_dff_B_XJFTwsvg8_2;
	wire w_dff_B_qzN7AVFu1_2;
	wire w_dff_B_RHCQOPhW4_2;
	wire w_dff_B_4yo4dVHH8_2;
	wire w_dff_B_vSoP8dTC1_2;
	wire w_dff_B_3mftr2mb9_2;
	wire w_dff_B_uV4YDR5P6_2;
	wire w_dff_B_35pUyFmV2_2;
	wire w_dff_B_oE49qvc90_2;
	wire w_dff_B_HtFINoEQ4_2;
	wire w_dff_B_UJncnEO08_2;
	wire w_dff_B_r7iq2aZb3_2;
	wire w_dff_B_2HkC6nbC5_2;
	wire w_dff_B_1mu5OWs52_1;
	wire w_dff_B_fx9haq3O3_2;
	wire w_dff_B_YfMA7yYg6_2;
	wire w_dff_B_jztVFGoW9_2;
	wire w_dff_B_UtV1uj8u9_2;
	wire w_dff_B_ZebFH1Ax8_2;
	wire w_dff_B_G50801TZ8_2;
	wire w_dff_B_94tuSiRp4_2;
	wire w_dff_B_TIMERHmp5_2;
	wire w_dff_B_Echx574a5_2;
	wire w_dff_B_tRKm64bN8_2;
	wire w_dff_B_ajetV92m8_2;
	wire w_dff_B_5r6tFA737_2;
	wire w_dff_B_37MzKY7l3_2;
	wire w_dff_B_V51WLoZA6_2;
	wire w_dff_B_Bk0ZjsuH0_2;
	wire w_dff_B_vggDPlZB8_2;
	wire w_dff_B_jrMZqvoa6_2;
	wire w_dff_B_oZRJ3UTB2_2;
	wire w_dff_B_8n0VR7Yz7_2;
	wire w_dff_B_mLwm33GN1_2;
	wire w_dff_B_EN0qF3oE4_2;
	wire w_dff_B_rMNk3DzX1_2;
	wire w_dff_B_AF4cXdQd9_2;
	wire w_dff_B_XMVHqsc73_2;
	wire w_dff_B_z1VVwp4Y0_2;
	wire w_dff_B_IIYiEoRg0_2;
	wire w_dff_B_wb5hKJfC2_2;
	wire w_dff_B_3KyRdlSd7_2;
	wire w_dff_B_cEzJSqq35_2;
	wire w_dff_B_tiFV97GI2_2;
	wire w_dff_B_59BGuEmy0_2;
	wire w_dff_B_tWUDG0Vs2_2;
	wire w_dff_B_UiR0cI807_2;
	wire w_dff_B_08ESIBcq8_2;
	wire w_dff_B_vAIYuKNk3_2;
	wire w_dff_B_6AUDhgD76_2;
	wire w_dff_B_4vd5f4yR0_2;
	wire w_dff_B_oHs6fx5U7_2;
	wire w_dff_B_q7UVgjRl9_2;
	wire w_dff_B_aP3utOCb8_2;
	wire w_dff_B_IzhBC1Of2_2;
	wire w_dff_B_crzB92Gp2_2;
	wire w_dff_B_TbklrleN4_2;
	wire w_dff_B_wvGEp2xp2_2;
	wire w_dff_B_A4pjQGCK7_1;
	wire w_dff_B_FnXJUlif7_2;
	wire w_dff_B_u0Jv3aqi7_2;
	wire w_dff_B_b6lgS73J8_2;
	wire w_dff_B_AbhwuB7d4_2;
	wire w_dff_B_W11WnIzr4_2;
	wire w_dff_B_veHGK0tW9_2;
	wire w_dff_B_LCDF74L72_2;
	wire w_dff_B_dWltNYjq9_2;
	wire w_dff_B_3yihavyc2_2;
	wire w_dff_B_f7VucrrQ7_2;
	wire w_dff_B_dPb9Go098_2;
	wire w_dff_B_xsBvHCo94_2;
	wire w_dff_B_h0cos4mL5_2;
	wire w_dff_B_xIJW41TO3_2;
	wire w_dff_B_9rXEMFgp1_2;
	wire w_dff_B_ZxEWPVTO8_2;
	wire w_dff_B_46TE9PDf6_2;
	wire w_dff_B_kCQksZOY7_2;
	wire w_dff_B_yp6xNKAH8_2;
	wire w_dff_B_Iz8mMGtd4_2;
	wire w_dff_B_5CXB30p35_2;
	wire w_dff_B_WFpXvUFk3_2;
	wire w_dff_B_LsTKBciX4_2;
	wire w_dff_B_lxdCiglv5_2;
	wire w_dff_B_tUBomGYf4_2;
	wire w_dff_B_CDUf4V7V9_2;
	wire w_dff_B_xObiIz8G8_2;
	wire w_dff_B_xVzciGid0_2;
	wire w_dff_B_MU6FulMD7_2;
	wire w_dff_B_JNPVonrv8_2;
	wire w_dff_B_2bmkkxQE5_2;
	wire w_dff_B_oXNII3Wb9_2;
	wire w_dff_B_783TQtc27_2;
	wire w_dff_B_9fTZuK665_2;
	wire w_dff_B_CB8uP2Fw9_2;
	wire w_dff_B_1ldaiBDb7_2;
	wire w_dff_B_PkKDIW489_2;
	wire w_dff_B_02l0st186_2;
	wire w_dff_B_Vw0RU65l8_2;
	wire w_dff_B_V4twCLF92_2;
	wire w_dff_B_Z7ZDwvJ80_1;
	wire w_dff_B_woEOB4hB1_2;
	wire w_dff_B_mDLFQIFL5_2;
	wire w_dff_B_dJ6203jA6_2;
	wire w_dff_B_lKymu9Lv4_2;
	wire w_dff_B_JPkCIFal8_2;
	wire w_dff_B_DbfqoEeI1_2;
	wire w_dff_B_U91YbclF1_2;
	wire w_dff_B_fXLij1Mx7_2;
	wire w_dff_B_qOOmlspL1_2;
	wire w_dff_B_VlyAqOLq8_2;
	wire w_dff_B_rE80ocvs4_2;
	wire w_dff_B_RyLxkEpr5_2;
	wire w_dff_B_xfO8Phnw0_2;
	wire w_dff_B_tm6IjM5W7_2;
	wire w_dff_B_joA427e71_2;
	wire w_dff_B_jtNb9Dqs1_2;
	wire w_dff_B_d2Bicvdq8_2;
	wire w_dff_B_Xy2KueEx5_2;
	wire w_dff_B_p5eCBVpM5_2;
	wire w_dff_B_8r2l9ORy4_2;
	wire w_dff_B_899Nl0u35_2;
	wire w_dff_B_Xskf7ANf0_2;
	wire w_dff_B_srHJoi8r6_2;
	wire w_dff_B_XrxUk0ap3_2;
	wire w_dff_B_8tBkrL922_2;
	wire w_dff_B_bNnqb7Ur8_2;
	wire w_dff_B_dOpIcEEJ1_2;
	wire w_dff_B_3TquZD4L8_2;
	wire w_dff_B_uzVvRaG98_2;
	wire w_dff_B_I5PyVKJE5_2;
	wire w_dff_B_V4WBCfy56_2;
	wire w_dff_B_0PjtLUVy8_2;
	wire w_dff_B_ddjO5ckY1_2;
	wire w_dff_B_ULlziK0B4_2;
	wire w_dff_B_fKPvmQG84_2;
	wire w_dff_B_bkzLefRO7_2;
	wire w_dff_B_tB5h44mQ6_1;
	wire w_dff_B_Y6Lt9qFR1_2;
	wire w_dff_B_sdmIJJiy6_2;
	wire w_dff_B_e0JaXbkX8_2;
	wire w_dff_B_Z5IoM4KV9_2;
	wire w_dff_B_l7b6rMQt2_2;
	wire w_dff_B_VIi6iYqQ0_2;
	wire w_dff_B_eQM7WvpS7_2;
	wire w_dff_B_yFjIxuYn2_2;
	wire w_dff_B_uLFsrxjJ0_2;
	wire w_dff_B_Nzz2xrKI9_2;
	wire w_dff_B_rto4OUmf2_2;
	wire w_dff_B_LB06HmON2_2;
	wire w_dff_B_Ns69LjTy3_2;
	wire w_dff_B_g8BCCC211_2;
	wire w_dff_B_wbnkx0T13_2;
	wire w_dff_B_id3uFHpD0_2;
	wire w_dff_B_usQTZ7oR4_2;
	wire w_dff_B_c6cJmcVJ2_2;
	wire w_dff_B_EvwR6gro0_2;
	wire w_dff_B_HoIrTVtM7_2;
	wire w_dff_B_DKo8EdJc7_2;
	wire w_dff_B_7mOIfWiO7_2;
	wire w_dff_B_h6fDJDHS9_2;
	wire w_dff_B_m92kKJL86_2;
	wire w_dff_B_XgZGUoUN4_2;
	wire w_dff_B_OHfZSjCa0_2;
	wire w_dff_B_X5Dacjfa3_2;
	wire w_dff_B_DllvmJjb1_2;
	wire w_dff_B_GRzYs9UU0_2;
	wire w_dff_B_f0pfmsU71_2;
	wire w_dff_B_OaNem0ST0_2;
	wire w_dff_B_72E2VBGY8_2;
	wire w_dff_B_JqiJPZgx9_1;
	wire w_dff_B_wz2j3OsE3_2;
	wire w_dff_B_x6OCiYCV3_2;
	wire w_dff_B_XizDq3wQ9_2;
	wire w_dff_B_l7w4yQkK1_2;
	wire w_dff_B_7zhnYyxv2_2;
	wire w_dff_B_aF4DWmiM4_2;
	wire w_dff_B_N5k7GIlI5_2;
	wire w_dff_B_9cIQunZl8_2;
	wire w_dff_B_rB0COoHL2_2;
	wire w_dff_B_8Z5bNeUv2_2;
	wire w_dff_B_I2nQITPJ1_2;
	wire w_dff_B_62UScHEs7_2;
	wire w_dff_B_nC8ZqM5K7_2;
	wire w_dff_B_ZoLICgUo6_2;
	wire w_dff_B_YLU3kOcs8_2;
	wire w_dff_B_baOsjY5c2_2;
	wire w_dff_B_mxpmkjTt4_2;
	wire w_dff_B_ciZMMJGM1_2;
	wire w_dff_B_Q2LiyG181_2;
	wire w_dff_B_rOQXuXeo8_2;
	wire w_dff_B_9Bg31B148_2;
	wire w_dff_B_I2zr3lj56_2;
	wire w_dff_B_vskFeLij2_2;
	wire w_dff_B_Aq76FbGq0_2;
	wire w_dff_B_Eb4qjR1P0_2;
	wire w_dff_B_nRKGAYik5_2;
	wire w_dff_B_NOQOgkWw8_2;
	wire w_dff_B_PNvyRkvI3_1;
	wire w_dff_B_94zjszsN3_2;
	wire w_dff_B_Ah8ScVZB7_2;
	wire w_dff_B_WqqXRcvh2_2;
	wire w_dff_B_mRZXVqgv4_2;
	wire w_dff_B_Pwa2BY1K2_2;
	wire w_dff_B_eCPEyWZa9_2;
	wire w_dff_B_mE27JYPy5_2;
	wire w_dff_B_BWCfL8cj3_2;
	wire w_dff_B_W6MVfBXk8_2;
	wire w_dff_B_LPcYtsBO0_2;
	wire w_dff_B_77y0nqge2_2;
	wire w_dff_B_ZHHbx8e05_2;
	wire w_dff_B_YF3wRVRy4_2;
	wire w_dff_B_yOVIrUnP1_2;
	wire w_dff_B_VWrr8tZA1_2;
	wire w_dff_B_TDPBBekm7_2;
	wire w_dff_B_Kx6zWY4F7_2;
	wire w_dff_B_EdVhn0Ov9_2;
	wire w_dff_B_0PwMVtqr8_2;
	wire w_dff_B_oyyZiBef2_2;
	wire w_dff_B_i6g2mmxq3_2;
	wire w_dff_B_t4pLYhXH6_2;
	wire w_dff_B_b0JCdIFC3_2;
	wire w_dff_B_rYzcXI5W9_2;
	wire w_dff_B_4LcJR0th3_2;
	wire w_dff_B_sMQcSNB69_1;
	wire w_dff_B_qiWnmlq81_2;
	wire w_dff_B_h0j2oLgh8_2;
	wire w_dff_B_ZDT7n5Hv1_2;
	wire w_dff_B_RlYLjQvk9_2;
	wire w_dff_B_jJrQumHY0_2;
	wire w_dff_B_nZoprrbN3_2;
	wire w_dff_B_l2NmkNVe2_2;
	wire w_dff_B_rtNthS4D2_2;
	wire w_dff_B_SXe0O2YX3_2;
	wire w_dff_B_LIFYLMSx8_2;
	wire w_dff_B_BY7AOyL14_2;
	wire w_dff_B_nhyMnMBl7_2;
	wire w_dff_B_YSv1apY30_2;
	wire w_dff_B_h4kWvDaG6_2;
	wire w_dff_B_KORiv8Ni3_2;
	wire w_dff_B_ZO7wDaH22_2;
	wire w_dff_B_IwsFy9vA6_2;
	wire w_dff_B_3hAzUktV8_2;
	wire w_dff_B_BMwuPzhD5_2;
	wire w_dff_B_Veom8jI67_2;
	wire w_dff_B_m6wpOOTX3_2;
	wire w_dff_B_9cKVxRGY2_2;
	wire w_dff_B_pdx9xkB96_1;
	wire w_dff_B_VxD0nNwJ2_2;
	wire w_dff_B_BXTyLVDb1_2;
	wire w_dff_B_haLYPqUp7_2;
	wire w_dff_B_ebf72IZ39_2;
	wire w_dff_B_nJzcCgIt2_2;
	wire w_dff_B_2l3WI0sp5_2;
	wire w_dff_B_Y4OTmPUh0_2;
	wire w_dff_B_xKW4vRda4_2;
	wire w_dff_B_CR9zV5al8_2;
	wire w_dff_B_s7EP1w689_2;
	wire w_dff_B_M51abpuQ7_2;
	wire w_dff_B_eIwrQVmt6_2;
	wire w_dff_B_NGhfny2I7_2;
	wire w_dff_B_bx12cM4l8_2;
	wire w_dff_B_w7SSzkEF1_2;
	wire w_dff_B_ylhBoDkU3_2;
	wire w_dff_B_XUlRkKmS3_2;
	wire w_dff_B_79Wcx5u26_2;
	wire w_dff_B_MqZfHPqe4_2;
	wire w_dff_B_qDrVah190_1;
	wire w_dff_B_bBHxkFfT2_2;
	wire w_dff_B_wqTWrfma3_2;
	wire w_dff_B_SJt05p5r3_2;
	wire w_dff_B_NumCiepD9_2;
	wire w_dff_B_Ig6YHL9A9_2;
	wire w_dff_B_iUJjc4pH5_2;
	wire w_dff_B_lmYmd38Z4_2;
	wire w_dff_B_Jjln5ErG9_2;
	wire w_dff_B_1OhHQiec1_2;
	wire w_dff_B_UldrICCv1_2;
	wire w_dff_B_RXC2QJlE3_2;
	wire w_dff_B_MBKh6QIq4_2;
	wire w_dff_B_Yz8IP7JI9_2;
	wire w_dff_B_bEmJq9Q26_2;
	wire w_dff_B_8iNnw4fd3_2;
	wire w_dff_B_dUlgKmam6_2;
	wire w_dff_B_OuzEvqxX7_1;
	wire w_dff_B_p575ndzE0_2;
	wire w_dff_B_4tIrRp6y3_2;
	wire w_dff_B_aJrelXs39_2;
	wire w_dff_B_yX0hV0zB7_2;
	wire w_dff_B_LLoECp1X8_2;
	wire w_dff_B_0TpDOiCf3_2;
	wire w_dff_B_8IhBZRR65_2;
	wire w_dff_B_blKFOxBF6_2;
	wire w_dff_B_QEGnW7u19_2;
	wire w_dff_B_L4wEvSvt2_2;
	wire w_dff_B_kweSgKqg4_2;
	wire w_dff_B_0l63gjYM2_2;
	wire w_dff_B_FMIx6HkA4_2;
	wire w_dff_B_Th5MwW257_1;
	wire w_dff_B_NcUp0Ci72_2;
	wire w_dff_B_c3TfShXe5_2;
	wire w_dff_B_fTBGaos44_2;
	wire w_dff_B_g2SpbvpB2_2;
	wire w_dff_B_OxVT2tcz6_2;
	wire w_dff_B_Rlhd1RZ53_2;
	wire w_dff_B_XFxrXvdU6_2;
	wire w_dff_B_0hucysWl5_2;
	wire w_dff_B_eylds8PW2_2;
	wire w_dff_B_r2tZCzxO0_2;
	wire w_dff_B_yseD4T131_2;
	wire w_dff_B_8UsONRXs4_1;
	wire w_dff_B_i5s3NL2W3_1;
	wire w_dff_B_UXBtV24U6_1;
	wire w_dff_B_yhLU7zb81_1;
	wire w_dff_B_z1IWhVkG5_1;
	wire w_dff_B_Z6o9Hakd3_1;
	wire w_dff_B_SJeyUxvo2_0;
	wire w_dff_B_wrk2j1G20_0;
	wire w_dff_A_MrsLvblf1_0;
	wire w_dff_A_R9Z5k56G0_0;
	wire w_dff_A_sw2PtKtX2_0;
	wire w_dff_B_2psNJ8Fq6_1;
	wire w_dff_A_vN8Ty6XF4_0;
	wire w_dff_A_Tru88F5E9_1;
	wire w_dff_A_srnRvMnm4_1;
	wire w_dff_A_z36lHbXL5_1;
	wire w_dff_A_Ib01DOzk8_1;
	wire w_dff_A_Ou5AVYtg3_1;
	wire w_dff_A_yDHm8PpD2_1;
	wire w_dff_A_F1pYYuP78_1;
	wire w_dff_A_04uEiypF3_1;
	wire w_dff_B_LOyfXsth5_1;
	wire w_dff_A_Hvb89mYh3_1;
	wire w_dff_B_mSbZR5nX4_1;
	wire w_dff_B_Ejj13FDg1_2;
	wire w_dff_B_umvEI9Vo6_2;
	wire w_dff_B_FUzfAqvL8_2;
	wire w_dff_B_ITm47nRE0_2;
	wire w_dff_B_IvY5Cxcl5_2;
	wire w_dff_B_xrEQa0iw9_2;
	wire w_dff_B_iB3dktwx3_2;
	wire w_dff_B_IcjrXihW5_2;
	wire w_dff_B_oCmQpDPh9_2;
	wire w_dff_B_j0oG0F0G4_2;
	wire w_dff_B_z8J6ruUG0_2;
	wire w_dff_B_pGJKsymL9_2;
	wire w_dff_B_L8IgM5Zy6_2;
	wire w_dff_B_8m2k3oyM8_2;
	wire w_dff_B_YwRopqfB3_2;
	wire w_dff_B_GEsXNV6y5_2;
	wire w_dff_B_p0xbA5Ai8_2;
	wire w_dff_B_q6XIlSm58_2;
	wire w_dff_B_Q5qOZsg61_2;
	wire w_dff_B_qh1sDJVQ2_2;
	wire w_dff_B_VuvW6dgs2_2;
	wire w_dff_B_IGKpHItS6_2;
	wire w_dff_B_cHEDTrUP0_2;
	wire w_dff_B_0YQkRkXF8_2;
	wire w_dff_B_Kj2OZhRL7_2;
	wire w_dff_B_OYx71PWU9_2;
	wire w_dff_B_V6KxGlsT4_2;
	wire w_dff_B_g9hd9jit8_2;
	wire w_dff_B_vXpvzYHM7_2;
	wire w_dff_B_UjGuASmA9_2;
	wire w_dff_B_WGXuEf7o3_2;
	wire w_dff_B_5nc5dami1_2;
	wire w_dff_B_lvsYMnRp1_2;
	wire w_dff_B_qWuLwY080_2;
	wire w_dff_B_oiOybrMn6_2;
	wire w_dff_B_r6KyqbrR0_2;
	wire w_dff_B_XnZgAs7f9_2;
	wire w_dff_B_NODFih3y9_2;
	wire w_dff_B_fLzc46Ce3_2;
	wire w_dff_B_42jNCee70_2;
	wire w_dff_B_yeWMj1072_2;
	wire w_dff_B_Aojw71c43_2;
	wire w_dff_B_mU5xv5Ij6_2;
	wire w_dff_B_srGj8NzH7_2;
	wire w_dff_B_4PXeIdUz4_2;
	wire w_dff_B_Ko9Gsvxi5_2;
	wire w_dff_B_wHB96kvt5_2;
	wire w_dff_B_ACndFeqS3_2;
	wire w_dff_B_ykurAHmU2_2;
	wire w_dff_B_fQEvWDZd2_2;
	wire w_dff_B_iwbOJypr8_2;
	wire w_dff_B_rXXBjKT04_2;
	wire w_dff_B_ZmG8bPWg0_2;
	wire w_dff_B_75PHjK6M9_2;
	wire w_dff_B_41ptGfqe8_1;
	wire w_dff_B_geUBvjFh7_2;
	wire w_dff_B_RZKNY6CS2_2;
	wire w_dff_B_pf1BbJ5J8_2;
	wire w_dff_B_EWnqIpaA8_2;
	wire w_dff_B_Li1A4bY65_2;
	wire w_dff_B_f6PjTMbV3_2;
	wire w_dff_B_0H3tDfsL7_2;
	wire w_dff_B_lwAyrWz72_2;
	wire w_dff_B_7HTn104q4_2;
	wire w_dff_B_z1vOFJ5q5_2;
	wire w_dff_B_WkGOZLW77_2;
	wire w_dff_B_BU0WOKZz5_2;
	wire w_dff_B_cyCdttq31_2;
	wire w_dff_B_m9MlvMKq4_2;
	wire w_dff_B_60oNfWN27_2;
	wire w_dff_B_XQV099jo4_2;
	wire w_dff_B_MHVfk0DL6_2;
	wire w_dff_B_Jnz2xk1V0_2;
	wire w_dff_B_41HSxumI2_2;
	wire w_dff_B_QhLlWjY38_2;
	wire w_dff_B_MqyGJm1L5_2;
	wire w_dff_B_r41UVl7Y9_2;
	wire w_dff_B_ELVGJrJk8_2;
	wire w_dff_B_e4tBWFxm6_2;
	wire w_dff_B_vPXOdMit6_2;
	wire w_dff_B_56FuqRwM2_2;
	wire w_dff_B_nIL7XCRY7_2;
	wire w_dff_B_SIZ9O1VG9_2;
	wire w_dff_B_k3WNy3345_2;
	wire w_dff_B_c75UBdPK7_2;
	wire w_dff_B_xmVdhNrQ0_2;
	wire w_dff_B_903JaLxB3_2;
	wire w_dff_B_0mrL5mLA8_2;
	wire w_dff_B_jYjJuIVq3_2;
	wire w_dff_B_g0jwsfyE0_2;
	wire w_dff_B_QFvel9269_2;
	wire w_dff_B_qogUaso08_2;
	wire w_dff_B_l8fT2krH8_2;
	wire w_dff_B_C7tR32BQ0_2;
	wire w_dff_B_76XomXZs9_2;
	wire w_dff_B_J0Ufhwpm7_2;
	wire w_dff_B_fTyxRqd77_2;
	wire w_dff_B_pj1VU2v43_2;
	wire w_dff_B_uHePrxfz2_2;
	wire w_dff_B_4r5AkvxC9_2;
	wire w_dff_B_U7wureC74_2;
	wire w_dff_B_gqDYvhZe3_2;
	wire w_dff_B_uF3q11ah9_2;
	wire w_dff_B_5oksoLxC0_2;
	wire w_dff_B_kfVdW4aC6_2;
	wire w_dff_B_gC3Rv0z41_1;
	wire w_dff_B_jT8LzB527_2;
	wire w_dff_B_W0ZmB8Ho4_2;
	wire w_dff_B_AmiSepg94_2;
	wire w_dff_B_3fgl0hCo3_2;
	wire w_dff_B_Qc5DzA5Q8_2;
	wire w_dff_B_sW3pWa7H3_2;
	wire w_dff_B_FJblDYcg0_2;
	wire w_dff_B_bIPXvJRG1_2;
	wire w_dff_B_gsznbvZ46_2;
	wire w_dff_B_5Fihdx7n4_2;
	wire w_dff_B_i0yZvowo8_2;
	wire w_dff_B_eWz0jVWp9_2;
	wire w_dff_B_ntf0nUQE3_2;
	wire w_dff_B_doikCE2z5_2;
	wire w_dff_B_ipaRpm2w1_2;
	wire w_dff_B_yyjjj4Qy8_2;
	wire w_dff_B_swsjroU35_2;
	wire w_dff_B_XQVhgTYB8_2;
	wire w_dff_B_XMIeaaOw0_2;
	wire w_dff_B_c8b6EEaw5_2;
	wire w_dff_B_4WMR2ZzK2_2;
	wire w_dff_B_YvCy8vvI3_2;
	wire w_dff_B_NtPpTp807_2;
	wire w_dff_B_ulFXfwZm0_2;
	wire w_dff_B_HtplOrIW4_2;
	wire w_dff_B_l1DokOau1_2;
	wire w_dff_B_E4SZPomJ6_2;
	wire w_dff_B_s6U3UHmG4_2;
	wire w_dff_B_cGHYqfnb2_2;
	wire w_dff_B_TnAnl9QO9_2;
	wire w_dff_B_3gfV9m352_2;
	wire w_dff_B_s1tnnurs4_2;
	wire w_dff_B_7PwPP5Cm1_2;
	wire w_dff_B_2tQ9lGuU8_2;
	wire w_dff_B_QmzEqv8E2_2;
	wire w_dff_B_AS7lg4Kf4_2;
	wire w_dff_B_whwD1eTk2_2;
	wire w_dff_B_LDEa0inY4_2;
	wire w_dff_B_4VzBaOai2_2;
	wire w_dff_B_hd3L1nA42_2;
	wire w_dff_B_ijvmdrRa9_2;
	wire w_dff_B_xu4GHzgO6_2;
	wire w_dff_B_Ibm9RoZ63_2;
	wire w_dff_B_NXJungvK4_2;
	wire w_dff_B_BGuYp3u05_2;
	wire w_dff_B_7bx0Xb2Q0_2;
	wire w_dff_B_bCY77S658_1;
	wire w_dff_B_V6RJLTFs0_2;
	wire w_dff_B_h2jtc9p91_2;
	wire w_dff_B_3ltZOvc64_2;
	wire w_dff_B_7S3PMFjP1_2;
	wire w_dff_B_88fwvHQb1_2;
	wire w_dff_B_sbClGWUO8_2;
	wire w_dff_B_SISSsBgx5_2;
	wire w_dff_B_FMlXwUqq6_2;
	wire w_dff_B_Cj8FaT1T8_2;
	wire w_dff_B_92FFWy2l9_2;
	wire w_dff_B_ylJbDdbT2_2;
	wire w_dff_B_TFaJemOH3_2;
	wire w_dff_B_O6SJOrJG9_2;
	wire w_dff_B_vOmZ0eok6_2;
	wire w_dff_B_IscFfvsp6_2;
	wire w_dff_B_r8LAgrPk4_2;
	wire w_dff_B_qoeSUkIe6_2;
	wire w_dff_B_mfI2KR4f3_2;
	wire w_dff_B_VGU6obil9_2;
	wire w_dff_B_foXoIVQb9_2;
	wire w_dff_B_OEHadiIT7_2;
	wire w_dff_B_uv7ME0AH9_2;
	wire w_dff_B_gbScNmri3_2;
	wire w_dff_B_fGgc8efR3_2;
	wire w_dff_B_7wAcj6WB8_2;
	wire w_dff_B_0cocnuP30_2;
	wire w_dff_B_ZJQ4THPG5_2;
	wire w_dff_B_ZBK0Ce3x0_2;
	wire w_dff_B_V08ECaFc4_2;
	wire w_dff_B_rMaAlsfY6_2;
	wire w_dff_B_2bGgQ2qh5_2;
	wire w_dff_B_Xdt4naIX0_2;
	wire w_dff_B_p5vZOwmM8_2;
	wire w_dff_B_QCKbahQL3_2;
	wire w_dff_B_MGN1ipDK0_2;
	wire w_dff_B_H4YxNmQo7_2;
	wire w_dff_B_XkRIf8Hz2_2;
	wire w_dff_B_Mp2ifXT79_2;
	wire w_dff_B_MquMrvv39_2;
	wire w_dff_B_U0h6fLI23_2;
	wire w_dff_B_3rVbqRBO3_2;
	wire w_dff_B_hHfKE0vn2_2;
	wire w_dff_B_8uuf1NPF9_1;
	wire w_dff_B_8W0a4QFq5_2;
	wire w_dff_B_Zzr90bZu7_2;
	wire w_dff_B_oCpmkZgS4_2;
	wire w_dff_B_cSpuQyeN8_2;
	wire w_dff_B_czLHytWY8_2;
	wire w_dff_B_Od2bjCmf6_2;
	wire w_dff_B_y7pZWHVO9_2;
	wire w_dff_B_upvZbSKu0_2;
	wire w_dff_B_ajmSSkjV0_2;
	wire w_dff_B_G1OcHUp34_2;
	wire w_dff_B_8jcfrtjq0_2;
	wire w_dff_B_FdIi7iov8_2;
	wire w_dff_B_8dYf9r8b4_2;
	wire w_dff_B_kSqZamUx9_2;
	wire w_dff_B_a6ufy1Un4_2;
	wire w_dff_B_XmwejyP26_2;
	wire w_dff_B_rllJl9KP3_2;
	wire w_dff_B_G2fqfeIo8_2;
	wire w_dff_B_jKMgF7Qh3_2;
	wire w_dff_B_o1VfcBMx8_2;
	wire w_dff_B_gMCmfg1B0_2;
	wire w_dff_B_xlvvTZfE2_2;
	wire w_dff_B_BWvDlSpP4_2;
	wire w_dff_B_vVK2PL6q3_2;
	wire w_dff_B_TV50pzx35_2;
	wire w_dff_B_vhoxp4Az4_2;
	wire w_dff_B_wayJIXNz8_2;
	wire w_dff_B_K2Xhf19H5_2;
	wire w_dff_B_25U39w9H4_2;
	wire w_dff_B_Cus5OcBd0_2;
	wire w_dff_B_Q9jgfP202_2;
	wire w_dff_B_Dccwno3t9_2;
	wire w_dff_B_7Nhz5uH56_2;
	wire w_dff_B_UOCWkoL34_2;
	wire w_dff_B_aWQQDVVC9_2;
	wire w_dff_B_OGKro7M29_2;
	wire w_dff_B_uxlbT8043_2;
	wire w_dff_B_niD869Mu6_2;
	wire w_dff_B_AjoZInzR4_1;
	wire w_dff_B_pIjbyzw96_2;
	wire w_dff_B_n5eLjJz29_2;
	wire w_dff_B_tZuXqGTK5_2;
	wire w_dff_B_Ibq5R8j12_2;
	wire w_dff_B_Jvq2UC8s7_2;
	wire w_dff_B_Rt1K60Na5_2;
	wire w_dff_B_BkDZH8WR6_2;
	wire w_dff_B_tWaOV1KK1_2;
	wire w_dff_B_CJMzdSok6_2;
	wire w_dff_B_ztQmL6nz0_2;
	wire w_dff_B_9mqc3Ao92_2;
	wire w_dff_B_O3W17pQ15_2;
	wire w_dff_B_J4Zz7LsP4_2;
	wire w_dff_B_2KWcHWup0_2;
	wire w_dff_B_QUmbG9yf1_2;
	wire w_dff_B_hla1cY9Y8_2;
	wire w_dff_B_GEzHCmKz5_2;
	wire w_dff_B_auESlpph5_2;
	wire w_dff_B_4f3I6soJ2_2;
	wire w_dff_B_95CPVkjc1_2;
	wire w_dff_B_Lvfo8yf86_2;
	wire w_dff_B_GzjYyes91_2;
	wire w_dff_B_FEuV478o9_2;
	wire w_dff_B_0YoGJYha3_2;
	wire w_dff_B_a09rMzAG5_2;
	wire w_dff_B_EzDJem7c1_2;
	wire w_dff_B_wCBlYzyR4_2;
	wire w_dff_B_IzqOz8po1_2;
	wire w_dff_B_u9zubPfy8_2;
	wire w_dff_B_UtBZzhJt2_2;
	wire w_dff_B_n0ikSsPP2_2;
	wire w_dff_B_4GVukgXr0_2;
	wire w_dff_B_8pMa8pGJ1_2;
	wire w_dff_B_wZRVoe8d1_2;
	wire w_dff_B_CPSDcxeo0_1;
	wire w_dff_B_pkIXgoCW0_2;
	wire w_dff_B_qL122ReC9_2;
	wire w_dff_B_CEfFlcDu0_2;
	wire w_dff_B_OaUVFtHj8_2;
	wire w_dff_B_m5Xpi6ss2_2;
	wire w_dff_B_Gu7VTcKj0_2;
	wire w_dff_B_MmVG5Zm49_2;
	wire w_dff_B_SY2MVKr11_2;
	wire w_dff_B_SvmLfalu9_2;
	wire w_dff_B_DPx3AT5T9_2;
	wire w_dff_B_FhunLZ0A9_2;
	wire w_dff_B_D7zCsoZQ5_2;
	wire w_dff_B_6YSeV2Bq1_2;
	wire w_dff_B_WSKAjr3g2_2;
	wire w_dff_B_R7UFBQkP5_2;
	wire w_dff_B_r2PpmB2L5_2;
	wire w_dff_B_D4DvMUMe3_2;
	wire w_dff_B_bThkq4ZT6_2;
	wire w_dff_B_7giKRh5M5_2;
	wire w_dff_B_YVUhQyBk8_2;
	wire w_dff_B_JOFnZy7U4_2;
	wire w_dff_B_yjMxemBL2_2;
	wire w_dff_B_YQvke0zO7_2;
	wire w_dff_B_5iujL0oo1_2;
	wire w_dff_B_eE3jrWdx9_2;
	wire w_dff_B_J1uBbdG53_2;
	wire w_dff_B_kUxMpTmz3_2;
	wire w_dff_B_zzFGn0zt8_2;
	wire w_dff_B_PgDjnd6z1_2;
	wire w_dff_B_L7rgudxM0_2;
	wire w_dff_B_2eWKUzzW9_1;
	wire w_dff_B_91JATJxl9_2;
	wire w_dff_B_AQSNkDys5_2;
	wire w_dff_B_J3129anV8_2;
	wire w_dff_B_YYa7I4iS4_2;
	wire w_dff_B_RqZR2cBd7_2;
	wire w_dff_B_anPhin0E3_2;
	wire w_dff_B_Fi8zziLH7_2;
	wire w_dff_B_7YMmdHuy7_2;
	wire w_dff_B_oH0vbbef6_2;
	wire w_dff_B_XkDJSfbK4_2;
	wire w_dff_B_MlgJ31f45_2;
	wire w_dff_B_EUG5hBs56_2;
	wire w_dff_B_HjeZR5zt2_2;
	wire w_dff_B_tob1Cp0L5_2;
	wire w_dff_B_SSKae8cT4_2;
	wire w_dff_B_oKdZxUj41_2;
	wire w_dff_B_DjMOWeJy8_2;
	wire w_dff_B_XstjE5572_2;
	wire w_dff_B_SdX8df405_2;
	wire w_dff_B_d6OQDYRy6_2;
	wire w_dff_B_p0SDXEes4_2;
	wire w_dff_B_3rnfloFZ3_2;
	wire w_dff_B_FH9w0fmJ4_2;
	wire w_dff_B_Wx7Efk4F4_2;
	wire w_dff_B_XlOikqK90_2;
	wire w_dff_B_TmNOlf9n0_2;
	wire w_dff_B_RtdkC2mD4_1;
	wire w_dff_B_6PfcSkGz6_2;
	wire w_dff_B_oBviVAW80_2;
	wire w_dff_B_PQN2gM129_2;
	wire w_dff_B_NHsx9DbZ8_2;
	wire w_dff_B_Hu68tsAF5_2;
	wire w_dff_B_fz7Cus5n0_2;
	wire w_dff_B_x06G9Chp7_2;
	wire w_dff_B_swhybO3A6_2;
	wire w_dff_B_fy4x7IpU2_2;
	wire w_dff_B_GT8MMnUN9_2;
	wire w_dff_B_R8GnHqlY7_2;
	wire w_dff_B_BmKcjgLl8_2;
	wire w_dff_B_KvB2Wl8E0_2;
	wire w_dff_B_n0CsZ01L3_2;
	wire w_dff_B_KK4ApRKM8_2;
	wire w_dff_B_7gxUUBDR9_2;
	wire w_dff_B_4f0ajlLY9_2;
	wire w_dff_B_ILKuVmAd9_2;
	wire w_dff_B_QRIHWUsw8_2;
	wire w_dff_B_HnGLTB9O7_2;
	wire w_dff_B_GP9JAZhC8_2;
	wire w_dff_B_Fo72BbEF4_1;
	wire w_dff_B_LVlIYL3C2_2;
	wire w_dff_B_ZWCw7MDQ5_2;
	wire w_dff_B_faN7JA1a0_2;
	wire w_dff_B_zjF7C7RV7_2;
	wire w_dff_B_rfzX121o4_2;
	wire w_dff_B_Kxrdym9R8_2;
	wire w_dff_B_HIpDGStJ0_2;
	wire w_dff_B_8366iCDu3_2;
	wire w_dff_B_8YZY78lu5_2;
	wire w_dff_B_9NA4N8Lp3_2;
	wire w_dff_B_aLLSB5Lk2_2;
	wire w_dff_B_4hhFZWI41_2;
	wire w_dff_B_0fFqT3866_2;
	wire w_dff_B_6kwJyHEd0_2;
	wire w_dff_B_c4BHIpOz5_2;
	wire w_dff_B_vcEkbXEZ7_2;
	wire w_dff_B_LMs7POFQ8_2;
	wire w_dff_B_5p8CRa7h9_2;
	wire w_dff_B_vZPtaRWA8_2;
	wire w_dff_B_VX0TK40R4_1;
	wire w_dff_B_cz58degP2_2;
	wire w_dff_B_vrSXT5b96_2;
	wire w_dff_B_sHe4B7qA3_2;
	wire w_dff_B_aIdpIA1u1_2;
	wire w_dff_B_I0EmQrU52_2;
	wire w_dff_B_tLuahK4X4_2;
	wire w_dff_B_0BatgX1U8_2;
	wire w_dff_B_5TX5zvkd6_2;
	wire w_dff_B_poBBREZb0_2;
	wire w_dff_B_bsSzjpNN0_2;
	wire w_dff_B_EXJcq01N7_2;
	wire w_dff_B_kctEHTof3_2;
	wire w_dff_B_TqhesGzM8_2;
	wire w_dff_B_Q8XWme3d4_2;
	wire w_dff_B_Y8OjuYp30_2;
	wire w_dff_B_0cS1Hx3N3_2;
	wire w_dff_B_bu33HQNV7_2;
	wire w_dff_B_fD5g9lbL1_1;
	wire w_dff_B_MTQAPdOR2_2;
	wire w_dff_B_jtQ8Y7GX4_2;
	wire w_dff_B_10TE86aF9_2;
	wire w_dff_B_ncnuwJ2E3_2;
	wire w_dff_B_bzuIbQoh6_2;
	wire w_dff_B_21e51WDS9_2;
	wire w_dff_B_ERTz4txs2_2;
	wire w_dff_B_VxRWLuUO7_2;
	wire w_dff_B_O1ZusvBL0_2;
	wire w_dff_B_TDCgQw3H6_2;
	wire w_dff_B_9XHbzvvr1_2;
	wire w_dff_B_chRGbMx43_2;
	wire w_dff_B_a4v49fP78_2;
	wire w_dff_B_wXiLleDA8_2;
	wire w_dff_B_UFwAyNCv0_1;
	wire w_dff_B_MEHfKbew9_2;
	wire w_dff_B_LrNxf9oc7_2;
	wire w_dff_B_EGze31uY3_2;
	wire w_dff_B_X647aHxM6_2;
	wire w_dff_B_MSQ59Pwh8_2;
	wire w_dff_B_RuXvByrj7_2;
	wire w_dff_B_Ps3ZqFUD9_2;
	wire w_dff_B_f3mfKWtz7_2;
	wire w_dff_B_l1f4Eccm7_2;
	wire w_dff_B_XzPR8iDa5_2;
	wire w_dff_B_AJXfXcpy5_2;
	wire w_dff_B_RKXxBQcS6_2;
	wire w_dff_B_VCOEMQuA2_1;
	wire w_dff_B_yqtwYyqE3_1;
	wire w_dff_B_oh5YNsE37_1;
	wire w_dff_B_Fnn0jdrm6_1;
	wire w_dff_B_A27aPuPb3_1;
	wire w_dff_B_t0DlR4tB3_1;
	wire w_dff_B_wIvBc2Ns2_0;
	wire w_dff_B_zSHMYozx7_0;
	wire w_dff_A_p4yOhTTZ4_0;
	wire w_dff_A_MqQUNCDP0_0;
	wire w_dff_A_gsSunOMy6_0;
	wire w_dff_B_mzYTa5E69_1;
	wire w_dff_A_xi5AQlVt6_0;
	wire w_dff_A_MZXWqFtS9_1;
	wire w_dff_A_UfhNzngE2_1;
	wire w_dff_A_my0qZSVl3_1;
	wire w_dff_A_hE7lVLGO5_1;
	wire w_dff_A_71TKbdsM7_1;
	wire w_dff_A_DKvQaQ6L6_1;
	wire w_dff_A_LauM8jeY5_1;
	wire w_dff_A_AW1PADH56_1;
	wire w_dff_B_081Xrddf4_1;
	wire w_dff_B_PELpkZGR6_1;
	wire w_dff_B_UPlWjVfl7_1;
	wire w_dff_B_5v7Cwybu6_2;
	wire w_dff_B_f1OG74Oz3_2;
	wire w_dff_B_qdN04MBe9_2;
	wire w_dff_B_3dV18AZc7_2;
	wire w_dff_B_J0pmaD6N1_2;
	wire w_dff_B_ZMIiXKNE4_2;
	wire w_dff_B_r5Zq5X2H7_2;
	wire w_dff_B_frcr2BQ58_2;
	wire w_dff_B_6VN7LgEd2_2;
	wire w_dff_B_mPJKC1FO5_2;
	wire w_dff_B_3ufNL6YE1_2;
	wire w_dff_B_G0gLPMY86_2;
	wire w_dff_B_CMuiVO743_2;
	wire w_dff_B_jbWSueBK0_2;
	wire w_dff_B_rnx8ihFa0_2;
	wire w_dff_B_lkEdDCNd5_2;
	wire w_dff_B_5Kqjs0H78_2;
	wire w_dff_B_yTlv3t160_2;
	wire w_dff_B_eP7KzkAU1_2;
	wire w_dff_B_zHfpANWv3_2;
	wire w_dff_B_2VKmsVJD1_2;
	wire w_dff_B_pDgrJjwb8_2;
	wire w_dff_B_NCEZoyRg9_2;
	wire w_dff_B_hpRTIMEf5_2;
	wire w_dff_B_uw15CJv09_2;
	wire w_dff_B_7SqJUegL5_2;
	wire w_dff_B_fsTo1ptP8_2;
	wire w_dff_B_pFdLz4Cc4_2;
	wire w_dff_B_nGEyyGEa8_2;
	wire w_dff_B_kkk8bx8y7_2;
	wire w_dff_B_oXHz3RBJ8_2;
	wire w_dff_B_4cTCC7kT1_2;
	wire w_dff_B_pSZ7TYnB4_2;
	wire w_dff_B_pB83XQWe5_2;
	wire w_dff_B_d64f9uoR8_2;
	wire w_dff_B_U1DOPePd6_2;
	wire w_dff_B_LMq2bu8i3_2;
	wire w_dff_B_TcZANVD60_2;
	wire w_dff_B_tcfZoO6z3_2;
	wire w_dff_B_S2lf0fWp3_2;
	wire w_dff_B_3CAGL5ax6_2;
	wire w_dff_B_ljXJ2ynj2_2;
	wire w_dff_B_665JCJru3_2;
	wire w_dff_B_zOTBCFUP3_2;
	wire w_dff_B_CVk7hsi26_2;
	wire w_dff_B_pddNHisA9_2;
	wire w_dff_B_OsphWy6H8_2;
	wire w_dff_B_lhckDvac9_2;
	wire w_dff_B_mWv5pILD7_2;
	wire w_dff_B_nBofrBcW4_2;
	wire w_dff_B_bSDy59976_2;
	wire w_dff_B_JLr79cM30_2;
	wire w_dff_B_T26zHkVu5_2;
	wire w_dff_B_r62pziid6_2;
	wire w_dff_B_dLkIvAW73_2;
	wire w_dff_B_DWU7mLRu5_2;
	wire w_dff_B_v6oMuJO42_2;
	wire w_dff_B_Rm6MhEQf4_2;
	wire w_dff_B_HtVBoJV96_2;
	wire w_dff_B_PVvCbUy14_2;
	wire w_dff_B_KmfJV7hs9_2;
	wire w_dff_B_kXzCZgBD6_2;
	wire w_dff_B_fwUUWTIM0_2;
	wire w_dff_B_OHFUtWk27_2;
	wire w_dff_B_Of0j8XoX2_2;
	wire w_dff_B_JORh3Z2K5_2;
	wire w_dff_B_kKn3i41J6_2;
	wire w_dff_B_NkkRH9ZQ8_2;
	wire w_dff_B_2GkZ8hpD9_2;
	wire w_dff_B_eujWYkjA4_2;
	wire w_dff_B_KRbT3pt91_2;
	wire w_dff_B_JhzzV94S2_2;
	wire w_dff_B_hz98RGvz8_2;
	wire w_dff_B_08fJ1fTh5_2;
	wire w_dff_B_d6Hgq5M18_2;
	wire w_dff_B_f0vzKlBO2_2;
	wire w_dff_B_cZyrIjHG1_2;
	wire w_dff_B_KbZiRDfg4_2;
	wire w_dff_B_NSWvBMA29_2;
	wire w_dff_B_1oX7jY9N5_2;
	wire w_dff_B_ajKvOeor9_2;
	wire w_dff_B_hRclBnZW3_2;
	wire w_dff_B_vlt6mRqO8_2;
	wire w_dff_B_CQ4DIJ6n0_2;
	wire w_dff_B_O0ZoKvlz7_2;
	wire w_dff_B_xMIDyI3U4_2;
	wire w_dff_B_qLMiArfw7_2;
	wire w_dff_B_zwtG02J54_2;
	wire w_dff_B_YaN0fOWd5_2;
	wire w_dff_B_lysFEHkd7_2;
	wire w_dff_B_VMaSCxnd1_2;
	wire w_dff_B_pVXkeNhE4_2;
	wire w_dff_B_IuMVvph68_2;
	wire w_dff_B_GekZBews5_2;
	wire w_dff_B_fEGvgOtp1_2;
	wire w_dff_B_UapzPCYt3_2;
	wire w_dff_B_0DBgrgZV6_2;
	wire w_dff_B_Ui2zdgbZ5_2;
	wire w_dff_B_robcFZAe6_2;
	wire w_dff_B_3ITGfKaW9_2;
	wire w_dff_B_BDOogQE10_2;
	wire w_dff_B_6B4Ao2BR9_2;
	wire w_dff_B_H35qfwNg9_2;
	wire w_dff_B_FyEso6WK7_2;
	wire w_dff_B_yBtzNJ2J0_2;
	wire w_dff_B_S0RrCZ7l0_2;
	wire w_dff_B_ylm2zTC42_2;
	wire w_dff_B_jTuo7NQI0_2;
	wire w_dff_B_he1rIc3I5_2;
	wire w_dff_B_836wzKpd8_2;
	wire w_dff_B_7dGqTvEF8_2;
	wire w_dff_B_3QhjI9FW5_2;
	wire w_dff_B_KwmOwAnj1_2;
	wire w_dff_B_fosja2Hu4_2;
	wire w_dff_A_aQrQ35x31_1;
	wire w_dff_B_C92hqvgL8_1;
	wire w_dff_B_grHPxLff2_2;
	wire w_dff_B_2t0uBdcP6_2;
	wire w_dff_B_Agovedgy2_2;
	wire w_dff_B_XnFqnkd55_2;
	wire w_dff_B_nRECSmre3_2;
	wire w_dff_B_Gbg1xO0r7_2;
	wire w_dff_B_dLnvZYU03_2;
	wire w_dff_B_mGjCruk43_2;
	wire w_dff_B_Ds66a7Zk9_2;
	wire w_dff_B_4NHEN7pu4_2;
	wire w_dff_B_pzRuHHUT5_2;
	wire w_dff_B_dIIfp8xh6_2;
	wire w_dff_B_jWvrj71G7_2;
	wire w_dff_B_Ja1ABzjF7_2;
	wire w_dff_B_5CoJBZyy4_2;
	wire w_dff_B_S15C6HcH4_2;
	wire w_dff_B_lyuZzVzM8_2;
	wire w_dff_B_yPAyk9lF2_2;
	wire w_dff_B_lk2w28Fo1_2;
	wire w_dff_B_sV5fIFD98_2;
	wire w_dff_B_6zrt42610_2;
	wire w_dff_B_jtnQ4U8k3_2;
	wire w_dff_B_SZvDbafQ3_2;
	wire w_dff_B_SDNxZN1g3_2;
	wire w_dff_B_dhSrtEEv9_2;
	wire w_dff_B_IBTHqlCX4_2;
	wire w_dff_B_FYvFNWhv6_2;
	wire w_dff_B_NPGUVlxb0_2;
	wire w_dff_B_MWl8q4I98_2;
	wire w_dff_B_kMgM8Tg71_2;
	wire w_dff_B_LSOUMlfv1_2;
	wire w_dff_B_G4BYq1t22_2;
	wire w_dff_B_StOvbnaR9_2;
	wire w_dff_B_or6V7SCe8_2;
	wire w_dff_B_5XqyY2eQ6_2;
	wire w_dff_B_1dDZwQAr9_2;
	wire w_dff_B_sD0CfKGj3_2;
	wire w_dff_B_YjL7x2uR4_2;
	wire w_dff_B_uAUcWnL02_2;
	wire w_dff_B_vRsIJSpv7_2;
	wire w_dff_B_42mpVIHe2_2;
	wire w_dff_B_yl0REqCP3_2;
	wire w_dff_B_CvoZ9Ung1_2;
	wire w_dff_B_ml8z6I3A4_2;
	wire w_dff_B_4blErXlR5_2;
	wire w_dff_B_7EkaFK5e0_2;
	wire w_dff_B_A1ZfeXeZ0_2;
	wire w_dff_B_U8JkEi1S5_2;
	wire w_dff_B_J7GcF8Kw5_2;
	wire w_dff_B_woChbYS79_2;
	wire w_dff_B_EjCfjk3d5_2;
	wire w_dff_B_kb8mRVRf4_2;
	wire w_dff_B_66jx00kP9_2;
	wire w_dff_B_p3eyB6Cd5_2;
	wire w_dff_B_eIaXRKAC9_2;
	wire w_dff_B_3ETeiOUN6_1;
	wire w_dff_B_4p6E7E1O0_1;
	wire w_dff_B_r5DEL3wF3_2;
	wire w_dff_B_41nrji832_2;
	wire w_dff_B_8F8cbYSV3_2;
	wire w_dff_B_BsFOJEvq2_2;
	wire w_dff_B_RMjv8qhD2_2;
	wire w_dff_B_Xefi5GXi6_2;
	wire w_dff_B_ZiS5HXpC5_2;
	wire w_dff_B_UcpOn7Jw3_2;
	wire w_dff_B_GRDGAL5z3_2;
	wire w_dff_B_DkiRuxjS4_2;
	wire w_dff_B_JmQDMNcD6_2;
	wire w_dff_B_40TCthHB3_2;
	wire w_dff_B_HLiXnyRE4_2;
	wire w_dff_B_J4o6ukSd5_2;
	wire w_dff_B_5NfzmMAL4_2;
	wire w_dff_B_bT8o41Ha4_2;
	wire w_dff_B_hCVkK3CI6_2;
	wire w_dff_B_Nn5HNoY04_2;
	wire w_dff_B_jGjPlxOJ2_2;
	wire w_dff_B_sioFT1Gn2_2;
	wire w_dff_B_s7w2bqc97_2;
	wire w_dff_B_m5vN53pR8_2;
	wire w_dff_B_1ajmfdsi1_2;
	wire w_dff_B_ZVb7hnVn9_2;
	wire w_dff_B_kTg5F5Uw8_2;
	wire w_dff_B_BfAL3iO21_2;
	wire w_dff_B_vlYk47kL3_2;
	wire w_dff_B_m8yavwcg5_2;
	wire w_dff_B_HvUKYcwq5_2;
	wire w_dff_B_mnqqvzLX5_2;
	wire w_dff_B_XJOE9A6E5_2;
	wire w_dff_B_PVsj90Kj4_2;
	wire w_dff_B_6B4ijnv61_2;
	wire w_dff_B_JJ7eaP0L2_2;
	wire w_dff_B_OaljYqE97_2;
	wire w_dff_B_Ydaoss7M1_2;
	wire w_dff_B_h6yxs8or0_2;
	wire w_dff_B_KjWYSJ7N2_2;
	wire w_dff_B_HqwWS43L9_2;
	wire w_dff_B_YyNfbTiP0_2;
	wire w_dff_B_N9BA0jPQ2_2;
	wire w_dff_B_noWhhSHy3_2;
	wire w_dff_B_BCpTLhAm0_2;
	wire w_dff_B_zRJPFy7l0_2;
	wire w_dff_B_1DRiESHt5_2;
	wire w_dff_B_PgG3sjmQ2_2;
	wire w_dff_B_gZWKAKOx8_2;
	wire w_dff_B_Lh3Q3shL4_2;
	wire w_dff_B_lUCdtiE86_2;
	wire w_dff_B_Nozv5TuX6_2;
	wire w_dff_B_AmTbGDv35_2;
	wire w_dff_B_ow1ACzzW2_2;
	wire w_dff_B_HFGdEqMT4_2;
	wire w_dff_B_FNKI545q1_2;
	wire w_dff_B_KrnCxEr38_2;
	wire w_dff_B_DauTOFYo8_2;
	wire w_dff_B_IV5fNUIQ2_2;
	wire w_dff_B_ho4FAEGm2_2;
	wire w_dff_B_cY8mQqxw9_2;
	wire w_dff_B_D1La8O7d4_2;
	wire w_dff_B_mSswtA1x9_2;
	wire w_dff_B_owMSigKX4_2;
	wire w_dff_B_4QbQ19Db6_2;
	wire w_dff_B_8XDFSGgI4_2;
	wire w_dff_B_ViWPzmuD8_2;
	wire w_dff_B_5y5s0Fwa5_2;
	wire w_dff_B_AROnbn3k2_2;
	wire w_dff_B_Mg6T2Yox1_2;
	wire w_dff_B_AFIxo8Gk2_2;
	wire w_dff_B_rylRi0Fa8_2;
	wire w_dff_B_wbsNyRlg3_2;
	wire w_dff_B_VIYIXzl65_2;
	wire w_dff_B_H0yJlRON3_2;
	wire w_dff_B_JmeE15He0_2;
	wire w_dff_B_N4uAV5mt4_2;
	wire w_dff_B_hFx8PE626_2;
	wire w_dff_B_R9P3XLvI8_2;
	wire w_dff_B_GcIMSQIs1_2;
	wire w_dff_B_RSrqNa6d8_2;
	wire w_dff_B_I3e2HnSc6_2;
	wire w_dff_B_6v8dgnx22_2;
	wire w_dff_B_VhYtEGdF0_2;
	wire w_dff_B_Zk5GAJos8_2;
	wire w_dff_B_TQuqQPn63_2;
	wire w_dff_B_GItCAx1e5_2;
	wire w_dff_B_Q7WRgSCv3_2;
	wire w_dff_B_mqDfCepF3_2;
	wire w_dff_B_w5f0Zlpc7_2;
	wire w_dff_B_M4Scfoab0_2;
	wire w_dff_B_YzKK4ROU9_2;
	wire w_dff_B_8p4IIfyw3_2;
	wire w_dff_B_JVjmycqe6_2;
	wire w_dff_B_h8pzWNGf7_2;
	wire w_dff_B_Xdq2iI6f7_2;
	wire w_dff_B_M0uDOyqm7_2;
	wire w_dff_B_wYU0PGcR7_2;
	wire w_dff_B_wn0HOENM2_2;
	wire w_dff_B_pG2N7egd5_2;
	wire w_dff_B_UsXC6kDV5_2;
	wire w_dff_B_8DaWnkuS7_2;
	wire w_dff_B_yBGWBQQ73_2;
	wire w_dff_B_HMAyniji3_2;
	wire w_dff_B_qj2Sy5ei5_2;
	wire w_dff_B_kHRFU87x7_2;
	wire w_dff_B_TSuX6jo15_2;
	wire w_dff_B_NjmfjCyy8_2;
	wire w_dff_B_hqG9jUJl5_2;
	wire w_dff_B_HZcRA8yf1_1;
	wire w_dff_B_DBvI3FUx2_2;
	wire w_dff_B_0bcAbLjy1_2;
	wire w_dff_B_pLM2oyV69_2;
	wire w_dff_B_QyA5ih9P2_2;
	wire w_dff_B_tlYb8Ct29_2;
	wire w_dff_B_GUWN96WQ5_2;
	wire w_dff_B_XE9YeepA2_2;
	wire w_dff_B_QeLZ2IJi2_2;
	wire w_dff_B_FBoJmY6D3_2;
	wire w_dff_B_cNUbaqCd4_2;
	wire w_dff_B_BzgW8faj8_2;
	wire w_dff_B_cGdMyVA66_2;
	wire w_dff_B_A7Xjo4ef8_2;
	wire w_dff_B_0tvM4rOw1_2;
	wire w_dff_B_0MFJM3tm7_2;
	wire w_dff_B_9QnjixyN7_2;
	wire w_dff_B_u6xCdFJu4_2;
	wire w_dff_B_zmE3oj9M0_2;
	wire w_dff_B_WtUrwfds3_2;
	wire w_dff_B_4wu9n1Mw6_2;
	wire w_dff_B_nDrme8X40_2;
	wire w_dff_B_6YbSQnxc5_2;
	wire w_dff_B_j9s88Kr50_2;
	wire w_dff_B_n5MbotQ47_2;
	wire w_dff_B_QdihqDre8_2;
	wire w_dff_B_VrAU1dhq1_2;
	wire w_dff_B_fixnhraI4_2;
	wire w_dff_B_XJFtRB5M8_2;
	wire w_dff_B_qOCNdoRj7_2;
	wire w_dff_B_AnMfmTVn5_2;
	wire w_dff_B_cznM22t16_2;
	wire w_dff_B_bynwQf8f8_2;
	wire w_dff_B_PoecEloe9_2;
	wire w_dff_B_YEvfCuoy8_2;
	wire w_dff_B_rnrDXxx41_2;
	wire w_dff_B_OECkqqyE4_2;
	wire w_dff_B_1b1BGJsA9_2;
	wire w_dff_B_TvnV2T2i9_2;
	wire w_dff_B_wiJHOoZ48_2;
	wire w_dff_B_SzOkO6av7_2;
	wire w_dff_B_Uxw2Ipnu7_2;
	wire w_dff_B_blLPoyJI9_2;
	wire w_dff_B_yE1wnOeW0_2;
	wire w_dff_B_FtgpU8QG4_2;
	wire w_dff_B_OoBrKVxl6_2;
	wire w_dff_B_b5X33vDF0_2;
	wire w_dff_B_mS5tJWfv6_2;
	wire w_dff_B_lk55Bam87_2;
	wire w_dff_B_KS0wfYEv8_2;
	wire w_dff_B_Dvayqm2X9_2;
	wire w_dff_B_fpdTFUYa8_2;
	wire w_dff_B_IRqDxaMe2_1;
	wire w_dff_B_hxknXZrK4_1;
	wire w_dff_B_5KS1wJEA4_2;
	wire w_dff_B_kywnD8D52_2;
	wire w_dff_B_JA8KGkvM4_2;
	wire w_dff_B_HbnxkMWh2_2;
	wire w_dff_B_P0esF45n4_2;
	wire w_dff_B_XCEmDejO7_2;
	wire w_dff_B_YEiDr6lP2_2;
	wire w_dff_B_1AgA72WP7_2;
	wire w_dff_B_BgpCTGJ53_2;
	wire w_dff_B_WfNCh4uI6_2;
	wire w_dff_B_gH4EAu6N1_2;
	wire w_dff_B_YvK5si3a3_2;
	wire w_dff_B_pGSOdx9c0_2;
	wire w_dff_B_YVHKVAro5_2;
	wire w_dff_B_ybRAsPRh1_2;
	wire w_dff_B_dpliggGD8_2;
	wire w_dff_B_SYalu5ew7_2;
	wire w_dff_B_JPK31wup3_2;
	wire w_dff_B_2pjFRDFr0_2;
	wire w_dff_B_b2UZ6BZj7_2;
	wire w_dff_B_W8ek7kr86_2;
	wire w_dff_B_aUo1xKZw6_2;
	wire w_dff_B_ZqZfp8yf8_2;
	wire w_dff_B_ZfTsfHxK5_2;
	wire w_dff_B_Jxaxbwb33_2;
	wire w_dff_B_pyyKvmwy2_2;
	wire w_dff_B_L7Fcjvbs8_2;
	wire w_dff_B_PnLBA0UL6_2;
	wire w_dff_B_pYvE194M6_2;
	wire w_dff_B_Ei8ldF8G1_2;
	wire w_dff_B_1PeOV0S97_2;
	wire w_dff_B_1dCMWeoB6_2;
	wire w_dff_B_7PZTt0Nl6_2;
	wire w_dff_B_Nixu45cg7_2;
	wire w_dff_B_o9BeNMxs4_2;
	wire w_dff_B_dPjRhudc3_2;
	wire w_dff_B_I18DbIgU8_2;
	wire w_dff_B_fl6qs6778_2;
	wire w_dff_B_ryPWfqGa6_2;
	wire w_dff_B_9pQwhCmg7_2;
	wire w_dff_B_WMqxo3Es3_2;
	wire w_dff_B_kYVTeL8l2_2;
	wire w_dff_B_ok5uJN1p7_2;
	wire w_dff_B_siBtAxSY7_2;
	wire w_dff_B_qWczEMzF2_2;
	wire w_dff_B_TIO3sbTp7_2;
	wire w_dff_B_swwn3wE48_2;
	wire w_dff_B_BsNym0BD6_2;
	wire w_dff_B_ealXpbdV2_2;
	wire w_dff_B_8iza5Kt46_2;
	wire w_dff_B_GXbmv8rY9_2;
	wire w_dff_B_XOeGf7qs7_2;
	wire w_dff_B_v6Cgo9NB8_2;
	wire w_dff_B_wSEXmgPU0_2;
	wire w_dff_B_hBHke2de9_2;
	wire w_dff_B_UNMbelaW4_2;
	wire w_dff_B_kobvEVYX1_2;
	wire w_dff_B_UnQM4R7c6_2;
	wire w_dff_B_LCbHCw8t7_2;
	wire w_dff_B_HzALTBaN4_2;
	wire w_dff_B_tysyyMfp0_2;
	wire w_dff_B_m5zu1xe02_2;
	wire w_dff_B_qQP2INB56_2;
	wire w_dff_B_u60CNJ896_2;
	wire w_dff_B_PHrOfp9n6_2;
	wire w_dff_B_QJ3luVGO8_2;
	wire w_dff_B_HAjFXVIc1_2;
	wire w_dff_B_PMh6y69q2_2;
	wire w_dff_B_xmGpfmcz5_2;
	wire w_dff_B_Lk5xmkvt5_2;
	wire w_dff_B_8AoPRLl48_2;
	wire w_dff_B_VSxlUXr04_2;
	wire w_dff_B_yTOMP64G7_2;
	wire w_dff_B_Df3n2kFg9_2;
	wire w_dff_B_sg3UA50U7_2;
	wire w_dff_B_oq90p8J44_2;
	wire w_dff_B_5u973HIt0_2;
	wire w_dff_B_D8vfNS1L9_2;
	wire w_dff_B_Lac3mYhn1_2;
	wire w_dff_B_iJYaALo58_2;
	wire w_dff_B_hxm3uO8t9_2;
	wire w_dff_B_w41tatFL0_2;
	wire w_dff_B_nh76Sbsk4_2;
	wire w_dff_B_SldmnIo06_2;
	wire w_dff_B_JJZvrVZY7_2;
	wire w_dff_B_qSktLfQv8_2;
	wire w_dff_B_xROvHceJ8_2;
	wire w_dff_B_dRrEVYHj5_2;
	wire w_dff_B_8F4mGf0c5_2;
	wire w_dff_B_rAZiex4m4_2;
	wire w_dff_B_LzIUIt3x7_2;
	wire w_dff_B_HfomW0Ed8_2;
	wire w_dff_B_md8JpPnn8_2;
	wire w_dff_B_SOKTh8qq0_2;
	wire w_dff_B_eZk0nAOL2_2;
	wire w_dff_B_7r3JzWwv3_2;
	wire w_dff_B_UyeOzMud5_2;
	wire w_dff_B_ZgDUxRu08_2;
	wire w_dff_B_jQz8xYvG9_2;
	wire w_dff_B_4H58eYGh5_1;
	wire w_dff_B_iK0CLIKr8_2;
	wire w_dff_B_gJhXQPSx6_2;
	wire w_dff_B_clkvx3ng3_2;
	wire w_dff_B_HUTX4Mc65_2;
	wire w_dff_B_ICUFsK3n1_2;
	wire w_dff_B_A4EuyVaJ1_2;
	wire w_dff_B_BT39IYJk7_2;
	wire w_dff_B_iHUdGvY64_2;
	wire w_dff_B_Vkybx9sd6_2;
	wire w_dff_B_2hR0JXpz0_2;
	wire w_dff_B_BONtfjYJ0_2;
	wire w_dff_B_S5PEcgqK1_2;
	wire w_dff_B_EIshArMQ8_2;
	wire w_dff_B_oKJfnPyo3_2;
	wire w_dff_B_7MRlVLlA9_2;
	wire w_dff_B_IxnnyTHG6_2;
	wire w_dff_B_qtsZK9MU1_2;
	wire w_dff_B_aNBclOXF6_2;
	wire w_dff_B_Kak0d9OD3_2;
	wire w_dff_B_KeMCybJm5_2;
	wire w_dff_B_81SBDW203_2;
	wire w_dff_B_1V6OoTMh3_2;
	wire w_dff_B_RaGXJgGj1_2;
	wire w_dff_B_o8GRixEZ3_2;
	wire w_dff_B_pLjPmnNs7_2;
	wire w_dff_B_5yyJ8P2h7_2;
	wire w_dff_B_uyht0P7T4_2;
	wire w_dff_B_gOzMkHVW5_2;
	wire w_dff_B_oQjzj1si8_2;
	wire w_dff_B_hlNPSmZN2_2;
	wire w_dff_B_hNyIm47R4_2;
	wire w_dff_B_7IPpYafO4_2;
	wire w_dff_B_lX9rPIp45_2;
	wire w_dff_B_akycZ8pd1_2;
	wire w_dff_B_Xrqzdsys4_2;
	wire w_dff_B_plqKYCF24_2;
	wire w_dff_B_p29naSmn1_2;
	wire w_dff_B_HP8VGHm88_2;
	wire w_dff_B_HdqSspbk1_2;
	wire w_dff_B_r0mf3nj57_2;
	wire w_dff_B_HIEjp3Vf1_2;
	wire w_dff_B_KZMw3vOh0_2;
	wire w_dff_B_dJDkOySD7_2;
	wire w_dff_B_GgSrqpV50_2;
	wire w_dff_B_aoa3D9JD2_2;
	wire w_dff_B_wSk8cq3o3_2;
	wire w_dff_B_DI2GWMrx8_2;
	wire w_dff_B_Ywyy6tRh3_1;
	wire w_dff_B_yr9DqX8w2_1;
	wire w_dff_B_ZBHDNJzt6_2;
	wire w_dff_B_RmLoZWni9_2;
	wire w_dff_B_yjM5zYcU9_2;
	wire w_dff_B_n3A0exga1_2;
	wire w_dff_B_QtAb0TbW6_2;
	wire w_dff_B_0dSs4GBc5_2;
	wire w_dff_B_hC7cbqva6_2;
	wire w_dff_B_gUP1Vrog7_2;
	wire w_dff_B_xIHU875o3_2;
	wire w_dff_B_BZ5gUWDc3_2;
	wire w_dff_B_SduZHkGW3_2;
	wire w_dff_B_rY42VeaF9_2;
	wire w_dff_B_JpIlw6kJ2_2;
	wire w_dff_B_Req1KuG09_2;
	wire w_dff_B_1u2LQapE3_2;
	wire w_dff_B_Um9K5SFx7_2;
	wire w_dff_B_00UchqWP0_2;
	wire w_dff_B_YxL4j6fr9_2;
	wire w_dff_B_jmYPMs3A7_2;
	wire w_dff_B_KTaYiATc4_2;
	wire w_dff_B_GT5CY0NJ1_2;
	wire w_dff_B_uPnJlxGY6_2;
	wire w_dff_B_4TfFEFmg9_2;
	wire w_dff_B_bCnXdMgz3_2;
	wire w_dff_B_HzCfA7cZ8_2;
	wire w_dff_B_BFKUpc1U5_2;
	wire w_dff_B_0LRMnEKd8_2;
	wire w_dff_B_uglbfiYX0_2;
	wire w_dff_B_QGDZ9MTw1_2;
	wire w_dff_B_5Meo4a0n4_2;
	wire w_dff_B_SA7uSTSo8_2;
	wire w_dff_B_azP34OCt8_2;
	wire w_dff_B_pX9ORayd2_2;
	wire w_dff_B_Me2PQC3N9_2;
	wire w_dff_B_OxvjDJ3p1_2;
	wire w_dff_B_BwER6cLT9_2;
	wire w_dff_B_sXh5Bkkm4_2;
	wire w_dff_B_deZ7pzqU8_2;
	wire w_dff_B_TvISKjQx3_2;
	wire w_dff_B_lr0asqRj2_2;
	wire w_dff_B_WYGTdMM76_2;
	wire w_dff_B_U2e5r6Nl9_2;
	wire w_dff_B_JvU7r4pt9_2;
	wire w_dff_B_DfVGyMBd9_2;
	wire w_dff_B_dmwKZURY8_2;
	wire w_dff_B_SXHO6v2R8_2;
	wire w_dff_B_AXoFbq769_2;
	wire w_dff_B_A6m6aOKY2_2;
	wire w_dff_B_bgIJkmEK1_2;
	wire w_dff_B_KTE7Lz235_2;
	wire w_dff_B_gmtkPaLR3_2;
	wire w_dff_B_LhX2oZAg1_2;
	wire w_dff_B_rXEFJwjP6_2;
	wire w_dff_B_GJZ9DoLp6_2;
	wire w_dff_B_VebLElUT1_2;
	wire w_dff_B_J01WigQ02_2;
	wire w_dff_B_XJU5Cm8H4_2;
	wire w_dff_B_UcD1Ktzn3_2;
	wire w_dff_B_8PvWckt09_2;
	wire w_dff_B_xnWoSRgK2_2;
	wire w_dff_B_v3seb3v67_2;
	wire w_dff_B_PFm7VDJ03_2;
	wire w_dff_B_H8JqCsWv3_2;
	wire w_dff_B_s5hRRsaH8_2;
	wire w_dff_B_XIEIcuha0_2;
	wire w_dff_B_Qx86ozSY4_2;
	wire w_dff_B_YWkvLIPl9_2;
	wire w_dff_B_Qlte1brX2_2;
	wire w_dff_B_qZScaye56_2;
	wire w_dff_B_PQjzMQKF6_2;
	wire w_dff_B_IaYODAFQ0_2;
	wire w_dff_B_EB9xEaQh4_2;
	wire w_dff_B_ik7VVAML4_2;
	wire w_dff_B_WFEwjM4p7_2;
	wire w_dff_B_BzHw6BKf6_2;
	wire w_dff_B_c1Yp6nVe7_2;
	wire w_dff_B_kENMhCXh5_2;
	wire w_dff_B_fw8qvMm93_2;
	wire w_dff_B_hQUSD2Ng3_2;
	wire w_dff_B_u5CPnxKk6_2;
	wire w_dff_B_hO2WXrgp2_2;
	wire w_dff_B_0BPhTIYv2_2;
	wire w_dff_B_qq5oRZqx1_2;
	wire w_dff_B_n31KSzgu9_2;
	wire w_dff_B_0jfTam7d6_2;
	wire w_dff_B_CEhtiWqJ5_2;
	wire w_dff_B_14UZf4QF2_2;
	wire w_dff_B_S55qrRp56_2;
	wire w_dff_B_YlIqJLc14_2;
	wire w_dff_B_o76WopWf3_2;
	wire w_dff_B_AdJXDMSH1_2;
	wire w_dff_B_15EDfjX83_1;
	wire w_dff_B_hw018sdB4_2;
	wire w_dff_B_w1GA6uHh1_2;
	wire w_dff_B_WUq4pdFE3_2;
	wire w_dff_B_nl0jVKUQ3_2;
	wire w_dff_B_5qBng3mg5_2;
	wire w_dff_B_KdTJFGpu1_2;
	wire w_dff_B_eAEFeRr96_2;
	wire w_dff_B_UQQ4umHl8_2;
	wire w_dff_B_MNn7b7Xs9_2;
	wire w_dff_B_LqY1PsdG1_2;
	wire w_dff_B_G9ctXz6g4_2;
	wire w_dff_B_npYuCtBM9_2;
	wire w_dff_B_zvV1A57O7_2;
	wire w_dff_B_MRy8ADoc4_2;
	wire w_dff_B_BpPjR14f1_2;
	wire w_dff_B_oUISqR6o9_2;
	wire w_dff_B_36X7dkTJ0_2;
	wire w_dff_B_cAQL9vEU0_2;
	wire w_dff_B_Jong7ev57_2;
	wire w_dff_B_EkqaA7YN8_2;
	wire w_dff_B_CEDnOjeO9_2;
	wire w_dff_B_UE83noeL6_2;
	wire w_dff_B_ORLXTgM02_2;
	wire w_dff_B_NPDXFtjq4_2;
	wire w_dff_B_webvFmka7_2;
	wire w_dff_B_35URPWFz7_2;
	wire w_dff_B_JeGnx6XI0_2;
	wire w_dff_B_IuYgknc22_2;
	wire w_dff_B_5bA0Ij1U2_2;
	wire w_dff_B_AooL0T7V5_2;
	wire w_dff_B_4pYvItSK8_2;
	wire w_dff_B_f2FJ0NOx6_2;
	wire w_dff_B_uEmygJSJ5_2;
	wire w_dff_B_JFA7JtGe1_2;
	wire w_dff_B_3rzeB9eI1_2;
	wire w_dff_B_tcYRE7Kr5_2;
	wire w_dff_B_JJ2X8Wkx6_2;
	wire w_dff_B_5O9OFVnQ4_2;
	wire w_dff_B_250ee1ss1_2;
	wire w_dff_B_eXC6rSt59_2;
	wire w_dff_B_YYr8HkEN2_2;
	wire w_dff_B_ELxEnowF3_2;
	wire w_dff_B_Jq1IKcFg1_2;
	wire w_dff_B_fcbH6VQR2_1;
	wire w_dff_B_bI5IHVx85_1;
	wire w_dff_B_lteTwQdY1_2;
	wire w_dff_B_iLcR157s8_2;
	wire w_dff_B_eZMmiQCN8_2;
	wire w_dff_B_S5naS7Vj3_2;
	wire w_dff_B_RZeVmmhQ4_2;
	wire w_dff_B_fxRrV9pX4_2;
	wire w_dff_B_X8NUlGL60_2;
	wire w_dff_B_xgQOqUCw7_2;
	wire w_dff_B_fC2WItM03_2;
	wire w_dff_B_EGZFkNvT4_2;
	wire w_dff_B_DDLyHUMJ9_2;
	wire w_dff_B_wfJQxeM52_2;
	wire w_dff_B_dTSHe7BF0_2;
	wire w_dff_B_z2yU9exO5_2;
	wire w_dff_B_2sssUxLd8_2;
	wire w_dff_B_awshfGlE6_2;
	wire w_dff_B_LNURQio10_2;
	wire w_dff_B_ByZzTT6o7_2;
	wire w_dff_B_XnHKelct7_2;
	wire w_dff_B_A3VL9cYM8_2;
	wire w_dff_B_gyfyoaY33_2;
	wire w_dff_B_PX5SqSWe1_2;
	wire w_dff_B_SmpGvvSq4_2;
	wire w_dff_B_S3tmkxzO9_2;
	wire w_dff_B_d8v3CkdT2_2;
	wire w_dff_B_jkyGrMiy0_2;
	wire w_dff_B_UmyfR7cI8_2;
	wire w_dff_B_0gsQyXWp5_2;
	wire w_dff_B_46xgBcQX6_2;
	wire w_dff_B_mj1QzL3k1_2;
	wire w_dff_B_bI7ElMqh7_2;
	wire w_dff_B_g6H5fklB8_2;
	wire w_dff_B_BGr92eYH7_2;
	wire w_dff_B_gT91Cokv4_2;
	wire w_dff_B_891SdkNe1_2;
	wire w_dff_B_D53wKc4P8_2;
	wire w_dff_B_9zP7aAPd5_2;
	wire w_dff_B_BpSotqvJ2_2;
	wire w_dff_B_MwHRYxnq2_2;
	wire w_dff_B_io3x0prC6_2;
	wire w_dff_B_Hbpoq7ZI9_2;
	wire w_dff_B_4K9zM5Yz5_2;
	wire w_dff_B_GFpIGppL7_2;
	wire w_dff_B_uxbj7PjQ9_2;
	wire w_dff_B_aMkKiomu6_2;
	wire w_dff_B_3LSiX3WJ0_2;
	wire w_dff_B_WRnF1dbG2_2;
	wire w_dff_B_YpoexdLl1_2;
	wire w_dff_B_ONCPzIwO2_2;
	wire w_dff_B_fAufSgq51_2;
	wire w_dff_B_l0RKTsTW7_2;
	wire w_dff_B_Z1c9yUfT4_2;
	wire w_dff_B_uhLlVpYw7_2;
	wire w_dff_B_PqVieLC61_2;
	wire w_dff_B_XDL8dbcl6_2;
	wire w_dff_B_INqlzx837_2;
	wire w_dff_B_Hb9zzTJE2_2;
	wire w_dff_B_56KtMsJx4_2;
	wire w_dff_B_cvKGoKbM4_2;
	wire w_dff_B_ZZCrM4em0_2;
	wire w_dff_B_YaQLFveC0_2;
	wire w_dff_B_8UFTCT2L5_2;
	wire w_dff_B_GICkqN6N8_2;
	wire w_dff_B_6mlta9xD4_2;
	wire w_dff_B_d9rEHVlX3_2;
	wire w_dff_B_NrsRAcI75_2;
	wire w_dff_B_azmRlFvL6_2;
	wire w_dff_B_K0NkzhIB2_2;
	wire w_dff_B_l6rcGCcK6_2;
	wire w_dff_B_8NaDjJ7R7_2;
	wire w_dff_B_LEyHWSU28_2;
	wire w_dff_B_kwg80eUZ5_2;
	wire w_dff_B_1raf0HVA7_2;
	wire w_dff_B_290cngb96_2;
	wire w_dff_B_UrUNSdwe0_2;
	wire w_dff_B_qX66UXMo7_2;
	wire w_dff_B_tPxFV14z8_2;
	wire w_dff_B_Qd9CJMmI7_2;
	wire w_dff_B_1BzwHCJs7_2;
	wire w_dff_B_x4Wou5S19_2;
	wire w_dff_B_XXPJS6kv8_2;
	wire w_dff_B_PBFYhsH57_2;
	wire w_dff_B_vpqxp1Kb7_2;
	wire w_dff_B_9ydfEmg55_1;
	wire w_dff_B_ZMS2Vlgh3_2;
	wire w_dff_B_SqCleVKN9_2;
	wire w_dff_B_vK3Zz64v9_2;
	wire w_dff_B_fXarcyMf0_2;
	wire w_dff_B_Se9J04Kq3_2;
	wire w_dff_B_zFJDWkud6_2;
	wire w_dff_B_jJShNd7i2_2;
	wire w_dff_B_toKTsgxP8_2;
	wire w_dff_B_d9j0DKPJ6_2;
	wire w_dff_B_Nl3ZX58E8_2;
	wire w_dff_B_gIEUCPnm6_2;
	wire w_dff_B_DRaPI8Wl7_2;
	wire w_dff_B_kwuV2xiU5_2;
	wire w_dff_B_Xk6vgI0U5_2;
	wire w_dff_B_hq6ZSFrN0_2;
	wire w_dff_B_F3EP3AeZ4_2;
	wire w_dff_B_LAizMQ1M0_2;
	wire w_dff_B_9F0VmLuT0_2;
	wire w_dff_B_njGHyIku0_2;
	wire w_dff_B_2xhwFLI90_2;
	wire w_dff_B_s1obosXv1_2;
	wire w_dff_B_E3TtFOE52_2;
	wire w_dff_B_mGGnLoVQ7_2;
	wire w_dff_B_lJggEX4b9_2;
	wire w_dff_B_OaSbouYj8_2;
	wire w_dff_B_HLrOsYkm2_2;
	wire w_dff_B_lTtlyRh95_2;
	wire w_dff_B_crmkhb9j1_2;
	wire w_dff_B_AmQhiB013_2;
	wire w_dff_B_iZLbhxoo7_2;
	wire w_dff_B_qwtc29Jh7_2;
	wire w_dff_B_nC1IgaNQ6_2;
	wire w_dff_B_OpapyPtB9_2;
	wire w_dff_B_tILYIIsp6_2;
	wire w_dff_B_sQjQBrpf0_2;
	wire w_dff_B_OG30zOvl3_2;
	wire w_dff_B_2NPYnQza8_2;
	wire w_dff_B_qEOmvMIj2_2;
	wire w_dff_B_ICMzF6Jr6_2;
	wire w_dff_B_X7xodnwm1_1;
	wire w_dff_B_nlXGNjIF6_1;
	wire w_dff_B_0NPQCha60_2;
	wire w_dff_B_n18SuO5a3_2;
	wire w_dff_B_t43B5j8c5_2;
	wire w_dff_B_F84NreC82_2;
	wire w_dff_B_AOkS4PYT5_2;
	wire w_dff_B_SmYUXrUs2_2;
	wire w_dff_B_AnSy7udP7_2;
	wire w_dff_B_S0RfVLwC6_2;
	wire w_dff_B_BDYfIA1O9_2;
	wire w_dff_B_haaLgri37_2;
	wire w_dff_B_cL3Pn4GH0_2;
	wire w_dff_B_J0Z3k1ML2_2;
	wire w_dff_B_EJoyquFC8_2;
	wire w_dff_B_ZDL4Brfd7_2;
	wire w_dff_B_TETDjt7T8_2;
	wire w_dff_B_knKaKNxA8_2;
	wire w_dff_B_9roTWaUf2_2;
	wire w_dff_B_EKtsm1xm8_2;
	wire w_dff_B_Z3xbjfB47_2;
	wire w_dff_B_8xkb2ZLw7_2;
	wire w_dff_B_29d2u9qo9_2;
	wire w_dff_B_irvvmkuX2_2;
	wire w_dff_B_oX2YHHF74_2;
	wire w_dff_B_uHYM0hIk7_2;
	wire w_dff_B_swMWQBmI5_2;
	wire w_dff_B_bogDKblD1_2;
	wire w_dff_B_WnXDne0P8_2;
	wire w_dff_B_gT2D0SUk3_2;
	wire w_dff_B_TgMPwA4Q2_2;
	wire w_dff_B_2yjlCh1N1_2;
	wire w_dff_B_rbD5szq79_2;
	wire w_dff_B_15H3kabV2_2;
	wire w_dff_B_fIMasrvF3_2;
	wire w_dff_B_0hxaG8rN4_2;
	wire w_dff_B_pwCNOjhA3_2;
	wire w_dff_B_ef7mrUa07_2;
	wire w_dff_B_D0bcy96T8_2;
	wire w_dff_B_7eP7DN1Y4_2;
	wire w_dff_B_rCVC8Nrv3_2;
	wire w_dff_B_SMQlLS9G7_2;
	wire w_dff_B_KwZlrEUg5_2;
	wire w_dff_B_8sU7tmQn6_2;
	wire w_dff_B_bUJCqNGF9_2;
	wire w_dff_B_wTpbPT1U3_2;
	wire w_dff_B_hvL0KFLo6_2;
	wire w_dff_B_tYBrYaQC0_2;
	wire w_dff_B_Q6sD4Qeb5_2;
	wire w_dff_B_wff3Dzjk0_2;
	wire w_dff_B_al9gX4Yh0_2;
	wire w_dff_B_0asvR0wp9_2;
	wire w_dff_B_D7XTMrYT5_2;
	wire w_dff_B_4zdIWGLF7_2;
	wire w_dff_B_mV09WgCd9_2;
	wire w_dff_B_OZxWyJjY5_2;
	wire w_dff_B_ExYSN7yU2_2;
	wire w_dff_B_OGkyOXb97_2;
	wire w_dff_B_bCIaheV48_2;
	wire w_dff_B_cAWOpRNm5_2;
	wire w_dff_B_ZtgcNjdf2_2;
	wire w_dff_B_PK76ddSN5_2;
	wire w_dff_B_rl7TjIv99_2;
	wire w_dff_B_lR7Wf5kq2_2;
	wire w_dff_B_EkuLaFIM1_2;
	wire w_dff_B_GLbYpbuX3_2;
	wire w_dff_B_QuGF6xXi6_2;
	wire w_dff_B_BR0o74Rc7_2;
	wire w_dff_B_Ktywyk4b1_2;
	wire w_dff_B_yK91rIF66_2;
	wire w_dff_B_Q9QehKZ13_2;
	wire w_dff_B_QohVCJko7_2;
	wire w_dff_B_bHbVmv3S5_2;
	wire w_dff_B_pPjyttP71_2;
	wire w_dff_B_UBiOOzAm4_2;
	wire w_dff_B_O76LVzGe3_2;
	wire w_dff_B_7ewJLvDw1_2;
	wire w_dff_B_ZKC0WEWM3_1;
	wire w_dff_B_BNC8kMfX0_2;
	wire w_dff_B_2AFvZx8t7_2;
	wire w_dff_B_vdvEouQM7_2;
	wire w_dff_B_hoio2uhr0_2;
	wire w_dff_B_iOV2Hjtg3_2;
	wire w_dff_B_IXm6Ny388_2;
	wire w_dff_B_2ukPKuky7_2;
	wire w_dff_B_tSSubhgk2_2;
	wire w_dff_B_Rc69CJUn5_2;
	wire w_dff_B_Xu3So4dr6_2;
	wire w_dff_B_DItVifN45_2;
	wire w_dff_B_eyvana3L5_2;
	wire w_dff_B_HLyMGbqo1_2;
	wire w_dff_B_O1tkoqEf2_2;
	wire w_dff_B_EfE2ysZA5_2;
	wire w_dff_B_0dS5CT4o2_2;
	wire w_dff_B_wXc8zhX84_2;
	wire w_dff_B_clctTt8x1_2;
	wire w_dff_B_WWG48nvQ1_2;
	wire w_dff_B_ez0DO1L38_2;
	wire w_dff_B_2CWKtBYO2_2;
	wire w_dff_B_oCquieuX0_2;
	wire w_dff_B_6yu15raF8_2;
	wire w_dff_B_nsPbGACH3_2;
	wire w_dff_B_4HnGiibP4_2;
	wire w_dff_B_B62lF1dI8_2;
	wire w_dff_B_cGkTm7iv7_2;
	wire w_dff_B_I1xc5ct55_2;
	wire w_dff_B_2h7iqjcF0_2;
	wire w_dff_B_0ZHmcmaX0_2;
	wire w_dff_B_FmNj1nCT7_2;
	wire w_dff_B_nGKmKZuY9_2;
	wire w_dff_B_2JtS07gc5_2;
	wire w_dff_B_pzdKgBdT1_2;
	wire w_dff_B_rdWGEVfD7_2;
	wire w_dff_B_4zw2Wckk3_1;
	wire w_dff_B_jpgEFxr40_1;
	wire w_dff_B_7FcKe92B1_2;
	wire w_dff_B_gt0Mjkak6_2;
	wire w_dff_B_6T9qt8P13_2;
	wire w_dff_B_NcJYkPxn7_2;
	wire w_dff_B_VDJSfolT0_2;
	wire w_dff_B_s9LaQPmQ2_2;
	wire w_dff_B_8tIsUzxP2_2;
	wire w_dff_B_7tuKtVzO5_2;
	wire w_dff_B_r6x1NBrr6_2;
	wire w_dff_B_08WEnwmU5_2;
	wire w_dff_B_Gcelk3Ma2_2;
	wire w_dff_B_UDEQTZPQ9_2;
	wire w_dff_B_S9xv1bjO3_2;
	wire w_dff_B_NFUzX4r40_2;
	wire w_dff_B_RC8upy0Y3_2;
	wire w_dff_B_UH0dkvVo6_2;
	wire w_dff_B_2dZ8ulhM2_2;
	wire w_dff_B_KyfxT94a6_2;
	wire w_dff_B_vVeQjTaB7_2;
	wire w_dff_B_fHdOZAZR9_2;
	wire w_dff_B_aQQlbn8U9_2;
	wire w_dff_B_Pemg0udW0_2;
	wire w_dff_B_gQLaWQFL5_2;
	wire w_dff_B_CUdGUCs62_2;
	wire w_dff_B_6RuOt6mp1_2;
	wire w_dff_B_AmNTbTcf3_2;
	wire w_dff_B_G0a8hd3Z7_2;
	wire w_dff_B_hYWoXIzD2_2;
	wire w_dff_B_tCIblQOO6_2;
	wire w_dff_B_zxD86mAu4_2;
	wire w_dff_B_5k0XQMr77_2;
	wire w_dff_B_j3hSLS2j5_2;
	wire w_dff_B_bvtdjLpj9_2;
	wire w_dff_B_hCIdtIQp0_2;
	wire w_dff_B_c9LG3Gxg3_2;
	wire w_dff_B_TBEWTNIU2_2;
	wire w_dff_B_9mjOgcBi6_2;
	wire w_dff_B_b8GU8LQn6_2;
	wire w_dff_B_055S17Mu4_2;
	wire w_dff_B_nglLsSAt2_2;
	wire w_dff_B_hs6kqYo93_2;
	wire w_dff_B_hcVUC0IR4_2;
	wire w_dff_B_1PL7pokc7_2;
	wire w_dff_B_Qf8KEaym9_2;
	wire w_dff_B_2jSFyZfJ7_2;
	wire w_dff_B_gZOxMbrp7_2;
	wire w_dff_B_v0vdtG773_2;
	wire w_dff_B_tvge0oW91_2;
	wire w_dff_B_sFk0Ya3X5_2;
	wire w_dff_B_rZVCU9z56_2;
	wire w_dff_B_YOGAjIAm8_2;
	wire w_dff_B_qwYDQuNE9_2;
	wire w_dff_B_3JTkb7hs3_2;
	wire w_dff_B_V4sVBbUs0_2;
	wire w_dff_B_iKiZRmR45_2;
	wire w_dff_B_7bkktzIr1_2;
	wire w_dff_B_5rD8c5gv0_2;
	wire w_dff_B_11dv5sD72_2;
	wire w_dff_B_4CrBkHdb8_2;
	wire w_dff_B_OMidsCf33_2;
	wire w_dff_B_BDBFFa2H9_2;
	wire w_dff_B_9wfcP7qg3_2;
	wire w_dff_B_9DcX31kt0_2;
	wire w_dff_B_SrBj10tN2_2;
	wire w_dff_B_M25pG8lK2_2;
	wire w_dff_B_kHchIEaa6_2;
	wire w_dff_B_UnfEEObK3_2;
	wire w_dff_B_5Ib0KJ6z6_1;
	wire w_dff_B_6mDeWR194_2;
	wire w_dff_B_e6VEtXIN7_2;
	wire w_dff_B_UCsQuMDI3_2;
	wire w_dff_B_JRcnFvYy4_2;
	wire w_dff_B_MFX8Wkw83_2;
	wire w_dff_B_mzGL6Rjl6_2;
	wire w_dff_B_WFH46CMZ3_2;
	wire w_dff_B_ge74TO3H0_2;
	wire w_dff_B_9nAkBgvF4_2;
	wire w_dff_B_tEkRrEQx5_2;
	wire w_dff_B_eYeKBaxX4_2;
	wire w_dff_B_shl8RVuo8_2;
	wire w_dff_B_vW9Omg9Y5_2;
	wire w_dff_B_mZFqtfPm4_2;
	wire w_dff_B_khDeRDKf5_2;
	wire w_dff_B_lLYUcJ0l3_2;
	wire w_dff_B_nDEpZeTr1_2;
	wire w_dff_B_oRanvpB28_2;
	wire w_dff_B_Xg6cKKdn8_2;
	wire w_dff_B_rUxF75Gh1_2;
	wire w_dff_B_lATFeJ7o8_2;
	wire w_dff_B_n1s3b0gx8_2;
	wire w_dff_B_xyvqGlYi3_2;
	wire w_dff_B_ZViB0PM44_2;
	wire w_dff_B_mzIA7bHb1_2;
	wire w_dff_B_LMxFCVxi2_2;
	wire w_dff_B_lKy1rCvA4_2;
	wire w_dff_B_MA7Um7Op1_2;
	wire w_dff_B_onbLRaAG6_2;
	wire w_dff_B_N7kavOKX5_2;
	wire w_dff_B_jdG9VyKO9_2;
	wire w_dff_B_LSNcCxB14_1;
	wire w_dff_B_vQjzTvuR7_1;
	wire w_dff_B_ibLykyi51_2;
	wire w_dff_B_s9QbUPPy4_2;
	wire w_dff_B_JkBdRdHn1_2;
	wire w_dff_B_4Jorb95c9_2;
	wire w_dff_B_1TCjGsp41_2;
	wire w_dff_B_mRbUQ3g31_2;
	wire w_dff_B_azAAQTRp2_2;
	wire w_dff_B_rzrCC7gD0_2;
	wire w_dff_B_Ruytk1vZ0_2;
	wire w_dff_B_XUH9uMB30_2;
	wire w_dff_B_MroiVKSx5_2;
	wire w_dff_B_Ta7dHKfX4_2;
	wire w_dff_B_pTwgOsb36_2;
	wire w_dff_B_DNcvXVLo1_2;
	wire w_dff_B_EYpDFgBa6_2;
	wire w_dff_B_do05VpS64_2;
	wire w_dff_B_VRyluxtt1_2;
	wire w_dff_B_TlAaYFG82_2;
	wire w_dff_B_Str4OJXp6_2;
	wire w_dff_B_JtTlxIsj9_2;
	wire w_dff_B_Pp8lzc4Y1_2;
	wire w_dff_B_RVJo6Cox1_2;
	wire w_dff_B_O5zsZdx58_2;
	wire w_dff_B_on58kIbA4_2;
	wire w_dff_B_mdLUZads8_2;
	wire w_dff_B_Y63PJbbi7_2;
	wire w_dff_B_dwipn1rX2_2;
	wire w_dff_B_GkoW1heP5_2;
	wire w_dff_B_3a0ws0L71_2;
	wire w_dff_B_6GyjjIVl4_2;
	wire w_dff_B_IGZpL0219_2;
	wire w_dff_B_XEpzRJvB0_2;
	wire w_dff_B_6sXv0xHP5_2;
	wire w_dff_B_A9yybFE71_2;
	wire w_dff_B_8k5jswkw5_2;
	wire w_dff_B_J8DRx8WX8_2;
	wire w_dff_B_eyLxlTuN3_2;
	wire w_dff_B_IF5onHPo3_2;
	wire w_dff_B_ULKHogEp3_2;
	wire w_dff_B_o5MC7lmz3_2;
	wire w_dff_B_Egf9GCyA2_2;
	wire w_dff_B_Wp0eq3h40_2;
	wire w_dff_B_UTino0ZK6_2;
	wire w_dff_B_xNTmY2ne4_2;
	wire w_dff_B_mt0QN3742_2;
	wire w_dff_B_RU52QQuH0_2;
	wire w_dff_B_6Ccp02qV8_2;
	wire w_dff_B_zVrLvjrx1_2;
	wire w_dff_B_hPaFveAv8_2;
	wire w_dff_B_lTKs7F450_2;
	wire w_dff_B_4fYwJyMx9_2;
	wire w_dff_B_cVcvy8Hg7_2;
	wire w_dff_B_KIGlNau69_2;
	wire w_dff_B_1PfSOphx1_2;
	wire w_dff_B_g8nA3w162_2;
	wire w_dff_B_QT5HnJV77_2;
	wire w_dff_B_ounjcS661_2;
	wire w_dff_B_irSCcU5R7_2;
	wire w_dff_B_24k6eYsp4_2;
	wire w_dff_B_eVn4YkX40_1;
	wire w_dff_B_bcA32Be96_2;
	wire w_dff_B_12jGT5iy4_2;
	wire w_dff_B_mXjMtn4r1_2;
	wire w_dff_B_zEStQkLn0_2;
	wire w_dff_B_Oju0jybA7_2;
	wire w_dff_B_kZEymnYy2_2;
	wire w_dff_B_9Kv2D6ss0_2;
	wire w_dff_B_To2LDRTW2_2;
	wire w_dff_B_DRh7zhKd8_2;
	wire w_dff_B_ZrLYkahn4_2;
	wire w_dff_B_7om8xK6W1_2;
	wire w_dff_B_juQnec570_2;
	wire w_dff_B_llXl76rH8_2;
	wire w_dff_B_nczVXYaZ6_2;
	wire w_dff_B_CgQ9lM237_2;
	wire w_dff_B_H4rYk0z34_2;
	wire w_dff_B_MtpIjnst4_2;
	wire w_dff_B_d2bQqD3o7_2;
	wire w_dff_B_c0lx2f367_2;
	wire w_dff_B_VnXblzEc8_2;
	wire w_dff_B_acjOKS6m0_2;
	wire w_dff_B_OKCdYD7p1_2;
	wire w_dff_B_6pmO231M2_2;
	wire w_dff_B_11lJgs1H3_2;
	wire w_dff_B_7htPfhn37_2;
	wire w_dff_B_MEA4sZFM7_2;
	wire w_dff_B_cqr3P2Ay4_2;
	wire w_dff_B_mGTa7ymT7_1;
	wire w_dff_B_meQsglwa0_1;
	wire w_dff_B_WyQdZu1G7_2;
	wire w_dff_B_oBi0Ul3v7_2;
	wire w_dff_B_10I6NcpG1_2;
	wire w_dff_B_dAoGwnK16_2;
	wire w_dff_B_llaNNY9k5_2;
	wire w_dff_B_0yrPQEYH1_2;
	wire w_dff_B_S8UkZmQP4_2;
	wire w_dff_B_yCnypHLG3_2;
	wire w_dff_B_zAvpxqvI1_2;
	wire w_dff_B_q98XcGyK4_2;
	wire w_dff_B_swfoPuTx3_2;
	wire w_dff_B_eAFofZcY0_2;
	wire w_dff_B_n1LLCpb47_2;
	wire w_dff_B_swi9ghk14_2;
	wire w_dff_B_Rs0wV5UK9_2;
	wire w_dff_B_99iUJNDd3_2;
	wire w_dff_B_3fH8X0Og1_2;
	wire w_dff_B_I6TdlgN36_2;
	wire w_dff_B_hmCv5Pzt1_2;
	wire w_dff_B_Dq9MvurV8_2;
	wire w_dff_B_3xe1moFK4_2;
	wire w_dff_B_zKPuNROK4_2;
	wire w_dff_B_OQdcmkcf5_2;
	wire w_dff_B_x0NmA8Gt4_2;
	wire w_dff_B_1yjvzkdL5_2;
	wire w_dff_B_Ijjsn1bS6_2;
	wire w_dff_B_p0bRLz0k3_2;
	wire w_dff_B_wrgEB7nz3_2;
	wire w_dff_B_8VbBVnmX6_2;
	wire w_dff_B_6kBtE20E3_2;
	wire w_dff_B_CW53KMFZ8_2;
	wire w_dff_B_UsQPoqyH9_2;
	wire w_dff_B_XO43nQfU9_2;
	wire w_dff_B_Y4MTR1hm7_2;
	wire w_dff_B_nu9ZHmxk8_2;
	wire w_dff_B_Xg0YCQo83_2;
	wire w_dff_B_JFMTEVnT9_2;
	wire w_dff_B_MZkzplGT3_2;
	wire w_dff_B_tMWkEoQz2_2;
	wire w_dff_B_JOlqMAD76_2;
	wire w_dff_B_TW2E4hbb8_2;
	wire w_dff_B_7r5Qeh8O9_2;
	wire w_dff_B_ZXZrfq8x5_2;
	wire w_dff_B_f18JwbVl1_2;
	wire w_dff_B_XNgtLl0o0_2;
	wire w_dff_B_erCkOw5d8_2;
	wire w_dff_B_VVeSMAgY2_2;
	wire w_dff_B_0XNddVoS8_2;
	wire w_dff_B_6N6dtyd68_2;
	wire w_dff_B_zZeO24ZO9_2;
	wire w_dff_B_mAl5mvvM9_2;
	wire w_dff_B_MiHFayT22_1;
	wire w_dff_B_6zRCsN5I2_2;
	wire w_dff_B_hmc8dgcw6_2;
	wire w_dff_B_siPT53r59_2;
	wire w_dff_B_M5VmMrFx9_2;
	wire w_dff_B_MSfkfmxL6_2;
	wire w_dff_B_AqV1lGGE3_2;
	wire w_dff_B_IwUBOxKk4_2;
	wire w_dff_B_QxY2O6uL2_2;
	wire w_dff_B_pnjtYi0U3_2;
	wire w_dff_B_GQwWV3tM8_2;
	wire w_dff_B_2FJrH1991_2;
	wire w_dff_B_53qjY3DZ7_2;
	wire w_dff_B_tWS8GqNM7_2;
	wire w_dff_B_Ncememkz1_2;
	wire w_dff_B_H27Ncgy10_2;
	wire w_dff_B_Zu0aLVpB7_2;
	wire w_dff_B_cBJZNKeD1_2;
	wire w_dff_B_R0xnnk9L3_2;
	wire w_dff_B_QYyFxlef0_2;
	wire w_dff_B_AFaUlWWF0_2;
	wire w_dff_B_NeAUwhoJ1_2;
	wire w_dff_B_YBQHYPJ85_2;
	wire w_dff_B_N0Tsv9Tp0_2;
	wire w_dff_B_5LwBCvTA9_1;
	wire w_dff_B_2UYJmSWs0_1;
	wire w_dff_B_yBjCL9c09_2;
	wire w_dff_B_WiLuKK9K3_2;
	wire w_dff_B_QAyQGM3A2_2;
	wire w_dff_B_wqT00hx83_2;
	wire w_dff_B_fBfICTYq0_2;
	wire w_dff_B_6HAJBTrF0_2;
	wire w_dff_B_FBM7TZ6n2_2;
	wire w_dff_B_3kmW9Kiy3_2;
	wire w_dff_B_4ikPSIaQ3_2;
	wire w_dff_B_udyCn42C1_2;
	wire w_dff_B_ocRjkFt70_2;
	wire w_dff_B_bPEcba2J5_2;
	wire w_dff_B_CTYdPjno3_2;
	wire w_dff_B_tMLHx8p98_2;
	wire w_dff_B_A0wU6i6D4_2;
	wire w_dff_B_mHjUDGzn5_2;
	wire w_dff_B_1nUWKe6m7_2;
	wire w_dff_B_6Li8uaB89_2;
	wire w_dff_B_AGZPkQLo8_2;
	wire w_dff_B_Lwcvv2XE9_2;
	wire w_dff_B_Y5Gh3Yym8_2;
	wire w_dff_B_zXbVV5OP3_2;
	wire w_dff_B_ls6NnuRX6_2;
	wire w_dff_B_wVoB6uRS9_2;
	wire w_dff_B_iirIfLG89_2;
	wire w_dff_B_IXb9wSKN3_2;
	wire w_dff_B_Igk4Mib62_2;
	wire w_dff_B_ZjaErCCv8_2;
	wire w_dff_B_bcPIvtUJ4_2;
	wire w_dff_B_hvdYaCEX5_2;
	wire w_dff_B_gW63nihM1_2;
	wire w_dff_B_fpEvUovD7_2;
	wire w_dff_B_SksLlSMZ9_2;
	wire w_dff_B_SSuJn0qK5_2;
	wire w_dff_B_aV4EAW3S3_2;
	wire w_dff_B_uM4aMKp82_2;
	wire w_dff_B_hAc2qsIN2_2;
	wire w_dff_B_Hy3qaCsF0_2;
	wire w_dff_B_IEPpiw0e2_2;
	wire w_dff_B_CMeRreZc7_2;
	wire w_dff_B_H42GKPi99_2;
	wire w_dff_B_lQleofwo6_2;
	wire w_dff_B_mB60qQA78_2;
	wire w_dff_B_7k9iJ5tT6_1;
	wire w_dff_B_SK7ixJDL3_2;
	wire w_dff_B_sR0uFpe75_2;
	wire w_dff_B_WGOTq29G5_2;
	wire w_dff_B_iDHRGbm33_2;
	wire w_dff_B_c6Mhr2Ba4_2;
	wire w_dff_B_zAsTsVJR7_2;
	wire w_dff_B_rp6kxHkv3_2;
	wire w_dff_B_mzWakkxk3_2;
	wire w_dff_B_azXYWqpz2_2;
	wire w_dff_B_nb8owcxN6_2;
	wire w_dff_B_PHbfqBnV0_2;
	wire w_dff_B_Cn08fwCC5_2;
	wire w_dff_B_IiyBCTar5_2;
	wire w_dff_B_ne1Iznhr2_2;
	wire w_dff_B_BFgKVyXo3_2;
	wire w_dff_B_U0JDzBCI0_2;
	wire w_dff_B_HPMWVqFw8_2;
	wire w_dff_B_gZGtd2Gi4_2;
	wire w_dff_B_rOjuu2xq3_2;
	wire w_dff_B_YPFpbhph5_1;
	wire w_dff_B_DCPQC2Kw1_1;
	wire w_dff_B_WEHEShuh7_2;
	wire w_dff_B_t7WOkIAn1_2;
	wire w_dff_B_TBKjdZve0_2;
	wire w_dff_B_mZJxy1Tw7_2;
	wire w_dff_B_7GGeUX2V7_2;
	wire w_dff_B_itFfMoP16_2;
	wire w_dff_B_N6cZe30a7_2;
	wire w_dff_B_8RBPbisT3_2;
	wire w_dff_B_tqzRjAZo4_2;
	wire w_dff_B_0h8o1GjY6_2;
	wire w_dff_B_puAnTaMN9_2;
	wire w_dff_B_nJi0isK64_2;
	wire w_dff_B_iMRQ4lTU9_2;
	wire w_dff_B_gM7jwQeG7_2;
	wire w_dff_B_eIEwx81R7_2;
	wire w_dff_B_WTdmoGjV0_2;
	wire w_dff_B_Hhmpk3g62_2;
	wire w_dff_B_AKrMBL1h4_2;
	wire w_dff_B_fBgfm8bz8_2;
	wire w_dff_B_AdgTnOUt5_2;
	wire w_dff_B_dFoGbecY3_2;
	wire w_dff_B_qX1pOQzH7_2;
	wire w_dff_B_ZMKitu0y7_2;
	wire w_dff_B_9iVniqH93_2;
	wire w_dff_B_s7Y9Kv6W2_2;
	wire w_dff_B_fxrp6rHV6_2;
	wire w_dff_B_6soAIcis3_2;
	wire w_dff_B_EFZBgCdr0_2;
	wire w_dff_B_MK3I8beV8_2;
	wire w_dff_B_EBLi6mFi8_2;
	wire w_dff_B_UIuPmVgr4_2;
	wire w_dff_B_osNrJkuP9_2;
	wire w_dff_B_Uptxipqr6_2;
	wire w_dff_B_aWfsZ3VJ7_2;
	wire w_dff_B_RvqdFM2d3_2;
	wire w_dff_B_0Gb9Fong5_1;
	wire w_dff_B_g3Irwatn0_2;
	wire w_dff_B_S0Gbhlc82_2;
	wire w_dff_B_gU5NsR8t5_2;
	wire w_dff_B_b35qg5Y62_2;
	wire w_dff_B_aEIJ8oQw6_2;
	wire w_dff_B_yzTLXsOn9_2;
	wire w_dff_B_lMm3TnGF6_2;
	wire w_dff_B_saLKSXE94_2;
	wire w_dff_B_G6WDknzh2_2;
	wire w_dff_B_PQySZ21H7_2;
	wire w_dff_B_ud3fYL8c4_2;
	wire w_dff_B_iaSJi1CZ6_2;
	wire w_dff_B_6asxB7TE8_2;
	wire w_dff_B_y7WuCpIE4_2;
	wire w_dff_B_FD98udlP0_2;
	wire w_dff_B_d372Oo5A1_2;
	wire w_dff_B_hyelq2598_2;
	wire w_dff_B_JYpE4nrd8_2;
	wire w_dff_B_jjdl1HXT5_2;
	wire w_dff_B_1JzSWLQv2_2;
	wire w_dff_B_JtxHj3i14_2;
	wire w_dff_B_AahmCqvJ0_2;
	wire w_dff_B_igypnapb5_2;
	wire w_dff_B_w3A1wWQ14_2;
	wire w_dff_B_tweRq4vJ5_2;
	wire w_dff_B_Mi5d83Fo4_2;
	wire w_dff_B_0sA4WOD92_2;
	wire w_dff_B_XVO8klnG6_2;
	wire w_dff_B_T5A98wyQ2_2;
	wire w_dff_B_95UCo4TK0_2;
	wire w_dff_B_KQWddzh79_2;
	wire w_dff_B_sjtr7rUO1_2;
	wire w_dff_B_L7oXhL0G3_2;
	wire w_dff_B_38xMc8u08_2;
	wire w_dff_B_26EDGsq77_2;
	wire w_dff_B_xYulOIww0_2;
	wire w_dff_B_TV9oSqo39_2;
	wire w_dff_B_lnBUZir81_2;
	wire w_dff_B_f4sHwQoT5_2;
	wire w_dff_B_rHvJMzyq5_2;
	wire w_dff_B_fr1DhGc09_2;
	wire w_dff_B_lu06mhQM1_2;
	wire w_dff_B_eYIqDh9G5_1;
	wire w_dff_B_lPV6Fhfl4_2;
	wire w_dff_B_ixrbUdjT3_2;
	wire w_dff_B_HtZglrRJ8_2;
	wire w_dff_B_ZSq65Qju7_2;
	wire w_dff_B_CbjeNfc21_2;
	wire w_dff_B_dl6SEOlw9_2;
	wire w_dff_B_thHIcPAa4_2;
	wire w_dff_B_7vDaRG5I2_2;
	wire w_dff_B_Wg7xHT2A3_2;
	wire w_dff_B_f3hvHBZV4_2;
	wire w_dff_B_fsycHxs66_2;
	wire w_dff_A_RhDR8iYU1_0;
	wire w_dff_A_MC7RPwqJ2_0;
	wire w_dff_A_WmXhKVT75_0;
	wire w_dff_B_qHewBVZt4_2;
	wire w_dff_B_V60rxirR2_1;
	wire w_dff_B_kbzGUNAt3_1;
	wire w_dff_B_suLSGBXS0_1;
	wire w_dff_B_ML2YcFrR7_1;
	wire w_dff_B_wgj4zyG66_1;
	wire w_dff_B_rP85qQ8J0_1;
	wire w_dff_B_NVAwxQ8j6_1;
	wire w_dff_B_hodFMUDZ4_1;
	wire w_dff_A_WKPsJg287_1;
	wire w_dff_A_tI8ZURF34_1;
	wire w_dff_A_xPZGakul1_1;
	wire w_dff_A_MEwpgw3j7_1;
	wire w_dff_A_d5cPW0z26_1;
	wire w_dff_A_uPuFJxVi0_1;
	wire w_dff_A_RSjd2ENx5_1;
	wire w_dff_B_VdZF60TW4_2;
	wire w_dff_B_k1MB6W6t7_2;
	wire w_dff_B_gRaz6dBT7_2;
	wire w_dff_B_H79v9Uq58_2;
	wire w_dff_B_Imlk7Eki1_2;
	wire w_dff_B_hxtgEtn99_2;
	wire w_dff_B_S1QBbm186_2;
	wire w_dff_B_pkHOALHt4_2;
	wire w_dff_B_hlGenjoK5_2;
	wire w_dff_B_jaHXtSYv4_2;
	wire w_dff_B_BFY5D3Vg9_1;
	wire w_dff_B_m910XB5j8_2;
	wire w_dff_B_vzdzVgz41_2;
	wire w_dff_B_20BlkzZ02_2;
	wire w_dff_B_z58mmzRV5_2;
	wire w_dff_B_KocCuaqj5_2;
	wire w_dff_B_Y3yudIDv2_2;
	wire w_dff_B_hgcUEBts6_2;
	wire w_dff_B_N8ucdRpL4_2;
	wire w_dff_B_rjpJ8Lqi1_2;
	wire w_dff_B_S3wHjT2K0_2;
	wire w_dff_B_7hsdjXtW4_2;
	wire w_dff_B_9vzWDEwn2_2;
	wire w_dff_B_l45lPUQS4_2;
	wire w_dff_A_08zg0qyi5_0;
	wire w_dff_A_pMFqqMNj9_0;
	wire w_dff_A_8xMT58BS1_0;
	wire w_dff_A_SZgnYqYp9_0;
	wire w_dff_A_tkYEQ15O7_1;
	wire w_dff_A_RxpTO1Zh9_1;
	wire w_dff_B_0mee9hQv7_1;
	wire w_dff_B_l0KD2s4z2_1;
	wire w_dff_B_oZbFmwUg7_1;
	wire w_dff_B_DCx1VC6Y7_1;
	wire w_dff_B_rf367TDu7_1;
	wire w_dff_A_mlAWXDW60_0;
	wire w_dff_A_rfFuhg8h4_0;
	wire w_dff_A_YjJMEe3C2_0;
	wire w_dff_A_a9Fc5BLn6_0;
	wire w_dff_A_bmzQ5Z6I6_0;
	wire w_dff_A_reLcFVwy2_0;
	wire w_dff_B_9nAcROIB4_2;
	wire w_dff_A_465exy0V6_1;
	wire w_dff_A_lZyKX5BD7_1;
	wire w_dff_A_Tg2TvWQO4_1;
	wire w_dff_A_TuVbJBvl8_1;
	wire w_dff_A_8hSQ65zN0_1;
	wire w_dff_A_OnSTmqyq1_1;
	wire w_dff_A_u8sRXF6f7_0;
	wire w_dff_A_O7IBO4CG5_0;
	wire w_dff_A_uBqUbjxD5_0;
	wire w_dff_A_QnjCtdwm1_0;
	wire w_dff_A_aRGGjZYo6_0;
	wire w_dff_A_RjIseovg1_0;
	wire w_dff_A_wERotExv1_0;
	wire w_dff_A_0gYpOujG3_0;
	wire w_dff_A_dyyIoITs1_0;
	wire w_dff_A_IRObgaE56_0;
	wire w_dff_A_nQZ1IWK35_0;
	wire w_dff_A_TZ2Sz1g82_0;
	wire w_dff_A_IjEeqSlc8_0;
	wire w_dff_A_a5zOXXRW9_0;
	wire w_dff_A_UgOeq3E74_0;
	wire w_dff_A_YhIT9Jj34_0;
	wire w_dff_A_vpMQtO4F4_0;
	wire w_dff_A_ipGv5gIj3_0;
	wire w_dff_A_FbGLY1V18_0;
	wire w_dff_A_7DRm5FfY8_0;
	wire w_dff_A_kbvrLwRX2_0;
	wire w_dff_A_Wkw9DGp21_0;
	wire w_dff_A_UvEGBe7f5_0;
	wire w_dff_A_nRvBmrCg1_0;
	wire w_dff_A_SPsbKPKH1_0;
	wire w_dff_A_eVTDbam93_0;
	wire w_dff_A_Wt9gVfJI8_0;
	wire w_dff_A_Eiz2eeZs1_0;
	wire w_dff_A_R3afGlWJ6_0;
	wire w_dff_A_CdI7CRYe4_0;
	wire w_dff_A_KkAMD7Cx9_0;
	wire w_dff_A_li4NKrln5_0;
	wire w_dff_A_oqjCF0In6_0;
	wire w_dff_A_FE5wqB124_0;
	wire w_dff_A_4R16xZrH7_0;
	wire w_dff_A_LJOV3Lxx9_0;
	wire w_dff_A_MGOwzsVF3_0;
	wire w_dff_A_lyksgwbU2_0;
	wire w_dff_A_86477Pek7_0;
	wire w_dff_A_c54GyUP38_0;
	wire w_dff_A_mASEeWWt9_0;
	wire w_dff_A_mj9Fs4110_0;
	wire w_dff_A_0Jazty1V2_0;
	wire w_dff_A_WHN79rNy5_0;
	wire w_dff_A_4lCsJIWU6_0;
	wire w_dff_A_dE0hqBcc4_0;
	wire w_dff_A_Ls5lsSD16_0;
	wire w_dff_A_vwyglYq09_0;
	wire w_dff_A_kFViTijJ7_0;
	wire w_dff_A_vPsWXsLZ0_0;
	wire w_dff_A_is7H95T40_0;
	wire w_dff_A_mXrHs79t9_0;
	wire w_dff_A_hKa7peHF0_0;
	wire w_dff_A_8dxI3AM84_0;
	wire w_dff_A_iuYQRbip0_0;
	wire w_dff_A_KnGhanup8_0;
	wire w_dff_A_qEq9LsPR5_0;
	wire w_dff_A_hIjfV8Al0_0;
	wire w_dff_A_I3bJZEvu1_0;
	wire w_dff_A_VJfYeyLo8_0;
	wire w_dff_A_rR5XOtlX0_0;
	wire w_dff_A_P7RDMqrv4_0;
	wire w_dff_A_Yw1rUEkr6_0;
	wire w_dff_A_8pWPZ5so7_0;
	wire w_dff_A_TCKFPob91_0;
	wire w_dff_A_iXOKyWzx4_0;
	wire w_dff_A_y4qfZ9Im3_0;
	wire w_dff_A_ZaDG8Mq34_0;
	wire w_dff_A_W1qK3Myh1_0;
	wire w_dff_A_MbeK9Jcu1_0;
	wire w_dff_A_54b37qpb1_0;
	wire w_dff_A_2Efcu3yJ9_0;
	wire w_dff_A_JQbFPgSh8_0;
	wire w_dff_A_nW1ypwyI6_0;
	wire w_dff_A_7d1LhOvD7_2;
	wire w_dff_A_rvczDX1L2_0;
	wire w_dff_A_sLsmbTZ66_0;
	wire w_dff_A_Wg7qmMMc2_0;
	wire w_dff_A_QWAcJONC2_0;
	wire w_dff_A_NXbXGzJ11_0;
	wire w_dff_A_LNGtkm7A0_0;
	wire w_dff_A_v03aTqCa8_0;
	wire w_dff_A_PvXQ8A7N6_0;
	wire w_dff_A_Rg34ntno7_0;
	wire w_dff_A_tJHxOajH5_0;
	wire w_dff_A_b9E0guGl5_0;
	wire w_dff_A_lw1IlMQZ0_0;
	wire w_dff_A_mYcqDf071_0;
	wire w_dff_A_RiVu5ex30_0;
	wire w_dff_A_IL7RVIdG0_0;
	wire w_dff_A_Goycacxx8_0;
	wire w_dff_A_opmy3WvA4_0;
	wire w_dff_A_jVbglBum3_0;
	wire w_dff_A_Ac8D5KiO0_0;
	wire w_dff_A_RZowy2XY7_0;
	wire w_dff_A_KqatYKAM2_0;
	wire w_dff_A_iI9MGEWT4_0;
	wire w_dff_A_wHGDIevi8_0;
	wire w_dff_A_wKkHWfzP7_0;
	wire w_dff_A_kUIoZqy33_0;
	wire w_dff_A_A78dhmsf1_0;
	wire w_dff_A_gIJTDeFf4_0;
	wire w_dff_A_RiCB1H3h2_0;
	wire w_dff_A_lOI8om2V0_0;
	wire w_dff_A_bNW4aXBV0_0;
	wire w_dff_A_K3xSEreo1_0;
	wire w_dff_A_dVCcKt8d7_0;
	wire w_dff_A_3C7lMoD16_0;
	wire w_dff_A_8iyDK62l3_0;
	wire w_dff_A_TB05FPcS2_0;
	wire w_dff_A_YY1ktvQR6_0;
	wire w_dff_A_8xwuFCjV3_0;
	wire w_dff_A_8TjjNzAq3_0;
	wire w_dff_A_H1WrmOOh5_0;
	wire w_dff_A_F1bXCwum3_0;
	wire w_dff_A_czNI0Agy8_0;
	wire w_dff_A_SE8FeqzN4_0;
	wire w_dff_A_CWiZwwt58_0;
	wire w_dff_A_i7kBb1Zc1_0;
	wire w_dff_A_3OHjbTN80_0;
	wire w_dff_A_nhDOU8Jb7_0;
	wire w_dff_A_80FsTp2J1_0;
	wire w_dff_A_bu4DrZPu4_0;
	wire w_dff_A_AyJjQC3H0_0;
	wire w_dff_A_8EacnzDo2_0;
	wire w_dff_A_wB3jjJIo3_0;
	wire w_dff_A_oR9lj3Cj3_0;
	wire w_dff_A_NjBX5f7n4_0;
	wire w_dff_A_6d6rJqBF1_0;
	wire w_dff_A_NrdAXYeZ4_0;
	wire w_dff_A_8bGzGdwd0_0;
	wire w_dff_A_o2tMKMkp2_0;
	wire w_dff_A_8jEqjpPQ3_0;
	wire w_dff_A_w3gmyqSr3_0;
	wire w_dff_A_NFynntpd8_0;
	wire w_dff_A_1lAAMchZ3_0;
	wire w_dff_A_Ne5boROJ6_0;
	wire w_dff_A_dGOd6PBg2_0;
	wire w_dff_A_S0SUIxPg2_0;
	wire w_dff_A_jRb1ubOH0_0;
	wire w_dff_A_IInP2Buv4_0;
	wire w_dff_A_eOqaNz979_0;
	wire w_dff_A_p7U3kNJM0_0;
	wire w_dff_A_jtKUE8BM5_0;
	wire w_dff_A_BkkyqPNt8_0;
	wire w_dff_A_bZQbIqBj5_0;
	wire w_dff_A_e8HaFF4D6_2;
	wire w_dff_A_ZZg83iRK9_0;
	wire w_dff_A_1ELkWDTe3_0;
	wire w_dff_A_vnFrLtHI5_0;
	wire w_dff_A_oDQXVNpp3_0;
	wire w_dff_A_mdfKnGhh8_0;
	wire w_dff_A_O3K9QHJD2_0;
	wire w_dff_A_2BX4wbWT0_0;
	wire w_dff_A_ixwumU436_0;
	wire w_dff_A_tR5rl26t7_0;
	wire w_dff_A_AH08WWq24_0;
	wire w_dff_A_dX3eqge23_0;
	wire w_dff_A_zVugR1mv3_0;
	wire w_dff_A_JiBEC2kq1_0;
	wire w_dff_A_DSkflptN6_0;
	wire w_dff_A_1cydg5nh3_0;
	wire w_dff_A_KD3R02fk3_0;
	wire w_dff_A_Ntnv9MjG3_0;
	wire w_dff_A_NWqy4acc9_0;
	wire w_dff_A_i4GF1qP82_0;
	wire w_dff_A_lIzvw1CS9_0;
	wire w_dff_A_JwLov5Xj2_0;
	wire w_dff_A_zL6EUY6B3_0;
	wire w_dff_A_sACBSGvS2_0;
	wire w_dff_A_rObrAbyh5_0;
	wire w_dff_A_F8mBgC9n2_0;
	wire w_dff_A_Pzjv24El2_0;
	wire w_dff_A_Aif2BL8Q7_0;
	wire w_dff_A_WDTI2AWs7_0;
	wire w_dff_A_QMehkqT62_0;
	wire w_dff_A_Y8lwrufa9_0;
	wire w_dff_A_2nP9Ufdi4_0;
	wire w_dff_A_9ftYyt6u2_0;
	wire w_dff_A_kWSAGsnT8_0;
	wire w_dff_A_32jPwhUT7_0;
	wire w_dff_A_fkZe9YOD5_0;
	wire w_dff_A_dimGw5UX6_0;
	wire w_dff_A_kW56nKPb5_0;
	wire w_dff_A_lyDQ4kJU5_0;
	wire w_dff_A_eh7A5qZo0_0;
	wire w_dff_A_c3Pnpf1J1_0;
	wire w_dff_A_VDThfbob4_0;
	wire w_dff_A_3GIsObAc5_0;
	wire w_dff_A_9YWWJm5T3_0;
	wire w_dff_A_ZXVFgdLK3_0;
	wire w_dff_A_o4gPJLkS2_0;
	wire w_dff_A_FNTkhPLx7_0;
	wire w_dff_A_1dfbKyYl6_0;
	wire w_dff_A_NkXw6eyl4_0;
	wire w_dff_A_LhDLpsCR0_0;
	wire w_dff_A_kR2dOtYY0_0;
	wire w_dff_A_NmTd3ng58_0;
	wire w_dff_A_ApbI0e9z0_0;
	wire w_dff_A_nj1SBpVm6_0;
	wire w_dff_A_7OoIpG8y9_0;
	wire w_dff_A_pXZbzZkY2_0;
	wire w_dff_A_fNoTmXkC1_0;
	wire w_dff_A_vnDR5rbC2_0;
	wire w_dff_A_SbuqzeQm8_0;
	wire w_dff_A_gVE3prvY1_0;
	wire w_dff_A_fVXq8srf3_0;
	wire w_dff_A_6ZPVnYmI2_0;
	wire w_dff_A_wpIIYxmW6_0;
	wire w_dff_A_IJVHL4aj9_0;
	wire w_dff_A_2xVWeuRV3_0;
	wire w_dff_A_W3WCDQQi3_0;
	wire w_dff_A_A7eHw9W44_0;
	wire w_dff_A_pgrOyBBg0_0;
	wire w_dff_A_DmqY5Xux5_0;
	wire w_dff_A_Q4wViHZO3_2;
	wire w_dff_A_UKGyNndE4_0;
	wire w_dff_A_qUeEvSGB0_0;
	wire w_dff_A_uUFbC5Eb7_0;
	wire w_dff_A_ABV271t69_0;
	wire w_dff_A_LhK1w2Fz8_0;
	wire w_dff_A_0xGoPeYp4_0;
	wire w_dff_A_LbJY9ZJz3_0;
	wire w_dff_A_rO1PLAT97_0;
	wire w_dff_A_Rn1PcijY6_0;
	wire w_dff_A_VbOZqn9n0_0;
	wire w_dff_A_Kqcb5LSI4_0;
	wire w_dff_A_IE7xaUEc8_0;
	wire w_dff_A_QsSa10gD7_0;
	wire w_dff_A_CemuLbpo5_0;
	wire w_dff_A_cYpjudqf8_0;
	wire w_dff_A_uS62HLbT8_0;
	wire w_dff_A_aAITNGHM8_0;
	wire w_dff_A_c7WM03iH2_0;
	wire w_dff_A_VMVN8ZTE0_0;
	wire w_dff_A_edAnMSk69_0;
	wire w_dff_A_5bGqQTTI1_0;
	wire w_dff_A_qxJQYNKX9_0;
	wire w_dff_A_zqH6VjWv6_0;
	wire w_dff_A_fFlxY9z75_0;
	wire w_dff_A_lVbwfm9p1_0;
	wire w_dff_A_wIgw8zl50_0;
	wire w_dff_A_VyzX67HB0_0;
	wire w_dff_A_YZXJXWSo8_0;
	wire w_dff_A_oPgPigwE1_0;
	wire w_dff_A_l47orzlV2_0;
	wire w_dff_A_CTRyvGVw5_0;
	wire w_dff_A_wy5wa6GW2_0;
	wire w_dff_A_FJ4FBgg43_0;
	wire w_dff_A_wWjU7aGC3_0;
	wire w_dff_A_pnMt5kN98_0;
	wire w_dff_A_Z0KSpMFG3_0;
	wire w_dff_A_k9nttZJ53_0;
	wire w_dff_A_8oN7L5TL1_0;
	wire w_dff_A_KQvu6Vn18_0;
	wire w_dff_A_mO4b9Xv36_0;
	wire w_dff_A_Gqpo25ko8_0;
	wire w_dff_A_OiJChVz76_0;
	wire w_dff_A_0oUw4awM1_0;
	wire w_dff_A_BUIBv3MN7_0;
	wire w_dff_A_510i0Ffj1_0;
	wire w_dff_A_63jS389e1_0;
	wire w_dff_A_jK0spGO02_0;
	wire w_dff_A_PylGZhxj8_0;
	wire w_dff_A_OLtjmGcU0_0;
	wire w_dff_A_wCqrIRxR5_0;
	wire w_dff_A_ByPe0qEa0_0;
	wire w_dff_A_NzPsVdYV3_0;
	wire w_dff_A_Ld4GxZ712_0;
	wire w_dff_A_Jio3chGL5_0;
	wire w_dff_A_Evu8NZnU2_0;
	wire w_dff_A_FnrptbQf6_0;
	wire w_dff_A_GcCGrIZl5_0;
	wire w_dff_A_jZ55oJcH8_0;
	wire w_dff_A_PyPE5ikt1_0;
	wire w_dff_A_E5PSy3W04_0;
	wire w_dff_A_bm2wDxTQ4_0;
	wire w_dff_A_BK8ocyvE5_0;
	wire w_dff_A_gJzrV2Jq6_0;
	wire w_dff_A_2eqOwn7e3_0;
	wire w_dff_A_0zBuhWTA2_0;
	wire w_dff_A_b8H84EUd8_2;
	wire w_dff_A_TfOUa18I0_0;
	wire w_dff_A_kOYBWUmp5_0;
	wire w_dff_A_OsZUU0qz7_0;
	wire w_dff_A_EnPSnzTH3_0;
	wire w_dff_A_p5HfxFzY9_0;
	wire w_dff_A_R6DcDzhx9_0;
	wire w_dff_A_TBEkWVCz0_0;
	wire w_dff_A_mjo7B4Fa6_0;
	wire w_dff_A_DOHeVL7p1_0;
	wire w_dff_A_jTxufXdv3_0;
	wire w_dff_A_PrAnHZNC9_0;
	wire w_dff_A_hgyb57m38_0;
	wire w_dff_A_1yimvYdx1_0;
	wire w_dff_A_pq0AN4Bz7_0;
	wire w_dff_A_S5TbOQHk3_0;
	wire w_dff_A_tE7M3Alx8_0;
	wire w_dff_A_a9cnZ2ms4_0;
	wire w_dff_A_H1HuJkNV0_0;
	wire w_dff_A_cmwQA2G10_0;
	wire w_dff_A_AjzvMHCx6_0;
	wire w_dff_A_EbAumOFk7_0;
	wire w_dff_A_ysdZlWv88_0;
	wire w_dff_A_Bbez2tlE5_0;
	wire w_dff_A_6XLO7Fw82_0;
	wire w_dff_A_hKh6lD7L9_0;
	wire w_dff_A_cGkyTB5W4_0;
	wire w_dff_A_fMIrfBBI8_0;
	wire w_dff_A_JYUNmNKE9_0;
	wire w_dff_A_CvHAEX0k4_0;
	wire w_dff_A_Gv4SL5FF2_0;
	wire w_dff_A_zfun9FGi9_0;
	wire w_dff_A_9NU0YyFk1_0;
	wire w_dff_A_G2j0uwhU0_0;
	wire w_dff_A_PdFBEcAu9_0;
	wire w_dff_A_0WdiCdjO4_0;
	wire w_dff_A_HCUgIoKA0_0;
	wire w_dff_A_rfFoVhDr4_0;
	wire w_dff_A_hyB6LONs5_0;
	wire w_dff_A_ltjay0QD0_0;
	wire w_dff_A_LvphP0BZ5_0;
	wire w_dff_A_J2kPCyek1_0;
	wire w_dff_A_yTJRrLgV9_0;
	wire w_dff_A_qu3U2GnF7_0;
	wire w_dff_A_G2UL7Bd80_0;
	wire w_dff_A_wNcBxNYb8_0;
	wire w_dff_A_bDySrMfT6_0;
	wire w_dff_A_d8Rc8Dj91_0;
	wire w_dff_A_PP7L8aRr7_0;
	wire w_dff_A_RHkARyY51_0;
	wire w_dff_A_oh4qkzh30_0;
	wire w_dff_A_vb6UVT9T2_0;
	wire w_dff_A_a6ahhC4d8_0;
	wire w_dff_A_LgnjWNqr0_0;
	wire w_dff_A_b9I6DdCh8_0;
	wire w_dff_A_v8BwIdj35_0;
	wire w_dff_A_tGAEwy2j6_0;
	wire w_dff_A_NUWJri9V5_0;
	wire w_dff_A_zIXL6pBc1_0;
	wire w_dff_A_204SQmAl0_0;
	wire w_dff_A_P1U7JFDu8_0;
	wire w_dff_A_GOGGinFG4_0;
	wire w_dff_A_sWpZw6D99_0;
	wire w_dff_A_8Uk1cOcq0_2;
	wire w_dff_A_ZNdjjxTJ1_0;
	wire w_dff_A_GtvGFjjC7_0;
	wire w_dff_A_ghWEGvCc2_0;
	wire w_dff_A_FLSV3KvY3_0;
	wire w_dff_A_Bb4iMqSI9_0;
	wire w_dff_A_5BoyWzza5_0;
	wire w_dff_A_Hu7weckT3_0;
	wire w_dff_A_nPGEJE8D5_0;
	wire w_dff_A_2lmtdOzz6_0;
	wire w_dff_A_1xOC7Avq8_0;
	wire w_dff_A_i7Sdlbpb2_0;
	wire w_dff_A_HSvDHkDo9_0;
	wire w_dff_A_k7SyHhOQ6_0;
	wire w_dff_A_kJpWwXy29_0;
	wire w_dff_A_UWTEAV8C2_0;
	wire w_dff_A_6gvOMjes6_0;
	wire w_dff_A_de6d6Jpu2_0;
	wire w_dff_A_d7DrD2qF3_0;
	wire w_dff_A_VpcXFAxc1_0;
	wire w_dff_A_lzvGUfaV5_0;
	wire w_dff_A_0DNugwJW1_0;
	wire w_dff_A_LAuOrVh08_0;
	wire w_dff_A_of0dPu3C3_0;
	wire w_dff_A_tJKfD2rm2_0;
	wire w_dff_A_V36l25ax3_0;
	wire w_dff_A_anlxOSS95_0;
	wire w_dff_A_fF1kcHot1_0;
	wire w_dff_A_CzeJ0s053_0;
	wire w_dff_A_31htIorp6_0;
	wire w_dff_A_Ie903EKS2_0;
	wire w_dff_A_vyUY25xC3_0;
	wire w_dff_A_JwsDxDiU1_0;
	wire w_dff_A_xUjGRNrk5_0;
	wire w_dff_A_FjjpXrAd0_0;
	wire w_dff_A_zS849JfP3_0;
	wire w_dff_A_2A6zkH867_0;
	wire w_dff_A_m2Xk6hNZ6_0;
	wire w_dff_A_FRFGGGmw2_0;
	wire w_dff_A_t040DJOD7_0;
	wire w_dff_A_luahPP6e8_0;
	wire w_dff_A_jT8CVY1H6_0;
	wire w_dff_A_hDcxsap11_0;
	wire w_dff_A_TdIJKXMH6_0;
	wire w_dff_A_CEm9jKnO4_0;
	wire w_dff_A_2zrtAXyg6_0;
	wire w_dff_A_If2MmPWx1_0;
	wire w_dff_A_DKdcllYN9_0;
	wire w_dff_A_Ikoz8JaA7_0;
	wire w_dff_A_Qh5t4D9u8_0;
	wire w_dff_A_ICyzaWu23_0;
	wire w_dff_A_F0fqGvBY9_0;
	wire w_dff_A_rS0FBamH3_0;
	wire w_dff_A_JGJ9vYXy5_0;
	wire w_dff_A_uIBqQaBQ8_0;
	wire w_dff_A_Uqvkm0sU2_0;
	wire w_dff_A_kKTB73Rd6_0;
	wire w_dff_A_wFRSiLAG9_0;
	wire w_dff_A_DBujhYrI0_0;
	wire w_dff_A_8D78vdMV3_0;
	wire w_dff_A_5EPJFSK63_2;
	wire w_dff_A_DOExoYER6_0;
	wire w_dff_A_tFuCoYJZ8_0;
	wire w_dff_A_znDc7feD8_0;
	wire w_dff_A_hf6uyi5n3_0;
	wire w_dff_A_EhYx15uM5_0;
	wire w_dff_A_yctUxyfm9_0;
	wire w_dff_A_qAeChpos2_0;
	wire w_dff_A_7G5BdfF69_0;
	wire w_dff_A_hkBNqklD3_0;
	wire w_dff_A_Ca6reP3d4_0;
	wire w_dff_A_ujVpV9dA3_0;
	wire w_dff_A_PODTHDFB5_0;
	wire w_dff_A_maef2V9b2_0;
	wire w_dff_A_5RtaVRdA0_0;
	wire w_dff_A_GP2sS9ak0_0;
	wire w_dff_A_htKBQqzB2_0;
	wire w_dff_A_NPTNKuUW0_0;
	wire w_dff_A_bDOonGCq8_0;
	wire w_dff_A_TJbWIYZT1_0;
	wire w_dff_A_CvGGnXvv3_0;
	wire w_dff_A_cplFvibM7_0;
	wire w_dff_A_mUEyJ9456_0;
	wire w_dff_A_Ntkvz3F21_0;
	wire w_dff_A_XuGkLMtx1_0;
	wire w_dff_A_c8kEqfk06_0;
	wire w_dff_A_gtTQ0BmB3_0;
	wire w_dff_A_yud3cl7S4_0;
	wire w_dff_A_OXLZpy2o2_0;
	wire w_dff_A_XaMmCvE16_0;
	wire w_dff_A_zjPs8UHG2_0;
	wire w_dff_A_9YE8RIk48_0;
	wire w_dff_A_OucV5Ba50_0;
	wire w_dff_A_wXqAISRH6_0;
	wire w_dff_A_BE9GZZZM2_0;
	wire w_dff_A_MgWkUPIG2_0;
	wire w_dff_A_BfX6LqHl6_0;
	wire w_dff_A_XWMywfCp9_0;
	wire w_dff_A_VDjwOVe88_0;
	wire w_dff_A_z9SvHDb44_0;
	wire w_dff_A_Ivyi9z878_0;
	wire w_dff_A_XACCBGIh2_0;
	wire w_dff_A_C8moW3nw2_0;
	wire w_dff_A_OmSf8ubk7_0;
	wire w_dff_A_0kAqH5D97_0;
	wire w_dff_A_3CnDak9C2_0;
	wire w_dff_A_ER9dLIIt3_0;
	wire w_dff_A_BHu30DB33_0;
	wire w_dff_A_d3pgP1Ip1_0;
	wire w_dff_A_BWQHLhiv4_0;
	wire w_dff_A_FKtdbGcd0_0;
	wire w_dff_A_R0HwiVEl2_0;
	wire w_dff_A_lQAtHQA38_0;
	wire w_dff_A_706FWQ9x8_0;
	wire w_dff_A_lB78BTCY6_0;
	wire w_dff_A_R3LZrqqa6_0;
	wire w_dff_A_HxYS5P9r5_0;
	wire w_dff_A_zuCOQdnm3_2;
	wire w_dff_A_qOywLTmq5_0;
	wire w_dff_A_obdsjDGW8_0;
	wire w_dff_A_xlJxa8Vb2_0;
	wire w_dff_A_0bgbmw1u7_0;
	wire w_dff_A_ILkNZUoq5_0;
	wire w_dff_A_6eI363v60_0;
	wire w_dff_A_uA1SrmJJ7_0;
	wire w_dff_A_WNXOlrTT4_0;
	wire w_dff_A_YSD7njIx0_0;
	wire w_dff_A_Zqxssgrr2_0;
	wire w_dff_A_Akfrz6Km5_0;
	wire w_dff_A_fKmMWVFy6_0;
	wire w_dff_A_IweDFsLr9_0;
	wire w_dff_A_zQP5IMQI2_0;
	wire w_dff_A_2lCCdQtA1_0;
	wire w_dff_A_I5Rk9tDT0_0;
	wire w_dff_A_IRbZlG1X4_0;
	wire w_dff_A_unJmHk0G7_0;
	wire w_dff_A_1jJQ6CmA6_0;
	wire w_dff_A_xYVOu8Jh1_0;
	wire w_dff_A_WDrDF0rk5_0;
	wire w_dff_A_Edd5FS4Z2_0;
	wire w_dff_A_lZxAB5FU0_0;
	wire w_dff_A_k8jVv6X26_0;
	wire w_dff_A_8SPu4LWF3_0;
	wire w_dff_A_7K4dkvlQ1_0;
	wire w_dff_A_PrJMawVA5_0;
	wire w_dff_A_FC40UmaC4_0;
	wire w_dff_A_RmGkp7WL1_0;
	wire w_dff_A_rEhQd5jb2_0;
	wire w_dff_A_80r88e0W0_0;
	wire w_dff_A_h4QrjZNp1_0;
	wire w_dff_A_121wZNT26_0;
	wire w_dff_A_uU3aGcZC1_0;
	wire w_dff_A_aGe0Gktb9_0;
	wire w_dff_A_WzXfX8em9_0;
	wire w_dff_A_8f80AzCn1_0;
	wire w_dff_A_wmo9AFjC0_0;
	wire w_dff_A_pYmXnEHf3_0;
	wire w_dff_A_0NJjoHbh9_0;
	wire w_dff_A_3a2wgAyG2_0;
	wire w_dff_A_P8qjI5I76_0;
	wire w_dff_A_JgVGlE3Y2_0;
	wire w_dff_A_IbaDT5Bz6_0;
	wire w_dff_A_xVbIfwN30_0;
	wire w_dff_A_bw9XVCDf6_0;
	wire w_dff_A_9LKUqm8Z1_0;
	wire w_dff_A_3z8tURqP9_0;
	wire w_dff_A_l3by0rJL6_0;
	wire w_dff_A_AAdKUJSg5_0;
	wire w_dff_A_pt1GigVO4_0;
	wire w_dff_A_NS9ytCAQ5_0;
	wire w_dff_A_nT6kWBI53_0;
	wire w_dff_A_uq7HrGud8_2;
	wire w_dff_A_TMxT9gq27_0;
	wire w_dff_A_PsjvmN2d9_0;
	wire w_dff_A_vXdKlroq6_0;
	wire w_dff_A_qfwb87hp9_0;
	wire w_dff_A_L07fzR2f8_0;
	wire w_dff_A_971nGRUg1_0;
	wire w_dff_A_SxVku1ct4_0;
	wire w_dff_A_V3tVN4Im0_0;
	wire w_dff_A_73MxvM4L4_0;
	wire w_dff_A_Qr2dQSRe8_0;
	wire w_dff_A_6AuDajus5_0;
	wire w_dff_A_KBSfT7WF8_0;
	wire w_dff_A_rN9DevVI5_0;
	wire w_dff_A_rDKvsiUw2_0;
	wire w_dff_A_db6qlW7L2_0;
	wire w_dff_A_AjWnCn5s5_0;
	wire w_dff_A_v6P0995l6_0;
	wire w_dff_A_HleEHpDh9_0;
	wire w_dff_A_WVxaPR7a4_0;
	wire w_dff_A_rsIb9tsD8_0;
	wire w_dff_A_MHvAQU5z9_0;
	wire w_dff_A_9XflZ5wp0_0;
	wire w_dff_A_UEueVxvp1_0;
	wire w_dff_A_OIPmpoyZ1_0;
	wire w_dff_A_vImvgJRu9_0;
	wire w_dff_A_8h1GZ9yV9_0;
	wire w_dff_A_JHZmJGuN9_0;
	wire w_dff_A_e3anqOcU8_0;
	wire w_dff_A_NUDoO1gp9_0;
	wire w_dff_A_BdB3dXRQ4_0;
	wire w_dff_A_Y72CWuER7_0;
	wire w_dff_A_4KZaRmfv3_0;
	wire w_dff_A_vAhxgl6A1_0;
	wire w_dff_A_tgqErB8D2_0;
	wire w_dff_A_w1tZIuUt0_0;
	wire w_dff_A_bXXoCxit5_0;
	wire w_dff_A_RIUOzydE8_0;
	wire w_dff_A_uZT6NxH66_0;
	wire w_dff_A_6PVFqrjo6_0;
	wire w_dff_A_mVpMqK286_0;
	wire w_dff_A_5ooabH5y0_0;
	wire w_dff_A_LFHCtNum7_0;
	wire w_dff_A_mIL0jEPn8_0;
	wire w_dff_A_srqtGN0P2_0;
	wire w_dff_A_TAGBjDXW2_0;
	wire w_dff_A_DY96cPWi0_0;
	wire w_dff_A_vnoVe3jP8_0;
	wire w_dff_A_VVtpKOgZ7_0;
	wire w_dff_A_pw87yFbv8_0;
	wire w_dff_A_OubrqH7L0_0;
	wire w_dff_A_tHOt4IdH3_2;
	wire w_dff_A_7MZ2mz0k9_0;
	wire w_dff_A_b53s00F83_0;
	wire w_dff_A_ON4f8Xev3_0;
	wire w_dff_A_rcV7KJvx1_0;
	wire w_dff_A_jiCQ3TVQ2_0;
	wire w_dff_A_YYc3vBDR8_0;
	wire w_dff_A_jxbKZIqH0_0;
	wire w_dff_A_L1AwM1XF7_0;
	wire w_dff_A_dW5p6cFb7_0;
	wire w_dff_A_mCOWp0Dz3_0;
	wire w_dff_A_BpcZKrht8_0;
	wire w_dff_A_UVpQz22G2_0;
	wire w_dff_A_ez836HoA6_0;
	wire w_dff_A_RXF2V9y21_0;
	wire w_dff_A_esYAQnNT3_0;
	wire w_dff_A_E7bdT8Qd7_0;
	wire w_dff_A_tWqpCV4W5_0;
	wire w_dff_A_Bt6CXAh35_0;
	wire w_dff_A_KMM8obS68_0;
	wire w_dff_A_Er8mGpZx7_0;
	wire w_dff_A_GUNE9TJG3_0;
	wire w_dff_A_Hy7srK5u6_0;
	wire w_dff_A_ooQDCWvY6_0;
	wire w_dff_A_PjHqxL2c7_0;
	wire w_dff_A_Nm06FgkS6_0;
	wire w_dff_A_ukDWKzIP0_0;
	wire w_dff_A_psb2gkeg9_0;
	wire w_dff_A_oqhmc8u12_0;
	wire w_dff_A_WhpULsPz1_0;
	wire w_dff_A_FFeUrgin0_0;
	wire w_dff_A_KtR2M6lK4_0;
	wire w_dff_A_3GKXB7wb8_0;
	wire w_dff_A_OwuJQKDl3_0;
	wire w_dff_A_XSDVcXWM2_0;
	wire w_dff_A_LGv7DrxZ3_0;
	wire w_dff_A_1RQp3Hw82_0;
	wire w_dff_A_k7OETGIC4_0;
	wire w_dff_A_jmvKePer1_0;
	wire w_dff_A_CoEy92EC6_0;
	wire w_dff_A_wfgYk0t26_0;
	wire w_dff_A_v0I5MAlB2_0;
	wire w_dff_A_pud9JJYd8_0;
	wire w_dff_A_thm4pJLX7_0;
	wire w_dff_A_o77bWtWN7_0;
	wire w_dff_A_tQlpkEYN5_0;
	wire w_dff_A_DIG3mYDe4_0;
	wire w_dff_A_H5p053tj6_0;
	wire w_dff_A_c2Mb5ZJa8_2;
	wire w_dff_A_2QtLixsD2_0;
	wire w_dff_A_uuvaZpmj0_0;
	wire w_dff_A_mYaJyjgA8_0;
	wire w_dff_A_mufysFVm3_0;
	wire w_dff_A_2OdettXL0_0;
	wire w_dff_A_a7kqf7gA5_0;
	wire w_dff_A_SHPEgKHV2_0;
	wire w_dff_A_FF0HUAtC9_0;
	wire w_dff_A_AIuHiakr5_0;
	wire w_dff_A_XmEka2YI7_0;
	wire w_dff_A_NLUI8hMV8_0;
	wire w_dff_A_Bml7fNx51_0;
	wire w_dff_A_OmdLPao80_0;
	wire w_dff_A_wOHgARtJ1_0;
	wire w_dff_A_1uVmMeJY5_0;
	wire w_dff_A_MCQdHX6S4_0;
	wire w_dff_A_e6nGIGsS4_0;
	wire w_dff_A_GvN2DDQe0_0;
	wire w_dff_A_6cqk7zSv7_0;
	wire w_dff_A_IG0gKjKu3_0;
	wire w_dff_A_fVajJqO53_0;
	wire w_dff_A_VX9jnV2g5_0;
	wire w_dff_A_T05j5q9S7_0;
	wire w_dff_A_O8KAUTFA7_0;
	wire w_dff_A_30WMGuhX5_0;
	wire w_dff_A_qTIIqKoI4_0;
	wire w_dff_A_C2fTUw5T8_0;
	wire w_dff_A_ZGz6OgcM6_0;
	wire w_dff_A_Adb92XRc7_0;
	wire w_dff_A_VkDvRo3x6_0;
	wire w_dff_A_edGDrP0i1_0;
	wire w_dff_A_LyBLZUL77_0;
	wire w_dff_A_KSp9iXih7_0;
	wire w_dff_A_CqboO7gP9_0;
	wire w_dff_A_wTqkJNrg5_0;
	wire w_dff_A_SUDamReS7_0;
	wire w_dff_A_xMWb35Nh5_0;
	wire w_dff_A_FX2pFjiI5_0;
	wire w_dff_A_YgLFpDns5_0;
	wire w_dff_A_OBDpYuvZ6_0;
	wire w_dff_A_4fkCDQ9o1_0;
	wire w_dff_A_FxMM6J437_0;
	wire w_dff_A_kqZzRckG2_0;
	wire w_dff_A_VKpCHKDA0_0;
	wire w_dff_A_BoBfaVd45_2;
	wire w_dff_A_HUwlSYhX6_0;
	wire w_dff_A_oIUR6dqM9_0;
	wire w_dff_A_CzJaNVTa4_0;
	wire w_dff_A_9sacLv096_0;
	wire w_dff_A_0ZElR9Dc1_0;
	wire w_dff_A_HIkn0sTv5_0;
	wire w_dff_A_wbvpgRiS7_0;
	wire w_dff_A_xAdwfQ3B9_0;
	wire w_dff_A_deja45NH0_0;
	wire w_dff_A_BwkW8nvS9_0;
	wire w_dff_A_x2m5ql8I9_0;
	wire w_dff_A_mKLxjuKN6_0;
	wire w_dff_A_MFDQ4FUW7_0;
	wire w_dff_A_gz2DMb8F5_0;
	wire w_dff_A_JXtw0OmZ1_0;
	wire w_dff_A_nrJ9HFnl9_0;
	wire w_dff_A_1m26w6zd1_0;
	wire w_dff_A_1r3QkQAT1_0;
	wire w_dff_A_uC2UPu4F6_0;
	wire w_dff_A_oxskycKV2_0;
	wire w_dff_A_p6BT5YFx8_0;
	wire w_dff_A_6JPh4bs26_0;
	wire w_dff_A_wnTXVRLI8_0;
	wire w_dff_A_v6j4jcbP7_0;
	wire w_dff_A_jOoIs8z15_0;
	wire w_dff_A_kS8S7GOY8_0;
	wire w_dff_A_EztnLaan4_0;
	wire w_dff_A_qgEKCMsP4_0;
	wire w_dff_A_daTCcLCA0_0;
	wire w_dff_A_UTAKWyje5_0;
	wire w_dff_A_hT4eIrcv5_0;
	wire w_dff_A_wIV3bZsk2_0;
	wire w_dff_A_1Vw0DgM69_0;
	wire w_dff_A_dFckzMtr4_0;
	wire w_dff_A_5BEBlbZ29_0;
	wire w_dff_A_PN0c7vH34_0;
	wire w_dff_A_DhitR4bT0_0;
	wire w_dff_A_PbYHS0fY7_0;
	wire w_dff_A_x8gxo9aW4_0;
	wire w_dff_A_y0Hedgor8_0;
	wire w_dff_A_4FbZpWqa9_0;
	wire w_dff_A_KgRkqf0R7_2;
	wire w_dff_A_57TOYDhe0_0;
	wire w_dff_A_fQwaJS1I2_0;
	wire w_dff_A_eMsrY0Yu1_0;
	wire w_dff_A_tahyBwYu3_0;
	wire w_dff_A_VMzGH1sg5_0;
	wire w_dff_A_QaHnpNmE9_0;
	wire w_dff_A_eoRusGuQ0_0;
	wire w_dff_A_E2a54sDe0_0;
	wire w_dff_A_sQMCH4ZL4_0;
	wire w_dff_A_yCGMJXXz7_0;
	wire w_dff_A_7o0AS5ii1_0;
	wire w_dff_A_0xDEqeb50_0;
	wire w_dff_A_wwATG9FF7_0;
	wire w_dff_A_HnjsgwUJ7_0;
	wire w_dff_A_TONDlJX68_0;
	wire w_dff_A_4EGW1fdJ4_0;
	wire w_dff_A_wnSFTbd79_0;
	wire w_dff_A_gMyykVh03_0;
	wire w_dff_A_wenZNzJ06_0;
	wire w_dff_A_VzdA0mXs9_0;
	wire w_dff_A_F4832aG50_0;
	wire w_dff_A_RbuTCF7e5_0;
	wire w_dff_A_Bgt5IYUY9_0;
	wire w_dff_A_Ssko7M8N9_0;
	wire w_dff_A_lXMPsd2B7_0;
	wire w_dff_A_at9SIGRH3_0;
	wire w_dff_A_MxziXfO06_0;
	wire w_dff_A_E9eGopf17_0;
	wire w_dff_A_T8eY0KiG9_0;
	wire w_dff_A_5mKPFMY43_0;
	wire w_dff_A_bCXUs6fO8_0;
	wire w_dff_A_5gQRNCgM9_0;
	wire w_dff_A_qk7Gvbf94_0;
	wire w_dff_A_lrigsKGL7_0;
	wire w_dff_A_i8B0Knw88_0;
	wire w_dff_A_yGXwLH0h1_0;
	wire w_dff_A_liBpevxS9_0;
	wire w_dff_A_LGhsnsmq0_0;
	wire w_dff_A_WOK9KqFE4_2;
	wire w_dff_A_ndBKPnsb5_0;
	wire w_dff_A_9FPoiyZj3_0;
	wire w_dff_A_MWTCJmFJ4_0;
	wire w_dff_A_1ZDy1A874_0;
	wire w_dff_A_ZZO9IYEu9_0;
	wire w_dff_A_qduycNea2_0;
	wire w_dff_A_2spqaFr38_0;
	wire w_dff_A_ole6pWoS9_0;
	wire w_dff_A_KBiPeFWu1_0;
	wire w_dff_A_ijdeybMF7_0;
	wire w_dff_A_d622vyQJ8_0;
	wire w_dff_A_gCXp2lHf5_0;
	wire w_dff_A_j0ID7f9B8_0;
	wire w_dff_A_ueqchTOU7_0;
	wire w_dff_A_MBwDEREv2_0;
	wire w_dff_A_74Iev9hV4_0;
	wire w_dff_A_OWYvHwqG4_0;
	wire w_dff_A_v62q8RnP2_0;
	wire w_dff_A_Dw4O4psQ2_0;
	wire w_dff_A_xrq29jW81_0;
	wire w_dff_A_GCfYRd367_0;
	wire w_dff_A_5R800uff2_0;
	wire w_dff_A_iGcAk4P08_0;
	wire w_dff_A_TN8vkqXp6_0;
	wire w_dff_A_CwtW7hEU5_0;
	wire w_dff_A_zRjZBrFB2_0;
	wire w_dff_A_tnAyMi1B7_0;
	wire w_dff_A_yi6Rjdes2_0;
	wire w_dff_A_fnskD6jX3_0;
	wire w_dff_A_sgerVUJA3_0;
	wire w_dff_A_p9kkbE3G7_0;
	wire w_dff_A_Ms9amRbX0_0;
	wire w_dff_A_X6YQEXw06_0;
	wire w_dff_A_XJaLv4NV8_0;
	wire w_dff_A_lH8qR5tA7_0;
	wire w_dff_A_Mc6r1u771_2;
	wire w_dff_A_dX7JRheo4_0;
	wire w_dff_A_OUzDuztl7_0;
	wire w_dff_A_iJoGHwXF7_0;
	wire w_dff_A_x3YpxVtV3_0;
	wire w_dff_A_ee2Zi4Ac3_0;
	wire w_dff_A_xlpeibEP4_0;
	wire w_dff_A_j8VdFpOx2_0;
	wire w_dff_A_6WjwWCuz3_0;
	wire w_dff_A_GJ3arNn35_0;
	wire w_dff_A_w8sfpaRZ1_0;
	wire w_dff_A_cZz6kNqm6_0;
	wire w_dff_A_QmjvM2kS7_0;
	wire w_dff_A_7gsmhxh15_0;
	wire w_dff_A_5ENBYldk3_0;
	wire w_dff_A_q4x1fN763_0;
	wire w_dff_A_tpSB7hXw1_0;
	wire w_dff_A_sZ23K3yj8_0;
	wire w_dff_A_HA3tr5Lf5_0;
	wire w_dff_A_CFnht59b9_0;
	wire w_dff_A_afBxeI4K3_0;
	wire w_dff_A_Fu7jvWCu8_0;
	wire w_dff_A_XOdfpkN27_0;
	wire w_dff_A_q744yOYU7_0;
	wire w_dff_A_fopuVnDL1_0;
	wire w_dff_A_BUCk9ajE2_0;
	wire w_dff_A_eccZzo577_0;
	wire w_dff_A_Dpn8PgxM3_0;
	wire w_dff_A_IIoy88BV9_0;
	wire w_dff_A_fm2Dkq923_0;
	wire w_dff_A_9lpUHn895_0;
	wire w_dff_A_yESDubGW9_0;
	wire w_dff_A_moQNCgH28_0;
	wire w_dff_A_jiWzWt4L4_2;
	wire w_dff_A_dIDqiBOl1_0;
	wire w_dff_A_rSzBirvM6_0;
	wire w_dff_A_O4pnc5ZF8_0;
	wire w_dff_A_yOzwVeDO3_0;
	wire w_dff_A_BvvWRKY71_0;
	wire w_dff_A_gZca098h3_0;
	wire w_dff_A_6QztLE7t8_0;
	wire w_dff_A_i4VIAhdq7_0;
	wire w_dff_A_L3JheTda3_0;
	wire w_dff_A_xh6BYOtE9_0;
	wire w_dff_A_Djx1k5t62_0;
	wire w_dff_A_lslRqdRj0_0;
	wire w_dff_A_0fggVyqM5_0;
	wire w_dff_A_ysXlWTMC6_0;
	wire w_dff_A_jWZOckRJ8_0;
	wire w_dff_A_1429AVg40_0;
	wire w_dff_A_v59ynbEa8_0;
	wire w_dff_A_i2nvBmoI1_0;
	wire w_dff_A_CPDVvugB0_0;
	wire w_dff_A_ib6BZRE60_0;
	wire w_dff_A_99663i0F7_0;
	wire w_dff_A_wVoIObD59_0;
	wire w_dff_A_dQtWPCFS9_0;
	wire w_dff_A_Vo73PJKF6_0;
	wire w_dff_A_m75zSvps6_0;
	wire w_dff_A_iMMfIQ1a0_0;
	wire w_dff_A_iNE2THiY9_0;
	wire w_dff_A_MukCaABT9_0;
	wire w_dff_A_tBYGjeYF6_0;
	wire w_dff_A_9rj7sGa51_2;
	wire w_dff_A_2rGyWqxD3_0;
	wire w_dff_A_khaU6VDl5_0;
	wire w_dff_A_Oh9wJ5Ih3_0;
	wire w_dff_A_tjVsJESb1_0;
	wire w_dff_A_6pAtnv5w4_0;
	wire w_dff_A_5UoN3ttN7_0;
	wire w_dff_A_NuwQXmk26_0;
	wire w_dff_A_3s7FdnUw9_0;
	wire w_dff_A_i4t0viAy5_0;
	wire w_dff_A_ir5fzIHe6_0;
	wire w_dff_A_5qOx8dTl2_0;
	wire w_dff_A_rshkanSd1_0;
	wire w_dff_A_ORGcrKS00_0;
	wire w_dff_A_sfQRTK811_0;
	wire w_dff_A_X6zOP7RR0_0;
	wire w_dff_A_DOx1sjIz1_0;
	wire w_dff_A_Ibzrda5f4_0;
	wire w_dff_A_VOZsTIRo4_0;
	wire w_dff_A_RPMMjNOU7_0;
	wire w_dff_A_fQGSJnZe1_0;
	wire w_dff_A_cZDEOagL6_0;
	wire w_dff_A_2RcTKpIL0_0;
	wire w_dff_A_cxaeQwDO2_0;
	wire w_dff_A_54QgSaxP3_0;
	wire w_dff_A_nLkAw5aV9_0;
	wire w_dff_A_QGqAXeGI1_0;
	wire w_dff_A_uL2v6ct47_0;
	wire w_dff_A_BV07xd3i5_2;
	wire w_dff_A_Xje03yDQ2_0;
	wire w_dff_A_h3zk6Jrn3_0;
	wire w_dff_A_E7uRVTQs3_0;
	wire w_dff_A_78bz6EeU3_0;
	wire w_dff_A_rk42nJcK8_0;
	wire w_dff_A_AuAcb4qo2_0;
	wire w_dff_A_yCzpgHmG8_0;
	wire w_dff_A_PzbMTrsG7_0;
	wire w_dff_A_6ilraf8U8_0;
	wire w_dff_A_ERJQ2PEi7_0;
	wire w_dff_A_Xglk7kj67_0;
	wire w_dff_A_0VlsmHk84_0;
	wire w_dff_A_XQCPMD2T6_0;
	wire w_dff_A_WvWgsSb78_0;
	wire w_dff_A_tiDfvPNe3_0;
	wire w_dff_A_jAU90iYK9_0;
	wire w_dff_A_bhup45yS8_0;
	wire w_dff_A_TON4qgDI1_0;
	wire w_dff_A_ALIL2MM26_0;
	wire w_dff_A_tpE6xbK47_0;
	wire w_dff_A_lQsRyypa8_0;
	wire w_dff_A_345vOSOY1_0;
	wire w_dff_A_yrkWl3Vk0_0;
	wire w_dff_A_mmVyKzX16_0;
	wire w_dff_A_3h3AmvJd6_0;
	wire w_dff_A_9g6kPTWT1_2;
	wire w_dff_A_yYzAMPrF3_0;
	wire w_dff_A_FIQC2Vn73_0;
	wire w_dff_A_2hVNT5ue5_0;
	wire w_dff_A_IpiW9ErK0_0;
	wire w_dff_A_X7b5pT8H5_0;
	wire w_dff_A_KSLVvw7z9_0;
	wire w_dff_A_rQpk7rlt3_0;
	wire w_dff_A_PhxBhS2G7_0;
	wire w_dff_A_ywX332KF8_0;
	wire w_dff_A_cV7qit4H8_0;
	wire w_dff_A_1Gzg5Pmu1_0;
	wire w_dff_A_OrmdwKwG3_0;
	wire w_dff_A_kzCWQrg84_0;
	wire w_dff_A_jgz46Cau5_0;
	wire w_dff_A_XuK0fD9s2_0;
	wire w_dff_A_PioRJHem1_0;
	wire w_dff_A_Q8l92rz44_0;
	wire w_dff_A_zJnz07Xw2_0;
	wire w_dff_A_lmS6NKWW0_0;
	wire w_dff_A_2aZ1pcVh3_0;
	wire w_dff_A_pCuekJw62_0;
	wire w_dff_A_08N4RNqu0_0;
	wire w_dff_A_bQNov0F77_0;
	wire w_dff_A_ZwLS8Cc48_0;
	wire w_dff_A_fM5Zpmhi3_2;
	wire w_dff_A_LW1HRYzu7_0;
	wire w_dff_A_bML1SCrV3_0;
	wire w_dff_A_KkdrC1ro0_0;
	wire w_dff_A_nOBiBduh0_0;
	wire w_dff_A_tff23dYW3_0;
	wire w_dff_A_Pk9lk0Yd8_0;
	wire w_dff_A_Wxs6fsYc3_0;
	wire w_dff_A_ZEZOWqKD0_0;
	wire w_dff_A_rKRik5gr8_0;
	wire w_dff_A_C5cdIUN94_0;
	wire w_dff_A_z9CzoWJW0_0;
	wire w_dff_A_oOn6l4V28_0;
	wire w_dff_A_Xw7WBAyt0_0;
	wire w_dff_A_wgknJs2g1_0;
	wire w_dff_A_7yNV4YqP2_0;
	wire w_dff_A_fcAL6fWU0_0;
	wire w_dff_A_EDALEDbp9_0;
	wire w_dff_A_xzFzyeM54_0;
	wire w_dff_A_sQmwGAnI9_0;
	wire w_dff_A_bFpczJJL5_0;
	wire w_dff_A_mLs2v7d82_0;
	wire w_dff_A_Aa8iMiQH0_0;
	wire w_dff_A_ErYJJyU15_2;
	wire w_dff_A_oWT8ksqJ6_0;
	wire w_dff_A_2T3mfj314_0;
	wire w_dff_A_djmyjo4D4_0;
	wire w_dff_A_lVAzPl6C8_0;
	wire w_dff_A_lFx7YcLt3_0;
	wire w_dff_A_zRZgQr203_0;
	wire w_dff_A_1vdkRwWs1_0;
	wire w_dff_A_2d2Tid294_0;
	wire w_dff_A_PoSyKR9j0_0;
	wire w_dff_A_5Xz4HYIk4_0;
	wire w_dff_A_8aKbN7V35_0;
	wire w_dff_A_MdfagJWI4_0;
	wire w_dff_A_LooAqoFO0_0;
	wire w_dff_A_lmTmNccP0_0;
	wire w_dff_A_Ro6I1P4M6_0;
	wire w_dff_A_0Uy8eLJh2_0;
	wire w_dff_A_TDBduI0B3_0;
	wire w_dff_A_GbBGdva52_0;
	wire w_dff_A_sPKB2ABh1_0;
	wire w_dff_A_lkA1ZPkL1_0;
	wire w_dff_A_AzVrOdhu4_2;
	wire w_dff_A_uWjJLX7o1_0;
	wire w_dff_A_1mrElvGu7_0;
	wire w_dff_A_rCc925j66_0;
	wire w_dff_A_x6hk4h9o8_0;
	wire w_dff_A_IlsXXzrE7_0;
	wire w_dff_A_WGstDMbS8_0;
	wire w_dff_A_uKI2OQuO0_0;
	wire w_dff_A_cpKHbzom4_0;
	wire w_dff_A_A7fIhCAC5_0;
	wire w_dff_A_ivY0gT9Z9_0;
	wire w_dff_A_T7xeaIm81_0;
	wire w_dff_A_W3a0RCIO4_0;
	wire w_dff_A_odJUDopP1_0;
	wire w_dff_A_Yqy7GRQy4_0;
	wire w_dff_A_2YDdMQ9S2_0;
	wire w_dff_A_1BOzJxMq6_0;
	wire w_dff_A_1B5UmdWk3_0;
	wire w_dff_A_jAJg68wu4_0;
	wire w_dff_A_bjPY08b41_2;
	wire w_dff_A_2jBrYvVK0_0;
	wire w_dff_A_sa08IdHG5_0;
	wire w_dff_A_3TWzhnyY7_0;
	wire w_dff_A_tCf1CIk89_0;
	wire w_dff_A_2zFm7QTR3_0;
	wire w_dff_A_LkHqktZR0_0;
	wire w_dff_A_nRIk1TJg3_0;
	wire w_dff_A_ncE8H9nG1_0;
	wire w_dff_A_LVRb8WOa1_0;
	wire w_dff_A_XedGkZsb1_0;
	wire w_dff_A_ucfMcgXy8_0;
	wire w_dff_A_H3XSbEDj4_0;
	wire w_dff_A_vgVmitma8_0;
	wire w_dff_A_o7EufxxD1_0;
	wire w_dff_A_0I8W9pMw5_0;
	wire w_dff_A_19jiXv2I0_0;
	wire w_dff_A_DmqhRz3o5_2;
	wire w_dff_A_DgWwyF5U2_0;
	wire w_dff_A_SAeZcok29_0;
	wire w_dff_A_zxbBAUMZ4_0;
	wire w_dff_A_nmTVdO7T7_0;
	wire w_dff_A_FDfXMotY6_0;
	wire w_dff_A_dBCUMnWG3_0;
	wire w_dff_A_m4crRSXh5_0;
	wire w_dff_A_vJ6qf8iR8_0;
	wire w_dff_A_95jBNy331_0;
	wire w_dff_A_dcPMNw3X9_0;
	wire w_dff_A_yFIo1lZg7_0;
	wire w_dff_A_aNlcE4804_0;
	wire w_dff_A_39Q1XvvA2_0;
	wire w_dff_A_U0Pke4dh7_0;
	wire w_dff_A_Gu5QXbuJ7_2;
	wire w_dff_A_kFYN7hz33_0;
	wire w_dff_A_emrWU3Oz4_0;
	wire w_dff_A_LdM5n9v23_0;
	wire w_dff_A_x07z2FN34_0;
	wire w_dff_A_BzDGGaaP5_0;
	wire w_dff_A_WoQ0EsWS5_0;
	wire w_dff_A_9KzTNYGp0_0;
	wire w_dff_A_WiLPlZry6_0;
	wire w_dff_A_9g4tYXBj5_0;
	wire w_dff_A_aqwKUeEP2_0;
	wire w_dff_A_37BxLqwc4_0;
	wire w_dff_A_TkdbBbfy6_0;
	wire w_dff_A_TOoGb41g9_2;
	wire w_dff_A_OeQAHLUb8_0;
	wire w_dff_A_IGYDdBTf8_0;
	wire w_dff_A_qc1UiXSs2_0;
	wire w_dff_A_aGtVqjBI9_0;
	wire w_dff_A_cXTYmrrz6_0;
	wire w_dff_A_U4Fj0e5N2_0;
	wire w_dff_A_KSiVsY284_0;
	wire w_dff_A_M1cFi3QN5_0;
	wire w_dff_A_Yk6xc5Rb3_0;
	wire w_dff_A_2HGFNCac5_0;
	wire w_dff_A_CFydfasb0_2;
	wire w_dff_A_6gjinRhx1_0;
	wire w_dff_A_ItJXiioD4_0;
	wire w_dff_A_QN6EevqU0_0;
	wire w_dff_A_YXvjz82R3_0;
	wire w_dff_A_j5ZdIJbF2_0;
	wire w_dff_A_WpW4oPeJ4_0;
	wire w_dff_A_UteeaXOf7_0;
	wire w_dff_A_bL2kAIyG7_0;
	wire w_dff_A_J0Xe6gJm8_2;
	wire w_dff_A_7w5cS6BW1_0;
	wire w_dff_A_4bAsWJVA0_0;
	wire w_dff_A_gwJiPMT72_0;
	wire w_dff_A_hFKyAnbg6_0;
	wire w_dff_A_KKdOJg614_0;
	wire w_dff_A_N4F2ehqO5_0;
	wire w_dff_A_kkcMHLRb7_2;
	wire w_dff_A_tvTGKUOh1_0;
	wire w_dff_A_SVrbNEq45_0;
	wire w_dff_A_zOepyAGb0_0;
	wire w_dff_A_txUfsu520_0;
	wire w_dff_A_2YEfK94H7_2;
	wire w_dff_A_XH2YOm5t7_0;
	wire w_dff_A_TVk2CzHW5_0;
	wire w_dff_A_rdgwxBzJ1_2;
	jand g0000(.dina(w_G273gat_7[2]),.dinb(w_G1gat_7[1]),.dout(G545gat_fa_),.clk(gclk));
	jand g0001(.dina(w_G273gat_7[1]),.dinb(w_G18gat_7[2]),.dout(n65),.clk(gclk));
	jand g0002(.dina(w_G290gat_7[2]),.dinb(w_G1gat_7[0]),.dout(n66),.clk(gclk));
	jor g0003(.dina(n66),.dinb(w_n65_0[1]),.dout(n67),.clk(gclk));
	jand g0004(.dina(w_G290gat_7[1]),.dinb(w_G18gat_7[1]),.dout(n68),.clk(gclk));
	jand g0005(.dina(n68),.dinb(w_G545gat_0),.dout(n69),.clk(gclk));
	jnot g0006(.din(w_n69_0[1]),.dout(n70),.clk(gclk));
	jand g0007(.dina(w_n70_0[1]),.dinb(w_dff_B_3FRV3OSY1_1),.dout(w_dff_A_7d1LhOvD7_2),.clk(gclk));
	jand g0008(.dina(w_G307gat_7[2]),.dinb(w_G1gat_6[2]),.dout(n72),.clk(gclk));
	jnot g0009(.din(w_n72_0[1]),.dout(n73),.clk(gclk));
	jnot g0010(.din(w_G18gat_7[0]),.dout(n74),.clk(gclk));
	jnot g0011(.din(w_G290gat_7[0]),.dout(n75),.clk(gclk));
	jor g0012(.dina(w_n75_0[1]),.dinb(n74),.dout(n76),.clk(gclk));
	jnot g0013(.din(w_G35gat_7[2]),.dout(n77),.clk(gclk));
	jnot g0014(.din(w_G273gat_7[0]),.dout(n78),.clk(gclk));
	jor g0015(.dina(w_n78_0[1]),.dinb(w_n77_0[1]),.dout(n79),.clk(gclk));
	jand g0016(.dina(n79),.dinb(n76),.dout(n80),.clk(gclk));
	jand g0017(.dina(w_G290gat_6[2]),.dinb(w_G35gat_7[1]),.dout(n81),.clk(gclk));
	jand g0018(.dina(w_n81_0[1]),.dinb(w_n65_0[0]),.dout(n82),.clk(gclk));
	jor g0019(.dina(w_n82_1[1]),.dinb(n80),.dout(n83),.clk(gclk));
	jand g0020(.dina(n83),.dinb(w_n70_0[0]),.dout(n84),.clk(gclk));
	jnot g0021(.din(w_n82_1[0]),.dout(n85),.clk(gclk));
	jand g0022(.dina(w_n85_0[1]),.dinb(w_n69_0[0]),.dout(n86),.clk(gclk));
	jor g0023(.dina(w_dff_B_PSo8MNph8_0),.dinb(w_n84_0[1]),.dout(n87),.clk(gclk));
	jxor g0024(.dina(w_n87_0[1]),.dinb(w_dff_B_jMMSq32A1_1),.dout(w_dff_A_e8HaFF4D6_2),.clk(gclk));
	jand g0025(.dina(w_G324gat_7[1]),.dinb(w_G1gat_6[1]),.dout(n89),.clk(gclk));
	jnot g0026(.din(w_n89_0[1]),.dout(n90),.clk(gclk));
	jnot g0027(.din(w_n84_0[0]),.dout(n91),.clk(gclk));
	jor g0028(.dina(w_n87_0[0]),.dinb(w_n72_0[0]),.dout(n92),.clk(gclk));
	jand g0029(.dina(n92),.dinb(w_dff_B_s2BIrOrl5_1),.dout(n93),.clk(gclk));
	jand g0030(.dina(w_G307gat_7[1]),.dinb(w_G18gat_6[2]),.dout(n94),.clk(gclk));
	jnot g0031(.din(w_n94_0[1]),.dout(n95),.clk(gclk));
	jand g0032(.dina(w_G273gat_6[2]),.dinb(w_G52gat_7[2]),.dout(n96),.clk(gclk));
	jor g0033(.dina(w_n96_0[1]),.dinb(w_n81_0[0]),.dout(n97),.clk(gclk));
	jand g0034(.dina(w_G273gat_6[1]),.dinb(w_G35gat_7[0]),.dout(n98),.clk(gclk));
	jand g0035(.dina(w_G290gat_6[1]),.dinb(w_G52gat_7[1]),.dout(n99),.clk(gclk));
	jand g0036(.dina(w_n99_0[1]),.dinb(n98),.dout(n100),.clk(gclk));
	jnot g0037(.din(w_n100_1[1]),.dout(n101),.clk(gclk));
	jand g0038(.dina(w_n101_0[2]),.dinb(w_dff_B_OcM2U1nk7_1),.dout(n102),.clk(gclk));
	jor g0039(.dina(n102),.dinb(w_n82_0[2]),.dout(n103),.clk(gclk));
	jand g0040(.dina(w_n101_0[1]),.dinb(w_n82_0[1]),.dout(n104),.clk(gclk));
	jnot g0041(.din(w_n104_0[1]),.dout(n105),.clk(gclk));
	jand g0042(.dina(n105),.dinb(w_n103_0[1]),.dout(n106),.clk(gclk));
	jxor g0043(.dina(n106),.dinb(w_dff_B_Mc0qdUx74_1),.dout(n107),.clk(gclk));
	jxor g0044(.dina(w_n107_0[1]),.dinb(w_n93_0[1]),.dout(n108),.clk(gclk));
	jxor g0045(.dina(w_n108_0[1]),.dinb(w_dff_B_cSsKQ9UH7_1),.dout(w_dff_A_Q4wViHZO3_2),.clk(gclk));
	jand g0046(.dina(w_G341gat_7[1]),.dinb(w_G1gat_6[0]),.dout(n110),.clk(gclk));
	jnot g0047(.din(w_n110_0[1]),.dout(n111),.clk(gclk));
	jnot g0048(.din(w_n107_0[0]),.dout(n112),.clk(gclk));
	jor g0049(.dina(n112),.dinb(w_n93_0[0]),.dout(n113),.clk(gclk));
	jor g0050(.dina(w_n108_0[0]),.dinb(w_n89_0[0]),.dout(n114),.clk(gclk));
	jand g0051(.dina(n114),.dinb(w_dff_B_xBBblVJN9_1),.dout(n115),.clk(gclk));
	jand g0052(.dina(w_G324gat_7[0]),.dinb(w_G18gat_6[1]),.dout(n116),.clk(gclk));
	jnot g0053(.din(w_n116_0[1]),.dout(n117),.clk(gclk));
	jor g0054(.dina(w_n75_0[0]),.dinb(w_n77_0[0]),.dout(n118),.clk(gclk));
	jnot g0055(.din(w_G52gat_7[0]),.dout(n119),.clk(gclk));
	jor g0056(.dina(w_n78_0[0]),.dinb(n119),.dout(n120),.clk(gclk));
	jand g0057(.dina(n120),.dinb(n118),.dout(n121),.clk(gclk));
	jor g0058(.dina(w_n100_1[0]),.dinb(n121),.dout(n122),.clk(gclk));
	jand g0059(.dina(n122),.dinb(w_n85_0[0]),.dout(n123),.clk(gclk));
	jor g0060(.dina(w_n104_0[0]),.dinb(n123),.dout(n124),.clk(gclk));
	jor g0061(.dina(n124),.dinb(w_n94_0[0]),.dout(n125),.clk(gclk));
	jand g0062(.dina(n125),.dinb(w_n103_0[0]),.dout(n126),.clk(gclk));
	jand g0063(.dina(w_G307gat_7[0]),.dinb(w_G35gat_6[2]),.dout(n127),.clk(gclk));
	jnot g0064(.din(n127),.dout(n128),.clk(gclk));
	jand g0065(.dina(w_G273gat_6[0]),.dinb(w_G69gat_7[1]),.dout(n129),.clk(gclk));
	jor g0066(.dina(w_n129_0[1]),.dinb(w_n99_0[0]),.dout(n130),.clk(gclk));
	jand g0067(.dina(w_G290gat_6[0]),.dinb(w_G69gat_7[0]),.dout(n131),.clk(gclk));
	jand g0068(.dina(w_n131_0[1]),.dinb(w_n96_0[0]),.dout(n132),.clk(gclk));
	jnot g0069(.din(w_n132_0[2]),.dout(n133),.clk(gclk));
	jand g0070(.dina(w_n133_0[2]),.dinb(w_n130_0[1]),.dout(n134),.clk(gclk));
	jor g0071(.dina(n134),.dinb(w_n100_0[2]),.dout(n135),.clk(gclk));
	jand g0072(.dina(w_n133_0[1]),.dinb(w_n100_0[1]),.dout(n136),.clk(gclk));
	jnot g0073(.din(n136),.dout(n137),.clk(gclk));
	jand g0074(.dina(n137),.dinb(n135),.dout(n138),.clk(gclk));
	jxor g0075(.dina(w_n138_0[1]),.dinb(w_n128_0[1]),.dout(n139),.clk(gclk));
	jnot g0076(.din(w_n139_0[1]),.dout(n140),.clk(gclk));
	jxor g0077(.dina(w_n140_0[1]),.dinb(w_n126_0[2]),.dout(n141),.clk(gclk));
	jxor g0078(.dina(n141),.dinb(w_dff_B_z5yrB3Ls7_1),.dout(n142),.clk(gclk));
	jxor g0079(.dina(w_n142_0[1]),.dinb(w_n115_0[1]),.dout(n143),.clk(gclk));
	jxor g0080(.dina(w_n143_0[1]),.dinb(w_dff_B_8JplcJiB0_1),.dout(w_dff_A_b8H84EUd8_2),.clk(gclk));
	jand g0081(.dina(w_G358gat_7[1]),.dinb(w_G1gat_5[2]),.dout(n145),.clk(gclk));
	jnot g0082(.din(w_n145_0[1]),.dout(n146),.clk(gclk));
	jnot g0083(.din(w_n142_0[0]),.dout(n147),.clk(gclk));
	jor g0084(.dina(n147),.dinb(w_n115_0[0]),.dout(n148),.clk(gclk));
	jor g0085(.dina(w_n143_0[0]),.dinb(w_n110_0[0]),.dout(n149),.clk(gclk));
	jand g0086(.dina(n149),.dinb(w_dff_B_3eb8cAjZ3_1),.dout(n150),.clk(gclk));
	jand g0087(.dina(w_G341gat_7[0]),.dinb(w_G18gat_6[0]),.dout(n151),.clk(gclk));
	jnot g0088(.din(w_n151_0[1]),.dout(n152),.clk(gclk));
	jor g0089(.dina(w_n140_0[0]),.dinb(w_n126_0[1]),.dout(n153),.clk(gclk));
	jxor g0090(.dina(w_n139_0[0]),.dinb(w_n126_0[0]),.dout(n154),.clk(gclk));
	jor g0091(.dina(n154),.dinb(w_n116_0[0]),.dout(n155),.clk(gclk));
	jand g0092(.dina(n155),.dinb(w_dff_B_1ANJNn590_1),.dout(n156),.clk(gclk));
	jand g0093(.dina(w_G324gat_6[2]),.dinb(w_G35gat_6[1]),.dout(n157),.clk(gclk));
	jnot g0094(.din(n157),.dout(n158),.clk(gclk));
	jnot g0095(.din(w_n130_0[0]),.dout(n159),.clk(gclk));
	jor g0096(.dina(w_n132_0[1]),.dinb(n159),.dout(n160),.clk(gclk));
	jand g0097(.dina(n160),.dinb(w_n101_0[0]),.dout(n161),.clk(gclk));
	jand g0098(.dina(w_n138_0[0]),.dinb(w_n128_0[0]),.dout(n162),.clk(gclk));
	jor g0099(.dina(n162),.dinb(w_dff_B_xBFu5Phx7_1),.dout(n163),.clk(gclk));
	jand g0100(.dina(w_G307gat_6[2]),.dinb(w_G52gat_6[2]),.dout(n164),.clk(gclk));
	jnot g0101(.din(n164),.dout(n165),.clk(gclk));
	jand g0102(.dina(w_G273gat_5[2]),.dinb(w_G86gat_7[1]),.dout(n166),.clk(gclk));
	jor g0103(.dina(w_n166_0[1]),.dinb(w_n131_0[0]),.dout(n167),.clk(gclk));
	jand g0104(.dina(w_G290gat_5[2]),.dinb(w_G86gat_7[0]),.dout(n168),.clk(gclk));
	jand g0105(.dina(w_n168_0[1]),.dinb(w_n129_0[0]),.dout(n169),.clk(gclk));
	jnot g0106(.din(w_n169_0[2]),.dout(n170),.clk(gclk));
	jand g0107(.dina(w_n170_0[1]),.dinb(w_dff_B_KKHmuLIX0_1),.dout(n171),.clk(gclk));
	jor g0108(.dina(n171),.dinb(w_n132_0[0]),.dout(n172),.clk(gclk));
	jor g0109(.dina(w_n169_0[1]),.dinb(w_n133_0[0]),.dout(n173),.clk(gclk));
	jand g0110(.dina(w_dff_B_y5d7qXEA7_0),.dinb(w_n172_0[1]),.dout(n174),.clk(gclk));
	jxor g0111(.dina(w_n174_0[1]),.dinb(w_n165_0[1]),.dout(n175),.clk(gclk));
	jxor g0112(.dina(w_n175_0[1]),.dinb(w_n163_0[1]),.dout(n176),.clk(gclk));
	jxor g0113(.dina(w_n176_0[1]),.dinb(w_n158_0[1]),.dout(n177),.clk(gclk));
	jnot g0114(.din(w_n177_0[1]),.dout(n178),.clk(gclk));
	jxor g0115(.dina(w_n178_0[1]),.dinb(w_n156_0[2]),.dout(n179),.clk(gclk));
	jxor g0116(.dina(n179),.dinb(w_dff_B_Y8lCDkCI6_1),.dout(n180),.clk(gclk));
	jxor g0117(.dina(w_n180_0[1]),.dinb(w_n150_0[1]),.dout(n181),.clk(gclk));
	jxor g0118(.dina(w_n181_0[1]),.dinb(w_dff_B_QcEJJi5q5_1),.dout(w_dff_A_8Uk1cOcq0_2),.clk(gclk));
	jand g0119(.dina(w_G375gat_7[1]),.dinb(w_G1gat_5[1]),.dout(n183),.clk(gclk));
	jnot g0120(.din(w_n183_0[1]),.dout(n184),.clk(gclk));
	jnot g0121(.din(w_n180_0[0]),.dout(n185),.clk(gclk));
	jor g0122(.dina(n185),.dinb(w_n150_0[0]),.dout(n186),.clk(gclk));
	jor g0123(.dina(w_n181_0[0]),.dinb(w_n145_0[0]),.dout(n187),.clk(gclk));
	jand g0124(.dina(n187),.dinb(w_dff_B_pbsMynBF6_1),.dout(n188),.clk(gclk));
	jand g0125(.dina(w_G358gat_7[0]),.dinb(w_G18gat_5[2]),.dout(n189),.clk(gclk));
	jnot g0126(.din(w_n189_0[1]),.dout(n190),.clk(gclk));
	jor g0127(.dina(w_n178_0[0]),.dinb(w_n156_0[1]),.dout(n191),.clk(gclk));
	jxor g0128(.dina(w_n177_0[0]),.dinb(w_n156_0[0]),.dout(n192),.clk(gclk));
	jor g0129(.dina(n192),.dinb(w_n151_0[0]),.dout(n193),.clk(gclk));
	jand g0130(.dina(n193),.dinb(w_dff_B_eeFZZLUH4_1),.dout(n194),.clk(gclk));
	jand g0131(.dina(w_G341gat_6[2]),.dinb(w_G35gat_6[0]),.dout(n195),.clk(gclk));
	jnot g0132(.din(n195),.dout(n196),.clk(gclk));
	jand g0133(.dina(w_n175_0[0]),.dinb(w_n163_0[0]),.dout(n197),.clk(gclk));
	jand g0134(.dina(w_n176_0[0]),.dinb(w_n158_0[0]),.dout(n198),.clk(gclk));
	jor g0135(.dina(n198),.dinb(w_dff_B_5TW31LH74_1),.dout(n199),.clk(gclk));
	jand g0136(.dina(w_G324gat_6[1]),.dinb(w_G52gat_6[1]),.dout(n200),.clk(gclk));
	jnot g0137(.din(n200),.dout(n201),.clk(gclk));
	jnot g0138(.din(w_n172_0[0]),.dout(n202),.clk(gclk));
	jand g0139(.dina(w_n174_0[0]),.dinb(w_n165_0[0]),.dout(n203),.clk(gclk));
	jor g0140(.dina(n203),.dinb(w_dff_B_840c3GDk4_1),.dout(n204),.clk(gclk));
	jand g0141(.dina(w_G307gat_6[1]),.dinb(w_G69gat_6[2]),.dout(n205),.clk(gclk));
	jnot g0142(.din(n205),.dout(n206),.clk(gclk));
	jand g0143(.dina(w_G273gat_5[1]),.dinb(w_G103gat_7[1]),.dout(n207),.clk(gclk));
	jor g0144(.dina(w_n207_0[1]),.dinb(w_n168_0[0]),.dout(n208),.clk(gclk));
	jand g0145(.dina(w_G290gat_5[1]),.dinb(w_G103gat_7[0]),.dout(n209),.clk(gclk));
	jand g0146(.dina(w_n209_0[1]),.dinb(w_n166_0[0]),.dout(n210),.clk(gclk));
	jnot g0147(.din(w_n210_1[1]),.dout(n211),.clk(gclk));
	jand g0148(.dina(n211),.dinb(w_dff_B_4EFGqvCf7_1),.dout(n212),.clk(gclk));
	jor g0149(.dina(n212),.dinb(w_n169_0[0]),.dout(n213),.clk(gclk));
	jor g0150(.dina(w_n210_1[0]),.dinb(w_n170_0[0]),.dout(n214),.clk(gclk));
	jand g0151(.dina(w_dff_B_K5WYOovD9_0),.dinb(w_n213_0[1]),.dout(n215),.clk(gclk));
	jxor g0152(.dina(w_n215_0[1]),.dinb(w_n206_0[1]),.dout(n216),.clk(gclk));
	jxor g0153(.dina(w_n216_0[1]),.dinb(w_n204_0[1]),.dout(n217),.clk(gclk));
	jxor g0154(.dina(w_n217_0[1]),.dinb(w_n201_0[1]),.dout(n218),.clk(gclk));
	jxor g0155(.dina(w_n218_0[1]),.dinb(w_n199_0[1]),.dout(n219),.clk(gclk));
	jxor g0156(.dina(w_n219_0[1]),.dinb(w_n196_0[1]),.dout(n220),.clk(gclk));
	jnot g0157(.din(w_n220_0[1]),.dout(n221),.clk(gclk));
	jxor g0158(.dina(w_n221_0[1]),.dinb(w_n194_0[2]),.dout(n222),.clk(gclk));
	jxor g0159(.dina(n222),.dinb(w_dff_B_TzMqASIS7_1),.dout(n223),.clk(gclk));
	jxor g0160(.dina(w_n223_0[1]),.dinb(w_n188_0[1]),.dout(n224),.clk(gclk));
	jxor g0161(.dina(w_n224_0[1]),.dinb(w_dff_B_kiwggGnl5_1),.dout(w_dff_A_5EPJFSK63_2),.clk(gclk));
	jand g0162(.dina(w_G392gat_7[1]),.dinb(w_G1gat_5[0]),.dout(n226),.clk(gclk));
	jnot g0163(.din(w_n226_0[1]),.dout(n227),.clk(gclk));
	jnot g0164(.din(w_n223_0[0]),.dout(n228),.clk(gclk));
	jor g0165(.dina(n228),.dinb(w_n188_0[0]),.dout(n229),.clk(gclk));
	jor g0166(.dina(w_n224_0[0]),.dinb(w_n183_0[0]),.dout(n230),.clk(gclk));
	jand g0167(.dina(n230),.dinb(w_dff_B_MLjx4sMy3_1),.dout(n231),.clk(gclk));
	jand g0168(.dina(w_G375gat_7[0]),.dinb(w_G18gat_5[1]),.dout(n232),.clk(gclk));
	jnot g0169(.din(w_n232_0[1]),.dout(n233),.clk(gclk));
	jor g0170(.dina(w_n221_0[0]),.dinb(w_n194_0[1]),.dout(n234),.clk(gclk));
	jxor g0171(.dina(w_n220_0[0]),.dinb(w_n194_0[0]),.dout(n235),.clk(gclk));
	jor g0172(.dina(n235),.dinb(w_n189_0[0]),.dout(n236),.clk(gclk));
	jand g0173(.dina(n236),.dinb(w_dff_B_cbtQ91dg3_1),.dout(n237),.clk(gclk));
	jand g0174(.dina(w_G358gat_6[2]),.dinb(w_G35gat_5[2]),.dout(n238),.clk(gclk));
	jnot g0175(.din(n238),.dout(n239),.clk(gclk));
	jand g0176(.dina(w_n218_0[0]),.dinb(w_n199_0[0]),.dout(n240),.clk(gclk));
	jand g0177(.dina(w_n219_0[0]),.dinb(w_n196_0[0]),.dout(n241),.clk(gclk));
	jor g0178(.dina(n241),.dinb(w_dff_B_2fcWdJM90_1),.dout(n242),.clk(gclk));
	jand g0179(.dina(w_G341gat_6[1]),.dinb(w_G52gat_6[0]),.dout(n243),.clk(gclk));
	jnot g0180(.din(n243),.dout(n244),.clk(gclk));
	jand g0181(.dina(w_n216_0[0]),.dinb(w_n204_0[0]),.dout(n245),.clk(gclk));
	jand g0182(.dina(w_n217_0[0]),.dinb(w_n201_0[0]),.dout(n246),.clk(gclk));
	jor g0183(.dina(n246),.dinb(w_dff_B_63xYh7mI9_1),.dout(n247),.clk(gclk));
	jand g0184(.dina(w_G324gat_6[0]),.dinb(w_G69gat_6[1]),.dout(n248),.clk(gclk));
	jnot g0185(.din(n248),.dout(n249),.clk(gclk));
	jnot g0186(.din(w_n213_0[0]),.dout(n250),.clk(gclk));
	jand g0187(.dina(w_n215_0[0]),.dinb(w_n206_0[0]),.dout(n251),.clk(gclk));
	jor g0188(.dina(n251),.dinb(w_dff_B_KmYDFXAP3_1),.dout(n252),.clk(gclk));
	jand g0189(.dina(w_G307gat_6[0]),.dinb(w_G86gat_6[2]),.dout(n253),.clk(gclk));
	jnot g0190(.din(n253),.dout(n254),.clk(gclk));
	jand g0191(.dina(w_G273gat_5[0]),.dinb(w_G120gat_7[1]),.dout(n255),.clk(gclk));
	jor g0192(.dina(w_n255_0[1]),.dinb(w_n209_0[0]),.dout(n256),.clk(gclk));
	jand g0193(.dina(w_G290gat_5[0]),.dinb(w_G120gat_7[0]),.dout(n257),.clk(gclk));
	jand g0194(.dina(w_n257_0[1]),.dinb(w_n207_0[0]),.dout(n258),.clk(gclk));
	jnot g0195(.din(w_n258_0[2]),.dout(n259),.clk(gclk));
	jand g0196(.dina(w_n259_0[1]),.dinb(w_dff_B_9hPIJqTT8_1),.dout(n260),.clk(gclk));
	jor g0197(.dina(n260),.dinb(w_n210_0[2]),.dout(n261),.clk(gclk));
	jand g0198(.dina(w_n259_0[0]),.dinb(w_n210_0[1]),.dout(n262),.clk(gclk));
	jnot g0199(.din(n262),.dout(n263),.clk(gclk));
	jand g0200(.dina(n263),.dinb(w_n261_0[1]),.dout(n264),.clk(gclk));
	jxor g0201(.dina(w_n264_0[1]),.dinb(w_n254_0[1]),.dout(n265),.clk(gclk));
	jxor g0202(.dina(w_n265_0[1]),.dinb(w_n252_0[1]),.dout(n266),.clk(gclk));
	jxor g0203(.dina(w_n266_0[1]),.dinb(w_n249_0[1]),.dout(n267),.clk(gclk));
	jxor g0204(.dina(w_n267_0[1]),.dinb(w_n247_0[1]),.dout(n268),.clk(gclk));
	jxor g0205(.dina(w_n268_0[1]),.dinb(w_n244_0[1]),.dout(n269),.clk(gclk));
	jxor g0206(.dina(w_n269_0[1]),.dinb(w_n242_0[1]),.dout(n270),.clk(gclk));
	jxor g0207(.dina(w_n270_0[1]),.dinb(w_n239_0[1]),.dout(n271),.clk(gclk));
	jnot g0208(.din(w_n271_0[1]),.dout(n272),.clk(gclk));
	jxor g0209(.dina(w_n272_0[1]),.dinb(w_n237_0[2]),.dout(n273),.clk(gclk));
	jxor g0210(.dina(n273),.dinb(w_dff_B_2sGGj5117_1),.dout(n274),.clk(gclk));
	jxor g0211(.dina(w_n274_0[1]),.dinb(w_n231_0[1]),.dout(n275),.clk(gclk));
	jxor g0212(.dina(w_n275_0[1]),.dinb(w_dff_B_TAGRaUJf0_1),.dout(w_dff_A_zuCOQdnm3_2),.clk(gclk));
	jand g0213(.dina(w_G409gat_7[1]),.dinb(w_G1gat_4[2]),.dout(n277),.clk(gclk));
	jnot g0214(.din(w_n277_0[1]),.dout(n278),.clk(gclk));
	jnot g0215(.din(w_n274_0[0]),.dout(n279),.clk(gclk));
	jor g0216(.dina(n279),.dinb(w_n231_0[0]),.dout(n280),.clk(gclk));
	jor g0217(.dina(w_n275_0[0]),.dinb(w_n226_0[0]),.dout(n281),.clk(gclk));
	jand g0218(.dina(n281),.dinb(w_dff_B_EtRKUMoM0_1),.dout(n282),.clk(gclk));
	jand g0219(.dina(w_G392gat_7[0]),.dinb(w_G18gat_5[0]),.dout(n283),.clk(gclk));
	jnot g0220(.din(w_n283_0[1]),.dout(n284),.clk(gclk));
	jor g0221(.dina(w_n272_0[0]),.dinb(w_n237_0[1]),.dout(n285),.clk(gclk));
	jxor g0222(.dina(w_n271_0[0]),.dinb(w_n237_0[0]),.dout(n286),.clk(gclk));
	jor g0223(.dina(n286),.dinb(w_n232_0[0]),.dout(n287),.clk(gclk));
	jand g0224(.dina(n287),.dinb(w_dff_B_O8JHUWz01_1),.dout(n288),.clk(gclk));
	jand g0225(.dina(w_G375gat_6[2]),.dinb(w_G35gat_5[1]),.dout(n289),.clk(gclk));
	jnot g0226(.din(n289),.dout(n290),.clk(gclk));
	jand g0227(.dina(w_n269_0[0]),.dinb(w_n242_0[0]),.dout(n291),.clk(gclk));
	jand g0228(.dina(w_n270_0[0]),.dinb(w_n239_0[0]),.dout(n292),.clk(gclk));
	jor g0229(.dina(n292),.dinb(w_dff_B_al8aNhS70_1),.dout(n293),.clk(gclk));
	jand g0230(.dina(w_G358gat_6[1]),.dinb(w_G52gat_5[2]),.dout(n294),.clk(gclk));
	jnot g0231(.din(n294),.dout(n295),.clk(gclk));
	jand g0232(.dina(w_n267_0[0]),.dinb(w_n247_0[0]),.dout(n296),.clk(gclk));
	jand g0233(.dina(w_n268_0[0]),.dinb(w_n244_0[0]),.dout(n297),.clk(gclk));
	jor g0234(.dina(n297),.dinb(w_dff_B_TaolNwSg5_1),.dout(n298),.clk(gclk));
	jand g0235(.dina(w_G341gat_6[0]),.dinb(w_G69gat_6[0]),.dout(n299),.clk(gclk));
	jnot g0236(.din(n299),.dout(n300),.clk(gclk));
	jand g0237(.dina(w_n265_0[0]),.dinb(w_n252_0[0]),.dout(n301),.clk(gclk));
	jand g0238(.dina(w_n266_0[0]),.dinb(w_n249_0[0]),.dout(n302),.clk(gclk));
	jor g0239(.dina(n302),.dinb(w_dff_B_4pUskhmR3_1),.dout(n303),.clk(gclk));
	jand g0240(.dina(w_G324gat_5[2]),.dinb(w_G86gat_6[1]),.dout(n304),.clk(gclk));
	jnot g0241(.din(n304),.dout(n305),.clk(gclk));
	jnot g0242(.din(w_n261_0[0]),.dout(n306),.clk(gclk));
	jand g0243(.dina(w_n264_0[0]),.dinb(w_n254_0[0]),.dout(n307),.clk(gclk));
	jor g0244(.dina(n307),.dinb(w_dff_B_zXRprNEB1_1),.dout(n308),.clk(gclk));
	jand g0245(.dina(w_G307gat_5[2]),.dinb(w_G103gat_6[2]),.dout(n309),.clk(gclk));
	jnot g0246(.din(n309),.dout(n310),.clk(gclk));
	jand g0247(.dina(w_G273gat_4[2]),.dinb(w_G137gat_7[1]),.dout(n311),.clk(gclk));
	jor g0248(.dina(w_n311_0[1]),.dinb(w_n257_0[0]),.dout(n312),.clk(gclk));
	jand g0249(.dina(w_G290gat_4[2]),.dinb(w_G137gat_7[0]),.dout(n313),.clk(gclk));
	jand g0250(.dina(w_n313_0[1]),.dinb(w_n255_0[0]),.dout(n314),.clk(gclk));
	jnot g0251(.din(w_n314_0[2]),.dout(n315),.clk(gclk));
	jand g0252(.dina(w_n315_0[1]),.dinb(w_dff_B_oBTVm2AH7_1),.dout(n316),.clk(gclk));
	jor g0253(.dina(n316),.dinb(w_n258_0[1]),.dout(n317),.clk(gclk));
	jand g0254(.dina(w_n315_0[0]),.dinb(w_n258_0[0]),.dout(n318),.clk(gclk));
	jnot g0255(.din(n318),.dout(n319),.clk(gclk));
	jand g0256(.dina(n319),.dinb(w_n317_0[1]),.dout(n320),.clk(gclk));
	jxor g0257(.dina(w_n320_0[1]),.dinb(w_n310_0[1]),.dout(n321),.clk(gclk));
	jxor g0258(.dina(w_n321_0[1]),.dinb(w_n308_0[1]),.dout(n322),.clk(gclk));
	jxor g0259(.dina(w_n322_0[1]),.dinb(w_n305_0[1]),.dout(n323),.clk(gclk));
	jxor g0260(.dina(w_n323_0[1]),.dinb(w_n303_0[1]),.dout(n324),.clk(gclk));
	jxor g0261(.dina(w_n324_0[1]),.dinb(w_n300_0[1]),.dout(n325),.clk(gclk));
	jxor g0262(.dina(w_n325_0[1]),.dinb(w_n298_0[1]),.dout(n326),.clk(gclk));
	jxor g0263(.dina(w_n326_0[1]),.dinb(w_n295_0[1]),.dout(n327),.clk(gclk));
	jxor g0264(.dina(w_n327_0[1]),.dinb(w_n293_0[1]),.dout(n328),.clk(gclk));
	jxor g0265(.dina(w_n328_0[1]),.dinb(w_n290_0[1]),.dout(n329),.clk(gclk));
	jnot g0266(.din(w_n329_0[1]),.dout(n330),.clk(gclk));
	jxor g0267(.dina(w_n330_0[1]),.dinb(w_n288_0[2]),.dout(n331),.clk(gclk));
	jxor g0268(.dina(n331),.dinb(w_dff_B_1NeGTeA62_1),.dout(n332),.clk(gclk));
	jxor g0269(.dina(w_n332_0[1]),.dinb(w_n282_0[1]),.dout(n333),.clk(gclk));
	jxor g0270(.dina(w_n333_0[1]),.dinb(w_dff_B_NtzpAMMQ5_1),.dout(w_dff_A_uq7HrGud8_2),.clk(gclk));
	jand g0271(.dina(w_G426gat_7[1]),.dinb(w_G1gat_4[1]),.dout(n335),.clk(gclk));
	jnot g0272(.din(w_n335_0[1]),.dout(n336),.clk(gclk));
	jnot g0273(.din(w_n332_0[0]),.dout(n337),.clk(gclk));
	jor g0274(.dina(n337),.dinb(w_n282_0[0]),.dout(n338),.clk(gclk));
	jor g0275(.dina(w_n333_0[0]),.dinb(w_n277_0[0]),.dout(n339),.clk(gclk));
	jand g0276(.dina(n339),.dinb(w_dff_B_G2a9mku59_1),.dout(n340),.clk(gclk));
	jand g0277(.dina(w_G409gat_7[0]),.dinb(w_G18gat_4[2]),.dout(n341),.clk(gclk));
	jnot g0278(.din(w_n341_0[1]),.dout(n342),.clk(gclk));
	jor g0279(.dina(w_n330_0[0]),.dinb(w_n288_0[1]),.dout(n343),.clk(gclk));
	jxor g0280(.dina(w_n329_0[0]),.dinb(w_n288_0[0]),.dout(n344),.clk(gclk));
	jor g0281(.dina(n344),.dinb(w_n283_0[0]),.dout(n345),.clk(gclk));
	jand g0282(.dina(n345),.dinb(w_dff_B_fe1ABSNx2_1),.dout(n346),.clk(gclk));
	jand g0283(.dina(w_G392gat_6[2]),.dinb(w_G35gat_5[0]),.dout(n347),.clk(gclk));
	jnot g0284(.din(n347),.dout(n348),.clk(gclk));
	jand g0285(.dina(w_n327_0[0]),.dinb(w_n293_0[0]),.dout(n349),.clk(gclk));
	jand g0286(.dina(w_n328_0[0]),.dinb(w_n290_0[0]),.dout(n350),.clk(gclk));
	jor g0287(.dina(n350),.dinb(w_dff_B_jDbqou9V2_1),.dout(n351),.clk(gclk));
	jand g0288(.dina(w_G375gat_6[1]),.dinb(w_G52gat_5[1]),.dout(n352),.clk(gclk));
	jnot g0289(.din(n352),.dout(n353),.clk(gclk));
	jand g0290(.dina(w_n325_0[0]),.dinb(w_n298_0[0]),.dout(n354),.clk(gclk));
	jand g0291(.dina(w_n326_0[0]),.dinb(w_n295_0[0]),.dout(n355),.clk(gclk));
	jor g0292(.dina(n355),.dinb(w_dff_B_xT0WLZwq2_1),.dout(n356),.clk(gclk));
	jand g0293(.dina(w_G358gat_6[0]),.dinb(w_G69gat_5[2]),.dout(n357),.clk(gclk));
	jnot g0294(.din(n357),.dout(n358),.clk(gclk));
	jand g0295(.dina(w_n323_0[0]),.dinb(w_n303_0[0]),.dout(n359),.clk(gclk));
	jand g0296(.dina(w_n324_0[0]),.dinb(w_n300_0[0]),.dout(n360),.clk(gclk));
	jor g0297(.dina(n360),.dinb(w_dff_B_wBflJaNu9_1),.dout(n361),.clk(gclk));
	jand g0298(.dina(w_G341gat_5[2]),.dinb(w_G86gat_6[0]),.dout(n362),.clk(gclk));
	jnot g0299(.din(n362),.dout(n363),.clk(gclk));
	jand g0300(.dina(w_n321_0[0]),.dinb(w_n308_0[0]),.dout(n364),.clk(gclk));
	jand g0301(.dina(w_n322_0[0]),.dinb(w_n305_0[0]),.dout(n365),.clk(gclk));
	jor g0302(.dina(n365),.dinb(w_dff_B_BRvDgPUz5_1),.dout(n366),.clk(gclk));
	jand g0303(.dina(w_G324gat_5[1]),.dinb(w_G103gat_6[1]),.dout(n367),.clk(gclk));
	jnot g0304(.din(n367),.dout(n368),.clk(gclk));
	jnot g0305(.din(w_n317_0[0]),.dout(n369),.clk(gclk));
	jand g0306(.dina(w_n320_0[0]),.dinb(w_n310_0[0]),.dout(n370),.clk(gclk));
	jor g0307(.dina(n370),.dinb(w_dff_B_frfc0sZl2_1),.dout(n371),.clk(gclk));
	jand g0308(.dina(w_G307gat_5[1]),.dinb(w_G120gat_6[2]),.dout(n372),.clk(gclk));
	jand g0309(.dina(w_G273gat_4[1]),.dinb(w_G154gat_7[1]),.dout(n373),.clk(gclk));
	jor g0310(.dina(w_n373_0[1]),.dinb(w_n313_0[0]),.dout(n374),.clk(gclk));
	jand g0311(.dina(w_G290gat_4[1]),.dinb(w_G154gat_7[0]),.dout(n375),.clk(gclk));
	jand g0312(.dina(w_n375_0[1]),.dinb(w_n311_0[0]),.dout(n376),.clk(gclk));
	jnot g0313(.din(w_n376_0[2]),.dout(n377),.clk(gclk));
	jand g0314(.dina(w_n377_0[1]),.dinb(w_dff_B_wP9WFB291_1),.dout(n378),.clk(gclk));
	jor g0315(.dina(n378),.dinb(w_n314_0[1]),.dout(n379),.clk(gclk));
	jnot g0316(.din(n379),.dout(n380),.clk(gclk));
	jand g0317(.dina(w_n377_0[0]),.dinb(w_n314_0[0]),.dout(n381),.clk(gclk));
	jor g0318(.dina(w_dff_B_KMrHkR3x1_0),.dinb(w_n380_0[1]),.dout(n382),.clk(gclk));
	jxor g0319(.dina(w_n382_0[1]),.dinb(w_n372_0[1]),.dout(n383),.clk(gclk));
	jxor g0320(.dina(w_n383_0[1]),.dinb(w_n371_0[1]),.dout(n384),.clk(gclk));
	jxor g0321(.dina(w_n384_0[1]),.dinb(w_n368_0[1]),.dout(n385),.clk(gclk));
	jxor g0322(.dina(w_n385_0[1]),.dinb(w_n366_0[1]),.dout(n386),.clk(gclk));
	jxor g0323(.dina(w_n386_0[1]),.dinb(w_n363_0[1]),.dout(n387),.clk(gclk));
	jxor g0324(.dina(w_n387_0[1]),.dinb(w_n361_0[1]),.dout(n388),.clk(gclk));
	jxor g0325(.dina(w_n388_0[1]),.dinb(w_n358_0[1]),.dout(n389),.clk(gclk));
	jxor g0326(.dina(w_n389_0[1]),.dinb(w_n356_0[1]),.dout(n390),.clk(gclk));
	jxor g0327(.dina(w_n390_0[1]),.dinb(w_n353_0[1]),.dout(n391),.clk(gclk));
	jxor g0328(.dina(w_n391_0[1]),.dinb(w_n351_0[1]),.dout(n392),.clk(gclk));
	jxor g0329(.dina(w_n392_0[1]),.dinb(w_n348_0[1]),.dout(n393),.clk(gclk));
	jnot g0330(.din(w_n393_0[1]),.dout(n394),.clk(gclk));
	jxor g0331(.dina(w_n394_0[1]),.dinb(w_n346_0[2]),.dout(n395),.clk(gclk));
	jxor g0332(.dina(n395),.dinb(w_dff_B_9zhxnigc6_1),.dout(n396),.clk(gclk));
	jxor g0333(.dina(w_n396_0[1]),.dinb(w_n340_0[1]),.dout(n397),.clk(gclk));
	jxor g0334(.dina(w_n397_0[1]),.dinb(w_dff_B_7PYVdMoG0_1),.dout(w_dff_A_tHOt4IdH3_2),.clk(gclk));
	jand g0335(.dina(w_G443gat_7[1]),.dinb(w_G1gat_4[0]),.dout(n399),.clk(gclk));
	jnot g0336(.din(w_n399_0[1]),.dout(n400),.clk(gclk));
	jnot g0337(.din(w_n396_0[0]),.dout(n401),.clk(gclk));
	jor g0338(.dina(n401),.dinb(w_n340_0[0]),.dout(n402),.clk(gclk));
	jor g0339(.dina(w_n397_0[0]),.dinb(w_n335_0[0]),.dout(n403),.clk(gclk));
	jand g0340(.dina(n403),.dinb(w_dff_B_r79Ag4N17_1),.dout(n404),.clk(gclk));
	jand g0341(.dina(w_G426gat_7[0]),.dinb(w_G18gat_4[1]),.dout(n405),.clk(gclk));
	jnot g0342(.din(w_n405_0[1]),.dout(n406),.clk(gclk));
	jor g0343(.dina(w_n394_0[0]),.dinb(w_n346_0[1]),.dout(n407),.clk(gclk));
	jxor g0344(.dina(w_n393_0[0]),.dinb(w_n346_0[0]),.dout(n408),.clk(gclk));
	jor g0345(.dina(n408),.dinb(w_n341_0[0]),.dout(n409),.clk(gclk));
	jand g0346(.dina(n409),.dinb(w_dff_B_kPMvTxiM2_1),.dout(n410),.clk(gclk));
	jand g0347(.dina(w_G409gat_6[2]),.dinb(w_G35gat_4[2]),.dout(n411),.clk(gclk));
	jnot g0348(.din(n411),.dout(n412),.clk(gclk));
	jand g0349(.dina(w_n391_0[0]),.dinb(w_n351_0[0]),.dout(n413),.clk(gclk));
	jand g0350(.dina(w_n392_0[0]),.dinb(w_n348_0[0]),.dout(n414),.clk(gclk));
	jor g0351(.dina(n414),.dinb(w_dff_B_NdpLZSRB4_1),.dout(n415),.clk(gclk));
	jand g0352(.dina(w_G392gat_6[1]),.dinb(w_G52gat_5[0]),.dout(n416),.clk(gclk));
	jnot g0353(.din(n416),.dout(n417),.clk(gclk));
	jand g0354(.dina(w_n389_0[0]),.dinb(w_n356_0[0]),.dout(n418),.clk(gclk));
	jand g0355(.dina(w_n390_0[0]),.dinb(w_n353_0[0]),.dout(n419),.clk(gclk));
	jor g0356(.dina(n419),.dinb(w_dff_B_6lk4vICq9_1),.dout(n420),.clk(gclk));
	jand g0357(.dina(w_G375gat_6[0]),.dinb(w_G69gat_5[1]),.dout(n421),.clk(gclk));
	jnot g0358(.din(n421),.dout(n422),.clk(gclk));
	jand g0359(.dina(w_n387_0[0]),.dinb(w_n361_0[0]),.dout(n423),.clk(gclk));
	jand g0360(.dina(w_n388_0[0]),.dinb(w_n358_0[0]),.dout(n424),.clk(gclk));
	jor g0361(.dina(n424),.dinb(w_dff_B_VavVFlVG0_1),.dout(n425),.clk(gclk));
	jand g0362(.dina(w_G358gat_5[2]),.dinb(w_G86gat_5[2]),.dout(n426),.clk(gclk));
	jnot g0363(.din(n426),.dout(n427),.clk(gclk));
	jand g0364(.dina(w_n385_0[0]),.dinb(w_n366_0[0]),.dout(n428),.clk(gclk));
	jand g0365(.dina(w_n386_0[0]),.dinb(w_n363_0[0]),.dout(n429),.clk(gclk));
	jor g0366(.dina(n429),.dinb(w_dff_B_WEau1fSs0_1),.dout(n430),.clk(gclk));
	jand g0367(.dina(w_G341gat_5[1]),.dinb(w_G103gat_6[0]),.dout(n431),.clk(gclk));
	jnot g0368(.din(n431),.dout(n432),.clk(gclk));
	jand g0369(.dina(w_n383_0[0]),.dinb(w_n371_0[0]),.dout(n433),.clk(gclk));
	jand g0370(.dina(w_n384_0[0]),.dinb(w_n368_0[0]),.dout(n434),.clk(gclk));
	jor g0371(.dina(n434),.dinb(w_dff_B_Q5Fcfau46_1),.dout(n435),.clk(gclk));
	jand g0372(.dina(w_G324gat_5[0]),.dinb(w_G120gat_6[1]),.dout(n436),.clk(gclk));
	jnot g0373(.din(n436),.dout(n437),.clk(gclk));
	jnot g0374(.din(w_n372_0[0]),.dout(n438),.clk(gclk));
	jnot g0375(.din(w_n382_0[0]),.dout(n439),.clk(gclk));
	jand g0376(.dina(n439),.dinb(w_dff_B_aSZoaJ0K5_1),.dout(n440),.clk(gclk));
	jor g0377(.dina(n440),.dinb(w_n380_0[0]),.dout(n441),.clk(gclk));
	jand g0378(.dina(w_G307gat_5[0]),.dinb(w_G137gat_6[2]),.dout(n442),.clk(gclk));
	jand g0379(.dina(w_G273gat_4[0]),.dinb(w_G171gat_7[1]),.dout(n443),.clk(gclk));
	jor g0380(.dina(w_n443_0[1]),.dinb(w_n375_0[0]),.dout(n444),.clk(gclk));
	jand g0381(.dina(w_G290gat_4[0]),.dinb(w_G171gat_7[0]),.dout(n445),.clk(gclk));
	jand g0382(.dina(w_n445_0[1]),.dinb(w_n373_0[0]),.dout(n446),.clk(gclk));
	jnot g0383(.din(w_n446_0[2]),.dout(n447),.clk(gclk));
	jand g0384(.dina(w_n447_0[1]),.dinb(w_dff_B_B7uYD8kd4_1),.dout(n448),.clk(gclk));
	jor g0385(.dina(n448),.dinb(w_n376_0[1]),.dout(n449),.clk(gclk));
	jnot g0386(.din(n449),.dout(n450),.clk(gclk));
	jand g0387(.dina(w_n447_0[0]),.dinb(w_n376_0[0]),.dout(n451),.clk(gclk));
	jor g0388(.dina(w_dff_B_UK5oVL1A8_0),.dinb(w_n450_0[1]),.dout(n452),.clk(gclk));
	jxor g0389(.dina(w_n452_0[1]),.dinb(w_n442_0[1]),.dout(n453),.clk(gclk));
	jxor g0390(.dina(w_n453_0[1]),.dinb(w_n441_0[1]),.dout(n454),.clk(gclk));
	jxor g0391(.dina(w_n454_0[1]),.dinb(w_n437_0[1]),.dout(n455),.clk(gclk));
	jxor g0392(.dina(w_n455_0[1]),.dinb(w_n435_0[1]),.dout(n456),.clk(gclk));
	jxor g0393(.dina(w_n456_0[1]),.dinb(w_n432_0[1]),.dout(n457),.clk(gclk));
	jxor g0394(.dina(w_n457_0[1]),.dinb(w_n430_0[1]),.dout(n458),.clk(gclk));
	jxor g0395(.dina(w_n458_0[1]),.dinb(w_n427_0[1]),.dout(n459),.clk(gclk));
	jxor g0396(.dina(w_n459_0[1]),.dinb(w_n425_0[1]),.dout(n460),.clk(gclk));
	jxor g0397(.dina(w_n460_0[1]),.dinb(w_n422_0[1]),.dout(n461),.clk(gclk));
	jxor g0398(.dina(w_n461_0[1]),.dinb(w_n420_0[1]),.dout(n462),.clk(gclk));
	jxor g0399(.dina(w_n462_0[1]),.dinb(w_n417_0[1]),.dout(n463),.clk(gclk));
	jxor g0400(.dina(w_n463_0[1]),.dinb(w_n415_0[1]),.dout(n464),.clk(gclk));
	jxor g0401(.dina(w_n464_0[1]),.dinb(w_n412_0[1]),.dout(n465),.clk(gclk));
	jnot g0402(.din(w_n465_0[1]),.dout(n466),.clk(gclk));
	jxor g0403(.dina(w_n466_0[1]),.dinb(w_n410_0[2]),.dout(n467),.clk(gclk));
	jxor g0404(.dina(n467),.dinb(w_dff_B_vfMFIONK9_1),.dout(n468),.clk(gclk));
	jxor g0405(.dina(w_n468_0[1]),.dinb(w_n404_0[1]),.dout(n469),.clk(gclk));
	jxor g0406(.dina(w_n469_0[1]),.dinb(w_dff_B_N82dfrYa9_1),.dout(w_dff_A_c2Mb5ZJa8_2),.clk(gclk));
	jand g0407(.dina(w_G460gat_7[1]),.dinb(w_G1gat_3[2]),.dout(n471),.clk(gclk));
	jnot g0408(.din(w_n471_0[1]),.dout(n472),.clk(gclk));
	jnot g0409(.din(w_n468_0[0]),.dout(n473),.clk(gclk));
	jor g0410(.dina(n473),.dinb(w_n404_0[0]),.dout(n474),.clk(gclk));
	jor g0411(.dina(w_n469_0[0]),.dinb(w_n399_0[0]),.dout(n475),.clk(gclk));
	jand g0412(.dina(n475),.dinb(w_dff_B_Sas486Fy7_1),.dout(n476),.clk(gclk));
	jand g0413(.dina(w_G443gat_7[0]),.dinb(w_G18gat_4[0]),.dout(n477),.clk(gclk));
	jnot g0414(.din(w_n477_0[1]),.dout(n478),.clk(gclk));
	jor g0415(.dina(w_n466_0[0]),.dinb(w_n410_0[1]),.dout(n479),.clk(gclk));
	jxor g0416(.dina(w_n465_0[0]),.dinb(w_n410_0[0]),.dout(n480),.clk(gclk));
	jor g0417(.dina(n480),.dinb(w_n405_0[0]),.dout(n481),.clk(gclk));
	jand g0418(.dina(n481),.dinb(w_dff_B_FEoRVAiC6_1),.dout(n482),.clk(gclk));
	jand g0419(.dina(w_G426gat_6[2]),.dinb(w_G35gat_4[1]),.dout(n483),.clk(gclk));
	jnot g0420(.din(n483),.dout(n484),.clk(gclk));
	jand g0421(.dina(w_n463_0[0]),.dinb(w_n415_0[0]),.dout(n485),.clk(gclk));
	jand g0422(.dina(w_n464_0[0]),.dinb(w_n412_0[0]),.dout(n486),.clk(gclk));
	jor g0423(.dina(n486),.dinb(w_dff_B_Voqlg2Yh1_1),.dout(n487),.clk(gclk));
	jand g0424(.dina(w_G409gat_6[1]),.dinb(w_G52gat_4[2]),.dout(n488),.clk(gclk));
	jnot g0425(.din(n488),.dout(n489),.clk(gclk));
	jand g0426(.dina(w_n461_0[0]),.dinb(w_n420_0[0]),.dout(n490),.clk(gclk));
	jand g0427(.dina(w_n462_0[0]),.dinb(w_n417_0[0]),.dout(n491),.clk(gclk));
	jor g0428(.dina(n491),.dinb(w_dff_B_o0IytErQ1_1),.dout(n492),.clk(gclk));
	jand g0429(.dina(w_G392gat_6[0]),.dinb(w_G69gat_5[0]),.dout(n493),.clk(gclk));
	jnot g0430(.din(n493),.dout(n494),.clk(gclk));
	jand g0431(.dina(w_n459_0[0]),.dinb(w_n425_0[0]),.dout(n495),.clk(gclk));
	jand g0432(.dina(w_n460_0[0]),.dinb(w_n422_0[0]),.dout(n496),.clk(gclk));
	jor g0433(.dina(n496),.dinb(w_dff_B_0ub2UGTJ6_1),.dout(n497),.clk(gclk));
	jand g0434(.dina(w_G375gat_5[2]),.dinb(w_G86gat_5[1]),.dout(n498),.clk(gclk));
	jnot g0435(.din(n498),.dout(n499),.clk(gclk));
	jand g0436(.dina(w_n457_0[0]),.dinb(w_n430_0[0]),.dout(n500),.clk(gclk));
	jand g0437(.dina(w_n458_0[0]),.dinb(w_n427_0[0]),.dout(n501),.clk(gclk));
	jor g0438(.dina(n501),.dinb(w_dff_B_6mIyvaqr8_1),.dout(n502),.clk(gclk));
	jand g0439(.dina(w_G358gat_5[1]),.dinb(w_G103gat_5[2]),.dout(n503),.clk(gclk));
	jnot g0440(.din(n503),.dout(n504),.clk(gclk));
	jand g0441(.dina(w_n455_0[0]),.dinb(w_n435_0[0]),.dout(n505),.clk(gclk));
	jand g0442(.dina(w_n456_0[0]),.dinb(w_n432_0[0]),.dout(n506),.clk(gclk));
	jor g0443(.dina(n506),.dinb(w_dff_B_Vf2dWUQs7_1),.dout(n507),.clk(gclk));
	jand g0444(.dina(w_G341gat_5[0]),.dinb(w_G120gat_6[0]),.dout(n508),.clk(gclk));
	jnot g0445(.din(n508),.dout(n509),.clk(gclk));
	jand g0446(.dina(w_n453_0[0]),.dinb(w_n441_0[0]),.dout(n510),.clk(gclk));
	jand g0447(.dina(w_n454_0[0]),.dinb(w_n437_0[0]),.dout(n511),.clk(gclk));
	jor g0448(.dina(n511),.dinb(w_dff_B_NrstpOeQ0_1),.dout(n512),.clk(gclk));
	jand g0449(.dina(w_G324gat_4[2]),.dinb(w_G137gat_6[1]),.dout(n513),.clk(gclk));
	jnot g0450(.din(n513),.dout(n514),.clk(gclk));
	jnot g0451(.din(w_n442_0[0]),.dout(n515),.clk(gclk));
	jnot g0452(.din(w_n452_0[0]),.dout(n516),.clk(gclk));
	jand g0453(.dina(n516),.dinb(w_dff_B_7b9zcMbq5_1),.dout(n517),.clk(gclk));
	jor g0454(.dina(n517),.dinb(w_n450_0[0]),.dout(n518),.clk(gclk));
	jand g0455(.dina(w_G307gat_4[2]),.dinb(w_G154gat_6[2]),.dout(n519),.clk(gclk));
	jand g0456(.dina(w_G273gat_3[2]),.dinb(w_G188gat_7[1]),.dout(n520),.clk(gclk));
	jor g0457(.dina(w_n520_0[1]),.dinb(w_n445_0[0]),.dout(n521),.clk(gclk));
	jand g0458(.dina(w_G290gat_3[2]),.dinb(w_G188gat_7[0]),.dout(n522),.clk(gclk));
	jand g0459(.dina(w_n522_0[1]),.dinb(w_n443_0[0]),.dout(n523),.clk(gclk));
	jnot g0460(.din(w_n523_0[2]),.dout(n524),.clk(gclk));
	jand g0461(.dina(w_n524_0[1]),.dinb(w_dff_B_O5bHpvuc3_1),.dout(n525),.clk(gclk));
	jor g0462(.dina(n525),.dinb(w_n446_0[1]),.dout(n526),.clk(gclk));
	jnot g0463(.din(n526),.dout(n527),.clk(gclk));
	jand g0464(.dina(w_n524_0[0]),.dinb(w_n446_0[0]),.dout(n528),.clk(gclk));
	jor g0465(.dina(w_dff_B_BR1rDjUz4_0),.dinb(w_n527_0[1]),.dout(n529),.clk(gclk));
	jxor g0466(.dina(w_n529_0[1]),.dinb(w_n519_0[1]),.dout(n530),.clk(gclk));
	jxor g0467(.dina(w_n530_0[1]),.dinb(w_n518_0[1]),.dout(n531),.clk(gclk));
	jxor g0468(.dina(w_n531_0[1]),.dinb(w_n514_0[1]),.dout(n532),.clk(gclk));
	jxor g0469(.dina(w_n532_0[1]),.dinb(w_n512_0[1]),.dout(n533),.clk(gclk));
	jxor g0470(.dina(w_n533_0[1]),.dinb(w_n509_0[1]),.dout(n534),.clk(gclk));
	jxor g0471(.dina(w_n534_0[1]),.dinb(w_n507_0[1]),.dout(n535),.clk(gclk));
	jxor g0472(.dina(w_n535_0[1]),.dinb(w_n504_0[1]),.dout(n536),.clk(gclk));
	jxor g0473(.dina(w_n536_0[1]),.dinb(w_n502_0[1]),.dout(n537),.clk(gclk));
	jxor g0474(.dina(w_n537_0[1]),.dinb(w_n499_0[1]),.dout(n538),.clk(gclk));
	jxor g0475(.dina(w_n538_0[1]),.dinb(w_n497_0[1]),.dout(n539),.clk(gclk));
	jxor g0476(.dina(w_n539_0[1]),.dinb(w_n494_0[1]),.dout(n540),.clk(gclk));
	jxor g0477(.dina(w_n540_0[1]),.dinb(w_n492_0[1]),.dout(n541),.clk(gclk));
	jxor g0478(.dina(w_n541_0[1]),.dinb(w_n489_0[1]),.dout(n542),.clk(gclk));
	jxor g0479(.dina(w_n542_0[1]),.dinb(w_n487_0[1]),.dout(n543),.clk(gclk));
	jxor g0480(.dina(w_n543_0[1]),.dinb(w_n484_0[1]),.dout(n544),.clk(gclk));
	jnot g0481(.din(w_n544_0[1]),.dout(n545),.clk(gclk));
	jxor g0482(.dina(w_n545_0[1]),.dinb(w_n482_0[2]),.dout(n546),.clk(gclk));
	jxor g0483(.dina(n546),.dinb(w_dff_B_i7Y5QUbp9_1),.dout(n547),.clk(gclk));
	jxor g0484(.dina(w_n547_0[1]),.dinb(w_n476_0[1]),.dout(n548),.clk(gclk));
	jxor g0485(.dina(w_n548_0[1]),.dinb(w_dff_B_rp1raYfx8_1),.dout(w_dff_A_BoBfaVd45_2),.clk(gclk));
	jand g0486(.dina(w_G477gat_7[1]),.dinb(w_G1gat_3[1]),.dout(n550),.clk(gclk));
	jnot g0487(.din(w_n550_0[1]),.dout(n551),.clk(gclk));
	jnot g0488(.din(w_n547_0[0]),.dout(n552),.clk(gclk));
	jor g0489(.dina(n552),.dinb(w_n476_0[0]),.dout(n553),.clk(gclk));
	jor g0490(.dina(w_n548_0[0]),.dinb(w_n471_0[0]),.dout(n554),.clk(gclk));
	jand g0491(.dina(n554),.dinb(w_dff_B_XVNnUZs48_1),.dout(n555),.clk(gclk));
	jand g0492(.dina(w_G460gat_7[0]),.dinb(w_G18gat_3[2]),.dout(n556),.clk(gclk));
	jnot g0493(.din(w_n556_0[1]),.dout(n557),.clk(gclk));
	jor g0494(.dina(w_n545_0[0]),.dinb(w_n482_0[1]),.dout(n558),.clk(gclk));
	jxor g0495(.dina(w_n544_0[0]),.dinb(w_n482_0[0]),.dout(n559),.clk(gclk));
	jor g0496(.dina(n559),.dinb(w_n477_0[0]),.dout(n560),.clk(gclk));
	jand g0497(.dina(n560),.dinb(w_dff_B_wMbzty9e4_1),.dout(n561),.clk(gclk));
	jand g0498(.dina(w_G443gat_6[2]),.dinb(w_G35gat_4[0]),.dout(n562),.clk(gclk));
	jnot g0499(.din(n562),.dout(n563),.clk(gclk));
	jand g0500(.dina(w_n542_0[0]),.dinb(w_n487_0[0]),.dout(n564),.clk(gclk));
	jand g0501(.dina(w_n543_0[0]),.dinb(w_n484_0[0]),.dout(n565),.clk(gclk));
	jor g0502(.dina(n565),.dinb(w_dff_B_qm7W71SE7_1),.dout(n566),.clk(gclk));
	jand g0503(.dina(w_G426gat_6[1]),.dinb(w_G52gat_4[1]),.dout(n567),.clk(gclk));
	jnot g0504(.din(n567),.dout(n568),.clk(gclk));
	jand g0505(.dina(w_n540_0[0]),.dinb(w_n492_0[0]),.dout(n569),.clk(gclk));
	jand g0506(.dina(w_n541_0[0]),.dinb(w_n489_0[0]),.dout(n570),.clk(gclk));
	jor g0507(.dina(n570),.dinb(w_dff_B_T5RspWwv6_1),.dout(n571),.clk(gclk));
	jand g0508(.dina(w_G409gat_6[0]),.dinb(w_G69gat_4[2]),.dout(n572),.clk(gclk));
	jnot g0509(.din(n572),.dout(n573),.clk(gclk));
	jand g0510(.dina(w_n538_0[0]),.dinb(w_n497_0[0]),.dout(n574),.clk(gclk));
	jand g0511(.dina(w_n539_0[0]),.dinb(w_n494_0[0]),.dout(n575),.clk(gclk));
	jor g0512(.dina(n575),.dinb(w_dff_B_7S1vnxda9_1),.dout(n576),.clk(gclk));
	jand g0513(.dina(w_G392gat_5[2]),.dinb(w_G86gat_5[0]),.dout(n577),.clk(gclk));
	jnot g0514(.din(n577),.dout(n578),.clk(gclk));
	jand g0515(.dina(w_n536_0[0]),.dinb(w_n502_0[0]),.dout(n579),.clk(gclk));
	jand g0516(.dina(w_n537_0[0]),.dinb(w_n499_0[0]),.dout(n580),.clk(gclk));
	jor g0517(.dina(n580),.dinb(w_dff_B_mt15VX7D5_1),.dout(n581),.clk(gclk));
	jand g0518(.dina(w_G375gat_5[1]),.dinb(w_G103gat_5[1]),.dout(n582),.clk(gclk));
	jnot g0519(.din(n582),.dout(n583),.clk(gclk));
	jand g0520(.dina(w_n534_0[0]),.dinb(w_n507_0[0]),.dout(n584),.clk(gclk));
	jand g0521(.dina(w_n535_0[0]),.dinb(w_n504_0[0]),.dout(n585),.clk(gclk));
	jor g0522(.dina(n585),.dinb(w_dff_B_fglGzeOF8_1),.dout(n586),.clk(gclk));
	jand g0523(.dina(w_G358gat_5[0]),.dinb(w_G120gat_5[2]),.dout(n587),.clk(gclk));
	jnot g0524(.din(n587),.dout(n588),.clk(gclk));
	jand g0525(.dina(w_n532_0[0]),.dinb(w_n512_0[0]),.dout(n589),.clk(gclk));
	jand g0526(.dina(w_n533_0[0]),.dinb(w_n509_0[0]),.dout(n590),.clk(gclk));
	jor g0527(.dina(n590),.dinb(w_dff_B_TXZvMaLp9_1),.dout(n591),.clk(gclk));
	jand g0528(.dina(w_G341gat_4[2]),.dinb(w_G137gat_6[0]),.dout(n592),.clk(gclk));
	jnot g0529(.din(n592),.dout(n593),.clk(gclk));
	jand g0530(.dina(w_n530_0[0]),.dinb(w_n518_0[0]),.dout(n594),.clk(gclk));
	jand g0531(.dina(w_n531_0[0]),.dinb(w_n514_0[0]),.dout(n595),.clk(gclk));
	jor g0532(.dina(n595),.dinb(w_dff_B_0hhdmz5A7_1),.dout(n596),.clk(gclk));
	jand g0533(.dina(w_G324gat_4[1]),.dinb(w_G154gat_6[1]),.dout(n597),.clk(gclk));
	jnot g0534(.din(n597),.dout(n598),.clk(gclk));
	jnot g0535(.din(w_n519_0[0]),.dout(n599),.clk(gclk));
	jnot g0536(.din(w_n529_0[0]),.dout(n600),.clk(gclk));
	jand g0537(.dina(n600),.dinb(w_dff_B_bUtnm8xz7_1),.dout(n601),.clk(gclk));
	jor g0538(.dina(n601),.dinb(w_n527_0[0]),.dout(n602),.clk(gclk));
	jand g0539(.dina(w_G307gat_4[1]),.dinb(w_G171gat_6[2]),.dout(n603),.clk(gclk));
	jand g0540(.dina(w_G273gat_3[1]),.dinb(w_G205gat_7[1]),.dout(n604),.clk(gclk));
	jor g0541(.dina(w_n604_0[1]),.dinb(w_n522_0[0]),.dout(n605),.clk(gclk));
	jand g0542(.dina(w_G290gat_3[1]),.dinb(w_G205gat_7[0]),.dout(n606),.clk(gclk));
	jand g0543(.dina(w_n606_0[1]),.dinb(w_n520_0[0]),.dout(n607),.clk(gclk));
	jnot g0544(.din(w_n607_0[2]),.dout(n608),.clk(gclk));
	jand g0545(.dina(w_n608_0[1]),.dinb(w_dff_B_8Jm3I2aR8_1),.dout(n609),.clk(gclk));
	jor g0546(.dina(n609),.dinb(w_n523_0[1]),.dout(n610),.clk(gclk));
	jnot g0547(.din(n610),.dout(n611),.clk(gclk));
	jand g0548(.dina(w_n608_0[0]),.dinb(w_n523_0[0]),.dout(n612),.clk(gclk));
	jor g0549(.dina(w_dff_B_EekNaYkb0_0),.dinb(w_n611_0[1]),.dout(n613),.clk(gclk));
	jxor g0550(.dina(w_n613_0[1]),.dinb(w_n603_0[1]),.dout(n614),.clk(gclk));
	jxor g0551(.dina(w_n614_0[1]),.dinb(w_n602_0[1]),.dout(n615),.clk(gclk));
	jxor g0552(.dina(w_n615_0[1]),.dinb(w_n598_0[1]),.dout(n616),.clk(gclk));
	jxor g0553(.dina(w_n616_0[1]),.dinb(w_n596_0[1]),.dout(n617),.clk(gclk));
	jxor g0554(.dina(w_n617_0[1]),.dinb(w_n593_0[1]),.dout(n618),.clk(gclk));
	jxor g0555(.dina(w_n618_0[1]),.dinb(w_n591_0[1]),.dout(n619),.clk(gclk));
	jxor g0556(.dina(w_n619_0[1]),.dinb(w_n588_0[1]),.dout(n620),.clk(gclk));
	jxor g0557(.dina(w_n620_0[1]),.dinb(w_n586_0[1]),.dout(n621),.clk(gclk));
	jxor g0558(.dina(w_n621_0[1]),.dinb(w_n583_0[1]),.dout(n622),.clk(gclk));
	jxor g0559(.dina(w_n622_0[1]),.dinb(w_n581_0[1]),.dout(n623),.clk(gclk));
	jxor g0560(.dina(w_n623_0[1]),.dinb(w_n578_0[1]),.dout(n624),.clk(gclk));
	jxor g0561(.dina(w_n624_0[1]),.dinb(w_n576_0[1]),.dout(n625),.clk(gclk));
	jxor g0562(.dina(w_n625_0[1]),.dinb(w_n573_0[1]),.dout(n626),.clk(gclk));
	jxor g0563(.dina(w_n626_0[1]),.dinb(w_n571_0[1]),.dout(n627),.clk(gclk));
	jxor g0564(.dina(w_n627_0[1]),.dinb(w_n568_0[1]),.dout(n628),.clk(gclk));
	jxor g0565(.dina(w_n628_0[1]),.dinb(w_n566_0[1]),.dout(n629),.clk(gclk));
	jxor g0566(.dina(w_n629_0[1]),.dinb(w_n563_0[1]),.dout(n630),.clk(gclk));
	jnot g0567(.din(w_n630_0[1]),.dout(n631),.clk(gclk));
	jxor g0568(.dina(w_n631_0[1]),.dinb(w_n561_0[2]),.dout(n632),.clk(gclk));
	jxor g0569(.dina(n632),.dinb(w_dff_B_Ga7CVoxM6_1),.dout(n633),.clk(gclk));
	jxor g0570(.dina(w_n633_0[1]),.dinb(w_n555_0[1]),.dout(n634),.clk(gclk));
	jxor g0571(.dina(w_n634_0[1]),.dinb(w_dff_B_3CG9xstA3_1),.dout(w_dff_A_KgRkqf0R7_2),.clk(gclk));
	jand g0572(.dina(w_G494gat_7[1]),.dinb(w_G1gat_3[0]),.dout(n636),.clk(gclk));
	jnot g0573(.din(w_n636_0[1]),.dout(n637),.clk(gclk));
	jnot g0574(.din(w_n633_0[0]),.dout(n638),.clk(gclk));
	jor g0575(.dina(n638),.dinb(w_n555_0[0]),.dout(n639),.clk(gclk));
	jor g0576(.dina(w_n634_0[0]),.dinb(w_n550_0[0]),.dout(n640),.clk(gclk));
	jand g0577(.dina(n640),.dinb(w_dff_B_y1OoywVh9_1),.dout(n641),.clk(gclk));
	jand g0578(.dina(w_G477gat_7[0]),.dinb(w_G18gat_3[1]),.dout(n642),.clk(gclk));
	jnot g0579(.din(w_n642_0[1]),.dout(n643),.clk(gclk));
	jor g0580(.dina(w_n631_0[0]),.dinb(w_n561_0[1]),.dout(n644),.clk(gclk));
	jxor g0581(.dina(w_n630_0[0]),.dinb(w_n561_0[0]),.dout(n645),.clk(gclk));
	jor g0582(.dina(n645),.dinb(w_n556_0[0]),.dout(n646),.clk(gclk));
	jand g0583(.dina(n646),.dinb(w_dff_B_BZtiQIGW5_1),.dout(n647),.clk(gclk));
	jand g0584(.dina(w_G460gat_6[2]),.dinb(w_G35gat_3[2]),.dout(n648),.clk(gclk));
	jnot g0585(.din(n648),.dout(n649),.clk(gclk));
	jand g0586(.dina(w_n628_0[0]),.dinb(w_n566_0[0]),.dout(n650),.clk(gclk));
	jand g0587(.dina(w_n629_0[0]),.dinb(w_n563_0[0]),.dout(n651),.clk(gclk));
	jor g0588(.dina(n651),.dinb(w_dff_B_mEGkhFkZ1_1),.dout(n652),.clk(gclk));
	jand g0589(.dina(w_G443gat_6[1]),.dinb(w_G52gat_4[0]),.dout(n653),.clk(gclk));
	jnot g0590(.din(n653),.dout(n654),.clk(gclk));
	jand g0591(.dina(w_n626_0[0]),.dinb(w_n571_0[0]),.dout(n655),.clk(gclk));
	jand g0592(.dina(w_n627_0[0]),.dinb(w_n568_0[0]),.dout(n656),.clk(gclk));
	jor g0593(.dina(n656),.dinb(w_dff_B_oNQaC9jL0_1),.dout(n657),.clk(gclk));
	jand g0594(.dina(w_G426gat_6[0]),.dinb(w_G69gat_4[1]),.dout(n658),.clk(gclk));
	jnot g0595(.din(n658),.dout(n659),.clk(gclk));
	jand g0596(.dina(w_n624_0[0]),.dinb(w_n576_0[0]),.dout(n660),.clk(gclk));
	jand g0597(.dina(w_n625_0[0]),.dinb(w_n573_0[0]),.dout(n661),.clk(gclk));
	jor g0598(.dina(n661),.dinb(w_dff_B_ambeZDru3_1),.dout(n662),.clk(gclk));
	jand g0599(.dina(w_G409gat_5[2]),.dinb(w_G86gat_4[2]),.dout(n663),.clk(gclk));
	jnot g0600(.din(n663),.dout(n664),.clk(gclk));
	jand g0601(.dina(w_n622_0[0]),.dinb(w_n581_0[0]),.dout(n665),.clk(gclk));
	jand g0602(.dina(w_n623_0[0]),.dinb(w_n578_0[0]),.dout(n666),.clk(gclk));
	jor g0603(.dina(n666),.dinb(w_dff_B_URPxwRpp9_1),.dout(n667),.clk(gclk));
	jand g0604(.dina(w_G392gat_5[1]),.dinb(w_G103gat_5[0]),.dout(n668),.clk(gclk));
	jnot g0605(.din(n668),.dout(n669),.clk(gclk));
	jand g0606(.dina(w_n620_0[0]),.dinb(w_n586_0[0]),.dout(n670),.clk(gclk));
	jand g0607(.dina(w_n621_0[0]),.dinb(w_n583_0[0]),.dout(n671),.clk(gclk));
	jor g0608(.dina(n671),.dinb(w_dff_B_wUqJfUUX3_1),.dout(n672),.clk(gclk));
	jand g0609(.dina(w_G375gat_5[0]),.dinb(w_G120gat_5[1]),.dout(n673),.clk(gclk));
	jnot g0610(.din(n673),.dout(n674),.clk(gclk));
	jand g0611(.dina(w_n618_0[0]),.dinb(w_n591_0[0]),.dout(n675),.clk(gclk));
	jand g0612(.dina(w_n619_0[0]),.dinb(w_n588_0[0]),.dout(n676),.clk(gclk));
	jor g0613(.dina(n676),.dinb(w_dff_B_50KEP5WD7_1),.dout(n677),.clk(gclk));
	jand g0614(.dina(w_G358gat_4[2]),.dinb(w_G137gat_5[2]),.dout(n678),.clk(gclk));
	jnot g0615(.din(n678),.dout(n679),.clk(gclk));
	jand g0616(.dina(w_n616_0[0]),.dinb(w_n596_0[0]),.dout(n680),.clk(gclk));
	jand g0617(.dina(w_n617_0[0]),.dinb(w_n593_0[0]),.dout(n681),.clk(gclk));
	jor g0618(.dina(n681),.dinb(w_dff_B_ylrELTML5_1),.dout(n682),.clk(gclk));
	jand g0619(.dina(w_G341gat_4[1]),.dinb(w_G154gat_6[0]),.dout(n683),.clk(gclk));
	jnot g0620(.din(n683),.dout(n684),.clk(gclk));
	jand g0621(.dina(w_n614_0[0]),.dinb(w_n602_0[0]),.dout(n685),.clk(gclk));
	jand g0622(.dina(w_n615_0[0]),.dinb(w_n598_0[0]),.dout(n686),.clk(gclk));
	jor g0623(.dina(n686),.dinb(w_dff_B_Lv9VvjLv5_1),.dout(n687),.clk(gclk));
	jand g0624(.dina(w_G324gat_4[0]),.dinb(w_G171gat_6[1]),.dout(n688),.clk(gclk));
	jnot g0625(.din(n688),.dout(n689),.clk(gclk));
	jnot g0626(.din(w_n603_0[0]),.dout(n690),.clk(gclk));
	jnot g0627(.din(w_n613_0[0]),.dout(n691),.clk(gclk));
	jand g0628(.dina(n691),.dinb(w_dff_B_zSBRfi7M7_1),.dout(n692),.clk(gclk));
	jor g0629(.dina(n692),.dinb(w_n611_0[0]),.dout(n693),.clk(gclk));
	jand g0630(.dina(w_G307gat_4[0]),.dinb(w_G188gat_6[2]),.dout(n694),.clk(gclk));
	jand g0631(.dina(w_G273gat_3[0]),.dinb(w_G222gat_7[1]),.dout(n695),.clk(gclk));
	jor g0632(.dina(w_n695_0[2]),.dinb(w_n606_0[0]),.dout(n696),.clk(gclk));
	jand g0633(.dina(w_G290gat_3[0]),.dinb(w_G222gat_7[0]),.dout(n697),.clk(gclk));
	jand g0634(.dina(w_n697_0[1]),.dinb(w_n604_0[0]),.dout(n698),.clk(gclk));
	jnot g0635(.din(w_n698_0[2]),.dout(n699),.clk(gclk));
	jand g0636(.dina(w_n699_0[1]),.dinb(w_dff_B_2psNJ8Fq6_1),.dout(n700),.clk(gclk));
	jor g0637(.dina(n700),.dinb(w_n607_0[1]),.dout(n701),.clk(gclk));
	jnot g0638(.din(n701),.dout(n702),.clk(gclk));
	jand g0639(.dina(w_n699_0[0]),.dinb(w_n607_0[0]),.dout(n703),.clk(gclk));
	jor g0640(.dina(w_dff_B_wrk2j1G20_0),.dinb(w_n702_0[1]),.dout(n704),.clk(gclk));
	jxor g0641(.dina(w_n704_0[1]),.dinb(w_n694_0[1]),.dout(n705),.clk(gclk));
	jxor g0642(.dina(w_n705_0[1]),.dinb(w_n693_0[1]),.dout(n706),.clk(gclk));
	jxor g0643(.dina(w_n706_0[1]),.dinb(w_n689_0[1]),.dout(n707),.clk(gclk));
	jxor g0644(.dina(w_n707_0[1]),.dinb(w_n687_0[1]),.dout(n708),.clk(gclk));
	jxor g0645(.dina(w_n708_0[1]),.dinb(w_n684_0[1]),.dout(n709),.clk(gclk));
	jxor g0646(.dina(w_n709_0[1]),.dinb(w_n682_0[1]),.dout(n710),.clk(gclk));
	jxor g0647(.dina(w_n710_0[1]),.dinb(w_n679_0[1]),.dout(n711),.clk(gclk));
	jxor g0648(.dina(w_n711_0[1]),.dinb(w_n677_0[1]),.dout(n712),.clk(gclk));
	jxor g0649(.dina(w_n712_0[1]),.dinb(w_n674_0[1]),.dout(n713),.clk(gclk));
	jxor g0650(.dina(w_n713_0[1]),.dinb(w_n672_0[1]),.dout(n714),.clk(gclk));
	jxor g0651(.dina(w_n714_0[1]),.dinb(w_n669_0[1]),.dout(n715),.clk(gclk));
	jxor g0652(.dina(w_n715_0[1]),.dinb(w_n667_0[1]),.dout(n716),.clk(gclk));
	jxor g0653(.dina(w_n716_0[1]),.dinb(w_n664_0[1]),.dout(n717),.clk(gclk));
	jxor g0654(.dina(w_n717_0[1]),.dinb(w_n662_0[1]),.dout(n718),.clk(gclk));
	jxor g0655(.dina(w_n718_0[1]),.dinb(w_n659_0[1]),.dout(n719),.clk(gclk));
	jxor g0656(.dina(w_n719_0[1]),.dinb(w_n657_0[1]),.dout(n720),.clk(gclk));
	jxor g0657(.dina(w_n720_0[1]),.dinb(w_n654_0[1]),.dout(n721),.clk(gclk));
	jxor g0658(.dina(w_n721_0[1]),.dinb(w_n652_0[1]),.dout(n722),.clk(gclk));
	jxor g0659(.dina(w_n722_0[1]),.dinb(w_n649_0[1]),.dout(n723),.clk(gclk));
	jnot g0660(.din(w_n723_0[1]),.dout(n724),.clk(gclk));
	jxor g0661(.dina(w_n724_0[1]),.dinb(w_n647_0[2]),.dout(n725),.clk(gclk));
	jxor g0662(.dina(n725),.dinb(w_dff_B_ecnqGgPb9_1),.dout(n726),.clk(gclk));
	jxor g0663(.dina(w_n726_0[1]),.dinb(w_n641_0[1]),.dout(n727),.clk(gclk));
	jxor g0664(.dina(w_n727_0[1]),.dinb(w_dff_B_tPTGsLaV0_1),.dout(w_dff_A_WOK9KqFE4_2),.clk(gclk));
	jand g0665(.dina(w_G511gat_7[1]),.dinb(w_G1gat_2[2]),.dout(n729),.clk(gclk));
	jnot g0666(.din(w_n729_0[1]),.dout(n730),.clk(gclk));
	jnot g0667(.din(w_n726_0[0]),.dout(n731),.clk(gclk));
	jor g0668(.dina(n731),.dinb(w_n641_0[0]),.dout(n732),.clk(gclk));
	jor g0669(.dina(w_n727_0[0]),.dinb(w_n636_0[0]),.dout(n733),.clk(gclk));
	jand g0670(.dina(n733),.dinb(w_dff_B_DpzuuPns0_1),.dout(n734),.clk(gclk));
	jand g0671(.dina(w_G494gat_7[0]),.dinb(w_G18gat_3[0]),.dout(n735),.clk(gclk));
	jnot g0672(.din(w_n735_0[1]),.dout(n736),.clk(gclk));
	jor g0673(.dina(w_n724_0[0]),.dinb(w_n647_0[1]),.dout(n737),.clk(gclk));
	jxor g0674(.dina(w_n723_0[0]),.dinb(w_n647_0[0]),.dout(n738),.clk(gclk));
	jor g0675(.dina(n738),.dinb(w_n642_0[0]),.dout(n739),.clk(gclk));
	jand g0676(.dina(n739),.dinb(w_dff_B_EyD3ZNz90_1),.dout(n740),.clk(gclk));
	jand g0677(.dina(w_G477gat_6[2]),.dinb(w_G35gat_3[1]),.dout(n741),.clk(gclk));
	jnot g0678(.din(n741),.dout(n742),.clk(gclk));
	jand g0679(.dina(w_n721_0[0]),.dinb(w_n652_0[0]),.dout(n743),.clk(gclk));
	jand g0680(.dina(w_n722_0[0]),.dinb(w_n649_0[0]),.dout(n744),.clk(gclk));
	jor g0681(.dina(n744),.dinb(w_dff_B_oSL6BcdO5_1),.dout(n745),.clk(gclk));
	jand g0682(.dina(w_G460gat_6[1]),.dinb(w_G52gat_3[2]),.dout(n746),.clk(gclk));
	jnot g0683(.din(n746),.dout(n747),.clk(gclk));
	jand g0684(.dina(w_n719_0[0]),.dinb(w_n657_0[0]),.dout(n748),.clk(gclk));
	jand g0685(.dina(w_n720_0[0]),.dinb(w_n654_0[0]),.dout(n749),.clk(gclk));
	jor g0686(.dina(n749),.dinb(w_dff_B_HCj8WZ5M8_1),.dout(n750),.clk(gclk));
	jand g0687(.dina(w_G443gat_6[0]),.dinb(w_G69gat_4[0]),.dout(n751),.clk(gclk));
	jnot g0688(.din(n751),.dout(n752),.clk(gclk));
	jand g0689(.dina(w_n717_0[0]),.dinb(w_n662_0[0]),.dout(n753),.clk(gclk));
	jand g0690(.dina(w_n718_0[0]),.dinb(w_n659_0[0]),.dout(n754),.clk(gclk));
	jor g0691(.dina(n754),.dinb(w_dff_B_ScF5DwwC9_1),.dout(n755),.clk(gclk));
	jand g0692(.dina(w_G426gat_5[2]),.dinb(w_G86gat_4[1]),.dout(n756),.clk(gclk));
	jnot g0693(.din(n756),.dout(n757),.clk(gclk));
	jand g0694(.dina(w_n715_0[0]),.dinb(w_n667_0[0]),.dout(n758),.clk(gclk));
	jand g0695(.dina(w_n716_0[0]),.dinb(w_n664_0[0]),.dout(n759),.clk(gclk));
	jor g0696(.dina(n759),.dinb(w_dff_B_bcO87PmO5_1),.dout(n760),.clk(gclk));
	jand g0697(.dina(w_G409gat_5[1]),.dinb(w_G103gat_4[2]),.dout(n761),.clk(gclk));
	jnot g0698(.din(n761),.dout(n762),.clk(gclk));
	jand g0699(.dina(w_n713_0[0]),.dinb(w_n672_0[0]),.dout(n763),.clk(gclk));
	jand g0700(.dina(w_n714_0[0]),.dinb(w_n669_0[0]),.dout(n764),.clk(gclk));
	jor g0701(.dina(n764),.dinb(w_dff_B_OItvkCtj8_1),.dout(n765),.clk(gclk));
	jand g0702(.dina(w_G392gat_5[0]),.dinb(w_G120gat_5[0]),.dout(n766),.clk(gclk));
	jnot g0703(.din(n766),.dout(n767),.clk(gclk));
	jand g0704(.dina(w_n711_0[0]),.dinb(w_n677_0[0]),.dout(n768),.clk(gclk));
	jand g0705(.dina(w_n712_0[0]),.dinb(w_n674_0[0]),.dout(n769),.clk(gclk));
	jor g0706(.dina(n769),.dinb(w_dff_B_akapbC7f5_1),.dout(n770),.clk(gclk));
	jand g0707(.dina(w_G375gat_4[2]),.dinb(w_G137gat_5[1]),.dout(n771),.clk(gclk));
	jnot g0708(.din(n771),.dout(n772),.clk(gclk));
	jand g0709(.dina(w_n709_0[0]),.dinb(w_n682_0[0]),.dout(n773),.clk(gclk));
	jand g0710(.dina(w_n710_0[0]),.dinb(w_n679_0[0]),.dout(n774),.clk(gclk));
	jor g0711(.dina(n774),.dinb(w_dff_B_X2359Wtm1_1),.dout(n775),.clk(gclk));
	jand g0712(.dina(w_G358gat_4[1]),.dinb(w_G154gat_5[2]),.dout(n776),.clk(gclk));
	jnot g0713(.din(n776),.dout(n777),.clk(gclk));
	jand g0714(.dina(w_n707_0[0]),.dinb(w_n687_0[0]),.dout(n778),.clk(gclk));
	jand g0715(.dina(w_n708_0[0]),.dinb(w_n684_0[0]),.dout(n779),.clk(gclk));
	jor g0716(.dina(n779),.dinb(w_dff_B_AAYbOxiG6_1),.dout(n780),.clk(gclk));
	jand g0717(.dina(w_G341gat_4[0]),.dinb(w_G171gat_6[0]),.dout(n781),.clk(gclk));
	jnot g0718(.din(n781),.dout(n782),.clk(gclk));
	jand g0719(.dina(w_n705_0[0]),.dinb(w_n693_0[0]),.dout(n783),.clk(gclk));
	jand g0720(.dina(w_n706_0[0]),.dinb(w_n689_0[0]),.dout(n784),.clk(gclk));
	jor g0721(.dina(n784),.dinb(w_dff_B_5vWzdcRT7_1),.dout(n785),.clk(gclk));
	jand g0722(.dina(w_G324gat_3[2]),.dinb(w_G188gat_6[1]),.dout(n786),.clk(gclk));
	jnot g0723(.din(n786),.dout(n787),.clk(gclk));
	jnot g0724(.din(w_n694_0[0]),.dout(n788),.clk(gclk));
	jnot g0725(.din(w_n704_0[0]),.dout(n789),.clk(gclk));
	jand g0726(.dina(n789),.dinb(w_dff_B_Z6o9Hakd3_1),.dout(n790),.clk(gclk));
	jor g0727(.dina(n790),.dinb(w_n702_0[0]),.dout(n791),.clk(gclk));
	jand g0728(.dina(w_G307gat_3[2]),.dinb(w_G205gat_6[2]),.dout(n792),.clk(gclk));
	jand g0729(.dina(w_G273gat_2[2]),.dinb(w_G239gat_7[1]),.dout(n793),.clk(gclk));
	jor g0730(.dina(w_n793_0[1]),.dinb(w_n697_0[0]),.dout(n794),.clk(gclk));
	jand g0731(.dina(w_G290gat_2[2]),.dinb(w_G239gat_7[0]),.dout(n795),.clk(gclk));
	jand g0732(.dina(w_n795_0[1]),.dinb(w_n695_0[1]),.dout(n796),.clk(gclk));
	jnot g0733(.din(n796),.dout(n797),.clk(gclk));
	jand g0734(.dina(w_n797_0[2]),.dinb(w_dff_B_mzYTa5E69_1),.dout(n798),.clk(gclk));
	jor g0735(.dina(n798),.dinb(w_n698_0[1]),.dout(n799),.clk(gclk));
	jnot g0736(.din(n799),.dout(n800),.clk(gclk));
	jand g0737(.dina(w_n797_0[1]),.dinb(w_n698_0[0]),.dout(n801),.clk(gclk));
	jor g0738(.dina(w_dff_B_zSHMYozx7_0),.dinb(w_n800_0[1]),.dout(n802),.clk(gclk));
	jxor g0739(.dina(w_n802_0[1]),.dinb(w_n792_0[1]),.dout(n803),.clk(gclk));
	jxor g0740(.dina(w_n803_0[1]),.dinb(w_n791_0[1]),.dout(n804),.clk(gclk));
	jxor g0741(.dina(w_n804_0[1]),.dinb(w_n787_0[1]),.dout(n805),.clk(gclk));
	jxor g0742(.dina(w_n805_0[1]),.dinb(w_n785_0[1]),.dout(n806),.clk(gclk));
	jxor g0743(.dina(w_n806_0[1]),.dinb(w_n782_0[1]),.dout(n807),.clk(gclk));
	jxor g0744(.dina(w_n807_0[1]),.dinb(w_n780_0[1]),.dout(n808),.clk(gclk));
	jxor g0745(.dina(w_n808_0[1]),.dinb(w_n777_0[1]),.dout(n809),.clk(gclk));
	jxor g0746(.dina(w_n809_0[1]),.dinb(w_n775_0[1]),.dout(n810),.clk(gclk));
	jxor g0747(.dina(w_n810_0[1]),.dinb(w_n772_0[1]),.dout(n811),.clk(gclk));
	jxor g0748(.dina(w_n811_0[1]),.dinb(w_n770_0[1]),.dout(n812),.clk(gclk));
	jxor g0749(.dina(w_n812_0[1]),.dinb(w_n767_0[1]),.dout(n813),.clk(gclk));
	jxor g0750(.dina(w_n813_0[1]),.dinb(w_n765_0[1]),.dout(n814),.clk(gclk));
	jxor g0751(.dina(w_n814_0[1]),.dinb(w_n762_0[1]),.dout(n815),.clk(gclk));
	jxor g0752(.dina(w_n815_0[1]),.dinb(w_n760_0[1]),.dout(n816),.clk(gclk));
	jxor g0753(.dina(w_n816_0[1]),.dinb(w_n757_0[1]),.dout(n817),.clk(gclk));
	jxor g0754(.dina(w_n817_0[1]),.dinb(w_n755_0[1]),.dout(n818),.clk(gclk));
	jxor g0755(.dina(w_n818_0[1]),.dinb(w_n752_0[1]),.dout(n819),.clk(gclk));
	jxor g0756(.dina(w_n819_0[1]),.dinb(w_n750_0[1]),.dout(n820),.clk(gclk));
	jxor g0757(.dina(w_n820_0[1]),.dinb(w_n747_0[1]),.dout(n821),.clk(gclk));
	jxor g0758(.dina(w_n821_0[1]),.dinb(w_n745_0[1]),.dout(n822),.clk(gclk));
	jxor g0759(.dina(w_n822_0[1]),.dinb(w_n742_0[1]),.dout(n823),.clk(gclk));
	jnot g0760(.din(w_n823_0[1]),.dout(n824),.clk(gclk));
	jxor g0761(.dina(w_n824_0[1]),.dinb(w_n740_0[2]),.dout(n825),.clk(gclk));
	jxor g0762(.dina(n825),.dinb(w_dff_B_xjv428pr0_1),.dout(n826),.clk(gclk));
	jxor g0763(.dina(w_n826_0[1]),.dinb(w_n734_0[1]),.dout(n827),.clk(gclk));
	jxor g0764(.dina(w_n827_0[1]),.dinb(w_dff_B_xMYa2SRa8_1),.dout(w_dff_A_Mc6r1u771_2),.clk(gclk));
	jand g0765(.dina(w_G528gat_7[1]),.dinb(w_G1gat_2[1]),.dout(n829),.clk(gclk));
	jnot g0766(.din(w_n829_0[1]),.dout(n830),.clk(gclk));
	jnot g0767(.din(w_n826_0[0]),.dout(n831),.clk(gclk));
	jor g0768(.dina(n831),.dinb(w_n734_0[0]),.dout(n832),.clk(gclk));
	jor g0769(.dina(w_n827_0[0]),.dinb(w_n729_0[0]),.dout(n833),.clk(gclk));
	jand g0770(.dina(n833),.dinb(w_dff_B_WgXmBxuA8_1),.dout(n834),.clk(gclk));
	jand g0771(.dina(w_G511gat_7[0]),.dinb(w_G18gat_2[2]),.dout(n835),.clk(gclk));
	jor g0772(.dina(w_n824_0[0]),.dinb(w_n740_0[1]),.dout(n836),.clk(gclk));
	jxor g0773(.dina(w_n823_0[0]),.dinb(w_n740_0[0]),.dout(n837),.clk(gclk));
	jor g0774(.dina(n837),.dinb(w_n735_0[0]),.dout(n838),.clk(gclk));
	jand g0775(.dina(n838),.dinb(w_dff_B_ovdRJMmp2_1),.dout(n839),.clk(gclk));
	jand g0776(.dina(w_G494gat_6[2]),.dinb(w_G35gat_3[0]),.dout(n840),.clk(gclk));
	jnot g0777(.din(w_n840_0[1]),.dout(n841),.clk(gclk));
	jand g0778(.dina(w_n821_0[0]),.dinb(w_n745_0[0]),.dout(n842),.clk(gclk));
	jand g0779(.dina(w_n822_0[0]),.dinb(w_n742_0[0]),.dout(n843),.clk(gclk));
	jor g0780(.dina(n843),.dinb(w_dff_B_fW2vjjGI2_1),.dout(n844),.clk(gclk));
	jand g0781(.dina(w_G477gat_6[1]),.dinb(w_G52gat_3[1]),.dout(n845),.clk(gclk));
	jnot g0782(.din(n845),.dout(n846),.clk(gclk));
	jand g0783(.dina(w_n819_0[0]),.dinb(w_n750_0[0]),.dout(n847),.clk(gclk));
	jand g0784(.dina(w_n820_0[0]),.dinb(w_n747_0[0]),.dout(n848),.clk(gclk));
	jor g0785(.dina(n848),.dinb(w_dff_B_zMMYx8m05_1),.dout(n849),.clk(gclk));
	jand g0786(.dina(w_G460gat_6[0]),.dinb(w_G69gat_3[2]),.dout(n850),.clk(gclk));
	jnot g0787(.din(n850),.dout(n851),.clk(gclk));
	jand g0788(.dina(w_n817_0[0]),.dinb(w_n755_0[0]),.dout(n852),.clk(gclk));
	jand g0789(.dina(w_n818_0[0]),.dinb(w_n752_0[0]),.dout(n853),.clk(gclk));
	jor g0790(.dina(n853),.dinb(w_dff_B_ts1N6ri07_1),.dout(n854),.clk(gclk));
	jand g0791(.dina(w_G443gat_5[2]),.dinb(w_G86gat_4[0]),.dout(n855),.clk(gclk));
	jnot g0792(.din(n855),.dout(n856),.clk(gclk));
	jand g0793(.dina(w_n815_0[0]),.dinb(w_n760_0[0]),.dout(n857),.clk(gclk));
	jand g0794(.dina(w_n816_0[0]),.dinb(w_n757_0[0]),.dout(n858),.clk(gclk));
	jor g0795(.dina(n858),.dinb(w_dff_B_ejihLi905_1),.dout(n859),.clk(gclk));
	jand g0796(.dina(w_G426gat_5[1]),.dinb(w_G103gat_4[1]),.dout(n860),.clk(gclk));
	jnot g0797(.din(n860),.dout(n861),.clk(gclk));
	jand g0798(.dina(w_n813_0[0]),.dinb(w_n765_0[0]),.dout(n862),.clk(gclk));
	jand g0799(.dina(w_n814_0[0]),.dinb(w_n762_0[0]),.dout(n863),.clk(gclk));
	jor g0800(.dina(n863),.dinb(w_dff_B_BjPK4aKx5_1),.dout(n864),.clk(gclk));
	jand g0801(.dina(w_G409gat_5[0]),.dinb(w_G120gat_4[2]),.dout(n865),.clk(gclk));
	jnot g0802(.din(n865),.dout(n866),.clk(gclk));
	jand g0803(.dina(w_n811_0[0]),.dinb(w_n770_0[0]),.dout(n867),.clk(gclk));
	jand g0804(.dina(w_n812_0[0]),.dinb(w_n767_0[0]),.dout(n868),.clk(gclk));
	jor g0805(.dina(n868),.dinb(w_dff_B_PslMiuzK5_1),.dout(n869),.clk(gclk));
	jand g0806(.dina(w_G392gat_4[2]),.dinb(w_G137gat_5[0]),.dout(n870),.clk(gclk));
	jnot g0807(.din(n870),.dout(n871),.clk(gclk));
	jand g0808(.dina(w_n809_0[0]),.dinb(w_n775_0[0]),.dout(n872),.clk(gclk));
	jand g0809(.dina(w_n810_0[0]),.dinb(w_n772_0[0]),.dout(n873),.clk(gclk));
	jor g0810(.dina(n873),.dinb(w_dff_B_jyFNJZ921_1),.dout(n874),.clk(gclk));
	jand g0811(.dina(w_G375gat_4[1]),.dinb(w_G154gat_5[1]),.dout(n875),.clk(gclk));
	jnot g0812(.din(n875),.dout(n876),.clk(gclk));
	jand g0813(.dina(w_n807_0[0]),.dinb(w_n780_0[0]),.dout(n877),.clk(gclk));
	jand g0814(.dina(w_n808_0[0]),.dinb(w_n777_0[0]),.dout(n878),.clk(gclk));
	jor g0815(.dina(n878),.dinb(w_dff_B_I2zCEZrO8_1),.dout(n879),.clk(gclk));
	jand g0816(.dina(w_G358gat_4[0]),.dinb(w_G171gat_5[2]),.dout(n880),.clk(gclk));
	jnot g0817(.din(n880),.dout(n881),.clk(gclk));
	jand g0818(.dina(w_n805_0[0]),.dinb(w_n785_0[0]),.dout(n882),.clk(gclk));
	jand g0819(.dina(w_n806_0[0]),.dinb(w_n782_0[0]),.dout(n883),.clk(gclk));
	jor g0820(.dina(n883),.dinb(w_dff_B_mzUSu3Sl6_1),.dout(n884),.clk(gclk));
	jand g0821(.dina(w_G341gat_3[2]),.dinb(w_G188gat_6[0]),.dout(n885),.clk(gclk));
	jnot g0822(.din(n885),.dout(n886),.clk(gclk));
	jand g0823(.dina(w_n803_0[0]),.dinb(w_n791_0[0]),.dout(n887),.clk(gclk));
	jand g0824(.dina(w_n804_0[0]),.dinb(w_n787_0[0]),.dout(n888),.clk(gclk));
	jor g0825(.dina(n888),.dinb(w_dff_B_Th5MwW257_1),.dout(n889),.clk(gclk));
	jand g0826(.dina(w_G324gat_3[1]),.dinb(w_G205gat_6[1]),.dout(n890),.clk(gclk));
	jnot g0827(.din(n890),.dout(n891),.clk(gclk));
	jnot g0828(.din(w_n792_0[0]),.dout(n892),.clk(gclk));
	jnot g0829(.din(w_n802_0[0]),.dout(n893),.clk(gclk));
	jand g0830(.dina(n893),.dinb(w_dff_B_t0DlR4tB3_1),.dout(n894),.clk(gclk));
	jor g0831(.dina(n894),.dinb(w_n800_0[0]),.dout(n895),.clk(gclk));
	jand g0832(.dina(w_G307gat_3[1]),.dinb(w_G222gat_6[2]),.dout(n896),.clk(gclk));
	jnot g0833(.din(w_n795_0[0]),.dout(n897),.clk(gclk));
	jand g0834(.dina(w_G273gat_2[1]),.dinb(w_G256gat_7[1]),.dout(n898),.clk(gclk));
	jand g0835(.dina(w_n898_0[1]),.dinb(w_n897_0[1]),.dout(n899),.clk(gclk));
	jnot g0836(.din(n899),.dout(n900),.clk(gclk));
	jor g0837(.dina(w_n898_0[0]),.dinb(w_n897_0[0]),.dout(n901),.clk(gclk));
	jand g0838(.dina(w_n901_0[1]),.dinb(w_n797_0[0]),.dout(n902),.clk(gclk));
	jand g0839(.dina(n902),.dinb(n900),.dout(n903),.clk(gclk));
	jnot g0840(.din(w_n901_0[0]),.dout(n904),.clk(gclk));
	jand g0841(.dina(n904),.dinb(w_n695_0[0]),.dout(n905),.clk(gclk));
	jor g0842(.dina(n905),.dinb(w_n903_0[1]),.dout(n906),.clk(gclk));
	jxor g0843(.dina(w_n906_0[1]),.dinb(w_n896_0[1]),.dout(n907),.clk(gclk));
	jxor g0844(.dina(w_n907_0[1]),.dinb(w_n895_0[1]),.dout(n908),.clk(gclk));
	jxor g0845(.dina(w_n908_0[1]),.dinb(w_n891_0[1]),.dout(n909),.clk(gclk));
	jxor g0846(.dina(w_n909_0[1]),.dinb(w_n889_0[1]),.dout(n910),.clk(gclk));
	jxor g0847(.dina(w_n910_0[1]),.dinb(w_n886_0[1]),.dout(n911),.clk(gclk));
	jxor g0848(.dina(w_n911_0[1]),.dinb(w_n884_0[1]),.dout(n912),.clk(gclk));
	jxor g0849(.dina(w_n912_0[1]),.dinb(w_n881_0[1]),.dout(n913),.clk(gclk));
	jxor g0850(.dina(w_n913_0[1]),.dinb(w_n879_0[1]),.dout(n914),.clk(gclk));
	jxor g0851(.dina(w_n914_0[1]),.dinb(w_n876_0[1]),.dout(n915),.clk(gclk));
	jxor g0852(.dina(w_n915_0[1]),.dinb(w_n874_0[1]),.dout(n916),.clk(gclk));
	jxor g0853(.dina(w_n916_0[1]),.dinb(w_n871_0[1]),.dout(n917),.clk(gclk));
	jxor g0854(.dina(w_n917_0[1]),.dinb(w_n869_0[1]),.dout(n918),.clk(gclk));
	jxor g0855(.dina(w_n918_0[1]),.dinb(w_n866_0[1]),.dout(n919),.clk(gclk));
	jxor g0856(.dina(w_n919_0[1]),.dinb(w_n864_0[1]),.dout(n920),.clk(gclk));
	jxor g0857(.dina(w_n920_0[1]),.dinb(w_n861_0[1]),.dout(n921),.clk(gclk));
	jxor g0858(.dina(w_n921_0[1]),.dinb(w_n859_0[1]),.dout(n922),.clk(gclk));
	jxor g0859(.dina(w_n922_0[1]),.dinb(w_n856_0[1]),.dout(n923),.clk(gclk));
	jxor g0860(.dina(w_n923_0[1]),.dinb(w_n854_0[1]),.dout(n924),.clk(gclk));
	jxor g0861(.dina(w_n924_0[1]),.dinb(w_n851_0[1]),.dout(n925),.clk(gclk));
	jxor g0862(.dina(w_n925_0[1]),.dinb(w_n849_0[1]),.dout(n926),.clk(gclk));
	jxor g0863(.dina(w_n926_0[1]),.dinb(w_n846_0[1]),.dout(n927),.clk(gclk));
	jxor g0864(.dina(w_n927_0[2]),.dinb(w_n844_0[2]),.dout(n928),.clk(gclk));
	jxor g0865(.dina(n928),.dinb(w_dff_B_7RVIsGbA0_1),.dout(n929),.clk(gclk));
	jxor g0866(.dina(w_n929_0[1]),.dinb(w_n839_0[1]),.dout(n930),.clk(gclk));
	jxor g0867(.dina(w_n930_0[1]),.dinb(w_n835_0[1]),.dout(n931),.clk(gclk));
	jxor g0868(.dina(w_n931_0[1]),.dinb(w_n834_0[1]),.dout(n932),.clk(gclk));
	jxor g0869(.dina(w_n932_0[1]),.dinb(w_dff_B_eG6R2dfb6_1),.dout(w_dff_A_jiWzWt4L4_2),.clk(gclk));
	jnot g0870(.din(w_n931_0[0]),.dout(n934),.clk(gclk));
	jor g0871(.dina(n934),.dinb(w_n834_0[0]),.dout(n935),.clk(gclk));
	jor g0872(.dina(w_n932_0[0]),.dinb(w_n829_0[0]),.dout(n936),.clk(gclk));
	jand g0873(.dina(n936),.dinb(w_dff_B_2Jd0iHVW5_1),.dout(n937),.clk(gclk));
	jand g0874(.dina(w_G528gat_7[0]),.dinb(w_G18gat_2[1]),.dout(n938),.clk(gclk));
	jnot g0875(.din(w_n929_0[0]),.dout(n939),.clk(gclk));
	jor g0876(.dina(n939),.dinb(w_n839_0[0]),.dout(n940),.clk(gclk));
	jor g0877(.dina(w_n930_0[0]),.dinb(w_n835_0[0]),.dout(n941),.clk(gclk));
	jand g0878(.dina(n941),.dinb(w_dff_B_sU9bcwMw6_1),.dout(n942),.clk(gclk));
	jand g0879(.dina(w_G511gat_6[2]),.dinb(w_G35gat_2[2]),.dout(n943),.clk(gclk));
	jand g0880(.dina(w_n927_0[1]),.dinb(w_n844_0[1]),.dout(n944),.clk(gclk));
	jnot g0881(.din(n944),.dout(n945),.clk(gclk));
	jnot g0882(.din(w_n927_0[0]),.dout(n946),.clk(gclk));
	jxor g0883(.dina(n946),.dinb(w_n844_0[0]),.dout(n947),.clk(gclk));
	jor g0884(.dina(n947),.dinb(w_n840_0[0]),.dout(n948),.clk(gclk));
	jand g0885(.dina(n948),.dinb(n945),.dout(n949),.clk(gclk));
	jand g0886(.dina(w_G494gat_6[1]),.dinb(w_G52gat_3[0]),.dout(n950),.clk(gclk));
	jnot g0887(.din(n950),.dout(n951),.clk(gclk));
	jand g0888(.dina(w_n925_0[0]),.dinb(w_n849_0[0]),.dout(n952),.clk(gclk));
	jand g0889(.dina(w_n926_0[0]),.dinb(w_n846_0[0]),.dout(n953),.clk(gclk));
	jor g0890(.dina(n953),.dinb(w_dff_B_veTUZf680_1),.dout(n954),.clk(gclk));
	jand g0891(.dina(w_G477gat_6[0]),.dinb(w_G69gat_3[1]),.dout(n955),.clk(gclk));
	jnot g0892(.din(n955),.dout(n956),.clk(gclk));
	jand g0893(.dina(w_n923_0[0]),.dinb(w_n854_0[0]),.dout(n957),.clk(gclk));
	jand g0894(.dina(w_n924_0[0]),.dinb(w_n851_0[0]),.dout(n958),.clk(gclk));
	jor g0895(.dina(n958),.dinb(w_dff_B_pBI9Lvgg8_1),.dout(n959),.clk(gclk));
	jand g0896(.dina(w_G460gat_5[2]),.dinb(w_G86gat_3[2]),.dout(n960),.clk(gclk));
	jnot g0897(.din(n960),.dout(n961),.clk(gclk));
	jand g0898(.dina(w_n921_0[0]),.dinb(w_n859_0[0]),.dout(n962),.clk(gclk));
	jand g0899(.dina(w_n922_0[0]),.dinb(w_n856_0[0]),.dout(n963),.clk(gclk));
	jor g0900(.dina(n963),.dinb(w_dff_B_hgj8ijXl0_1),.dout(n964),.clk(gclk));
	jand g0901(.dina(w_G443gat_5[1]),.dinb(w_G103gat_4[0]),.dout(n965),.clk(gclk));
	jnot g0902(.din(n965),.dout(n966),.clk(gclk));
	jand g0903(.dina(w_n919_0[0]),.dinb(w_n864_0[0]),.dout(n967),.clk(gclk));
	jand g0904(.dina(w_n920_0[0]),.dinb(w_n861_0[0]),.dout(n968),.clk(gclk));
	jor g0905(.dina(n968),.dinb(w_dff_B_E28e5hOE1_1),.dout(n969),.clk(gclk));
	jand g0906(.dina(w_G426gat_5[0]),.dinb(w_G120gat_4[1]),.dout(n970),.clk(gclk));
	jnot g0907(.din(n970),.dout(n971),.clk(gclk));
	jand g0908(.dina(w_n917_0[0]),.dinb(w_n869_0[0]),.dout(n972),.clk(gclk));
	jand g0909(.dina(w_n918_0[0]),.dinb(w_n866_0[0]),.dout(n973),.clk(gclk));
	jor g0910(.dina(n973),.dinb(w_dff_B_EmgwCGB41_1),.dout(n974),.clk(gclk));
	jand g0911(.dina(w_G409gat_4[2]),.dinb(w_G137gat_4[2]),.dout(n975),.clk(gclk));
	jnot g0912(.din(n975),.dout(n976),.clk(gclk));
	jand g0913(.dina(w_n915_0[0]),.dinb(w_n874_0[0]),.dout(n977),.clk(gclk));
	jand g0914(.dina(w_n916_0[0]),.dinb(w_n871_0[0]),.dout(n978),.clk(gclk));
	jor g0915(.dina(n978),.dinb(w_dff_B_nncCmUwm5_1),.dout(n979),.clk(gclk));
	jand g0916(.dina(w_G392gat_4[1]),.dinb(w_G154gat_5[0]),.dout(n980),.clk(gclk));
	jnot g0917(.din(n980),.dout(n981),.clk(gclk));
	jand g0918(.dina(w_n913_0[0]),.dinb(w_n879_0[0]),.dout(n982),.clk(gclk));
	jand g0919(.dina(w_n914_0[0]),.dinb(w_n876_0[0]),.dout(n983),.clk(gclk));
	jor g0920(.dina(n983),.dinb(w_dff_B_og15hhse0_1),.dout(n984),.clk(gclk));
	jand g0921(.dina(w_G375gat_4[0]),.dinb(w_G171gat_5[1]),.dout(n985),.clk(gclk));
	jnot g0922(.din(n985),.dout(n986),.clk(gclk));
	jand g0923(.dina(w_n911_0[0]),.dinb(w_n884_0[0]),.dout(n987),.clk(gclk));
	jand g0924(.dina(w_n912_0[0]),.dinb(w_n881_0[0]),.dout(n988),.clk(gclk));
	jor g0925(.dina(n988),.dinb(w_dff_B_qeu9lj3P5_1),.dout(n989),.clk(gclk));
	jand g0926(.dina(w_G358gat_3[2]),.dinb(w_G188gat_5[2]),.dout(n990),.clk(gclk));
	jnot g0927(.din(n990),.dout(n991),.clk(gclk));
	jand g0928(.dina(w_n909_0[0]),.dinb(w_n889_0[0]),.dout(n992),.clk(gclk));
	jand g0929(.dina(w_n910_0[0]),.dinb(w_n886_0[0]),.dout(n993),.clk(gclk));
	jor g0930(.dina(n993),.dinb(w_dff_B_OuzEvqxX7_1),.dout(n994),.clk(gclk));
	jand g0931(.dina(w_G341gat_3[1]),.dinb(w_G205gat_6[0]),.dout(n995),.clk(gclk));
	jnot g0932(.din(n995),.dout(n996),.clk(gclk));
	jand g0933(.dina(w_n907_0[0]),.dinb(w_n895_0[0]),.dout(n997),.clk(gclk));
	jand g0934(.dina(w_n908_0[0]),.dinb(w_n891_0[0]),.dout(n998),.clk(gclk));
	jor g0935(.dina(n998),.dinb(w_dff_B_UFwAyNCv0_1),.dout(n999),.clk(gclk));
	jand g0936(.dina(w_G324gat_3[0]),.dinb(w_G222gat_6[1]),.dout(n1000),.clk(gclk));
	jnot g0937(.din(n1000),.dout(n1001),.clk(gclk));
	jnot g0938(.din(w_n896_0[0]),.dout(n1002),.clk(gclk));
	jnot g0939(.din(w_n906_0[0]),.dout(n1003),.clk(gclk));
	jand g0940(.dina(n1003),.dinb(w_dff_B_rf367TDu7_1),.dout(n1004),.clk(gclk));
	jor g0941(.dina(n1004),.dinb(w_n903_0[0]),.dout(n1005),.clk(gclk));
	jand g0942(.dina(w_G307gat_3[0]),.dinb(w_G239gat_6[2]),.dout(n1006),.clk(gclk));
	jand g0943(.dina(w_G290gat_2[1]),.dinb(w_G256gat_7[0]),.dout(n1007),.clk(gclk));
	jnot g0944(.din(n1007),.dout(n1008),.clk(gclk));
	jor g0945(.dina(w_n1008_0[1]),.dinb(w_n793_0[0]),.dout(n1009),.clk(gclk));
	jxor g0946(.dina(w_n1009_0[1]),.dinb(w_n1006_0[1]),.dout(n1010),.clk(gclk));
	jxor g0947(.dina(w_n1010_0[1]),.dinb(w_n1005_0[1]),.dout(n1011),.clk(gclk));
	jxor g0948(.dina(w_n1011_0[1]),.dinb(w_n1001_0[1]),.dout(n1012),.clk(gclk));
	jxor g0949(.dina(w_n1012_0[1]),.dinb(w_n999_0[1]),.dout(n1013),.clk(gclk));
	jxor g0950(.dina(w_n1013_0[1]),.dinb(w_n996_0[1]),.dout(n1014),.clk(gclk));
	jxor g0951(.dina(w_n1014_0[1]),.dinb(w_n994_0[1]),.dout(n1015),.clk(gclk));
	jxor g0952(.dina(w_n1015_0[1]),.dinb(w_n991_0[1]),.dout(n1016),.clk(gclk));
	jxor g0953(.dina(w_n1016_0[1]),.dinb(w_n989_0[1]),.dout(n1017),.clk(gclk));
	jxor g0954(.dina(w_n1017_0[1]),.dinb(w_n986_0[1]),.dout(n1018),.clk(gclk));
	jxor g0955(.dina(w_n1018_0[1]),.dinb(w_n984_0[1]),.dout(n1019),.clk(gclk));
	jxor g0956(.dina(w_n1019_0[1]),.dinb(w_n981_0[1]),.dout(n1020),.clk(gclk));
	jxor g0957(.dina(w_n1020_0[1]),.dinb(w_n979_0[1]),.dout(n1021),.clk(gclk));
	jxor g0958(.dina(w_n1021_0[1]),.dinb(w_n976_0[1]),.dout(n1022),.clk(gclk));
	jxor g0959(.dina(w_n1022_0[1]),.dinb(w_n974_0[1]),.dout(n1023),.clk(gclk));
	jxor g0960(.dina(w_n1023_0[1]),.dinb(w_n971_0[1]),.dout(n1024),.clk(gclk));
	jxor g0961(.dina(w_n1024_0[1]),.dinb(w_n969_0[1]),.dout(n1025),.clk(gclk));
	jxor g0962(.dina(w_n1025_0[1]),.dinb(w_n966_0[1]),.dout(n1026),.clk(gclk));
	jxor g0963(.dina(w_n1026_0[1]),.dinb(w_n964_0[1]),.dout(n1027),.clk(gclk));
	jxor g0964(.dina(w_n1027_0[1]),.dinb(w_n961_0[1]),.dout(n1028),.clk(gclk));
	jxor g0965(.dina(w_n1028_0[1]),.dinb(w_n959_0[1]),.dout(n1029),.clk(gclk));
	jxor g0966(.dina(w_n1029_0[1]),.dinb(w_n956_0[1]),.dout(n1030),.clk(gclk));
	jxor g0967(.dina(w_n1030_0[1]),.dinb(w_n954_0[1]),.dout(n1031),.clk(gclk));
	jxor g0968(.dina(w_n1031_0[1]),.dinb(w_n951_0[1]),.dout(n1032),.clk(gclk));
	jxor g0969(.dina(w_n1032_0[1]),.dinb(w_n949_0[1]),.dout(n1033),.clk(gclk));
	jxor g0970(.dina(w_n1033_0[1]),.dinb(w_n943_0[1]),.dout(n1034),.clk(gclk));
	jnot g0971(.din(w_n1034_0[1]),.dout(n1035),.clk(gclk));
	jxor g0972(.dina(w_n1035_0[1]),.dinb(w_n942_0[2]),.dout(n1036),.clk(gclk));
	jxor g0973(.dina(n1036),.dinb(w_n938_0[1]),.dout(n1037),.clk(gclk));
	jxor g0974(.dina(w_n1037_0[1]),.dinb(w_n937_0[1]),.dout(w_dff_A_9rj7sGa51_2),.clk(gclk));
	jand g0975(.dina(w_n1037_0[0]),.dinb(w_n937_0[0]),.dout(n1039),.clk(gclk));
	jor g0976(.dina(w_n1035_0[0]),.dinb(w_n942_0[1]),.dout(n1040),.clk(gclk));
	jxor g0977(.dina(w_n1034_0[0]),.dinb(w_n942_0[0]),.dout(n1041),.clk(gclk));
	jor g0978(.dina(n1041),.dinb(w_n938_0[0]),.dout(n1042),.clk(gclk));
	jand g0979(.dina(n1042),.dinb(w_dff_B_RiwhK7vq5_1),.dout(n1043),.clk(gclk));
	jand g0980(.dina(w_G528gat_6[2]),.dinb(w_G35gat_2[1]),.dout(n1044),.clk(gclk));
	jnot g0981(.din(w_n1032_0[0]),.dout(n1045),.clk(gclk));
	jor g0982(.dina(n1045),.dinb(w_n949_0[0]),.dout(n1046),.clk(gclk));
	jor g0983(.dina(w_n1033_0[0]),.dinb(w_n943_0[0]),.dout(n1047),.clk(gclk));
	jand g0984(.dina(n1047),.dinb(w_dff_B_C5C6vHsw0_1),.dout(n1048),.clk(gclk));
	jand g0985(.dina(w_G511gat_6[1]),.dinb(w_G52gat_2[2]),.dout(n1049),.clk(gclk));
	jand g0986(.dina(w_n1030_0[0]),.dinb(w_n954_0[0]),.dout(n1050),.clk(gclk));
	jand g0987(.dina(w_n1031_0[0]),.dinb(w_n951_0[0]),.dout(n1051),.clk(gclk));
	jor g0988(.dina(n1051),.dinb(w_dff_B_ReanFiuq9_1),.dout(n1052),.clk(gclk));
	jand g0989(.dina(w_G494gat_6[0]),.dinb(w_G69gat_3[0]),.dout(n1053),.clk(gclk));
	jnot g0990(.din(n1053),.dout(n1054),.clk(gclk));
	jand g0991(.dina(w_n1028_0[0]),.dinb(w_n959_0[0]),.dout(n1055),.clk(gclk));
	jand g0992(.dina(w_n1029_0[0]),.dinb(w_n956_0[0]),.dout(n1056),.clk(gclk));
	jor g0993(.dina(n1056),.dinb(w_dff_B_e7fGPhgE3_1),.dout(n1057),.clk(gclk));
	jand g0994(.dina(w_G477gat_5[2]),.dinb(w_G86gat_3[1]),.dout(n1058),.clk(gclk));
	jnot g0995(.din(n1058),.dout(n1059),.clk(gclk));
	jand g0996(.dina(w_n1026_0[0]),.dinb(w_n964_0[0]),.dout(n1060),.clk(gclk));
	jand g0997(.dina(w_n1027_0[0]),.dinb(w_n961_0[0]),.dout(n1061),.clk(gclk));
	jor g0998(.dina(n1061),.dinb(w_dff_B_5UvB3LGI1_1),.dout(n1062),.clk(gclk));
	jand g0999(.dina(w_G460gat_5[1]),.dinb(w_G103gat_3[2]),.dout(n1063),.clk(gclk));
	jnot g1000(.din(n1063),.dout(n1064),.clk(gclk));
	jand g1001(.dina(w_n1024_0[0]),.dinb(w_n969_0[0]),.dout(n1065),.clk(gclk));
	jand g1002(.dina(w_n1025_0[0]),.dinb(w_n966_0[0]),.dout(n1066),.clk(gclk));
	jor g1003(.dina(n1066),.dinb(w_dff_B_oBxkf0G21_1),.dout(n1067),.clk(gclk));
	jand g1004(.dina(w_G443gat_5[0]),.dinb(w_G120gat_4[0]),.dout(n1068),.clk(gclk));
	jnot g1005(.din(n1068),.dout(n1069),.clk(gclk));
	jand g1006(.dina(w_n1022_0[0]),.dinb(w_n974_0[0]),.dout(n1070),.clk(gclk));
	jand g1007(.dina(w_n1023_0[0]),.dinb(w_n971_0[0]),.dout(n1071),.clk(gclk));
	jor g1008(.dina(n1071),.dinb(w_dff_B_Te2DMkeV2_1),.dout(n1072),.clk(gclk));
	jand g1009(.dina(w_G426gat_4[2]),.dinb(w_G137gat_4[1]),.dout(n1073),.clk(gclk));
	jnot g1010(.din(n1073),.dout(n1074),.clk(gclk));
	jand g1011(.dina(w_n1020_0[0]),.dinb(w_n979_0[0]),.dout(n1075),.clk(gclk));
	jand g1012(.dina(w_n1021_0[0]),.dinb(w_n976_0[0]),.dout(n1076),.clk(gclk));
	jor g1013(.dina(n1076),.dinb(w_dff_B_EkaceZ4V3_1),.dout(n1077),.clk(gclk));
	jand g1014(.dina(w_G409gat_4[1]),.dinb(w_G154gat_4[2]),.dout(n1078),.clk(gclk));
	jnot g1015(.din(n1078),.dout(n1079),.clk(gclk));
	jand g1016(.dina(w_n1018_0[0]),.dinb(w_n984_0[0]),.dout(n1080),.clk(gclk));
	jand g1017(.dina(w_n1019_0[0]),.dinb(w_n981_0[0]),.dout(n1081),.clk(gclk));
	jor g1018(.dina(n1081),.dinb(w_dff_B_RJaWybtq6_1),.dout(n1082),.clk(gclk));
	jand g1019(.dina(w_G392gat_4[0]),.dinb(w_G171gat_5[0]),.dout(n1083),.clk(gclk));
	jnot g1020(.din(n1083),.dout(n1084),.clk(gclk));
	jand g1021(.dina(w_n1016_0[0]),.dinb(w_n989_0[0]),.dout(n1085),.clk(gclk));
	jand g1022(.dina(w_n1017_0[0]),.dinb(w_n986_0[0]),.dout(n1086),.clk(gclk));
	jor g1023(.dina(n1086),.dinb(w_dff_B_gCRseKSX3_1),.dout(n1087),.clk(gclk));
	jand g1024(.dina(w_G375gat_3[2]),.dinb(w_G188gat_5[1]),.dout(n1088),.clk(gclk));
	jnot g1025(.din(n1088),.dout(n1089),.clk(gclk));
	jand g1026(.dina(w_n1014_0[0]),.dinb(w_n994_0[0]),.dout(n1090),.clk(gclk));
	jand g1027(.dina(w_n1015_0[0]),.dinb(w_n991_0[0]),.dout(n1091),.clk(gclk));
	jor g1028(.dina(n1091),.dinb(w_dff_B_qDrVah190_1),.dout(n1092),.clk(gclk));
	jand g1029(.dina(w_G358gat_3[1]),.dinb(w_G205gat_5[2]),.dout(n1093),.clk(gclk));
	jnot g1030(.din(n1093),.dout(n1094),.clk(gclk));
	jand g1031(.dina(w_n1012_0[0]),.dinb(w_n999_0[0]),.dout(n1095),.clk(gclk));
	jand g1032(.dina(w_n1013_0[0]),.dinb(w_n996_0[0]),.dout(n1096),.clk(gclk));
	jor g1033(.dina(n1096),.dinb(w_dff_B_fD5g9lbL1_1),.dout(n1097),.clk(gclk));
	jand g1034(.dina(w_G341gat_3[0]),.dinb(w_G222gat_6[0]),.dout(n1098),.clk(gclk));
	jnot g1035(.din(n1098),.dout(n1099),.clk(gclk));
	jand g1036(.dina(w_n1010_0[0]),.dinb(w_n1005_0[0]),.dout(n1100),.clk(gclk));
	jand g1037(.dina(w_n1011_0[0]),.dinb(w_n1001_0[0]),.dout(n1101),.clk(gclk));
	jor g1038(.dina(n1101),.dinb(w_dff_B_BFY5D3Vg9_1),.dout(n1102),.clk(gclk));
	jand g1039(.dina(w_G324gat_2[2]),.dinb(w_G239gat_6[1]),.dout(n1103),.clk(gclk));
	jand g1040(.dina(w_G307gat_2[2]),.dinb(w_G256gat_6[2]),.dout(n1104),.clk(gclk));
	jnot g1041(.din(w_n1006_0[0]),.dout(n1105),.clk(gclk));
	jnot g1042(.din(w_n1009_0[0]),.dout(n1106),.clk(gclk));
	jand g1043(.dina(n1106),.dinb(w_dff_B_hodFMUDZ4_1),.dout(n1107),.clk(gclk));
	jor g1044(.dina(n1107),.dinb(w_n1008_0[0]),.dout(n1108),.clk(gclk));
	jnot g1045(.din(n1108),.dout(n1109),.clk(gclk));
	jor g1046(.dina(w_n1109_0[1]),.dinb(w_dff_B_rP85qQ8J0_1),.dout(n1110),.clk(gclk));
	jand g1047(.dina(w_n1109_0[0]),.dinb(w_G307gat_2[1]),.dout(n1111),.clk(gclk));
	jnot g1048(.din(n1111),.dout(n1112),.clk(gclk));
	jand g1049(.dina(n1112),.dinb(w_n1110_0[1]),.dout(n1113),.clk(gclk));
	jnot g1050(.din(n1113),.dout(n1114),.clk(gclk));
	jxor g1051(.dina(w_n1114_0[1]),.dinb(w_n1103_0[1]),.dout(n1115),.clk(gclk));
	jxor g1052(.dina(w_n1115_0[1]),.dinb(w_n1102_0[1]),.dout(n1116),.clk(gclk));
	jxor g1053(.dina(w_n1116_0[1]),.dinb(w_n1099_0[1]),.dout(n1117),.clk(gclk));
	jxor g1054(.dina(w_n1117_0[1]),.dinb(w_n1097_0[1]),.dout(n1118),.clk(gclk));
	jxor g1055(.dina(w_n1118_0[1]),.dinb(w_n1094_0[1]),.dout(n1119),.clk(gclk));
	jxor g1056(.dina(w_n1119_0[1]),.dinb(w_n1092_0[1]),.dout(n1120),.clk(gclk));
	jxor g1057(.dina(w_n1120_0[1]),.dinb(w_n1089_0[1]),.dout(n1121),.clk(gclk));
	jxor g1058(.dina(w_n1121_0[1]),.dinb(w_n1087_0[1]),.dout(n1122),.clk(gclk));
	jxor g1059(.dina(w_n1122_0[1]),.dinb(w_n1084_0[1]),.dout(n1123),.clk(gclk));
	jxor g1060(.dina(w_n1123_0[1]),.dinb(w_n1082_0[1]),.dout(n1124),.clk(gclk));
	jxor g1061(.dina(w_n1124_0[1]),.dinb(w_n1079_0[1]),.dout(n1125),.clk(gclk));
	jxor g1062(.dina(w_n1125_0[1]),.dinb(w_n1077_0[1]),.dout(n1126),.clk(gclk));
	jxor g1063(.dina(w_n1126_0[1]),.dinb(w_n1074_0[1]),.dout(n1127),.clk(gclk));
	jxor g1064(.dina(w_n1127_0[1]),.dinb(w_n1072_0[1]),.dout(n1128),.clk(gclk));
	jxor g1065(.dina(w_n1128_0[1]),.dinb(w_n1069_0[1]),.dout(n1129),.clk(gclk));
	jxor g1066(.dina(w_n1129_0[1]),.dinb(w_n1067_0[1]),.dout(n1130),.clk(gclk));
	jxor g1067(.dina(w_n1130_0[1]),.dinb(w_n1064_0[1]),.dout(n1131),.clk(gclk));
	jxor g1068(.dina(w_n1131_0[1]),.dinb(w_n1062_0[1]),.dout(n1132),.clk(gclk));
	jxor g1069(.dina(w_n1132_0[1]),.dinb(w_n1059_0[1]),.dout(n1133),.clk(gclk));
	jxor g1070(.dina(w_n1133_0[1]),.dinb(w_n1057_0[1]),.dout(n1134),.clk(gclk));
	jxor g1071(.dina(w_n1134_0[1]),.dinb(w_n1054_0[1]),.dout(n1135),.clk(gclk));
	jxor g1072(.dina(w_n1135_0[1]),.dinb(w_n1052_0[1]),.dout(n1136),.clk(gclk));
	jnot g1073(.din(n1136),.dout(n1137),.clk(gclk));
	jxor g1074(.dina(w_n1137_0[1]),.dinb(w_n1049_0[1]),.dout(n1138),.clk(gclk));
	jxor g1075(.dina(w_n1138_0[1]),.dinb(w_n1048_0[1]),.dout(n1139),.clk(gclk));
	jxor g1076(.dina(w_n1139_0[1]),.dinb(w_n1044_0[1]),.dout(n1140),.clk(gclk));
	jxor g1077(.dina(w_n1140_0[1]),.dinb(w_n1043_0[1]),.dout(n1141),.clk(gclk));
	jnot g1078(.din(w_n1141_0[1]),.dout(n1142),.clk(gclk));
	jxor g1079(.dina(n1142),.dinb(w_n1039_0[1]),.dout(w_dff_A_BV07xd3i5_2),.clk(gclk));
	jnot g1080(.din(w_n1140_0[0]),.dout(n1144),.clk(gclk));
	jor g1081(.dina(n1144),.dinb(w_n1043_0[0]),.dout(n1145),.clk(gclk));
	jor g1082(.dina(w_n1141_0[0]),.dinb(w_n1039_0[0]),.dout(n1146),.clk(gclk));
	jand g1083(.dina(n1146),.dinb(w_dff_B_OmGa2UCE3_1),.dout(n1147),.clk(gclk));
	jnot g1084(.din(w_n1138_0[0]),.dout(n1148),.clk(gclk));
	jor g1085(.dina(n1148),.dinb(w_n1048_0[0]),.dout(n1149),.clk(gclk));
	jor g1086(.dina(w_n1139_0[0]),.dinb(w_n1044_0[0]),.dout(n1150),.clk(gclk));
	jand g1087(.dina(n1150),.dinb(n1149),.dout(n1151),.clk(gclk));
	jand g1088(.dina(w_G528gat_6[1]),.dinb(w_G52gat_2[1]),.dout(n1152),.clk(gclk));
	jand g1089(.dina(w_n1135_0[0]),.dinb(w_n1052_0[0]),.dout(n1153),.clk(gclk));
	jnot g1090(.din(n1153),.dout(n1154),.clk(gclk));
	jor g1091(.dina(w_n1137_0[0]),.dinb(w_n1049_0[0]),.dout(n1155),.clk(gclk));
	jand g1092(.dina(n1155),.dinb(w_dff_B_DOH2dNe61_1),.dout(n1156),.clk(gclk));
	jand g1093(.dina(w_G511gat_6[0]),.dinb(w_G69gat_2[2]),.dout(n1157),.clk(gclk));
	jnot g1094(.din(n1157),.dout(n1158),.clk(gclk));
	jand g1095(.dina(w_n1133_0[0]),.dinb(w_n1057_0[0]),.dout(n1159),.clk(gclk));
	jand g1096(.dina(w_n1134_0[0]),.dinb(w_n1054_0[0]),.dout(n1160),.clk(gclk));
	jor g1097(.dina(n1160),.dinb(w_dff_B_1FdTulTQ5_1),.dout(n1161),.clk(gclk));
	jand g1098(.dina(w_G494gat_5[2]),.dinb(w_G86gat_3[0]),.dout(n1162),.clk(gclk));
	jnot g1099(.din(n1162),.dout(n1163),.clk(gclk));
	jand g1100(.dina(w_n1131_0[0]),.dinb(w_n1062_0[0]),.dout(n1164),.clk(gclk));
	jand g1101(.dina(w_n1132_0[0]),.dinb(w_n1059_0[0]),.dout(n1165),.clk(gclk));
	jor g1102(.dina(n1165),.dinb(w_dff_B_adC3VRFf2_1),.dout(n1166),.clk(gclk));
	jand g1103(.dina(w_G477gat_5[1]),.dinb(w_G103gat_3[1]),.dout(n1167),.clk(gclk));
	jnot g1104(.din(n1167),.dout(n1168),.clk(gclk));
	jand g1105(.dina(w_n1129_0[0]),.dinb(w_n1067_0[0]),.dout(n1169),.clk(gclk));
	jand g1106(.dina(w_n1130_0[0]),.dinb(w_n1064_0[0]),.dout(n1170),.clk(gclk));
	jor g1107(.dina(n1170),.dinb(w_dff_B_XCy6AqqE0_1),.dout(n1171),.clk(gclk));
	jand g1108(.dina(w_G460gat_5[0]),.dinb(w_G120gat_3[2]),.dout(n1172),.clk(gclk));
	jnot g1109(.din(n1172),.dout(n1173),.clk(gclk));
	jand g1110(.dina(w_n1127_0[0]),.dinb(w_n1072_0[0]),.dout(n1174),.clk(gclk));
	jand g1111(.dina(w_n1128_0[0]),.dinb(w_n1069_0[0]),.dout(n1175),.clk(gclk));
	jor g1112(.dina(n1175),.dinb(w_dff_B_G4BLumyx3_1),.dout(n1176),.clk(gclk));
	jand g1113(.dina(w_G443gat_4[2]),.dinb(w_G137gat_4[0]),.dout(n1177),.clk(gclk));
	jnot g1114(.din(n1177),.dout(n1178),.clk(gclk));
	jand g1115(.dina(w_n1125_0[0]),.dinb(w_n1077_0[0]),.dout(n1179),.clk(gclk));
	jand g1116(.dina(w_n1126_0[0]),.dinb(w_n1074_0[0]),.dout(n1180),.clk(gclk));
	jor g1117(.dina(n1180),.dinb(w_dff_B_buQPiXvj6_1),.dout(n1181),.clk(gclk));
	jand g1118(.dina(w_G426gat_4[1]),.dinb(w_G154gat_4[1]),.dout(n1182),.clk(gclk));
	jnot g1119(.din(n1182),.dout(n1183),.clk(gclk));
	jand g1120(.dina(w_n1123_0[0]),.dinb(w_n1082_0[0]),.dout(n1184),.clk(gclk));
	jand g1121(.dina(w_n1124_0[0]),.dinb(w_n1079_0[0]),.dout(n1185),.clk(gclk));
	jor g1122(.dina(n1185),.dinb(w_dff_B_fvxKhTZJ1_1),.dout(n1186),.clk(gclk));
	jand g1123(.dina(w_G409gat_4[0]),.dinb(w_G171gat_4[2]),.dout(n1187),.clk(gclk));
	jnot g1124(.din(n1187),.dout(n1188),.clk(gclk));
	jand g1125(.dina(w_n1121_0[0]),.dinb(w_n1087_0[0]),.dout(n1189),.clk(gclk));
	jand g1126(.dina(w_n1122_0[0]),.dinb(w_n1084_0[0]),.dout(n1190),.clk(gclk));
	jor g1127(.dina(n1190),.dinb(w_dff_B_OGayP6UF0_1),.dout(n1191),.clk(gclk));
	jand g1128(.dina(w_G392gat_3[2]),.dinb(w_G188gat_5[0]),.dout(n1192),.clk(gclk));
	jnot g1129(.din(n1192),.dout(n1193),.clk(gclk));
	jand g1130(.dina(w_n1119_0[0]),.dinb(w_n1092_0[0]),.dout(n1194),.clk(gclk));
	jand g1131(.dina(w_n1120_0[0]),.dinb(w_n1089_0[0]),.dout(n1195),.clk(gclk));
	jor g1132(.dina(n1195),.dinb(w_dff_B_pdx9xkB96_1),.dout(n1196),.clk(gclk));
	jand g1133(.dina(w_G375gat_3[1]),.dinb(w_G205gat_5[1]),.dout(n1197),.clk(gclk));
	jnot g1134(.din(n1197),.dout(n1198),.clk(gclk));
	jand g1135(.dina(w_n1117_0[0]),.dinb(w_n1097_0[0]),.dout(n1199),.clk(gclk));
	jand g1136(.dina(w_n1118_0[0]),.dinb(w_n1094_0[0]),.dout(n1200),.clk(gclk));
	jor g1137(.dina(n1200),.dinb(w_dff_B_VX0TK40R4_1),.dout(n1201),.clk(gclk));
	jand g1138(.dina(w_G358gat_3[0]),.dinb(w_G222gat_5[2]),.dout(n1202),.clk(gclk));
	jnot g1139(.din(n1202),.dout(n1203),.clk(gclk));
	jand g1140(.dina(w_n1115_0[0]),.dinb(w_n1102_0[0]),.dout(n1204),.clk(gclk));
	jand g1141(.dina(w_n1116_0[0]),.dinb(w_n1099_0[0]),.dout(n1205),.clk(gclk));
	jor g1142(.dina(n1205),.dinb(w_dff_B_eYIqDh9G5_1),.dout(n1206),.clk(gclk));
	jand g1143(.dina(w_G341gat_2[2]),.dinb(w_G239gat_6[0]),.dout(n1207),.clk(gclk));
	jand g1144(.dina(w_G324gat_2[1]),.dinb(w_G256gat_6[1]),.dout(n1208),.clk(gclk));
	jor g1145(.dina(w_n1114_0[0]),.dinb(w_n1103_0[0]),.dout(n1209),.clk(gclk));
	jand g1146(.dina(n1209),.dinb(w_n1110_0[0]),.dout(n1210),.clk(gclk));
	jxor g1147(.dina(w_n1210_0[1]),.dinb(w_n1208_0[1]),.dout(n1211),.clk(gclk));
	jnot g1148(.din(n1211),.dout(n1212),.clk(gclk));
	jxor g1149(.dina(w_n1212_0[1]),.dinb(w_n1207_0[1]),.dout(n1213),.clk(gclk));
	jxor g1150(.dina(w_n1213_0[1]),.dinb(w_n1206_0[1]),.dout(n1214),.clk(gclk));
	jxor g1151(.dina(w_n1214_0[1]),.dinb(w_n1203_0[1]),.dout(n1215),.clk(gclk));
	jxor g1152(.dina(w_n1215_0[1]),.dinb(w_n1201_0[1]),.dout(n1216),.clk(gclk));
	jxor g1153(.dina(w_n1216_0[1]),.dinb(w_n1198_0[1]),.dout(n1217),.clk(gclk));
	jxor g1154(.dina(w_n1217_0[1]),.dinb(w_n1196_0[1]),.dout(n1218),.clk(gclk));
	jxor g1155(.dina(w_n1218_0[1]),.dinb(w_n1193_0[1]),.dout(n1219),.clk(gclk));
	jxor g1156(.dina(w_n1219_0[1]),.dinb(w_n1191_0[1]),.dout(n1220),.clk(gclk));
	jxor g1157(.dina(w_n1220_0[1]),.dinb(w_n1188_0[1]),.dout(n1221),.clk(gclk));
	jxor g1158(.dina(w_n1221_0[1]),.dinb(w_n1186_0[1]),.dout(n1222),.clk(gclk));
	jxor g1159(.dina(w_n1222_0[1]),.dinb(w_n1183_0[1]),.dout(n1223),.clk(gclk));
	jxor g1160(.dina(w_n1223_0[1]),.dinb(w_n1181_0[1]),.dout(n1224),.clk(gclk));
	jxor g1161(.dina(w_n1224_0[1]),.dinb(w_n1178_0[1]),.dout(n1225),.clk(gclk));
	jxor g1162(.dina(w_n1225_0[1]),.dinb(w_n1176_0[1]),.dout(n1226),.clk(gclk));
	jxor g1163(.dina(w_n1226_0[1]),.dinb(w_n1173_0[1]),.dout(n1227),.clk(gclk));
	jxor g1164(.dina(w_n1227_0[1]),.dinb(w_n1171_0[1]),.dout(n1228),.clk(gclk));
	jxor g1165(.dina(w_n1228_0[1]),.dinb(w_n1168_0[1]),.dout(n1229),.clk(gclk));
	jxor g1166(.dina(w_n1229_0[1]),.dinb(w_n1166_0[1]),.dout(n1230),.clk(gclk));
	jxor g1167(.dina(w_n1230_0[1]),.dinb(w_n1163_0[1]),.dout(n1231),.clk(gclk));
	jxor g1168(.dina(w_n1231_0[1]),.dinb(w_n1161_0[1]),.dout(n1232),.clk(gclk));
	jxor g1169(.dina(w_n1232_0[1]),.dinb(w_n1158_0[1]),.dout(n1233),.clk(gclk));
	jnot g1170(.din(n1233),.dout(n1234),.clk(gclk));
	jxor g1171(.dina(w_n1234_0[1]),.dinb(w_n1156_0[1]),.dout(n1235),.clk(gclk));
	jnot g1172(.din(n1235),.dout(n1236),.clk(gclk));
	jxor g1173(.dina(w_n1236_0[1]),.dinb(w_n1152_0[1]),.dout(n1237),.clk(gclk));
	jxor g1174(.dina(w_n1237_0[1]),.dinb(w_n1151_0[1]),.dout(n1238),.clk(gclk));
	jnot g1175(.din(w_n1238_0[1]),.dout(n1239),.clk(gclk));
	jxor g1176(.dina(n1239),.dinb(w_n1147_0[1]),.dout(w_dff_A_9g6kPTWT1_2),.clk(gclk));
	jnot g1177(.din(w_n1237_0[0]),.dout(n1241),.clk(gclk));
	jor g1178(.dina(n1241),.dinb(w_n1151_0[0]),.dout(n1242),.clk(gclk));
	jor g1179(.dina(w_n1238_0[0]),.dinb(w_n1147_0[0]),.dout(n1243),.clk(gclk));
	jand g1180(.dina(n1243),.dinb(w_dff_B_BBetNlil1_1),.dout(n1244),.clk(gclk));
	jor g1181(.dina(w_n1234_0[0]),.dinb(w_n1156_0[0]),.dout(n1245),.clk(gclk));
	jor g1182(.dina(w_n1236_0[0]),.dinb(w_n1152_0[0]),.dout(n1246),.clk(gclk));
	jand g1183(.dina(n1246),.dinb(w_dff_B_JNPv3mIo9_1),.dout(n1247),.clk(gclk));
	jand g1184(.dina(w_G528gat_6[0]),.dinb(w_G69gat_2[1]),.dout(n1248),.clk(gclk));
	jand g1185(.dina(w_n1231_0[0]),.dinb(w_n1161_0[0]),.dout(n1249),.clk(gclk));
	jand g1186(.dina(w_n1232_0[0]),.dinb(w_n1158_0[0]),.dout(n1250),.clk(gclk));
	jor g1187(.dina(n1250),.dinb(w_dff_B_PO12R7st0_1),.dout(n1251),.clk(gclk));
	jand g1188(.dina(w_G511gat_5[2]),.dinb(w_G86gat_2[2]),.dout(n1252),.clk(gclk));
	jnot g1189(.din(n1252),.dout(n1253),.clk(gclk));
	jand g1190(.dina(w_n1229_0[0]),.dinb(w_n1166_0[0]),.dout(n1254),.clk(gclk));
	jand g1191(.dina(w_n1230_0[0]),.dinb(w_n1163_0[0]),.dout(n1255),.clk(gclk));
	jor g1192(.dina(n1255),.dinb(w_dff_B_lpCrGuqL4_1),.dout(n1256),.clk(gclk));
	jand g1193(.dina(w_G494gat_5[1]),.dinb(w_G103gat_3[0]),.dout(n1257),.clk(gclk));
	jnot g1194(.din(n1257),.dout(n1258),.clk(gclk));
	jand g1195(.dina(w_n1227_0[0]),.dinb(w_n1171_0[0]),.dout(n1259),.clk(gclk));
	jand g1196(.dina(w_n1228_0[0]),.dinb(w_n1168_0[0]),.dout(n1260),.clk(gclk));
	jor g1197(.dina(n1260),.dinb(w_dff_B_zK7yrA7e2_1),.dout(n1261),.clk(gclk));
	jand g1198(.dina(w_G477gat_5[0]),.dinb(w_G120gat_3[1]),.dout(n1262),.clk(gclk));
	jnot g1199(.din(n1262),.dout(n1263),.clk(gclk));
	jand g1200(.dina(w_n1225_0[0]),.dinb(w_n1176_0[0]),.dout(n1264),.clk(gclk));
	jand g1201(.dina(w_n1226_0[0]),.dinb(w_n1173_0[0]),.dout(n1265),.clk(gclk));
	jor g1202(.dina(n1265),.dinb(w_dff_B_pso4BWIG7_1),.dout(n1266),.clk(gclk));
	jand g1203(.dina(w_G460gat_4[2]),.dinb(w_G137gat_3[2]),.dout(n1267),.clk(gclk));
	jnot g1204(.din(n1267),.dout(n1268),.clk(gclk));
	jand g1205(.dina(w_n1223_0[0]),.dinb(w_n1181_0[0]),.dout(n1269),.clk(gclk));
	jand g1206(.dina(w_n1224_0[0]),.dinb(w_n1178_0[0]),.dout(n1270),.clk(gclk));
	jor g1207(.dina(n1270),.dinb(w_dff_B_ScPyrVF34_1),.dout(n1271),.clk(gclk));
	jand g1208(.dina(w_G443gat_4[1]),.dinb(w_G154gat_4[0]),.dout(n1272),.clk(gclk));
	jnot g1209(.din(n1272),.dout(n1273),.clk(gclk));
	jand g1210(.dina(w_n1221_0[0]),.dinb(w_n1186_0[0]),.dout(n1274),.clk(gclk));
	jand g1211(.dina(w_n1222_0[0]),.dinb(w_n1183_0[0]),.dout(n1275),.clk(gclk));
	jor g1212(.dina(n1275),.dinb(w_dff_B_2pzKa2wU6_1),.dout(n1276),.clk(gclk));
	jand g1213(.dina(w_G426gat_4[0]),.dinb(w_G171gat_4[1]),.dout(n1277),.clk(gclk));
	jnot g1214(.din(n1277),.dout(n1278),.clk(gclk));
	jand g1215(.dina(w_n1219_0[0]),.dinb(w_n1191_0[0]),.dout(n1279),.clk(gclk));
	jand g1216(.dina(w_n1220_0[0]),.dinb(w_n1188_0[0]),.dout(n1280),.clk(gclk));
	jor g1217(.dina(n1280),.dinb(w_dff_B_GEWdfR901_1),.dout(n1281),.clk(gclk));
	jand g1218(.dina(w_G409gat_3[2]),.dinb(w_G188gat_4[2]),.dout(n1282),.clk(gclk));
	jnot g1219(.din(n1282),.dout(n1283),.clk(gclk));
	jand g1220(.dina(w_n1217_0[0]),.dinb(w_n1196_0[0]),.dout(n1284),.clk(gclk));
	jand g1221(.dina(w_n1218_0[0]),.dinb(w_n1193_0[0]),.dout(n1285),.clk(gclk));
	jor g1222(.dina(n1285),.dinb(w_dff_B_sMQcSNB69_1),.dout(n1286),.clk(gclk));
	jand g1223(.dina(w_G392gat_3[1]),.dinb(w_G205gat_5[0]),.dout(n1287),.clk(gclk));
	jnot g1224(.din(n1287),.dout(n1288),.clk(gclk));
	jand g1225(.dina(w_n1215_0[0]),.dinb(w_n1201_0[0]),.dout(n1289),.clk(gclk));
	jand g1226(.dina(w_n1216_0[0]),.dinb(w_n1198_0[0]),.dout(n1290),.clk(gclk));
	jor g1227(.dina(n1290),.dinb(w_dff_B_Fo72BbEF4_1),.dout(n1291),.clk(gclk));
	jand g1228(.dina(w_G375gat_3[0]),.dinb(w_G222gat_5[1]),.dout(n1292),.clk(gclk));
	jnot g1229(.din(n1292),.dout(n1293),.clk(gclk));
	jand g1230(.dina(w_n1213_0[0]),.dinb(w_n1206_0[0]),.dout(n1294),.clk(gclk));
	jand g1231(.dina(w_n1214_0[0]),.dinb(w_n1203_0[0]),.dout(n1295),.clk(gclk));
	jor g1232(.dina(n1295),.dinb(w_dff_B_0Gb9Fong5_1),.dout(n1296),.clk(gclk));
	jand g1233(.dina(w_G358gat_2[2]),.dinb(w_G239gat_5[2]),.dout(n1297),.clk(gclk));
	jand g1234(.dina(w_G341gat_2[1]),.dinb(w_G256gat_6[0]),.dout(n1298),.clk(gclk));
	jor g1235(.dina(w_n1210_0[0]),.dinb(w_n1208_0[0]),.dout(n1299),.clk(gclk));
	jor g1236(.dina(w_n1212_0[0]),.dinb(w_n1207_0[0]),.dout(n1300),.clk(gclk));
	jand g1237(.dina(n1300),.dinb(w_dff_B_DCPQC2Kw1_1),.dout(n1301),.clk(gclk));
	jxor g1238(.dina(w_n1301_0[1]),.dinb(w_n1298_0[1]),.dout(n1302),.clk(gclk));
	jnot g1239(.din(n1302),.dout(n1303),.clk(gclk));
	jxor g1240(.dina(w_n1303_0[1]),.dinb(w_n1297_0[1]),.dout(n1304),.clk(gclk));
	jxor g1241(.dina(w_n1304_0[1]),.dinb(w_n1296_0[1]),.dout(n1305),.clk(gclk));
	jxor g1242(.dina(w_n1305_0[1]),.dinb(w_n1293_0[1]),.dout(n1306),.clk(gclk));
	jxor g1243(.dina(w_n1306_0[1]),.dinb(w_n1291_0[1]),.dout(n1307),.clk(gclk));
	jxor g1244(.dina(w_n1307_0[1]),.dinb(w_n1288_0[1]),.dout(n1308),.clk(gclk));
	jxor g1245(.dina(w_n1308_0[1]),.dinb(w_n1286_0[1]),.dout(n1309),.clk(gclk));
	jxor g1246(.dina(w_n1309_0[1]),.dinb(w_n1283_0[1]),.dout(n1310),.clk(gclk));
	jxor g1247(.dina(w_n1310_0[1]),.dinb(w_n1281_0[1]),.dout(n1311),.clk(gclk));
	jxor g1248(.dina(w_n1311_0[1]),.dinb(w_n1278_0[1]),.dout(n1312),.clk(gclk));
	jxor g1249(.dina(w_n1312_0[1]),.dinb(w_n1276_0[1]),.dout(n1313),.clk(gclk));
	jxor g1250(.dina(w_n1313_0[1]),.dinb(w_n1273_0[1]),.dout(n1314),.clk(gclk));
	jxor g1251(.dina(w_n1314_0[1]),.dinb(w_n1271_0[1]),.dout(n1315),.clk(gclk));
	jxor g1252(.dina(w_n1315_0[1]),.dinb(w_n1268_0[1]),.dout(n1316),.clk(gclk));
	jxor g1253(.dina(w_n1316_0[1]),.dinb(w_n1266_0[1]),.dout(n1317),.clk(gclk));
	jxor g1254(.dina(w_n1317_0[1]),.dinb(w_n1263_0[1]),.dout(n1318),.clk(gclk));
	jxor g1255(.dina(w_n1318_0[1]),.dinb(w_n1261_0[1]),.dout(n1319),.clk(gclk));
	jxor g1256(.dina(w_n1319_0[1]),.dinb(w_n1258_0[1]),.dout(n1320),.clk(gclk));
	jxor g1257(.dina(w_n1320_0[1]),.dinb(w_n1256_0[1]),.dout(n1321),.clk(gclk));
	jxor g1258(.dina(w_n1321_0[1]),.dinb(w_n1253_0[1]),.dout(n1322),.clk(gclk));
	jxor g1259(.dina(w_n1322_0[1]),.dinb(w_n1251_0[1]),.dout(n1323),.clk(gclk));
	jnot g1260(.din(n1323),.dout(n1324),.clk(gclk));
	jxor g1261(.dina(w_n1324_0[1]),.dinb(w_n1248_0[1]),.dout(n1325),.clk(gclk));
	jxor g1262(.dina(w_n1325_0[1]),.dinb(w_n1247_0[1]),.dout(n1326),.clk(gclk));
	jnot g1263(.din(w_n1326_0[1]),.dout(n1327),.clk(gclk));
	jxor g1264(.dina(w_dff_B_nYPmOVXp3_0),.dinb(w_n1244_0[1]),.dout(w_dff_A_fM5Zpmhi3_2),.clk(gclk));
	jnot g1265(.din(w_n1325_0[0]),.dout(n1329),.clk(gclk));
	jor g1266(.dina(w_dff_B_yOr46Oam9_0),.dinb(w_n1247_0[0]),.dout(n1330),.clk(gclk));
	jor g1267(.dina(w_n1326_0[0]),.dinb(w_n1244_0[0]),.dout(n1331),.clk(gclk));
	jand g1268(.dina(n1331),.dinb(w_dff_B_W6JW4JY46_1),.dout(n1332),.clk(gclk));
	jnot g1269(.din(w_n1251_0[0]),.dout(n1333),.clk(gclk));
	jnot g1270(.din(w_n1322_0[0]),.dout(n1334),.clk(gclk));
	jor g1271(.dina(w_dff_B_ErSGtDO89_0),.dinb(n1333),.dout(n1335),.clk(gclk));
	jor g1272(.dina(w_n1324_0[0]),.dinb(w_n1248_0[0]),.dout(n1336),.clk(gclk));
	jand g1273(.dina(n1336),.dinb(w_dff_B_FYr4FdfB3_1),.dout(n1337),.clk(gclk));
	jand g1274(.dina(w_G528gat_5[2]),.dinb(w_G86gat_2[1]),.dout(n1338),.clk(gclk));
	jand g1275(.dina(w_n1320_0[0]),.dinb(w_n1256_0[0]),.dout(n1339),.clk(gclk));
	jand g1276(.dina(w_n1321_0[0]),.dinb(w_n1253_0[0]),.dout(n1340),.clk(gclk));
	jor g1277(.dina(n1340),.dinb(w_dff_B_pdJuQq7B8_1),.dout(n1341),.clk(gclk));
	jand g1278(.dina(w_G511gat_5[1]),.dinb(w_G103gat_2[2]),.dout(n1342),.clk(gclk));
	jnot g1279(.din(n1342),.dout(n1343),.clk(gclk));
	jand g1280(.dina(w_n1318_0[0]),.dinb(w_n1261_0[0]),.dout(n1344),.clk(gclk));
	jand g1281(.dina(w_n1319_0[0]),.dinb(w_n1258_0[0]),.dout(n1345),.clk(gclk));
	jor g1282(.dina(n1345),.dinb(w_dff_B_bDocydhb6_1),.dout(n1346),.clk(gclk));
	jand g1283(.dina(w_G494gat_5[0]),.dinb(w_G120gat_3[0]),.dout(n1347),.clk(gclk));
	jnot g1284(.din(n1347),.dout(n1348),.clk(gclk));
	jand g1285(.dina(w_n1316_0[0]),.dinb(w_n1266_0[0]),.dout(n1349),.clk(gclk));
	jand g1286(.dina(w_n1317_0[0]),.dinb(w_n1263_0[0]),.dout(n1350),.clk(gclk));
	jor g1287(.dina(n1350),.dinb(w_dff_B_wy76JoGg3_1),.dout(n1351),.clk(gclk));
	jand g1288(.dina(w_G477gat_4[2]),.dinb(w_G137gat_3[1]),.dout(n1352),.clk(gclk));
	jnot g1289(.din(n1352),.dout(n1353),.clk(gclk));
	jand g1290(.dina(w_n1314_0[0]),.dinb(w_n1271_0[0]),.dout(n1354),.clk(gclk));
	jand g1291(.dina(w_n1315_0[0]),.dinb(w_n1268_0[0]),.dout(n1355),.clk(gclk));
	jor g1292(.dina(n1355),.dinb(w_dff_B_FzF9b9Ge7_1),.dout(n1356),.clk(gclk));
	jand g1293(.dina(w_G460gat_4[1]),.dinb(w_G154gat_3[2]),.dout(n1357),.clk(gclk));
	jnot g1294(.din(n1357),.dout(n1358),.clk(gclk));
	jand g1295(.dina(w_n1312_0[0]),.dinb(w_n1276_0[0]),.dout(n1359),.clk(gclk));
	jand g1296(.dina(w_n1313_0[0]),.dinb(w_n1273_0[0]),.dout(n1360),.clk(gclk));
	jor g1297(.dina(n1360),.dinb(w_dff_B_CE7lS43i5_1),.dout(n1361),.clk(gclk));
	jand g1298(.dina(w_G443gat_4[0]),.dinb(w_G171gat_4[0]),.dout(n1362),.clk(gclk));
	jnot g1299(.din(n1362),.dout(n1363),.clk(gclk));
	jand g1300(.dina(w_n1310_0[0]),.dinb(w_n1281_0[0]),.dout(n1364),.clk(gclk));
	jand g1301(.dina(w_n1311_0[0]),.dinb(w_n1278_0[0]),.dout(n1365),.clk(gclk));
	jor g1302(.dina(n1365),.dinb(w_dff_B_3PqYq3sP3_1),.dout(n1366),.clk(gclk));
	jand g1303(.dina(w_G426gat_3[2]),.dinb(w_G188gat_4[1]),.dout(n1367),.clk(gclk));
	jnot g1304(.din(n1367),.dout(n1368),.clk(gclk));
	jand g1305(.dina(w_n1308_0[0]),.dinb(w_n1286_0[0]),.dout(n1369),.clk(gclk));
	jand g1306(.dina(w_n1309_0[0]),.dinb(w_n1283_0[0]),.dout(n1370),.clk(gclk));
	jor g1307(.dina(n1370),.dinb(w_dff_B_PNvyRkvI3_1),.dout(n1371),.clk(gclk));
	jand g1308(.dina(w_G409gat_3[1]),.dinb(w_G205gat_4[2]),.dout(n1372),.clk(gclk));
	jnot g1309(.din(n1372),.dout(n1373),.clk(gclk));
	jand g1310(.dina(w_n1306_0[0]),.dinb(w_n1291_0[0]),.dout(n1374),.clk(gclk));
	jand g1311(.dina(w_n1307_0[0]),.dinb(w_n1288_0[0]),.dout(n1375),.clk(gclk));
	jor g1312(.dina(n1375),.dinb(w_dff_B_RtdkC2mD4_1),.dout(n1376),.clk(gclk));
	jand g1313(.dina(w_G392gat_3[0]),.dinb(w_G222gat_5[0]),.dout(n1377),.clk(gclk));
	jnot g1314(.din(n1377),.dout(n1378),.clk(gclk));
	jand g1315(.dina(w_n1304_0[0]),.dinb(w_n1296_0[0]),.dout(n1379),.clk(gclk));
	jand g1316(.dina(w_n1305_0[0]),.dinb(w_n1293_0[0]),.dout(n1380),.clk(gclk));
	jor g1317(.dina(n1380),.dinb(w_dff_B_7k9iJ5tT6_1),.dout(n1381),.clk(gclk));
	jand g1318(.dina(w_G375gat_2[2]),.dinb(w_G239gat_5[1]),.dout(n1382),.clk(gclk));
	jand g1319(.dina(w_G358gat_2[1]),.dinb(w_G256gat_5[2]),.dout(n1383),.clk(gclk));
	jor g1320(.dina(w_n1301_0[0]),.dinb(w_n1298_0[0]),.dout(n1384),.clk(gclk));
	jor g1321(.dina(w_n1303_0[0]),.dinb(w_n1297_0[0]),.dout(n1385),.clk(gclk));
	jand g1322(.dina(n1385),.dinb(w_dff_B_2UYJmSWs0_1),.dout(n1386),.clk(gclk));
	jxor g1323(.dina(w_n1386_0[1]),.dinb(w_n1383_0[1]),.dout(n1387),.clk(gclk));
	jnot g1324(.din(n1387),.dout(n1388),.clk(gclk));
	jxor g1325(.dina(w_n1388_0[1]),.dinb(w_n1382_0[1]),.dout(n1389),.clk(gclk));
	jxor g1326(.dina(w_n1389_0[1]),.dinb(w_n1381_0[1]),.dout(n1390),.clk(gclk));
	jxor g1327(.dina(w_n1390_0[1]),.dinb(w_n1378_0[1]),.dout(n1391),.clk(gclk));
	jxor g1328(.dina(w_n1391_0[1]),.dinb(w_n1376_0[1]),.dout(n1392),.clk(gclk));
	jxor g1329(.dina(w_n1392_0[1]),.dinb(w_n1373_0[1]),.dout(n1393),.clk(gclk));
	jxor g1330(.dina(w_n1393_0[1]),.dinb(w_n1371_0[1]),.dout(n1394),.clk(gclk));
	jxor g1331(.dina(w_n1394_0[1]),.dinb(w_n1368_0[1]),.dout(n1395),.clk(gclk));
	jxor g1332(.dina(w_n1395_0[1]),.dinb(w_n1366_0[1]),.dout(n1396),.clk(gclk));
	jxor g1333(.dina(w_n1396_0[1]),.dinb(w_n1363_0[1]),.dout(n1397),.clk(gclk));
	jxor g1334(.dina(w_n1397_0[1]),.dinb(w_n1361_0[1]),.dout(n1398),.clk(gclk));
	jxor g1335(.dina(w_n1398_0[1]),.dinb(w_n1358_0[1]),.dout(n1399),.clk(gclk));
	jxor g1336(.dina(w_n1399_0[1]),.dinb(w_n1356_0[1]),.dout(n1400),.clk(gclk));
	jxor g1337(.dina(w_n1400_0[1]),.dinb(w_n1353_0[1]),.dout(n1401),.clk(gclk));
	jxor g1338(.dina(w_n1401_0[1]),.dinb(w_n1351_0[1]),.dout(n1402),.clk(gclk));
	jxor g1339(.dina(w_n1402_0[1]),.dinb(w_n1348_0[1]),.dout(n1403),.clk(gclk));
	jxor g1340(.dina(w_n1403_0[1]),.dinb(w_n1346_0[1]),.dout(n1404),.clk(gclk));
	jxor g1341(.dina(w_n1404_0[1]),.dinb(w_n1343_0[1]),.dout(n1405),.clk(gclk));
	jxor g1342(.dina(w_n1405_0[1]),.dinb(w_n1341_0[1]),.dout(n1406),.clk(gclk));
	jnot g1343(.din(n1406),.dout(n1407),.clk(gclk));
	jxor g1344(.dina(w_n1407_0[1]),.dinb(w_n1338_0[1]),.dout(n1408),.clk(gclk));
	jnot g1345(.din(n1408),.dout(n1409),.clk(gclk));
	jxor g1346(.dina(w_n1409_0[1]),.dinb(w_n1337_0[1]),.dout(n1410),.clk(gclk));
	jxor g1347(.dina(w_n1410_0[1]),.dinb(w_n1332_0[1]),.dout(w_dff_A_ErYJJyU15_2),.clk(gclk));
	jor g1348(.dina(w_n1409_0[0]),.dinb(w_n1337_0[0]),.dout(n1412),.clk(gclk));
	jnot g1349(.din(w_n1410_0[0]),.dout(n1413),.clk(gclk));
	jor g1350(.dina(w_dff_B_w6qGUp2q7_0),.dinb(w_n1332_0[0]),.dout(n1414),.clk(gclk));
	jand g1351(.dina(n1414),.dinb(w_dff_B_0wQXfKuk2_1),.dout(n1415),.clk(gclk));
	jnot g1352(.din(w_n1341_0[0]),.dout(n1416),.clk(gclk));
	jnot g1353(.din(w_n1405_0[0]),.dout(n1417),.clk(gclk));
	jor g1354(.dina(n1417),.dinb(n1416),.dout(n1418),.clk(gclk));
	jor g1355(.dina(w_n1407_0[0]),.dinb(w_n1338_0[0]),.dout(n1419),.clk(gclk));
	jand g1356(.dina(n1419),.dinb(w_dff_B_LlyAvuTl5_1),.dout(n1420),.clk(gclk));
	jand g1357(.dina(w_G528gat_5[1]),.dinb(w_G103gat_2[1]),.dout(n1421),.clk(gclk));
	jand g1358(.dina(w_n1403_0[0]),.dinb(w_n1346_0[0]),.dout(n1422),.clk(gclk));
	jand g1359(.dina(w_n1404_0[0]),.dinb(w_n1343_0[0]),.dout(n1423),.clk(gclk));
	jor g1360(.dina(n1423),.dinb(w_dff_B_0sLmQqVT3_1),.dout(n1424),.clk(gclk));
	jand g1361(.dina(w_G511gat_5[0]),.dinb(w_G120gat_2[2]),.dout(n1425),.clk(gclk));
	jnot g1362(.din(n1425),.dout(n1426),.clk(gclk));
	jand g1363(.dina(w_n1401_0[0]),.dinb(w_n1351_0[0]),.dout(n1427),.clk(gclk));
	jand g1364(.dina(w_n1402_0[0]),.dinb(w_n1348_0[0]),.dout(n1428),.clk(gclk));
	jor g1365(.dina(n1428),.dinb(w_dff_B_ZSPAhZlk1_1),.dout(n1429),.clk(gclk));
	jand g1366(.dina(w_G494gat_4[2]),.dinb(w_G137gat_3[0]),.dout(n1430),.clk(gclk));
	jnot g1367(.din(n1430),.dout(n1431),.clk(gclk));
	jand g1368(.dina(w_n1399_0[0]),.dinb(w_n1356_0[0]),.dout(n1432),.clk(gclk));
	jand g1369(.dina(w_n1400_0[0]),.dinb(w_n1353_0[0]),.dout(n1433),.clk(gclk));
	jor g1370(.dina(n1433),.dinb(w_dff_B_BlR6EJkB2_1),.dout(n1434),.clk(gclk));
	jand g1371(.dina(w_G477gat_4[1]),.dinb(w_G154gat_3[1]),.dout(n1435),.clk(gclk));
	jnot g1372(.din(n1435),.dout(n1436),.clk(gclk));
	jand g1373(.dina(w_n1397_0[0]),.dinb(w_n1361_0[0]),.dout(n1437),.clk(gclk));
	jand g1374(.dina(w_n1398_0[0]),.dinb(w_n1358_0[0]),.dout(n1438),.clk(gclk));
	jor g1375(.dina(n1438),.dinb(w_dff_B_0zbkiSiI3_1),.dout(n1439),.clk(gclk));
	jand g1376(.dina(w_G460gat_4[0]),.dinb(w_G171gat_3[2]),.dout(n1440),.clk(gclk));
	jnot g1377(.din(n1440),.dout(n1441),.clk(gclk));
	jand g1378(.dina(w_n1395_0[0]),.dinb(w_n1366_0[0]),.dout(n1442),.clk(gclk));
	jand g1379(.dina(w_n1396_0[0]),.dinb(w_n1363_0[0]),.dout(n1443),.clk(gclk));
	jor g1380(.dina(n1443),.dinb(w_dff_B_ZYR8bUcq9_1),.dout(n1444),.clk(gclk));
	jand g1381(.dina(w_G443gat_3[2]),.dinb(w_G188gat_4[0]),.dout(n1445),.clk(gclk));
	jnot g1382(.din(n1445),.dout(n1446),.clk(gclk));
	jand g1383(.dina(w_n1393_0[0]),.dinb(w_n1371_0[0]),.dout(n1447),.clk(gclk));
	jand g1384(.dina(w_n1394_0[0]),.dinb(w_n1368_0[0]),.dout(n1448),.clk(gclk));
	jor g1385(.dina(n1448),.dinb(w_dff_B_JqiJPZgx9_1),.dout(n1449),.clk(gclk));
	jand g1386(.dina(w_G426gat_3[1]),.dinb(w_G205gat_4[1]),.dout(n1450),.clk(gclk));
	jnot g1387(.din(n1450),.dout(n1451),.clk(gclk));
	jand g1388(.dina(w_n1391_0[0]),.dinb(w_n1376_0[0]),.dout(n1452),.clk(gclk));
	jand g1389(.dina(w_n1392_0[0]),.dinb(w_n1373_0[0]),.dout(n1453),.clk(gclk));
	jor g1390(.dina(n1453),.dinb(w_dff_B_2eWKUzzW9_1),.dout(n1454),.clk(gclk));
	jand g1391(.dina(w_G409gat_3[0]),.dinb(w_G222gat_4[2]),.dout(n1455),.clk(gclk));
	jnot g1392(.din(n1455),.dout(n1456),.clk(gclk));
	jand g1393(.dina(w_n1389_0[0]),.dinb(w_n1381_0[0]),.dout(n1457),.clk(gclk));
	jand g1394(.dina(w_n1390_0[0]),.dinb(w_n1378_0[0]),.dout(n1458),.clk(gclk));
	jor g1395(.dina(n1458),.dinb(w_dff_B_MiHFayT22_1),.dout(n1459),.clk(gclk));
	jand g1396(.dina(w_G392gat_2[2]),.dinb(w_G239gat_5[0]),.dout(n1460),.clk(gclk));
	jand g1397(.dina(w_G375gat_2[1]),.dinb(w_G256gat_5[1]),.dout(n1461),.clk(gclk));
	jor g1398(.dina(w_n1386_0[0]),.dinb(w_n1383_0[0]),.dout(n1462),.clk(gclk));
	jor g1399(.dina(w_n1388_0[0]),.dinb(w_n1382_0[0]),.dout(n1463),.clk(gclk));
	jand g1400(.dina(n1463),.dinb(w_dff_B_meQsglwa0_1),.dout(n1464),.clk(gclk));
	jxor g1401(.dina(w_n1464_0[1]),.dinb(w_n1461_0[1]),.dout(n1465),.clk(gclk));
	jnot g1402(.din(n1465),.dout(n1466),.clk(gclk));
	jxor g1403(.dina(w_n1466_0[1]),.dinb(w_n1460_0[1]),.dout(n1467),.clk(gclk));
	jxor g1404(.dina(w_n1467_0[1]),.dinb(w_n1459_0[1]),.dout(n1468),.clk(gclk));
	jxor g1405(.dina(w_n1468_0[1]),.dinb(w_n1456_0[1]),.dout(n1469),.clk(gclk));
	jxor g1406(.dina(w_n1469_0[1]),.dinb(w_n1454_0[1]),.dout(n1470),.clk(gclk));
	jxor g1407(.dina(w_n1470_0[1]),.dinb(w_n1451_0[1]),.dout(n1471),.clk(gclk));
	jxor g1408(.dina(w_n1471_0[1]),.dinb(w_n1449_0[1]),.dout(n1472),.clk(gclk));
	jxor g1409(.dina(w_n1472_0[1]),.dinb(w_n1446_0[1]),.dout(n1473),.clk(gclk));
	jxor g1410(.dina(w_n1473_0[1]),.dinb(w_n1444_0[1]),.dout(n1474),.clk(gclk));
	jxor g1411(.dina(w_n1474_0[1]),.dinb(w_n1441_0[1]),.dout(n1475),.clk(gclk));
	jxor g1412(.dina(w_n1475_0[1]),.dinb(w_n1439_0[1]),.dout(n1476),.clk(gclk));
	jxor g1413(.dina(w_n1476_0[1]),.dinb(w_n1436_0[1]),.dout(n1477),.clk(gclk));
	jxor g1414(.dina(w_n1477_0[1]),.dinb(w_n1434_0[1]),.dout(n1478),.clk(gclk));
	jxor g1415(.dina(w_n1478_0[1]),.dinb(w_n1431_0[1]),.dout(n1479),.clk(gclk));
	jxor g1416(.dina(w_n1479_0[1]),.dinb(w_n1429_0[1]),.dout(n1480),.clk(gclk));
	jxor g1417(.dina(w_n1480_0[1]),.dinb(w_n1426_0[1]),.dout(n1481),.clk(gclk));
	jxor g1418(.dina(w_n1481_0[1]),.dinb(w_n1424_0[1]),.dout(n1482),.clk(gclk));
	jnot g1419(.din(n1482),.dout(n1483),.clk(gclk));
	jxor g1420(.dina(w_n1483_0[1]),.dinb(w_n1421_0[1]),.dout(n1484),.clk(gclk));
	jnot g1421(.din(n1484),.dout(n1485),.clk(gclk));
	jxor g1422(.dina(w_n1485_0[1]),.dinb(w_n1420_0[1]),.dout(n1486),.clk(gclk));
	jxor g1423(.dina(w_n1486_0[1]),.dinb(w_n1415_0[1]),.dout(w_dff_A_AzVrOdhu4_2),.clk(gclk));
	jor g1424(.dina(w_n1485_0[0]),.dinb(w_n1420_0[0]),.dout(n1488),.clk(gclk));
	jnot g1425(.din(w_n1486_0[0]),.dout(n1489),.clk(gclk));
	jor g1426(.dina(w_dff_B_cotjRpX83_0),.dinb(w_n1415_0[0]),.dout(n1490),.clk(gclk));
	jand g1427(.dina(n1490),.dinb(w_dff_B_KasjwAkM9_1),.dout(n1491),.clk(gclk));
	jnot g1428(.din(w_n1424_0[0]),.dout(n1492),.clk(gclk));
	jnot g1429(.din(w_n1481_0[0]),.dout(n1493),.clk(gclk));
	jor g1430(.dina(n1493),.dinb(n1492),.dout(n1494),.clk(gclk));
	jor g1431(.dina(w_n1483_0[0]),.dinb(w_n1421_0[0]),.dout(n1495),.clk(gclk));
	jand g1432(.dina(n1495),.dinb(w_dff_B_lyPa9dUU4_1),.dout(n1496),.clk(gclk));
	jand g1433(.dina(w_G528gat_5[0]),.dinb(w_G120gat_2[1]),.dout(n1497),.clk(gclk));
	jand g1434(.dina(w_n1479_0[0]),.dinb(w_n1429_0[0]),.dout(n1498),.clk(gclk));
	jand g1435(.dina(w_n1480_0[0]),.dinb(w_n1426_0[0]),.dout(n1499),.clk(gclk));
	jor g1436(.dina(n1499),.dinb(w_dff_B_e2bwT7h06_1),.dout(n1500),.clk(gclk));
	jand g1437(.dina(w_G511gat_4[2]),.dinb(w_G137gat_2[2]),.dout(n1501),.clk(gclk));
	jnot g1438(.din(n1501),.dout(n1502),.clk(gclk));
	jand g1439(.dina(w_n1477_0[0]),.dinb(w_n1434_0[0]),.dout(n1503),.clk(gclk));
	jand g1440(.dina(w_n1478_0[0]),.dinb(w_n1431_0[0]),.dout(n1504),.clk(gclk));
	jor g1441(.dina(n1504),.dinb(w_dff_B_aRK956Io7_1),.dout(n1505),.clk(gclk));
	jand g1442(.dina(w_G494gat_4[1]),.dinb(w_G154gat_3[0]),.dout(n1506),.clk(gclk));
	jnot g1443(.din(n1506),.dout(n1507),.clk(gclk));
	jand g1444(.dina(w_n1475_0[0]),.dinb(w_n1439_0[0]),.dout(n1508),.clk(gclk));
	jand g1445(.dina(w_n1476_0[0]),.dinb(w_n1436_0[0]),.dout(n1509),.clk(gclk));
	jor g1446(.dina(n1509),.dinb(w_dff_B_6NaOW2oA3_1),.dout(n1510),.clk(gclk));
	jand g1447(.dina(w_G477gat_4[0]),.dinb(w_G171gat_3[1]),.dout(n1511),.clk(gclk));
	jnot g1448(.din(n1511),.dout(n1512),.clk(gclk));
	jand g1449(.dina(w_n1473_0[0]),.dinb(w_n1444_0[0]),.dout(n1513),.clk(gclk));
	jand g1450(.dina(w_n1474_0[0]),.dinb(w_n1441_0[0]),.dout(n1514),.clk(gclk));
	jor g1451(.dina(n1514),.dinb(w_dff_B_yhcxjPXC0_1),.dout(n1515),.clk(gclk));
	jand g1452(.dina(w_G460gat_3[2]),.dinb(w_G188gat_3[2]),.dout(n1516),.clk(gclk));
	jnot g1453(.din(n1516),.dout(n1517),.clk(gclk));
	jand g1454(.dina(w_n1471_0[0]),.dinb(w_n1449_0[0]),.dout(n1518),.clk(gclk));
	jand g1455(.dina(w_n1472_0[0]),.dinb(w_n1446_0[0]),.dout(n1519),.clk(gclk));
	jor g1456(.dina(n1519),.dinb(w_dff_B_tB5h44mQ6_1),.dout(n1520),.clk(gclk));
	jand g1457(.dina(w_G443gat_3[1]),.dinb(w_G205gat_4[0]),.dout(n1521),.clk(gclk));
	jnot g1458(.din(n1521),.dout(n1522),.clk(gclk));
	jand g1459(.dina(w_n1469_0[0]),.dinb(w_n1454_0[0]),.dout(n1523),.clk(gclk));
	jand g1460(.dina(w_n1470_0[0]),.dinb(w_n1451_0[0]),.dout(n1524),.clk(gclk));
	jor g1461(.dina(n1524),.dinb(w_dff_B_CPSDcxeo0_1),.dout(n1525),.clk(gclk));
	jand g1462(.dina(w_G426gat_3[0]),.dinb(w_G222gat_4[1]),.dout(n1526),.clk(gclk));
	jnot g1463(.din(n1526),.dout(n1527),.clk(gclk));
	jand g1464(.dina(w_n1467_0[0]),.dinb(w_n1459_0[0]),.dout(n1528),.clk(gclk));
	jand g1465(.dina(w_n1468_0[0]),.dinb(w_n1456_0[0]),.dout(n1529),.clk(gclk));
	jor g1466(.dina(n1529),.dinb(w_dff_B_eVn4YkX40_1),.dout(n1530),.clk(gclk));
	jand g1467(.dina(w_G409gat_2[2]),.dinb(w_G239gat_4[2]),.dout(n1531),.clk(gclk));
	jand g1468(.dina(w_G392gat_2[1]),.dinb(w_G256gat_5[0]),.dout(n1532),.clk(gclk));
	jor g1469(.dina(w_n1464_0[0]),.dinb(w_n1461_0[0]),.dout(n1533),.clk(gclk));
	jor g1470(.dina(w_n1466_0[0]),.dinb(w_n1460_0[0]),.dout(n1534),.clk(gclk));
	jand g1471(.dina(n1534),.dinb(w_dff_B_vQjzTvuR7_1),.dout(n1535),.clk(gclk));
	jxor g1472(.dina(w_n1535_0[1]),.dinb(w_n1532_0[1]),.dout(n1536),.clk(gclk));
	jnot g1473(.din(n1536),.dout(n1537),.clk(gclk));
	jxor g1474(.dina(w_n1537_0[1]),.dinb(w_n1531_0[1]),.dout(n1538),.clk(gclk));
	jxor g1475(.dina(w_n1538_0[1]),.dinb(w_n1530_0[1]),.dout(n1539),.clk(gclk));
	jxor g1476(.dina(w_n1539_0[1]),.dinb(w_n1527_0[1]),.dout(n1540),.clk(gclk));
	jxor g1477(.dina(w_n1540_0[1]),.dinb(w_n1525_0[1]),.dout(n1541),.clk(gclk));
	jxor g1478(.dina(w_n1541_0[1]),.dinb(w_n1522_0[1]),.dout(n1542),.clk(gclk));
	jxor g1479(.dina(w_n1542_0[1]),.dinb(w_n1520_0[1]),.dout(n1543),.clk(gclk));
	jxor g1480(.dina(w_n1543_0[1]),.dinb(w_n1517_0[1]),.dout(n1544),.clk(gclk));
	jxor g1481(.dina(w_n1544_0[1]),.dinb(w_n1515_0[1]),.dout(n1545),.clk(gclk));
	jxor g1482(.dina(w_n1545_0[1]),.dinb(w_n1512_0[1]),.dout(n1546),.clk(gclk));
	jxor g1483(.dina(w_n1546_0[1]),.dinb(w_n1510_0[1]),.dout(n1547),.clk(gclk));
	jxor g1484(.dina(w_n1547_0[1]),.dinb(w_n1507_0[1]),.dout(n1548),.clk(gclk));
	jxor g1485(.dina(w_n1548_0[1]),.dinb(w_n1505_0[1]),.dout(n1549),.clk(gclk));
	jxor g1486(.dina(w_n1549_0[1]),.dinb(w_n1502_0[1]),.dout(n1550),.clk(gclk));
	jxor g1487(.dina(w_n1550_0[1]),.dinb(w_n1500_0[1]),.dout(n1551),.clk(gclk));
	jnot g1488(.din(n1551),.dout(n1552),.clk(gclk));
	jxor g1489(.dina(w_n1552_0[1]),.dinb(w_n1497_0[1]),.dout(n1553),.clk(gclk));
	jnot g1490(.din(n1553),.dout(n1554),.clk(gclk));
	jxor g1491(.dina(w_n1554_0[1]),.dinb(w_n1496_0[1]),.dout(n1555),.clk(gclk));
	jxor g1492(.dina(w_n1555_0[1]),.dinb(w_n1491_0[1]),.dout(w_dff_A_bjPY08b41_2),.clk(gclk));
	jor g1493(.dina(w_n1554_0[0]),.dinb(w_n1496_0[0]),.dout(n1557),.clk(gclk));
	jnot g1494(.din(w_n1555_0[0]),.dout(n1558),.clk(gclk));
	jor g1495(.dina(w_dff_B_m0hmfefD1_0),.dinb(w_n1491_0[0]),.dout(n1559),.clk(gclk));
	jand g1496(.dina(n1559),.dinb(w_dff_B_EAv8BngY7_1),.dout(n1560),.clk(gclk));
	jnot g1497(.din(w_n1500_0[0]),.dout(n1561),.clk(gclk));
	jnot g1498(.din(w_n1550_0[0]),.dout(n1562),.clk(gclk));
	jor g1499(.dina(w_dff_B_s9pv34mm5_0),.dinb(n1561),.dout(n1563),.clk(gclk));
	jor g1500(.dina(w_n1552_0[0]),.dinb(w_n1497_0[0]),.dout(n1564),.clk(gclk));
	jand g1501(.dina(n1564),.dinb(w_dff_B_a7Ek4TkY8_1),.dout(n1565),.clk(gclk));
	jand g1502(.dina(w_G528gat_4[2]),.dinb(w_G137gat_2[1]),.dout(n1566),.clk(gclk));
	jand g1503(.dina(w_n1548_0[0]),.dinb(w_n1505_0[0]),.dout(n1567),.clk(gclk));
	jand g1504(.dina(w_n1549_0[0]),.dinb(w_n1502_0[0]),.dout(n1568),.clk(gclk));
	jor g1505(.dina(n1568),.dinb(w_dff_B_CdmtuydS5_1),.dout(n1569),.clk(gclk));
	jand g1506(.dina(w_G511gat_4[1]),.dinb(w_G154gat_2[2]),.dout(n1570),.clk(gclk));
	jnot g1507(.din(n1570),.dout(n1571),.clk(gclk));
	jand g1508(.dina(w_n1546_0[0]),.dinb(w_n1510_0[0]),.dout(n1572),.clk(gclk));
	jand g1509(.dina(w_n1547_0[0]),.dinb(w_n1507_0[0]),.dout(n1573),.clk(gclk));
	jor g1510(.dina(n1573),.dinb(w_dff_B_tX56hz7o5_1),.dout(n1574),.clk(gclk));
	jand g1511(.dina(w_G494gat_4[0]),.dinb(w_G171gat_3[0]),.dout(n1575),.clk(gclk));
	jnot g1512(.din(n1575),.dout(n1576),.clk(gclk));
	jand g1513(.dina(w_n1544_0[0]),.dinb(w_n1515_0[0]),.dout(n1577),.clk(gclk));
	jand g1514(.dina(w_n1545_0[0]),.dinb(w_n1512_0[0]),.dout(n1578),.clk(gclk));
	jor g1515(.dina(n1578),.dinb(w_dff_B_T6U1i5sD6_1),.dout(n1579),.clk(gclk));
	jand g1516(.dina(w_G477gat_3[2]),.dinb(w_G188gat_3[1]),.dout(n1580),.clk(gclk));
	jnot g1517(.din(n1580),.dout(n1581),.clk(gclk));
	jand g1518(.dina(w_n1542_0[0]),.dinb(w_n1520_0[0]),.dout(n1582),.clk(gclk));
	jand g1519(.dina(w_n1543_0[0]),.dinb(w_n1517_0[0]),.dout(n1583),.clk(gclk));
	jor g1520(.dina(n1583),.dinb(w_dff_B_Z7ZDwvJ80_1),.dout(n1584),.clk(gclk));
	jand g1521(.dina(w_G460gat_3[1]),.dinb(w_G205gat_3[2]),.dout(n1585),.clk(gclk));
	jnot g1522(.din(n1585),.dout(n1586),.clk(gclk));
	jand g1523(.dina(w_n1540_0[0]),.dinb(w_n1525_0[0]),.dout(n1587),.clk(gclk));
	jand g1524(.dina(w_n1541_0[0]),.dinb(w_n1522_0[0]),.dout(n1588),.clk(gclk));
	jor g1525(.dina(n1588),.dinb(w_dff_B_AjoZInzR4_1),.dout(n1589),.clk(gclk));
	jand g1526(.dina(w_G443gat_3[0]),.dinb(w_G222gat_4[0]),.dout(n1590),.clk(gclk));
	jnot g1527(.din(n1590),.dout(n1591),.clk(gclk));
	jand g1528(.dina(w_n1538_0[0]),.dinb(w_n1530_0[0]),.dout(n1592),.clk(gclk));
	jand g1529(.dina(w_n1539_0[0]),.dinb(w_n1527_0[0]),.dout(n1593),.clk(gclk));
	jor g1530(.dina(n1593),.dinb(w_dff_B_5Ib0KJ6z6_1),.dout(n1594),.clk(gclk));
	jand g1531(.dina(w_G426gat_2[2]),.dinb(w_G239gat_4[1]),.dout(n1595),.clk(gclk));
	jand g1532(.dina(w_G409gat_2[1]),.dinb(w_G256gat_4[2]),.dout(n1596),.clk(gclk));
	jor g1533(.dina(w_n1535_0[0]),.dinb(w_n1532_0[0]),.dout(n1597),.clk(gclk));
	jor g1534(.dina(w_n1537_0[0]),.dinb(w_n1531_0[0]),.dout(n1598),.clk(gclk));
	jand g1535(.dina(n1598),.dinb(w_dff_B_jpgEFxr40_1),.dout(n1599),.clk(gclk));
	jxor g1536(.dina(w_n1599_0[1]),.dinb(w_n1596_0[1]),.dout(n1600),.clk(gclk));
	jnot g1537(.din(n1600),.dout(n1601),.clk(gclk));
	jxor g1538(.dina(w_n1601_0[1]),.dinb(w_n1595_0[1]),.dout(n1602),.clk(gclk));
	jxor g1539(.dina(w_n1602_0[1]),.dinb(w_n1594_0[1]),.dout(n1603),.clk(gclk));
	jxor g1540(.dina(w_n1603_0[1]),.dinb(w_n1591_0[1]),.dout(n1604),.clk(gclk));
	jxor g1541(.dina(w_n1604_0[1]),.dinb(w_n1589_0[1]),.dout(n1605),.clk(gclk));
	jxor g1542(.dina(w_n1605_0[1]),.dinb(w_n1586_0[1]),.dout(n1606),.clk(gclk));
	jxor g1543(.dina(w_n1606_0[1]),.dinb(w_n1584_0[1]),.dout(n1607),.clk(gclk));
	jxor g1544(.dina(w_n1607_0[1]),.dinb(w_n1581_0[1]),.dout(n1608),.clk(gclk));
	jxor g1545(.dina(w_n1608_0[1]),.dinb(w_n1579_0[1]),.dout(n1609),.clk(gclk));
	jxor g1546(.dina(w_n1609_0[1]),.dinb(w_n1576_0[1]),.dout(n1610),.clk(gclk));
	jxor g1547(.dina(w_n1610_0[1]),.dinb(w_n1574_0[1]),.dout(n1611),.clk(gclk));
	jxor g1548(.dina(w_n1611_0[1]),.dinb(w_n1571_0[1]),.dout(n1612),.clk(gclk));
	jxor g1549(.dina(w_n1612_0[1]),.dinb(w_n1569_0[1]),.dout(n1613),.clk(gclk));
	jnot g1550(.din(n1613),.dout(n1614),.clk(gclk));
	jxor g1551(.dina(w_n1614_0[1]),.dinb(w_n1566_0[1]),.dout(n1615),.clk(gclk));
	jnot g1552(.din(n1615),.dout(n1616),.clk(gclk));
	jxor g1553(.dina(w_n1616_0[1]),.dinb(w_n1565_0[1]),.dout(n1617),.clk(gclk));
	jxor g1554(.dina(w_n1617_0[1]),.dinb(w_n1560_0[1]),.dout(w_dff_A_DmqhRz3o5_2),.clk(gclk));
	jor g1555(.dina(w_n1616_0[0]),.dinb(w_n1565_0[0]),.dout(n1619),.clk(gclk));
	jnot g1556(.din(w_n1617_0[0]),.dout(n1620),.clk(gclk));
	jor g1557(.dina(w_dff_B_6YQoVxFh5_0),.dinb(w_n1560_0[0]),.dout(n1621),.clk(gclk));
	jand g1558(.dina(n1621),.dinb(w_dff_B_ARhsUsw33_1),.dout(n1622),.clk(gclk));
	jnot g1559(.din(w_n1569_0[0]),.dout(n1623),.clk(gclk));
	jnot g1560(.din(w_n1612_0[0]),.dout(n1624),.clk(gclk));
	jor g1561(.dina(n1624),.dinb(n1623),.dout(n1625),.clk(gclk));
	jor g1562(.dina(w_n1614_0[0]),.dinb(w_n1566_0[0]),.dout(n1626),.clk(gclk));
	jand g1563(.dina(n1626),.dinb(w_dff_B_EkZtMXUx2_1),.dout(n1627),.clk(gclk));
	jand g1564(.dina(w_G528gat_4[1]),.dinb(w_G154gat_2[1]),.dout(n1628),.clk(gclk));
	jand g1565(.dina(w_n1610_0[0]),.dinb(w_n1574_0[0]),.dout(n1629),.clk(gclk));
	jand g1566(.dina(w_n1611_0[0]),.dinb(w_n1571_0[0]),.dout(n1630),.clk(gclk));
	jor g1567(.dina(n1630),.dinb(w_dff_B_8piwo4me2_1),.dout(n1631),.clk(gclk));
	jand g1568(.dina(w_G511gat_4[0]),.dinb(w_G171gat_2[2]),.dout(n1632),.clk(gclk));
	jnot g1569(.din(n1632),.dout(n1633),.clk(gclk));
	jand g1570(.dina(w_n1608_0[0]),.dinb(w_n1579_0[0]),.dout(n1634),.clk(gclk));
	jand g1571(.dina(w_n1609_0[0]),.dinb(w_n1576_0[0]),.dout(n1635),.clk(gclk));
	jor g1572(.dina(n1635),.dinb(w_dff_B_QKibgKDa8_1),.dout(n1636),.clk(gclk));
	jand g1573(.dina(w_G494gat_3[2]),.dinb(w_G188gat_3[0]),.dout(n1637),.clk(gclk));
	jnot g1574(.din(n1637),.dout(n1638),.clk(gclk));
	jand g1575(.dina(w_n1606_0[0]),.dinb(w_n1584_0[0]),.dout(n1639),.clk(gclk));
	jand g1576(.dina(w_n1607_0[0]),.dinb(w_n1581_0[0]),.dout(n1640),.clk(gclk));
	jor g1577(.dina(n1640),.dinb(w_dff_B_A4pjQGCK7_1),.dout(n1641),.clk(gclk));
	jand g1578(.dina(w_G477gat_3[1]),.dinb(w_G205gat_3[1]),.dout(n1642),.clk(gclk));
	jnot g1579(.din(n1642),.dout(n1643),.clk(gclk));
	jand g1580(.dina(w_n1604_0[0]),.dinb(w_n1589_0[0]),.dout(n1644),.clk(gclk));
	jand g1581(.dina(w_n1605_0[0]),.dinb(w_n1586_0[0]),.dout(n1645),.clk(gclk));
	jor g1582(.dina(n1645),.dinb(w_dff_B_8uuf1NPF9_1),.dout(n1646),.clk(gclk));
	jand g1583(.dina(w_G460gat_3[0]),.dinb(w_G222gat_3[2]),.dout(n1647),.clk(gclk));
	jnot g1584(.din(n1647),.dout(n1648),.clk(gclk));
	jand g1585(.dina(w_n1602_0[0]),.dinb(w_n1594_0[0]),.dout(n1649),.clk(gclk));
	jand g1586(.dina(w_n1603_0[0]),.dinb(w_n1591_0[0]),.dout(n1650),.clk(gclk));
	jor g1587(.dina(n1650),.dinb(w_dff_B_ZKC0WEWM3_1),.dout(n1651),.clk(gclk));
	jand g1588(.dina(w_G443gat_2[2]),.dinb(w_G239gat_4[0]),.dout(n1652),.clk(gclk));
	jand g1589(.dina(w_G426gat_2[1]),.dinb(w_G256gat_4[1]),.dout(n1653),.clk(gclk));
	jor g1590(.dina(w_n1599_0[0]),.dinb(w_n1596_0[0]),.dout(n1654),.clk(gclk));
	jor g1591(.dina(w_n1601_0[0]),.dinb(w_n1595_0[0]),.dout(n1655),.clk(gclk));
	jand g1592(.dina(n1655),.dinb(w_dff_B_nlXGNjIF6_1),.dout(n1656),.clk(gclk));
	jxor g1593(.dina(w_n1656_0[1]),.dinb(w_n1653_0[1]),.dout(n1657),.clk(gclk));
	jnot g1594(.din(n1657),.dout(n1658),.clk(gclk));
	jxor g1595(.dina(w_n1658_0[1]),.dinb(w_n1652_0[1]),.dout(n1659),.clk(gclk));
	jxor g1596(.dina(w_n1659_0[1]),.dinb(w_n1651_0[1]),.dout(n1660),.clk(gclk));
	jxor g1597(.dina(w_n1660_0[1]),.dinb(w_n1648_0[1]),.dout(n1661),.clk(gclk));
	jxor g1598(.dina(w_n1661_0[1]),.dinb(w_n1646_0[1]),.dout(n1662),.clk(gclk));
	jxor g1599(.dina(w_n1662_0[1]),.dinb(w_n1643_0[1]),.dout(n1663),.clk(gclk));
	jxor g1600(.dina(w_n1663_0[1]),.dinb(w_n1641_0[1]),.dout(n1664),.clk(gclk));
	jxor g1601(.dina(w_n1664_0[1]),.dinb(w_n1638_0[1]),.dout(n1665),.clk(gclk));
	jxor g1602(.dina(w_n1665_0[1]),.dinb(w_n1636_0[1]),.dout(n1666),.clk(gclk));
	jxor g1603(.dina(w_n1666_0[1]),.dinb(w_n1633_0[1]),.dout(n1667),.clk(gclk));
	jxor g1604(.dina(w_n1667_0[1]),.dinb(w_n1631_0[1]),.dout(n1668),.clk(gclk));
	jnot g1605(.din(n1668),.dout(n1669),.clk(gclk));
	jxor g1606(.dina(w_n1669_0[1]),.dinb(w_n1628_0[1]),.dout(n1670),.clk(gclk));
	jnot g1607(.din(n1670),.dout(n1671),.clk(gclk));
	jxor g1608(.dina(w_n1671_0[1]),.dinb(w_n1627_0[1]),.dout(n1672),.clk(gclk));
	jxor g1609(.dina(w_n1672_0[1]),.dinb(w_n1622_0[1]),.dout(w_dff_A_Gu5QXbuJ7_2),.clk(gclk));
	jor g1610(.dina(w_n1671_0[0]),.dinb(w_n1627_0[0]),.dout(n1674),.clk(gclk));
	jnot g1611(.din(w_n1672_0[0]),.dout(n1675),.clk(gclk));
	jor g1612(.dina(w_dff_B_Tze7IZDs2_0),.dinb(w_n1622_0[0]),.dout(n1676),.clk(gclk));
	jand g1613(.dina(n1676),.dinb(w_dff_B_mtlvViN33_1),.dout(n1677),.clk(gclk));
	jnot g1614(.din(w_n1631_0[0]),.dout(n1678),.clk(gclk));
	jnot g1615(.din(w_n1667_0[0]),.dout(n1679),.clk(gclk));
	jor g1616(.dina(n1679),.dinb(w_dff_B_1uK7f00G7_1),.dout(n1680),.clk(gclk));
	jor g1617(.dina(w_n1669_0[0]),.dinb(w_n1628_0[0]),.dout(n1681),.clk(gclk));
	jand g1618(.dina(n1681),.dinb(w_dff_B_lVy3GB6O5_1),.dout(n1682),.clk(gclk));
	jand g1619(.dina(w_G528gat_4[0]),.dinb(w_G171gat_2[1]),.dout(n1683),.clk(gclk));
	jnot g1620(.din(n1683),.dout(n1684),.clk(gclk));
	jand g1621(.dina(w_n1665_0[0]),.dinb(w_n1636_0[0]),.dout(n1685),.clk(gclk));
	jand g1622(.dina(w_n1666_0[0]),.dinb(w_n1633_0[0]),.dout(n1686),.clk(gclk));
	jor g1623(.dina(n1686),.dinb(w_dff_B_6E1WzGAH5_1),.dout(n1687),.clk(gclk));
	jand g1624(.dina(w_G511gat_3[2]),.dinb(w_G188gat_2[2]),.dout(n1688),.clk(gclk));
	jnot g1625(.din(n1688),.dout(n1689),.clk(gclk));
	jand g1626(.dina(w_n1663_0[0]),.dinb(w_n1641_0[0]),.dout(n1690),.clk(gclk));
	jand g1627(.dina(w_n1664_0[0]),.dinb(w_n1638_0[0]),.dout(n1691),.clk(gclk));
	jor g1628(.dina(n1691),.dinb(w_dff_B_1mu5OWs52_1),.dout(n1692),.clk(gclk));
	jand g1629(.dina(w_G494gat_3[1]),.dinb(w_G205gat_3[0]),.dout(n1693),.clk(gclk));
	jnot g1630(.din(n1693),.dout(n1694),.clk(gclk));
	jand g1631(.dina(w_n1661_0[0]),.dinb(w_n1646_0[0]),.dout(n1695),.clk(gclk));
	jand g1632(.dina(w_n1662_0[0]),.dinb(w_n1643_0[0]),.dout(n1696),.clk(gclk));
	jor g1633(.dina(n1696),.dinb(w_dff_B_bCY77S658_1),.dout(n1697),.clk(gclk));
	jand g1634(.dina(w_G477gat_3[0]),.dinb(w_G222gat_3[1]),.dout(n1698),.clk(gclk));
	jnot g1635(.din(n1698),.dout(n1699),.clk(gclk));
	jand g1636(.dina(w_n1659_0[0]),.dinb(w_n1651_0[0]),.dout(n1700),.clk(gclk));
	jand g1637(.dina(w_n1660_0[0]),.dinb(w_n1648_0[0]),.dout(n1701),.clk(gclk));
	jor g1638(.dina(n1701),.dinb(w_dff_B_9ydfEmg55_1),.dout(n1702),.clk(gclk));
	jand g1639(.dina(w_G460gat_2[2]),.dinb(w_G239gat_3[2]),.dout(n1703),.clk(gclk));
	jand g1640(.dina(w_G443gat_2[1]),.dinb(w_G256gat_4[0]),.dout(n1704),.clk(gclk));
	jor g1641(.dina(w_n1656_0[0]),.dinb(w_n1653_0[0]),.dout(n1705),.clk(gclk));
	jor g1642(.dina(w_n1658_0[0]),.dinb(w_n1652_0[0]),.dout(n1706),.clk(gclk));
	jand g1643(.dina(n1706),.dinb(w_dff_B_bI5IHVx85_1),.dout(n1707),.clk(gclk));
	jxor g1644(.dina(w_n1707_0[1]),.dinb(w_n1704_0[1]),.dout(n1708),.clk(gclk));
	jnot g1645(.din(n1708),.dout(n1709),.clk(gclk));
	jxor g1646(.dina(w_n1709_0[1]),.dinb(w_n1703_0[1]),.dout(n1710),.clk(gclk));
	jxor g1647(.dina(w_n1710_0[1]),.dinb(w_n1702_0[1]),.dout(n1711),.clk(gclk));
	jxor g1648(.dina(w_n1711_0[1]),.dinb(w_n1699_0[1]),.dout(n1712),.clk(gclk));
	jxor g1649(.dina(w_n1712_0[1]),.dinb(w_n1697_0[1]),.dout(n1713),.clk(gclk));
	jxor g1650(.dina(w_n1713_0[1]),.dinb(w_n1694_0[1]),.dout(n1714),.clk(gclk));
	jxor g1651(.dina(w_n1714_0[1]),.dinb(w_n1692_0[1]),.dout(n1715),.clk(gclk));
	jxor g1652(.dina(w_n1715_0[1]),.dinb(w_n1689_0[1]),.dout(n1716),.clk(gclk));
	jxor g1653(.dina(w_n1716_0[1]),.dinb(w_n1687_0[1]),.dout(n1717),.clk(gclk));
	jxor g1654(.dina(w_n1717_0[1]),.dinb(w_n1684_0[1]),.dout(n1718),.clk(gclk));
	jnot g1655(.din(n1718),.dout(n1719),.clk(gclk));
	jxor g1656(.dina(w_n1719_0[1]),.dinb(w_n1682_0[1]),.dout(n1720),.clk(gclk));
	jxor g1657(.dina(w_n1720_0[1]),.dinb(w_n1677_0[1]),.dout(w_dff_A_TOoGb41g9_2),.clk(gclk));
	jor g1658(.dina(w_n1719_0[0]),.dinb(w_n1682_0[0]),.dout(n1722),.clk(gclk));
	jnot g1659(.din(w_n1720_0[0]),.dout(n1723),.clk(gclk));
	jor g1660(.dina(w_dff_B_5CmIey8H7_0),.dinb(w_n1677_0[0]),.dout(n1724),.clk(gclk));
	jand g1661(.dina(n1724),.dinb(w_dff_B_XjLyrqrv9_1),.dout(n1725),.clk(gclk));
	jand g1662(.dina(w_n1716_0[0]),.dinb(w_n1687_0[0]),.dout(n1726),.clk(gclk));
	jand g1663(.dina(w_n1717_0[0]),.dinb(w_n1684_0[0]),.dout(n1727),.clk(gclk));
	jor g1664(.dina(n1727),.dinb(w_dff_B_2R8ssFfu8_1),.dout(n1728),.clk(gclk));
	jand g1665(.dina(w_G528gat_3[2]),.dinb(w_G188gat_2[1]),.dout(n1729),.clk(gclk));
	jnot g1666(.din(n1729),.dout(n1730),.clk(gclk));
	jand g1667(.dina(w_n1714_0[0]),.dinb(w_n1692_0[0]),.dout(n1731),.clk(gclk));
	jand g1668(.dina(w_n1715_0[0]),.dinb(w_n1689_0[0]),.dout(n1732),.clk(gclk));
	jor g1669(.dina(n1732),.dinb(w_dff_B_gNgsEzPQ0_1),.dout(n1733),.clk(gclk));
	jand g1670(.dina(w_G511gat_3[1]),.dinb(w_G205gat_2[2]),.dout(n1734),.clk(gclk));
	jnot g1671(.din(n1734),.dout(n1735),.clk(gclk));
	jand g1672(.dina(w_n1712_0[0]),.dinb(w_n1697_0[0]),.dout(n1736),.clk(gclk));
	jand g1673(.dina(w_n1713_0[0]),.dinb(w_n1694_0[0]),.dout(n1737),.clk(gclk));
	jor g1674(.dina(n1737),.dinb(w_dff_B_gC3Rv0z41_1),.dout(n1738),.clk(gclk));
	jand g1675(.dina(w_G494gat_3[0]),.dinb(w_G222gat_3[0]),.dout(n1739),.clk(gclk));
	jnot g1676(.din(n1739),.dout(n1740),.clk(gclk));
	jand g1677(.dina(w_n1710_0[0]),.dinb(w_n1702_0[0]),.dout(n1741),.clk(gclk));
	jand g1678(.dina(w_n1711_0[0]),.dinb(w_n1699_0[0]),.dout(n1742),.clk(gclk));
	jor g1679(.dina(n1742),.dinb(w_dff_B_15EDfjX83_1),.dout(n1743),.clk(gclk));
	jand g1680(.dina(w_G477gat_2[2]),.dinb(w_G239gat_3[1]),.dout(n1744),.clk(gclk));
	jand g1681(.dina(w_G460gat_2[1]),.dinb(w_G256gat_3[2]),.dout(n1745),.clk(gclk));
	jor g1682(.dina(w_n1707_0[0]),.dinb(w_n1704_0[0]),.dout(n1746),.clk(gclk));
	jor g1683(.dina(w_n1709_0[0]),.dinb(w_n1703_0[0]),.dout(n1747),.clk(gclk));
	jand g1684(.dina(n1747),.dinb(w_dff_B_yr9DqX8w2_1),.dout(n1748),.clk(gclk));
	jxor g1685(.dina(w_n1748_0[1]),.dinb(w_n1745_0[1]),.dout(n1749),.clk(gclk));
	jnot g1686(.din(n1749),.dout(n1750),.clk(gclk));
	jxor g1687(.dina(w_n1750_0[1]),.dinb(w_n1744_0[1]),.dout(n1751),.clk(gclk));
	jxor g1688(.dina(w_n1751_0[1]),.dinb(w_n1743_0[1]),.dout(n1752),.clk(gclk));
	jxor g1689(.dina(w_n1752_0[1]),.dinb(w_n1740_0[1]),.dout(n1753),.clk(gclk));
	jxor g1690(.dina(w_n1753_0[1]),.dinb(w_n1738_0[1]),.dout(n1754),.clk(gclk));
	jxor g1691(.dina(w_n1754_0[1]),.dinb(w_n1735_0[1]),.dout(n1755),.clk(gclk));
	jxor g1692(.dina(w_n1755_0[1]),.dinb(w_n1733_0[1]),.dout(n1756),.clk(gclk));
	jxor g1693(.dina(w_n1756_0[1]),.dinb(w_n1730_0[1]),.dout(n1757),.clk(gclk));
	jxor g1694(.dina(w_n1757_0[1]),.dinb(w_n1728_0[1]),.dout(n1758),.clk(gclk));
	jxor g1695(.dina(w_n1758_0[1]),.dinb(w_n1725_0[1]),.dout(w_dff_A_CFydfasb0_2),.clk(gclk));
	jnot g1696(.din(w_n1728_0[0]),.dout(n1760),.clk(gclk));
	jnot g1697(.din(w_n1757_0[0]),.dout(n1761),.clk(gclk));
	jor g1698(.dina(n1761),.dinb(w_dff_B_e7rQmgAM9_1),.dout(n1762),.clk(gclk));
	jnot g1699(.din(w_n1758_0[0]),.dout(n1763),.clk(gclk));
	jor g1700(.dina(w_dff_B_W6zUBB6O9_0),.dinb(w_n1725_0[0]),.dout(n1764),.clk(gclk));
	jand g1701(.dina(n1764),.dinb(w_dff_B_yshrl5Ud5_1),.dout(n1765),.clk(gclk));
	jand g1702(.dina(w_n1755_0[0]),.dinb(w_n1733_0[0]),.dout(n1766),.clk(gclk));
	jand g1703(.dina(w_n1756_0[0]),.dinb(w_n1730_0[0]),.dout(n1767),.clk(gclk));
	jor g1704(.dina(n1767),.dinb(w_dff_B_GY0AmhZ59_1),.dout(n1768),.clk(gclk));
	jand g1705(.dina(w_G528gat_3[1]),.dinb(w_G205gat_2[1]),.dout(n1769),.clk(gclk));
	jnot g1706(.din(n1769),.dout(n1770),.clk(gclk));
	jand g1707(.dina(w_n1753_0[0]),.dinb(w_n1738_0[0]),.dout(n1771),.clk(gclk));
	jand g1708(.dina(w_n1754_0[0]),.dinb(w_n1735_0[0]),.dout(n1772),.clk(gclk));
	jor g1709(.dina(n1772),.dinb(w_dff_B_41ptGfqe8_1),.dout(n1773),.clk(gclk));
	jand g1710(.dina(w_G511gat_3[0]),.dinb(w_G222gat_2[2]),.dout(n1774),.clk(gclk));
	jnot g1711(.din(n1774),.dout(n1775),.clk(gclk));
	jand g1712(.dina(w_n1751_0[0]),.dinb(w_n1743_0[0]),.dout(n1776),.clk(gclk));
	jand g1713(.dina(w_n1752_0[0]),.dinb(w_n1740_0[0]),.dout(n1777),.clk(gclk));
	jor g1714(.dina(n1777),.dinb(w_dff_B_4H58eYGh5_1),.dout(n1778),.clk(gclk));
	jand g1715(.dina(w_G494gat_2[2]),.dinb(w_G239gat_3[0]),.dout(n1779),.clk(gclk));
	jand g1716(.dina(w_G477gat_2[1]),.dinb(w_G256gat_3[1]),.dout(n1780),.clk(gclk));
	jor g1717(.dina(w_n1748_0[0]),.dinb(w_n1745_0[0]),.dout(n1781),.clk(gclk));
	jor g1718(.dina(w_n1750_0[0]),.dinb(w_n1744_0[0]),.dout(n1782),.clk(gclk));
	jand g1719(.dina(n1782),.dinb(w_dff_B_hxknXZrK4_1),.dout(n1783),.clk(gclk));
	jxor g1720(.dina(w_n1783_0[1]),.dinb(w_n1780_0[1]),.dout(n1784),.clk(gclk));
	jnot g1721(.din(n1784),.dout(n1785),.clk(gclk));
	jxor g1722(.dina(w_n1785_0[1]),.dinb(w_n1779_0[1]),.dout(n1786),.clk(gclk));
	jxor g1723(.dina(w_n1786_0[1]),.dinb(w_n1778_0[1]),.dout(n1787),.clk(gclk));
	jxor g1724(.dina(w_n1787_0[1]),.dinb(w_n1775_0[1]),.dout(n1788),.clk(gclk));
	jxor g1725(.dina(w_n1788_0[1]),.dinb(w_n1773_0[1]),.dout(n1789),.clk(gclk));
	jxor g1726(.dina(w_n1789_0[1]),.dinb(w_n1770_0[1]),.dout(n1790),.clk(gclk));
	jxor g1727(.dina(w_n1790_0[1]),.dinb(w_n1768_0[1]),.dout(n1791),.clk(gclk));
	jxor g1728(.dina(w_n1791_0[1]),.dinb(w_n1765_0[1]),.dout(w_dff_A_J0Xe6gJm8_2),.clk(gclk));
	jnot g1729(.din(w_n1768_0[0]),.dout(n1793),.clk(gclk));
	jnot g1730(.din(w_n1790_0[0]),.dout(n1794),.clk(gclk));
	jor g1731(.dina(n1794),.dinb(w_dff_B_r5DeWLnr2_1),.dout(n1795),.clk(gclk));
	jnot g1732(.din(w_n1791_0[0]),.dout(n1796),.clk(gclk));
	jor g1733(.dina(w_dff_B_sqeRZOro5_0),.dinb(w_n1765_0[0]),.dout(n1797),.clk(gclk));
	jand g1734(.dina(n1797),.dinb(w_dff_B_7um8b3989_1),.dout(n1798),.clk(gclk));
	jand g1735(.dina(w_n1788_0[0]),.dinb(w_n1773_0[0]),.dout(n1799),.clk(gclk));
	jand g1736(.dina(w_n1789_0[0]),.dinb(w_n1770_0[0]),.dout(n1800),.clk(gclk));
	jor g1737(.dina(n1800),.dinb(w_dff_B_mSbZR5nX4_1),.dout(n1801),.clk(gclk));
	jand g1738(.dina(w_G528gat_3[0]),.dinb(w_G222gat_2[1]),.dout(n1802),.clk(gclk));
	jnot g1739(.din(n1802),.dout(n1803),.clk(gclk));
	jand g1740(.dina(w_n1786_0[0]),.dinb(w_n1778_0[0]),.dout(n1804),.clk(gclk));
	jand g1741(.dina(w_n1787_0[0]),.dinb(w_n1775_0[0]),.dout(n1805),.clk(gclk));
	jor g1742(.dina(n1805),.dinb(w_dff_B_HZcRA8yf1_1),.dout(n1806),.clk(gclk));
	jand g1743(.dina(w_G511gat_2[2]),.dinb(w_G239gat_2[2]),.dout(n1807),.clk(gclk));
	jand g1744(.dina(w_G494gat_2[1]),.dinb(w_G256gat_3[0]),.dout(n1808),.clk(gclk));
	jor g1745(.dina(w_n1783_0[0]),.dinb(w_n1780_0[0]),.dout(n1809),.clk(gclk));
	jor g1746(.dina(w_n1785_0[0]),.dinb(w_n1779_0[0]),.dout(n1810),.clk(gclk));
	jand g1747(.dina(n1810),.dinb(w_dff_B_4p6E7E1O0_1),.dout(n1811),.clk(gclk));
	jxor g1748(.dina(w_n1811_0[1]),.dinb(w_n1808_0[1]),.dout(n1812),.clk(gclk));
	jnot g1749(.din(n1812),.dout(n1813),.clk(gclk));
	jxor g1750(.dina(w_n1813_0[1]),.dinb(w_n1807_0[1]),.dout(n1814),.clk(gclk));
	jxor g1751(.dina(w_n1814_0[1]),.dinb(w_n1806_0[1]),.dout(n1815),.clk(gclk));
	jxor g1752(.dina(w_n1815_0[1]),.dinb(w_n1803_0[1]),.dout(n1816),.clk(gclk));
	jxor g1753(.dina(w_n1816_0[1]),.dinb(w_n1801_0[1]),.dout(n1817),.clk(gclk));
	jxor g1754(.dina(w_n1817_0[1]),.dinb(w_n1798_0[1]),.dout(w_dff_A_kkcMHLRb7_2),.clk(gclk));
	jnot g1755(.din(w_n1801_0[0]),.dout(n1819),.clk(gclk));
	jnot g1756(.din(w_n1816_0[0]),.dout(n1820),.clk(gclk));
	jor g1757(.dina(n1820),.dinb(w_dff_B_LOyfXsth5_1),.dout(n1821),.clk(gclk));
	jnot g1758(.din(w_n1817_0[0]),.dout(n1822),.clk(gclk));
	jor g1759(.dina(w_dff_B_E29MaRkv1_0),.dinb(w_n1798_0[0]),.dout(n1823),.clk(gclk));
	jand g1760(.dina(n1823),.dinb(w_dff_B_bXC1YG0R2_1),.dout(n1824),.clk(gclk));
	jand g1761(.dina(w_n1814_0[0]),.dinb(w_n1806_0[0]),.dout(n1825),.clk(gclk));
	jand g1762(.dina(w_n1815_0[0]),.dinb(w_n1803_0[0]),.dout(n1826),.clk(gclk));
	jor g1763(.dina(n1826),.dinb(w_dff_B_C92hqvgL8_1),.dout(n1827),.clk(gclk));
	jand g1764(.dina(w_G528gat_2[2]),.dinb(w_G239gat_2[1]),.dout(n1828),.clk(gclk));
	jand g1765(.dina(w_G511gat_2[1]),.dinb(w_G256gat_2[2]),.dout(n1829),.clk(gclk));
	jor g1766(.dina(w_n1811_0[0]),.dinb(w_n1808_0[0]),.dout(n1830),.clk(gclk));
	jor g1767(.dina(w_n1813_0[0]),.dinb(w_n1807_0[0]),.dout(n1831),.clk(gclk));
	jand g1768(.dina(n1831),.dinb(w_dff_B_UPlWjVfl7_1),.dout(n1832),.clk(gclk));
	jxor g1769(.dina(w_n1832_0[1]),.dinb(w_n1829_0[1]),.dout(n1833),.clk(gclk));
	jnot g1770(.din(n1833),.dout(n1834),.clk(gclk));
	jxor g1771(.dina(w_n1834_0[1]),.dinb(w_n1828_0[1]),.dout(n1835),.clk(gclk));
	jxor g1772(.dina(w_n1835_0[1]),.dinb(w_n1827_0[1]),.dout(n1836),.clk(gclk));
	jxor g1773(.dina(w_n1836_0[1]),.dinb(w_n1824_0[1]),.dout(w_dff_A_2YEfK94H7_2),.clk(gclk));
	jand g1774(.dina(w_G528gat_2[1]),.dinb(w_G256gat_2[1]),.dout(n1838),.clk(gclk));
	jor g1775(.dina(w_n1832_0[0]),.dinb(w_n1829_0[0]),.dout(n1839),.clk(gclk));
	jor g1776(.dina(w_n1834_0[0]),.dinb(w_n1828_0[0]),.dout(n1840),.clk(gclk));
	jand g1777(.dina(n1840),.dinb(w_dff_B_WeG7aV7r0_1),.dout(n1841),.clk(gclk));
	jor g1778(.dina(w_n1841_0[1]),.dinb(w_n1838_0[1]),.dout(n1842),.clk(gclk));
	jnot g1779(.din(w_n1827_0[0]),.dout(n1843),.clk(gclk));
	jnot g1780(.din(w_n1835_0[0]),.dout(n1844),.clk(gclk));
	jor g1781(.dina(n1844),.dinb(w_dff_B_081Xrddf4_1),.dout(n1845),.clk(gclk));
	jnot g1782(.din(w_n1836_0[0]),.dout(n1846),.clk(gclk));
	jor g1783(.dina(w_dff_B_SRiaM2L53_0),.dinb(w_n1824_0[0]),.dout(n1847),.clk(gclk));
	jand g1784(.dina(n1847),.dinb(w_dff_B_axl2M9jY6_1),.dout(n1848),.clk(gclk));
	jxor g1785(.dina(w_n1841_0[0]),.dinb(w_n1838_0[0]),.dout(n1849),.clk(gclk));
	jnot g1786(.din(w_n1849_0[1]),.dout(n1850),.clk(gclk));
	jor g1787(.dina(w_dff_B_6I7wTHAp0_0),.dinb(w_n1848_0[1]),.dout(n1851),.clk(gclk));
	jand g1788(.dina(n1851),.dinb(w_dff_B_AJQXN7UJ4_1),.dout(G6287gat),.clk(gclk));
	jxor g1789(.dina(w_n1849_0[0]),.dinb(w_n1848_0[0]),.dout(w_dff_A_rdgwxBzJ1_2),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_G1gat_0[0]),.doutb(w_G1gat_0[1]),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G1gat_1(.douta(w_G1gat_1[0]),.doutb(w_G1gat_1[1]),.doutc(w_G1gat_1[2]),.din(w_G1gat_0[0]));
	jspl3 jspl3_w_G1gat_2(.douta(w_G1gat_2[0]),.doutb(w_G1gat_2[1]),.doutc(w_G1gat_2[2]),.din(w_G1gat_0[1]));
	jspl3 jspl3_w_G1gat_3(.douta(w_G1gat_3[0]),.doutb(w_G1gat_3[1]),.doutc(w_G1gat_3[2]),.din(w_G1gat_0[2]));
	jspl3 jspl3_w_G1gat_4(.douta(w_G1gat_4[0]),.doutb(w_G1gat_4[1]),.doutc(w_G1gat_4[2]),.din(w_G1gat_1[0]));
	jspl3 jspl3_w_G1gat_5(.douta(w_G1gat_5[0]),.doutb(w_G1gat_5[1]),.doutc(w_G1gat_5[2]),.din(w_G1gat_1[1]));
	jspl3 jspl3_w_G1gat_6(.douta(w_G1gat_6[0]),.doutb(w_G1gat_6[1]),.doutc(w_G1gat_6[2]),.din(w_G1gat_1[2]));
	jspl jspl_w_G1gat_7(.douta(w_G1gat_7[0]),.doutb(w_G1gat_7[1]),.din(w_G1gat_2[0]));
	jspl3 jspl3_w_G18gat_0(.douta(w_G18gat_0[0]),.doutb(w_G18gat_0[1]),.doutc(w_G18gat_0[2]),.din(G18gat));
	jspl3 jspl3_w_G18gat_1(.douta(w_G18gat_1[0]),.doutb(w_G18gat_1[1]),.doutc(w_G18gat_1[2]),.din(w_G18gat_0[0]));
	jspl3 jspl3_w_G18gat_2(.douta(w_G18gat_2[0]),.doutb(w_G18gat_2[1]),.doutc(w_G18gat_2[2]),.din(w_G18gat_0[1]));
	jspl3 jspl3_w_G18gat_3(.douta(w_G18gat_3[0]),.doutb(w_G18gat_3[1]),.doutc(w_G18gat_3[2]),.din(w_G18gat_0[2]));
	jspl3 jspl3_w_G18gat_4(.douta(w_G18gat_4[0]),.doutb(w_G18gat_4[1]),.doutc(w_G18gat_4[2]),.din(w_G18gat_1[0]));
	jspl3 jspl3_w_G18gat_5(.douta(w_G18gat_5[0]),.doutb(w_G18gat_5[1]),.doutc(w_G18gat_5[2]),.din(w_G18gat_1[1]));
	jspl3 jspl3_w_G18gat_6(.douta(w_G18gat_6[0]),.doutb(w_G18gat_6[1]),.doutc(w_G18gat_6[2]),.din(w_G18gat_1[2]));
	jspl3 jspl3_w_G18gat_7(.douta(w_G18gat_7[0]),.doutb(w_G18gat_7[1]),.doutc(w_G18gat_7[2]),.din(w_G18gat_2[0]));
	jspl3 jspl3_w_G35gat_0(.douta(w_G35gat_0[0]),.doutb(w_G35gat_0[1]),.doutc(w_G35gat_0[2]),.din(G35gat));
	jspl3 jspl3_w_G35gat_1(.douta(w_G35gat_1[0]),.doutb(w_G35gat_1[1]),.doutc(w_G35gat_1[2]),.din(w_G35gat_0[0]));
	jspl3 jspl3_w_G35gat_2(.douta(w_G35gat_2[0]),.doutb(w_G35gat_2[1]),.doutc(w_G35gat_2[2]),.din(w_G35gat_0[1]));
	jspl3 jspl3_w_G35gat_3(.douta(w_G35gat_3[0]),.doutb(w_G35gat_3[1]),.doutc(w_G35gat_3[2]),.din(w_G35gat_0[2]));
	jspl3 jspl3_w_G35gat_4(.douta(w_G35gat_4[0]),.doutb(w_G35gat_4[1]),.doutc(w_G35gat_4[2]),.din(w_G35gat_1[0]));
	jspl3 jspl3_w_G35gat_5(.douta(w_G35gat_5[0]),.doutb(w_G35gat_5[1]),.doutc(w_G35gat_5[2]),.din(w_G35gat_1[1]));
	jspl3 jspl3_w_G35gat_6(.douta(w_G35gat_6[0]),.doutb(w_G35gat_6[1]),.doutc(w_G35gat_6[2]),.din(w_G35gat_1[2]));
	jspl3 jspl3_w_G35gat_7(.douta(w_G35gat_7[0]),.doutb(w_G35gat_7[1]),.doutc(w_G35gat_7[2]),.din(w_G35gat_2[0]));
	jspl3 jspl3_w_G52gat_0(.douta(w_G52gat_0[0]),.doutb(w_G52gat_0[1]),.doutc(w_G52gat_0[2]),.din(G52gat));
	jspl3 jspl3_w_G52gat_1(.douta(w_G52gat_1[0]),.doutb(w_G52gat_1[1]),.doutc(w_G52gat_1[2]),.din(w_G52gat_0[0]));
	jspl3 jspl3_w_G52gat_2(.douta(w_G52gat_2[0]),.doutb(w_G52gat_2[1]),.doutc(w_G52gat_2[2]),.din(w_G52gat_0[1]));
	jspl3 jspl3_w_G52gat_3(.douta(w_G52gat_3[0]),.doutb(w_G52gat_3[1]),.doutc(w_G52gat_3[2]),.din(w_G52gat_0[2]));
	jspl3 jspl3_w_G52gat_4(.douta(w_G52gat_4[0]),.doutb(w_G52gat_4[1]),.doutc(w_G52gat_4[2]),.din(w_G52gat_1[0]));
	jspl3 jspl3_w_G52gat_5(.douta(w_G52gat_5[0]),.doutb(w_G52gat_5[1]),.doutc(w_G52gat_5[2]),.din(w_G52gat_1[1]));
	jspl3 jspl3_w_G52gat_6(.douta(w_G52gat_6[0]),.doutb(w_G52gat_6[1]),.doutc(w_G52gat_6[2]),.din(w_G52gat_1[2]));
	jspl3 jspl3_w_G52gat_7(.douta(w_G52gat_7[0]),.doutb(w_G52gat_7[1]),.doutc(w_G52gat_7[2]),.din(w_G52gat_2[0]));
	jspl3 jspl3_w_G69gat_0(.douta(w_G69gat_0[0]),.doutb(w_G69gat_0[1]),.doutc(w_G69gat_0[2]),.din(G69gat));
	jspl3 jspl3_w_G69gat_1(.douta(w_G69gat_1[0]),.doutb(w_G69gat_1[1]),.doutc(w_G69gat_1[2]),.din(w_G69gat_0[0]));
	jspl3 jspl3_w_G69gat_2(.douta(w_G69gat_2[0]),.doutb(w_G69gat_2[1]),.doutc(w_G69gat_2[2]),.din(w_G69gat_0[1]));
	jspl3 jspl3_w_G69gat_3(.douta(w_G69gat_3[0]),.doutb(w_G69gat_3[1]),.doutc(w_G69gat_3[2]),.din(w_G69gat_0[2]));
	jspl3 jspl3_w_G69gat_4(.douta(w_G69gat_4[0]),.doutb(w_G69gat_4[1]),.doutc(w_G69gat_4[2]),.din(w_G69gat_1[0]));
	jspl3 jspl3_w_G69gat_5(.douta(w_G69gat_5[0]),.doutb(w_G69gat_5[1]),.doutc(w_G69gat_5[2]),.din(w_G69gat_1[1]));
	jspl3 jspl3_w_G69gat_6(.douta(w_G69gat_6[0]),.doutb(w_G69gat_6[1]),.doutc(w_G69gat_6[2]),.din(w_G69gat_1[2]));
	jspl jspl_w_G69gat_7(.douta(w_G69gat_7[0]),.doutb(w_G69gat_7[1]),.din(w_G69gat_2[0]));
	jspl3 jspl3_w_G86gat_0(.douta(w_G86gat_0[0]),.doutb(w_G86gat_0[1]),.doutc(w_G86gat_0[2]),.din(G86gat));
	jspl3 jspl3_w_G86gat_1(.douta(w_G86gat_1[0]),.doutb(w_G86gat_1[1]),.doutc(w_G86gat_1[2]),.din(w_G86gat_0[0]));
	jspl3 jspl3_w_G86gat_2(.douta(w_G86gat_2[0]),.doutb(w_G86gat_2[1]),.doutc(w_G86gat_2[2]),.din(w_G86gat_0[1]));
	jspl3 jspl3_w_G86gat_3(.douta(w_G86gat_3[0]),.doutb(w_G86gat_3[1]),.doutc(w_G86gat_3[2]),.din(w_G86gat_0[2]));
	jspl3 jspl3_w_G86gat_4(.douta(w_G86gat_4[0]),.doutb(w_G86gat_4[1]),.doutc(w_G86gat_4[2]),.din(w_G86gat_1[0]));
	jspl3 jspl3_w_G86gat_5(.douta(w_G86gat_5[0]),.doutb(w_G86gat_5[1]),.doutc(w_G86gat_5[2]),.din(w_G86gat_1[1]));
	jspl3 jspl3_w_G86gat_6(.douta(w_G86gat_6[0]),.doutb(w_G86gat_6[1]),.doutc(w_G86gat_6[2]),.din(w_G86gat_1[2]));
	jspl jspl_w_G86gat_7(.douta(w_G86gat_7[0]),.doutb(w_G86gat_7[1]),.din(w_G86gat_2[0]));
	jspl3 jspl3_w_G103gat_0(.douta(w_G103gat_0[0]),.doutb(w_G103gat_0[1]),.doutc(w_G103gat_0[2]),.din(G103gat));
	jspl3 jspl3_w_G103gat_1(.douta(w_G103gat_1[0]),.doutb(w_G103gat_1[1]),.doutc(w_G103gat_1[2]),.din(w_G103gat_0[0]));
	jspl3 jspl3_w_G103gat_2(.douta(w_G103gat_2[0]),.doutb(w_G103gat_2[1]),.doutc(w_G103gat_2[2]),.din(w_G103gat_0[1]));
	jspl3 jspl3_w_G103gat_3(.douta(w_G103gat_3[0]),.doutb(w_G103gat_3[1]),.doutc(w_G103gat_3[2]),.din(w_G103gat_0[2]));
	jspl3 jspl3_w_G103gat_4(.douta(w_G103gat_4[0]),.doutb(w_G103gat_4[1]),.doutc(w_G103gat_4[2]),.din(w_G103gat_1[0]));
	jspl3 jspl3_w_G103gat_5(.douta(w_G103gat_5[0]),.doutb(w_G103gat_5[1]),.doutc(w_G103gat_5[2]),.din(w_G103gat_1[1]));
	jspl3 jspl3_w_G103gat_6(.douta(w_G103gat_6[0]),.doutb(w_G103gat_6[1]),.doutc(w_G103gat_6[2]),.din(w_G103gat_1[2]));
	jspl jspl_w_G103gat_7(.douta(w_G103gat_7[0]),.doutb(w_G103gat_7[1]),.din(w_G103gat_2[0]));
	jspl3 jspl3_w_G120gat_0(.douta(w_G120gat_0[0]),.doutb(w_G120gat_0[1]),.doutc(w_G120gat_0[2]),.din(G120gat));
	jspl3 jspl3_w_G120gat_1(.douta(w_G120gat_1[0]),.doutb(w_G120gat_1[1]),.doutc(w_G120gat_1[2]),.din(w_G120gat_0[0]));
	jspl3 jspl3_w_G120gat_2(.douta(w_G120gat_2[0]),.doutb(w_G120gat_2[1]),.doutc(w_G120gat_2[2]),.din(w_G120gat_0[1]));
	jspl3 jspl3_w_G120gat_3(.douta(w_G120gat_3[0]),.doutb(w_G120gat_3[1]),.doutc(w_G120gat_3[2]),.din(w_G120gat_0[2]));
	jspl3 jspl3_w_G120gat_4(.douta(w_G120gat_4[0]),.doutb(w_G120gat_4[1]),.doutc(w_G120gat_4[2]),.din(w_G120gat_1[0]));
	jspl3 jspl3_w_G120gat_5(.douta(w_G120gat_5[0]),.doutb(w_G120gat_5[1]),.doutc(w_G120gat_5[2]),.din(w_G120gat_1[1]));
	jspl3 jspl3_w_G120gat_6(.douta(w_G120gat_6[0]),.doutb(w_G120gat_6[1]),.doutc(w_G120gat_6[2]),.din(w_G120gat_1[2]));
	jspl jspl_w_G120gat_7(.douta(w_G120gat_7[0]),.doutb(w_G120gat_7[1]),.din(w_G120gat_2[0]));
	jspl3 jspl3_w_G137gat_0(.douta(w_G137gat_0[0]),.doutb(w_G137gat_0[1]),.doutc(w_G137gat_0[2]),.din(G137gat));
	jspl3 jspl3_w_G137gat_1(.douta(w_G137gat_1[0]),.doutb(w_G137gat_1[1]),.doutc(w_G137gat_1[2]),.din(w_G137gat_0[0]));
	jspl3 jspl3_w_G137gat_2(.douta(w_G137gat_2[0]),.doutb(w_G137gat_2[1]),.doutc(w_G137gat_2[2]),.din(w_G137gat_0[1]));
	jspl3 jspl3_w_G137gat_3(.douta(w_G137gat_3[0]),.doutb(w_G137gat_3[1]),.doutc(w_G137gat_3[2]),.din(w_G137gat_0[2]));
	jspl3 jspl3_w_G137gat_4(.douta(w_G137gat_4[0]),.doutb(w_G137gat_4[1]),.doutc(w_G137gat_4[2]),.din(w_G137gat_1[0]));
	jspl3 jspl3_w_G137gat_5(.douta(w_G137gat_5[0]),.doutb(w_G137gat_5[1]),.doutc(w_G137gat_5[2]),.din(w_G137gat_1[1]));
	jspl3 jspl3_w_G137gat_6(.douta(w_G137gat_6[0]),.doutb(w_G137gat_6[1]),.doutc(w_G137gat_6[2]),.din(w_G137gat_1[2]));
	jspl jspl_w_G137gat_7(.douta(w_G137gat_7[0]),.doutb(w_G137gat_7[1]),.din(w_G137gat_2[0]));
	jspl3 jspl3_w_G154gat_0(.douta(w_G154gat_0[0]),.doutb(w_G154gat_0[1]),.doutc(w_G154gat_0[2]),.din(G154gat));
	jspl3 jspl3_w_G154gat_1(.douta(w_G154gat_1[0]),.doutb(w_G154gat_1[1]),.doutc(w_G154gat_1[2]),.din(w_G154gat_0[0]));
	jspl3 jspl3_w_G154gat_2(.douta(w_G154gat_2[0]),.doutb(w_G154gat_2[1]),.doutc(w_G154gat_2[2]),.din(w_G154gat_0[1]));
	jspl3 jspl3_w_G154gat_3(.douta(w_G154gat_3[0]),.doutb(w_G154gat_3[1]),.doutc(w_G154gat_3[2]),.din(w_G154gat_0[2]));
	jspl3 jspl3_w_G154gat_4(.douta(w_G154gat_4[0]),.doutb(w_G154gat_4[1]),.doutc(w_G154gat_4[2]),.din(w_G154gat_1[0]));
	jspl3 jspl3_w_G154gat_5(.douta(w_G154gat_5[0]),.doutb(w_G154gat_5[1]),.doutc(w_G154gat_5[2]),.din(w_G154gat_1[1]));
	jspl3 jspl3_w_G154gat_6(.douta(w_G154gat_6[0]),.doutb(w_G154gat_6[1]),.doutc(w_G154gat_6[2]),.din(w_G154gat_1[2]));
	jspl jspl_w_G154gat_7(.douta(w_G154gat_7[0]),.doutb(w_G154gat_7[1]),.din(w_G154gat_2[0]));
	jspl3 jspl3_w_G171gat_0(.douta(w_G171gat_0[0]),.doutb(w_G171gat_0[1]),.doutc(w_G171gat_0[2]),.din(G171gat));
	jspl3 jspl3_w_G171gat_1(.douta(w_G171gat_1[0]),.doutb(w_G171gat_1[1]),.doutc(w_G171gat_1[2]),.din(w_G171gat_0[0]));
	jspl3 jspl3_w_G171gat_2(.douta(w_G171gat_2[0]),.doutb(w_G171gat_2[1]),.doutc(w_G171gat_2[2]),.din(w_G171gat_0[1]));
	jspl3 jspl3_w_G171gat_3(.douta(w_G171gat_3[0]),.doutb(w_G171gat_3[1]),.doutc(w_G171gat_3[2]),.din(w_G171gat_0[2]));
	jspl3 jspl3_w_G171gat_4(.douta(w_G171gat_4[0]),.doutb(w_G171gat_4[1]),.doutc(w_G171gat_4[2]),.din(w_G171gat_1[0]));
	jspl3 jspl3_w_G171gat_5(.douta(w_G171gat_5[0]),.doutb(w_G171gat_5[1]),.doutc(w_G171gat_5[2]),.din(w_G171gat_1[1]));
	jspl3 jspl3_w_G171gat_6(.douta(w_G171gat_6[0]),.doutb(w_G171gat_6[1]),.doutc(w_G171gat_6[2]),.din(w_G171gat_1[2]));
	jspl jspl_w_G171gat_7(.douta(w_G171gat_7[0]),.doutb(w_G171gat_7[1]),.din(w_G171gat_2[0]));
	jspl3 jspl3_w_G188gat_0(.douta(w_G188gat_0[0]),.doutb(w_G188gat_0[1]),.doutc(w_G188gat_0[2]),.din(G188gat));
	jspl3 jspl3_w_G188gat_1(.douta(w_G188gat_1[0]),.doutb(w_G188gat_1[1]),.doutc(w_G188gat_1[2]),.din(w_G188gat_0[0]));
	jspl3 jspl3_w_G188gat_2(.douta(w_G188gat_2[0]),.doutb(w_G188gat_2[1]),.doutc(w_G188gat_2[2]),.din(w_G188gat_0[1]));
	jspl3 jspl3_w_G188gat_3(.douta(w_G188gat_3[0]),.doutb(w_G188gat_3[1]),.doutc(w_G188gat_3[2]),.din(w_G188gat_0[2]));
	jspl3 jspl3_w_G188gat_4(.douta(w_G188gat_4[0]),.doutb(w_G188gat_4[1]),.doutc(w_G188gat_4[2]),.din(w_G188gat_1[0]));
	jspl3 jspl3_w_G188gat_5(.douta(w_G188gat_5[0]),.doutb(w_G188gat_5[1]),.doutc(w_G188gat_5[2]),.din(w_G188gat_1[1]));
	jspl3 jspl3_w_G188gat_6(.douta(w_G188gat_6[0]),.doutb(w_G188gat_6[1]),.doutc(w_G188gat_6[2]),.din(w_G188gat_1[2]));
	jspl jspl_w_G188gat_7(.douta(w_G188gat_7[0]),.doutb(w_G188gat_7[1]),.din(w_G188gat_2[0]));
	jspl3 jspl3_w_G205gat_0(.douta(w_G205gat_0[0]),.doutb(w_G205gat_0[1]),.doutc(w_G205gat_0[2]),.din(G205gat));
	jspl3 jspl3_w_G205gat_1(.douta(w_G205gat_1[0]),.doutb(w_G205gat_1[1]),.doutc(w_G205gat_1[2]),.din(w_G205gat_0[0]));
	jspl3 jspl3_w_G205gat_2(.douta(w_G205gat_2[0]),.doutb(w_G205gat_2[1]),.doutc(w_G205gat_2[2]),.din(w_G205gat_0[1]));
	jspl3 jspl3_w_G205gat_3(.douta(w_G205gat_3[0]),.doutb(w_G205gat_3[1]),.doutc(w_G205gat_3[2]),.din(w_G205gat_0[2]));
	jspl3 jspl3_w_G205gat_4(.douta(w_G205gat_4[0]),.doutb(w_G205gat_4[1]),.doutc(w_G205gat_4[2]),.din(w_G205gat_1[0]));
	jspl3 jspl3_w_G205gat_5(.douta(w_G205gat_5[0]),.doutb(w_G205gat_5[1]),.doutc(w_G205gat_5[2]),.din(w_G205gat_1[1]));
	jspl3 jspl3_w_G205gat_6(.douta(w_G205gat_6[0]),.doutb(w_G205gat_6[1]),.doutc(w_G205gat_6[2]),.din(w_G205gat_1[2]));
	jspl jspl_w_G205gat_7(.douta(w_G205gat_7[0]),.doutb(w_G205gat_7[1]),.din(w_G205gat_2[0]));
	jspl3 jspl3_w_G222gat_0(.douta(w_G222gat_0[0]),.doutb(w_G222gat_0[1]),.doutc(w_G222gat_0[2]),.din(G222gat));
	jspl3 jspl3_w_G222gat_1(.douta(w_G222gat_1[0]),.doutb(w_G222gat_1[1]),.doutc(w_G222gat_1[2]),.din(w_G222gat_0[0]));
	jspl3 jspl3_w_G222gat_2(.douta(w_G222gat_2[0]),.doutb(w_G222gat_2[1]),.doutc(w_G222gat_2[2]),.din(w_G222gat_0[1]));
	jspl3 jspl3_w_G222gat_3(.douta(w_G222gat_3[0]),.doutb(w_G222gat_3[1]),.doutc(w_G222gat_3[2]),.din(w_G222gat_0[2]));
	jspl3 jspl3_w_G222gat_4(.douta(w_G222gat_4[0]),.doutb(w_G222gat_4[1]),.doutc(w_G222gat_4[2]),.din(w_G222gat_1[0]));
	jspl3 jspl3_w_G222gat_5(.douta(w_G222gat_5[0]),.doutb(w_G222gat_5[1]),.doutc(w_G222gat_5[2]),.din(w_G222gat_1[1]));
	jspl3 jspl3_w_G222gat_6(.douta(w_G222gat_6[0]),.doutb(w_G222gat_6[1]),.doutc(w_G222gat_6[2]),.din(w_G222gat_1[2]));
	jspl jspl_w_G222gat_7(.douta(w_G222gat_7[0]),.doutb(w_G222gat_7[1]),.din(w_G222gat_2[0]));
	jspl3 jspl3_w_G239gat_0(.douta(w_G239gat_0[0]),.doutb(w_G239gat_0[1]),.doutc(w_G239gat_0[2]),.din(G239gat));
	jspl3 jspl3_w_G239gat_1(.douta(w_G239gat_1[0]),.doutb(w_G239gat_1[1]),.doutc(w_G239gat_1[2]),.din(w_G239gat_0[0]));
	jspl3 jspl3_w_G239gat_2(.douta(w_G239gat_2[0]),.doutb(w_G239gat_2[1]),.doutc(w_G239gat_2[2]),.din(w_G239gat_0[1]));
	jspl3 jspl3_w_G239gat_3(.douta(w_G239gat_3[0]),.doutb(w_G239gat_3[1]),.doutc(w_G239gat_3[2]),.din(w_G239gat_0[2]));
	jspl3 jspl3_w_G239gat_4(.douta(w_G239gat_4[0]),.doutb(w_G239gat_4[1]),.doutc(w_G239gat_4[2]),.din(w_G239gat_1[0]));
	jspl3 jspl3_w_G239gat_5(.douta(w_G239gat_5[0]),.doutb(w_G239gat_5[1]),.doutc(w_G239gat_5[2]),.din(w_G239gat_1[1]));
	jspl3 jspl3_w_G239gat_6(.douta(w_G239gat_6[0]),.doutb(w_G239gat_6[1]),.doutc(w_G239gat_6[2]),.din(w_G239gat_1[2]));
	jspl jspl_w_G239gat_7(.douta(w_G239gat_7[0]),.doutb(w_G239gat_7[1]),.din(w_G239gat_2[0]));
	jspl3 jspl3_w_G256gat_0(.douta(w_G256gat_0[0]),.doutb(w_G256gat_0[1]),.doutc(w_G256gat_0[2]),.din(G256gat));
	jspl3 jspl3_w_G256gat_1(.douta(w_G256gat_1[0]),.doutb(w_G256gat_1[1]),.doutc(w_G256gat_1[2]),.din(w_G256gat_0[0]));
	jspl3 jspl3_w_G256gat_2(.douta(w_G256gat_2[0]),.doutb(w_G256gat_2[1]),.doutc(w_G256gat_2[2]),.din(w_G256gat_0[1]));
	jspl3 jspl3_w_G256gat_3(.douta(w_G256gat_3[0]),.doutb(w_G256gat_3[1]),.doutc(w_G256gat_3[2]),.din(w_G256gat_0[2]));
	jspl3 jspl3_w_G256gat_4(.douta(w_G256gat_4[0]),.doutb(w_G256gat_4[1]),.doutc(w_G256gat_4[2]),.din(w_G256gat_1[0]));
	jspl3 jspl3_w_G256gat_5(.douta(w_G256gat_5[0]),.doutb(w_G256gat_5[1]),.doutc(w_G256gat_5[2]),.din(w_G256gat_1[1]));
	jspl3 jspl3_w_G256gat_6(.douta(w_G256gat_6[0]),.doutb(w_G256gat_6[1]),.doutc(w_G256gat_6[2]),.din(w_G256gat_1[2]));
	jspl jspl_w_G256gat_7(.douta(w_G256gat_7[0]),.doutb(w_G256gat_7[1]),.din(w_G256gat_2[0]));
	jspl3 jspl3_w_G273gat_0(.douta(w_G273gat_0[0]),.doutb(w_G273gat_0[1]),.doutc(w_G273gat_0[2]),.din(G273gat));
	jspl3 jspl3_w_G273gat_1(.douta(w_G273gat_1[0]),.doutb(w_G273gat_1[1]),.doutc(w_G273gat_1[2]),.din(w_G273gat_0[0]));
	jspl3 jspl3_w_G273gat_2(.douta(w_G273gat_2[0]),.doutb(w_G273gat_2[1]),.doutc(w_G273gat_2[2]),.din(w_G273gat_0[1]));
	jspl3 jspl3_w_G273gat_3(.douta(w_G273gat_3[0]),.doutb(w_G273gat_3[1]),.doutc(w_G273gat_3[2]),.din(w_G273gat_0[2]));
	jspl3 jspl3_w_G273gat_4(.douta(w_G273gat_4[0]),.doutb(w_G273gat_4[1]),.doutc(w_G273gat_4[2]),.din(w_G273gat_1[0]));
	jspl3 jspl3_w_G273gat_5(.douta(w_G273gat_5[0]),.doutb(w_G273gat_5[1]),.doutc(w_G273gat_5[2]),.din(w_G273gat_1[1]));
	jspl3 jspl3_w_G273gat_6(.douta(w_G273gat_6[0]),.doutb(w_G273gat_6[1]),.doutc(w_G273gat_6[2]),.din(w_G273gat_1[2]));
	jspl3 jspl3_w_G273gat_7(.douta(w_G273gat_7[0]),.doutb(w_G273gat_7[1]),.doutc(w_G273gat_7[2]),.din(w_G273gat_2[0]));
	jspl3 jspl3_w_G290gat_0(.douta(w_G290gat_0[0]),.doutb(w_G290gat_0[1]),.doutc(w_G290gat_0[2]),.din(G290gat));
	jspl3 jspl3_w_G290gat_1(.douta(w_G290gat_1[0]),.doutb(w_G290gat_1[1]),.doutc(w_G290gat_1[2]),.din(w_G290gat_0[0]));
	jspl3 jspl3_w_G290gat_2(.douta(w_G290gat_2[0]),.doutb(w_G290gat_2[1]),.doutc(w_G290gat_2[2]),.din(w_G290gat_0[1]));
	jspl3 jspl3_w_G290gat_3(.douta(w_G290gat_3[0]),.doutb(w_G290gat_3[1]),.doutc(w_G290gat_3[2]),.din(w_G290gat_0[2]));
	jspl3 jspl3_w_G290gat_4(.douta(w_G290gat_4[0]),.doutb(w_G290gat_4[1]),.doutc(w_G290gat_4[2]),.din(w_G290gat_1[0]));
	jspl3 jspl3_w_G290gat_5(.douta(w_G290gat_5[0]),.doutb(w_G290gat_5[1]),.doutc(w_G290gat_5[2]),.din(w_G290gat_1[1]));
	jspl3 jspl3_w_G290gat_6(.douta(w_G290gat_6[0]),.doutb(w_G290gat_6[1]),.doutc(w_G290gat_6[2]),.din(w_G290gat_1[2]));
	jspl3 jspl3_w_G290gat_7(.douta(w_G290gat_7[0]),.doutb(w_G290gat_7[1]),.doutc(w_G290gat_7[2]),.din(w_G290gat_2[0]));
	jspl3 jspl3_w_G307gat_0(.douta(w_G307gat_0[0]),.doutb(w_G307gat_0[1]),.doutc(w_G307gat_0[2]),.din(G307gat));
	jspl3 jspl3_w_G307gat_1(.douta(w_G307gat_1[0]),.doutb(w_G307gat_1[1]),.doutc(w_G307gat_1[2]),.din(w_G307gat_0[0]));
	jspl3 jspl3_w_G307gat_2(.douta(w_G307gat_2[0]),.doutb(w_dff_A_RSjd2ENx5_1),.doutc(w_G307gat_2[2]),.din(w_G307gat_0[1]));
	jspl3 jspl3_w_G307gat_3(.douta(w_G307gat_3[0]),.doutb(w_G307gat_3[1]),.doutc(w_G307gat_3[2]),.din(w_G307gat_0[2]));
	jspl3 jspl3_w_G307gat_4(.douta(w_G307gat_4[0]),.doutb(w_G307gat_4[1]),.doutc(w_G307gat_4[2]),.din(w_G307gat_1[0]));
	jspl3 jspl3_w_G307gat_5(.douta(w_G307gat_5[0]),.doutb(w_G307gat_5[1]),.doutc(w_G307gat_5[2]),.din(w_G307gat_1[1]));
	jspl3 jspl3_w_G307gat_6(.douta(w_G307gat_6[0]),.doutb(w_G307gat_6[1]),.doutc(w_G307gat_6[2]),.din(w_G307gat_1[2]));
	jspl3 jspl3_w_G307gat_7(.douta(w_G307gat_7[0]),.doutb(w_G307gat_7[1]),.doutc(w_G307gat_7[2]),.din(w_G307gat_2[0]));
	jspl3 jspl3_w_G324gat_0(.douta(w_G324gat_0[0]),.doutb(w_G324gat_0[1]),.doutc(w_G324gat_0[2]),.din(G324gat));
	jspl3 jspl3_w_G324gat_1(.douta(w_G324gat_1[0]),.doutb(w_G324gat_1[1]),.doutc(w_G324gat_1[2]),.din(w_G324gat_0[0]));
	jspl3 jspl3_w_G324gat_2(.douta(w_G324gat_2[0]),.doutb(w_G324gat_2[1]),.doutc(w_G324gat_2[2]),.din(w_G324gat_0[1]));
	jspl3 jspl3_w_G324gat_3(.douta(w_G324gat_3[0]),.doutb(w_G324gat_3[1]),.doutc(w_G324gat_3[2]),.din(w_G324gat_0[2]));
	jspl3 jspl3_w_G324gat_4(.douta(w_G324gat_4[0]),.doutb(w_G324gat_4[1]),.doutc(w_G324gat_4[2]),.din(w_G324gat_1[0]));
	jspl3 jspl3_w_G324gat_5(.douta(w_G324gat_5[0]),.doutb(w_G324gat_5[1]),.doutc(w_G324gat_5[2]),.din(w_G324gat_1[1]));
	jspl3 jspl3_w_G324gat_6(.douta(w_G324gat_6[0]),.doutb(w_G324gat_6[1]),.doutc(w_G324gat_6[2]),.din(w_G324gat_1[2]));
	jspl jspl_w_G324gat_7(.douta(w_G324gat_7[0]),.doutb(w_G324gat_7[1]),.din(w_G324gat_2[0]));
	jspl3 jspl3_w_G341gat_0(.douta(w_G341gat_0[0]),.doutb(w_G341gat_0[1]),.doutc(w_G341gat_0[2]),.din(G341gat));
	jspl3 jspl3_w_G341gat_1(.douta(w_G341gat_1[0]),.doutb(w_G341gat_1[1]),.doutc(w_G341gat_1[2]),.din(w_G341gat_0[0]));
	jspl3 jspl3_w_G341gat_2(.douta(w_G341gat_2[0]),.doutb(w_G341gat_2[1]),.doutc(w_G341gat_2[2]),.din(w_G341gat_0[1]));
	jspl3 jspl3_w_G341gat_3(.douta(w_G341gat_3[0]),.doutb(w_G341gat_3[1]),.doutc(w_G341gat_3[2]),.din(w_G341gat_0[2]));
	jspl3 jspl3_w_G341gat_4(.douta(w_G341gat_4[0]),.doutb(w_G341gat_4[1]),.doutc(w_G341gat_4[2]),.din(w_G341gat_1[0]));
	jspl3 jspl3_w_G341gat_5(.douta(w_G341gat_5[0]),.doutb(w_G341gat_5[1]),.doutc(w_G341gat_5[2]),.din(w_G341gat_1[1]));
	jspl3 jspl3_w_G341gat_6(.douta(w_G341gat_6[0]),.doutb(w_G341gat_6[1]),.doutc(w_G341gat_6[2]),.din(w_G341gat_1[2]));
	jspl jspl_w_G341gat_7(.douta(w_G341gat_7[0]),.doutb(w_G341gat_7[1]),.din(w_G341gat_2[0]));
	jspl3 jspl3_w_G358gat_0(.douta(w_G358gat_0[0]),.doutb(w_G358gat_0[1]),.doutc(w_G358gat_0[2]),.din(G358gat));
	jspl3 jspl3_w_G358gat_1(.douta(w_G358gat_1[0]),.doutb(w_G358gat_1[1]),.doutc(w_G358gat_1[2]),.din(w_G358gat_0[0]));
	jspl3 jspl3_w_G358gat_2(.douta(w_G358gat_2[0]),.doutb(w_G358gat_2[1]),.doutc(w_G358gat_2[2]),.din(w_G358gat_0[1]));
	jspl3 jspl3_w_G358gat_3(.douta(w_G358gat_3[0]),.doutb(w_G358gat_3[1]),.doutc(w_G358gat_3[2]),.din(w_G358gat_0[2]));
	jspl3 jspl3_w_G358gat_4(.douta(w_G358gat_4[0]),.doutb(w_G358gat_4[1]),.doutc(w_G358gat_4[2]),.din(w_G358gat_1[0]));
	jspl3 jspl3_w_G358gat_5(.douta(w_G358gat_5[0]),.doutb(w_G358gat_5[1]),.doutc(w_G358gat_5[2]),.din(w_G358gat_1[1]));
	jspl3 jspl3_w_G358gat_6(.douta(w_G358gat_6[0]),.doutb(w_G358gat_6[1]),.doutc(w_G358gat_6[2]),.din(w_G358gat_1[2]));
	jspl jspl_w_G358gat_7(.douta(w_G358gat_7[0]),.doutb(w_G358gat_7[1]),.din(w_G358gat_2[0]));
	jspl3 jspl3_w_G375gat_0(.douta(w_G375gat_0[0]),.doutb(w_G375gat_0[1]),.doutc(w_G375gat_0[2]),.din(G375gat));
	jspl3 jspl3_w_G375gat_1(.douta(w_G375gat_1[0]),.doutb(w_G375gat_1[1]),.doutc(w_G375gat_1[2]),.din(w_G375gat_0[0]));
	jspl3 jspl3_w_G375gat_2(.douta(w_G375gat_2[0]),.doutb(w_G375gat_2[1]),.doutc(w_G375gat_2[2]),.din(w_G375gat_0[1]));
	jspl3 jspl3_w_G375gat_3(.douta(w_G375gat_3[0]),.doutb(w_G375gat_3[1]),.doutc(w_G375gat_3[2]),.din(w_G375gat_0[2]));
	jspl3 jspl3_w_G375gat_4(.douta(w_G375gat_4[0]),.doutb(w_G375gat_4[1]),.doutc(w_G375gat_4[2]),.din(w_G375gat_1[0]));
	jspl3 jspl3_w_G375gat_5(.douta(w_G375gat_5[0]),.doutb(w_G375gat_5[1]),.doutc(w_G375gat_5[2]),.din(w_G375gat_1[1]));
	jspl3 jspl3_w_G375gat_6(.douta(w_G375gat_6[0]),.doutb(w_G375gat_6[1]),.doutc(w_G375gat_6[2]),.din(w_G375gat_1[2]));
	jspl jspl_w_G375gat_7(.douta(w_G375gat_7[0]),.doutb(w_G375gat_7[1]),.din(w_G375gat_2[0]));
	jspl3 jspl3_w_G392gat_0(.douta(w_G392gat_0[0]),.doutb(w_G392gat_0[1]),.doutc(w_G392gat_0[2]),.din(G392gat));
	jspl3 jspl3_w_G392gat_1(.douta(w_G392gat_1[0]),.doutb(w_G392gat_1[1]),.doutc(w_G392gat_1[2]),.din(w_G392gat_0[0]));
	jspl3 jspl3_w_G392gat_2(.douta(w_G392gat_2[0]),.doutb(w_G392gat_2[1]),.doutc(w_G392gat_2[2]),.din(w_G392gat_0[1]));
	jspl3 jspl3_w_G392gat_3(.douta(w_G392gat_3[0]),.doutb(w_G392gat_3[1]),.doutc(w_G392gat_3[2]),.din(w_G392gat_0[2]));
	jspl3 jspl3_w_G392gat_4(.douta(w_G392gat_4[0]),.doutb(w_G392gat_4[1]),.doutc(w_G392gat_4[2]),.din(w_G392gat_1[0]));
	jspl3 jspl3_w_G392gat_5(.douta(w_G392gat_5[0]),.doutb(w_G392gat_5[1]),.doutc(w_G392gat_5[2]),.din(w_G392gat_1[1]));
	jspl3 jspl3_w_G392gat_6(.douta(w_G392gat_6[0]),.doutb(w_G392gat_6[1]),.doutc(w_G392gat_6[2]),.din(w_G392gat_1[2]));
	jspl jspl_w_G392gat_7(.douta(w_G392gat_7[0]),.doutb(w_G392gat_7[1]),.din(w_G392gat_2[0]));
	jspl3 jspl3_w_G409gat_0(.douta(w_G409gat_0[0]),.doutb(w_G409gat_0[1]),.doutc(w_G409gat_0[2]),.din(G409gat));
	jspl3 jspl3_w_G409gat_1(.douta(w_G409gat_1[0]),.doutb(w_G409gat_1[1]),.doutc(w_G409gat_1[2]),.din(w_G409gat_0[0]));
	jspl3 jspl3_w_G409gat_2(.douta(w_G409gat_2[0]),.doutb(w_G409gat_2[1]),.doutc(w_G409gat_2[2]),.din(w_G409gat_0[1]));
	jspl3 jspl3_w_G409gat_3(.douta(w_G409gat_3[0]),.doutb(w_G409gat_3[1]),.doutc(w_G409gat_3[2]),.din(w_G409gat_0[2]));
	jspl3 jspl3_w_G409gat_4(.douta(w_G409gat_4[0]),.doutb(w_G409gat_4[1]),.doutc(w_G409gat_4[2]),.din(w_G409gat_1[0]));
	jspl3 jspl3_w_G409gat_5(.douta(w_G409gat_5[0]),.doutb(w_G409gat_5[1]),.doutc(w_G409gat_5[2]),.din(w_G409gat_1[1]));
	jspl3 jspl3_w_G409gat_6(.douta(w_G409gat_6[0]),.doutb(w_G409gat_6[1]),.doutc(w_G409gat_6[2]),.din(w_G409gat_1[2]));
	jspl jspl_w_G409gat_7(.douta(w_G409gat_7[0]),.doutb(w_G409gat_7[1]),.din(w_G409gat_2[0]));
	jspl3 jspl3_w_G426gat_0(.douta(w_G426gat_0[0]),.doutb(w_G426gat_0[1]),.doutc(w_G426gat_0[2]),.din(G426gat));
	jspl3 jspl3_w_G426gat_1(.douta(w_G426gat_1[0]),.doutb(w_G426gat_1[1]),.doutc(w_G426gat_1[2]),.din(w_G426gat_0[0]));
	jspl3 jspl3_w_G426gat_2(.douta(w_G426gat_2[0]),.doutb(w_G426gat_2[1]),.doutc(w_G426gat_2[2]),.din(w_G426gat_0[1]));
	jspl3 jspl3_w_G426gat_3(.douta(w_G426gat_3[0]),.doutb(w_G426gat_3[1]),.doutc(w_G426gat_3[2]),.din(w_G426gat_0[2]));
	jspl3 jspl3_w_G426gat_4(.douta(w_G426gat_4[0]),.doutb(w_G426gat_4[1]),.doutc(w_G426gat_4[2]),.din(w_G426gat_1[0]));
	jspl3 jspl3_w_G426gat_5(.douta(w_G426gat_5[0]),.doutb(w_G426gat_5[1]),.doutc(w_G426gat_5[2]),.din(w_G426gat_1[1]));
	jspl3 jspl3_w_G426gat_6(.douta(w_G426gat_6[0]),.doutb(w_G426gat_6[1]),.doutc(w_G426gat_6[2]),.din(w_G426gat_1[2]));
	jspl jspl_w_G426gat_7(.douta(w_G426gat_7[0]),.doutb(w_G426gat_7[1]),.din(w_G426gat_2[0]));
	jspl3 jspl3_w_G443gat_0(.douta(w_G443gat_0[0]),.doutb(w_G443gat_0[1]),.doutc(w_G443gat_0[2]),.din(G443gat));
	jspl3 jspl3_w_G443gat_1(.douta(w_G443gat_1[0]),.doutb(w_G443gat_1[1]),.doutc(w_G443gat_1[2]),.din(w_G443gat_0[0]));
	jspl3 jspl3_w_G443gat_2(.douta(w_G443gat_2[0]),.doutb(w_G443gat_2[1]),.doutc(w_G443gat_2[2]),.din(w_G443gat_0[1]));
	jspl3 jspl3_w_G443gat_3(.douta(w_G443gat_3[0]),.doutb(w_G443gat_3[1]),.doutc(w_G443gat_3[2]),.din(w_G443gat_0[2]));
	jspl3 jspl3_w_G443gat_4(.douta(w_G443gat_4[0]),.doutb(w_G443gat_4[1]),.doutc(w_G443gat_4[2]),.din(w_G443gat_1[0]));
	jspl3 jspl3_w_G443gat_5(.douta(w_G443gat_5[0]),.doutb(w_G443gat_5[1]),.doutc(w_G443gat_5[2]),.din(w_G443gat_1[1]));
	jspl3 jspl3_w_G443gat_6(.douta(w_G443gat_6[0]),.doutb(w_G443gat_6[1]),.doutc(w_G443gat_6[2]),.din(w_G443gat_1[2]));
	jspl jspl_w_G443gat_7(.douta(w_G443gat_7[0]),.doutb(w_G443gat_7[1]),.din(w_G443gat_2[0]));
	jspl3 jspl3_w_G460gat_0(.douta(w_G460gat_0[0]),.doutb(w_G460gat_0[1]),.doutc(w_G460gat_0[2]),.din(G460gat));
	jspl3 jspl3_w_G460gat_1(.douta(w_G460gat_1[0]),.doutb(w_G460gat_1[1]),.doutc(w_G460gat_1[2]),.din(w_G460gat_0[0]));
	jspl3 jspl3_w_G460gat_2(.douta(w_G460gat_2[0]),.doutb(w_G460gat_2[1]),.doutc(w_G460gat_2[2]),.din(w_G460gat_0[1]));
	jspl3 jspl3_w_G460gat_3(.douta(w_G460gat_3[0]),.doutb(w_G460gat_3[1]),.doutc(w_G460gat_3[2]),.din(w_G460gat_0[2]));
	jspl3 jspl3_w_G460gat_4(.douta(w_G460gat_4[0]),.doutb(w_G460gat_4[1]),.doutc(w_G460gat_4[2]),.din(w_G460gat_1[0]));
	jspl3 jspl3_w_G460gat_5(.douta(w_G460gat_5[0]),.doutb(w_G460gat_5[1]),.doutc(w_G460gat_5[2]),.din(w_G460gat_1[1]));
	jspl3 jspl3_w_G460gat_6(.douta(w_G460gat_6[0]),.doutb(w_G460gat_6[1]),.doutc(w_G460gat_6[2]),.din(w_G460gat_1[2]));
	jspl jspl_w_G460gat_7(.douta(w_G460gat_7[0]),.doutb(w_G460gat_7[1]),.din(w_G460gat_2[0]));
	jspl3 jspl3_w_G477gat_0(.douta(w_G477gat_0[0]),.doutb(w_G477gat_0[1]),.doutc(w_G477gat_0[2]),.din(G477gat));
	jspl3 jspl3_w_G477gat_1(.douta(w_G477gat_1[0]),.doutb(w_G477gat_1[1]),.doutc(w_G477gat_1[2]),.din(w_G477gat_0[0]));
	jspl3 jspl3_w_G477gat_2(.douta(w_G477gat_2[0]),.doutb(w_G477gat_2[1]),.doutc(w_G477gat_2[2]),.din(w_G477gat_0[1]));
	jspl3 jspl3_w_G477gat_3(.douta(w_G477gat_3[0]),.doutb(w_G477gat_3[1]),.doutc(w_G477gat_3[2]),.din(w_G477gat_0[2]));
	jspl3 jspl3_w_G477gat_4(.douta(w_G477gat_4[0]),.doutb(w_G477gat_4[1]),.doutc(w_G477gat_4[2]),.din(w_G477gat_1[0]));
	jspl3 jspl3_w_G477gat_5(.douta(w_G477gat_5[0]),.doutb(w_G477gat_5[1]),.doutc(w_G477gat_5[2]),.din(w_G477gat_1[1]));
	jspl3 jspl3_w_G477gat_6(.douta(w_G477gat_6[0]),.doutb(w_G477gat_6[1]),.doutc(w_G477gat_6[2]),.din(w_G477gat_1[2]));
	jspl jspl_w_G477gat_7(.douta(w_G477gat_7[0]),.doutb(w_G477gat_7[1]),.din(w_G477gat_2[0]));
	jspl3 jspl3_w_G494gat_0(.douta(w_G494gat_0[0]),.doutb(w_G494gat_0[1]),.doutc(w_G494gat_0[2]),.din(G494gat));
	jspl3 jspl3_w_G494gat_1(.douta(w_G494gat_1[0]),.doutb(w_G494gat_1[1]),.doutc(w_G494gat_1[2]),.din(w_G494gat_0[0]));
	jspl3 jspl3_w_G494gat_2(.douta(w_G494gat_2[0]),.doutb(w_G494gat_2[1]),.doutc(w_G494gat_2[2]),.din(w_G494gat_0[1]));
	jspl3 jspl3_w_G494gat_3(.douta(w_G494gat_3[0]),.doutb(w_G494gat_3[1]),.doutc(w_G494gat_3[2]),.din(w_G494gat_0[2]));
	jspl3 jspl3_w_G494gat_4(.douta(w_G494gat_4[0]),.doutb(w_G494gat_4[1]),.doutc(w_G494gat_4[2]),.din(w_G494gat_1[0]));
	jspl3 jspl3_w_G494gat_5(.douta(w_G494gat_5[0]),.doutb(w_G494gat_5[1]),.doutc(w_G494gat_5[2]),.din(w_G494gat_1[1]));
	jspl3 jspl3_w_G494gat_6(.douta(w_G494gat_6[0]),.doutb(w_G494gat_6[1]),.doutc(w_G494gat_6[2]),.din(w_G494gat_1[2]));
	jspl jspl_w_G494gat_7(.douta(w_G494gat_7[0]),.doutb(w_G494gat_7[1]),.din(w_G494gat_2[0]));
	jspl3 jspl3_w_G511gat_0(.douta(w_G511gat_0[0]),.doutb(w_G511gat_0[1]),.doutc(w_G511gat_0[2]),.din(G511gat));
	jspl3 jspl3_w_G511gat_1(.douta(w_G511gat_1[0]),.doutb(w_G511gat_1[1]),.doutc(w_G511gat_1[2]),.din(w_G511gat_0[0]));
	jspl3 jspl3_w_G511gat_2(.douta(w_G511gat_2[0]),.doutb(w_G511gat_2[1]),.doutc(w_G511gat_2[2]),.din(w_G511gat_0[1]));
	jspl3 jspl3_w_G511gat_3(.douta(w_G511gat_3[0]),.doutb(w_G511gat_3[1]),.doutc(w_G511gat_3[2]),.din(w_G511gat_0[2]));
	jspl3 jspl3_w_G511gat_4(.douta(w_G511gat_4[0]),.doutb(w_G511gat_4[1]),.doutc(w_G511gat_4[2]),.din(w_G511gat_1[0]));
	jspl3 jspl3_w_G511gat_5(.douta(w_G511gat_5[0]),.doutb(w_G511gat_5[1]),.doutc(w_G511gat_5[2]),.din(w_G511gat_1[1]));
	jspl3 jspl3_w_G511gat_6(.douta(w_G511gat_6[0]),.doutb(w_G511gat_6[1]),.doutc(w_G511gat_6[2]),.din(w_G511gat_1[2]));
	jspl jspl_w_G511gat_7(.douta(w_G511gat_7[0]),.doutb(w_G511gat_7[1]),.din(w_G511gat_2[0]));
	jspl3 jspl3_w_G528gat_0(.douta(w_G528gat_0[0]),.doutb(w_G528gat_0[1]),.doutc(w_G528gat_0[2]),.din(G528gat));
	jspl3 jspl3_w_G528gat_1(.douta(w_G528gat_1[0]),.doutb(w_G528gat_1[1]),.doutc(w_G528gat_1[2]),.din(w_G528gat_0[0]));
	jspl3 jspl3_w_G528gat_2(.douta(w_G528gat_2[0]),.doutb(w_G528gat_2[1]),.doutc(w_G528gat_2[2]),.din(w_G528gat_0[1]));
	jspl3 jspl3_w_G528gat_3(.douta(w_G528gat_3[0]),.doutb(w_G528gat_3[1]),.doutc(w_G528gat_3[2]),.din(w_G528gat_0[2]));
	jspl3 jspl3_w_G528gat_4(.douta(w_G528gat_4[0]),.doutb(w_G528gat_4[1]),.doutc(w_G528gat_4[2]),.din(w_G528gat_1[0]));
	jspl3 jspl3_w_G528gat_5(.douta(w_G528gat_5[0]),.doutb(w_G528gat_5[1]),.doutc(w_G528gat_5[2]),.din(w_G528gat_1[1]));
	jspl3 jspl3_w_G528gat_6(.douta(w_G528gat_6[0]),.doutb(w_G528gat_6[1]),.doutc(w_G528gat_6[2]),.din(w_G528gat_1[2]));
	jspl jspl_w_G528gat_7(.douta(w_G528gat_7[0]),.doutb(w_G528gat_7[1]),.din(w_G528gat_2[0]));
	jspl jspl_w_G545gat_0(.douta(w_G545gat_0),.doutb(w_dff_A_OnSTmqyq1_1),.din(G545gat_fa_));
	jspl jspl_w_n65_0(.douta(w_n65_0[0]),.doutb(w_n65_0[1]),.din(n65));
	jspl jspl_w_n69_0(.douta(w_dff_A_YDMEMreQ6_0),.doutb(w_n69_0[1]),.din(n69));
	jspl jspl_w_n70_0(.douta(w_dff_A_x31Ir6Po7_0),.doutb(w_n70_0[1]),.din(n70));
	jspl jspl_w_n72_0(.douta(w_dff_A_OX7nFsGl7_0),.doutb(w_n72_0[1]),.din(n72));
	jspl jspl_w_n75_0(.douta(w_n75_0[0]),.doutb(w_n75_0[1]),.din(n75));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl jspl_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.din(n78));
	jspl jspl_w_n81_0(.douta(w_n81_0[0]),.doutb(w_n81_0[1]),.din(n81));
	jspl3 jspl3_w_n82_0(.douta(w_n82_0[0]),.doutb(w_dff_A_balw0lKA6_1),.doutc(w_dff_A_jO2YVfKU2_2),.din(n82));
	jspl jspl_w_n82_1(.douta(w_n82_1[0]),.doutb(w_dff_A_latRsa6l4_1),.din(w_n82_0[0]));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n85_0(.douta(w_dff_A_MmWWRJ4h6_0),.doutb(w_n85_0[1]),.din(n85));
	jspl jspl_w_n87_0(.douta(w_n87_0[0]),.doutb(w_n87_0[1]),.din(n87));
	jspl jspl_w_n89_0(.douta(w_dff_A_kiy2BO7f5_0),.doutb(w_n89_0[1]),.din(n89));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl jspl_w_n94_0(.douta(w_dff_A_GfrnQwgt6_0),.doutb(w_n94_0[1]),.din(n94));
	jspl jspl_w_n96_0(.douta(w_n96_0[0]),.doutb(w_n96_0[1]),.din(n96));
	jspl jspl_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.din(n99));
	jspl3 jspl3_w_n100_0(.douta(w_n100_0[0]),.doutb(w_dff_A_8BlzFoWF9_1),.doutc(w_dff_A_ZXYPmR2t3_2),.din(n100));
	jspl jspl_w_n100_1(.douta(w_dff_A_9S0is7Qi5_0),.doutb(w_n100_1[1]),.din(w_n100_0[0]));
	jspl3 jspl3_w_n101_0(.douta(w_dff_A_D2IVofeZ1_0),.doutb(w_n101_0[1]),.doutc(w_n101_0[2]),.din(n101));
	jspl jspl_w_n103_0(.douta(w_dff_A_nDVYqqP91_0),.doutb(w_n103_0[1]),.din(n103));
	jspl jspl_w_n104_0(.douta(w_dff_A_tW1bCqem0_0),.doutb(w_n104_0[1]),.din(n104));
	jspl jspl_w_n107_0(.douta(w_n107_0[0]),.doutb(w_dff_A_4iAploSe2_1),.din(n107));
	jspl jspl_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n110_0(.douta(w_dff_A_EVKqHyce1_0),.doutb(w_n110_0[1]),.din(n110));
	jspl jspl_w_n115_0(.douta(w_n115_0[0]),.doutb(w_n115_0[1]),.din(n115));
	jspl jspl_w_n116_0(.douta(w_dff_A_NiDcVqga0_0),.doutb(w_n116_0[1]),.din(n116));
	jspl3 jspl3_w_n126_0(.douta(w_n126_0[0]),.doutb(w_n126_0[1]),.doutc(w_n126_0[2]),.din(n126));
	jspl jspl_w_n128_0(.douta(w_n128_0[0]),.doutb(w_n128_0[1]),.din(w_dff_B_s8Xsddgu1_2));
	jspl jspl_w_n129_0(.douta(w_n129_0[0]),.doutb(w_n129_0[1]),.din(n129));
	jspl jspl_w_n130_0(.douta(w_n130_0[0]),.doutb(w_dff_A_R32qMOHF2_1),.din(n130));
	jspl jspl_w_n131_0(.douta(w_n131_0[0]),.doutb(w_n131_0[1]),.din(n131));
	jspl3 jspl3_w_n132_0(.douta(w_dff_A_kW5i3c4R9_0),.doutb(w_dff_A_fhzCCFL74_1),.doutc(w_n132_0[2]),.din(n132));
	jspl3 jspl3_w_n133_0(.douta(w_n133_0[0]),.doutb(w_n133_0[1]),.doutc(w_n133_0[2]),.din(n133));
	jspl jspl_w_n138_0(.douta(w_n138_0[0]),.doutb(w_n138_0[1]),.din(n138));
	jspl jspl_w_n139_0(.douta(w_dff_A_SwFztyXO9_0),.doutb(w_n139_0[1]),.din(n139));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl jspl_w_n142_0(.douta(w_n142_0[0]),.doutb(w_dff_A_Bw9625kf4_1),.din(n142));
	jspl jspl_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.din(n143));
	jspl jspl_w_n145_0(.douta(w_dff_A_vuvYPKsd0_0),.doutb(w_n145_0[1]),.din(n145));
	jspl jspl_w_n150_0(.douta(w_n150_0[0]),.doutb(w_n150_0[1]),.din(n150));
	jspl jspl_w_n151_0(.douta(w_dff_A_HWEN1MZi5_0),.doutb(w_n151_0[1]),.din(n151));
	jspl3 jspl3_w_n156_0(.douta(w_n156_0[0]),.doutb(w_n156_0[1]),.doutc(w_n156_0[2]),.din(n156));
	jspl jspl_w_n158_0(.douta(w_n158_0[0]),.doutb(w_n158_0[1]),.din(w_dff_B_p6mphz8N5_2));
	jspl jspl_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.din(n163));
	jspl jspl_w_n165_0(.douta(w_n165_0[0]),.doutb(w_n165_0[1]),.din(w_dff_B_MwjjekUY8_2));
	jspl jspl_w_n166_0(.douta(w_n166_0[0]),.doutb(w_n166_0[1]),.din(n166));
	jspl jspl_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.din(n168));
	jspl3 jspl3_w_n169_0(.douta(w_dff_A_S5jpLcNQ9_0),.doutb(w_dff_A_0436c07I2_1),.doutc(w_n169_0[2]),.din(n169));
	jspl jspl_w_n170_0(.douta(w_n170_0[0]),.doutb(w_n170_0[1]),.din(n170));
	jspl jspl_w_n172_0(.douta(w_n172_0[0]),.doutb(w_n172_0[1]),.din(n172));
	jspl jspl_w_n174_0(.douta(w_n174_0[0]),.doutb(w_n174_0[1]),.din(n174));
	jspl jspl_w_n175_0(.douta(w_n175_0[0]),.doutb(w_n175_0[1]),.din(w_dff_B_JHKovzKr2_2));
	jspl jspl_w_n176_0(.douta(w_n176_0[0]),.doutb(w_n176_0[1]),.din(n176));
	jspl jspl_w_n177_0(.douta(w_dff_A_AQPO0Rr33_0),.doutb(w_n177_0[1]),.din(n177));
	jspl jspl_w_n178_0(.douta(w_n178_0[0]),.doutb(w_n178_0[1]),.din(n178));
	jspl jspl_w_n180_0(.douta(w_n180_0[0]),.doutb(w_dff_A_abjFZba61_1),.din(n180));
	jspl jspl_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.din(n181));
	jspl jspl_w_n183_0(.douta(w_dff_A_wIZmNCxX4_0),.doutb(w_n183_0[1]),.din(n183));
	jspl jspl_w_n188_0(.douta(w_n188_0[0]),.doutb(w_n188_0[1]),.din(n188));
	jspl jspl_w_n189_0(.douta(w_dff_A_4hwEkcxO6_0),.doutb(w_n189_0[1]),.din(n189));
	jspl3 jspl3_w_n194_0(.douta(w_n194_0[0]),.doutb(w_n194_0[1]),.doutc(w_n194_0[2]),.din(n194));
	jspl jspl_w_n196_0(.douta(w_n196_0[0]),.doutb(w_n196_0[1]),.din(w_dff_B_tViMIGoP6_2));
	jspl jspl_w_n199_0(.douta(w_n199_0[0]),.doutb(w_n199_0[1]),.din(n199));
	jspl jspl_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.din(w_dff_B_8cqyc2hd9_2));
	jspl jspl_w_n204_0(.douta(w_n204_0[0]),.doutb(w_n204_0[1]),.din(n204));
	jspl jspl_w_n206_0(.douta(w_n206_0[0]),.doutb(w_n206_0[1]),.din(w_dff_B_sgCcalFI4_2));
	jspl jspl_w_n207_0(.douta(w_n207_0[0]),.doutb(w_n207_0[1]),.din(n207));
	jspl jspl_w_n209_0(.douta(w_n209_0[0]),.doutb(w_n209_0[1]),.din(n209));
	jspl3 jspl3_w_n210_0(.douta(w_n210_0[0]),.doutb(w_dff_A_mTvMtSiG7_1),.doutc(w_dff_A_Y3Yw9DWj9_2),.din(n210));
	jspl jspl_w_n210_1(.douta(w_dff_A_1dikcfgM7_0),.doutb(w_n210_1[1]),.din(w_n210_0[0]));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_n213_0[1]),.din(n213));
	jspl jspl_w_n215_0(.douta(w_n215_0[0]),.doutb(w_n215_0[1]),.din(n215));
	jspl jspl_w_n216_0(.douta(w_n216_0[0]),.doutb(w_n216_0[1]),.din(w_dff_B_NuTfgCbl3_2));
	jspl jspl_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.din(n217));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.din(w_dff_B_LYxRxdqy1_2));
	jspl jspl_w_n219_0(.douta(w_n219_0[0]),.doutb(w_n219_0[1]),.din(n219));
	jspl jspl_w_n220_0(.douta(w_dff_A_UvMWN99Q9_0),.doutb(w_n220_0[1]),.din(n220));
	jspl jspl_w_n221_0(.douta(w_n221_0[0]),.doutb(w_n221_0[1]),.din(n221));
	jspl jspl_w_n223_0(.douta(w_n223_0[0]),.doutb(w_dff_A_G11zUqc14_1),.din(n223));
	jspl jspl_w_n224_0(.douta(w_n224_0[0]),.doutb(w_n224_0[1]),.din(n224));
	jspl jspl_w_n226_0(.douta(w_dff_A_JPXdPWUu5_0),.doutb(w_n226_0[1]),.din(n226));
	jspl jspl_w_n231_0(.douta(w_n231_0[0]),.doutb(w_n231_0[1]),.din(n231));
	jspl jspl_w_n232_0(.douta(w_dff_A_9rl5Eyhd7_0),.doutb(w_n232_0[1]),.din(n232));
	jspl3 jspl3_w_n237_0(.douta(w_n237_0[0]),.doutb(w_n237_0[1]),.doutc(w_n237_0[2]),.din(n237));
	jspl jspl_w_n239_0(.douta(w_n239_0[0]),.doutb(w_n239_0[1]),.din(w_dff_B_psODmytO6_2));
	jspl jspl_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.din(n242));
	jspl jspl_w_n244_0(.douta(w_n244_0[0]),.doutb(w_n244_0[1]),.din(w_dff_B_kXxIFRYn3_2));
	jspl jspl_w_n247_0(.douta(w_n247_0[0]),.doutb(w_n247_0[1]),.din(n247));
	jspl jspl_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.din(w_dff_B_NzaK6og78_2));
	jspl jspl_w_n252_0(.douta(w_n252_0[0]),.doutb(w_n252_0[1]),.din(n252));
	jspl jspl_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.din(w_dff_B_u3Vi490M7_2));
	jspl jspl_w_n255_0(.douta(w_n255_0[0]),.doutb(w_n255_0[1]),.din(n255));
	jspl jspl_w_n257_0(.douta(w_n257_0[0]),.doutb(w_n257_0[1]),.din(n257));
	jspl3 jspl3_w_n258_0(.douta(w_dff_A_AvuFHgdL3_0),.doutb(w_dff_A_jWxdfK7Z8_1),.doutc(w_n258_0[2]),.din(n258));
	jspl jspl_w_n259_0(.douta(w_n259_0[0]),.doutb(w_n259_0[1]),.din(n259));
	jspl jspl_w_n261_0(.douta(w_n261_0[0]),.doutb(w_n261_0[1]),.din(n261));
	jspl jspl_w_n264_0(.douta(w_n264_0[0]),.doutb(w_n264_0[1]),.din(n264));
	jspl jspl_w_n265_0(.douta(w_n265_0[0]),.doutb(w_n265_0[1]),.din(w_dff_B_2ZFijG8y4_2));
	jspl jspl_w_n266_0(.douta(w_n266_0[0]),.doutb(w_n266_0[1]),.din(n266));
	jspl jspl_w_n267_0(.douta(w_n267_0[0]),.doutb(w_n267_0[1]),.din(w_dff_B_LhM19GdE6_2));
	jspl jspl_w_n268_0(.douta(w_n268_0[0]),.doutb(w_n268_0[1]),.din(n268));
	jspl jspl_w_n269_0(.douta(w_n269_0[0]),.doutb(w_n269_0[1]),.din(w_dff_B_DveKxQYH6_2));
	jspl jspl_w_n270_0(.douta(w_n270_0[0]),.doutb(w_n270_0[1]),.din(n270));
	jspl jspl_w_n271_0(.douta(w_dff_A_MysAQcee9_0),.doutb(w_n271_0[1]),.din(n271));
	jspl jspl_w_n272_0(.douta(w_n272_0[0]),.doutb(w_n272_0[1]),.din(n272));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_dff_A_dd2KuOew4_1),.din(n274));
	jspl jspl_w_n275_0(.douta(w_n275_0[0]),.doutb(w_n275_0[1]),.din(n275));
	jspl jspl_w_n277_0(.douta(w_dff_A_NzASmWdC1_0),.doutb(w_n277_0[1]),.din(n277));
	jspl jspl_w_n282_0(.douta(w_n282_0[0]),.doutb(w_n282_0[1]),.din(n282));
	jspl jspl_w_n283_0(.douta(w_dff_A_fWFkXRlH4_0),.doutb(w_n283_0[1]),.din(n283));
	jspl3 jspl3_w_n288_0(.douta(w_n288_0[0]),.doutb(w_n288_0[1]),.doutc(w_n288_0[2]),.din(n288));
	jspl jspl_w_n290_0(.douta(w_n290_0[0]),.doutb(w_n290_0[1]),.din(w_dff_B_9vo0u5m23_2));
	jspl jspl_w_n293_0(.douta(w_n293_0[0]),.doutb(w_n293_0[1]),.din(n293));
	jspl jspl_w_n295_0(.douta(w_n295_0[0]),.doutb(w_n295_0[1]),.din(w_dff_B_zfj2YvDS8_2));
	jspl jspl_w_n298_0(.douta(w_n298_0[0]),.doutb(w_n298_0[1]),.din(n298));
	jspl jspl_w_n300_0(.douta(w_n300_0[0]),.doutb(w_n300_0[1]),.din(w_dff_B_Fh9L8oXW3_2));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.din(n303));
	jspl jspl_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.din(w_dff_B_6rTgYPtY9_2));
	jspl jspl_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.din(n308));
	jspl jspl_w_n310_0(.douta(w_n310_0[0]),.doutb(w_n310_0[1]),.din(w_dff_B_Vr0RTiuP0_2));
	jspl jspl_w_n311_0(.douta(w_n311_0[0]),.doutb(w_n311_0[1]),.din(n311));
	jspl jspl_w_n313_0(.douta(w_n313_0[0]),.doutb(w_n313_0[1]),.din(n313));
	jspl3 jspl3_w_n314_0(.douta(w_dff_A_ahOAYgm48_0),.doutb(w_dff_A_N92C5aQQ8_1),.doutc(w_n314_0[2]),.din(n314));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl jspl_w_n317_0(.douta(w_n317_0[0]),.doutb(w_n317_0[1]),.din(n317));
	jspl jspl_w_n320_0(.douta(w_n320_0[0]),.doutb(w_n320_0[1]),.din(n320));
	jspl jspl_w_n321_0(.douta(w_n321_0[0]),.doutb(w_n321_0[1]),.din(w_dff_B_VPsceqs67_2));
	jspl jspl_w_n322_0(.douta(w_n322_0[0]),.doutb(w_n322_0[1]),.din(n322));
	jspl jspl_w_n323_0(.douta(w_n323_0[0]),.doutb(w_n323_0[1]),.din(w_dff_B_3l4SKcDE9_2));
	jspl jspl_w_n324_0(.douta(w_n324_0[0]),.doutb(w_n324_0[1]),.din(n324));
	jspl jspl_w_n325_0(.douta(w_n325_0[0]),.doutb(w_n325_0[1]),.din(w_dff_B_nj6Se62c5_2));
	jspl jspl_w_n326_0(.douta(w_n326_0[0]),.doutb(w_n326_0[1]),.din(n326));
	jspl jspl_w_n327_0(.douta(w_n327_0[0]),.doutb(w_n327_0[1]),.din(w_dff_B_3RE2EL7P0_2));
	jspl jspl_w_n328_0(.douta(w_n328_0[0]),.doutb(w_n328_0[1]),.din(n328));
	jspl jspl_w_n329_0(.douta(w_dff_A_QRKEAwBf9_0),.doutb(w_n329_0[1]),.din(n329));
	jspl jspl_w_n330_0(.douta(w_n330_0[0]),.doutb(w_n330_0[1]),.din(n330));
	jspl jspl_w_n332_0(.douta(w_n332_0[0]),.doutb(w_dff_A_ZBNkQBen1_1),.din(n332));
	jspl jspl_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.din(n333));
	jspl jspl_w_n335_0(.douta(w_dff_A_KQ2O2otq9_0),.doutb(w_n335_0[1]),.din(n335));
	jspl jspl_w_n340_0(.douta(w_n340_0[0]),.doutb(w_n340_0[1]),.din(n340));
	jspl jspl_w_n341_0(.douta(w_dff_A_4O2bYNf23_0),.doutb(w_n341_0[1]),.din(n341));
	jspl3 jspl3_w_n346_0(.douta(w_n346_0[0]),.doutb(w_n346_0[1]),.doutc(w_n346_0[2]),.din(n346));
	jspl jspl_w_n348_0(.douta(w_n348_0[0]),.doutb(w_n348_0[1]),.din(w_dff_B_o72n8RB88_2));
	jspl jspl_w_n351_0(.douta(w_n351_0[0]),.doutb(w_n351_0[1]),.din(n351));
	jspl jspl_w_n353_0(.douta(w_n353_0[0]),.doutb(w_n353_0[1]),.din(w_dff_B_odjSL4HC4_2));
	jspl jspl_w_n356_0(.douta(w_n356_0[0]),.doutb(w_n356_0[1]),.din(n356));
	jspl jspl_w_n358_0(.douta(w_n358_0[0]),.doutb(w_n358_0[1]),.din(w_dff_B_z3z38aMv1_2));
	jspl jspl_w_n361_0(.douta(w_n361_0[0]),.doutb(w_n361_0[1]),.din(n361));
	jspl jspl_w_n363_0(.douta(w_n363_0[0]),.doutb(w_n363_0[1]),.din(w_dff_B_21WflzzA2_2));
	jspl jspl_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.din(n366));
	jspl jspl_w_n368_0(.douta(w_n368_0[0]),.doutb(w_n368_0[1]),.din(w_dff_B_BeecgaRi2_2));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(n371));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_dff_A_evwGOEkL4_1),.din(n372));
	jspl jspl_w_n373_0(.douta(w_n373_0[0]),.doutb(w_n373_0[1]),.din(n373));
	jspl jspl_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.din(n375));
	jspl3 jspl3_w_n376_0(.douta(w_dff_A_xQ8IgenW8_0),.doutb(w_dff_A_xriyLzyx7_1),.doutc(w_n376_0[2]),.din(n376));
	jspl jspl_w_n377_0(.douta(w_n377_0[0]),.doutb(w_n377_0[1]),.din(n377));
	jspl jspl_w_n380_0(.douta(w_dff_A_wYtxhkNR9_0),.doutb(w_n380_0[1]),.din(n380));
	jspl jspl_w_n382_0(.douta(w_n382_0[0]),.doutb(w_n382_0[1]),.din(n382));
	jspl jspl_w_n383_0(.douta(w_n383_0[0]),.doutb(w_n383_0[1]),.din(n383));
	jspl jspl_w_n384_0(.douta(w_n384_0[0]),.doutb(w_n384_0[1]),.din(n384));
	jspl jspl_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.din(w_dff_B_hGv4qMwx9_2));
	jspl jspl_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.din(n386));
	jspl jspl_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.din(w_dff_B_mh08k7Jk4_2));
	jspl jspl_w_n388_0(.douta(w_n388_0[0]),.doutb(w_n388_0[1]),.din(n388));
	jspl jspl_w_n389_0(.douta(w_n389_0[0]),.doutb(w_n389_0[1]),.din(w_dff_B_CqLjs5BL4_2));
	jspl jspl_w_n390_0(.douta(w_n390_0[0]),.doutb(w_n390_0[1]),.din(n390));
	jspl jspl_w_n391_0(.douta(w_n391_0[0]),.doutb(w_n391_0[1]),.din(w_dff_B_ce9XI3zW7_2));
	jspl jspl_w_n392_0(.douta(w_n392_0[0]),.doutb(w_n392_0[1]),.din(n392));
	jspl jspl_w_n393_0(.douta(w_dff_A_f6dTGFVx1_0),.doutb(w_n393_0[1]),.din(n393));
	jspl jspl_w_n394_0(.douta(w_n394_0[0]),.doutb(w_n394_0[1]),.din(n394));
	jspl jspl_w_n396_0(.douta(w_n396_0[0]),.doutb(w_dff_A_pdtZY1cb0_1),.din(n396));
	jspl jspl_w_n397_0(.douta(w_n397_0[0]),.doutb(w_n397_0[1]),.din(n397));
	jspl jspl_w_n399_0(.douta(w_dff_A_R4ZeTc807_0),.doutb(w_n399_0[1]),.din(n399));
	jspl jspl_w_n404_0(.douta(w_n404_0[0]),.doutb(w_n404_0[1]),.din(n404));
	jspl jspl_w_n405_0(.douta(w_dff_A_ymql107S1_0),.doutb(w_n405_0[1]),.din(n405));
	jspl3 jspl3_w_n410_0(.douta(w_n410_0[0]),.doutb(w_n410_0[1]),.doutc(w_n410_0[2]),.din(n410));
	jspl jspl_w_n412_0(.douta(w_n412_0[0]),.doutb(w_n412_0[1]),.din(w_dff_B_m3egyPwj4_2));
	jspl jspl_w_n415_0(.douta(w_n415_0[0]),.doutb(w_n415_0[1]),.din(n415));
	jspl jspl_w_n417_0(.douta(w_n417_0[0]),.doutb(w_n417_0[1]),.din(w_dff_B_NH7vxheQ8_2));
	jspl jspl_w_n420_0(.douta(w_n420_0[0]),.doutb(w_n420_0[1]),.din(n420));
	jspl jspl_w_n422_0(.douta(w_n422_0[0]),.doutb(w_n422_0[1]),.din(w_dff_B_DMYriVf68_2));
	jspl jspl_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.din(n425));
	jspl jspl_w_n427_0(.douta(w_n427_0[0]),.doutb(w_n427_0[1]),.din(w_dff_B_7NIX7gzS4_2));
	jspl jspl_w_n430_0(.douta(w_n430_0[0]),.doutb(w_n430_0[1]),.din(n430));
	jspl jspl_w_n432_0(.douta(w_n432_0[0]),.doutb(w_n432_0[1]),.din(w_dff_B_mcltNOjw8_2));
	jspl jspl_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.din(w_dff_B_qWfI2QVG8_2));
	jspl jspl_w_n437_0(.douta(w_n437_0[0]),.doutb(w_n437_0[1]),.din(w_dff_B_45LVaV9I9_2));
	jspl jspl_w_n441_0(.douta(w_n441_0[0]),.doutb(w_n441_0[1]),.din(n441));
	jspl jspl_w_n442_0(.douta(w_n442_0[0]),.doutb(w_dff_A_BbMEquCd0_1),.din(n442));
	jspl jspl_w_n443_0(.douta(w_n443_0[0]),.doutb(w_n443_0[1]),.din(n443));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl3 jspl3_w_n446_0(.douta(w_dff_A_B9LfuwoA9_0),.doutb(w_dff_A_KPFWeGym0_1),.doutc(w_n446_0[2]),.din(n446));
	jspl jspl_w_n447_0(.douta(w_n447_0[0]),.doutb(w_n447_0[1]),.din(n447));
	jspl jspl_w_n450_0(.douta(w_dff_A_PLejDV5i4_0),.doutb(w_n450_0[1]),.din(n450));
	jspl jspl_w_n452_0(.douta(w_n452_0[0]),.doutb(w_n452_0[1]),.din(n452));
	jspl jspl_w_n453_0(.douta(w_n453_0[0]),.doutb(w_n453_0[1]),.din(w_dff_B_lYkQHvFO0_2));
	jspl jspl_w_n454_0(.douta(w_n454_0[0]),.doutb(w_n454_0[1]),.din(n454));
	jspl jspl_w_n455_0(.douta(w_n455_0[0]),.doutb(w_n455_0[1]),.din(n455));
	jspl jspl_w_n456_0(.douta(w_n456_0[0]),.doutb(w_n456_0[1]),.din(n456));
	jspl jspl_w_n457_0(.douta(w_n457_0[0]),.doutb(w_n457_0[1]),.din(n457));
	jspl jspl_w_n458_0(.douta(w_n458_0[0]),.doutb(w_n458_0[1]),.din(n458));
	jspl jspl_w_n459_0(.douta(w_n459_0[0]),.doutb(w_n459_0[1]),.din(w_dff_B_99G06CEw4_2));
	jspl jspl_w_n460_0(.douta(w_n460_0[0]),.doutb(w_n460_0[1]),.din(n460));
	jspl jspl_w_n461_0(.douta(w_n461_0[0]),.doutb(w_n461_0[1]),.din(w_dff_B_PUBqbE3j7_2));
	jspl jspl_w_n462_0(.douta(w_n462_0[0]),.doutb(w_n462_0[1]),.din(n462));
	jspl jspl_w_n463_0(.douta(w_n463_0[0]),.doutb(w_n463_0[1]),.din(w_dff_B_A822Pj3E2_2));
	jspl jspl_w_n464_0(.douta(w_n464_0[0]),.doutb(w_n464_0[1]),.din(n464));
	jspl jspl_w_n465_0(.douta(w_dff_A_14eYYD6s0_0),.doutb(w_n465_0[1]),.din(n465));
	jspl jspl_w_n466_0(.douta(w_n466_0[0]),.doutb(w_n466_0[1]),.din(n466));
	jspl jspl_w_n468_0(.douta(w_n468_0[0]),.doutb(w_dff_A_q8tDLDGG5_1),.din(n468));
	jspl jspl_w_n469_0(.douta(w_n469_0[0]),.doutb(w_n469_0[1]),.din(n469));
	jspl jspl_w_n471_0(.douta(w_dff_A_YKx6JKpo5_0),.doutb(w_n471_0[1]),.din(n471));
	jspl jspl_w_n476_0(.douta(w_n476_0[0]),.doutb(w_n476_0[1]),.din(n476));
	jspl jspl_w_n477_0(.douta(w_dff_A_VqxSOFmS0_0),.doutb(w_n477_0[1]),.din(n477));
	jspl3 jspl3_w_n482_0(.douta(w_n482_0[0]),.doutb(w_n482_0[1]),.doutc(w_n482_0[2]),.din(n482));
	jspl jspl_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.din(w_dff_B_CCND9ubK0_2));
	jspl jspl_w_n487_0(.douta(w_n487_0[0]),.doutb(w_n487_0[1]),.din(n487));
	jspl jspl_w_n489_0(.douta(w_n489_0[0]),.doutb(w_n489_0[1]),.din(w_dff_B_lXtCB2Gg5_2));
	jspl jspl_w_n492_0(.douta(w_n492_0[0]),.doutb(w_n492_0[1]),.din(n492));
	jspl jspl_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.din(w_dff_B_6D0AnOxI9_2));
	jspl jspl_w_n497_0(.douta(w_n497_0[0]),.doutb(w_n497_0[1]),.din(n497));
	jspl jspl_w_n499_0(.douta(w_n499_0[0]),.doutb(w_n499_0[1]),.din(w_dff_B_En3EkI4x6_2));
	jspl jspl_w_n502_0(.douta(w_n502_0[0]),.doutb(w_n502_0[1]),.din(n502));
	jspl jspl_w_n504_0(.douta(w_n504_0[0]),.doutb(w_n504_0[1]),.din(w_dff_B_teV2fcSQ9_2));
	jspl jspl_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.din(n507));
	jspl jspl_w_n509_0(.douta(w_n509_0[0]),.doutb(w_n509_0[1]),.din(w_dff_B_FoTdDfnG1_2));
	jspl jspl_w_n512_0(.douta(w_n512_0[0]),.doutb(w_n512_0[1]),.din(n512));
	jspl jspl_w_n514_0(.douta(w_n514_0[0]),.doutb(w_n514_0[1]),.din(w_dff_B_aESPuByd0_2));
	jspl jspl_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.din(n518));
	jspl jspl_w_n519_0(.douta(w_n519_0[0]),.doutb(w_dff_A_fhhOmcMR1_1),.din(n519));
	jspl jspl_w_n520_0(.douta(w_n520_0[0]),.doutb(w_n520_0[1]),.din(n520));
	jspl jspl_w_n522_0(.douta(w_n522_0[0]),.doutb(w_n522_0[1]),.din(n522));
	jspl3 jspl3_w_n523_0(.douta(w_dff_A_dGQ0nULC2_0),.doutb(w_dff_A_KSo3umKP5_1),.doutc(w_n523_0[2]),.din(n523));
	jspl jspl_w_n524_0(.douta(w_n524_0[0]),.doutb(w_n524_0[1]),.din(n524));
	jspl jspl_w_n527_0(.douta(w_dff_A_FLv3uGPk2_0),.doutb(w_n527_0[1]),.din(n527));
	jspl jspl_w_n529_0(.douta(w_n529_0[0]),.doutb(w_n529_0[1]),.din(n529));
	jspl jspl_w_n530_0(.douta(w_n530_0[0]),.doutb(w_n530_0[1]),.din(w_dff_B_0jqNEiRK1_2));
	jspl jspl_w_n531_0(.douta(w_n531_0[0]),.doutb(w_n531_0[1]),.din(n531));
	jspl jspl_w_n532_0(.douta(w_n532_0[0]),.doutb(w_n532_0[1]),.din(w_dff_B_HiolJOlV9_2));
	jspl jspl_w_n533_0(.douta(w_n533_0[0]),.doutb(w_n533_0[1]),.din(n533));
	jspl jspl_w_n534_0(.douta(w_n534_0[0]),.doutb(w_n534_0[1]),.din(n534));
	jspl jspl_w_n535_0(.douta(w_n535_0[0]),.doutb(w_n535_0[1]),.din(n535));
	jspl jspl_w_n536_0(.douta(w_n536_0[0]),.doutb(w_n536_0[1]),.din(n536));
	jspl jspl_w_n537_0(.douta(w_n537_0[0]),.doutb(w_n537_0[1]),.din(n537));
	jspl jspl_w_n538_0(.douta(w_n538_0[0]),.doutb(w_n538_0[1]),.din(w_dff_B_60jCzz1X6_2));
	jspl jspl_w_n539_0(.douta(w_n539_0[0]),.doutb(w_n539_0[1]),.din(n539));
	jspl jspl_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.din(w_dff_B_y0jHMrmq7_2));
	jspl jspl_w_n541_0(.douta(w_n541_0[0]),.doutb(w_n541_0[1]),.din(n541));
	jspl jspl_w_n542_0(.douta(w_n542_0[0]),.doutb(w_n542_0[1]),.din(w_dff_B_WcIQi2vz7_2));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_n543_0[1]),.din(n543));
	jspl jspl_w_n544_0(.douta(w_dff_A_2N5I4kY78_0),.doutb(w_n544_0[1]),.din(n544));
	jspl jspl_w_n545_0(.douta(w_n545_0[0]),.doutb(w_n545_0[1]),.din(n545));
	jspl jspl_w_n547_0(.douta(w_n547_0[0]),.doutb(w_dff_A_J8sheeoS5_1),.din(n547));
	jspl jspl_w_n548_0(.douta(w_n548_0[0]),.doutb(w_n548_0[1]),.din(n548));
	jspl jspl_w_n550_0(.douta(w_dff_A_aYONlrSn6_0),.doutb(w_n550_0[1]),.din(n550));
	jspl jspl_w_n555_0(.douta(w_n555_0[0]),.doutb(w_n555_0[1]),.din(n555));
	jspl jspl_w_n556_0(.douta(w_dff_A_Jpe6BBw50_0),.doutb(w_n556_0[1]),.din(n556));
	jspl3 jspl3_w_n561_0(.douta(w_n561_0[0]),.doutb(w_n561_0[1]),.doutc(w_n561_0[2]),.din(n561));
	jspl jspl_w_n563_0(.douta(w_n563_0[0]),.doutb(w_n563_0[1]),.din(w_dff_B_S0rXoPdI4_2));
	jspl jspl_w_n566_0(.douta(w_n566_0[0]),.doutb(w_n566_0[1]),.din(n566));
	jspl jspl_w_n568_0(.douta(w_n568_0[0]),.doutb(w_n568_0[1]),.din(w_dff_B_w04eOjon8_2));
	jspl jspl_w_n571_0(.douta(w_n571_0[0]),.doutb(w_n571_0[1]),.din(n571));
	jspl jspl_w_n573_0(.douta(w_n573_0[0]),.doutb(w_n573_0[1]),.din(w_dff_B_YtxsDGOU2_2));
	jspl jspl_w_n576_0(.douta(w_n576_0[0]),.doutb(w_n576_0[1]),.din(n576));
	jspl jspl_w_n578_0(.douta(w_n578_0[0]),.doutb(w_n578_0[1]),.din(w_dff_B_36Zt8hAt2_2));
	jspl jspl_w_n581_0(.douta(w_n581_0[0]),.doutb(w_n581_0[1]),.din(n581));
	jspl jspl_w_n583_0(.douta(w_n583_0[0]),.doutb(w_n583_0[1]),.din(w_dff_B_FnvGQ8Bn4_2));
	jspl jspl_w_n586_0(.douta(w_n586_0[0]),.doutb(w_n586_0[1]),.din(n586));
	jspl jspl_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.din(w_dff_B_8pJGz1xv6_2));
	jspl jspl_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.din(n591));
	jspl jspl_w_n593_0(.douta(w_n593_0[0]),.doutb(w_n593_0[1]),.din(w_dff_B_T57MD6st6_2));
	jspl jspl_w_n596_0(.douta(w_n596_0[0]),.doutb(w_n596_0[1]),.din(n596));
	jspl jspl_w_n598_0(.douta(w_n598_0[0]),.doutb(w_n598_0[1]),.din(w_dff_B_aiLqEprQ5_2));
	jspl jspl_w_n602_0(.douta(w_n602_0[0]),.doutb(w_n602_0[1]),.din(n602));
	jspl jspl_w_n603_0(.douta(w_n603_0[0]),.doutb(w_dff_A_zum0rnsQ5_1),.din(n603));
	jspl jspl_w_n604_0(.douta(w_n604_0[0]),.doutb(w_n604_0[1]),.din(n604));
	jspl jspl_w_n606_0(.douta(w_n606_0[0]),.doutb(w_n606_0[1]),.din(n606));
	jspl3 jspl3_w_n607_0(.douta(w_dff_A_vN8Ty6XF4_0),.doutb(w_dff_A_srnRvMnm4_1),.doutc(w_n607_0[2]),.din(n607));
	jspl jspl_w_n608_0(.douta(w_n608_0[0]),.doutb(w_n608_0[1]),.din(n608));
	jspl jspl_w_n611_0(.douta(w_dff_A_uWveNDfc0_0),.doutb(w_n611_0[1]),.din(n611));
	jspl jspl_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.din(n613));
	jspl jspl_w_n614_0(.douta(w_n614_0[0]),.doutb(w_n614_0[1]),.din(w_dff_B_2FQMyY2l4_2));
	jspl jspl_w_n615_0(.douta(w_n615_0[0]),.doutb(w_n615_0[1]),.din(n615));
	jspl jspl_w_n616_0(.douta(w_n616_0[0]),.doutb(w_n616_0[1]),.din(w_dff_B_HPEZ81tM1_2));
	jspl jspl_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.din(n617));
	jspl jspl_w_n618_0(.douta(w_n618_0[0]),.doutb(w_n618_0[1]),.din(w_dff_B_hOcmHsaa3_2));
	jspl jspl_w_n619_0(.douta(w_n619_0[0]),.doutb(w_n619_0[1]),.din(n619));
	jspl jspl_w_n620_0(.douta(w_n620_0[0]),.doutb(w_n620_0[1]),.din(n620));
	jspl jspl_w_n621_0(.douta(w_n621_0[0]),.doutb(w_n621_0[1]),.din(n621));
	jspl jspl_w_n622_0(.douta(w_n622_0[0]),.doutb(w_n622_0[1]),.din(n622));
	jspl jspl_w_n623_0(.douta(w_n623_0[0]),.doutb(w_n623_0[1]),.din(n623));
	jspl jspl_w_n624_0(.douta(w_n624_0[0]),.doutb(w_n624_0[1]),.din(w_dff_B_smBEFrpg5_2));
	jspl jspl_w_n625_0(.douta(w_n625_0[0]),.doutb(w_n625_0[1]),.din(n625));
	jspl jspl_w_n626_0(.douta(w_n626_0[0]),.doutb(w_n626_0[1]),.din(w_dff_B_TPz8dDkP1_2));
	jspl jspl_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.din(n627));
	jspl jspl_w_n628_0(.douta(w_n628_0[0]),.doutb(w_n628_0[1]),.din(w_dff_B_9FCmbrcm4_2));
	jspl jspl_w_n629_0(.douta(w_n629_0[0]),.doutb(w_n629_0[1]),.din(n629));
	jspl jspl_w_n630_0(.douta(w_dff_A_XG0hYoUi2_0),.doutb(w_n630_0[1]),.din(n630));
	jspl jspl_w_n631_0(.douta(w_n631_0[0]),.doutb(w_n631_0[1]),.din(n631));
	jspl jspl_w_n633_0(.douta(w_n633_0[0]),.doutb(w_dff_A_XitmDLyL7_1),.din(n633));
	jspl jspl_w_n634_0(.douta(w_n634_0[0]),.doutb(w_n634_0[1]),.din(n634));
	jspl jspl_w_n636_0(.douta(w_dff_A_evevrTmx4_0),.doutb(w_n636_0[1]),.din(n636));
	jspl jspl_w_n641_0(.douta(w_n641_0[0]),.doutb(w_n641_0[1]),.din(n641));
	jspl jspl_w_n642_0(.douta(w_dff_A_KkeADDaJ8_0),.doutb(w_n642_0[1]),.din(n642));
	jspl3 jspl3_w_n647_0(.douta(w_n647_0[0]),.doutb(w_n647_0[1]),.doutc(w_n647_0[2]),.din(n647));
	jspl jspl_w_n649_0(.douta(w_n649_0[0]),.doutb(w_n649_0[1]),.din(w_dff_B_53epCT4a7_2));
	jspl jspl_w_n652_0(.douta(w_n652_0[0]),.doutb(w_n652_0[1]),.din(n652));
	jspl jspl_w_n654_0(.douta(w_n654_0[0]),.doutb(w_n654_0[1]),.din(w_dff_B_za3ROloz1_2));
	jspl jspl_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.din(n657));
	jspl jspl_w_n659_0(.douta(w_n659_0[0]),.doutb(w_n659_0[1]),.din(w_dff_B_2n9qfHGe5_2));
	jspl jspl_w_n662_0(.douta(w_n662_0[0]),.doutb(w_n662_0[1]),.din(n662));
	jspl jspl_w_n664_0(.douta(w_n664_0[0]),.doutb(w_n664_0[1]),.din(w_dff_B_aetrGM480_2));
	jspl jspl_w_n667_0(.douta(w_n667_0[0]),.doutb(w_n667_0[1]),.din(n667));
	jspl jspl_w_n669_0(.douta(w_n669_0[0]),.doutb(w_n669_0[1]),.din(w_dff_B_gvaO9FrA4_2));
	jspl jspl_w_n672_0(.douta(w_n672_0[0]),.doutb(w_n672_0[1]),.din(n672));
	jspl jspl_w_n674_0(.douta(w_n674_0[0]),.doutb(w_n674_0[1]),.din(w_dff_B_CsMAmuPH7_2));
	jspl jspl_w_n677_0(.douta(w_n677_0[0]),.doutb(w_n677_0[1]),.din(n677));
	jspl jspl_w_n679_0(.douta(w_n679_0[0]),.doutb(w_n679_0[1]),.din(w_dff_B_RJPkQgDR3_2));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.din(n682));
	jspl jspl_w_n684_0(.douta(w_n684_0[0]),.doutb(w_n684_0[1]),.din(w_dff_B_1XoMUMZI6_2));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_n687_0[1]),.din(n687));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(w_dff_B_kW0xO70A7_2));
	jspl jspl_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.din(n693));
	jspl jspl_w_n694_0(.douta(w_n694_0[0]),.doutb(w_dff_A_04uEiypF3_1),.din(n694));
	jspl3 jspl3_w_n695_0(.douta(w_dff_A_reLcFVwy2_0),.doutb(w_n695_0[1]),.doutc(w_n695_0[2]),.din(n695));
	jspl jspl_w_n697_0(.douta(w_n697_0[0]),.doutb(w_n697_0[1]),.din(n697));
	jspl3 jspl3_w_n698_0(.douta(w_dff_A_xi5AQlVt6_0),.doutb(w_dff_A_UfhNzngE2_1),.doutc(w_n698_0[2]),.din(n698));
	jspl jspl_w_n699_0(.douta(w_n699_0[0]),.doutb(w_n699_0[1]),.din(n699));
	jspl jspl_w_n702_0(.douta(w_dff_A_sw2PtKtX2_0),.doutb(w_n702_0[1]),.din(n702));
	jspl jspl_w_n704_0(.douta(w_n704_0[0]),.doutb(w_n704_0[1]),.din(n704));
	jspl jspl_w_n705_0(.douta(w_n705_0[0]),.doutb(w_n705_0[1]),.din(w_dff_B_Q9usjkEE9_2));
	jspl jspl_w_n706_0(.douta(w_n706_0[0]),.doutb(w_n706_0[1]),.din(n706));
	jspl jspl_w_n707_0(.douta(w_n707_0[0]),.doutb(w_n707_0[1]),.din(w_dff_B_3ZxVpABO3_2));
	jspl jspl_w_n708_0(.douta(w_n708_0[0]),.doutb(w_n708_0[1]),.din(n708));
	jspl jspl_w_n709_0(.douta(w_n709_0[0]),.doutb(w_n709_0[1]),.din(w_dff_B_hrRlyOSk0_2));
	jspl jspl_w_n710_0(.douta(w_n710_0[0]),.doutb(w_n710_0[1]),.din(n710));
	jspl jspl_w_n711_0(.douta(w_n711_0[0]),.doutb(w_n711_0[1]),.din(w_dff_B_TlpexhRO4_2));
	jspl jspl_w_n712_0(.douta(w_n712_0[0]),.doutb(w_n712_0[1]),.din(n712));
	jspl jspl_w_n713_0(.douta(w_n713_0[0]),.doutb(w_n713_0[1]),.din(n713));
	jspl jspl_w_n714_0(.douta(w_n714_0[0]),.doutb(w_n714_0[1]),.din(n714));
	jspl jspl_w_n715_0(.douta(w_n715_0[0]),.doutb(w_n715_0[1]),.din(n715));
	jspl jspl_w_n716_0(.douta(w_n716_0[0]),.doutb(w_n716_0[1]),.din(n716));
	jspl jspl_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.din(w_dff_B_Jf9q3FuV5_2));
	jspl jspl_w_n718_0(.douta(w_n718_0[0]),.doutb(w_n718_0[1]),.din(n718));
	jspl jspl_w_n719_0(.douta(w_n719_0[0]),.doutb(w_n719_0[1]),.din(w_dff_B_fkjO06sJ2_2));
	jspl jspl_w_n720_0(.douta(w_n720_0[0]),.doutb(w_n720_0[1]),.din(n720));
	jspl jspl_w_n721_0(.douta(w_n721_0[0]),.doutb(w_n721_0[1]),.din(w_dff_B_ZBEN2qtH8_2));
	jspl jspl_w_n722_0(.douta(w_n722_0[0]),.doutb(w_n722_0[1]),.din(n722));
	jspl jspl_w_n723_0(.douta(w_dff_A_TUptm82n2_0),.doutb(w_n723_0[1]),.din(n723));
	jspl jspl_w_n724_0(.douta(w_n724_0[0]),.doutb(w_n724_0[1]),.din(n724));
	jspl jspl_w_n726_0(.douta(w_n726_0[0]),.doutb(w_dff_A_90iIDhbQ1_1),.din(n726));
	jspl jspl_w_n727_0(.douta(w_n727_0[0]),.doutb(w_n727_0[1]),.din(n727));
	jspl jspl_w_n729_0(.douta(w_dff_A_v4PrTfen7_0),.doutb(w_n729_0[1]),.din(n729));
	jspl jspl_w_n734_0(.douta(w_n734_0[0]),.doutb(w_n734_0[1]),.din(n734));
	jspl jspl_w_n735_0(.douta(w_dff_A_gv2XXJR31_0),.doutb(w_n735_0[1]),.din(n735));
	jspl3 jspl3_w_n740_0(.douta(w_n740_0[0]),.doutb(w_n740_0[1]),.doutc(w_n740_0[2]),.din(n740));
	jspl jspl_w_n742_0(.douta(w_n742_0[0]),.doutb(w_n742_0[1]),.din(w_dff_B_XHgoh4ZN7_2));
	jspl jspl_w_n745_0(.douta(w_n745_0[0]),.doutb(w_n745_0[1]),.din(n745));
	jspl jspl_w_n747_0(.douta(w_n747_0[0]),.doutb(w_n747_0[1]),.din(w_dff_B_MZeffkU02_2));
	jspl jspl_w_n750_0(.douta(w_n750_0[0]),.doutb(w_n750_0[1]),.din(n750));
	jspl jspl_w_n752_0(.douta(w_n752_0[0]),.doutb(w_n752_0[1]),.din(w_dff_B_vREFlxaq6_2));
	jspl jspl_w_n755_0(.douta(w_n755_0[0]),.doutb(w_n755_0[1]),.din(n755));
	jspl jspl_w_n757_0(.douta(w_n757_0[0]),.doutb(w_n757_0[1]),.din(w_dff_B_kRNE0XN38_2));
	jspl jspl_w_n760_0(.douta(w_n760_0[0]),.doutb(w_n760_0[1]),.din(n760));
	jspl jspl_w_n762_0(.douta(w_n762_0[0]),.doutb(w_n762_0[1]),.din(w_dff_B_ZHXhiKye4_2));
	jspl jspl_w_n765_0(.douta(w_n765_0[0]),.doutb(w_n765_0[1]),.din(n765));
	jspl jspl_w_n767_0(.douta(w_n767_0[0]),.doutb(w_n767_0[1]),.din(w_dff_B_AjlORad90_2));
	jspl jspl_w_n770_0(.douta(w_n770_0[0]),.doutb(w_n770_0[1]),.din(n770));
	jspl jspl_w_n772_0(.douta(w_n772_0[0]),.doutb(w_n772_0[1]),.din(w_dff_B_IgHq9uxs3_2));
	jspl jspl_w_n775_0(.douta(w_n775_0[0]),.doutb(w_n775_0[1]),.din(n775));
	jspl jspl_w_n777_0(.douta(w_n777_0[0]),.doutb(w_n777_0[1]),.din(w_dff_B_e9sc4Qcq2_2));
	jspl jspl_w_n780_0(.douta(w_n780_0[0]),.doutb(w_n780_0[1]),.din(n780));
	jspl jspl_w_n782_0(.douta(w_n782_0[0]),.doutb(w_n782_0[1]),.din(w_dff_B_qZbZfeDP3_2));
	jspl jspl_w_n785_0(.douta(w_n785_0[0]),.doutb(w_n785_0[1]),.din(n785));
	jspl jspl_w_n787_0(.douta(w_n787_0[0]),.doutb(w_n787_0[1]),.din(w_dff_B_eylds8PW2_2));
	jspl jspl_w_n791_0(.douta(w_n791_0[0]),.doutb(w_n791_0[1]),.din(n791));
	jspl jspl_w_n792_0(.douta(w_n792_0[0]),.doutb(w_dff_A_AW1PADH56_1),.din(n792));
	jspl jspl_w_n793_0(.douta(w_dff_A_SZgnYqYp9_0),.doutb(w_n793_0[1]),.din(n793));
	jspl jspl_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.din(n795));
	jspl3 jspl3_w_n797_0(.douta(w_n797_0[0]),.doutb(w_n797_0[1]),.doutc(w_n797_0[2]),.din(n797));
	jspl jspl_w_n800_0(.douta(w_dff_A_gsSunOMy6_0),.doutb(w_n800_0[1]),.din(n800));
	jspl jspl_w_n802_0(.douta(w_n802_0[0]),.doutb(w_n802_0[1]),.din(n802));
	jspl jspl_w_n803_0(.douta(w_n803_0[0]),.doutb(w_n803_0[1]),.din(w_dff_B_yseD4T131_2));
	jspl jspl_w_n804_0(.douta(w_n804_0[0]),.doutb(w_n804_0[1]),.din(n804));
	jspl jspl_w_n805_0(.douta(w_n805_0[0]),.doutb(w_n805_0[1]),.din(w_dff_B_fwDr6czM6_2));
	jspl jspl_w_n806_0(.douta(w_n806_0[0]),.doutb(w_n806_0[1]),.din(n806));
	jspl jspl_w_n807_0(.douta(w_n807_0[0]),.doutb(w_n807_0[1]),.din(w_dff_B_3AHQoFUj2_2));
	jspl jspl_w_n808_0(.douta(w_n808_0[0]),.doutb(w_n808_0[1]),.din(n808));
	jspl jspl_w_n809_0(.douta(w_n809_0[0]),.doutb(w_n809_0[1]),.din(w_dff_B_Z9zB7At31_2));
	jspl jspl_w_n810_0(.douta(w_n810_0[0]),.doutb(w_n810_0[1]),.din(n810));
	jspl jspl_w_n811_0(.douta(w_n811_0[0]),.doutb(w_n811_0[1]),.din(w_dff_B_wXnEFDJP0_2));
	jspl jspl_w_n812_0(.douta(w_n812_0[0]),.doutb(w_n812_0[1]),.din(n812));
	jspl jspl_w_n813_0(.douta(w_n813_0[0]),.doutb(w_n813_0[1]),.din(n813));
	jspl jspl_w_n814_0(.douta(w_n814_0[0]),.doutb(w_n814_0[1]),.din(n814));
	jspl jspl_w_n815_0(.douta(w_n815_0[0]),.doutb(w_n815_0[1]),.din(n815));
	jspl jspl_w_n816_0(.douta(w_n816_0[0]),.doutb(w_n816_0[1]),.din(n816));
	jspl jspl_w_n817_0(.douta(w_n817_0[0]),.doutb(w_n817_0[1]),.din(w_dff_B_6ugO9nhT4_2));
	jspl jspl_w_n818_0(.douta(w_n818_0[0]),.doutb(w_n818_0[1]),.din(n818));
	jspl jspl_w_n819_0(.douta(w_n819_0[0]),.doutb(w_n819_0[1]),.din(w_dff_B_NrvwmNJd9_2));
	jspl jspl_w_n820_0(.douta(w_n820_0[0]),.doutb(w_n820_0[1]),.din(n820));
	jspl jspl_w_n821_0(.douta(w_n821_0[0]),.doutb(w_n821_0[1]),.din(w_dff_B_xlzt7Jp13_2));
	jspl jspl_w_n822_0(.douta(w_n822_0[0]),.doutb(w_n822_0[1]),.din(n822));
	jspl jspl_w_n823_0(.douta(w_dff_A_pNJ353jV9_0),.doutb(w_n823_0[1]),.din(n823));
	jspl jspl_w_n824_0(.douta(w_n824_0[0]),.doutb(w_n824_0[1]),.din(n824));
	jspl jspl_w_n826_0(.douta(w_n826_0[0]),.doutb(w_dff_A_ls7XPJqC5_1),.din(n826));
	jspl jspl_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.din(n827));
	jspl jspl_w_n829_0(.douta(w_dff_A_UeowzV526_0),.doutb(w_n829_0[1]),.din(n829));
	jspl jspl_w_n834_0(.douta(w_n834_0[0]),.doutb(w_n834_0[1]),.din(n834));
	jspl jspl_w_n835_0(.douta(w_n835_0[0]),.doutb(w_n835_0[1]),.din(w_dff_B_AQetBEn90_2));
	jspl jspl_w_n839_0(.douta(w_n839_0[0]),.doutb(w_n839_0[1]),.din(n839));
	jspl jspl_w_n840_0(.douta(w_dff_A_rddEyTe76_0),.doutb(w_n840_0[1]),.din(n840));
	jspl3 jspl3_w_n844_0(.douta(w_n844_0[0]),.doutb(w_n844_0[1]),.doutc(w_n844_0[2]),.din(n844));
	jspl jspl_w_n846_0(.douta(w_n846_0[0]),.doutb(w_n846_0[1]),.din(w_dff_B_oW3OI4Cm9_2));
	jspl jspl_w_n849_0(.douta(w_n849_0[0]),.doutb(w_n849_0[1]),.din(n849));
	jspl jspl_w_n851_0(.douta(w_n851_0[0]),.doutb(w_n851_0[1]),.din(w_dff_B_FvJ5VlAH2_2));
	jspl jspl_w_n854_0(.douta(w_n854_0[0]),.doutb(w_n854_0[1]),.din(n854));
	jspl jspl_w_n856_0(.douta(w_n856_0[0]),.doutb(w_n856_0[1]),.din(w_dff_B_lyf6aRnj3_2));
	jspl jspl_w_n859_0(.douta(w_n859_0[0]),.doutb(w_n859_0[1]),.din(n859));
	jspl jspl_w_n861_0(.douta(w_n861_0[0]),.doutb(w_n861_0[1]),.din(w_dff_B_OIsxnejw5_2));
	jspl jspl_w_n864_0(.douta(w_n864_0[0]),.doutb(w_n864_0[1]),.din(n864));
	jspl jspl_w_n866_0(.douta(w_n866_0[0]),.doutb(w_n866_0[1]),.din(w_dff_B_krEo57156_2));
	jspl jspl_w_n869_0(.douta(w_n869_0[0]),.doutb(w_n869_0[1]),.din(n869));
	jspl jspl_w_n871_0(.douta(w_n871_0[0]),.doutb(w_n871_0[1]),.din(w_dff_B_6nbRevOp8_2));
	jspl jspl_w_n874_0(.douta(w_n874_0[0]),.doutb(w_n874_0[1]),.din(n874));
	jspl jspl_w_n876_0(.douta(w_n876_0[0]),.doutb(w_n876_0[1]),.din(w_dff_B_TXHiw2xj9_2));
	jspl jspl_w_n879_0(.douta(w_n879_0[0]),.doutb(w_n879_0[1]),.din(n879));
	jspl jspl_w_n881_0(.douta(w_n881_0[0]),.doutb(w_n881_0[1]),.din(w_dff_B_hZonOQGc3_2));
	jspl jspl_w_n884_0(.douta(w_n884_0[0]),.doutb(w_n884_0[1]),.din(n884));
	jspl jspl_w_n886_0(.douta(w_n886_0[0]),.doutb(w_n886_0[1]),.din(w_dff_B_0l63gjYM2_2));
	jspl jspl_w_n889_0(.douta(w_n889_0[0]),.doutb(w_n889_0[1]),.din(n889));
	jspl jspl_w_n891_0(.douta(w_n891_0[0]),.doutb(w_n891_0[1]),.din(w_dff_B_l1f4Eccm7_2));
	jspl jspl_w_n895_0(.douta(w_n895_0[0]),.doutb(w_n895_0[1]),.din(n895));
	jspl jspl_w_n896_0(.douta(w_n896_0[0]),.doutb(w_dff_A_8hSQ65zN0_1),.din(n896));
	jspl jspl_w_n897_0(.douta(w_n897_0[0]),.doutb(w_n897_0[1]),.din(n897));
	jspl jspl_w_n898_0(.douta(w_n898_0[0]),.doutb(w_n898_0[1]),.din(w_dff_B_9nAcROIB4_2));
	jspl jspl_w_n901_0(.douta(w_n901_0[0]),.doutb(w_n901_0[1]),.din(n901));
	jspl jspl_w_n903_0(.douta(w_dff_A_YjJMEe3C2_0),.doutb(w_n903_0[1]),.din(n903));
	jspl jspl_w_n906_0(.douta(w_n906_0[0]),.doutb(w_n906_0[1]),.din(n906));
	jspl jspl_w_n907_0(.douta(w_n907_0[0]),.doutb(w_n907_0[1]),.din(w_dff_B_RKXxBQcS6_2));
	jspl jspl_w_n908_0(.douta(w_n908_0[0]),.doutb(w_n908_0[1]),.din(n908));
	jspl jspl_w_n909_0(.douta(w_n909_0[0]),.doutb(w_n909_0[1]),.din(w_dff_B_FMIx6HkA4_2));
	jspl jspl_w_n910_0(.douta(w_n910_0[0]),.doutb(w_n910_0[1]),.din(n910));
	jspl jspl_w_n911_0(.douta(w_n911_0[0]),.doutb(w_n911_0[1]),.din(w_dff_B_VPqAJya48_2));
	jspl jspl_w_n912_0(.douta(w_n912_0[0]),.doutb(w_n912_0[1]),.din(n912));
	jspl jspl_w_n913_0(.douta(w_n913_0[0]),.doutb(w_n913_0[1]),.din(w_dff_B_C2tPhRZm2_2));
	jspl jspl_w_n914_0(.douta(w_n914_0[0]),.doutb(w_n914_0[1]),.din(n914));
	jspl jspl_w_n915_0(.douta(w_n915_0[0]),.doutb(w_n915_0[1]),.din(w_dff_B_4QWmYAAQ7_2));
	jspl jspl_w_n916_0(.douta(w_n916_0[0]),.doutb(w_n916_0[1]),.din(n916));
	jspl jspl_w_n917_0(.douta(w_n917_0[0]),.doutb(w_n917_0[1]),.din(w_dff_B_KJRKARdL5_2));
	jspl jspl_w_n918_0(.douta(w_n918_0[0]),.doutb(w_n918_0[1]),.din(n918));
	jspl jspl_w_n919_0(.douta(w_n919_0[0]),.doutb(w_n919_0[1]),.din(n919));
	jspl jspl_w_n920_0(.douta(w_n920_0[0]),.doutb(w_n920_0[1]),.din(n920));
	jspl jspl_w_n921_0(.douta(w_n921_0[0]),.doutb(w_n921_0[1]),.din(n921));
	jspl jspl_w_n922_0(.douta(w_n922_0[0]),.doutb(w_n922_0[1]),.din(n922));
	jspl jspl_w_n923_0(.douta(w_n923_0[0]),.doutb(w_n923_0[1]),.din(w_dff_B_r0eWN7pX6_2));
	jspl jspl_w_n924_0(.douta(w_n924_0[0]),.doutb(w_n924_0[1]),.din(n924));
	jspl jspl_w_n925_0(.douta(w_n925_0[0]),.doutb(w_n925_0[1]),.din(w_dff_B_k1sYNB9t6_2));
	jspl jspl_w_n926_0(.douta(w_n926_0[0]),.doutb(w_n926_0[1]),.din(n926));
	jspl3 jspl3_w_n927_0(.douta(w_n927_0[0]),.doutb(w_dff_A_wALpsxUl8_1),.doutc(w_dff_A_9OrlJGK70_2),.din(n927));
	jspl jspl_w_n929_0(.douta(w_n929_0[0]),.doutb(w_dff_A_cONBtyJ46_1),.din(n929));
	jspl jspl_w_n930_0(.douta(w_n930_0[0]),.doutb(w_n930_0[1]),.din(n930));
	jspl jspl_w_n931_0(.douta(w_n931_0[0]),.doutb(w_dff_A_hQoEVyXq2_1),.din(n931));
	jspl jspl_w_n932_0(.douta(w_n932_0[0]),.doutb(w_n932_0[1]),.din(n932));
	jspl jspl_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.din(n937));
	jspl jspl_w_n938_0(.douta(w_n938_0[0]),.doutb(w_n938_0[1]),.din(w_dff_B_wKqaqs3V7_2));
	jspl3 jspl3_w_n942_0(.douta(w_n942_0[0]),.doutb(w_n942_0[1]),.doutc(w_n942_0[2]),.din(n942));
	jspl jspl_w_n943_0(.douta(w_n943_0[0]),.doutb(w_n943_0[1]),.din(w_dff_B_YoBgo9Qz8_2));
	jspl jspl_w_n949_0(.douta(w_n949_0[0]),.doutb(w_n949_0[1]),.din(n949));
	jspl jspl_w_n951_0(.douta(w_n951_0[0]),.doutb(w_n951_0[1]),.din(w_dff_B_NQ7tOS5e6_2));
	jspl jspl_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.din(n954));
	jspl jspl_w_n956_0(.douta(w_n956_0[0]),.doutb(w_n956_0[1]),.din(w_dff_B_65svk5wf5_2));
	jspl jspl_w_n959_0(.douta(w_n959_0[0]),.doutb(w_n959_0[1]),.din(n959));
	jspl jspl_w_n961_0(.douta(w_n961_0[0]),.doutb(w_n961_0[1]),.din(w_dff_B_9hb6a1Uh9_2));
	jspl jspl_w_n964_0(.douta(w_n964_0[0]),.doutb(w_n964_0[1]),.din(n964));
	jspl jspl_w_n966_0(.douta(w_n966_0[0]),.doutb(w_n966_0[1]),.din(w_dff_B_JKhRRn0h9_2));
	jspl jspl_w_n969_0(.douta(w_n969_0[0]),.doutb(w_n969_0[1]),.din(n969));
	jspl jspl_w_n971_0(.douta(w_n971_0[0]),.doutb(w_n971_0[1]),.din(w_dff_B_0GgBGg4k2_2));
	jspl jspl_w_n974_0(.douta(w_n974_0[0]),.doutb(w_n974_0[1]),.din(n974));
	jspl jspl_w_n976_0(.douta(w_n976_0[0]),.doutb(w_n976_0[1]),.din(w_dff_B_5gsdl4R01_2));
	jspl jspl_w_n979_0(.douta(w_n979_0[0]),.doutb(w_n979_0[1]),.din(n979));
	jspl jspl_w_n981_0(.douta(w_n981_0[0]),.doutb(w_n981_0[1]),.din(w_dff_B_L1lMMz1t6_2));
	jspl jspl_w_n984_0(.douta(w_n984_0[0]),.doutb(w_n984_0[1]),.din(n984));
	jspl jspl_w_n986_0(.douta(w_n986_0[0]),.doutb(w_n986_0[1]),.din(w_dff_B_SYNboMum6_2));
	jspl jspl_w_n989_0(.douta(w_n989_0[0]),.doutb(w_n989_0[1]),.din(n989));
	jspl jspl_w_n991_0(.douta(w_n991_0[0]),.doutb(w_n991_0[1]),.din(w_dff_B_8iNnw4fd3_2));
	jspl jspl_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.din(n994));
	jspl jspl_w_n996_0(.douta(w_n996_0[0]),.doutb(w_n996_0[1]),.din(w_dff_B_chRGbMx43_2));
	jspl jspl_w_n999_0(.douta(w_n999_0[0]),.doutb(w_n999_0[1]),.din(n999));
	jspl jspl_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.din(w_dff_B_N8ucdRpL4_2));
	jspl jspl_w_n1005_0(.douta(w_n1005_0[0]),.doutb(w_n1005_0[1]),.din(n1005));
	jspl jspl_w_n1006_0(.douta(w_n1006_0[0]),.doutb(w_dff_A_RxpTO1Zh9_1),.din(n1006));
	jspl jspl_w_n1008_0(.douta(w_dff_A_8xMT58BS1_0),.doutb(w_n1008_0[1]),.din(n1008));
	jspl jspl_w_n1009_0(.douta(w_n1009_0[0]),.doutb(w_n1009_0[1]),.din(n1009));
	jspl jspl_w_n1010_0(.douta(w_n1010_0[0]),.doutb(w_n1010_0[1]),.din(w_dff_B_l45lPUQS4_2));
	jspl jspl_w_n1011_0(.douta(w_n1011_0[0]),.doutb(w_n1011_0[1]),.din(n1011));
	jspl jspl_w_n1012_0(.douta(w_n1012_0[0]),.doutb(w_n1012_0[1]),.din(w_dff_B_wXiLleDA8_2));
	jspl jspl_w_n1013_0(.douta(w_n1013_0[0]),.doutb(w_n1013_0[1]),.din(n1013));
	jspl jspl_w_n1014_0(.douta(w_n1014_0[0]),.doutb(w_n1014_0[1]),.din(w_dff_B_dUlgKmam6_2));
	jspl jspl_w_n1015_0(.douta(w_n1015_0[0]),.doutb(w_n1015_0[1]),.din(n1015));
	jspl jspl_w_n1016_0(.douta(w_n1016_0[0]),.doutb(w_n1016_0[1]),.din(w_dff_B_xixEthtw6_2));
	jspl jspl_w_n1017_0(.douta(w_n1017_0[0]),.doutb(w_n1017_0[1]),.din(n1017));
	jspl jspl_w_n1018_0(.douta(w_n1018_0[0]),.doutb(w_n1018_0[1]),.din(w_dff_B_TUzQBg6C0_2));
	jspl jspl_w_n1019_0(.douta(w_n1019_0[0]),.doutb(w_n1019_0[1]),.din(n1019));
	jspl jspl_w_n1020_0(.douta(w_n1020_0[0]),.doutb(w_n1020_0[1]),.din(w_dff_B_CuRktE837_2));
	jspl jspl_w_n1021_0(.douta(w_n1021_0[0]),.doutb(w_n1021_0[1]),.din(n1021));
	jspl jspl_w_n1022_0(.douta(w_n1022_0[0]),.doutb(w_n1022_0[1]),.din(w_dff_B_zSTRPc7K1_2));
	jspl jspl_w_n1023_0(.douta(w_n1023_0[0]),.doutb(w_n1023_0[1]),.din(n1023));
	jspl jspl_w_n1024_0(.douta(w_n1024_0[0]),.doutb(w_n1024_0[1]),.din(n1024));
	jspl jspl_w_n1025_0(.douta(w_n1025_0[0]),.doutb(w_n1025_0[1]),.din(n1025));
	jspl jspl_w_n1026_0(.douta(w_n1026_0[0]),.doutb(w_n1026_0[1]),.din(n1026));
	jspl jspl_w_n1027_0(.douta(w_n1027_0[0]),.doutb(w_n1027_0[1]),.din(n1027));
	jspl jspl_w_n1028_0(.douta(w_n1028_0[0]),.doutb(w_n1028_0[1]),.din(w_dff_B_j5PCsBuH8_2));
	jspl jspl_w_n1029_0(.douta(w_n1029_0[0]),.doutb(w_n1029_0[1]),.din(n1029));
	jspl jspl_w_n1030_0(.douta(w_n1030_0[0]),.doutb(w_n1030_0[1]),.din(w_dff_B_7fn1wqLK1_2));
	jspl jspl_w_n1031_0(.douta(w_n1031_0[0]),.doutb(w_n1031_0[1]),.din(n1031));
	jspl jspl_w_n1032_0(.douta(w_n1032_0[0]),.doutb(w_dff_A_Voa2nWZi3_1),.din(n1032));
	jspl jspl_w_n1033_0(.douta(w_n1033_0[0]),.doutb(w_n1033_0[1]),.din(n1033));
	jspl jspl_w_n1034_0(.douta(w_dff_A_oCU1WYQG2_0),.doutb(w_n1034_0[1]),.din(n1034));
	jspl jspl_w_n1035_0(.douta(w_n1035_0[0]),.doutb(w_n1035_0[1]),.din(n1035));
	jspl jspl_w_n1037_0(.douta(w_n1037_0[0]),.doutb(w_n1037_0[1]),.din(w_dff_B_k77NgaMe2_2));
	jspl jspl_w_n1039_0(.douta(w_n1039_0[0]),.doutb(w_dff_A_hrBreWcA4_1),.din(n1039));
	jspl jspl_w_n1043_0(.douta(w_n1043_0[0]),.doutb(w_n1043_0[1]),.din(n1043));
	jspl jspl_w_n1044_0(.douta(w_n1044_0[0]),.doutb(w_n1044_0[1]),.din(w_dff_B_RMjRo5a85_2));
	jspl jspl_w_n1048_0(.douta(w_dff_A_Gr7HxICE1_0),.doutb(w_n1048_0[1]),.din(n1048));
	jspl jspl_w_n1049_0(.douta(w_n1049_0[0]),.doutb(w_n1049_0[1]),.din(w_dff_B_9Ia7o4WF4_2));
	jspl jspl_w_n1052_0(.douta(w_n1052_0[0]),.doutb(w_n1052_0[1]),.din(n1052));
	jspl jspl_w_n1054_0(.douta(w_n1054_0[0]),.doutb(w_n1054_0[1]),.din(w_dff_B_SPEl12Do8_2));
	jspl jspl_w_n1057_0(.douta(w_n1057_0[0]),.doutb(w_n1057_0[1]),.din(n1057));
	jspl jspl_w_n1059_0(.douta(w_n1059_0[0]),.doutb(w_n1059_0[1]),.din(w_dff_B_hezCouQL0_2));
	jspl jspl_w_n1062_0(.douta(w_n1062_0[0]),.doutb(w_n1062_0[1]),.din(n1062));
	jspl jspl_w_n1064_0(.douta(w_n1064_0[0]),.doutb(w_n1064_0[1]),.din(w_dff_B_NrD0JuhJ0_2));
	jspl jspl_w_n1067_0(.douta(w_n1067_0[0]),.doutb(w_n1067_0[1]),.din(n1067));
	jspl jspl_w_n1069_0(.douta(w_n1069_0[0]),.doutb(w_n1069_0[1]),.din(w_dff_B_GJjsYhnp3_2));
	jspl jspl_w_n1072_0(.douta(w_n1072_0[0]),.doutb(w_n1072_0[1]),.din(n1072));
	jspl jspl_w_n1074_0(.douta(w_n1074_0[0]),.doutb(w_n1074_0[1]),.din(w_dff_B_2OVZiyHD6_2));
	jspl jspl_w_n1077_0(.douta(w_n1077_0[0]),.doutb(w_n1077_0[1]),.din(n1077));
	jspl jspl_w_n1079_0(.douta(w_n1079_0[0]),.doutb(w_n1079_0[1]),.din(w_dff_B_RiuwrtiS3_2));
	jspl jspl_w_n1082_0(.douta(w_n1082_0[0]),.doutb(w_n1082_0[1]),.din(n1082));
	jspl jspl_w_n1084_0(.douta(w_n1084_0[0]),.doutb(w_n1084_0[1]),.din(w_dff_B_7bZcCXZS1_2));
	jspl jspl_w_n1087_0(.douta(w_n1087_0[0]),.doutb(w_n1087_0[1]),.din(n1087));
	jspl jspl_w_n1089_0(.douta(w_n1089_0[0]),.doutb(w_n1089_0[1]),.din(w_dff_B_79Wcx5u26_2));
	jspl jspl_w_n1092_0(.douta(w_n1092_0[0]),.doutb(w_n1092_0[1]),.din(n1092));
	jspl jspl_w_n1094_0(.douta(w_n1094_0[0]),.doutb(w_n1094_0[1]),.din(w_dff_B_Y8OjuYp30_2));
	jspl jspl_w_n1097_0(.douta(w_n1097_0[0]),.doutb(w_n1097_0[1]),.din(n1097));
	jspl jspl_w_n1099_0(.douta(w_n1099_0[0]),.doutb(w_n1099_0[1]),.din(w_dff_B_fsycHxs66_2));
	jspl jspl_w_n1102_0(.douta(w_n1102_0[0]),.doutb(w_n1102_0[1]),.din(n1102));
	jspl jspl_w_n1103_0(.douta(w_n1103_0[0]),.doutb(w_n1103_0[1]),.din(w_dff_B_jaHXtSYv4_2));
	jspl jspl_w_n1109_0(.douta(w_n1109_0[0]),.doutb(w_n1109_0[1]),.din(n1109));
	jspl jspl_w_n1110_0(.douta(w_dff_A_WmXhKVT75_0),.doutb(w_n1110_0[1]),.din(w_dff_B_qHewBVZt4_2));
	jspl jspl_w_n1114_0(.douta(w_n1114_0[0]),.doutb(w_n1114_0[1]),.din(n1114));
	jspl jspl_w_n1115_0(.douta(w_n1115_0[0]),.doutb(w_n1115_0[1]),.din(n1115));
	jspl jspl_w_n1116_0(.douta(w_n1116_0[0]),.doutb(w_n1116_0[1]),.din(n1116));
	jspl jspl_w_n1117_0(.douta(w_n1117_0[0]),.doutb(w_n1117_0[1]),.din(w_dff_B_bu33HQNV7_2));
	jspl jspl_w_n1118_0(.douta(w_n1118_0[0]),.doutb(w_n1118_0[1]),.din(n1118));
	jspl jspl_w_n1119_0(.douta(w_n1119_0[0]),.doutb(w_n1119_0[1]),.din(w_dff_B_MqZfHPqe4_2));
	jspl jspl_w_n1120_0(.douta(w_n1120_0[0]),.doutb(w_n1120_0[1]),.din(n1120));
	jspl jspl_w_n1121_0(.douta(w_n1121_0[0]),.doutb(w_n1121_0[1]),.din(w_dff_B_GbmpGLAX9_2));
	jspl jspl_w_n1122_0(.douta(w_n1122_0[0]),.doutb(w_n1122_0[1]),.din(n1122));
	jspl jspl_w_n1123_0(.douta(w_n1123_0[0]),.doutb(w_n1123_0[1]),.din(w_dff_B_CcpcWgtq1_2));
	jspl jspl_w_n1124_0(.douta(w_n1124_0[0]),.doutb(w_n1124_0[1]),.din(n1124));
	jspl jspl_w_n1125_0(.douta(w_n1125_0[0]),.doutb(w_n1125_0[1]),.din(w_dff_B_o0s09aK91_2));
	jspl jspl_w_n1126_0(.douta(w_n1126_0[0]),.doutb(w_n1126_0[1]),.din(n1126));
	jspl jspl_w_n1127_0(.douta(w_n1127_0[0]),.doutb(w_n1127_0[1]),.din(w_dff_B_kDDcdUhh8_2));
	jspl jspl_w_n1128_0(.douta(w_n1128_0[0]),.doutb(w_n1128_0[1]),.din(n1128));
	jspl jspl_w_n1129_0(.douta(w_n1129_0[0]),.doutb(w_n1129_0[1]),.din(n1129));
	jspl jspl_w_n1130_0(.douta(w_n1130_0[0]),.doutb(w_n1130_0[1]),.din(n1130));
	jspl jspl_w_n1131_0(.douta(w_n1131_0[0]),.doutb(w_n1131_0[1]),.din(n1131));
	jspl jspl_w_n1132_0(.douta(w_n1132_0[0]),.doutb(w_n1132_0[1]),.din(n1132));
	jspl jspl_w_n1133_0(.douta(w_n1133_0[0]),.doutb(w_n1133_0[1]),.din(w_dff_B_dwHvenCd1_2));
	jspl jspl_w_n1134_0(.douta(w_n1134_0[0]),.doutb(w_n1134_0[1]),.din(n1134));
	jspl jspl_w_n1135_0(.douta(w_n1135_0[0]),.doutb(w_n1135_0[1]),.din(w_dff_B_xK3sLJvh1_2));
	jspl jspl_w_n1137_0(.douta(w_n1137_0[0]),.doutb(w_n1137_0[1]),.din(n1137));
	jspl jspl_w_n1138_0(.douta(w_n1138_0[0]),.doutb(w_n1138_0[1]),.din(n1138));
	jspl jspl_w_n1139_0(.douta(w_n1139_0[0]),.doutb(w_n1139_0[1]),.din(n1139));
	jspl jspl_w_n1140_0(.douta(w_n1140_0[0]),.doutb(w_dff_A_ZxkjIyrc9_1),.din(n1140));
	jspl jspl_w_n1141_0(.douta(w_n1141_0[0]),.doutb(w_n1141_0[1]),.din(n1141));
	jspl jspl_w_n1147_0(.douta(w_n1147_0[0]),.doutb(w_n1147_0[1]),.din(n1147));
	jspl jspl_w_n1151_0(.douta(w_dff_A_NPQRlaQD6_0),.doutb(w_n1151_0[1]),.din(w_dff_B_QGHX3ctl8_2));
	jspl jspl_w_n1152_0(.douta(w_n1152_0[0]),.doutb(w_n1152_0[1]),.din(w_dff_B_Ycu9g66M0_2));
	jspl jspl_w_n1156_0(.douta(w_n1156_0[0]),.doutb(w_n1156_0[1]),.din(n1156));
	jspl jspl_w_n1158_0(.douta(w_n1158_0[0]),.doutb(w_n1158_0[1]),.din(w_dff_B_C1CopPj13_2));
	jspl jspl_w_n1161_0(.douta(w_n1161_0[0]),.doutb(w_n1161_0[1]),.din(n1161));
	jspl jspl_w_n1163_0(.douta(w_n1163_0[0]),.doutb(w_n1163_0[1]),.din(w_dff_B_8aqOsc927_2));
	jspl jspl_w_n1166_0(.douta(w_n1166_0[0]),.doutb(w_n1166_0[1]),.din(n1166));
	jspl jspl_w_n1168_0(.douta(w_n1168_0[0]),.doutb(w_n1168_0[1]),.din(w_dff_B_E2OoLQUy0_2));
	jspl jspl_w_n1171_0(.douta(w_n1171_0[0]),.doutb(w_n1171_0[1]),.din(n1171));
	jspl jspl_w_n1173_0(.douta(w_n1173_0[0]),.doutb(w_n1173_0[1]),.din(w_dff_B_j1oyz5BA5_2));
	jspl jspl_w_n1176_0(.douta(w_n1176_0[0]),.doutb(w_n1176_0[1]),.din(n1176));
	jspl jspl_w_n1178_0(.douta(w_n1178_0[0]),.doutb(w_n1178_0[1]),.din(w_dff_B_2l75t1df1_2));
	jspl jspl_w_n1181_0(.douta(w_n1181_0[0]),.doutb(w_n1181_0[1]),.din(n1181));
	jspl jspl_w_n1183_0(.douta(w_n1183_0[0]),.doutb(w_n1183_0[1]),.din(w_dff_B_UAI8SVqq1_2));
	jspl jspl_w_n1186_0(.douta(w_n1186_0[0]),.doutb(w_n1186_0[1]),.din(n1186));
	jspl jspl_w_n1188_0(.douta(w_n1188_0[0]),.doutb(w_n1188_0[1]),.din(w_dff_B_OX7pxmD05_2));
	jspl jspl_w_n1191_0(.douta(w_n1191_0[0]),.doutb(w_n1191_0[1]),.din(n1191));
	jspl jspl_w_n1193_0(.douta(w_n1193_0[0]),.doutb(w_n1193_0[1]),.din(w_dff_B_m6wpOOTX3_2));
	jspl jspl_w_n1196_0(.douta(w_n1196_0[0]),.doutb(w_n1196_0[1]),.din(n1196));
	jspl jspl_w_n1198_0(.douta(w_n1198_0[0]),.doutb(w_n1198_0[1]),.din(w_dff_B_5p8CRa7h9_2));
	jspl jspl_w_n1201_0(.douta(w_n1201_0[0]),.doutb(w_n1201_0[1]),.din(n1201));
	jspl jspl_w_n1203_0(.douta(w_n1203_0[0]),.doutb(w_n1203_0[1]),.din(w_dff_B_FD98udlP0_2));
	jspl jspl_w_n1206_0(.douta(w_n1206_0[0]),.doutb(w_n1206_0[1]),.din(w_dff_B_lu06mhQM1_2));
	jspl jspl_w_n1207_0(.douta(w_n1207_0[0]),.doutb(w_n1207_0[1]),.din(w_dff_B_fr1DhGc09_2));
	jspl jspl_w_n1208_0(.douta(w_n1208_0[0]),.doutb(w_n1208_0[1]),.din(w_dff_B_0sA4WOD92_2));
	jspl jspl_w_n1210_0(.douta(w_n1210_0[0]),.doutb(w_n1210_0[1]),.din(n1210));
	jspl jspl_w_n1212_0(.douta(w_n1212_0[0]),.doutb(w_n1212_0[1]),.din(n1212));
	jspl jspl_w_n1213_0(.douta(w_n1213_0[0]),.doutb(w_n1213_0[1]),.din(n1213));
	jspl jspl_w_n1214_0(.douta(w_n1214_0[0]),.doutb(w_n1214_0[1]),.din(n1214));
	jspl jspl_w_n1215_0(.douta(w_n1215_0[0]),.doutb(w_n1215_0[1]),.din(w_dff_B_vZPtaRWA8_2));
	jspl jspl_w_n1216_0(.douta(w_n1216_0[0]),.doutb(w_n1216_0[1]),.din(n1216));
	jspl jspl_w_n1217_0(.douta(w_n1217_0[0]),.doutb(w_n1217_0[1]),.din(w_dff_B_9cKVxRGY2_2));
	jspl jspl_w_n1218_0(.douta(w_n1218_0[0]),.doutb(w_n1218_0[1]),.din(n1218));
	jspl jspl_w_n1219_0(.douta(w_n1219_0[0]),.doutb(w_n1219_0[1]),.din(w_dff_B_D9ufeY0w9_2));
	jspl jspl_w_n1220_0(.douta(w_n1220_0[0]),.doutb(w_n1220_0[1]),.din(n1220));
	jspl jspl_w_n1221_0(.douta(w_n1221_0[0]),.doutb(w_n1221_0[1]),.din(w_dff_B_Z0a9KuK07_2));
	jspl jspl_w_n1222_0(.douta(w_n1222_0[0]),.doutb(w_n1222_0[1]),.din(n1222));
	jspl jspl_w_n1223_0(.douta(w_n1223_0[0]),.doutb(w_n1223_0[1]),.din(w_dff_B_06mQNvWb6_2));
	jspl jspl_w_n1224_0(.douta(w_n1224_0[0]),.doutb(w_n1224_0[1]),.din(n1224));
	jspl jspl_w_n1225_0(.douta(w_n1225_0[0]),.doutb(w_n1225_0[1]),.din(w_dff_B_9lJINcr55_2));
	jspl jspl_w_n1226_0(.douta(w_n1226_0[0]),.doutb(w_n1226_0[1]),.din(n1226));
	jspl jspl_w_n1227_0(.douta(w_n1227_0[0]),.doutb(w_n1227_0[1]),.din(n1227));
	jspl jspl_w_n1228_0(.douta(w_n1228_0[0]),.doutb(w_n1228_0[1]),.din(n1228));
	jspl jspl_w_n1229_0(.douta(w_n1229_0[0]),.doutb(w_n1229_0[1]),.din(n1229));
	jspl jspl_w_n1230_0(.douta(w_n1230_0[0]),.doutb(w_n1230_0[1]),.din(n1230));
	jspl jspl_w_n1231_0(.douta(w_n1231_0[0]),.doutb(w_n1231_0[1]),.din(w_dff_B_yl0l0a1u5_2));
	jspl jspl_w_n1232_0(.douta(w_n1232_0[0]),.doutb(w_n1232_0[1]),.din(n1232));
	jspl jspl_w_n1234_0(.douta(w_n1234_0[0]),.doutb(w_n1234_0[1]),.din(w_dff_B_DxnsUaBS1_2));
	jspl jspl_w_n1236_0(.douta(w_n1236_0[0]),.doutb(w_n1236_0[1]),.din(n1236));
	jspl jspl_w_n1237_0(.douta(w_n1237_0[0]),.doutb(w_n1237_0[1]),.din(n1237));
	jspl jspl_w_n1238_0(.douta(w_dff_A_3F2qeiCQ3_0),.doutb(w_n1238_0[1]),.din(n1238));
	jspl jspl_w_n1244_0(.douta(w_n1244_0[0]),.doutb(w_n1244_0[1]),.din(n1244));
	jspl jspl_w_n1247_0(.douta(w_n1247_0[0]),.doutb(w_n1247_0[1]),.din(n1247));
	jspl jspl_w_n1248_0(.douta(w_n1248_0[0]),.doutb(w_n1248_0[1]),.din(w_dff_B_TkXN03tm1_2));
	jspl jspl_w_n1251_0(.douta(w_n1251_0[0]),.doutb(w_n1251_0[1]),.din(n1251));
	jspl jspl_w_n1253_0(.douta(w_n1253_0[0]),.doutb(w_n1253_0[1]),.din(w_dff_B_ohmRqlak2_2));
	jspl jspl_w_n1256_0(.douta(w_n1256_0[0]),.doutb(w_n1256_0[1]),.din(n1256));
	jspl jspl_w_n1258_0(.douta(w_n1258_0[0]),.doutb(w_n1258_0[1]),.din(w_dff_B_jqkbv9TZ6_2));
	jspl jspl_w_n1261_0(.douta(w_n1261_0[0]),.doutb(w_n1261_0[1]),.din(n1261));
	jspl jspl_w_n1263_0(.douta(w_n1263_0[0]),.doutb(w_n1263_0[1]),.din(w_dff_B_xJ4lo3gy1_2));
	jspl jspl_w_n1266_0(.douta(w_n1266_0[0]),.doutb(w_n1266_0[1]),.din(n1266));
	jspl jspl_w_n1268_0(.douta(w_n1268_0[0]),.doutb(w_n1268_0[1]),.din(w_dff_B_20xgkSPY9_2));
	jspl jspl_w_n1271_0(.douta(w_n1271_0[0]),.doutb(w_n1271_0[1]),.din(n1271));
	jspl jspl_w_n1273_0(.douta(w_n1273_0[0]),.doutb(w_n1273_0[1]),.din(w_dff_B_w0rM8Gjh0_2));
	jspl jspl_w_n1276_0(.douta(w_n1276_0[0]),.doutb(w_n1276_0[1]),.din(n1276));
	jspl jspl_w_n1278_0(.douta(w_n1278_0[0]),.doutb(w_n1278_0[1]),.din(w_dff_B_rCZSACc71_2));
	jspl jspl_w_n1281_0(.douta(w_n1281_0[0]),.doutb(w_n1281_0[1]),.din(n1281));
	jspl jspl_w_n1283_0(.douta(w_n1283_0[0]),.doutb(w_n1283_0[1]),.din(w_dff_B_rYzcXI5W9_2));
	jspl jspl_w_n1286_0(.douta(w_n1286_0[0]),.doutb(w_n1286_0[1]),.din(n1286));
	jspl jspl_w_n1288_0(.douta(w_n1288_0[0]),.doutb(w_n1288_0[1]),.din(w_dff_B_GP9JAZhC8_2));
	jspl jspl_w_n1291_0(.douta(w_n1291_0[0]),.doutb(w_n1291_0[1]),.din(n1291));
	jspl jspl_w_n1293_0(.douta(w_n1293_0[0]),.doutb(w_n1293_0[1]),.din(w_dff_B_rOjuu2xq3_2));
	jspl jspl_w_n1296_0(.douta(w_n1296_0[0]),.doutb(w_n1296_0[1]),.din(w_dff_B_RvqdFM2d3_2));
	jspl jspl_w_n1297_0(.douta(w_n1297_0[0]),.doutb(w_n1297_0[1]),.din(w_dff_B_aWfsZ3VJ7_2));
	jspl jspl_w_n1298_0(.douta(w_n1298_0[0]),.doutb(w_n1298_0[1]),.din(w_dff_B_WTdmoGjV0_2));
	jspl jspl_w_n1301_0(.douta(w_n1301_0[0]),.doutb(w_n1301_0[1]),.din(n1301));
	jspl jspl_w_n1303_0(.douta(w_n1303_0[0]),.doutb(w_n1303_0[1]),.din(n1303));
	jspl jspl_w_n1304_0(.douta(w_n1304_0[0]),.doutb(w_n1304_0[1]),.din(n1304));
	jspl jspl_w_n1305_0(.douta(w_n1305_0[0]),.doutb(w_n1305_0[1]),.din(n1305));
	jspl jspl_w_n1306_0(.douta(w_n1306_0[0]),.doutb(w_n1306_0[1]),.din(n1306));
	jspl jspl_w_n1307_0(.douta(w_n1307_0[0]),.doutb(w_n1307_0[1]),.din(n1307));
	jspl jspl_w_n1308_0(.douta(w_n1308_0[0]),.doutb(w_n1308_0[1]),.din(w_dff_B_4LcJR0th3_2));
	jspl jspl_w_n1309_0(.douta(w_n1309_0[0]),.doutb(w_n1309_0[1]),.din(n1309));
	jspl jspl_w_n1310_0(.douta(w_n1310_0[0]),.doutb(w_n1310_0[1]),.din(w_dff_B_JzaWxUPK5_2));
	jspl jspl_w_n1311_0(.douta(w_n1311_0[0]),.doutb(w_n1311_0[1]),.din(n1311));
	jspl jspl_w_n1312_0(.douta(w_n1312_0[0]),.doutb(w_n1312_0[1]),.din(w_dff_B_rTBOuZFw4_2));
	jspl jspl_w_n1313_0(.douta(w_n1313_0[0]),.doutb(w_n1313_0[1]),.din(n1313));
	jspl jspl_w_n1314_0(.douta(w_n1314_0[0]),.doutb(w_n1314_0[1]),.din(w_dff_B_xSk7omfA1_2));
	jspl jspl_w_n1315_0(.douta(w_n1315_0[0]),.doutb(w_n1315_0[1]),.din(n1315));
	jspl jspl_w_n1316_0(.douta(w_n1316_0[0]),.doutb(w_n1316_0[1]),.din(w_dff_B_j4ccORpw4_2));
	jspl jspl_w_n1317_0(.douta(w_n1317_0[0]),.doutb(w_n1317_0[1]),.din(n1317));
	jspl jspl_w_n1318_0(.douta(w_n1318_0[0]),.doutb(w_n1318_0[1]),.din(n1318));
	jspl jspl_w_n1319_0(.douta(w_n1319_0[0]),.doutb(w_n1319_0[1]),.din(n1319));
	jspl jspl_w_n1320_0(.douta(w_n1320_0[0]),.doutb(w_n1320_0[1]),.din(n1320));
	jspl jspl_w_n1321_0(.douta(w_n1321_0[0]),.doutb(w_n1321_0[1]),.din(n1321));
	jspl jspl_w_n1322_0(.douta(w_n1322_0[0]),.doutb(w_dff_A_kYtAJoyj3_1),.din(n1322));
	jspl jspl_w_n1324_0(.douta(w_n1324_0[0]),.doutb(w_n1324_0[1]),.din(n1324));
	jspl jspl_w_n1325_0(.douta(w_n1325_0[0]),.doutb(w_dff_A_IPnXeFHN0_1),.din(n1325));
	jspl jspl_w_n1326_0(.douta(w_dff_A_GY0tRlvX7_0),.doutb(w_n1326_0[1]),.din(n1326));
	jspl jspl_w_n1332_0(.douta(w_n1332_0[0]),.doutb(w_n1332_0[1]),.din(n1332));
	jspl jspl_w_n1337_0(.douta(w_n1337_0[0]),.doutb(w_n1337_0[1]),.din(n1337));
	jspl jspl_w_n1338_0(.douta(w_n1338_0[0]),.doutb(w_n1338_0[1]),.din(w_dff_B_CAjFbE2G4_2));
	jspl jspl_w_n1341_0(.douta(w_n1341_0[0]),.doutb(w_n1341_0[1]),.din(n1341));
	jspl jspl_w_n1343_0(.douta(w_n1343_0[0]),.doutb(w_n1343_0[1]),.din(w_dff_B_y92mo1M43_2));
	jspl jspl_w_n1346_0(.douta(w_n1346_0[0]),.doutb(w_n1346_0[1]),.din(n1346));
	jspl jspl_w_n1348_0(.douta(w_n1348_0[0]),.doutb(w_n1348_0[1]),.din(w_dff_B_1mUiIhGD0_2));
	jspl jspl_w_n1351_0(.douta(w_n1351_0[0]),.doutb(w_n1351_0[1]),.din(n1351));
	jspl jspl_w_n1353_0(.douta(w_n1353_0[0]),.doutb(w_n1353_0[1]),.din(w_dff_B_Patk0o6B2_2));
	jspl jspl_w_n1356_0(.douta(w_n1356_0[0]),.doutb(w_n1356_0[1]),.din(n1356));
	jspl jspl_w_n1358_0(.douta(w_n1358_0[0]),.doutb(w_n1358_0[1]),.din(w_dff_B_ZKhslv1z7_2));
	jspl jspl_w_n1361_0(.douta(w_n1361_0[0]),.doutb(w_n1361_0[1]),.din(n1361));
	jspl jspl_w_n1363_0(.douta(w_n1363_0[0]),.doutb(w_n1363_0[1]),.din(w_dff_B_7yT6s86O9_2));
	jspl jspl_w_n1366_0(.douta(w_n1366_0[0]),.doutb(w_n1366_0[1]),.din(n1366));
	jspl jspl_w_n1368_0(.douta(w_n1368_0[0]),.doutb(w_n1368_0[1]),.din(w_dff_B_NOQOgkWw8_2));
	jspl jspl_w_n1371_0(.douta(w_n1371_0[0]),.doutb(w_n1371_0[1]),.din(n1371));
	jspl jspl_w_n1373_0(.douta(w_n1373_0[0]),.doutb(w_n1373_0[1]),.din(w_dff_B_XlOikqK90_2));
	jspl jspl_w_n1376_0(.douta(w_n1376_0[0]),.doutb(w_n1376_0[1]),.din(w_dff_B_TmNOlf9n0_2));
	jspl jspl_w_n1378_0(.douta(w_n1378_0[0]),.doutb(w_n1378_0[1]),.din(w_dff_B_N0Tsv9Tp0_2));
	jspl jspl_w_n1381_0(.douta(w_n1381_0[0]),.doutb(w_n1381_0[1]),.din(w_dff_B_mB60qQA78_2));
	jspl jspl_w_n1382_0(.douta(w_n1382_0[0]),.doutb(w_n1382_0[1]),.din(w_dff_B_lQleofwo6_2));
	jspl jspl_w_n1383_0(.douta(w_n1383_0[0]),.doutb(w_n1383_0[1]),.din(w_dff_B_Lwcvv2XE9_2));
	jspl jspl_w_n1386_0(.douta(w_n1386_0[0]),.doutb(w_n1386_0[1]),.din(n1386));
	jspl jspl_w_n1388_0(.douta(w_n1388_0[0]),.doutb(w_n1388_0[1]),.din(n1388));
	jspl jspl_w_n1389_0(.douta(w_n1389_0[0]),.doutb(w_n1389_0[1]),.din(n1389));
	jspl jspl_w_n1390_0(.douta(w_n1390_0[0]),.doutb(w_n1390_0[1]),.din(n1390));
	jspl jspl_w_n1391_0(.douta(w_n1391_0[0]),.doutb(w_n1391_0[1]),.din(n1391));
	jspl jspl_w_n1392_0(.douta(w_n1392_0[0]),.doutb(w_n1392_0[1]),.din(n1392));
	jspl jspl_w_n1393_0(.douta(w_n1393_0[0]),.doutb(w_n1393_0[1]),.din(n1393));
	jspl jspl_w_n1394_0(.douta(w_n1394_0[0]),.doutb(w_n1394_0[1]),.din(n1394));
	jspl jspl_w_n1395_0(.douta(w_n1395_0[0]),.doutb(w_n1395_0[1]),.din(w_dff_B_N7HFNmL51_2));
	jspl jspl_w_n1396_0(.douta(w_n1396_0[0]),.doutb(w_n1396_0[1]),.din(n1396));
	jspl jspl_w_n1397_0(.douta(w_n1397_0[0]),.doutb(w_n1397_0[1]),.din(w_dff_B_wETVknfo3_2));
	jspl jspl_w_n1398_0(.douta(w_n1398_0[0]),.doutb(w_n1398_0[1]),.din(n1398));
	jspl jspl_w_n1399_0(.douta(w_n1399_0[0]),.doutb(w_n1399_0[1]),.din(w_dff_B_PpKZCrKf2_2));
	jspl jspl_w_n1400_0(.douta(w_n1400_0[0]),.doutb(w_n1400_0[1]),.din(n1400));
	jspl jspl_w_n1401_0(.douta(w_n1401_0[0]),.doutb(w_n1401_0[1]),.din(w_dff_B_h43tcy7G1_2));
	jspl jspl_w_n1402_0(.douta(w_n1402_0[0]),.doutb(w_n1402_0[1]),.din(n1402));
	jspl jspl_w_n1403_0(.douta(w_n1403_0[0]),.doutb(w_n1403_0[1]),.din(n1403));
	jspl jspl_w_n1404_0(.douta(w_n1404_0[0]),.doutb(w_n1404_0[1]),.din(n1404));
	jspl jspl_w_n1405_0(.douta(w_n1405_0[0]),.doutb(w_n1405_0[1]),.din(n1405));
	jspl jspl_w_n1407_0(.douta(w_n1407_0[0]),.doutb(w_n1407_0[1]),.din(n1407));
	jspl jspl_w_n1409_0(.douta(w_n1409_0[0]),.doutb(w_n1409_0[1]),.din(n1409));
	jspl jspl_w_n1410_0(.douta(w_n1410_0[0]),.doutb(w_dff_A_vT4dEFkO3_1),.din(n1410));
	jspl jspl_w_n1415_0(.douta(w_n1415_0[0]),.doutb(w_n1415_0[1]),.din(n1415));
	jspl jspl_w_n1420_0(.douta(w_n1420_0[0]),.doutb(w_n1420_0[1]),.din(w_dff_B_16GkUzZv0_2));
	jspl jspl_w_n1421_0(.douta(w_n1421_0[0]),.doutb(w_n1421_0[1]),.din(w_dff_B_mHXheFJ27_2));
	jspl jspl_w_n1424_0(.douta(w_n1424_0[0]),.doutb(w_n1424_0[1]),.din(n1424));
	jspl jspl_w_n1426_0(.douta(w_n1426_0[0]),.doutb(w_n1426_0[1]),.din(w_dff_B_EZtOMoZi1_2));
	jspl jspl_w_n1429_0(.douta(w_n1429_0[0]),.doutb(w_n1429_0[1]),.din(n1429));
	jspl jspl_w_n1431_0(.douta(w_n1431_0[0]),.doutb(w_n1431_0[1]),.din(w_dff_B_xqaVoTr96_2));
	jspl jspl_w_n1434_0(.douta(w_n1434_0[0]),.doutb(w_n1434_0[1]),.din(n1434));
	jspl jspl_w_n1436_0(.douta(w_n1436_0[0]),.doutb(w_n1436_0[1]),.din(w_dff_B_apora1Ov2_2));
	jspl jspl_w_n1439_0(.douta(w_n1439_0[0]),.doutb(w_n1439_0[1]),.din(n1439));
	jspl jspl_w_n1441_0(.douta(w_n1441_0[0]),.doutb(w_n1441_0[1]),.din(w_dff_B_eriIFOdA8_2));
	jspl jspl_w_n1444_0(.douta(w_n1444_0[0]),.doutb(w_n1444_0[1]),.din(n1444));
	jspl jspl_w_n1446_0(.douta(w_n1446_0[0]),.doutb(w_n1446_0[1]),.din(w_dff_B_OaNem0ST0_2));
	jspl jspl_w_n1449_0(.douta(w_n1449_0[0]),.doutb(w_n1449_0[1]),.din(w_dff_B_72E2VBGY8_2));
	jspl jspl_w_n1451_0(.douta(w_n1451_0[0]),.doutb(w_n1451_0[1]),.din(w_dff_B_PgDjnd6z1_2));
	jspl jspl_w_n1454_0(.douta(w_n1454_0[0]),.doutb(w_n1454_0[1]),.din(w_dff_B_L7rgudxM0_2));
	jspl jspl_w_n1456_0(.douta(w_n1456_0[0]),.doutb(w_n1456_0[1]),.din(w_dff_B_cqr3P2Ay4_2));
	jspl jspl_w_n1459_0(.douta(w_n1459_0[0]),.doutb(w_n1459_0[1]),.din(w_dff_B_mAl5mvvM9_2));
	jspl jspl_w_n1460_0(.douta(w_n1460_0[0]),.doutb(w_n1460_0[1]),.din(w_dff_B_zZeO24ZO9_2));
	jspl jspl_w_n1461_0(.douta(w_n1461_0[0]),.doutb(w_n1461_0[1]),.din(w_dff_B_x0NmA8Gt4_2));
	jspl jspl_w_n1464_0(.douta(w_n1464_0[0]),.doutb(w_n1464_0[1]),.din(n1464));
	jspl jspl_w_n1466_0(.douta(w_n1466_0[0]),.doutb(w_n1466_0[1]),.din(n1466));
	jspl jspl_w_n1467_0(.douta(w_n1467_0[0]),.doutb(w_n1467_0[1]),.din(n1467));
	jspl jspl_w_n1468_0(.douta(w_n1468_0[0]),.doutb(w_n1468_0[1]),.din(n1468));
	jspl jspl_w_n1469_0(.douta(w_n1469_0[0]),.doutb(w_n1469_0[1]),.din(n1469));
	jspl jspl_w_n1470_0(.douta(w_n1470_0[0]),.doutb(w_n1470_0[1]),.din(n1470));
	jspl jspl_w_n1471_0(.douta(w_n1471_0[0]),.doutb(w_n1471_0[1]),.din(n1471));
	jspl jspl_w_n1472_0(.douta(w_n1472_0[0]),.doutb(w_n1472_0[1]),.din(n1472));
	jspl jspl_w_n1473_0(.douta(w_n1473_0[0]),.doutb(w_n1473_0[1]),.din(n1473));
	jspl jspl_w_n1474_0(.douta(w_n1474_0[0]),.doutb(w_n1474_0[1]),.din(n1474));
	jspl jspl_w_n1475_0(.douta(w_n1475_0[0]),.doutb(w_n1475_0[1]),.din(w_dff_B_Jmxx0iWk6_2));
	jspl jspl_w_n1476_0(.douta(w_n1476_0[0]),.doutb(w_n1476_0[1]),.din(n1476));
	jspl jspl_w_n1477_0(.douta(w_n1477_0[0]),.doutb(w_n1477_0[1]),.din(w_dff_B_gCURn5tp9_2));
	jspl jspl_w_n1478_0(.douta(w_n1478_0[0]),.doutb(w_n1478_0[1]),.din(n1478));
	jspl jspl_w_n1479_0(.douta(w_n1479_0[0]),.doutb(w_n1479_0[1]),.din(w_dff_B_tAhCEUVg1_2));
	jspl jspl_w_n1480_0(.douta(w_n1480_0[0]),.doutb(w_n1480_0[1]),.din(n1480));
	jspl jspl_w_n1481_0(.douta(w_n1481_0[0]),.doutb(w_n1481_0[1]),.din(n1481));
	jspl jspl_w_n1483_0(.douta(w_n1483_0[0]),.doutb(w_n1483_0[1]),.din(n1483));
	jspl jspl_w_n1485_0(.douta(w_n1485_0[0]),.doutb(w_n1485_0[1]),.din(n1485));
	jspl jspl_w_n1486_0(.douta(w_n1486_0[0]),.doutb(w_dff_A_njEHyu7l3_1),.din(n1486));
	jspl jspl_w_n1491_0(.douta(w_n1491_0[0]),.doutb(w_n1491_0[1]),.din(n1491));
	jspl jspl_w_n1496_0(.douta(w_n1496_0[0]),.doutb(w_n1496_0[1]),.din(w_dff_B_af4nwA5n9_2));
	jspl jspl_w_n1497_0(.douta(w_n1497_0[0]),.doutb(w_n1497_0[1]),.din(w_dff_B_tUghYg4N8_2));
	jspl jspl_w_n1500_0(.douta(w_n1500_0[0]),.doutb(w_n1500_0[1]),.din(n1500));
	jspl jspl_w_n1502_0(.douta(w_n1502_0[0]),.doutb(w_n1502_0[1]),.din(w_dff_B_TLbaPM3u0_2));
	jspl jspl_w_n1505_0(.douta(w_n1505_0[0]),.doutb(w_n1505_0[1]),.din(n1505));
	jspl jspl_w_n1507_0(.douta(w_n1507_0[0]),.doutb(w_n1507_0[1]),.din(w_dff_B_k7ju0uw85_2));
	jspl jspl_w_n1510_0(.douta(w_n1510_0[0]),.doutb(w_n1510_0[1]),.din(n1510));
	jspl jspl_w_n1512_0(.douta(w_n1512_0[0]),.doutb(w_n1512_0[1]),.din(w_dff_B_64mFQgHf1_2));
	jspl jspl_w_n1515_0(.douta(w_n1515_0[0]),.doutb(w_n1515_0[1]),.din(w_dff_B_a5IKWAgM2_2));
	jspl jspl_w_n1517_0(.douta(w_n1517_0[0]),.doutb(w_n1517_0[1]),.din(w_dff_B_fKPvmQG84_2));
	jspl jspl_w_n1520_0(.douta(w_n1520_0[0]),.doutb(w_n1520_0[1]),.din(w_dff_B_bkzLefRO7_2));
	jspl jspl_w_n1522_0(.douta(w_n1522_0[0]),.doutb(w_n1522_0[1]),.din(w_dff_B_8pMa8pGJ1_2));
	jspl jspl_w_n1525_0(.douta(w_n1525_0[0]),.doutb(w_n1525_0[1]),.din(w_dff_B_wZRVoe8d1_2));
	jspl jspl_w_n1527_0(.douta(w_n1527_0[0]),.doutb(w_n1527_0[1]),.din(w_dff_B_jdG9VyKO9_2));
	jspl jspl_w_n1530_0(.douta(w_n1530_0[0]),.doutb(w_n1530_0[1]),.din(w_dff_B_24k6eYsp4_2));
	jspl jspl_w_n1531_0(.douta(w_n1531_0[0]),.doutb(w_n1531_0[1]),.din(w_dff_B_irSCcU5R7_2));
	jspl jspl_w_n1532_0(.douta(w_n1532_0[0]),.doutb(w_n1532_0[1]),.din(w_dff_B_GkoW1heP5_2));
	jspl jspl_w_n1535_0(.douta(w_n1535_0[0]),.doutb(w_n1535_0[1]),.din(n1535));
	jspl jspl_w_n1537_0(.douta(w_n1537_0[0]),.doutb(w_n1537_0[1]),.din(n1537));
	jspl jspl_w_n1538_0(.douta(w_n1538_0[0]),.doutb(w_n1538_0[1]),.din(n1538));
	jspl jspl_w_n1539_0(.douta(w_n1539_0[0]),.doutb(w_n1539_0[1]),.din(n1539));
	jspl jspl_w_n1540_0(.douta(w_n1540_0[0]),.doutb(w_n1540_0[1]),.din(n1540));
	jspl jspl_w_n1541_0(.douta(w_n1541_0[0]),.doutb(w_n1541_0[1]),.din(n1541));
	jspl jspl_w_n1542_0(.douta(w_n1542_0[0]),.doutb(w_n1542_0[1]),.din(n1542));
	jspl jspl_w_n1543_0(.douta(w_n1543_0[0]),.doutb(w_n1543_0[1]),.din(n1543));
	jspl jspl_w_n1544_0(.douta(w_n1544_0[0]),.doutb(w_n1544_0[1]),.din(n1544));
	jspl jspl_w_n1545_0(.douta(w_n1545_0[0]),.doutb(w_n1545_0[1]),.din(n1545));
	jspl jspl_w_n1546_0(.douta(w_n1546_0[0]),.doutb(w_n1546_0[1]),.din(n1546));
	jspl jspl_w_n1547_0(.douta(w_n1547_0[0]),.doutb(w_n1547_0[1]),.din(n1547));
	jspl jspl_w_n1548_0(.douta(w_n1548_0[0]),.doutb(w_n1548_0[1]),.din(w_dff_B_OzTc8R7Z8_2));
	jspl jspl_w_n1549_0(.douta(w_n1549_0[0]),.doutb(w_n1549_0[1]),.din(n1549));
	jspl jspl_w_n1550_0(.douta(w_n1550_0[0]),.doutb(w_dff_A_F5DGNIku5_1),.din(n1550));
	jspl jspl_w_n1552_0(.douta(w_n1552_0[0]),.doutb(w_n1552_0[1]),.din(n1552));
	jspl jspl_w_n1554_0(.douta(w_n1554_0[0]),.doutb(w_n1554_0[1]),.din(n1554));
	jspl jspl_w_n1555_0(.douta(w_n1555_0[0]),.doutb(w_dff_A_xmslFCKQ7_1),.din(n1555));
	jspl jspl_w_n1560_0(.douta(w_n1560_0[0]),.doutb(w_n1560_0[1]),.din(n1560));
	jspl jspl_w_n1565_0(.douta(w_n1565_0[0]),.doutb(w_n1565_0[1]),.din(n1565));
	jspl jspl_w_n1566_0(.douta(w_n1566_0[0]),.doutb(w_n1566_0[1]),.din(w_dff_B_EVsqjVM83_2));
	jspl jspl_w_n1569_0(.douta(w_n1569_0[0]),.doutb(w_n1569_0[1]),.din(n1569));
	jspl jspl_w_n1571_0(.douta(w_n1571_0[0]),.doutb(w_n1571_0[1]),.din(w_dff_B_wG1Npweu9_2));
	jspl jspl_w_n1574_0(.douta(w_n1574_0[0]),.doutb(w_n1574_0[1]),.din(w_dff_B_Noqgof8s2_2));
	jspl jspl_w_n1576_0(.douta(w_n1576_0[0]),.doutb(w_n1576_0[1]),.din(w_dff_B_gEEO3E7I5_2));
	jspl jspl_w_n1579_0(.douta(w_n1579_0[0]),.doutb(w_n1579_0[1]),.din(w_dff_B_cPxo96Ll1_2));
	jspl jspl_w_n1581_0(.douta(w_n1581_0[0]),.doutb(w_n1581_0[1]),.din(w_dff_B_Vw0RU65l8_2));
	jspl jspl_w_n1584_0(.douta(w_n1584_0[0]),.doutb(w_n1584_0[1]),.din(w_dff_B_V4twCLF92_2));
	jspl jspl_w_n1586_0(.douta(w_n1586_0[0]),.doutb(w_n1586_0[1]),.din(w_dff_B_uxlbT8043_2));
	jspl jspl_w_n1589_0(.douta(w_n1589_0[0]),.doutb(w_n1589_0[1]),.din(w_dff_B_niD869Mu6_2));
	jspl jspl_w_n1591_0(.douta(w_n1591_0[0]),.doutb(w_n1591_0[1]),.din(w_dff_B_rdWGEVfD7_2));
	jspl jspl_w_n1594_0(.douta(w_n1594_0[0]),.doutb(w_n1594_0[1]),.din(w_dff_B_UnfEEObK3_2));
	jspl jspl_w_n1595_0(.douta(w_n1595_0[0]),.doutb(w_n1595_0[1]),.din(w_dff_B_kHchIEaa6_2));
	jspl jspl_w_n1596_0(.douta(w_n1596_0[0]),.doutb(w_n1596_0[1]),.din(w_dff_B_j3hSLS2j5_2));
	jspl jspl_w_n1599_0(.douta(w_n1599_0[0]),.doutb(w_n1599_0[1]),.din(n1599));
	jspl jspl_w_n1601_0(.douta(w_n1601_0[0]),.doutb(w_n1601_0[1]),.din(n1601));
	jspl jspl_w_n1602_0(.douta(w_n1602_0[0]),.doutb(w_n1602_0[1]),.din(n1602));
	jspl jspl_w_n1603_0(.douta(w_n1603_0[0]),.doutb(w_n1603_0[1]),.din(n1603));
	jspl jspl_w_n1604_0(.douta(w_n1604_0[0]),.doutb(w_n1604_0[1]),.din(n1604));
	jspl jspl_w_n1605_0(.douta(w_n1605_0[0]),.doutb(w_n1605_0[1]),.din(n1605));
	jspl jspl_w_n1606_0(.douta(w_n1606_0[0]),.doutb(w_n1606_0[1]),.din(n1606));
	jspl jspl_w_n1607_0(.douta(w_n1607_0[0]),.doutb(w_n1607_0[1]),.din(n1607));
	jspl jspl_w_n1608_0(.douta(w_n1608_0[0]),.doutb(w_n1608_0[1]),.din(n1608));
	jspl jspl_w_n1609_0(.douta(w_n1609_0[0]),.doutb(w_n1609_0[1]),.din(n1609));
	jspl jspl_w_n1610_0(.douta(w_n1610_0[0]),.doutb(w_n1610_0[1]),.din(n1610));
	jspl jspl_w_n1611_0(.douta(w_n1611_0[0]),.doutb(w_n1611_0[1]),.din(n1611));
	jspl jspl_w_n1612_0(.douta(w_n1612_0[0]),.doutb(w_n1612_0[1]),.din(n1612));
	jspl jspl_w_n1614_0(.douta(w_n1614_0[0]),.doutb(w_n1614_0[1]),.din(n1614));
	jspl jspl_w_n1616_0(.douta(w_n1616_0[0]),.doutb(w_n1616_0[1]),.din(n1616));
	jspl jspl_w_n1617_0(.douta(w_n1617_0[0]),.doutb(w_dff_A_9NTLJcnU8_1),.din(n1617));
	jspl jspl_w_n1622_0(.douta(w_n1622_0[0]),.doutb(w_n1622_0[1]),.din(n1622));
	jspl jspl_w_n1627_0(.douta(w_n1627_0[0]),.doutb(w_n1627_0[1]),.din(w_dff_B_DlNTa9EC7_2));
	jspl jspl_w_n1628_0(.douta(w_n1628_0[0]),.doutb(w_n1628_0[1]),.din(w_dff_B_Zcxv3EB42_2));
	jspl jspl_w_n1631_0(.douta(w_n1631_0[0]),.doutb(w_dff_A_zzjBz9dq1_1),.din(n1631));
	jspl jspl_w_n1633_0(.douta(w_n1633_0[0]),.doutb(w_n1633_0[1]),.din(w_dff_B_oltETmjT9_2));
	jspl jspl_w_n1636_0(.douta(w_n1636_0[0]),.doutb(w_n1636_0[1]),.din(w_dff_B_dpZfKvVX0_2));
	jspl jspl_w_n1638_0(.douta(w_n1638_0[0]),.doutb(w_n1638_0[1]),.din(w_dff_B_TbklrleN4_2));
	jspl jspl_w_n1641_0(.douta(w_n1641_0[0]),.doutb(w_n1641_0[1]),.din(w_dff_B_wvGEp2xp2_2));
	jspl jspl_w_n1643_0(.douta(w_n1643_0[0]),.doutb(w_n1643_0[1]),.din(w_dff_B_3rVbqRBO3_2));
	jspl jspl_w_n1646_0(.douta(w_n1646_0[0]),.doutb(w_n1646_0[1]),.din(w_dff_B_hHfKE0vn2_2));
	jspl jspl_w_n1648_0(.douta(w_n1648_0[0]),.doutb(w_n1648_0[1]),.din(w_dff_B_ICMzF6Jr6_2));
	jspl jspl_w_n1651_0(.douta(w_n1651_0[0]),.doutb(w_n1651_0[1]),.din(w_dff_B_7ewJLvDw1_2));
	jspl jspl_w_n1652_0(.douta(w_n1652_0[0]),.doutb(w_n1652_0[1]),.din(w_dff_B_O76LVzGe3_2));
	jspl jspl_w_n1653_0(.douta(w_n1653_0[0]),.doutb(w_n1653_0[1]),.din(w_dff_B_ef7mrUa07_2));
	jspl jspl_w_n1656_0(.douta(w_n1656_0[0]),.doutb(w_n1656_0[1]),.din(n1656));
	jspl jspl_w_n1658_0(.douta(w_n1658_0[0]),.doutb(w_n1658_0[1]),.din(n1658));
	jspl jspl_w_n1659_0(.douta(w_n1659_0[0]),.doutb(w_n1659_0[1]),.din(n1659));
	jspl jspl_w_n1660_0(.douta(w_n1660_0[0]),.doutb(w_n1660_0[1]),.din(n1660));
	jspl jspl_w_n1661_0(.douta(w_n1661_0[0]),.doutb(w_n1661_0[1]),.din(n1661));
	jspl jspl_w_n1662_0(.douta(w_n1662_0[0]),.doutb(w_n1662_0[1]),.din(n1662));
	jspl jspl_w_n1663_0(.douta(w_n1663_0[0]),.doutb(w_n1663_0[1]),.din(n1663));
	jspl jspl_w_n1664_0(.douta(w_n1664_0[0]),.doutb(w_n1664_0[1]),.din(n1664));
	jspl jspl_w_n1665_0(.douta(w_n1665_0[0]),.doutb(w_n1665_0[1]),.din(n1665));
	jspl jspl_w_n1666_0(.douta(w_n1666_0[0]),.doutb(w_n1666_0[1]),.din(n1666));
	jspl jspl_w_n1667_0(.douta(w_n1667_0[0]),.doutb(w_n1667_0[1]),.din(n1667));
	jspl jspl_w_n1669_0(.douta(w_n1669_0[0]),.doutb(w_n1669_0[1]),.din(n1669));
	jspl jspl_w_n1671_0(.douta(w_n1671_0[0]),.doutb(w_n1671_0[1]),.din(n1671));
	jspl jspl_w_n1672_0(.douta(w_n1672_0[0]),.doutb(w_dff_A_PseeWV7o8_1),.din(n1672));
	jspl jspl_w_n1677_0(.douta(w_n1677_0[0]),.doutb(w_n1677_0[1]),.din(n1677));
	jspl jspl_w_n1682_0(.douta(w_n1682_0[0]),.doutb(w_n1682_0[1]),.din(w_dff_B_HeUhQdQa6_2));
	jspl jspl_w_n1684_0(.douta(w_n1684_0[0]),.doutb(w_n1684_0[1]),.din(w_dff_B_eRWRvYFs0_2));
	jspl jspl_w_n1687_0(.douta(w_n1687_0[0]),.doutb(w_n1687_0[1]),.din(w_dff_B_vidOmM8E0_2));
	jspl jspl_w_n1689_0(.douta(w_n1689_0[0]),.doutb(w_n1689_0[1]),.din(w_dff_B_r7iq2aZb3_2));
	jspl jspl_w_n1692_0(.douta(w_n1692_0[0]),.doutb(w_n1692_0[1]),.din(w_dff_B_2HkC6nbC5_2));
	jspl jspl_w_n1694_0(.douta(w_n1694_0[0]),.doutb(w_n1694_0[1]),.din(w_dff_B_BGuYp3u05_2));
	jspl jspl_w_n1697_0(.douta(w_n1697_0[0]),.doutb(w_n1697_0[1]),.din(w_dff_B_7bx0Xb2Q0_2));
	jspl jspl_w_n1699_0(.douta(w_n1699_0[0]),.doutb(w_n1699_0[1]),.din(w_dff_B_Jq1IKcFg1_2));
	jspl jspl_w_n1702_0(.douta(w_n1702_0[0]),.doutb(w_n1702_0[1]),.din(w_dff_B_vpqxp1Kb7_2));
	jspl jspl_w_n1703_0(.douta(w_n1703_0[0]),.doutb(w_n1703_0[1]),.din(w_dff_B_PBFYhsH57_2));
	jspl jspl_w_n1704_0(.douta(w_n1704_0[0]),.doutb(w_n1704_0[1]),.din(w_dff_B_io3x0prC6_2));
	jspl jspl_w_n1707_0(.douta(w_n1707_0[0]),.doutb(w_n1707_0[1]),.din(n1707));
	jspl jspl_w_n1709_0(.douta(w_n1709_0[0]),.doutb(w_n1709_0[1]),.din(n1709));
	jspl jspl_w_n1710_0(.douta(w_n1710_0[0]),.doutb(w_n1710_0[1]),.din(n1710));
	jspl jspl_w_n1711_0(.douta(w_n1711_0[0]),.doutb(w_n1711_0[1]),.din(n1711));
	jspl jspl_w_n1712_0(.douta(w_n1712_0[0]),.doutb(w_n1712_0[1]),.din(n1712));
	jspl jspl_w_n1713_0(.douta(w_n1713_0[0]),.doutb(w_n1713_0[1]),.din(n1713));
	jspl jspl_w_n1714_0(.douta(w_n1714_0[0]),.doutb(w_n1714_0[1]),.din(n1714));
	jspl jspl_w_n1715_0(.douta(w_n1715_0[0]),.doutb(w_n1715_0[1]),.din(n1715));
	jspl jspl_w_n1716_0(.douta(w_n1716_0[0]),.doutb(w_n1716_0[1]),.din(n1716));
	jspl jspl_w_n1717_0(.douta(w_n1717_0[0]),.doutb(w_n1717_0[1]),.din(n1717));
	jspl jspl_w_n1719_0(.douta(w_n1719_0[0]),.doutb(w_n1719_0[1]),.din(n1719));
	jspl jspl_w_n1720_0(.douta(w_n1720_0[0]),.doutb(w_dff_A_4SVq3Cyq9_1),.din(n1720));
	jspl jspl_w_n1725_0(.douta(w_n1725_0[0]),.doutb(w_n1725_0[1]),.din(n1725));
	jspl jspl_w_n1728_0(.douta(w_n1728_0[0]),.doutb(w_dff_A_KDTpLwao3_1),.din(n1728));
	jspl jspl_w_n1730_0(.douta(w_n1730_0[0]),.doutb(w_n1730_0[1]),.din(w_dff_B_9RcW6zgb1_2));
	jspl jspl_w_n1733_0(.douta(w_n1733_0[0]),.doutb(w_n1733_0[1]),.din(w_dff_B_xqDSkUBz5_2));
	jspl jspl_w_n1735_0(.douta(w_n1735_0[0]),.doutb(w_n1735_0[1]),.din(w_dff_B_5oksoLxC0_2));
	jspl jspl_w_n1738_0(.douta(w_n1738_0[0]),.doutb(w_n1738_0[1]),.din(w_dff_B_kfVdW4aC6_2));
	jspl jspl_w_n1740_0(.douta(w_n1740_0[0]),.doutb(w_n1740_0[1]),.din(w_dff_B_DI2GWMrx8_2));
	jspl jspl_w_n1743_0(.douta(w_n1743_0[0]),.doutb(w_n1743_0[1]),.din(w_dff_B_AdJXDMSH1_2));
	jspl jspl_w_n1744_0(.douta(w_n1744_0[0]),.doutb(w_n1744_0[1]),.din(w_dff_B_o76WopWf3_2));
	jspl jspl_w_n1745_0(.douta(w_n1745_0[0]),.doutb(w_n1745_0[1]),.din(w_dff_B_DfVGyMBd9_2));
	jspl jspl_w_n1748_0(.douta(w_n1748_0[0]),.doutb(w_n1748_0[1]),.din(n1748));
	jspl jspl_w_n1750_0(.douta(w_n1750_0[0]),.doutb(w_n1750_0[1]),.din(n1750));
	jspl jspl_w_n1751_0(.douta(w_n1751_0[0]),.doutb(w_n1751_0[1]),.din(n1751));
	jspl jspl_w_n1752_0(.douta(w_n1752_0[0]),.doutb(w_n1752_0[1]),.din(n1752));
	jspl jspl_w_n1753_0(.douta(w_n1753_0[0]),.doutb(w_n1753_0[1]),.din(n1753));
	jspl jspl_w_n1754_0(.douta(w_n1754_0[0]),.doutb(w_n1754_0[1]),.din(n1754));
	jspl jspl_w_n1755_0(.douta(w_n1755_0[0]),.doutb(w_n1755_0[1]),.din(n1755));
	jspl jspl_w_n1756_0(.douta(w_n1756_0[0]),.doutb(w_n1756_0[1]),.din(n1756));
	jspl jspl_w_n1757_0(.douta(w_n1757_0[0]),.doutb(w_n1757_0[1]),.din(n1757));
	jspl jspl_w_n1758_0(.douta(w_n1758_0[0]),.doutb(w_dff_A_3bR1yH9e9_1),.din(n1758));
	jspl jspl_w_n1765_0(.douta(w_n1765_0[0]),.doutb(w_n1765_0[1]),.din(n1765));
	jspl jspl_w_n1768_0(.douta(w_n1768_0[0]),.doutb(w_dff_A_NXdfcoJP4_1),.din(n1768));
	jspl jspl_w_n1770_0(.douta(w_n1770_0[0]),.doutb(w_n1770_0[1]),.din(w_dff_B_ZmG8bPWg0_2));
	jspl jspl_w_n1773_0(.douta(w_n1773_0[0]),.doutb(w_n1773_0[1]),.din(w_dff_B_75PHjK6M9_2));
	jspl jspl_w_n1775_0(.douta(w_n1775_0[0]),.doutb(w_n1775_0[1]),.din(w_dff_B_fpdTFUYa8_2));
	jspl jspl_w_n1778_0(.douta(w_n1778_0[0]),.doutb(w_n1778_0[1]),.din(w_dff_B_jQz8xYvG9_2));
	jspl jspl_w_n1779_0(.douta(w_n1779_0[0]),.doutb(w_n1779_0[1]),.din(w_dff_B_ZgDUxRu08_2));
	jspl jspl_w_n1780_0(.douta(w_n1780_0[0]),.doutb(w_n1780_0[1]),.din(w_dff_B_BsNym0BD6_2));
	jspl jspl_w_n1783_0(.douta(w_n1783_0[0]),.doutb(w_n1783_0[1]),.din(n1783));
	jspl jspl_w_n1785_0(.douta(w_n1785_0[0]),.doutb(w_n1785_0[1]),.din(n1785));
	jspl jspl_w_n1786_0(.douta(w_n1786_0[0]),.doutb(w_n1786_0[1]),.din(n1786));
	jspl jspl_w_n1787_0(.douta(w_n1787_0[0]),.doutb(w_n1787_0[1]),.din(n1787));
	jspl jspl_w_n1788_0(.douta(w_n1788_0[0]),.doutb(w_n1788_0[1]),.din(n1788));
	jspl jspl_w_n1789_0(.douta(w_n1789_0[0]),.doutb(w_n1789_0[1]),.din(n1789));
	jspl jspl_w_n1790_0(.douta(w_n1790_0[0]),.doutb(w_n1790_0[1]),.din(n1790));
	jspl jspl_w_n1791_0(.douta(w_n1791_0[0]),.doutb(w_dff_A_IoAnXfgU6_1),.din(n1791));
	jspl jspl_w_n1798_0(.douta(w_n1798_0[0]),.doutb(w_n1798_0[1]),.din(n1798));
	jspl jspl_w_n1801_0(.douta(w_n1801_0[0]),.doutb(w_dff_A_Hvb89mYh3_1),.din(n1801));
	jspl jspl_w_n1803_0(.douta(w_n1803_0[0]),.doutb(w_n1803_0[1]),.din(w_dff_B_eIaXRKAC9_2));
	jspl jspl_w_n1806_0(.douta(w_n1806_0[0]),.doutb(w_n1806_0[1]),.din(w_dff_B_hqG9jUJl5_2));
	jspl jspl_w_n1807_0(.douta(w_n1807_0[0]),.doutb(w_n1807_0[1]),.din(w_dff_B_NjmfjCyy8_2));
	jspl jspl_w_n1808_0(.douta(w_n1808_0[0]),.doutb(w_n1808_0[1]),.din(w_dff_B_ow1ACzzW2_2));
	jspl jspl_w_n1811_0(.douta(w_n1811_0[0]),.doutb(w_n1811_0[1]),.din(n1811));
	jspl jspl_w_n1813_0(.douta(w_n1813_0[0]),.doutb(w_n1813_0[1]),.din(n1813));
	jspl jspl_w_n1814_0(.douta(w_n1814_0[0]),.doutb(w_n1814_0[1]),.din(n1814));
	jspl jspl_w_n1815_0(.douta(w_n1815_0[0]),.doutb(w_n1815_0[1]),.din(n1815));
	jspl jspl_w_n1816_0(.douta(w_n1816_0[0]),.doutb(w_n1816_0[1]),.din(n1816));
	jspl jspl_w_n1817_0(.douta(w_n1817_0[0]),.doutb(w_dff_A_eIaV6tH83_1),.din(n1817));
	jspl jspl_w_n1824_0(.douta(w_n1824_0[0]),.doutb(w_n1824_0[1]),.din(n1824));
	jspl jspl_w_n1827_0(.douta(w_n1827_0[0]),.doutb(w_dff_A_aQrQ35x31_1),.din(n1827));
	jspl jspl_w_n1828_0(.douta(w_n1828_0[0]),.doutb(w_n1828_0[1]),.din(w_dff_B_fosja2Hu4_2));
	jspl jspl_w_n1829_0(.douta(w_n1829_0[0]),.doutb(w_n1829_0[1]),.din(w_dff_B_DWU7mLRu5_2));
	jspl jspl_w_n1832_0(.douta(w_n1832_0[0]),.doutb(w_n1832_0[1]),.din(n1832));
	jspl jspl_w_n1834_0(.douta(w_n1834_0[0]),.doutb(w_n1834_0[1]),.din(n1834));
	jspl jspl_w_n1835_0(.douta(w_n1835_0[0]),.doutb(w_n1835_0[1]),.din(n1835));
	jspl jspl_w_n1836_0(.douta(w_n1836_0[0]),.doutb(w_dff_A_0qrSNxvr5_1),.din(n1836));
	jspl jspl_w_n1838_0(.douta(w_n1838_0[0]),.doutb(w_n1838_0[1]),.din(w_dff_B_Z1zRk0uY1_2));
	jspl jspl_w_n1841_0(.douta(w_n1841_0[0]),.doutb(w_n1841_0[1]),.din(n1841));
	jspl jspl_w_n1848_0(.douta(w_n1848_0[0]),.doutb(w_n1848_0[1]),.din(n1848));
	jspl jspl_w_n1849_0(.douta(w_dff_A_QBk0R33Z3_0),.doutb(w_n1849_0[1]),.din(n1849));
	jdff dff_B_3FRV3OSY1_1(.din(n67),.dout(w_dff_B_3FRV3OSY1_1),.clk(gclk));
	jdff dff_B_tzS6DnrW4_1(.din(n73),.dout(w_dff_B_tzS6DnrW4_1),.clk(gclk));
	jdff dff_B_VxIDHxam6_1(.din(w_dff_B_tzS6DnrW4_1),.dout(w_dff_B_VxIDHxam6_1),.clk(gclk));
	jdff dff_B_ha9tIQWA4_1(.din(w_dff_B_VxIDHxam6_1),.dout(w_dff_B_ha9tIQWA4_1),.clk(gclk));
	jdff dff_B_jMMSq32A1_1(.din(w_dff_B_ha9tIQWA4_1),.dout(w_dff_B_jMMSq32A1_1),.clk(gclk));
	jdff dff_B_ZlFNlmzc9_1(.din(n90),.dout(w_dff_B_ZlFNlmzc9_1),.clk(gclk));
	jdff dff_B_6XD066jy3_1(.din(w_dff_B_ZlFNlmzc9_1),.dout(w_dff_B_6XD066jy3_1),.clk(gclk));
	jdff dff_B_9OzVm5of4_1(.din(w_dff_B_6XD066jy3_1),.dout(w_dff_B_9OzVm5of4_1),.clk(gclk));
	jdff dff_B_veTJQclE4_1(.din(w_dff_B_9OzVm5of4_1),.dout(w_dff_B_veTJQclE4_1),.clk(gclk));
	jdff dff_B_x5apiaGv1_1(.din(w_dff_B_veTJQclE4_1),.dout(w_dff_B_x5apiaGv1_1),.clk(gclk));
	jdff dff_B_1mlkccCS3_1(.din(w_dff_B_x5apiaGv1_1),.dout(w_dff_B_1mlkccCS3_1),.clk(gclk));
	jdff dff_B_cSsKQ9UH7_1(.din(w_dff_B_1mlkccCS3_1),.dout(w_dff_B_cSsKQ9UH7_1),.clk(gclk));
	jdff dff_B_TqF3Kyx21_1(.din(n111),.dout(w_dff_B_TqF3Kyx21_1),.clk(gclk));
	jdff dff_B_YjBbOTB80_1(.din(w_dff_B_TqF3Kyx21_1),.dout(w_dff_B_YjBbOTB80_1),.clk(gclk));
	jdff dff_B_BOxqgtoR5_1(.din(w_dff_B_YjBbOTB80_1),.dout(w_dff_B_BOxqgtoR5_1),.clk(gclk));
	jdff dff_B_Xxmuud8I0_1(.din(w_dff_B_BOxqgtoR5_1),.dout(w_dff_B_Xxmuud8I0_1),.clk(gclk));
	jdff dff_B_b1tBh9bS4_1(.din(w_dff_B_Xxmuud8I0_1),.dout(w_dff_B_b1tBh9bS4_1),.clk(gclk));
	jdff dff_B_UsYlwApm6_1(.din(w_dff_B_b1tBh9bS4_1),.dout(w_dff_B_UsYlwApm6_1),.clk(gclk));
	jdff dff_B_DsS1jNqW1_1(.din(w_dff_B_UsYlwApm6_1),.dout(w_dff_B_DsS1jNqW1_1),.clk(gclk));
	jdff dff_B_8wetMZx70_1(.din(w_dff_B_DsS1jNqW1_1),.dout(w_dff_B_8wetMZx70_1),.clk(gclk));
	jdff dff_B_l6ggz8262_1(.din(w_dff_B_8wetMZx70_1),.dout(w_dff_B_l6ggz8262_1),.clk(gclk));
	jdff dff_B_8JplcJiB0_1(.din(w_dff_B_l6ggz8262_1),.dout(w_dff_B_8JplcJiB0_1),.clk(gclk));
	jdff dff_B_XbHPK9DO3_1(.din(n146),.dout(w_dff_B_XbHPK9DO3_1),.clk(gclk));
	jdff dff_B_e6cgpSpf1_1(.din(w_dff_B_XbHPK9DO3_1),.dout(w_dff_B_e6cgpSpf1_1),.clk(gclk));
	jdff dff_B_2KBjygSb8_1(.din(w_dff_B_e6cgpSpf1_1),.dout(w_dff_B_2KBjygSb8_1),.clk(gclk));
	jdff dff_B_8yoM9yav3_1(.din(w_dff_B_2KBjygSb8_1),.dout(w_dff_B_8yoM9yav3_1),.clk(gclk));
	jdff dff_B_tlcf4OLo2_1(.din(w_dff_B_8yoM9yav3_1),.dout(w_dff_B_tlcf4OLo2_1),.clk(gclk));
	jdff dff_B_4imTgWz93_1(.din(w_dff_B_tlcf4OLo2_1),.dout(w_dff_B_4imTgWz93_1),.clk(gclk));
	jdff dff_B_jb3PVe8J8_1(.din(w_dff_B_4imTgWz93_1),.dout(w_dff_B_jb3PVe8J8_1),.clk(gclk));
	jdff dff_B_3BUodJPE9_1(.din(w_dff_B_jb3PVe8J8_1),.dout(w_dff_B_3BUodJPE9_1),.clk(gclk));
	jdff dff_B_0574HHts2_1(.din(w_dff_B_3BUodJPE9_1),.dout(w_dff_B_0574HHts2_1),.clk(gclk));
	jdff dff_B_1mRT852b6_1(.din(w_dff_B_0574HHts2_1),.dout(w_dff_B_1mRT852b6_1),.clk(gclk));
	jdff dff_B_r5OIKcNp3_1(.din(w_dff_B_1mRT852b6_1),.dout(w_dff_B_r5OIKcNp3_1),.clk(gclk));
	jdff dff_B_ywNGUkGh3_1(.din(w_dff_B_r5OIKcNp3_1),.dout(w_dff_B_ywNGUkGh3_1),.clk(gclk));
	jdff dff_B_QcEJJi5q5_1(.din(w_dff_B_ywNGUkGh3_1),.dout(w_dff_B_QcEJJi5q5_1),.clk(gclk));
	jdff dff_B_2sZeV0CD3_1(.din(n184),.dout(w_dff_B_2sZeV0CD3_1),.clk(gclk));
	jdff dff_B_ghT6ytBR1_1(.din(w_dff_B_2sZeV0CD3_1),.dout(w_dff_B_ghT6ytBR1_1),.clk(gclk));
	jdff dff_B_ysQBawSr4_1(.din(w_dff_B_ghT6ytBR1_1),.dout(w_dff_B_ysQBawSr4_1),.clk(gclk));
	jdff dff_B_pveCeIwn2_1(.din(w_dff_B_ysQBawSr4_1),.dout(w_dff_B_pveCeIwn2_1),.clk(gclk));
	jdff dff_B_VObvQZJ06_1(.din(w_dff_B_pveCeIwn2_1),.dout(w_dff_B_VObvQZJ06_1),.clk(gclk));
	jdff dff_B_ExXvj7BS1_1(.din(w_dff_B_VObvQZJ06_1),.dout(w_dff_B_ExXvj7BS1_1),.clk(gclk));
	jdff dff_B_j1cevLAF1_1(.din(w_dff_B_ExXvj7BS1_1),.dout(w_dff_B_j1cevLAF1_1),.clk(gclk));
	jdff dff_B_GxfvPRXo7_1(.din(w_dff_B_j1cevLAF1_1),.dout(w_dff_B_GxfvPRXo7_1),.clk(gclk));
	jdff dff_B_HhQvWPrz0_1(.din(w_dff_B_GxfvPRXo7_1),.dout(w_dff_B_HhQvWPrz0_1),.clk(gclk));
	jdff dff_B_mnqfQLlW2_1(.din(w_dff_B_HhQvWPrz0_1),.dout(w_dff_B_mnqfQLlW2_1),.clk(gclk));
	jdff dff_B_z9VEiMmP8_1(.din(w_dff_B_mnqfQLlW2_1),.dout(w_dff_B_z9VEiMmP8_1),.clk(gclk));
	jdff dff_B_xMn0ITae1_1(.din(w_dff_B_z9VEiMmP8_1),.dout(w_dff_B_xMn0ITae1_1),.clk(gclk));
	jdff dff_B_ewCwHZCZ0_1(.din(w_dff_B_xMn0ITae1_1),.dout(w_dff_B_ewCwHZCZ0_1),.clk(gclk));
	jdff dff_B_QoLFz0zf3_1(.din(w_dff_B_ewCwHZCZ0_1),.dout(w_dff_B_QoLFz0zf3_1),.clk(gclk));
	jdff dff_B_l86IBcNm1_1(.din(w_dff_B_QoLFz0zf3_1),.dout(w_dff_B_l86IBcNm1_1),.clk(gclk));
	jdff dff_B_kiwggGnl5_1(.din(w_dff_B_l86IBcNm1_1),.dout(w_dff_B_kiwggGnl5_1),.clk(gclk));
	jdff dff_B_abxSj8tI2_1(.din(n227),.dout(w_dff_B_abxSj8tI2_1),.clk(gclk));
	jdff dff_B_fmM58jD45_1(.din(w_dff_B_abxSj8tI2_1),.dout(w_dff_B_fmM58jD45_1),.clk(gclk));
	jdff dff_B_SVDUn8oa2_1(.din(w_dff_B_fmM58jD45_1),.dout(w_dff_B_SVDUn8oa2_1),.clk(gclk));
	jdff dff_B_j3ONxwAh5_1(.din(w_dff_B_SVDUn8oa2_1),.dout(w_dff_B_j3ONxwAh5_1),.clk(gclk));
	jdff dff_B_aw7WoDnN4_1(.din(w_dff_B_j3ONxwAh5_1),.dout(w_dff_B_aw7WoDnN4_1),.clk(gclk));
	jdff dff_B_7GY3ZO541_1(.din(w_dff_B_aw7WoDnN4_1),.dout(w_dff_B_7GY3ZO541_1),.clk(gclk));
	jdff dff_B_lOjagvgO9_1(.din(w_dff_B_7GY3ZO541_1),.dout(w_dff_B_lOjagvgO9_1),.clk(gclk));
	jdff dff_B_vYASkG8n9_1(.din(w_dff_B_lOjagvgO9_1),.dout(w_dff_B_vYASkG8n9_1),.clk(gclk));
	jdff dff_B_U1Pd7OVs7_1(.din(w_dff_B_vYASkG8n9_1),.dout(w_dff_B_U1Pd7OVs7_1),.clk(gclk));
	jdff dff_B_5zUAPdQo9_1(.din(w_dff_B_U1Pd7OVs7_1),.dout(w_dff_B_5zUAPdQo9_1),.clk(gclk));
	jdff dff_B_GsaYMcr60_1(.din(w_dff_B_5zUAPdQo9_1),.dout(w_dff_B_GsaYMcr60_1),.clk(gclk));
	jdff dff_B_cknEWKCP9_1(.din(w_dff_B_GsaYMcr60_1),.dout(w_dff_B_cknEWKCP9_1),.clk(gclk));
	jdff dff_B_RTzxDbo07_1(.din(w_dff_B_cknEWKCP9_1),.dout(w_dff_B_RTzxDbo07_1),.clk(gclk));
	jdff dff_B_tfuvyd3x2_1(.din(w_dff_B_RTzxDbo07_1),.dout(w_dff_B_tfuvyd3x2_1),.clk(gclk));
	jdff dff_B_AF5hPx0J7_1(.din(w_dff_B_tfuvyd3x2_1),.dout(w_dff_B_AF5hPx0J7_1),.clk(gclk));
	jdff dff_B_uXxDI9bO5_1(.din(w_dff_B_AF5hPx0J7_1),.dout(w_dff_B_uXxDI9bO5_1),.clk(gclk));
	jdff dff_B_rjvlO9LX2_1(.din(w_dff_B_uXxDI9bO5_1),.dout(w_dff_B_rjvlO9LX2_1),.clk(gclk));
	jdff dff_B_LDGGGVfw2_1(.din(w_dff_B_rjvlO9LX2_1),.dout(w_dff_B_LDGGGVfw2_1),.clk(gclk));
	jdff dff_B_TAGRaUJf0_1(.din(w_dff_B_LDGGGVfw2_1),.dout(w_dff_B_TAGRaUJf0_1),.clk(gclk));
	jdff dff_B_m3IXWPoE5_1(.din(n278),.dout(w_dff_B_m3IXWPoE5_1),.clk(gclk));
	jdff dff_B_fq4LRnHV2_1(.din(w_dff_B_m3IXWPoE5_1),.dout(w_dff_B_fq4LRnHV2_1),.clk(gclk));
	jdff dff_B_P0aUQM8E8_1(.din(w_dff_B_fq4LRnHV2_1),.dout(w_dff_B_P0aUQM8E8_1),.clk(gclk));
	jdff dff_B_RyggImi25_1(.din(w_dff_B_P0aUQM8E8_1),.dout(w_dff_B_RyggImi25_1),.clk(gclk));
	jdff dff_B_s5qXbtjj8_1(.din(w_dff_B_RyggImi25_1),.dout(w_dff_B_s5qXbtjj8_1),.clk(gclk));
	jdff dff_B_yarOBbtK5_1(.din(w_dff_B_s5qXbtjj8_1),.dout(w_dff_B_yarOBbtK5_1),.clk(gclk));
	jdff dff_B_4iVZKolt8_1(.din(w_dff_B_yarOBbtK5_1),.dout(w_dff_B_4iVZKolt8_1),.clk(gclk));
	jdff dff_B_i7QAnRf78_1(.din(w_dff_B_4iVZKolt8_1),.dout(w_dff_B_i7QAnRf78_1),.clk(gclk));
	jdff dff_B_L4G8jCl37_1(.din(w_dff_B_i7QAnRf78_1),.dout(w_dff_B_L4G8jCl37_1),.clk(gclk));
	jdff dff_B_eGvjOvZb0_1(.din(w_dff_B_L4G8jCl37_1),.dout(w_dff_B_eGvjOvZb0_1),.clk(gclk));
	jdff dff_B_OEpOfUij9_1(.din(w_dff_B_eGvjOvZb0_1),.dout(w_dff_B_OEpOfUij9_1),.clk(gclk));
	jdff dff_B_LpCIXDfk1_1(.din(w_dff_B_OEpOfUij9_1),.dout(w_dff_B_LpCIXDfk1_1),.clk(gclk));
	jdff dff_B_f7FUm4Yq4_1(.din(w_dff_B_LpCIXDfk1_1),.dout(w_dff_B_f7FUm4Yq4_1),.clk(gclk));
	jdff dff_B_LgnLW0fG9_1(.din(w_dff_B_f7FUm4Yq4_1),.dout(w_dff_B_LgnLW0fG9_1),.clk(gclk));
	jdff dff_B_OdqFMnh06_1(.din(w_dff_B_LgnLW0fG9_1),.dout(w_dff_B_OdqFMnh06_1),.clk(gclk));
	jdff dff_B_nB35EGLw1_1(.din(w_dff_B_OdqFMnh06_1),.dout(w_dff_B_nB35EGLw1_1),.clk(gclk));
	jdff dff_B_IUKdWtAb3_1(.din(w_dff_B_nB35EGLw1_1),.dout(w_dff_B_IUKdWtAb3_1),.clk(gclk));
	jdff dff_B_0GZO3Pon4_1(.din(w_dff_B_IUKdWtAb3_1),.dout(w_dff_B_0GZO3Pon4_1),.clk(gclk));
	jdff dff_B_MCKfq1186_1(.din(w_dff_B_0GZO3Pon4_1),.dout(w_dff_B_MCKfq1186_1),.clk(gclk));
	jdff dff_B_VND7Ereb9_1(.din(w_dff_B_MCKfq1186_1),.dout(w_dff_B_VND7Ereb9_1),.clk(gclk));
	jdff dff_B_WDv7auJn1_1(.din(w_dff_B_VND7Ereb9_1),.dout(w_dff_B_WDv7auJn1_1),.clk(gclk));
	jdff dff_B_NtzpAMMQ5_1(.din(w_dff_B_WDv7auJn1_1),.dout(w_dff_B_NtzpAMMQ5_1),.clk(gclk));
	jdff dff_B_tM6B2SdG8_1(.din(n336),.dout(w_dff_B_tM6B2SdG8_1),.clk(gclk));
	jdff dff_B_hxb9EYi46_1(.din(w_dff_B_tM6B2SdG8_1),.dout(w_dff_B_hxb9EYi46_1),.clk(gclk));
	jdff dff_B_HAvgtCbm0_1(.din(w_dff_B_hxb9EYi46_1),.dout(w_dff_B_HAvgtCbm0_1),.clk(gclk));
	jdff dff_B_xlDvBJx33_1(.din(w_dff_B_HAvgtCbm0_1),.dout(w_dff_B_xlDvBJx33_1),.clk(gclk));
	jdff dff_B_I3fXIWZ77_1(.din(w_dff_B_xlDvBJx33_1),.dout(w_dff_B_I3fXIWZ77_1),.clk(gclk));
	jdff dff_B_mnw3fniH1_1(.din(w_dff_B_I3fXIWZ77_1),.dout(w_dff_B_mnw3fniH1_1),.clk(gclk));
	jdff dff_B_zvg1jZKl6_1(.din(w_dff_B_mnw3fniH1_1),.dout(w_dff_B_zvg1jZKl6_1),.clk(gclk));
	jdff dff_B_dluCOjUp9_1(.din(w_dff_B_zvg1jZKl6_1),.dout(w_dff_B_dluCOjUp9_1),.clk(gclk));
	jdff dff_B_U0UsSENG4_1(.din(w_dff_B_dluCOjUp9_1),.dout(w_dff_B_U0UsSENG4_1),.clk(gclk));
	jdff dff_B_NyKtFR510_1(.din(w_dff_B_U0UsSENG4_1),.dout(w_dff_B_NyKtFR510_1),.clk(gclk));
	jdff dff_B_jj6fPb5s9_1(.din(w_dff_B_NyKtFR510_1),.dout(w_dff_B_jj6fPb5s9_1),.clk(gclk));
	jdff dff_B_emUqo5MA2_1(.din(w_dff_B_jj6fPb5s9_1),.dout(w_dff_B_emUqo5MA2_1),.clk(gclk));
	jdff dff_B_09jwJg3T4_1(.din(w_dff_B_emUqo5MA2_1),.dout(w_dff_B_09jwJg3T4_1),.clk(gclk));
	jdff dff_B_QI2QzpDT6_1(.din(w_dff_B_09jwJg3T4_1),.dout(w_dff_B_QI2QzpDT6_1),.clk(gclk));
	jdff dff_B_AJT4CnW13_1(.din(w_dff_B_QI2QzpDT6_1),.dout(w_dff_B_AJT4CnW13_1),.clk(gclk));
	jdff dff_B_emjodvUZ5_1(.din(w_dff_B_AJT4CnW13_1),.dout(w_dff_B_emjodvUZ5_1),.clk(gclk));
	jdff dff_B_LVmnjLSK7_1(.din(w_dff_B_emjodvUZ5_1),.dout(w_dff_B_LVmnjLSK7_1),.clk(gclk));
	jdff dff_B_HMddPGFz1_1(.din(w_dff_B_LVmnjLSK7_1),.dout(w_dff_B_HMddPGFz1_1),.clk(gclk));
	jdff dff_B_xCTg7QvE2_1(.din(w_dff_B_HMddPGFz1_1),.dout(w_dff_B_xCTg7QvE2_1),.clk(gclk));
	jdff dff_B_d8mlmS3d1_1(.din(w_dff_B_xCTg7QvE2_1),.dout(w_dff_B_d8mlmS3d1_1),.clk(gclk));
	jdff dff_B_6rj66GPP9_1(.din(w_dff_B_d8mlmS3d1_1),.dout(w_dff_B_6rj66GPP9_1),.clk(gclk));
	jdff dff_B_BegVnqY61_1(.din(w_dff_B_6rj66GPP9_1),.dout(w_dff_B_BegVnqY61_1),.clk(gclk));
	jdff dff_B_nlzDf3JQ8_1(.din(w_dff_B_BegVnqY61_1),.dout(w_dff_B_nlzDf3JQ8_1),.clk(gclk));
	jdff dff_B_p5ZFmHRw7_1(.din(w_dff_B_nlzDf3JQ8_1),.dout(w_dff_B_p5ZFmHRw7_1),.clk(gclk));
	jdff dff_B_7PYVdMoG0_1(.din(w_dff_B_p5ZFmHRw7_1),.dout(w_dff_B_7PYVdMoG0_1),.clk(gclk));
	jdff dff_B_f7ERvtf70_1(.din(n400),.dout(w_dff_B_f7ERvtf70_1),.clk(gclk));
	jdff dff_B_wiUZgfzF6_1(.din(w_dff_B_f7ERvtf70_1),.dout(w_dff_B_wiUZgfzF6_1),.clk(gclk));
	jdff dff_B_HhkEzole3_1(.din(w_dff_B_wiUZgfzF6_1),.dout(w_dff_B_HhkEzole3_1),.clk(gclk));
	jdff dff_B_ClOxpV8b1_1(.din(w_dff_B_HhkEzole3_1),.dout(w_dff_B_ClOxpV8b1_1),.clk(gclk));
	jdff dff_B_fAWMF5Wi6_1(.din(w_dff_B_ClOxpV8b1_1),.dout(w_dff_B_fAWMF5Wi6_1),.clk(gclk));
	jdff dff_B_j4ubxkx71_1(.din(w_dff_B_fAWMF5Wi6_1),.dout(w_dff_B_j4ubxkx71_1),.clk(gclk));
	jdff dff_B_g0qfZzsD4_1(.din(w_dff_B_j4ubxkx71_1),.dout(w_dff_B_g0qfZzsD4_1),.clk(gclk));
	jdff dff_B_7qAExO8r4_1(.din(w_dff_B_g0qfZzsD4_1),.dout(w_dff_B_7qAExO8r4_1),.clk(gclk));
	jdff dff_B_2qeprMuU1_1(.din(w_dff_B_7qAExO8r4_1),.dout(w_dff_B_2qeprMuU1_1),.clk(gclk));
	jdff dff_B_YTgH9Afm7_1(.din(w_dff_B_2qeprMuU1_1),.dout(w_dff_B_YTgH9Afm7_1),.clk(gclk));
	jdff dff_B_zcqFA8Wl0_1(.din(w_dff_B_YTgH9Afm7_1),.dout(w_dff_B_zcqFA8Wl0_1),.clk(gclk));
	jdff dff_B_zOMgdbVA7_1(.din(w_dff_B_zcqFA8Wl0_1),.dout(w_dff_B_zOMgdbVA7_1),.clk(gclk));
	jdff dff_B_lVWfBE479_1(.din(w_dff_B_zOMgdbVA7_1),.dout(w_dff_B_lVWfBE479_1),.clk(gclk));
	jdff dff_B_rWv6YpuE1_1(.din(w_dff_B_lVWfBE479_1),.dout(w_dff_B_rWv6YpuE1_1),.clk(gclk));
	jdff dff_B_slmxmLJT8_1(.din(w_dff_B_rWv6YpuE1_1),.dout(w_dff_B_slmxmLJT8_1),.clk(gclk));
	jdff dff_B_JoeVYMHM5_1(.din(w_dff_B_slmxmLJT8_1),.dout(w_dff_B_JoeVYMHM5_1),.clk(gclk));
	jdff dff_B_zSendvSt1_1(.din(w_dff_B_JoeVYMHM5_1),.dout(w_dff_B_zSendvSt1_1),.clk(gclk));
	jdff dff_B_S15Yp8XT0_1(.din(w_dff_B_zSendvSt1_1),.dout(w_dff_B_S15Yp8XT0_1),.clk(gclk));
	jdff dff_B_ot8aqExn0_1(.din(w_dff_B_S15Yp8XT0_1),.dout(w_dff_B_ot8aqExn0_1),.clk(gclk));
	jdff dff_B_CFn3SMXg3_1(.din(w_dff_B_ot8aqExn0_1),.dout(w_dff_B_CFn3SMXg3_1),.clk(gclk));
	jdff dff_B_mn1cQTSZ7_1(.din(w_dff_B_CFn3SMXg3_1),.dout(w_dff_B_mn1cQTSZ7_1),.clk(gclk));
	jdff dff_B_fb82xcaX4_1(.din(w_dff_B_mn1cQTSZ7_1),.dout(w_dff_B_fb82xcaX4_1),.clk(gclk));
	jdff dff_B_oU3W5YhB5_1(.din(w_dff_B_fb82xcaX4_1),.dout(w_dff_B_oU3W5YhB5_1),.clk(gclk));
	jdff dff_B_mBXNtslG7_1(.din(w_dff_B_oU3W5YhB5_1),.dout(w_dff_B_mBXNtslG7_1),.clk(gclk));
	jdff dff_B_f2vFp1tY3_1(.din(w_dff_B_mBXNtslG7_1),.dout(w_dff_B_f2vFp1tY3_1),.clk(gclk));
	jdff dff_B_0TqlkH5f5_1(.din(w_dff_B_f2vFp1tY3_1),.dout(w_dff_B_0TqlkH5f5_1),.clk(gclk));
	jdff dff_B_KpMIxvXc7_1(.din(w_dff_B_0TqlkH5f5_1),.dout(w_dff_B_KpMIxvXc7_1),.clk(gclk));
	jdff dff_B_N82dfrYa9_1(.din(w_dff_B_KpMIxvXc7_1),.dout(w_dff_B_N82dfrYa9_1),.clk(gclk));
	jdff dff_B_vV4gSXGs0_1(.din(n472),.dout(w_dff_B_vV4gSXGs0_1),.clk(gclk));
	jdff dff_B_o8lrPJoM1_1(.din(w_dff_B_vV4gSXGs0_1),.dout(w_dff_B_o8lrPJoM1_1),.clk(gclk));
	jdff dff_B_r0o7HmVf9_1(.din(w_dff_B_o8lrPJoM1_1),.dout(w_dff_B_r0o7HmVf9_1),.clk(gclk));
	jdff dff_B_bjGuhllO6_1(.din(w_dff_B_r0o7HmVf9_1),.dout(w_dff_B_bjGuhllO6_1),.clk(gclk));
	jdff dff_B_T1AUH2Ff3_1(.din(w_dff_B_bjGuhllO6_1),.dout(w_dff_B_T1AUH2Ff3_1),.clk(gclk));
	jdff dff_B_5aQGEkCr3_1(.din(w_dff_B_T1AUH2Ff3_1),.dout(w_dff_B_5aQGEkCr3_1),.clk(gclk));
	jdff dff_B_atN5qAza3_1(.din(w_dff_B_5aQGEkCr3_1),.dout(w_dff_B_atN5qAza3_1),.clk(gclk));
	jdff dff_B_x6V5G3zo2_1(.din(w_dff_B_atN5qAza3_1),.dout(w_dff_B_x6V5G3zo2_1),.clk(gclk));
	jdff dff_B_6mRlSyiG1_1(.din(w_dff_B_x6V5G3zo2_1),.dout(w_dff_B_6mRlSyiG1_1),.clk(gclk));
	jdff dff_B_2HrLUCD95_1(.din(w_dff_B_6mRlSyiG1_1),.dout(w_dff_B_2HrLUCD95_1),.clk(gclk));
	jdff dff_B_SAwXU5909_1(.din(w_dff_B_2HrLUCD95_1),.dout(w_dff_B_SAwXU5909_1),.clk(gclk));
	jdff dff_B_alzmbQ5D8_1(.din(w_dff_B_SAwXU5909_1),.dout(w_dff_B_alzmbQ5D8_1),.clk(gclk));
	jdff dff_B_uos9j3hj8_1(.din(w_dff_B_alzmbQ5D8_1),.dout(w_dff_B_uos9j3hj8_1),.clk(gclk));
	jdff dff_B_p6s9f53C7_1(.din(w_dff_B_uos9j3hj8_1),.dout(w_dff_B_p6s9f53C7_1),.clk(gclk));
	jdff dff_B_23sqyV4G0_1(.din(w_dff_B_p6s9f53C7_1),.dout(w_dff_B_23sqyV4G0_1),.clk(gclk));
	jdff dff_B_tmRTLLGG7_1(.din(w_dff_B_23sqyV4G0_1),.dout(w_dff_B_tmRTLLGG7_1),.clk(gclk));
	jdff dff_B_LdNvkQAU9_1(.din(w_dff_B_tmRTLLGG7_1),.dout(w_dff_B_LdNvkQAU9_1),.clk(gclk));
	jdff dff_B_ksqaA3H48_1(.din(w_dff_B_LdNvkQAU9_1),.dout(w_dff_B_ksqaA3H48_1),.clk(gclk));
	jdff dff_B_n4wnCgRt3_1(.din(w_dff_B_ksqaA3H48_1),.dout(w_dff_B_n4wnCgRt3_1),.clk(gclk));
	jdff dff_B_tHAqzUIO9_1(.din(w_dff_B_n4wnCgRt3_1),.dout(w_dff_B_tHAqzUIO9_1),.clk(gclk));
	jdff dff_B_LiPwz7S20_1(.din(w_dff_B_tHAqzUIO9_1),.dout(w_dff_B_LiPwz7S20_1),.clk(gclk));
	jdff dff_B_fS7HDFdk1_1(.din(w_dff_B_LiPwz7S20_1),.dout(w_dff_B_fS7HDFdk1_1),.clk(gclk));
	jdff dff_B_vd6OvMni6_1(.din(w_dff_B_fS7HDFdk1_1),.dout(w_dff_B_vd6OvMni6_1),.clk(gclk));
	jdff dff_B_X402efUH3_1(.din(w_dff_B_vd6OvMni6_1),.dout(w_dff_B_X402efUH3_1),.clk(gclk));
	jdff dff_B_YBmjWnM61_1(.din(w_dff_B_X402efUH3_1),.dout(w_dff_B_YBmjWnM61_1),.clk(gclk));
	jdff dff_B_wttfy1U82_1(.din(w_dff_B_YBmjWnM61_1),.dout(w_dff_B_wttfy1U82_1),.clk(gclk));
	jdff dff_B_DBNqSZ240_1(.din(w_dff_B_wttfy1U82_1),.dout(w_dff_B_DBNqSZ240_1),.clk(gclk));
	jdff dff_B_d8wE2Uer4_1(.din(w_dff_B_DBNqSZ240_1),.dout(w_dff_B_d8wE2Uer4_1),.clk(gclk));
	jdff dff_B_QZdtZDCn1_1(.din(w_dff_B_d8wE2Uer4_1),.dout(w_dff_B_QZdtZDCn1_1),.clk(gclk));
	jdff dff_B_Yr1vIQ269_1(.din(w_dff_B_QZdtZDCn1_1),.dout(w_dff_B_Yr1vIQ269_1),.clk(gclk));
	jdff dff_B_rp1raYfx8_1(.din(w_dff_B_Yr1vIQ269_1),.dout(w_dff_B_rp1raYfx8_1),.clk(gclk));
	jdff dff_B_kCXG7ccs1_1(.din(n551),.dout(w_dff_B_kCXG7ccs1_1),.clk(gclk));
	jdff dff_B_tfPxnPeR4_1(.din(w_dff_B_kCXG7ccs1_1),.dout(w_dff_B_tfPxnPeR4_1),.clk(gclk));
	jdff dff_B_KyjXoe9I9_1(.din(w_dff_B_tfPxnPeR4_1),.dout(w_dff_B_KyjXoe9I9_1),.clk(gclk));
	jdff dff_B_WXo3Jx9S1_1(.din(w_dff_B_KyjXoe9I9_1),.dout(w_dff_B_WXo3Jx9S1_1),.clk(gclk));
	jdff dff_B_CQWxuADi2_1(.din(w_dff_B_WXo3Jx9S1_1),.dout(w_dff_B_CQWxuADi2_1),.clk(gclk));
	jdff dff_B_ewuybWPi6_1(.din(w_dff_B_CQWxuADi2_1),.dout(w_dff_B_ewuybWPi6_1),.clk(gclk));
	jdff dff_B_nFucVkYg9_1(.din(w_dff_B_ewuybWPi6_1),.dout(w_dff_B_nFucVkYg9_1),.clk(gclk));
	jdff dff_B_OEPrANys4_1(.din(w_dff_B_nFucVkYg9_1),.dout(w_dff_B_OEPrANys4_1),.clk(gclk));
	jdff dff_B_3FMTbEV32_1(.din(w_dff_B_OEPrANys4_1),.dout(w_dff_B_3FMTbEV32_1),.clk(gclk));
	jdff dff_B_cVsX0Vlq1_1(.din(w_dff_B_3FMTbEV32_1),.dout(w_dff_B_cVsX0Vlq1_1),.clk(gclk));
	jdff dff_B_7yipnxMK4_1(.din(w_dff_B_cVsX0Vlq1_1),.dout(w_dff_B_7yipnxMK4_1),.clk(gclk));
	jdff dff_B_mZLm2enn4_1(.din(w_dff_B_7yipnxMK4_1),.dout(w_dff_B_mZLm2enn4_1),.clk(gclk));
	jdff dff_B_Mld6iIyQ6_1(.din(w_dff_B_mZLm2enn4_1),.dout(w_dff_B_Mld6iIyQ6_1),.clk(gclk));
	jdff dff_B_alg5Gp4J8_1(.din(w_dff_B_Mld6iIyQ6_1),.dout(w_dff_B_alg5Gp4J8_1),.clk(gclk));
	jdff dff_B_M7md7Umi8_1(.din(w_dff_B_alg5Gp4J8_1),.dout(w_dff_B_M7md7Umi8_1),.clk(gclk));
	jdff dff_B_4VdDZshB9_1(.din(w_dff_B_M7md7Umi8_1),.dout(w_dff_B_4VdDZshB9_1),.clk(gclk));
	jdff dff_B_kqR09lbr4_1(.din(w_dff_B_4VdDZshB9_1),.dout(w_dff_B_kqR09lbr4_1),.clk(gclk));
	jdff dff_B_QPegivjI8_1(.din(w_dff_B_kqR09lbr4_1),.dout(w_dff_B_QPegivjI8_1),.clk(gclk));
	jdff dff_B_SDOqiyuU7_1(.din(w_dff_B_QPegivjI8_1),.dout(w_dff_B_SDOqiyuU7_1),.clk(gclk));
	jdff dff_B_oBlrIWPA2_1(.din(w_dff_B_SDOqiyuU7_1),.dout(w_dff_B_oBlrIWPA2_1),.clk(gclk));
	jdff dff_B_B5qQ1p6k5_1(.din(w_dff_B_oBlrIWPA2_1),.dout(w_dff_B_B5qQ1p6k5_1),.clk(gclk));
	jdff dff_B_GYsVnjmm1_1(.din(w_dff_B_B5qQ1p6k5_1),.dout(w_dff_B_GYsVnjmm1_1),.clk(gclk));
	jdff dff_B_be6zHySW2_1(.din(w_dff_B_GYsVnjmm1_1),.dout(w_dff_B_be6zHySW2_1),.clk(gclk));
	jdff dff_B_SWoxspAq3_1(.din(w_dff_B_be6zHySW2_1),.dout(w_dff_B_SWoxspAq3_1),.clk(gclk));
	jdff dff_B_6m5zXTgz9_1(.din(w_dff_B_SWoxspAq3_1),.dout(w_dff_B_6m5zXTgz9_1),.clk(gclk));
	jdff dff_B_DAUafqyZ5_1(.din(w_dff_B_6m5zXTgz9_1),.dout(w_dff_B_DAUafqyZ5_1),.clk(gclk));
	jdff dff_B_hZnynIeh0_1(.din(w_dff_B_DAUafqyZ5_1),.dout(w_dff_B_hZnynIeh0_1),.clk(gclk));
	jdff dff_B_ifkqVlaJ3_1(.din(w_dff_B_hZnynIeh0_1),.dout(w_dff_B_ifkqVlaJ3_1),.clk(gclk));
	jdff dff_B_29WaMTkW6_1(.din(w_dff_B_ifkqVlaJ3_1),.dout(w_dff_B_29WaMTkW6_1),.clk(gclk));
	jdff dff_B_QUYCBp1w1_1(.din(w_dff_B_29WaMTkW6_1),.dout(w_dff_B_QUYCBp1w1_1),.clk(gclk));
	jdff dff_B_MYLIJuEe3_1(.din(w_dff_B_QUYCBp1w1_1),.dout(w_dff_B_MYLIJuEe3_1),.clk(gclk));
	jdff dff_B_pAA7W6Lg1_1(.din(w_dff_B_MYLIJuEe3_1),.dout(w_dff_B_pAA7W6Lg1_1),.clk(gclk));
	jdff dff_B_gL4nA4Lz8_1(.din(w_dff_B_pAA7W6Lg1_1),.dout(w_dff_B_gL4nA4Lz8_1),.clk(gclk));
	jdff dff_B_3CG9xstA3_1(.din(w_dff_B_gL4nA4Lz8_1),.dout(w_dff_B_3CG9xstA3_1),.clk(gclk));
	jdff dff_B_1Qz7w2UC3_1(.din(n637),.dout(w_dff_B_1Qz7w2UC3_1),.clk(gclk));
	jdff dff_B_8vGu5hgd2_1(.din(w_dff_B_1Qz7w2UC3_1),.dout(w_dff_B_8vGu5hgd2_1),.clk(gclk));
	jdff dff_B_rOZ0ysnI4_1(.din(w_dff_B_8vGu5hgd2_1),.dout(w_dff_B_rOZ0ysnI4_1),.clk(gclk));
	jdff dff_B_8NtzV6A68_1(.din(w_dff_B_rOZ0ysnI4_1),.dout(w_dff_B_8NtzV6A68_1),.clk(gclk));
	jdff dff_B_Yb6stWZa1_1(.din(w_dff_B_8NtzV6A68_1),.dout(w_dff_B_Yb6stWZa1_1),.clk(gclk));
	jdff dff_B_Uv0qjueR9_1(.din(w_dff_B_Yb6stWZa1_1),.dout(w_dff_B_Uv0qjueR9_1),.clk(gclk));
	jdff dff_B_evmr8apB2_1(.din(w_dff_B_Uv0qjueR9_1),.dout(w_dff_B_evmr8apB2_1),.clk(gclk));
	jdff dff_B_Q0tinFuv6_1(.din(w_dff_B_evmr8apB2_1),.dout(w_dff_B_Q0tinFuv6_1),.clk(gclk));
	jdff dff_B_PmDzMrum9_1(.din(w_dff_B_Q0tinFuv6_1),.dout(w_dff_B_PmDzMrum9_1),.clk(gclk));
	jdff dff_B_gE6BLSiU0_1(.din(w_dff_B_PmDzMrum9_1),.dout(w_dff_B_gE6BLSiU0_1),.clk(gclk));
	jdff dff_B_ZYRBFtCg1_1(.din(w_dff_B_gE6BLSiU0_1),.dout(w_dff_B_ZYRBFtCg1_1),.clk(gclk));
	jdff dff_B_6M1Gccuy5_1(.din(w_dff_B_ZYRBFtCg1_1),.dout(w_dff_B_6M1Gccuy5_1),.clk(gclk));
	jdff dff_B_c4FUp6yr5_1(.din(w_dff_B_6M1Gccuy5_1),.dout(w_dff_B_c4FUp6yr5_1),.clk(gclk));
	jdff dff_B_9uueaT3B7_1(.din(w_dff_B_c4FUp6yr5_1),.dout(w_dff_B_9uueaT3B7_1),.clk(gclk));
	jdff dff_B_n74dByiy5_1(.din(w_dff_B_9uueaT3B7_1),.dout(w_dff_B_n74dByiy5_1),.clk(gclk));
	jdff dff_B_i5xs0pLM2_1(.din(w_dff_B_n74dByiy5_1),.dout(w_dff_B_i5xs0pLM2_1),.clk(gclk));
	jdff dff_B_D8QHiqNG5_1(.din(w_dff_B_i5xs0pLM2_1),.dout(w_dff_B_D8QHiqNG5_1),.clk(gclk));
	jdff dff_B_WEtqzBk58_1(.din(w_dff_B_D8QHiqNG5_1),.dout(w_dff_B_WEtqzBk58_1),.clk(gclk));
	jdff dff_B_XxrgRmDw6_1(.din(w_dff_B_WEtqzBk58_1),.dout(w_dff_B_XxrgRmDw6_1),.clk(gclk));
	jdff dff_B_ux8VR4h52_1(.din(w_dff_B_XxrgRmDw6_1),.dout(w_dff_B_ux8VR4h52_1),.clk(gclk));
	jdff dff_B_0FWt9EOj8_1(.din(w_dff_B_ux8VR4h52_1),.dout(w_dff_B_0FWt9EOj8_1),.clk(gclk));
	jdff dff_B_OeLgFibZ7_1(.din(w_dff_B_0FWt9EOj8_1),.dout(w_dff_B_OeLgFibZ7_1),.clk(gclk));
	jdff dff_B_8gitHIJ50_1(.din(w_dff_B_OeLgFibZ7_1),.dout(w_dff_B_8gitHIJ50_1),.clk(gclk));
	jdff dff_B_3WcVn7vX6_1(.din(w_dff_B_8gitHIJ50_1),.dout(w_dff_B_3WcVn7vX6_1),.clk(gclk));
	jdff dff_B_rEOHq21o6_1(.din(w_dff_B_3WcVn7vX6_1),.dout(w_dff_B_rEOHq21o6_1),.clk(gclk));
	jdff dff_B_6NhvmuVH1_1(.din(w_dff_B_rEOHq21o6_1),.dout(w_dff_B_6NhvmuVH1_1),.clk(gclk));
	jdff dff_B_RWn2bz0N6_1(.din(w_dff_B_6NhvmuVH1_1),.dout(w_dff_B_RWn2bz0N6_1),.clk(gclk));
	jdff dff_B_EWMTpNai1_1(.din(w_dff_B_RWn2bz0N6_1),.dout(w_dff_B_EWMTpNai1_1),.clk(gclk));
	jdff dff_B_MerO0PB70_1(.din(w_dff_B_EWMTpNai1_1),.dout(w_dff_B_MerO0PB70_1),.clk(gclk));
	jdff dff_B_kFLXeI0q6_1(.din(w_dff_B_MerO0PB70_1),.dout(w_dff_B_kFLXeI0q6_1),.clk(gclk));
	jdff dff_B_cyMf9eUe5_1(.din(w_dff_B_kFLXeI0q6_1),.dout(w_dff_B_cyMf9eUe5_1),.clk(gclk));
	jdff dff_B_1ZEggp9p7_1(.din(w_dff_B_cyMf9eUe5_1),.dout(w_dff_B_1ZEggp9p7_1),.clk(gclk));
	jdff dff_B_xLb88RAj3_1(.din(w_dff_B_1ZEggp9p7_1),.dout(w_dff_B_xLb88RAj3_1),.clk(gclk));
	jdff dff_B_mtv59oc30_1(.din(w_dff_B_xLb88RAj3_1),.dout(w_dff_B_mtv59oc30_1),.clk(gclk));
	jdff dff_B_Isi4F8E74_1(.din(w_dff_B_mtv59oc30_1),.dout(w_dff_B_Isi4F8E74_1),.clk(gclk));
	jdff dff_B_Qcd02HFj4_1(.din(w_dff_B_Isi4F8E74_1),.dout(w_dff_B_Qcd02HFj4_1),.clk(gclk));
	jdff dff_B_tPTGsLaV0_1(.din(w_dff_B_Qcd02HFj4_1),.dout(w_dff_B_tPTGsLaV0_1),.clk(gclk));
	jdff dff_B_sFUxrmKn2_1(.din(n730),.dout(w_dff_B_sFUxrmKn2_1),.clk(gclk));
	jdff dff_B_a9lb9UVr0_1(.din(w_dff_B_sFUxrmKn2_1),.dout(w_dff_B_a9lb9UVr0_1),.clk(gclk));
	jdff dff_B_hCoDeQjV6_1(.din(w_dff_B_a9lb9UVr0_1),.dout(w_dff_B_hCoDeQjV6_1),.clk(gclk));
	jdff dff_B_gzVFP90e4_1(.din(w_dff_B_hCoDeQjV6_1),.dout(w_dff_B_gzVFP90e4_1),.clk(gclk));
	jdff dff_B_0WQxg2FI6_1(.din(w_dff_B_gzVFP90e4_1),.dout(w_dff_B_0WQxg2FI6_1),.clk(gclk));
	jdff dff_B_7NcIjERV3_1(.din(w_dff_B_0WQxg2FI6_1),.dout(w_dff_B_7NcIjERV3_1),.clk(gclk));
	jdff dff_B_nKF7123N6_1(.din(w_dff_B_7NcIjERV3_1),.dout(w_dff_B_nKF7123N6_1),.clk(gclk));
	jdff dff_B_Ll9sTDLV6_1(.din(w_dff_B_nKF7123N6_1),.dout(w_dff_B_Ll9sTDLV6_1),.clk(gclk));
	jdff dff_B_UiPn8pnG6_1(.din(w_dff_B_Ll9sTDLV6_1),.dout(w_dff_B_UiPn8pnG6_1),.clk(gclk));
	jdff dff_B_B3QeUWtN6_1(.din(w_dff_B_UiPn8pnG6_1),.dout(w_dff_B_B3QeUWtN6_1),.clk(gclk));
	jdff dff_B_jjvuWWT53_1(.din(w_dff_B_B3QeUWtN6_1),.dout(w_dff_B_jjvuWWT53_1),.clk(gclk));
	jdff dff_B_Cy24TzKo4_1(.din(w_dff_B_jjvuWWT53_1),.dout(w_dff_B_Cy24TzKo4_1),.clk(gclk));
	jdff dff_B_AvrJc9Fh3_1(.din(w_dff_B_Cy24TzKo4_1),.dout(w_dff_B_AvrJc9Fh3_1),.clk(gclk));
	jdff dff_B_7P7v1f2R5_1(.din(w_dff_B_AvrJc9Fh3_1),.dout(w_dff_B_7P7v1f2R5_1),.clk(gclk));
	jdff dff_B_Ftur8imG0_1(.din(w_dff_B_7P7v1f2R5_1),.dout(w_dff_B_Ftur8imG0_1),.clk(gclk));
	jdff dff_B_EuNF3oqt9_1(.din(w_dff_B_Ftur8imG0_1),.dout(w_dff_B_EuNF3oqt9_1),.clk(gclk));
	jdff dff_B_ROre4ehw0_1(.din(w_dff_B_EuNF3oqt9_1),.dout(w_dff_B_ROre4ehw0_1),.clk(gclk));
	jdff dff_B_Icv5Cas06_1(.din(w_dff_B_ROre4ehw0_1),.dout(w_dff_B_Icv5Cas06_1),.clk(gclk));
	jdff dff_B_6C3O9f618_1(.din(w_dff_B_Icv5Cas06_1),.dout(w_dff_B_6C3O9f618_1),.clk(gclk));
	jdff dff_B_rtFAHHBq0_1(.din(w_dff_B_6C3O9f618_1),.dout(w_dff_B_rtFAHHBq0_1),.clk(gclk));
	jdff dff_B_SUPdgmT26_1(.din(w_dff_B_rtFAHHBq0_1),.dout(w_dff_B_SUPdgmT26_1),.clk(gclk));
	jdff dff_B_HWA83ljg1_1(.din(w_dff_B_SUPdgmT26_1),.dout(w_dff_B_HWA83ljg1_1),.clk(gclk));
	jdff dff_B_3tb95YT87_1(.din(w_dff_B_HWA83ljg1_1),.dout(w_dff_B_3tb95YT87_1),.clk(gclk));
	jdff dff_B_QlWV5ZWu3_1(.din(w_dff_B_3tb95YT87_1),.dout(w_dff_B_QlWV5ZWu3_1),.clk(gclk));
	jdff dff_B_QYVvlqZl4_1(.din(w_dff_B_QlWV5ZWu3_1),.dout(w_dff_B_QYVvlqZl4_1),.clk(gclk));
	jdff dff_B_tPk13MuO0_1(.din(w_dff_B_QYVvlqZl4_1),.dout(w_dff_B_tPk13MuO0_1),.clk(gclk));
	jdff dff_B_NoJYw5590_1(.din(w_dff_B_tPk13MuO0_1),.dout(w_dff_B_NoJYw5590_1),.clk(gclk));
	jdff dff_B_NfP8PkSF3_1(.din(w_dff_B_NoJYw5590_1),.dout(w_dff_B_NfP8PkSF3_1),.clk(gclk));
	jdff dff_B_tQwdKdFd9_1(.din(w_dff_B_NfP8PkSF3_1),.dout(w_dff_B_tQwdKdFd9_1),.clk(gclk));
	jdff dff_B_t68SnBns4_1(.din(w_dff_B_tQwdKdFd9_1),.dout(w_dff_B_t68SnBns4_1),.clk(gclk));
	jdff dff_B_5eOFGvez3_1(.din(w_dff_B_t68SnBns4_1),.dout(w_dff_B_5eOFGvez3_1),.clk(gclk));
	jdff dff_B_EiwBf9Ie5_1(.din(w_dff_B_5eOFGvez3_1),.dout(w_dff_B_EiwBf9Ie5_1),.clk(gclk));
	jdff dff_B_cp3TvIVf9_1(.din(w_dff_B_EiwBf9Ie5_1),.dout(w_dff_B_cp3TvIVf9_1),.clk(gclk));
	jdff dff_B_YUC97WWG0_1(.din(w_dff_B_cp3TvIVf9_1),.dout(w_dff_B_YUC97WWG0_1),.clk(gclk));
	jdff dff_B_PXBcDd5b3_1(.din(w_dff_B_YUC97WWG0_1),.dout(w_dff_B_PXBcDd5b3_1),.clk(gclk));
	jdff dff_B_hsZqMFhJ3_1(.din(w_dff_B_PXBcDd5b3_1),.dout(w_dff_B_hsZqMFhJ3_1),.clk(gclk));
	jdff dff_B_bqNHNd9T7_1(.din(w_dff_B_hsZqMFhJ3_1),.dout(w_dff_B_bqNHNd9T7_1),.clk(gclk));
	jdff dff_B_R6d7TecP0_1(.din(w_dff_B_bqNHNd9T7_1),.dout(w_dff_B_R6d7TecP0_1),.clk(gclk));
	jdff dff_B_IFujLWY08_1(.din(w_dff_B_R6d7TecP0_1),.dout(w_dff_B_IFujLWY08_1),.clk(gclk));
	jdff dff_B_xMYa2SRa8_1(.din(w_dff_B_IFujLWY08_1),.dout(w_dff_B_xMYa2SRa8_1),.clk(gclk));
	jdff dff_B_oCldZxq23_1(.din(n830),.dout(w_dff_B_oCldZxq23_1),.clk(gclk));
	jdff dff_B_IGGrZXnp3_1(.din(w_dff_B_oCldZxq23_1),.dout(w_dff_B_IGGrZXnp3_1),.clk(gclk));
	jdff dff_B_CTGbThQI0_1(.din(w_dff_B_IGGrZXnp3_1),.dout(w_dff_B_CTGbThQI0_1),.clk(gclk));
	jdff dff_B_s79fFjKv1_1(.din(w_dff_B_CTGbThQI0_1),.dout(w_dff_B_s79fFjKv1_1),.clk(gclk));
	jdff dff_B_REH0IWYZ2_1(.din(w_dff_B_s79fFjKv1_1),.dout(w_dff_B_REH0IWYZ2_1),.clk(gclk));
	jdff dff_B_083CD5wE9_1(.din(w_dff_B_REH0IWYZ2_1),.dout(w_dff_B_083CD5wE9_1),.clk(gclk));
	jdff dff_B_VSl1wgOi2_1(.din(w_dff_B_083CD5wE9_1),.dout(w_dff_B_VSl1wgOi2_1),.clk(gclk));
	jdff dff_B_aIONJ2mi4_1(.din(w_dff_B_VSl1wgOi2_1),.dout(w_dff_B_aIONJ2mi4_1),.clk(gclk));
	jdff dff_B_abvVIJ2j0_1(.din(w_dff_B_aIONJ2mi4_1),.dout(w_dff_B_abvVIJ2j0_1),.clk(gclk));
	jdff dff_B_0Y8Nd7JK9_1(.din(w_dff_B_abvVIJ2j0_1),.dout(w_dff_B_0Y8Nd7JK9_1),.clk(gclk));
	jdff dff_B_vwbuSnOT1_1(.din(w_dff_B_0Y8Nd7JK9_1),.dout(w_dff_B_vwbuSnOT1_1),.clk(gclk));
	jdff dff_B_7le6HbYy0_1(.din(w_dff_B_vwbuSnOT1_1),.dout(w_dff_B_7le6HbYy0_1),.clk(gclk));
	jdff dff_B_UMLSg4MG9_1(.din(w_dff_B_7le6HbYy0_1),.dout(w_dff_B_UMLSg4MG9_1),.clk(gclk));
	jdff dff_B_Js5upuCB5_1(.din(w_dff_B_UMLSg4MG9_1),.dout(w_dff_B_Js5upuCB5_1),.clk(gclk));
	jdff dff_B_xsZlMiFw6_1(.din(w_dff_B_Js5upuCB5_1),.dout(w_dff_B_xsZlMiFw6_1),.clk(gclk));
	jdff dff_B_tCrQe8HZ1_1(.din(w_dff_B_xsZlMiFw6_1),.dout(w_dff_B_tCrQe8HZ1_1),.clk(gclk));
	jdff dff_B_JboN2GVL0_1(.din(w_dff_B_tCrQe8HZ1_1),.dout(w_dff_B_JboN2GVL0_1),.clk(gclk));
	jdff dff_B_VyhYR3BZ3_1(.din(w_dff_B_JboN2GVL0_1),.dout(w_dff_B_VyhYR3BZ3_1),.clk(gclk));
	jdff dff_B_aHGbkyCo1_1(.din(w_dff_B_VyhYR3BZ3_1),.dout(w_dff_B_aHGbkyCo1_1),.clk(gclk));
	jdff dff_B_3QxYAQfJ2_1(.din(w_dff_B_aHGbkyCo1_1),.dout(w_dff_B_3QxYAQfJ2_1),.clk(gclk));
	jdff dff_B_zLHK66928_1(.din(w_dff_B_3QxYAQfJ2_1),.dout(w_dff_B_zLHK66928_1),.clk(gclk));
	jdff dff_B_3BYEE1pX4_1(.din(w_dff_B_zLHK66928_1),.dout(w_dff_B_3BYEE1pX4_1),.clk(gclk));
	jdff dff_B_9BFhlPnb4_1(.din(w_dff_B_3BYEE1pX4_1),.dout(w_dff_B_9BFhlPnb4_1),.clk(gclk));
	jdff dff_B_AP6uzT607_1(.din(w_dff_B_9BFhlPnb4_1),.dout(w_dff_B_AP6uzT607_1),.clk(gclk));
	jdff dff_B_DnPi3aFF2_1(.din(w_dff_B_AP6uzT607_1),.dout(w_dff_B_DnPi3aFF2_1),.clk(gclk));
	jdff dff_B_jUOIzjKU2_1(.din(w_dff_B_DnPi3aFF2_1),.dout(w_dff_B_jUOIzjKU2_1),.clk(gclk));
	jdff dff_B_EUCmrPbZ2_1(.din(w_dff_B_jUOIzjKU2_1),.dout(w_dff_B_EUCmrPbZ2_1),.clk(gclk));
	jdff dff_B_RdmUctx22_1(.din(w_dff_B_EUCmrPbZ2_1),.dout(w_dff_B_RdmUctx22_1),.clk(gclk));
	jdff dff_B_oZkFp8qa8_1(.din(w_dff_B_RdmUctx22_1),.dout(w_dff_B_oZkFp8qa8_1),.clk(gclk));
	jdff dff_B_pWo908Su2_1(.din(w_dff_B_oZkFp8qa8_1),.dout(w_dff_B_pWo908Su2_1),.clk(gclk));
	jdff dff_B_hTbA170c1_1(.din(w_dff_B_pWo908Su2_1),.dout(w_dff_B_hTbA170c1_1),.clk(gclk));
	jdff dff_B_4aWxsDc90_1(.din(w_dff_B_hTbA170c1_1),.dout(w_dff_B_4aWxsDc90_1),.clk(gclk));
	jdff dff_B_91vhNdIB6_1(.din(w_dff_B_4aWxsDc90_1),.dout(w_dff_B_91vhNdIB6_1),.clk(gclk));
	jdff dff_B_94Tj5YPh4_1(.din(w_dff_B_91vhNdIB6_1),.dout(w_dff_B_94Tj5YPh4_1),.clk(gclk));
	jdff dff_B_UQjdE8xZ5_1(.din(w_dff_B_94Tj5YPh4_1),.dout(w_dff_B_UQjdE8xZ5_1),.clk(gclk));
	jdff dff_B_VnsM0W395_1(.din(w_dff_B_UQjdE8xZ5_1),.dout(w_dff_B_VnsM0W395_1),.clk(gclk));
	jdff dff_B_wdDfIAoD4_1(.din(w_dff_B_VnsM0W395_1),.dout(w_dff_B_wdDfIAoD4_1),.clk(gclk));
	jdff dff_B_Ni3DAazg6_1(.din(w_dff_B_wdDfIAoD4_1),.dout(w_dff_B_Ni3DAazg6_1),.clk(gclk));
	jdff dff_B_AcOt0G3U1_1(.din(w_dff_B_Ni3DAazg6_1),.dout(w_dff_B_AcOt0G3U1_1),.clk(gclk));
	jdff dff_B_Njn7T5vJ0_1(.din(w_dff_B_AcOt0G3U1_1),.dout(w_dff_B_Njn7T5vJ0_1),.clk(gclk));
	jdff dff_B_FDPn5Wpe1_1(.din(w_dff_B_Njn7T5vJ0_1),.dout(w_dff_B_FDPn5Wpe1_1),.clk(gclk));
	jdff dff_B_DFYNvs9J6_1(.din(w_dff_B_FDPn5Wpe1_1),.dout(w_dff_B_DFYNvs9J6_1),.clk(gclk));
	jdff dff_B_eG6R2dfb6_1(.din(w_dff_B_DFYNvs9J6_1),.dout(w_dff_B_eG6R2dfb6_1),.clk(gclk));
	jdff dff_B_nYPmOVXp3_0(.din(n1327),.dout(w_dff_B_nYPmOVXp3_0),.clk(gclk));
	jdff dff_B_h2NQdNi83_1(.din(n1842),.dout(w_dff_B_h2NQdNi83_1),.clk(gclk));
	jdff dff_B_w6xAud9Y6_1(.din(w_dff_B_h2NQdNi83_1),.dout(w_dff_B_w6xAud9Y6_1),.clk(gclk));
	jdff dff_B_j1HUws5y5_1(.din(w_dff_B_w6xAud9Y6_1),.dout(w_dff_B_j1HUws5y5_1),.clk(gclk));
	jdff dff_B_weuFHwps7_1(.din(w_dff_B_j1HUws5y5_1),.dout(w_dff_B_weuFHwps7_1),.clk(gclk));
	jdff dff_B_K4gMSjdJ2_1(.din(w_dff_B_weuFHwps7_1),.dout(w_dff_B_K4gMSjdJ2_1),.clk(gclk));
	jdff dff_B_UK1pMBul3_1(.din(w_dff_B_K4gMSjdJ2_1),.dout(w_dff_B_UK1pMBul3_1),.clk(gclk));
	jdff dff_B_dpAYw9U66_1(.din(w_dff_B_UK1pMBul3_1),.dout(w_dff_B_dpAYw9U66_1),.clk(gclk));
	jdff dff_B_3FPqNqRg6_1(.din(w_dff_B_dpAYw9U66_1),.dout(w_dff_B_3FPqNqRg6_1),.clk(gclk));
	jdff dff_B_RMgXq30i1_1(.din(w_dff_B_3FPqNqRg6_1),.dout(w_dff_B_RMgXq30i1_1),.clk(gclk));
	jdff dff_B_GuIkOsrU9_1(.din(w_dff_B_RMgXq30i1_1),.dout(w_dff_B_GuIkOsrU9_1),.clk(gclk));
	jdff dff_B_eOPWVIyh9_1(.din(w_dff_B_GuIkOsrU9_1),.dout(w_dff_B_eOPWVIyh9_1),.clk(gclk));
	jdff dff_B_98YfWaMd6_1(.din(w_dff_B_eOPWVIyh9_1),.dout(w_dff_B_98YfWaMd6_1),.clk(gclk));
	jdff dff_B_AJQXN7UJ4_1(.din(w_dff_B_98YfWaMd6_1),.dout(w_dff_B_AJQXN7UJ4_1),.clk(gclk));
	jdff dff_B_39OHMP0W1_0(.din(n1850),.dout(w_dff_B_39OHMP0W1_0),.clk(gclk));
	jdff dff_B_OUfenZMD6_0(.din(w_dff_B_39OHMP0W1_0),.dout(w_dff_B_OUfenZMD6_0),.clk(gclk));
	jdff dff_B_L6Be0ODT9_0(.din(w_dff_B_OUfenZMD6_0),.dout(w_dff_B_L6Be0ODT9_0),.clk(gclk));
	jdff dff_B_Zy4gqZv55_0(.din(w_dff_B_L6Be0ODT9_0),.dout(w_dff_B_Zy4gqZv55_0),.clk(gclk));
	jdff dff_B_15S0DRQx3_0(.din(w_dff_B_Zy4gqZv55_0),.dout(w_dff_B_15S0DRQx3_0),.clk(gclk));
	jdff dff_B_NGHghf4S2_0(.din(w_dff_B_15S0DRQx3_0),.dout(w_dff_B_NGHghf4S2_0),.clk(gclk));
	jdff dff_B_yATPcVva5_0(.din(w_dff_B_NGHghf4S2_0),.dout(w_dff_B_yATPcVva5_0),.clk(gclk));
	jdff dff_B_P11wpji41_0(.din(w_dff_B_yATPcVva5_0),.dout(w_dff_B_P11wpji41_0),.clk(gclk));
	jdff dff_B_xYQC0U1N6_0(.din(w_dff_B_P11wpji41_0),.dout(w_dff_B_xYQC0U1N6_0),.clk(gclk));
	jdff dff_B_r8nRu9jp0_0(.din(w_dff_B_xYQC0U1N6_0),.dout(w_dff_B_r8nRu9jp0_0),.clk(gclk));
	jdff dff_B_6I7wTHAp0_0(.din(w_dff_B_r8nRu9jp0_0),.dout(w_dff_B_6I7wTHAp0_0),.clk(gclk));
	jdff dff_A_ut6G07172_0(.dout(w_n1849_0[0]),.din(w_dff_A_ut6G07172_0),.clk(gclk));
	jdff dff_A_j8oWk5Pk2_0(.dout(w_dff_A_ut6G07172_0),.din(w_dff_A_j8oWk5Pk2_0),.clk(gclk));
	jdff dff_A_4eV7sBfX8_0(.dout(w_dff_A_j8oWk5Pk2_0),.din(w_dff_A_4eV7sBfX8_0),.clk(gclk));
	jdff dff_A_2MoJfxAt0_0(.dout(w_dff_A_4eV7sBfX8_0),.din(w_dff_A_2MoJfxAt0_0),.clk(gclk));
	jdff dff_A_VCXPxjPL6_0(.dout(w_dff_A_2MoJfxAt0_0),.din(w_dff_A_VCXPxjPL6_0),.clk(gclk));
	jdff dff_A_EwPuKEHs2_0(.dout(w_dff_A_VCXPxjPL6_0),.din(w_dff_A_EwPuKEHs2_0),.clk(gclk));
	jdff dff_A_zj2c6nf41_0(.dout(w_dff_A_EwPuKEHs2_0),.din(w_dff_A_zj2c6nf41_0),.clk(gclk));
	jdff dff_A_ZhxcM4KJ4_0(.dout(w_dff_A_zj2c6nf41_0),.din(w_dff_A_ZhxcM4KJ4_0),.clk(gclk));
	jdff dff_A_lugix02b7_0(.dout(w_dff_A_ZhxcM4KJ4_0),.din(w_dff_A_lugix02b7_0),.clk(gclk));
	jdff dff_A_IPF9IkbT3_0(.dout(w_dff_A_lugix02b7_0),.din(w_dff_A_IPF9IkbT3_0),.clk(gclk));
	jdff dff_A_284Si4af7_0(.dout(w_dff_A_IPF9IkbT3_0),.din(w_dff_A_284Si4af7_0),.clk(gclk));
	jdff dff_A_QBk0R33Z3_0(.dout(w_dff_A_284Si4af7_0),.din(w_dff_A_QBk0R33Z3_0),.clk(gclk));
	jdff dff_B_xVnw1T4P0_1(.din(n1839),.dout(w_dff_B_xVnw1T4P0_1),.clk(gclk));
	jdff dff_B_WeG7aV7r0_1(.din(w_dff_B_xVnw1T4P0_1),.dout(w_dff_B_WeG7aV7r0_1),.clk(gclk));
	jdff dff_B_ge5YKwtn3_2(.din(n1838),.dout(w_dff_B_ge5YKwtn3_2),.clk(gclk));
	jdff dff_B_uOnjh6FF0_2(.din(w_dff_B_ge5YKwtn3_2),.dout(w_dff_B_uOnjh6FF0_2),.clk(gclk));
	jdff dff_B_7dltARmO9_2(.din(w_dff_B_uOnjh6FF0_2),.dout(w_dff_B_7dltARmO9_2),.clk(gclk));
	jdff dff_B_dYqFSJCv4_2(.din(w_dff_B_7dltARmO9_2),.dout(w_dff_B_dYqFSJCv4_2),.clk(gclk));
	jdff dff_B_hDWLPYSj5_2(.din(w_dff_B_dYqFSJCv4_2),.dout(w_dff_B_hDWLPYSj5_2),.clk(gclk));
	jdff dff_B_ktoieRTt7_2(.din(w_dff_B_hDWLPYSj5_2),.dout(w_dff_B_ktoieRTt7_2),.clk(gclk));
	jdff dff_B_eGcA9lNu1_2(.din(w_dff_B_ktoieRTt7_2),.dout(w_dff_B_eGcA9lNu1_2),.clk(gclk));
	jdff dff_B_GLCtRJhO2_2(.din(w_dff_B_eGcA9lNu1_2),.dout(w_dff_B_GLCtRJhO2_2),.clk(gclk));
	jdff dff_B_UhUHDKJs4_2(.din(w_dff_B_GLCtRJhO2_2),.dout(w_dff_B_UhUHDKJs4_2),.clk(gclk));
	jdff dff_B_v8rodcin4_2(.din(w_dff_B_UhUHDKJs4_2),.dout(w_dff_B_v8rodcin4_2),.clk(gclk));
	jdff dff_B_9D2a0kP39_2(.din(w_dff_B_v8rodcin4_2),.dout(w_dff_B_9D2a0kP39_2),.clk(gclk));
	jdff dff_B_IRruBjsc7_2(.din(w_dff_B_9D2a0kP39_2),.dout(w_dff_B_IRruBjsc7_2),.clk(gclk));
	jdff dff_B_9SBKtdGh8_2(.din(w_dff_B_IRruBjsc7_2),.dout(w_dff_B_9SBKtdGh8_2),.clk(gclk));
	jdff dff_B_MCcCQBYY6_2(.din(w_dff_B_9SBKtdGh8_2),.dout(w_dff_B_MCcCQBYY6_2),.clk(gclk));
	jdff dff_B_HZ0SNEbB3_2(.din(w_dff_B_MCcCQBYY6_2),.dout(w_dff_B_HZ0SNEbB3_2),.clk(gclk));
	jdff dff_B_xsA2ur2w2_2(.din(w_dff_B_HZ0SNEbB3_2),.dout(w_dff_B_xsA2ur2w2_2),.clk(gclk));
	jdff dff_B_ZfUXriGL6_2(.din(w_dff_B_xsA2ur2w2_2),.dout(w_dff_B_ZfUXriGL6_2),.clk(gclk));
	jdff dff_B_ZyGa1XKK1_2(.din(w_dff_B_ZfUXriGL6_2),.dout(w_dff_B_ZyGa1XKK1_2),.clk(gclk));
	jdff dff_B_noLV7L8v9_2(.din(w_dff_B_ZyGa1XKK1_2),.dout(w_dff_B_noLV7L8v9_2),.clk(gclk));
	jdff dff_B_pwctVWsi5_2(.din(w_dff_B_noLV7L8v9_2),.dout(w_dff_B_pwctVWsi5_2),.clk(gclk));
	jdff dff_B_ALlT3D7p5_2(.din(w_dff_B_pwctVWsi5_2),.dout(w_dff_B_ALlT3D7p5_2),.clk(gclk));
	jdff dff_B_9zlQwrjG4_2(.din(w_dff_B_ALlT3D7p5_2),.dout(w_dff_B_9zlQwrjG4_2),.clk(gclk));
	jdff dff_B_5Hh2I43g5_2(.din(w_dff_B_9zlQwrjG4_2),.dout(w_dff_B_5Hh2I43g5_2),.clk(gclk));
	jdff dff_B_3Z2Abyrm9_2(.din(w_dff_B_5Hh2I43g5_2),.dout(w_dff_B_3Z2Abyrm9_2),.clk(gclk));
	jdff dff_B_QVE63Xpr3_2(.din(w_dff_B_3Z2Abyrm9_2),.dout(w_dff_B_QVE63Xpr3_2),.clk(gclk));
	jdff dff_B_gMekOidd8_2(.din(w_dff_B_QVE63Xpr3_2),.dout(w_dff_B_gMekOidd8_2),.clk(gclk));
	jdff dff_B_WlBOIRCB2_2(.din(w_dff_B_gMekOidd8_2),.dout(w_dff_B_WlBOIRCB2_2),.clk(gclk));
	jdff dff_B_bi5BQzpe5_2(.din(w_dff_B_WlBOIRCB2_2),.dout(w_dff_B_bi5BQzpe5_2),.clk(gclk));
	jdff dff_B_P91ieAHo2_2(.din(w_dff_B_bi5BQzpe5_2),.dout(w_dff_B_P91ieAHo2_2),.clk(gclk));
	jdff dff_B_wilyBuqr6_2(.din(w_dff_B_P91ieAHo2_2),.dout(w_dff_B_wilyBuqr6_2),.clk(gclk));
	jdff dff_B_ERYonw4I7_2(.din(w_dff_B_wilyBuqr6_2),.dout(w_dff_B_ERYonw4I7_2),.clk(gclk));
	jdff dff_B_Lr5wXo5p7_2(.din(w_dff_B_ERYonw4I7_2),.dout(w_dff_B_Lr5wXo5p7_2),.clk(gclk));
	jdff dff_B_P9xRXVrX5_2(.din(w_dff_B_Lr5wXo5p7_2),.dout(w_dff_B_P9xRXVrX5_2),.clk(gclk));
	jdff dff_B_ilDlmYak6_2(.din(w_dff_B_P9xRXVrX5_2),.dout(w_dff_B_ilDlmYak6_2),.clk(gclk));
	jdff dff_B_WwsrPN2o0_2(.din(w_dff_B_ilDlmYak6_2),.dout(w_dff_B_WwsrPN2o0_2),.clk(gclk));
	jdff dff_B_13jMJ3xx1_2(.din(w_dff_B_WwsrPN2o0_2),.dout(w_dff_B_13jMJ3xx1_2),.clk(gclk));
	jdff dff_B_JRJiaY1R1_2(.din(w_dff_B_13jMJ3xx1_2),.dout(w_dff_B_JRJiaY1R1_2),.clk(gclk));
	jdff dff_B_yH53UUPr2_2(.din(w_dff_B_JRJiaY1R1_2),.dout(w_dff_B_yH53UUPr2_2),.clk(gclk));
	jdff dff_B_2m82q0HC0_2(.din(w_dff_B_yH53UUPr2_2),.dout(w_dff_B_2m82q0HC0_2),.clk(gclk));
	jdff dff_B_uQcGInwi9_2(.din(w_dff_B_2m82q0HC0_2),.dout(w_dff_B_uQcGInwi9_2),.clk(gclk));
	jdff dff_B_nZrOZltL0_2(.din(w_dff_B_uQcGInwi9_2),.dout(w_dff_B_nZrOZltL0_2),.clk(gclk));
	jdff dff_B_etKkFuI77_2(.din(w_dff_B_nZrOZltL0_2),.dout(w_dff_B_etKkFuI77_2),.clk(gclk));
	jdff dff_B_1fFlJiSp1_2(.din(w_dff_B_etKkFuI77_2),.dout(w_dff_B_1fFlJiSp1_2),.clk(gclk));
	jdff dff_B_Ttqu1gge7_2(.din(w_dff_B_1fFlJiSp1_2),.dout(w_dff_B_Ttqu1gge7_2),.clk(gclk));
	jdff dff_B_P0vgnwCv1_2(.din(w_dff_B_Ttqu1gge7_2),.dout(w_dff_B_P0vgnwCv1_2),.clk(gclk));
	jdff dff_B_voaJivia8_2(.din(w_dff_B_P0vgnwCv1_2),.dout(w_dff_B_voaJivia8_2),.clk(gclk));
	jdff dff_B_Kk9wTNeM2_2(.din(w_dff_B_voaJivia8_2),.dout(w_dff_B_Kk9wTNeM2_2),.clk(gclk));
	jdff dff_B_18GxfdaB7_2(.din(w_dff_B_Kk9wTNeM2_2),.dout(w_dff_B_18GxfdaB7_2),.clk(gclk));
	jdff dff_B_LyHkaUR49_2(.din(w_dff_B_18GxfdaB7_2),.dout(w_dff_B_LyHkaUR49_2),.clk(gclk));
	jdff dff_B_oIOR0dmo3_2(.din(w_dff_B_LyHkaUR49_2),.dout(w_dff_B_oIOR0dmo3_2),.clk(gclk));
	jdff dff_B_Iz8tKzEp8_2(.din(w_dff_B_oIOR0dmo3_2),.dout(w_dff_B_Iz8tKzEp8_2),.clk(gclk));
	jdff dff_B_shPZTjE78_2(.din(w_dff_B_Iz8tKzEp8_2),.dout(w_dff_B_shPZTjE78_2),.clk(gclk));
	jdff dff_B_A68aUUPC3_2(.din(w_dff_B_shPZTjE78_2),.dout(w_dff_B_A68aUUPC3_2),.clk(gclk));
	jdff dff_B_jhc8pLKm4_2(.din(w_dff_B_A68aUUPC3_2),.dout(w_dff_B_jhc8pLKm4_2),.clk(gclk));
	jdff dff_B_U9JniUaH8_2(.din(w_dff_B_jhc8pLKm4_2),.dout(w_dff_B_U9JniUaH8_2),.clk(gclk));
	jdff dff_B_oJdtqV5z9_2(.din(w_dff_B_U9JniUaH8_2),.dout(w_dff_B_oJdtqV5z9_2),.clk(gclk));
	jdff dff_B_aYCWcGSM8_2(.din(w_dff_B_oJdtqV5z9_2),.dout(w_dff_B_aYCWcGSM8_2),.clk(gclk));
	jdff dff_B_COra2qfM4_2(.din(w_dff_B_aYCWcGSM8_2),.dout(w_dff_B_COra2qfM4_2),.clk(gclk));
	jdff dff_B_7UCxlYQc8_2(.din(w_dff_B_COra2qfM4_2),.dout(w_dff_B_7UCxlYQc8_2),.clk(gclk));
	jdff dff_B_Z1zRk0uY1_2(.din(w_dff_B_7UCxlYQc8_2),.dout(w_dff_B_Z1zRk0uY1_2),.clk(gclk));
	jdff dff_B_o9ACfJgY0_1(.din(n1845),.dout(w_dff_B_o9ACfJgY0_1),.clk(gclk));
	jdff dff_B_cPOEvITt8_1(.din(w_dff_B_o9ACfJgY0_1),.dout(w_dff_B_cPOEvITt8_1),.clk(gclk));
	jdff dff_B_XGwvc5G29_1(.din(w_dff_B_cPOEvITt8_1),.dout(w_dff_B_XGwvc5G29_1),.clk(gclk));
	jdff dff_B_o8h1KEpz0_1(.din(w_dff_B_XGwvc5G29_1),.dout(w_dff_B_o8h1KEpz0_1),.clk(gclk));
	jdff dff_B_FhFui9Xf6_1(.din(w_dff_B_o8h1KEpz0_1),.dout(w_dff_B_FhFui9Xf6_1),.clk(gclk));
	jdff dff_B_3RwaW1OU2_1(.din(w_dff_B_FhFui9Xf6_1),.dout(w_dff_B_3RwaW1OU2_1),.clk(gclk));
	jdff dff_B_qiqCAw8V7_1(.din(w_dff_B_3RwaW1OU2_1),.dout(w_dff_B_qiqCAw8V7_1),.clk(gclk));
	jdff dff_B_KkPLgnen0_1(.din(w_dff_B_qiqCAw8V7_1),.dout(w_dff_B_KkPLgnen0_1),.clk(gclk));
	jdff dff_B_Z9C3wXrT3_1(.din(w_dff_B_KkPLgnen0_1),.dout(w_dff_B_Z9C3wXrT3_1),.clk(gclk));
	jdff dff_B_cQs5ZD5z6_1(.din(w_dff_B_Z9C3wXrT3_1),.dout(w_dff_B_cQs5ZD5z6_1),.clk(gclk));
	jdff dff_B_axl2M9jY6_1(.din(w_dff_B_cQs5ZD5z6_1),.dout(w_dff_B_axl2M9jY6_1),.clk(gclk));
	jdff dff_B_d8alS8uA0_0(.din(n1846),.dout(w_dff_B_d8alS8uA0_0),.clk(gclk));
	jdff dff_B_5sHni9tO0_0(.din(w_dff_B_d8alS8uA0_0),.dout(w_dff_B_5sHni9tO0_0),.clk(gclk));
	jdff dff_B_1SUwnsbX8_0(.din(w_dff_B_5sHni9tO0_0),.dout(w_dff_B_1SUwnsbX8_0),.clk(gclk));
	jdff dff_B_mLEFg69p4_0(.din(w_dff_B_1SUwnsbX8_0),.dout(w_dff_B_mLEFg69p4_0),.clk(gclk));
	jdff dff_B_j4DcIPp68_0(.din(w_dff_B_mLEFg69p4_0),.dout(w_dff_B_j4DcIPp68_0),.clk(gclk));
	jdff dff_B_R1K5cPig8_0(.din(w_dff_B_j4DcIPp68_0),.dout(w_dff_B_R1K5cPig8_0),.clk(gclk));
	jdff dff_B_so0dxkMW6_0(.din(w_dff_B_R1K5cPig8_0),.dout(w_dff_B_so0dxkMW6_0),.clk(gclk));
	jdff dff_B_iEzwuLDR8_0(.din(w_dff_B_so0dxkMW6_0),.dout(w_dff_B_iEzwuLDR8_0),.clk(gclk));
	jdff dff_B_3jds2xVB2_0(.din(w_dff_B_iEzwuLDR8_0),.dout(w_dff_B_3jds2xVB2_0),.clk(gclk));
	jdff dff_B_SRiaM2L53_0(.din(w_dff_B_3jds2xVB2_0),.dout(w_dff_B_SRiaM2L53_0),.clk(gclk));
	jdff dff_A_7VKAsHle8_1(.dout(w_n1836_0[1]),.din(w_dff_A_7VKAsHle8_1),.clk(gclk));
	jdff dff_A_UZY1CrhJ1_1(.dout(w_dff_A_7VKAsHle8_1),.din(w_dff_A_UZY1CrhJ1_1),.clk(gclk));
	jdff dff_A_ViV3GljL8_1(.dout(w_dff_A_UZY1CrhJ1_1),.din(w_dff_A_ViV3GljL8_1),.clk(gclk));
	jdff dff_A_bcsj0KjH5_1(.dout(w_dff_A_ViV3GljL8_1),.din(w_dff_A_bcsj0KjH5_1),.clk(gclk));
	jdff dff_A_ijZFIdMx3_1(.dout(w_dff_A_bcsj0KjH5_1),.din(w_dff_A_ijZFIdMx3_1),.clk(gclk));
	jdff dff_A_0YRQSRgp9_1(.dout(w_dff_A_ijZFIdMx3_1),.din(w_dff_A_0YRQSRgp9_1),.clk(gclk));
	jdff dff_A_guFOqtuK1_1(.dout(w_dff_A_0YRQSRgp9_1),.din(w_dff_A_guFOqtuK1_1),.clk(gclk));
	jdff dff_A_87hGvDmh0_1(.dout(w_dff_A_guFOqtuK1_1),.din(w_dff_A_87hGvDmh0_1),.clk(gclk));
	jdff dff_A_Y9aOEV3y0_1(.dout(w_dff_A_87hGvDmh0_1),.din(w_dff_A_Y9aOEV3y0_1),.clk(gclk));
	jdff dff_A_YWfTYHQ56_1(.dout(w_dff_A_Y9aOEV3y0_1),.din(w_dff_A_YWfTYHQ56_1),.clk(gclk));
	jdff dff_A_0qrSNxvr5_1(.dout(w_dff_A_YWfTYHQ56_1),.din(w_dff_A_0qrSNxvr5_1),.clk(gclk));
	jdff dff_B_YEAzskLF4_1(.din(n1821),.dout(w_dff_B_YEAzskLF4_1),.clk(gclk));
	jdff dff_B_rMusndVY0_1(.din(w_dff_B_YEAzskLF4_1),.dout(w_dff_B_rMusndVY0_1),.clk(gclk));
	jdff dff_B_5gi6yClv4_1(.din(w_dff_B_rMusndVY0_1),.dout(w_dff_B_5gi6yClv4_1),.clk(gclk));
	jdff dff_B_ZmqVvHfH9_1(.din(w_dff_B_5gi6yClv4_1),.dout(w_dff_B_ZmqVvHfH9_1),.clk(gclk));
	jdff dff_B_V4WhLO7C5_1(.din(w_dff_B_ZmqVvHfH9_1),.dout(w_dff_B_V4WhLO7C5_1),.clk(gclk));
	jdff dff_B_BQPEx8m24_1(.din(w_dff_B_V4WhLO7C5_1),.dout(w_dff_B_BQPEx8m24_1),.clk(gclk));
	jdff dff_B_3kphcJ8Y9_1(.din(w_dff_B_BQPEx8m24_1),.dout(w_dff_B_3kphcJ8Y9_1),.clk(gclk));
	jdff dff_B_LZt5y3kR9_1(.din(w_dff_B_3kphcJ8Y9_1),.dout(w_dff_B_LZt5y3kR9_1),.clk(gclk));
	jdff dff_B_YEMg0A4Q4_1(.din(w_dff_B_LZt5y3kR9_1),.dout(w_dff_B_YEMg0A4Q4_1),.clk(gclk));
	jdff dff_B_6Hr1ygcP3_1(.din(w_dff_B_YEMg0A4Q4_1),.dout(w_dff_B_6Hr1ygcP3_1),.clk(gclk));
	jdff dff_B_bXC1YG0R2_1(.din(w_dff_B_6Hr1ygcP3_1),.dout(w_dff_B_bXC1YG0R2_1),.clk(gclk));
	jdff dff_B_ianbkAXR0_0(.din(n1822),.dout(w_dff_B_ianbkAXR0_0),.clk(gclk));
	jdff dff_B_BwzHQZTA6_0(.din(w_dff_B_ianbkAXR0_0),.dout(w_dff_B_BwzHQZTA6_0),.clk(gclk));
	jdff dff_B_0fFYEaoK5_0(.din(w_dff_B_BwzHQZTA6_0),.dout(w_dff_B_0fFYEaoK5_0),.clk(gclk));
	jdff dff_B_pdEzTE1M5_0(.din(w_dff_B_0fFYEaoK5_0),.dout(w_dff_B_pdEzTE1M5_0),.clk(gclk));
	jdff dff_B_EvVAsKtu6_0(.din(w_dff_B_pdEzTE1M5_0),.dout(w_dff_B_EvVAsKtu6_0),.clk(gclk));
	jdff dff_B_7A4DT3zN2_0(.din(w_dff_B_EvVAsKtu6_0),.dout(w_dff_B_7A4DT3zN2_0),.clk(gclk));
	jdff dff_B_qB0lheFZ7_0(.din(w_dff_B_7A4DT3zN2_0),.dout(w_dff_B_qB0lheFZ7_0),.clk(gclk));
	jdff dff_B_SoNZnL051_0(.din(w_dff_B_qB0lheFZ7_0),.dout(w_dff_B_SoNZnL051_0),.clk(gclk));
	jdff dff_B_67VTckUz2_0(.din(w_dff_B_SoNZnL051_0),.dout(w_dff_B_67VTckUz2_0),.clk(gclk));
	jdff dff_B_E29MaRkv1_0(.din(w_dff_B_67VTckUz2_0),.dout(w_dff_B_E29MaRkv1_0),.clk(gclk));
	jdff dff_A_Mj40EOBe6_1(.dout(w_n1817_0[1]),.din(w_dff_A_Mj40EOBe6_1),.clk(gclk));
	jdff dff_A_bsSvo46Y5_1(.dout(w_dff_A_Mj40EOBe6_1),.din(w_dff_A_bsSvo46Y5_1),.clk(gclk));
	jdff dff_A_HkR7Ylcm6_1(.dout(w_dff_A_bsSvo46Y5_1),.din(w_dff_A_HkR7Ylcm6_1),.clk(gclk));
	jdff dff_A_F3AxsMFG9_1(.dout(w_dff_A_HkR7Ylcm6_1),.din(w_dff_A_F3AxsMFG9_1),.clk(gclk));
	jdff dff_A_U20mPH2w6_1(.dout(w_dff_A_F3AxsMFG9_1),.din(w_dff_A_U20mPH2w6_1),.clk(gclk));
	jdff dff_A_H8pWA1CF4_1(.dout(w_dff_A_U20mPH2w6_1),.din(w_dff_A_H8pWA1CF4_1),.clk(gclk));
	jdff dff_A_yAmQbFP07_1(.dout(w_dff_A_H8pWA1CF4_1),.din(w_dff_A_yAmQbFP07_1),.clk(gclk));
	jdff dff_A_sKtmNH8T0_1(.dout(w_dff_A_yAmQbFP07_1),.din(w_dff_A_sKtmNH8T0_1),.clk(gclk));
	jdff dff_A_xDVMtuT66_1(.dout(w_dff_A_sKtmNH8T0_1),.din(w_dff_A_xDVMtuT66_1),.clk(gclk));
	jdff dff_A_ScOg4b7Q9_1(.dout(w_dff_A_xDVMtuT66_1),.din(w_dff_A_ScOg4b7Q9_1),.clk(gclk));
	jdff dff_A_eIaV6tH83_1(.dout(w_dff_A_ScOg4b7Q9_1),.din(w_dff_A_eIaV6tH83_1),.clk(gclk));
	jdff dff_B_5YvjGBAs8_1(.din(n1795),.dout(w_dff_B_5YvjGBAs8_1),.clk(gclk));
	jdff dff_B_8UiDUOn22_1(.din(w_dff_B_5YvjGBAs8_1),.dout(w_dff_B_8UiDUOn22_1),.clk(gclk));
	jdff dff_B_bZ1rNLCr2_1(.din(w_dff_B_8UiDUOn22_1),.dout(w_dff_B_bZ1rNLCr2_1),.clk(gclk));
	jdff dff_B_ONt2Z9LH7_1(.din(w_dff_B_bZ1rNLCr2_1),.dout(w_dff_B_ONt2Z9LH7_1),.clk(gclk));
	jdff dff_B_t39CgGCb0_1(.din(w_dff_B_ONt2Z9LH7_1),.dout(w_dff_B_t39CgGCb0_1),.clk(gclk));
	jdff dff_B_zL86rSCx0_1(.din(w_dff_B_t39CgGCb0_1),.dout(w_dff_B_zL86rSCx0_1),.clk(gclk));
	jdff dff_B_q5XuGfCR8_1(.din(w_dff_B_zL86rSCx0_1),.dout(w_dff_B_q5XuGfCR8_1),.clk(gclk));
	jdff dff_B_G55bmCv26_1(.din(w_dff_B_q5XuGfCR8_1),.dout(w_dff_B_G55bmCv26_1),.clk(gclk));
	jdff dff_B_Eh9dYSzZ7_1(.din(w_dff_B_G55bmCv26_1),.dout(w_dff_B_Eh9dYSzZ7_1),.clk(gclk));
	jdff dff_B_d9jDqZ8E4_1(.din(w_dff_B_Eh9dYSzZ7_1),.dout(w_dff_B_d9jDqZ8E4_1),.clk(gclk));
	jdff dff_B_7um8b3989_1(.din(w_dff_B_d9jDqZ8E4_1),.dout(w_dff_B_7um8b3989_1),.clk(gclk));
	jdff dff_B_749dpsfz8_0(.din(n1796),.dout(w_dff_B_749dpsfz8_0),.clk(gclk));
	jdff dff_B_skbY2O4v8_0(.din(w_dff_B_749dpsfz8_0),.dout(w_dff_B_skbY2O4v8_0),.clk(gclk));
	jdff dff_B_DMlJozVD5_0(.din(w_dff_B_skbY2O4v8_0),.dout(w_dff_B_DMlJozVD5_0),.clk(gclk));
	jdff dff_B_fhmqYWYx6_0(.din(w_dff_B_DMlJozVD5_0),.dout(w_dff_B_fhmqYWYx6_0),.clk(gclk));
	jdff dff_B_GzG1hbKr7_0(.din(w_dff_B_fhmqYWYx6_0),.dout(w_dff_B_GzG1hbKr7_0),.clk(gclk));
	jdff dff_B_UidKZxkQ4_0(.din(w_dff_B_GzG1hbKr7_0),.dout(w_dff_B_UidKZxkQ4_0),.clk(gclk));
	jdff dff_B_1dzjzpZw2_0(.din(w_dff_B_UidKZxkQ4_0),.dout(w_dff_B_1dzjzpZw2_0),.clk(gclk));
	jdff dff_B_e3bYoBsL9_0(.din(w_dff_B_1dzjzpZw2_0),.dout(w_dff_B_e3bYoBsL9_0),.clk(gclk));
	jdff dff_B_MMAW9hxB9_0(.din(w_dff_B_e3bYoBsL9_0),.dout(w_dff_B_MMAW9hxB9_0),.clk(gclk));
	jdff dff_B_sqeRZOro5_0(.din(w_dff_B_MMAW9hxB9_0),.dout(w_dff_B_sqeRZOro5_0),.clk(gclk));
	jdff dff_A_mswBxS1X9_1(.dout(w_n1791_0[1]),.din(w_dff_A_mswBxS1X9_1),.clk(gclk));
	jdff dff_A_UeLFYQ4b1_1(.dout(w_dff_A_mswBxS1X9_1),.din(w_dff_A_UeLFYQ4b1_1),.clk(gclk));
	jdff dff_A_TYKipJmp5_1(.dout(w_dff_A_UeLFYQ4b1_1),.din(w_dff_A_TYKipJmp5_1),.clk(gclk));
	jdff dff_A_YL9q3rcN2_1(.dout(w_dff_A_TYKipJmp5_1),.din(w_dff_A_YL9q3rcN2_1),.clk(gclk));
	jdff dff_A_b5X0aJG49_1(.dout(w_dff_A_YL9q3rcN2_1),.din(w_dff_A_b5X0aJG49_1),.clk(gclk));
	jdff dff_A_Ok1SW55K5_1(.dout(w_dff_A_b5X0aJG49_1),.din(w_dff_A_Ok1SW55K5_1),.clk(gclk));
	jdff dff_A_t08ZGmFO9_1(.dout(w_dff_A_Ok1SW55K5_1),.din(w_dff_A_t08ZGmFO9_1),.clk(gclk));
	jdff dff_A_xhE2jIkx8_1(.dout(w_dff_A_t08ZGmFO9_1),.din(w_dff_A_xhE2jIkx8_1),.clk(gclk));
	jdff dff_A_xAT2xVsN4_1(.dout(w_dff_A_xhE2jIkx8_1),.din(w_dff_A_xAT2xVsN4_1),.clk(gclk));
	jdff dff_A_drFri1Aq6_1(.dout(w_dff_A_xAT2xVsN4_1),.din(w_dff_A_drFri1Aq6_1),.clk(gclk));
	jdff dff_A_IoAnXfgU6_1(.dout(w_dff_A_drFri1Aq6_1),.din(w_dff_A_IoAnXfgU6_1),.clk(gclk));
	jdff dff_B_arrQLrjA0_1(.din(n1762),.dout(w_dff_B_arrQLrjA0_1),.clk(gclk));
	jdff dff_B_wdj2zzep9_1(.din(w_dff_B_arrQLrjA0_1),.dout(w_dff_B_wdj2zzep9_1),.clk(gclk));
	jdff dff_B_cv8hbwiA3_1(.din(w_dff_B_wdj2zzep9_1),.dout(w_dff_B_cv8hbwiA3_1),.clk(gclk));
	jdff dff_B_mBMwSrKI0_1(.din(w_dff_B_cv8hbwiA3_1),.dout(w_dff_B_mBMwSrKI0_1),.clk(gclk));
	jdff dff_B_ZNrIb3Ob7_1(.din(w_dff_B_mBMwSrKI0_1),.dout(w_dff_B_ZNrIb3Ob7_1),.clk(gclk));
	jdff dff_B_62OmB0kE6_1(.din(w_dff_B_ZNrIb3Ob7_1),.dout(w_dff_B_62OmB0kE6_1),.clk(gclk));
	jdff dff_B_TC6QIwv07_1(.din(w_dff_B_62OmB0kE6_1),.dout(w_dff_B_TC6QIwv07_1),.clk(gclk));
	jdff dff_B_yQECvr7t1_1(.din(w_dff_B_TC6QIwv07_1),.dout(w_dff_B_yQECvr7t1_1),.clk(gclk));
	jdff dff_B_DYxvsUTe6_1(.din(w_dff_B_yQECvr7t1_1),.dout(w_dff_B_DYxvsUTe6_1),.clk(gclk));
	jdff dff_B_bg5QWs855_1(.din(w_dff_B_DYxvsUTe6_1),.dout(w_dff_B_bg5QWs855_1),.clk(gclk));
	jdff dff_B_yshrl5Ud5_1(.din(w_dff_B_bg5QWs855_1),.dout(w_dff_B_yshrl5Ud5_1),.clk(gclk));
	jdff dff_B_2rU6hWhb0_0(.din(n1763),.dout(w_dff_B_2rU6hWhb0_0),.clk(gclk));
	jdff dff_B_gCDpAbbi9_0(.din(w_dff_B_2rU6hWhb0_0),.dout(w_dff_B_gCDpAbbi9_0),.clk(gclk));
	jdff dff_B_4h9QGvdW3_0(.din(w_dff_B_gCDpAbbi9_0),.dout(w_dff_B_4h9QGvdW3_0),.clk(gclk));
	jdff dff_B_syhtqtz50_0(.din(w_dff_B_4h9QGvdW3_0),.dout(w_dff_B_syhtqtz50_0),.clk(gclk));
	jdff dff_B_DhS074Qe9_0(.din(w_dff_B_syhtqtz50_0),.dout(w_dff_B_DhS074Qe9_0),.clk(gclk));
	jdff dff_B_rfxAJ5Yw9_0(.din(w_dff_B_DhS074Qe9_0),.dout(w_dff_B_rfxAJ5Yw9_0),.clk(gclk));
	jdff dff_B_OkSZCMOR4_0(.din(w_dff_B_rfxAJ5Yw9_0),.dout(w_dff_B_OkSZCMOR4_0),.clk(gclk));
	jdff dff_B_OCfgNTLu2_0(.din(w_dff_B_OkSZCMOR4_0),.dout(w_dff_B_OCfgNTLu2_0),.clk(gclk));
	jdff dff_B_61oQJSTp8_0(.din(w_dff_B_OCfgNTLu2_0),.dout(w_dff_B_61oQJSTp8_0),.clk(gclk));
	jdff dff_B_W6zUBB6O9_0(.din(w_dff_B_61oQJSTp8_0),.dout(w_dff_B_W6zUBB6O9_0),.clk(gclk));
	jdff dff_A_mxwr8UYm7_1(.dout(w_n1758_0[1]),.din(w_dff_A_mxwr8UYm7_1),.clk(gclk));
	jdff dff_A_IFCPKTSb9_1(.dout(w_dff_A_mxwr8UYm7_1),.din(w_dff_A_IFCPKTSb9_1),.clk(gclk));
	jdff dff_A_t0TQDQ423_1(.dout(w_dff_A_IFCPKTSb9_1),.din(w_dff_A_t0TQDQ423_1),.clk(gclk));
	jdff dff_A_Btn4SYhf5_1(.dout(w_dff_A_t0TQDQ423_1),.din(w_dff_A_Btn4SYhf5_1),.clk(gclk));
	jdff dff_A_4uPoGXNf8_1(.dout(w_dff_A_Btn4SYhf5_1),.din(w_dff_A_4uPoGXNf8_1),.clk(gclk));
	jdff dff_A_kps6M7715_1(.dout(w_dff_A_4uPoGXNf8_1),.din(w_dff_A_kps6M7715_1),.clk(gclk));
	jdff dff_A_tqWCwPQ50_1(.dout(w_dff_A_kps6M7715_1),.din(w_dff_A_tqWCwPQ50_1),.clk(gclk));
	jdff dff_A_aFTLbqF16_1(.dout(w_dff_A_tqWCwPQ50_1),.din(w_dff_A_aFTLbqF16_1),.clk(gclk));
	jdff dff_A_B98nMDlS7_1(.dout(w_dff_A_aFTLbqF16_1),.din(w_dff_A_B98nMDlS7_1),.clk(gclk));
	jdff dff_A_cOOiRZiJ6_1(.dout(w_dff_A_B98nMDlS7_1),.din(w_dff_A_cOOiRZiJ6_1),.clk(gclk));
	jdff dff_A_3bR1yH9e9_1(.dout(w_dff_A_cOOiRZiJ6_1),.din(w_dff_A_3bR1yH9e9_1),.clk(gclk));
	jdff dff_B_WnJUfAew8_1(.din(n1722),.dout(w_dff_B_WnJUfAew8_1),.clk(gclk));
	jdff dff_B_Kj1H0aPJ0_1(.din(w_dff_B_WnJUfAew8_1),.dout(w_dff_B_Kj1H0aPJ0_1),.clk(gclk));
	jdff dff_B_L7PzYaCk1_1(.din(w_dff_B_Kj1H0aPJ0_1),.dout(w_dff_B_L7PzYaCk1_1),.clk(gclk));
	jdff dff_B_TYZClh2K1_1(.din(w_dff_B_L7PzYaCk1_1),.dout(w_dff_B_TYZClh2K1_1),.clk(gclk));
	jdff dff_B_0u6ciJRm1_1(.din(w_dff_B_TYZClh2K1_1),.dout(w_dff_B_0u6ciJRm1_1),.clk(gclk));
	jdff dff_B_2lCvsLXn6_1(.din(w_dff_B_0u6ciJRm1_1),.dout(w_dff_B_2lCvsLXn6_1),.clk(gclk));
	jdff dff_B_DjyO0dHN9_1(.din(w_dff_B_2lCvsLXn6_1),.dout(w_dff_B_DjyO0dHN9_1),.clk(gclk));
	jdff dff_B_UJGNFLuM7_1(.din(w_dff_B_DjyO0dHN9_1),.dout(w_dff_B_UJGNFLuM7_1),.clk(gclk));
	jdff dff_B_fWiL7Xtt8_1(.din(w_dff_B_UJGNFLuM7_1),.dout(w_dff_B_fWiL7Xtt8_1),.clk(gclk));
	jdff dff_B_q2RjPvxV1_1(.din(w_dff_B_fWiL7Xtt8_1),.dout(w_dff_B_q2RjPvxV1_1),.clk(gclk));
	jdff dff_B_XjLyrqrv9_1(.din(w_dff_B_q2RjPvxV1_1),.dout(w_dff_B_XjLyrqrv9_1),.clk(gclk));
	jdff dff_B_dC54bDG36_0(.din(n1723),.dout(w_dff_B_dC54bDG36_0),.clk(gclk));
	jdff dff_B_YhLA8U5Y5_0(.din(w_dff_B_dC54bDG36_0),.dout(w_dff_B_YhLA8U5Y5_0),.clk(gclk));
	jdff dff_B_EOwbEmdX9_0(.din(w_dff_B_YhLA8U5Y5_0),.dout(w_dff_B_EOwbEmdX9_0),.clk(gclk));
	jdff dff_B_XE0L8f0U6_0(.din(w_dff_B_EOwbEmdX9_0),.dout(w_dff_B_XE0L8f0U6_0),.clk(gclk));
	jdff dff_B_5gv2pbhi4_0(.din(w_dff_B_XE0L8f0U6_0),.dout(w_dff_B_5gv2pbhi4_0),.clk(gclk));
	jdff dff_B_cekxpdly7_0(.din(w_dff_B_5gv2pbhi4_0),.dout(w_dff_B_cekxpdly7_0),.clk(gclk));
	jdff dff_B_pL8ykWlX0_0(.din(w_dff_B_cekxpdly7_0),.dout(w_dff_B_pL8ykWlX0_0),.clk(gclk));
	jdff dff_B_46e03LDC6_0(.din(w_dff_B_pL8ykWlX0_0),.dout(w_dff_B_46e03LDC6_0),.clk(gclk));
	jdff dff_B_5CmIey8H7_0(.din(w_dff_B_46e03LDC6_0),.dout(w_dff_B_5CmIey8H7_0),.clk(gclk));
	jdff dff_A_u380fZG16_1(.dout(w_n1720_0[1]),.din(w_dff_A_u380fZG16_1),.clk(gclk));
	jdff dff_A_dayGIxwK3_1(.dout(w_dff_A_u380fZG16_1),.din(w_dff_A_dayGIxwK3_1),.clk(gclk));
	jdff dff_A_nnaOHHwf3_1(.dout(w_dff_A_dayGIxwK3_1),.din(w_dff_A_nnaOHHwf3_1),.clk(gclk));
	jdff dff_A_RLPkLiQf4_1(.dout(w_dff_A_nnaOHHwf3_1),.din(w_dff_A_RLPkLiQf4_1),.clk(gclk));
	jdff dff_A_mF3z3wDM0_1(.dout(w_dff_A_RLPkLiQf4_1),.din(w_dff_A_mF3z3wDM0_1),.clk(gclk));
	jdff dff_A_gtl5zLcf6_1(.dout(w_dff_A_mF3z3wDM0_1),.din(w_dff_A_gtl5zLcf6_1),.clk(gclk));
	jdff dff_A_rEqRhFPT8_1(.dout(w_dff_A_gtl5zLcf6_1),.din(w_dff_A_rEqRhFPT8_1),.clk(gclk));
	jdff dff_A_KnR9i2lp7_1(.dout(w_dff_A_rEqRhFPT8_1),.din(w_dff_A_KnR9i2lp7_1),.clk(gclk));
	jdff dff_A_FDqqWS4F2_1(.dout(w_dff_A_KnR9i2lp7_1),.din(w_dff_A_FDqqWS4F2_1),.clk(gclk));
	jdff dff_A_4SVq3Cyq9_1(.dout(w_dff_A_FDqqWS4F2_1),.din(w_dff_A_4SVq3Cyq9_1),.clk(gclk));
	jdff dff_B_MsVoWa3L2_1(.din(n1674),.dout(w_dff_B_MsVoWa3L2_1),.clk(gclk));
	jdff dff_B_60a7kRpr4_1(.din(w_dff_B_MsVoWa3L2_1),.dout(w_dff_B_60a7kRpr4_1),.clk(gclk));
	jdff dff_B_Np9BxNl36_1(.din(w_dff_B_60a7kRpr4_1),.dout(w_dff_B_Np9BxNl36_1),.clk(gclk));
	jdff dff_B_XlZxtOUp8_1(.din(w_dff_B_Np9BxNl36_1),.dout(w_dff_B_XlZxtOUp8_1),.clk(gclk));
	jdff dff_B_aAK0I0uV1_1(.din(w_dff_B_XlZxtOUp8_1),.dout(w_dff_B_aAK0I0uV1_1),.clk(gclk));
	jdff dff_B_YioF7NQx9_1(.din(w_dff_B_aAK0I0uV1_1),.dout(w_dff_B_YioF7NQx9_1),.clk(gclk));
	jdff dff_B_0Px2zpau2_1(.din(w_dff_B_YioF7NQx9_1),.dout(w_dff_B_0Px2zpau2_1),.clk(gclk));
	jdff dff_B_vY0YaZ6a4_1(.din(w_dff_B_0Px2zpau2_1),.dout(w_dff_B_vY0YaZ6a4_1),.clk(gclk));
	jdff dff_B_4qelXxch3_1(.din(w_dff_B_vY0YaZ6a4_1),.dout(w_dff_B_4qelXxch3_1),.clk(gclk));
	jdff dff_B_mtlvViN33_1(.din(w_dff_B_4qelXxch3_1),.dout(w_dff_B_mtlvViN33_1),.clk(gclk));
	jdff dff_B_liyKuP360_0(.din(n1675),.dout(w_dff_B_liyKuP360_0),.clk(gclk));
	jdff dff_B_szUbbBuD2_0(.din(w_dff_B_liyKuP360_0),.dout(w_dff_B_szUbbBuD2_0),.clk(gclk));
	jdff dff_B_sQKoR2ul9_0(.din(w_dff_B_szUbbBuD2_0),.dout(w_dff_B_sQKoR2ul9_0),.clk(gclk));
	jdff dff_B_jsPi28bt0_0(.din(w_dff_B_sQKoR2ul9_0),.dout(w_dff_B_jsPi28bt0_0),.clk(gclk));
	jdff dff_B_n3mW5Eo46_0(.din(w_dff_B_jsPi28bt0_0),.dout(w_dff_B_n3mW5Eo46_0),.clk(gclk));
	jdff dff_B_BlcJPBFe0_0(.din(w_dff_B_n3mW5Eo46_0),.dout(w_dff_B_BlcJPBFe0_0),.clk(gclk));
	jdff dff_B_6UsnmYeN3_0(.din(w_dff_B_BlcJPBFe0_0),.dout(w_dff_B_6UsnmYeN3_0),.clk(gclk));
	jdff dff_B_Tze7IZDs2_0(.din(w_dff_B_6UsnmYeN3_0),.dout(w_dff_B_Tze7IZDs2_0),.clk(gclk));
	jdff dff_A_hkeAjjSB2_1(.dout(w_n1672_0[1]),.din(w_dff_A_hkeAjjSB2_1),.clk(gclk));
	jdff dff_A_8YjD7zZi1_1(.dout(w_dff_A_hkeAjjSB2_1),.din(w_dff_A_8YjD7zZi1_1),.clk(gclk));
	jdff dff_A_5lkyAW9x8_1(.dout(w_dff_A_8YjD7zZi1_1),.din(w_dff_A_5lkyAW9x8_1),.clk(gclk));
	jdff dff_A_xBHAMgpt6_1(.dout(w_dff_A_5lkyAW9x8_1),.din(w_dff_A_xBHAMgpt6_1),.clk(gclk));
	jdff dff_A_HDJofp8d4_1(.dout(w_dff_A_xBHAMgpt6_1),.din(w_dff_A_HDJofp8d4_1),.clk(gclk));
	jdff dff_A_KwCiN0Sy0_1(.dout(w_dff_A_HDJofp8d4_1),.din(w_dff_A_KwCiN0Sy0_1),.clk(gclk));
	jdff dff_A_Hhxneuyj6_1(.dout(w_dff_A_KwCiN0Sy0_1),.din(w_dff_A_Hhxneuyj6_1),.clk(gclk));
	jdff dff_A_hzYJS89d0_1(.dout(w_dff_A_Hhxneuyj6_1),.din(w_dff_A_hzYJS89d0_1),.clk(gclk));
	jdff dff_A_PseeWV7o8_1(.dout(w_dff_A_hzYJS89d0_1),.din(w_dff_A_PseeWV7o8_1),.clk(gclk));
	jdff dff_B_a7YIOk8M8_1(.din(n1619),.dout(w_dff_B_a7YIOk8M8_1),.clk(gclk));
	jdff dff_B_dZbbqaue6_1(.din(w_dff_B_a7YIOk8M8_1),.dout(w_dff_B_dZbbqaue6_1),.clk(gclk));
	jdff dff_B_o19TEuSk0_1(.din(w_dff_B_dZbbqaue6_1),.dout(w_dff_B_o19TEuSk0_1),.clk(gclk));
	jdff dff_B_LU2YWc9d6_1(.din(w_dff_B_o19TEuSk0_1),.dout(w_dff_B_LU2YWc9d6_1),.clk(gclk));
	jdff dff_B_SAjuZs1F7_1(.din(w_dff_B_LU2YWc9d6_1),.dout(w_dff_B_SAjuZs1F7_1),.clk(gclk));
	jdff dff_B_kAZFaCcr0_1(.din(w_dff_B_SAjuZs1F7_1),.dout(w_dff_B_kAZFaCcr0_1),.clk(gclk));
	jdff dff_B_dhgKUgDp9_1(.din(w_dff_B_kAZFaCcr0_1),.dout(w_dff_B_dhgKUgDp9_1),.clk(gclk));
	jdff dff_B_vZYIiGeW8_1(.din(w_dff_B_dhgKUgDp9_1),.dout(w_dff_B_vZYIiGeW8_1),.clk(gclk));
	jdff dff_B_osgi03YI5_1(.din(w_dff_B_vZYIiGeW8_1),.dout(w_dff_B_osgi03YI5_1),.clk(gclk));
	jdff dff_B_ARhsUsw33_1(.din(w_dff_B_osgi03YI5_1),.dout(w_dff_B_ARhsUsw33_1),.clk(gclk));
	jdff dff_B_eqChqEf42_0(.din(n1620),.dout(w_dff_B_eqChqEf42_0),.clk(gclk));
	jdff dff_B_9xaitLE90_0(.din(w_dff_B_eqChqEf42_0),.dout(w_dff_B_9xaitLE90_0),.clk(gclk));
	jdff dff_B_5vca0cLj1_0(.din(w_dff_B_9xaitLE90_0),.dout(w_dff_B_5vca0cLj1_0),.clk(gclk));
	jdff dff_B_hxYnyNWb0_0(.din(w_dff_B_5vca0cLj1_0),.dout(w_dff_B_hxYnyNWb0_0),.clk(gclk));
	jdff dff_B_inrFCRUM7_0(.din(w_dff_B_hxYnyNWb0_0),.dout(w_dff_B_inrFCRUM7_0),.clk(gclk));
	jdff dff_B_eOcvstmW6_0(.din(w_dff_B_inrFCRUM7_0),.dout(w_dff_B_eOcvstmW6_0),.clk(gclk));
	jdff dff_B_32WcYKRw9_0(.din(w_dff_B_eOcvstmW6_0),.dout(w_dff_B_32WcYKRw9_0),.clk(gclk));
	jdff dff_B_6YQoVxFh5_0(.din(w_dff_B_32WcYKRw9_0),.dout(w_dff_B_6YQoVxFh5_0),.clk(gclk));
	jdff dff_A_mA5lx3FM3_1(.dout(w_n1617_0[1]),.din(w_dff_A_mA5lx3FM3_1),.clk(gclk));
	jdff dff_A_taLSbNYm3_1(.dout(w_dff_A_mA5lx3FM3_1),.din(w_dff_A_taLSbNYm3_1),.clk(gclk));
	jdff dff_A_DRq3fT7G6_1(.dout(w_dff_A_taLSbNYm3_1),.din(w_dff_A_DRq3fT7G6_1),.clk(gclk));
	jdff dff_A_dofAhVII2_1(.dout(w_dff_A_DRq3fT7G6_1),.din(w_dff_A_dofAhVII2_1),.clk(gclk));
	jdff dff_A_hfR7aPfM0_1(.dout(w_dff_A_dofAhVII2_1),.din(w_dff_A_hfR7aPfM0_1),.clk(gclk));
	jdff dff_A_SkuTR7Ef7_1(.dout(w_dff_A_hfR7aPfM0_1),.din(w_dff_A_SkuTR7Ef7_1),.clk(gclk));
	jdff dff_A_FJjl9Pkl0_1(.dout(w_dff_A_SkuTR7Ef7_1),.din(w_dff_A_FJjl9Pkl0_1),.clk(gclk));
	jdff dff_A_uRC3vwxj8_1(.dout(w_dff_A_FJjl9Pkl0_1),.din(w_dff_A_uRC3vwxj8_1),.clk(gclk));
	jdff dff_A_9NTLJcnU8_1(.dout(w_dff_A_uRC3vwxj8_1),.din(w_dff_A_9NTLJcnU8_1),.clk(gclk));
	jdff dff_B_H92v0Rrm3_1(.din(n1557),.dout(w_dff_B_H92v0Rrm3_1),.clk(gclk));
	jdff dff_B_8B6yT9DT0_1(.din(w_dff_B_H92v0Rrm3_1),.dout(w_dff_B_8B6yT9DT0_1),.clk(gclk));
	jdff dff_B_kG9W971c6_1(.din(w_dff_B_8B6yT9DT0_1),.dout(w_dff_B_kG9W971c6_1),.clk(gclk));
	jdff dff_B_ezsMz3ps2_1(.din(w_dff_B_kG9W971c6_1),.dout(w_dff_B_ezsMz3ps2_1),.clk(gclk));
	jdff dff_B_bQtBB8yb6_1(.din(w_dff_B_ezsMz3ps2_1),.dout(w_dff_B_bQtBB8yb6_1),.clk(gclk));
	jdff dff_B_N1gPcbpr7_1(.din(w_dff_B_bQtBB8yb6_1),.dout(w_dff_B_N1gPcbpr7_1),.clk(gclk));
	jdff dff_B_Xd7nkYJJ5_1(.din(w_dff_B_N1gPcbpr7_1),.dout(w_dff_B_Xd7nkYJJ5_1),.clk(gclk));
	jdff dff_B_EAv8BngY7_1(.din(w_dff_B_Xd7nkYJJ5_1),.dout(w_dff_B_EAv8BngY7_1),.clk(gclk));
	jdff dff_B_hhXVJfRN7_0(.din(n1558),.dout(w_dff_B_hhXVJfRN7_0),.clk(gclk));
	jdff dff_B_jOg8jmyr1_0(.din(w_dff_B_hhXVJfRN7_0),.dout(w_dff_B_jOg8jmyr1_0),.clk(gclk));
	jdff dff_B_ASlbXrhA5_0(.din(w_dff_B_jOg8jmyr1_0),.dout(w_dff_B_ASlbXrhA5_0),.clk(gclk));
	jdff dff_B_XW7fl4cO5_0(.din(w_dff_B_ASlbXrhA5_0),.dout(w_dff_B_XW7fl4cO5_0),.clk(gclk));
	jdff dff_B_htQ0YOcZ4_0(.din(w_dff_B_XW7fl4cO5_0),.dout(w_dff_B_htQ0YOcZ4_0),.clk(gclk));
	jdff dff_B_m0hmfefD1_0(.din(w_dff_B_htQ0YOcZ4_0),.dout(w_dff_B_m0hmfefD1_0),.clk(gclk));
	jdff dff_A_GarCRriD1_1(.dout(w_n1555_0[1]),.din(w_dff_A_GarCRriD1_1),.clk(gclk));
	jdff dff_A_TA1hEKgS4_1(.dout(w_dff_A_GarCRriD1_1),.din(w_dff_A_TA1hEKgS4_1),.clk(gclk));
	jdff dff_A_Qn41WNQI1_1(.dout(w_dff_A_TA1hEKgS4_1),.din(w_dff_A_Qn41WNQI1_1),.clk(gclk));
	jdff dff_A_IsTiWrYf3_1(.dout(w_dff_A_Qn41WNQI1_1),.din(w_dff_A_IsTiWrYf3_1),.clk(gclk));
	jdff dff_A_daiH8hST4_1(.dout(w_dff_A_IsTiWrYf3_1),.din(w_dff_A_daiH8hST4_1),.clk(gclk));
	jdff dff_A_OWyDLyKj7_1(.dout(w_dff_A_daiH8hST4_1),.din(w_dff_A_OWyDLyKj7_1),.clk(gclk));
	jdff dff_A_xmslFCKQ7_1(.dout(w_dff_A_OWyDLyKj7_1),.din(w_dff_A_xmslFCKQ7_1),.clk(gclk));
	jdff dff_B_atpQrkQn9_1(.din(n1488),.dout(w_dff_B_atpQrkQn9_1),.clk(gclk));
	jdff dff_B_s36uqheW1_1(.din(w_dff_B_atpQrkQn9_1),.dout(w_dff_B_s36uqheW1_1),.clk(gclk));
	jdff dff_B_JFKjl0bP0_1(.din(w_dff_B_s36uqheW1_1),.dout(w_dff_B_JFKjl0bP0_1),.clk(gclk));
	jdff dff_B_mcZUAll60_1(.din(w_dff_B_JFKjl0bP0_1),.dout(w_dff_B_mcZUAll60_1),.clk(gclk));
	jdff dff_B_FnujWyla8_1(.din(w_dff_B_mcZUAll60_1),.dout(w_dff_B_FnujWyla8_1),.clk(gclk));
	jdff dff_B_D2ZhCCaW9_1(.din(w_dff_B_FnujWyla8_1),.dout(w_dff_B_D2ZhCCaW9_1),.clk(gclk));
	jdff dff_B_KasjwAkM9_1(.din(w_dff_B_D2ZhCCaW9_1),.dout(w_dff_B_KasjwAkM9_1),.clk(gclk));
	jdff dff_B_6kN2imgs3_0(.din(n1489),.dout(w_dff_B_6kN2imgs3_0),.clk(gclk));
	jdff dff_B_EiultIJq1_0(.din(w_dff_B_6kN2imgs3_0),.dout(w_dff_B_EiultIJq1_0),.clk(gclk));
	jdff dff_B_aE74eXWs0_0(.din(w_dff_B_EiultIJq1_0),.dout(w_dff_B_aE74eXWs0_0),.clk(gclk));
	jdff dff_B_23oOUYVq6_0(.din(w_dff_B_aE74eXWs0_0),.dout(w_dff_B_23oOUYVq6_0),.clk(gclk));
	jdff dff_B_cotjRpX83_0(.din(w_dff_B_23oOUYVq6_0),.dout(w_dff_B_cotjRpX83_0),.clk(gclk));
	jdff dff_A_rMpQbARe6_1(.dout(w_n1486_0[1]),.din(w_dff_A_rMpQbARe6_1),.clk(gclk));
	jdff dff_A_HBMx0F6Y6_1(.dout(w_dff_A_rMpQbARe6_1),.din(w_dff_A_HBMx0F6Y6_1),.clk(gclk));
	jdff dff_A_acFAoB715_1(.dout(w_dff_A_HBMx0F6Y6_1),.din(w_dff_A_acFAoB715_1),.clk(gclk));
	jdff dff_A_gELSl4NY6_1(.dout(w_dff_A_acFAoB715_1),.din(w_dff_A_gELSl4NY6_1),.clk(gclk));
	jdff dff_A_pc60ZrUb1_1(.dout(w_dff_A_gELSl4NY6_1),.din(w_dff_A_pc60ZrUb1_1),.clk(gclk));
	jdff dff_A_njEHyu7l3_1(.dout(w_dff_A_pc60ZrUb1_1),.din(w_dff_A_njEHyu7l3_1),.clk(gclk));
	jdff dff_B_q05ACBSj4_1(.din(n1412),.dout(w_dff_B_q05ACBSj4_1),.clk(gclk));
	jdff dff_B_xZx0QW7B2_1(.din(w_dff_B_q05ACBSj4_1),.dout(w_dff_B_xZx0QW7B2_1),.clk(gclk));
	jdff dff_B_fWrkI66s4_1(.din(w_dff_B_xZx0QW7B2_1),.dout(w_dff_B_fWrkI66s4_1),.clk(gclk));
	jdff dff_B_GlgzqquN0_1(.din(w_dff_B_fWrkI66s4_1),.dout(w_dff_B_GlgzqquN0_1),.clk(gclk));
	jdff dff_B_w0BcUHRx3_1(.din(w_dff_B_GlgzqquN0_1),.dout(w_dff_B_w0BcUHRx3_1),.clk(gclk));
	jdff dff_B_0wQXfKuk2_1(.din(w_dff_B_w0BcUHRx3_1),.dout(w_dff_B_0wQXfKuk2_1),.clk(gclk));
	jdff dff_B_d1g90P6Y5_0(.din(n1413),.dout(w_dff_B_d1g90P6Y5_0),.clk(gclk));
	jdff dff_B_CpLBWBme5_0(.din(w_dff_B_d1g90P6Y5_0),.dout(w_dff_B_CpLBWBme5_0),.clk(gclk));
	jdff dff_B_YpiA6JQf3_0(.din(w_dff_B_CpLBWBme5_0),.dout(w_dff_B_YpiA6JQf3_0),.clk(gclk));
	jdff dff_B_w6qGUp2q7_0(.din(w_dff_B_YpiA6JQf3_0),.dout(w_dff_B_w6qGUp2q7_0),.clk(gclk));
	jdff dff_A_qRWrLJHO5_1(.dout(w_n1410_0[1]),.din(w_dff_A_qRWrLJHO5_1),.clk(gclk));
	jdff dff_A_rLQ3MIbx8_1(.dout(w_dff_A_qRWrLJHO5_1),.din(w_dff_A_rLQ3MIbx8_1),.clk(gclk));
	jdff dff_A_wshycQhA0_1(.dout(w_dff_A_rLQ3MIbx8_1),.din(w_dff_A_wshycQhA0_1),.clk(gclk));
	jdff dff_A_PZSan8Hh2_1(.dout(w_dff_A_wshycQhA0_1),.din(w_dff_A_PZSan8Hh2_1),.clk(gclk));
	jdff dff_A_vT4dEFkO3_1(.dout(w_dff_A_PZSan8Hh2_1),.din(w_dff_A_vT4dEFkO3_1),.clk(gclk));
	jdff dff_B_TneMuxcJ0_1(.din(n1330),.dout(w_dff_B_TneMuxcJ0_1),.clk(gclk));
	jdff dff_B_R5r31NiQ5_1(.din(w_dff_B_TneMuxcJ0_1),.dout(w_dff_B_R5r31NiQ5_1),.clk(gclk));
	jdff dff_B_W6JW4JY46_1(.din(w_dff_B_R5r31NiQ5_1),.dout(w_dff_B_W6JW4JY46_1),.clk(gclk));
	jdff dff_A_hPDweS9h2_0(.dout(w_n1326_0[0]),.din(w_dff_A_hPDweS9h2_0),.clk(gclk));
	jdff dff_A_GY0tRlvX7_0(.dout(w_dff_A_hPDweS9h2_0),.din(w_dff_A_GY0tRlvX7_0),.clk(gclk));
	jdff dff_B_BBetNlil1_1(.din(n1242),.dout(w_dff_B_BBetNlil1_1),.clk(gclk));
	jdff dff_A_3F2qeiCQ3_0(.dout(w_n1238_0[0]),.din(w_dff_A_3F2qeiCQ3_0),.clk(gclk));
	jdff dff_B_OmGa2UCE3_1(.din(n1145),.dout(w_dff_B_OmGa2UCE3_1),.clk(gclk));
	jdff dff_A_hrBreWcA4_1(.dout(w_n1039_0[1]),.din(w_dff_A_hrBreWcA4_1),.clk(gclk));
	jdff dff_B_k77NgaMe2_2(.din(n1037),.dout(w_dff_B_k77NgaMe2_2),.clk(gclk));
	jdff dff_B_2Jd0iHVW5_1(.din(n935),.dout(w_dff_B_2Jd0iHVW5_1),.clk(gclk));
	jdff dff_A_XztLsaWI3_0(.dout(w_n829_0[0]),.din(w_dff_A_XztLsaWI3_0),.clk(gclk));
	jdff dff_A_xnlAbdHd7_0(.dout(w_dff_A_XztLsaWI3_0),.din(w_dff_A_xnlAbdHd7_0),.clk(gclk));
	jdff dff_A_IZBE0o1x6_0(.dout(w_dff_A_xnlAbdHd7_0),.din(w_dff_A_IZBE0o1x6_0),.clk(gclk));
	jdff dff_A_WYzqc2nb3_0(.dout(w_dff_A_IZBE0o1x6_0),.din(w_dff_A_WYzqc2nb3_0),.clk(gclk));
	jdff dff_A_rMekzOQB9_0(.dout(w_dff_A_WYzqc2nb3_0),.din(w_dff_A_rMekzOQB9_0),.clk(gclk));
	jdff dff_A_2uvANXjR1_0(.dout(w_dff_A_rMekzOQB9_0),.din(w_dff_A_2uvANXjR1_0),.clk(gclk));
	jdff dff_A_GKRicQKM4_0(.dout(w_dff_A_2uvANXjR1_0),.din(w_dff_A_GKRicQKM4_0),.clk(gclk));
	jdff dff_A_iK5LrSOU7_0(.dout(w_dff_A_GKRicQKM4_0),.din(w_dff_A_iK5LrSOU7_0),.clk(gclk));
	jdff dff_A_HtoL1htq2_0(.dout(w_dff_A_iK5LrSOU7_0),.din(w_dff_A_HtoL1htq2_0),.clk(gclk));
	jdff dff_A_giro5rPs9_0(.dout(w_dff_A_HtoL1htq2_0),.din(w_dff_A_giro5rPs9_0),.clk(gclk));
	jdff dff_A_TNBabMUo3_0(.dout(w_dff_A_giro5rPs9_0),.din(w_dff_A_TNBabMUo3_0),.clk(gclk));
	jdff dff_A_UQiFp3kU6_0(.dout(w_dff_A_TNBabMUo3_0),.din(w_dff_A_UQiFp3kU6_0),.clk(gclk));
	jdff dff_A_YxTF7zei4_0(.dout(w_dff_A_UQiFp3kU6_0),.din(w_dff_A_YxTF7zei4_0),.clk(gclk));
	jdff dff_A_uQYrV3Kw3_0(.dout(w_dff_A_YxTF7zei4_0),.din(w_dff_A_uQYrV3Kw3_0),.clk(gclk));
	jdff dff_A_dzzTosjp0_0(.dout(w_dff_A_uQYrV3Kw3_0),.din(w_dff_A_dzzTosjp0_0),.clk(gclk));
	jdff dff_A_lJw1AJoj7_0(.dout(w_dff_A_dzzTosjp0_0),.din(w_dff_A_lJw1AJoj7_0),.clk(gclk));
	jdff dff_A_uCWYDUEs9_0(.dout(w_dff_A_lJw1AJoj7_0),.din(w_dff_A_uCWYDUEs9_0),.clk(gclk));
	jdff dff_A_UrefqLHB0_0(.dout(w_dff_A_uCWYDUEs9_0),.din(w_dff_A_UrefqLHB0_0),.clk(gclk));
	jdff dff_A_QqBQw9H95_0(.dout(w_dff_A_UrefqLHB0_0),.din(w_dff_A_QqBQw9H95_0),.clk(gclk));
	jdff dff_A_iUYgljVi1_0(.dout(w_dff_A_QqBQw9H95_0),.din(w_dff_A_iUYgljVi1_0),.clk(gclk));
	jdff dff_A_tQvnKtQ70_0(.dout(w_dff_A_iUYgljVi1_0),.din(w_dff_A_tQvnKtQ70_0),.clk(gclk));
	jdff dff_A_oPVbxvsv2_0(.dout(w_dff_A_tQvnKtQ70_0),.din(w_dff_A_oPVbxvsv2_0),.clk(gclk));
	jdff dff_A_itqnddGD8_0(.dout(w_dff_A_oPVbxvsv2_0),.din(w_dff_A_itqnddGD8_0),.clk(gclk));
	jdff dff_A_3JlSNcIc5_0(.dout(w_dff_A_itqnddGD8_0),.din(w_dff_A_3JlSNcIc5_0),.clk(gclk));
	jdff dff_A_raRNB5ki5_0(.dout(w_dff_A_3JlSNcIc5_0),.din(w_dff_A_raRNB5ki5_0),.clk(gclk));
	jdff dff_A_5WqZGXYg5_0(.dout(w_dff_A_raRNB5ki5_0),.din(w_dff_A_5WqZGXYg5_0),.clk(gclk));
	jdff dff_A_dewhXr0h6_0(.dout(w_dff_A_5WqZGXYg5_0),.din(w_dff_A_dewhXr0h6_0),.clk(gclk));
	jdff dff_A_QSqF0f3R4_0(.dout(w_dff_A_dewhXr0h6_0),.din(w_dff_A_QSqF0f3R4_0),.clk(gclk));
	jdff dff_A_cXIP6Qxb4_0(.dout(w_dff_A_QSqF0f3R4_0),.din(w_dff_A_cXIP6Qxb4_0),.clk(gclk));
	jdff dff_A_veMi3zVL4_0(.dout(w_dff_A_cXIP6Qxb4_0),.din(w_dff_A_veMi3zVL4_0),.clk(gclk));
	jdff dff_A_W5I2SHU40_0(.dout(w_dff_A_veMi3zVL4_0),.din(w_dff_A_W5I2SHU40_0),.clk(gclk));
	jdff dff_A_W8t6BoxU0_0(.dout(w_dff_A_W5I2SHU40_0),.din(w_dff_A_W8t6BoxU0_0),.clk(gclk));
	jdff dff_A_1fyNjCk01_0(.dout(w_dff_A_W8t6BoxU0_0),.din(w_dff_A_1fyNjCk01_0),.clk(gclk));
	jdff dff_A_9PvjUJ8f1_0(.dout(w_dff_A_1fyNjCk01_0),.din(w_dff_A_9PvjUJ8f1_0),.clk(gclk));
	jdff dff_A_qYzi9ijr9_0(.dout(w_dff_A_9PvjUJ8f1_0),.din(w_dff_A_qYzi9ijr9_0),.clk(gclk));
	jdff dff_A_M1TmlG254_0(.dout(w_dff_A_qYzi9ijr9_0),.din(w_dff_A_M1TmlG254_0),.clk(gclk));
	jdff dff_A_5G5kckfl5_0(.dout(w_dff_A_M1TmlG254_0),.din(w_dff_A_5G5kckfl5_0),.clk(gclk));
	jdff dff_A_mPZQ5b8e5_0(.dout(w_dff_A_5G5kckfl5_0),.din(w_dff_A_mPZQ5b8e5_0),.clk(gclk));
	jdff dff_A_MqVzcWX48_0(.dout(w_dff_A_mPZQ5b8e5_0),.din(w_dff_A_MqVzcWX48_0),.clk(gclk));
	jdff dff_A_Iu5dIaPF2_0(.dout(w_dff_A_MqVzcWX48_0),.din(w_dff_A_Iu5dIaPF2_0),.clk(gclk));
	jdff dff_A_bqv7GY0M5_0(.dout(w_dff_A_Iu5dIaPF2_0),.din(w_dff_A_bqv7GY0M5_0),.clk(gclk));
	jdff dff_A_S72Wv5Nx9_0(.dout(w_dff_A_bqv7GY0M5_0),.din(w_dff_A_S72Wv5Nx9_0),.clk(gclk));
	jdff dff_A_z6gwAQrs2_0(.dout(w_dff_A_S72Wv5Nx9_0),.din(w_dff_A_z6gwAQrs2_0),.clk(gclk));
	jdff dff_A_UeowzV526_0(.dout(w_dff_A_z6gwAQrs2_0),.din(w_dff_A_UeowzV526_0),.clk(gclk));
	jdff dff_A_hQoEVyXq2_1(.dout(w_n931_0[1]),.din(w_dff_A_hQoEVyXq2_1),.clk(gclk));
	jdff dff_B_WgXmBxuA8_1(.din(n832),.dout(w_dff_B_WgXmBxuA8_1),.clk(gclk));
	jdff dff_A_PiiIzt3R8_0(.dout(w_n729_0[0]),.din(w_dff_A_PiiIzt3R8_0),.clk(gclk));
	jdff dff_A_I6e6MBN94_0(.dout(w_dff_A_PiiIzt3R8_0),.din(w_dff_A_I6e6MBN94_0),.clk(gclk));
	jdff dff_A_DI0hUnOy4_0(.dout(w_dff_A_I6e6MBN94_0),.din(w_dff_A_DI0hUnOy4_0),.clk(gclk));
	jdff dff_A_j2gyYtOg8_0(.dout(w_dff_A_DI0hUnOy4_0),.din(w_dff_A_j2gyYtOg8_0),.clk(gclk));
	jdff dff_A_FUuFRAB05_0(.dout(w_dff_A_j2gyYtOg8_0),.din(w_dff_A_FUuFRAB05_0),.clk(gclk));
	jdff dff_A_PC4p1H1m1_0(.dout(w_dff_A_FUuFRAB05_0),.din(w_dff_A_PC4p1H1m1_0),.clk(gclk));
	jdff dff_A_ff5HL2R95_0(.dout(w_dff_A_PC4p1H1m1_0),.din(w_dff_A_ff5HL2R95_0),.clk(gclk));
	jdff dff_A_Ed77mGnc4_0(.dout(w_dff_A_ff5HL2R95_0),.din(w_dff_A_Ed77mGnc4_0),.clk(gclk));
	jdff dff_A_BJEJ6zXE4_0(.dout(w_dff_A_Ed77mGnc4_0),.din(w_dff_A_BJEJ6zXE4_0),.clk(gclk));
	jdff dff_A_Rw5MsoPp1_0(.dout(w_dff_A_BJEJ6zXE4_0),.din(w_dff_A_Rw5MsoPp1_0),.clk(gclk));
	jdff dff_A_vt7VItj09_0(.dout(w_dff_A_Rw5MsoPp1_0),.din(w_dff_A_vt7VItj09_0),.clk(gclk));
	jdff dff_A_2ikhUUUE6_0(.dout(w_dff_A_vt7VItj09_0),.din(w_dff_A_2ikhUUUE6_0),.clk(gclk));
	jdff dff_A_9vdDxUv13_0(.dout(w_dff_A_2ikhUUUE6_0),.din(w_dff_A_9vdDxUv13_0),.clk(gclk));
	jdff dff_A_B3Q9oF6k0_0(.dout(w_dff_A_9vdDxUv13_0),.din(w_dff_A_B3Q9oF6k0_0),.clk(gclk));
	jdff dff_A_bKwww85G7_0(.dout(w_dff_A_B3Q9oF6k0_0),.din(w_dff_A_bKwww85G7_0),.clk(gclk));
	jdff dff_A_2b9e82EN5_0(.dout(w_dff_A_bKwww85G7_0),.din(w_dff_A_2b9e82EN5_0),.clk(gclk));
	jdff dff_A_P19Sqdo77_0(.dout(w_dff_A_2b9e82EN5_0),.din(w_dff_A_P19Sqdo77_0),.clk(gclk));
	jdff dff_A_SZzxIYQ15_0(.dout(w_dff_A_P19Sqdo77_0),.din(w_dff_A_SZzxIYQ15_0),.clk(gclk));
	jdff dff_A_cB4yQMR73_0(.dout(w_dff_A_SZzxIYQ15_0),.din(w_dff_A_cB4yQMR73_0),.clk(gclk));
	jdff dff_A_c0vytwfD9_0(.dout(w_dff_A_cB4yQMR73_0),.din(w_dff_A_c0vytwfD9_0),.clk(gclk));
	jdff dff_A_c8KSx1ND0_0(.dout(w_dff_A_c0vytwfD9_0),.din(w_dff_A_c8KSx1ND0_0),.clk(gclk));
	jdff dff_A_JiHQIVAM4_0(.dout(w_dff_A_c8KSx1ND0_0),.din(w_dff_A_JiHQIVAM4_0),.clk(gclk));
	jdff dff_A_kYty4V296_0(.dout(w_dff_A_JiHQIVAM4_0),.din(w_dff_A_kYty4V296_0),.clk(gclk));
	jdff dff_A_RojqhZIA9_0(.dout(w_dff_A_kYty4V296_0),.din(w_dff_A_RojqhZIA9_0),.clk(gclk));
	jdff dff_A_wP5F6fzZ2_0(.dout(w_dff_A_RojqhZIA9_0),.din(w_dff_A_wP5F6fzZ2_0),.clk(gclk));
	jdff dff_A_QZY8CUOS1_0(.dout(w_dff_A_wP5F6fzZ2_0),.din(w_dff_A_QZY8CUOS1_0),.clk(gclk));
	jdff dff_A_jGHnAh5L7_0(.dout(w_dff_A_QZY8CUOS1_0),.din(w_dff_A_jGHnAh5L7_0),.clk(gclk));
	jdff dff_A_nXyRtF1i2_0(.dout(w_dff_A_jGHnAh5L7_0),.din(w_dff_A_nXyRtF1i2_0),.clk(gclk));
	jdff dff_A_XwPGBhfq3_0(.dout(w_dff_A_nXyRtF1i2_0),.din(w_dff_A_XwPGBhfq3_0),.clk(gclk));
	jdff dff_A_222ylpW08_0(.dout(w_dff_A_XwPGBhfq3_0),.din(w_dff_A_222ylpW08_0),.clk(gclk));
	jdff dff_A_NuBlYdaU7_0(.dout(w_dff_A_222ylpW08_0),.din(w_dff_A_NuBlYdaU7_0),.clk(gclk));
	jdff dff_A_iqjfqWP06_0(.dout(w_dff_A_NuBlYdaU7_0),.din(w_dff_A_iqjfqWP06_0),.clk(gclk));
	jdff dff_A_6NZ3krYe9_0(.dout(w_dff_A_iqjfqWP06_0),.din(w_dff_A_6NZ3krYe9_0),.clk(gclk));
	jdff dff_A_3pOUc97J3_0(.dout(w_dff_A_6NZ3krYe9_0),.din(w_dff_A_3pOUc97J3_0),.clk(gclk));
	jdff dff_A_dp2Y069B6_0(.dout(w_dff_A_3pOUc97J3_0),.din(w_dff_A_dp2Y069B6_0),.clk(gclk));
	jdff dff_A_t8XThZsf8_0(.dout(w_dff_A_dp2Y069B6_0),.din(w_dff_A_t8XThZsf8_0),.clk(gclk));
	jdff dff_A_oz8NCmJL2_0(.dout(w_dff_A_t8XThZsf8_0),.din(w_dff_A_oz8NCmJL2_0),.clk(gclk));
	jdff dff_A_9CdNR69I7_0(.dout(w_dff_A_oz8NCmJL2_0),.din(w_dff_A_9CdNR69I7_0),.clk(gclk));
	jdff dff_A_L1XzuGHU3_0(.dout(w_dff_A_9CdNR69I7_0),.din(w_dff_A_L1XzuGHU3_0),.clk(gclk));
	jdff dff_A_WhIZKAjF7_0(.dout(w_dff_A_L1XzuGHU3_0),.din(w_dff_A_WhIZKAjF7_0),.clk(gclk));
	jdff dff_A_v4PrTfen7_0(.dout(w_dff_A_WhIZKAjF7_0),.din(w_dff_A_v4PrTfen7_0),.clk(gclk));
	jdff dff_A_ls7XPJqC5_1(.dout(w_n826_0[1]),.din(w_dff_A_ls7XPJqC5_1),.clk(gclk));
	jdff dff_B_8VzzC10B8_1(.din(n736),.dout(w_dff_B_8VzzC10B8_1),.clk(gclk));
	jdff dff_B_lW2Bhz3d1_1(.din(w_dff_B_8VzzC10B8_1),.dout(w_dff_B_lW2Bhz3d1_1),.clk(gclk));
	jdff dff_B_GszznvkK5_1(.din(w_dff_B_lW2Bhz3d1_1),.dout(w_dff_B_GszznvkK5_1),.clk(gclk));
	jdff dff_B_dIqA0EZB7_1(.din(w_dff_B_GszznvkK5_1),.dout(w_dff_B_dIqA0EZB7_1),.clk(gclk));
	jdff dff_B_IjjNUSPc6_1(.din(w_dff_B_dIqA0EZB7_1),.dout(w_dff_B_IjjNUSPc6_1),.clk(gclk));
	jdff dff_B_kNGsYjop5_1(.din(w_dff_B_IjjNUSPc6_1),.dout(w_dff_B_kNGsYjop5_1),.clk(gclk));
	jdff dff_B_B1YHmoVt1_1(.din(w_dff_B_kNGsYjop5_1),.dout(w_dff_B_B1YHmoVt1_1),.clk(gclk));
	jdff dff_B_Bblgcefy8_1(.din(w_dff_B_B1YHmoVt1_1),.dout(w_dff_B_Bblgcefy8_1),.clk(gclk));
	jdff dff_B_5op6F0yd7_1(.din(w_dff_B_Bblgcefy8_1),.dout(w_dff_B_5op6F0yd7_1),.clk(gclk));
	jdff dff_B_m0G09LZF4_1(.din(w_dff_B_5op6F0yd7_1),.dout(w_dff_B_m0G09LZF4_1),.clk(gclk));
	jdff dff_B_Qi8aYOEC6_1(.din(w_dff_B_m0G09LZF4_1),.dout(w_dff_B_Qi8aYOEC6_1),.clk(gclk));
	jdff dff_B_kCqh92Sm3_1(.din(w_dff_B_Qi8aYOEC6_1),.dout(w_dff_B_kCqh92Sm3_1),.clk(gclk));
	jdff dff_B_qPkrqY9x8_1(.din(w_dff_B_kCqh92Sm3_1),.dout(w_dff_B_qPkrqY9x8_1),.clk(gclk));
	jdff dff_B_Df7brTSZ1_1(.din(w_dff_B_qPkrqY9x8_1),.dout(w_dff_B_Df7brTSZ1_1),.clk(gclk));
	jdff dff_B_dsPxwSMv0_1(.din(w_dff_B_Df7brTSZ1_1),.dout(w_dff_B_dsPxwSMv0_1),.clk(gclk));
	jdff dff_B_1aRYIuQ52_1(.din(w_dff_B_dsPxwSMv0_1),.dout(w_dff_B_1aRYIuQ52_1),.clk(gclk));
	jdff dff_B_A610nrWP2_1(.din(w_dff_B_1aRYIuQ52_1),.dout(w_dff_B_A610nrWP2_1),.clk(gclk));
	jdff dff_B_gGKQdiBh5_1(.din(w_dff_B_A610nrWP2_1),.dout(w_dff_B_gGKQdiBh5_1),.clk(gclk));
	jdff dff_B_qEuix4A42_1(.din(w_dff_B_gGKQdiBh5_1),.dout(w_dff_B_qEuix4A42_1),.clk(gclk));
	jdff dff_B_d1zF20rF8_1(.din(w_dff_B_qEuix4A42_1),.dout(w_dff_B_d1zF20rF8_1),.clk(gclk));
	jdff dff_B_gf3e94Nk0_1(.din(w_dff_B_d1zF20rF8_1),.dout(w_dff_B_gf3e94Nk0_1),.clk(gclk));
	jdff dff_B_e084yyqQ9_1(.din(w_dff_B_gf3e94Nk0_1),.dout(w_dff_B_e084yyqQ9_1),.clk(gclk));
	jdff dff_B_pKqFTqWp9_1(.din(w_dff_B_e084yyqQ9_1),.dout(w_dff_B_pKqFTqWp9_1),.clk(gclk));
	jdff dff_B_9pu5oilm6_1(.din(w_dff_B_pKqFTqWp9_1),.dout(w_dff_B_9pu5oilm6_1),.clk(gclk));
	jdff dff_B_7q7EsWDB4_1(.din(w_dff_B_9pu5oilm6_1),.dout(w_dff_B_7q7EsWDB4_1),.clk(gclk));
	jdff dff_B_idov8ouX8_1(.din(w_dff_B_7q7EsWDB4_1),.dout(w_dff_B_idov8ouX8_1),.clk(gclk));
	jdff dff_B_anLHWe976_1(.din(w_dff_B_idov8ouX8_1),.dout(w_dff_B_anLHWe976_1),.clk(gclk));
	jdff dff_B_XJxIqut58_1(.din(w_dff_B_anLHWe976_1),.dout(w_dff_B_XJxIqut58_1),.clk(gclk));
	jdff dff_B_0oEBqDHD6_1(.din(w_dff_B_XJxIqut58_1),.dout(w_dff_B_0oEBqDHD6_1),.clk(gclk));
	jdff dff_B_5uNkM3F92_1(.din(w_dff_B_0oEBqDHD6_1),.dout(w_dff_B_5uNkM3F92_1),.clk(gclk));
	jdff dff_B_Y3RneUl01_1(.din(w_dff_B_5uNkM3F92_1),.dout(w_dff_B_Y3RneUl01_1),.clk(gclk));
	jdff dff_B_z0sf1KzW4_1(.din(w_dff_B_Y3RneUl01_1),.dout(w_dff_B_z0sf1KzW4_1),.clk(gclk));
	jdff dff_B_uHKisNI68_1(.din(w_dff_B_z0sf1KzW4_1),.dout(w_dff_B_uHKisNI68_1),.clk(gclk));
	jdff dff_B_YMFs8YlH7_1(.din(w_dff_B_uHKisNI68_1),.dout(w_dff_B_YMFs8YlH7_1),.clk(gclk));
	jdff dff_B_hkwLdqAe5_1(.din(w_dff_B_YMFs8YlH7_1),.dout(w_dff_B_hkwLdqAe5_1),.clk(gclk));
	jdff dff_B_sig7arG82_1(.din(w_dff_B_hkwLdqAe5_1),.dout(w_dff_B_sig7arG82_1),.clk(gclk));
	jdff dff_B_xjv428pr0_1(.din(w_dff_B_sig7arG82_1),.dout(w_dff_B_xjv428pr0_1),.clk(gclk));
	jdff dff_B_DpzuuPns0_1(.din(n732),.dout(w_dff_B_DpzuuPns0_1),.clk(gclk));
	jdff dff_A_nA9jw31B6_0(.dout(w_n636_0[0]),.din(w_dff_A_nA9jw31B6_0),.clk(gclk));
	jdff dff_A_23tyB7qe4_0(.dout(w_dff_A_nA9jw31B6_0),.din(w_dff_A_23tyB7qe4_0),.clk(gclk));
	jdff dff_A_XwaEOSLh7_0(.dout(w_dff_A_23tyB7qe4_0),.din(w_dff_A_XwaEOSLh7_0),.clk(gclk));
	jdff dff_A_vE5fslys9_0(.dout(w_dff_A_XwaEOSLh7_0),.din(w_dff_A_vE5fslys9_0),.clk(gclk));
	jdff dff_A_6YvIlmwi6_0(.dout(w_dff_A_vE5fslys9_0),.din(w_dff_A_6YvIlmwi6_0),.clk(gclk));
	jdff dff_A_YYyqgfnK7_0(.dout(w_dff_A_6YvIlmwi6_0),.din(w_dff_A_YYyqgfnK7_0),.clk(gclk));
	jdff dff_A_2EN1hU2K0_0(.dout(w_dff_A_YYyqgfnK7_0),.din(w_dff_A_2EN1hU2K0_0),.clk(gclk));
	jdff dff_A_hzwtpl9Z3_0(.dout(w_dff_A_2EN1hU2K0_0),.din(w_dff_A_hzwtpl9Z3_0),.clk(gclk));
	jdff dff_A_90gH4jFa1_0(.dout(w_dff_A_hzwtpl9Z3_0),.din(w_dff_A_90gH4jFa1_0),.clk(gclk));
	jdff dff_A_FgzVbrpY4_0(.dout(w_dff_A_90gH4jFa1_0),.din(w_dff_A_FgzVbrpY4_0),.clk(gclk));
	jdff dff_A_1XcERHTm8_0(.dout(w_dff_A_FgzVbrpY4_0),.din(w_dff_A_1XcERHTm8_0),.clk(gclk));
	jdff dff_A_wBvetjQi4_0(.dout(w_dff_A_1XcERHTm8_0),.din(w_dff_A_wBvetjQi4_0),.clk(gclk));
	jdff dff_A_ZgbRKsPe0_0(.dout(w_dff_A_wBvetjQi4_0),.din(w_dff_A_ZgbRKsPe0_0),.clk(gclk));
	jdff dff_A_fjrB3MRu2_0(.dout(w_dff_A_ZgbRKsPe0_0),.din(w_dff_A_fjrB3MRu2_0),.clk(gclk));
	jdff dff_A_4viJ7sGW2_0(.dout(w_dff_A_fjrB3MRu2_0),.din(w_dff_A_4viJ7sGW2_0),.clk(gclk));
	jdff dff_A_ZWMKS3Hy3_0(.dout(w_dff_A_4viJ7sGW2_0),.din(w_dff_A_ZWMKS3Hy3_0),.clk(gclk));
	jdff dff_A_mjQvio0T8_0(.dout(w_dff_A_ZWMKS3Hy3_0),.din(w_dff_A_mjQvio0T8_0),.clk(gclk));
	jdff dff_A_kLFRzyFN5_0(.dout(w_dff_A_mjQvio0T8_0),.din(w_dff_A_kLFRzyFN5_0),.clk(gclk));
	jdff dff_A_mWy1c4T31_0(.dout(w_dff_A_kLFRzyFN5_0),.din(w_dff_A_mWy1c4T31_0),.clk(gclk));
	jdff dff_A_HCg9oAAy7_0(.dout(w_dff_A_mWy1c4T31_0),.din(w_dff_A_HCg9oAAy7_0),.clk(gclk));
	jdff dff_A_djxzIVmo4_0(.dout(w_dff_A_HCg9oAAy7_0),.din(w_dff_A_djxzIVmo4_0),.clk(gclk));
	jdff dff_A_R5abQt844_0(.dout(w_dff_A_djxzIVmo4_0),.din(w_dff_A_R5abQt844_0),.clk(gclk));
	jdff dff_A_CmWCl49J9_0(.dout(w_dff_A_R5abQt844_0),.din(w_dff_A_CmWCl49J9_0),.clk(gclk));
	jdff dff_A_z0bjo0uP4_0(.dout(w_dff_A_CmWCl49J9_0),.din(w_dff_A_z0bjo0uP4_0),.clk(gclk));
	jdff dff_A_JXVj8edD7_0(.dout(w_dff_A_z0bjo0uP4_0),.din(w_dff_A_JXVj8edD7_0),.clk(gclk));
	jdff dff_A_fyaOQ5gL1_0(.dout(w_dff_A_JXVj8edD7_0),.din(w_dff_A_fyaOQ5gL1_0),.clk(gclk));
	jdff dff_A_i7Zvo5oI9_0(.dout(w_dff_A_fyaOQ5gL1_0),.din(w_dff_A_i7Zvo5oI9_0),.clk(gclk));
	jdff dff_A_1t8sO5HL6_0(.dout(w_dff_A_i7Zvo5oI9_0),.din(w_dff_A_1t8sO5HL6_0),.clk(gclk));
	jdff dff_A_q8C2996N9_0(.dout(w_dff_A_1t8sO5HL6_0),.din(w_dff_A_q8C2996N9_0),.clk(gclk));
	jdff dff_A_WzsIyWS02_0(.dout(w_dff_A_q8C2996N9_0),.din(w_dff_A_WzsIyWS02_0),.clk(gclk));
	jdff dff_A_UKKkdDDR4_0(.dout(w_dff_A_WzsIyWS02_0),.din(w_dff_A_UKKkdDDR4_0),.clk(gclk));
	jdff dff_A_LVFMzPm42_0(.dout(w_dff_A_UKKkdDDR4_0),.din(w_dff_A_LVFMzPm42_0),.clk(gclk));
	jdff dff_A_5IrwuyqO3_0(.dout(w_dff_A_LVFMzPm42_0),.din(w_dff_A_5IrwuyqO3_0),.clk(gclk));
	jdff dff_A_LXmC66Bo0_0(.dout(w_dff_A_5IrwuyqO3_0),.din(w_dff_A_LXmC66Bo0_0),.clk(gclk));
	jdff dff_A_WusR1u5e7_0(.dout(w_dff_A_LXmC66Bo0_0),.din(w_dff_A_WusR1u5e7_0),.clk(gclk));
	jdff dff_A_gSX6UWhN7_0(.dout(w_dff_A_WusR1u5e7_0),.din(w_dff_A_gSX6UWhN7_0),.clk(gclk));
	jdff dff_A_Jb2z1ag75_0(.dout(w_dff_A_gSX6UWhN7_0),.din(w_dff_A_Jb2z1ag75_0),.clk(gclk));
	jdff dff_A_evevrTmx4_0(.dout(w_dff_A_Jb2z1ag75_0),.din(w_dff_A_evevrTmx4_0),.clk(gclk));
	jdff dff_A_90iIDhbQ1_1(.dout(w_n726_0[1]),.din(w_dff_A_90iIDhbQ1_1),.clk(gclk));
	jdff dff_B_8GwMWOwi5_1(.din(n643),.dout(w_dff_B_8GwMWOwi5_1),.clk(gclk));
	jdff dff_B_wjSGixRt4_1(.din(w_dff_B_8GwMWOwi5_1),.dout(w_dff_B_wjSGixRt4_1),.clk(gclk));
	jdff dff_B_PfTadJ1a7_1(.din(w_dff_B_wjSGixRt4_1),.dout(w_dff_B_PfTadJ1a7_1),.clk(gclk));
	jdff dff_B_xbIpS5bo9_1(.din(w_dff_B_PfTadJ1a7_1),.dout(w_dff_B_xbIpS5bo9_1),.clk(gclk));
	jdff dff_B_rjAWUfle1_1(.din(w_dff_B_xbIpS5bo9_1),.dout(w_dff_B_rjAWUfle1_1),.clk(gclk));
	jdff dff_B_3hSQSrmw5_1(.din(w_dff_B_rjAWUfle1_1),.dout(w_dff_B_3hSQSrmw5_1),.clk(gclk));
	jdff dff_B_IGCzFkC48_1(.din(w_dff_B_3hSQSrmw5_1),.dout(w_dff_B_IGCzFkC48_1),.clk(gclk));
	jdff dff_B_TTqoxdy02_1(.din(w_dff_B_IGCzFkC48_1),.dout(w_dff_B_TTqoxdy02_1),.clk(gclk));
	jdff dff_B_EbOVk6836_1(.din(w_dff_B_TTqoxdy02_1),.dout(w_dff_B_EbOVk6836_1),.clk(gclk));
	jdff dff_B_Nd3oec7e5_1(.din(w_dff_B_EbOVk6836_1),.dout(w_dff_B_Nd3oec7e5_1),.clk(gclk));
	jdff dff_B_aK7nwTNr0_1(.din(w_dff_B_Nd3oec7e5_1),.dout(w_dff_B_aK7nwTNr0_1),.clk(gclk));
	jdff dff_B_mBYciLTO1_1(.din(w_dff_B_aK7nwTNr0_1),.dout(w_dff_B_mBYciLTO1_1),.clk(gclk));
	jdff dff_B_LZfPGB4O3_1(.din(w_dff_B_mBYciLTO1_1),.dout(w_dff_B_LZfPGB4O3_1),.clk(gclk));
	jdff dff_B_PkFReVkE7_1(.din(w_dff_B_LZfPGB4O3_1),.dout(w_dff_B_PkFReVkE7_1),.clk(gclk));
	jdff dff_B_8E8txXkl3_1(.din(w_dff_B_PkFReVkE7_1),.dout(w_dff_B_8E8txXkl3_1),.clk(gclk));
	jdff dff_B_rk4MerAO0_1(.din(w_dff_B_8E8txXkl3_1),.dout(w_dff_B_rk4MerAO0_1),.clk(gclk));
	jdff dff_B_1B0G0wJu3_1(.din(w_dff_B_rk4MerAO0_1),.dout(w_dff_B_1B0G0wJu3_1),.clk(gclk));
	jdff dff_B_Ypa3paFi0_1(.din(w_dff_B_1B0G0wJu3_1),.dout(w_dff_B_Ypa3paFi0_1),.clk(gclk));
	jdff dff_B_BepEl4gS3_1(.din(w_dff_B_Ypa3paFi0_1),.dout(w_dff_B_BepEl4gS3_1),.clk(gclk));
	jdff dff_B_zw0CxJy35_1(.din(w_dff_B_BepEl4gS3_1),.dout(w_dff_B_zw0CxJy35_1),.clk(gclk));
	jdff dff_B_XCArx3YC5_1(.din(w_dff_B_zw0CxJy35_1),.dout(w_dff_B_XCArx3YC5_1),.clk(gclk));
	jdff dff_B_Tfpplh7L3_1(.din(w_dff_B_XCArx3YC5_1),.dout(w_dff_B_Tfpplh7L3_1),.clk(gclk));
	jdff dff_B_npfMN3jQ8_1(.din(w_dff_B_Tfpplh7L3_1),.dout(w_dff_B_npfMN3jQ8_1),.clk(gclk));
	jdff dff_B_zcm2AJ8X1_1(.din(w_dff_B_npfMN3jQ8_1),.dout(w_dff_B_zcm2AJ8X1_1),.clk(gclk));
	jdff dff_B_TJysLcki0_1(.din(w_dff_B_zcm2AJ8X1_1),.dout(w_dff_B_TJysLcki0_1),.clk(gclk));
	jdff dff_B_ATal7wO17_1(.din(w_dff_B_TJysLcki0_1),.dout(w_dff_B_ATal7wO17_1),.clk(gclk));
	jdff dff_B_V5qXykAA4_1(.din(w_dff_B_ATal7wO17_1),.dout(w_dff_B_V5qXykAA4_1),.clk(gclk));
	jdff dff_B_AwxioecJ7_1(.din(w_dff_B_V5qXykAA4_1),.dout(w_dff_B_AwxioecJ7_1),.clk(gclk));
	jdff dff_B_m0V5luZO3_1(.din(w_dff_B_AwxioecJ7_1),.dout(w_dff_B_m0V5luZO3_1),.clk(gclk));
	jdff dff_B_G3AF7vZ51_1(.din(w_dff_B_m0V5luZO3_1),.dout(w_dff_B_G3AF7vZ51_1),.clk(gclk));
	jdff dff_B_FhKe6taQ1_1(.din(w_dff_B_G3AF7vZ51_1),.dout(w_dff_B_FhKe6taQ1_1),.clk(gclk));
	jdff dff_B_FxSvqxgM2_1(.din(w_dff_B_FhKe6taQ1_1),.dout(w_dff_B_FxSvqxgM2_1),.clk(gclk));
	jdff dff_B_0FnM0RF66_1(.din(w_dff_B_FxSvqxgM2_1),.dout(w_dff_B_0FnM0RF66_1),.clk(gclk));
	jdff dff_B_ecnqGgPb9_1(.din(w_dff_B_0FnM0RF66_1),.dout(w_dff_B_ecnqGgPb9_1),.clk(gclk));
	jdff dff_B_y1OoywVh9_1(.din(n639),.dout(w_dff_B_y1OoywVh9_1),.clk(gclk));
	jdff dff_A_wjHhreBH5_0(.dout(w_n550_0[0]),.din(w_dff_A_wjHhreBH5_0),.clk(gclk));
	jdff dff_A_kHIIfzcz3_0(.dout(w_dff_A_wjHhreBH5_0),.din(w_dff_A_kHIIfzcz3_0),.clk(gclk));
	jdff dff_A_pNw3Vfkk7_0(.dout(w_dff_A_kHIIfzcz3_0),.din(w_dff_A_pNw3Vfkk7_0),.clk(gclk));
	jdff dff_A_CuI1nMiy9_0(.dout(w_dff_A_pNw3Vfkk7_0),.din(w_dff_A_CuI1nMiy9_0),.clk(gclk));
	jdff dff_A_WjdbFQ856_0(.dout(w_dff_A_CuI1nMiy9_0),.din(w_dff_A_WjdbFQ856_0),.clk(gclk));
	jdff dff_A_8FPxcX2V4_0(.dout(w_dff_A_WjdbFQ856_0),.din(w_dff_A_8FPxcX2V4_0),.clk(gclk));
	jdff dff_A_6V0mvtf37_0(.dout(w_dff_A_8FPxcX2V4_0),.din(w_dff_A_6V0mvtf37_0),.clk(gclk));
	jdff dff_A_eCAGxrrg2_0(.dout(w_dff_A_6V0mvtf37_0),.din(w_dff_A_eCAGxrrg2_0),.clk(gclk));
	jdff dff_A_ltU7wmsA2_0(.dout(w_dff_A_eCAGxrrg2_0),.din(w_dff_A_ltU7wmsA2_0),.clk(gclk));
	jdff dff_A_2xJ5iN1W9_0(.dout(w_dff_A_ltU7wmsA2_0),.din(w_dff_A_2xJ5iN1W9_0),.clk(gclk));
	jdff dff_A_sSc3NPIN9_0(.dout(w_dff_A_2xJ5iN1W9_0),.din(w_dff_A_sSc3NPIN9_0),.clk(gclk));
	jdff dff_A_vbGXJaMS9_0(.dout(w_dff_A_sSc3NPIN9_0),.din(w_dff_A_vbGXJaMS9_0),.clk(gclk));
	jdff dff_A_CMML3V2z0_0(.dout(w_dff_A_vbGXJaMS9_0),.din(w_dff_A_CMML3V2z0_0),.clk(gclk));
	jdff dff_A_ka4veQaB0_0(.dout(w_dff_A_CMML3V2z0_0),.din(w_dff_A_ka4veQaB0_0),.clk(gclk));
	jdff dff_A_uBByO3HM8_0(.dout(w_dff_A_ka4veQaB0_0),.din(w_dff_A_uBByO3HM8_0),.clk(gclk));
	jdff dff_A_pWQUe7gN1_0(.dout(w_dff_A_uBByO3HM8_0),.din(w_dff_A_pWQUe7gN1_0),.clk(gclk));
	jdff dff_A_rw4GaEQf6_0(.dout(w_dff_A_pWQUe7gN1_0),.din(w_dff_A_rw4GaEQf6_0),.clk(gclk));
	jdff dff_A_asnyFLVr1_0(.dout(w_dff_A_rw4GaEQf6_0),.din(w_dff_A_asnyFLVr1_0),.clk(gclk));
	jdff dff_A_Iwagun5z0_0(.dout(w_dff_A_asnyFLVr1_0),.din(w_dff_A_Iwagun5z0_0),.clk(gclk));
	jdff dff_A_QjD8yeB65_0(.dout(w_dff_A_Iwagun5z0_0),.din(w_dff_A_QjD8yeB65_0),.clk(gclk));
	jdff dff_A_i8nJWRvf8_0(.dout(w_dff_A_QjD8yeB65_0),.din(w_dff_A_i8nJWRvf8_0),.clk(gclk));
	jdff dff_A_XOYjXaGu2_0(.dout(w_dff_A_i8nJWRvf8_0),.din(w_dff_A_XOYjXaGu2_0),.clk(gclk));
	jdff dff_A_Efev6IZb6_0(.dout(w_dff_A_XOYjXaGu2_0),.din(w_dff_A_Efev6IZb6_0),.clk(gclk));
	jdff dff_A_oRSD7Bg98_0(.dout(w_dff_A_Efev6IZb6_0),.din(w_dff_A_oRSD7Bg98_0),.clk(gclk));
	jdff dff_A_4Ew5CFO26_0(.dout(w_dff_A_oRSD7Bg98_0),.din(w_dff_A_4Ew5CFO26_0),.clk(gclk));
	jdff dff_A_s9G4wvIg4_0(.dout(w_dff_A_4Ew5CFO26_0),.din(w_dff_A_s9G4wvIg4_0),.clk(gclk));
	jdff dff_A_rfCgWFzs2_0(.dout(w_dff_A_s9G4wvIg4_0),.din(w_dff_A_rfCgWFzs2_0),.clk(gclk));
	jdff dff_A_GCa1fvs20_0(.dout(w_dff_A_rfCgWFzs2_0),.din(w_dff_A_GCa1fvs20_0),.clk(gclk));
	jdff dff_A_6ZEIhEwW2_0(.dout(w_dff_A_GCa1fvs20_0),.din(w_dff_A_6ZEIhEwW2_0),.clk(gclk));
	jdff dff_A_H1nUe7rP0_0(.dout(w_dff_A_6ZEIhEwW2_0),.din(w_dff_A_H1nUe7rP0_0),.clk(gclk));
	jdff dff_A_jSl38lnw2_0(.dout(w_dff_A_H1nUe7rP0_0),.din(w_dff_A_jSl38lnw2_0),.clk(gclk));
	jdff dff_A_SP3GChog1_0(.dout(w_dff_A_jSl38lnw2_0),.din(w_dff_A_SP3GChog1_0),.clk(gclk));
	jdff dff_A_S0GLViYs8_0(.dout(w_dff_A_SP3GChog1_0),.din(w_dff_A_S0GLViYs8_0),.clk(gclk));
	jdff dff_A_hrtsktC32_0(.dout(w_dff_A_S0GLViYs8_0),.din(w_dff_A_hrtsktC32_0),.clk(gclk));
	jdff dff_A_aYONlrSn6_0(.dout(w_dff_A_hrtsktC32_0),.din(w_dff_A_aYONlrSn6_0),.clk(gclk));
	jdff dff_A_XitmDLyL7_1(.dout(w_n633_0[1]),.din(w_dff_A_XitmDLyL7_1),.clk(gclk));
	jdff dff_B_bQKhF1F47_1(.din(n557),.dout(w_dff_B_bQKhF1F47_1),.clk(gclk));
	jdff dff_B_vjuSIyUB2_1(.din(w_dff_B_bQKhF1F47_1),.dout(w_dff_B_vjuSIyUB2_1),.clk(gclk));
	jdff dff_B_PcHPSCLQ2_1(.din(w_dff_B_vjuSIyUB2_1),.dout(w_dff_B_PcHPSCLQ2_1),.clk(gclk));
	jdff dff_B_QdtqTTb28_1(.din(w_dff_B_PcHPSCLQ2_1),.dout(w_dff_B_QdtqTTb28_1),.clk(gclk));
	jdff dff_B_qXnzfyTX4_1(.din(w_dff_B_QdtqTTb28_1),.dout(w_dff_B_qXnzfyTX4_1),.clk(gclk));
	jdff dff_B_qIzEorvX0_1(.din(w_dff_B_qXnzfyTX4_1),.dout(w_dff_B_qIzEorvX0_1),.clk(gclk));
	jdff dff_B_nL0F2n6x6_1(.din(w_dff_B_qIzEorvX0_1),.dout(w_dff_B_nL0F2n6x6_1),.clk(gclk));
	jdff dff_B_yvW3kLcj1_1(.din(w_dff_B_nL0F2n6x6_1),.dout(w_dff_B_yvW3kLcj1_1),.clk(gclk));
	jdff dff_B_fFf8iiWK8_1(.din(w_dff_B_yvW3kLcj1_1),.dout(w_dff_B_fFf8iiWK8_1),.clk(gclk));
	jdff dff_B_RLagDZks1_1(.din(w_dff_B_fFf8iiWK8_1),.dout(w_dff_B_RLagDZks1_1),.clk(gclk));
	jdff dff_B_Ut3jzycM5_1(.din(w_dff_B_RLagDZks1_1),.dout(w_dff_B_Ut3jzycM5_1),.clk(gclk));
	jdff dff_B_doUVHaHM0_1(.din(w_dff_B_Ut3jzycM5_1),.dout(w_dff_B_doUVHaHM0_1),.clk(gclk));
	jdff dff_B_p50seZT68_1(.din(w_dff_B_doUVHaHM0_1),.dout(w_dff_B_p50seZT68_1),.clk(gclk));
	jdff dff_B_U9Ml2wZm5_1(.din(w_dff_B_p50seZT68_1),.dout(w_dff_B_U9Ml2wZm5_1),.clk(gclk));
	jdff dff_B_MREcElIB3_1(.din(w_dff_B_U9Ml2wZm5_1),.dout(w_dff_B_MREcElIB3_1),.clk(gclk));
	jdff dff_B_YW9BFBrY3_1(.din(w_dff_B_MREcElIB3_1),.dout(w_dff_B_YW9BFBrY3_1),.clk(gclk));
	jdff dff_B_mHPEN9Xj0_1(.din(w_dff_B_YW9BFBrY3_1),.dout(w_dff_B_mHPEN9Xj0_1),.clk(gclk));
	jdff dff_B_5br7u1YE9_1(.din(w_dff_B_mHPEN9Xj0_1),.dout(w_dff_B_5br7u1YE9_1),.clk(gclk));
	jdff dff_B_rW3gkcug8_1(.din(w_dff_B_5br7u1YE9_1),.dout(w_dff_B_rW3gkcug8_1),.clk(gclk));
	jdff dff_B_VpOX9ND18_1(.din(w_dff_B_rW3gkcug8_1),.dout(w_dff_B_VpOX9ND18_1),.clk(gclk));
	jdff dff_B_RnKFdvZv0_1(.din(w_dff_B_VpOX9ND18_1),.dout(w_dff_B_RnKFdvZv0_1),.clk(gclk));
	jdff dff_B_4BS9jKbC4_1(.din(w_dff_B_RnKFdvZv0_1),.dout(w_dff_B_4BS9jKbC4_1),.clk(gclk));
	jdff dff_B_tOPjf5nt5_1(.din(w_dff_B_4BS9jKbC4_1),.dout(w_dff_B_tOPjf5nt5_1),.clk(gclk));
	jdff dff_B_hblLleH77_1(.din(w_dff_B_tOPjf5nt5_1),.dout(w_dff_B_hblLleH77_1),.clk(gclk));
	jdff dff_B_6OcBKw6m0_1(.din(w_dff_B_hblLleH77_1),.dout(w_dff_B_6OcBKw6m0_1),.clk(gclk));
	jdff dff_B_buaxEEK13_1(.din(w_dff_B_6OcBKw6m0_1),.dout(w_dff_B_buaxEEK13_1),.clk(gclk));
	jdff dff_B_rFvh3htF3_1(.din(w_dff_B_buaxEEK13_1),.dout(w_dff_B_rFvh3htF3_1),.clk(gclk));
	jdff dff_B_9Yvcven91_1(.din(w_dff_B_rFvh3htF3_1),.dout(w_dff_B_9Yvcven91_1),.clk(gclk));
	jdff dff_B_8cNmkGp30_1(.din(w_dff_B_9Yvcven91_1),.dout(w_dff_B_8cNmkGp30_1),.clk(gclk));
	jdff dff_B_M7jHNoC75_1(.din(w_dff_B_8cNmkGp30_1),.dout(w_dff_B_M7jHNoC75_1),.clk(gclk));
	jdff dff_B_Ga7CVoxM6_1(.din(w_dff_B_M7jHNoC75_1),.dout(w_dff_B_Ga7CVoxM6_1),.clk(gclk));
	jdff dff_B_XVNnUZs48_1(.din(n553),.dout(w_dff_B_XVNnUZs48_1),.clk(gclk));
	jdff dff_A_cup175MQ3_0(.dout(w_n471_0[0]),.din(w_dff_A_cup175MQ3_0),.clk(gclk));
	jdff dff_A_VGGhTwsL0_0(.dout(w_dff_A_cup175MQ3_0),.din(w_dff_A_VGGhTwsL0_0),.clk(gclk));
	jdff dff_A_8JxtuMRC3_0(.dout(w_dff_A_VGGhTwsL0_0),.din(w_dff_A_8JxtuMRC3_0),.clk(gclk));
	jdff dff_A_p7tuihX95_0(.dout(w_dff_A_8JxtuMRC3_0),.din(w_dff_A_p7tuihX95_0),.clk(gclk));
	jdff dff_A_PbganX0l8_0(.dout(w_dff_A_p7tuihX95_0),.din(w_dff_A_PbganX0l8_0),.clk(gclk));
	jdff dff_A_WDaqGhkC0_0(.dout(w_dff_A_PbganX0l8_0),.din(w_dff_A_WDaqGhkC0_0),.clk(gclk));
	jdff dff_A_f0j3Hkkh9_0(.dout(w_dff_A_WDaqGhkC0_0),.din(w_dff_A_f0j3Hkkh9_0),.clk(gclk));
	jdff dff_A_9hW3Rs4c1_0(.dout(w_dff_A_f0j3Hkkh9_0),.din(w_dff_A_9hW3Rs4c1_0),.clk(gclk));
	jdff dff_A_pAF6pTS79_0(.dout(w_dff_A_9hW3Rs4c1_0),.din(w_dff_A_pAF6pTS79_0),.clk(gclk));
	jdff dff_A_SJTcTBc30_0(.dout(w_dff_A_pAF6pTS79_0),.din(w_dff_A_SJTcTBc30_0),.clk(gclk));
	jdff dff_A_68QkYdto2_0(.dout(w_dff_A_SJTcTBc30_0),.din(w_dff_A_68QkYdto2_0),.clk(gclk));
	jdff dff_A_ILiET0zh3_0(.dout(w_dff_A_68QkYdto2_0),.din(w_dff_A_ILiET0zh3_0),.clk(gclk));
	jdff dff_A_ZO5bSGG75_0(.dout(w_dff_A_ILiET0zh3_0),.din(w_dff_A_ZO5bSGG75_0),.clk(gclk));
	jdff dff_A_3u8TvXnr2_0(.dout(w_dff_A_ZO5bSGG75_0),.din(w_dff_A_3u8TvXnr2_0),.clk(gclk));
	jdff dff_A_H2nB6pCw4_0(.dout(w_dff_A_3u8TvXnr2_0),.din(w_dff_A_H2nB6pCw4_0),.clk(gclk));
	jdff dff_A_RZTEJqO27_0(.dout(w_dff_A_H2nB6pCw4_0),.din(w_dff_A_RZTEJqO27_0),.clk(gclk));
	jdff dff_A_JoNuCgjT2_0(.dout(w_dff_A_RZTEJqO27_0),.din(w_dff_A_JoNuCgjT2_0),.clk(gclk));
	jdff dff_A_qL8ypbtA8_0(.dout(w_dff_A_JoNuCgjT2_0),.din(w_dff_A_qL8ypbtA8_0),.clk(gclk));
	jdff dff_A_2aoblbmy5_0(.dout(w_dff_A_qL8ypbtA8_0),.din(w_dff_A_2aoblbmy5_0),.clk(gclk));
	jdff dff_A_OhyDLvdh6_0(.dout(w_dff_A_2aoblbmy5_0),.din(w_dff_A_OhyDLvdh6_0),.clk(gclk));
	jdff dff_A_iSskpdNs3_0(.dout(w_dff_A_OhyDLvdh6_0),.din(w_dff_A_iSskpdNs3_0),.clk(gclk));
	jdff dff_A_hQfPfrTh2_0(.dout(w_dff_A_iSskpdNs3_0),.din(w_dff_A_hQfPfrTh2_0),.clk(gclk));
	jdff dff_A_u0aQlJdh3_0(.dout(w_dff_A_hQfPfrTh2_0),.din(w_dff_A_u0aQlJdh3_0),.clk(gclk));
	jdff dff_A_DOmuxUPB5_0(.dout(w_dff_A_u0aQlJdh3_0),.din(w_dff_A_DOmuxUPB5_0),.clk(gclk));
	jdff dff_A_GuuIyRFy5_0(.dout(w_dff_A_DOmuxUPB5_0),.din(w_dff_A_GuuIyRFy5_0),.clk(gclk));
	jdff dff_A_1DyrCIQR3_0(.dout(w_dff_A_GuuIyRFy5_0),.din(w_dff_A_1DyrCIQR3_0),.clk(gclk));
	jdff dff_A_Sz2mTKNr3_0(.dout(w_dff_A_1DyrCIQR3_0),.din(w_dff_A_Sz2mTKNr3_0),.clk(gclk));
	jdff dff_A_7RPHRJMB6_0(.dout(w_dff_A_Sz2mTKNr3_0),.din(w_dff_A_7RPHRJMB6_0),.clk(gclk));
	jdff dff_A_Yngj7ojn7_0(.dout(w_dff_A_7RPHRJMB6_0),.din(w_dff_A_Yngj7ojn7_0),.clk(gclk));
	jdff dff_A_VegrjOOJ0_0(.dout(w_dff_A_Yngj7ojn7_0),.din(w_dff_A_VegrjOOJ0_0),.clk(gclk));
	jdff dff_A_GpCWbGKG9_0(.dout(w_dff_A_VegrjOOJ0_0),.din(w_dff_A_GpCWbGKG9_0),.clk(gclk));
	jdff dff_A_YKx6JKpo5_0(.dout(w_dff_A_GpCWbGKG9_0),.din(w_dff_A_YKx6JKpo5_0),.clk(gclk));
	jdff dff_A_J8sheeoS5_1(.dout(w_n547_0[1]),.din(w_dff_A_J8sheeoS5_1),.clk(gclk));
	jdff dff_B_jrF5iNMt4_1(.din(n478),.dout(w_dff_B_jrF5iNMt4_1),.clk(gclk));
	jdff dff_B_hMXa6umq4_1(.din(w_dff_B_jrF5iNMt4_1),.dout(w_dff_B_hMXa6umq4_1),.clk(gclk));
	jdff dff_B_33VFdYq93_1(.din(w_dff_B_hMXa6umq4_1),.dout(w_dff_B_33VFdYq93_1),.clk(gclk));
	jdff dff_B_CqaD6UHH1_1(.din(w_dff_B_33VFdYq93_1),.dout(w_dff_B_CqaD6UHH1_1),.clk(gclk));
	jdff dff_B_UfUEr0xq4_1(.din(w_dff_B_CqaD6UHH1_1),.dout(w_dff_B_UfUEr0xq4_1),.clk(gclk));
	jdff dff_B_pQzfiOQg9_1(.din(w_dff_B_UfUEr0xq4_1),.dout(w_dff_B_pQzfiOQg9_1),.clk(gclk));
	jdff dff_B_D8CY7Prf3_1(.din(w_dff_B_pQzfiOQg9_1),.dout(w_dff_B_D8CY7Prf3_1),.clk(gclk));
	jdff dff_B_iQni8Os93_1(.din(w_dff_B_D8CY7Prf3_1),.dout(w_dff_B_iQni8Os93_1),.clk(gclk));
	jdff dff_B_4JPkIfmu0_1(.din(w_dff_B_iQni8Os93_1),.dout(w_dff_B_4JPkIfmu0_1),.clk(gclk));
	jdff dff_B_gPMIkARU2_1(.din(w_dff_B_4JPkIfmu0_1),.dout(w_dff_B_gPMIkARU2_1),.clk(gclk));
	jdff dff_B_jv1RGV173_1(.din(w_dff_B_gPMIkARU2_1),.dout(w_dff_B_jv1RGV173_1),.clk(gclk));
	jdff dff_B_uskEw4QF4_1(.din(w_dff_B_jv1RGV173_1),.dout(w_dff_B_uskEw4QF4_1),.clk(gclk));
	jdff dff_B_NIyWbGYb4_1(.din(w_dff_B_uskEw4QF4_1),.dout(w_dff_B_NIyWbGYb4_1),.clk(gclk));
	jdff dff_B_mpsZPCTS8_1(.din(w_dff_B_NIyWbGYb4_1),.dout(w_dff_B_mpsZPCTS8_1),.clk(gclk));
	jdff dff_B_66iPT5vT4_1(.din(w_dff_B_mpsZPCTS8_1),.dout(w_dff_B_66iPT5vT4_1),.clk(gclk));
	jdff dff_B_m0XG0Q223_1(.din(w_dff_B_66iPT5vT4_1),.dout(w_dff_B_m0XG0Q223_1),.clk(gclk));
	jdff dff_B_1TFWPF3C5_1(.din(w_dff_B_m0XG0Q223_1),.dout(w_dff_B_1TFWPF3C5_1),.clk(gclk));
	jdff dff_B_a6UUGYvC2_1(.din(w_dff_B_1TFWPF3C5_1),.dout(w_dff_B_a6UUGYvC2_1),.clk(gclk));
	jdff dff_B_zTNQmmtu5_1(.din(w_dff_B_a6UUGYvC2_1),.dout(w_dff_B_zTNQmmtu5_1),.clk(gclk));
	jdff dff_B_TfPXk9OU3_1(.din(w_dff_B_zTNQmmtu5_1),.dout(w_dff_B_TfPXk9OU3_1),.clk(gclk));
	jdff dff_B_wkDuxIzr9_1(.din(w_dff_B_TfPXk9OU3_1),.dout(w_dff_B_wkDuxIzr9_1),.clk(gclk));
	jdff dff_B_ds9l8EH26_1(.din(w_dff_B_wkDuxIzr9_1),.dout(w_dff_B_ds9l8EH26_1),.clk(gclk));
	jdff dff_B_nbv2E0wK9_1(.din(w_dff_B_ds9l8EH26_1),.dout(w_dff_B_nbv2E0wK9_1),.clk(gclk));
	jdff dff_B_7sfGItpL4_1(.din(w_dff_B_nbv2E0wK9_1),.dout(w_dff_B_7sfGItpL4_1),.clk(gclk));
	jdff dff_B_lkAEWT7l6_1(.din(w_dff_B_7sfGItpL4_1),.dout(w_dff_B_lkAEWT7l6_1),.clk(gclk));
	jdff dff_B_9MUXxqf55_1(.din(w_dff_B_lkAEWT7l6_1),.dout(w_dff_B_9MUXxqf55_1),.clk(gclk));
	jdff dff_B_IwBOIOfu2_1(.din(w_dff_B_9MUXxqf55_1),.dout(w_dff_B_IwBOIOfu2_1),.clk(gclk));
	jdff dff_B_i7Y5QUbp9_1(.din(w_dff_B_IwBOIOfu2_1),.dout(w_dff_B_i7Y5QUbp9_1),.clk(gclk));
	jdff dff_B_Sas486Fy7_1(.din(n474),.dout(w_dff_B_Sas486Fy7_1),.clk(gclk));
	jdff dff_A_clNM4O544_0(.dout(w_n399_0[0]),.din(w_dff_A_clNM4O544_0),.clk(gclk));
	jdff dff_A_FRDKW83e5_0(.dout(w_dff_A_clNM4O544_0),.din(w_dff_A_FRDKW83e5_0),.clk(gclk));
	jdff dff_A_2pubCDBU9_0(.dout(w_dff_A_FRDKW83e5_0),.din(w_dff_A_2pubCDBU9_0),.clk(gclk));
	jdff dff_A_u6cC8iEo2_0(.dout(w_dff_A_2pubCDBU9_0),.din(w_dff_A_u6cC8iEo2_0),.clk(gclk));
	jdff dff_A_bihMRFSc1_0(.dout(w_dff_A_u6cC8iEo2_0),.din(w_dff_A_bihMRFSc1_0),.clk(gclk));
	jdff dff_A_Tp5ukWrU6_0(.dout(w_dff_A_bihMRFSc1_0),.din(w_dff_A_Tp5ukWrU6_0),.clk(gclk));
	jdff dff_A_PQHBQeQ88_0(.dout(w_dff_A_Tp5ukWrU6_0),.din(w_dff_A_PQHBQeQ88_0),.clk(gclk));
	jdff dff_A_6hKGXp2n6_0(.dout(w_dff_A_PQHBQeQ88_0),.din(w_dff_A_6hKGXp2n6_0),.clk(gclk));
	jdff dff_A_2hLXjuSt9_0(.dout(w_dff_A_6hKGXp2n6_0),.din(w_dff_A_2hLXjuSt9_0),.clk(gclk));
	jdff dff_A_VT9uk01s8_0(.dout(w_dff_A_2hLXjuSt9_0),.din(w_dff_A_VT9uk01s8_0),.clk(gclk));
	jdff dff_A_ba218ma79_0(.dout(w_dff_A_VT9uk01s8_0),.din(w_dff_A_ba218ma79_0),.clk(gclk));
	jdff dff_A_LH6i8iDf7_0(.dout(w_dff_A_ba218ma79_0),.din(w_dff_A_LH6i8iDf7_0),.clk(gclk));
	jdff dff_A_k0fnviVx3_0(.dout(w_dff_A_LH6i8iDf7_0),.din(w_dff_A_k0fnviVx3_0),.clk(gclk));
	jdff dff_A_pcNzs3g52_0(.dout(w_dff_A_k0fnviVx3_0),.din(w_dff_A_pcNzs3g52_0),.clk(gclk));
	jdff dff_A_SKeRgjCD9_0(.dout(w_dff_A_pcNzs3g52_0),.din(w_dff_A_SKeRgjCD9_0),.clk(gclk));
	jdff dff_A_DlXmu2b54_0(.dout(w_dff_A_SKeRgjCD9_0),.din(w_dff_A_DlXmu2b54_0),.clk(gclk));
	jdff dff_A_IcQ1nQXP5_0(.dout(w_dff_A_DlXmu2b54_0),.din(w_dff_A_IcQ1nQXP5_0),.clk(gclk));
	jdff dff_A_9j7mjvKU0_0(.dout(w_dff_A_IcQ1nQXP5_0),.din(w_dff_A_9j7mjvKU0_0),.clk(gclk));
	jdff dff_A_isWUtwEk6_0(.dout(w_dff_A_9j7mjvKU0_0),.din(w_dff_A_isWUtwEk6_0),.clk(gclk));
	jdff dff_A_c2KFI1wt8_0(.dout(w_dff_A_isWUtwEk6_0),.din(w_dff_A_c2KFI1wt8_0),.clk(gclk));
	jdff dff_A_zUYihYQ72_0(.dout(w_dff_A_c2KFI1wt8_0),.din(w_dff_A_zUYihYQ72_0),.clk(gclk));
	jdff dff_A_S80ML2T33_0(.dout(w_dff_A_zUYihYQ72_0),.din(w_dff_A_S80ML2T33_0),.clk(gclk));
	jdff dff_A_2kzZNoJ95_0(.dout(w_dff_A_S80ML2T33_0),.din(w_dff_A_2kzZNoJ95_0),.clk(gclk));
	jdff dff_A_uwNEA9JR7_0(.dout(w_dff_A_2kzZNoJ95_0),.din(w_dff_A_uwNEA9JR7_0),.clk(gclk));
	jdff dff_A_zMfLwwtg2_0(.dout(w_dff_A_uwNEA9JR7_0),.din(w_dff_A_zMfLwwtg2_0),.clk(gclk));
	jdff dff_A_MKBp2C5v8_0(.dout(w_dff_A_zMfLwwtg2_0),.din(w_dff_A_MKBp2C5v8_0),.clk(gclk));
	jdff dff_A_nLBL5pzN6_0(.dout(w_dff_A_MKBp2C5v8_0),.din(w_dff_A_nLBL5pzN6_0),.clk(gclk));
	jdff dff_A_YLBwudag3_0(.dout(w_dff_A_nLBL5pzN6_0),.din(w_dff_A_YLBwudag3_0),.clk(gclk));
	jdff dff_A_R4ZeTc807_0(.dout(w_dff_A_YLBwudag3_0),.din(w_dff_A_R4ZeTc807_0),.clk(gclk));
	jdff dff_A_q8tDLDGG5_1(.dout(w_n468_0[1]),.din(w_dff_A_q8tDLDGG5_1),.clk(gclk));
	jdff dff_B_ZL5VaW9n3_1(.din(n406),.dout(w_dff_B_ZL5VaW9n3_1),.clk(gclk));
	jdff dff_B_JsJNkWNH7_1(.din(w_dff_B_ZL5VaW9n3_1),.dout(w_dff_B_JsJNkWNH7_1),.clk(gclk));
	jdff dff_B_dEhn0jED6_1(.din(w_dff_B_JsJNkWNH7_1),.dout(w_dff_B_dEhn0jED6_1),.clk(gclk));
	jdff dff_B_7dYbH2lr6_1(.din(w_dff_B_dEhn0jED6_1),.dout(w_dff_B_7dYbH2lr6_1),.clk(gclk));
	jdff dff_B_WAvn0rNU6_1(.din(w_dff_B_7dYbH2lr6_1),.dout(w_dff_B_WAvn0rNU6_1),.clk(gclk));
	jdff dff_B_2qcrzXlP2_1(.din(w_dff_B_WAvn0rNU6_1),.dout(w_dff_B_2qcrzXlP2_1),.clk(gclk));
	jdff dff_B_qqCwWwgw5_1(.din(w_dff_B_2qcrzXlP2_1),.dout(w_dff_B_qqCwWwgw5_1),.clk(gclk));
	jdff dff_B_D7WDdV4b2_1(.din(w_dff_B_qqCwWwgw5_1),.dout(w_dff_B_D7WDdV4b2_1),.clk(gclk));
	jdff dff_B_Vfe8ybqM6_1(.din(w_dff_B_D7WDdV4b2_1),.dout(w_dff_B_Vfe8ybqM6_1),.clk(gclk));
	jdff dff_B_Vm90iu193_1(.din(w_dff_B_Vfe8ybqM6_1),.dout(w_dff_B_Vm90iu193_1),.clk(gclk));
	jdff dff_B_gplyiiRe7_1(.din(w_dff_B_Vm90iu193_1),.dout(w_dff_B_gplyiiRe7_1),.clk(gclk));
	jdff dff_B_tPqXlddp7_1(.din(w_dff_B_gplyiiRe7_1),.dout(w_dff_B_tPqXlddp7_1),.clk(gclk));
	jdff dff_B_KIn84tUX8_1(.din(w_dff_B_tPqXlddp7_1),.dout(w_dff_B_KIn84tUX8_1),.clk(gclk));
	jdff dff_B_gdAerqbx6_1(.din(w_dff_B_KIn84tUX8_1),.dout(w_dff_B_gdAerqbx6_1),.clk(gclk));
	jdff dff_B_X6cvKOX49_1(.din(w_dff_B_gdAerqbx6_1),.dout(w_dff_B_X6cvKOX49_1),.clk(gclk));
	jdff dff_B_QauYEzdS0_1(.din(w_dff_B_X6cvKOX49_1),.dout(w_dff_B_QauYEzdS0_1),.clk(gclk));
	jdff dff_B_dftS0TZo7_1(.din(w_dff_B_QauYEzdS0_1),.dout(w_dff_B_dftS0TZo7_1),.clk(gclk));
	jdff dff_B_1q90oM0k9_1(.din(w_dff_B_dftS0TZo7_1),.dout(w_dff_B_1q90oM0k9_1),.clk(gclk));
	jdff dff_B_AoFvBdpB5_1(.din(w_dff_B_1q90oM0k9_1),.dout(w_dff_B_AoFvBdpB5_1),.clk(gclk));
	jdff dff_B_KFqcFrUX6_1(.din(w_dff_B_AoFvBdpB5_1),.dout(w_dff_B_KFqcFrUX6_1),.clk(gclk));
	jdff dff_B_RRU6Zs145_1(.din(w_dff_B_KFqcFrUX6_1),.dout(w_dff_B_RRU6Zs145_1),.clk(gclk));
	jdff dff_B_WPcY44fS0_1(.din(w_dff_B_RRU6Zs145_1),.dout(w_dff_B_WPcY44fS0_1),.clk(gclk));
	jdff dff_B_UlbgQ8MC5_1(.din(w_dff_B_WPcY44fS0_1),.dout(w_dff_B_UlbgQ8MC5_1),.clk(gclk));
	jdff dff_B_gzwSsxYP3_1(.din(w_dff_B_UlbgQ8MC5_1),.dout(w_dff_B_gzwSsxYP3_1),.clk(gclk));
	jdff dff_B_vfMFIONK9_1(.din(w_dff_B_gzwSsxYP3_1),.dout(w_dff_B_vfMFIONK9_1),.clk(gclk));
	jdff dff_B_r79Ag4N17_1(.din(n402),.dout(w_dff_B_r79Ag4N17_1),.clk(gclk));
	jdff dff_A_07XvEf3d4_0(.dout(w_n335_0[0]),.din(w_dff_A_07XvEf3d4_0),.clk(gclk));
	jdff dff_A_S71DeJ4S7_0(.dout(w_dff_A_07XvEf3d4_0),.din(w_dff_A_S71DeJ4S7_0),.clk(gclk));
	jdff dff_A_AyP7AboR5_0(.dout(w_dff_A_S71DeJ4S7_0),.din(w_dff_A_AyP7AboR5_0),.clk(gclk));
	jdff dff_A_1RfPkj7S2_0(.dout(w_dff_A_AyP7AboR5_0),.din(w_dff_A_1RfPkj7S2_0),.clk(gclk));
	jdff dff_A_3JrGAypj5_0(.dout(w_dff_A_1RfPkj7S2_0),.din(w_dff_A_3JrGAypj5_0),.clk(gclk));
	jdff dff_A_SGAlmRUy8_0(.dout(w_dff_A_3JrGAypj5_0),.din(w_dff_A_SGAlmRUy8_0),.clk(gclk));
	jdff dff_A_vRWkMEVA7_0(.dout(w_dff_A_SGAlmRUy8_0),.din(w_dff_A_vRWkMEVA7_0),.clk(gclk));
	jdff dff_A_eYZc56bQ0_0(.dout(w_dff_A_vRWkMEVA7_0),.din(w_dff_A_eYZc56bQ0_0),.clk(gclk));
	jdff dff_A_AL1Jq1aZ1_0(.dout(w_dff_A_eYZc56bQ0_0),.din(w_dff_A_AL1Jq1aZ1_0),.clk(gclk));
	jdff dff_A_tiCsG0FA5_0(.dout(w_dff_A_AL1Jq1aZ1_0),.din(w_dff_A_tiCsG0FA5_0),.clk(gclk));
	jdff dff_A_ZM8KHHC41_0(.dout(w_dff_A_tiCsG0FA5_0),.din(w_dff_A_ZM8KHHC41_0),.clk(gclk));
	jdff dff_A_yG9RquUF1_0(.dout(w_dff_A_ZM8KHHC41_0),.din(w_dff_A_yG9RquUF1_0),.clk(gclk));
	jdff dff_A_BQAGjrTr2_0(.dout(w_dff_A_yG9RquUF1_0),.din(w_dff_A_BQAGjrTr2_0),.clk(gclk));
	jdff dff_A_VKyZLDAL4_0(.dout(w_dff_A_BQAGjrTr2_0),.din(w_dff_A_VKyZLDAL4_0),.clk(gclk));
	jdff dff_A_sXRZKFtq1_0(.dout(w_dff_A_VKyZLDAL4_0),.din(w_dff_A_sXRZKFtq1_0),.clk(gclk));
	jdff dff_A_WcV7LFru5_0(.dout(w_dff_A_sXRZKFtq1_0),.din(w_dff_A_WcV7LFru5_0),.clk(gclk));
	jdff dff_A_KyVO6UQE1_0(.dout(w_dff_A_WcV7LFru5_0),.din(w_dff_A_KyVO6UQE1_0),.clk(gclk));
	jdff dff_A_bADsdaOd3_0(.dout(w_dff_A_KyVO6UQE1_0),.din(w_dff_A_bADsdaOd3_0),.clk(gclk));
	jdff dff_A_VaKaZm7P5_0(.dout(w_dff_A_bADsdaOd3_0),.din(w_dff_A_VaKaZm7P5_0),.clk(gclk));
	jdff dff_A_iQtCWTZW2_0(.dout(w_dff_A_VaKaZm7P5_0),.din(w_dff_A_iQtCWTZW2_0),.clk(gclk));
	jdff dff_A_9rJU7ldF3_0(.dout(w_dff_A_iQtCWTZW2_0),.din(w_dff_A_9rJU7ldF3_0),.clk(gclk));
	jdff dff_A_BOGCJ2fr5_0(.dout(w_dff_A_9rJU7ldF3_0),.din(w_dff_A_BOGCJ2fr5_0),.clk(gclk));
	jdff dff_A_3yB3pTCZ0_0(.dout(w_dff_A_BOGCJ2fr5_0),.din(w_dff_A_3yB3pTCZ0_0),.clk(gclk));
	jdff dff_A_pedVWmIY0_0(.dout(w_dff_A_3yB3pTCZ0_0),.din(w_dff_A_pedVWmIY0_0),.clk(gclk));
	jdff dff_A_rxJ6Gxda0_0(.dout(w_dff_A_pedVWmIY0_0),.din(w_dff_A_rxJ6Gxda0_0),.clk(gclk));
	jdff dff_A_KQ2O2otq9_0(.dout(w_dff_A_rxJ6Gxda0_0),.din(w_dff_A_KQ2O2otq9_0),.clk(gclk));
	jdff dff_A_pdtZY1cb0_1(.dout(w_n396_0[1]),.din(w_dff_A_pdtZY1cb0_1),.clk(gclk));
	jdff dff_B_uaji9XrL9_1(.din(n342),.dout(w_dff_B_uaji9XrL9_1),.clk(gclk));
	jdff dff_B_V2XGEC8k2_1(.din(w_dff_B_uaji9XrL9_1),.dout(w_dff_B_V2XGEC8k2_1),.clk(gclk));
	jdff dff_B_8ddoDOuH7_1(.din(w_dff_B_V2XGEC8k2_1),.dout(w_dff_B_8ddoDOuH7_1),.clk(gclk));
	jdff dff_B_MzbcbGUO3_1(.din(w_dff_B_8ddoDOuH7_1),.dout(w_dff_B_MzbcbGUO3_1),.clk(gclk));
	jdff dff_B_3nXnYQNm5_1(.din(w_dff_B_MzbcbGUO3_1),.dout(w_dff_B_3nXnYQNm5_1),.clk(gclk));
	jdff dff_B_3DZjDbuJ3_1(.din(w_dff_B_3nXnYQNm5_1),.dout(w_dff_B_3DZjDbuJ3_1),.clk(gclk));
	jdff dff_B_zEBeWXrs6_1(.din(w_dff_B_3DZjDbuJ3_1),.dout(w_dff_B_zEBeWXrs6_1),.clk(gclk));
	jdff dff_B_7u9uNGiF4_1(.din(w_dff_B_zEBeWXrs6_1),.dout(w_dff_B_7u9uNGiF4_1),.clk(gclk));
	jdff dff_B_iC2ahARG7_1(.din(w_dff_B_7u9uNGiF4_1),.dout(w_dff_B_iC2ahARG7_1),.clk(gclk));
	jdff dff_B_B77UuNaF2_1(.din(w_dff_B_iC2ahARG7_1),.dout(w_dff_B_B77UuNaF2_1),.clk(gclk));
	jdff dff_B_7NcS5zV68_1(.din(w_dff_B_B77UuNaF2_1),.dout(w_dff_B_7NcS5zV68_1),.clk(gclk));
	jdff dff_B_6n4SH0qe0_1(.din(w_dff_B_7NcS5zV68_1),.dout(w_dff_B_6n4SH0qe0_1),.clk(gclk));
	jdff dff_B_z1Jwm19L5_1(.din(w_dff_B_6n4SH0qe0_1),.dout(w_dff_B_z1Jwm19L5_1),.clk(gclk));
	jdff dff_B_DNVYFIAU3_1(.din(w_dff_B_z1Jwm19L5_1),.dout(w_dff_B_DNVYFIAU3_1),.clk(gclk));
	jdff dff_B_T3LTlcff9_1(.din(w_dff_B_DNVYFIAU3_1),.dout(w_dff_B_T3LTlcff9_1),.clk(gclk));
	jdff dff_B_LHX2JYat5_1(.din(w_dff_B_T3LTlcff9_1),.dout(w_dff_B_LHX2JYat5_1),.clk(gclk));
	jdff dff_B_48TZ66Tv1_1(.din(w_dff_B_LHX2JYat5_1),.dout(w_dff_B_48TZ66Tv1_1),.clk(gclk));
	jdff dff_B_RnpQ5oW77_1(.din(w_dff_B_48TZ66Tv1_1),.dout(w_dff_B_RnpQ5oW77_1),.clk(gclk));
	jdff dff_B_KQtljAQK4_1(.din(w_dff_B_RnpQ5oW77_1),.dout(w_dff_B_KQtljAQK4_1),.clk(gclk));
	jdff dff_B_0kHpSL6g5_1(.din(w_dff_B_KQtljAQK4_1),.dout(w_dff_B_0kHpSL6g5_1),.clk(gclk));
	jdff dff_B_cwlt9MPQ2_1(.din(w_dff_B_0kHpSL6g5_1),.dout(w_dff_B_cwlt9MPQ2_1),.clk(gclk));
	jdff dff_B_9zhxnigc6_1(.din(w_dff_B_cwlt9MPQ2_1),.dout(w_dff_B_9zhxnigc6_1),.clk(gclk));
	jdff dff_B_G2a9mku59_1(.din(n338),.dout(w_dff_B_G2a9mku59_1),.clk(gclk));
	jdff dff_A_WNAubkdK7_0(.dout(w_n277_0[0]),.din(w_dff_A_WNAubkdK7_0),.clk(gclk));
	jdff dff_A_Gko9mBMh7_0(.dout(w_dff_A_WNAubkdK7_0),.din(w_dff_A_Gko9mBMh7_0),.clk(gclk));
	jdff dff_A_PnNbR9Vs1_0(.dout(w_dff_A_Gko9mBMh7_0),.din(w_dff_A_PnNbR9Vs1_0),.clk(gclk));
	jdff dff_A_4tqugQMX6_0(.dout(w_dff_A_PnNbR9Vs1_0),.din(w_dff_A_4tqugQMX6_0),.clk(gclk));
	jdff dff_A_VOBEbYy45_0(.dout(w_dff_A_4tqugQMX6_0),.din(w_dff_A_VOBEbYy45_0),.clk(gclk));
	jdff dff_A_PKufTHoC4_0(.dout(w_dff_A_VOBEbYy45_0),.din(w_dff_A_PKufTHoC4_0),.clk(gclk));
	jdff dff_A_pOyXgVy32_0(.dout(w_dff_A_PKufTHoC4_0),.din(w_dff_A_pOyXgVy32_0),.clk(gclk));
	jdff dff_A_EiDPqxd47_0(.dout(w_dff_A_pOyXgVy32_0),.din(w_dff_A_EiDPqxd47_0),.clk(gclk));
	jdff dff_A_onxi8iqR4_0(.dout(w_dff_A_EiDPqxd47_0),.din(w_dff_A_onxi8iqR4_0),.clk(gclk));
	jdff dff_A_36dRa3KG5_0(.dout(w_dff_A_onxi8iqR4_0),.din(w_dff_A_36dRa3KG5_0),.clk(gclk));
	jdff dff_A_HQNQH4wm9_0(.dout(w_dff_A_36dRa3KG5_0),.din(w_dff_A_HQNQH4wm9_0),.clk(gclk));
	jdff dff_A_1utdlHDO5_0(.dout(w_dff_A_HQNQH4wm9_0),.din(w_dff_A_1utdlHDO5_0),.clk(gclk));
	jdff dff_A_TOHpIvxF1_0(.dout(w_dff_A_1utdlHDO5_0),.din(w_dff_A_TOHpIvxF1_0),.clk(gclk));
	jdff dff_A_Kujq2QhY2_0(.dout(w_dff_A_TOHpIvxF1_0),.din(w_dff_A_Kujq2QhY2_0),.clk(gclk));
	jdff dff_A_kKiCe1CS3_0(.dout(w_dff_A_Kujq2QhY2_0),.din(w_dff_A_kKiCe1CS3_0),.clk(gclk));
	jdff dff_A_AyFQGTNA1_0(.dout(w_dff_A_kKiCe1CS3_0),.din(w_dff_A_AyFQGTNA1_0),.clk(gclk));
	jdff dff_A_gIufiRDE7_0(.dout(w_dff_A_AyFQGTNA1_0),.din(w_dff_A_gIufiRDE7_0),.clk(gclk));
	jdff dff_A_YDtrAI5W8_0(.dout(w_dff_A_gIufiRDE7_0),.din(w_dff_A_YDtrAI5W8_0),.clk(gclk));
	jdff dff_A_yoD1KkwS9_0(.dout(w_dff_A_YDtrAI5W8_0),.din(w_dff_A_yoD1KkwS9_0),.clk(gclk));
	jdff dff_A_61wkXLfz2_0(.dout(w_dff_A_yoD1KkwS9_0),.din(w_dff_A_61wkXLfz2_0),.clk(gclk));
	jdff dff_A_M9Vj75ie0_0(.dout(w_dff_A_61wkXLfz2_0),.din(w_dff_A_M9Vj75ie0_0),.clk(gclk));
	jdff dff_A_Yi0R7pV94_0(.dout(w_dff_A_M9Vj75ie0_0),.din(w_dff_A_Yi0R7pV94_0),.clk(gclk));
	jdff dff_A_NzASmWdC1_0(.dout(w_dff_A_Yi0R7pV94_0),.din(w_dff_A_NzASmWdC1_0),.clk(gclk));
	jdff dff_A_ZBNkQBen1_1(.dout(w_n332_0[1]),.din(w_dff_A_ZBNkQBen1_1),.clk(gclk));
	jdff dff_B_sQHggNVV2_1(.din(n284),.dout(w_dff_B_sQHggNVV2_1),.clk(gclk));
	jdff dff_B_0a2EIjzn2_1(.din(w_dff_B_sQHggNVV2_1),.dout(w_dff_B_0a2EIjzn2_1),.clk(gclk));
	jdff dff_B_g74iP5qI6_1(.din(w_dff_B_0a2EIjzn2_1),.dout(w_dff_B_g74iP5qI6_1),.clk(gclk));
	jdff dff_B_mgLSvAeH6_1(.din(w_dff_B_g74iP5qI6_1),.dout(w_dff_B_mgLSvAeH6_1),.clk(gclk));
	jdff dff_B_TpEiFXiZ6_1(.din(w_dff_B_mgLSvAeH6_1),.dout(w_dff_B_TpEiFXiZ6_1),.clk(gclk));
	jdff dff_B_tDN3qfWj5_1(.din(w_dff_B_TpEiFXiZ6_1),.dout(w_dff_B_tDN3qfWj5_1),.clk(gclk));
	jdff dff_B_3JPPXOvh9_1(.din(w_dff_B_tDN3qfWj5_1),.dout(w_dff_B_3JPPXOvh9_1),.clk(gclk));
	jdff dff_B_UtoxWck83_1(.din(w_dff_B_3JPPXOvh9_1),.dout(w_dff_B_UtoxWck83_1),.clk(gclk));
	jdff dff_B_2yGWQ7121_1(.din(w_dff_B_UtoxWck83_1),.dout(w_dff_B_2yGWQ7121_1),.clk(gclk));
	jdff dff_B_jB9nM9qL7_1(.din(w_dff_B_2yGWQ7121_1),.dout(w_dff_B_jB9nM9qL7_1),.clk(gclk));
	jdff dff_B_FARCtiGb1_1(.din(w_dff_B_jB9nM9qL7_1),.dout(w_dff_B_FARCtiGb1_1),.clk(gclk));
	jdff dff_B_giBP00WZ2_1(.din(w_dff_B_FARCtiGb1_1),.dout(w_dff_B_giBP00WZ2_1),.clk(gclk));
	jdff dff_B_VwapzuL72_1(.din(w_dff_B_giBP00WZ2_1),.dout(w_dff_B_VwapzuL72_1),.clk(gclk));
	jdff dff_B_HmBmlcBA0_1(.din(w_dff_B_VwapzuL72_1),.dout(w_dff_B_HmBmlcBA0_1),.clk(gclk));
	jdff dff_B_mrciLR6N7_1(.din(w_dff_B_HmBmlcBA0_1),.dout(w_dff_B_mrciLR6N7_1),.clk(gclk));
	jdff dff_B_GSMkC0mH3_1(.din(w_dff_B_mrciLR6N7_1),.dout(w_dff_B_GSMkC0mH3_1),.clk(gclk));
	jdff dff_B_guxh1W8Y9_1(.din(w_dff_B_GSMkC0mH3_1),.dout(w_dff_B_guxh1W8Y9_1),.clk(gclk));
	jdff dff_B_RVtFTpM18_1(.din(w_dff_B_guxh1W8Y9_1),.dout(w_dff_B_RVtFTpM18_1),.clk(gclk));
	jdff dff_B_1NeGTeA62_1(.din(w_dff_B_RVtFTpM18_1),.dout(w_dff_B_1NeGTeA62_1),.clk(gclk));
	jdff dff_B_EtRKUMoM0_1(.din(n280),.dout(w_dff_B_EtRKUMoM0_1),.clk(gclk));
	jdff dff_A_yd2wSgOJ3_0(.dout(w_n226_0[0]),.din(w_dff_A_yd2wSgOJ3_0),.clk(gclk));
	jdff dff_A_dTud4PkE8_0(.dout(w_dff_A_yd2wSgOJ3_0),.din(w_dff_A_dTud4PkE8_0),.clk(gclk));
	jdff dff_A_16Otk0LG3_0(.dout(w_dff_A_dTud4PkE8_0),.din(w_dff_A_16Otk0LG3_0),.clk(gclk));
	jdff dff_A_VrZ2eqAD3_0(.dout(w_dff_A_16Otk0LG3_0),.din(w_dff_A_VrZ2eqAD3_0),.clk(gclk));
	jdff dff_A_394mG6D45_0(.dout(w_dff_A_VrZ2eqAD3_0),.din(w_dff_A_394mG6D45_0),.clk(gclk));
	jdff dff_A_CcPw8DQa1_0(.dout(w_dff_A_394mG6D45_0),.din(w_dff_A_CcPw8DQa1_0),.clk(gclk));
	jdff dff_A_8zxqr1RF4_0(.dout(w_dff_A_CcPw8DQa1_0),.din(w_dff_A_8zxqr1RF4_0),.clk(gclk));
	jdff dff_A_8INlV0gl9_0(.dout(w_dff_A_8zxqr1RF4_0),.din(w_dff_A_8INlV0gl9_0),.clk(gclk));
	jdff dff_A_B8Ldhac90_0(.dout(w_dff_A_8INlV0gl9_0),.din(w_dff_A_B8Ldhac90_0),.clk(gclk));
	jdff dff_A_KQZqEpd62_0(.dout(w_dff_A_B8Ldhac90_0),.din(w_dff_A_KQZqEpd62_0),.clk(gclk));
	jdff dff_A_PSu4PeRC0_0(.dout(w_dff_A_KQZqEpd62_0),.din(w_dff_A_PSu4PeRC0_0),.clk(gclk));
	jdff dff_A_MxZaryhj4_0(.dout(w_dff_A_PSu4PeRC0_0),.din(w_dff_A_MxZaryhj4_0),.clk(gclk));
	jdff dff_A_PaFBBoOj8_0(.dout(w_dff_A_MxZaryhj4_0),.din(w_dff_A_PaFBBoOj8_0),.clk(gclk));
	jdff dff_A_2Vf80ylI8_0(.dout(w_dff_A_PaFBBoOj8_0),.din(w_dff_A_2Vf80ylI8_0),.clk(gclk));
	jdff dff_A_gFaHzqXF3_0(.dout(w_dff_A_2Vf80ylI8_0),.din(w_dff_A_gFaHzqXF3_0),.clk(gclk));
	jdff dff_A_rsFsgka31_0(.dout(w_dff_A_gFaHzqXF3_0),.din(w_dff_A_rsFsgka31_0),.clk(gclk));
	jdff dff_A_47xJSKVp3_0(.dout(w_dff_A_rsFsgka31_0),.din(w_dff_A_47xJSKVp3_0),.clk(gclk));
	jdff dff_A_EbhXl6AE0_0(.dout(w_dff_A_47xJSKVp3_0),.din(w_dff_A_EbhXl6AE0_0),.clk(gclk));
	jdff dff_A_mADN9N8V2_0(.dout(w_dff_A_EbhXl6AE0_0),.din(w_dff_A_mADN9N8V2_0),.clk(gclk));
	jdff dff_A_JPXdPWUu5_0(.dout(w_dff_A_mADN9N8V2_0),.din(w_dff_A_JPXdPWUu5_0),.clk(gclk));
	jdff dff_A_dd2KuOew4_1(.dout(w_n274_0[1]),.din(w_dff_A_dd2KuOew4_1),.clk(gclk));
	jdff dff_B_F1mXoP8m7_1(.din(n233),.dout(w_dff_B_F1mXoP8m7_1),.clk(gclk));
	jdff dff_B_cnK0nCHN4_1(.din(w_dff_B_F1mXoP8m7_1),.dout(w_dff_B_cnK0nCHN4_1),.clk(gclk));
	jdff dff_B_mtYEvDP34_1(.din(w_dff_B_cnK0nCHN4_1),.dout(w_dff_B_mtYEvDP34_1),.clk(gclk));
	jdff dff_B_qzSAt64H2_1(.din(w_dff_B_mtYEvDP34_1),.dout(w_dff_B_qzSAt64H2_1),.clk(gclk));
	jdff dff_B_InDJSpJP6_1(.din(w_dff_B_qzSAt64H2_1),.dout(w_dff_B_InDJSpJP6_1),.clk(gclk));
	jdff dff_B_e9LzUf0S0_1(.din(w_dff_B_InDJSpJP6_1),.dout(w_dff_B_e9LzUf0S0_1),.clk(gclk));
	jdff dff_B_yttmxCRk8_1(.din(w_dff_B_e9LzUf0S0_1),.dout(w_dff_B_yttmxCRk8_1),.clk(gclk));
	jdff dff_B_3JdfAORd1_1(.din(w_dff_B_yttmxCRk8_1),.dout(w_dff_B_3JdfAORd1_1),.clk(gclk));
	jdff dff_B_fpJaDYb26_1(.din(w_dff_B_3JdfAORd1_1),.dout(w_dff_B_fpJaDYb26_1),.clk(gclk));
	jdff dff_B_RU9jkWQh0_1(.din(w_dff_B_fpJaDYb26_1),.dout(w_dff_B_RU9jkWQh0_1),.clk(gclk));
	jdff dff_B_9u5QYrI36_1(.din(w_dff_B_RU9jkWQh0_1),.dout(w_dff_B_9u5QYrI36_1),.clk(gclk));
	jdff dff_B_A51qYh7k0_1(.din(w_dff_B_9u5QYrI36_1),.dout(w_dff_B_A51qYh7k0_1),.clk(gclk));
	jdff dff_B_5wXpyIlb9_1(.din(w_dff_B_A51qYh7k0_1),.dout(w_dff_B_5wXpyIlb9_1),.clk(gclk));
	jdff dff_B_n6hjHG9P8_1(.din(w_dff_B_5wXpyIlb9_1),.dout(w_dff_B_n6hjHG9P8_1),.clk(gclk));
	jdff dff_B_ghI2TLLK7_1(.din(w_dff_B_n6hjHG9P8_1),.dout(w_dff_B_ghI2TLLK7_1),.clk(gclk));
	jdff dff_B_2sGGj5117_1(.din(w_dff_B_ghI2TLLK7_1),.dout(w_dff_B_2sGGj5117_1),.clk(gclk));
	jdff dff_B_MLjx4sMy3_1(.din(n229),.dout(w_dff_B_MLjx4sMy3_1),.clk(gclk));
	jdff dff_A_jIPo6DQn7_0(.dout(w_n183_0[0]),.din(w_dff_A_jIPo6DQn7_0),.clk(gclk));
	jdff dff_A_BEoNHnEm8_0(.dout(w_dff_A_jIPo6DQn7_0),.din(w_dff_A_BEoNHnEm8_0),.clk(gclk));
	jdff dff_A_UoeXRQNw2_0(.dout(w_dff_A_BEoNHnEm8_0),.din(w_dff_A_UoeXRQNw2_0),.clk(gclk));
	jdff dff_A_jgtar52N4_0(.dout(w_dff_A_UoeXRQNw2_0),.din(w_dff_A_jgtar52N4_0),.clk(gclk));
	jdff dff_A_qSSw6ntj5_0(.dout(w_dff_A_jgtar52N4_0),.din(w_dff_A_qSSw6ntj5_0),.clk(gclk));
	jdff dff_A_T7JiqPbL0_0(.dout(w_dff_A_qSSw6ntj5_0),.din(w_dff_A_T7JiqPbL0_0),.clk(gclk));
	jdff dff_A_tgdsUr972_0(.dout(w_dff_A_T7JiqPbL0_0),.din(w_dff_A_tgdsUr972_0),.clk(gclk));
	jdff dff_A_MYKZjBnC5_0(.dout(w_dff_A_tgdsUr972_0),.din(w_dff_A_MYKZjBnC5_0),.clk(gclk));
	jdff dff_A_X2TWBBO39_0(.dout(w_dff_A_MYKZjBnC5_0),.din(w_dff_A_X2TWBBO39_0),.clk(gclk));
	jdff dff_A_tdEjQUA01_0(.dout(w_dff_A_X2TWBBO39_0),.din(w_dff_A_tdEjQUA01_0),.clk(gclk));
	jdff dff_A_rkvro7cG4_0(.dout(w_dff_A_tdEjQUA01_0),.din(w_dff_A_rkvro7cG4_0),.clk(gclk));
	jdff dff_A_ckoPgMau3_0(.dout(w_dff_A_rkvro7cG4_0),.din(w_dff_A_ckoPgMau3_0),.clk(gclk));
	jdff dff_A_FghHqTZj2_0(.dout(w_dff_A_ckoPgMau3_0),.din(w_dff_A_FghHqTZj2_0),.clk(gclk));
	jdff dff_A_J97Nnlbp0_0(.dout(w_dff_A_FghHqTZj2_0),.din(w_dff_A_J97Nnlbp0_0),.clk(gclk));
	jdff dff_A_JJYQDiXV5_0(.dout(w_dff_A_J97Nnlbp0_0),.din(w_dff_A_JJYQDiXV5_0),.clk(gclk));
	jdff dff_A_6zj07BYk5_0(.dout(w_dff_A_JJYQDiXV5_0),.din(w_dff_A_6zj07BYk5_0),.clk(gclk));
	jdff dff_A_wIZmNCxX4_0(.dout(w_dff_A_6zj07BYk5_0),.din(w_dff_A_wIZmNCxX4_0),.clk(gclk));
	jdff dff_A_G11zUqc14_1(.dout(w_n223_0[1]),.din(w_dff_A_G11zUqc14_1),.clk(gclk));
	jdff dff_B_msPiOmBT6_1(.din(n190),.dout(w_dff_B_msPiOmBT6_1),.clk(gclk));
	jdff dff_B_9K8Fc5g41_1(.din(w_dff_B_msPiOmBT6_1),.dout(w_dff_B_9K8Fc5g41_1),.clk(gclk));
	jdff dff_B_7Y8ID8hz4_1(.din(w_dff_B_9K8Fc5g41_1),.dout(w_dff_B_7Y8ID8hz4_1),.clk(gclk));
	jdff dff_B_m7TJb8T42_1(.din(w_dff_B_7Y8ID8hz4_1),.dout(w_dff_B_m7TJb8T42_1),.clk(gclk));
	jdff dff_B_KjcKKkyc3_1(.din(w_dff_B_m7TJb8T42_1),.dout(w_dff_B_KjcKKkyc3_1),.clk(gclk));
	jdff dff_B_XOmIvBiT7_1(.din(w_dff_B_KjcKKkyc3_1),.dout(w_dff_B_XOmIvBiT7_1),.clk(gclk));
	jdff dff_B_b4BIqd5J5_1(.din(w_dff_B_XOmIvBiT7_1),.dout(w_dff_B_b4BIqd5J5_1),.clk(gclk));
	jdff dff_B_QlSxxFjz7_1(.din(w_dff_B_b4BIqd5J5_1),.dout(w_dff_B_QlSxxFjz7_1),.clk(gclk));
	jdff dff_B_uMAiGIYJ8_1(.din(w_dff_B_QlSxxFjz7_1),.dout(w_dff_B_uMAiGIYJ8_1),.clk(gclk));
	jdff dff_B_FUD1bpmc2_1(.din(w_dff_B_uMAiGIYJ8_1),.dout(w_dff_B_FUD1bpmc2_1),.clk(gclk));
	jdff dff_B_whOG2x2d8_1(.din(w_dff_B_FUD1bpmc2_1),.dout(w_dff_B_whOG2x2d8_1),.clk(gclk));
	jdff dff_B_5vO4kvi22_1(.din(w_dff_B_whOG2x2d8_1),.dout(w_dff_B_5vO4kvi22_1),.clk(gclk));
	jdff dff_B_TzMqASIS7_1(.din(w_dff_B_5vO4kvi22_1),.dout(w_dff_B_TzMqASIS7_1),.clk(gclk));
	jdff dff_B_pbsMynBF6_1(.din(n186),.dout(w_dff_B_pbsMynBF6_1),.clk(gclk));
	jdff dff_A_1zRpXd2X4_0(.dout(w_n145_0[0]),.din(w_dff_A_1zRpXd2X4_0),.clk(gclk));
	jdff dff_A_rMclxszd8_0(.dout(w_dff_A_1zRpXd2X4_0),.din(w_dff_A_rMclxszd8_0),.clk(gclk));
	jdff dff_A_X7OvdmMJ0_0(.dout(w_dff_A_rMclxszd8_0),.din(w_dff_A_X7OvdmMJ0_0),.clk(gclk));
	jdff dff_A_pOInmols4_0(.dout(w_dff_A_X7OvdmMJ0_0),.din(w_dff_A_pOInmols4_0),.clk(gclk));
	jdff dff_A_LydU78NP4_0(.dout(w_dff_A_pOInmols4_0),.din(w_dff_A_LydU78NP4_0),.clk(gclk));
	jdff dff_A_fgn7zzmi1_0(.dout(w_dff_A_LydU78NP4_0),.din(w_dff_A_fgn7zzmi1_0),.clk(gclk));
	jdff dff_A_3UFqp5xG1_0(.dout(w_dff_A_fgn7zzmi1_0),.din(w_dff_A_3UFqp5xG1_0),.clk(gclk));
	jdff dff_A_rbqVl4It0_0(.dout(w_dff_A_3UFqp5xG1_0),.din(w_dff_A_rbqVl4It0_0),.clk(gclk));
	jdff dff_A_Ve2xpuXI7_0(.dout(w_dff_A_rbqVl4It0_0),.din(w_dff_A_Ve2xpuXI7_0),.clk(gclk));
	jdff dff_A_bIJGbnrZ6_0(.dout(w_dff_A_Ve2xpuXI7_0),.din(w_dff_A_bIJGbnrZ6_0),.clk(gclk));
	jdff dff_A_R8xzFM1X6_0(.dout(w_dff_A_bIJGbnrZ6_0),.din(w_dff_A_R8xzFM1X6_0),.clk(gclk));
	jdff dff_A_WbyxWmyk1_0(.dout(w_dff_A_R8xzFM1X6_0),.din(w_dff_A_WbyxWmyk1_0),.clk(gclk));
	jdff dff_A_c8emaS972_0(.dout(w_dff_A_WbyxWmyk1_0),.din(w_dff_A_c8emaS972_0),.clk(gclk));
	jdff dff_A_vuvYPKsd0_0(.dout(w_dff_A_c8emaS972_0),.din(w_dff_A_vuvYPKsd0_0),.clk(gclk));
	jdff dff_A_abjFZba61_1(.dout(w_n180_0[1]),.din(w_dff_A_abjFZba61_1),.clk(gclk));
	jdff dff_B_znPVCf3g9_1(.din(n152),.dout(w_dff_B_znPVCf3g9_1),.clk(gclk));
	jdff dff_B_uTY9VtKv1_1(.din(w_dff_B_znPVCf3g9_1),.dout(w_dff_B_uTY9VtKv1_1),.clk(gclk));
	jdff dff_B_QvttyXg92_1(.din(w_dff_B_uTY9VtKv1_1),.dout(w_dff_B_QvttyXg92_1),.clk(gclk));
	jdff dff_B_ow2AcIkY8_1(.din(w_dff_B_QvttyXg92_1),.dout(w_dff_B_ow2AcIkY8_1),.clk(gclk));
	jdff dff_B_VsT4Cj7R0_1(.din(w_dff_B_ow2AcIkY8_1),.dout(w_dff_B_VsT4Cj7R0_1),.clk(gclk));
	jdff dff_B_kPhGAsQz8_1(.din(w_dff_B_VsT4Cj7R0_1),.dout(w_dff_B_kPhGAsQz8_1),.clk(gclk));
	jdff dff_B_sephocXF6_1(.din(w_dff_B_kPhGAsQz8_1),.dout(w_dff_B_sephocXF6_1),.clk(gclk));
	jdff dff_B_7IqEQ2Rw3_1(.din(w_dff_B_sephocXF6_1),.dout(w_dff_B_7IqEQ2Rw3_1),.clk(gclk));
	jdff dff_B_R7Ngk5aT2_1(.din(w_dff_B_7IqEQ2Rw3_1),.dout(w_dff_B_R7Ngk5aT2_1),.clk(gclk));
	jdff dff_B_Y8lCDkCI6_1(.din(w_dff_B_R7Ngk5aT2_1),.dout(w_dff_B_Y8lCDkCI6_1),.clk(gclk));
	jdff dff_B_3eb8cAjZ3_1(.din(n148),.dout(w_dff_B_3eb8cAjZ3_1),.clk(gclk));
	jdff dff_A_1yPGyo8y2_0(.dout(w_n110_0[0]),.din(w_dff_A_1yPGyo8y2_0),.clk(gclk));
	jdff dff_A_EjRqAhi79_0(.dout(w_dff_A_1yPGyo8y2_0),.din(w_dff_A_EjRqAhi79_0),.clk(gclk));
	jdff dff_A_JIpqIlhj3_0(.dout(w_dff_A_EjRqAhi79_0),.din(w_dff_A_JIpqIlhj3_0),.clk(gclk));
	jdff dff_A_tzommCdL5_0(.dout(w_dff_A_JIpqIlhj3_0),.din(w_dff_A_tzommCdL5_0),.clk(gclk));
	jdff dff_A_LIEnoCqY8_0(.dout(w_dff_A_tzommCdL5_0),.din(w_dff_A_LIEnoCqY8_0),.clk(gclk));
	jdff dff_A_gHrsytin8_0(.dout(w_dff_A_LIEnoCqY8_0),.din(w_dff_A_gHrsytin8_0),.clk(gclk));
	jdff dff_A_fT46BE4Z8_0(.dout(w_dff_A_gHrsytin8_0),.din(w_dff_A_fT46BE4Z8_0),.clk(gclk));
	jdff dff_A_aFpAwGkv1_0(.dout(w_dff_A_fT46BE4Z8_0),.din(w_dff_A_aFpAwGkv1_0),.clk(gclk));
	jdff dff_A_K3J3VhNi6_0(.dout(w_dff_A_aFpAwGkv1_0),.din(w_dff_A_K3J3VhNi6_0),.clk(gclk));
	jdff dff_A_jdGnuqf83_0(.dout(w_dff_A_K3J3VhNi6_0),.din(w_dff_A_jdGnuqf83_0),.clk(gclk));
	jdff dff_A_EVKqHyce1_0(.dout(w_dff_A_jdGnuqf83_0),.din(w_dff_A_EVKqHyce1_0),.clk(gclk));
	jdff dff_A_Bw9625kf4_1(.dout(w_n142_0[1]),.din(w_dff_A_Bw9625kf4_1),.clk(gclk));
	jdff dff_B_5lTOWi381_1(.din(n117),.dout(w_dff_B_5lTOWi381_1),.clk(gclk));
	jdff dff_B_nKOywrTp7_1(.din(w_dff_B_5lTOWi381_1),.dout(w_dff_B_nKOywrTp7_1),.clk(gclk));
	jdff dff_B_ivFGV6Zl1_1(.din(w_dff_B_nKOywrTp7_1),.dout(w_dff_B_ivFGV6Zl1_1),.clk(gclk));
	jdff dff_B_Oeuj6ZRK6_1(.din(w_dff_B_ivFGV6Zl1_1),.dout(w_dff_B_Oeuj6ZRK6_1),.clk(gclk));
	jdff dff_B_YknQjzgM1_1(.din(w_dff_B_Oeuj6ZRK6_1),.dout(w_dff_B_YknQjzgM1_1),.clk(gclk));
	jdff dff_B_4ez6oAxy9_1(.din(w_dff_B_YknQjzgM1_1),.dout(w_dff_B_4ez6oAxy9_1),.clk(gclk));
	jdff dff_B_z5yrB3Ls7_1(.din(w_dff_B_4ez6oAxy9_1),.dout(w_dff_B_z5yrB3Ls7_1),.clk(gclk));
	jdff dff_B_xBBblVJN9_1(.din(n113),.dout(w_dff_B_xBBblVJN9_1),.clk(gclk));
	jdff dff_A_O17b2fkp1_0(.dout(w_n89_0[0]),.din(w_dff_A_O17b2fkp1_0),.clk(gclk));
	jdff dff_A_Y4F5XlY71_0(.dout(w_dff_A_O17b2fkp1_0),.din(w_dff_A_Y4F5XlY71_0),.clk(gclk));
	jdff dff_A_fUs8N7ld7_0(.dout(w_dff_A_Y4F5XlY71_0),.din(w_dff_A_fUs8N7ld7_0),.clk(gclk));
	jdff dff_A_MMsPaLNi4_0(.dout(w_dff_A_fUs8N7ld7_0),.din(w_dff_A_MMsPaLNi4_0),.clk(gclk));
	jdff dff_A_OVUgk53k2_0(.dout(w_dff_A_MMsPaLNi4_0),.din(w_dff_A_OVUgk53k2_0),.clk(gclk));
	jdff dff_A_R6l0TgAt6_0(.dout(w_dff_A_OVUgk53k2_0),.din(w_dff_A_R6l0TgAt6_0),.clk(gclk));
	jdff dff_A_VzizVc8V0_0(.dout(w_dff_A_R6l0TgAt6_0),.din(w_dff_A_VzizVc8V0_0),.clk(gclk));
	jdff dff_A_kiy2BO7f5_0(.dout(w_dff_A_VzizVc8V0_0),.din(w_dff_A_kiy2BO7f5_0),.clk(gclk));
	jdff dff_A_4iAploSe2_1(.dout(w_n107_0[1]),.din(w_dff_A_4iAploSe2_1),.clk(gclk));
	jdff dff_B_xhEpL6TF3_1(.din(n95),.dout(w_dff_B_xhEpL6TF3_1),.clk(gclk));
	jdff dff_B_G4j0ydwA7_1(.din(w_dff_B_xhEpL6TF3_1),.dout(w_dff_B_G4j0ydwA7_1),.clk(gclk));
	jdff dff_B_KJVIe0q63_1(.din(w_dff_B_G4j0ydwA7_1),.dout(w_dff_B_KJVIe0q63_1),.clk(gclk));
	jdff dff_B_Mc0qdUx74_1(.din(w_dff_B_KJVIe0q63_1),.dout(w_dff_B_Mc0qdUx74_1),.clk(gclk));
	jdff dff_B_s2BIrOrl5_1(.din(n91),.dout(w_dff_B_s2BIrOrl5_1),.clk(gclk));
	jdff dff_B_PSo8MNph8_0(.din(n86),.dout(w_dff_B_PSo8MNph8_0),.clk(gclk));
	jdff dff_A_TcIp6Mog2_0(.dout(w_n72_0[0]),.din(w_dff_A_TcIp6Mog2_0),.clk(gclk));
	jdff dff_A_sRvmt9jy6_0(.dout(w_dff_A_TcIp6Mog2_0),.din(w_dff_A_sRvmt9jy6_0),.clk(gclk));
	jdff dff_A_butF18JX5_0(.dout(w_dff_A_sRvmt9jy6_0),.din(w_dff_A_butF18JX5_0),.clk(gclk));
	jdff dff_A_1Eby9pJV6_0(.dout(w_dff_A_butF18JX5_0),.din(w_dff_A_1Eby9pJV6_0),.clk(gclk));
	jdff dff_A_OX7nFsGl7_0(.dout(w_dff_A_1Eby9pJV6_0),.din(w_dff_A_OX7nFsGl7_0),.clk(gclk));
	jdff dff_A_x31Ir6Po7_0(.dout(w_n70_0[0]),.din(w_dff_A_x31Ir6Po7_0),.clk(gclk));
	jdff dff_A_YDMEMreQ6_0(.dout(w_n69_0[0]),.din(w_dff_A_YDMEMreQ6_0),.clk(gclk));
	jdff dff_A_ZxkjIyrc9_1(.dout(w_n1140_0[1]),.din(w_dff_A_ZxkjIyrc9_1),.clk(gclk));
	jdff dff_B_RiwhK7vq5_1(.din(n1040),.dout(w_dff_B_RiwhK7vq5_1),.clk(gclk));
	jdff dff_B_wlm8K5mf0_2(.din(n938),.dout(w_dff_B_wlm8K5mf0_2),.clk(gclk));
	jdff dff_B_9DyEIpxU0_2(.din(w_dff_B_wlm8K5mf0_2),.dout(w_dff_B_9DyEIpxU0_2),.clk(gclk));
	jdff dff_B_QOBEJ13A7_2(.din(w_dff_B_9DyEIpxU0_2),.dout(w_dff_B_QOBEJ13A7_2),.clk(gclk));
	jdff dff_B_eKOMNCZY4_2(.din(w_dff_B_QOBEJ13A7_2),.dout(w_dff_B_eKOMNCZY4_2),.clk(gclk));
	jdff dff_B_IHNDThLe2_2(.din(w_dff_B_eKOMNCZY4_2),.dout(w_dff_B_IHNDThLe2_2),.clk(gclk));
	jdff dff_B_DO2laoWd9_2(.din(w_dff_B_IHNDThLe2_2),.dout(w_dff_B_DO2laoWd9_2),.clk(gclk));
	jdff dff_B_3ILXNG2K0_2(.din(w_dff_B_DO2laoWd9_2),.dout(w_dff_B_3ILXNG2K0_2),.clk(gclk));
	jdff dff_B_XwxPcHRt9_2(.din(w_dff_B_3ILXNG2K0_2),.dout(w_dff_B_XwxPcHRt9_2),.clk(gclk));
	jdff dff_B_cWQYjVO54_2(.din(w_dff_B_XwxPcHRt9_2),.dout(w_dff_B_cWQYjVO54_2),.clk(gclk));
	jdff dff_B_u4zv1JeY5_2(.din(w_dff_B_cWQYjVO54_2),.dout(w_dff_B_u4zv1JeY5_2),.clk(gclk));
	jdff dff_B_Mfvhq5wL2_2(.din(w_dff_B_u4zv1JeY5_2),.dout(w_dff_B_Mfvhq5wL2_2),.clk(gclk));
	jdff dff_B_7k9eOmYL7_2(.din(w_dff_B_Mfvhq5wL2_2),.dout(w_dff_B_7k9eOmYL7_2),.clk(gclk));
	jdff dff_B_zqDm2X7C0_2(.din(w_dff_B_7k9eOmYL7_2),.dout(w_dff_B_zqDm2X7C0_2),.clk(gclk));
	jdff dff_B_bsSSdUYK4_2(.din(w_dff_B_zqDm2X7C0_2),.dout(w_dff_B_bsSSdUYK4_2),.clk(gclk));
	jdff dff_B_fAI1qAow0_2(.din(w_dff_B_bsSSdUYK4_2),.dout(w_dff_B_fAI1qAow0_2),.clk(gclk));
	jdff dff_B_pDPQ9iTi9_2(.din(w_dff_B_fAI1qAow0_2),.dout(w_dff_B_pDPQ9iTi9_2),.clk(gclk));
	jdff dff_B_JjtxkxWH7_2(.din(w_dff_B_pDPQ9iTi9_2),.dout(w_dff_B_JjtxkxWH7_2),.clk(gclk));
	jdff dff_B_TrlfOvVw6_2(.din(w_dff_B_JjtxkxWH7_2),.dout(w_dff_B_TrlfOvVw6_2),.clk(gclk));
	jdff dff_B_mxlSVfqZ6_2(.din(w_dff_B_TrlfOvVw6_2),.dout(w_dff_B_mxlSVfqZ6_2),.clk(gclk));
	jdff dff_B_p0eQka6R1_2(.din(w_dff_B_mxlSVfqZ6_2),.dout(w_dff_B_p0eQka6R1_2),.clk(gclk));
	jdff dff_B_nuCChVu33_2(.din(w_dff_B_p0eQka6R1_2),.dout(w_dff_B_nuCChVu33_2),.clk(gclk));
	jdff dff_B_M68hpCGC0_2(.din(w_dff_B_nuCChVu33_2),.dout(w_dff_B_M68hpCGC0_2),.clk(gclk));
	jdff dff_B_3EgGeu4s0_2(.din(w_dff_B_M68hpCGC0_2),.dout(w_dff_B_3EgGeu4s0_2),.clk(gclk));
	jdff dff_B_TBLieZRy2_2(.din(w_dff_B_3EgGeu4s0_2),.dout(w_dff_B_TBLieZRy2_2),.clk(gclk));
	jdff dff_B_u2iHJdBs5_2(.din(w_dff_B_TBLieZRy2_2),.dout(w_dff_B_u2iHJdBs5_2),.clk(gclk));
	jdff dff_B_BMsMvpkg9_2(.din(w_dff_B_u2iHJdBs5_2),.dout(w_dff_B_BMsMvpkg9_2),.clk(gclk));
	jdff dff_B_LvuS2iwE2_2(.din(w_dff_B_BMsMvpkg9_2),.dout(w_dff_B_LvuS2iwE2_2),.clk(gclk));
	jdff dff_B_2I2ldc0Q1_2(.din(w_dff_B_LvuS2iwE2_2),.dout(w_dff_B_2I2ldc0Q1_2),.clk(gclk));
	jdff dff_B_ZT3XjHeo4_2(.din(w_dff_B_2I2ldc0Q1_2),.dout(w_dff_B_ZT3XjHeo4_2),.clk(gclk));
	jdff dff_B_bvi7awdg8_2(.din(w_dff_B_ZT3XjHeo4_2),.dout(w_dff_B_bvi7awdg8_2),.clk(gclk));
	jdff dff_B_rocixNWt1_2(.din(w_dff_B_bvi7awdg8_2),.dout(w_dff_B_rocixNWt1_2),.clk(gclk));
	jdff dff_B_Su9B3HDt0_2(.din(w_dff_B_rocixNWt1_2),.dout(w_dff_B_Su9B3HDt0_2),.clk(gclk));
	jdff dff_B_RJTu95gr9_2(.din(w_dff_B_Su9B3HDt0_2),.dout(w_dff_B_RJTu95gr9_2),.clk(gclk));
	jdff dff_B_vuVW65hV3_2(.din(w_dff_B_RJTu95gr9_2),.dout(w_dff_B_vuVW65hV3_2),.clk(gclk));
	jdff dff_B_GpdtCDhE0_2(.din(w_dff_B_vuVW65hV3_2),.dout(w_dff_B_GpdtCDhE0_2),.clk(gclk));
	jdff dff_B_EtbdMEIt7_2(.din(w_dff_B_GpdtCDhE0_2),.dout(w_dff_B_EtbdMEIt7_2),.clk(gclk));
	jdff dff_B_gL9dlKkl5_2(.din(w_dff_B_EtbdMEIt7_2),.dout(w_dff_B_gL9dlKkl5_2),.clk(gclk));
	jdff dff_B_wbzRpzcA5_2(.din(w_dff_B_gL9dlKkl5_2),.dout(w_dff_B_wbzRpzcA5_2),.clk(gclk));
	jdff dff_B_iVbP97Cc2_2(.din(w_dff_B_wbzRpzcA5_2),.dout(w_dff_B_iVbP97Cc2_2),.clk(gclk));
	jdff dff_B_NNZxI4Y85_2(.din(w_dff_B_iVbP97Cc2_2),.dout(w_dff_B_NNZxI4Y85_2),.clk(gclk));
	jdff dff_B_zO54pNgP7_2(.din(w_dff_B_NNZxI4Y85_2),.dout(w_dff_B_zO54pNgP7_2),.clk(gclk));
	jdff dff_B_zxiSrnG13_2(.din(w_dff_B_zO54pNgP7_2),.dout(w_dff_B_zxiSrnG13_2),.clk(gclk));
	jdff dff_B_Vlr8Yz1X6_2(.din(w_dff_B_zxiSrnG13_2),.dout(w_dff_B_Vlr8Yz1X6_2),.clk(gclk));
	jdff dff_B_wKqaqs3V7_2(.din(w_dff_B_Vlr8Yz1X6_2),.dout(w_dff_B_wKqaqs3V7_2),.clk(gclk));
	jdff dff_A_oCU1WYQG2_0(.dout(w_n1034_0[0]),.din(w_dff_A_oCU1WYQG2_0),.clk(gclk));
	jdff dff_B_sU9bcwMw6_1(.din(n940),.dout(w_dff_B_sU9bcwMw6_1),.clk(gclk));
	jdff dff_B_VJypzdYV9_2(.din(n835),.dout(w_dff_B_VJypzdYV9_2),.clk(gclk));
	jdff dff_B_Y2k4OLYn9_2(.din(w_dff_B_VJypzdYV9_2),.dout(w_dff_B_Y2k4OLYn9_2),.clk(gclk));
	jdff dff_B_BjMOCRay1_2(.din(w_dff_B_Y2k4OLYn9_2),.dout(w_dff_B_BjMOCRay1_2),.clk(gclk));
	jdff dff_B_imY2ErmR9_2(.din(w_dff_B_BjMOCRay1_2),.dout(w_dff_B_imY2ErmR9_2),.clk(gclk));
	jdff dff_B_TY4unhCk6_2(.din(w_dff_B_imY2ErmR9_2),.dout(w_dff_B_TY4unhCk6_2),.clk(gclk));
	jdff dff_B_7gY5SbKn7_2(.din(w_dff_B_TY4unhCk6_2),.dout(w_dff_B_7gY5SbKn7_2),.clk(gclk));
	jdff dff_B_7WMmc1Q55_2(.din(w_dff_B_7gY5SbKn7_2),.dout(w_dff_B_7WMmc1Q55_2),.clk(gclk));
	jdff dff_B_Z7pnereq8_2(.din(w_dff_B_7WMmc1Q55_2),.dout(w_dff_B_Z7pnereq8_2),.clk(gclk));
	jdff dff_B_uky2RO3m1_2(.din(w_dff_B_Z7pnereq8_2),.dout(w_dff_B_uky2RO3m1_2),.clk(gclk));
	jdff dff_B_WCkNCACs6_2(.din(w_dff_B_uky2RO3m1_2),.dout(w_dff_B_WCkNCACs6_2),.clk(gclk));
	jdff dff_B_skYH6HWA4_2(.din(w_dff_B_WCkNCACs6_2),.dout(w_dff_B_skYH6HWA4_2),.clk(gclk));
	jdff dff_B_DDRNHVOi9_2(.din(w_dff_B_skYH6HWA4_2),.dout(w_dff_B_DDRNHVOi9_2),.clk(gclk));
	jdff dff_B_IfW36s7h2_2(.din(w_dff_B_DDRNHVOi9_2),.dout(w_dff_B_IfW36s7h2_2),.clk(gclk));
	jdff dff_B_wZmO0LWb3_2(.din(w_dff_B_IfW36s7h2_2),.dout(w_dff_B_wZmO0LWb3_2),.clk(gclk));
	jdff dff_B_CfzwRqWY3_2(.din(w_dff_B_wZmO0LWb3_2),.dout(w_dff_B_CfzwRqWY3_2),.clk(gclk));
	jdff dff_B_tqabiXk82_2(.din(w_dff_B_CfzwRqWY3_2),.dout(w_dff_B_tqabiXk82_2),.clk(gclk));
	jdff dff_B_Y9CPakYO9_2(.din(w_dff_B_tqabiXk82_2),.dout(w_dff_B_Y9CPakYO9_2),.clk(gclk));
	jdff dff_B_v9p8bOxX9_2(.din(w_dff_B_Y9CPakYO9_2),.dout(w_dff_B_v9p8bOxX9_2),.clk(gclk));
	jdff dff_B_haKXbpP99_2(.din(w_dff_B_v9p8bOxX9_2),.dout(w_dff_B_haKXbpP99_2),.clk(gclk));
	jdff dff_B_udy1DNGD2_2(.din(w_dff_B_haKXbpP99_2),.dout(w_dff_B_udy1DNGD2_2),.clk(gclk));
	jdff dff_B_WKiDCyR22_2(.din(w_dff_B_udy1DNGD2_2),.dout(w_dff_B_WKiDCyR22_2),.clk(gclk));
	jdff dff_B_WlRhaTgl7_2(.din(w_dff_B_WKiDCyR22_2),.dout(w_dff_B_WlRhaTgl7_2),.clk(gclk));
	jdff dff_B_t5Hj2OAO4_2(.din(w_dff_B_WlRhaTgl7_2),.dout(w_dff_B_t5Hj2OAO4_2),.clk(gclk));
	jdff dff_B_4NhvaBxW3_2(.din(w_dff_B_t5Hj2OAO4_2),.dout(w_dff_B_4NhvaBxW3_2),.clk(gclk));
	jdff dff_B_UbmjPo4v2_2(.din(w_dff_B_4NhvaBxW3_2),.dout(w_dff_B_UbmjPo4v2_2),.clk(gclk));
	jdff dff_B_VczT7VEE2_2(.din(w_dff_B_UbmjPo4v2_2),.dout(w_dff_B_VczT7VEE2_2),.clk(gclk));
	jdff dff_B_cB3JZs4O7_2(.din(w_dff_B_VczT7VEE2_2),.dout(w_dff_B_cB3JZs4O7_2),.clk(gclk));
	jdff dff_B_2xd6d1XP0_2(.din(w_dff_B_cB3JZs4O7_2),.dout(w_dff_B_2xd6d1XP0_2),.clk(gclk));
	jdff dff_B_tOKVNuNH8_2(.din(w_dff_B_2xd6d1XP0_2),.dout(w_dff_B_tOKVNuNH8_2),.clk(gclk));
	jdff dff_B_LYhKJWIc2_2(.din(w_dff_B_tOKVNuNH8_2),.dout(w_dff_B_LYhKJWIc2_2),.clk(gclk));
	jdff dff_B_nBqCEzFN0_2(.din(w_dff_B_LYhKJWIc2_2),.dout(w_dff_B_nBqCEzFN0_2),.clk(gclk));
	jdff dff_B_84Bzju1Y5_2(.din(w_dff_B_nBqCEzFN0_2),.dout(w_dff_B_84Bzju1Y5_2),.clk(gclk));
	jdff dff_B_ynuEwP5C3_2(.din(w_dff_B_84Bzju1Y5_2),.dout(w_dff_B_ynuEwP5C3_2),.clk(gclk));
	jdff dff_B_k8s1KtEa8_2(.din(w_dff_B_ynuEwP5C3_2),.dout(w_dff_B_k8s1KtEa8_2),.clk(gclk));
	jdff dff_B_ayWRMvj83_2(.din(w_dff_B_k8s1KtEa8_2),.dout(w_dff_B_ayWRMvj83_2),.clk(gclk));
	jdff dff_B_sLv6jA1Q2_2(.din(w_dff_B_ayWRMvj83_2),.dout(w_dff_B_sLv6jA1Q2_2),.clk(gclk));
	jdff dff_B_p0TIb4wo2_2(.din(w_dff_B_sLv6jA1Q2_2),.dout(w_dff_B_p0TIb4wo2_2),.clk(gclk));
	jdff dff_B_PKqJBaaX4_2(.din(w_dff_B_p0TIb4wo2_2),.dout(w_dff_B_PKqJBaaX4_2),.clk(gclk));
	jdff dff_B_PuUXjBx90_2(.din(w_dff_B_PKqJBaaX4_2),.dout(w_dff_B_PuUXjBx90_2),.clk(gclk));
	jdff dff_B_ihQYhirz0_2(.din(w_dff_B_PuUXjBx90_2),.dout(w_dff_B_ihQYhirz0_2),.clk(gclk));
	jdff dff_B_AQetBEn90_2(.din(w_dff_B_ihQYhirz0_2),.dout(w_dff_B_AQetBEn90_2),.clk(gclk));
	jdff dff_A_cONBtyJ46_1(.dout(w_n929_0[1]),.din(w_dff_A_cONBtyJ46_1),.clk(gclk));
	jdff dff_B_AvjPNMHL6_1(.din(n841),.dout(w_dff_B_AvjPNMHL6_1),.clk(gclk));
	jdff dff_B_mqiQvk0p7_1(.din(w_dff_B_AvjPNMHL6_1),.dout(w_dff_B_mqiQvk0p7_1),.clk(gclk));
	jdff dff_B_acdaogRU1_1(.din(w_dff_B_mqiQvk0p7_1),.dout(w_dff_B_acdaogRU1_1),.clk(gclk));
	jdff dff_B_qgxLf77o2_1(.din(w_dff_B_acdaogRU1_1),.dout(w_dff_B_qgxLf77o2_1),.clk(gclk));
	jdff dff_B_fFsmRr6I2_1(.din(w_dff_B_qgxLf77o2_1),.dout(w_dff_B_fFsmRr6I2_1),.clk(gclk));
	jdff dff_B_jcUMisnA9_1(.din(w_dff_B_fFsmRr6I2_1),.dout(w_dff_B_jcUMisnA9_1),.clk(gclk));
	jdff dff_B_2eOApgTo6_1(.din(w_dff_B_jcUMisnA9_1),.dout(w_dff_B_2eOApgTo6_1),.clk(gclk));
	jdff dff_B_6scP1DdX7_1(.din(w_dff_B_2eOApgTo6_1),.dout(w_dff_B_6scP1DdX7_1),.clk(gclk));
	jdff dff_B_TSPbQ89E1_1(.din(w_dff_B_6scP1DdX7_1),.dout(w_dff_B_TSPbQ89E1_1),.clk(gclk));
	jdff dff_B_fGWUI9Tp2_1(.din(w_dff_B_TSPbQ89E1_1),.dout(w_dff_B_fGWUI9Tp2_1),.clk(gclk));
	jdff dff_B_M3u0kNba0_1(.din(w_dff_B_fGWUI9Tp2_1),.dout(w_dff_B_M3u0kNba0_1),.clk(gclk));
	jdff dff_B_VIQCteMv2_1(.din(w_dff_B_M3u0kNba0_1),.dout(w_dff_B_VIQCteMv2_1),.clk(gclk));
	jdff dff_B_SRQYIHw39_1(.din(w_dff_B_VIQCteMv2_1),.dout(w_dff_B_SRQYIHw39_1),.clk(gclk));
	jdff dff_B_MmkCkwgi4_1(.din(w_dff_B_SRQYIHw39_1),.dout(w_dff_B_MmkCkwgi4_1),.clk(gclk));
	jdff dff_B_lxBhCIgM5_1(.din(w_dff_B_MmkCkwgi4_1),.dout(w_dff_B_lxBhCIgM5_1),.clk(gclk));
	jdff dff_B_6ED25RvQ3_1(.din(w_dff_B_lxBhCIgM5_1),.dout(w_dff_B_6ED25RvQ3_1),.clk(gclk));
	jdff dff_B_WBldEzQT6_1(.din(w_dff_B_6ED25RvQ3_1),.dout(w_dff_B_WBldEzQT6_1),.clk(gclk));
	jdff dff_B_CPlagn032_1(.din(w_dff_B_WBldEzQT6_1),.dout(w_dff_B_CPlagn032_1),.clk(gclk));
	jdff dff_B_2DjvS6QV6_1(.din(w_dff_B_CPlagn032_1),.dout(w_dff_B_2DjvS6QV6_1),.clk(gclk));
	jdff dff_B_jmOwVMch1_1(.din(w_dff_B_2DjvS6QV6_1),.dout(w_dff_B_jmOwVMch1_1),.clk(gclk));
	jdff dff_B_MLvqnb6r0_1(.din(w_dff_B_jmOwVMch1_1),.dout(w_dff_B_MLvqnb6r0_1),.clk(gclk));
	jdff dff_B_xZtk7he16_1(.din(w_dff_B_MLvqnb6r0_1),.dout(w_dff_B_xZtk7he16_1),.clk(gclk));
	jdff dff_B_D1HSzlMy5_1(.din(w_dff_B_xZtk7he16_1),.dout(w_dff_B_D1HSzlMy5_1),.clk(gclk));
	jdff dff_B_USsH6uLG6_1(.din(w_dff_B_D1HSzlMy5_1),.dout(w_dff_B_USsH6uLG6_1),.clk(gclk));
	jdff dff_B_63BIwxNr4_1(.din(w_dff_B_USsH6uLG6_1),.dout(w_dff_B_63BIwxNr4_1),.clk(gclk));
	jdff dff_B_MkaGDmVJ4_1(.din(w_dff_B_63BIwxNr4_1),.dout(w_dff_B_MkaGDmVJ4_1),.clk(gclk));
	jdff dff_B_fzUX9pqF2_1(.din(w_dff_B_MkaGDmVJ4_1),.dout(w_dff_B_fzUX9pqF2_1),.clk(gclk));
	jdff dff_B_ZEqeuxXy8_1(.din(w_dff_B_fzUX9pqF2_1),.dout(w_dff_B_ZEqeuxXy8_1),.clk(gclk));
	jdff dff_B_YH8ylwvq8_1(.din(w_dff_B_ZEqeuxXy8_1),.dout(w_dff_B_YH8ylwvq8_1),.clk(gclk));
	jdff dff_B_bOLYBQKJ0_1(.din(w_dff_B_YH8ylwvq8_1),.dout(w_dff_B_bOLYBQKJ0_1),.clk(gclk));
	jdff dff_B_adV0flcJ0_1(.din(w_dff_B_bOLYBQKJ0_1),.dout(w_dff_B_adV0flcJ0_1),.clk(gclk));
	jdff dff_B_DPKHiAnn9_1(.din(w_dff_B_adV0flcJ0_1),.dout(w_dff_B_DPKHiAnn9_1),.clk(gclk));
	jdff dff_B_9NcFDRM84_1(.din(w_dff_B_DPKHiAnn9_1),.dout(w_dff_B_9NcFDRM84_1),.clk(gclk));
	jdff dff_B_n67DSODH3_1(.din(w_dff_B_9NcFDRM84_1),.dout(w_dff_B_n67DSODH3_1),.clk(gclk));
	jdff dff_B_7l2d7zuR9_1(.din(w_dff_B_n67DSODH3_1),.dout(w_dff_B_7l2d7zuR9_1),.clk(gclk));
	jdff dff_B_6DCynWGq4_1(.din(w_dff_B_7l2d7zuR9_1),.dout(w_dff_B_6DCynWGq4_1),.clk(gclk));
	jdff dff_B_7RVIsGbA0_1(.din(w_dff_B_6DCynWGq4_1),.dout(w_dff_B_7RVIsGbA0_1),.clk(gclk));
	jdff dff_B_ovdRJMmp2_1(.din(n836),.dout(w_dff_B_ovdRJMmp2_1),.clk(gclk));
	jdff dff_A_UVdQvCkA8_0(.dout(w_n735_0[0]),.din(w_dff_A_UVdQvCkA8_0),.clk(gclk));
	jdff dff_A_04aJCo1j7_0(.dout(w_dff_A_UVdQvCkA8_0),.din(w_dff_A_04aJCo1j7_0),.clk(gclk));
	jdff dff_A_UxLiuMz43_0(.dout(w_dff_A_04aJCo1j7_0),.din(w_dff_A_UxLiuMz43_0),.clk(gclk));
	jdff dff_A_KhvWNSVw3_0(.dout(w_dff_A_UxLiuMz43_0),.din(w_dff_A_KhvWNSVw3_0),.clk(gclk));
	jdff dff_A_ms6nHWDr4_0(.dout(w_dff_A_KhvWNSVw3_0),.din(w_dff_A_ms6nHWDr4_0),.clk(gclk));
	jdff dff_A_CIWGLgWw2_0(.dout(w_dff_A_ms6nHWDr4_0),.din(w_dff_A_CIWGLgWw2_0),.clk(gclk));
	jdff dff_A_xkzRNhBk4_0(.dout(w_dff_A_CIWGLgWw2_0),.din(w_dff_A_xkzRNhBk4_0),.clk(gclk));
	jdff dff_A_xTzD6xi55_0(.dout(w_dff_A_xkzRNhBk4_0),.din(w_dff_A_xTzD6xi55_0),.clk(gclk));
	jdff dff_A_lszBqshw8_0(.dout(w_dff_A_xTzD6xi55_0),.din(w_dff_A_lszBqshw8_0),.clk(gclk));
	jdff dff_A_BQj4aOpR2_0(.dout(w_dff_A_lszBqshw8_0),.din(w_dff_A_BQj4aOpR2_0),.clk(gclk));
	jdff dff_A_0xU5GpCO3_0(.dout(w_dff_A_BQj4aOpR2_0),.din(w_dff_A_0xU5GpCO3_0),.clk(gclk));
	jdff dff_A_Qv7ZXBIv3_0(.dout(w_dff_A_0xU5GpCO3_0),.din(w_dff_A_Qv7ZXBIv3_0),.clk(gclk));
	jdff dff_A_k7Df8nbQ4_0(.dout(w_dff_A_Qv7ZXBIv3_0),.din(w_dff_A_k7Df8nbQ4_0),.clk(gclk));
	jdff dff_A_QQiiX0Vu0_0(.dout(w_dff_A_k7Df8nbQ4_0),.din(w_dff_A_QQiiX0Vu0_0),.clk(gclk));
	jdff dff_A_9piMC1ul0_0(.dout(w_dff_A_QQiiX0Vu0_0),.din(w_dff_A_9piMC1ul0_0),.clk(gclk));
	jdff dff_A_6AQH89uj8_0(.dout(w_dff_A_9piMC1ul0_0),.din(w_dff_A_6AQH89uj8_0),.clk(gclk));
	jdff dff_A_4xNyVkIb0_0(.dout(w_dff_A_6AQH89uj8_0),.din(w_dff_A_4xNyVkIb0_0),.clk(gclk));
	jdff dff_A_6WqT3W6u4_0(.dout(w_dff_A_4xNyVkIb0_0),.din(w_dff_A_6WqT3W6u4_0),.clk(gclk));
	jdff dff_A_kiUOKrWm1_0(.dout(w_dff_A_6WqT3W6u4_0),.din(w_dff_A_kiUOKrWm1_0),.clk(gclk));
	jdff dff_A_AeuFT1PZ5_0(.dout(w_dff_A_kiUOKrWm1_0),.din(w_dff_A_AeuFT1PZ5_0),.clk(gclk));
	jdff dff_A_oa8WIHar6_0(.dout(w_dff_A_AeuFT1PZ5_0),.din(w_dff_A_oa8WIHar6_0),.clk(gclk));
	jdff dff_A_Fd0sMzLa5_0(.dout(w_dff_A_oa8WIHar6_0),.din(w_dff_A_Fd0sMzLa5_0),.clk(gclk));
	jdff dff_A_vOuxIzFn3_0(.dout(w_dff_A_Fd0sMzLa5_0),.din(w_dff_A_vOuxIzFn3_0),.clk(gclk));
	jdff dff_A_VdoUm5ic5_0(.dout(w_dff_A_vOuxIzFn3_0),.din(w_dff_A_VdoUm5ic5_0),.clk(gclk));
	jdff dff_A_WTkvgKrv1_0(.dout(w_dff_A_VdoUm5ic5_0),.din(w_dff_A_WTkvgKrv1_0),.clk(gclk));
	jdff dff_A_bp7H5e9c0_0(.dout(w_dff_A_WTkvgKrv1_0),.din(w_dff_A_bp7H5e9c0_0),.clk(gclk));
	jdff dff_A_u6MW3VeA7_0(.dout(w_dff_A_bp7H5e9c0_0),.din(w_dff_A_u6MW3VeA7_0),.clk(gclk));
	jdff dff_A_wMp9Fyq01_0(.dout(w_dff_A_u6MW3VeA7_0),.din(w_dff_A_wMp9Fyq01_0),.clk(gclk));
	jdff dff_A_qyK09UQA0_0(.dout(w_dff_A_wMp9Fyq01_0),.din(w_dff_A_qyK09UQA0_0),.clk(gclk));
	jdff dff_A_Vvrmtr2d3_0(.dout(w_dff_A_qyK09UQA0_0),.din(w_dff_A_Vvrmtr2d3_0),.clk(gclk));
	jdff dff_A_phSzcfPN8_0(.dout(w_dff_A_Vvrmtr2d3_0),.din(w_dff_A_phSzcfPN8_0),.clk(gclk));
	jdff dff_A_tDjoEEd31_0(.dout(w_dff_A_phSzcfPN8_0),.din(w_dff_A_tDjoEEd31_0),.clk(gclk));
	jdff dff_A_W39d1HSr2_0(.dout(w_dff_A_tDjoEEd31_0),.din(w_dff_A_W39d1HSr2_0),.clk(gclk));
	jdff dff_A_Amm4FCpX8_0(.dout(w_dff_A_W39d1HSr2_0),.din(w_dff_A_Amm4FCpX8_0),.clk(gclk));
	jdff dff_A_vqcRHNxM6_0(.dout(w_dff_A_Amm4FCpX8_0),.din(w_dff_A_vqcRHNxM6_0),.clk(gclk));
	jdff dff_A_r8hunF2l9_0(.dout(w_dff_A_vqcRHNxM6_0),.din(w_dff_A_r8hunF2l9_0),.clk(gclk));
	jdff dff_A_Mz91aW7g2_0(.dout(w_dff_A_r8hunF2l9_0),.din(w_dff_A_Mz91aW7g2_0),.clk(gclk));
	jdff dff_A_gv2XXJR31_0(.dout(w_dff_A_Mz91aW7g2_0),.din(w_dff_A_gv2XXJR31_0),.clk(gclk));
	jdff dff_A_pNJ353jV9_0(.dout(w_n823_0[0]),.din(w_dff_A_pNJ353jV9_0),.clk(gclk));
	jdff dff_B_EyD3ZNz90_1(.din(n737),.dout(w_dff_B_EyD3ZNz90_1),.clk(gclk));
	jdff dff_A_HuXg3usU8_0(.dout(w_n642_0[0]),.din(w_dff_A_HuXg3usU8_0),.clk(gclk));
	jdff dff_A_VhUgFByC0_0(.dout(w_dff_A_HuXg3usU8_0),.din(w_dff_A_VhUgFByC0_0),.clk(gclk));
	jdff dff_A_T8OBfhSl4_0(.dout(w_dff_A_VhUgFByC0_0),.din(w_dff_A_T8OBfhSl4_0),.clk(gclk));
	jdff dff_A_ZTw5wOAj9_0(.dout(w_dff_A_T8OBfhSl4_0),.din(w_dff_A_ZTw5wOAj9_0),.clk(gclk));
	jdff dff_A_Iq7nWvCZ3_0(.dout(w_dff_A_ZTw5wOAj9_0),.din(w_dff_A_Iq7nWvCZ3_0),.clk(gclk));
	jdff dff_A_yAVt7SLb7_0(.dout(w_dff_A_Iq7nWvCZ3_0),.din(w_dff_A_yAVt7SLb7_0),.clk(gclk));
	jdff dff_A_3T4qwT0d2_0(.dout(w_dff_A_yAVt7SLb7_0),.din(w_dff_A_3T4qwT0d2_0),.clk(gclk));
	jdff dff_A_tloxYKW44_0(.dout(w_dff_A_3T4qwT0d2_0),.din(w_dff_A_tloxYKW44_0),.clk(gclk));
	jdff dff_A_ICBfhIee0_0(.dout(w_dff_A_tloxYKW44_0),.din(w_dff_A_ICBfhIee0_0),.clk(gclk));
	jdff dff_A_6pWsmhI01_0(.dout(w_dff_A_ICBfhIee0_0),.din(w_dff_A_6pWsmhI01_0),.clk(gclk));
	jdff dff_A_OMfI1VVd3_0(.dout(w_dff_A_6pWsmhI01_0),.din(w_dff_A_OMfI1VVd3_0),.clk(gclk));
	jdff dff_A_31gBrAmU9_0(.dout(w_dff_A_OMfI1VVd3_0),.din(w_dff_A_31gBrAmU9_0),.clk(gclk));
	jdff dff_A_KYey5Sve1_0(.dout(w_dff_A_31gBrAmU9_0),.din(w_dff_A_KYey5Sve1_0),.clk(gclk));
	jdff dff_A_HVEucIQN2_0(.dout(w_dff_A_KYey5Sve1_0),.din(w_dff_A_HVEucIQN2_0),.clk(gclk));
	jdff dff_A_rkunZU9h1_0(.dout(w_dff_A_HVEucIQN2_0),.din(w_dff_A_rkunZU9h1_0),.clk(gclk));
	jdff dff_A_j1oYindC5_0(.dout(w_dff_A_rkunZU9h1_0),.din(w_dff_A_j1oYindC5_0),.clk(gclk));
	jdff dff_A_VYrKM87F3_0(.dout(w_dff_A_j1oYindC5_0),.din(w_dff_A_VYrKM87F3_0),.clk(gclk));
	jdff dff_A_EKz6TQDI9_0(.dout(w_dff_A_VYrKM87F3_0),.din(w_dff_A_EKz6TQDI9_0),.clk(gclk));
	jdff dff_A_f2mVVxbV6_0(.dout(w_dff_A_EKz6TQDI9_0),.din(w_dff_A_f2mVVxbV6_0),.clk(gclk));
	jdff dff_A_jLXU7hEw3_0(.dout(w_dff_A_f2mVVxbV6_0),.din(w_dff_A_jLXU7hEw3_0),.clk(gclk));
	jdff dff_A_Dh7TuOOs1_0(.dout(w_dff_A_jLXU7hEw3_0),.din(w_dff_A_Dh7TuOOs1_0),.clk(gclk));
	jdff dff_A_gee1VQJY0_0(.dout(w_dff_A_Dh7TuOOs1_0),.din(w_dff_A_gee1VQJY0_0),.clk(gclk));
	jdff dff_A_UiBaxkEB2_0(.dout(w_dff_A_gee1VQJY0_0),.din(w_dff_A_UiBaxkEB2_0),.clk(gclk));
	jdff dff_A_gF0DgSDn7_0(.dout(w_dff_A_UiBaxkEB2_0),.din(w_dff_A_gF0DgSDn7_0),.clk(gclk));
	jdff dff_A_5nJP6kj45_0(.dout(w_dff_A_gF0DgSDn7_0),.din(w_dff_A_5nJP6kj45_0),.clk(gclk));
	jdff dff_A_5YlSKAyw2_0(.dout(w_dff_A_5nJP6kj45_0),.din(w_dff_A_5YlSKAyw2_0),.clk(gclk));
	jdff dff_A_9UrDpWcG8_0(.dout(w_dff_A_5YlSKAyw2_0),.din(w_dff_A_9UrDpWcG8_0),.clk(gclk));
	jdff dff_A_0xb8Nnld4_0(.dout(w_dff_A_9UrDpWcG8_0),.din(w_dff_A_0xb8Nnld4_0),.clk(gclk));
	jdff dff_A_b0OUSrwL9_0(.dout(w_dff_A_0xb8Nnld4_0),.din(w_dff_A_b0OUSrwL9_0),.clk(gclk));
	jdff dff_A_tKVgjKau1_0(.dout(w_dff_A_b0OUSrwL9_0),.din(w_dff_A_tKVgjKau1_0),.clk(gclk));
	jdff dff_A_NhYBq0aE6_0(.dout(w_dff_A_tKVgjKau1_0),.din(w_dff_A_NhYBq0aE6_0),.clk(gclk));
	jdff dff_A_294attYK5_0(.dout(w_dff_A_NhYBq0aE6_0),.din(w_dff_A_294attYK5_0),.clk(gclk));
	jdff dff_A_tGA5ayuD0_0(.dout(w_dff_A_294attYK5_0),.din(w_dff_A_tGA5ayuD0_0),.clk(gclk));
	jdff dff_A_1U8j3zsV2_0(.dout(w_dff_A_tGA5ayuD0_0),.din(w_dff_A_1U8j3zsV2_0),.clk(gclk));
	jdff dff_A_KkeADDaJ8_0(.dout(w_dff_A_1U8j3zsV2_0),.din(w_dff_A_KkeADDaJ8_0),.clk(gclk));
	jdff dff_A_TUptm82n2_0(.dout(w_n723_0[0]),.din(w_dff_A_TUptm82n2_0),.clk(gclk));
	jdff dff_B_BZtiQIGW5_1(.din(n644),.dout(w_dff_B_BZtiQIGW5_1),.clk(gclk));
	jdff dff_A_YmDAWMXy9_0(.dout(w_n556_0[0]),.din(w_dff_A_YmDAWMXy9_0),.clk(gclk));
	jdff dff_A_3sjevCOi3_0(.dout(w_dff_A_YmDAWMXy9_0),.din(w_dff_A_3sjevCOi3_0),.clk(gclk));
	jdff dff_A_LuA94Ww84_0(.dout(w_dff_A_3sjevCOi3_0),.din(w_dff_A_LuA94Ww84_0),.clk(gclk));
	jdff dff_A_ZEFFbOkh0_0(.dout(w_dff_A_LuA94Ww84_0),.din(w_dff_A_ZEFFbOkh0_0),.clk(gclk));
	jdff dff_A_36Ksepbw6_0(.dout(w_dff_A_ZEFFbOkh0_0),.din(w_dff_A_36Ksepbw6_0),.clk(gclk));
	jdff dff_A_BqwJaW1i7_0(.dout(w_dff_A_36Ksepbw6_0),.din(w_dff_A_BqwJaW1i7_0),.clk(gclk));
	jdff dff_A_WV7QDBiF0_0(.dout(w_dff_A_BqwJaW1i7_0),.din(w_dff_A_WV7QDBiF0_0),.clk(gclk));
	jdff dff_A_Q9VywNaz5_0(.dout(w_dff_A_WV7QDBiF0_0),.din(w_dff_A_Q9VywNaz5_0),.clk(gclk));
	jdff dff_A_dRGyk5DL1_0(.dout(w_dff_A_Q9VywNaz5_0),.din(w_dff_A_dRGyk5DL1_0),.clk(gclk));
	jdff dff_A_a6JJmDOB4_0(.dout(w_dff_A_dRGyk5DL1_0),.din(w_dff_A_a6JJmDOB4_0),.clk(gclk));
	jdff dff_A_8sF6Pv531_0(.dout(w_dff_A_a6JJmDOB4_0),.din(w_dff_A_8sF6Pv531_0),.clk(gclk));
	jdff dff_A_PVGlaclK5_0(.dout(w_dff_A_8sF6Pv531_0),.din(w_dff_A_PVGlaclK5_0),.clk(gclk));
	jdff dff_A_AVHr9Sag9_0(.dout(w_dff_A_PVGlaclK5_0),.din(w_dff_A_AVHr9Sag9_0),.clk(gclk));
	jdff dff_A_9yEu5N526_0(.dout(w_dff_A_AVHr9Sag9_0),.din(w_dff_A_9yEu5N526_0),.clk(gclk));
	jdff dff_A_FFbwqjPf7_0(.dout(w_dff_A_9yEu5N526_0),.din(w_dff_A_FFbwqjPf7_0),.clk(gclk));
	jdff dff_A_BN9ZPw1b9_0(.dout(w_dff_A_FFbwqjPf7_0),.din(w_dff_A_BN9ZPw1b9_0),.clk(gclk));
	jdff dff_A_d622n9di5_0(.dout(w_dff_A_BN9ZPw1b9_0),.din(w_dff_A_d622n9di5_0),.clk(gclk));
	jdff dff_A_xxYF6zzz1_0(.dout(w_dff_A_d622n9di5_0),.din(w_dff_A_xxYF6zzz1_0),.clk(gclk));
	jdff dff_A_LwGpTb137_0(.dout(w_dff_A_xxYF6zzz1_0),.din(w_dff_A_LwGpTb137_0),.clk(gclk));
	jdff dff_A_B31UjaJ41_0(.dout(w_dff_A_LwGpTb137_0),.din(w_dff_A_B31UjaJ41_0),.clk(gclk));
	jdff dff_A_umLnOgFL4_0(.dout(w_dff_A_B31UjaJ41_0),.din(w_dff_A_umLnOgFL4_0),.clk(gclk));
	jdff dff_A_sjVppoKo5_0(.dout(w_dff_A_umLnOgFL4_0),.din(w_dff_A_sjVppoKo5_0),.clk(gclk));
	jdff dff_A_oGxl3qyH6_0(.dout(w_dff_A_sjVppoKo5_0),.din(w_dff_A_oGxl3qyH6_0),.clk(gclk));
	jdff dff_A_uK2dd1MW6_0(.dout(w_dff_A_oGxl3qyH6_0),.din(w_dff_A_uK2dd1MW6_0),.clk(gclk));
	jdff dff_A_og1RfghJ3_0(.dout(w_dff_A_uK2dd1MW6_0),.din(w_dff_A_og1RfghJ3_0),.clk(gclk));
	jdff dff_A_NBSdpVgE9_0(.dout(w_dff_A_og1RfghJ3_0),.din(w_dff_A_NBSdpVgE9_0),.clk(gclk));
	jdff dff_A_X2au5xLe7_0(.dout(w_dff_A_NBSdpVgE9_0),.din(w_dff_A_X2au5xLe7_0),.clk(gclk));
	jdff dff_A_faA1aRbu0_0(.dout(w_dff_A_X2au5xLe7_0),.din(w_dff_A_faA1aRbu0_0),.clk(gclk));
	jdff dff_A_uorRZza72_0(.dout(w_dff_A_faA1aRbu0_0),.din(w_dff_A_uorRZza72_0),.clk(gclk));
	jdff dff_A_sOpgKyRl1_0(.dout(w_dff_A_uorRZza72_0),.din(w_dff_A_sOpgKyRl1_0),.clk(gclk));
	jdff dff_A_HnJjiojV1_0(.dout(w_dff_A_sOpgKyRl1_0),.din(w_dff_A_HnJjiojV1_0),.clk(gclk));
	jdff dff_A_Jpe6BBw50_0(.dout(w_dff_A_HnJjiojV1_0),.din(w_dff_A_Jpe6BBw50_0),.clk(gclk));
	jdff dff_A_XG0hYoUi2_0(.dout(w_n630_0[0]),.din(w_dff_A_XG0hYoUi2_0),.clk(gclk));
	jdff dff_B_wMbzty9e4_1(.din(n558),.dout(w_dff_B_wMbzty9e4_1),.clk(gclk));
	jdff dff_A_KaHITHHw3_0(.dout(w_n477_0[0]),.din(w_dff_A_KaHITHHw3_0),.clk(gclk));
	jdff dff_A_YHcdlSYS8_0(.dout(w_dff_A_KaHITHHw3_0),.din(w_dff_A_YHcdlSYS8_0),.clk(gclk));
	jdff dff_A_71bnE8T27_0(.dout(w_dff_A_YHcdlSYS8_0),.din(w_dff_A_71bnE8T27_0),.clk(gclk));
	jdff dff_A_IcYZhxDj6_0(.dout(w_dff_A_71bnE8T27_0),.din(w_dff_A_IcYZhxDj6_0),.clk(gclk));
	jdff dff_A_MeUppa0m2_0(.dout(w_dff_A_IcYZhxDj6_0),.din(w_dff_A_MeUppa0m2_0),.clk(gclk));
	jdff dff_A_vDoUtolz6_0(.dout(w_dff_A_MeUppa0m2_0),.din(w_dff_A_vDoUtolz6_0),.clk(gclk));
	jdff dff_A_FtzTPT0R4_0(.dout(w_dff_A_vDoUtolz6_0),.din(w_dff_A_FtzTPT0R4_0),.clk(gclk));
	jdff dff_A_qkDOJSN16_0(.dout(w_dff_A_FtzTPT0R4_0),.din(w_dff_A_qkDOJSN16_0),.clk(gclk));
	jdff dff_A_Exg6Qtis6_0(.dout(w_dff_A_qkDOJSN16_0),.din(w_dff_A_Exg6Qtis6_0),.clk(gclk));
	jdff dff_A_w2w9PQBI8_0(.dout(w_dff_A_Exg6Qtis6_0),.din(w_dff_A_w2w9PQBI8_0),.clk(gclk));
	jdff dff_A_J2LgcBq67_0(.dout(w_dff_A_w2w9PQBI8_0),.din(w_dff_A_J2LgcBq67_0),.clk(gclk));
	jdff dff_A_DeMBVa2p6_0(.dout(w_dff_A_J2LgcBq67_0),.din(w_dff_A_DeMBVa2p6_0),.clk(gclk));
	jdff dff_A_dzqe0GZw0_0(.dout(w_dff_A_DeMBVa2p6_0),.din(w_dff_A_dzqe0GZw0_0),.clk(gclk));
	jdff dff_A_IcvYiBy34_0(.dout(w_dff_A_dzqe0GZw0_0),.din(w_dff_A_IcvYiBy34_0),.clk(gclk));
	jdff dff_A_t5ToewZA2_0(.dout(w_dff_A_IcvYiBy34_0),.din(w_dff_A_t5ToewZA2_0),.clk(gclk));
	jdff dff_A_5CZrI5LA4_0(.dout(w_dff_A_t5ToewZA2_0),.din(w_dff_A_5CZrI5LA4_0),.clk(gclk));
	jdff dff_A_AxmcDDgY1_0(.dout(w_dff_A_5CZrI5LA4_0),.din(w_dff_A_AxmcDDgY1_0),.clk(gclk));
	jdff dff_A_K7y1rP592_0(.dout(w_dff_A_AxmcDDgY1_0),.din(w_dff_A_K7y1rP592_0),.clk(gclk));
	jdff dff_A_MVOJowLq9_0(.dout(w_dff_A_K7y1rP592_0),.din(w_dff_A_MVOJowLq9_0),.clk(gclk));
	jdff dff_A_IAsHkHwr8_0(.dout(w_dff_A_MVOJowLq9_0),.din(w_dff_A_IAsHkHwr8_0),.clk(gclk));
	jdff dff_A_6Z8LPAIr1_0(.dout(w_dff_A_IAsHkHwr8_0),.din(w_dff_A_6Z8LPAIr1_0),.clk(gclk));
	jdff dff_A_rT5Ohd2b5_0(.dout(w_dff_A_6Z8LPAIr1_0),.din(w_dff_A_rT5Ohd2b5_0),.clk(gclk));
	jdff dff_A_zfIy0Op68_0(.dout(w_dff_A_rT5Ohd2b5_0),.din(w_dff_A_zfIy0Op68_0),.clk(gclk));
	jdff dff_A_z2sX11c36_0(.dout(w_dff_A_zfIy0Op68_0),.din(w_dff_A_z2sX11c36_0),.clk(gclk));
	jdff dff_A_XVEZyGxX8_0(.dout(w_dff_A_z2sX11c36_0),.din(w_dff_A_XVEZyGxX8_0),.clk(gclk));
	jdff dff_A_6oUrGpVr9_0(.dout(w_dff_A_XVEZyGxX8_0),.din(w_dff_A_6oUrGpVr9_0),.clk(gclk));
	jdff dff_A_vozhl1db5_0(.dout(w_dff_A_6oUrGpVr9_0),.din(w_dff_A_vozhl1db5_0),.clk(gclk));
	jdff dff_A_AX55zDq92_0(.dout(w_dff_A_vozhl1db5_0),.din(w_dff_A_AX55zDq92_0),.clk(gclk));
	jdff dff_A_VqxSOFmS0_0(.dout(w_dff_A_AX55zDq92_0),.din(w_dff_A_VqxSOFmS0_0),.clk(gclk));
	jdff dff_A_2N5I4kY78_0(.dout(w_n544_0[0]),.din(w_dff_A_2N5I4kY78_0),.clk(gclk));
	jdff dff_B_FEoRVAiC6_1(.din(n479),.dout(w_dff_B_FEoRVAiC6_1),.clk(gclk));
	jdff dff_A_rSSfFkGL7_0(.dout(w_n405_0[0]),.din(w_dff_A_rSSfFkGL7_0),.clk(gclk));
	jdff dff_A_2P6IX7Vy4_0(.dout(w_dff_A_rSSfFkGL7_0),.din(w_dff_A_2P6IX7Vy4_0),.clk(gclk));
	jdff dff_A_jZ0Pp9hB4_0(.dout(w_dff_A_2P6IX7Vy4_0),.din(w_dff_A_jZ0Pp9hB4_0),.clk(gclk));
	jdff dff_A_FuL9DUHR5_0(.dout(w_dff_A_jZ0Pp9hB4_0),.din(w_dff_A_FuL9DUHR5_0),.clk(gclk));
	jdff dff_A_nFAIsQCq7_0(.dout(w_dff_A_FuL9DUHR5_0),.din(w_dff_A_nFAIsQCq7_0),.clk(gclk));
	jdff dff_A_gcJcQK3r4_0(.dout(w_dff_A_nFAIsQCq7_0),.din(w_dff_A_gcJcQK3r4_0),.clk(gclk));
	jdff dff_A_eUkOJ6RB7_0(.dout(w_dff_A_gcJcQK3r4_0),.din(w_dff_A_eUkOJ6RB7_0),.clk(gclk));
	jdff dff_A_Bzw9U4m02_0(.dout(w_dff_A_eUkOJ6RB7_0),.din(w_dff_A_Bzw9U4m02_0),.clk(gclk));
	jdff dff_A_mf73h0d85_0(.dout(w_dff_A_Bzw9U4m02_0),.din(w_dff_A_mf73h0d85_0),.clk(gclk));
	jdff dff_A_OhHNfjlm2_0(.dout(w_dff_A_mf73h0d85_0),.din(w_dff_A_OhHNfjlm2_0),.clk(gclk));
	jdff dff_A_B2Fb4YMo2_0(.dout(w_dff_A_OhHNfjlm2_0),.din(w_dff_A_B2Fb4YMo2_0),.clk(gclk));
	jdff dff_A_u6twTcmm9_0(.dout(w_dff_A_B2Fb4YMo2_0),.din(w_dff_A_u6twTcmm9_0),.clk(gclk));
	jdff dff_A_wAzQ8J249_0(.dout(w_dff_A_u6twTcmm9_0),.din(w_dff_A_wAzQ8J249_0),.clk(gclk));
	jdff dff_A_apdojfAh8_0(.dout(w_dff_A_wAzQ8J249_0),.din(w_dff_A_apdojfAh8_0),.clk(gclk));
	jdff dff_A_VGhAByjY6_0(.dout(w_dff_A_apdojfAh8_0),.din(w_dff_A_VGhAByjY6_0),.clk(gclk));
	jdff dff_A_VM7tfSf83_0(.dout(w_dff_A_VGhAByjY6_0),.din(w_dff_A_VM7tfSf83_0),.clk(gclk));
	jdff dff_A_J7xDq3NS9_0(.dout(w_dff_A_VM7tfSf83_0),.din(w_dff_A_J7xDq3NS9_0),.clk(gclk));
	jdff dff_A_GMkWIvKo6_0(.dout(w_dff_A_J7xDq3NS9_0),.din(w_dff_A_GMkWIvKo6_0),.clk(gclk));
	jdff dff_A_plhgGVHr5_0(.dout(w_dff_A_GMkWIvKo6_0),.din(w_dff_A_plhgGVHr5_0),.clk(gclk));
	jdff dff_A_PXn4uhnT1_0(.dout(w_dff_A_plhgGVHr5_0),.din(w_dff_A_PXn4uhnT1_0),.clk(gclk));
	jdff dff_A_tBZUMiHN1_0(.dout(w_dff_A_PXn4uhnT1_0),.din(w_dff_A_tBZUMiHN1_0),.clk(gclk));
	jdff dff_A_16NOPfRQ9_0(.dout(w_dff_A_tBZUMiHN1_0),.din(w_dff_A_16NOPfRQ9_0),.clk(gclk));
	jdff dff_A_zmfxMyyQ8_0(.dout(w_dff_A_16NOPfRQ9_0),.din(w_dff_A_zmfxMyyQ8_0),.clk(gclk));
	jdff dff_A_CNh7Nu3u2_0(.dout(w_dff_A_zmfxMyyQ8_0),.din(w_dff_A_CNh7Nu3u2_0),.clk(gclk));
	jdff dff_A_gtpigkUz9_0(.dout(w_dff_A_CNh7Nu3u2_0),.din(w_dff_A_gtpigkUz9_0),.clk(gclk));
	jdff dff_A_ymql107S1_0(.dout(w_dff_A_gtpigkUz9_0),.din(w_dff_A_ymql107S1_0),.clk(gclk));
	jdff dff_A_14eYYD6s0_0(.dout(w_n465_0[0]),.din(w_dff_A_14eYYD6s0_0),.clk(gclk));
	jdff dff_B_kPMvTxiM2_1(.din(n407),.dout(w_dff_B_kPMvTxiM2_1),.clk(gclk));
	jdff dff_A_YeJVYQXg0_0(.dout(w_n341_0[0]),.din(w_dff_A_YeJVYQXg0_0),.clk(gclk));
	jdff dff_A_R38Uz8Qr5_0(.dout(w_dff_A_YeJVYQXg0_0),.din(w_dff_A_R38Uz8Qr5_0),.clk(gclk));
	jdff dff_A_YeDyhrtn7_0(.dout(w_dff_A_R38Uz8Qr5_0),.din(w_dff_A_YeDyhrtn7_0),.clk(gclk));
	jdff dff_A_JRTqZJJi4_0(.dout(w_dff_A_YeDyhrtn7_0),.din(w_dff_A_JRTqZJJi4_0),.clk(gclk));
	jdff dff_A_GppyQCC35_0(.dout(w_dff_A_JRTqZJJi4_0),.din(w_dff_A_GppyQCC35_0),.clk(gclk));
	jdff dff_A_ZVfjUG6W6_0(.dout(w_dff_A_GppyQCC35_0),.din(w_dff_A_ZVfjUG6W6_0),.clk(gclk));
	jdff dff_A_HUEjaspn9_0(.dout(w_dff_A_ZVfjUG6W6_0),.din(w_dff_A_HUEjaspn9_0),.clk(gclk));
	jdff dff_A_Eycn70NM7_0(.dout(w_dff_A_HUEjaspn9_0),.din(w_dff_A_Eycn70NM7_0),.clk(gclk));
	jdff dff_A_1dG69cYp3_0(.dout(w_dff_A_Eycn70NM7_0),.din(w_dff_A_1dG69cYp3_0),.clk(gclk));
	jdff dff_A_LEBvhOVo8_0(.dout(w_dff_A_1dG69cYp3_0),.din(w_dff_A_LEBvhOVo8_0),.clk(gclk));
	jdff dff_A_um5d6ucm7_0(.dout(w_dff_A_LEBvhOVo8_0),.din(w_dff_A_um5d6ucm7_0),.clk(gclk));
	jdff dff_A_yDEYgugP7_0(.dout(w_dff_A_um5d6ucm7_0),.din(w_dff_A_yDEYgugP7_0),.clk(gclk));
	jdff dff_A_fFN5noq34_0(.dout(w_dff_A_yDEYgugP7_0),.din(w_dff_A_fFN5noq34_0),.clk(gclk));
	jdff dff_A_th0X1hPA4_0(.dout(w_dff_A_fFN5noq34_0),.din(w_dff_A_th0X1hPA4_0),.clk(gclk));
	jdff dff_A_xENboy8f2_0(.dout(w_dff_A_th0X1hPA4_0),.din(w_dff_A_xENboy8f2_0),.clk(gclk));
	jdff dff_A_uP4UVEoX6_0(.dout(w_dff_A_xENboy8f2_0),.din(w_dff_A_uP4UVEoX6_0),.clk(gclk));
	jdff dff_A_SdN53j033_0(.dout(w_dff_A_uP4UVEoX6_0),.din(w_dff_A_SdN53j033_0),.clk(gclk));
	jdff dff_A_uud2UxEa9_0(.dout(w_dff_A_SdN53j033_0),.din(w_dff_A_uud2UxEa9_0),.clk(gclk));
	jdff dff_A_6rdpdBqO0_0(.dout(w_dff_A_uud2UxEa9_0),.din(w_dff_A_6rdpdBqO0_0),.clk(gclk));
	jdff dff_A_AFdo8ZFi4_0(.dout(w_dff_A_6rdpdBqO0_0),.din(w_dff_A_AFdo8ZFi4_0),.clk(gclk));
	jdff dff_A_arRcaiPL9_0(.dout(w_dff_A_AFdo8ZFi4_0),.din(w_dff_A_arRcaiPL9_0),.clk(gclk));
	jdff dff_A_wNODA5kc9_0(.dout(w_dff_A_arRcaiPL9_0),.din(w_dff_A_wNODA5kc9_0),.clk(gclk));
	jdff dff_A_4O2bYNf23_0(.dout(w_dff_A_wNODA5kc9_0),.din(w_dff_A_4O2bYNf23_0),.clk(gclk));
	jdff dff_A_f6dTGFVx1_0(.dout(w_n393_0[0]),.din(w_dff_A_f6dTGFVx1_0),.clk(gclk));
	jdff dff_B_fe1ABSNx2_1(.din(n343),.dout(w_dff_B_fe1ABSNx2_1),.clk(gclk));
	jdff dff_A_v4h6FCT37_0(.dout(w_n283_0[0]),.din(w_dff_A_v4h6FCT37_0),.clk(gclk));
	jdff dff_A_xurBvHRF2_0(.dout(w_dff_A_v4h6FCT37_0),.din(w_dff_A_xurBvHRF2_0),.clk(gclk));
	jdff dff_A_thaJ0oX79_0(.dout(w_dff_A_xurBvHRF2_0),.din(w_dff_A_thaJ0oX79_0),.clk(gclk));
	jdff dff_A_3J2MmRBC0_0(.dout(w_dff_A_thaJ0oX79_0),.din(w_dff_A_3J2MmRBC0_0),.clk(gclk));
	jdff dff_A_EoRG3Vju7_0(.dout(w_dff_A_3J2MmRBC0_0),.din(w_dff_A_EoRG3Vju7_0),.clk(gclk));
	jdff dff_A_fPKf6J8R7_0(.dout(w_dff_A_EoRG3Vju7_0),.din(w_dff_A_fPKf6J8R7_0),.clk(gclk));
	jdff dff_A_HfWU2cp27_0(.dout(w_dff_A_fPKf6J8R7_0),.din(w_dff_A_HfWU2cp27_0),.clk(gclk));
	jdff dff_A_S3sF77xW4_0(.dout(w_dff_A_HfWU2cp27_0),.din(w_dff_A_S3sF77xW4_0),.clk(gclk));
	jdff dff_A_qnzCvVW00_0(.dout(w_dff_A_S3sF77xW4_0),.din(w_dff_A_qnzCvVW00_0),.clk(gclk));
	jdff dff_A_Oo8rQiay1_0(.dout(w_dff_A_qnzCvVW00_0),.din(w_dff_A_Oo8rQiay1_0),.clk(gclk));
	jdff dff_A_aZ8uug2N0_0(.dout(w_dff_A_Oo8rQiay1_0),.din(w_dff_A_aZ8uug2N0_0),.clk(gclk));
	jdff dff_A_O9TNbANi8_0(.dout(w_dff_A_aZ8uug2N0_0),.din(w_dff_A_O9TNbANi8_0),.clk(gclk));
	jdff dff_A_UsrYieBD6_0(.dout(w_dff_A_O9TNbANi8_0),.din(w_dff_A_UsrYieBD6_0),.clk(gclk));
	jdff dff_A_LxWqcRCL8_0(.dout(w_dff_A_UsrYieBD6_0),.din(w_dff_A_LxWqcRCL8_0),.clk(gclk));
	jdff dff_A_LhjZQx3V7_0(.dout(w_dff_A_LxWqcRCL8_0),.din(w_dff_A_LhjZQx3V7_0),.clk(gclk));
	jdff dff_A_xp19xgGk1_0(.dout(w_dff_A_LhjZQx3V7_0),.din(w_dff_A_xp19xgGk1_0),.clk(gclk));
	jdff dff_A_6wr8L5QS8_0(.dout(w_dff_A_xp19xgGk1_0),.din(w_dff_A_6wr8L5QS8_0),.clk(gclk));
	jdff dff_A_Il3ZipLs2_0(.dout(w_dff_A_6wr8L5QS8_0),.din(w_dff_A_Il3ZipLs2_0),.clk(gclk));
	jdff dff_A_W4SPQo6p9_0(.dout(w_dff_A_Il3ZipLs2_0),.din(w_dff_A_W4SPQo6p9_0),.clk(gclk));
	jdff dff_A_fWFkXRlH4_0(.dout(w_dff_A_W4SPQo6p9_0),.din(w_dff_A_fWFkXRlH4_0),.clk(gclk));
	jdff dff_A_QRKEAwBf9_0(.dout(w_n329_0[0]),.din(w_dff_A_QRKEAwBf9_0),.clk(gclk));
	jdff dff_B_O8JHUWz01_1(.din(n285),.dout(w_dff_B_O8JHUWz01_1),.clk(gclk));
	jdff dff_A_9POCDiGY1_0(.dout(w_n232_0[0]),.din(w_dff_A_9POCDiGY1_0),.clk(gclk));
	jdff dff_A_ZCHKqSSI1_0(.dout(w_dff_A_9POCDiGY1_0),.din(w_dff_A_ZCHKqSSI1_0),.clk(gclk));
	jdff dff_A_0S0TpdwX1_0(.dout(w_dff_A_ZCHKqSSI1_0),.din(w_dff_A_0S0TpdwX1_0),.clk(gclk));
	jdff dff_A_Mdz7uxmj4_0(.dout(w_dff_A_0S0TpdwX1_0),.din(w_dff_A_Mdz7uxmj4_0),.clk(gclk));
	jdff dff_A_I4W6y1b86_0(.dout(w_dff_A_Mdz7uxmj4_0),.din(w_dff_A_I4W6y1b86_0),.clk(gclk));
	jdff dff_A_w9YcuNlA4_0(.dout(w_dff_A_I4W6y1b86_0),.din(w_dff_A_w9YcuNlA4_0),.clk(gclk));
	jdff dff_A_4Yyi2UMC7_0(.dout(w_dff_A_w9YcuNlA4_0),.din(w_dff_A_4Yyi2UMC7_0),.clk(gclk));
	jdff dff_A_m6OJCe4J6_0(.dout(w_dff_A_4Yyi2UMC7_0),.din(w_dff_A_m6OJCe4J6_0),.clk(gclk));
	jdff dff_A_T10kneES8_0(.dout(w_dff_A_m6OJCe4J6_0),.din(w_dff_A_T10kneES8_0),.clk(gclk));
	jdff dff_A_LY7tWZne4_0(.dout(w_dff_A_T10kneES8_0),.din(w_dff_A_LY7tWZne4_0),.clk(gclk));
	jdff dff_A_ixXQUpog3_0(.dout(w_dff_A_LY7tWZne4_0),.din(w_dff_A_ixXQUpog3_0),.clk(gclk));
	jdff dff_A_JesL3Qq71_0(.dout(w_dff_A_ixXQUpog3_0),.din(w_dff_A_JesL3Qq71_0),.clk(gclk));
	jdff dff_A_RwR5CIS09_0(.dout(w_dff_A_JesL3Qq71_0),.din(w_dff_A_RwR5CIS09_0),.clk(gclk));
	jdff dff_A_awMZdQbR4_0(.dout(w_dff_A_RwR5CIS09_0),.din(w_dff_A_awMZdQbR4_0),.clk(gclk));
	jdff dff_A_wdugtVvB2_0(.dout(w_dff_A_awMZdQbR4_0),.din(w_dff_A_wdugtVvB2_0),.clk(gclk));
	jdff dff_A_4J1mDx4A8_0(.dout(w_dff_A_wdugtVvB2_0),.din(w_dff_A_4J1mDx4A8_0),.clk(gclk));
	jdff dff_A_9rl5Eyhd7_0(.dout(w_dff_A_4J1mDx4A8_0),.din(w_dff_A_9rl5Eyhd7_0),.clk(gclk));
	jdff dff_A_MysAQcee9_0(.dout(w_n271_0[0]),.din(w_dff_A_MysAQcee9_0),.clk(gclk));
	jdff dff_B_cbtQ91dg3_1(.din(n234),.dout(w_dff_B_cbtQ91dg3_1),.clk(gclk));
	jdff dff_A_4IDSjOmg1_0(.dout(w_n189_0[0]),.din(w_dff_A_4IDSjOmg1_0),.clk(gclk));
	jdff dff_A_yeXiaizK6_0(.dout(w_dff_A_4IDSjOmg1_0),.din(w_dff_A_yeXiaizK6_0),.clk(gclk));
	jdff dff_A_BRa5oHz15_0(.dout(w_dff_A_yeXiaizK6_0),.din(w_dff_A_BRa5oHz15_0),.clk(gclk));
	jdff dff_A_8A3KkQU06_0(.dout(w_dff_A_BRa5oHz15_0),.din(w_dff_A_8A3KkQU06_0),.clk(gclk));
	jdff dff_A_dKFWCrB36_0(.dout(w_dff_A_8A3KkQU06_0),.din(w_dff_A_dKFWCrB36_0),.clk(gclk));
	jdff dff_A_GbwxdbAl8_0(.dout(w_dff_A_dKFWCrB36_0),.din(w_dff_A_GbwxdbAl8_0),.clk(gclk));
	jdff dff_A_wxEnhyk05_0(.dout(w_dff_A_GbwxdbAl8_0),.din(w_dff_A_wxEnhyk05_0),.clk(gclk));
	jdff dff_A_SxUNq4le0_0(.dout(w_dff_A_wxEnhyk05_0),.din(w_dff_A_SxUNq4le0_0),.clk(gclk));
	jdff dff_A_vx89NLt18_0(.dout(w_dff_A_SxUNq4le0_0),.din(w_dff_A_vx89NLt18_0),.clk(gclk));
	jdff dff_A_TS2dk8aB6_0(.dout(w_dff_A_vx89NLt18_0),.din(w_dff_A_TS2dk8aB6_0),.clk(gclk));
	jdff dff_A_Ft1061mu7_0(.dout(w_dff_A_TS2dk8aB6_0),.din(w_dff_A_Ft1061mu7_0),.clk(gclk));
	jdff dff_A_CO63azFW2_0(.dout(w_dff_A_Ft1061mu7_0),.din(w_dff_A_CO63azFW2_0),.clk(gclk));
	jdff dff_A_sbQXxpaQ1_0(.dout(w_dff_A_CO63azFW2_0),.din(w_dff_A_sbQXxpaQ1_0),.clk(gclk));
	jdff dff_A_4hwEkcxO6_0(.dout(w_dff_A_sbQXxpaQ1_0),.din(w_dff_A_4hwEkcxO6_0),.clk(gclk));
	jdff dff_A_UvMWN99Q9_0(.dout(w_n220_0[0]),.din(w_dff_A_UvMWN99Q9_0),.clk(gclk));
	jdff dff_B_eeFZZLUH4_1(.din(n191),.dout(w_dff_B_eeFZZLUH4_1),.clk(gclk));
	jdff dff_A_dkxWOv9F3_0(.dout(w_n151_0[0]),.din(w_dff_A_dkxWOv9F3_0),.clk(gclk));
	jdff dff_A_2T6ae3xM2_0(.dout(w_dff_A_dkxWOv9F3_0),.din(w_dff_A_2T6ae3xM2_0),.clk(gclk));
	jdff dff_A_ma8HyiPD1_0(.dout(w_dff_A_2T6ae3xM2_0),.din(w_dff_A_ma8HyiPD1_0),.clk(gclk));
	jdff dff_A_U2wuna6b7_0(.dout(w_dff_A_ma8HyiPD1_0),.din(w_dff_A_U2wuna6b7_0),.clk(gclk));
	jdff dff_A_UpQ6p02F9_0(.dout(w_dff_A_U2wuna6b7_0),.din(w_dff_A_UpQ6p02F9_0),.clk(gclk));
	jdff dff_A_deECsCTN8_0(.dout(w_dff_A_UpQ6p02F9_0),.din(w_dff_A_deECsCTN8_0),.clk(gclk));
	jdff dff_A_SK85NqZm4_0(.dout(w_dff_A_deECsCTN8_0),.din(w_dff_A_SK85NqZm4_0),.clk(gclk));
	jdff dff_A_yIvN9eRV9_0(.dout(w_dff_A_SK85NqZm4_0),.din(w_dff_A_yIvN9eRV9_0),.clk(gclk));
	jdff dff_A_ibvQb0Gk5_0(.dout(w_dff_A_yIvN9eRV9_0),.din(w_dff_A_ibvQb0Gk5_0),.clk(gclk));
	jdff dff_A_LjPZjcXj8_0(.dout(w_dff_A_ibvQb0Gk5_0),.din(w_dff_A_LjPZjcXj8_0),.clk(gclk));
	jdff dff_A_HWEN1MZi5_0(.dout(w_dff_A_LjPZjcXj8_0),.din(w_dff_A_HWEN1MZi5_0),.clk(gclk));
	jdff dff_A_AQPO0Rr33_0(.dout(w_n177_0[0]),.din(w_dff_A_AQPO0Rr33_0),.clk(gclk));
	jdff dff_B_1ANJNn590_1(.din(n153),.dout(w_dff_B_1ANJNn590_1),.clk(gclk));
	jdff dff_A_zrNSo0n93_0(.dout(w_n116_0[0]),.din(w_dff_A_zrNSo0n93_0),.clk(gclk));
	jdff dff_A_lOpvbmHH4_0(.dout(w_dff_A_zrNSo0n93_0),.din(w_dff_A_lOpvbmHH4_0),.clk(gclk));
	jdff dff_A_AntLwJ2t4_0(.dout(w_dff_A_lOpvbmHH4_0),.din(w_dff_A_AntLwJ2t4_0),.clk(gclk));
	jdff dff_A_gk6giD027_0(.dout(w_dff_A_AntLwJ2t4_0),.din(w_dff_A_gk6giD027_0),.clk(gclk));
	jdff dff_A_sCloH9aA0_0(.dout(w_dff_A_gk6giD027_0),.din(w_dff_A_sCloH9aA0_0),.clk(gclk));
	jdff dff_A_IBKEFPBT2_0(.dout(w_dff_A_sCloH9aA0_0),.din(w_dff_A_IBKEFPBT2_0),.clk(gclk));
	jdff dff_A_7Xa03SXm3_0(.dout(w_dff_A_IBKEFPBT2_0),.din(w_dff_A_7Xa03SXm3_0),.clk(gclk));
	jdff dff_A_NiDcVqga0_0(.dout(w_dff_A_7Xa03SXm3_0),.din(w_dff_A_NiDcVqga0_0),.clk(gclk));
	jdff dff_A_SwFztyXO9_0(.dout(w_n139_0[0]),.din(w_dff_A_SwFztyXO9_0),.clk(gclk));
	jdff dff_A_tW1bCqem0_0(.dout(w_n104_0[0]),.din(w_dff_A_tW1bCqem0_0),.clk(gclk));
	jdff dff_A_MmWWRJ4h6_0(.dout(w_n85_0[0]),.din(w_dff_A_MmWWRJ4h6_0),.clk(gclk));
	jdff dff_A_latRsa6l4_1(.dout(w_n82_1[1]),.din(w_dff_A_latRsa6l4_1),.clk(gclk));
	jdff dff_A_tARccCuP3_0(.dout(w_n94_0[0]),.din(w_dff_A_tARccCuP3_0),.clk(gclk));
	jdff dff_A_2FdPF67W0_0(.dout(w_dff_A_tARccCuP3_0),.din(w_dff_A_2FdPF67W0_0),.clk(gclk));
	jdff dff_A_4pnYCnEO6_0(.dout(w_dff_A_2FdPF67W0_0),.din(w_dff_A_4pnYCnEO6_0),.clk(gclk));
	jdff dff_A_kb4H3JFE0_0(.dout(w_dff_A_4pnYCnEO6_0),.din(w_dff_A_kb4H3JFE0_0),.clk(gclk));
	jdff dff_A_GfrnQwgt6_0(.dout(w_dff_A_kb4H3JFE0_0),.din(w_dff_A_GfrnQwgt6_0),.clk(gclk));
	jdff dff_A_dAinsZSM4_0(.dout(w_n103_0[0]),.din(w_dff_A_dAinsZSM4_0),.clk(gclk));
	jdff dff_A_nDVYqqP91_0(.dout(w_dff_A_dAinsZSM4_0),.din(w_dff_A_nDVYqqP91_0),.clk(gclk));
	jdff dff_B_OcM2U1nk7_1(.din(n97),.dout(w_dff_B_OcM2U1nk7_1),.clk(gclk));
	jdff dff_A_balw0lKA6_1(.dout(w_n82_0[1]),.din(w_dff_A_balw0lKA6_1),.clk(gclk));
	jdff dff_A_z69XGoAz2_2(.dout(w_n82_0[2]),.din(w_dff_A_z69XGoAz2_2),.clk(gclk));
	jdff dff_A_jO2YVfKU2_2(.dout(w_dff_A_z69XGoAz2_2),.din(w_dff_A_jO2YVfKU2_2),.clk(gclk));
	jdff dff_A_NPQRlaQD6_0(.dout(w_n1151_0[0]),.din(w_dff_A_NPQRlaQD6_0),.clk(gclk));
	jdff dff_B_QGHX3ctl8_2(.din(n1151),.dout(w_dff_B_QGHX3ctl8_2),.clk(gclk));
	jdff dff_B_MHoeFrk23_2(.din(n1044),.dout(w_dff_B_MHoeFrk23_2),.clk(gclk));
	jdff dff_B_gws117dq8_2(.din(w_dff_B_MHoeFrk23_2),.dout(w_dff_B_gws117dq8_2),.clk(gclk));
	jdff dff_B_tifPlCMi5_2(.din(w_dff_B_gws117dq8_2),.dout(w_dff_B_tifPlCMi5_2),.clk(gclk));
	jdff dff_B_Rj64qouw7_2(.din(w_dff_B_tifPlCMi5_2),.dout(w_dff_B_Rj64qouw7_2),.clk(gclk));
	jdff dff_B_kQlaz3Tw8_2(.din(w_dff_B_Rj64qouw7_2),.dout(w_dff_B_kQlaz3Tw8_2),.clk(gclk));
	jdff dff_B_rRtv8xqQ1_2(.din(w_dff_B_kQlaz3Tw8_2),.dout(w_dff_B_rRtv8xqQ1_2),.clk(gclk));
	jdff dff_B_ey2UuyBs2_2(.din(w_dff_B_rRtv8xqQ1_2),.dout(w_dff_B_ey2UuyBs2_2),.clk(gclk));
	jdff dff_B_F0p8rIpF7_2(.din(w_dff_B_ey2UuyBs2_2),.dout(w_dff_B_F0p8rIpF7_2),.clk(gclk));
	jdff dff_B_Br6ydx2a0_2(.din(w_dff_B_F0p8rIpF7_2),.dout(w_dff_B_Br6ydx2a0_2),.clk(gclk));
	jdff dff_B_2zzmWZYw0_2(.din(w_dff_B_Br6ydx2a0_2),.dout(w_dff_B_2zzmWZYw0_2),.clk(gclk));
	jdff dff_B_vp6DkEgp1_2(.din(w_dff_B_2zzmWZYw0_2),.dout(w_dff_B_vp6DkEgp1_2),.clk(gclk));
	jdff dff_B_MDnTEYkg5_2(.din(w_dff_B_vp6DkEgp1_2),.dout(w_dff_B_MDnTEYkg5_2),.clk(gclk));
	jdff dff_B_F3di0N1X6_2(.din(w_dff_B_MDnTEYkg5_2),.dout(w_dff_B_F3di0N1X6_2),.clk(gclk));
	jdff dff_B_GAOlDm706_2(.din(w_dff_B_F3di0N1X6_2),.dout(w_dff_B_GAOlDm706_2),.clk(gclk));
	jdff dff_B_7jCxRxhH3_2(.din(w_dff_B_GAOlDm706_2),.dout(w_dff_B_7jCxRxhH3_2),.clk(gclk));
	jdff dff_B_ifmk5Njb2_2(.din(w_dff_B_7jCxRxhH3_2),.dout(w_dff_B_ifmk5Njb2_2),.clk(gclk));
	jdff dff_B_aIOg3fAo8_2(.din(w_dff_B_ifmk5Njb2_2),.dout(w_dff_B_aIOg3fAo8_2),.clk(gclk));
	jdff dff_B_0ATg7qQP5_2(.din(w_dff_B_aIOg3fAo8_2),.dout(w_dff_B_0ATg7qQP5_2),.clk(gclk));
	jdff dff_B_7H3zKe8G2_2(.din(w_dff_B_0ATg7qQP5_2),.dout(w_dff_B_7H3zKe8G2_2),.clk(gclk));
	jdff dff_B_k910qDAn8_2(.din(w_dff_B_7H3zKe8G2_2),.dout(w_dff_B_k910qDAn8_2),.clk(gclk));
	jdff dff_B_Xxr9HxW06_2(.din(w_dff_B_k910qDAn8_2),.dout(w_dff_B_Xxr9HxW06_2),.clk(gclk));
	jdff dff_B_wOXhzEnW7_2(.din(w_dff_B_Xxr9HxW06_2),.dout(w_dff_B_wOXhzEnW7_2),.clk(gclk));
	jdff dff_B_d1jkG5A91_2(.din(w_dff_B_wOXhzEnW7_2),.dout(w_dff_B_d1jkG5A91_2),.clk(gclk));
	jdff dff_B_Zvy5EmfT8_2(.din(w_dff_B_d1jkG5A91_2),.dout(w_dff_B_Zvy5EmfT8_2),.clk(gclk));
	jdff dff_B_M7Dc5XBP8_2(.din(w_dff_B_Zvy5EmfT8_2),.dout(w_dff_B_M7Dc5XBP8_2),.clk(gclk));
	jdff dff_B_18qI0mSA0_2(.din(w_dff_B_M7Dc5XBP8_2),.dout(w_dff_B_18qI0mSA0_2),.clk(gclk));
	jdff dff_B_uUHLfI278_2(.din(w_dff_B_18qI0mSA0_2),.dout(w_dff_B_uUHLfI278_2),.clk(gclk));
	jdff dff_B_idxkNm928_2(.din(w_dff_B_uUHLfI278_2),.dout(w_dff_B_idxkNm928_2),.clk(gclk));
	jdff dff_B_icSfbRwi4_2(.din(w_dff_B_idxkNm928_2),.dout(w_dff_B_icSfbRwi4_2),.clk(gclk));
	jdff dff_B_LcGvbYJG9_2(.din(w_dff_B_icSfbRwi4_2),.dout(w_dff_B_LcGvbYJG9_2),.clk(gclk));
	jdff dff_B_RupLQkck6_2(.din(w_dff_B_LcGvbYJG9_2),.dout(w_dff_B_RupLQkck6_2),.clk(gclk));
	jdff dff_B_SqA6HFO79_2(.din(w_dff_B_RupLQkck6_2),.dout(w_dff_B_SqA6HFO79_2),.clk(gclk));
	jdff dff_B_8ZUQ4tkS4_2(.din(w_dff_B_SqA6HFO79_2),.dout(w_dff_B_8ZUQ4tkS4_2),.clk(gclk));
	jdff dff_B_ag5IAlUv0_2(.din(w_dff_B_8ZUQ4tkS4_2),.dout(w_dff_B_ag5IAlUv0_2),.clk(gclk));
	jdff dff_B_PNcUOeWy6_2(.din(w_dff_B_ag5IAlUv0_2),.dout(w_dff_B_PNcUOeWy6_2),.clk(gclk));
	jdff dff_B_FY9qpg459_2(.din(w_dff_B_PNcUOeWy6_2),.dout(w_dff_B_FY9qpg459_2),.clk(gclk));
	jdff dff_B_OeklvmLV9_2(.din(w_dff_B_FY9qpg459_2),.dout(w_dff_B_OeklvmLV9_2),.clk(gclk));
	jdff dff_B_XWAljari1_2(.din(w_dff_B_OeklvmLV9_2),.dout(w_dff_B_XWAljari1_2),.clk(gclk));
	jdff dff_B_iJHGWhC59_2(.din(w_dff_B_XWAljari1_2),.dout(w_dff_B_iJHGWhC59_2),.clk(gclk));
	jdff dff_B_Qrjc45HK0_2(.din(w_dff_B_iJHGWhC59_2),.dout(w_dff_B_Qrjc45HK0_2),.clk(gclk));
	jdff dff_B_RrNwMvPl4_2(.din(w_dff_B_Qrjc45HK0_2),.dout(w_dff_B_RrNwMvPl4_2),.clk(gclk));
	jdff dff_B_ObwdBbpI9_2(.din(w_dff_B_RrNwMvPl4_2),.dout(w_dff_B_ObwdBbpI9_2),.clk(gclk));
	jdff dff_B_V7ssezCX9_2(.din(w_dff_B_ObwdBbpI9_2),.dout(w_dff_B_V7ssezCX9_2),.clk(gclk));
	jdff dff_B_RMjRo5a85_2(.din(w_dff_B_V7ssezCX9_2),.dout(w_dff_B_RMjRo5a85_2),.clk(gclk));
	jdff dff_A_Gr7HxICE1_0(.dout(w_n1048_0[0]),.din(w_dff_A_Gr7HxICE1_0),.clk(gclk));
	jdff dff_B_C5C6vHsw0_1(.din(n1046),.dout(w_dff_B_C5C6vHsw0_1),.clk(gclk));
	jdff dff_B_iaZRAhFW6_2(.din(n943),.dout(w_dff_B_iaZRAhFW6_2),.clk(gclk));
	jdff dff_B_2TDY65Zz8_2(.din(w_dff_B_iaZRAhFW6_2),.dout(w_dff_B_2TDY65Zz8_2),.clk(gclk));
	jdff dff_B_0fhOpMHw5_2(.din(w_dff_B_2TDY65Zz8_2),.dout(w_dff_B_0fhOpMHw5_2),.clk(gclk));
	jdff dff_B_vvzU0n9K2_2(.din(w_dff_B_0fhOpMHw5_2),.dout(w_dff_B_vvzU0n9K2_2),.clk(gclk));
	jdff dff_B_10vFc8aT8_2(.din(w_dff_B_vvzU0n9K2_2),.dout(w_dff_B_10vFc8aT8_2),.clk(gclk));
	jdff dff_B_SMvp4JlQ5_2(.din(w_dff_B_10vFc8aT8_2),.dout(w_dff_B_SMvp4JlQ5_2),.clk(gclk));
	jdff dff_B_tP7UwAxs3_2(.din(w_dff_B_SMvp4JlQ5_2),.dout(w_dff_B_tP7UwAxs3_2),.clk(gclk));
	jdff dff_B_JfNg4S6k6_2(.din(w_dff_B_tP7UwAxs3_2),.dout(w_dff_B_JfNg4S6k6_2),.clk(gclk));
	jdff dff_B_bYrUj9De7_2(.din(w_dff_B_JfNg4S6k6_2),.dout(w_dff_B_bYrUj9De7_2),.clk(gclk));
	jdff dff_B_Cgosjsxv6_2(.din(w_dff_B_bYrUj9De7_2),.dout(w_dff_B_Cgosjsxv6_2),.clk(gclk));
	jdff dff_B_Aml9V9434_2(.din(w_dff_B_Cgosjsxv6_2),.dout(w_dff_B_Aml9V9434_2),.clk(gclk));
	jdff dff_B_a7R85p2m3_2(.din(w_dff_B_Aml9V9434_2),.dout(w_dff_B_a7R85p2m3_2),.clk(gclk));
	jdff dff_B_5xuTbzze6_2(.din(w_dff_B_a7R85p2m3_2),.dout(w_dff_B_5xuTbzze6_2),.clk(gclk));
	jdff dff_B_V0r0Cty86_2(.din(w_dff_B_5xuTbzze6_2),.dout(w_dff_B_V0r0Cty86_2),.clk(gclk));
	jdff dff_B_wbkapKat3_2(.din(w_dff_B_V0r0Cty86_2),.dout(w_dff_B_wbkapKat3_2),.clk(gclk));
	jdff dff_B_X0QoIk4I0_2(.din(w_dff_B_wbkapKat3_2),.dout(w_dff_B_X0QoIk4I0_2),.clk(gclk));
	jdff dff_B_ika6nGXW6_2(.din(w_dff_B_X0QoIk4I0_2),.dout(w_dff_B_ika6nGXW6_2),.clk(gclk));
	jdff dff_B_wyaMoXPG7_2(.din(w_dff_B_ika6nGXW6_2),.dout(w_dff_B_wyaMoXPG7_2),.clk(gclk));
	jdff dff_B_JNFVLx476_2(.din(w_dff_B_wyaMoXPG7_2),.dout(w_dff_B_JNFVLx476_2),.clk(gclk));
	jdff dff_B_x6WgiwO93_2(.din(w_dff_B_JNFVLx476_2),.dout(w_dff_B_x6WgiwO93_2),.clk(gclk));
	jdff dff_B_JMVRf94X0_2(.din(w_dff_B_x6WgiwO93_2),.dout(w_dff_B_JMVRf94X0_2),.clk(gclk));
	jdff dff_B_BoPQ9V3g4_2(.din(w_dff_B_JMVRf94X0_2),.dout(w_dff_B_BoPQ9V3g4_2),.clk(gclk));
	jdff dff_B_ZYOlnaYm7_2(.din(w_dff_B_BoPQ9V3g4_2),.dout(w_dff_B_ZYOlnaYm7_2),.clk(gclk));
	jdff dff_B_4jhnZ5ka0_2(.din(w_dff_B_ZYOlnaYm7_2),.dout(w_dff_B_4jhnZ5ka0_2),.clk(gclk));
	jdff dff_B_eIRitcNo3_2(.din(w_dff_B_4jhnZ5ka0_2),.dout(w_dff_B_eIRitcNo3_2),.clk(gclk));
	jdff dff_B_TvqE9uf95_2(.din(w_dff_B_eIRitcNo3_2),.dout(w_dff_B_TvqE9uf95_2),.clk(gclk));
	jdff dff_B_3bKDlMsj1_2(.din(w_dff_B_TvqE9uf95_2),.dout(w_dff_B_3bKDlMsj1_2),.clk(gclk));
	jdff dff_B_DcS1Cs1W5_2(.din(w_dff_B_3bKDlMsj1_2),.dout(w_dff_B_DcS1Cs1W5_2),.clk(gclk));
	jdff dff_B_fonBbvhv6_2(.din(w_dff_B_DcS1Cs1W5_2),.dout(w_dff_B_fonBbvhv6_2),.clk(gclk));
	jdff dff_B_y1KNow2p2_2(.din(w_dff_B_fonBbvhv6_2),.dout(w_dff_B_y1KNow2p2_2),.clk(gclk));
	jdff dff_B_BIs2VB3x1_2(.din(w_dff_B_y1KNow2p2_2),.dout(w_dff_B_BIs2VB3x1_2),.clk(gclk));
	jdff dff_B_Czt5w7if6_2(.din(w_dff_B_BIs2VB3x1_2),.dout(w_dff_B_Czt5w7if6_2),.clk(gclk));
	jdff dff_B_9GKbfECR6_2(.din(w_dff_B_Czt5w7if6_2),.dout(w_dff_B_9GKbfECR6_2),.clk(gclk));
	jdff dff_B_0VfGIVGN6_2(.din(w_dff_B_9GKbfECR6_2),.dout(w_dff_B_0VfGIVGN6_2),.clk(gclk));
	jdff dff_B_0bHdgDPC4_2(.din(w_dff_B_0VfGIVGN6_2),.dout(w_dff_B_0bHdgDPC4_2),.clk(gclk));
	jdff dff_B_spyQcbM83_2(.din(w_dff_B_0bHdgDPC4_2),.dout(w_dff_B_spyQcbM83_2),.clk(gclk));
	jdff dff_B_QJYOa0LS2_2(.din(w_dff_B_spyQcbM83_2),.dout(w_dff_B_QJYOa0LS2_2),.clk(gclk));
	jdff dff_B_CF9HbN4S9_2(.din(w_dff_B_QJYOa0LS2_2),.dout(w_dff_B_CF9HbN4S9_2),.clk(gclk));
	jdff dff_B_cPZGtjOu4_2(.din(w_dff_B_CF9HbN4S9_2),.dout(w_dff_B_cPZGtjOu4_2),.clk(gclk));
	jdff dff_B_IJd8LxC51_2(.din(w_dff_B_cPZGtjOu4_2),.dout(w_dff_B_IJd8LxC51_2),.clk(gclk));
	jdff dff_B_YoBgo9Qz8_2(.din(w_dff_B_IJd8LxC51_2),.dout(w_dff_B_YoBgo9Qz8_2),.clk(gclk));
	jdff dff_A_Voa2nWZi3_1(.dout(w_n1032_0[1]),.din(w_dff_A_Voa2nWZi3_1),.clk(gclk));
	jdff dff_A_wffRyLGQ2_0(.dout(w_n840_0[0]),.din(w_dff_A_wffRyLGQ2_0),.clk(gclk));
	jdff dff_A_Jiev30sR6_0(.dout(w_dff_A_wffRyLGQ2_0),.din(w_dff_A_Jiev30sR6_0),.clk(gclk));
	jdff dff_A_yRzzr99x9_0(.dout(w_dff_A_Jiev30sR6_0),.din(w_dff_A_yRzzr99x9_0),.clk(gclk));
	jdff dff_A_okwQI6dM4_0(.dout(w_dff_A_yRzzr99x9_0),.din(w_dff_A_okwQI6dM4_0),.clk(gclk));
	jdff dff_A_WlfA4e3J1_0(.dout(w_dff_A_okwQI6dM4_0),.din(w_dff_A_WlfA4e3J1_0),.clk(gclk));
	jdff dff_A_9izv6p7Q0_0(.dout(w_dff_A_WlfA4e3J1_0),.din(w_dff_A_9izv6p7Q0_0),.clk(gclk));
	jdff dff_A_oG2l49pI2_0(.dout(w_dff_A_9izv6p7Q0_0),.din(w_dff_A_oG2l49pI2_0),.clk(gclk));
	jdff dff_A_JrvRMgIl1_0(.dout(w_dff_A_oG2l49pI2_0),.din(w_dff_A_JrvRMgIl1_0),.clk(gclk));
	jdff dff_A_o6Cj6fUe2_0(.dout(w_dff_A_JrvRMgIl1_0),.din(w_dff_A_o6Cj6fUe2_0),.clk(gclk));
	jdff dff_A_AZb03TZg5_0(.dout(w_dff_A_o6Cj6fUe2_0),.din(w_dff_A_AZb03TZg5_0),.clk(gclk));
	jdff dff_A_AYp5yxnn5_0(.dout(w_dff_A_AZb03TZg5_0),.din(w_dff_A_AYp5yxnn5_0),.clk(gclk));
	jdff dff_A_M83VFdcT0_0(.dout(w_dff_A_AYp5yxnn5_0),.din(w_dff_A_M83VFdcT0_0),.clk(gclk));
	jdff dff_A_vgfgNsFQ8_0(.dout(w_dff_A_M83VFdcT0_0),.din(w_dff_A_vgfgNsFQ8_0),.clk(gclk));
	jdff dff_A_AbLuLFGa1_0(.dout(w_dff_A_vgfgNsFQ8_0),.din(w_dff_A_AbLuLFGa1_0),.clk(gclk));
	jdff dff_A_0enXMpnx4_0(.dout(w_dff_A_AbLuLFGa1_0),.din(w_dff_A_0enXMpnx4_0),.clk(gclk));
	jdff dff_A_2SNGlnfv3_0(.dout(w_dff_A_0enXMpnx4_0),.din(w_dff_A_2SNGlnfv3_0),.clk(gclk));
	jdff dff_A_DuIUZFrL8_0(.dout(w_dff_A_2SNGlnfv3_0),.din(w_dff_A_DuIUZFrL8_0),.clk(gclk));
	jdff dff_A_8fEtIe8F0_0(.dout(w_dff_A_DuIUZFrL8_0),.din(w_dff_A_8fEtIe8F0_0),.clk(gclk));
	jdff dff_A_NIK03Wgq9_0(.dout(w_dff_A_8fEtIe8F0_0),.din(w_dff_A_NIK03Wgq9_0),.clk(gclk));
	jdff dff_A_QjXnEzaT1_0(.dout(w_dff_A_NIK03Wgq9_0),.din(w_dff_A_QjXnEzaT1_0),.clk(gclk));
	jdff dff_A_bzEBMzYu8_0(.dout(w_dff_A_QjXnEzaT1_0),.din(w_dff_A_bzEBMzYu8_0),.clk(gclk));
	jdff dff_A_oa3qovs33_0(.dout(w_dff_A_bzEBMzYu8_0),.din(w_dff_A_oa3qovs33_0),.clk(gclk));
	jdff dff_A_j22LvmOX9_0(.dout(w_dff_A_oa3qovs33_0),.din(w_dff_A_j22LvmOX9_0),.clk(gclk));
	jdff dff_A_WO8fjwTM6_0(.dout(w_dff_A_j22LvmOX9_0),.din(w_dff_A_WO8fjwTM6_0),.clk(gclk));
	jdff dff_A_k4v5EosN3_0(.dout(w_dff_A_WO8fjwTM6_0),.din(w_dff_A_k4v5EosN3_0),.clk(gclk));
	jdff dff_A_bvLb5Hwb9_0(.dout(w_dff_A_k4v5EosN3_0),.din(w_dff_A_bvLb5Hwb9_0),.clk(gclk));
	jdff dff_A_gl2Xkir28_0(.dout(w_dff_A_bvLb5Hwb9_0),.din(w_dff_A_gl2Xkir28_0),.clk(gclk));
	jdff dff_A_cKB4c44g8_0(.dout(w_dff_A_gl2Xkir28_0),.din(w_dff_A_cKB4c44g8_0),.clk(gclk));
	jdff dff_A_fIXzMqHS5_0(.dout(w_dff_A_cKB4c44g8_0),.din(w_dff_A_fIXzMqHS5_0),.clk(gclk));
	jdff dff_A_DtHx8EY68_0(.dout(w_dff_A_fIXzMqHS5_0),.din(w_dff_A_DtHx8EY68_0),.clk(gclk));
	jdff dff_A_8PxlBvTy6_0(.dout(w_dff_A_DtHx8EY68_0),.din(w_dff_A_8PxlBvTy6_0),.clk(gclk));
	jdff dff_A_yC00dDdR2_0(.dout(w_dff_A_8PxlBvTy6_0),.din(w_dff_A_yC00dDdR2_0),.clk(gclk));
	jdff dff_A_DkrMaw6R4_0(.dout(w_dff_A_yC00dDdR2_0),.din(w_dff_A_DkrMaw6R4_0),.clk(gclk));
	jdff dff_A_PddTMFSd3_0(.dout(w_dff_A_DkrMaw6R4_0),.din(w_dff_A_PddTMFSd3_0),.clk(gclk));
	jdff dff_A_X1EWdI6e8_0(.dout(w_dff_A_PddTMFSd3_0),.din(w_dff_A_X1EWdI6e8_0),.clk(gclk));
	jdff dff_A_gEHaypot5_0(.dout(w_dff_A_X1EWdI6e8_0),.din(w_dff_A_gEHaypot5_0),.clk(gclk));
	jdff dff_A_aGBweFga6_0(.dout(w_dff_A_gEHaypot5_0),.din(w_dff_A_aGBweFga6_0),.clk(gclk));
	jdff dff_A_rddEyTe76_0(.dout(w_dff_A_aGBweFga6_0),.din(w_dff_A_rddEyTe76_0),.clk(gclk));
	jdff dff_A_wALpsxUl8_1(.dout(w_n927_0[1]),.din(w_dff_A_wALpsxUl8_1),.clk(gclk));
	jdff dff_A_9OrlJGK70_2(.dout(w_n927_0[2]),.din(w_dff_A_9OrlJGK70_2),.clk(gclk));
	jdff dff_B_fW2vjjGI2_1(.din(n842),.dout(w_dff_B_fW2vjjGI2_1),.clk(gclk));
	jdff dff_B_IJ5OlnYO2_2(.din(n742),.dout(w_dff_B_IJ5OlnYO2_2),.clk(gclk));
	jdff dff_B_8IgOr1vF2_2(.din(w_dff_B_IJ5OlnYO2_2),.dout(w_dff_B_8IgOr1vF2_2),.clk(gclk));
	jdff dff_B_rl6nwMBb7_2(.din(w_dff_B_8IgOr1vF2_2),.dout(w_dff_B_rl6nwMBb7_2),.clk(gclk));
	jdff dff_B_TStHV4gC1_2(.din(w_dff_B_rl6nwMBb7_2),.dout(w_dff_B_TStHV4gC1_2),.clk(gclk));
	jdff dff_B_VS3KmYDs1_2(.din(w_dff_B_TStHV4gC1_2),.dout(w_dff_B_VS3KmYDs1_2),.clk(gclk));
	jdff dff_B_RDOWJLpY9_2(.din(w_dff_B_VS3KmYDs1_2),.dout(w_dff_B_RDOWJLpY9_2),.clk(gclk));
	jdff dff_B_F4WPU77a4_2(.din(w_dff_B_RDOWJLpY9_2),.dout(w_dff_B_F4WPU77a4_2),.clk(gclk));
	jdff dff_B_MsPTZtWX0_2(.din(w_dff_B_F4WPU77a4_2),.dout(w_dff_B_MsPTZtWX0_2),.clk(gclk));
	jdff dff_B_N7hLyVMd8_2(.din(w_dff_B_MsPTZtWX0_2),.dout(w_dff_B_N7hLyVMd8_2),.clk(gclk));
	jdff dff_B_UaRHLEQh0_2(.din(w_dff_B_N7hLyVMd8_2),.dout(w_dff_B_UaRHLEQh0_2),.clk(gclk));
	jdff dff_B_KKTM7mhX0_2(.din(w_dff_B_UaRHLEQh0_2),.dout(w_dff_B_KKTM7mhX0_2),.clk(gclk));
	jdff dff_B_eFNfMcul8_2(.din(w_dff_B_KKTM7mhX0_2),.dout(w_dff_B_eFNfMcul8_2),.clk(gclk));
	jdff dff_B_CGWKM9Es8_2(.din(w_dff_B_eFNfMcul8_2),.dout(w_dff_B_CGWKM9Es8_2),.clk(gclk));
	jdff dff_B_SKRDRi1s4_2(.din(w_dff_B_CGWKM9Es8_2),.dout(w_dff_B_SKRDRi1s4_2),.clk(gclk));
	jdff dff_B_gSelskiQ9_2(.din(w_dff_B_SKRDRi1s4_2),.dout(w_dff_B_gSelskiQ9_2),.clk(gclk));
	jdff dff_B_O39CEEfe2_2(.din(w_dff_B_gSelskiQ9_2),.dout(w_dff_B_O39CEEfe2_2),.clk(gclk));
	jdff dff_B_Hn0InsQg1_2(.din(w_dff_B_O39CEEfe2_2),.dout(w_dff_B_Hn0InsQg1_2),.clk(gclk));
	jdff dff_B_CE985Xd50_2(.din(w_dff_B_Hn0InsQg1_2),.dout(w_dff_B_CE985Xd50_2),.clk(gclk));
	jdff dff_B_GtU9kTDA0_2(.din(w_dff_B_CE985Xd50_2),.dout(w_dff_B_GtU9kTDA0_2),.clk(gclk));
	jdff dff_B_OB8Bx5xK2_2(.din(w_dff_B_GtU9kTDA0_2),.dout(w_dff_B_OB8Bx5xK2_2),.clk(gclk));
	jdff dff_B_GLYUIhhM4_2(.din(w_dff_B_OB8Bx5xK2_2),.dout(w_dff_B_GLYUIhhM4_2),.clk(gclk));
	jdff dff_B_kYmFj8NL4_2(.din(w_dff_B_GLYUIhhM4_2),.dout(w_dff_B_kYmFj8NL4_2),.clk(gclk));
	jdff dff_B_LatTYkkC1_2(.din(w_dff_B_kYmFj8NL4_2),.dout(w_dff_B_LatTYkkC1_2),.clk(gclk));
	jdff dff_B_dQMelPoN9_2(.din(w_dff_B_LatTYkkC1_2),.dout(w_dff_B_dQMelPoN9_2),.clk(gclk));
	jdff dff_B_RGqQmZMC8_2(.din(w_dff_B_dQMelPoN9_2),.dout(w_dff_B_RGqQmZMC8_2),.clk(gclk));
	jdff dff_B_oOjENsPs8_2(.din(w_dff_B_RGqQmZMC8_2),.dout(w_dff_B_oOjENsPs8_2),.clk(gclk));
	jdff dff_B_rkcCQZ1A9_2(.din(w_dff_B_oOjENsPs8_2),.dout(w_dff_B_rkcCQZ1A9_2),.clk(gclk));
	jdff dff_B_QOlkaEfQ8_2(.din(w_dff_B_rkcCQZ1A9_2),.dout(w_dff_B_QOlkaEfQ8_2),.clk(gclk));
	jdff dff_B_1IeHQctC1_2(.din(w_dff_B_QOlkaEfQ8_2),.dout(w_dff_B_1IeHQctC1_2),.clk(gclk));
	jdff dff_B_HeUSRud13_2(.din(w_dff_B_1IeHQctC1_2),.dout(w_dff_B_HeUSRud13_2),.clk(gclk));
	jdff dff_B_SaltxAMU0_2(.din(w_dff_B_HeUSRud13_2),.dout(w_dff_B_SaltxAMU0_2),.clk(gclk));
	jdff dff_B_9V9GPrAc5_2(.din(w_dff_B_SaltxAMU0_2),.dout(w_dff_B_9V9GPrAc5_2),.clk(gclk));
	jdff dff_B_YFh1Hbc80_2(.din(w_dff_B_9V9GPrAc5_2),.dout(w_dff_B_YFh1Hbc80_2),.clk(gclk));
	jdff dff_B_XHgoh4ZN7_2(.din(w_dff_B_YFh1Hbc80_2),.dout(w_dff_B_XHgoh4ZN7_2),.clk(gclk));
	jdff dff_B_xlzt7Jp13_2(.din(n821),.dout(w_dff_B_xlzt7Jp13_2),.clk(gclk));
	jdff dff_B_oSL6BcdO5_1(.din(n743),.dout(w_dff_B_oSL6BcdO5_1),.clk(gclk));
	jdff dff_B_iMdscc0W2_2(.din(n649),.dout(w_dff_B_iMdscc0W2_2),.clk(gclk));
	jdff dff_B_jFQW4TTe5_2(.din(w_dff_B_iMdscc0W2_2),.dout(w_dff_B_jFQW4TTe5_2),.clk(gclk));
	jdff dff_B_tGPVsApc9_2(.din(w_dff_B_jFQW4TTe5_2),.dout(w_dff_B_tGPVsApc9_2),.clk(gclk));
	jdff dff_B_pGsXkn8C9_2(.din(w_dff_B_tGPVsApc9_2),.dout(w_dff_B_pGsXkn8C9_2),.clk(gclk));
	jdff dff_B_057dNnmj0_2(.din(w_dff_B_pGsXkn8C9_2),.dout(w_dff_B_057dNnmj0_2),.clk(gclk));
	jdff dff_B_OY10Ofyj4_2(.din(w_dff_B_057dNnmj0_2),.dout(w_dff_B_OY10Ofyj4_2),.clk(gclk));
	jdff dff_B_rbpXlvB25_2(.din(w_dff_B_OY10Ofyj4_2),.dout(w_dff_B_rbpXlvB25_2),.clk(gclk));
	jdff dff_B_Bqq1RtNr1_2(.din(w_dff_B_rbpXlvB25_2),.dout(w_dff_B_Bqq1RtNr1_2),.clk(gclk));
	jdff dff_B_liNTPTn07_2(.din(w_dff_B_Bqq1RtNr1_2),.dout(w_dff_B_liNTPTn07_2),.clk(gclk));
	jdff dff_B_ZgOedF5v2_2(.din(w_dff_B_liNTPTn07_2),.dout(w_dff_B_ZgOedF5v2_2),.clk(gclk));
	jdff dff_B_UTHrbvr56_2(.din(w_dff_B_ZgOedF5v2_2),.dout(w_dff_B_UTHrbvr56_2),.clk(gclk));
	jdff dff_B_Z1kbUkjJ4_2(.din(w_dff_B_UTHrbvr56_2),.dout(w_dff_B_Z1kbUkjJ4_2),.clk(gclk));
	jdff dff_B_r2aTpHtA9_2(.din(w_dff_B_Z1kbUkjJ4_2),.dout(w_dff_B_r2aTpHtA9_2),.clk(gclk));
	jdff dff_B_TQBDAibS2_2(.din(w_dff_B_r2aTpHtA9_2),.dout(w_dff_B_TQBDAibS2_2),.clk(gclk));
	jdff dff_B_UFo8eQQv2_2(.din(w_dff_B_TQBDAibS2_2),.dout(w_dff_B_UFo8eQQv2_2),.clk(gclk));
	jdff dff_B_Zmc2OscO3_2(.din(w_dff_B_UFo8eQQv2_2),.dout(w_dff_B_Zmc2OscO3_2),.clk(gclk));
	jdff dff_B_QroViJCe0_2(.din(w_dff_B_Zmc2OscO3_2),.dout(w_dff_B_QroViJCe0_2),.clk(gclk));
	jdff dff_B_5vHej5g29_2(.din(w_dff_B_QroViJCe0_2),.dout(w_dff_B_5vHej5g29_2),.clk(gclk));
	jdff dff_B_balQTqqz3_2(.din(w_dff_B_5vHej5g29_2),.dout(w_dff_B_balQTqqz3_2),.clk(gclk));
	jdff dff_B_3sTWP1yL3_2(.din(w_dff_B_balQTqqz3_2),.dout(w_dff_B_3sTWP1yL3_2),.clk(gclk));
	jdff dff_B_YT72ouv26_2(.din(w_dff_B_3sTWP1yL3_2),.dout(w_dff_B_YT72ouv26_2),.clk(gclk));
	jdff dff_B_5ODYHuU70_2(.din(w_dff_B_YT72ouv26_2),.dout(w_dff_B_5ODYHuU70_2),.clk(gclk));
	jdff dff_B_BigxqMvF8_2(.din(w_dff_B_5ODYHuU70_2),.dout(w_dff_B_BigxqMvF8_2),.clk(gclk));
	jdff dff_B_AVo9YrBg9_2(.din(w_dff_B_BigxqMvF8_2),.dout(w_dff_B_AVo9YrBg9_2),.clk(gclk));
	jdff dff_B_GcNonWx66_2(.din(w_dff_B_AVo9YrBg9_2),.dout(w_dff_B_GcNonWx66_2),.clk(gclk));
	jdff dff_B_UKi28Gol0_2(.din(w_dff_B_GcNonWx66_2),.dout(w_dff_B_UKi28Gol0_2),.clk(gclk));
	jdff dff_B_zOMFcPxr4_2(.din(w_dff_B_UKi28Gol0_2),.dout(w_dff_B_zOMFcPxr4_2),.clk(gclk));
	jdff dff_B_bZJxbUq97_2(.din(w_dff_B_zOMFcPxr4_2),.dout(w_dff_B_bZJxbUq97_2),.clk(gclk));
	jdff dff_B_CVPIZxQW3_2(.din(w_dff_B_bZJxbUq97_2),.dout(w_dff_B_CVPIZxQW3_2),.clk(gclk));
	jdff dff_B_mWtJKION0_2(.din(w_dff_B_CVPIZxQW3_2),.dout(w_dff_B_mWtJKION0_2),.clk(gclk));
	jdff dff_B_53epCT4a7_2(.din(w_dff_B_mWtJKION0_2),.dout(w_dff_B_53epCT4a7_2),.clk(gclk));
	jdff dff_B_ZBEN2qtH8_2(.din(n721),.dout(w_dff_B_ZBEN2qtH8_2),.clk(gclk));
	jdff dff_B_mEGkhFkZ1_1(.din(n650),.dout(w_dff_B_mEGkhFkZ1_1),.clk(gclk));
	jdff dff_B_QNY9H9gw2_2(.din(n563),.dout(w_dff_B_QNY9H9gw2_2),.clk(gclk));
	jdff dff_B_qMXoEl3D7_2(.din(w_dff_B_QNY9H9gw2_2),.dout(w_dff_B_qMXoEl3D7_2),.clk(gclk));
	jdff dff_B_FInI1Q5Q0_2(.din(w_dff_B_qMXoEl3D7_2),.dout(w_dff_B_FInI1Q5Q0_2),.clk(gclk));
	jdff dff_B_Hj0o3xIa6_2(.din(w_dff_B_FInI1Q5Q0_2),.dout(w_dff_B_Hj0o3xIa6_2),.clk(gclk));
	jdff dff_B_PpNK2lKF5_2(.din(w_dff_B_Hj0o3xIa6_2),.dout(w_dff_B_PpNK2lKF5_2),.clk(gclk));
	jdff dff_B_6ruxRVpm7_2(.din(w_dff_B_PpNK2lKF5_2),.dout(w_dff_B_6ruxRVpm7_2),.clk(gclk));
	jdff dff_B_l1sk7anW1_2(.din(w_dff_B_6ruxRVpm7_2),.dout(w_dff_B_l1sk7anW1_2),.clk(gclk));
	jdff dff_B_0LpA89Jc7_2(.din(w_dff_B_l1sk7anW1_2),.dout(w_dff_B_0LpA89Jc7_2),.clk(gclk));
	jdff dff_B_1XyAd6jb9_2(.din(w_dff_B_0LpA89Jc7_2),.dout(w_dff_B_1XyAd6jb9_2),.clk(gclk));
	jdff dff_B_roRoidhf6_2(.din(w_dff_B_1XyAd6jb9_2),.dout(w_dff_B_roRoidhf6_2),.clk(gclk));
	jdff dff_B_Vh5jt5Ez2_2(.din(w_dff_B_roRoidhf6_2),.dout(w_dff_B_Vh5jt5Ez2_2),.clk(gclk));
	jdff dff_B_hZMrdm1s0_2(.din(w_dff_B_Vh5jt5Ez2_2),.dout(w_dff_B_hZMrdm1s0_2),.clk(gclk));
	jdff dff_B_bt2OBplg4_2(.din(w_dff_B_hZMrdm1s0_2),.dout(w_dff_B_bt2OBplg4_2),.clk(gclk));
	jdff dff_B_2CCavDMt0_2(.din(w_dff_B_bt2OBplg4_2),.dout(w_dff_B_2CCavDMt0_2),.clk(gclk));
	jdff dff_B_pAgxNNHr2_2(.din(w_dff_B_2CCavDMt0_2),.dout(w_dff_B_pAgxNNHr2_2),.clk(gclk));
	jdff dff_B_uTiVbRAA8_2(.din(w_dff_B_pAgxNNHr2_2),.dout(w_dff_B_uTiVbRAA8_2),.clk(gclk));
	jdff dff_B_Zbqh0ZSs0_2(.din(w_dff_B_uTiVbRAA8_2),.dout(w_dff_B_Zbqh0ZSs0_2),.clk(gclk));
	jdff dff_B_w5XslQ6o1_2(.din(w_dff_B_Zbqh0ZSs0_2),.dout(w_dff_B_w5XslQ6o1_2),.clk(gclk));
	jdff dff_B_5DNGVSKm0_2(.din(w_dff_B_w5XslQ6o1_2),.dout(w_dff_B_5DNGVSKm0_2),.clk(gclk));
	jdff dff_B_EewqZM6m7_2(.din(w_dff_B_5DNGVSKm0_2),.dout(w_dff_B_EewqZM6m7_2),.clk(gclk));
	jdff dff_B_KnMiODfg2_2(.din(w_dff_B_EewqZM6m7_2),.dout(w_dff_B_KnMiODfg2_2),.clk(gclk));
	jdff dff_B_ptY0swbn7_2(.din(w_dff_B_KnMiODfg2_2),.dout(w_dff_B_ptY0swbn7_2),.clk(gclk));
	jdff dff_B_kjBbuBWi9_2(.din(w_dff_B_ptY0swbn7_2),.dout(w_dff_B_kjBbuBWi9_2),.clk(gclk));
	jdff dff_B_D96xFsyD7_2(.din(w_dff_B_kjBbuBWi9_2),.dout(w_dff_B_D96xFsyD7_2),.clk(gclk));
	jdff dff_B_LoGBgwd11_2(.din(w_dff_B_D96xFsyD7_2),.dout(w_dff_B_LoGBgwd11_2),.clk(gclk));
	jdff dff_B_XYasrhLl9_2(.din(w_dff_B_LoGBgwd11_2),.dout(w_dff_B_XYasrhLl9_2),.clk(gclk));
	jdff dff_B_xk4ibRrF9_2(.din(w_dff_B_XYasrhLl9_2),.dout(w_dff_B_xk4ibRrF9_2),.clk(gclk));
	jdff dff_B_S0rXoPdI4_2(.din(w_dff_B_xk4ibRrF9_2),.dout(w_dff_B_S0rXoPdI4_2),.clk(gclk));
	jdff dff_B_9FCmbrcm4_2(.din(n628),.dout(w_dff_B_9FCmbrcm4_2),.clk(gclk));
	jdff dff_B_qm7W71SE7_1(.din(n564),.dout(w_dff_B_qm7W71SE7_1),.clk(gclk));
	jdff dff_B_UJCveD5s6_2(.din(n484),.dout(w_dff_B_UJCveD5s6_2),.clk(gclk));
	jdff dff_B_XhEtsp7o1_2(.din(w_dff_B_UJCveD5s6_2),.dout(w_dff_B_XhEtsp7o1_2),.clk(gclk));
	jdff dff_B_7TDTOO5L2_2(.din(w_dff_B_XhEtsp7o1_2),.dout(w_dff_B_7TDTOO5L2_2),.clk(gclk));
	jdff dff_B_j6oRqiWS4_2(.din(w_dff_B_7TDTOO5L2_2),.dout(w_dff_B_j6oRqiWS4_2),.clk(gclk));
	jdff dff_B_2GhB4nT59_2(.din(w_dff_B_j6oRqiWS4_2),.dout(w_dff_B_2GhB4nT59_2),.clk(gclk));
	jdff dff_B_ccEB6Pcf4_2(.din(w_dff_B_2GhB4nT59_2),.dout(w_dff_B_ccEB6Pcf4_2),.clk(gclk));
	jdff dff_B_oBomMU8s7_2(.din(w_dff_B_ccEB6Pcf4_2),.dout(w_dff_B_oBomMU8s7_2),.clk(gclk));
	jdff dff_B_KNKsVjQm0_2(.din(w_dff_B_oBomMU8s7_2),.dout(w_dff_B_KNKsVjQm0_2),.clk(gclk));
	jdff dff_B_nt40BZEQ4_2(.din(w_dff_B_KNKsVjQm0_2),.dout(w_dff_B_nt40BZEQ4_2),.clk(gclk));
	jdff dff_B_Rwy0X4qp1_2(.din(w_dff_B_nt40BZEQ4_2),.dout(w_dff_B_Rwy0X4qp1_2),.clk(gclk));
	jdff dff_B_k9NhsHdL9_2(.din(w_dff_B_Rwy0X4qp1_2),.dout(w_dff_B_k9NhsHdL9_2),.clk(gclk));
	jdff dff_B_OgDnLGtX7_2(.din(w_dff_B_k9NhsHdL9_2),.dout(w_dff_B_OgDnLGtX7_2),.clk(gclk));
	jdff dff_B_pPJF5NhR9_2(.din(w_dff_B_OgDnLGtX7_2),.dout(w_dff_B_pPJF5NhR9_2),.clk(gclk));
	jdff dff_B_kc4KIVQx5_2(.din(w_dff_B_pPJF5NhR9_2),.dout(w_dff_B_kc4KIVQx5_2),.clk(gclk));
	jdff dff_B_IC22vasF6_2(.din(w_dff_B_kc4KIVQx5_2),.dout(w_dff_B_IC22vasF6_2),.clk(gclk));
	jdff dff_B_f1wTeq276_2(.din(w_dff_B_IC22vasF6_2),.dout(w_dff_B_f1wTeq276_2),.clk(gclk));
	jdff dff_B_vBVb1UCN5_2(.din(w_dff_B_f1wTeq276_2),.dout(w_dff_B_vBVb1UCN5_2),.clk(gclk));
	jdff dff_B_BhBeVO2I9_2(.din(w_dff_B_vBVb1UCN5_2),.dout(w_dff_B_BhBeVO2I9_2),.clk(gclk));
	jdff dff_B_FSxNYMdQ9_2(.din(w_dff_B_BhBeVO2I9_2),.dout(w_dff_B_FSxNYMdQ9_2),.clk(gclk));
	jdff dff_B_N8DuCpGu2_2(.din(w_dff_B_FSxNYMdQ9_2),.dout(w_dff_B_N8DuCpGu2_2),.clk(gclk));
	jdff dff_B_kiSpnneP1_2(.din(w_dff_B_N8DuCpGu2_2),.dout(w_dff_B_kiSpnneP1_2),.clk(gclk));
	jdff dff_B_YPdz383g3_2(.din(w_dff_B_kiSpnneP1_2),.dout(w_dff_B_YPdz383g3_2),.clk(gclk));
	jdff dff_B_GgPbChkp9_2(.din(w_dff_B_YPdz383g3_2),.dout(w_dff_B_GgPbChkp9_2),.clk(gclk));
	jdff dff_B_I8e2cYpL6_2(.din(w_dff_B_GgPbChkp9_2),.dout(w_dff_B_I8e2cYpL6_2),.clk(gclk));
	jdff dff_B_CCND9ubK0_2(.din(w_dff_B_I8e2cYpL6_2),.dout(w_dff_B_CCND9ubK0_2),.clk(gclk));
	jdff dff_B_WcIQi2vz7_2(.din(n542),.dout(w_dff_B_WcIQi2vz7_2),.clk(gclk));
	jdff dff_B_Voqlg2Yh1_1(.din(n485),.dout(w_dff_B_Voqlg2Yh1_1),.clk(gclk));
	jdff dff_B_sdAh0Vr59_2(.din(n412),.dout(w_dff_B_sdAh0Vr59_2),.clk(gclk));
	jdff dff_B_HWYeEN6q5_2(.din(w_dff_B_sdAh0Vr59_2),.dout(w_dff_B_HWYeEN6q5_2),.clk(gclk));
	jdff dff_B_EbCUtrqW3_2(.din(w_dff_B_HWYeEN6q5_2),.dout(w_dff_B_EbCUtrqW3_2),.clk(gclk));
	jdff dff_B_pybQll3U4_2(.din(w_dff_B_EbCUtrqW3_2),.dout(w_dff_B_pybQll3U4_2),.clk(gclk));
	jdff dff_B_F7jBQweO7_2(.din(w_dff_B_pybQll3U4_2),.dout(w_dff_B_F7jBQweO7_2),.clk(gclk));
	jdff dff_B_2vXrbfAh1_2(.din(w_dff_B_F7jBQweO7_2),.dout(w_dff_B_2vXrbfAh1_2),.clk(gclk));
	jdff dff_B_0YqPQxRO0_2(.din(w_dff_B_2vXrbfAh1_2),.dout(w_dff_B_0YqPQxRO0_2),.clk(gclk));
	jdff dff_B_o4abx7OD4_2(.din(w_dff_B_0YqPQxRO0_2),.dout(w_dff_B_o4abx7OD4_2),.clk(gclk));
	jdff dff_B_BbHWM7GS3_2(.din(w_dff_B_o4abx7OD4_2),.dout(w_dff_B_BbHWM7GS3_2),.clk(gclk));
	jdff dff_B_O3NBLQHP3_2(.din(w_dff_B_BbHWM7GS3_2),.dout(w_dff_B_O3NBLQHP3_2),.clk(gclk));
	jdff dff_B_HfLyjiRQ8_2(.din(w_dff_B_O3NBLQHP3_2),.dout(w_dff_B_HfLyjiRQ8_2),.clk(gclk));
	jdff dff_B_GlUM8oqM5_2(.din(w_dff_B_HfLyjiRQ8_2),.dout(w_dff_B_GlUM8oqM5_2),.clk(gclk));
	jdff dff_B_6HUbN8uF2_2(.din(w_dff_B_GlUM8oqM5_2),.dout(w_dff_B_6HUbN8uF2_2),.clk(gclk));
	jdff dff_B_nkT76NXQ8_2(.din(w_dff_B_6HUbN8uF2_2),.dout(w_dff_B_nkT76NXQ8_2),.clk(gclk));
	jdff dff_B_fX5wZIZn9_2(.din(w_dff_B_nkT76NXQ8_2),.dout(w_dff_B_fX5wZIZn9_2),.clk(gclk));
	jdff dff_B_rvPz3zkP7_2(.din(w_dff_B_fX5wZIZn9_2),.dout(w_dff_B_rvPz3zkP7_2),.clk(gclk));
	jdff dff_B_ljo04jbn2_2(.din(w_dff_B_rvPz3zkP7_2),.dout(w_dff_B_ljo04jbn2_2),.clk(gclk));
	jdff dff_B_V1ZSVRvV4_2(.din(w_dff_B_ljo04jbn2_2),.dout(w_dff_B_V1ZSVRvV4_2),.clk(gclk));
	jdff dff_B_YvxezPYK2_2(.din(w_dff_B_V1ZSVRvV4_2),.dout(w_dff_B_YvxezPYK2_2),.clk(gclk));
	jdff dff_B_M3KLAOSb8_2(.din(w_dff_B_YvxezPYK2_2),.dout(w_dff_B_M3KLAOSb8_2),.clk(gclk));
	jdff dff_B_QdKVDZSg5_2(.din(w_dff_B_M3KLAOSb8_2),.dout(w_dff_B_QdKVDZSg5_2),.clk(gclk));
	jdff dff_B_m3egyPwj4_2(.din(w_dff_B_QdKVDZSg5_2),.dout(w_dff_B_m3egyPwj4_2),.clk(gclk));
	jdff dff_B_A822Pj3E2_2(.din(n463),.dout(w_dff_B_A822Pj3E2_2),.clk(gclk));
	jdff dff_B_NdpLZSRB4_1(.din(n413),.dout(w_dff_B_NdpLZSRB4_1),.clk(gclk));
	jdff dff_B_XUqUdk527_2(.din(n348),.dout(w_dff_B_XUqUdk527_2),.clk(gclk));
	jdff dff_B_mfiIfL1c9_2(.din(w_dff_B_XUqUdk527_2),.dout(w_dff_B_mfiIfL1c9_2),.clk(gclk));
	jdff dff_B_CaB7WW3i5_2(.din(w_dff_B_mfiIfL1c9_2),.dout(w_dff_B_CaB7WW3i5_2),.clk(gclk));
	jdff dff_B_a7SQIuAl9_2(.din(w_dff_B_CaB7WW3i5_2),.dout(w_dff_B_a7SQIuAl9_2),.clk(gclk));
	jdff dff_B_i1YtFsae0_2(.din(w_dff_B_a7SQIuAl9_2),.dout(w_dff_B_i1YtFsae0_2),.clk(gclk));
	jdff dff_B_LgQKcvdf3_2(.din(w_dff_B_i1YtFsae0_2),.dout(w_dff_B_LgQKcvdf3_2),.clk(gclk));
	jdff dff_B_iHry2Aq55_2(.din(w_dff_B_LgQKcvdf3_2),.dout(w_dff_B_iHry2Aq55_2),.clk(gclk));
	jdff dff_B_mMgSrYur5_2(.din(w_dff_B_iHry2Aq55_2),.dout(w_dff_B_mMgSrYur5_2),.clk(gclk));
	jdff dff_B_eNYHndts9_2(.din(w_dff_B_mMgSrYur5_2),.dout(w_dff_B_eNYHndts9_2),.clk(gclk));
	jdff dff_B_L2PolUdN0_2(.din(w_dff_B_eNYHndts9_2),.dout(w_dff_B_L2PolUdN0_2),.clk(gclk));
	jdff dff_B_ajjNMWC26_2(.din(w_dff_B_L2PolUdN0_2),.dout(w_dff_B_ajjNMWC26_2),.clk(gclk));
	jdff dff_B_zfI7wkQw6_2(.din(w_dff_B_ajjNMWC26_2),.dout(w_dff_B_zfI7wkQw6_2),.clk(gclk));
	jdff dff_B_qCWSYLrs6_2(.din(w_dff_B_zfI7wkQw6_2),.dout(w_dff_B_qCWSYLrs6_2),.clk(gclk));
	jdff dff_B_1wvC4odU9_2(.din(w_dff_B_qCWSYLrs6_2),.dout(w_dff_B_1wvC4odU9_2),.clk(gclk));
	jdff dff_B_PUpj6HfG9_2(.din(w_dff_B_1wvC4odU9_2),.dout(w_dff_B_PUpj6HfG9_2),.clk(gclk));
	jdff dff_B_LMGXKl6t7_2(.din(w_dff_B_PUpj6HfG9_2),.dout(w_dff_B_LMGXKl6t7_2),.clk(gclk));
	jdff dff_B_5BpYIurk2_2(.din(w_dff_B_LMGXKl6t7_2),.dout(w_dff_B_5BpYIurk2_2),.clk(gclk));
	jdff dff_B_ag9VBo1Y6_2(.din(w_dff_B_5BpYIurk2_2),.dout(w_dff_B_ag9VBo1Y6_2),.clk(gclk));
	jdff dff_B_o72n8RB88_2(.din(w_dff_B_ag9VBo1Y6_2),.dout(w_dff_B_o72n8RB88_2),.clk(gclk));
	jdff dff_B_ce9XI3zW7_2(.din(n391),.dout(w_dff_B_ce9XI3zW7_2),.clk(gclk));
	jdff dff_B_jDbqou9V2_1(.din(n349),.dout(w_dff_B_jDbqou9V2_1),.clk(gclk));
	jdff dff_B_7GHg35vR0_2(.din(n290),.dout(w_dff_B_7GHg35vR0_2),.clk(gclk));
	jdff dff_B_oCDg3lK08_2(.din(w_dff_B_7GHg35vR0_2),.dout(w_dff_B_oCDg3lK08_2),.clk(gclk));
	jdff dff_B_TcUJFPef2_2(.din(w_dff_B_oCDg3lK08_2),.dout(w_dff_B_TcUJFPef2_2),.clk(gclk));
	jdff dff_B_HzEkmRhg0_2(.din(w_dff_B_TcUJFPef2_2),.dout(w_dff_B_HzEkmRhg0_2),.clk(gclk));
	jdff dff_B_LWuWehQz4_2(.din(w_dff_B_HzEkmRhg0_2),.dout(w_dff_B_LWuWehQz4_2),.clk(gclk));
	jdff dff_B_5P0B3daq3_2(.din(w_dff_B_LWuWehQz4_2),.dout(w_dff_B_5P0B3daq3_2),.clk(gclk));
	jdff dff_B_QLyzIFN62_2(.din(w_dff_B_5P0B3daq3_2),.dout(w_dff_B_QLyzIFN62_2),.clk(gclk));
	jdff dff_B_QWjgs8c67_2(.din(w_dff_B_QLyzIFN62_2),.dout(w_dff_B_QWjgs8c67_2),.clk(gclk));
	jdff dff_B_snrHGHww9_2(.din(w_dff_B_QWjgs8c67_2),.dout(w_dff_B_snrHGHww9_2),.clk(gclk));
	jdff dff_B_NXZQbBGI2_2(.din(w_dff_B_snrHGHww9_2),.dout(w_dff_B_NXZQbBGI2_2),.clk(gclk));
	jdff dff_B_uvL3rfcW6_2(.din(w_dff_B_NXZQbBGI2_2),.dout(w_dff_B_uvL3rfcW6_2),.clk(gclk));
	jdff dff_B_m7NKtxLp4_2(.din(w_dff_B_uvL3rfcW6_2),.dout(w_dff_B_m7NKtxLp4_2),.clk(gclk));
	jdff dff_B_EYmoJy0P8_2(.din(w_dff_B_m7NKtxLp4_2),.dout(w_dff_B_EYmoJy0P8_2),.clk(gclk));
	jdff dff_B_oXEPrpvp0_2(.din(w_dff_B_EYmoJy0P8_2),.dout(w_dff_B_oXEPrpvp0_2),.clk(gclk));
	jdff dff_B_B8d0Foqb2_2(.din(w_dff_B_oXEPrpvp0_2),.dout(w_dff_B_B8d0Foqb2_2),.clk(gclk));
	jdff dff_B_9vo0u5m23_2(.din(w_dff_B_B8d0Foqb2_2),.dout(w_dff_B_9vo0u5m23_2),.clk(gclk));
	jdff dff_B_3RE2EL7P0_2(.din(n327),.dout(w_dff_B_3RE2EL7P0_2),.clk(gclk));
	jdff dff_B_al8aNhS70_1(.din(n291),.dout(w_dff_B_al8aNhS70_1),.clk(gclk));
	jdff dff_B_k6V0TNG19_2(.din(n239),.dout(w_dff_B_k6V0TNG19_2),.clk(gclk));
	jdff dff_B_MXawkFPT4_2(.din(w_dff_B_k6V0TNG19_2),.dout(w_dff_B_MXawkFPT4_2),.clk(gclk));
	jdff dff_B_1othvyRy4_2(.din(w_dff_B_MXawkFPT4_2),.dout(w_dff_B_1othvyRy4_2),.clk(gclk));
	jdff dff_B_r2xHZHD81_2(.din(w_dff_B_1othvyRy4_2),.dout(w_dff_B_r2xHZHD81_2),.clk(gclk));
	jdff dff_B_mO3HnqJG0_2(.din(w_dff_B_r2xHZHD81_2),.dout(w_dff_B_mO3HnqJG0_2),.clk(gclk));
	jdff dff_B_D7ZVLqB92_2(.din(w_dff_B_mO3HnqJG0_2),.dout(w_dff_B_D7ZVLqB92_2),.clk(gclk));
	jdff dff_B_N433o7ZI4_2(.din(w_dff_B_D7ZVLqB92_2),.dout(w_dff_B_N433o7ZI4_2),.clk(gclk));
	jdff dff_B_BdcSgprP4_2(.din(w_dff_B_N433o7ZI4_2),.dout(w_dff_B_BdcSgprP4_2),.clk(gclk));
	jdff dff_B_qRGWIEP82_2(.din(w_dff_B_BdcSgprP4_2),.dout(w_dff_B_qRGWIEP82_2),.clk(gclk));
	jdff dff_B_22AIujaK0_2(.din(w_dff_B_qRGWIEP82_2),.dout(w_dff_B_22AIujaK0_2),.clk(gclk));
	jdff dff_B_03nXaE3f7_2(.din(w_dff_B_22AIujaK0_2),.dout(w_dff_B_03nXaE3f7_2),.clk(gclk));
	jdff dff_B_UjOpp8Dk8_2(.din(w_dff_B_03nXaE3f7_2),.dout(w_dff_B_UjOpp8Dk8_2),.clk(gclk));
	jdff dff_B_psODmytO6_2(.din(w_dff_B_UjOpp8Dk8_2),.dout(w_dff_B_psODmytO6_2),.clk(gclk));
	jdff dff_B_DveKxQYH6_2(.din(n269),.dout(w_dff_B_DveKxQYH6_2),.clk(gclk));
	jdff dff_B_2fcWdJM90_1(.din(n240),.dout(w_dff_B_2fcWdJM90_1),.clk(gclk));
	jdff dff_B_v1Z9jLdn7_2(.din(n196),.dout(w_dff_B_v1Z9jLdn7_2),.clk(gclk));
	jdff dff_B_OGDdeCCB7_2(.din(w_dff_B_v1Z9jLdn7_2),.dout(w_dff_B_OGDdeCCB7_2),.clk(gclk));
	jdff dff_B_G8xzG6C29_2(.din(w_dff_B_OGDdeCCB7_2),.dout(w_dff_B_G8xzG6C29_2),.clk(gclk));
	jdff dff_B_UERly8ar0_2(.din(w_dff_B_G8xzG6C29_2),.dout(w_dff_B_UERly8ar0_2),.clk(gclk));
	jdff dff_B_2xCgGoC53_2(.din(w_dff_B_UERly8ar0_2),.dout(w_dff_B_2xCgGoC53_2),.clk(gclk));
	jdff dff_B_Yrxj0Kgk9_2(.din(w_dff_B_2xCgGoC53_2),.dout(w_dff_B_Yrxj0Kgk9_2),.clk(gclk));
	jdff dff_B_4WYVfu2E8_2(.din(w_dff_B_Yrxj0Kgk9_2),.dout(w_dff_B_4WYVfu2E8_2),.clk(gclk));
	jdff dff_B_vMZ5OOKg0_2(.din(w_dff_B_4WYVfu2E8_2),.dout(w_dff_B_vMZ5OOKg0_2),.clk(gclk));
	jdff dff_B_d8kcAuRM0_2(.din(w_dff_B_vMZ5OOKg0_2),.dout(w_dff_B_d8kcAuRM0_2),.clk(gclk));
	jdff dff_B_tViMIGoP6_2(.din(w_dff_B_d8kcAuRM0_2),.dout(w_dff_B_tViMIGoP6_2),.clk(gclk));
	jdff dff_B_LYxRxdqy1_2(.din(n218),.dout(w_dff_B_LYxRxdqy1_2),.clk(gclk));
	jdff dff_B_5TW31LH74_1(.din(n197),.dout(w_dff_B_5TW31LH74_1),.clk(gclk));
	jdff dff_B_pklqfeAD2_2(.din(n158),.dout(w_dff_B_pklqfeAD2_2),.clk(gclk));
	jdff dff_B_VIApfomQ3_2(.din(w_dff_B_pklqfeAD2_2),.dout(w_dff_B_VIApfomQ3_2),.clk(gclk));
	jdff dff_B_znQYor7B9_2(.din(w_dff_B_VIApfomQ3_2),.dout(w_dff_B_znQYor7B9_2),.clk(gclk));
	jdff dff_B_kDZqI6jJ4_2(.din(w_dff_B_znQYor7B9_2),.dout(w_dff_B_kDZqI6jJ4_2),.clk(gclk));
	jdff dff_B_q4MDs3Rk9_2(.din(w_dff_B_kDZqI6jJ4_2),.dout(w_dff_B_q4MDs3Rk9_2),.clk(gclk));
	jdff dff_B_dCnCZZZE5_2(.din(w_dff_B_q4MDs3Rk9_2),.dout(w_dff_B_dCnCZZZE5_2),.clk(gclk));
	jdff dff_B_p6mphz8N5_2(.din(w_dff_B_dCnCZZZE5_2),.dout(w_dff_B_p6mphz8N5_2),.clk(gclk));
	jdff dff_B_JHKovzKr2_2(.din(n175),.dout(w_dff_B_JHKovzKr2_2),.clk(gclk));
	jdff dff_B_Lo1si02i0_1(.din(n161),.dout(w_dff_B_Lo1si02i0_1),.clk(gclk));
	jdff dff_B_xBFu5Phx7_1(.din(w_dff_B_Lo1si02i0_1),.dout(w_dff_B_xBFu5Phx7_1),.clk(gclk));
	jdff dff_B_98WjUXC83_2(.din(n128),.dout(w_dff_B_98WjUXC83_2),.clk(gclk));
	jdff dff_B_cZeyvtrC4_2(.din(w_dff_B_98WjUXC83_2),.dout(w_dff_B_cZeyvtrC4_2),.clk(gclk));
	jdff dff_B_fODRA8fO1_2(.din(w_dff_B_cZeyvtrC4_2),.dout(w_dff_B_fODRA8fO1_2),.clk(gclk));
	jdff dff_B_s8Xsddgu1_2(.din(w_dff_B_fODRA8fO1_2),.dout(w_dff_B_s8Xsddgu1_2),.clk(gclk));
	jdff dff_A_R32qMOHF2_1(.dout(w_n130_0[1]),.din(w_dff_A_R32qMOHF2_1),.clk(gclk));
	jdff dff_A_D2IVofeZ1_0(.dout(w_n101_0[0]),.din(w_dff_A_D2IVofeZ1_0),.clk(gclk));
	jdff dff_A_9S0is7Qi5_0(.dout(w_n100_1[0]),.din(w_dff_A_9S0is7Qi5_0),.clk(gclk));
	jdff dff_A_8BlzFoWF9_1(.dout(w_n100_0[1]),.din(w_dff_A_8BlzFoWF9_1),.clk(gclk));
	jdff dff_A_NwSCs7bj4_2(.dout(w_n100_0[2]),.din(w_dff_A_NwSCs7bj4_2),.clk(gclk));
	jdff dff_A_ZXYPmR2t3_2(.dout(w_dff_A_NwSCs7bj4_2),.din(w_dff_A_ZXYPmR2t3_2),.clk(gclk));
	jdff dff_B_yOr46Oam9_0(.din(n1329),.dout(w_dff_B_yOr46Oam9_0),.clk(gclk));
	jdff dff_A_U692QmXf8_1(.dout(w_n1325_0[1]),.din(w_dff_A_U692QmXf8_1),.clk(gclk));
	jdff dff_A_IPnXeFHN0_1(.dout(w_dff_A_U692QmXf8_1),.din(w_dff_A_IPnXeFHN0_1),.clk(gclk));
	jdff dff_B_i5Q5GgX24_1(.din(n1245),.dout(w_dff_B_i5Q5GgX24_1),.clk(gclk));
	jdff dff_B_JNPv3mIo9_1(.din(w_dff_B_i5Q5GgX24_1),.dout(w_dff_B_JNPv3mIo9_1),.clk(gclk));
	jdff dff_B_jAaslnVt5_2(.din(n1152),.dout(w_dff_B_jAaslnVt5_2),.clk(gclk));
	jdff dff_B_WDRKdxAH1_2(.din(w_dff_B_jAaslnVt5_2),.dout(w_dff_B_WDRKdxAH1_2),.clk(gclk));
	jdff dff_B_f9uoqLHw5_2(.din(w_dff_B_WDRKdxAH1_2),.dout(w_dff_B_f9uoqLHw5_2),.clk(gclk));
	jdff dff_B_AMSHqjDG7_2(.din(w_dff_B_f9uoqLHw5_2),.dout(w_dff_B_AMSHqjDG7_2),.clk(gclk));
	jdff dff_B_o9VwloPg3_2(.din(w_dff_B_AMSHqjDG7_2),.dout(w_dff_B_o9VwloPg3_2),.clk(gclk));
	jdff dff_B_ay0dwz2M9_2(.din(w_dff_B_o9VwloPg3_2),.dout(w_dff_B_ay0dwz2M9_2),.clk(gclk));
	jdff dff_B_rkuvduRC8_2(.din(w_dff_B_ay0dwz2M9_2),.dout(w_dff_B_rkuvduRC8_2),.clk(gclk));
	jdff dff_B_SxoeFFU92_2(.din(w_dff_B_rkuvduRC8_2),.dout(w_dff_B_SxoeFFU92_2),.clk(gclk));
	jdff dff_B_nrRDnhYj9_2(.din(w_dff_B_SxoeFFU92_2),.dout(w_dff_B_nrRDnhYj9_2),.clk(gclk));
	jdff dff_B_P9wYd6x00_2(.din(w_dff_B_nrRDnhYj9_2),.dout(w_dff_B_P9wYd6x00_2),.clk(gclk));
	jdff dff_B_u1Gkuo0E9_2(.din(w_dff_B_P9wYd6x00_2),.dout(w_dff_B_u1Gkuo0E9_2),.clk(gclk));
	jdff dff_B_TiZHioho0_2(.din(w_dff_B_u1Gkuo0E9_2),.dout(w_dff_B_TiZHioho0_2),.clk(gclk));
	jdff dff_B_xicjWSWt0_2(.din(w_dff_B_TiZHioho0_2),.dout(w_dff_B_xicjWSWt0_2),.clk(gclk));
	jdff dff_B_Z9PyoSK47_2(.din(w_dff_B_xicjWSWt0_2),.dout(w_dff_B_Z9PyoSK47_2),.clk(gclk));
	jdff dff_B_2ifOi42V8_2(.din(w_dff_B_Z9PyoSK47_2),.dout(w_dff_B_2ifOi42V8_2),.clk(gclk));
	jdff dff_B_XhAMf2eX6_2(.din(w_dff_B_2ifOi42V8_2),.dout(w_dff_B_XhAMf2eX6_2),.clk(gclk));
	jdff dff_B_eaDWm4203_2(.din(w_dff_B_XhAMf2eX6_2),.dout(w_dff_B_eaDWm4203_2),.clk(gclk));
	jdff dff_B_6vWy6wCL8_2(.din(w_dff_B_eaDWm4203_2),.dout(w_dff_B_6vWy6wCL8_2),.clk(gclk));
	jdff dff_B_qxi5hrBP4_2(.din(w_dff_B_6vWy6wCL8_2),.dout(w_dff_B_qxi5hrBP4_2),.clk(gclk));
	jdff dff_B_VyECjBLD2_2(.din(w_dff_B_qxi5hrBP4_2),.dout(w_dff_B_VyECjBLD2_2),.clk(gclk));
	jdff dff_B_e6XjtRon2_2(.din(w_dff_B_VyECjBLD2_2),.dout(w_dff_B_e6XjtRon2_2),.clk(gclk));
	jdff dff_B_CrYiwVtH3_2(.din(w_dff_B_e6XjtRon2_2),.dout(w_dff_B_CrYiwVtH3_2),.clk(gclk));
	jdff dff_B_kCnhktvL1_2(.din(w_dff_B_CrYiwVtH3_2),.dout(w_dff_B_kCnhktvL1_2),.clk(gclk));
	jdff dff_B_fqGu5zJg1_2(.din(w_dff_B_kCnhktvL1_2),.dout(w_dff_B_fqGu5zJg1_2),.clk(gclk));
	jdff dff_B_scwyyet63_2(.din(w_dff_B_fqGu5zJg1_2),.dout(w_dff_B_scwyyet63_2),.clk(gclk));
	jdff dff_B_0guQVbUe6_2(.din(w_dff_B_scwyyet63_2),.dout(w_dff_B_0guQVbUe6_2),.clk(gclk));
	jdff dff_B_h1VlblDI5_2(.din(w_dff_B_0guQVbUe6_2),.dout(w_dff_B_h1VlblDI5_2),.clk(gclk));
	jdff dff_B_EA0GKumX9_2(.din(w_dff_B_h1VlblDI5_2),.dout(w_dff_B_EA0GKumX9_2),.clk(gclk));
	jdff dff_B_uP1G5RxD5_2(.din(w_dff_B_EA0GKumX9_2),.dout(w_dff_B_uP1G5RxD5_2),.clk(gclk));
	jdff dff_B_WVF5oxW86_2(.din(w_dff_B_uP1G5RxD5_2),.dout(w_dff_B_WVF5oxW86_2),.clk(gclk));
	jdff dff_B_RU3lt3cc7_2(.din(w_dff_B_WVF5oxW86_2),.dout(w_dff_B_RU3lt3cc7_2),.clk(gclk));
	jdff dff_B_u0KFp77y1_2(.din(w_dff_B_RU3lt3cc7_2),.dout(w_dff_B_u0KFp77y1_2),.clk(gclk));
	jdff dff_B_S09I4NAK0_2(.din(w_dff_B_u0KFp77y1_2),.dout(w_dff_B_S09I4NAK0_2),.clk(gclk));
	jdff dff_B_1iXi2EKq2_2(.din(w_dff_B_S09I4NAK0_2),.dout(w_dff_B_1iXi2EKq2_2),.clk(gclk));
	jdff dff_B_We1EybXJ2_2(.din(w_dff_B_1iXi2EKq2_2),.dout(w_dff_B_We1EybXJ2_2),.clk(gclk));
	jdff dff_B_wAilYS1r5_2(.din(w_dff_B_We1EybXJ2_2),.dout(w_dff_B_wAilYS1r5_2),.clk(gclk));
	jdff dff_B_ChOaTK1q7_2(.din(w_dff_B_wAilYS1r5_2),.dout(w_dff_B_ChOaTK1q7_2),.clk(gclk));
	jdff dff_B_seCLvjU91_2(.din(w_dff_B_ChOaTK1q7_2),.dout(w_dff_B_seCLvjU91_2),.clk(gclk));
	jdff dff_B_zhzxnqSk0_2(.din(w_dff_B_seCLvjU91_2),.dout(w_dff_B_zhzxnqSk0_2),.clk(gclk));
	jdff dff_B_Od0HTU9o4_2(.din(w_dff_B_zhzxnqSk0_2),.dout(w_dff_B_Od0HTU9o4_2),.clk(gclk));
	jdff dff_B_BITHYmtq6_2(.din(w_dff_B_Od0HTU9o4_2),.dout(w_dff_B_BITHYmtq6_2),.clk(gclk));
	jdff dff_B_efLQbOd50_2(.din(w_dff_B_BITHYmtq6_2),.dout(w_dff_B_efLQbOd50_2),.clk(gclk));
	jdff dff_B_u5obT7YS6_2(.din(w_dff_B_efLQbOd50_2),.dout(w_dff_B_u5obT7YS6_2),.clk(gclk));
	jdff dff_B_K0dT0OMv0_2(.din(w_dff_B_u5obT7YS6_2),.dout(w_dff_B_K0dT0OMv0_2),.clk(gclk));
	jdff dff_B_OtPzkkDJ3_2(.din(w_dff_B_K0dT0OMv0_2),.dout(w_dff_B_OtPzkkDJ3_2),.clk(gclk));
	jdff dff_B_Ycu9g66M0_2(.din(w_dff_B_OtPzkkDJ3_2),.dout(w_dff_B_Ycu9g66M0_2),.clk(gclk));
	jdff dff_B_DxnsUaBS1_2(.din(n1234),.dout(w_dff_B_DxnsUaBS1_2),.clk(gclk));
	jdff dff_B_DOH2dNe61_1(.din(n1154),.dout(w_dff_B_DOH2dNe61_1),.clk(gclk));
	jdff dff_B_Dm35Epxf3_2(.din(n1049),.dout(w_dff_B_Dm35Epxf3_2),.clk(gclk));
	jdff dff_B_spdaXV6m5_2(.din(w_dff_B_Dm35Epxf3_2),.dout(w_dff_B_spdaXV6m5_2),.clk(gclk));
	jdff dff_B_6FcRjeyT7_2(.din(w_dff_B_spdaXV6m5_2),.dout(w_dff_B_6FcRjeyT7_2),.clk(gclk));
	jdff dff_B_Eab1VxWV3_2(.din(w_dff_B_6FcRjeyT7_2),.dout(w_dff_B_Eab1VxWV3_2),.clk(gclk));
	jdff dff_B_XEXLONgk2_2(.din(w_dff_B_Eab1VxWV3_2),.dout(w_dff_B_XEXLONgk2_2),.clk(gclk));
	jdff dff_B_y8ZMA8v00_2(.din(w_dff_B_XEXLONgk2_2),.dout(w_dff_B_y8ZMA8v00_2),.clk(gclk));
	jdff dff_B_WHEhknZP7_2(.din(w_dff_B_y8ZMA8v00_2),.dout(w_dff_B_WHEhknZP7_2),.clk(gclk));
	jdff dff_B_PwaeNsOc6_2(.din(w_dff_B_WHEhknZP7_2),.dout(w_dff_B_PwaeNsOc6_2),.clk(gclk));
	jdff dff_B_PKsSXaIl1_2(.din(w_dff_B_PwaeNsOc6_2),.dout(w_dff_B_PKsSXaIl1_2),.clk(gclk));
	jdff dff_B_M81eb61a7_2(.din(w_dff_B_PKsSXaIl1_2),.dout(w_dff_B_M81eb61a7_2),.clk(gclk));
	jdff dff_B_scetwMPr7_2(.din(w_dff_B_M81eb61a7_2),.dout(w_dff_B_scetwMPr7_2),.clk(gclk));
	jdff dff_B_X7d9ZqKg6_2(.din(w_dff_B_scetwMPr7_2),.dout(w_dff_B_X7d9ZqKg6_2),.clk(gclk));
	jdff dff_B_B5jRDPeS3_2(.din(w_dff_B_X7d9ZqKg6_2),.dout(w_dff_B_B5jRDPeS3_2),.clk(gclk));
	jdff dff_B_dCPPhaFI7_2(.din(w_dff_B_B5jRDPeS3_2),.dout(w_dff_B_dCPPhaFI7_2),.clk(gclk));
	jdff dff_B_J3QBwTyD9_2(.din(w_dff_B_dCPPhaFI7_2),.dout(w_dff_B_J3QBwTyD9_2),.clk(gclk));
	jdff dff_B_KtSpz4A72_2(.din(w_dff_B_J3QBwTyD9_2),.dout(w_dff_B_KtSpz4A72_2),.clk(gclk));
	jdff dff_B_X7xx28KV1_2(.din(w_dff_B_KtSpz4A72_2),.dout(w_dff_B_X7xx28KV1_2),.clk(gclk));
	jdff dff_B_20jGAzNF7_2(.din(w_dff_B_X7xx28KV1_2),.dout(w_dff_B_20jGAzNF7_2),.clk(gclk));
	jdff dff_B_dH5f8ZMy5_2(.din(w_dff_B_20jGAzNF7_2),.dout(w_dff_B_dH5f8ZMy5_2),.clk(gclk));
	jdff dff_B_92asM1Ah7_2(.din(w_dff_B_dH5f8ZMy5_2),.dout(w_dff_B_92asM1Ah7_2),.clk(gclk));
	jdff dff_B_nRLOAZKs0_2(.din(w_dff_B_92asM1Ah7_2),.dout(w_dff_B_nRLOAZKs0_2),.clk(gclk));
	jdff dff_B_2Mjul4hS6_2(.din(w_dff_B_nRLOAZKs0_2),.dout(w_dff_B_2Mjul4hS6_2),.clk(gclk));
	jdff dff_B_OUHK7XmR8_2(.din(w_dff_B_2Mjul4hS6_2),.dout(w_dff_B_OUHK7XmR8_2),.clk(gclk));
	jdff dff_B_QLKb3DCw2_2(.din(w_dff_B_OUHK7XmR8_2),.dout(w_dff_B_QLKb3DCw2_2),.clk(gclk));
	jdff dff_B_kbi6UYoJ0_2(.din(w_dff_B_QLKb3DCw2_2),.dout(w_dff_B_kbi6UYoJ0_2),.clk(gclk));
	jdff dff_B_W9BWA3aT2_2(.din(w_dff_B_kbi6UYoJ0_2),.dout(w_dff_B_W9BWA3aT2_2),.clk(gclk));
	jdff dff_B_p8H4l33e3_2(.din(w_dff_B_W9BWA3aT2_2),.dout(w_dff_B_p8H4l33e3_2),.clk(gclk));
	jdff dff_B_DhC8iWBV8_2(.din(w_dff_B_p8H4l33e3_2),.dout(w_dff_B_DhC8iWBV8_2),.clk(gclk));
	jdff dff_B_MHEttRoN0_2(.din(w_dff_B_DhC8iWBV8_2),.dout(w_dff_B_MHEttRoN0_2),.clk(gclk));
	jdff dff_B_YjRiMxhe4_2(.din(w_dff_B_MHEttRoN0_2),.dout(w_dff_B_YjRiMxhe4_2),.clk(gclk));
	jdff dff_B_kpnditTe6_2(.din(w_dff_B_YjRiMxhe4_2),.dout(w_dff_B_kpnditTe6_2),.clk(gclk));
	jdff dff_B_eN0tyKXH9_2(.din(w_dff_B_kpnditTe6_2),.dout(w_dff_B_eN0tyKXH9_2),.clk(gclk));
	jdff dff_B_p2tJ8tsJ5_2(.din(w_dff_B_eN0tyKXH9_2),.dout(w_dff_B_p2tJ8tsJ5_2),.clk(gclk));
	jdff dff_B_5AH076gK6_2(.din(w_dff_B_p2tJ8tsJ5_2),.dout(w_dff_B_5AH076gK6_2),.clk(gclk));
	jdff dff_B_Bf1i3PuS7_2(.din(w_dff_B_5AH076gK6_2),.dout(w_dff_B_Bf1i3PuS7_2),.clk(gclk));
	jdff dff_B_6y5Is34i5_2(.din(w_dff_B_Bf1i3PuS7_2),.dout(w_dff_B_6y5Is34i5_2),.clk(gclk));
	jdff dff_B_2NieMKZc8_2(.din(w_dff_B_6y5Is34i5_2),.dout(w_dff_B_2NieMKZc8_2),.clk(gclk));
	jdff dff_B_VUAU0JZs5_2(.din(w_dff_B_2NieMKZc8_2),.dout(w_dff_B_VUAU0JZs5_2),.clk(gclk));
	jdff dff_B_NBxWaCyk3_2(.din(w_dff_B_VUAU0JZs5_2),.dout(w_dff_B_NBxWaCyk3_2),.clk(gclk));
	jdff dff_B_fsZIy8ab7_2(.din(w_dff_B_NBxWaCyk3_2),.dout(w_dff_B_fsZIy8ab7_2),.clk(gclk));
	jdff dff_B_Lk7lfpJo0_2(.din(w_dff_B_fsZIy8ab7_2),.dout(w_dff_B_Lk7lfpJo0_2),.clk(gclk));
	jdff dff_B_9Ia7o4WF4_2(.din(w_dff_B_Lk7lfpJo0_2),.dout(w_dff_B_9Ia7o4WF4_2),.clk(gclk));
	jdff dff_B_xK3sLJvh1_2(.din(n1135),.dout(w_dff_B_xK3sLJvh1_2),.clk(gclk));
	jdff dff_B_ReanFiuq9_1(.din(n1050),.dout(w_dff_B_ReanFiuq9_1),.clk(gclk));
	jdff dff_B_kd5W7eq48_2(.din(n951),.dout(w_dff_B_kd5W7eq48_2),.clk(gclk));
	jdff dff_B_bSqiJIAL2_2(.din(w_dff_B_kd5W7eq48_2),.dout(w_dff_B_bSqiJIAL2_2),.clk(gclk));
	jdff dff_B_s9AVR4QJ7_2(.din(w_dff_B_bSqiJIAL2_2),.dout(w_dff_B_s9AVR4QJ7_2),.clk(gclk));
	jdff dff_B_uOvxAZgz8_2(.din(w_dff_B_s9AVR4QJ7_2),.dout(w_dff_B_uOvxAZgz8_2),.clk(gclk));
	jdff dff_B_yCNIsvPl7_2(.din(w_dff_B_uOvxAZgz8_2),.dout(w_dff_B_yCNIsvPl7_2),.clk(gclk));
	jdff dff_B_4gRAYFMp6_2(.din(w_dff_B_yCNIsvPl7_2),.dout(w_dff_B_4gRAYFMp6_2),.clk(gclk));
	jdff dff_B_1HFBDYUU6_2(.din(w_dff_B_4gRAYFMp6_2),.dout(w_dff_B_1HFBDYUU6_2),.clk(gclk));
	jdff dff_B_p5h5Y9lv0_2(.din(w_dff_B_1HFBDYUU6_2),.dout(w_dff_B_p5h5Y9lv0_2),.clk(gclk));
	jdff dff_B_n8BAi0lj0_2(.din(w_dff_B_p5h5Y9lv0_2),.dout(w_dff_B_n8BAi0lj0_2),.clk(gclk));
	jdff dff_B_IZZl6UlQ7_2(.din(w_dff_B_n8BAi0lj0_2),.dout(w_dff_B_IZZl6UlQ7_2),.clk(gclk));
	jdff dff_B_TtO1xaW49_2(.din(w_dff_B_IZZl6UlQ7_2),.dout(w_dff_B_TtO1xaW49_2),.clk(gclk));
	jdff dff_B_L92VncoI1_2(.din(w_dff_B_TtO1xaW49_2),.dout(w_dff_B_L92VncoI1_2),.clk(gclk));
	jdff dff_B_knM46jCd4_2(.din(w_dff_B_L92VncoI1_2),.dout(w_dff_B_knM46jCd4_2),.clk(gclk));
	jdff dff_B_k9r9QfiP1_2(.din(w_dff_B_knM46jCd4_2),.dout(w_dff_B_k9r9QfiP1_2),.clk(gclk));
	jdff dff_B_i9B2Xl7L9_2(.din(w_dff_B_k9r9QfiP1_2),.dout(w_dff_B_i9B2Xl7L9_2),.clk(gclk));
	jdff dff_B_077RMbcc9_2(.din(w_dff_B_i9B2Xl7L9_2),.dout(w_dff_B_077RMbcc9_2),.clk(gclk));
	jdff dff_B_z9sBgvdy8_2(.din(w_dff_B_077RMbcc9_2),.dout(w_dff_B_z9sBgvdy8_2),.clk(gclk));
	jdff dff_B_jVRchJe06_2(.din(w_dff_B_z9sBgvdy8_2),.dout(w_dff_B_jVRchJe06_2),.clk(gclk));
	jdff dff_B_ZMeHh2362_2(.din(w_dff_B_jVRchJe06_2),.dout(w_dff_B_ZMeHh2362_2),.clk(gclk));
	jdff dff_B_0vpAugcX0_2(.din(w_dff_B_ZMeHh2362_2),.dout(w_dff_B_0vpAugcX0_2),.clk(gclk));
	jdff dff_B_RlEOiPQl5_2(.din(w_dff_B_0vpAugcX0_2),.dout(w_dff_B_RlEOiPQl5_2),.clk(gclk));
	jdff dff_B_JJxAOLQ72_2(.din(w_dff_B_RlEOiPQl5_2),.dout(w_dff_B_JJxAOLQ72_2),.clk(gclk));
	jdff dff_B_VflyZQf91_2(.din(w_dff_B_JJxAOLQ72_2),.dout(w_dff_B_VflyZQf91_2),.clk(gclk));
	jdff dff_B_3GwdQ9y38_2(.din(w_dff_B_VflyZQf91_2),.dout(w_dff_B_3GwdQ9y38_2),.clk(gclk));
	jdff dff_B_NYtYSTII0_2(.din(w_dff_B_3GwdQ9y38_2),.dout(w_dff_B_NYtYSTII0_2),.clk(gclk));
	jdff dff_B_A2GR43w15_2(.din(w_dff_B_NYtYSTII0_2),.dout(w_dff_B_A2GR43w15_2),.clk(gclk));
	jdff dff_B_bh7xWzCl8_2(.din(w_dff_B_A2GR43w15_2),.dout(w_dff_B_bh7xWzCl8_2),.clk(gclk));
	jdff dff_B_rV1Cd45P9_2(.din(w_dff_B_bh7xWzCl8_2),.dout(w_dff_B_rV1Cd45P9_2),.clk(gclk));
	jdff dff_B_FPPMKExE6_2(.din(w_dff_B_rV1Cd45P9_2),.dout(w_dff_B_FPPMKExE6_2),.clk(gclk));
	jdff dff_B_M8ZdatmK8_2(.din(w_dff_B_FPPMKExE6_2),.dout(w_dff_B_M8ZdatmK8_2),.clk(gclk));
	jdff dff_B_FqWQonU96_2(.din(w_dff_B_M8ZdatmK8_2),.dout(w_dff_B_FqWQonU96_2),.clk(gclk));
	jdff dff_B_PakFZR2O0_2(.din(w_dff_B_FqWQonU96_2),.dout(w_dff_B_PakFZR2O0_2),.clk(gclk));
	jdff dff_B_mkgt8N1q3_2(.din(w_dff_B_PakFZR2O0_2),.dout(w_dff_B_mkgt8N1q3_2),.clk(gclk));
	jdff dff_B_tJknHRp68_2(.din(w_dff_B_mkgt8N1q3_2),.dout(w_dff_B_tJknHRp68_2),.clk(gclk));
	jdff dff_B_yzHuByxt2_2(.din(w_dff_B_tJknHRp68_2),.dout(w_dff_B_yzHuByxt2_2),.clk(gclk));
	jdff dff_B_7ojqKWlw1_2(.din(w_dff_B_yzHuByxt2_2),.dout(w_dff_B_7ojqKWlw1_2),.clk(gclk));
	jdff dff_B_NQ7tOS5e6_2(.din(w_dff_B_7ojqKWlw1_2),.dout(w_dff_B_NQ7tOS5e6_2),.clk(gclk));
	jdff dff_B_7fn1wqLK1_2(.din(n1030),.dout(w_dff_B_7fn1wqLK1_2),.clk(gclk));
	jdff dff_B_veTUZf680_1(.din(n952),.dout(w_dff_B_veTUZf680_1),.clk(gclk));
	jdff dff_B_1MFlNQlG1_2(.din(n846),.dout(w_dff_B_1MFlNQlG1_2),.clk(gclk));
	jdff dff_B_0eN4ZT366_2(.din(w_dff_B_1MFlNQlG1_2),.dout(w_dff_B_0eN4ZT366_2),.clk(gclk));
	jdff dff_B_4ojSBjCe6_2(.din(w_dff_B_0eN4ZT366_2),.dout(w_dff_B_4ojSBjCe6_2),.clk(gclk));
	jdff dff_B_zo6D3ETH3_2(.din(w_dff_B_4ojSBjCe6_2),.dout(w_dff_B_zo6D3ETH3_2),.clk(gclk));
	jdff dff_B_KruONTMx9_2(.din(w_dff_B_zo6D3ETH3_2),.dout(w_dff_B_KruONTMx9_2),.clk(gclk));
	jdff dff_B_o0qIjMcI0_2(.din(w_dff_B_KruONTMx9_2),.dout(w_dff_B_o0qIjMcI0_2),.clk(gclk));
	jdff dff_B_WiooH75D1_2(.din(w_dff_B_o0qIjMcI0_2),.dout(w_dff_B_WiooH75D1_2),.clk(gclk));
	jdff dff_B_J5bK2PNU9_2(.din(w_dff_B_WiooH75D1_2),.dout(w_dff_B_J5bK2PNU9_2),.clk(gclk));
	jdff dff_B_8mZNg4Bt8_2(.din(w_dff_B_J5bK2PNU9_2),.dout(w_dff_B_8mZNg4Bt8_2),.clk(gclk));
	jdff dff_B_sPXgLBGy4_2(.din(w_dff_B_8mZNg4Bt8_2),.dout(w_dff_B_sPXgLBGy4_2),.clk(gclk));
	jdff dff_B_RljsrN7P1_2(.din(w_dff_B_sPXgLBGy4_2),.dout(w_dff_B_RljsrN7P1_2),.clk(gclk));
	jdff dff_B_4kslgDHs2_2(.din(w_dff_B_RljsrN7P1_2),.dout(w_dff_B_4kslgDHs2_2),.clk(gclk));
	jdff dff_B_iL4uqpSt0_2(.din(w_dff_B_4kslgDHs2_2),.dout(w_dff_B_iL4uqpSt0_2),.clk(gclk));
	jdff dff_B_lSTVk3zs6_2(.din(w_dff_B_iL4uqpSt0_2),.dout(w_dff_B_lSTVk3zs6_2),.clk(gclk));
	jdff dff_B_bndFLteT9_2(.din(w_dff_B_lSTVk3zs6_2),.dout(w_dff_B_bndFLteT9_2),.clk(gclk));
	jdff dff_B_XFXya9ej0_2(.din(w_dff_B_bndFLteT9_2),.dout(w_dff_B_XFXya9ej0_2),.clk(gclk));
	jdff dff_B_7UGjaJmc3_2(.din(w_dff_B_XFXya9ej0_2),.dout(w_dff_B_7UGjaJmc3_2),.clk(gclk));
	jdff dff_B_NyH3w9a65_2(.din(w_dff_B_7UGjaJmc3_2),.dout(w_dff_B_NyH3w9a65_2),.clk(gclk));
	jdff dff_B_Cfij2J5D3_2(.din(w_dff_B_NyH3w9a65_2),.dout(w_dff_B_Cfij2J5D3_2),.clk(gclk));
	jdff dff_B_hxt3pRNb1_2(.din(w_dff_B_Cfij2J5D3_2),.dout(w_dff_B_hxt3pRNb1_2),.clk(gclk));
	jdff dff_B_iZ9qV8Xy0_2(.din(w_dff_B_hxt3pRNb1_2),.dout(w_dff_B_iZ9qV8Xy0_2),.clk(gclk));
	jdff dff_B_lRQXa5jr7_2(.din(w_dff_B_iZ9qV8Xy0_2),.dout(w_dff_B_lRQXa5jr7_2),.clk(gclk));
	jdff dff_B_Mp2o1zNl5_2(.din(w_dff_B_lRQXa5jr7_2),.dout(w_dff_B_Mp2o1zNl5_2),.clk(gclk));
	jdff dff_B_oRPwrnrs1_2(.din(w_dff_B_Mp2o1zNl5_2),.dout(w_dff_B_oRPwrnrs1_2),.clk(gclk));
	jdff dff_B_SNSed7v20_2(.din(w_dff_B_oRPwrnrs1_2),.dout(w_dff_B_SNSed7v20_2),.clk(gclk));
	jdff dff_B_ilCQwkt75_2(.din(w_dff_B_SNSed7v20_2),.dout(w_dff_B_ilCQwkt75_2),.clk(gclk));
	jdff dff_B_rdJAEZub9_2(.din(w_dff_B_ilCQwkt75_2),.dout(w_dff_B_rdJAEZub9_2),.clk(gclk));
	jdff dff_B_SOy1ZkQG2_2(.din(w_dff_B_rdJAEZub9_2),.dout(w_dff_B_SOy1ZkQG2_2),.clk(gclk));
	jdff dff_B_Ucw9Lnho8_2(.din(w_dff_B_SOy1ZkQG2_2),.dout(w_dff_B_Ucw9Lnho8_2),.clk(gclk));
	jdff dff_B_xpm8tpan2_2(.din(w_dff_B_Ucw9Lnho8_2),.dout(w_dff_B_xpm8tpan2_2),.clk(gclk));
	jdff dff_B_bbJOOXCc6_2(.din(w_dff_B_xpm8tpan2_2),.dout(w_dff_B_bbJOOXCc6_2),.clk(gclk));
	jdff dff_B_qHtDA7VN9_2(.din(w_dff_B_bbJOOXCc6_2),.dout(w_dff_B_qHtDA7VN9_2),.clk(gclk));
	jdff dff_B_j4Sgkr0I9_2(.din(w_dff_B_qHtDA7VN9_2),.dout(w_dff_B_j4Sgkr0I9_2),.clk(gclk));
	jdff dff_B_oW3OI4Cm9_2(.din(w_dff_B_j4Sgkr0I9_2),.dout(w_dff_B_oW3OI4Cm9_2),.clk(gclk));
	jdff dff_B_k1sYNB9t6_2(.din(n925),.dout(w_dff_B_k1sYNB9t6_2),.clk(gclk));
	jdff dff_B_zMMYx8m05_1(.din(n847),.dout(w_dff_B_zMMYx8m05_1),.clk(gclk));
	jdff dff_B_hLjqSoFN7_2(.din(n747),.dout(w_dff_B_hLjqSoFN7_2),.clk(gclk));
	jdff dff_B_APoPfVjO3_2(.din(w_dff_B_hLjqSoFN7_2),.dout(w_dff_B_APoPfVjO3_2),.clk(gclk));
	jdff dff_B_Bra40SYJ4_2(.din(w_dff_B_APoPfVjO3_2),.dout(w_dff_B_Bra40SYJ4_2),.clk(gclk));
	jdff dff_B_uHVFLnpZ9_2(.din(w_dff_B_Bra40SYJ4_2),.dout(w_dff_B_uHVFLnpZ9_2),.clk(gclk));
	jdff dff_B_JYAUm4iW2_2(.din(w_dff_B_uHVFLnpZ9_2),.dout(w_dff_B_JYAUm4iW2_2),.clk(gclk));
	jdff dff_B_LCVNXzDv4_2(.din(w_dff_B_JYAUm4iW2_2),.dout(w_dff_B_LCVNXzDv4_2),.clk(gclk));
	jdff dff_B_kjKg7emo8_2(.din(w_dff_B_LCVNXzDv4_2),.dout(w_dff_B_kjKg7emo8_2),.clk(gclk));
	jdff dff_B_51pMvQNO7_2(.din(w_dff_B_kjKg7emo8_2),.dout(w_dff_B_51pMvQNO7_2),.clk(gclk));
	jdff dff_B_jd3hHe7a2_2(.din(w_dff_B_51pMvQNO7_2),.dout(w_dff_B_jd3hHe7a2_2),.clk(gclk));
	jdff dff_B_ggBOShHj9_2(.din(w_dff_B_jd3hHe7a2_2),.dout(w_dff_B_ggBOShHj9_2),.clk(gclk));
	jdff dff_B_HwbKrmSb1_2(.din(w_dff_B_ggBOShHj9_2),.dout(w_dff_B_HwbKrmSb1_2),.clk(gclk));
	jdff dff_B_EET26NwP6_2(.din(w_dff_B_HwbKrmSb1_2),.dout(w_dff_B_EET26NwP6_2),.clk(gclk));
	jdff dff_B_bgYwDUoa3_2(.din(w_dff_B_EET26NwP6_2),.dout(w_dff_B_bgYwDUoa3_2),.clk(gclk));
	jdff dff_B_ELpMcuE14_2(.din(w_dff_B_bgYwDUoa3_2),.dout(w_dff_B_ELpMcuE14_2),.clk(gclk));
	jdff dff_B_KcuxWioZ5_2(.din(w_dff_B_ELpMcuE14_2),.dout(w_dff_B_KcuxWioZ5_2),.clk(gclk));
	jdff dff_B_0dGhzTqP6_2(.din(w_dff_B_KcuxWioZ5_2),.dout(w_dff_B_0dGhzTqP6_2),.clk(gclk));
	jdff dff_B_7ghHuPuN3_2(.din(w_dff_B_0dGhzTqP6_2),.dout(w_dff_B_7ghHuPuN3_2),.clk(gclk));
	jdff dff_B_ebQO4LoM7_2(.din(w_dff_B_7ghHuPuN3_2),.dout(w_dff_B_ebQO4LoM7_2),.clk(gclk));
	jdff dff_B_o0GDCZ3h2_2(.din(w_dff_B_ebQO4LoM7_2),.dout(w_dff_B_o0GDCZ3h2_2),.clk(gclk));
	jdff dff_B_xDjETYky4_2(.din(w_dff_B_o0GDCZ3h2_2),.dout(w_dff_B_xDjETYky4_2),.clk(gclk));
	jdff dff_B_AsUrr5bl6_2(.din(w_dff_B_xDjETYky4_2),.dout(w_dff_B_AsUrr5bl6_2),.clk(gclk));
	jdff dff_B_NqiSNVvD0_2(.din(w_dff_B_AsUrr5bl6_2),.dout(w_dff_B_NqiSNVvD0_2),.clk(gclk));
	jdff dff_B_9x5qZPpR0_2(.din(w_dff_B_NqiSNVvD0_2),.dout(w_dff_B_9x5qZPpR0_2),.clk(gclk));
	jdff dff_B_Pu9DKG484_2(.din(w_dff_B_9x5qZPpR0_2),.dout(w_dff_B_Pu9DKG484_2),.clk(gclk));
	jdff dff_B_8LSz4q5N1_2(.din(w_dff_B_Pu9DKG484_2),.dout(w_dff_B_8LSz4q5N1_2),.clk(gclk));
	jdff dff_B_uHWOdmql1_2(.din(w_dff_B_8LSz4q5N1_2),.dout(w_dff_B_uHWOdmql1_2),.clk(gclk));
	jdff dff_B_mlwlzIqc9_2(.din(w_dff_B_uHWOdmql1_2),.dout(w_dff_B_mlwlzIqc9_2),.clk(gclk));
	jdff dff_B_w0kTrk9X0_2(.din(w_dff_B_mlwlzIqc9_2),.dout(w_dff_B_w0kTrk9X0_2),.clk(gclk));
	jdff dff_B_GtifgqIH0_2(.din(w_dff_B_w0kTrk9X0_2),.dout(w_dff_B_GtifgqIH0_2),.clk(gclk));
	jdff dff_B_9lXJlrPk0_2(.din(w_dff_B_GtifgqIH0_2),.dout(w_dff_B_9lXJlrPk0_2),.clk(gclk));
	jdff dff_B_MZeffkU02_2(.din(w_dff_B_9lXJlrPk0_2),.dout(w_dff_B_MZeffkU02_2),.clk(gclk));
	jdff dff_B_NrvwmNJd9_2(.din(n819),.dout(w_dff_B_NrvwmNJd9_2),.clk(gclk));
	jdff dff_B_HCj8WZ5M8_1(.din(n748),.dout(w_dff_B_HCj8WZ5M8_1),.clk(gclk));
	jdff dff_B_1nUfeMI19_2(.din(n654),.dout(w_dff_B_1nUfeMI19_2),.clk(gclk));
	jdff dff_B_r4TgFsLg4_2(.din(w_dff_B_1nUfeMI19_2),.dout(w_dff_B_r4TgFsLg4_2),.clk(gclk));
	jdff dff_B_U7eK7ras0_2(.din(w_dff_B_r4TgFsLg4_2),.dout(w_dff_B_U7eK7ras0_2),.clk(gclk));
	jdff dff_B_zrvC81M98_2(.din(w_dff_B_U7eK7ras0_2),.dout(w_dff_B_zrvC81M98_2),.clk(gclk));
	jdff dff_B_27TquYjo6_2(.din(w_dff_B_zrvC81M98_2),.dout(w_dff_B_27TquYjo6_2),.clk(gclk));
	jdff dff_B_TRzeehci4_2(.din(w_dff_B_27TquYjo6_2),.dout(w_dff_B_TRzeehci4_2),.clk(gclk));
	jdff dff_B_FADVWIPW6_2(.din(w_dff_B_TRzeehci4_2),.dout(w_dff_B_FADVWIPW6_2),.clk(gclk));
	jdff dff_B_owwTMn0U6_2(.din(w_dff_B_FADVWIPW6_2),.dout(w_dff_B_owwTMn0U6_2),.clk(gclk));
	jdff dff_B_6k6UJhV44_2(.din(w_dff_B_owwTMn0U6_2),.dout(w_dff_B_6k6UJhV44_2),.clk(gclk));
	jdff dff_B_wf9KYBtm9_2(.din(w_dff_B_6k6UJhV44_2),.dout(w_dff_B_wf9KYBtm9_2),.clk(gclk));
	jdff dff_B_dpSXt6cN0_2(.din(w_dff_B_wf9KYBtm9_2),.dout(w_dff_B_dpSXt6cN0_2),.clk(gclk));
	jdff dff_B_WmjDN2X53_2(.din(w_dff_B_dpSXt6cN0_2),.dout(w_dff_B_WmjDN2X53_2),.clk(gclk));
	jdff dff_B_9rOUK7gv4_2(.din(w_dff_B_WmjDN2X53_2),.dout(w_dff_B_9rOUK7gv4_2),.clk(gclk));
	jdff dff_B_0ntmxdeh9_2(.din(w_dff_B_9rOUK7gv4_2),.dout(w_dff_B_0ntmxdeh9_2),.clk(gclk));
	jdff dff_B_IYb19NAp3_2(.din(w_dff_B_0ntmxdeh9_2),.dout(w_dff_B_IYb19NAp3_2),.clk(gclk));
	jdff dff_B_BNwk8ty04_2(.din(w_dff_B_IYb19NAp3_2),.dout(w_dff_B_BNwk8ty04_2),.clk(gclk));
	jdff dff_B_SVIbwp204_2(.din(w_dff_B_BNwk8ty04_2),.dout(w_dff_B_SVIbwp204_2),.clk(gclk));
	jdff dff_B_7TVy182l6_2(.din(w_dff_B_SVIbwp204_2),.dout(w_dff_B_7TVy182l6_2),.clk(gclk));
	jdff dff_B_BdpKSbg85_2(.din(w_dff_B_7TVy182l6_2),.dout(w_dff_B_BdpKSbg85_2),.clk(gclk));
	jdff dff_B_3E69npys3_2(.din(w_dff_B_BdpKSbg85_2),.dout(w_dff_B_3E69npys3_2),.clk(gclk));
	jdff dff_B_gUBw3JOx5_2(.din(w_dff_B_3E69npys3_2),.dout(w_dff_B_gUBw3JOx5_2),.clk(gclk));
	jdff dff_B_pQ6i6UA62_2(.din(w_dff_B_gUBw3JOx5_2),.dout(w_dff_B_pQ6i6UA62_2),.clk(gclk));
	jdff dff_B_OcfXnWdd8_2(.din(w_dff_B_pQ6i6UA62_2),.dout(w_dff_B_OcfXnWdd8_2),.clk(gclk));
	jdff dff_B_VJgSELb14_2(.din(w_dff_B_OcfXnWdd8_2),.dout(w_dff_B_VJgSELb14_2),.clk(gclk));
	jdff dff_B_67gh5KcN0_2(.din(w_dff_B_VJgSELb14_2),.dout(w_dff_B_67gh5KcN0_2),.clk(gclk));
	jdff dff_B_NrHTQXjL7_2(.din(w_dff_B_67gh5KcN0_2),.dout(w_dff_B_NrHTQXjL7_2),.clk(gclk));
	jdff dff_B_UzLe5UKv6_2(.din(w_dff_B_NrHTQXjL7_2),.dout(w_dff_B_UzLe5UKv6_2),.clk(gclk));
	jdff dff_B_za3ROloz1_2(.din(w_dff_B_UzLe5UKv6_2),.dout(w_dff_B_za3ROloz1_2),.clk(gclk));
	jdff dff_B_fkjO06sJ2_2(.din(n719),.dout(w_dff_B_fkjO06sJ2_2),.clk(gclk));
	jdff dff_B_oNQaC9jL0_1(.din(n655),.dout(w_dff_B_oNQaC9jL0_1),.clk(gclk));
	jdff dff_B_JhXoKu6z7_2(.din(n568),.dout(w_dff_B_JhXoKu6z7_2),.clk(gclk));
	jdff dff_B_Cch5dsic8_2(.din(w_dff_B_JhXoKu6z7_2),.dout(w_dff_B_Cch5dsic8_2),.clk(gclk));
	jdff dff_B_LFIHne1m0_2(.din(w_dff_B_Cch5dsic8_2),.dout(w_dff_B_LFIHne1m0_2),.clk(gclk));
	jdff dff_B_u9d8O3ND9_2(.din(w_dff_B_LFIHne1m0_2),.dout(w_dff_B_u9d8O3ND9_2),.clk(gclk));
	jdff dff_B_Ov5TIUFx9_2(.din(w_dff_B_u9d8O3ND9_2),.dout(w_dff_B_Ov5TIUFx9_2),.clk(gclk));
	jdff dff_B_RqyCoBIX2_2(.din(w_dff_B_Ov5TIUFx9_2),.dout(w_dff_B_RqyCoBIX2_2),.clk(gclk));
	jdff dff_B_OFcUnF6F3_2(.din(w_dff_B_RqyCoBIX2_2),.dout(w_dff_B_OFcUnF6F3_2),.clk(gclk));
	jdff dff_B_0zouLgnG1_2(.din(w_dff_B_OFcUnF6F3_2),.dout(w_dff_B_0zouLgnG1_2),.clk(gclk));
	jdff dff_B_toc16hBi5_2(.din(w_dff_B_0zouLgnG1_2),.dout(w_dff_B_toc16hBi5_2),.clk(gclk));
	jdff dff_B_TXI1F9mV5_2(.din(w_dff_B_toc16hBi5_2),.dout(w_dff_B_TXI1F9mV5_2),.clk(gclk));
	jdff dff_B_btvoys767_2(.din(w_dff_B_TXI1F9mV5_2),.dout(w_dff_B_btvoys767_2),.clk(gclk));
	jdff dff_B_ubAH73YH1_2(.din(w_dff_B_btvoys767_2),.dout(w_dff_B_ubAH73YH1_2),.clk(gclk));
	jdff dff_B_WKnDMv1C8_2(.din(w_dff_B_ubAH73YH1_2),.dout(w_dff_B_WKnDMv1C8_2),.clk(gclk));
	jdff dff_B_WbdYm6aS0_2(.din(w_dff_B_WKnDMv1C8_2),.dout(w_dff_B_WbdYm6aS0_2),.clk(gclk));
	jdff dff_B_CPeD9D6j4_2(.din(w_dff_B_WbdYm6aS0_2),.dout(w_dff_B_CPeD9D6j4_2),.clk(gclk));
	jdff dff_B_OkSrRGy12_2(.din(w_dff_B_CPeD9D6j4_2),.dout(w_dff_B_OkSrRGy12_2),.clk(gclk));
	jdff dff_B_RUrXO1uE5_2(.din(w_dff_B_OkSrRGy12_2),.dout(w_dff_B_RUrXO1uE5_2),.clk(gclk));
	jdff dff_B_OpurLFzk8_2(.din(w_dff_B_RUrXO1uE5_2),.dout(w_dff_B_OpurLFzk8_2),.clk(gclk));
	jdff dff_B_6k1b1P5b2_2(.din(w_dff_B_OpurLFzk8_2),.dout(w_dff_B_6k1b1P5b2_2),.clk(gclk));
	jdff dff_B_qcQUQ9rg3_2(.din(w_dff_B_6k1b1P5b2_2),.dout(w_dff_B_qcQUQ9rg3_2),.clk(gclk));
	jdff dff_B_4Cjcde9o2_2(.din(w_dff_B_qcQUQ9rg3_2),.dout(w_dff_B_4Cjcde9o2_2),.clk(gclk));
	jdff dff_B_OyySodQ52_2(.din(w_dff_B_4Cjcde9o2_2),.dout(w_dff_B_OyySodQ52_2),.clk(gclk));
	jdff dff_B_Ni0jIFDv4_2(.din(w_dff_B_OyySodQ52_2),.dout(w_dff_B_Ni0jIFDv4_2),.clk(gclk));
	jdff dff_B_jtDwDZT59_2(.din(w_dff_B_Ni0jIFDv4_2),.dout(w_dff_B_jtDwDZT59_2),.clk(gclk));
	jdff dff_B_w04eOjon8_2(.din(w_dff_B_jtDwDZT59_2),.dout(w_dff_B_w04eOjon8_2),.clk(gclk));
	jdff dff_B_TPz8dDkP1_2(.din(n626),.dout(w_dff_B_TPz8dDkP1_2),.clk(gclk));
	jdff dff_B_T5RspWwv6_1(.din(n569),.dout(w_dff_B_T5RspWwv6_1),.clk(gclk));
	jdff dff_B_fSNe4Gi35_2(.din(n489),.dout(w_dff_B_fSNe4Gi35_2),.clk(gclk));
	jdff dff_B_MGVDY3nQ9_2(.din(w_dff_B_fSNe4Gi35_2),.dout(w_dff_B_MGVDY3nQ9_2),.clk(gclk));
	jdff dff_B_LKhWCFMS9_2(.din(w_dff_B_MGVDY3nQ9_2),.dout(w_dff_B_LKhWCFMS9_2),.clk(gclk));
	jdff dff_B_JvBHsJIQ3_2(.din(w_dff_B_LKhWCFMS9_2),.dout(w_dff_B_JvBHsJIQ3_2),.clk(gclk));
	jdff dff_B_os76MLwk6_2(.din(w_dff_B_JvBHsJIQ3_2),.dout(w_dff_B_os76MLwk6_2),.clk(gclk));
	jdff dff_B_tUa7eqWR4_2(.din(w_dff_B_os76MLwk6_2),.dout(w_dff_B_tUa7eqWR4_2),.clk(gclk));
	jdff dff_B_R9yK3csS1_2(.din(w_dff_B_tUa7eqWR4_2),.dout(w_dff_B_R9yK3csS1_2),.clk(gclk));
	jdff dff_B_eqDiBzSp9_2(.din(w_dff_B_R9yK3csS1_2),.dout(w_dff_B_eqDiBzSp9_2),.clk(gclk));
	jdff dff_B_XwtrnRCF6_2(.din(w_dff_B_eqDiBzSp9_2),.dout(w_dff_B_XwtrnRCF6_2),.clk(gclk));
	jdff dff_B_hsqfgo138_2(.din(w_dff_B_XwtrnRCF6_2),.dout(w_dff_B_hsqfgo138_2),.clk(gclk));
	jdff dff_B_lkSsZcwb9_2(.din(w_dff_B_hsqfgo138_2),.dout(w_dff_B_lkSsZcwb9_2),.clk(gclk));
	jdff dff_B_fYJXpoVy8_2(.din(w_dff_B_lkSsZcwb9_2),.dout(w_dff_B_fYJXpoVy8_2),.clk(gclk));
	jdff dff_B_8kgu35s13_2(.din(w_dff_B_fYJXpoVy8_2),.dout(w_dff_B_8kgu35s13_2),.clk(gclk));
	jdff dff_B_AWLHZFl22_2(.din(w_dff_B_8kgu35s13_2),.dout(w_dff_B_AWLHZFl22_2),.clk(gclk));
	jdff dff_B_NNc4Skoq2_2(.din(w_dff_B_AWLHZFl22_2),.dout(w_dff_B_NNc4Skoq2_2),.clk(gclk));
	jdff dff_B_UnMGkXVj1_2(.din(w_dff_B_NNc4Skoq2_2),.dout(w_dff_B_UnMGkXVj1_2),.clk(gclk));
	jdff dff_B_Oa8tzeVT3_2(.din(w_dff_B_UnMGkXVj1_2),.dout(w_dff_B_Oa8tzeVT3_2),.clk(gclk));
	jdff dff_B_y4oUdMDz2_2(.din(w_dff_B_Oa8tzeVT3_2),.dout(w_dff_B_y4oUdMDz2_2),.clk(gclk));
	jdff dff_B_j68deaQ98_2(.din(w_dff_B_y4oUdMDz2_2),.dout(w_dff_B_j68deaQ98_2),.clk(gclk));
	jdff dff_B_mBouTcgA7_2(.din(w_dff_B_j68deaQ98_2),.dout(w_dff_B_mBouTcgA7_2),.clk(gclk));
	jdff dff_B_HU2a7Mqb4_2(.din(w_dff_B_mBouTcgA7_2),.dout(w_dff_B_HU2a7Mqb4_2),.clk(gclk));
	jdff dff_B_lXtCB2Gg5_2(.din(w_dff_B_HU2a7Mqb4_2),.dout(w_dff_B_lXtCB2Gg5_2),.clk(gclk));
	jdff dff_B_y0jHMrmq7_2(.din(n540),.dout(w_dff_B_y0jHMrmq7_2),.clk(gclk));
	jdff dff_B_o0IytErQ1_1(.din(n490),.dout(w_dff_B_o0IytErQ1_1),.clk(gclk));
	jdff dff_B_ucXkrZDx5_2(.din(n417),.dout(w_dff_B_ucXkrZDx5_2),.clk(gclk));
	jdff dff_B_ydJOXd4d9_2(.din(w_dff_B_ucXkrZDx5_2),.dout(w_dff_B_ydJOXd4d9_2),.clk(gclk));
	jdff dff_B_LWpnIXHO7_2(.din(w_dff_B_ydJOXd4d9_2),.dout(w_dff_B_LWpnIXHO7_2),.clk(gclk));
	jdff dff_B_Bcbw6A0V4_2(.din(w_dff_B_LWpnIXHO7_2),.dout(w_dff_B_Bcbw6A0V4_2),.clk(gclk));
	jdff dff_B_qoT6i7rj0_2(.din(w_dff_B_Bcbw6A0V4_2),.dout(w_dff_B_qoT6i7rj0_2),.clk(gclk));
	jdff dff_B_LDqagPD31_2(.din(w_dff_B_qoT6i7rj0_2),.dout(w_dff_B_LDqagPD31_2),.clk(gclk));
	jdff dff_B_WAjYjVyj0_2(.din(w_dff_B_LDqagPD31_2),.dout(w_dff_B_WAjYjVyj0_2),.clk(gclk));
	jdff dff_B_C9xGoUl13_2(.din(w_dff_B_WAjYjVyj0_2),.dout(w_dff_B_C9xGoUl13_2),.clk(gclk));
	jdff dff_B_qmBgromb0_2(.din(w_dff_B_C9xGoUl13_2),.dout(w_dff_B_qmBgromb0_2),.clk(gclk));
	jdff dff_B_PYnyeRYe8_2(.din(w_dff_B_qmBgromb0_2),.dout(w_dff_B_PYnyeRYe8_2),.clk(gclk));
	jdff dff_B_F3Z9RT8L7_2(.din(w_dff_B_PYnyeRYe8_2),.dout(w_dff_B_F3Z9RT8L7_2),.clk(gclk));
	jdff dff_B_9LT574Eg5_2(.din(w_dff_B_F3Z9RT8L7_2),.dout(w_dff_B_9LT574Eg5_2),.clk(gclk));
	jdff dff_B_y8MtH8ep3_2(.din(w_dff_B_9LT574Eg5_2),.dout(w_dff_B_y8MtH8ep3_2),.clk(gclk));
	jdff dff_B_7NlvxpPL2_2(.din(w_dff_B_y8MtH8ep3_2),.dout(w_dff_B_7NlvxpPL2_2),.clk(gclk));
	jdff dff_B_XPNeS3VR2_2(.din(w_dff_B_7NlvxpPL2_2),.dout(w_dff_B_XPNeS3VR2_2),.clk(gclk));
	jdff dff_B_wEMM3LnP6_2(.din(w_dff_B_XPNeS3VR2_2),.dout(w_dff_B_wEMM3LnP6_2),.clk(gclk));
	jdff dff_B_YWnGqG0v9_2(.din(w_dff_B_wEMM3LnP6_2),.dout(w_dff_B_YWnGqG0v9_2),.clk(gclk));
	jdff dff_B_w8wLh6XU3_2(.din(w_dff_B_YWnGqG0v9_2),.dout(w_dff_B_w8wLh6XU3_2),.clk(gclk));
	jdff dff_B_NH7vxheQ8_2(.din(w_dff_B_w8wLh6XU3_2),.dout(w_dff_B_NH7vxheQ8_2),.clk(gclk));
	jdff dff_B_PUBqbE3j7_2(.din(n461),.dout(w_dff_B_PUBqbE3j7_2),.clk(gclk));
	jdff dff_B_6lk4vICq9_1(.din(n418),.dout(w_dff_B_6lk4vICq9_1),.clk(gclk));
	jdff dff_B_u2ild03L2_2(.din(n353),.dout(w_dff_B_u2ild03L2_2),.clk(gclk));
	jdff dff_B_ZeVZeRrl4_2(.din(w_dff_B_u2ild03L2_2),.dout(w_dff_B_ZeVZeRrl4_2),.clk(gclk));
	jdff dff_B_W4FDz4uA4_2(.din(w_dff_B_ZeVZeRrl4_2),.dout(w_dff_B_W4FDz4uA4_2),.clk(gclk));
	jdff dff_B_STI5qzlE4_2(.din(w_dff_B_W4FDz4uA4_2),.dout(w_dff_B_STI5qzlE4_2),.clk(gclk));
	jdff dff_B_HPYReZu66_2(.din(w_dff_B_STI5qzlE4_2),.dout(w_dff_B_HPYReZu66_2),.clk(gclk));
	jdff dff_B_jdO8fL5H8_2(.din(w_dff_B_HPYReZu66_2),.dout(w_dff_B_jdO8fL5H8_2),.clk(gclk));
	jdff dff_B_fKNculjk0_2(.din(w_dff_B_jdO8fL5H8_2),.dout(w_dff_B_fKNculjk0_2),.clk(gclk));
	jdff dff_B_J7DP4vnD7_2(.din(w_dff_B_fKNculjk0_2),.dout(w_dff_B_J7DP4vnD7_2),.clk(gclk));
	jdff dff_B_oUbEnMrs0_2(.din(w_dff_B_J7DP4vnD7_2),.dout(w_dff_B_oUbEnMrs0_2),.clk(gclk));
	jdff dff_B_x8DoXHst6_2(.din(w_dff_B_oUbEnMrs0_2),.dout(w_dff_B_x8DoXHst6_2),.clk(gclk));
	jdff dff_B_7PvO9cLP0_2(.din(w_dff_B_x8DoXHst6_2),.dout(w_dff_B_7PvO9cLP0_2),.clk(gclk));
	jdff dff_B_RPRND2GF9_2(.din(w_dff_B_7PvO9cLP0_2),.dout(w_dff_B_RPRND2GF9_2),.clk(gclk));
	jdff dff_B_JI98W9DV0_2(.din(w_dff_B_RPRND2GF9_2),.dout(w_dff_B_JI98W9DV0_2),.clk(gclk));
	jdff dff_B_wWwjP0kI7_2(.din(w_dff_B_JI98W9DV0_2),.dout(w_dff_B_wWwjP0kI7_2),.clk(gclk));
	jdff dff_B_g8Jwdm8a4_2(.din(w_dff_B_wWwjP0kI7_2),.dout(w_dff_B_g8Jwdm8a4_2),.clk(gclk));
	jdff dff_B_odjSL4HC4_2(.din(w_dff_B_g8Jwdm8a4_2),.dout(w_dff_B_odjSL4HC4_2),.clk(gclk));
	jdff dff_B_CqLjs5BL4_2(.din(n389),.dout(w_dff_B_CqLjs5BL4_2),.clk(gclk));
	jdff dff_B_xT0WLZwq2_1(.din(n354),.dout(w_dff_B_xT0WLZwq2_1),.clk(gclk));
	jdff dff_B_RKKdMgNN3_2(.din(n295),.dout(w_dff_B_RKKdMgNN3_2),.clk(gclk));
	jdff dff_B_0DpLjLmY6_2(.din(w_dff_B_RKKdMgNN3_2),.dout(w_dff_B_0DpLjLmY6_2),.clk(gclk));
	jdff dff_B_v29ksKNL0_2(.din(w_dff_B_0DpLjLmY6_2),.dout(w_dff_B_v29ksKNL0_2),.clk(gclk));
	jdff dff_B_G98R3u7e8_2(.din(w_dff_B_v29ksKNL0_2),.dout(w_dff_B_G98R3u7e8_2),.clk(gclk));
	jdff dff_B_gXyykDV45_2(.din(w_dff_B_G98R3u7e8_2),.dout(w_dff_B_gXyykDV45_2),.clk(gclk));
	jdff dff_B_oCySopo13_2(.din(w_dff_B_gXyykDV45_2),.dout(w_dff_B_oCySopo13_2),.clk(gclk));
	jdff dff_B_BdqtUJ2l9_2(.din(w_dff_B_oCySopo13_2),.dout(w_dff_B_BdqtUJ2l9_2),.clk(gclk));
	jdff dff_B_tT89ZdvF9_2(.din(w_dff_B_BdqtUJ2l9_2),.dout(w_dff_B_tT89ZdvF9_2),.clk(gclk));
	jdff dff_B_3oAWeIJS4_2(.din(w_dff_B_tT89ZdvF9_2),.dout(w_dff_B_3oAWeIJS4_2),.clk(gclk));
	jdff dff_B_AQuR4vss1_2(.din(w_dff_B_3oAWeIJS4_2),.dout(w_dff_B_AQuR4vss1_2),.clk(gclk));
	jdff dff_B_hBQ9ltan8_2(.din(w_dff_B_AQuR4vss1_2),.dout(w_dff_B_hBQ9ltan8_2),.clk(gclk));
	jdff dff_B_vYU6pmby5_2(.din(w_dff_B_hBQ9ltan8_2),.dout(w_dff_B_vYU6pmby5_2),.clk(gclk));
	jdff dff_B_zfj2YvDS8_2(.din(w_dff_B_vYU6pmby5_2),.dout(w_dff_B_zfj2YvDS8_2),.clk(gclk));
	jdff dff_B_nj6Se62c5_2(.din(n325),.dout(w_dff_B_nj6Se62c5_2),.clk(gclk));
	jdff dff_B_TaolNwSg5_1(.din(n296),.dout(w_dff_B_TaolNwSg5_1),.clk(gclk));
	jdff dff_B_XOMwYQ1g5_2(.din(n244),.dout(w_dff_B_XOMwYQ1g5_2),.clk(gclk));
	jdff dff_B_RjhhO5uD1_2(.din(w_dff_B_XOMwYQ1g5_2),.dout(w_dff_B_RjhhO5uD1_2),.clk(gclk));
	jdff dff_B_aOsYWP852_2(.din(w_dff_B_RjhhO5uD1_2),.dout(w_dff_B_aOsYWP852_2),.clk(gclk));
	jdff dff_B_faJLiB5J2_2(.din(w_dff_B_aOsYWP852_2),.dout(w_dff_B_faJLiB5J2_2),.clk(gclk));
	jdff dff_B_GLqZUqOV1_2(.din(w_dff_B_faJLiB5J2_2),.dout(w_dff_B_GLqZUqOV1_2),.clk(gclk));
	jdff dff_B_XGMTY2iG4_2(.din(w_dff_B_GLqZUqOV1_2),.dout(w_dff_B_XGMTY2iG4_2),.clk(gclk));
	jdff dff_B_cT7NVXqe5_2(.din(w_dff_B_XGMTY2iG4_2),.dout(w_dff_B_cT7NVXqe5_2),.clk(gclk));
	jdff dff_B_5TKpctYA4_2(.din(w_dff_B_cT7NVXqe5_2),.dout(w_dff_B_5TKpctYA4_2),.clk(gclk));
	jdff dff_B_VsouEbG68_2(.din(w_dff_B_5TKpctYA4_2),.dout(w_dff_B_VsouEbG68_2),.clk(gclk));
	jdff dff_B_kXxIFRYn3_2(.din(w_dff_B_VsouEbG68_2),.dout(w_dff_B_kXxIFRYn3_2),.clk(gclk));
	jdff dff_B_LhM19GdE6_2(.din(n267),.dout(w_dff_B_LhM19GdE6_2),.clk(gclk));
	jdff dff_B_63xYh7mI9_1(.din(n245),.dout(w_dff_B_63xYh7mI9_1),.clk(gclk));
	jdff dff_B_lUvToWTD5_2(.din(n201),.dout(w_dff_B_lUvToWTD5_2),.clk(gclk));
	jdff dff_B_nT9XyHk90_2(.din(w_dff_B_lUvToWTD5_2),.dout(w_dff_B_nT9XyHk90_2),.clk(gclk));
	jdff dff_B_fAvqAzWA9_2(.din(w_dff_B_nT9XyHk90_2),.dout(w_dff_B_fAvqAzWA9_2),.clk(gclk));
	jdff dff_B_ziFl5Luj2_2(.din(w_dff_B_fAvqAzWA9_2),.dout(w_dff_B_ziFl5Luj2_2),.clk(gclk));
	jdff dff_B_0jAIa8Ra8_2(.din(w_dff_B_ziFl5Luj2_2),.dout(w_dff_B_0jAIa8Ra8_2),.clk(gclk));
	jdff dff_B_nOvOlYwI9_2(.din(w_dff_B_0jAIa8Ra8_2),.dout(w_dff_B_nOvOlYwI9_2),.clk(gclk));
	jdff dff_B_8cqyc2hd9_2(.din(w_dff_B_nOvOlYwI9_2),.dout(w_dff_B_8cqyc2hd9_2),.clk(gclk));
	jdff dff_B_NuTfgCbl3_2(.din(n216),.dout(w_dff_B_NuTfgCbl3_2),.clk(gclk));
	jdff dff_B_840c3GDk4_1(.din(n202),.dout(w_dff_B_840c3GDk4_1),.clk(gclk));
	jdff dff_B_y5d7qXEA7_0(.din(n173),.dout(w_dff_B_y5d7qXEA7_0),.clk(gclk));
	jdff dff_B_MvKZ4hK44_2(.din(n165),.dout(w_dff_B_MvKZ4hK44_2),.clk(gclk));
	jdff dff_B_i0AiXt3t0_2(.din(w_dff_B_MvKZ4hK44_2),.dout(w_dff_B_i0AiXt3t0_2),.clk(gclk));
	jdff dff_B_bLePfPt96_2(.din(w_dff_B_i0AiXt3t0_2),.dout(w_dff_B_bLePfPt96_2),.clk(gclk));
	jdff dff_B_MwjjekUY8_2(.din(w_dff_B_bLePfPt96_2),.dout(w_dff_B_MwjjekUY8_2),.clk(gclk));
	jdff dff_B_KKHmuLIX0_1(.din(n167),.dout(w_dff_B_KKHmuLIX0_1),.clk(gclk));
	jdff dff_A_8E5w6H2V9_0(.dout(w_n132_0[0]),.din(w_dff_A_8E5w6H2V9_0),.clk(gclk));
	jdff dff_A_kW5i3c4R9_0(.dout(w_dff_A_8E5w6H2V9_0),.din(w_dff_A_kW5i3c4R9_0),.clk(gclk));
	jdff dff_A_fhzCCFL74_1(.dout(w_n132_0[1]),.din(w_dff_A_fhzCCFL74_1),.clk(gclk));
	jdff dff_B_FYr4FdfB3_1(.din(n1335),.dout(w_dff_B_FYr4FdfB3_1),.clk(gclk));
	jdff dff_B_97dahFt13_2(.din(n1248),.dout(w_dff_B_97dahFt13_2),.clk(gclk));
	jdff dff_B_kM2w0pJj4_2(.din(w_dff_B_97dahFt13_2),.dout(w_dff_B_kM2w0pJj4_2),.clk(gclk));
	jdff dff_B_sdvDUFMH0_2(.din(w_dff_B_kM2w0pJj4_2),.dout(w_dff_B_sdvDUFMH0_2),.clk(gclk));
	jdff dff_B_ye70Y0S27_2(.din(w_dff_B_sdvDUFMH0_2),.dout(w_dff_B_ye70Y0S27_2),.clk(gclk));
	jdff dff_B_tOA5M8gj2_2(.din(w_dff_B_ye70Y0S27_2),.dout(w_dff_B_tOA5M8gj2_2),.clk(gclk));
	jdff dff_B_canzLa4y0_2(.din(w_dff_B_tOA5M8gj2_2),.dout(w_dff_B_canzLa4y0_2),.clk(gclk));
	jdff dff_B_z2WiqUud6_2(.din(w_dff_B_canzLa4y0_2),.dout(w_dff_B_z2WiqUud6_2),.clk(gclk));
	jdff dff_B_wb7ixjfM7_2(.din(w_dff_B_z2WiqUud6_2),.dout(w_dff_B_wb7ixjfM7_2),.clk(gclk));
	jdff dff_B_KOEcrsUM2_2(.din(w_dff_B_wb7ixjfM7_2),.dout(w_dff_B_KOEcrsUM2_2),.clk(gclk));
	jdff dff_B_eZqMxb2o3_2(.din(w_dff_B_KOEcrsUM2_2),.dout(w_dff_B_eZqMxb2o3_2),.clk(gclk));
	jdff dff_B_lxWqMd960_2(.din(w_dff_B_eZqMxb2o3_2),.dout(w_dff_B_lxWqMd960_2),.clk(gclk));
	jdff dff_B_Vzi2AMkV3_2(.din(w_dff_B_lxWqMd960_2),.dout(w_dff_B_Vzi2AMkV3_2),.clk(gclk));
	jdff dff_B_yjBAKb3p0_2(.din(w_dff_B_Vzi2AMkV3_2),.dout(w_dff_B_yjBAKb3p0_2),.clk(gclk));
	jdff dff_B_1QmP0zAE6_2(.din(w_dff_B_yjBAKb3p0_2),.dout(w_dff_B_1QmP0zAE6_2),.clk(gclk));
	jdff dff_B_Clfefpkr0_2(.din(w_dff_B_1QmP0zAE6_2),.dout(w_dff_B_Clfefpkr0_2),.clk(gclk));
	jdff dff_B_wvS48xXe8_2(.din(w_dff_B_Clfefpkr0_2),.dout(w_dff_B_wvS48xXe8_2),.clk(gclk));
	jdff dff_B_FMFdajSE8_2(.din(w_dff_B_wvS48xXe8_2),.dout(w_dff_B_FMFdajSE8_2),.clk(gclk));
	jdff dff_B_F0U9BQuG0_2(.din(w_dff_B_FMFdajSE8_2),.dout(w_dff_B_F0U9BQuG0_2),.clk(gclk));
	jdff dff_B_jp4O6DnO3_2(.din(w_dff_B_F0U9BQuG0_2),.dout(w_dff_B_jp4O6DnO3_2),.clk(gclk));
	jdff dff_B_NpJKpymw5_2(.din(w_dff_B_jp4O6DnO3_2),.dout(w_dff_B_NpJKpymw5_2),.clk(gclk));
	jdff dff_B_NWlGvxaR1_2(.din(w_dff_B_NpJKpymw5_2),.dout(w_dff_B_NWlGvxaR1_2),.clk(gclk));
	jdff dff_B_BRLxfiIB6_2(.din(w_dff_B_NWlGvxaR1_2),.dout(w_dff_B_BRLxfiIB6_2),.clk(gclk));
	jdff dff_B_Xnznz3Hc7_2(.din(w_dff_B_BRLxfiIB6_2),.dout(w_dff_B_Xnznz3Hc7_2),.clk(gclk));
	jdff dff_B_IkTFQmgJ4_2(.din(w_dff_B_Xnznz3Hc7_2),.dout(w_dff_B_IkTFQmgJ4_2),.clk(gclk));
	jdff dff_B_xfdBIZhg2_2(.din(w_dff_B_IkTFQmgJ4_2),.dout(w_dff_B_xfdBIZhg2_2),.clk(gclk));
	jdff dff_B_zHvjn4iN1_2(.din(w_dff_B_xfdBIZhg2_2),.dout(w_dff_B_zHvjn4iN1_2),.clk(gclk));
	jdff dff_B_Vsu5ghWg6_2(.din(w_dff_B_zHvjn4iN1_2),.dout(w_dff_B_Vsu5ghWg6_2),.clk(gclk));
	jdff dff_B_daI5tDWJ4_2(.din(w_dff_B_Vsu5ghWg6_2),.dout(w_dff_B_daI5tDWJ4_2),.clk(gclk));
	jdff dff_B_tqj6Turq9_2(.din(w_dff_B_daI5tDWJ4_2),.dout(w_dff_B_tqj6Turq9_2),.clk(gclk));
	jdff dff_B_yWe4buxL1_2(.din(w_dff_B_tqj6Turq9_2),.dout(w_dff_B_yWe4buxL1_2),.clk(gclk));
	jdff dff_B_ojg5zu0o8_2(.din(w_dff_B_yWe4buxL1_2),.dout(w_dff_B_ojg5zu0o8_2),.clk(gclk));
	jdff dff_B_tvYn0OcY7_2(.din(w_dff_B_ojg5zu0o8_2),.dout(w_dff_B_tvYn0OcY7_2),.clk(gclk));
	jdff dff_B_pfHaJ1on5_2(.din(w_dff_B_tvYn0OcY7_2),.dout(w_dff_B_pfHaJ1on5_2),.clk(gclk));
	jdff dff_B_eFlPGGgw9_2(.din(w_dff_B_pfHaJ1on5_2),.dout(w_dff_B_eFlPGGgw9_2),.clk(gclk));
	jdff dff_B_wTqoOGBS9_2(.din(w_dff_B_eFlPGGgw9_2),.dout(w_dff_B_wTqoOGBS9_2),.clk(gclk));
	jdff dff_B_1w1TVNSQ3_2(.din(w_dff_B_wTqoOGBS9_2),.dout(w_dff_B_1w1TVNSQ3_2),.clk(gclk));
	jdff dff_B_SN7CToZX4_2(.din(w_dff_B_1w1TVNSQ3_2),.dout(w_dff_B_SN7CToZX4_2),.clk(gclk));
	jdff dff_B_2azUBcUx4_2(.din(w_dff_B_SN7CToZX4_2),.dout(w_dff_B_2azUBcUx4_2),.clk(gclk));
	jdff dff_B_Uh8vgPYg3_2(.din(w_dff_B_2azUBcUx4_2),.dout(w_dff_B_Uh8vgPYg3_2),.clk(gclk));
	jdff dff_B_UjghNXSM2_2(.din(w_dff_B_Uh8vgPYg3_2),.dout(w_dff_B_UjghNXSM2_2),.clk(gclk));
	jdff dff_B_Vl97vaTn6_2(.din(w_dff_B_UjghNXSM2_2),.dout(w_dff_B_Vl97vaTn6_2),.clk(gclk));
	jdff dff_B_P26eiy1G5_2(.din(w_dff_B_Vl97vaTn6_2),.dout(w_dff_B_P26eiy1G5_2),.clk(gclk));
	jdff dff_B_NO15k2Oc6_2(.din(w_dff_B_P26eiy1G5_2),.dout(w_dff_B_NO15k2Oc6_2),.clk(gclk));
	jdff dff_B_QNpmEh2r7_2(.din(w_dff_B_NO15k2Oc6_2),.dout(w_dff_B_QNpmEh2r7_2),.clk(gclk));
	jdff dff_B_TkXN03tm1_2(.din(w_dff_B_QNpmEh2r7_2),.dout(w_dff_B_TkXN03tm1_2),.clk(gclk));
	jdff dff_B_ErSGtDO89_0(.din(n1334),.dout(w_dff_B_ErSGtDO89_0),.clk(gclk));
	jdff dff_A_kYtAJoyj3_1(.dout(w_n1322_0[1]),.din(w_dff_A_kYtAJoyj3_1),.clk(gclk));
	jdff dff_B_PO12R7st0_1(.din(n1249),.dout(w_dff_B_PO12R7st0_1),.clk(gclk));
	jdff dff_B_G1maRCRW3_2(.din(n1158),.dout(w_dff_B_G1maRCRW3_2),.clk(gclk));
	jdff dff_B_Q64g7U0e7_2(.din(w_dff_B_G1maRCRW3_2),.dout(w_dff_B_Q64g7U0e7_2),.clk(gclk));
	jdff dff_B_UbQ2xhCw9_2(.din(w_dff_B_Q64g7U0e7_2),.dout(w_dff_B_UbQ2xhCw9_2),.clk(gclk));
	jdff dff_B_GchuL2Ck6_2(.din(w_dff_B_UbQ2xhCw9_2),.dout(w_dff_B_GchuL2Ck6_2),.clk(gclk));
	jdff dff_B_Y2h6OELG8_2(.din(w_dff_B_GchuL2Ck6_2),.dout(w_dff_B_Y2h6OELG8_2),.clk(gclk));
	jdff dff_B_SmnIKM9c9_2(.din(w_dff_B_Y2h6OELG8_2),.dout(w_dff_B_SmnIKM9c9_2),.clk(gclk));
	jdff dff_B_T6OUy6Wr5_2(.din(w_dff_B_SmnIKM9c9_2),.dout(w_dff_B_T6OUy6Wr5_2),.clk(gclk));
	jdff dff_B_MAVHHYY07_2(.din(w_dff_B_T6OUy6Wr5_2),.dout(w_dff_B_MAVHHYY07_2),.clk(gclk));
	jdff dff_B_nI5hRsFM4_2(.din(w_dff_B_MAVHHYY07_2),.dout(w_dff_B_nI5hRsFM4_2),.clk(gclk));
	jdff dff_B_VPiU3bUU2_2(.din(w_dff_B_nI5hRsFM4_2),.dout(w_dff_B_VPiU3bUU2_2),.clk(gclk));
	jdff dff_B_VO0rdYS86_2(.din(w_dff_B_VPiU3bUU2_2),.dout(w_dff_B_VO0rdYS86_2),.clk(gclk));
	jdff dff_B_xnIqzth18_2(.din(w_dff_B_VO0rdYS86_2),.dout(w_dff_B_xnIqzth18_2),.clk(gclk));
	jdff dff_B_PHhCAjey3_2(.din(w_dff_B_xnIqzth18_2),.dout(w_dff_B_PHhCAjey3_2),.clk(gclk));
	jdff dff_B_gYLMXeYr0_2(.din(w_dff_B_PHhCAjey3_2),.dout(w_dff_B_gYLMXeYr0_2),.clk(gclk));
	jdff dff_B_sfVftEcX5_2(.din(w_dff_B_gYLMXeYr0_2),.dout(w_dff_B_sfVftEcX5_2),.clk(gclk));
	jdff dff_B_iHWmKDPY2_2(.din(w_dff_B_sfVftEcX5_2),.dout(w_dff_B_iHWmKDPY2_2),.clk(gclk));
	jdff dff_B_lWA7B3iK7_2(.din(w_dff_B_iHWmKDPY2_2),.dout(w_dff_B_lWA7B3iK7_2),.clk(gclk));
	jdff dff_B_G23HMgzn4_2(.din(w_dff_B_lWA7B3iK7_2),.dout(w_dff_B_G23HMgzn4_2),.clk(gclk));
	jdff dff_B_ucLvddoU5_2(.din(w_dff_B_G23HMgzn4_2),.dout(w_dff_B_ucLvddoU5_2),.clk(gclk));
	jdff dff_B_nvPwtDLH3_2(.din(w_dff_B_ucLvddoU5_2),.dout(w_dff_B_nvPwtDLH3_2),.clk(gclk));
	jdff dff_B_XMI1GGMD8_2(.din(w_dff_B_nvPwtDLH3_2),.dout(w_dff_B_XMI1GGMD8_2),.clk(gclk));
	jdff dff_B_dj8YkQ9B8_2(.din(w_dff_B_XMI1GGMD8_2),.dout(w_dff_B_dj8YkQ9B8_2),.clk(gclk));
	jdff dff_B_neCjZH8g0_2(.din(w_dff_B_dj8YkQ9B8_2),.dout(w_dff_B_neCjZH8g0_2),.clk(gclk));
	jdff dff_B_mwiq29ZP1_2(.din(w_dff_B_neCjZH8g0_2),.dout(w_dff_B_mwiq29ZP1_2),.clk(gclk));
	jdff dff_B_oWVLYtYp5_2(.din(w_dff_B_mwiq29ZP1_2),.dout(w_dff_B_oWVLYtYp5_2),.clk(gclk));
	jdff dff_B_2ph7WAf20_2(.din(w_dff_B_oWVLYtYp5_2),.dout(w_dff_B_2ph7WAf20_2),.clk(gclk));
	jdff dff_B_To9WhxcV1_2(.din(w_dff_B_2ph7WAf20_2),.dout(w_dff_B_To9WhxcV1_2),.clk(gclk));
	jdff dff_B_xPwgAhsL9_2(.din(w_dff_B_To9WhxcV1_2),.dout(w_dff_B_xPwgAhsL9_2),.clk(gclk));
	jdff dff_B_uXZKAVL43_2(.din(w_dff_B_xPwgAhsL9_2),.dout(w_dff_B_uXZKAVL43_2),.clk(gclk));
	jdff dff_B_nfefX84y6_2(.din(w_dff_B_uXZKAVL43_2),.dout(w_dff_B_nfefX84y6_2),.clk(gclk));
	jdff dff_B_bLHxjmhz6_2(.din(w_dff_B_nfefX84y6_2),.dout(w_dff_B_bLHxjmhz6_2),.clk(gclk));
	jdff dff_B_yBHXCI0G8_2(.din(w_dff_B_bLHxjmhz6_2),.dout(w_dff_B_yBHXCI0G8_2),.clk(gclk));
	jdff dff_B_6Xd9MZD60_2(.din(w_dff_B_yBHXCI0G8_2),.dout(w_dff_B_6Xd9MZD60_2),.clk(gclk));
	jdff dff_B_xHJA97rU7_2(.din(w_dff_B_6Xd9MZD60_2),.dout(w_dff_B_xHJA97rU7_2),.clk(gclk));
	jdff dff_B_O3NERh0V7_2(.din(w_dff_B_xHJA97rU7_2),.dout(w_dff_B_O3NERh0V7_2),.clk(gclk));
	jdff dff_B_VeJfhk6p7_2(.din(w_dff_B_O3NERh0V7_2),.dout(w_dff_B_VeJfhk6p7_2),.clk(gclk));
	jdff dff_B_w5VGHhFp4_2(.din(w_dff_B_VeJfhk6p7_2),.dout(w_dff_B_w5VGHhFp4_2),.clk(gclk));
	jdff dff_B_hcXKlHQ22_2(.din(w_dff_B_w5VGHhFp4_2),.dout(w_dff_B_hcXKlHQ22_2),.clk(gclk));
	jdff dff_B_x3gphihD4_2(.din(w_dff_B_hcXKlHQ22_2),.dout(w_dff_B_x3gphihD4_2),.clk(gclk));
	jdff dff_B_C1CopPj13_2(.din(w_dff_B_x3gphihD4_2),.dout(w_dff_B_C1CopPj13_2),.clk(gclk));
	jdff dff_B_yl0l0a1u5_2(.din(n1231),.dout(w_dff_B_yl0l0a1u5_2),.clk(gclk));
	jdff dff_B_1FdTulTQ5_1(.din(n1159),.dout(w_dff_B_1FdTulTQ5_1),.clk(gclk));
	jdff dff_B_WDUMuBKs2_2(.din(n1054),.dout(w_dff_B_WDUMuBKs2_2),.clk(gclk));
	jdff dff_B_tHPoC6bH8_2(.din(w_dff_B_WDUMuBKs2_2),.dout(w_dff_B_tHPoC6bH8_2),.clk(gclk));
	jdff dff_B_iuPXHBei1_2(.din(w_dff_B_tHPoC6bH8_2),.dout(w_dff_B_iuPXHBei1_2),.clk(gclk));
	jdff dff_B_wOLEZ0023_2(.din(w_dff_B_iuPXHBei1_2),.dout(w_dff_B_wOLEZ0023_2),.clk(gclk));
	jdff dff_B_3CbNm7mZ3_2(.din(w_dff_B_wOLEZ0023_2),.dout(w_dff_B_3CbNm7mZ3_2),.clk(gclk));
	jdff dff_B_33K1CaVa9_2(.din(w_dff_B_3CbNm7mZ3_2),.dout(w_dff_B_33K1CaVa9_2),.clk(gclk));
	jdff dff_B_NuYLS1BX4_2(.din(w_dff_B_33K1CaVa9_2),.dout(w_dff_B_NuYLS1BX4_2),.clk(gclk));
	jdff dff_B_NG9JutYO9_2(.din(w_dff_B_NuYLS1BX4_2),.dout(w_dff_B_NG9JutYO9_2),.clk(gclk));
	jdff dff_B_tMct18bU3_2(.din(w_dff_B_NG9JutYO9_2),.dout(w_dff_B_tMct18bU3_2),.clk(gclk));
	jdff dff_B_6ytrvTXf3_2(.din(w_dff_B_tMct18bU3_2),.dout(w_dff_B_6ytrvTXf3_2),.clk(gclk));
	jdff dff_B_J0a2xsRx4_2(.din(w_dff_B_6ytrvTXf3_2),.dout(w_dff_B_J0a2xsRx4_2),.clk(gclk));
	jdff dff_B_qOZOIK6A6_2(.din(w_dff_B_J0a2xsRx4_2),.dout(w_dff_B_qOZOIK6A6_2),.clk(gclk));
	jdff dff_B_FrL6L2WZ9_2(.din(w_dff_B_qOZOIK6A6_2),.dout(w_dff_B_FrL6L2WZ9_2),.clk(gclk));
	jdff dff_B_1Hhp8gWr8_2(.din(w_dff_B_FrL6L2WZ9_2),.dout(w_dff_B_1Hhp8gWr8_2),.clk(gclk));
	jdff dff_B_wybK3zaP9_2(.din(w_dff_B_1Hhp8gWr8_2),.dout(w_dff_B_wybK3zaP9_2),.clk(gclk));
	jdff dff_B_e4Ywqcf42_2(.din(w_dff_B_wybK3zaP9_2),.dout(w_dff_B_e4Ywqcf42_2),.clk(gclk));
	jdff dff_B_T4vBLDra3_2(.din(w_dff_B_e4Ywqcf42_2),.dout(w_dff_B_T4vBLDra3_2),.clk(gclk));
	jdff dff_B_vVwrYBw38_2(.din(w_dff_B_T4vBLDra3_2),.dout(w_dff_B_vVwrYBw38_2),.clk(gclk));
	jdff dff_B_Bb3YooaZ9_2(.din(w_dff_B_vVwrYBw38_2),.dout(w_dff_B_Bb3YooaZ9_2),.clk(gclk));
	jdff dff_B_J64LuYsM8_2(.din(w_dff_B_Bb3YooaZ9_2),.dout(w_dff_B_J64LuYsM8_2),.clk(gclk));
	jdff dff_B_pcviOWKM5_2(.din(w_dff_B_J64LuYsM8_2),.dout(w_dff_B_pcviOWKM5_2),.clk(gclk));
	jdff dff_B_YSQZGqYA8_2(.din(w_dff_B_pcviOWKM5_2),.dout(w_dff_B_YSQZGqYA8_2),.clk(gclk));
	jdff dff_B_LTyKT05K8_2(.din(w_dff_B_YSQZGqYA8_2),.dout(w_dff_B_LTyKT05K8_2),.clk(gclk));
	jdff dff_B_ZbNZszgQ1_2(.din(w_dff_B_LTyKT05K8_2),.dout(w_dff_B_ZbNZszgQ1_2),.clk(gclk));
	jdff dff_B_xCevtBru7_2(.din(w_dff_B_ZbNZszgQ1_2),.dout(w_dff_B_xCevtBru7_2),.clk(gclk));
	jdff dff_B_Z1Yh5kcX9_2(.din(w_dff_B_xCevtBru7_2),.dout(w_dff_B_Z1Yh5kcX9_2),.clk(gclk));
	jdff dff_B_zYtxJ5f01_2(.din(w_dff_B_Z1Yh5kcX9_2),.dout(w_dff_B_zYtxJ5f01_2),.clk(gclk));
	jdff dff_B_pSBAOqev4_2(.din(w_dff_B_zYtxJ5f01_2),.dout(w_dff_B_pSBAOqev4_2),.clk(gclk));
	jdff dff_B_qjoQU56g2_2(.din(w_dff_B_pSBAOqev4_2),.dout(w_dff_B_qjoQU56g2_2),.clk(gclk));
	jdff dff_B_doZPJe446_2(.din(w_dff_B_qjoQU56g2_2),.dout(w_dff_B_doZPJe446_2),.clk(gclk));
	jdff dff_B_fBFLnPRJ9_2(.din(w_dff_B_doZPJe446_2),.dout(w_dff_B_fBFLnPRJ9_2),.clk(gclk));
	jdff dff_B_R8Mu0ulb9_2(.din(w_dff_B_fBFLnPRJ9_2),.dout(w_dff_B_R8Mu0ulb9_2),.clk(gclk));
	jdff dff_B_xcIS3Db01_2(.din(w_dff_B_R8Mu0ulb9_2),.dout(w_dff_B_xcIS3Db01_2),.clk(gclk));
	jdff dff_B_LDj1WWAe8_2(.din(w_dff_B_xcIS3Db01_2),.dout(w_dff_B_LDj1WWAe8_2),.clk(gclk));
	jdff dff_B_eQ3WmxFV6_2(.din(w_dff_B_LDj1WWAe8_2),.dout(w_dff_B_eQ3WmxFV6_2),.clk(gclk));
	jdff dff_B_50d97sJh9_2(.din(w_dff_B_eQ3WmxFV6_2),.dout(w_dff_B_50d97sJh9_2),.clk(gclk));
	jdff dff_B_SPEl12Do8_2(.din(w_dff_B_50d97sJh9_2),.dout(w_dff_B_SPEl12Do8_2),.clk(gclk));
	jdff dff_B_dwHvenCd1_2(.din(n1133),.dout(w_dff_B_dwHvenCd1_2),.clk(gclk));
	jdff dff_B_e7fGPhgE3_1(.din(n1055),.dout(w_dff_B_e7fGPhgE3_1),.clk(gclk));
	jdff dff_B_LmsiQImZ3_2(.din(n956),.dout(w_dff_B_LmsiQImZ3_2),.clk(gclk));
	jdff dff_B_8CLIK6zu7_2(.din(w_dff_B_LmsiQImZ3_2),.dout(w_dff_B_8CLIK6zu7_2),.clk(gclk));
	jdff dff_B_4bWhRPM23_2(.din(w_dff_B_8CLIK6zu7_2),.dout(w_dff_B_4bWhRPM23_2),.clk(gclk));
	jdff dff_B_6YuIOJ1G8_2(.din(w_dff_B_4bWhRPM23_2),.dout(w_dff_B_6YuIOJ1G8_2),.clk(gclk));
	jdff dff_B_OuAbxXVj7_2(.din(w_dff_B_6YuIOJ1G8_2),.dout(w_dff_B_OuAbxXVj7_2),.clk(gclk));
	jdff dff_B_rTGNjhvs5_2(.din(w_dff_B_OuAbxXVj7_2),.dout(w_dff_B_rTGNjhvs5_2),.clk(gclk));
	jdff dff_B_IzYZFxIU4_2(.din(w_dff_B_rTGNjhvs5_2),.dout(w_dff_B_IzYZFxIU4_2),.clk(gclk));
	jdff dff_B_1h37I6P49_2(.din(w_dff_B_IzYZFxIU4_2),.dout(w_dff_B_1h37I6P49_2),.clk(gclk));
	jdff dff_B_b7RuuJtX6_2(.din(w_dff_B_1h37I6P49_2),.dout(w_dff_B_b7RuuJtX6_2),.clk(gclk));
	jdff dff_B_rq5qyBfF8_2(.din(w_dff_B_b7RuuJtX6_2),.dout(w_dff_B_rq5qyBfF8_2),.clk(gclk));
	jdff dff_B_WNWLDnI84_2(.din(w_dff_B_rq5qyBfF8_2),.dout(w_dff_B_WNWLDnI84_2),.clk(gclk));
	jdff dff_B_cO8QrZAa1_2(.din(w_dff_B_WNWLDnI84_2),.dout(w_dff_B_cO8QrZAa1_2),.clk(gclk));
	jdff dff_B_msLjvfIU6_2(.din(w_dff_B_cO8QrZAa1_2),.dout(w_dff_B_msLjvfIU6_2),.clk(gclk));
	jdff dff_B_MGLBF5eC1_2(.din(w_dff_B_msLjvfIU6_2),.dout(w_dff_B_MGLBF5eC1_2),.clk(gclk));
	jdff dff_B_lDkGGy7K7_2(.din(w_dff_B_MGLBF5eC1_2),.dout(w_dff_B_lDkGGy7K7_2),.clk(gclk));
	jdff dff_B_TeVGVNDj4_2(.din(w_dff_B_lDkGGy7K7_2),.dout(w_dff_B_TeVGVNDj4_2),.clk(gclk));
	jdff dff_B_cwoCL9eg1_2(.din(w_dff_B_TeVGVNDj4_2),.dout(w_dff_B_cwoCL9eg1_2),.clk(gclk));
	jdff dff_B_GQukG6X37_2(.din(w_dff_B_cwoCL9eg1_2),.dout(w_dff_B_GQukG6X37_2),.clk(gclk));
	jdff dff_B_J239FyPX1_2(.din(w_dff_B_GQukG6X37_2),.dout(w_dff_B_J239FyPX1_2),.clk(gclk));
	jdff dff_B_sA8k7kSF3_2(.din(w_dff_B_J239FyPX1_2),.dout(w_dff_B_sA8k7kSF3_2),.clk(gclk));
	jdff dff_B_RDMpURB99_2(.din(w_dff_B_sA8k7kSF3_2),.dout(w_dff_B_RDMpURB99_2),.clk(gclk));
	jdff dff_B_5iE0CbGz1_2(.din(w_dff_B_RDMpURB99_2),.dout(w_dff_B_5iE0CbGz1_2),.clk(gclk));
	jdff dff_B_PX3zf5Gz8_2(.din(w_dff_B_5iE0CbGz1_2),.dout(w_dff_B_PX3zf5Gz8_2),.clk(gclk));
	jdff dff_B_IhNFsn7B3_2(.din(w_dff_B_PX3zf5Gz8_2),.dout(w_dff_B_IhNFsn7B3_2),.clk(gclk));
	jdff dff_B_pORJCIuw4_2(.din(w_dff_B_IhNFsn7B3_2),.dout(w_dff_B_pORJCIuw4_2),.clk(gclk));
	jdff dff_B_wGuVFKaH5_2(.din(w_dff_B_pORJCIuw4_2),.dout(w_dff_B_wGuVFKaH5_2),.clk(gclk));
	jdff dff_B_3uCZmPoo8_2(.din(w_dff_B_wGuVFKaH5_2),.dout(w_dff_B_3uCZmPoo8_2),.clk(gclk));
	jdff dff_B_gPlS9qr43_2(.din(w_dff_B_3uCZmPoo8_2),.dout(w_dff_B_gPlS9qr43_2),.clk(gclk));
	jdff dff_B_ktyEjLTY7_2(.din(w_dff_B_gPlS9qr43_2),.dout(w_dff_B_ktyEjLTY7_2),.clk(gclk));
	jdff dff_B_9CtZTChJ3_2(.din(w_dff_B_ktyEjLTY7_2),.dout(w_dff_B_9CtZTChJ3_2),.clk(gclk));
	jdff dff_B_Fhb1x64I8_2(.din(w_dff_B_9CtZTChJ3_2),.dout(w_dff_B_Fhb1x64I8_2),.clk(gclk));
	jdff dff_B_5hKuInnK9_2(.din(w_dff_B_Fhb1x64I8_2),.dout(w_dff_B_5hKuInnK9_2),.clk(gclk));
	jdff dff_B_hws0KtPy6_2(.din(w_dff_B_5hKuInnK9_2),.dout(w_dff_B_hws0KtPy6_2),.clk(gclk));
	jdff dff_B_65svk5wf5_2(.din(w_dff_B_hws0KtPy6_2),.dout(w_dff_B_65svk5wf5_2),.clk(gclk));
	jdff dff_B_j5PCsBuH8_2(.din(n1028),.dout(w_dff_B_j5PCsBuH8_2),.clk(gclk));
	jdff dff_B_pBI9Lvgg8_1(.din(n957),.dout(w_dff_B_pBI9Lvgg8_1),.clk(gclk));
	jdff dff_B_wzDJ8GCf6_2(.din(n851),.dout(w_dff_B_wzDJ8GCf6_2),.clk(gclk));
	jdff dff_B_OpDI0DFm5_2(.din(w_dff_B_wzDJ8GCf6_2),.dout(w_dff_B_OpDI0DFm5_2),.clk(gclk));
	jdff dff_B_IvLQERmA4_2(.din(w_dff_B_OpDI0DFm5_2),.dout(w_dff_B_IvLQERmA4_2),.clk(gclk));
	jdff dff_B_TOp3wvWf0_2(.din(w_dff_B_IvLQERmA4_2),.dout(w_dff_B_TOp3wvWf0_2),.clk(gclk));
	jdff dff_B_A3nHQHCi0_2(.din(w_dff_B_TOp3wvWf0_2),.dout(w_dff_B_A3nHQHCi0_2),.clk(gclk));
	jdff dff_B_B3ko1R7p6_2(.din(w_dff_B_A3nHQHCi0_2),.dout(w_dff_B_B3ko1R7p6_2),.clk(gclk));
	jdff dff_B_fNYjTCIu3_2(.din(w_dff_B_B3ko1R7p6_2),.dout(w_dff_B_fNYjTCIu3_2),.clk(gclk));
	jdff dff_B_SOwTlDjF2_2(.din(w_dff_B_fNYjTCIu3_2),.dout(w_dff_B_SOwTlDjF2_2),.clk(gclk));
	jdff dff_B_TCvgAghv5_2(.din(w_dff_B_SOwTlDjF2_2),.dout(w_dff_B_TCvgAghv5_2),.clk(gclk));
	jdff dff_B_iyMBxWQQ9_2(.din(w_dff_B_TCvgAghv5_2),.dout(w_dff_B_iyMBxWQQ9_2),.clk(gclk));
	jdff dff_B_D5ACEWdk6_2(.din(w_dff_B_iyMBxWQQ9_2),.dout(w_dff_B_D5ACEWdk6_2),.clk(gclk));
	jdff dff_B_IHkhM8kn8_2(.din(w_dff_B_D5ACEWdk6_2),.dout(w_dff_B_IHkhM8kn8_2),.clk(gclk));
	jdff dff_B_ZhaEjqcn4_2(.din(w_dff_B_IHkhM8kn8_2),.dout(w_dff_B_ZhaEjqcn4_2),.clk(gclk));
	jdff dff_B_8eldP4aa5_2(.din(w_dff_B_ZhaEjqcn4_2),.dout(w_dff_B_8eldP4aa5_2),.clk(gclk));
	jdff dff_B_UAtNCGJR1_2(.din(w_dff_B_8eldP4aa5_2),.dout(w_dff_B_UAtNCGJR1_2),.clk(gclk));
	jdff dff_B_Pb1SEEpV5_2(.din(w_dff_B_UAtNCGJR1_2),.dout(w_dff_B_Pb1SEEpV5_2),.clk(gclk));
	jdff dff_B_VZjmkF8E2_2(.din(w_dff_B_Pb1SEEpV5_2),.dout(w_dff_B_VZjmkF8E2_2),.clk(gclk));
	jdff dff_B_SQ1korkG5_2(.din(w_dff_B_VZjmkF8E2_2),.dout(w_dff_B_SQ1korkG5_2),.clk(gclk));
	jdff dff_B_rKvf5muT9_2(.din(w_dff_B_SQ1korkG5_2),.dout(w_dff_B_rKvf5muT9_2),.clk(gclk));
	jdff dff_B_Zjp6PeYn3_2(.din(w_dff_B_rKvf5muT9_2),.dout(w_dff_B_Zjp6PeYn3_2),.clk(gclk));
	jdff dff_B_8iRFxlKX4_2(.din(w_dff_B_Zjp6PeYn3_2),.dout(w_dff_B_8iRFxlKX4_2),.clk(gclk));
	jdff dff_B_bPyhQSOP4_2(.din(w_dff_B_8iRFxlKX4_2),.dout(w_dff_B_bPyhQSOP4_2),.clk(gclk));
	jdff dff_B_Wtx5tA226_2(.din(w_dff_B_bPyhQSOP4_2),.dout(w_dff_B_Wtx5tA226_2),.clk(gclk));
	jdff dff_B_Vh4MYR6s0_2(.din(w_dff_B_Wtx5tA226_2),.dout(w_dff_B_Vh4MYR6s0_2),.clk(gclk));
	jdff dff_B_UBhSE7YF7_2(.din(w_dff_B_Vh4MYR6s0_2),.dout(w_dff_B_UBhSE7YF7_2),.clk(gclk));
	jdff dff_B_Q9jpslpw3_2(.din(w_dff_B_UBhSE7YF7_2),.dout(w_dff_B_Q9jpslpw3_2),.clk(gclk));
	jdff dff_B_L2o0Hqbn7_2(.din(w_dff_B_Q9jpslpw3_2),.dout(w_dff_B_L2o0Hqbn7_2),.clk(gclk));
	jdff dff_B_8bwieWx31_2(.din(w_dff_B_L2o0Hqbn7_2),.dout(w_dff_B_8bwieWx31_2),.clk(gclk));
	jdff dff_B_lL1GPZWx1_2(.din(w_dff_B_8bwieWx31_2),.dout(w_dff_B_lL1GPZWx1_2),.clk(gclk));
	jdff dff_B_d5zoKY9j2_2(.din(w_dff_B_lL1GPZWx1_2),.dout(w_dff_B_d5zoKY9j2_2),.clk(gclk));
	jdff dff_B_FvJ5VlAH2_2(.din(w_dff_B_d5zoKY9j2_2),.dout(w_dff_B_FvJ5VlAH2_2),.clk(gclk));
	jdff dff_B_r0eWN7pX6_2(.din(n923),.dout(w_dff_B_r0eWN7pX6_2),.clk(gclk));
	jdff dff_B_ts1N6ri07_1(.din(n852),.dout(w_dff_B_ts1N6ri07_1),.clk(gclk));
	jdff dff_B_YqdZnYp53_2(.din(n752),.dout(w_dff_B_YqdZnYp53_2),.clk(gclk));
	jdff dff_B_kmMz4Gf42_2(.din(w_dff_B_YqdZnYp53_2),.dout(w_dff_B_kmMz4Gf42_2),.clk(gclk));
	jdff dff_B_43mAdFk75_2(.din(w_dff_B_kmMz4Gf42_2),.dout(w_dff_B_43mAdFk75_2),.clk(gclk));
	jdff dff_B_6i7Y3gjJ6_2(.din(w_dff_B_43mAdFk75_2),.dout(w_dff_B_6i7Y3gjJ6_2),.clk(gclk));
	jdff dff_B_TPqjHbOt1_2(.din(w_dff_B_6i7Y3gjJ6_2),.dout(w_dff_B_TPqjHbOt1_2),.clk(gclk));
	jdff dff_B_gPv13XMD8_2(.din(w_dff_B_TPqjHbOt1_2),.dout(w_dff_B_gPv13XMD8_2),.clk(gclk));
	jdff dff_B_JDbgwmlQ8_2(.din(w_dff_B_gPv13XMD8_2),.dout(w_dff_B_JDbgwmlQ8_2),.clk(gclk));
	jdff dff_B_nxTYpnUK8_2(.din(w_dff_B_JDbgwmlQ8_2),.dout(w_dff_B_nxTYpnUK8_2),.clk(gclk));
	jdff dff_B_bRG6w92b1_2(.din(w_dff_B_nxTYpnUK8_2),.dout(w_dff_B_bRG6w92b1_2),.clk(gclk));
	jdff dff_B_uullTJNc3_2(.din(w_dff_B_bRG6w92b1_2),.dout(w_dff_B_uullTJNc3_2),.clk(gclk));
	jdff dff_B_Vchd5S709_2(.din(w_dff_B_uullTJNc3_2),.dout(w_dff_B_Vchd5S709_2),.clk(gclk));
	jdff dff_B_lYzj0mSx3_2(.din(w_dff_B_Vchd5S709_2),.dout(w_dff_B_lYzj0mSx3_2),.clk(gclk));
	jdff dff_B_OTVnSV1y4_2(.din(w_dff_B_lYzj0mSx3_2),.dout(w_dff_B_OTVnSV1y4_2),.clk(gclk));
	jdff dff_B_X9qIEM6a7_2(.din(w_dff_B_OTVnSV1y4_2),.dout(w_dff_B_X9qIEM6a7_2),.clk(gclk));
	jdff dff_B_jyz3z9Kz0_2(.din(w_dff_B_X9qIEM6a7_2),.dout(w_dff_B_jyz3z9Kz0_2),.clk(gclk));
	jdff dff_B_Zq7N5mJb5_2(.din(w_dff_B_jyz3z9Kz0_2),.dout(w_dff_B_Zq7N5mJb5_2),.clk(gclk));
	jdff dff_B_VCjJqEBn3_2(.din(w_dff_B_Zq7N5mJb5_2),.dout(w_dff_B_VCjJqEBn3_2),.clk(gclk));
	jdff dff_B_yenbJd053_2(.din(w_dff_B_VCjJqEBn3_2),.dout(w_dff_B_yenbJd053_2),.clk(gclk));
	jdff dff_B_xulcjw5X0_2(.din(w_dff_B_yenbJd053_2),.dout(w_dff_B_xulcjw5X0_2),.clk(gclk));
	jdff dff_B_evc9jos05_2(.din(w_dff_B_xulcjw5X0_2),.dout(w_dff_B_evc9jos05_2),.clk(gclk));
	jdff dff_B_5SfTaJ0x0_2(.din(w_dff_B_evc9jos05_2),.dout(w_dff_B_5SfTaJ0x0_2),.clk(gclk));
	jdff dff_B_QUB7MmDY1_2(.din(w_dff_B_5SfTaJ0x0_2),.dout(w_dff_B_QUB7MmDY1_2),.clk(gclk));
	jdff dff_B_aOnfFLsY0_2(.din(w_dff_B_QUB7MmDY1_2),.dout(w_dff_B_aOnfFLsY0_2),.clk(gclk));
	jdff dff_B_WLQ1ZuIR2_2(.din(w_dff_B_aOnfFLsY0_2),.dout(w_dff_B_WLQ1ZuIR2_2),.clk(gclk));
	jdff dff_B_jAPbVsbm7_2(.din(w_dff_B_WLQ1ZuIR2_2),.dout(w_dff_B_jAPbVsbm7_2),.clk(gclk));
	jdff dff_B_E0p2adVD9_2(.din(w_dff_B_jAPbVsbm7_2),.dout(w_dff_B_E0p2adVD9_2),.clk(gclk));
	jdff dff_B_ZNy59xiD0_2(.din(w_dff_B_E0p2adVD9_2),.dout(w_dff_B_ZNy59xiD0_2),.clk(gclk));
	jdff dff_B_vREFlxaq6_2(.din(w_dff_B_ZNy59xiD0_2),.dout(w_dff_B_vREFlxaq6_2),.clk(gclk));
	jdff dff_B_6ugO9nhT4_2(.din(n817),.dout(w_dff_B_6ugO9nhT4_2),.clk(gclk));
	jdff dff_B_ScF5DwwC9_1(.din(n753),.dout(w_dff_B_ScF5DwwC9_1),.clk(gclk));
	jdff dff_B_PvOC5jrK0_2(.din(n659),.dout(w_dff_B_PvOC5jrK0_2),.clk(gclk));
	jdff dff_B_4tPRFRgg6_2(.din(w_dff_B_PvOC5jrK0_2),.dout(w_dff_B_4tPRFRgg6_2),.clk(gclk));
	jdff dff_B_kudyrlO27_2(.din(w_dff_B_4tPRFRgg6_2),.dout(w_dff_B_kudyrlO27_2),.clk(gclk));
	jdff dff_B_qfalpslK9_2(.din(w_dff_B_kudyrlO27_2),.dout(w_dff_B_qfalpslK9_2),.clk(gclk));
	jdff dff_B_V3HQj16c1_2(.din(w_dff_B_qfalpslK9_2),.dout(w_dff_B_V3HQj16c1_2),.clk(gclk));
	jdff dff_B_QDyQD9Zb0_2(.din(w_dff_B_V3HQj16c1_2),.dout(w_dff_B_QDyQD9Zb0_2),.clk(gclk));
	jdff dff_B_DaCLurpc9_2(.din(w_dff_B_QDyQD9Zb0_2),.dout(w_dff_B_DaCLurpc9_2),.clk(gclk));
	jdff dff_B_6QTSgAb25_2(.din(w_dff_B_DaCLurpc9_2),.dout(w_dff_B_6QTSgAb25_2),.clk(gclk));
	jdff dff_B_2euEQrjF8_2(.din(w_dff_B_6QTSgAb25_2),.dout(w_dff_B_2euEQrjF8_2),.clk(gclk));
	jdff dff_B_paSe0hMp1_2(.din(w_dff_B_2euEQrjF8_2),.dout(w_dff_B_paSe0hMp1_2),.clk(gclk));
	jdff dff_B_n5Tgybgr7_2(.din(w_dff_B_paSe0hMp1_2),.dout(w_dff_B_n5Tgybgr7_2),.clk(gclk));
	jdff dff_B_xsJ9fH2c7_2(.din(w_dff_B_n5Tgybgr7_2),.dout(w_dff_B_xsJ9fH2c7_2),.clk(gclk));
	jdff dff_B_oXKF7KbU7_2(.din(w_dff_B_xsJ9fH2c7_2),.dout(w_dff_B_oXKF7KbU7_2),.clk(gclk));
	jdff dff_B_uEedBUuE2_2(.din(w_dff_B_oXKF7KbU7_2),.dout(w_dff_B_uEedBUuE2_2),.clk(gclk));
	jdff dff_B_iKwcjPnB7_2(.din(w_dff_B_uEedBUuE2_2),.dout(w_dff_B_iKwcjPnB7_2),.clk(gclk));
	jdff dff_B_ou0gdfKh1_2(.din(w_dff_B_iKwcjPnB7_2),.dout(w_dff_B_ou0gdfKh1_2),.clk(gclk));
	jdff dff_B_myqiBtY24_2(.din(w_dff_B_ou0gdfKh1_2),.dout(w_dff_B_myqiBtY24_2),.clk(gclk));
	jdff dff_B_SKuD2mDk0_2(.din(w_dff_B_myqiBtY24_2),.dout(w_dff_B_SKuD2mDk0_2),.clk(gclk));
	jdff dff_B_oDNeadf12_2(.din(w_dff_B_SKuD2mDk0_2),.dout(w_dff_B_oDNeadf12_2),.clk(gclk));
	jdff dff_B_IPPejWRp4_2(.din(w_dff_B_oDNeadf12_2),.dout(w_dff_B_IPPejWRp4_2),.clk(gclk));
	jdff dff_B_3TBBLLiv7_2(.din(w_dff_B_IPPejWRp4_2),.dout(w_dff_B_3TBBLLiv7_2),.clk(gclk));
	jdff dff_B_KRrt0mCn7_2(.din(w_dff_B_3TBBLLiv7_2),.dout(w_dff_B_KRrt0mCn7_2),.clk(gclk));
	jdff dff_B_v7HP5egH3_2(.din(w_dff_B_KRrt0mCn7_2),.dout(w_dff_B_v7HP5egH3_2),.clk(gclk));
	jdff dff_B_l2K1yHub2_2(.din(w_dff_B_v7HP5egH3_2),.dout(w_dff_B_l2K1yHub2_2),.clk(gclk));
	jdff dff_B_2n9qfHGe5_2(.din(w_dff_B_l2K1yHub2_2),.dout(w_dff_B_2n9qfHGe5_2),.clk(gclk));
	jdff dff_B_Jf9q3FuV5_2(.din(n717),.dout(w_dff_B_Jf9q3FuV5_2),.clk(gclk));
	jdff dff_B_ambeZDru3_1(.din(n660),.dout(w_dff_B_ambeZDru3_1),.clk(gclk));
	jdff dff_B_pT211enw6_2(.din(n573),.dout(w_dff_B_pT211enw6_2),.clk(gclk));
	jdff dff_B_5RbJpCSr5_2(.din(w_dff_B_pT211enw6_2),.dout(w_dff_B_5RbJpCSr5_2),.clk(gclk));
	jdff dff_B_BnSh8e9n1_2(.din(w_dff_B_5RbJpCSr5_2),.dout(w_dff_B_BnSh8e9n1_2),.clk(gclk));
	jdff dff_B_Oa3AfMKN1_2(.din(w_dff_B_BnSh8e9n1_2),.dout(w_dff_B_Oa3AfMKN1_2),.clk(gclk));
	jdff dff_B_FUq7BMzz2_2(.din(w_dff_B_Oa3AfMKN1_2),.dout(w_dff_B_FUq7BMzz2_2),.clk(gclk));
	jdff dff_B_69ytwXJt8_2(.din(w_dff_B_FUq7BMzz2_2),.dout(w_dff_B_69ytwXJt8_2),.clk(gclk));
	jdff dff_B_kAl9rvsN4_2(.din(w_dff_B_69ytwXJt8_2),.dout(w_dff_B_kAl9rvsN4_2),.clk(gclk));
	jdff dff_B_4ccqOJDd4_2(.din(w_dff_B_kAl9rvsN4_2),.dout(w_dff_B_4ccqOJDd4_2),.clk(gclk));
	jdff dff_B_Shtvuj1w8_2(.din(w_dff_B_4ccqOJDd4_2),.dout(w_dff_B_Shtvuj1w8_2),.clk(gclk));
	jdff dff_B_4irAzCcn9_2(.din(w_dff_B_Shtvuj1w8_2),.dout(w_dff_B_4irAzCcn9_2),.clk(gclk));
	jdff dff_B_cc4iG2Le1_2(.din(w_dff_B_4irAzCcn9_2),.dout(w_dff_B_cc4iG2Le1_2),.clk(gclk));
	jdff dff_B_Acxl081n6_2(.din(w_dff_B_cc4iG2Le1_2),.dout(w_dff_B_Acxl081n6_2),.clk(gclk));
	jdff dff_B_fWheg23y9_2(.din(w_dff_B_Acxl081n6_2),.dout(w_dff_B_fWheg23y9_2),.clk(gclk));
	jdff dff_B_NKNkC2Cm6_2(.din(w_dff_B_fWheg23y9_2),.dout(w_dff_B_NKNkC2Cm6_2),.clk(gclk));
	jdff dff_B_GS2PR2bm7_2(.din(w_dff_B_NKNkC2Cm6_2),.dout(w_dff_B_GS2PR2bm7_2),.clk(gclk));
	jdff dff_B_rV9VqsnX6_2(.din(w_dff_B_GS2PR2bm7_2),.dout(w_dff_B_rV9VqsnX6_2),.clk(gclk));
	jdff dff_B_WGkWsx5q0_2(.din(w_dff_B_rV9VqsnX6_2),.dout(w_dff_B_WGkWsx5q0_2),.clk(gclk));
	jdff dff_B_u1wLJopG9_2(.din(w_dff_B_WGkWsx5q0_2),.dout(w_dff_B_u1wLJopG9_2),.clk(gclk));
	jdff dff_B_MwQPq3qX3_2(.din(w_dff_B_u1wLJopG9_2),.dout(w_dff_B_MwQPq3qX3_2),.clk(gclk));
	jdff dff_B_F2UjT6mZ9_2(.din(w_dff_B_MwQPq3qX3_2),.dout(w_dff_B_F2UjT6mZ9_2),.clk(gclk));
	jdff dff_B_j4WSWt6l8_2(.din(w_dff_B_F2UjT6mZ9_2),.dout(w_dff_B_j4WSWt6l8_2),.clk(gclk));
	jdff dff_B_YtxsDGOU2_2(.din(w_dff_B_j4WSWt6l8_2),.dout(w_dff_B_YtxsDGOU2_2),.clk(gclk));
	jdff dff_B_smBEFrpg5_2(.din(n624),.dout(w_dff_B_smBEFrpg5_2),.clk(gclk));
	jdff dff_B_7S1vnxda9_1(.din(n574),.dout(w_dff_B_7S1vnxda9_1),.clk(gclk));
	jdff dff_B_uWHYvu380_2(.din(n494),.dout(w_dff_B_uWHYvu380_2),.clk(gclk));
	jdff dff_B_LJhkuRgl3_2(.din(w_dff_B_uWHYvu380_2),.dout(w_dff_B_LJhkuRgl3_2),.clk(gclk));
	jdff dff_B_mvKh69Z53_2(.din(w_dff_B_LJhkuRgl3_2),.dout(w_dff_B_mvKh69Z53_2),.clk(gclk));
	jdff dff_B_F6qK8rmi9_2(.din(w_dff_B_mvKh69Z53_2),.dout(w_dff_B_F6qK8rmi9_2),.clk(gclk));
	jdff dff_B_cwclJGCG1_2(.din(w_dff_B_F6qK8rmi9_2),.dout(w_dff_B_cwclJGCG1_2),.clk(gclk));
	jdff dff_B_izOQKGti7_2(.din(w_dff_B_cwclJGCG1_2),.dout(w_dff_B_izOQKGti7_2),.clk(gclk));
	jdff dff_B_FS2E4zBV6_2(.din(w_dff_B_izOQKGti7_2),.dout(w_dff_B_FS2E4zBV6_2),.clk(gclk));
	jdff dff_B_9SNvCuRv9_2(.din(w_dff_B_FS2E4zBV6_2),.dout(w_dff_B_9SNvCuRv9_2),.clk(gclk));
	jdff dff_B_xQyJCR9W3_2(.din(w_dff_B_9SNvCuRv9_2),.dout(w_dff_B_xQyJCR9W3_2),.clk(gclk));
	jdff dff_B_RgON4shO5_2(.din(w_dff_B_xQyJCR9W3_2),.dout(w_dff_B_RgON4shO5_2),.clk(gclk));
	jdff dff_B_XmO9pUmN1_2(.din(w_dff_B_RgON4shO5_2),.dout(w_dff_B_XmO9pUmN1_2),.clk(gclk));
	jdff dff_B_rIKw22Tb8_2(.din(w_dff_B_XmO9pUmN1_2),.dout(w_dff_B_rIKw22Tb8_2),.clk(gclk));
	jdff dff_B_zCITm22H5_2(.din(w_dff_B_rIKw22Tb8_2),.dout(w_dff_B_zCITm22H5_2),.clk(gclk));
	jdff dff_B_u899r1GP3_2(.din(w_dff_B_zCITm22H5_2),.dout(w_dff_B_u899r1GP3_2),.clk(gclk));
	jdff dff_B_UVKIPfSg1_2(.din(w_dff_B_u899r1GP3_2),.dout(w_dff_B_UVKIPfSg1_2),.clk(gclk));
	jdff dff_B_uhNwhAlK3_2(.din(w_dff_B_UVKIPfSg1_2),.dout(w_dff_B_uhNwhAlK3_2),.clk(gclk));
	jdff dff_B_zq1Xb35I2_2(.din(w_dff_B_uhNwhAlK3_2),.dout(w_dff_B_zq1Xb35I2_2),.clk(gclk));
	jdff dff_B_TryxKBJx8_2(.din(w_dff_B_zq1Xb35I2_2),.dout(w_dff_B_TryxKBJx8_2),.clk(gclk));
	jdff dff_B_6D0AnOxI9_2(.din(w_dff_B_TryxKBJx8_2),.dout(w_dff_B_6D0AnOxI9_2),.clk(gclk));
	jdff dff_B_60jCzz1X6_2(.din(n538),.dout(w_dff_B_60jCzz1X6_2),.clk(gclk));
	jdff dff_B_0ub2UGTJ6_1(.din(n495),.dout(w_dff_B_0ub2UGTJ6_1),.clk(gclk));
	jdff dff_B_hZP5Pcea3_2(.din(n422),.dout(w_dff_B_hZP5Pcea3_2),.clk(gclk));
	jdff dff_B_xaF7K1LR1_2(.din(w_dff_B_hZP5Pcea3_2),.dout(w_dff_B_xaF7K1LR1_2),.clk(gclk));
	jdff dff_B_6NBxfdrw1_2(.din(w_dff_B_xaF7K1LR1_2),.dout(w_dff_B_6NBxfdrw1_2),.clk(gclk));
	jdff dff_B_DzFcIKYo9_2(.din(w_dff_B_6NBxfdrw1_2),.dout(w_dff_B_DzFcIKYo9_2),.clk(gclk));
	jdff dff_B_cIXviL1N7_2(.din(w_dff_B_DzFcIKYo9_2),.dout(w_dff_B_cIXviL1N7_2),.clk(gclk));
	jdff dff_B_GKUwsO8n9_2(.din(w_dff_B_cIXviL1N7_2),.dout(w_dff_B_GKUwsO8n9_2),.clk(gclk));
	jdff dff_B_zQ5YPaKt5_2(.din(w_dff_B_GKUwsO8n9_2),.dout(w_dff_B_zQ5YPaKt5_2),.clk(gclk));
	jdff dff_B_A8lGErrZ9_2(.din(w_dff_B_zQ5YPaKt5_2),.dout(w_dff_B_A8lGErrZ9_2),.clk(gclk));
	jdff dff_B_7PCCRPQf4_2(.din(w_dff_B_A8lGErrZ9_2),.dout(w_dff_B_7PCCRPQf4_2),.clk(gclk));
	jdff dff_B_XFS9fUwq4_2(.din(w_dff_B_7PCCRPQf4_2),.dout(w_dff_B_XFS9fUwq4_2),.clk(gclk));
	jdff dff_B_04UenHlJ6_2(.din(w_dff_B_XFS9fUwq4_2),.dout(w_dff_B_04UenHlJ6_2),.clk(gclk));
	jdff dff_B_VJuDTfFt3_2(.din(w_dff_B_04UenHlJ6_2),.dout(w_dff_B_VJuDTfFt3_2),.clk(gclk));
	jdff dff_B_Lh6ghqtr8_2(.din(w_dff_B_VJuDTfFt3_2),.dout(w_dff_B_Lh6ghqtr8_2),.clk(gclk));
	jdff dff_B_BkLOlcoO5_2(.din(w_dff_B_Lh6ghqtr8_2),.dout(w_dff_B_BkLOlcoO5_2),.clk(gclk));
	jdff dff_B_GoYdnHUq3_2(.din(w_dff_B_BkLOlcoO5_2),.dout(w_dff_B_GoYdnHUq3_2),.clk(gclk));
	jdff dff_B_DMYriVf68_2(.din(w_dff_B_GoYdnHUq3_2),.dout(w_dff_B_DMYriVf68_2),.clk(gclk));
	jdff dff_B_99G06CEw4_2(.din(n459),.dout(w_dff_B_99G06CEw4_2),.clk(gclk));
	jdff dff_B_VavVFlVG0_1(.din(n423),.dout(w_dff_B_VavVFlVG0_1),.clk(gclk));
	jdff dff_B_l6lJxTBy4_2(.din(n358),.dout(w_dff_B_l6lJxTBy4_2),.clk(gclk));
	jdff dff_B_Zu9RzIMr3_2(.din(w_dff_B_l6lJxTBy4_2),.dout(w_dff_B_Zu9RzIMr3_2),.clk(gclk));
	jdff dff_B_meauC6jk3_2(.din(w_dff_B_Zu9RzIMr3_2),.dout(w_dff_B_meauC6jk3_2),.clk(gclk));
	jdff dff_B_F4RgRU7D9_2(.din(w_dff_B_meauC6jk3_2),.dout(w_dff_B_F4RgRU7D9_2),.clk(gclk));
	jdff dff_B_XRQJSKkf0_2(.din(w_dff_B_F4RgRU7D9_2),.dout(w_dff_B_XRQJSKkf0_2),.clk(gclk));
	jdff dff_B_bzJFWsZ66_2(.din(w_dff_B_XRQJSKkf0_2),.dout(w_dff_B_bzJFWsZ66_2),.clk(gclk));
	jdff dff_B_2Rga0I6R9_2(.din(w_dff_B_bzJFWsZ66_2),.dout(w_dff_B_2Rga0I6R9_2),.clk(gclk));
	jdff dff_B_Q8fkGh5e6_2(.din(w_dff_B_2Rga0I6R9_2),.dout(w_dff_B_Q8fkGh5e6_2),.clk(gclk));
	jdff dff_B_y92OjV0m5_2(.din(w_dff_B_Q8fkGh5e6_2),.dout(w_dff_B_y92OjV0m5_2),.clk(gclk));
	jdff dff_B_Z2uRmlb57_2(.din(w_dff_B_y92OjV0m5_2),.dout(w_dff_B_Z2uRmlb57_2),.clk(gclk));
	jdff dff_B_ENARae1N1_2(.din(w_dff_B_Z2uRmlb57_2),.dout(w_dff_B_ENARae1N1_2),.clk(gclk));
	jdff dff_B_BW0Xlbkn2_2(.din(w_dff_B_ENARae1N1_2),.dout(w_dff_B_BW0Xlbkn2_2),.clk(gclk));
	jdff dff_B_z3z38aMv1_2(.din(w_dff_B_BW0Xlbkn2_2),.dout(w_dff_B_z3z38aMv1_2),.clk(gclk));
	jdff dff_B_mh08k7Jk4_2(.din(n387),.dout(w_dff_B_mh08k7Jk4_2),.clk(gclk));
	jdff dff_B_wBflJaNu9_1(.din(n359),.dout(w_dff_B_wBflJaNu9_1),.clk(gclk));
	jdff dff_B_Hg4HGYb48_2(.din(n300),.dout(w_dff_B_Hg4HGYb48_2),.clk(gclk));
	jdff dff_B_EGYQy1GI8_2(.din(w_dff_B_Hg4HGYb48_2),.dout(w_dff_B_EGYQy1GI8_2),.clk(gclk));
	jdff dff_B_wtoysNb52_2(.din(w_dff_B_EGYQy1GI8_2),.dout(w_dff_B_wtoysNb52_2),.clk(gclk));
	jdff dff_B_nnmYLzoN4_2(.din(w_dff_B_wtoysNb52_2),.dout(w_dff_B_nnmYLzoN4_2),.clk(gclk));
	jdff dff_B_BgbXiQmy6_2(.din(w_dff_B_nnmYLzoN4_2),.dout(w_dff_B_BgbXiQmy6_2),.clk(gclk));
	jdff dff_B_5DaD8okL6_2(.din(w_dff_B_BgbXiQmy6_2),.dout(w_dff_B_5DaD8okL6_2),.clk(gclk));
	jdff dff_B_1qb0wsjc3_2(.din(w_dff_B_5DaD8okL6_2),.dout(w_dff_B_1qb0wsjc3_2),.clk(gclk));
	jdff dff_B_2OvjnneS9_2(.din(w_dff_B_1qb0wsjc3_2),.dout(w_dff_B_2OvjnneS9_2),.clk(gclk));
	jdff dff_B_MOR0XDjc2_2(.din(w_dff_B_2OvjnneS9_2),.dout(w_dff_B_MOR0XDjc2_2),.clk(gclk));
	jdff dff_B_Fh9L8oXW3_2(.din(w_dff_B_MOR0XDjc2_2),.dout(w_dff_B_Fh9L8oXW3_2),.clk(gclk));
	jdff dff_B_3l4SKcDE9_2(.din(n323),.dout(w_dff_B_3l4SKcDE9_2),.clk(gclk));
	jdff dff_B_4pUskhmR3_1(.din(n301),.dout(w_dff_B_4pUskhmR3_1),.clk(gclk));
	jdff dff_B_Zffz6OVe5_2(.din(n249),.dout(w_dff_B_Zffz6OVe5_2),.clk(gclk));
	jdff dff_B_mqFqbXDs5_2(.din(w_dff_B_Zffz6OVe5_2),.dout(w_dff_B_mqFqbXDs5_2),.clk(gclk));
	jdff dff_B_eDp7MZDI5_2(.din(w_dff_B_mqFqbXDs5_2),.dout(w_dff_B_eDp7MZDI5_2),.clk(gclk));
	jdff dff_B_90Go2Bhy0_2(.din(w_dff_B_eDp7MZDI5_2),.dout(w_dff_B_90Go2Bhy0_2),.clk(gclk));
	jdff dff_B_8ojogRrX5_2(.din(w_dff_B_90Go2Bhy0_2),.dout(w_dff_B_8ojogRrX5_2),.clk(gclk));
	jdff dff_B_i3BNk4I12_2(.din(w_dff_B_8ojogRrX5_2),.dout(w_dff_B_i3BNk4I12_2),.clk(gclk));
	jdff dff_B_NzaK6og78_2(.din(w_dff_B_i3BNk4I12_2),.dout(w_dff_B_NzaK6og78_2),.clk(gclk));
	jdff dff_B_2ZFijG8y4_2(.din(n265),.dout(w_dff_B_2ZFijG8y4_2),.clk(gclk));
	jdff dff_B_KmYDFXAP3_1(.din(n250),.dout(w_dff_B_KmYDFXAP3_1),.clk(gclk));
	jdff dff_B_K5WYOovD9_0(.din(n214),.dout(w_dff_B_K5WYOovD9_0),.clk(gclk));
	jdff dff_B_NYY6r2fA2_2(.din(n206),.dout(w_dff_B_NYY6r2fA2_2),.clk(gclk));
	jdff dff_B_e0vTI1iP1_2(.din(w_dff_B_NYY6r2fA2_2),.dout(w_dff_B_e0vTI1iP1_2),.clk(gclk));
	jdff dff_B_tnEQxkZm4_2(.din(w_dff_B_e0vTI1iP1_2),.dout(w_dff_B_tnEQxkZm4_2),.clk(gclk));
	jdff dff_B_sgCcalFI4_2(.din(w_dff_B_tnEQxkZm4_2),.dout(w_dff_B_sgCcalFI4_2),.clk(gclk));
	jdff dff_B_4EFGqvCf7_1(.din(n208),.dout(w_dff_B_4EFGqvCf7_1),.clk(gclk));
	jdff dff_A_1dikcfgM7_0(.dout(w_n210_1[0]),.din(w_dff_A_1dikcfgM7_0),.clk(gclk));
	jdff dff_A_vdeHAEpJ2_0(.dout(w_n169_0[0]),.din(w_dff_A_vdeHAEpJ2_0),.clk(gclk));
	jdff dff_A_S5jpLcNQ9_0(.dout(w_dff_A_vdeHAEpJ2_0),.din(w_dff_A_S5jpLcNQ9_0),.clk(gclk));
	jdff dff_A_0436c07I2_1(.dout(w_n169_0[1]),.din(w_dff_A_0436c07I2_1),.clk(gclk));
	jdff dff_B_16GkUzZv0_2(.din(n1420),.dout(w_dff_B_16GkUzZv0_2),.clk(gclk));
	jdff dff_B_LlyAvuTl5_1(.din(n1418),.dout(w_dff_B_LlyAvuTl5_1),.clk(gclk));
	jdff dff_B_oEuP862p2_2(.din(n1338),.dout(w_dff_B_oEuP862p2_2),.clk(gclk));
	jdff dff_B_2FCJ6bpK1_2(.din(w_dff_B_oEuP862p2_2),.dout(w_dff_B_2FCJ6bpK1_2),.clk(gclk));
	jdff dff_B_qXX7wsY90_2(.din(w_dff_B_2FCJ6bpK1_2),.dout(w_dff_B_qXX7wsY90_2),.clk(gclk));
	jdff dff_B_MnL8R5MZ8_2(.din(w_dff_B_qXX7wsY90_2),.dout(w_dff_B_MnL8R5MZ8_2),.clk(gclk));
	jdff dff_B_rmY4Ptp70_2(.din(w_dff_B_MnL8R5MZ8_2),.dout(w_dff_B_rmY4Ptp70_2),.clk(gclk));
	jdff dff_B_8ctsjS5W8_2(.din(w_dff_B_rmY4Ptp70_2),.dout(w_dff_B_8ctsjS5W8_2),.clk(gclk));
	jdff dff_B_BoSfgg6J1_2(.din(w_dff_B_8ctsjS5W8_2),.dout(w_dff_B_BoSfgg6J1_2),.clk(gclk));
	jdff dff_B_QdedzU871_2(.din(w_dff_B_BoSfgg6J1_2),.dout(w_dff_B_QdedzU871_2),.clk(gclk));
	jdff dff_B_0UnuHLDC7_2(.din(w_dff_B_QdedzU871_2),.dout(w_dff_B_0UnuHLDC7_2),.clk(gclk));
	jdff dff_B_eNHY3aZ41_2(.din(w_dff_B_0UnuHLDC7_2),.dout(w_dff_B_eNHY3aZ41_2),.clk(gclk));
	jdff dff_B_OYthKwP47_2(.din(w_dff_B_eNHY3aZ41_2),.dout(w_dff_B_OYthKwP47_2),.clk(gclk));
	jdff dff_B_N22Abqi71_2(.din(w_dff_B_OYthKwP47_2),.dout(w_dff_B_N22Abqi71_2),.clk(gclk));
	jdff dff_B_nS1bcpwc5_2(.din(w_dff_B_N22Abqi71_2),.dout(w_dff_B_nS1bcpwc5_2),.clk(gclk));
	jdff dff_B_zVmWG6I28_2(.din(w_dff_B_nS1bcpwc5_2),.dout(w_dff_B_zVmWG6I28_2),.clk(gclk));
	jdff dff_B_aWVtrNGj7_2(.din(w_dff_B_zVmWG6I28_2),.dout(w_dff_B_aWVtrNGj7_2),.clk(gclk));
	jdff dff_B_zyJ1kUiO0_2(.din(w_dff_B_aWVtrNGj7_2),.dout(w_dff_B_zyJ1kUiO0_2),.clk(gclk));
	jdff dff_B_j02usAVa0_2(.din(w_dff_B_zyJ1kUiO0_2),.dout(w_dff_B_j02usAVa0_2),.clk(gclk));
	jdff dff_B_4SqEQTPA9_2(.din(w_dff_B_j02usAVa0_2),.dout(w_dff_B_4SqEQTPA9_2),.clk(gclk));
	jdff dff_B_Ur1Yvhqh7_2(.din(w_dff_B_4SqEQTPA9_2),.dout(w_dff_B_Ur1Yvhqh7_2),.clk(gclk));
	jdff dff_B_ttgQNeSP6_2(.din(w_dff_B_Ur1Yvhqh7_2),.dout(w_dff_B_ttgQNeSP6_2),.clk(gclk));
	jdff dff_B_RTUYvkxv7_2(.din(w_dff_B_ttgQNeSP6_2),.dout(w_dff_B_RTUYvkxv7_2),.clk(gclk));
	jdff dff_B_VChcbkYF1_2(.din(w_dff_B_RTUYvkxv7_2),.dout(w_dff_B_VChcbkYF1_2),.clk(gclk));
	jdff dff_B_Mymb4dbm0_2(.din(w_dff_B_VChcbkYF1_2),.dout(w_dff_B_Mymb4dbm0_2),.clk(gclk));
	jdff dff_B_MRo1fH5Q9_2(.din(w_dff_B_Mymb4dbm0_2),.dout(w_dff_B_MRo1fH5Q9_2),.clk(gclk));
	jdff dff_B_Cad5qNF82_2(.din(w_dff_B_MRo1fH5Q9_2),.dout(w_dff_B_Cad5qNF82_2),.clk(gclk));
	jdff dff_B_b1nxdM0V6_2(.din(w_dff_B_Cad5qNF82_2),.dout(w_dff_B_b1nxdM0V6_2),.clk(gclk));
	jdff dff_B_NwW9LOgV5_2(.din(w_dff_B_b1nxdM0V6_2),.dout(w_dff_B_NwW9LOgV5_2),.clk(gclk));
	jdff dff_B_BunGjR6r7_2(.din(w_dff_B_NwW9LOgV5_2),.dout(w_dff_B_BunGjR6r7_2),.clk(gclk));
	jdff dff_B_FsOwk66u3_2(.din(w_dff_B_BunGjR6r7_2),.dout(w_dff_B_FsOwk66u3_2),.clk(gclk));
	jdff dff_B_uNqCDQEp1_2(.din(w_dff_B_FsOwk66u3_2),.dout(w_dff_B_uNqCDQEp1_2),.clk(gclk));
	jdff dff_B_uhVxvnRV0_2(.din(w_dff_B_uNqCDQEp1_2),.dout(w_dff_B_uhVxvnRV0_2),.clk(gclk));
	jdff dff_B_8jOKIvXi1_2(.din(w_dff_B_uhVxvnRV0_2),.dout(w_dff_B_8jOKIvXi1_2),.clk(gclk));
	jdff dff_B_7N7nnwl53_2(.din(w_dff_B_8jOKIvXi1_2),.dout(w_dff_B_7N7nnwl53_2),.clk(gclk));
	jdff dff_B_DVINhr4B0_2(.din(w_dff_B_7N7nnwl53_2),.dout(w_dff_B_DVINhr4B0_2),.clk(gclk));
	jdff dff_B_4hZRj11s0_2(.din(w_dff_B_DVINhr4B0_2),.dout(w_dff_B_4hZRj11s0_2),.clk(gclk));
	jdff dff_B_eFxfwSUJ7_2(.din(w_dff_B_4hZRj11s0_2),.dout(w_dff_B_eFxfwSUJ7_2),.clk(gclk));
	jdff dff_B_aiTdjmL76_2(.din(w_dff_B_eFxfwSUJ7_2),.dout(w_dff_B_aiTdjmL76_2),.clk(gclk));
	jdff dff_B_K0232ANi8_2(.din(w_dff_B_aiTdjmL76_2),.dout(w_dff_B_K0232ANi8_2),.clk(gclk));
	jdff dff_B_te5GG3Dy5_2(.din(w_dff_B_K0232ANi8_2),.dout(w_dff_B_te5GG3Dy5_2),.clk(gclk));
	jdff dff_B_F2cji9dj0_2(.din(w_dff_B_te5GG3Dy5_2),.dout(w_dff_B_F2cji9dj0_2),.clk(gclk));
	jdff dff_B_1AcWBykD1_2(.din(w_dff_B_F2cji9dj0_2),.dout(w_dff_B_1AcWBykD1_2),.clk(gclk));
	jdff dff_B_3WeEeyUq7_2(.din(w_dff_B_1AcWBykD1_2),.dout(w_dff_B_3WeEeyUq7_2),.clk(gclk));
	jdff dff_B_nP6Q6lid7_2(.din(w_dff_B_3WeEeyUq7_2),.dout(w_dff_B_nP6Q6lid7_2),.clk(gclk));
	jdff dff_B_HBO5oRPH1_2(.din(w_dff_B_nP6Q6lid7_2),.dout(w_dff_B_HBO5oRPH1_2),.clk(gclk));
	jdff dff_B_CAjFbE2G4_2(.din(w_dff_B_HBO5oRPH1_2),.dout(w_dff_B_CAjFbE2G4_2),.clk(gclk));
	jdff dff_B_pdJuQq7B8_1(.din(n1339),.dout(w_dff_B_pdJuQq7B8_1),.clk(gclk));
	jdff dff_B_chTdOyU17_2(.din(n1253),.dout(w_dff_B_chTdOyU17_2),.clk(gclk));
	jdff dff_B_Z2Q8o9qI7_2(.din(w_dff_B_chTdOyU17_2),.dout(w_dff_B_Z2Q8o9qI7_2),.clk(gclk));
	jdff dff_B_N4xaF1I83_2(.din(w_dff_B_Z2Q8o9qI7_2),.dout(w_dff_B_N4xaF1I83_2),.clk(gclk));
	jdff dff_B_fnokAywJ5_2(.din(w_dff_B_N4xaF1I83_2),.dout(w_dff_B_fnokAywJ5_2),.clk(gclk));
	jdff dff_B_NM8bVZpu9_2(.din(w_dff_B_fnokAywJ5_2),.dout(w_dff_B_NM8bVZpu9_2),.clk(gclk));
	jdff dff_B_2liClNdT1_2(.din(w_dff_B_NM8bVZpu9_2),.dout(w_dff_B_2liClNdT1_2),.clk(gclk));
	jdff dff_B_6NSKfvJq5_2(.din(w_dff_B_2liClNdT1_2),.dout(w_dff_B_6NSKfvJq5_2),.clk(gclk));
	jdff dff_B_Gvfcs4qJ3_2(.din(w_dff_B_6NSKfvJq5_2),.dout(w_dff_B_Gvfcs4qJ3_2),.clk(gclk));
	jdff dff_B_aB3ZMS1L8_2(.din(w_dff_B_Gvfcs4qJ3_2),.dout(w_dff_B_aB3ZMS1L8_2),.clk(gclk));
	jdff dff_B_u9npDKRN6_2(.din(w_dff_B_aB3ZMS1L8_2),.dout(w_dff_B_u9npDKRN6_2),.clk(gclk));
	jdff dff_B_B9aHE3oi2_2(.din(w_dff_B_u9npDKRN6_2),.dout(w_dff_B_B9aHE3oi2_2),.clk(gclk));
	jdff dff_B_Ei6sL0dE9_2(.din(w_dff_B_B9aHE3oi2_2),.dout(w_dff_B_Ei6sL0dE9_2),.clk(gclk));
	jdff dff_B_oo9UdODz6_2(.din(w_dff_B_Ei6sL0dE9_2),.dout(w_dff_B_oo9UdODz6_2),.clk(gclk));
	jdff dff_B_tBI6EE1Q0_2(.din(w_dff_B_oo9UdODz6_2),.dout(w_dff_B_tBI6EE1Q0_2),.clk(gclk));
	jdff dff_B_tZzyRcw01_2(.din(w_dff_B_tBI6EE1Q0_2),.dout(w_dff_B_tZzyRcw01_2),.clk(gclk));
	jdff dff_B_A5maOp4O6_2(.din(w_dff_B_tZzyRcw01_2),.dout(w_dff_B_A5maOp4O6_2),.clk(gclk));
	jdff dff_B_j1UCzGsH7_2(.din(w_dff_B_A5maOp4O6_2),.dout(w_dff_B_j1UCzGsH7_2),.clk(gclk));
	jdff dff_B_iSYxG9pj5_2(.din(w_dff_B_j1UCzGsH7_2),.dout(w_dff_B_iSYxG9pj5_2),.clk(gclk));
	jdff dff_B_UMJ4k9Yu1_2(.din(w_dff_B_iSYxG9pj5_2),.dout(w_dff_B_UMJ4k9Yu1_2),.clk(gclk));
	jdff dff_B_ZDpuUfWg8_2(.din(w_dff_B_UMJ4k9Yu1_2),.dout(w_dff_B_ZDpuUfWg8_2),.clk(gclk));
	jdff dff_B_BRKGf0Ev2_2(.din(w_dff_B_ZDpuUfWg8_2),.dout(w_dff_B_BRKGf0Ev2_2),.clk(gclk));
	jdff dff_B_7l7sEoCG9_2(.din(w_dff_B_BRKGf0Ev2_2),.dout(w_dff_B_7l7sEoCG9_2),.clk(gclk));
	jdff dff_B_nOgqgypv4_2(.din(w_dff_B_7l7sEoCG9_2),.dout(w_dff_B_nOgqgypv4_2),.clk(gclk));
	jdff dff_B_YclXjoTc9_2(.din(w_dff_B_nOgqgypv4_2),.dout(w_dff_B_YclXjoTc9_2),.clk(gclk));
	jdff dff_B_xatqhX4U5_2(.din(w_dff_B_YclXjoTc9_2),.dout(w_dff_B_xatqhX4U5_2),.clk(gclk));
	jdff dff_B_M7p0NrRz6_2(.din(w_dff_B_xatqhX4U5_2),.dout(w_dff_B_M7p0NrRz6_2),.clk(gclk));
	jdff dff_B_0TSKVTvp0_2(.din(w_dff_B_M7p0NrRz6_2),.dout(w_dff_B_0TSKVTvp0_2),.clk(gclk));
	jdff dff_B_SCIfQhJ49_2(.din(w_dff_B_0TSKVTvp0_2),.dout(w_dff_B_SCIfQhJ49_2),.clk(gclk));
	jdff dff_B_gq05zGsY8_2(.din(w_dff_B_SCIfQhJ49_2),.dout(w_dff_B_gq05zGsY8_2),.clk(gclk));
	jdff dff_B_LtheA07r3_2(.din(w_dff_B_gq05zGsY8_2),.dout(w_dff_B_LtheA07r3_2),.clk(gclk));
	jdff dff_B_ojVqX1w55_2(.din(w_dff_B_LtheA07r3_2),.dout(w_dff_B_ojVqX1w55_2),.clk(gclk));
	jdff dff_B_wSZW6EuG9_2(.din(w_dff_B_ojVqX1w55_2),.dout(w_dff_B_wSZW6EuG9_2),.clk(gclk));
	jdff dff_B_At1IcBmn8_2(.din(w_dff_B_wSZW6EuG9_2),.dout(w_dff_B_At1IcBmn8_2),.clk(gclk));
	jdff dff_B_iGi0t4qg6_2(.din(w_dff_B_At1IcBmn8_2),.dout(w_dff_B_iGi0t4qg6_2),.clk(gclk));
	jdff dff_B_lkkK2CV79_2(.din(w_dff_B_iGi0t4qg6_2),.dout(w_dff_B_lkkK2CV79_2),.clk(gclk));
	jdff dff_B_6ObnPa4j5_2(.din(w_dff_B_lkkK2CV79_2),.dout(w_dff_B_6ObnPa4j5_2),.clk(gclk));
	jdff dff_B_hn6oqsic3_2(.din(w_dff_B_6ObnPa4j5_2),.dout(w_dff_B_hn6oqsic3_2),.clk(gclk));
	jdff dff_B_pzi2CGvT6_2(.din(w_dff_B_hn6oqsic3_2),.dout(w_dff_B_pzi2CGvT6_2),.clk(gclk));
	jdff dff_B_PnKzv59X5_2(.din(w_dff_B_pzi2CGvT6_2),.dout(w_dff_B_PnKzv59X5_2),.clk(gclk));
	jdff dff_B_ohmRqlak2_2(.din(w_dff_B_PnKzv59X5_2),.dout(w_dff_B_ohmRqlak2_2),.clk(gclk));
	jdff dff_B_lpCrGuqL4_1(.din(n1254),.dout(w_dff_B_lpCrGuqL4_1),.clk(gclk));
	jdff dff_B_xMSg6Pv57_2(.din(n1163),.dout(w_dff_B_xMSg6Pv57_2),.clk(gclk));
	jdff dff_B_E9U3GXRQ5_2(.din(w_dff_B_xMSg6Pv57_2),.dout(w_dff_B_E9U3GXRQ5_2),.clk(gclk));
	jdff dff_B_CP7JYHcq8_2(.din(w_dff_B_E9U3GXRQ5_2),.dout(w_dff_B_CP7JYHcq8_2),.clk(gclk));
	jdff dff_B_L9GOE1g96_2(.din(w_dff_B_CP7JYHcq8_2),.dout(w_dff_B_L9GOE1g96_2),.clk(gclk));
	jdff dff_B_NoW9bIoI4_2(.din(w_dff_B_L9GOE1g96_2),.dout(w_dff_B_NoW9bIoI4_2),.clk(gclk));
	jdff dff_B_YFVVYW8j0_2(.din(w_dff_B_NoW9bIoI4_2),.dout(w_dff_B_YFVVYW8j0_2),.clk(gclk));
	jdff dff_B_a0Rvi3PB2_2(.din(w_dff_B_YFVVYW8j0_2),.dout(w_dff_B_a0Rvi3PB2_2),.clk(gclk));
	jdff dff_B_LBrZgVoU5_2(.din(w_dff_B_a0Rvi3PB2_2),.dout(w_dff_B_LBrZgVoU5_2),.clk(gclk));
	jdff dff_B_tk3aPc7C7_2(.din(w_dff_B_LBrZgVoU5_2),.dout(w_dff_B_tk3aPc7C7_2),.clk(gclk));
	jdff dff_B_u9ssFZvA8_2(.din(w_dff_B_tk3aPc7C7_2),.dout(w_dff_B_u9ssFZvA8_2),.clk(gclk));
	jdff dff_B_Fl0OUili8_2(.din(w_dff_B_u9ssFZvA8_2),.dout(w_dff_B_Fl0OUili8_2),.clk(gclk));
	jdff dff_B_hYDrS2Ux9_2(.din(w_dff_B_Fl0OUili8_2),.dout(w_dff_B_hYDrS2Ux9_2),.clk(gclk));
	jdff dff_B_DfHYd1zE0_2(.din(w_dff_B_hYDrS2Ux9_2),.dout(w_dff_B_DfHYd1zE0_2),.clk(gclk));
	jdff dff_B_jqxNP8hZ4_2(.din(w_dff_B_DfHYd1zE0_2),.dout(w_dff_B_jqxNP8hZ4_2),.clk(gclk));
	jdff dff_B_kuYCNlZG7_2(.din(w_dff_B_jqxNP8hZ4_2),.dout(w_dff_B_kuYCNlZG7_2),.clk(gclk));
	jdff dff_B_Px6qQJVb1_2(.din(w_dff_B_kuYCNlZG7_2),.dout(w_dff_B_Px6qQJVb1_2),.clk(gclk));
	jdff dff_B_VV58nyGG9_2(.din(w_dff_B_Px6qQJVb1_2),.dout(w_dff_B_VV58nyGG9_2),.clk(gclk));
	jdff dff_B_8eEwJLS32_2(.din(w_dff_B_VV58nyGG9_2),.dout(w_dff_B_8eEwJLS32_2),.clk(gclk));
	jdff dff_B_z2gX4LoL0_2(.din(w_dff_B_8eEwJLS32_2),.dout(w_dff_B_z2gX4LoL0_2),.clk(gclk));
	jdff dff_B_tZ7WiEt35_2(.din(w_dff_B_z2gX4LoL0_2),.dout(w_dff_B_tZ7WiEt35_2),.clk(gclk));
	jdff dff_B_kTUwXg5W8_2(.din(w_dff_B_tZ7WiEt35_2),.dout(w_dff_B_kTUwXg5W8_2),.clk(gclk));
	jdff dff_B_tTmRNDrj0_2(.din(w_dff_B_kTUwXg5W8_2),.dout(w_dff_B_tTmRNDrj0_2),.clk(gclk));
	jdff dff_B_LKiUVsHw3_2(.din(w_dff_B_tTmRNDrj0_2),.dout(w_dff_B_LKiUVsHw3_2),.clk(gclk));
	jdff dff_B_LnJBXjGF4_2(.din(w_dff_B_LKiUVsHw3_2),.dout(w_dff_B_LnJBXjGF4_2),.clk(gclk));
	jdff dff_B_8ymCK2S00_2(.din(w_dff_B_LnJBXjGF4_2),.dout(w_dff_B_8ymCK2S00_2),.clk(gclk));
	jdff dff_B_l0TVVT9J5_2(.din(w_dff_B_8ymCK2S00_2),.dout(w_dff_B_l0TVVT9J5_2),.clk(gclk));
	jdff dff_B_lnSV6onm5_2(.din(w_dff_B_l0TVVT9J5_2),.dout(w_dff_B_lnSV6onm5_2),.clk(gclk));
	jdff dff_B_oIsHcuvu5_2(.din(w_dff_B_lnSV6onm5_2),.dout(w_dff_B_oIsHcuvu5_2),.clk(gclk));
	jdff dff_B_TD1EOJbO4_2(.din(w_dff_B_oIsHcuvu5_2),.dout(w_dff_B_TD1EOJbO4_2),.clk(gclk));
	jdff dff_B_GTscYVNi9_2(.din(w_dff_B_TD1EOJbO4_2),.dout(w_dff_B_GTscYVNi9_2),.clk(gclk));
	jdff dff_B_0Pyrvwmj5_2(.din(w_dff_B_GTscYVNi9_2),.dout(w_dff_B_0Pyrvwmj5_2),.clk(gclk));
	jdff dff_B_ReYYuzyW9_2(.din(w_dff_B_0Pyrvwmj5_2),.dout(w_dff_B_ReYYuzyW9_2),.clk(gclk));
	jdff dff_B_QzHvZwvc8_2(.din(w_dff_B_ReYYuzyW9_2),.dout(w_dff_B_QzHvZwvc8_2),.clk(gclk));
	jdff dff_B_nBE31lqW3_2(.din(w_dff_B_QzHvZwvc8_2),.dout(w_dff_B_nBE31lqW3_2),.clk(gclk));
	jdff dff_B_M6j72Ivz5_2(.din(w_dff_B_nBE31lqW3_2),.dout(w_dff_B_M6j72Ivz5_2),.clk(gclk));
	jdff dff_B_tsGImOhK0_2(.din(w_dff_B_M6j72Ivz5_2),.dout(w_dff_B_tsGImOhK0_2),.clk(gclk));
	jdff dff_B_8aqOsc927_2(.din(w_dff_B_tsGImOhK0_2),.dout(w_dff_B_8aqOsc927_2),.clk(gclk));
	jdff dff_B_adC3VRFf2_1(.din(n1164),.dout(w_dff_B_adC3VRFf2_1),.clk(gclk));
	jdff dff_B_nZwFZUuS8_2(.din(n1059),.dout(w_dff_B_nZwFZUuS8_2),.clk(gclk));
	jdff dff_B_fghC81nT8_2(.din(w_dff_B_nZwFZUuS8_2),.dout(w_dff_B_fghC81nT8_2),.clk(gclk));
	jdff dff_B_W84BEZuG4_2(.din(w_dff_B_fghC81nT8_2),.dout(w_dff_B_W84BEZuG4_2),.clk(gclk));
	jdff dff_B_Q9Kvb8bM8_2(.din(w_dff_B_W84BEZuG4_2),.dout(w_dff_B_Q9Kvb8bM8_2),.clk(gclk));
	jdff dff_B_n8tv2Y4G5_2(.din(w_dff_B_Q9Kvb8bM8_2),.dout(w_dff_B_n8tv2Y4G5_2),.clk(gclk));
	jdff dff_B_MQ79rhWR4_2(.din(w_dff_B_n8tv2Y4G5_2),.dout(w_dff_B_MQ79rhWR4_2),.clk(gclk));
	jdff dff_B_CLBbNLD51_2(.din(w_dff_B_MQ79rhWR4_2),.dout(w_dff_B_CLBbNLD51_2),.clk(gclk));
	jdff dff_B_HeqE217R7_2(.din(w_dff_B_CLBbNLD51_2),.dout(w_dff_B_HeqE217R7_2),.clk(gclk));
	jdff dff_B_vID76VdG3_2(.din(w_dff_B_HeqE217R7_2),.dout(w_dff_B_vID76VdG3_2),.clk(gclk));
	jdff dff_B_ND2md9je1_2(.din(w_dff_B_vID76VdG3_2),.dout(w_dff_B_ND2md9je1_2),.clk(gclk));
	jdff dff_B_a5u4UEfa0_2(.din(w_dff_B_ND2md9je1_2),.dout(w_dff_B_a5u4UEfa0_2),.clk(gclk));
	jdff dff_B_gb6uSkQw7_2(.din(w_dff_B_a5u4UEfa0_2),.dout(w_dff_B_gb6uSkQw7_2),.clk(gclk));
	jdff dff_B_PIyZ6Yf77_2(.din(w_dff_B_gb6uSkQw7_2),.dout(w_dff_B_PIyZ6Yf77_2),.clk(gclk));
	jdff dff_B_Q9uXNTZf7_2(.din(w_dff_B_PIyZ6Yf77_2),.dout(w_dff_B_Q9uXNTZf7_2),.clk(gclk));
	jdff dff_B_eEQSogE30_2(.din(w_dff_B_Q9uXNTZf7_2),.dout(w_dff_B_eEQSogE30_2),.clk(gclk));
	jdff dff_B_rCIWTCVw9_2(.din(w_dff_B_eEQSogE30_2),.dout(w_dff_B_rCIWTCVw9_2),.clk(gclk));
	jdff dff_B_C3Y2j74P1_2(.din(w_dff_B_rCIWTCVw9_2),.dout(w_dff_B_C3Y2j74P1_2),.clk(gclk));
	jdff dff_B_hNCZ22lm5_2(.din(w_dff_B_C3Y2j74P1_2),.dout(w_dff_B_hNCZ22lm5_2),.clk(gclk));
	jdff dff_B_r7At73XZ7_2(.din(w_dff_B_hNCZ22lm5_2),.dout(w_dff_B_r7At73XZ7_2),.clk(gclk));
	jdff dff_B_at497RtK3_2(.din(w_dff_B_r7At73XZ7_2),.dout(w_dff_B_at497RtK3_2),.clk(gclk));
	jdff dff_B_oIaN6k833_2(.din(w_dff_B_at497RtK3_2),.dout(w_dff_B_oIaN6k833_2),.clk(gclk));
	jdff dff_B_z4ZJdOQc2_2(.din(w_dff_B_oIaN6k833_2),.dout(w_dff_B_z4ZJdOQc2_2),.clk(gclk));
	jdff dff_B_Z3NA1rv65_2(.din(w_dff_B_z4ZJdOQc2_2),.dout(w_dff_B_Z3NA1rv65_2),.clk(gclk));
	jdff dff_B_O8QjDOkw8_2(.din(w_dff_B_Z3NA1rv65_2),.dout(w_dff_B_O8QjDOkw8_2),.clk(gclk));
	jdff dff_B_JSWpm2pQ9_2(.din(w_dff_B_O8QjDOkw8_2),.dout(w_dff_B_JSWpm2pQ9_2),.clk(gclk));
	jdff dff_B_P6ywCwKw3_2(.din(w_dff_B_JSWpm2pQ9_2),.dout(w_dff_B_P6ywCwKw3_2),.clk(gclk));
	jdff dff_B_tgNWZzZ02_2(.din(w_dff_B_P6ywCwKw3_2),.dout(w_dff_B_tgNWZzZ02_2),.clk(gclk));
	jdff dff_B_NB4urrU51_2(.din(w_dff_B_tgNWZzZ02_2),.dout(w_dff_B_NB4urrU51_2),.clk(gclk));
	jdff dff_B_5GDDgcpi7_2(.din(w_dff_B_NB4urrU51_2),.dout(w_dff_B_5GDDgcpi7_2),.clk(gclk));
	jdff dff_B_IxXY4A5c0_2(.din(w_dff_B_5GDDgcpi7_2),.dout(w_dff_B_IxXY4A5c0_2),.clk(gclk));
	jdff dff_B_b8TbJFpE6_2(.din(w_dff_B_IxXY4A5c0_2),.dout(w_dff_B_b8TbJFpE6_2),.clk(gclk));
	jdff dff_B_7E5RzLfs3_2(.din(w_dff_B_b8TbJFpE6_2),.dout(w_dff_B_7E5RzLfs3_2),.clk(gclk));
	jdff dff_B_Gx4FnGt11_2(.din(w_dff_B_7E5RzLfs3_2),.dout(w_dff_B_Gx4FnGt11_2),.clk(gclk));
	jdff dff_B_hezCouQL0_2(.din(w_dff_B_Gx4FnGt11_2),.dout(w_dff_B_hezCouQL0_2),.clk(gclk));
	jdff dff_B_5UvB3LGI1_1(.din(n1060),.dout(w_dff_B_5UvB3LGI1_1),.clk(gclk));
	jdff dff_B_mCXEI6MU7_2(.din(n961),.dout(w_dff_B_mCXEI6MU7_2),.clk(gclk));
	jdff dff_B_O0VDQWk33_2(.din(w_dff_B_mCXEI6MU7_2),.dout(w_dff_B_O0VDQWk33_2),.clk(gclk));
	jdff dff_B_CzGRzmdV8_2(.din(w_dff_B_O0VDQWk33_2),.dout(w_dff_B_CzGRzmdV8_2),.clk(gclk));
	jdff dff_B_Zy6iEuIS8_2(.din(w_dff_B_CzGRzmdV8_2),.dout(w_dff_B_Zy6iEuIS8_2),.clk(gclk));
	jdff dff_B_Rzq0WHkh1_2(.din(w_dff_B_Zy6iEuIS8_2),.dout(w_dff_B_Rzq0WHkh1_2),.clk(gclk));
	jdff dff_B_3jIJbPnN8_2(.din(w_dff_B_Rzq0WHkh1_2),.dout(w_dff_B_3jIJbPnN8_2),.clk(gclk));
	jdff dff_B_vSRM9jtN1_2(.din(w_dff_B_3jIJbPnN8_2),.dout(w_dff_B_vSRM9jtN1_2),.clk(gclk));
	jdff dff_B_C064Ldx37_2(.din(w_dff_B_vSRM9jtN1_2),.dout(w_dff_B_C064Ldx37_2),.clk(gclk));
	jdff dff_B_UqCfUbbl0_2(.din(w_dff_B_C064Ldx37_2),.dout(w_dff_B_UqCfUbbl0_2),.clk(gclk));
	jdff dff_B_4gNqZQ6U3_2(.din(w_dff_B_UqCfUbbl0_2),.dout(w_dff_B_4gNqZQ6U3_2),.clk(gclk));
	jdff dff_B_a3Pynn9J5_2(.din(w_dff_B_4gNqZQ6U3_2),.dout(w_dff_B_a3Pynn9J5_2),.clk(gclk));
	jdff dff_B_c7KDfeEO5_2(.din(w_dff_B_a3Pynn9J5_2),.dout(w_dff_B_c7KDfeEO5_2),.clk(gclk));
	jdff dff_B_gBzgjfyH6_2(.din(w_dff_B_c7KDfeEO5_2),.dout(w_dff_B_gBzgjfyH6_2),.clk(gclk));
	jdff dff_B_5SEIbU7t3_2(.din(w_dff_B_gBzgjfyH6_2),.dout(w_dff_B_5SEIbU7t3_2),.clk(gclk));
	jdff dff_B_415qIkVG1_2(.din(w_dff_B_5SEIbU7t3_2),.dout(w_dff_B_415qIkVG1_2),.clk(gclk));
	jdff dff_B_v3rUocvQ8_2(.din(w_dff_B_415qIkVG1_2),.dout(w_dff_B_v3rUocvQ8_2),.clk(gclk));
	jdff dff_B_3haXmg0g8_2(.din(w_dff_B_v3rUocvQ8_2),.dout(w_dff_B_3haXmg0g8_2),.clk(gclk));
	jdff dff_B_KNCiGKZ97_2(.din(w_dff_B_3haXmg0g8_2),.dout(w_dff_B_KNCiGKZ97_2),.clk(gclk));
	jdff dff_B_rf24kMxm6_2(.din(w_dff_B_KNCiGKZ97_2),.dout(w_dff_B_rf24kMxm6_2),.clk(gclk));
	jdff dff_B_lNUudiTQ0_2(.din(w_dff_B_rf24kMxm6_2),.dout(w_dff_B_lNUudiTQ0_2),.clk(gclk));
	jdff dff_B_2UpIYckQ7_2(.din(w_dff_B_lNUudiTQ0_2),.dout(w_dff_B_2UpIYckQ7_2),.clk(gclk));
	jdff dff_B_QQtLohz15_2(.din(w_dff_B_2UpIYckQ7_2),.dout(w_dff_B_QQtLohz15_2),.clk(gclk));
	jdff dff_B_aYNdfhs14_2(.din(w_dff_B_QQtLohz15_2),.dout(w_dff_B_aYNdfhs14_2),.clk(gclk));
	jdff dff_B_L1fuHQAh4_2(.din(w_dff_B_aYNdfhs14_2),.dout(w_dff_B_L1fuHQAh4_2),.clk(gclk));
	jdff dff_B_MTCZ4dim3_2(.din(w_dff_B_L1fuHQAh4_2),.dout(w_dff_B_MTCZ4dim3_2),.clk(gclk));
	jdff dff_B_qt7G1FVR1_2(.din(w_dff_B_MTCZ4dim3_2),.dout(w_dff_B_qt7G1FVR1_2),.clk(gclk));
	jdff dff_B_NP9hEVwk7_2(.din(w_dff_B_qt7G1FVR1_2),.dout(w_dff_B_NP9hEVwk7_2),.clk(gclk));
	jdff dff_B_U4zjTHIe6_2(.din(w_dff_B_NP9hEVwk7_2),.dout(w_dff_B_U4zjTHIe6_2),.clk(gclk));
	jdff dff_B_dYxUp4ZZ2_2(.din(w_dff_B_U4zjTHIe6_2),.dout(w_dff_B_dYxUp4ZZ2_2),.clk(gclk));
	jdff dff_B_ftWiGBnT3_2(.din(w_dff_B_dYxUp4ZZ2_2),.dout(w_dff_B_ftWiGBnT3_2),.clk(gclk));
	jdff dff_B_9hb6a1Uh9_2(.din(w_dff_B_ftWiGBnT3_2),.dout(w_dff_B_9hb6a1Uh9_2),.clk(gclk));
	jdff dff_B_hgj8ijXl0_1(.din(n962),.dout(w_dff_B_hgj8ijXl0_1),.clk(gclk));
	jdff dff_B_SVC12NAg3_2(.din(n856),.dout(w_dff_B_SVC12NAg3_2),.clk(gclk));
	jdff dff_B_T8Zumf2g3_2(.din(w_dff_B_SVC12NAg3_2),.dout(w_dff_B_T8Zumf2g3_2),.clk(gclk));
	jdff dff_B_6qLkuQYL8_2(.din(w_dff_B_T8Zumf2g3_2),.dout(w_dff_B_6qLkuQYL8_2),.clk(gclk));
	jdff dff_B_fqbulSk57_2(.din(w_dff_B_6qLkuQYL8_2),.dout(w_dff_B_fqbulSk57_2),.clk(gclk));
	jdff dff_B_iDJaM1gZ3_2(.din(w_dff_B_fqbulSk57_2),.dout(w_dff_B_iDJaM1gZ3_2),.clk(gclk));
	jdff dff_B_KGVodRJG6_2(.din(w_dff_B_iDJaM1gZ3_2),.dout(w_dff_B_KGVodRJG6_2),.clk(gclk));
	jdff dff_B_Ranb23lH1_2(.din(w_dff_B_KGVodRJG6_2),.dout(w_dff_B_Ranb23lH1_2),.clk(gclk));
	jdff dff_B_T7WTgaHo4_2(.din(w_dff_B_Ranb23lH1_2),.dout(w_dff_B_T7WTgaHo4_2),.clk(gclk));
	jdff dff_B_NuDEaQ5W8_2(.din(w_dff_B_T7WTgaHo4_2),.dout(w_dff_B_NuDEaQ5W8_2),.clk(gclk));
	jdff dff_B_USGlNJi82_2(.din(w_dff_B_NuDEaQ5W8_2),.dout(w_dff_B_USGlNJi82_2),.clk(gclk));
	jdff dff_B_r1SfLcPh4_2(.din(w_dff_B_USGlNJi82_2),.dout(w_dff_B_r1SfLcPh4_2),.clk(gclk));
	jdff dff_B_rlHly6nH8_2(.din(w_dff_B_r1SfLcPh4_2),.dout(w_dff_B_rlHly6nH8_2),.clk(gclk));
	jdff dff_B_E0ZwuUQ76_2(.din(w_dff_B_rlHly6nH8_2),.dout(w_dff_B_E0ZwuUQ76_2),.clk(gclk));
	jdff dff_B_Wd3YRfVH6_2(.din(w_dff_B_E0ZwuUQ76_2),.dout(w_dff_B_Wd3YRfVH6_2),.clk(gclk));
	jdff dff_B_USoAhaje4_2(.din(w_dff_B_Wd3YRfVH6_2),.dout(w_dff_B_USoAhaje4_2),.clk(gclk));
	jdff dff_B_1A3IAvez5_2(.din(w_dff_B_USoAhaje4_2),.dout(w_dff_B_1A3IAvez5_2),.clk(gclk));
	jdff dff_B_uwKaJnVk3_2(.din(w_dff_B_1A3IAvez5_2),.dout(w_dff_B_uwKaJnVk3_2),.clk(gclk));
	jdff dff_B_52vhSuAy0_2(.din(w_dff_B_uwKaJnVk3_2),.dout(w_dff_B_52vhSuAy0_2),.clk(gclk));
	jdff dff_B_MzU2Z5P66_2(.din(w_dff_B_52vhSuAy0_2),.dout(w_dff_B_MzU2Z5P66_2),.clk(gclk));
	jdff dff_B_rFlLrsM89_2(.din(w_dff_B_MzU2Z5P66_2),.dout(w_dff_B_rFlLrsM89_2),.clk(gclk));
	jdff dff_B_FoivV4FK2_2(.din(w_dff_B_rFlLrsM89_2),.dout(w_dff_B_FoivV4FK2_2),.clk(gclk));
	jdff dff_B_1lSY83kJ5_2(.din(w_dff_B_FoivV4FK2_2),.dout(w_dff_B_1lSY83kJ5_2),.clk(gclk));
	jdff dff_B_U6pn8MCV0_2(.din(w_dff_B_1lSY83kJ5_2),.dout(w_dff_B_U6pn8MCV0_2),.clk(gclk));
	jdff dff_B_FRwaVpTt6_2(.din(w_dff_B_U6pn8MCV0_2),.dout(w_dff_B_FRwaVpTt6_2),.clk(gclk));
	jdff dff_B_YbsbpVBo5_2(.din(w_dff_B_FRwaVpTt6_2),.dout(w_dff_B_YbsbpVBo5_2),.clk(gclk));
	jdff dff_B_DogKVEKI8_2(.din(w_dff_B_YbsbpVBo5_2),.dout(w_dff_B_DogKVEKI8_2),.clk(gclk));
	jdff dff_B_EvPQsQTx9_2(.din(w_dff_B_DogKVEKI8_2),.dout(w_dff_B_EvPQsQTx9_2),.clk(gclk));
	jdff dff_B_lyf6aRnj3_2(.din(w_dff_B_EvPQsQTx9_2),.dout(w_dff_B_lyf6aRnj3_2),.clk(gclk));
	jdff dff_B_ejihLi905_1(.din(n857),.dout(w_dff_B_ejihLi905_1),.clk(gclk));
	jdff dff_B_8tmlnGSw0_2(.din(n757),.dout(w_dff_B_8tmlnGSw0_2),.clk(gclk));
	jdff dff_B_jYs3cOUC2_2(.din(w_dff_B_8tmlnGSw0_2),.dout(w_dff_B_jYs3cOUC2_2),.clk(gclk));
	jdff dff_B_rnlV4XhB4_2(.din(w_dff_B_jYs3cOUC2_2),.dout(w_dff_B_rnlV4XhB4_2),.clk(gclk));
	jdff dff_B_5bgru6wk6_2(.din(w_dff_B_rnlV4XhB4_2),.dout(w_dff_B_5bgru6wk6_2),.clk(gclk));
	jdff dff_B_5FJUSTER4_2(.din(w_dff_B_5bgru6wk6_2),.dout(w_dff_B_5FJUSTER4_2),.clk(gclk));
	jdff dff_B_TgHwNfGx5_2(.din(w_dff_B_5FJUSTER4_2),.dout(w_dff_B_TgHwNfGx5_2),.clk(gclk));
	jdff dff_B_BIfroLRr4_2(.din(w_dff_B_TgHwNfGx5_2),.dout(w_dff_B_BIfroLRr4_2),.clk(gclk));
	jdff dff_B_KLTNwEvz7_2(.din(w_dff_B_BIfroLRr4_2),.dout(w_dff_B_KLTNwEvz7_2),.clk(gclk));
	jdff dff_B_A9JB9CBx1_2(.din(w_dff_B_KLTNwEvz7_2),.dout(w_dff_B_A9JB9CBx1_2),.clk(gclk));
	jdff dff_B_B79SkSOP5_2(.din(w_dff_B_A9JB9CBx1_2),.dout(w_dff_B_B79SkSOP5_2),.clk(gclk));
	jdff dff_B_kVzTENRN5_2(.din(w_dff_B_B79SkSOP5_2),.dout(w_dff_B_kVzTENRN5_2),.clk(gclk));
	jdff dff_B_HOolG97J3_2(.din(w_dff_B_kVzTENRN5_2),.dout(w_dff_B_HOolG97J3_2),.clk(gclk));
	jdff dff_B_ub6LlqDt7_2(.din(w_dff_B_HOolG97J3_2),.dout(w_dff_B_ub6LlqDt7_2),.clk(gclk));
	jdff dff_B_rXfaiVXV7_2(.din(w_dff_B_ub6LlqDt7_2),.dout(w_dff_B_rXfaiVXV7_2),.clk(gclk));
	jdff dff_B_OmLrzGUh4_2(.din(w_dff_B_rXfaiVXV7_2),.dout(w_dff_B_OmLrzGUh4_2),.clk(gclk));
	jdff dff_B_rVcu2sb88_2(.din(w_dff_B_OmLrzGUh4_2),.dout(w_dff_B_rVcu2sb88_2),.clk(gclk));
	jdff dff_B_tiC8XncD4_2(.din(w_dff_B_rVcu2sb88_2),.dout(w_dff_B_tiC8XncD4_2),.clk(gclk));
	jdff dff_B_NFzBo2b02_2(.din(w_dff_B_tiC8XncD4_2),.dout(w_dff_B_NFzBo2b02_2),.clk(gclk));
	jdff dff_B_4oNoGlTu0_2(.din(w_dff_B_NFzBo2b02_2),.dout(w_dff_B_4oNoGlTu0_2),.clk(gclk));
	jdff dff_B_zkskbeVv0_2(.din(w_dff_B_4oNoGlTu0_2),.dout(w_dff_B_zkskbeVv0_2),.clk(gclk));
	jdff dff_B_DBALOCue2_2(.din(w_dff_B_zkskbeVv0_2),.dout(w_dff_B_DBALOCue2_2),.clk(gclk));
	jdff dff_B_exPGFf5H8_2(.din(w_dff_B_DBALOCue2_2),.dout(w_dff_B_exPGFf5H8_2),.clk(gclk));
	jdff dff_B_X27X6G9E4_2(.din(w_dff_B_exPGFf5H8_2),.dout(w_dff_B_X27X6G9E4_2),.clk(gclk));
	jdff dff_B_rVdzUtEe9_2(.din(w_dff_B_X27X6G9E4_2),.dout(w_dff_B_rVdzUtEe9_2),.clk(gclk));
	jdff dff_B_kRNE0XN38_2(.din(w_dff_B_rVdzUtEe9_2),.dout(w_dff_B_kRNE0XN38_2),.clk(gclk));
	jdff dff_B_bcO87PmO5_1(.din(n758),.dout(w_dff_B_bcO87PmO5_1),.clk(gclk));
	jdff dff_B_15o0CNIv7_2(.din(n664),.dout(w_dff_B_15o0CNIv7_2),.clk(gclk));
	jdff dff_B_xDZqN6vV3_2(.din(w_dff_B_15o0CNIv7_2),.dout(w_dff_B_xDZqN6vV3_2),.clk(gclk));
	jdff dff_B_WxaKVyv42_2(.din(w_dff_B_xDZqN6vV3_2),.dout(w_dff_B_WxaKVyv42_2),.clk(gclk));
	jdff dff_B_1oUppQOW7_2(.din(w_dff_B_WxaKVyv42_2),.dout(w_dff_B_1oUppQOW7_2),.clk(gclk));
	jdff dff_B_RTD3wpxT4_2(.din(w_dff_B_1oUppQOW7_2),.dout(w_dff_B_RTD3wpxT4_2),.clk(gclk));
	jdff dff_B_O6tY3K6D3_2(.din(w_dff_B_RTD3wpxT4_2),.dout(w_dff_B_O6tY3K6D3_2),.clk(gclk));
	jdff dff_B_VIM8IrZv5_2(.din(w_dff_B_O6tY3K6D3_2),.dout(w_dff_B_VIM8IrZv5_2),.clk(gclk));
	jdff dff_B_zZP8cuCn5_2(.din(w_dff_B_VIM8IrZv5_2),.dout(w_dff_B_zZP8cuCn5_2),.clk(gclk));
	jdff dff_B_SggYFhFN6_2(.din(w_dff_B_zZP8cuCn5_2),.dout(w_dff_B_SggYFhFN6_2),.clk(gclk));
	jdff dff_B_w3hIOeJM8_2(.din(w_dff_B_SggYFhFN6_2),.dout(w_dff_B_w3hIOeJM8_2),.clk(gclk));
	jdff dff_B_bgnhEpoc2_2(.din(w_dff_B_w3hIOeJM8_2),.dout(w_dff_B_bgnhEpoc2_2),.clk(gclk));
	jdff dff_B_9aT2FqOb2_2(.din(w_dff_B_bgnhEpoc2_2),.dout(w_dff_B_9aT2FqOb2_2),.clk(gclk));
	jdff dff_B_XF7sNaeb1_2(.din(w_dff_B_9aT2FqOb2_2),.dout(w_dff_B_XF7sNaeb1_2),.clk(gclk));
	jdff dff_B_g8ZFeTXx7_2(.din(w_dff_B_XF7sNaeb1_2),.dout(w_dff_B_g8ZFeTXx7_2),.clk(gclk));
	jdff dff_B_juyLj4hL1_2(.din(w_dff_B_g8ZFeTXx7_2),.dout(w_dff_B_juyLj4hL1_2),.clk(gclk));
	jdff dff_B_VoESLRuS1_2(.din(w_dff_B_juyLj4hL1_2),.dout(w_dff_B_VoESLRuS1_2),.clk(gclk));
	jdff dff_B_AqrnZTjL2_2(.din(w_dff_B_VoESLRuS1_2),.dout(w_dff_B_AqrnZTjL2_2),.clk(gclk));
	jdff dff_B_RZYSF6Ie9_2(.din(w_dff_B_AqrnZTjL2_2),.dout(w_dff_B_RZYSF6Ie9_2),.clk(gclk));
	jdff dff_B_zu2LB1KE1_2(.din(w_dff_B_RZYSF6Ie9_2),.dout(w_dff_B_zu2LB1KE1_2),.clk(gclk));
	jdff dff_B_bwquSfY57_2(.din(w_dff_B_zu2LB1KE1_2),.dout(w_dff_B_bwquSfY57_2),.clk(gclk));
	jdff dff_B_sOd524Ka7_2(.din(w_dff_B_bwquSfY57_2),.dout(w_dff_B_sOd524Ka7_2),.clk(gclk));
	jdff dff_B_aetrGM480_2(.din(w_dff_B_sOd524Ka7_2),.dout(w_dff_B_aetrGM480_2),.clk(gclk));
	jdff dff_B_URPxwRpp9_1(.din(n665),.dout(w_dff_B_URPxwRpp9_1),.clk(gclk));
	jdff dff_B_JX1JPsH39_2(.din(n578),.dout(w_dff_B_JX1JPsH39_2),.clk(gclk));
	jdff dff_B_LzIMJpeT5_2(.din(w_dff_B_JX1JPsH39_2),.dout(w_dff_B_LzIMJpeT5_2),.clk(gclk));
	jdff dff_B_RHRCl1m07_2(.din(w_dff_B_LzIMJpeT5_2),.dout(w_dff_B_RHRCl1m07_2),.clk(gclk));
	jdff dff_B_kVRLkMIe7_2(.din(w_dff_B_RHRCl1m07_2),.dout(w_dff_B_kVRLkMIe7_2),.clk(gclk));
	jdff dff_B_JrghY2dp3_2(.din(w_dff_B_kVRLkMIe7_2),.dout(w_dff_B_JrghY2dp3_2),.clk(gclk));
	jdff dff_B_VIqPRXn84_2(.din(w_dff_B_JrghY2dp3_2),.dout(w_dff_B_VIqPRXn84_2),.clk(gclk));
	jdff dff_B_86Mvjovt1_2(.din(w_dff_B_VIqPRXn84_2),.dout(w_dff_B_86Mvjovt1_2),.clk(gclk));
	jdff dff_B_tJqfScUJ3_2(.din(w_dff_B_86Mvjovt1_2),.dout(w_dff_B_tJqfScUJ3_2),.clk(gclk));
	jdff dff_B_pHeX8w844_2(.din(w_dff_B_tJqfScUJ3_2),.dout(w_dff_B_pHeX8w844_2),.clk(gclk));
	jdff dff_B_gxYV5lXF4_2(.din(w_dff_B_pHeX8w844_2),.dout(w_dff_B_gxYV5lXF4_2),.clk(gclk));
	jdff dff_B_j4FeBo5q3_2(.din(w_dff_B_gxYV5lXF4_2),.dout(w_dff_B_j4FeBo5q3_2),.clk(gclk));
	jdff dff_B_A4h8XyKt2_2(.din(w_dff_B_j4FeBo5q3_2),.dout(w_dff_B_A4h8XyKt2_2),.clk(gclk));
	jdff dff_B_fxIZkuyq5_2(.din(w_dff_B_A4h8XyKt2_2),.dout(w_dff_B_fxIZkuyq5_2),.clk(gclk));
	jdff dff_B_OVMCcV4M9_2(.din(w_dff_B_fxIZkuyq5_2),.dout(w_dff_B_OVMCcV4M9_2),.clk(gclk));
	jdff dff_B_d4lPeMhm0_2(.din(w_dff_B_OVMCcV4M9_2),.dout(w_dff_B_d4lPeMhm0_2),.clk(gclk));
	jdff dff_B_gxhFJIEX7_2(.din(w_dff_B_d4lPeMhm0_2),.dout(w_dff_B_gxhFJIEX7_2),.clk(gclk));
	jdff dff_B_PfbytpzH3_2(.din(w_dff_B_gxhFJIEX7_2),.dout(w_dff_B_PfbytpzH3_2),.clk(gclk));
	jdff dff_B_9p9WPMGU1_2(.din(w_dff_B_PfbytpzH3_2),.dout(w_dff_B_9p9WPMGU1_2),.clk(gclk));
	jdff dff_B_36Zt8hAt2_2(.din(w_dff_B_9p9WPMGU1_2),.dout(w_dff_B_36Zt8hAt2_2),.clk(gclk));
	jdff dff_B_mt15VX7D5_1(.din(n579),.dout(w_dff_B_mt15VX7D5_1),.clk(gclk));
	jdff dff_B_QDVq3hhf5_2(.din(n499),.dout(w_dff_B_QDVq3hhf5_2),.clk(gclk));
	jdff dff_B_laVjKb8a7_2(.din(w_dff_B_QDVq3hhf5_2),.dout(w_dff_B_laVjKb8a7_2),.clk(gclk));
	jdff dff_B_13uV7ovM8_2(.din(w_dff_B_laVjKb8a7_2),.dout(w_dff_B_13uV7ovM8_2),.clk(gclk));
	jdff dff_B_TWvCCRVY6_2(.din(w_dff_B_13uV7ovM8_2),.dout(w_dff_B_TWvCCRVY6_2),.clk(gclk));
	jdff dff_B_SV5xxY753_2(.din(w_dff_B_TWvCCRVY6_2),.dout(w_dff_B_SV5xxY753_2),.clk(gclk));
	jdff dff_B_5Vk9CDUZ0_2(.din(w_dff_B_SV5xxY753_2),.dout(w_dff_B_5Vk9CDUZ0_2),.clk(gclk));
	jdff dff_B_sqsRiXlB5_2(.din(w_dff_B_5Vk9CDUZ0_2),.dout(w_dff_B_sqsRiXlB5_2),.clk(gclk));
	jdff dff_B_HsnvKVp48_2(.din(w_dff_B_sqsRiXlB5_2),.dout(w_dff_B_HsnvKVp48_2),.clk(gclk));
	jdff dff_B_m50m7EFJ1_2(.din(w_dff_B_HsnvKVp48_2),.dout(w_dff_B_m50m7EFJ1_2),.clk(gclk));
	jdff dff_B_CLPglvEP6_2(.din(w_dff_B_m50m7EFJ1_2),.dout(w_dff_B_CLPglvEP6_2),.clk(gclk));
	jdff dff_B_41jZgiFH2_2(.din(w_dff_B_CLPglvEP6_2),.dout(w_dff_B_41jZgiFH2_2),.clk(gclk));
	jdff dff_B_iWxlPfgi3_2(.din(w_dff_B_41jZgiFH2_2),.dout(w_dff_B_iWxlPfgi3_2),.clk(gclk));
	jdff dff_B_VzJY0HY34_2(.din(w_dff_B_iWxlPfgi3_2),.dout(w_dff_B_VzJY0HY34_2),.clk(gclk));
	jdff dff_B_BtmYRip35_2(.din(w_dff_B_VzJY0HY34_2),.dout(w_dff_B_BtmYRip35_2),.clk(gclk));
	jdff dff_B_NiKik2ow3_2(.din(w_dff_B_BtmYRip35_2),.dout(w_dff_B_NiKik2ow3_2),.clk(gclk));
	jdff dff_B_En3EkI4x6_2(.din(w_dff_B_NiKik2ow3_2),.dout(w_dff_B_En3EkI4x6_2),.clk(gclk));
	jdff dff_B_6mIyvaqr8_1(.din(n500),.dout(w_dff_B_6mIyvaqr8_1),.clk(gclk));
	jdff dff_B_ZkG2sCKQ3_2(.din(n427),.dout(w_dff_B_ZkG2sCKQ3_2),.clk(gclk));
	jdff dff_B_yz6FXYRl2_2(.din(w_dff_B_ZkG2sCKQ3_2),.dout(w_dff_B_yz6FXYRl2_2),.clk(gclk));
	jdff dff_B_PvE48pp64_2(.din(w_dff_B_yz6FXYRl2_2),.dout(w_dff_B_PvE48pp64_2),.clk(gclk));
	jdff dff_B_RzRloISO6_2(.din(w_dff_B_PvE48pp64_2),.dout(w_dff_B_RzRloISO6_2),.clk(gclk));
	jdff dff_B_DpzYwDeu2_2(.din(w_dff_B_RzRloISO6_2),.dout(w_dff_B_DpzYwDeu2_2),.clk(gclk));
	jdff dff_B_auSHm8h75_2(.din(w_dff_B_DpzYwDeu2_2),.dout(w_dff_B_auSHm8h75_2),.clk(gclk));
	jdff dff_B_UTZuA6aA1_2(.din(w_dff_B_auSHm8h75_2),.dout(w_dff_B_UTZuA6aA1_2),.clk(gclk));
	jdff dff_B_aLw4IxKS5_2(.din(w_dff_B_UTZuA6aA1_2),.dout(w_dff_B_aLw4IxKS5_2),.clk(gclk));
	jdff dff_B_a5EYDvMD5_2(.din(w_dff_B_aLw4IxKS5_2),.dout(w_dff_B_a5EYDvMD5_2),.clk(gclk));
	jdff dff_B_jCqgFF7T6_2(.din(w_dff_B_a5EYDvMD5_2),.dout(w_dff_B_jCqgFF7T6_2),.clk(gclk));
	jdff dff_B_bbkjXoID6_2(.din(w_dff_B_jCqgFF7T6_2),.dout(w_dff_B_bbkjXoID6_2),.clk(gclk));
	jdff dff_B_B72SyqhR8_2(.din(w_dff_B_bbkjXoID6_2),.dout(w_dff_B_B72SyqhR8_2),.clk(gclk));
	jdff dff_B_7NIX7gzS4_2(.din(w_dff_B_B72SyqhR8_2),.dout(w_dff_B_7NIX7gzS4_2),.clk(gclk));
	jdff dff_B_WEau1fSs0_1(.din(n428),.dout(w_dff_B_WEau1fSs0_1),.clk(gclk));
	jdff dff_B_o8LENZfH4_2(.din(n363),.dout(w_dff_B_o8LENZfH4_2),.clk(gclk));
	jdff dff_B_mYcDDcaN1_2(.din(w_dff_B_o8LENZfH4_2),.dout(w_dff_B_mYcDDcaN1_2),.clk(gclk));
	jdff dff_B_3xPx2mjP2_2(.din(w_dff_B_mYcDDcaN1_2),.dout(w_dff_B_3xPx2mjP2_2),.clk(gclk));
	jdff dff_B_EU0XWfQ37_2(.din(w_dff_B_3xPx2mjP2_2),.dout(w_dff_B_EU0XWfQ37_2),.clk(gclk));
	jdff dff_B_1WI1LxuM9_2(.din(w_dff_B_EU0XWfQ37_2),.dout(w_dff_B_1WI1LxuM9_2),.clk(gclk));
	jdff dff_B_Mq67UBh45_2(.din(w_dff_B_1WI1LxuM9_2),.dout(w_dff_B_Mq67UBh45_2),.clk(gclk));
	jdff dff_B_GkKC40wH3_2(.din(w_dff_B_Mq67UBh45_2),.dout(w_dff_B_GkKC40wH3_2),.clk(gclk));
	jdff dff_B_Vd9qOpJS2_2(.din(w_dff_B_GkKC40wH3_2),.dout(w_dff_B_Vd9qOpJS2_2),.clk(gclk));
	jdff dff_B_1I7m3Dei3_2(.din(w_dff_B_Vd9qOpJS2_2),.dout(w_dff_B_1I7m3Dei3_2),.clk(gclk));
	jdff dff_B_21WflzzA2_2(.din(w_dff_B_1I7m3Dei3_2),.dout(w_dff_B_21WflzzA2_2),.clk(gclk));
	jdff dff_B_hGv4qMwx9_2(.din(n385),.dout(w_dff_B_hGv4qMwx9_2),.clk(gclk));
	jdff dff_B_BRvDgPUz5_1(.din(n364),.dout(w_dff_B_BRvDgPUz5_1),.clk(gclk));
	jdff dff_B_gkTAIXDB4_2(.din(n305),.dout(w_dff_B_gkTAIXDB4_2),.clk(gclk));
	jdff dff_B_5AEfshf03_2(.din(w_dff_B_gkTAIXDB4_2),.dout(w_dff_B_5AEfshf03_2),.clk(gclk));
	jdff dff_B_sn5xgl242_2(.din(w_dff_B_5AEfshf03_2),.dout(w_dff_B_sn5xgl242_2),.clk(gclk));
	jdff dff_B_StLJC8py1_2(.din(w_dff_B_sn5xgl242_2),.dout(w_dff_B_StLJC8py1_2),.clk(gclk));
	jdff dff_B_3aGprczc4_2(.din(w_dff_B_StLJC8py1_2),.dout(w_dff_B_3aGprczc4_2),.clk(gclk));
	jdff dff_B_BuSQx6z12_2(.din(w_dff_B_3aGprczc4_2),.dout(w_dff_B_BuSQx6z12_2),.clk(gclk));
	jdff dff_B_6rTgYPtY9_2(.din(w_dff_B_BuSQx6z12_2),.dout(w_dff_B_6rTgYPtY9_2),.clk(gclk));
	jdff dff_B_VPsceqs67_2(.din(n321),.dout(w_dff_B_VPsceqs67_2),.clk(gclk));
	jdff dff_B_zXRprNEB1_1(.din(n306),.dout(w_dff_B_zXRprNEB1_1),.clk(gclk));
	jdff dff_B_pfL42Ayq3_2(.din(n254),.dout(w_dff_B_pfL42Ayq3_2),.clk(gclk));
	jdff dff_B_qx0OKX9I8_2(.din(w_dff_B_pfL42Ayq3_2),.dout(w_dff_B_qx0OKX9I8_2),.clk(gclk));
	jdff dff_B_DPBQgWQQ8_2(.din(w_dff_B_qx0OKX9I8_2),.dout(w_dff_B_DPBQgWQQ8_2),.clk(gclk));
	jdff dff_B_u3Vi490M7_2(.din(w_dff_B_DPBQgWQQ8_2),.dout(w_dff_B_u3Vi490M7_2),.clk(gclk));
	jdff dff_B_9hPIJqTT8_1(.din(n256),.dout(w_dff_B_9hPIJqTT8_1),.clk(gclk));
	jdff dff_A_mTvMtSiG7_1(.dout(w_n210_0[1]),.din(w_dff_A_mTvMtSiG7_1),.clk(gclk));
	jdff dff_A_9AFadnxN6_2(.dout(w_n210_0[2]),.din(w_dff_A_9AFadnxN6_2),.clk(gclk));
	jdff dff_A_Y3Yw9DWj9_2(.dout(w_dff_A_9AFadnxN6_2),.din(w_dff_A_Y3Yw9DWj9_2),.clk(gclk));
	jdff dff_B_af4nwA5n9_2(.din(n1496),.dout(w_dff_B_af4nwA5n9_2),.clk(gclk));
	jdff dff_B_lyPa9dUU4_1(.din(n1494),.dout(w_dff_B_lyPa9dUU4_1),.clk(gclk));
	jdff dff_B_b91cSgik3_2(.din(n1421),.dout(w_dff_B_b91cSgik3_2),.clk(gclk));
	jdff dff_B_oSg7x4ko5_2(.din(w_dff_B_b91cSgik3_2),.dout(w_dff_B_oSg7x4ko5_2),.clk(gclk));
	jdff dff_B_qjZqg0KE8_2(.din(w_dff_B_oSg7x4ko5_2),.dout(w_dff_B_qjZqg0KE8_2),.clk(gclk));
	jdff dff_B_u7AMRP7r4_2(.din(w_dff_B_qjZqg0KE8_2),.dout(w_dff_B_u7AMRP7r4_2),.clk(gclk));
	jdff dff_B_FCrRxCp12_2(.din(w_dff_B_u7AMRP7r4_2),.dout(w_dff_B_FCrRxCp12_2),.clk(gclk));
	jdff dff_B_e9lWhaMh6_2(.din(w_dff_B_FCrRxCp12_2),.dout(w_dff_B_e9lWhaMh6_2),.clk(gclk));
	jdff dff_B_2Jin6f3F3_2(.din(w_dff_B_e9lWhaMh6_2),.dout(w_dff_B_2Jin6f3F3_2),.clk(gclk));
	jdff dff_B_8JFB5qkn8_2(.din(w_dff_B_2Jin6f3F3_2),.dout(w_dff_B_8JFB5qkn8_2),.clk(gclk));
	jdff dff_B_0EMXC8208_2(.din(w_dff_B_8JFB5qkn8_2),.dout(w_dff_B_0EMXC8208_2),.clk(gclk));
	jdff dff_B_NuzJ0KOO9_2(.din(w_dff_B_0EMXC8208_2),.dout(w_dff_B_NuzJ0KOO9_2),.clk(gclk));
	jdff dff_B_u46PCaA40_2(.din(w_dff_B_NuzJ0KOO9_2),.dout(w_dff_B_u46PCaA40_2),.clk(gclk));
	jdff dff_B_0ErCbtZ50_2(.din(w_dff_B_u46PCaA40_2),.dout(w_dff_B_0ErCbtZ50_2),.clk(gclk));
	jdff dff_B_uM9twtl81_2(.din(w_dff_B_0ErCbtZ50_2),.dout(w_dff_B_uM9twtl81_2),.clk(gclk));
	jdff dff_B_3LU7KrCG1_2(.din(w_dff_B_uM9twtl81_2),.dout(w_dff_B_3LU7KrCG1_2),.clk(gclk));
	jdff dff_B_Ql0WrQ9X9_2(.din(w_dff_B_3LU7KrCG1_2),.dout(w_dff_B_Ql0WrQ9X9_2),.clk(gclk));
	jdff dff_B_RkAULWx05_2(.din(w_dff_B_Ql0WrQ9X9_2),.dout(w_dff_B_RkAULWx05_2),.clk(gclk));
	jdff dff_B_6vocVvua1_2(.din(w_dff_B_RkAULWx05_2),.dout(w_dff_B_6vocVvua1_2),.clk(gclk));
	jdff dff_B_tW9KBL286_2(.din(w_dff_B_6vocVvua1_2),.dout(w_dff_B_tW9KBL286_2),.clk(gclk));
	jdff dff_B_ZyUpNRHt8_2(.din(w_dff_B_tW9KBL286_2),.dout(w_dff_B_ZyUpNRHt8_2),.clk(gclk));
	jdff dff_B_biC251xL4_2(.din(w_dff_B_ZyUpNRHt8_2),.dout(w_dff_B_biC251xL4_2),.clk(gclk));
	jdff dff_B_e92ZTNfs3_2(.din(w_dff_B_biC251xL4_2),.dout(w_dff_B_e92ZTNfs3_2),.clk(gclk));
	jdff dff_B_bNC18lju6_2(.din(w_dff_B_e92ZTNfs3_2),.dout(w_dff_B_bNC18lju6_2),.clk(gclk));
	jdff dff_B_cRmE4bC50_2(.din(w_dff_B_bNC18lju6_2),.dout(w_dff_B_cRmE4bC50_2),.clk(gclk));
	jdff dff_B_lfOlE06q1_2(.din(w_dff_B_cRmE4bC50_2),.dout(w_dff_B_lfOlE06q1_2),.clk(gclk));
	jdff dff_B_eoX6Bakl1_2(.din(w_dff_B_lfOlE06q1_2),.dout(w_dff_B_eoX6Bakl1_2),.clk(gclk));
	jdff dff_B_9TVjwXdf9_2(.din(w_dff_B_eoX6Bakl1_2),.dout(w_dff_B_9TVjwXdf9_2),.clk(gclk));
	jdff dff_B_YTqThHKS5_2(.din(w_dff_B_9TVjwXdf9_2),.dout(w_dff_B_YTqThHKS5_2),.clk(gclk));
	jdff dff_B_xlThTkhQ4_2(.din(w_dff_B_YTqThHKS5_2),.dout(w_dff_B_xlThTkhQ4_2),.clk(gclk));
	jdff dff_B_Nx0zpbCt3_2(.din(w_dff_B_xlThTkhQ4_2),.dout(w_dff_B_Nx0zpbCt3_2),.clk(gclk));
	jdff dff_B_bij20Ba39_2(.din(w_dff_B_Nx0zpbCt3_2),.dout(w_dff_B_bij20Ba39_2),.clk(gclk));
	jdff dff_B_C8CaNbL76_2(.din(w_dff_B_bij20Ba39_2),.dout(w_dff_B_C8CaNbL76_2),.clk(gclk));
	jdff dff_B_N5WoFur92_2(.din(w_dff_B_C8CaNbL76_2),.dout(w_dff_B_N5WoFur92_2),.clk(gclk));
	jdff dff_B_mZ5Xmqrh6_2(.din(w_dff_B_N5WoFur92_2),.dout(w_dff_B_mZ5Xmqrh6_2),.clk(gclk));
	jdff dff_B_0Ag6xAvX4_2(.din(w_dff_B_mZ5Xmqrh6_2),.dout(w_dff_B_0Ag6xAvX4_2),.clk(gclk));
	jdff dff_B_U0zwXmFV7_2(.din(w_dff_B_0Ag6xAvX4_2),.dout(w_dff_B_U0zwXmFV7_2),.clk(gclk));
	jdff dff_B_CuCPYtPz5_2(.din(w_dff_B_U0zwXmFV7_2),.dout(w_dff_B_CuCPYtPz5_2),.clk(gclk));
	jdff dff_B_pxy1iGAq9_2(.din(w_dff_B_CuCPYtPz5_2),.dout(w_dff_B_pxy1iGAq9_2),.clk(gclk));
	jdff dff_B_jR0iFg8K1_2(.din(w_dff_B_pxy1iGAq9_2),.dout(w_dff_B_jR0iFg8K1_2),.clk(gclk));
	jdff dff_B_1J0Cuqgg8_2(.din(w_dff_B_jR0iFg8K1_2),.dout(w_dff_B_1J0Cuqgg8_2),.clk(gclk));
	jdff dff_B_apvSUipR6_2(.din(w_dff_B_1J0Cuqgg8_2),.dout(w_dff_B_apvSUipR6_2),.clk(gclk));
	jdff dff_B_q7suo3Om0_2(.din(w_dff_B_apvSUipR6_2),.dout(w_dff_B_q7suo3Om0_2),.clk(gclk));
	jdff dff_B_So1lJT9J4_2(.din(w_dff_B_q7suo3Om0_2),.dout(w_dff_B_So1lJT9J4_2),.clk(gclk));
	jdff dff_B_UMZT43dn0_2(.din(w_dff_B_So1lJT9J4_2),.dout(w_dff_B_UMZT43dn0_2),.clk(gclk));
	jdff dff_B_KtAuF9hr8_2(.din(w_dff_B_UMZT43dn0_2),.dout(w_dff_B_KtAuF9hr8_2),.clk(gclk));
	jdff dff_B_yHuuOPrg8_2(.din(w_dff_B_KtAuF9hr8_2),.dout(w_dff_B_yHuuOPrg8_2),.clk(gclk));
	jdff dff_B_mHXheFJ27_2(.din(w_dff_B_yHuuOPrg8_2),.dout(w_dff_B_mHXheFJ27_2),.clk(gclk));
	jdff dff_B_0sLmQqVT3_1(.din(n1422),.dout(w_dff_B_0sLmQqVT3_1),.clk(gclk));
	jdff dff_B_5tJmI57P5_2(.din(n1343),.dout(w_dff_B_5tJmI57P5_2),.clk(gclk));
	jdff dff_B_9QME0q2B4_2(.din(w_dff_B_5tJmI57P5_2),.dout(w_dff_B_9QME0q2B4_2),.clk(gclk));
	jdff dff_B_7xhXWA223_2(.din(w_dff_B_9QME0q2B4_2),.dout(w_dff_B_7xhXWA223_2),.clk(gclk));
	jdff dff_B_dJOUgNBE3_2(.din(w_dff_B_7xhXWA223_2),.dout(w_dff_B_dJOUgNBE3_2),.clk(gclk));
	jdff dff_B_TwqBUNJx6_2(.din(w_dff_B_dJOUgNBE3_2),.dout(w_dff_B_TwqBUNJx6_2),.clk(gclk));
	jdff dff_B_OT7Snrp47_2(.din(w_dff_B_TwqBUNJx6_2),.dout(w_dff_B_OT7Snrp47_2),.clk(gclk));
	jdff dff_B_pDi4Wbia3_2(.din(w_dff_B_OT7Snrp47_2),.dout(w_dff_B_pDi4Wbia3_2),.clk(gclk));
	jdff dff_B_AUAjYsRO8_2(.din(w_dff_B_pDi4Wbia3_2),.dout(w_dff_B_AUAjYsRO8_2),.clk(gclk));
	jdff dff_B_2HlyQ3Bq3_2(.din(w_dff_B_AUAjYsRO8_2),.dout(w_dff_B_2HlyQ3Bq3_2),.clk(gclk));
	jdff dff_B_QDoAMHQW1_2(.din(w_dff_B_2HlyQ3Bq3_2),.dout(w_dff_B_QDoAMHQW1_2),.clk(gclk));
	jdff dff_B_kNc6j2k42_2(.din(w_dff_B_QDoAMHQW1_2),.dout(w_dff_B_kNc6j2k42_2),.clk(gclk));
	jdff dff_B_S9UkJYeo5_2(.din(w_dff_B_kNc6j2k42_2),.dout(w_dff_B_S9UkJYeo5_2),.clk(gclk));
	jdff dff_B_ullc4rfi4_2(.din(w_dff_B_S9UkJYeo5_2),.dout(w_dff_B_ullc4rfi4_2),.clk(gclk));
	jdff dff_B_IQtjO9Gk3_2(.din(w_dff_B_ullc4rfi4_2),.dout(w_dff_B_IQtjO9Gk3_2),.clk(gclk));
	jdff dff_B_wMJgVePA9_2(.din(w_dff_B_IQtjO9Gk3_2),.dout(w_dff_B_wMJgVePA9_2),.clk(gclk));
	jdff dff_B_z3dhxdxZ4_2(.din(w_dff_B_wMJgVePA9_2),.dout(w_dff_B_z3dhxdxZ4_2),.clk(gclk));
	jdff dff_B_h61JaaDv8_2(.din(w_dff_B_z3dhxdxZ4_2),.dout(w_dff_B_h61JaaDv8_2),.clk(gclk));
	jdff dff_B_2UEESRfr9_2(.din(w_dff_B_h61JaaDv8_2),.dout(w_dff_B_2UEESRfr9_2),.clk(gclk));
	jdff dff_B_tyLtbAUh7_2(.din(w_dff_B_2UEESRfr9_2),.dout(w_dff_B_tyLtbAUh7_2),.clk(gclk));
	jdff dff_B_ign3mPvn2_2(.din(w_dff_B_tyLtbAUh7_2),.dout(w_dff_B_ign3mPvn2_2),.clk(gclk));
	jdff dff_B_BKmplsR23_2(.din(w_dff_B_ign3mPvn2_2),.dout(w_dff_B_BKmplsR23_2),.clk(gclk));
	jdff dff_B_ACE7mfZj3_2(.din(w_dff_B_BKmplsR23_2),.dout(w_dff_B_ACE7mfZj3_2),.clk(gclk));
	jdff dff_B_7ilA3YS45_2(.din(w_dff_B_ACE7mfZj3_2),.dout(w_dff_B_7ilA3YS45_2),.clk(gclk));
	jdff dff_B_w5rh1REM0_2(.din(w_dff_B_7ilA3YS45_2),.dout(w_dff_B_w5rh1REM0_2),.clk(gclk));
	jdff dff_B_k3j7mOcY8_2(.din(w_dff_B_w5rh1REM0_2),.dout(w_dff_B_k3j7mOcY8_2),.clk(gclk));
	jdff dff_B_z5EWQJTw5_2(.din(w_dff_B_k3j7mOcY8_2),.dout(w_dff_B_z5EWQJTw5_2),.clk(gclk));
	jdff dff_B_FXUl9Wqj3_2(.din(w_dff_B_z5EWQJTw5_2),.dout(w_dff_B_FXUl9Wqj3_2),.clk(gclk));
	jdff dff_B_lt5yDCXU4_2(.din(w_dff_B_FXUl9Wqj3_2),.dout(w_dff_B_lt5yDCXU4_2),.clk(gclk));
	jdff dff_B_VAv23shb7_2(.din(w_dff_B_lt5yDCXU4_2),.dout(w_dff_B_VAv23shb7_2),.clk(gclk));
	jdff dff_B_iHuUAZne0_2(.din(w_dff_B_VAv23shb7_2),.dout(w_dff_B_iHuUAZne0_2),.clk(gclk));
	jdff dff_B_gHdQwUYq2_2(.din(w_dff_B_iHuUAZne0_2),.dout(w_dff_B_gHdQwUYq2_2),.clk(gclk));
	jdff dff_B_nQBWvc5R7_2(.din(w_dff_B_gHdQwUYq2_2),.dout(w_dff_B_nQBWvc5R7_2),.clk(gclk));
	jdff dff_B_10SL5MYS1_2(.din(w_dff_B_nQBWvc5R7_2),.dout(w_dff_B_10SL5MYS1_2),.clk(gclk));
	jdff dff_B_LWPKLSUN0_2(.din(w_dff_B_10SL5MYS1_2),.dout(w_dff_B_LWPKLSUN0_2),.clk(gclk));
	jdff dff_B_OOad25P37_2(.din(w_dff_B_LWPKLSUN0_2),.dout(w_dff_B_OOad25P37_2),.clk(gclk));
	jdff dff_B_RZEtVhtQ4_2(.din(w_dff_B_OOad25P37_2),.dout(w_dff_B_RZEtVhtQ4_2),.clk(gclk));
	jdff dff_B_Ayb7RcQF5_2(.din(w_dff_B_RZEtVhtQ4_2),.dout(w_dff_B_Ayb7RcQF5_2),.clk(gclk));
	jdff dff_B_GiRCWBgL6_2(.din(w_dff_B_Ayb7RcQF5_2),.dout(w_dff_B_GiRCWBgL6_2),.clk(gclk));
	jdff dff_B_GFOoJ2eq1_2(.din(w_dff_B_GiRCWBgL6_2),.dout(w_dff_B_GFOoJ2eq1_2),.clk(gclk));
	jdff dff_B_8QCyBW503_2(.din(w_dff_B_GFOoJ2eq1_2),.dout(w_dff_B_8QCyBW503_2),.clk(gclk));
	jdff dff_B_y92mo1M43_2(.din(w_dff_B_8QCyBW503_2),.dout(w_dff_B_y92mo1M43_2),.clk(gclk));
	jdff dff_B_bDocydhb6_1(.din(n1344),.dout(w_dff_B_bDocydhb6_1),.clk(gclk));
	jdff dff_B_Ail7x0LW9_2(.din(n1258),.dout(w_dff_B_Ail7x0LW9_2),.clk(gclk));
	jdff dff_B_xavbA5MR9_2(.din(w_dff_B_Ail7x0LW9_2),.dout(w_dff_B_xavbA5MR9_2),.clk(gclk));
	jdff dff_B_vHrddRzb8_2(.din(w_dff_B_xavbA5MR9_2),.dout(w_dff_B_vHrddRzb8_2),.clk(gclk));
	jdff dff_B_NJui82fM2_2(.din(w_dff_B_vHrddRzb8_2),.dout(w_dff_B_NJui82fM2_2),.clk(gclk));
	jdff dff_B_RskdySKq1_2(.din(w_dff_B_NJui82fM2_2),.dout(w_dff_B_RskdySKq1_2),.clk(gclk));
	jdff dff_B_hw3E776r6_2(.din(w_dff_B_RskdySKq1_2),.dout(w_dff_B_hw3E776r6_2),.clk(gclk));
	jdff dff_B_XIN9RZpx1_2(.din(w_dff_B_hw3E776r6_2),.dout(w_dff_B_XIN9RZpx1_2),.clk(gclk));
	jdff dff_B_d4Zgy1eJ0_2(.din(w_dff_B_XIN9RZpx1_2),.dout(w_dff_B_d4Zgy1eJ0_2),.clk(gclk));
	jdff dff_B_0NtEvgCP8_2(.din(w_dff_B_d4Zgy1eJ0_2),.dout(w_dff_B_0NtEvgCP8_2),.clk(gclk));
	jdff dff_B_RlnOtElS8_2(.din(w_dff_B_0NtEvgCP8_2),.dout(w_dff_B_RlnOtElS8_2),.clk(gclk));
	jdff dff_B_IfUQm2lL0_2(.din(w_dff_B_RlnOtElS8_2),.dout(w_dff_B_IfUQm2lL0_2),.clk(gclk));
	jdff dff_B_i5zHiUAi2_2(.din(w_dff_B_IfUQm2lL0_2),.dout(w_dff_B_i5zHiUAi2_2),.clk(gclk));
	jdff dff_B_KkSADCCF8_2(.din(w_dff_B_i5zHiUAi2_2),.dout(w_dff_B_KkSADCCF8_2),.clk(gclk));
	jdff dff_B_8g0Ewo7V6_2(.din(w_dff_B_KkSADCCF8_2),.dout(w_dff_B_8g0Ewo7V6_2),.clk(gclk));
	jdff dff_B_HSIJxpFC1_2(.din(w_dff_B_8g0Ewo7V6_2),.dout(w_dff_B_HSIJxpFC1_2),.clk(gclk));
	jdff dff_B_DAgV7bOd7_2(.din(w_dff_B_HSIJxpFC1_2),.dout(w_dff_B_DAgV7bOd7_2),.clk(gclk));
	jdff dff_B_dsajmSpj9_2(.din(w_dff_B_DAgV7bOd7_2),.dout(w_dff_B_dsajmSpj9_2),.clk(gclk));
	jdff dff_B_Pk4fXni59_2(.din(w_dff_B_dsajmSpj9_2),.dout(w_dff_B_Pk4fXni59_2),.clk(gclk));
	jdff dff_B_OVThfzDU0_2(.din(w_dff_B_Pk4fXni59_2),.dout(w_dff_B_OVThfzDU0_2),.clk(gclk));
	jdff dff_B_zWenA68s5_2(.din(w_dff_B_OVThfzDU0_2),.dout(w_dff_B_zWenA68s5_2),.clk(gclk));
	jdff dff_B_Eu3jSEHU6_2(.din(w_dff_B_zWenA68s5_2),.dout(w_dff_B_Eu3jSEHU6_2),.clk(gclk));
	jdff dff_B_RVVbgxur4_2(.din(w_dff_B_Eu3jSEHU6_2),.dout(w_dff_B_RVVbgxur4_2),.clk(gclk));
	jdff dff_B_DuuBdalP3_2(.din(w_dff_B_RVVbgxur4_2),.dout(w_dff_B_DuuBdalP3_2),.clk(gclk));
	jdff dff_B_REGAyUM73_2(.din(w_dff_B_DuuBdalP3_2),.dout(w_dff_B_REGAyUM73_2),.clk(gclk));
	jdff dff_B_a2ns7YfN0_2(.din(w_dff_B_REGAyUM73_2),.dout(w_dff_B_a2ns7YfN0_2),.clk(gclk));
	jdff dff_B_3fS8brj32_2(.din(w_dff_B_a2ns7YfN0_2),.dout(w_dff_B_3fS8brj32_2),.clk(gclk));
	jdff dff_B_Hgfq9Fns9_2(.din(w_dff_B_3fS8brj32_2),.dout(w_dff_B_Hgfq9Fns9_2),.clk(gclk));
	jdff dff_B_IOp36Eyd7_2(.din(w_dff_B_Hgfq9Fns9_2),.dout(w_dff_B_IOp36Eyd7_2),.clk(gclk));
	jdff dff_B_McR7QJ8w7_2(.din(w_dff_B_IOp36Eyd7_2),.dout(w_dff_B_McR7QJ8w7_2),.clk(gclk));
	jdff dff_B_xciPzj6d2_2(.din(w_dff_B_McR7QJ8w7_2),.dout(w_dff_B_xciPzj6d2_2),.clk(gclk));
	jdff dff_B_HCGnocdg4_2(.din(w_dff_B_xciPzj6d2_2),.dout(w_dff_B_HCGnocdg4_2),.clk(gclk));
	jdff dff_B_85Xw2VgO6_2(.din(w_dff_B_HCGnocdg4_2),.dout(w_dff_B_85Xw2VgO6_2),.clk(gclk));
	jdff dff_B_5voB3PvG2_2(.din(w_dff_B_85Xw2VgO6_2),.dout(w_dff_B_5voB3PvG2_2),.clk(gclk));
	jdff dff_B_mWk1ScFL8_2(.din(w_dff_B_5voB3PvG2_2),.dout(w_dff_B_mWk1ScFL8_2),.clk(gclk));
	jdff dff_B_Pg428fCG4_2(.din(w_dff_B_mWk1ScFL8_2),.dout(w_dff_B_Pg428fCG4_2),.clk(gclk));
	jdff dff_B_shBRayP63_2(.din(w_dff_B_Pg428fCG4_2),.dout(w_dff_B_shBRayP63_2),.clk(gclk));
	jdff dff_B_OTJVvwQm7_2(.din(w_dff_B_shBRayP63_2),.dout(w_dff_B_OTJVvwQm7_2),.clk(gclk));
	jdff dff_B_jqkbv9TZ6_2(.din(w_dff_B_OTJVvwQm7_2),.dout(w_dff_B_jqkbv9TZ6_2),.clk(gclk));
	jdff dff_B_zK7yrA7e2_1(.din(n1259),.dout(w_dff_B_zK7yrA7e2_1),.clk(gclk));
	jdff dff_B_7uyajVL02_2(.din(n1168),.dout(w_dff_B_7uyajVL02_2),.clk(gclk));
	jdff dff_B_aJI8Ek0i5_2(.din(w_dff_B_7uyajVL02_2),.dout(w_dff_B_aJI8Ek0i5_2),.clk(gclk));
	jdff dff_B_mlSvc89j3_2(.din(w_dff_B_aJI8Ek0i5_2),.dout(w_dff_B_mlSvc89j3_2),.clk(gclk));
	jdff dff_B_casXwag60_2(.din(w_dff_B_mlSvc89j3_2),.dout(w_dff_B_casXwag60_2),.clk(gclk));
	jdff dff_B_gtm8WN0E9_2(.din(w_dff_B_casXwag60_2),.dout(w_dff_B_gtm8WN0E9_2),.clk(gclk));
	jdff dff_B_8MCiHWbo3_2(.din(w_dff_B_gtm8WN0E9_2),.dout(w_dff_B_8MCiHWbo3_2),.clk(gclk));
	jdff dff_B_cYymuwiC9_2(.din(w_dff_B_8MCiHWbo3_2),.dout(w_dff_B_cYymuwiC9_2),.clk(gclk));
	jdff dff_B_9iBaMvuu7_2(.din(w_dff_B_cYymuwiC9_2),.dout(w_dff_B_9iBaMvuu7_2),.clk(gclk));
	jdff dff_B_PFTMqEUl0_2(.din(w_dff_B_9iBaMvuu7_2),.dout(w_dff_B_PFTMqEUl0_2),.clk(gclk));
	jdff dff_B_M8nr22Pk2_2(.din(w_dff_B_PFTMqEUl0_2),.dout(w_dff_B_M8nr22Pk2_2),.clk(gclk));
	jdff dff_B_D8TWBapD3_2(.din(w_dff_B_M8nr22Pk2_2),.dout(w_dff_B_D8TWBapD3_2),.clk(gclk));
	jdff dff_B_pbZqulTo2_2(.din(w_dff_B_D8TWBapD3_2),.dout(w_dff_B_pbZqulTo2_2),.clk(gclk));
	jdff dff_B_wMTcAZ8Y7_2(.din(w_dff_B_pbZqulTo2_2),.dout(w_dff_B_wMTcAZ8Y7_2),.clk(gclk));
	jdff dff_B_4tgce4Oe3_2(.din(w_dff_B_wMTcAZ8Y7_2),.dout(w_dff_B_4tgce4Oe3_2),.clk(gclk));
	jdff dff_B_B0kY7cIH1_2(.din(w_dff_B_4tgce4Oe3_2),.dout(w_dff_B_B0kY7cIH1_2),.clk(gclk));
	jdff dff_B_c076dEod8_2(.din(w_dff_B_B0kY7cIH1_2),.dout(w_dff_B_c076dEod8_2),.clk(gclk));
	jdff dff_B_5AyQ7Kps5_2(.din(w_dff_B_c076dEod8_2),.dout(w_dff_B_5AyQ7Kps5_2),.clk(gclk));
	jdff dff_B_zCdsglMz7_2(.din(w_dff_B_5AyQ7Kps5_2),.dout(w_dff_B_zCdsglMz7_2),.clk(gclk));
	jdff dff_B_7sk5J8Lk6_2(.din(w_dff_B_zCdsglMz7_2),.dout(w_dff_B_7sk5J8Lk6_2),.clk(gclk));
	jdff dff_B_3QNWTExY5_2(.din(w_dff_B_7sk5J8Lk6_2),.dout(w_dff_B_3QNWTExY5_2),.clk(gclk));
	jdff dff_B_CfXARsHa5_2(.din(w_dff_B_3QNWTExY5_2),.dout(w_dff_B_CfXARsHa5_2),.clk(gclk));
	jdff dff_B_UQzIMyu93_2(.din(w_dff_B_CfXARsHa5_2),.dout(w_dff_B_UQzIMyu93_2),.clk(gclk));
	jdff dff_B_I1spHyv23_2(.din(w_dff_B_UQzIMyu93_2),.dout(w_dff_B_I1spHyv23_2),.clk(gclk));
	jdff dff_B_iWjL12xB1_2(.din(w_dff_B_I1spHyv23_2),.dout(w_dff_B_iWjL12xB1_2),.clk(gclk));
	jdff dff_B_neoiNxse3_2(.din(w_dff_B_iWjL12xB1_2),.dout(w_dff_B_neoiNxse3_2),.clk(gclk));
	jdff dff_B_8FspEcO81_2(.din(w_dff_B_neoiNxse3_2),.dout(w_dff_B_8FspEcO81_2),.clk(gclk));
	jdff dff_B_8f7XQWKB3_2(.din(w_dff_B_8FspEcO81_2),.dout(w_dff_B_8f7XQWKB3_2),.clk(gclk));
	jdff dff_B_lALwfbKI4_2(.din(w_dff_B_8f7XQWKB3_2),.dout(w_dff_B_lALwfbKI4_2),.clk(gclk));
	jdff dff_B_m9RP6cwh6_2(.din(w_dff_B_lALwfbKI4_2),.dout(w_dff_B_m9RP6cwh6_2),.clk(gclk));
	jdff dff_B_SSSYWT8j9_2(.din(w_dff_B_m9RP6cwh6_2),.dout(w_dff_B_SSSYWT8j9_2),.clk(gclk));
	jdff dff_B_7VQRIbGZ3_2(.din(w_dff_B_SSSYWT8j9_2),.dout(w_dff_B_7VQRIbGZ3_2),.clk(gclk));
	jdff dff_B_V6QtCvTC6_2(.din(w_dff_B_7VQRIbGZ3_2),.dout(w_dff_B_V6QtCvTC6_2),.clk(gclk));
	jdff dff_B_WtOJPJKQ0_2(.din(w_dff_B_V6QtCvTC6_2),.dout(w_dff_B_WtOJPJKQ0_2),.clk(gclk));
	jdff dff_B_EDZ0dM3p1_2(.din(w_dff_B_WtOJPJKQ0_2),.dout(w_dff_B_EDZ0dM3p1_2),.clk(gclk));
	jdff dff_B_E2OoLQUy0_2(.din(w_dff_B_EDZ0dM3p1_2),.dout(w_dff_B_E2OoLQUy0_2),.clk(gclk));
	jdff dff_B_XCy6AqqE0_1(.din(n1169),.dout(w_dff_B_XCy6AqqE0_1),.clk(gclk));
	jdff dff_B_mOhtwAco6_2(.din(n1064),.dout(w_dff_B_mOhtwAco6_2),.clk(gclk));
	jdff dff_B_x0ipWgB22_2(.din(w_dff_B_mOhtwAco6_2),.dout(w_dff_B_x0ipWgB22_2),.clk(gclk));
	jdff dff_B_zf7ubohQ5_2(.din(w_dff_B_x0ipWgB22_2),.dout(w_dff_B_zf7ubohQ5_2),.clk(gclk));
	jdff dff_B_PeLc1mhz9_2(.din(w_dff_B_zf7ubohQ5_2),.dout(w_dff_B_PeLc1mhz9_2),.clk(gclk));
	jdff dff_B_whT14DNR7_2(.din(w_dff_B_PeLc1mhz9_2),.dout(w_dff_B_whT14DNR7_2),.clk(gclk));
	jdff dff_B_HWEOoNUW5_2(.din(w_dff_B_whT14DNR7_2),.dout(w_dff_B_HWEOoNUW5_2),.clk(gclk));
	jdff dff_B_VvaK21gh7_2(.din(w_dff_B_HWEOoNUW5_2),.dout(w_dff_B_VvaK21gh7_2),.clk(gclk));
	jdff dff_B_f7Ewsdfj0_2(.din(w_dff_B_VvaK21gh7_2),.dout(w_dff_B_f7Ewsdfj0_2),.clk(gclk));
	jdff dff_B_Uw2GXW670_2(.din(w_dff_B_f7Ewsdfj0_2),.dout(w_dff_B_Uw2GXW670_2),.clk(gclk));
	jdff dff_B_JoyZDAp41_2(.din(w_dff_B_Uw2GXW670_2),.dout(w_dff_B_JoyZDAp41_2),.clk(gclk));
	jdff dff_B_OKEVUuN66_2(.din(w_dff_B_JoyZDAp41_2),.dout(w_dff_B_OKEVUuN66_2),.clk(gclk));
	jdff dff_B_s2pdcjXa7_2(.din(w_dff_B_OKEVUuN66_2),.dout(w_dff_B_s2pdcjXa7_2),.clk(gclk));
	jdff dff_B_jPZTSIGX5_2(.din(w_dff_B_s2pdcjXa7_2),.dout(w_dff_B_jPZTSIGX5_2),.clk(gclk));
	jdff dff_B_sKgUjKXE1_2(.din(w_dff_B_jPZTSIGX5_2),.dout(w_dff_B_sKgUjKXE1_2),.clk(gclk));
	jdff dff_B_9PaQxmQP1_2(.din(w_dff_B_sKgUjKXE1_2),.dout(w_dff_B_9PaQxmQP1_2),.clk(gclk));
	jdff dff_B_ywhxro8M9_2(.din(w_dff_B_9PaQxmQP1_2),.dout(w_dff_B_ywhxro8M9_2),.clk(gclk));
	jdff dff_B_LptVu05a3_2(.din(w_dff_B_ywhxro8M9_2),.dout(w_dff_B_LptVu05a3_2),.clk(gclk));
	jdff dff_B_IuiQWMej4_2(.din(w_dff_B_LptVu05a3_2),.dout(w_dff_B_IuiQWMej4_2),.clk(gclk));
	jdff dff_B_fNhIjUJw6_2(.din(w_dff_B_IuiQWMej4_2),.dout(w_dff_B_fNhIjUJw6_2),.clk(gclk));
	jdff dff_B_OSaYeidp7_2(.din(w_dff_B_fNhIjUJw6_2),.dout(w_dff_B_OSaYeidp7_2),.clk(gclk));
	jdff dff_B_6Jqctgxu6_2(.din(w_dff_B_OSaYeidp7_2),.dout(w_dff_B_6Jqctgxu6_2),.clk(gclk));
	jdff dff_B_6vbSIVrz5_2(.din(w_dff_B_6Jqctgxu6_2),.dout(w_dff_B_6vbSIVrz5_2),.clk(gclk));
	jdff dff_B_hc25mcsi0_2(.din(w_dff_B_6vbSIVrz5_2),.dout(w_dff_B_hc25mcsi0_2),.clk(gclk));
	jdff dff_B_BHvM9pOO0_2(.din(w_dff_B_hc25mcsi0_2),.dout(w_dff_B_BHvM9pOO0_2),.clk(gclk));
	jdff dff_B_vZjccCfE4_2(.din(w_dff_B_BHvM9pOO0_2),.dout(w_dff_B_vZjccCfE4_2),.clk(gclk));
	jdff dff_B_KO3LgFCP8_2(.din(w_dff_B_vZjccCfE4_2),.dout(w_dff_B_KO3LgFCP8_2),.clk(gclk));
	jdff dff_B_K2se7K8b0_2(.din(w_dff_B_KO3LgFCP8_2),.dout(w_dff_B_K2se7K8b0_2),.clk(gclk));
	jdff dff_B_33bsCwZD8_2(.din(w_dff_B_K2se7K8b0_2),.dout(w_dff_B_33bsCwZD8_2),.clk(gclk));
	jdff dff_B_LPZAWkT82_2(.din(w_dff_B_33bsCwZD8_2),.dout(w_dff_B_LPZAWkT82_2),.clk(gclk));
	jdff dff_B_rdNKtdbr7_2(.din(w_dff_B_LPZAWkT82_2),.dout(w_dff_B_rdNKtdbr7_2),.clk(gclk));
	jdff dff_B_bzUD0DS71_2(.din(w_dff_B_rdNKtdbr7_2),.dout(w_dff_B_bzUD0DS71_2),.clk(gclk));
	jdff dff_B_NrD0JuhJ0_2(.din(w_dff_B_bzUD0DS71_2),.dout(w_dff_B_NrD0JuhJ0_2),.clk(gclk));
	jdff dff_B_oBxkf0G21_1(.din(n1065),.dout(w_dff_B_oBxkf0G21_1),.clk(gclk));
	jdff dff_B_nyQzncQx5_2(.din(n966),.dout(w_dff_B_nyQzncQx5_2),.clk(gclk));
	jdff dff_B_hENfEriK5_2(.din(w_dff_B_nyQzncQx5_2),.dout(w_dff_B_hENfEriK5_2),.clk(gclk));
	jdff dff_B_uC9fZBbf0_2(.din(w_dff_B_hENfEriK5_2),.dout(w_dff_B_uC9fZBbf0_2),.clk(gclk));
	jdff dff_B_95qiEZUQ9_2(.din(w_dff_B_uC9fZBbf0_2),.dout(w_dff_B_95qiEZUQ9_2),.clk(gclk));
	jdff dff_B_Q0983WCM7_2(.din(w_dff_B_95qiEZUQ9_2),.dout(w_dff_B_Q0983WCM7_2),.clk(gclk));
	jdff dff_B_t5DBuE1C2_2(.din(w_dff_B_Q0983WCM7_2),.dout(w_dff_B_t5DBuE1C2_2),.clk(gclk));
	jdff dff_B_xPq4QyHT7_2(.din(w_dff_B_t5DBuE1C2_2),.dout(w_dff_B_xPq4QyHT7_2),.clk(gclk));
	jdff dff_B_QnUdnQ4N2_2(.din(w_dff_B_xPq4QyHT7_2),.dout(w_dff_B_QnUdnQ4N2_2),.clk(gclk));
	jdff dff_B_DeNrO5LU5_2(.din(w_dff_B_QnUdnQ4N2_2),.dout(w_dff_B_DeNrO5LU5_2),.clk(gclk));
	jdff dff_B_lzcae39c3_2(.din(w_dff_B_DeNrO5LU5_2),.dout(w_dff_B_lzcae39c3_2),.clk(gclk));
	jdff dff_B_jjAg2ibS9_2(.din(w_dff_B_lzcae39c3_2),.dout(w_dff_B_jjAg2ibS9_2),.clk(gclk));
	jdff dff_B_HfQroRc54_2(.din(w_dff_B_jjAg2ibS9_2),.dout(w_dff_B_HfQroRc54_2),.clk(gclk));
	jdff dff_B_UnysazIq1_2(.din(w_dff_B_HfQroRc54_2),.dout(w_dff_B_UnysazIq1_2),.clk(gclk));
	jdff dff_B_B2BlSJOF6_2(.din(w_dff_B_UnysazIq1_2),.dout(w_dff_B_B2BlSJOF6_2),.clk(gclk));
	jdff dff_B_2ifCDld99_2(.din(w_dff_B_B2BlSJOF6_2),.dout(w_dff_B_2ifCDld99_2),.clk(gclk));
	jdff dff_B_KbyW8fFN2_2(.din(w_dff_B_2ifCDld99_2),.dout(w_dff_B_KbyW8fFN2_2),.clk(gclk));
	jdff dff_B_MPuTgbVK7_2(.din(w_dff_B_KbyW8fFN2_2),.dout(w_dff_B_MPuTgbVK7_2),.clk(gclk));
	jdff dff_B_tWotBzHZ0_2(.din(w_dff_B_MPuTgbVK7_2),.dout(w_dff_B_tWotBzHZ0_2),.clk(gclk));
	jdff dff_B_KeyjJanE4_2(.din(w_dff_B_tWotBzHZ0_2),.dout(w_dff_B_KeyjJanE4_2),.clk(gclk));
	jdff dff_B_zWDtDGxn6_2(.din(w_dff_B_KeyjJanE4_2),.dout(w_dff_B_zWDtDGxn6_2),.clk(gclk));
	jdff dff_B_DS3KBvOr0_2(.din(w_dff_B_zWDtDGxn6_2),.dout(w_dff_B_DS3KBvOr0_2),.clk(gclk));
	jdff dff_B_CG1L7VNh1_2(.din(w_dff_B_DS3KBvOr0_2),.dout(w_dff_B_CG1L7VNh1_2),.clk(gclk));
	jdff dff_B_zhuitS4c0_2(.din(w_dff_B_CG1L7VNh1_2),.dout(w_dff_B_zhuitS4c0_2),.clk(gclk));
	jdff dff_B_V8xvLMEC0_2(.din(w_dff_B_zhuitS4c0_2),.dout(w_dff_B_V8xvLMEC0_2),.clk(gclk));
	jdff dff_B_1mwnz31j4_2(.din(w_dff_B_V8xvLMEC0_2),.dout(w_dff_B_1mwnz31j4_2),.clk(gclk));
	jdff dff_B_o8JfBlew1_2(.din(w_dff_B_1mwnz31j4_2),.dout(w_dff_B_o8JfBlew1_2),.clk(gclk));
	jdff dff_B_NnywUvYP6_2(.din(w_dff_B_o8JfBlew1_2),.dout(w_dff_B_NnywUvYP6_2),.clk(gclk));
	jdff dff_B_AJzwcfb63_2(.din(w_dff_B_NnywUvYP6_2),.dout(w_dff_B_AJzwcfb63_2),.clk(gclk));
	jdff dff_B_JKhRRn0h9_2(.din(w_dff_B_AJzwcfb63_2),.dout(w_dff_B_JKhRRn0h9_2),.clk(gclk));
	jdff dff_B_E28e5hOE1_1(.din(n967),.dout(w_dff_B_E28e5hOE1_1),.clk(gclk));
	jdff dff_B_XOMImEQL4_2(.din(n861),.dout(w_dff_B_XOMImEQL4_2),.clk(gclk));
	jdff dff_B_qGKIcVa97_2(.din(w_dff_B_XOMImEQL4_2),.dout(w_dff_B_qGKIcVa97_2),.clk(gclk));
	jdff dff_B_HqFOYD4u0_2(.din(w_dff_B_qGKIcVa97_2),.dout(w_dff_B_HqFOYD4u0_2),.clk(gclk));
	jdff dff_B_lcSgrEP82_2(.din(w_dff_B_HqFOYD4u0_2),.dout(w_dff_B_lcSgrEP82_2),.clk(gclk));
	jdff dff_B_AljT9tO11_2(.din(w_dff_B_lcSgrEP82_2),.dout(w_dff_B_AljT9tO11_2),.clk(gclk));
	jdff dff_B_FruXNmDq8_2(.din(w_dff_B_AljT9tO11_2),.dout(w_dff_B_FruXNmDq8_2),.clk(gclk));
	jdff dff_B_3603w8rk5_2(.din(w_dff_B_FruXNmDq8_2),.dout(w_dff_B_3603w8rk5_2),.clk(gclk));
	jdff dff_B_OFuueyCD7_2(.din(w_dff_B_3603w8rk5_2),.dout(w_dff_B_OFuueyCD7_2),.clk(gclk));
	jdff dff_B_Oi6COfNE5_2(.din(w_dff_B_OFuueyCD7_2),.dout(w_dff_B_Oi6COfNE5_2),.clk(gclk));
	jdff dff_B_Ku37XT687_2(.din(w_dff_B_Oi6COfNE5_2),.dout(w_dff_B_Ku37XT687_2),.clk(gclk));
	jdff dff_B_5IOc2Odm5_2(.din(w_dff_B_Ku37XT687_2),.dout(w_dff_B_5IOc2Odm5_2),.clk(gclk));
	jdff dff_B_KSCjAnzz0_2(.din(w_dff_B_5IOc2Odm5_2),.dout(w_dff_B_KSCjAnzz0_2),.clk(gclk));
	jdff dff_B_k0txzxyL3_2(.din(w_dff_B_KSCjAnzz0_2),.dout(w_dff_B_k0txzxyL3_2),.clk(gclk));
	jdff dff_B_P8ezx6NU1_2(.din(w_dff_B_k0txzxyL3_2),.dout(w_dff_B_P8ezx6NU1_2),.clk(gclk));
	jdff dff_B_SaaKk0rA0_2(.din(w_dff_B_P8ezx6NU1_2),.dout(w_dff_B_SaaKk0rA0_2),.clk(gclk));
	jdff dff_B_B717Sm6c3_2(.din(w_dff_B_SaaKk0rA0_2),.dout(w_dff_B_B717Sm6c3_2),.clk(gclk));
	jdff dff_B_m7ZYFU6e0_2(.din(w_dff_B_B717Sm6c3_2),.dout(w_dff_B_m7ZYFU6e0_2),.clk(gclk));
	jdff dff_B_uAifJrff4_2(.din(w_dff_B_m7ZYFU6e0_2),.dout(w_dff_B_uAifJrff4_2),.clk(gclk));
	jdff dff_B_SGZ4B0SC9_2(.din(w_dff_B_uAifJrff4_2),.dout(w_dff_B_SGZ4B0SC9_2),.clk(gclk));
	jdff dff_B_Yl81yMHH5_2(.din(w_dff_B_SGZ4B0SC9_2),.dout(w_dff_B_Yl81yMHH5_2),.clk(gclk));
	jdff dff_B_pB7p2nKL1_2(.din(w_dff_B_Yl81yMHH5_2),.dout(w_dff_B_pB7p2nKL1_2),.clk(gclk));
	jdff dff_B_KtKs2P754_2(.din(w_dff_B_pB7p2nKL1_2),.dout(w_dff_B_KtKs2P754_2),.clk(gclk));
	jdff dff_B_Bdt25Oma6_2(.din(w_dff_B_KtKs2P754_2),.dout(w_dff_B_Bdt25Oma6_2),.clk(gclk));
	jdff dff_B_liaGK4Oh9_2(.din(w_dff_B_Bdt25Oma6_2),.dout(w_dff_B_liaGK4Oh9_2),.clk(gclk));
	jdff dff_B_753rPRre9_2(.din(w_dff_B_liaGK4Oh9_2),.dout(w_dff_B_753rPRre9_2),.clk(gclk));
	jdff dff_B_OIsxnejw5_2(.din(w_dff_B_753rPRre9_2),.dout(w_dff_B_OIsxnejw5_2),.clk(gclk));
	jdff dff_B_BjPK4aKx5_1(.din(n862),.dout(w_dff_B_BjPK4aKx5_1),.clk(gclk));
	jdff dff_B_DMqxYSwQ6_2(.din(n762),.dout(w_dff_B_DMqxYSwQ6_2),.clk(gclk));
	jdff dff_B_Z2s64YQC9_2(.din(w_dff_B_DMqxYSwQ6_2),.dout(w_dff_B_Z2s64YQC9_2),.clk(gclk));
	jdff dff_B_cuSyWlnS8_2(.din(w_dff_B_Z2s64YQC9_2),.dout(w_dff_B_cuSyWlnS8_2),.clk(gclk));
	jdff dff_B_Nbzw6ON34_2(.din(w_dff_B_cuSyWlnS8_2),.dout(w_dff_B_Nbzw6ON34_2),.clk(gclk));
	jdff dff_B_HH89iHAK3_2(.din(w_dff_B_Nbzw6ON34_2),.dout(w_dff_B_HH89iHAK3_2),.clk(gclk));
	jdff dff_B_C6LyLxPP1_2(.din(w_dff_B_HH89iHAK3_2),.dout(w_dff_B_C6LyLxPP1_2),.clk(gclk));
	jdff dff_B_hcv6tpdE9_2(.din(w_dff_B_C6LyLxPP1_2),.dout(w_dff_B_hcv6tpdE9_2),.clk(gclk));
	jdff dff_B_0szlR8g17_2(.din(w_dff_B_hcv6tpdE9_2),.dout(w_dff_B_0szlR8g17_2),.clk(gclk));
	jdff dff_B_ArXzfoTA0_2(.din(w_dff_B_0szlR8g17_2),.dout(w_dff_B_ArXzfoTA0_2),.clk(gclk));
	jdff dff_B_1B7dMboQ7_2(.din(w_dff_B_ArXzfoTA0_2),.dout(w_dff_B_1B7dMboQ7_2),.clk(gclk));
	jdff dff_B_a5FZGSEl5_2(.din(w_dff_B_1B7dMboQ7_2),.dout(w_dff_B_a5FZGSEl5_2),.clk(gclk));
	jdff dff_B_0Yhipu7D7_2(.din(w_dff_B_a5FZGSEl5_2),.dout(w_dff_B_0Yhipu7D7_2),.clk(gclk));
	jdff dff_B_1NUpT4y28_2(.din(w_dff_B_0Yhipu7D7_2),.dout(w_dff_B_1NUpT4y28_2),.clk(gclk));
	jdff dff_B_8xQEpUDT5_2(.din(w_dff_B_1NUpT4y28_2),.dout(w_dff_B_8xQEpUDT5_2),.clk(gclk));
	jdff dff_B_P6n3vYq81_2(.din(w_dff_B_8xQEpUDT5_2),.dout(w_dff_B_P6n3vYq81_2),.clk(gclk));
	jdff dff_B_p5tsQIBi6_2(.din(w_dff_B_P6n3vYq81_2),.dout(w_dff_B_p5tsQIBi6_2),.clk(gclk));
	jdff dff_B_LuONwujo3_2(.din(w_dff_B_p5tsQIBi6_2),.dout(w_dff_B_LuONwujo3_2),.clk(gclk));
	jdff dff_B_kvuIYBN82_2(.din(w_dff_B_LuONwujo3_2),.dout(w_dff_B_kvuIYBN82_2),.clk(gclk));
	jdff dff_B_B1AggMv63_2(.din(w_dff_B_kvuIYBN82_2),.dout(w_dff_B_B1AggMv63_2),.clk(gclk));
	jdff dff_B_6AdCB4FG6_2(.din(w_dff_B_B1AggMv63_2),.dout(w_dff_B_6AdCB4FG6_2),.clk(gclk));
	jdff dff_B_LLHzkkIu4_2(.din(w_dff_B_6AdCB4FG6_2),.dout(w_dff_B_LLHzkkIu4_2),.clk(gclk));
	jdff dff_B_xGKzri6L1_2(.din(w_dff_B_LLHzkkIu4_2),.dout(w_dff_B_xGKzri6L1_2),.clk(gclk));
	jdff dff_B_ZHXhiKye4_2(.din(w_dff_B_xGKzri6L1_2),.dout(w_dff_B_ZHXhiKye4_2),.clk(gclk));
	jdff dff_B_OItvkCtj8_1(.din(n763),.dout(w_dff_B_OItvkCtj8_1),.clk(gclk));
	jdff dff_B_9iip8WQh6_2(.din(n669),.dout(w_dff_B_9iip8WQh6_2),.clk(gclk));
	jdff dff_B_UZ6QsmhZ9_2(.din(w_dff_B_9iip8WQh6_2),.dout(w_dff_B_UZ6QsmhZ9_2),.clk(gclk));
	jdff dff_B_CN2r3IKi5_2(.din(w_dff_B_UZ6QsmhZ9_2),.dout(w_dff_B_CN2r3IKi5_2),.clk(gclk));
	jdff dff_B_55AyiywL1_2(.din(w_dff_B_CN2r3IKi5_2),.dout(w_dff_B_55AyiywL1_2),.clk(gclk));
	jdff dff_B_sR5FerlT7_2(.din(w_dff_B_55AyiywL1_2),.dout(w_dff_B_sR5FerlT7_2),.clk(gclk));
	jdff dff_B_8geRG4Xy3_2(.din(w_dff_B_sR5FerlT7_2),.dout(w_dff_B_8geRG4Xy3_2),.clk(gclk));
	jdff dff_B_DePmAgkt6_2(.din(w_dff_B_8geRG4Xy3_2),.dout(w_dff_B_DePmAgkt6_2),.clk(gclk));
	jdff dff_B_iU6G1aGu4_2(.din(w_dff_B_DePmAgkt6_2),.dout(w_dff_B_iU6G1aGu4_2),.clk(gclk));
	jdff dff_B_FqTiiNcf0_2(.din(w_dff_B_iU6G1aGu4_2),.dout(w_dff_B_FqTiiNcf0_2),.clk(gclk));
	jdff dff_B_QEpK86Ut0_2(.din(w_dff_B_FqTiiNcf0_2),.dout(w_dff_B_QEpK86Ut0_2),.clk(gclk));
	jdff dff_B_T56r6L5y9_2(.din(w_dff_B_QEpK86Ut0_2),.dout(w_dff_B_T56r6L5y9_2),.clk(gclk));
	jdff dff_B_P48ZY4Fs4_2(.din(w_dff_B_T56r6L5y9_2),.dout(w_dff_B_P48ZY4Fs4_2),.clk(gclk));
	jdff dff_B_Bjh8NZoH4_2(.din(w_dff_B_P48ZY4Fs4_2),.dout(w_dff_B_Bjh8NZoH4_2),.clk(gclk));
	jdff dff_B_BUMgbZW81_2(.din(w_dff_B_Bjh8NZoH4_2),.dout(w_dff_B_BUMgbZW81_2),.clk(gclk));
	jdff dff_B_Czt1wo8U3_2(.din(w_dff_B_BUMgbZW81_2),.dout(w_dff_B_Czt1wo8U3_2),.clk(gclk));
	jdff dff_B_YvoKr5Zw3_2(.din(w_dff_B_Czt1wo8U3_2),.dout(w_dff_B_YvoKr5Zw3_2),.clk(gclk));
	jdff dff_B_LcymxrAF2_2(.din(w_dff_B_YvoKr5Zw3_2),.dout(w_dff_B_LcymxrAF2_2),.clk(gclk));
	jdff dff_B_jrHV2jSQ8_2(.din(w_dff_B_LcymxrAF2_2),.dout(w_dff_B_jrHV2jSQ8_2),.clk(gclk));
	jdff dff_B_CPoqtNDM3_2(.din(w_dff_B_jrHV2jSQ8_2),.dout(w_dff_B_CPoqtNDM3_2),.clk(gclk));
	jdff dff_B_gvaO9FrA4_2(.din(w_dff_B_CPoqtNDM3_2),.dout(w_dff_B_gvaO9FrA4_2),.clk(gclk));
	jdff dff_B_wUqJfUUX3_1(.din(n670),.dout(w_dff_B_wUqJfUUX3_1),.clk(gclk));
	jdff dff_B_kFLC2GR77_2(.din(n583),.dout(w_dff_B_kFLC2GR77_2),.clk(gclk));
	jdff dff_B_TIqJxy468_2(.din(w_dff_B_kFLC2GR77_2),.dout(w_dff_B_TIqJxy468_2),.clk(gclk));
	jdff dff_B_68EIUyMI6_2(.din(w_dff_B_TIqJxy468_2),.dout(w_dff_B_68EIUyMI6_2),.clk(gclk));
	jdff dff_B_d73FkaNb1_2(.din(w_dff_B_68EIUyMI6_2),.dout(w_dff_B_d73FkaNb1_2),.clk(gclk));
	jdff dff_B_rswHVzdp1_2(.din(w_dff_B_d73FkaNb1_2),.dout(w_dff_B_rswHVzdp1_2),.clk(gclk));
	jdff dff_B_yGhtyHuM2_2(.din(w_dff_B_rswHVzdp1_2),.dout(w_dff_B_yGhtyHuM2_2),.clk(gclk));
	jdff dff_B_H36rjuGp4_2(.din(w_dff_B_yGhtyHuM2_2),.dout(w_dff_B_H36rjuGp4_2),.clk(gclk));
	jdff dff_B_NPyD8V6Q4_2(.din(w_dff_B_H36rjuGp4_2),.dout(w_dff_B_NPyD8V6Q4_2),.clk(gclk));
	jdff dff_B_kkvFLeXN6_2(.din(w_dff_B_NPyD8V6Q4_2),.dout(w_dff_B_kkvFLeXN6_2),.clk(gclk));
	jdff dff_B_MOs6bbNg7_2(.din(w_dff_B_kkvFLeXN6_2),.dout(w_dff_B_MOs6bbNg7_2),.clk(gclk));
	jdff dff_B_XgJLOM088_2(.din(w_dff_B_MOs6bbNg7_2),.dout(w_dff_B_XgJLOM088_2),.clk(gclk));
	jdff dff_B_Jqb2q0UQ9_2(.din(w_dff_B_XgJLOM088_2),.dout(w_dff_B_Jqb2q0UQ9_2),.clk(gclk));
	jdff dff_B_23u9yKB51_2(.din(w_dff_B_Jqb2q0UQ9_2),.dout(w_dff_B_23u9yKB51_2),.clk(gclk));
	jdff dff_B_vFV6DZay9_2(.din(w_dff_B_23u9yKB51_2),.dout(w_dff_B_vFV6DZay9_2),.clk(gclk));
	jdff dff_B_ljWA7UnI5_2(.din(w_dff_B_vFV6DZay9_2),.dout(w_dff_B_ljWA7UnI5_2),.clk(gclk));
	jdff dff_B_oIEOGCbR3_2(.din(w_dff_B_ljWA7UnI5_2),.dout(w_dff_B_oIEOGCbR3_2),.clk(gclk));
	jdff dff_B_FnvGQ8Bn4_2(.din(w_dff_B_oIEOGCbR3_2),.dout(w_dff_B_FnvGQ8Bn4_2),.clk(gclk));
	jdff dff_B_fglGzeOF8_1(.din(n584),.dout(w_dff_B_fglGzeOF8_1),.clk(gclk));
	jdff dff_B_GmEdFwzt9_2(.din(n504),.dout(w_dff_B_GmEdFwzt9_2),.clk(gclk));
	jdff dff_B_Wet41jYg8_2(.din(w_dff_B_GmEdFwzt9_2),.dout(w_dff_B_Wet41jYg8_2),.clk(gclk));
	jdff dff_B_0IM08Xhr6_2(.din(w_dff_B_Wet41jYg8_2),.dout(w_dff_B_0IM08Xhr6_2),.clk(gclk));
	jdff dff_B_Nm7ohPpE8_2(.din(w_dff_B_0IM08Xhr6_2),.dout(w_dff_B_Nm7ohPpE8_2),.clk(gclk));
	jdff dff_B_799TdZwW8_2(.din(w_dff_B_Nm7ohPpE8_2),.dout(w_dff_B_799TdZwW8_2),.clk(gclk));
	jdff dff_B_RCFvNIZR1_2(.din(w_dff_B_799TdZwW8_2),.dout(w_dff_B_RCFvNIZR1_2),.clk(gclk));
	jdff dff_B_FSi5VrUN6_2(.din(w_dff_B_RCFvNIZR1_2),.dout(w_dff_B_FSi5VrUN6_2),.clk(gclk));
	jdff dff_B_QZz8XZda1_2(.din(w_dff_B_FSi5VrUN6_2),.dout(w_dff_B_QZz8XZda1_2),.clk(gclk));
	jdff dff_B_WZuxoPR85_2(.din(w_dff_B_QZz8XZda1_2),.dout(w_dff_B_WZuxoPR85_2),.clk(gclk));
	jdff dff_B_PXzCCsIk5_2(.din(w_dff_B_WZuxoPR85_2),.dout(w_dff_B_PXzCCsIk5_2),.clk(gclk));
	jdff dff_B_IaG5tIM03_2(.din(w_dff_B_PXzCCsIk5_2),.dout(w_dff_B_IaG5tIM03_2),.clk(gclk));
	jdff dff_B_EZJV2KLH4_2(.din(w_dff_B_IaG5tIM03_2),.dout(w_dff_B_EZJV2KLH4_2),.clk(gclk));
	jdff dff_B_g1cfKTTf9_2(.din(w_dff_B_EZJV2KLH4_2),.dout(w_dff_B_g1cfKTTf9_2),.clk(gclk));
	jdff dff_B_teV2fcSQ9_2(.din(w_dff_B_g1cfKTTf9_2),.dout(w_dff_B_teV2fcSQ9_2),.clk(gclk));
	jdff dff_B_Vf2dWUQs7_1(.din(n505),.dout(w_dff_B_Vf2dWUQs7_1),.clk(gclk));
	jdff dff_B_cMyEysnW7_2(.din(n432),.dout(w_dff_B_cMyEysnW7_2),.clk(gclk));
	jdff dff_B_ZS1GBwxJ1_2(.din(w_dff_B_cMyEysnW7_2),.dout(w_dff_B_ZS1GBwxJ1_2),.clk(gclk));
	jdff dff_B_z8q1Xxtq9_2(.din(w_dff_B_ZS1GBwxJ1_2),.dout(w_dff_B_z8q1Xxtq9_2),.clk(gclk));
	jdff dff_B_88FlmuEy4_2(.din(w_dff_B_z8q1Xxtq9_2),.dout(w_dff_B_88FlmuEy4_2),.clk(gclk));
	jdff dff_B_C0jFK4sV5_2(.din(w_dff_B_88FlmuEy4_2),.dout(w_dff_B_C0jFK4sV5_2),.clk(gclk));
	jdff dff_B_A58XZpTV7_2(.din(w_dff_B_C0jFK4sV5_2),.dout(w_dff_B_A58XZpTV7_2),.clk(gclk));
	jdff dff_B_kPCrZGqh9_2(.din(w_dff_B_A58XZpTV7_2),.dout(w_dff_B_kPCrZGqh9_2),.clk(gclk));
	jdff dff_B_9eO8g0EC0_2(.din(w_dff_B_kPCrZGqh9_2),.dout(w_dff_B_9eO8g0EC0_2),.clk(gclk));
	jdff dff_B_Bb2lQgUJ4_2(.din(w_dff_B_9eO8g0EC0_2),.dout(w_dff_B_Bb2lQgUJ4_2),.clk(gclk));
	jdff dff_B_xj0jtopr1_2(.din(w_dff_B_Bb2lQgUJ4_2),.dout(w_dff_B_xj0jtopr1_2),.clk(gclk));
	jdff dff_B_mcltNOjw8_2(.din(w_dff_B_xj0jtopr1_2),.dout(w_dff_B_mcltNOjw8_2),.clk(gclk));
	jdff dff_B_qWfI2QVG8_2(.din(n435),.dout(w_dff_B_qWfI2QVG8_2),.clk(gclk));
	jdff dff_B_Q5Fcfau46_1(.din(n433),.dout(w_dff_B_Q5Fcfau46_1),.clk(gclk));
	jdff dff_B_U2vHbwWV2_2(.din(n368),.dout(w_dff_B_U2vHbwWV2_2),.clk(gclk));
	jdff dff_B_4MUSLB1k8_2(.din(w_dff_B_U2vHbwWV2_2),.dout(w_dff_B_4MUSLB1k8_2),.clk(gclk));
	jdff dff_B_cJrien2v6_2(.din(w_dff_B_4MUSLB1k8_2),.dout(w_dff_B_cJrien2v6_2),.clk(gclk));
	jdff dff_B_yGpplbgN8_2(.din(w_dff_B_cJrien2v6_2),.dout(w_dff_B_yGpplbgN8_2),.clk(gclk));
	jdff dff_B_oeqtDQfZ4_2(.din(w_dff_B_yGpplbgN8_2),.dout(w_dff_B_oeqtDQfZ4_2),.clk(gclk));
	jdff dff_B_P2HwkiEj0_2(.din(w_dff_B_oeqtDQfZ4_2),.dout(w_dff_B_P2HwkiEj0_2),.clk(gclk));
	jdff dff_B_BeecgaRi2_2(.din(w_dff_B_P2HwkiEj0_2),.dout(w_dff_B_BeecgaRi2_2),.clk(gclk));
	jdff dff_B_frfc0sZl2_1(.din(n369),.dout(w_dff_B_frfc0sZl2_1),.clk(gclk));
	jdff dff_B_kEXGgwSC7_2(.din(n310),.dout(w_dff_B_kEXGgwSC7_2),.clk(gclk));
	jdff dff_B_u817jq6I1_2(.din(w_dff_B_kEXGgwSC7_2),.dout(w_dff_B_u817jq6I1_2),.clk(gclk));
	jdff dff_B_hT7sTadY8_2(.din(w_dff_B_u817jq6I1_2),.dout(w_dff_B_hT7sTadY8_2),.clk(gclk));
	jdff dff_B_Vr0RTiuP0_2(.din(w_dff_B_hT7sTadY8_2),.dout(w_dff_B_Vr0RTiuP0_2),.clk(gclk));
	jdff dff_B_oBTVm2AH7_1(.din(n312),.dout(w_dff_B_oBTVm2AH7_1),.clk(gclk));
	jdff dff_A_AvuFHgdL3_0(.dout(w_n258_0[0]),.din(w_dff_A_AvuFHgdL3_0),.clk(gclk));
	jdff dff_A_7C2puQDr9_1(.dout(w_n258_0[1]),.din(w_dff_A_7C2puQDr9_1),.clk(gclk));
	jdff dff_A_jWxdfK7Z8_1(.dout(w_dff_A_7C2puQDr9_1),.din(w_dff_A_jWxdfK7Z8_1),.clk(gclk));
	jdff dff_B_a7Ek4TkY8_1(.din(n1563),.dout(w_dff_B_a7Ek4TkY8_1),.clk(gclk));
	jdff dff_B_6OiQ7KOP5_2(.din(n1497),.dout(w_dff_B_6OiQ7KOP5_2),.clk(gclk));
	jdff dff_B_VAkpoyWb1_2(.din(w_dff_B_6OiQ7KOP5_2),.dout(w_dff_B_VAkpoyWb1_2),.clk(gclk));
	jdff dff_B_JxIrZkrD4_2(.din(w_dff_B_VAkpoyWb1_2),.dout(w_dff_B_JxIrZkrD4_2),.clk(gclk));
	jdff dff_B_iQLfoj5c4_2(.din(w_dff_B_JxIrZkrD4_2),.dout(w_dff_B_iQLfoj5c4_2),.clk(gclk));
	jdff dff_B_YxIZrGR83_2(.din(w_dff_B_iQLfoj5c4_2),.dout(w_dff_B_YxIZrGR83_2),.clk(gclk));
	jdff dff_B_o6gtRhGj2_2(.din(w_dff_B_YxIZrGR83_2),.dout(w_dff_B_o6gtRhGj2_2),.clk(gclk));
	jdff dff_B_TW9KYJLO6_2(.din(w_dff_B_o6gtRhGj2_2),.dout(w_dff_B_TW9KYJLO6_2),.clk(gclk));
	jdff dff_B_k6VH2Q193_2(.din(w_dff_B_TW9KYJLO6_2),.dout(w_dff_B_k6VH2Q193_2),.clk(gclk));
	jdff dff_B_25UzyUww6_2(.din(w_dff_B_k6VH2Q193_2),.dout(w_dff_B_25UzyUww6_2),.clk(gclk));
	jdff dff_B_6km1JTS97_2(.din(w_dff_B_25UzyUww6_2),.dout(w_dff_B_6km1JTS97_2),.clk(gclk));
	jdff dff_B_VKnZfUOf9_2(.din(w_dff_B_6km1JTS97_2),.dout(w_dff_B_VKnZfUOf9_2),.clk(gclk));
	jdff dff_B_38KD7hC70_2(.din(w_dff_B_VKnZfUOf9_2),.dout(w_dff_B_38KD7hC70_2),.clk(gclk));
	jdff dff_B_b8etlaOw9_2(.din(w_dff_B_38KD7hC70_2),.dout(w_dff_B_b8etlaOw9_2),.clk(gclk));
	jdff dff_B_hjrHoEkS4_2(.din(w_dff_B_b8etlaOw9_2),.dout(w_dff_B_hjrHoEkS4_2),.clk(gclk));
	jdff dff_B_kEykrjUL0_2(.din(w_dff_B_hjrHoEkS4_2),.dout(w_dff_B_kEykrjUL0_2),.clk(gclk));
	jdff dff_B_vq3QEiX60_2(.din(w_dff_B_kEykrjUL0_2),.dout(w_dff_B_vq3QEiX60_2),.clk(gclk));
	jdff dff_B_EnuqSSC76_2(.din(w_dff_B_vq3QEiX60_2),.dout(w_dff_B_EnuqSSC76_2),.clk(gclk));
	jdff dff_B_RyGsuda15_2(.din(w_dff_B_EnuqSSC76_2),.dout(w_dff_B_RyGsuda15_2),.clk(gclk));
	jdff dff_B_gXBYITOv9_2(.din(w_dff_B_RyGsuda15_2),.dout(w_dff_B_gXBYITOv9_2),.clk(gclk));
	jdff dff_B_s8ONbQNv6_2(.din(w_dff_B_gXBYITOv9_2),.dout(w_dff_B_s8ONbQNv6_2),.clk(gclk));
	jdff dff_B_wGlfMzgV9_2(.din(w_dff_B_s8ONbQNv6_2),.dout(w_dff_B_wGlfMzgV9_2),.clk(gclk));
	jdff dff_B_zYRG2Gs04_2(.din(w_dff_B_wGlfMzgV9_2),.dout(w_dff_B_zYRG2Gs04_2),.clk(gclk));
	jdff dff_B_c91Sn8wm0_2(.din(w_dff_B_zYRG2Gs04_2),.dout(w_dff_B_c91Sn8wm0_2),.clk(gclk));
	jdff dff_B_eus8bNGi7_2(.din(w_dff_B_c91Sn8wm0_2),.dout(w_dff_B_eus8bNGi7_2),.clk(gclk));
	jdff dff_B_w9D4qMMB1_2(.din(w_dff_B_eus8bNGi7_2),.dout(w_dff_B_w9D4qMMB1_2),.clk(gclk));
	jdff dff_B_AxNKrLfK5_2(.din(w_dff_B_w9D4qMMB1_2),.dout(w_dff_B_AxNKrLfK5_2),.clk(gclk));
	jdff dff_B_j7ItMyId4_2(.din(w_dff_B_AxNKrLfK5_2),.dout(w_dff_B_j7ItMyId4_2),.clk(gclk));
	jdff dff_B_fiq6Y3Uz5_2(.din(w_dff_B_j7ItMyId4_2),.dout(w_dff_B_fiq6Y3Uz5_2),.clk(gclk));
	jdff dff_B_Ehj2jM1H8_2(.din(w_dff_B_fiq6Y3Uz5_2),.dout(w_dff_B_Ehj2jM1H8_2),.clk(gclk));
	jdff dff_B_XxuADOnt9_2(.din(w_dff_B_Ehj2jM1H8_2),.dout(w_dff_B_XxuADOnt9_2),.clk(gclk));
	jdff dff_B_suFlq2yO6_2(.din(w_dff_B_XxuADOnt9_2),.dout(w_dff_B_suFlq2yO6_2),.clk(gclk));
	jdff dff_B_9XRI0iW76_2(.din(w_dff_B_suFlq2yO6_2),.dout(w_dff_B_9XRI0iW76_2),.clk(gclk));
	jdff dff_B_DYWbz1V77_2(.din(w_dff_B_9XRI0iW76_2),.dout(w_dff_B_DYWbz1V77_2),.clk(gclk));
	jdff dff_B_t2OAjFSP9_2(.din(w_dff_B_DYWbz1V77_2),.dout(w_dff_B_t2OAjFSP9_2),.clk(gclk));
	jdff dff_B_rQhOI8dt1_2(.din(w_dff_B_t2OAjFSP9_2),.dout(w_dff_B_rQhOI8dt1_2),.clk(gclk));
	jdff dff_B_aXoHWW1L3_2(.din(w_dff_B_rQhOI8dt1_2),.dout(w_dff_B_aXoHWW1L3_2),.clk(gclk));
	jdff dff_B_bb8YBTnX9_2(.din(w_dff_B_aXoHWW1L3_2),.dout(w_dff_B_bb8YBTnX9_2),.clk(gclk));
	jdff dff_B_V0we07Ct8_2(.din(w_dff_B_bb8YBTnX9_2),.dout(w_dff_B_V0we07Ct8_2),.clk(gclk));
	jdff dff_B_4J5hfqI36_2(.din(w_dff_B_V0we07Ct8_2),.dout(w_dff_B_4J5hfqI36_2),.clk(gclk));
	jdff dff_B_gjALG9Sg6_2(.din(w_dff_B_4J5hfqI36_2),.dout(w_dff_B_gjALG9Sg6_2),.clk(gclk));
	jdff dff_B_vcd18Xy44_2(.din(w_dff_B_gjALG9Sg6_2),.dout(w_dff_B_vcd18Xy44_2),.clk(gclk));
	jdff dff_B_MaBGK2ZJ6_2(.din(w_dff_B_vcd18Xy44_2),.dout(w_dff_B_MaBGK2ZJ6_2),.clk(gclk));
	jdff dff_B_rdBsrFSB6_2(.din(w_dff_B_MaBGK2ZJ6_2),.dout(w_dff_B_rdBsrFSB6_2),.clk(gclk));
	jdff dff_B_fOTeTZGn3_2(.din(w_dff_B_rdBsrFSB6_2),.dout(w_dff_B_fOTeTZGn3_2),.clk(gclk));
	jdff dff_B_CglMBADb8_2(.din(w_dff_B_fOTeTZGn3_2),.dout(w_dff_B_CglMBADb8_2),.clk(gclk));
	jdff dff_B_tJOgbhkn2_2(.din(w_dff_B_CglMBADb8_2),.dout(w_dff_B_tJOgbhkn2_2),.clk(gclk));
	jdff dff_B_tUghYg4N8_2(.din(w_dff_B_tJOgbhkn2_2),.dout(w_dff_B_tUghYg4N8_2),.clk(gclk));
	jdff dff_B_s9pv34mm5_0(.din(n1562),.dout(w_dff_B_s9pv34mm5_0),.clk(gclk));
	jdff dff_A_F5DGNIku5_1(.dout(w_n1550_0[1]),.din(w_dff_A_F5DGNIku5_1),.clk(gclk));
	jdff dff_B_e2bwT7h06_1(.din(n1498),.dout(w_dff_B_e2bwT7h06_1),.clk(gclk));
	jdff dff_B_CRk1sifL2_2(.din(n1426),.dout(w_dff_B_CRk1sifL2_2),.clk(gclk));
	jdff dff_B_Ju8zlzNq1_2(.din(w_dff_B_CRk1sifL2_2),.dout(w_dff_B_Ju8zlzNq1_2),.clk(gclk));
	jdff dff_B_BY1FXfIO0_2(.din(w_dff_B_Ju8zlzNq1_2),.dout(w_dff_B_BY1FXfIO0_2),.clk(gclk));
	jdff dff_B_WfLnq02U3_2(.din(w_dff_B_BY1FXfIO0_2),.dout(w_dff_B_WfLnq02U3_2),.clk(gclk));
	jdff dff_B_ksq5eyME8_2(.din(w_dff_B_WfLnq02U3_2),.dout(w_dff_B_ksq5eyME8_2),.clk(gclk));
	jdff dff_B_l6MKBJQM9_2(.din(w_dff_B_ksq5eyME8_2),.dout(w_dff_B_l6MKBJQM9_2),.clk(gclk));
	jdff dff_B_930jjDuG8_2(.din(w_dff_B_l6MKBJQM9_2),.dout(w_dff_B_930jjDuG8_2),.clk(gclk));
	jdff dff_B_EsZfHCgp1_2(.din(w_dff_B_930jjDuG8_2),.dout(w_dff_B_EsZfHCgp1_2),.clk(gclk));
	jdff dff_B_JnaD8V9o0_2(.din(w_dff_B_EsZfHCgp1_2),.dout(w_dff_B_JnaD8V9o0_2),.clk(gclk));
	jdff dff_B_BjsTLkAz3_2(.din(w_dff_B_JnaD8V9o0_2),.dout(w_dff_B_BjsTLkAz3_2),.clk(gclk));
	jdff dff_B_RL6P5p603_2(.din(w_dff_B_BjsTLkAz3_2),.dout(w_dff_B_RL6P5p603_2),.clk(gclk));
	jdff dff_B_hIKrwDcf8_2(.din(w_dff_B_RL6P5p603_2),.dout(w_dff_B_hIKrwDcf8_2),.clk(gclk));
	jdff dff_B_ogz0763N5_2(.din(w_dff_B_hIKrwDcf8_2),.dout(w_dff_B_ogz0763N5_2),.clk(gclk));
	jdff dff_B_PfZnDpBT2_2(.din(w_dff_B_ogz0763N5_2),.dout(w_dff_B_PfZnDpBT2_2),.clk(gclk));
	jdff dff_B_tnuc2eg79_2(.din(w_dff_B_PfZnDpBT2_2),.dout(w_dff_B_tnuc2eg79_2),.clk(gclk));
	jdff dff_B_7k1bm7ej2_2(.din(w_dff_B_tnuc2eg79_2),.dout(w_dff_B_7k1bm7ej2_2),.clk(gclk));
	jdff dff_B_zvaQSFfi3_2(.din(w_dff_B_7k1bm7ej2_2),.dout(w_dff_B_zvaQSFfi3_2),.clk(gclk));
	jdff dff_B_cLNwiovw4_2(.din(w_dff_B_zvaQSFfi3_2),.dout(w_dff_B_cLNwiovw4_2),.clk(gclk));
	jdff dff_B_8wOJKZMX3_2(.din(w_dff_B_cLNwiovw4_2),.dout(w_dff_B_8wOJKZMX3_2),.clk(gclk));
	jdff dff_B_SLA6GgvG4_2(.din(w_dff_B_8wOJKZMX3_2),.dout(w_dff_B_SLA6GgvG4_2),.clk(gclk));
	jdff dff_B_amgcxnxY8_2(.din(w_dff_B_SLA6GgvG4_2),.dout(w_dff_B_amgcxnxY8_2),.clk(gclk));
	jdff dff_B_v4Dq6eWx9_2(.din(w_dff_B_amgcxnxY8_2),.dout(w_dff_B_v4Dq6eWx9_2),.clk(gclk));
	jdff dff_B_yNxQI4gv3_2(.din(w_dff_B_v4Dq6eWx9_2),.dout(w_dff_B_yNxQI4gv3_2),.clk(gclk));
	jdff dff_B_FGIvQC5V9_2(.din(w_dff_B_yNxQI4gv3_2),.dout(w_dff_B_FGIvQC5V9_2),.clk(gclk));
	jdff dff_B_FndKnCOF7_2(.din(w_dff_B_FGIvQC5V9_2),.dout(w_dff_B_FndKnCOF7_2),.clk(gclk));
	jdff dff_B_wIsyC8f90_2(.din(w_dff_B_FndKnCOF7_2),.dout(w_dff_B_wIsyC8f90_2),.clk(gclk));
	jdff dff_B_OuhIXG5k1_2(.din(w_dff_B_wIsyC8f90_2),.dout(w_dff_B_OuhIXG5k1_2),.clk(gclk));
	jdff dff_B_fM5tUCeI0_2(.din(w_dff_B_OuhIXG5k1_2),.dout(w_dff_B_fM5tUCeI0_2),.clk(gclk));
	jdff dff_B_cwCqhBH69_2(.din(w_dff_B_fM5tUCeI0_2),.dout(w_dff_B_cwCqhBH69_2),.clk(gclk));
	jdff dff_B_Pw1ZbvxO1_2(.din(w_dff_B_cwCqhBH69_2),.dout(w_dff_B_Pw1ZbvxO1_2),.clk(gclk));
	jdff dff_B_JyhtQZQO0_2(.din(w_dff_B_Pw1ZbvxO1_2),.dout(w_dff_B_JyhtQZQO0_2),.clk(gclk));
	jdff dff_B_5Dh4twdb5_2(.din(w_dff_B_JyhtQZQO0_2),.dout(w_dff_B_5Dh4twdb5_2),.clk(gclk));
	jdff dff_B_UfOpPLRJ1_2(.din(w_dff_B_5Dh4twdb5_2),.dout(w_dff_B_UfOpPLRJ1_2),.clk(gclk));
	jdff dff_B_g28XbUXD3_2(.din(w_dff_B_UfOpPLRJ1_2),.dout(w_dff_B_g28XbUXD3_2),.clk(gclk));
	jdff dff_B_zYdXWDBQ3_2(.din(w_dff_B_g28XbUXD3_2),.dout(w_dff_B_zYdXWDBQ3_2),.clk(gclk));
	jdff dff_B_uSFFYiaJ4_2(.din(w_dff_B_zYdXWDBQ3_2),.dout(w_dff_B_uSFFYiaJ4_2),.clk(gclk));
	jdff dff_B_j8gS4rYn5_2(.din(w_dff_B_uSFFYiaJ4_2),.dout(w_dff_B_j8gS4rYn5_2),.clk(gclk));
	jdff dff_B_cpus0BYS8_2(.din(w_dff_B_j8gS4rYn5_2),.dout(w_dff_B_cpus0BYS8_2),.clk(gclk));
	jdff dff_B_DnWkXHHD1_2(.din(w_dff_B_cpus0BYS8_2),.dout(w_dff_B_DnWkXHHD1_2),.clk(gclk));
	jdff dff_B_0UOEMpfM8_2(.din(w_dff_B_DnWkXHHD1_2),.dout(w_dff_B_0UOEMpfM8_2),.clk(gclk));
	jdff dff_B_HVbczsyo8_2(.din(w_dff_B_0UOEMpfM8_2),.dout(w_dff_B_HVbczsyo8_2),.clk(gclk));
	jdff dff_B_EZtOMoZi1_2(.din(w_dff_B_HVbczsyo8_2),.dout(w_dff_B_EZtOMoZi1_2),.clk(gclk));
	jdff dff_B_tAhCEUVg1_2(.din(n1479),.dout(w_dff_B_tAhCEUVg1_2),.clk(gclk));
	jdff dff_B_ZSPAhZlk1_1(.din(n1427),.dout(w_dff_B_ZSPAhZlk1_1),.clk(gclk));
	jdff dff_B_BBihBqEI5_2(.din(n1348),.dout(w_dff_B_BBihBqEI5_2),.clk(gclk));
	jdff dff_B_jDDh1dZe2_2(.din(w_dff_B_BBihBqEI5_2),.dout(w_dff_B_jDDh1dZe2_2),.clk(gclk));
	jdff dff_B_GgoR3HXw2_2(.din(w_dff_B_jDDh1dZe2_2),.dout(w_dff_B_GgoR3HXw2_2),.clk(gclk));
	jdff dff_B_HiHWYSxc4_2(.din(w_dff_B_GgoR3HXw2_2),.dout(w_dff_B_HiHWYSxc4_2),.clk(gclk));
	jdff dff_B_v3TXDpmH7_2(.din(w_dff_B_HiHWYSxc4_2),.dout(w_dff_B_v3TXDpmH7_2),.clk(gclk));
	jdff dff_B_9oJoUrMx1_2(.din(w_dff_B_v3TXDpmH7_2),.dout(w_dff_B_9oJoUrMx1_2),.clk(gclk));
	jdff dff_B_ISiofFKw6_2(.din(w_dff_B_9oJoUrMx1_2),.dout(w_dff_B_ISiofFKw6_2),.clk(gclk));
	jdff dff_B_xRZfEihv5_2(.din(w_dff_B_ISiofFKw6_2),.dout(w_dff_B_xRZfEihv5_2),.clk(gclk));
	jdff dff_B_hIyYMjOF2_2(.din(w_dff_B_xRZfEihv5_2),.dout(w_dff_B_hIyYMjOF2_2),.clk(gclk));
	jdff dff_B_X6nD6tSp8_2(.din(w_dff_B_hIyYMjOF2_2),.dout(w_dff_B_X6nD6tSp8_2),.clk(gclk));
	jdff dff_B_WKhHgbCe4_2(.din(w_dff_B_X6nD6tSp8_2),.dout(w_dff_B_WKhHgbCe4_2),.clk(gclk));
	jdff dff_B_kQ7EQnuO3_2(.din(w_dff_B_WKhHgbCe4_2),.dout(w_dff_B_kQ7EQnuO3_2),.clk(gclk));
	jdff dff_B_5zgnJw3n2_2(.din(w_dff_B_kQ7EQnuO3_2),.dout(w_dff_B_5zgnJw3n2_2),.clk(gclk));
	jdff dff_B_wHnUWgf08_2(.din(w_dff_B_5zgnJw3n2_2),.dout(w_dff_B_wHnUWgf08_2),.clk(gclk));
	jdff dff_B_VekJkxUo3_2(.din(w_dff_B_wHnUWgf08_2),.dout(w_dff_B_VekJkxUo3_2),.clk(gclk));
	jdff dff_B_DBhouzLf2_2(.din(w_dff_B_VekJkxUo3_2),.dout(w_dff_B_DBhouzLf2_2),.clk(gclk));
	jdff dff_B_Zfm53BT94_2(.din(w_dff_B_DBhouzLf2_2),.dout(w_dff_B_Zfm53BT94_2),.clk(gclk));
	jdff dff_B_IBqI79TY6_2(.din(w_dff_B_Zfm53BT94_2),.dout(w_dff_B_IBqI79TY6_2),.clk(gclk));
	jdff dff_B_68jk4Xgo4_2(.din(w_dff_B_IBqI79TY6_2),.dout(w_dff_B_68jk4Xgo4_2),.clk(gclk));
	jdff dff_B_sTWsASjY0_2(.din(w_dff_B_68jk4Xgo4_2),.dout(w_dff_B_sTWsASjY0_2),.clk(gclk));
	jdff dff_B_aGyb8gCw7_2(.din(w_dff_B_sTWsASjY0_2),.dout(w_dff_B_aGyb8gCw7_2),.clk(gclk));
	jdff dff_B_QVHn0I109_2(.din(w_dff_B_aGyb8gCw7_2),.dout(w_dff_B_QVHn0I109_2),.clk(gclk));
	jdff dff_B_79NxnVDp1_2(.din(w_dff_B_QVHn0I109_2),.dout(w_dff_B_79NxnVDp1_2),.clk(gclk));
	jdff dff_B_s7opvF8h8_2(.din(w_dff_B_79NxnVDp1_2),.dout(w_dff_B_s7opvF8h8_2),.clk(gclk));
	jdff dff_B_t78o9VrW6_2(.din(w_dff_B_s7opvF8h8_2),.dout(w_dff_B_t78o9VrW6_2),.clk(gclk));
	jdff dff_B_YrlfMDkA7_2(.din(w_dff_B_t78o9VrW6_2),.dout(w_dff_B_YrlfMDkA7_2),.clk(gclk));
	jdff dff_B_3PDqQoUz8_2(.din(w_dff_B_YrlfMDkA7_2),.dout(w_dff_B_3PDqQoUz8_2),.clk(gclk));
	jdff dff_B_6rpQnCHN7_2(.din(w_dff_B_3PDqQoUz8_2),.dout(w_dff_B_6rpQnCHN7_2),.clk(gclk));
	jdff dff_B_2JdcIaBd0_2(.din(w_dff_B_6rpQnCHN7_2),.dout(w_dff_B_2JdcIaBd0_2),.clk(gclk));
	jdff dff_B_eKtQYpni8_2(.din(w_dff_B_2JdcIaBd0_2),.dout(w_dff_B_eKtQYpni8_2),.clk(gclk));
	jdff dff_B_cIpnUKxG6_2(.din(w_dff_B_eKtQYpni8_2),.dout(w_dff_B_cIpnUKxG6_2),.clk(gclk));
	jdff dff_B_2EQaBGhu3_2(.din(w_dff_B_cIpnUKxG6_2),.dout(w_dff_B_2EQaBGhu3_2),.clk(gclk));
	jdff dff_B_TG6jqPYo9_2(.din(w_dff_B_2EQaBGhu3_2),.dout(w_dff_B_TG6jqPYo9_2),.clk(gclk));
	jdff dff_B_JIKEOoQC7_2(.din(w_dff_B_TG6jqPYo9_2),.dout(w_dff_B_JIKEOoQC7_2),.clk(gclk));
	jdff dff_B_dGFEP0HU9_2(.din(w_dff_B_JIKEOoQC7_2),.dout(w_dff_B_dGFEP0HU9_2),.clk(gclk));
	jdff dff_B_moFxXqUc3_2(.din(w_dff_B_dGFEP0HU9_2),.dout(w_dff_B_moFxXqUc3_2),.clk(gclk));
	jdff dff_B_zrGK7h9Q9_2(.din(w_dff_B_moFxXqUc3_2),.dout(w_dff_B_zrGK7h9Q9_2),.clk(gclk));
	jdff dff_B_yajQF2IL8_2(.din(w_dff_B_zrGK7h9Q9_2),.dout(w_dff_B_yajQF2IL8_2),.clk(gclk));
	jdff dff_B_1mUiIhGD0_2(.din(w_dff_B_yajQF2IL8_2),.dout(w_dff_B_1mUiIhGD0_2),.clk(gclk));
	jdff dff_B_h43tcy7G1_2(.din(n1401),.dout(w_dff_B_h43tcy7G1_2),.clk(gclk));
	jdff dff_B_wy76JoGg3_1(.din(n1349),.dout(w_dff_B_wy76JoGg3_1),.clk(gclk));
	jdff dff_B_NeX1hRvQ1_2(.din(n1263),.dout(w_dff_B_NeX1hRvQ1_2),.clk(gclk));
	jdff dff_B_RWBEAAdS1_2(.din(w_dff_B_NeX1hRvQ1_2),.dout(w_dff_B_RWBEAAdS1_2),.clk(gclk));
	jdff dff_B_RVTA9aVm7_2(.din(w_dff_B_RWBEAAdS1_2),.dout(w_dff_B_RVTA9aVm7_2),.clk(gclk));
	jdff dff_B_zf0beyWt6_2(.din(w_dff_B_RVTA9aVm7_2),.dout(w_dff_B_zf0beyWt6_2),.clk(gclk));
	jdff dff_B_ACwv2XYC1_2(.din(w_dff_B_zf0beyWt6_2),.dout(w_dff_B_ACwv2XYC1_2),.clk(gclk));
	jdff dff_B_ueVYOmkw0_2(.din(w_dff_B_ACwv2XYC1_2),.dout(w_dff_B_ueVYOmkw0_2),.clk(gclk));
	jdff dff_B_LgATYXHV8_2(.din(w_dff_B_ueVYOmkw0_2),.dout(w_dff_B_LgATYXHV8_2),.clk(gclk));
	jdff dff_B_uwK8qIgI7_2(.din(w_dff_B_LgATYXHV8_2),.dout(w_dff_B_uwK8qIgI7_2),.clk(gclk));
	jdff dff_B_u0jfZRod8_2(.din(w_dff_B_uwK8qIgI7_2),.dout(w_dff_B_u0jfZRod8_2),.clk(gclk));
	jdff dff_B_EHBcFeNq6_2(.din(w_dff_B_u0jfZRod8_2),.dout(w_dff_B_EHBcFeNq6_2),.clk(gclk));
	jdff dff_B_OJxLDOx33_2(.din(w_dff_B_EHBcFeNq6_2),.dout(w_dff_B_OJxLDOx33_2),.clk(gclk));
	jdff dff_B_rewFnKMG4_2(.din(w_dff_B_OJxLDOx33_2),.dout(w_dff_B_rewFnKMG4_2),.clk(gclk));
	jdff dff_B_4lNU28JW5_2(.din(w_dff_B_rewFnKMG4_2),.dout(w_dff_B_4lNU28JW5_2),.clk(gclk));
	jdff dff_B_8mQQWD5G9_2(.din(w_dff_B_4lNU28JW5_2),.dout(w_dff_B_8mQQWD5G9_2),.clk(gclk));
	jdff dff_B_ShnYhHWD6_2(.din(w_dff_B_8mQQWD5G9_2),.dout(w_dff_B_ShnYhHWD6_2),.clk(gclk));
	jdff dff_B_xlD0g9lO1_2(.din(w_dff_B_ShnYhHWD6_2),.dout(w_dff_B_xlD0g9lO1_2),.clk(gclk));
	jdff dff_B_fF2yctoZ7_2(.din(w_dff_B_xlD0g9lO1_2),.dout(w_dff_B_fF2yctoZ7_2),.clk(gclk));
	jdff dff_B_Y1wkKzun8_2(.din(w_dff_B_fF2yctoZ7_2),.dout(w_dff_B_Y1wkKzun8_2),.clk(gclk));
	jdff dff_B_dNSLuPXO6_2(.din(w_dff_B_Y1wkKzun8_2),.dout(w_dff_B_dNSLuPXO6_2),.clk(gclk));
	jdff dff_B_G8qqZ5KO9_2(.din(w_dff_B_dNSLuPXO6_2),.dout(w_dff_B_G8qqZ5KO9_2),.clk(gclk));
	jdff dff_B_OERPKPWq2_2(.din(w_dff_B_G8qqZ5KO9_2),.dout(w_dff_B_OERPKPWq2_2),.clk(gclk));
	jdff dff_B_Dueiev5m7_2(.din(w_dff_B_OERPKPWq2_2),.dout(w_dff_B_Dueiev5m7_2),.clk(gclk));
	jdff dff_B_G9m2nPnM6_2(.din(w_dff_B_Dueiev5m7_2),.dout(w_dff_B_G9m2nPnM6_2),.clk(gclk));
	jdff dff_B_P8kuslus2_2(.din(w_dff_B_G9m2nPnM6_2),.dout(w_dff_B_P8kuslus2_2),.clk(gclk));
	jdff dff_B_Lj7OmQTa2_2(.din(w_dff_B_P8kuslus2_2),.dout(w_dff_B_Lj7OmQTa2_2),.clk(gclk));
	jdff dff_B_DZv6EsN07_2(.din(w_dff_B_Lj7OmQTa2_2),.dout(w_dff_B_DZv6EsN07_2),.clk(gclk));
	jdff dff_B_08JtWV9c9_2(.din(w_dff_B_DZv6EsN07_2),.dout(w_dff_B_08JtWV9c9_2),.clk(gclk));
	jdff dff_B_4FmvezaM7_2(.din(w_dff_B_08JtWV9c9_2),.dout(w_dff_B_4FmvezaM7_2),.clk(gclk));
	jdff dff_B_ttAipD6f0_2(.din(w_dff_B_4FmvezaM7_2),.dout(w_dff_B_ttAipD6f0_2),.clk(gclk));
	jdff dff_B_c6VXBlo29_2(.din(w_dff_B_ttAipD6f0_2),.dout(w_dff_B_c6VXBlo29_2),.clk(gclk));
	jdff dff_B_sSyisVPl4_2(.din(w_dff_B_c6VXBlo29_2),.dout(w_dff_B_sSyisVPl4_2),.clk(gclk));
	jdff dff_B_XZx3L21p3_2(.din(w_dff_B_sSyisVPl4_2),.dout(w_dff_B_XZx3L21p3_2),.clk(gclk));
	jdff dff_B_BirgbWRu8_2(.din(w_dff_B_XZx3L21p3_2),.dout(w_dff_B_BirgbWRu8_2),.clk(gclk));
	jdff dff_B_HGNURKlE3_2(.din(w_dff_B_BirgbWRu8_2),.dout(w_dff_B_HGNURKlE3_2),.clk(gclk));
	jdff dff_B_7HTfMSpd3_2(.din(w_dff_B_HGNURKlE3_2),.dout(w_dff_B_7HTfMSpd3_2),.clk(gclk));
	jdff dff_B_xJ4lo3gy1_2(.din(w_dff_B_7HTfMSpd3_2),.dout(w_dff_B_xJ4lo3gy1_2),.clk(gclk));
	jdff dff_B_j4ccORpw4_2(.din(n1316),.dout(w_dff_B_j4ccORpw4_2),.clk(gclk));
	jdff dff_B_pso4BWIG7_1(.din(n1264),.dout(w_dff_B_pso4BWIG7_1),.clk(gclk));
	jdff dff_B_1358zHiR8_2(.din(n1173),.dout(w_dff_B_1358zHiR8_2),.clk(gclk));
	jdff dff_B_CYXUL9BU8_2(.din(w_dff_B_1358zHiR8_2),.dout(w_dff_B_CYXUL9BU8_2),.clk(gclk));
	jdff dff_B_ZSNxD25b5_2(.din(w_dff_B_CYXUL9BU8_2),.dout(w_dff_B_ZSNxD25b5_2),.clk(gclk));
	jdff dff_B_AYe82MC54_2(.din(w_dff_B_ZSNxD25b5_2),.dout(w_dff_B_AYe82MC54_2),.clk(gclk));
	jdff dff_B_UQRwkBIb4_2(.din(w_dff_B_AYe82MC54_2),.dout(w_dff_B_UQRwkBIb4_2),.clk(gclk));
	jdff dff_B_AdAe421E2_2(.din(w_dff_B_UQRwkBIb4_2),.dout(w_dff_B_AdAe421E2_2),.clk(gclk));
	jdff dff_B_6asGMBeO7_2(.din(w_dff_B_AdAe421E2_2),.dout(w_dff_B_6asGMBeO7_2),.clk(gclk));
	jdff dff_B_nKGYjs7M3_2(.din(w_dff_B_6asGMBeO7_2),.dout(w_dff_B_nKGYjs7M3_2),.clk(gclk));
	jdff dff_B_uPiQvcUB2_2(.din(w_dff_B_nKGYjs7M3_2),.dout(w_dff_B_uPiQvcUB2_2),.clk(gclk));
	jdff dff_B_MWdC6FJw8_2(.din(w_dff_B_uPiQvcUB2_2),.dout(w_dff_B_MWdC6FJw8_2),.clk(gclk));
	jdff dff_B_4OLM8gYH6_2(.din(w_dff_B_MWdC6FJw8_2),.dout(w_dff_B_4OLM8gYH6_2),.clk(gclk));
	jdff dff_B_YGzHT0Ke1_2(.din(w_dff_B_4OLM8gYH6_2),.dout(w_dff_B_YGzHT0Ke1_2),.clk(gclk));
	jdff dff_B_vcWwLAXK1_2(.din(w_dff_B_YGzHT0Ke1_2),.dout(w_dff_B_vcWwLAXK1_2),.clk(gclk));
	jdff dff_B_fzaBfLtr1_2(.din(w_dff_B_vcWwLAXK1_2),.dout(w_dff_B_fzaBfLtr1_2),.clk(gclk));
	jdff dff_B_MfQrkHRc2_2(.din(w_dff_B_fzaBfLtr1_2),.dout(w_dff_B_MfQrkHRc2_2),.clk(gclk));
	jdff dff_B_silPUtMO9_2(.din(w_dff_B_MfQrkHRc2_2),.dout(w_dff_B_silPUtMO9_2),.clk(gclk));
	jdff dff_B_S0Z2uyZL2_2(.din(w_dff_B_silPUtMO9_2),.dout(w_dff_B_S0Z2uyZL2_2),.clk(gclk));
	jdff dff_B_8yEk5SvW4_2(.din(w_dff_B_S0Z2uyZL2_2),.dout(w_dff_B_8yEk5SvW4_2),.clk(gclk));
	jdff dff_B_pEDkgknt9_2(.din(w_dff_B_8yEk5SvW4_2),.dout(w_dff_B_pEDkgknt9_2),.clk(gclk));
	jdff dff_B_OTlGUdHG2_2(.din(w_dff_B_pEDkgknt9_2),.dout(w_dff_B_OTlGUdHG2_2),.clk(gclk));
	jdff dff_B_uofPgif12_2(.din(w_dff_B_OTlGUdHG2_2),.dout(w_dff_B_uofPgif12_2),.clk(gclk));
	jdff dff_B_ChPGCqtO6_2(.din(w_dff_B_uofPgif12_2),.dout(w_dff_B_ChPGCqtO6_2),.clk(gclk));
	jdff dff_B_zcb7UaWP0_2(.din(w_dff_B_ChPGCqtO6_2),.dout(w_dff_B_zcb7UaWP0_2),.clk(gclk));
	jdff dff_B_GYbfLOCB6_2(.din(w_dff_B_zcb7UaWP0_2),.dout(w_dff_B_GYbfLOCB6_2),.clk(gclk));
	jdff dff_B_mqJNDizi8_2(.din(w_dff_B_GYbfLOCB6_2),.dout(w_dff_B_mqJNDizi8_2),.clk(gclk));
	jdff dff_B_YGE03wAb8_2(.din(w_dff_B_mqJNDizi8_2),.dout(w_dff_B_YGE03wAb8_2),.clk(gclk));
	jdff dff_B_Q292y9IC7_2(.din(w_dff_B_YGE03wAb8_2),.dout(w_dff_B_Q292y9IC7_2),.clk(gclk));
	jdff dff_B_WCye4B1L3_2(.din(w_dff_B_Q292y9IC7_2),.dout(w_dff_B_WCye4B1L3_2),.clk(gclk));
	jdff dff_B_B58ROhoa7_2(.din(w_dff_B_WCye4B1L3_2),.dout(w_dff_B_B58ROhoa7_2),.clk(gclk));
	jdff dff_B_MAo13koB8_2(.din(w_dff_B_B58ROhoa7_2),.dout(w_dff_B_MAo13koB8_2),.clk(gclk));
	jdff dff_B_Vcwkr3mJ5_2(.din(w_dff_B_MAo13koB8_2),.dout(w_dff_B_Vcwkr3mJ5_2),.clk(gclk));
	jdff dff_B_jX9rnMVy8_2(.din(w_dff_B_Vcwkr3mJ5_2),.dout(w_dff_B_jX9rnMVy8_2),.clk(gclk));
	jdff dff_B_j1oyz5BA5_2(.din(w_dff_B_jX9rnMVy8_2),.dout(w_dff_B_j1oyz5BA5_2),.clk(gclk));
	jdff dff_B_9lJINcr55_2(.din(n1225),.dout(w_dff_B_9lJINcr55_2),.clk(gclk));
	jdff dff_B_G4BLumyx3_1(.din(n1174),.dout(w_dff_B_G4BLumyx3_1),.clk(gclk));
	jdff dff_B_Q3jPNhJv6_2(.din(n1069),.dout(w_dff_B_Q3jPNhJv6_2),.clk(gclk));
	jdff dff_B_wbRrDhLM7_2(.din(w_dff_B_Q3jPNhJv6_2),.dout(w_dff_B_wbRrDhLM7_2),.clk(gclk));
	jdff dff_B_ZUZcUyXr0_2(.din(w_dff_B_wbRrDhLM7_2),.dout(w_dff_B_ZUZcUyXr0_2),.clk(gclk));
	jdff dff_B_gIIwQgTX3_2(.din(w_dff_B_ZUZcUyXr0_2),.dout(w_dff_B_gIIwQgTX3_2),.clk(gclk));
	jdff dff_B_xuS6p7uN6_2(.din(w_dff_B_gIIwQgTX3_2),.dout(w_dff_B_xuS6p7uN6_2),.clk(gclk));
	jdff dff_B_0iImqIBf5_2(.din(w_dff_B_xuS6p7uN6_2),.dout(w_dff_B_0iImqIBf5_2),.clk(gclk));
	jdff dff_B_vbz6hfqB8_2(.din(w_dff_B_0iImqIBf5_2),.dout(w_dff_B_vbz6hfqB8_2),.clk(gclk));
	jdff dff_B_qnixko3u2_2(.din(w_dff_B_vbz6hfqB8_2),.dout(w_dff_B_qnixko3u2_2),.clk(gclk));
	jdff dff_B_FTMFh1rF0_2(.din(w_dff_B_qnixko3u2_2),.dout(w_dff_B_FTMFh1rF0_2),.clk(gclk));
	jdff dff_B_AU68H9Ma6_2(.din(w_dff_B_FTMFh1rF0_2),.dout(w_dff_B_AU68H9Ma6_2),.clk(gclk));
	jdff dff_B_PXvKcBjt5_2(.din(w_dff_B_AU68H9Ma6_2),.dout(w_dff_B_PXvKcBjt5_2),.clk(gclk));
	jdff dff_B_KAXABrBD4_2(.din(w_dff_B_PXvKcBjt5_2),.dout(w_dff_B_KAXABrBD4_2),.clk(gclk));
	jdff dff_B_gdYoejx88_2(.din(w_dff_B_KAXABrBD4_2),.dout(w_dff_B_gdYoejx88_2),.clk(gclk));
	jdff dff_B_sVMqajT57_2(.din(w_dff_B_gdYoejx88_2),.dout(w_dff_B_sVMqajT57_2),.clk(gclk));
	jdff dff_B_wsJfr5GO5_2(.din(w_dff_B_sVMqajT57_2),.dout(w_dff_B_wsJfr5GO5_2),.clk(gclk));
	jdff dff_B_9QDL4fAG9_2(.din(w_dff_B_wsJfr5GO5_2),.dout(w_dff_B_9QDL4fAG9_2),.clk(gclk));
	jdff dff_B_kl0hNwtY1_2(.din(w_dff_B_9QDL4fAG9_2),.dout(w_dff_B_kl0hNwtY1_2),.clk(gclk));
	jdff dff_B_Moe8oQkM1_2(.din(w_dff_B_kl0hNwtY1_2),.dout(w_dff_B_Moe8oQkM1_2),.clk(gclk));
	jdff dff_B_Z0tkFoNr0_2(.din(w_dff_B_Moe8oQkM1_2),.dout(w_dff_B_Z0tkFoNr0_2),.clk(gclk));
	jdff dff_B_VGf10PbV4_2(.din(w_dff_B_Z0tkFoNr0_2),.dout(w_dff_B_VGf10PbV4_2),.clk(gclk));
	jdff dff_B_rQQEUbGa5_2(.din(w_dff_B_VGf10PbV4_2),.dout(w_dff_B_rQQEUbGa5_2),.clk(gclk));
	jdff dff_B_i4zFlsOZ1_2(.din(w_dff_B_rQQEUbGa5_2),.dout(w_dff_B_i4zFlsOZ1_2),.clk(gclk));
	jdff dff_B_UnitFUWO0_2(.din(w_dff_B_i4zFlsOZ1_2),.dout(w_dff_B_UnitFUWO0_2),.clk(gclk));
	jdff dff_B_xkZ4nLUA8_2(.din(w_dff_B_UnitFUWO0_2),.dout(w_dff_B_xkZ4nLUA8_2),.clk(gclk));
	jdff dff_B_Lgee2QSR6_2(.din(w_dff_B_xkZ4nLUA8_2),.dout(w_dff_B_Lgee2QSR6_2),.clk(gclk));
	jdff dff_B_yO2qVK7s6_2(.din(w_dff_B_Lgee2QSR6_2),.dout(w_dff_B_yO2qVK7s6_2),.clk(gclk));
	jdff dff_B_2NTOnvvt3_2(.din(w_dff_B_yO2qVK7s6_2),.dout(w_dff_B_2NTOnvvt3_2),.clk(gclk));
	jdff dff_B_doNzjmTP1_2(.din(w_dff_B_2NTOnvvt3_2),.dout(w_dff_B_doNzjmTP1_2),.clk(gclk));
	jdff dff_B_Dgg0nkJt3_2(.din(w_dff_B_doNzjmTP1_2),.dout(w_dff_B_Dgg0nkJt3_2),.clk(gclk));
	jdff dff_B_GJjsYhnp3_2(.din(w_dff_B_Dgg0nkJt3_2),.dout(w_dff_B_GJjsYhnp3_2),.clk(gclk));
	jdff dff_B_kDDcdUhh8_2(.din(n1127),.dout(w_dff_B_kDDcdUhh8_2),.clk(gclk));
	jdff dff_B_Te2DMkeV2_1(.din(n1070),.dout(w_dff_B_Te2DMkeV2_1),.clk(gclk));
	jdff dff_B_Jsa86ADT8_2(.din(n971),.dout(w_dff_B_Jsa86ADT8_2),.clk(gclk));
	jdff dff_B_WL9chbz29_2(.din(w_dff_B_Jsa86ADT8_2),.dout(w_dff_B_WL9chbz29_2),.clk(gclk));
	jdff dff_B_ULj5iaHx7_2(.din(w_dff_B_WL9chbz29_2),.dout(w_dff_B_ULj5iaHx7_2),.clk(gclk));
	jdff dff_B_DHBfNhz54_2(.din(w_dff_B_ULj5iaHx7_2),.dout(w_dff_B_DHBfNhz54_2),.clk(gclk));
	jdff dff_B_2qGWFMQl2_2(.din(w_dff_B_DHBfNhz54_2),.dout(w_dff_B_2qGWFMQl2_2),.clk(gclk));
	jdff dff_B_aQGaA4Za0_2(.din(w_dff_B_2qGWFMQl2_2),.dout(w_dff_B_aQGaA4Za0_2),.clk(gclk));
	jdff dff_B_mjHKD8rN8_2(.din(w_dff_B_aQGaA4Za0_2),.dout(w_dff_B_mjHKD8rN8_2),.clk(gclk));
	jdff dff_B_oBXeoxYE2_2(.din(w_dff_B_mjHKD8rN8_2),.dout(w_dff_B_oBXeoxYE2_2),.clk(gclk));
	jdff dff_B_UlvHVh8l3_2(.din(w_dff_B_oBXeoxYE2_2),.dout(w_dff_B_UlvHVh8l3_2),.clk(gclk));
	jdff dff_B_yrL2DVxN3_2(.din(w_dff_B_UlvHVh8l3_2),.dout(w_dff_B_yrL2DVxN3_2),.clk(gclk));
	jdff dff_B_NkKw86oq4_2(.din(w_dff_B_yrL2DVxN3_2),.dout(w_dff_B_NkKw86oq4_2),.clk(gclk));
	jdff dff_B_14l0rrfd8_2(.din(w_dff_B_NkKw86oq4_2),.dout(w_dff_B_14l0rrfd8_2),.clk(gclk));
	jdff dff_B_kXV8kFB23_2(.din(w_dff_B_14l0rrfd8_2),.dout(w_dff_B_kXV8kFB23_2),.clk(gclk));
	jdff dff_B_kSCqlgoC6_2(.din(w_dff_B_kXV8kFB23_2),.dout(w_dff_B_kSCqlgoC6_2),.clk(gclk));
	jdff dff_B_3iU9ar9N8_2(.din(w_dff_B_kSCqlgoC6_2),.dout(w_dff_B_3iU9ar9N8_2),.clk(gclk));
	jdff dff_B_Gw5pAFzS1_2(.din(w_dff_B_3iU9ar9N8_2),.dout(w_dff_B_Gw5pAFzS1_2),.clk(gclk));
	jdff dff_B_rVHpWqyr2_2(.din(w_dff_B_Gw5pAFzS1_2),.dout(w_dff_B_rVHpWqyr2_2),.clk(gclk));
	jdff dff_B_qrzvK4L54_2(.din(w_dff_B_rVHpWqyr2_2),.dout(w_dff_B_qrzvK4L54_2),.clk(gclk));
	jdff dff_B_kM7teKYt7_2(.din(w_dff_B_qrzvK4L54_2),.dout(w_dff_B_kM7teKYt7_2),.clk(gclk));
	jdff dff_B_ES7MMwfb4_2(.din(w_dff_B_kM7teKYt7_2),.dout(w_dff_B_ES7MMwfb4_2),.clk(gclk));
	jdff dff_B_yhxDzAL87_2(.din(w_dff_B_ES7MMwfb4_2),.dout(w_dff_B_yhxDzAL87_2),.clk(gclk));
	jdff dff_B_6vJfkKJo8_2(.din(w_dff_B_yhxDzAL87_2),.dout(w_dff_B_6vJfkKJo8_2),.clk(gclk));
	jdff dff_B_coBziEtT1_2(.din(w_dff_B_6vJfkKJo8_2),.dout(w_dff_B_coBziEtT1_2),.clk(gclk));
	jdff dff_B_9Hzk6QpC5_2(.din(w_dff_B_coBziEtT1_2),.dout(w_dff_B_9Hzk6QpC5_2),.clk(gclk));
	jdff dff_B_owkWELKf1_2(.din(w_dff_B_9Hzk6QpC5_2),.dout(w_dff_B_owkWELKf1_2),.clk(gclk));
	jdff dff_B_WJPbcDJ61_2(.din(w_dff_B_owkWELKf1_2),.dout(w_dff_B_WJPbcDJ61_2),.clk(gclk));
	jdff dff_B_0GgBGg4k2_2(.din(w_dff_B_WJPbcDJ61_2),.dout(w_dff_B_0GgBGg4k2_2),.clk(gclk));
	jdff dff_B_zSTRPc7K1_2(.din(n1022),.dout(w_dff_B_zSTRPc7K1_2),.clk(gclk));
	jdff dff_B_EmgwCGB41_1(.din(n972),.dout(w_dff_B_EmgwCGB41_1),.clk(gclk));
	jdff dff_B_3nxafNs61_2(.din(n866),.dout(w_dff_B_3nxafNs61_2),.clk(gclk));
	jdff dff_B_UVOgzU6u1_2(.din(w_dff_B_3nxafNs61_2),.dout(w_dff_B_UVOgzU6u1_2),.clk(gclk));
	jdff dff_B_GUrKVJXz2_2(.din(w_dff_B_UVOgzU6u1_2),.dout(w_dff_B_GUrKVJXz2_2),.clk(gclk));
	jdff dff_B_NJZcMozq2_2(.din(w_dff_B_GUrKVJXz2_2),.dout(w_dff_B_NJZcMozq2_2),.clk(gclk));
	jdff dff_B_NDV9Pm8I8_2(.din(w_dff_B_NJZcMozq2_2),.dout(w_dff_B_NDV9Pm8I8_2),.clk(gclk));
	jdff dff_B_o2j6B1N85_2(.din(w_dff_B_NDV9Pm8I8_2),.dout(w_dff_B_o2j6B1N85_2),.clk(gclk));
	jdff dff_B_vH3utIIh2_2(.din(w_dff_B_o2j6B1N85_2),.dout(w_dff_B_vH3utIIh2_2),.clk(gclk));
	jdff dff_B_wCKZoReK9_2(.din(w_dff_B_vH3utIIh2_2),.dout(w_dff_B_wCKZoReK9_2),.clk(gclk));
	jdff dff_B_UCXrvMmd6_2(.din(w_dff_B_wCKZoReK9_2),.dout(w_dff_B_UCXrvMmd6_2),.clk(gclk));
	jdff dff_B_ohqaDXTR8_2(.din(w_dff_B_UCXrvMmd6_2),.dout(w_dff_B_ohqaDXTR8_2),.clk(gclk));
	jdff dff_B_LdsytaWj7_2(.din(w_dff_B_ohqaDXTR8_2),.dout(w_dff_B_LdsytaWj7_2),.clk(gclk));
	jdff dff_B_0fx8rzbe7_2(.din(w_dff_B_LdsytaWj7_2),.dout(w_dff_B_0fx8rzbe7_2),.clk(gclk));
	jdff dff_B_6b4szKvX3_2(.din(w_dff_B_0fx8rzbe7_2),.dout(w_dff_B_6b4szKvX3_2),.clk(gclk));
	jdff dff_B_rUdwhUp44_2(.din(w_dff_B_6b4szKvX3_2),.dout(w_dff_B_rUdwhUp44_2),.clk(gclk));
	jdff dff_B_W7VYc7rs4_2(.din(w_dff_B_rUdwhUp44_2),.dout(w_dff_B_W7VYc7rs4_2),.clk(gclk));
	jdff dff_B_HGTTSMio6_2(.din(w_dff_B_W7VYc7rs4_2),.dout(w_dff_B_HGTTSMio6_2),.clk(gclk));
	jdff dff_B_aeVR1pgf9_2(.din(w_dff_B_HGTTSMio6_2),.dout(w_dff_B_aeVR1pgf9_2),.clk(gclk));
	jdff dff_B_GcMdokl36_2(.din(w_dff_B_aeVR1pgf9_2),.dout(w_dff_B_GcMdokl36_2),.clk(gclk));
	jdff dff_B_4LTIuvhI7_2(.din(w_dff_B_GcMdokl36_2),.dout(w_dff_B_4LTIuvhI7_2),.clk(gclk));
	jdff dff_B_bk8ANp4Q0_2(.din(w_dff_B_4LTIuvhI7_2),.dout(w_dff_B_bk8ANp4Q0_2),.clk(gclk));
	jdff dff_B_VkVesc1V1_2(.din(w_dff_B_bk8ANp4Q0_2),.dout(w_dff_B_VkVesc1V1_2),.clk(gclk));
	jdff dff_B_CCcb015G0_2(.din(w_dff_B_VkVesc1V1_2),.dout(w_dff_B_CCcb015G0_2),.clk(gclk));
	jdff dff_B_gPYa9o3J8_2(.din(w_dff_B_CCcb015G0_2),.dout(w_dff_B_gPYa9o3J8_2),.clk(gclk));
	jdff dff_B_krEo57156_2(.din(w_dff_B_gPYa9o3J8_2),.dout(w_dff_B_krEo57156_2),.clk(gclk));
	jdff dff_B_KJRKARdL5_2(.din(n917),.dout(w_dff_B_KJRKARdL5_2),.clk(gclk));
	jdff dff_B_PslMiuzK5_1(.din(n867),.dout(w_dff_B_PslMiuzK5_1),.clk(gclk));
	jdff dff_B_3wzpqXid2_2(.din(n767),.dout(w_dff_B_3wzpqXid2_2),.clk(gclk));
	jdff dff_B_ozkBiLVY8_2(.din(w_dff_B_3wzpqXid2_2),.dout(w_dff_B_ozkBiLVY8_2),.clk(gclk));
	jdff dff_B_eA6gvZl36_2(.din(w_dff_B_ozkBiLVY8_2),.dout(w_dff_B_eA6gvZl36_2),.clk(gclk));
	jdff dff_B_hsfvYqfn4_2(.din(w_dff_B_eA6gvZl36_2),.dout(w_dff_B_hsfvYqfn4_2),.clk(gclk));
	jdff dff_B_7IV9eM1K8_2(.din(w_dff_B_hsfvYqfn4_2),.dout(w_dff_B_7IV9eM1K8_2),.clk(gclk));
	jdff dff_B_3IQy30G14_2(.din(w_dff_B_7IV9eM1K8_2),.dout(w_dff_B_3IQy30G14_2),.clk(gclk));
	jdff dff_B_QF05wyeV8_2(.din(w_dff_B_3IQy30G14_2),.dout(w_dff_B_QF05wyeV8_2),.clk(gclk));
	jdff dff_B_6gY4hOPR1_2(.din(w_dff_B_QF05wyeV8_2),.dout(w_dff_B_6gY4hOPR1_2),.clk(gclk));
	jdff dff_B_hYDsCOy90_2(.din(w_dff_B_6gY4hOPR1_2),.dout(w_dff_B_hYDsCOy90_2),.clk(gclk));
	jdff dff_B_Iq8m2WdW3_2(.din(w_dff_B_hYDsCOy90_2),.dout(w_dff_B_Iq8m2WdW3_2),.clk(gclk));
	jdff dff_B_Fo6RKRtK0_2(.din(w_dff_B_Iq8m2WdW3_2),.dout(w_dff_B_Fo6RKRtK0_2),.clk(gclk));
	jdff dff_B_PPbiLaxP4_2(.din(w_dff_B_Fo6RKRtK0_2),.dout(w_dff_B_PPbiLaxP4_2),.clk(gclk));
	jdff dff_B_qfUqshtS3_2(.din(w_dff_B_PPbiLaxP4_2),.dout(w_dff_B_qfUqshtS3_2),.clk(gclk));
	jdff dff_B_HAn7BQya3_2(.din(w_dff_B_qfUqshtS3_2),.dout(w_dff_B_HAn7BQya3_2),.clk(gclk));
	jdff dff_B_o6nKKGqA4_2(.din(w_dff_B_HAn7BQya3_2),.dout(w_dff_B_o6nKKGqA4_2),.clk(gclk));
	jdff dff_B_W3KqP1vG5_2(.din(w_dff_B_o6nKKGqA4_2),.dout(w_dff_B_W3KqP1vG5_2),.clk(gclk));
	jdff dff_B_7HT5c9Ez2_2(.din(w_dff_B_W3KqP1vG5_2),.dout(w_dff_B_7HT5c9Ez2_2),.clk(gclk));
	jdff dff_B_P5rom5oU2_2(.din(w_dff_B_7HT5c9Ez2_2),.dout(w_dff_B_P5rom5oU2_2),.clk(gclk));
	jdff dff_B_aIRjaaT32_2(.din(w_dff_B_P5rom5oU2_2),.dout(w_dff_B_aIRjaaT32_2),.clk(gclk));
	jdff dff_B_qhDAxbfJ7_2(.din(w_dff_B_aIRjaaT32_2),.dout(w_dff_B_qhDAxbfJ7_2),.clk(gclk));
	jdff dff_B_AjlORad90_2(.din(w_dff_B_qhDAxbfJ7_2),.dout(w_dff_B_AjlORad90_2),.clk(gclk));
	jdff dff_B_wXnEFDJP0_2(.din(n811),.dout(w_dff_B_wXnEFDJP0_2),.clk(gclk));
	jdff dff_B_akapbC7f5_1(.din(n768),.dout(w_dff_B_akapbC7f5_1),.clk(gclk));
	jdff dff_B_Cdhe2alZ3_2(.din(n674),.dout(w_dff_B_Cdhe2alZ3_2),.clk(gclk));
	jdff dff_B_Xc8s8caI0_2(.din(w_dff_B_Cdhe2alZ3_2),.dout(w_dff_B_Xc8s8caI0_2),.clk(gclk));
	jdff dff_B_3urXrUrZ3_2(.din(w_dff_B_Xc8s8caI0_2),.dout(w_dff_B_3urXrUrZ3_2),.clk(gclk));
	jdff dff_B_56jTcQuB8_2(.din(w_dff_B_3urXrUrZ3_2),.dout(w_dff_B_56jTcQuB8_2),.clk(gclk));
	jdff dff_B_YA83Q8Oi2_2(.din(w_dff_B_56jTcQuB8_2),.dout(w_dff_B_YA83Q8Oi2_2),.clk(gclk));
	jdff dff_B_Ddzte2yZ6_2(.din(w_dff_B_YA83Q8Oi2_2),.dout(w_dff_B_Ddzte2yZ6_2),.clk(gclk));
	jdff dff_B_kcdaRHzb4_2(.din(w_dff_B_Ddzte2yZ6_2),.dout(w_dff_B_kcdaRHzb4_2),.clk(gclk));
	jdff dff_B_LDt8Pycl5_2(.din(w_dff_B_kcdaRHzb4_2),.dout(w_dff_B_LDt8Pycl5_2),.clk(gclk));
	jdff dff_B_8RBtMjv79_2(.din(w_dff_B_LDt8Pycl5_2),.dout(w_dff_B_8RBtMjv79_2),.clk(gclk));
	jdff dff_B_pZRsApnk2_2(.din(w_dff_B_8RBtMjv79_2),.dout(w_dff_B_pZRsApnk2_2),.clk(gclk));
	jdff dff_B_2j6luKJ57_2(.din(w_dff_B_pZRsApnk2_2),.dout(w_dff_B_2j6luKJ57_2),.clk(gclk));
	jdff dff_B_nCotYWDx6_2(.din(w_dff_B_2j6luKJ57_2),.dout(w_dff_B_nCotYWDx6_2),.clk(gclk));
	jdff dff_B_HBBJkLbV5_2(.din(w_dff_B_nCotYWDx6_2),.dout(w_dff_B_HBBJkLbV5_2),.clk(gclk));
	jdff dff_B_Zk2TiZMg6_2(.din(w_dff_B_HBBJkLbV5_2),.dout(w_dff_B_Zk2TiZMg6_2),.clk(gclk));
	jdff dff_B_Scitgxlo9_2(.din(w_dff_B_Zk2TiZMg6_2),.dout(w_dff_B_Scitgxlo9_2),.clk(gclk));
	jdff dff_B_zVYTE8Q64_2(.din(w_dff_B_Scitgxlo9_2),.dout(w_dff_B_zVYTE8Q64_2),.clk(gclk));
	jdff dff_B_htiST99C0_2(.din(w_dff_B_zVYTE8Q64_2),.dout(w_dff_B_htiST99C0_2),.clk(gclk));
	jdff dff_B_CsMAmuPH7_2(.din(w_dff_B_htiST99C0_2),.dout(w_dff_B_CsMAmuPH7_2),.clk(gclk));
	jdff dff_B_TlpexhRO4_2(.din(n711),.dout(w_dff_B_TlpexhRO4_2),.clk(gclk));
	jdff dff_B_50KEP5WD7_1(.din(n675),.dout(w_dff_B_50KEP5WD7_1),.clk(gclk));
	jdff dff_B_Z1TeaOf85_2(.din(n588),.dout(w_dff_B_Z1TeaOf85_2),.clk(gclk));
	jdff dff_B_fccJNTth2_2(.din(w_dff_B_Z1TeaOf85_2),.dout(w_dff_B_fccJNTth2_2),.clk(gclk));
	jdff dff_B_muVYIs6Z0_2(.din(w_dff_B_fccJNTth2_2),.dout(w_dff_B_muVYIs6Z0_2),.clk(gclk));
	jdff dff_B_2QHyCNqZ1_2(.din(w_dff_B_muVYIs6Z0_2),.dout(w_dff_B_2QHyCNqZ1_2),.clk(gclk));
	jdff dff_B_eEE9d9w62_2(.din(w_dff_B_2QHyCNqZ1_2),.dout(w_dff_B_eEE9d9w62_2),.clk(gclk));
	jdff dff_B_piToqil80_2(.din(w_dff_B_eEE9d9w62_2),.dout(w_dff_B_piToqil80_2),.clk(gclk));
	jdff dff_B_oQCZKjdf1_2(.din(w_dff_B_piToqil80_2),.dout(w_dff_B_oQCZKjdf1_2),.clk(gclk));
	jdff dff_B_xLwPjdD22_2(.din(w_dff_B_oQCZKjdf1_2),.dout(w_dff_B_xLwPjdD22_2),.clk(gclk));
	jdff dff_B_1LUUEQ075_2(.din(w_dff_B_xLwPjdD22_2),.dout(w_dff_B_1LUUEQ075_2),.clk(gclk));
	jdff dff_B_RAJxfbuE4_2(.din(w_dff_B_1LUUEQ075_2),.dout(w_dff_B_RAJxfbuE4_2),.clk(gclk));
	jdff dff_B_6uxPmr7A3_2(.din(w_dff_B_RAJxfbuE4_2),.dout(w_dff_B_6uxPmr7A3_2),.clk(gclk));
	jdff dff_B_92CiVAVv7_2(.din(w_dff_B_6uxPmr7A3_2),.dout(w_dff_B_92CiVAVv7_2),.clk(gclk));
	jdff dff_B_Zu1tM6Io1_2(.din(w_dff_B_92CiVAVv7_2),.dout(w_dff_B_Zu1tM6Io1_2),.clk(gclk));
	jdff dff_B_SucoWBa65_2(.din(w_dff_B_Zu1tM6Io1_2),.dout(w_dff_B_SucoWBa65_2),.clk(gclk));
	jdff dff_B_8pJGz1xv6_2(.din(w_dff_B_SucoWBa65_2),.dout(w_dff_B_8pJGz1xv6_2),.clk(gclk));
	jdff dff_B_hOcmHsaa3_2(.din(n618),.dout(w_dff_B_hOcmHsaa3_2),.clk(gclk));
	jdff dff_B_TXZvMaLp9_1(.din(n589),.dout(w_dff_B_TXZvMaLp9_1),.clk(gclk));
	jdff dff_B_hvmf0dpK5_2(.din(n509),.dout(w_dff_B_hvmf0dpK5_2),.clk(gclk));
	jdff dff_B_vc5hhF7P3_2(.din(w_dff_B_hvmf0dpK5_2),.dout(w_dff_B_vc5hhF7P3_2),.clk(gclk));
	jdff dff_B_vAboxJed7_2(.din(w_dff_B_vc5hhF7P3_2),.dout(w_dff_B_vAboxJed7_2),.clk(gclk));
	jdff dff_B_GDaAzkyS8_2(.din(w_dff_B_vAboxJed7_2),.dout(w_dff_B_GDaAzkyS8_2),.clk(gclk));
	jdff dff_B_gDNdf3p49_2(.din(w_dff_B_GDaAzkyS8_2),.dout(w_dff_B_gDNdf3p49_2),.clk(gclk));
	jdff dff_B_FxfT3svE7_2(.din(w_dff_B_gDNdf3p49_2),.dout(w_dff_B_FxfT3svE7_2),.clk(gclk));
	jdff dff_B_guMEdJmj5_2(.din(w_dff_B_FxfT3svE7_2),.dout(w_dff_B_guMEdJmj5_2),.clk(gclk));
	jdff dff_B_CtvSUjyT0_2(.din(w_dff_B_guMEdJmj5_2),.dout(w_dff_B_CtvSUjyT0_2),.clk(gclk));
	jdff dff_B_oO173jvh5_2(.din(w_dff_B_CtvSUjyT0_2),.dout(w_dff_B_oO173jvh5_2),.clk(gclk));
	jdff dff_B_gPYgbGhE7_2(.din(w_dff_B_oO173jvh5_2),.dout(w_dff_B_gPYgbGhE7_2),.clk(gclk));
	jdff dff_B_iZulZs0t8_2(.din(w_dff_B_gPYgbGhE7_2),.dout(w_dff_B_iZulZs0t8_2),.clk(gclk));
	jdff dff_B_FoTdDfnG1_2(.din(w_dff_B_iZulZs0t8_2),.dout(w_dff_B_FoTdDfnG1_2),.clk(gclk));
	jdff dff_B_HiolJOlV9_2(.din(n532),.dout(w_dff_B_HiolJOlV9_2),.clk(gclk));
	jdff dff_B_NrstpOeQ0_1(.din(n510),.dout(w_dff_B_NrstpOeQ0_1),.clk(gclk));
	jdff dff_B_GQeXlzud5_2(.din(n437),.dout(w_dff_B_GQeXlzud5_2),.clk(gclk));
	jdff dff_B_0beilgAt0_2(.din(w_dff_B_GQeXlzud5_2),.dout(w_dff_B_0beilgAt0_2),.clk(gclk));
	jdff dff_B_3ss2RhTb5_2(.din(w_dff_B_0beilgAt0_2),.dout(w_dff_B_3ss2RhTb5_2),.clk(gclk));
	jdff dff_B_Q3DYyzPh2_2(.din(w_dff_B_3ss2RhTb5_2),.dout(w_dff_B_Q3DYyzPh2_2),.clk(gclk));
	jdff dff_B_719WvJAH0_2(.din(w_dff_B_Q3DYyzPh2_2),.dout(w_dff_B_719WvJAH0_2),.clk(gclk));
	jdff dff_B_LQSDncny9_2(.din(w_dff_B_719WvJAH0_2),.dout(w_dff_B_LQSDncny9_2),.clk(gclk));
	jdff dff_B_7rBiztZi3_2(.din(w_dff_B_LQSDncny9_2),.dout(w_dff_B_7rBiztZi3_2),.clk(gclk));
	jdff dff_B_60wxpPpz4_2(.din(w_dff_B_7rBiztZi3_2),.dout(w_dff_B_60wxpPpz4_2),.clk(gclk));
	jdff dff_B_45LVaV9I9_2(.din(w_dff_B_60wxpPpz4_2),.dout(w_dff_B_45LVaV9I9_2),.clk(gclk));
	jdff dff_B_8C6irrye9_2(.din(n453),.dout(w_dff_B_8C6irrye9_2),.clk(gclk));
	jdff dff_B_lYkQHvFO0_2(.din(w_dff_B_8C6irrye9_2),.dout(w_dff_B_lYkQHvFO0_2),.clk(gclk));
	jdff dff_B_BsPgbHp52_1(.din(n438),.dout(w_dff_B_BsPgbHp52_1),.clk(gclk));
	jdff dff_B_ueJL4jap8_1(.din(w_dff_B_BsPgbHp52_1),.dout(w_dff_B_ueJL4jap8_1),.clk(gclk));
	jdff dff_B_QnoYSYpE9_1(.din(w_dff_B_ueJL4jap8_1),.dout(w_dff_B_QnoYSYpE9_1),.clk(gclk));
	jdff dff_B_O29eXEyM1_1(.din(w_dff_B_QnoYSYpE9_1),.dout(w_dff_B_O29eXEyM1_1),.clk(gclk));
	jdff dff_B_B5BTH9ym8_1(.din(w_dff_B_O29eXEyM1_1),.dout(w_dff_B_B5BTH9ym8_1),.clk(gclk));
	jdff dff_B_aSZoaJ0K5_1(.din(w_dff_B_B5BTH9ym8_1),.dout(w_dff_B_aSZoaJ0K5_1),.clk(gclk));
	jdff dff_B_rcbFvTAZ5_0(.din(n381),.dout(w_dff_B_rcbFvTAZ5_0),.clk(gclk));
	jdff dff_B_KMrHkR3x1_0(.din(w_dff_B_rcbFvTAZ5_0),.dout(w_dff_B_KMrHkR3x1_0),.clk(gclk));
	jdff dff_A_rRBiOC0i3_0(.dout(w_n380_0[0]),.din(w_dff_A_rRBiOC0i3_0),.clk(gclk));
	jdff dff_A_y1T94mrB0_0(.dout(w_dff_A_rRBiOC0i3_0),.din(w_dff_A_y1T94mrB0_0),.clk(gclk));
	jdff dff_A_wYtxhkNR9_0(.dout(w_dff_A_y1T94mrB0_0),.din(w_dff_A_wYtxhkNR9_0),.clk(gclk));
	jdff dff_B_wP9WFB291_1(.din(n374),.dout(w_dff_B_wP9WFB291_1),.clk(gclk));
	jdff dff_A_ahOAYgm48_0(.dout(w_n314_0[0]),.din(w_dff_A_ahOAYgm48_0),.clk(gclk));
	jdff dff_A_j98TKgFe4_1(.dout(w_n314_0[1]),.din(w_dff_A_j98TKgFe4_1),.clk(gclk));
	jdff dff_A_N92C5aQQ8_1(.dout(w_dff_A_j98TKgFe4_1),.din(w_dff_A_N92C5aQQ8_1),.clk(gclk));
	jdff dff_A_HgPoA1yu6_1(.dout(w_n372_0[1]),.din(w_dff_A_HgPoA1yu6_1),.clk(gclk));
	jdff dff_A_dolF8lSb0_1(.dout(w_dff_A_HgPoA1yu6_1),.din(w_dff_A_dolF8lSb0_1),.clk(gclk));
	jdff dff_A_0eUDpDWO3_1(.dout(w_dff_A_dolF8lSb0_1),.din(w_dff_A_0eUDpDWO3_1),.clk(gclk));
	jdff dff_A_YOjFMLg99_1(.dout(w_dff_A_0eUDpDWO3_1),.din(w_dff_A_YOjFMLg99_1),.clk(gclk));
	jdff dff_A_gnSkQPUF5_1(.dout(w_dff_A_YOjFMLg99_1),.din(w_dff_A_gnSkQPUF5_1),.clk(gclk));
	jdff dff_A_evwGOEkL4_1(.dout(w_dff_A_gnSkQPUF5_1),.din(w_dff_A_evwGOEkL4_1),.clk(gclk));
	jdff dff_B_6I2knGDc5_2(.din(n1627),.dout(w_dff_B_6I2knGDc5_2),.clk(gclk));
	jdff dff_B_DlNTa9EC7_2(.din(w_dff_B_6I2knGDc5_2),.dout(w_dff_B_DlNTa9EC7_2),.clk(gclk));
	jdff dff_B_EkZtMXUx2_1(.din(n1625),.dout(w_dff_B_EkZtMXUx2_1),.clk(gclk));
	jdff dff_B_ubP4Wdas1_2(.din(n1566),.dout(w_dff_B_ubP4Wdas1_2),.clk(gclk));
	jdff dff_B_dS7lo7wE7_2(.din(w_dff_B_ubP4Wdas1_2),.dout(w_dff_B_dS7lo7wE7_2),.clk(gclk));
	jdff dff_B_3lAGRwe02_2(.din(w_dff_B_dS7lo7wE7_2),.dout(w_dff_B_3lAGRwe02_2),.clk(gclk));
	jdff dff_B_DF2O6JJH6_2(.din(w_dff_B_3lAGRwe02_2),.dout(w_dff_B_DF2O6JJH6_2),.clk(gclk));
	jdff dff_B_z6aCkRW00_2(.din(w_dff_B_DF2O6JJH6_2),.dout(w_dff_B_z6aCkRW00_2),.clk(gclk));
	jdff dff_B_2etEtMpm6_2(.din(w_dff_B_z6aCkRW00_2),.dout(w_dff_B_2etEtMpm6_2),.clk(gclk));
	jdff dff_B_dM4QFiMw2_2(.din(w_dff_B_2etEtMpm6_2),.dout(w_dff_B_dM4QFiMw2_2),.clk(gclk));
	jdff dff_B_2yQ2y7g95_2(.din(w_dff_B_dM4QFiMw2_2),.dout(w_dff_B_2yQ2y7g95_2),.clk(gclk));
	jdff dff_B_wKWoGesb3_2(.din(w_dff_B_2yQ2y7g95_2),.dout(w_dff_B_wKWoGesb3_2),.clk(gclk));
	jdff dff_B_84NLMqOb9_2(.din(w_dff_B_wKWoGesb3_2),.dout(w_dff_B_84NLMqOb9_2),.clk(gclk));
	jdff dff_B_uf1EqLnv8_2(.din(w_dff_B_84NLMqOb9_2),.dout(w_dff_B_uf1EqLnv8_2),.clk(gclk));
	jdff dff_B_3QbwMOam5_2(.din(w_dff_B_uf1EqLnv8_2),.dout(w_dff_B_3QbwMOam5_2),.clk(gclk));
	jdff dff_B_SO8TDBDr4_2(.din(w_dff_B_3QbwMOam5_2),.dout(w_dff_B_SO8TDBDr4_2),.clk(gclk));
	jdff dff_B_4tgEq3PU0_2(.din(w_dff_B_SO8TDBDr4_2),.dout(w_dff_B_4tgEq3PU0_2),.clk(gclk));
	jdff dff_B_Spu0gkCn5_2(.din(w_dff_B_4tgEq3PU0_2),.dout(w_dff_B_Spu0gkCn5_2),.clk(gclk));
	jdff dff_B_NJAlfSUW4_2(.din(w_dff_B_Spu0gkCn5_2),.dout(w_dff_B_NJAlfSUW4_2),.clk(gclk));
	jdff dff_B_x5OsXYSJ8_2(.din(w_dff_B_NJAlfSUW4_2),.dout(w_dff_B_x5OsXYSJ8_2),.clk(gclk));
	jdff dff_B_KdhXDiYh3_2(.din(w_dff_B_x5OsXYSJ8_2),.dout(w_dff_B_KdhXDiYh3_2),.clk(gclk));
	jdff dff_B_CKwbgnXW0_2(.din(w_dff_B_KdhXDiYh3_2),.dout(w_dff_B_CKwbgnXW0_2),.clk(gclk));
	jdff dff_B_kcByU88V1_2(.din(w_dff_B_CKwbgnXW0_2),.dout(w_dff_B_kcByU88V1_2),.clk(gclk));
	jdff dff_B_heUYiaTb6_2(.din(w_dff_B_kcByU88V1_2),.dout(w_dff_B_heUYiaTb6_2),.clk(gclk));
	jdff dff_B_CWZPdP6U1_2(.din(w_dff_B_heUYiaTb6_2),.dout(w_dff_B_CWZPdP6U1_2),.clk(gclk));
	jdff dff_B_DUHs937k4_2(.din(w_dff_B_CWZPdP6U1_2),.dout(w_dff_B_DUHs937k4_2),.clk(gclk));
	jdff dff_B_IioNZuZc3_2(.din(w_dff_B_DUHs937k4_2),.dout(w_dff_B_IioNZuZc3_2),.clk(gclk));
	jdff dff_B_B9vIPMFR2_2(.din(w_dff_B_IioNZuZc3_2),.dout(w_dff_B_B9vIPMFR2_2),.clk(gclk));
	jdff dff_B_N80iKUl86_2(.din(w_dff_B_B9vIPMFR2_2),.dout(w_dff_B_N80iKUl86_2),.clk(gclk));
	jdff dff_B_ttFVcsjR6_2(.din(w_dff_B_N80iKUl86_2),.dout(w_dff_B_ttFVcsjR6_2),.clk(gclk));
	jdff dff_B_THKSeorq9_2(.din(w_dff_B_ttFVcsjR6_2),.dout(w_dff_B_THKSeorq9_2),.clk(gclk));
	jdff dff_B_w0GMMlyp1_2(.din(w_dff_B_THKSeorq9_2),.dout(w_dff_B_w0GMMlyp1_2),.clk(gclk));
	jdff dff_B_Yxrf35pC7_2(.din(w_dff_B_w0GMMlyp1_2),.dout(w_dff_B_Yxrf35pC7_2),.clk(gclk));
	jdff dff_B_4Il2zcGd3_2(.din(w_dff_B_Yxrf35pC7_2),.dout(w_dff_B_4Il2zcGd3_2),.clk(gclk));
	jdff dff_B_hS6HtJUS4_2(.din(w_dff_B_4Il2zcGd3_2),.dout(w_dff_B_hS6HtJUS4_2),.clk(gclk));
	jdff dff_B_OYsJtcii9_2(.din(w_dff_B_hS6HtJUS4_2),.dout(w_dff_B_OYsJtcii9_2),.clk(gclk));
	jdff dff_B_teUgY3HQ3_2(.din(w_dff_B_OYsJtcii9_2),.dout(w_dff_B_teUgY3HQ3_2),.clk(gclk));
	jdff dff_B_u5c6ACBd6_2(.din(w_dff_B_teUgY3HQ3_2),.dout(w_dff_B_u5c6ACBd6_2),.clk(gclk));
	jdff dff_B_3VTx7P0T4_2(.din(w_dff_B_u5c6ACBd6_2),.dout(w_dff_B_3VTx7P0T4_2),.clk(gclk));
	jdff dff_B_g0Tf01TQ6_2(.din(w_dff_B_3VTx7P0T4_2),.dout(w_dff_B_g0Tf01TQ6_2),.clk(gclk));
	jdff dff_B_WklhyrFh5_2(.din(w_dff_B_g0Tf01TQ6_2),.dout(w_dff_B_WklhyrFh5_2),.clk(gclk));
	jdff dff_B_31PN68Rk6_2(.din(w_dff_B_WklhyrFh5_2),.dout(w_dff_B_31PN68Rk6_2),.clk(gclk));
	jdff dff_B_TVlstJ6z2_2(.din(w_dff_B_31PN68Rk6_2),.dout(w_dff_B_TVlstJ6z2_2),.clk(gclk));
	jdff dff_B_AjfAb4Rw8_2(.din(w_dff_B_TVlstJ6z2_2),.dout(w_dff_B_AjfAb4Rw8_2),.clk(gclk));
	jdff dff_B_gBeuXSrg7_2(.din(w_dff_B_AjfAb4Rw8_2),.dout(w_dff_B_gBeuXSrg7_2),.clk(gclk));
	jdff dff_B_5W3R03Kh1_2(.din(w_dff_B_gBeuXSrg7_2),.dout(w_dff_B_5W3R03Kh1_2),.clk(gclk));
	jdff dff_B_1aagcxQJ3_2(.din(w_dff_B_5W3R03Kh1_2),.dout(w_dff_B_1aagcxQJ3_2),.clk(gclk));
	jdff dff_B_610dQHof7_2(.din(w_dff_B_1aagcxQJ3_2),.dout(w_dff_B_610dQHof7_2),.clk(gclk));
	jdff dff_B_ue8UUm0w1_2(.din(w_dff_B_610dQHof7_2),.dout(w_dff_B_ue8UUm0w1_2),.clk(gclk));
	jdff dff_B_EVsqjVM83_2(.din(w_dff_B_ue8UUm0w1_2),.dout(w_dff_B_EVsqjVM83_2),.clk(gclk));
	jdff dff_B_CdmtuydS5_1(.din(n1567),.dout(w_dff_B_CdmtuydS5_1),.clk(gclk));
	jdff dff_B_sxuDsbth0_2(.din(n1502),.dout(w_dff_B_sxuDsbth0_2),.clk(gclk));
	jdff dff_B_HzuHDBeP6_2(.din(w_dff_B_sxuDsbth0_2),.dout(w_dff_B_HzuHDBeP6_2),.clk(gclk));
	jdff dff_B_T7oGcoNR3_2(.din(w_dff_B_HzuHDBeP6_2),.dout(w_dff_B_T7oGcoNR3_2),.clk(gclk));
	jdff dff_B_VQjfX0IM0_2(.din(w_dff_B_T7oGcoNR3_2),.dout(w_dff_B_VQjfX0IM0_2),.clk(gclk));
	jdff dff_B_h9BWaBXz0_2(.din(w_dff_B_VQjfX0IM0_2),.dout(w_dff_B_h9BWaBXz0_2),.clk(gclk));
	jdff dff_B_bTqfafHR7_2(.din(w_dff_B_h9BWaBXz0_2),.dout(w_dff_B_bTqfafHR7_2),.clk(gclk));
	jdff dff_B_VMReU0S91_2(.din(w_dff_B_bTqfafHR7_2),.dout(w_dff_B_VMReU0S91_2),.clk(gclk));
	jdff dff_B_P0hUCw0P0_2(.din(w_dff_B_VMReU0S91_2),.dout(w_dff_B_P0hUCw0P0_2),.clk(gclk));
	jdff dff_B_1HrcFrfi5_2(.din(w_dff_B_P0hUCw0P0_2),.dout(w_dff_B_1HrcFrfi5_2),.clk(gclk));
	jdff dff_B_uesnWeIG6_2(.din(w_dff_B_1HrcFrfi5_2),.dout(w_dff_B_uesnWeIG6_2),.clk(gclk));
	jdff dff_B_vy6soyIt7_2(.din(w_dff_B_uesnWeIG6_2),.dout(w_dff_B_vy6soyIt7_2),.clk(gclk));
	jdff dff_B_2MKAJuKf8_2(.din(w_dff_B_vy6soyIt7_2),.dout(w_dff_B_2MKAJuKf8_2),.clk(gclk));
	jdff dff_B_kZu3kG5s9_2(.din(w_dff_B_2MKAJuKf8_2),.dout(w_dff_B_kZu3kG5s9_2),.clk(gclk));
	jdff dff_B_IXH8WcCY9_2(.din(w_dff_B_kZu3kG5s9_2),.dout(w_dff_B_IXH8WcCY9_2),.clk(gclk));
	jdff dff_B_WjKF1KD99_2(.din(w_dff_B_IXH8WcCY9_2),.dout(w_dff_B_WjKF1KD99_2),.clk(gclk));
	jdff dff_B_Dplf3ms51_2(.din(w_dff_B_WjKF1KD99_2),.dout(w_dff_B_Dplf3ms51_2),.clk(gclk));
	jdff dff_B_toTQhYKo8_2(.din(w_dff_B_Dplf3ms51_2),.dout(w_dff_B_toTQhYKo8_2),.clk(gclk));
	jdff dff_B_ibv82bX53_2(.din(w_dff_B_toTQhYKo8_2),.dout(w_dff_B_ibv82bX53_2),.clk(gclk));
	jdff dff_B_jfiRjN7D4_2(.din(w_dff_B_ibv82bX53_2),.dout(w_dff_B_jfiRjN7D4_2),.clk(gclk));
	jdff dff_B_u8pQr0sd9_2(.din(w_dff_B_jfiRjN7D4_2),.dout(w_dff_B_u8pQr0sd9_2),.clk(gclk));
	jdff dff_B_WzRyQTej3_2(.din(w_dff_B_u8pQr0sd9_2),.dout(w_dff_B_WzRyQTej3_2),.clk(gclk));
	jdff dff_B_ZqudcncV3_2(.din(w_dff_B_WzRyQTej3_2),.dout(w_dff_B_ZqudcncV3_2),.clk(gclk));
	jdff dff_B_Mv27uzwL3_2(.din(w_dff_B_ZqudcncV3_2),.dout(w_dff_B_Mv27uzwL3_2),.clk(gclk));
	jdff dff_B_9duGwFgx7_2(.din(w_dff_B_Mv27uzwL3_2),.dout(w_dff_B_9duGwFgx7_2),.clk(gclk));
	jdff dff_B_rVOXfMG23_2(.din(w_dff_B_9duGwFgx7_2),.dout(w_dff_B_rVOXfMG23_2),.clk(gclk));
	jdff dff_B_9zZnf4xZ4_2(.din(w_dff_B_rVOXfMG23_2),.dout(w_dff_B_9zZnf4xZ4_2),.clk(gclk));
	jdff dff_B_pICOT8mK6_2(.din(w_dff_B_9zZnf4xZ4_2),.dout(w_dff_B_pICOT8mK6_2),.clk(gclk));
	jdff dff_B_mZ2Pe8Zs1_2(.din(w_dff_B_pICOT8mK6_2),.dout(w_dff_B_mZ2Pe8Zs1_2),.clk(gclk));
	jdff dff_B_5VafzWNx4_2(.din(w_dff_B_mZ2Pe8Zs1_2),.dout(w_dff_B_5VafzWNx4_2),.clk(gclk));
	jdff dff_B_T20zpEtB5_2(.din(w_dff_B_5VafzWNx4_2),.dout(w_dff_B_T20zpEtB5_2),.clk(gclk));
	jdff dff_B_naGH2sfc0_2(.din(w_dff_B_T20zpEtB5_2),.dout(w_dff_B_naGH2sfc0_2),.clk(gclk));
	jdff dff_B_SmYMYUcR2_2(.din(w_dff_B_naGH2sfc0_2),.dout(w_dff_B_SmYMYUcR2_2),.clk(gclk));
	jdff dff_B_dfywWW1T7_2(.din(w_dff_B_SmYMYUcR2_2),.dout(w_dff_B_dfywWW1T7_2),.clk(gclk));
	jdff dff_B_FSTInDsE4_2(.din(w_dff_B_dfywWW1T7_2),.dout(w_dff_B_FSTInDsE4_2),.clk(gclk));
	jdff dff_B_oU7SjGEV6_2(.din(w_dff_B_FSTInDsE4_2),.dout(w_dff_B_oU7SjGEV6_2),.clk(gclk));
	jdff dff_B_DhItVa4b0_2(.din(w_dff_B_oU7SjGEV6_2),.dout(w_dff_B_DhItVa4b0_2),.clk(gclk));
	jdff dff_B_DM4qzMub8_2(.din(w_dff_B_DhItVa4b0_2),.dout(w_dff_B_DM4qzMub8_2),.clk(gclk));
	jdff dff_B_jr1AaHBJ1_2(.din(w_dff_B_DM4qzMub8_2),.dout(w_dff_B_jr1AaHBJ1_2),.clk(gclk));
	jdff dff_B_OBes7WtX2_2(.din(w_dff_B_jr1AaHBJ1_2),.dout(w_dff_B_OBes7WtX2_2),.clk(gclk));
	jdff dff_B_iJMIQNGM2_2(.din(w_dff_B_OBes7WtX2_2),.dout(w_dff_B_iJMIQNGM2_2),.clk(gclk));
	jdff dff_B_OgRPnqI63_2(.din(w_dff_B_iJMIQNGM2_2),.dout(w_dff_B_OgRPnqI63_2),.clk(gclk));
	jdff dff_B_TLbaPM3u0_2(.din(w_dff_B_OgRPnqI63_2),.dout(w_dff_B_TLbaPM3u0_2),.clk(gclk));
	jdff dff_B_OzTc8R7Z8_2(.din(n1548),.dout(w_dff_B_OzTc8R7Z8_2),.clk(gclk));
	jdff dff_B_aRK956Io7_1(.din(n1503),.dout(w_dff_B_aRK956Io7_1),.clk(gclk));
	jdff dff_B_7OEaWOFM5_2(.din(n1431),.dout(w_dff_B_7OEaWOFM5_2),.clk(gclk));
	jdff dff_B_vbdHOdD61_2(.din(w_dff_B_7OEaWOFM5_2),.dout(w_dff_B_vbdHOdD61_2),.clk(gclk));
	jdff dff_B_MgOg3O739_2(.din(w_dff_B_vbdHOdD61_2),.dout(w_dff_B_MgOg3O739_2),.clk(gclk));
	jdff dff_B_r3VCoTHa5_2(.din(w_dff_B_MgOg3O739_2),.dout(w_dff_B_r3VCoTHa5_2),.clk(gclk));
	jdff dff_B_4L3JdPvB6_2(.din(w_dff_B_r3VCoTHa5_2),.dout(w_dff_B_4L3JdPvB6_2),.clk(gclk));
	jdff dff_B_slHNYECG7_2(.din(w_dff_B_4L3JdPvB6_2),.dout(w_dff_B_slHNYECG7_2),.clk(gclk));
	jdff dff_B_xEOONrcV2_2(.din(w_dff_B_slHNYECG7_2),.dout(w_dff_B_xEOONrcV2_2),.clk(gclk));
	jdff dff_B_bwZdFMpz3_2(.din(w_dff_B_xEOONrcV2_2),.dout(w_dff_B_bwZdFMpz3_2),.clk(gclk));
	jdff dff_B_zrS0wVTp4_2(.din(w_dff_B_bwZdFMpz3_2),.dout(w_dff_B_zrS0wVTp4_2),.clk(gclk));
	jdff dff_B_BgugZ0gV1_2(.din(w_dff_B_zrS0wVTp4_2),.dout(w_dff_B_BgugZ0gV1_2),.clk(gclk));
	jdff dff_B_39Q4ytw93_2(.din(w_dff_B_BgugZ0gV1_2),.dout(w_dff_B_39Q4ytw93_2),.clk(gclk));
	jdff dff_B_Ir3EyOh10_2(.din(w_dff_B_39Q4ytw93_2),.dout(w_dff_B_Ir3EyOh10_2),.clk(gclk));
	jdff dff_B_x6LYUNE72_2(.din(w_dff_B_Ir3EyOh10_2),.dout(w_dff_B_x6LYUNE72_2),.clk(gclk));
	jdff dff_B_lNsOoBoq9_2(.din(w_dff_B_x6LYUNE72_2),.dout(w_dff_B_lNsOoBoq9_2),.clk(gclk));
	jdff dff_B_MK4LfCtl3_2(.din(w_dff_B_lNsOoBoq9_2),.dout(w_dff_B_MK4LfCtl3_2),.clk(gclk));
	jdff dff_B_nNNIllSw4_2(.din(w_dff_B_MK4LfCtl3_2),.dout(w_dff_B_nNNIllSw4_2),.clk(gclk));
	jdff dff_B_ORf6ql5j2_2(.din(w_dff_B_nNNIllSw4_2),.dout(w_dff_B_ORf6ql5j2_2),.clk(gclk));
	jdff dff_B_VpXoKOYz5_2(.din(w_dff_B_ORf6ql5j2_2),.dout(w_dff_B_VpXoKOYz5_2),.clk(gclk));
	jdff dff_B_praYt60y0_2(.din(w_dff_B_VpXoKOYz5_2),.dout(w_dff_B_praYt60y0_2),.clk(gclk));
	jdff dff_B_uUTCZeEs8_2(.din(w_dff_B_praYt60y0_2),.dout(w_dff_B_uUTCZeEs8_2),.clk(gclk));
	jdff dff_B_aAIaCyAP8_2(.din(w_dff_B_uUTCZeEs8_2),.dout(w_dff_B_aAIaCyAP8_2),.clk(gclk));
	jdff dff_B_l5uhyDoT0_2(.din(w_dff_B_aAIaCyAP8_2),.dout(w_dff_B_l5uhyDoT0_2),.clk(gclk));
	jdff dff_B_gUGeMuOa0_2(.din(w_dff_B_l5uhyDoT0_2),.dout(w_dff_B_gUGeMuOa0_2),.clk(gclk));
	jdff dff_B_0vH9r3UA2_2(.din(w_dff_B_gUGeMuOa0_2),.dout(w_dff_B_0vH9r3UA2_2),.clk(gclk));
	jdff dff_B_QPujcOcK3_2(.din(w_dff_B_0vH9r3UA2_2),.dout(w_dff_B_QPujcOcK3_2),.clk(gclk));
	jdff dff_B_uXk0qGrU1_2(.din(w_dff_B_QPujcOcK3_2),.dout(w_dff_B_uXk0qGrU1_2),.clk(gclk));
	jdff dff_B_Cd5vAkuo7_2(.din(w_dff_B_uXk0qGrU1_2),.dout(w_dff_B_Cd5vAkuo7_2),.clk(gclk));
	jdff dff_B_HrNndOAC0_2(.din(w_dff_B_Cd5vAkuo7_2),.dout(w_dff_B_HrNndOAC0_2),.clk(gclk));
	jdff dff_B_ZjZLhMMJ0_2(.din(w_dff_B_HrNndOAC0_2),.dout(w_dff_B_ZjZLhMMJ0_2),.clk(gclk));
	jdff dff_B_NA0zjnQs9_2(.din(w_dff_B_ZjZLhMMJ0_2),.dout(w_dff_B_NA0zjnQs9_2),.clk(gclk));
	jdff dff_B_bKvuNu7H1_2(.din(w_dff_B_NA0zjnQs9_2),.dout(w_dff_B_bKvuNu7H1_2),.clk(gclk));
	jdff dff_B_anbhfeed7_2(.din(w_dff_B_bKvuNu7H1_2),.dout(w_dff_B_anbhfeed7_2),.clk(gclk));
	jdff dff_B_TyEoFMTR6_2(.din(w_dff_B_anbhfeed7_2),.dout(w_dff_B_TyEoFMTR6_2),.clk(gclk));
	jdff dff_B_brb85nqy7_2(.din(w_dff_B_TyEoFMTR6_2),.dout(w_dff_B_brb85nqy7_2),.clk(gclk));
	jdff dff_B_t1hNhFKR7_2(.din(w_dff_B_brb85nqy7_2),.dout(w_dff_B_t1hNhFKR7_2),.clk(gclk));
	jdff dff_B_A552WBmt3_2(.din(w_dff_B_t1hNhFKR7_2),.dout(w_dff_B_A552WBmt3_2),.clk(gclk));
	jdff dff_B_0G3AblGa3_2(.din(w_dff_B_A552WBmt3_2),.dout(w_dff_B_0G3AblGa3_2),.clk(gclk));
	jdff dff_B_Lrp9Mhk18_2(.din(w_dff_B_0G3AblGa3_2),.dout(w_dff_B_Lrp9Mhk18_2),.clk(gclk));
	jdff dff_B_xqaVoTr96_2(.din(w_dff_B_Lrp9Mhk18_2),.dout(w_dff_B_xqaVoTr96_2),.clk(gclk));
	jdff dff_B_gCURn5tp9_2(.din(n1477),.dout(w_dff_B_gCURn5tp9_2),.clk(gclk));
	jdff dff_B_BlR6EJkB2_1(.din(n1432),.dout(w_dff_B_BlR6EJkB2_1),.clk(gclk));
	jdff dff_B_AZN01NqR1_2(.din(n1353),.dout(w_dff_B_AZN01NqR1_2),.clk(gclk));
	jdff dff_B_HarpwzLK1_2(.din(w_dff_B_AZN01NqR1_2),.dout(w_dff_B_HarpwzLK1_2),.clk(gclk));
	jdff dff_B_RRrPOGVW4_2(.din(w_dff_B_HarpwzLK1_2),.dout(w_dff_B_RRrPOGVW4_2),.clk(gclk));
	jdff dff_B_uXVhy4AP5_2(.din(w_dff_B_RRrPOGVW4_2),.dout(w_dff_B_uXVhy4AP5_2),.clk(gclk));
	jdff dff_B_CqD4oQ3g5_2(.din(w_dff_B_uXVhy4AP5_2),.dout(w_dff_B_CqD4oQ3g5_2),.clk(gclk));
	jdff dff_B_7EUXIAYI3_2(.din(w_dff_B_CqD4oQ3g5_2),.dout(w_dff_B_7EUXIAYI3_2),.clk(gclk));
	jdff dff_B_o1Nf8nId1_2(.din(w_dff_B_7EUXIAYI3_2),.dout(w_dff_B_o1Nf8nId1_2),.clk(gclk));
	jdff dff_B_XCXBjBFW6_2(.din(w_dff_B_o1Nf8nId1_2),.dout(w_dff_B_XCXBjBFW6_2),.clk(gclk));
	jdff dff_B_kmLVOZc66_2(.din(w_dff_B_XCXBjBFW6_2),.dout(w_dff_B_kmLVOZc66_2),.clk(gclk));
	jdff dff_B_aUlj0tMX7_2(.din(w_dff_B_kmLVOZc66_2),.dout(w_dff_B_aUlj0tMX7_2),.clk(gclk));
	jdff dff_B_VjgxiZoj7_2(.din(w_dff_B_aUlj0tMX7_2),.dout(w_dff_B_VjgxiZoj7_2),.clk(gclk));
	jdff dff_B_4AaBljX49_2(.din(w_dff_B_VjgxiZoj7_2),.dout(w_dff_B_4AaBljX49_2),.clk(gclk));
	jdff dff_B_FHdesKAm3_2(.din(w_dff_B_4AaBljX49_2),.dout(w_dff_B_FHdesKAm3_2),.clk(gclk));
	jdff dff_B_dkpHPHTX8_2(.din(w_dff_B_FHdesKAm3_2),.dout(w_dff_B_dkpHPHTX8_2),.clk(gclk));
	jdff dff_B_NSvE7o3u9_2(.din(w_dff_B_dkpHPHTX8_2),.dout(w_dff_B_NSvE7o3u9_2),.clk(gclk));
	jdff dff_B_Kvrrxyx49_2(.din(w_dff_B_NSvE7o3u9_2),.dout(w_dff_B_Kvrrxyx49_2),.clk(gclk));
	jdff dff_B_t3NzRcBg1_2(.din(w_dff_B_Kvrrxyx49_2),.dout(w_dff_B_t3NzRcBg1_2),.clk(gclk));
	jdff dff_B_5gohuiQp0_2(.din(w_dff_B_t3NzRcBg1_2),.dout(w_dff_B_5gohuiQp0_2),.clk(gclk));
	jdff dff_B_eCKb4z697_2(.din(w_dff_B_5gohuiQp0_2),.dout(w_dff_B_eCKb4z697_2),.clk(gclk));
	jdff dff_B_4T2rRRjW8_2(.din(w_dff_B_eCKb4z697_2),.dout(w_dff_B_4T2rRRjW8_2),.clk(gclk));
	jdff dff_B_v8jP46p51_2(.din(w_dff_B_4T2rRRjW8_2),.dout(w_dff_B_v8jP46p51_2),.clk(gclk));
	jdff dff_B_mQDVsplr8_2(.din(w_dff_B_v8jP46p51_2),.dout(w_dff_B_mQDVsplr8_2),.clk(gclk));
	jdff dff_B_XRcFEKP07_2(.din(w_dff_B_mQDVsplr8_2),.dout(w_dff_B_XRcFEKP07_2),.clk(gclk));
	jdff dff_B_miN0aHYX5_2(.din(w_dff_B_XRcFEKP07_2),.dout(w_dff_B_miN0aHYX5_2),.clk(gclk));
	jdff dff_B_f8tEK2dq2_2(.din(w_dff_B_miN0aHYX5_2),.dout(w_dff_B_f8tEK2dq2_2),.clk(gclk));
	jdff dff_B_KUJuGNsV2_2(.din(w_dff_B_f8tEK2dq2_2),.dout(w_dff_B_KUJuGNsV2_2),.clk(gclk));
	jdff dff_B_pHDRcmR51_2(.din(w_dff_B_KUJuGNsV2_2),.dout(w_dff_B_pHDRcmR51_2),.clk(gclk));
	jdff dff_B_YHtoN35Y2_2(.din(w_dff_B_pHDRcmR51_2),.dout(w_dff_B_YHtoN35Y2_2),.clk(gclk));
	jdff dff_B_nisqSuFC3_2(.din(w_dff_B_YHtoN35Y2_2),.dout(w_dff_B_nisqSuFC3_2),.clk(gclk));
	jdff dff_B_Vcs2YyyL3_2(.din(w_dff_B_nisqSuFC3_2),.dout(w_dff_B_Vcs2YyyL3_2),.clk(gclk));
	jdff dff_B_YRJXmm4d1_2(.din(w_dff_B_Vcs2YyyL3_2),.dout(w_dff_B_YRJXmm4d1_2),.clk(gclk));
	jdff dff_B_avE36V7U8_2(.din(w_dff_B_YRJXmm4d1_2),.dout(w_dff_B_avE36V7U8_2),.clk(gclk));
	jdff dff_B_gupLnxqX3_2(.din(w_dff_B_avE36V7U8_2),.dout(w_dff_B_gupLnxqX3_2),.clk(gclk));
	jdff dff_B_enY74l0d2_2(.din(w_dff_B_gupLnxqX3_2),.dout(w_dff_B_enY74l0d2_2),.clk(gclk));
	jdff dff_B_xEAcDscs6_2(.din(w_dff_B_enY74l0d2_2),.dout(w_dff_B_xEAcDscs6_2),.clk(gclk));
	jdff dff_B_Patk0o6B2_2(.din(w_dff_B_xEAcDscs6_2),.dout(w_dff_B_Patk0o6B2_2),.clk(gclk));
	jdff dff_B_PpKZCrKf2_2(.din(n1399),.dout(w_dff_B_PpKZCrKf2_2),.clk(gclk));
	jdff dff_B_FzF9b9Ge7_1(.din(n1354),.dout(w_dff_B_FzF9b9Ge7_1),.clk(gclk));
	jdff dff_B_lPFQZYYF1_2(.din(n1268),.dout(w_dff_B_lPFQZYYF1_2),.clk(gclk));
	jdff dff_B_iJQN5Sud1_2(.din(w_dff_B_lPFQZYYF1_2),.dout(w_dff_B_iJQN5Sud1_2),.clk(gclk));
	jdff dff_B_zSCAmNSA4_2(.din(w_dff_B_iJQN5Sud1_2),.dout(w_dff_B_zSCAmNSA4_2),.clk(gclk));
	jdff dff_B_TbaZtBKf4_2(.din(w_dff_B_zSCAmNSA4_2),.dout(w_dff_B_TbaZtBKf4_2),.clk(gclk));
	jdff dff_B_pgY9WjaR5_2(.din(w_dff_B_TbaZtBKf4_2),.dout(w_dff_B_pgY9WjaR5_2),.clk(gclk));
	jdff dff_B_i2miKn7D5_2(.din(w_dff_B_pgY9WjaR5_2),.dout(w_dff_B_i2miKn7D5_2),.clk(gclk));
	jdff dff_B_dwGCvwxX2_2(.din(w_dff_B_i2miKn7D5_2),.dout(w_dff_B_dwGCvwxX2_2),.clk(gclk));
	jdff dff_B_nCRjsMjQ9_2(.din(w_dff_B_dwGCvwxX2_2),.dout(w_dff_B_nCRjsMjQ9_2),.clk(gclk));
	jdff dff_B_tVoIQ5wF4_2(.din(w_dff_B_nCRjsMjQ9_2),.dout(w_dff_B_tVoIQ5wF4_2),.clk(gclk));
	jdff dff_B_I9YAnaHK0_2(.din(w_dff_B_tVoIQ5wF4_2),.dout(w_dff_B_I9YAnaHK0_2),.clk(gclk));
	jdff dff_B_FbkEBOwC4_2(.din(w_dff_B_I9YAnaHK0_2),.dout(w_dff_B_FbkEBOwC4_2),.clk(gclk));
	jdff dff_B_vaBNNtNn3_2(.din(w_dff_B_FbkEBOwC4_2),.dout(w_dff_B_vaBNNtNn3_2),.clk(gclk));
	jdff dff_B_LbtjHO9Z6_2(.din(w_dff_B_vaBNNtNn3_2),.dout(w_dff_B_LbtjHO9Z6_2),.clk(gclk));
	jdff dff_B_UHx5HpJW3_2(.din(w_dff_B_LbtjHO9Z6_2),.dout(w_dff_B_UHx5HpJW3_2),.clk(gclk));
	jdff dff_B_oMYBigI99_2(.din(w_dff_B_UHx5HpJW3_2),.dout(w_dff_B_oMYBigI99_2),.clk(gclk));
	jdff dff_B_0VTcO1vk3_2(.din(w_dff_B_oMYBigI99_2),.dout(w_dff_B_0VTcO1vk3_2),.clk(gclk));
	jdff dff_B_s0tQSQD75_2(.din(w_dff_B_0VTcO1vk3_2),.dout(w_dff_B_s0tQSQD75_2),.clk(gclk));
	jdff dff_B_cxYAnOAR4_2(.din(w_dff_B_s0tQSQD75_2),.dout(w_dff_B_cxYAnOAR4_2),.clk(gclk));
	jdff dff_B_Jc4RGxH64_2(.din(w_dff_B_cxYAnOAR4_2),.dout(w_dff_B_Jc4RGxH64_2),.clk(gclk));
	jdff dff_B_XfhYZyNu6_2(.din(w_dff_B_Jc4RGxH64_2),.dout(w_dff_B_XfhYZyNu6_2),.clk(gclk));
	jdff dff_B_YH5mPmX65_2(.din(w_dff_B_XfhYZyNu6_2),.dout(w_dff_B_YH5mPmX65_2),.clk(gclk));
	jdff dff_B_bZMqbk7c3_2(.din(w_dff_B_YH5mPmX65_2),.dout(w_dff_B_bZMqbk7c3_2),.clk(gclk));
	jdff dff_B_PKKC6atd7_2(.din(w_dff_B_bZMqbk7c3_2),.dout(w_dff_B_PKKC6atd7_2),.clk(gclk));
	jdff dff_B_wAHjK5OM4_2(.din(w_dff_B_PKKC6atd7_2),.dout(w_dff_B_wAHjK5OM4_2),.clk(gclk));
	jdff dff_B_Iw5ueGsH7_2(.din(w_dff_B_wAHjK5OM4_2),.dout(w_dff_B_Iw5ueGsH7_2),.clk(gclk));
	jdff dff_B_BOUJUf7R6_2(.din(w_dff_B_Iw5ueGsH7_2),.dout(w_dff_B_BOUJUf7R6_2),.clk(gclk));
	jdff dff_B_YeExXbwh8_2(.din(w_dff_B_BOUJUf7R6_2),.dout(w_dff_B_YeExXbwh8_2),.clk(gclk));
	jdff dff_B_lAYEKKoZ4_2(.din(w_dff_B_YeExXbwh8_2),.dout(w_dff_B_lAYEKKoZ4_2),.clk(gclk));
	jdff dff_B_mLTDj1ur8_2(.din(w_dff_B_lAYEKKoZ4_2),.dout(w_dff_B_mLTDj1ur8_2),.clk(gclk));
	jdff dff_B_8oYXsYGA1_2(.din(w_dff_B_mLTDj1ur8_2),.dout(w_dff_B_8oYXsYGA1_2),.clk(gclk));
	jdff dff_B_VggqWUL69_2(.din(w_dff_B_8oYXsYGA1_2),.dout(w_dff_B_VggqWUL69_2),.clk(gclk));
	jdff dff_B_swd6VmrS0_2(.din(w_dff_B_VggqWUL69_2),.dout(w_dff_B_swd6VmrS0_2),.clk(gclk));
	jdff dff_B_20xgkSPY9_2(.din(w_dff_B_swd6VmrS0_2),.dout(w_dff_B_20xgkSPY9_2),.clk(gclk));
	jdff dff_B_xSk7omfA1_2(.din(n1314),.dout(w_dff_B_xSk7omfA1_2),.clk(gclk));
	jdff dff_B_ScPyrVF34_1(.din(n1269),.dout(w_dff_B_ScPyrVF34_1),.clk(gclk));
	jdff dff_B_sFiR5tEY5_2(.din(n1178),.dout(w_dff_B_sFiR5tEY5_2),.clk(gclk));
	jdff dff_B_UnPw4Kie4_2(.din(w_dff_B_sFiR5tEY5_2),.dout(w_dff_B_UnPw4Kie4_2),.clk(gclk));
	jdff dff_B_ohWgRbZY0_2(.din(w_dff_B_UnPw4Kie4_2),.dout(w_dff_B_ohWgRbZY0_2),.clk(gclk));
	jdff dff_B_ZLwjlKpF3_2(.din(w_dff_B_ohWgRbZY0_2),.dout(w_dff_B_ZLwjlKpF3_2),.clk(gclk));
	jdff dff_B_6F7TUjP04_2(.din(w_dff_B_ZLwjlKpF3_2),.dout(w_dff_B_6F7TUjP04_2),.clk(gclk));
	jdff dff_B_HZv5SsZW7_2(.din(w_dff_B_6F7TUjP04_2),.dout(w_dff_B_HZv5SsZW7_2),.clk(gclk));
	jdff dff_B_1XqV9wbH1_2(.din(w_dff_B_HZv5SsZW7_2),.dout(w_dff_B_1XqV9wbH1_2),.clk(gclk));
	jdff dff_B_f92aTyxH2_2(.din(w_dff_B_1XqV9wbH1_2),.dout(w_dff_B_f92aTyxH2_2),.clk(gclk));
	jdff dff_B_3OWiSrvp2_2(.din(w_dff_B_f92aTyxH2_2),.dout(w_dff_B_3OWiSrvp2_2),.clk(gclk));
	jdff dff_B_DK6jW7Me2_2(.din(w_dff_B_3OWiSrvp2_2),.dout(w_dff_B_DK6jW7Me2_2),.clk(gclk));
	jdff dff_B_F2LSVmmD7_2(.din(w_dff_B_DK6jW7Me2_2),.dout(w_dff_B_F2LSVmmD7_2),.clk(gclk));
	jdff dff_B_3eVzFBCr0_2(.din(w_dff_B_F2LSVmmD7_2),.dout(w_dff_B_3eVzFBCr0_2),.clk(gclk));
	jdff dff_B_DdwjIYGD6_2(.din(w_dff_B_3eVzFBCr0_2),.dout(w_dff_B_DdwjIYGD6_2),.clk(gclk));
	jdff dff_B_h9UXEoPm3_2(.din(w_dff_B_DdwjIYGD6_2),.dout(w_dff_B_h9UXEoPm3_2),.clk(gclk));
	jdff dff_B_rs5s9YpB4_2(.din(w_dff_B_h9UXEoPm3_2),.dout(w_dff_B_rs5s9YpB4_2),.clk(gclk));
	jdff dff_B_SZ1YAXcV1_2(.din(w_dff_B_rs5s9YpB4_2),.dout(w_dff_B_SZ1YAXcV1_2),.clk(gclk));
	jdff dff_B_rDpriOgC5_2(.din(w_dff_B_SZ1YAXcV1_2),.dout(w_dff_B_rDpriOgC5_2),.clk(gclk));
	jdff dff_B_uqTahcw47_2(.din(w_dff_B_rDpriOgC5_2),.dout(w_dff_B_uqTahcw47_2),.clk(gclk));
	jdff dff_B_bsdKYveB5_2(.din(w_dff_B_uqTahcw47_2),.dout(w_dff_B_bsdKYveB5_2),.clk(gclk));
	jdff dff_B_ga8Y9ufL9_2(.din(w_dff_B_bsdKYveB5_2),.dout(w_dff_B_ga8Y9ufL9_2),.clk(gclk));
	jdff dff_B_IdXGlFdY1_2(.din(w_dff_B_ga8Y9ufL9_2),.dout(w_dff_B_IdXGlFdY1_2),.clk(gclk));
	jdff dff_B_jxx4Skw51_2(.din(w_dff_B_IdXGlFdY1_2),.dout(w_dff_B_jxx4Skw51_2),.clk(gclk));
	jdff dff_B_KDyzA9ow3_2(.din(w_dff_B_jxx4Skw51_2),.dout(w_dff_B_KDyzA9ow3_2),.clk(gclk));
	jdff dff_B_EApnyhfk6_2(.din(w_dff_B_KDyzA9ow3_2),.dout(w_dff_B_EApnyhfk6_2),.clk(gclk));
	jdff dff_B_I2hBWnyA5_2(.din(w_dff_B_EApnyhfk6_2),.dout(w_dff_B_I2hBWnyA5_2),.clk(gclk));
	jdff dff_B_7uvoe9dF3_2(.din(w_dff_B_I2hBWnyA5_2),.dout(w_dff_B_7uvoe9dF3_2),.clk(gclk));
	jdff dff_B_kwO31D1A2_2(.din(w_dff_B_7uvoe9dF3_2),.dout(w_dff_B_kwO31D1A2_2),.clk(gclk));
	jdff dff_B_g3DsQ5Nu8_2(.din(w_dff_B_kwO31D1A2_2),.dout(w_dff_B_g3DsQ5Nu8_2),.clk(gclk));
	jdff dff_B_Lnnx9r0k6_2(.din(w_dff_B_g3DsQ5Nu8_2),.dout(w_dff_B_Lnnx9r0k6_2),.clk(gclk));
	jdff dff_B_2l75t1df1_2(.din(w_dff_B_Lnnx9r0k6_2),.dout(w_dff_B_2l75t1df1_2),.clk(gclk));
	jdff dff_B_06mQNvWb6_2(.din(n1223),.dout(w_dff_B_06mQNvWb6_2),.clk(gclk));
	jdff dff_B_buQPiXvj6_1(.din(n1179),.dout(w_dff_B_buQPiXvj6_1),.clk(gclk));
	jdff dff_B_lKOzpYjF5_2(.din(n1074),.dout(w_dff_B_lKOzpYjF5_2),.clk(gclk));
	jdff dff_B_QtOqGyEj6_2(.din(w_dff_B_lKOzpYjF5_2),.dout(w_dff_B_QtOqGyEj6_2),.clk(gclk));
	jdff dff_B_vXbR900i4_2(.din(w_dff_B_QtOqGyEj6_2),.dout(w_dff_B_vXbR900i4_2),.clk(gclk));
	jdff dff_B_PJZ4Sj7W5_2(.din(w_dff_B_vXbR900i4_2),.dout(w_dff_B_PJZ4Sj7W5_2),.clk(gclk));
	jdff dff_B_5zxKD1uS1_2(.din(w_dff_B_PJZ4Sj7W5_2),.dout(w_dff_B_5zxKD1uS1_2),.clk(gclk));
	jdff dff_B_u5umJbrT3_2(.din(w_dff_B_5zxKD1uS1_2),.dout(w_dff_B_u5umJbrT3_2),.clk(gclk));
	jdff dff_B_4DbieKDR6_2(.din(w_dff_B_u5umJbrT3_2),.dout(w_dff_B_4DbieKDR6_2),.clk(gclk));
	jdff dff_B_8Xc0qH8Q7_2(.din(w_dff_B_4DbieKDR6_2),.dout(w_dff_B_8Xc0qH8Q7_2),.clk(gclk));
	jdff dff_B_3IwaWNBe9_2(.din(w_dff_B_8Xc0qH8Q7_2),.dout(w_dff_B_3IwaWNBe9_2),.clk(gclk));
	jdff dff_B_lstUPp760_2(.din(w_dff_B_3IwaWNBe9_2),.dout(w_dff_B_lstUPp760_2),.clk(gclk));
	jdff dff_B_ObUwMK1Z5_2(.din(w_dff_B_lstUPp760_2),.dout(w_dff_B_ObUwMK1Z5_2),.clk(gclk));
	jdff dff_B_SEy8Udo97_2(.din(w_dff_B_ObUwMK1Z5_2),.dout(w_dff_B_SEy8Udo97_2),.clk(gclk));
	jdff dff_B_E2Sd5Uo40_2(.din(w_dff_B_SEy8Udo97_2),.dout(w_dff_B_E2Sd5Uo40_2),.clk(gclk));
	jdff dff_B_hVoxkf8Y0_2(.din(w_dff_B_E2Sd5Uo40_2),.dout(w_dff_B_hVoxkf8Y0_2),.clk(gclk));
	jdff dff_B_uly6CBGn7_2(.din(w_dff_B_hVoxkf8Y0_2),.dout(w_dff_B_uly6CBGn7_2),.clk(gclk));
	jdff dff_B_VNy9mvCG3_2(.din(w_dff_B_uly6CBGn7_2),.dout(w_dff_B_VNy9mvCG3_2),.clk(gclk));
	jdff dff_B_osQLCnzQ4_2(.din(w_dff_B_VNy9mvCG3_2),.dout(w_dff_B_osQLCnzQ4_2),.clk(gclk));
	jdff dff_B_zV4r5tJg0_2(.din(w_dff_B_osQLCnzQ4_2),.dout(w_dff_B_zV4r5tJg0_2),.clk(gclk));
	jdff dff_B_V8ecpqJ66_2(.din(w_dff_B_zV4r5tJg0_2),.dout(w_dff_B_V8ecpqJ66_2),.clk(gclk));
	jdff dff_B_97GtppLO6_2(.din(w_dff_B_V8ecpqJ66_2),.dout(w_dff_B_97GtppLO6_2),.clk(gclk));
	jdff dff_B_cCGH2UfC9_2(.din(w_dff_B_97GtppLO6_2),.dout(w_dff_B_cCGH2UfC9_2),.clk(gclk));
	jdff dff_B_LegMgFmk3_2(.din(w_dff_B_cCGH2UfC9_2),.dout(w_dff_B_LegMgFmk3_2),.clk(gclk));
	jdff dff_B_ugYc6VgR7_2(.din(w_dff_B_LegMgFmk3_2),.dout(w_dff_B_ugYc6VgR7_2),.clk(gclk));
	jdff dff_B_IQpYjBsH7_2(.din(w_dff_B_ugYc6VgR7_2),.dout(w_dff_B_IQpYjBsH7_2),.clk(gclk));
	jdff dff_B_HSFqCjXr2_2(.din(w_dff_B_IQpYjBsH7_2),.dout(w_dff_B_HSFqCjXr2_2),.clk(gclk));
	jdff dff_B_vURq43Iq4_2(.din(w_dff_B_HSFqCjXr2_2),.dout(w_dff_B_vURq43Iq4_2),.clk(gclk));
	jdff dff_B_2OVZiyHD6_2(.din(w_dff_B_vURq43Iq4_2),.dout(w_dff_B_2OVZiyHD6_2),.clk(gclk));
	jdff dff_B_o0s09aK91_2(.din(n1125),.dout(w_dff_B_o0s09aK91_2),.clk(gclk));
	jdff dff_B_EkaceZ4V3_1(.din(n1075),.dout(w_dff_B_EkaceZ4V3_1),.clk(gclk));
	jdff dff_B_WZraOng41_2(.din(n976),.dout(w_dff_B_WZraOng41_2),.clk(gclk));
	jdff dff_B_tuXRDdq15_2(.din(w_dff_B_WZraOng41_2),.dout(w_dff_B_tuXRDdq15_2),.clk(gclk));
	jdff dff_B_aV6kqfA96_2(.din(w_dff_B_tuXRDdq15_2),.dout(w_dff_B_aV6kqfA96_2),.clk(gclk));
	jdff dff_B_kbbTU9Lb3_2(.din(w_dff_B_aV6kqfA96_2),.dout(w_dff_B_kbbTU9Lb3_2),.clk(gclk));
	jdff dff_B_rBBeuNnG8_2(.din(w_dff_B_kbbTU9Lb3_2),.dout(w_dff_B_rBBeuNnG8_2),.clk(gclk));
	jdff dff_B_4g6d9G5j8_2(.din(w_dff_B_rBBeuNnG8_2),.dout(w_dff_B_4g6d9G5j8_2),.clk(gclk));
	jdff dff_B_5f7ZHxoN4_2(.din(w_dff_B_4g6d9G5j8_2),.dout(w_dff_B_5f7ZHxoN4_2),.clk(gclk));
	jdff dff_B_2X1I82Bi2_2(.din(w_dff_B_5f7ZHxoN4_2),.dout(w_dff_B_2X1I82Bi2_2),.clk(gclk));
	jdff dff_B_O2ugICkc3_2(.din(w_dff_B_2X1I82Bi2_2),.dout(w_dff_B_O2ugICkc3_2),.clk(gclk));
	jdff dff_B_9aP4QBAP7_2(.din(w_dff_B_O2ugICkc3_2),.dout(w_dff_B_9aP4QBAP7_2),.clk(gclk));
	jdff dff_B_EqxxATn63_2(.din(w_dff_B_9aP4QBAP7_2),.dout(w_dff_B_EqxxATn63_2),.clk(gclk));
	jdff dff_B_aGWVTnKh6_2(.din(w_dff_B_EqxxATn63_2),.dout(w_dff_B_aGWVTnKh6_2),.clk(gclk));
	jdff dff_B_emYZGCaH5_2(.din(w_dff_B_aGWVTnKh6_2),.dout(w_dff_B_emYZGCaH5_2),.clk(gclk));
	jdff dff_B_QDRa7PTO6_2(.din(w_dff_B_emYZGCaH5_2),.dout(w_dff_B_QDRa7PTO6_2),.clk(gclk));
	jdff dff_B_AZXS3gTZ3_2(.din(w_dff_B_QDRa7PTO6_2),.dout(w_dff_B_AZXS3gTZ3_2),.clk(gclk));
	jdff dff_B_cXO8BBRn6_2(.din(w_dff_B_AZXS3gTZ3_2),.dout(w_dff_B_cXO8BBRn6_2),.clk(gclk));
	jdff dff_B_vmkl23lR7_2(.din(w_dff_B_cXO8BBRn6_2),.dout(w_dff_B_vmkl23lR7_2),.clk(gclk));
	jdff dff_B_cLXB7JSd8_2(.din(w_dff_B_vmkl23lR7_2),.dout(w_dff_B_cLXB7JSd8_2),.clk(gclk));
	jdff dff_B_e9xHyCbH4_2(.din(w_dff_B_cLXB7JSd8_2),.dout(w_dff_B_e9xHyCbH4_2),.clk(gclk));
	jdff dff_B_QXk2LXtD6_2(.din(w_dff_B_e9xHyCbH4_2),.dout(w_dff_B_QXk2LXtD6_2),.clk(gclk));
	jdff dff_B_sJ9jJqfW3_2(.din(w_dff_B_QXk2LXtD6_2),.dout(w_dff_B_sJ9jJqfW3_2),.clk(gclk));
	jdff dff_B_XsdUtOc81_2(.din(w_dff_B_sJ9jJqfW3_2),.dout(w_dff_B_XsdUtOc81_2),.clk(gclk));
	jdff dff_B_NIfLEVKF7_2(.din(w_dff_B_XsdUtOc81_2),.dout(w_dff_B_NIfLEVKF7_2),.clk(gclk));
	jdff dff_B_5gsdl4R01_2(.din(w_dff_B_NIfLEVKF7_2),.dout(w_dff_B_5gsdl4R01_2),.clk(gclk));
	jdff dff_B_CuRktE837_2(.din(n1020),.dout(w_dff_B_CuRktE837_2),.clk(gclk));
	jdff dff_B_nncCmUwm5_1(.din(n977),.dout(w_dff_B_nncCmUwm5_1),.clk(gclk));
	jdff dff_B_Wydq4k9Q5_2(.din(n871),.dout(w_dff_B_Wydq4k9Q5_2),.clk(gclk));
	jdff dff_B_QTUOfhUV6_2(.din(w_dff_B_Wydq4k9Q5_2),.dout(w_dff_B_QTUOfhUV6_2),.clk(gclk));
	jdff dff_B_ItN14GvT0_2(.din(w_dff_B_QTUOfhUV6_2),.dout(w_dff_B_ItN14GvT0_2),.clk(gclk));
	jdff dff_B_lJoiSbgk9_2(.din(w_dff_B_ItN14GvT0_2),.dout(w_dff_B_lJoiSbgk9_2),.clk(gclk));
	jdff dff_B_m18D4wSX1_2(.din(w_dff_B_lJoiSbgk9_2),.dout(w_dff_B_m18D4wSX1_2),.clk(gclk));
	jdff dff_B_zbnIlKzT9_2(.din(w_dff_B_m18D4wSX1_2),.dout(w_dff_B_zbnIlKzT9_2),.clk(gclk));
	jdff dff_B_3naIsnxH6_2(.din(w_dff_B_zbnIlKzT9_2),.dout(w_dff_B_3naIsnxH6_2),.clk(gclk));
	jdff dff_B_1CPGJZLE6_2(.din(w_dff_B_3naIsnxH6_2),.dout(w_dff_B_1CPGJZLE6_2),.clk(gclk));
	jdff dff_B_86oTyfjN9_2(.din(w_dff_B_1CPGJZLE6_2),.dout(w_dff_B_86oTyfjN9_2),.clk(gclk));
	jdff dff_B_xPyKY8817_2(.din(w_dff_B_86oTyfjN9_2),.dout(w_dff_B_xPyKY8817_2),.clk(gclk));
	jdff dff_B_9kAEL1bO5_2(.din(w_dff_B_xPyKY8817_2),.dout(w_dff_B_9kAEL1bO5_2),.clk(gclk));
	jdff dff_B_9b3RdcXm4_2(.din(w_dff_B_9kAEL1bO5_2),.dout(w_dff_B_9b3RdcXm4_2),.clk(gclk));
	jdff dff_B_3hpc6nPF2_2(.din(w_dff_B_9b3RdcXm4_2),.dout(w_dff_B_3hpc6nPF2_2),.clk(gclk));
	jdff dff_B_uMtkItIw9_2(.din(w_dff_B_3hpc6nPF2_2),.dout(w_dff_B_uMtkItIw9_2),.clk(gclk));
	jdff dff_B_MKmObVUb1_2(.din(w_dff_B_uMtkItIw9_2),.dout(w_dff_B_MKmObVUb1_2),.clk(gclk));
	jdff dff_B_VuzFrZNL5_2(.din(w_dff_B_MKmObVUb1_2),.dout(w_dff_B_VuzFrZNL5_2),.clk(gclk));
	jdff dff_B_pbb5q2Zf8_2(.din(w_dff_B_VuzFrZNL5_2),.dout(w_dff_B_pbb5q2Zf8_2),.clk(gclk));
	jdff dff_B_wkoLnsZ62_2(.din(w_dff_B_pbb5q2Zf8_2),.dout(w_dff_B_wkoLnsZ62_2),.clk(gclk));
	jdff dff_B_bi7cHT8i5_2(.din(w_dff_B_wkoLnsZ62_2),.dout(w_dff_B_bi7cHT8i5_2),.clk(gclk));
	jdff dff_B_4Kydrbx06_2(.din(w_dff_B_bi7cHT8i5_2),.dout(w_dff_B_4Kydrbx06_2),.clk(gclk));
	jdff dff_B_6nbRevOp8_2(.din(w_dff_B_4Kydrbx06_2),.dout(w_dff_B_6nbRevOp8_2),.clk(gclk));
	jdff dff_B_4QWmYAAQ7_2(.din(n915),.dout(w_dff_B_4QWmYAAQ7_2),.clk(gclk));
	jdff dff_B_jyFNJZ921_1(.din(n872),.dout(w_dff_B_jyFNJZ921_1),.clk(gclk));
	jdff dff_B_lcdzaeZM2_2(.din(n772),.dout(w_dff_B_lcdzaeZM2_2),.clk(gclk));
	jdff dff_B_qaTI2bvq7_2(.din(w_dff_B_lcdzaeZM2_2),.dout(w_dff_B_qaTI2bvq7_2),.clk(gclk));
	jdff dff_B_96YTQVBa9_2(.din(w_dff_B_qaTI2bvq7_2),.dout(w_dff_B_96YTQVBa9_2),.clk(gclk));
	jdff dff_B_TRZdrml47_2(.din(w_dff_B_96YTQVBa9_2),.dout(w_dff_B_TRZdrml47_2),.clk(gclk));
	jdff dff_B_6AYmfj6H6_2(.din(w_dff_B_TRZdrml47_2),.dout(w_dff_B_6AYmfj6H6_2),.clk(gclk));
	jdff dff_B_XuBtdsvm0_2(.din(w_dff_B_6AYmfj6H6_2),.dout(w_dff_B_XuBtdsvm0_2),.clk(gclk));
	jdff dff_B_R5pZwYaa1_2(.din(w_dff_B_XuBtdsvm0_2),.dout(w_dff_B_R5pZwYaa1_2),.clk(gclk));
	jdff dff_B_hBEez6Zn9_2(.din(w_dff_B_R5pZwYaa1_2),.dout(w_dff_B_hBEez6Zn9_2),.clk(gclk));
	jdff dff_B_FNz6hEYy3_2(.din(w_dff_B_hBEez6Zn9_2),.dout(w_dff_B_FNz6hEYy3_2),.clk(gclk));
	jdff dff_B_MuE07MkQ4_2(.din(w_dff_B_FNz6hEYy3_2),.dout(w_dff_B_MuE07MkQ4_2),.clk(gclk));
	jdff dff_B_Yc33j1h25_2(.din(w_dff_B_MuE07MkQ4_2),.dout(w_dff_B_Yc33j1h25_2),.clk(gclk));
	jdff dff_B_xjQuS2G13_2(.din(w_dff_B_Yc33j1h25_2),.dout(w_dff_B_xjQuS2G13_2),.clk(gclk));
	jdff dff_B_Mgmt5gov8_2(.din(w_dff_B_xjQuS2G13_2),.dout(w_dff_B_Mgmt5gov8_2),.clk(gclk));
	jdff dff_B_b5oeM0lI5_2(.din(w_dff_B_Mgmt5gov8_2),.dout(w_dff_B_b5oeM0lI5_2),.clk(gclk));
	jdff dff_B_qgLEczf59_2(.din(w_dff_B_b5oeM0lI5_2),.dout(w_dff_B_qgLEczf59_2),.clk(gclk));
	jdff dff_B_fT5eBe3o3_2(.din(w_dff_B_qgLEczf59_2),.dout(w_dff_B_fT5eBe3o3_2),.clk(gclk));
	jdff dff_B_BaqnRUWR7_2(.din(w_dff_B_fT5eBe3o3_2),.dout(w_dff_B_BaqnRUWR7_2),.clk(gclk));
	jdff dff_B_IgHq9uxs3_2(.din(w_dff_B_BaqnRUWR7_2),.dout(w_dff_B_IgHq9uxs3_2),.clk(gclk));
	jdff dff_B_Z9zB7At31_2(.din(n809),.dout(w_dff_B_Z9zB7At31_2),.clk(gclk));
	jdff dff_B_X2359Wtm1_1(.din(n773),.dout(w_dff_B_X2359Wtm1_1),.clk(gclk));
	jdff dff_B_wHreRi5L3_2(.din(n679),.dout(w_dff_B_wHreRi5L3_2),.clk(gclk));
	jdff dff_B_aF6BvOZO9_2(.din(w_dff_B_wHreRi5L3_2),.dout(w_dff_B_aF6BvOZO9_2),.clk(gclk));
	jdff dff_B_mY8Jb0KE5_2(.din(w_dff_B_aF6BvOZO9_2),.dout(w_dff_B_mY8Jb0KE5_2),.clk(gclk));
	jdff dff_B_6Q0BL26h6_2(.din(w_dff_B_mY8Jb0KE5_2),.dout(w_dff_B_6Q0BL26h6_2),.clk(gclk));
	jdff dff_B_KwP8AI9b1_2(.din(w_dff_B_6Q0BL26h6_2),.dout(w_dff_B_KwP8AI9b1_2),.clk(gclk));
	jdff dff_B_gXZ7ufps6_2(.din(w_dff_B_KwP8AI9b1_2),.dout(w_dff_B_gXZ7ufps6_2),.clk(gclk));
	jdff dff_B_SFGv87qC9_2(.din(w_dff_B_gXZ7ufps6_2),.dout(w_dff_B_SFGv87qC9_2),.clk(gclk));
	jdff dff_B_3SEij5VD0_2(.din(w_dff_B_SFGv87qC9_2),.dout(w_dff_B_3SEij5VD0_2),.clk(gclk));
	jdff dff_B_sME06cnY8_2(.din(w_dff_B_3SEij5VD0_2),.dout(w_dff_B_sME06cnY8_2),.clk(gclk));
	jdff dff_B_OD1yKOzs3_2(.din(w_dff_B_sME06cnY8_2),.dout(w_dff_B_OD1yKOzs3_2),.clk(gclk));
	jdff dff_B_TvCgD8ks9_2(.din(w_dff_B_OD1yKOzs3_2),.dout(w_dff_B_TvCgD8ks9_2),.clk(gclk));
	jdff dff_B_dmQnRqLb9_2(.din(w_dff_B_TvCgD8ks9_2),.dout(w_dff_B_dmQnRqLb9_2),.clk(gclk));
	jdff dff_B_rztMr0lF8_2(.din(w_dff_B_dmQnRqLb9_2),.dout(w_dff_B_rztMr0lF8_2),.clk(gclk));
	jdff dff_B_fzIesVWp9_2(.din(w_dff_B_rztMr0lF8_2),.dout(w_dff_B_fzIesVWp9_2),.clk(gclk));
	jdff dff_B_RJPkQgDR3_2(.din(w_dff_B_fzIesVWp9_2),.dout(w_dff_B_RJPkQgDR3_2),.clk(gclk));
	jdff dff_B_hrRlyOSk0_2(.din(n709),.dout(w_dff_B_hrRlyOSk0_2),.clk(gclk));
	jdff dff_B_ylrELTML5_1(.din(n680),.dout(w_dff_B_ylrELTML5_1),.clk(gclk));
	jdff dff_B_5WgVRk198_2(.din(n593),.dout(w_dff_B_5WgVRk198_2),.clk(gclk));
	jdff dff_B_9En3TXtx4_2(.din(w_dff_B_5WgVRk198_2),.dout(w_dff_B_9En3TXtx4_2),.clk(gclk));
	jdff dff_B_RC63I0fB5_2(.din(w_dff_B_9En3TXtx4_2),.dout(w_dff_B_RC63I0fB5_2),.clk(gclk));
	jdff dff_B_odALINGx2_2(.din(w_dff_B_RC63I0fB5_2),.dout(w_dff_B_odALINGx2_2),.clk(gclk));
	jdff dff_B_D1GKbF0c6_2(.din(w_dff_B_odALINGx2_2),.dout(w_dff_B_D1GKbF0c6_2),.clk(gclk));
	jdff dff_B_7sCYzbVI1_2(.din(w_dff_B_D1GKbF0c6_2),.dout(w_dff_B_7sCYzbVI1_2),.clk(gclk));
	jdff dff_B_si04EEu89_2(.din(w_dff_B_7sCYzbVI1_2),.dout(w_dff_B_si04EEu89_2),.clk(gclk));
	jdff dff_B_AiT3i1To3_2(.din(w_dff_B_si04EEu89_2),.dout(w_dff_B_AiT3i1To3_2),.clk(gclk));
	jdff dff_B_vMDhyFHi7_2(.din(w_dff_B_AiT3i1To3_2),.dout(w_dff_B_vMDhyFHi7_2),.clk(gclk));
	jdff dff_B_JU5pyfFM9_2(.din(w_dff_B_vMDhyFHi7_2),.dout(w_dff_B_JU5pyfFM9_2),.clk(gclk));
	jdff dff_B_ekup89cH3_2(.din(w_dff_B_JU5pyfFM9_2),.dout(w_dff_B_ekup89cH3_2),.clk(gclk));
	jdff dff_B_T57MD6st6_2(.din(w_dff_B_ekup89cH3_2),.dout(w_dff_B_T57MD6st6_2),.clk(gclk));
	jdff dff_B_HPEZ81tM1_2(.din(n616),.dout(w_dff_B_HPEZ81tM1_2),.clk(gclk));
	jdff dff_B_0hhdmz5A7_1(.din(n594),.dout(w_dff_B_0hhdmz5A7_1),.clk(gclk));
	jdff dff_B_GJ0sQQWE4_2(.din(n514),.dout(w_dff_B_GJ0sQQWE4_2),.clk(gclk));
	jdff dff_B_BMAXM5ca2_2(.din(w_dff_B_GJ0sQQWE4_2),.dout(w_dff_B_BMAXM5ca2_2),.clk(gclk));
	jdff dff_B_rgAEmIhb9_2(.din(w_dff_B_BMAXM5ca2_2),.dout(w_dff_B_rgAEmIhb9_2),.clk(gclk));
	jdff dff_B_z9jxILgS7_2(.din(w_dff_B_rgAEmIhb9_2),.dout(w_dff_B_z9jxILgS7_2),.clk(gclk));
	jdff dff_B_Yn1lVPN73_2(.din(w_dff_B_z9jxILgS7_2),.dout(w_dff_B_Yn1lVPN73_2),.clk(gclk));
	jdff dff_B_xELfyWBf3_2(.din(w_dff_B_Yn1lVPN73_2),.dout(w_dff_B_xELfyWBf3_2),.clk(gclk));
	jdff dff_B_7FJmKZb81_2(.din(w_dff_B_xELfyWBf3_2),.dout(w_dff_B_7FJmKZb81_2),.clk(gclk));
	jdff dff_B_PamvgK1M7_2(.din(w_dff_B_7FJmKZb81_2),.dout(w_dff_B_PamvgK1M7_2),.clk(gclk));
	jdff dff_B_aESPuByd0_2(.din(w_dff_B_PamvgK1M7_2),.dout(w_dff_B_aESPuByd0_2),.clk(gclk));
	jdff dff_B_dk64gEpf4_2(.din(n530),.dout(w_dff_B_dk64gEpf4_2),.clk(gclk));
	jdff dff_B_0jqNEiRK1_2(.din(w_dff_B_dk64gEpf4_2),.dout(w_dff_B_0jqNEiRK1_2),.clk(gclk));
	jdff dff_B_0cZVaPms4_1(.din(n515),.dout(w_dff_B_0cZVaPms4_1),.clk(gclk));
	jdff dff_B_J9N6v84s1_1(.din(w_dff_B_0cZVaPms4_1),.dout(w_dff_B_J9N6v84s1_1),.clk(gclk));
	jdff dff_B_ATxOrPEq5_1(.din(w_dff_B_J9N6v84s1_1),.dout(w_dff_B_ATxOrPEq5_1),.clk(gclk));
	jdff dff_B_Gp0urcmt4_1(.din(w_dff_B_ATxOrPEq5_1),.dout(w_dff_B_Gp0urcmt4_1),.clk(gclk));
	jdff dff_B_fKbhMkZJ9_1(.din(w_dff_B_Gp0urcmt4_1),.dout(w_dff_B_fKbhMkZJ9_1),.clk(gclk));
	jdff dff_B_7b9zcMbq5_1(.din(w_dff_B_fKbhMkZJ9_1),.dout(w_dff_B_7b9zcMbq5_1),.clk(gclk));
	jdff dff_B_qt3Ns1xz6_0(.din(n451),.dout(w_dff_B_qt3Ns1xz6_0),.clk(gclk));
	jdff dff_B_UK5oVL1A8_0(.din(w_dff_B_qt3Ns1xz6_0),.dout(w_dff_B_UK5oVL1A8_0),.clk(gclk));
	jdff dff_A_4mbiZx7q8_0(.dout(w_n450_0[0]),.din(w_dff_A_4mbiZx7q8_0),.clk(gclk));
	jdff dff_A_c7F6NGBy7_0(.dout(w_dff_A_4mbiZx7q8_0),.din(w_dff_A_c7F6NGBy7_0),.clk(gclk));
	jdff dff_A_PLejDV5i4_0(.dout(w_dff_A_c7F6NGBy7_0),.din(w_dff_A_PLejDV5i4_0),.clk(gclk));
	jdff dff_B_B7uYD8kd4_1(.din(n444),.dout(w_dff_B_B7uYD8kd4_1),.clk(gclk));
	jdff dff_A_xQ8IgenW8_0(.dout(w_n376_0[0]),.din(w_dff_A_xQ8IgenW8_0),.clk(gclk));
	jdff dff_A_gZ3zpvUA2_1(.dout(w_n376_0[1]),.din(w_dff_A_gZ3zpvUA2_1),.clk(gclk));
	jdff dff_A_xriyLzyx7_1(.dout(w_dff_A_gZ3zpvUA2_1),.din(w_dff_A_xriyLzyx7_1),.clk(gclk));
	jdff dff_A_oBtVO8qU7_1(.dout(w_n442_0[1]),.din(w_dff_A_oBtVO8qU7_1),.clk(gclk));
	jdff dff_A_wFrnZpCI9_1(.dout(w_dff_A_oBtVO8qU7_1),.din(w_dff_A_wFrnZpCI9_1),.clk(gclk));
	jdff dff_A_FU0O2HPX9_1(.dout(w_dff_A_wFrnZpCI9_1),.din(w_dff_A_FU0O2HPX9_1),.clk(gclk));
	jdff dff_A_PF47EiG56_1(.dout(w_dff_A_FU0O2HPX9_1),.din(w_dff_A_PF47EiG56_1),.clk(gclk));
	jdff dff_A_7OB2ckyA4_1(.dout(w_dff_A_PF47EiG56_1),.din(w_dff_A_7OB2ckyA4_1),.clk(gclk));
	jdff dff_A_BbMEquCd0_1(.dout(w_dff_A_7OB2ckyA4_1),.din(w_dff_A_BbMEquCd0_1),.clk(gclk));
	jdff dff_B_HeUhQdQa6_2(.din(n1682),.dout(w_dff_B_HeUhQdQa6_2),.clk(gclk));
	jdff dff_B_lVy3GB6O5_1(.din(n1680),.dout(w_dff_B_lVy3GB6O5_1),.clk(gclk));
	jdff dff_B_dQ3WJGGw7_2(.din(n1628),.dout(w_dff_B_dQ3WJGGw7_2),.clk(gclk));
	jdff dff_B_ldTcfqoU8_2(.din(w_dff_B_dQ3WJGGw7_2),.dout(w_dff_B_ldTcfqoU8_2),.clk(gclk));
	jdff dff_B_yZ6BmJrI4_2(.din(w_dff_B_ldTcfqoU8_2),.dout(w_dff_B_yZ6BmJrI4_2),.clk(gclk));
	jdff dff_B_xNLBdxsk3_2(.din(w_dff_B_yZ6BmJrI4_2),.dout(w_dff_B_xNLBdxsk3_2),.clk(gclk));
	jdff dff_B_qNahotcy8_2(.din(w_dff_B_xNLBdxsk3_2),.dout(w_dff_B_qNahotcy8_2),.clk(gclk));
	jdff dff_B_mOawhLJI5_2(.din(w_dff_B_qNahotcy8_2),.dout(w_dff_B_mOawhLJI5_2),.clk(gclk));
	jdff dff_B_TZUyEKTw9_2(.din(w_dff_B_mOawhLJI5_2),.dout(w_dff_B_TZUyEKTw9_2),.clk(gclk));
	jdff dff_B_wsvjI5u81_2(.din(w_dff_B_TZUyEKTw9_2),.dout(w_dff_B_wsvjI5u81_2),.clk(gclk));
	jdff dff_B_E6fgUefI1_2(.din(w_dff_B_wsvjI5u81_2),.dout(w_dff_B_E6fgUefI1_2),.clk(gclk));
	jdff dff_B_ktuDovzW2_2(.din(w_dff_B_E6fgUefI1_2),.dout(w_dff_B_ktuDovzW2_2),.clk(gclk));
	jdff dff_B_o1Wt4ZNl8_2(.din(w_dff_B_ktuDovzW2_2),.dout(w_dff_B_o1Wt4ZNl8_2),.clk(gclk));
	jdff dff_B_JehvfdXY1_2(.din(w_dff_B_o1Wt4ZNl8_2),.dout(w_dff_B_JehvfdXY1_2),.clk(gclk));
	jdff dff_B_pCYdOBkA6_2(.din(w_dff_B_JehvfdXY1_2),.dout(w_dff_B_pCYdOBkA6_2),.clk(gclk));
	jdff dff_B_aZ9m9OjY1_2(.din(w_dff_B_pCYdOBkA6_2),.dout(w_dff_B_aZ9m9OjY1_2),.clk(gclk));
	jdff dff_B_6GX5ZKiK9_2(.din(w_dff_B_aZ9m9OjY1_2),.dout(w_dff_B_6GX5ZKiK9_2),.clk(gclk));
	jdff dff_B_YS5Xjf8n2_2(.din(w_dff_B_6GX5ZKiK9_2),.dout(w_dff_B_YS5Xjf8n2_2),.clk(gclk));
	jdff dff_B_z459SVYz5_2(.din(w_dff_B_YS5Xjf8n2_2),.dout(w_dff_B_z459SVYz5_2),.clk(gclk));
	jdff dff_B_vZsySrL29_2(.din(w_dff_B_z459SVYz5_2),.dout(w_dff_B_vZsySrL29_2),.clk(gclk));
	jdff dff_B_Tp1rGKHW1_2(.din(w_dff_B_vZsySrL29_2),.dout(w_dff_B_Tp1rGKHW1_2),.clk(gclk));
	jdff dff_B_xxkAWJ7F4_2(.din(w_dff_B_Tp1rGKHW1_2),.dout(w_dff_B_xxkAWJ7F4_2),.clk(gclk));
	jdff dff_B_xHCqNPXw2_2(.din(w_dff_B_xxkAWJ7F4_2),.dout(w_dff_B_xHCqNPXw2_2),.clk(gclk));
	jdff dff_B_UE3jvtuC3_2(.din(w_dff_B_xHCqNPXw2_2),.dout(w_dff_B_UE3jvtuC3_2),.clk(gclk));
	jdff dff_B_EkKxvFEV9_2(.din(w_dff_B_UE3jvtuC3_2),.dout(w_dff_B_EkKxvFEV9_2),.clk(gclk));
	jdff dff_B_wIkZEgwB4_2(.din(w_dff_B_EkKxvFEV9_2),.dout(w_dff_B_wIkZEgwB4_2),.clk(gclk));
	jdff dff_B_cwMFckBl9_2(.din(w_dff_B_wIkZEgwB4_2),.dout(w_dff_B_cwMFckBl9_2),.clk(gclk));
	jdff dff_B_Lp9EeNir3_2(.din(w_dff_B_cwMFckBl9_2),.dout(w_dff_B_Lp9EeNir3_2),.clk(gclk));
	jdff dff_B_BddIGRgw3_2(.din(w_dff_B_Lp9EeNir3_2),.dout(w_dff_B_BddIGRgw3_2),.clk(gclk));
	jdff dff_B_JRcY3adb9_2(.din(w_dff_B_BddIGRgw3_2),.dout(w_dff_B_JRcY3adb9_2),.clk(gclk));
	jdff dff_B_Nmfldyfe3_2(.din(w_dff_B_JRcY3adb9_2),.dout(w_dff_B_Nmfldyfe3_2),.clk(gclk));
	jdff dff_B_4r3f1oaR5_2(.din(w_dff_B_Nmfldyfe3_2),.dout(w_dff_B_4r3f1oaR5_2),.clk(gclk));
	jdff dff_B_M1cAbZWF5_2(.din(w_dff_B_4r3f1oaR5_2),.dout(w_dff_B_M1cAbZWF5_2),.clk(gclk));
	jdff dff_B_bSafRusd4_2(.din(w_dff_B_M1cAbZWF5_2),.dout(w_dff_B_bSafRusd4_2),.clk(gclk));
	jdff dff_B_NTkWFEcR1_2(.din(w_dff_B_bSafRusd4_2),.dout(w_dff_B_NTkWFEcR1_2),.clk(gclk));
	jdff dff_B_mtWm4W9N8_2(.din(w_dff_B_NTkWFEcR1_2),.dout(w_dff_B_mtWm4W9N8_2),.clk(gclk));
	jdff dff_B_OBp95y760_2(.din(w_dff_B_mtWm4W9N8_2),.dout(w_dff_B_OBp95y760_2),.clk(gclk));
	jdff dff_B_yhdYSiQ66_2(.din(w_dff_B_OBp95y760_2),.dout(w_dff_B_yhdYSiQ66_2),.clk(gclk));
	jdff dff_B_zkNt7NFy7_2(.din(w_dff_B_yhdYSiQ66_2),.dout(w_dff_B_zkNt7NFy7_2),.clk(gclk));
	jdff dff_B_GxcqJDat1_2(.din(w_dff_B_zkNt7NFy7_2),.dout(w_dff_B_GxcqJDat1_2),.clk(gclk));
	jdff dff_B_ulZu1MnZ8_2(.din(w_dff_B_GxcqJDat1_2),.dout(w_dff_B_ulZu1MnZ8_2),.clk(gclk));
	jdff dff_B_GofV90ru9_2(.din(w_dff_B_ulZu1MnZ8_2),.dout(w_dff_B_GofV90ru9_2),.clk(gclk));
	jdff dff_B_Hk0erdO04_2(.din(w_dff_B_GofV90ru9_2),.dout(w_dff_B_Hk0erdO04_2),.clk(gclk));
	jdff dff_B_WQuHzJOg2_2(.din(w_dff_B_Hk0erdO04_2),.dout(w_dff_B_WQuHzJOg2_2),.clk(gclk));
	jdff dff_B_iLUMRCel7_2(.din(w_dff_B_WQuHzJOg2_2),.dout(w_dff_B_iLUMRCel7_2),.clk(gclk));
	jdff dff_B_Hp2dnVpw2_2(.din(w_dff_B_iLUMRCel7_2),.dout(w_dff_B_Hp2dnVpw2_2),.clk(gclk));
	jdff dff_B_6PCJZvOy1_2(.din(w_dff_B_Hp2dnVpw2_2),.dout(w_dff_B_6PCJZvOy1_2),.clk(gclk));
	jdff dff_B_vKAYiyDw8_2(.din(w_dff_B_6PCJZvOy1_2),.dout(w_dff_B_vKAYiyDw8_2),.clk(gclk));
	jdff dff_B_rkJpFx9l6_2(.din(w_dff_B_vKAYiyDw8_2),.dout(w_dff_B_rkJpFx9l6_2),.clk(gclk));
	jdff dff_B_FkJQaaKQ6_2(.din(w_dff_B_rkJpFx9l6_2),.dout(w_dff_B_FkJQaaKQ6_2),.clk(gclk));
	jdff dff_B_Zcxv3EB42_2(.din(w_dff_B_FkJQaaKQ6_2),.dout(w_dff_B_Zcxv3EB42_2),.clk(gclk));
	jdff dff_B_1uK7f00G7_1(.din(n1678),.dout(w_dff_B_1uK7f00G7_1),.clk(gclk));
	jdff dff_A_zzjBz9dq1_1(.dout(w_n1631_0[1]),.din(w_dff_A_zzjBz9dq1_1),.clk(gclk));
	jdff dff_B_8piwo4me2_1(.din(n1629),.dout(w_dff_B_8piwo4me2_1),.clk(gclk));
	jdff dff_B_GNtZnVvZ6_2(.din(n1571),.dout(w_dff_B_GNtZnVvZ6_2),.clk(gclk));
	jdff dff_B_BC58j5F35_2(.din(w_dff_B_GNtZnVvZ6_2),.dout(w_dff_B_BC58j5F35_2),.clk(gclk));
	jdff dff_B_tBUC1MJV0_2(.din(w_dff_B_BC58j5F35_2),.dout(w_dff_B_tBUC1MJV0_2),.clk(gclk));
	jdff dff_B_W3BlvzBt7_2(.din(w_dff_B_tBUC1MJV0_2),.dout(w_dff_B_W3BlvzBt7_2),.clk(gclk));
	jdff dff_B_fkrU0qgZ0_2(.din(w_dff_B_W3BlvzBt7_2),.dout(w_dff_B_fkrU0qgZ0_2),.clk(gclk));
	jdff dff_B_0IJ2MFpn8_2(.din(w_dff_B_fkrU0qgZ0_2),.dout(w_dff_B_0IJ2MFpn8_2),.clk(gclk));
	jdff dff_B_NtEEfmxq6_2(.din(w_dff_B_0IJ2MFpn8_2),.dout(w_dff_B_NtEEfmxq6_2),.clk(gclk));
	jdff dff_B_oDfhuqqw5_2(.din(w_dff_B_NtEEfmxq6_2),.dout(w_dff_B_oDfhuqqw5_2),.clk(gclk));
	jdff dff_B_O1v0LXH27_2(.din(w_dff_B_oDfhuqqw5_2),.dout(w_dff_B_O1v0LXH27_2),.clk(gclk));
	jdff dff_B_6hsAkfUT4_2(.din(w_dff_B_O1v0LXH27_2),.dout(w_dff_B_6hsAkfUT4_2),.clk(gclk));
	jdff dff_B_uKeW7jMU2_2(.din(w_dff_B_6hsAkfUT4_2),.dout(w_dff_B_uKeW7jMU2_2),.clk(gclk));
	jdff dff_B_telpEeq35_2(.din(w_dff_B_uKeW7jMU2_2),.dout(w_dff_B_telpEeq35_2),.clk(gclk));
	jdff dff_B_WjQ3XbRQ8_2(.din(w_dff_B_telpEeq35_2),.dout(w_dff_B_WjQ3XbRQ8_2),.clk(gclk));
	jdff dff_B_ljMxDcrC3_2(.din(w_dff_B_WjQ3XbRQ8_2),.dout(w_dff_B_ljMxDcrC3_2),.clk(gclk));
	jdff dff_B_LYdDuLik0_2(.din(w_dff_B_ljMxDcrC3_2),.dout(w_dff_B_LYdDuLik0_2),.clk(gclk));
	jdff dff_B_3bvJ530v8_2(.din(w_dff_B_LYdDuLik0_2),.dout(w_dff_B_3bvJ530v8_2),.clk(gclk));
	jdff dff_B_85rzEYy74_2(.din(w_dff_B_3bvJ530v8_2),.dout(w_dff_B_85rzEYy74_2),.clk(gclk));
	jdff dff_B_6bfBNvak7_2(.din(w_dff_B_85rzEYy74_2),.dout(w_dff_B_6bfBNvak7_2),.clk(gclk));
	jdff dff_B_nKxXDu9m9_2(.din(w_dff_B_6bfBNvak7_2),.dout(w_dff_B_nKxXDu9m9_2),.clk(gclk));
	jdff dff_B_ZK55cj8A1_2(.din(w_dff_B_nKxXDu9m9_2),.dout(w_dff_B_ZK55cj8A1_2),.clk(gclk));
	jdff dff_B_v7Jz1dQl8_2(.din(w_dff_B_ZK55cj8A1_2),.dout(w_dff_B_v7Jz1dQl8_2),.clk(gclk));
	jdff dff_B_GSQbuvq19_2(.din(w_dff_B_v7Jz1dQl8_2),.dout(w_dff_B_GSQbuvq19_2),.clk(gclk));
	jdff dff_B_BHwTPlm92_2(.din(w_dff_B_GSQbuvq19_2),.dout(w_dff_B_BHwTPlm92_2),.clk(gclk));
	jdff dff_B_0O5ul9Ub9_2(.din(w_dff_B_BHwTPlm92_2),.dout(w_dff_B_0O5ul9Ub9_2),.clk(gclk));
	jdff dff_B_T7aQKPFW2_2(.din(w_dff_B_0O5ul9Ub9_2),.dout(w_dff_B_T7aQKPFW2_2),.clk(gclk));
	jdff dff_B_pn3FhFV56_2(.din(w_dff_B_T7aQKPFW2_2),.dout(w_dff_B_pn3FhFV56_2),.clk(gclk));
	jdff dff_B_mWeyXP3g8_2(.din(w_dff_B_pn3FhFV56_2),.dout(w_dff_B_mWeyXP3g8_2),.clk(gclk));
	jdff dff_B_wuBXv44K0_2(.din(w_dff_B_mWeyXP3g8_2),.dout(w_dff_B_wuBXv44K0_2),.clk(gclk));
	jdff dff_B_RyPlMtWv9_2(.din(w_dff_B_wuBXv44K0_2),.dout(w_dff_B_RyPlMtWv9_2),.clk(gclk));
	jdff dff_B_euzJQrrl4_2(.din(w_dff_B_RyPlMtWv9_2),.dout(w_dff_B_euzJQrrl4_2),.clk(gclk));
	jdff dff_B_97zkkpKf2_2(.din(w_dff_B_euzJQrrl4_2),.dout(w_dff_B_97zkkpKf2_2),.clk(gclk));
	jdff dff_B_gA1ogjDf1_2(.din(w_dff_B_97zkkpKf2_2),.dout(w_dff_B_gA1ogjDf1_2),.clk(gclk));
	jdff dff_B_ZN5G2luJ2_2(.din(w_dff_B_gA1ogjDf1_2),.dout(w_dff_B_ZN5G2luJ2_2),.clk(gclk));
	jdff dff_B_sa8PHzss0_2(.din(w_dff_B_ZN5G2luJ2_2),.dout(w_dff_B_sa8PHzss0_2),.clk(gclk));
	jdff dff_B_1OPCSsHP9_2(.din(w_dff_B_sa8PHzss0_2),.dout(w_dff_B_1OPCSsHP9_2),.clk(gclk));
	jdff dff_B_HAPxhBxl3_2(.din(w_dff_B_1OPCSsHP9_2),.dout(w_dff_B_HAPxhBxl3_2),.clk(gclk));
	jdff dff_B_DKbrqyWa3_2(.din(w_dff_B_HAPxhBxl3_2),.dout(w_dff_B_DKbrqyWa3_2),.clk(gclk));
	jdff dff_B_9qOsFu9L6_2(.din(w_dff_B_DKbrqyWa3_2),.dout(w_dff_B_9qOsFu9L6_2),.clk(gclk));
	jdff dff_B_SKOBbt7E1_2(.din(w_dff_B_9qOsFu9L6_2),.dout(w_dff_B_SKOBbt7E1_2),.clk(gclk));
	jdff dff_B_Ylbd4SZn3_2(.din(w_dff_B_SKOBbt7E1_2),.dout(w_dff_B_Ylbd4SZn3_2),.clk(gclk));
	jdff dff_B_XCDLpu8W2_2(.din(w_dff_B_Ylbd4SZn3_2),.dout(w_dff_B_XCDLpu8W2_2),.clk(gclk));
	jdff dff_B_yCq2Ccq29_2(.din(w_dff_B_XCDLpu8W2_2),.dout(w_dff_B_yCq2Ccq29_2),.clk(gclk));
	jdff dff_B_wG1Npweu9_2(.din(w_dff_B_yCq2Ccq29_2),.dout(w_dff_B_wG1Npweu9_2),.clk(gclk));
	jdff dff_B_Noqgof8s2_2(.din(n1574),.dout(w_dff_B_Noqgof8s2_2),.clk(gclk));
	jdff dff_B_tX56hz7o5_1(.din(n1572),.dout(w_dff_B_tX56hz7o5_1),.clk(gclk));
	jdff dff_B_9FCnLDfC0_2(.din(n1507),.dout(w_dff_B_9FCnLDfC0_2),.clk(gclk));
	jdff dff_B_QILD84OU0_2(.din(w_dff_B_9FCnLDfC0_2),.dout(w_dff_B_QILD84OU0_2),.clk(gclk));
	jdff dff_B_SlzcR0VO9_2(.din(w_dff_B_QILD84OU0_2),.dout(w_dff_B_SlzcR0VO9_2),.clk(gclk));
	jdff dff_B_UBgjGxke7_2(.din(w_dff_B_SlzcR0VO9_2),.dout(w_dff_B_UBgjGxke7_2),.clk(gclk));
	jdff dff_B_0cXQYiqv7_2(.din(w_dff_B_UBgjGxke7_2),.dout(w_dff_B_0cXQYiqv7_2),.clk(gclk));
	jdff dff_B_DRzKXMe08_2(.din(w_dff_B_0cXQYiqv7_2),.dout(w_dff_B_DRzKXMe08_2),.clk(gclk));
	jdff dff_B_txBI72Yv5_2(.din(w_dff_B_DRzKXMe08_2),.dout(w_dff_B_txBI72Yv5_2),.clk(gclk));
	jdff dff_B_GtA5nQ8y6_2(.din(w_dff_B_txBI72Yv5_2),.dout(w_dff_B_GtA5nQ8y6_2),.clk(gclk));
	jdff dff_B_21a9CdXg4_2(.din(w_dff_B_GtA5nQ8y6_2),.dout(w_dff_B_21a9CdXg4_2),.clk(gclk));
	jdff dff_B_b3WqfLXW9_2(.din(w_dff_B_21a9CdXg4_2),.dout(w_dff_B_b3WqfLXW9_2),.clk(gclk));
	jdff dff_B_0R5jye7Y0_2(.din(w_dff_B_b3WqfLXW9_2),.dout(w_dff_B_0R5jye7Y0_2),.clk(gclk));
	jdff dff_B_qxEdKKvB9_2(.din(w_dff_B_0R5jye7Y0_2),.dout(w_dff_B_qxEdKKvB9_2),.clk(gclk));
	jdff dff_B_8FHL79Kr7_2(.din(w_dff_B_qxEdKKvB9_2),.dout(w_dff_B_8FHL79Kr7_2),.clk(gclk));
	jdff dff_B_lKwL8on02_2(.din(w_dff_B_8FHL79Kr7_2),.dout(w_dff_B_lKwL8on02_2),.clk(gclk));
	jdff dff_B_T6cuERnm2_2(.din(w_dff_B_lKwL8on02_2),.dout(w_dff_B_T6cuERnm2_2),.clk(gclk));
	jdff dff_B_hbNV5vVv1_2(.din(w_dff_B_T6cuERnm2_2),.dout(w_dff_B_hbNV5vVv1_2),.clk(gclk));
	jdff dff_B_V1usOsl04_2(.din(w_dff_B_hbNV5vVv1_2),.dout(w_dff_B_V1usOsl04_2),.clk(gclk));
	jdff dff_B_YNtdHl5H2_2(.din(w_dff_B_V1usOsl04_2),.dout(w_dff_B_YNtdHl5H2_2),.clk(gclk));
	jdff dff_B_41oDOv7S4_2(.din(w_dff_B_YNtdHl5H2_2),.dout(w_dff_B_41oDOv7S4_2),.clk(gclk));
	jdff dff_B_Av24EUB60_2(.din(w_dff_B_41oDOv7S4_2),.dout(w_dff_B_Av24EUB60_2),.clk(gclk));
	jdff dff_B_etygBPsg4_2(.din(w_dff_B_Av24EUB60_2),.dout(w_dff_B_etygBPsg4_2),.clk(gclk));
	jdff dff_B_37pUb7NC7_2(.din(w_dff_B_etygBPsg4_2),.dout(w_dff_B_37pUb7NC7_2),.clk(gclk));
	jdff dff_B_O76lKCOF6_2(.din(w_dff_B_37pUb7NC7_2),.dout(w_dff_B_O76lKCOF6_2),.clk(gclk));
	jdff dff_B_nORxJQ7s2_2(.din(w_dff_B_O76lKCOF6_2),.dout(w_dff_B_nORxJQ7s2_2),.clk(gclk));
	jdff dff_B_VzZVCbWW8_2(.din(w_dff_B_nORxJQ7s2_2),.dout(w_dff_B_VzZVCbWW8_2),.clk(gclk));
	jdff dff_B_mZa67PnZ2_2(.din(w_dff_B_VzZVCbWW8_2),.dout(w_dff_B_mZa67PnZ2_2),.clk(gclk));
	jdff dff_B_X6RWB88F6_2(.din(w_dff_B_mZa67PnZ2_2),.dout(w_dff_B_X6RWB88F6_2),.clk(gclk));
	jdff dff_B_CwGiKdgi9_2(.din(w_dff_B_X6RWB88F6_2),.dout(w_dff_B_CwGiKdgi9_2),.clk(gclk));
	jdff dff_B_4itIrE3x9_2(.din(w_dff_B_CwGiKdgi9_2),.dout(w_dff_B_4itIrE3x9_2),.clk(gclk));
	jdff dff_B_dTG4LYCM5_2(.din(w_dff_B_4itIrE3x9_2),.dout(w_dff_B_dTG4LYCM5_2),.clk(gclk));
	jdff dff_B_CuIpjjBq1_2(.din(w_dff_B_dTG4LYCM5_2),.dout(w_dff_B_CuIpjjBq1_2),.clk(gclk));
	jdff dff_B_jy9S97pJ4_2(.din(w_dff_B_CuIpjjBq1_2),.dout(w_dff_B_jy9S97pJ4_2),.clk(gclk));
	jdff dff_B_OuLfGXr64_2(.din(w_dff_B_jy9S97pJ4_2),.dout(w_dff_B_OuLfGXr64_2),.clk(gclk));
	jdff dff_B_vnVYfSRN1_2(.din(w_dff_B_OuLfGXr64_2),.dout(w_dff_B_vnVYfSRN1_2),.clk(gclk));
	jdff dff_B_0nkKLhek2_2(.din(w_dff_B_vnVYfSRN1_2),.dout(w_dff_B_0nkKLhek2_2),.clk(gclk));
	jdff dff_B_JKtBWnzS4_2(.din(w_dff_B_0nkKLhek2_2),.dout(w_dff_B_JKtBWnzS4_2),.clk(gclk));
	jdff dff_B_fkcq9az63_2(.din(w_dff_B_JKtBWnzS4_2),.dout(w_dff_B_fkcq9az63_2),.clk(gclk));
	jdff dff_B_kDxvW6Z86_2(.din(w_dff_B_fkcq9az63_2),.dout(w_dff_B_kDxvW6Z86_2),.clk(gclk));
	jdff dff_B_k7ju0uw85_2(.din(w_dff_B_kDxvW6Z86_2),.dout(w_dff_B_k7ju0uw85_2),.clk(gclk));
	jdff dff_B_6NaOW2oA3_1(.din(n1508),.dout(w_dff_B_6NaOW2oA3_1),.clk(gclk));
	jdff dff_B_nF1gvEjr2_2(.din(n1436),.dout(w_dff_B_nF1gvEjr2_2),.clk(gclk));
	jdff dff_B_CsWCo8Xl3_2(.din(w_dff_B_nF1gvEjr2_2),.dout(w_dff_B_CsWCo8Xl3_2),.clk(gclk));
	jdff dff_B_aR9Py4x91_2(.din(w_dff_B_CsWCo8Xl3_2),.dout(w_dff_B_aR9Py4x91_2),.clk(gclk));
	jdff dff_B_ZkldLel05_2(.din(w_dff_B_aR9Py4x91_2),.dout(w_dff_B_ZkldLel05_2),.clk(gclk));
	jdff dff_B_WmGppmAH4_2(.din(w_dff_B_ZkldLel05_2),.dout(w_dff_B_WmGppmAH4_2),.clk(gclk));
	jdff dff_B_83D1O2ez9_2(.din(w_dff_B_WmGppmAH4_2),.dout(w_dff_B_83D1O2ez9_2),.clk(gclk));
	jdff dff_B_V0QG3D9p3_2(.din(w_dff_B_83D1O2ez9_2),.dout(w_dff_B_V0QG3D9p3_2),.clk(gclk));
	jdff dff_B_d2eu5nKd1_2(.din(w_dff_B_V0QG3D9p3_2),.dout(w_dff_B_d2eu5nKd1_2),.clk(gclk));
	jdff dff_B_veuu8M036_2(.din(w_dff_B_d2eu5nKd1_2),.dout(w_dff_B_veuu8M036_2),.clk(gclk));
	jdff dff_B_yRRLMSK59_2(.din(w_dff_B_veuu8M036_2),.dout(w_dff_B_yRRLMSK59_2),.clk(gclk));
	jdff dff_B_8fR9fykw8_2(.din(w_dff_B_yRRLMSK59_2),.dout(w_dff_B_8fR9fykw8_2),.clk(gclk));
	jdff dff_B_epPw27jC9_2(.din(w_dff_B_8fR9fykw8_2),.dout(w_dff_B_epPw27jC9_2),.clk(gclk));
	jdff dff_B_l0jY552I6_2(.din(w_dff_B_epPw27jC9_2),.dout(w_dff_B_l0jY552I6_2),.clk(gclk));
	jdff dff_B_ulOYps4L6_2(.din(w_dff_B_l0jY552I6_2),.dout(w_dff_B_ulOYps4L6_2),.clk(gclk));
	jdff dff_B_RKaAF2Bz0_2(.din(w_dff_B_ulOYps4L6_2),.dout(w_dff_B_RKaAF2Bz0_2),.clk(gclk));
	jdff dff_B_hixJMzbZ9_2(.din(w_dff_B_RKaAF2Bz0_2),.dout(w_dff_B_hixJMzbZ9_2),.clk(gclk));
	jdff dff_B_SqpKesEp6_2(.din(w_dff_B_hixJMzbZ9_2),.dout(w_dff_B_SqpKesEp6_2),.clk(gclk));
	jdff dff_B_eVOb76Xz6_2(.din(w_dff_B_SqpKesEp6_2),.dout(w_dff_B_eVOb76Xz6_2),.clk(gclk));
	jdff dff_B_XCkHZtnd5_2(.din(w_dff_B_eVOb76Xz6_2),.dout(w_dff_B_XCkHZtnd5_2),.clk(gclk));
	jdff dff_B_TdGdLDEh4_2(.din(w_dff_B_XCkHZtnd5_2),.dout(w_dff_B_TdGdLDEh4_2),.clk(gclk));
	jdff dff_B_wyMWoNYX2_2(.din(w_dff_B_TdGdLDEh4_2),.dout(w_dff_B_wyMWoNYX2_2),.clk(gclk));
	jdff dff_B_mGxCDdZ50_2(.din(w_dff_B_wyMWoNYX2_2),.dout(w_dff_B_mGxCDdZ50_2),.clk(gclk));
	jdff dff_B_YEuEAVZI6_2(.din(w_dff_B_mGxCDdZ50_2),.dout(w_dff_B_YEuEAVZI6_2),.clk(gclk));
	jdff dff_B_WFzf4FDq0_2(.din(w_dff_B_YEuEAVZI6_2),.dout(w_dff_B_WFzf4FDq0_2),.clk(gclk));
	jdff dff_B_iRgy355T2_2(.din(w_dff_B_WFzf4FDq0_2),.dout(w_dff_B_iRgy355T2_2),.clk(gclk));
	jdff dff_B_dtcmYRqc6_2(.din(w_dff_B_iRgy355T2_2),.dout(w_dff_B_dtcmYRqc6_2),.clk(gclk));
	jdff dff_B_MOJ18p1E3_2(.din(w_dff_B_dtcmYRqc6_2),.dout(w_dff_B_MOJ18p1E3_2),.clk(gclk));
	jdff dff_B_KOtE8ltQ8_2(.din(w_dff_B_MOJ18p1E3_2),.dout(w_dff_B_KOtE8ltQ8_2),.clk(gclk));
	jdff dff_B_ghuSZZYC5_2(.din(w_dff_B_KOtE8ltQ8_2),.dout(w_dff_B_ghuSZZYC5_2),.clk(gclk));
	jdff dff_B_npqSoASv5_2(.din(w_dff_B_ghuSZZYC5_2),.dout(w_dff_B_npqSoASv5_2),.clk(gclk));
	jdff dff_B_jBDlSCiV5_2(.din(w_dff_B_npqSoASv5_2),.dout(w_dff_B_jBDlSCiV5_2),.clk(gclk));
	jdff dff_B_A3VBZ0HC6_2(.din(w_dff_B_jBDlSCiV5_2),.dout(w_dff_B_A3VBZ0HC6_2),.clk(gclk));
	jdff dff_B_t3u4FL7p9_2(.din(w_dff_B_A3VBZ0HC6_2),.dout(w_dff_B_t3u4FL7p9_2),.clk(gclk));
	jdff dff_B_TQfQi3H54_2(.din(w_dff_B_t3u4FL7p9_2),.dout(w_dff_B_TQfQi3H54_2),.clk(gclk));
	jdff dff_B_CFl6tAIv5_2(.din(w_dff_B_TQfQi3H54_2),.dout(w_dff_B_CFl6tAIv5_2),.clk(gclk));
	jdff dff_B_apora1Ov2_2(.din(w_dff_B_CFl6tAIv5_2),.dout(w_dff_B_apora1Ov2_2),.clk(gclk));
	jdff dff_B_Jmxx0iWk6_2(.din(n1475),.dout(w_dff_B_Jmxx0iWk6_2),.clk(gclk));
	jdff dff_B_0zbkiSiI3_1(.din(n1437),.dout(w_dff_B_0zbkiSiI3_1),.clk(gclk));
	jdff dff_B_ULwV9H8K6_2(.din(n1358),.dout(w_dff_B_ULwV9H8K6_2),.clk(gclk));
	jdff dff_B_xLGopkgf0_2(.din(w_dff_B_ULwV9H8K6_2),.dout(w_dff_B_xLGopkgf0_2),.clk(gclk));
	jdff dff_B_kNmXhQ9E1_2(.din(w_dff_B_xLGopkgf0_2),.dout(w_dff_B_kNmXhQ9E1_2),.clk(gclk));
	jdff dff_B_x645mFm42_2(.din(w_dff_B_kNmXhQ9E1_2),.dout(w_dff_B_x645mFm42_2),.clk(gclk));
	jdff dff_B_X4QKCLC96_2(.din(w_dff_B_x645mFm42_2),.dout(w_dff_B_X4QKCLC96_2),.clk(gclk));
	jdff dff_B_fz3qGhTS1_2(.din(w_dff_B_X4QKCLC96_2),.dout(w_dff_B_fz3qGhTS1_2),.clk(gclk));
	jdff dff_B_8zP02RlI7_2(.din(w_dff_B_fz3qGhTS1_2),.dout(w_dff_B_8zP02RlI7_2),.clk(gclk));
	jdff dff_B_logvZ88f8_2(.din(w_dff_B_8zP02RlI7_2),.dout(w_dff_B_logvZ88f8_2),.clk(gclk));
	jdff dff_B_Z2Id0T8t7_2(.din(w_dff_B_logvZ88f8_2),.dout(w_dff_B_Z2Id0T8t7_2),.clk(gclk));
	jdff dff_B_4V1y7eKD5_2(.din(w_dff_B_Z2Id0T8t7_2),.dout(w_dff_B_4V1y7eKD5_2),.clk(gclk));
	jdff dff_B_Ml2hwIKz8_2(.din(w_dff_B_4V1y7eKD5_2),.dout(w_dff_B_Ml2hwIKz8_2),.clk(gclk));
	jdff dff_B_zCSbThxH9_2(.din(w_dff_B_Ml2hwIKz8_2),.dout(w_dff_B_zCSbThxH9_2),.clk(gclk));
	jdff dff_B_jGWAjlyS7_2(.din(w_dff_B_zCSbThxH9_2),.dout(w_dff_B_jGWAjlyS7_2),.clk(gclk));
	jdff dff_B_zFz9ZT6K1_2(.din(w_dff_B_jGWAjlyS7_2),.dout(w_dff_B_zFz9ZT6K1_2),.clk(gclk));
	jdff dff_B_yuzxBeyp6_2(.din(w_dff_B_zFz9ZT6K1_2),.dout(w_dff_B_yuzxBeyp6_2),.clk(gclk));
	jdff dff_B_FawMs8CI6_2(.din(w_dff_B_yuzxBeyp6_2),.dout(w_dff_B_FawMs8CI6_2),.clk(gclk));
	jdff dff_B_4nMrm7rk6_2(.din(w_dff_B_FawMs8CI6_2),.dout(w_dff_B_4nMrm7rk6_2),.clk(gclk));
	jdff dff_B_O4o09TlU8_2(.din(w_dff_B_4nMrm7rk6_2),.dout(w_dff_B_O4o09TlU8_2),.clk(gclk));
	jdff dff_B_L130e9Lv0_2(.din(w_dff_B_O4o09TlU8_2),.dout(w_dff_B_L130e9Lv0_2),.clk(gclk));
	jdff dff_B_AgqRvNee2_2(.din(w_dff_B_L130e9Lv0_2),.dout(w_dff_B_AgqRvNee2_2),.clk(gclk));
	jdff dff_B_9gYvM1Gb5_2(.din(w_dff_B_AgqRvNee2_2),.dout(w_dff_B_9gYvM1Gb5_2),.clk(gclk));
	jdff dff_B_Gz9EnSyV9_2(.din(w_dff_B_9gYvM1Gb5_2),.dout(w_dff_B_Gz9EnSyV9_2),.clk(gclk));
	jdff dff_B_F2YcDJsJ5_2(.din(w_dff_B_Gz9EnSyV9_2),.dout(w_dff_B_F2YcDJsJ5_2),.clk(gclk));
	jdff dff_B_6Ous1wom8_2(.din(w_dff_B_F2YcDJsJ5_2),.dout(w_dff_B_6Ous1wom8_2),.clk(gclk));
	jdff dff_B_QMsrHuJN5_2(.din(w_dff_B_6Ous1wom8_2),.dout(w_dff_B_QMsrHuJN5_2),.clk(gclk));
	jdff dff_B_QXh3l63O4_2(.din(w_dff_B_QMsrHuJN5_2),.dout(w_dff_B_QXh3l63O4_2),.clk(gclk));
	jdff dff_B_V5mVErpJ3_2(.din(w_dff_B_QXh3l63O4_2),.dout(w_dff_B_V5mVErpJ3_2),.clk(gclk));
	jdff dff_B_Q9VBhwBD2_2(.din(w_dff_B_V5mVErpJ3_2),.dout(w_dff_B_Q9VBhwBD2_2),.clk(gclk));
	jdff dff_B_uXcl4qyC6_2(.din(w_dff_B_Q9VBhwBD2_2),.dout(w_dff_B_uXcl4qyC6_2),.clk(gclk));
	jdff dff_B_iGM9JZXL6_2(.din(w_dff_B_uXcl4qyC6_2),.dout(w_dff_B_iGM9JZXL6_2),.clk(gclk));
	jdff dff_B_NfLRQCCH1_2(.din(w_dff_B_iGM9JZXL6_2),.dout(w_dff_B_NfLRQCCH1_2),.clk(gclk));
	jdff dff_B_K4Osp7Zy8_2(.din(w_dff_B_NfLRQCCH1_2),.dout(w_dff_B_K4Osp7Zy8_2),.clk(gclk));
	jdff dff_B_ZKhslv1z7_2(.din(w_dff_B_K4Osp7Zy8_2),.dout(w_dff_B_ZKhslv1z7_2),.clk(gclk));
	jdff dff_B_wETVknfo3_2(.din(n1397),.dout(w_dff_B_wETVknfo3_2),.clk(gclk));
	jdff dff_B_CE7lS43i5_1(.din(n1359),.dout(w_dff_B_CE7lS43i5_1),.clk(gclk));
	jdff dff_B_oSkge1wz6_2(.din(n1273),.dout(w_dff_B_oSkge1wz6_2),.clk(gclk));
	jdff dff_B_OZNWplzX5_2(.din(w_dff_B_oSkge1wz6_2),.dout(w_dff_B_OZNWplzX5_2),.clk(gclk));
	jdff dff_B_i2w7qUCi6_2(.din(w_dff_B_OZNWplzX5_2),.dout(w_dff_B_i2w7qUCi6_2),.clk(gclk));
	jdff dff_B_WBafffGL1_2(.din(w_dff_B_i2w7qUCi6_2),.dout(w_dff_B_WBafffGL1_2),.clk(gclk));
	jdff dff_B_U9IasaPX0_2(.din(w_dff_B_WBafffGL1_2),.dout(w_dff_B_U9IasaPX0_2),.clk(gclk));
	jdff dff_B_7oxxEOqn1_2(.din(w_dff_B_U9IasaPX0_2),.dout(w_dff_B_7oxxEOqn1_2),.clk(gclk));
	jdff dff_B_hOVdS20Q4_2(.din(w_dff_B_7oxxEOqn1_2),.dout(w_dff_B_hOVdS20Q4_2),.clk(gclk));
	jdff dff_B_jzhZiZJb8_2(.din(w_dff_B_hOVdS20Q4_2),.dout(w_dff_B_jzhZiZJb8_2),.clk(gclk));
	jdff dff_B_jTONLOKF2_2(.din(w_dff_B_jzhZiZJb8_2),.dout(w_dff_B_jTONLOKF2_2),.clk(gclk));
	jdff dff_B_eAELwhp47_2(.din(w_dff_B_jTONLOKF2_2),.dout(w_dff_B_eAELwhp47_2),.clk(gclk));
	jdff dff_B_FB2ZC8Lh0_2(.din(w_dff_B_eAELwhp47_2),.dout(w_dff_B_FB2ZC8Lh0_2),.clk(gclk));
	jdff dff_B_hYGyFPaf4_2(.din(w_dff_B_FB2ZC8Lh0_2),.dout(w_dff_B_hYGyFPaf4_2),.clk(gclk));
	jdff dff_B_Ud8xlKNQ2_2(.din(w_dff_B_hYGyFPaf4_2),.dout(w_dff_B_Ud8xlKNQ2_2),.clk(gclk));
	jdff dff_B_ILOug0Gv0_2(.din(w_dff_B_Ud8xlKNQ2_2),.dout(w_dff_B_ILOug0Gv0_2),.clk(gclk));
	jdff dff_B_o7fHHtYa3_2(.din(w_dff_B_ILOug0Gv0_2),.dout(w_dff_B_o7fHHtYa3_2),.clk(gclk));
	jdff dff_B_e3JSNZto0_2(.din(w_dff_B_o7fHHtYa3_2),.dout(w_dff_B_e3JSNZto0_2),.clk(gclk));
	jdff dff_B_XkPs0ArA9_2(.din(w_dff_B_e3JSNZto0_2),.dout(w_dff_B_XkPs0ArA9_2),.clk(gclk));
	jdff dff_B_HZ29W4hh4_2(.din(w_dff_B_XkPs0ArA9_2),.dout(w_dff_B_HZ29W4hh4_2),.clk(gclk));
	jdff dff_B_ohXKGGyO3_2(.din(w_dff_B_HZ29W4hh4_2),.dout(w_dff_B_ohXKGGyO3_2),.clk(gclk));
	jdff dff_B_kHmhPEwo2_2(.din(w_dff_B_ohXKGGyO3_2),.dout(w_dff_B_kHmhPEwo2_2),.clk(gclk));
	jdff dff_B_P6WKDGfg9_2(.din(w_dff_B_kHmhPEwo2_2),.dout(w_dff_B_P6WKDGfg9_2),.clk(gclk));
	jdff dff_B_j2uuOPfn3_2(.din(w_dff_B_P6WKDGfg9_2),.dout(w_dff_B_j2uuOPfn3_2),.clk(gclk));
	jdff dff_B_MdQBCLTg5_2(.din(w_dff_B_j2uuOPfn3_2),.dout(w_dff_B_MdQBCLTg5_2),.clk(gclk));
	jdff dff_B_zthjBxNu4_2(.din(w_dff_B_MdQBCLTg5_2),.dout(w_dff_B_zthjBxNu4_2),.clk(gclk));
	jdff dff_B_nWdVCvXM9_2(.din(w_dff_B_zthjBxNu4_2),.dout(w_dff_B_nWdVCvXM9_2),.clk(gclk));
	jdff dff_B_2teXDn471_2(.din(w_dff_B_nWdVCvXM9_2),.dout(w_dff_B_2teXDn471_2),.clk(gclk));
	jdff dff_B_YVTNBWn52_2(.din(w_dff_B_2teXDn471_2),.dout(w_dff_B_YVTNBWn52_2),.clk(gclk));
	jdff dff_B_FOsclKzN3_2(.din(w_dff_B_YVTNBWn52_2),.dout(w_dff_B_FOsclKzN3_2),.clk(gclk));
	jdff dff_B_YSkeVL2d6_2(.din(w_dff_B_FOsclKzN3_2),.dout(w_dff_B_YSkeVL2d6_2),.clk(gclk));
	jdff dff_B_w0rM8Gjh0_2(.din(w_dff_B_YSkeVL2d6_2),.dout(w_dff_B_w0rM8Gjh0_2),.clk(gclk));
	jdff dff_B_rTBOuZFw4_2(.din(n1312),.dout(w_dff_B_rTBOuZFw4_2),.clk(gclk));
	jdff dff_B_2pzKa2wU6_1(.din(n1274),.dout(w_dff_B_2pzKa2wU6_1),.clk(gclk));
	jdff dff_B_ZUlZ66mh1_2(.din(n1183),.dout(w_dff_B_ZUlZ66mh1_2),.clk(gclk));
	jdff dff_B_X2hyDXX12_2(.din(w_dff_B_ZUlZ66mh1_2),.dout(w_dff_B_X2hyDXX12_2),.clk(gclk));
	jdff dff_B_lP4BmWsy2_2(.din(w_dff_B_X2hyDXX12_2),.dout(w_dff_B_lP4BmWsy2_2),.clk(gclk));
	jdff dff_B_gDpP7nfq6_2(.din(w_dff_B_lP4BmWsy2_2),.dout(w_dff_B_gDpP7nfq6_2),.clk(gclk));
	jdff dff_B_J5CRVO5y2_2(.din(w_dff_B_gDpP7nfq6_2),.dout(w_dff_B_J5CRVO5y2_2),.clk(gclk));
	jdff dff_B_glqvyk642_2(.din(w_dff_B_J5CRVO5y2_2),.dout(w_dff_B_glqvyk642_2),.clk(gclk));
	jdff dff_B_SxCFBQLJ0_2(.din(w_dff_B_glqvyk642_2),.dout(w_dff_B_SxCFBQLJ0_2),.clk(gclk));
	jdff dff_B_Yy3lo1wa7_2(.din(w_dff_B_SxCFBQLJ0_2),.dout(w_dff_B_Yy3lo1wa7_2),.clk(gclk));
	jdff dff_B_yV4xYn2e2_2(.din(w_dff_B_Yy3lo1wa7_2),.dout(w_dff_B_yV4xYn2e2_2),.clk(gclk));
	jdff dff_B_n3kDKDkW6_2(.din(w_dff_B_yV4xYn2e2_2),.dout(w_dff_B_n3kDKDkW6_2),.clk(gclk));
	jdff dff_B_OugAvdJv6_2(.din(w_dff_B_n3kDKDkW6_2),.dout(w_dff_B_OugAvdJv6_2),.clk(gclk));
	jdff dff_B_WwZaeYDE7_2(.din(w_dff_B_OugAvdJv6_2),.dout(w_dff_B_WwZaeYDE7_2),.clk(gclk));
	jdff dff_B_sSENcVUd2_2(.din(w_dff_B_WwZaeYDE7_2),.dout(w_dff_B_sSENcVUd2_2),.clk(gclk));
	jdff dff_B_drzbCvJF2_2(.din(w_dff_B_sSENcVUd2_2),.dout(w_dff_B_drzbCvJF2_2),.clk(gclk));
	jdff dff_B_6pnHQkNz0_2(.din(w_dff_B_drzbCvJF2_2),.dout(w_dff_B_6pnHQkNz0_2),.clk(gclk));
	jdff dff_B_GHGRV3z03_2(.din(w_dff_B_6pnHQkNz0_2),.dout(w_dff_B_GHGRV3z03_2),.clk(gclk));
	jdff dff_B_kx2W5BoE2_2(.din(w_dff_B_GHGRV3z03_2),.dout(w_dff_B_kx2W5BoE2_2),.clk(gclk));
	jdff dff_B_fCBQU8gt7_2(.din(w_dff_B_kx2W5BoE2_2),.dout(w_dff_B_fCBQU8gt7_2),.clk(gclk));
	jdff dff_B_Kwpo1Oyz0_2(.din(w_dff_B_fCBQU8gt7_2),.dout(w_dff_B_Kwpo1Oyz0_2),.clk(gclk));
	jdff dff_B_voDm8Txc9_2(.din(w_dff_B_Kwpo1Oyz0_2),.dout(w_dff_B_voDm8Txc9_2),.clk(gclk));
	jdff dff_B_GhN36jN26_2(.din(w_dff_B_voDm8Txc9_2),.dout(w_dff_B_GhN36jN26_2),.clk(gclk));
	jdff dff_B_jxzTPCt39_2(.din(w_dff_B_GhN36jN26_2),.dout(w_dff_B_jxzTPCt39_2),.clk(gclk));
	jdff dff_B_WX55OYxl8_2(.din(w_dff_B_jxzTPCt39_2),.dout(w_dff_B_WX55OYxl8_2),.clk(gclk));
	jdff dff_B_jQb6Iy5f1_2(.din(w_dff_B_WX55OYxl8_2),.dout(w_dff_B_jQb6Iy5f1_2),.clk(gclk));
	jdff dff_B_MUmWnAOJ1_2(.din(w_dff_B_jQb6Iy5f1_2),.dout(w_dff_B_MUmWnAOJ1_2),.clk(gclk));
	jdff dff_B_aLcJ985A1_2(.din(w_dff_B_MUmWnAOJ1_2),.dout(w_dff_B_aLcJ985A1_2),.clk(gclk));
	jdff dff_B_UAI8SVqq1_2(.din(w_dff_B_aLcJ985A1_2),.dout(w_dff_B_UAI8SVqq1_2),.clk(gclk));
	jdff dff_B_Z0a9KuK07_2(.din(n1221),.dout(w_dff_B_Z0a9KuK07_2),.clk(gclk));
	jdff dff_B_fvxKhTZJ1_1(.din(n1184),.dout(w_dff_B_fvxKhTZJ1_1),.clk(gclk));
	jdff dff_B_veLj3kF07_2(.din(n1079),.dout(w_dff_B_veLj3kF07_2),.clk(gclk));
	jdff dff_B_O7PMupaH6_2(.din(w_dff_B_veLj3kF07_2),.dout(w_dff_B_O7PMupaH6_2),.clk(gclk));
	jdff dff_B_YOWYBIXb8_2(.din(w_dff_B_O7PMupaH6_2),.dout(w_dff_B_YOWYBIXb8_2),.clk(gclk));
	jdff dff_B_DQTMxhKZ0_2(.din(w_dff_B_YOWYBIXb8_2),.dout(w_dff_B_DQTMxhKZ0_2),.clk(gclk));
	jdff dff_B_AMbMvFhE4_2(.din(w_dff_B_DQTMxhKZ0_2),.dout(w_dff_B_AMbMvFhE4_2),.clk(gclk));
	jdff dff_B_IbYMGAOT7_2(.din(w_dff_B_AMbMvFhE4_2),.dout(w_dff_B_IbYMGAOT7_2),.clk(gclk));
	jdff dff_B_yAzojypG2_2(.din(w_dff_B_IbYMGAOT7_2),.dout(w_dff_B_yAzojypG2_2),.clk(gclk));
	jdff dff_B_GDrmqKIT8_2(.din(w_dff_B_yAzojypG2_2),.dout(w_dff_B_GDrmqKIT8_2),.clk(gclk));
	jdff dff_B_z0gKijmK6_2(.din(w_dff_B_GDrmqKIT8_2),.dout(w_dff_B_z0gKijmK6_2),.clk(gclk));
	jdff dff_B_aQoWeWUe4_2(.din(w_dff_B_z0gKijmK6_2),.dout(w_dff_B_aQoWeWUe4_2),.clk(gclk));
	jdff dff_B_D00xBbtZ1_2(.din(w_dff_B_aQoWeWUe4_2),.dout(w_dff_B_D00xBbtZ1_2),.clk(gclk));
	jdff dff_B_AMRwQ9s03_2(.din(w_dff_B_D00xBbtZ1_2),.dout(w_dff_B_AMRwQ9s03_2),.clk(gclk));
	jdff dff_B_WYyPk8ze3_2(.din(w_dff_B_AMRwQ9s03_2),.dout(w_dff_B_WYyPk8ze3_2),.clk(gclk));
	jdff dff_B_6jHS5wNb1_2(.din(w_dff_B_WYyPk8ze3_2),.dout(w_dff_B_6jHS5wNb1_2),.clk(gclk));
	jdff dff_B_5aKXzY7B5_2(.din(w_dff_B_6jHS5wNb1_2),.dout(w_dff_B_5aKXzY7B5_2),.clk(gclk));
	jdff dff_B_O84dZUmr6_2(.din(w_dff_B_5aKXzY7B5_2),.dout(w_dff_B_O84dZUmr6_2),.clk(gclk));
	jdff dff_B_2CR7ZkHZ7_2(.din(w_dff_B_O84dZUmr6_2),.dout(w_dff_B_2CR7ZkHZ7_2),.clk(gclk));
	jdff dff_B_BjioOdj92_2(.din(w_dff_B_2CR7ZkHZ7_2),.dout(w_dff_B_BjioOdj92_2),.clk(gclk));
	jdff dff_B_iCCPp6X70_2(.din(w_dff_B_BjioOdj92_2),.dout(w_dff_B_iCCPp6X70_2),.clk(gclk));
	jdff dff_B_3f60c6z12_2(.din(w_dff_B_iCCPp6X70_2),.dout(w_dff_B_3f60c6z12_2),.clk(gclk));
	jdff dff_B_6XKfNODF8_2(.din(w_dff_B_3f60c6z12_2),.dout(w_dff_B_6XKfNODF8_2),.clk(gclk));
	jdff dff_B_QT9H3YyO9_2(.din(w_dff_B_6XKfNODF8_2),.dout(w_dff_B_QT9H3YyO9_2),.clk(gclk));
	jdff dff_B_WpwaJj4C1_2(.din(w_dff_B_QT9H3YyO9_2),.dout(w_dff_B_WpwaJj4C1_2),.clk(gclk));
	jdff dff_B_RiuwrtiS3_2(.din(w_dff_B_WpwaJj4C1_2),.dout(w_dff_B_RiuwrtiS3_2),.clk(gclk));
	jdff dff_B_CcpcWgtq1_2(.din(n1123),.dout(w_dff_B_CcpcWgtq1_2),.clk(gclk));
	jdff dff_B_RJaWybtq6_1(.din(n1080),.dout(w_dff_B_RJaWybtq6_1),.clk(gclk));
	jdff dff_B_gZBphBBI3_2(.din(n981),.dout(w_dff_B_gZBphBBI3_2),.clk(gclk));
	jdff dff_B_SR17P8wr8_2(.din(w_dff_B_gZBphBBI3_2),.dout(w_dff_B_SR17P8wr8_2),.clk(gclk));
	jdff dff_B_FxIyvZ0Q3_2(.din(w_dff_B_SR17P8wr8_2),.dout(w_dff_B_FxIyvZ0Q3_2),.clk(gclk));
	jdff dff_B_Rjvzmweo7_2(.din(w_dff_B_FxIyvZ0Q3_2),.dout(w_dff_B_Rjvzmweo7_2),.clk(gclk));
	jdff dff_B_dQXVGhtG9_2(.din(w_dff_B_Rjvzmweo7_2),.dout(w_dff_B_dQXVGhtG9_2),.clk(gclk));
	jdff dff_B_d6NWEL8l7_2(.din(w_dff_B_dQXVGhtG9_2),.dout(w_dff_B_d6NWEL8l7_2),.clk(gclk));
	jdff dff_B_qtRC3AJQ5_2(.din(w_dff_B_d6NWEL8l7_2),.dout(w_dff_B_qtRC3AJQ5_2),.clk(gclk));
	jdff dff_B_xPABRAl62_2(.din(w_dff_B_qtRC3AJQ5_2),.dout(w_dff_B_xPABRAl62_2),.clk(gclk));
	jdff dff_B_004D1zQR1_2(.din(w_dff_B_xPABRAl62_2),.dout(w_dff_B_004D1zQR1_2),.clk(gclk));
	jdff dff_B_sZxMmARE0_2(.din(w_dff_B_004D1zQR1_2),.dout(w_dff_B_sZxMmARE0_2),.clk(gclk));
	jdff dff_B_mDvlIhhp8_2(.din(w_dff_B_sZxMmARE0_2),.dout(w_dff_B_mDvlIhhp8_2),.clk(gclk));
	jdff dff_B_NItKVYYn2_2(.din(w_dff_B_mDvlIhhp8_2),.dout(w_dff_B_NItKVYYn2_2),.clk(gclk));
	jdff dff_B_rj8huoSf4_2(.din(w_dff_B_NItKVYYn2_2),.dout(w_dff_B_rj8huoSf4_2),.clk(gclk));
	jdff dff_B_blTyxex25_2(.din(w_dff_B_rj8huoSf4_2),.dout(w_dff_B_blTyxex25_2),.clk(gclk));
	jdff dff_B_yCObGZKb5_2(.din(w_dff_B_blTyxex25_2),.dout(w_dff_B_yCObGZKb5_2),.clk(gclk));
	jdff dff_B_mWNBCjqY6_2(.din(w_dff_B_yCObGZKb5_2),.dout(w_dff_B_mWNBCjqY6_2),.clk(gclk));
	jdff dff_B_XqvcoNFE0_2(.din(w_dff_B_mWNBCjqY6_2),.dout(w_dff_B_XqvcoNFE0_2),.clk(gclk));
	jdff dff_B_s3P77hdo3_2(.din(w_dff_B_XqvcoNFE0_2),.dout(w_dff_B_s3P77hdo3_2),.clk(gclk));
	jdff dff_B_hW4utQGO1_2(.din(w_dff_B_s3P77hdo3_2),.dout(w_dff_B_hW4utQGO1_2),.clk(gclk));
	jdff dff_B_7I4Blpxa0_2(.din(w_dff_B_hW4utQGO1_2),.dout(w_dff_B_7I4Blpxa0_2),.clk(gclk));
	jdff dff_B_L1lMMz1t6_2(.din(w_dff_B_7I4Blpxa0_2),.dout(w_dff_B_L1lMMz1t6_2),.clk(gclk));
	jdff dff_B_TUzQBg6C0_2(.din(n1018),.dout(w_dff_B_TUzQBg6C0_2),.clk(gclk));
	jdff dff_B_og15hhse0_1(.din(n982),.dout(w_dff_B_og15hhse0_1),.clk(gclk));
	jdff dff_B_NTBdzeu70_2(.din(n876),.dout(w_dff_B_NTBdzeu70_2),.clk(gclk));
	jdff dff_B_o8lAKN3h5_2(.din(w_dff_B_NTBdzeu70_2),.dout(w_dff_B_o8lAKN3h5_2),.clk(gclk));
	jdff dff_B_0JO8cvJI1_2(.din(w_dff_B_o8lAKN3h5_2),.dout(w_dff_B_0JO8cvJI1_2),.clk(gclk));
	jdff dff_B_apTJhYpV8_2(.din(w_dff_B_0JO8cvJI1_2),.dout(w_dff_B_apTJhYpV8_2),.clk(gclk));
	jdff dff_B_rgKonn0v0_2(.din(w_dff_B_apTJhYpV8_2),.dout(w_dff_B_rgKonn0v0_2),.clk(gclk));
	jdff dff_B_fApqZ5Nf5_2(.din(w_dff_B_rgKonn0v0_2),.dout(w_dff_B_fApqZ5Nf5_2),.clk(gclk));
	jdff dff_B_qOp703cz8_2(.din(w_dff_B_fApqZ5Nf5_2),.dout(w_dff_B_qOp703cz8_2),.clk(gclk));
	jdff dff_B_ylc0NLGw3_2(.din(w_dff_B_qOp703cz8_2),.dout(w_dff_B_ylc0NLGw3_2),.clk(gclk));
	jdff dff_B_IIPZQFjA2_2(.din(w_dff_B_ylc0NLGw3_2),.dout(w_dff_B_IIPZQFjA2_2),.clk(gclk));
	jdff dff_B_I3Y7cDo83_2(.din(w_dff_B_IIPZQFjA2_2),.dout(w_dff_B_I3Y7cDo83_2),.clk(gclk));
	jdff dff_B_JEheRk3y4_2(.din(w_dff_B_I3Y7cDo83_2),.dout(w_dff_B_JEheRk3y4_2),.clk(gclk));
	jdff dff_B_MNdHRZgK1_2(.din(w_dff_B_JEheRk3y4_2),.dout(w_dff_B_MNdHRZgK1_2),.clk(gclk));
	jdff dff_B_HuO5DTko5_2(.din(w_dff_B_MNdHRZgK1_2),.dout(w_dff_B_HuO5DTko5_2),.clk(gclk));
	jdff dff_B_5byUhrvB8_2(.din(w_dff_B_HuO5DTko5_2),.dout(w_dff_B_5byUhrvB8_2),.clk(gclk));
	jdff dff_B_TGNBIzIj4_2(.din(w_dff_B_5byUhrvB8_2),.dout(w_dff_B_TGNBIzIj4_2),.clk(gclk));
	jdff dff_B_iNOV77LL4_2(.din(w_dff_B_TGNBIzIj4_2),.dout(w_dff_B_iNOV77LL4_2),.clk(gclk));
	jdff dff_B_8OHwCIHs5_2(.din(w_dff_B_iNOV77LL4_2),.dout(w_dff_B_8OHwCIHs5_2),.clk(gclk));
	jdff dff_B_TXHiw2xj9_2(.din(w_dff_B_8OHwCIHs5_2),.dout(w_dff_B_TXHiw2xj9_2),.clk(gclk));
	jdff dff_B_C2tPhRZm2_2(.din(n913),.dout(w_dff_B_C2tPhRZm2_2),.clk(gclk));
	jdff dff_B_I2zCEZrO8_1(.din(n877),.dout(w_dff_B_I2zCEZrO8_1),.clk(gclk));
	jdff dff_B_3GSWQHF03_2(.din(n777),.dout(w_dff_B_3GSWQHF03_2),.clk(gclk));
	jdff dff_B_WzhtIyi69_2(.din(w_dff_B_3GSWQHF03_2),.dout(w_dff_B_WzhtIyi69_2),.clk(gclk));
	jdff dff_B_KNNWknm91_2(.din(w_dff_B_WzhtIyi69_2),.dout(w_dff_B_KNNWknm91_2),.clk(gclk));
	jdff dff_B_zXi14C1v5_2(.din(w_dff_B_KNNWknm91_2),.dout(w_dff_B_zXi14C1v5_2),.clk(gclk));
	jdff dff_B_u93RiUpC9_2(.din(w_dff_B_zXi14C1v5_2),.dout(w_dff_B_u93RiUpC9_2),.clk(gclk));
	jdff dff_B_DYSMGqam8_2(.din(w_dff_B_u93RiUpC9_2),.dout(w_dff_B_DYSMGqam8_2),.clk(gclk));
	jdff dff_B_pYaZClYR5_2(.din(w_dff_B_DYSMGqam8_2),.dout(w_dff_B_pYaZClYR5_2),.clk(gclk));
	jdff dff_B_lmerLkGA4_2(.din(w_dff_B_pYaZClYR5_2),.dout(w_dff_B_lmerLkGA4_2),.clk(gclk));
	jdff dff_B_hsQramjb0_2(.din(w_dff_B_lmerLkGA4_2),.dout(w_dff_B_hsQramjb0_2),.clk(gclk));
	jdff dff_B_ehVgmDyt9_2(.din(w_dff_B_hsQramjb0_2),.dout(w_dff_B_ehVgmDyt9_2),.clk(gclk));
	jdff dff_B_GvKI84w06_2(.din(w_dff_B_ehVgmDyt9_2),.dout(w_dff_B_GvKI84w06_2),.clk(gclk));
	jdff dff_B_33xAjp1R9_2(.din(w_dff_B_GvKI84w06_2),.dout(w_dff_B_33xAjp1R9_2),.clk(gclk));
	jdff dff_B_EQnXRH0y8_2(.din(w_dff_B_33xAjp1R9_2),.dout(w_dff_B_EQnXRH0y8_2),.clk(gclk));
	jdff dff_B_I8zPB7qr6_2(.din(w_dff_B_EQnXRH0y8_2),.dout(w_dff_B_I8zPB7qr6_2),.clk(gclk));
	jdff dff_B_e9sc4Qcq2_2(.din(w_dff_B_I8zPB7qr6_2),.dout(w_dff_B_e9sc4Qcq2_2),.clk(gclk));
	jdff dff_B_3AHQoFUj2_2(.din(n807),.dout(w_dff_B_3AHQoFUj2_2),.clk(gclk));
	jdff dff_B_AAYbOxiG6_1(.din(n778),.dout(w_dff_B_AAYbOxiG6_1),.clk(gclk));
	jdff dff_B_9BcOlL2r4_2(.din(n684),.dout(w_dff_B_9BcOlL2r4_2),.clk(gclk));
	jdff dff_B_G7qarGdR7_2(.din(w_dff_B_9BcOlL2r4_2),.dout(w_dff_B_G7qarGdR7_2),.clk(gclk));
	jdff dff_B_EIgsg5sb1_2(.din(w_dff_B_G7qarGdR7_2),.dout(w_dff_B_EIgsg5sb1_2),.clk(gclk));
	jdff dff_B_eouyq3bX3_2(.din(w_dff_B_EIgsg5sb1_2),.dout(w_dff_B_eouyq3bX3_2),.clk(gclk));
	jdff dff_B_BmKJk8Qk9_2(.din(w_dff_B_eouyq3bX3_2),.dout(w_dff_B_BmKJk8Qk9_2),.clk(gclk));
	jdff dff_B_16jA1Ug15_2(.din(w_dff_B_BmKJk8Qk9_2),.dout(w_dff_B_16jA1Ug15_2),.clk(gclk));
	jdff dff_B_wTA4GIow3_2(.din(w_dff_B_16jA1Ug15_2),.dout(w_dff_B_wTA4GIow3_2),.clk(gclk));
	jdff dff_B_VycL0m8f3_2(.din(w_dff_B_wTA4GIow3_2),.dout(w_dff_B_VycL0m8f3_2),.clk(gclk));
	jdff dff_B_hmV5wMXC0_2(.din(w_dff_B_VycL0m8f3_2),.dout(w_dff_B_hmV5wMXC0_2),.clk(gclk));
	jdff dff_B_SiwSrSmM3_2(.din(w_dff_B_hmV5wMXC0_2),.dout(w_dff_B_SiwSrSmM3_2),.clk(gclk));
	jdff dff_B_gxMSgUNz3_2(.din(w_dff_B_SiwSrSmM3_2),.dout(w_dff_B_gxMSgUNz3_2),.clk(gclk));
	jdff dff_B_1XoMUMZI6_2(.din(w_dff_B_gxMSgUNz3_2),.dout(w_dff_B_1XoMUMZI6_2),.clk(gclk));
	jdff dff_B_3ZxVpABO3_2(.din(n707),.dout(w_dff_B_3ZxVpABO3_2),.clk(gclk));
	jdff dff_B_Lv9VvjLv5_1(.din(n685),.dout(w_dff_B_Lv9VvjLv5_1),.clk(gclk));
	jdff dff_B_cUdok9yr9_2(.din(n598),.dout(w_dff_B_cUdok9yr9_2),.clk(gclk));
	jdff dff_B_sxjP9MWd4_2(.din(w_dff_B_cUdok9yr9_2),.dout(w_dff_B_sxjP9MWd4_2),.clk(gclk));
	jdff dff_B_e4GuuxXM5_2(.din(w_dff_B_sxjP9MWd4_2),.dout(w_dff_B_e4GuuxXM5_2),.clk(gclk));
	jdff dff_B_hcW5uvqd2_2(.din(w_dff_B_e4GuuxXM5_2),.dout(w_dff_B_hcW5uvqd2_2),.clk(gclk));
	jdff dff_B_nxG1Sv2Z9_2(.din(w_dff_B_hcW5uvqd2_2),.dout(w_dff_B_nxG1Sv2Z9_2),.clk(gclk));
	jdff dff_B_Lx6rwnjp9_2(.din(w_dff_B_nxG1Sv2Z9_2),.dout(w_dff_B_Lx6rwnjp9_2),.clk(gclk));
	jdff dff_B_uImVwb7e6_2(.din(w_dff_B_Lx6rwnjp9_2),.dout(w_dff_B_uImVwb7e6_2),.clk(gclk));
	jdff dff_B_mD5yxOv23_2(.din(w_dff_B_uImVwb7e6_2),.dout(w_dff_B_mD5yxOv23_2),.clk(gclk));
	jdff dff_B_aiLqEprQ5_2(.din(w_dff_B_mD5yxOv23_2),.dout(w_dff_B_aiLqEprQ5_2),.clk(gclk));
	jdff dff_B_k4hePdx60_2(.din(n614),.dout(w_dff_B_k4hePdx60_2),.clk(gclk));
	jdff dff_B_2FQMyY2l4_2(.din(w_dff_B_k4hePdx60_2),.dout(w_dff_B_2FQMyY2l4_2),.clk(gclk));
	jdff dff_B_kqE9i7Nb1_1(.din(n599),.dout(w_dff_B_kqE9i7Nb1_1),.clk(gclk));
	jdff dff_B_e5UcNpW79_1(.din(w_dff_B_kqE9i7Nb1_1),.dout(w_dff_B_e5UcNpW79_1),.clk(gclk));
	jdff dff_B_uhZNfmV57_1(.din(w_dff_B_e5UcNpW79_1),.dout(w_dff_B_uhZNfmV57_1),.clk(gclk));
	jdff dff_B_yUGuLAXp2_1(.din(w_dff_B_uhZNfmV57_1),.dout(w_dff_B_yUGuLAXp2_1),.clk(gclk));
	jdff dff_B_jAyon4UW6_1(.din(w_dff_B_yUGuLAXp2_1),.dout(w_dff_B_jAyon4UW6_1),.clk(gclk));
	jdff dff_B_bUtnm8xz7_1(.din(w_dff_B_jAyon4UW6_1),.dout(w_dff_B_bUtnm8xz7_1),.clk(gclk));
	jdff dff_B_jTeyabpQ6_0(.din(n528),.dout(w_dff_B_jTeyabpQ6_0),.clk(gclk));
	jdff dff_B_BR1rDjUz4_0(.din(w_dff_B_jTeyabpQ6_0),.dout(w_dff_B_BR1rDjUz4_0),.clk(gclk));
	jdff dff_A_v4WlWYID6_0(.dout(w_n527_0[0]),.din(w_dff_A_v4WlWYID6_0),.clk(gclk));
	jdff dff_A_j08K9JPj0_0(.dout(w_dff_A_v4WlWYID6_0),.din(w_dff_A_j08K9JPj0_0),.clk(gclk));
	jdff dff_A_FLv3uGPk2_0(.dout(w_dff_A_j08K9JPj0_0),.din(w_dff_A_FLv3uGPk2_0),.clk(gclk));
	jdff dff_B_O5bHpvuc3_1(.din(n521),.dout(w_dff_B_O5bHpvuc3_1),.clk(gclk));
	jdff dff_A_B9LfuwoA9_0(.dout(w_n446_0[0]),.din(w_dff_A_B9LfuwoA9_0),.clk(gclk));
	jdff dff_A_8Or30avU8_1(.dout(w_n446_0[1]),.din(w_dff_A_8Or30avU8_1),.clk(gclk));
	jdff dff_A_KPFWeGym0_1(.dout(w_dff_A_8Or30avU8_1),.din(w_dff_A_KPFWeGym0_1),.clk(gclk));
	jdff dff_A_nWoJEuQb5_1(.dout(w_n519_0[1]),.din(w_dff_A_nWoJEuQb5_1),.clk(gclk));
	jdff dff_A_fmU5U7Rz6_1(.dout(w_dff_A_nWoJEuQb5_1),.din(w_dff_A_fmU5U7Rz6_1),.clk(gclk));
	jdff dff_A_7n3N5W964_1(.dout(w_dff_A_fmU5U7Rz6_1),.din(w_dff_A_7n3N5W964_1),.clk(gclk));
	jdff dff_A_tLR7lvQq3_1(.dout(w_dff_A_7n3N5W964_1),.din(w_dff_A_tLR7lvQq3_1),.clk(gclk));
	jdff dff_A_YQ3K9KNn2_1(.dout(w_dff_A_tLR7lvQq3_1),.din(w_dff_A_YQ3K9KNn2_1),.clk(gclk));
	jdff dff_A_fhhOmcMR1_1(.dout(w_dff_A_YQ3K9KNn2_1),.din(w_dff_A_fhhOmcMR1_1),.clk(gclk));
	jdff dff_B_e7rQmgAM9_1(.din(n1760),.dout(w_dff_B_e7rQmgAM9_1),.clk(gclk));
	jdff dff_A_KDTpLwao3_1(.dout(w_n1728_0[1]),.din(w_dff_A_KDTpLwao3_1),.clk(gclk));
	jdff dff_B_2R8ssFfu8_1(.din(n1726),.dout(w_dff_B_2R8ssFfu8_1),.clk(gclk));
	jdff dff_B_4iEGNX4k6_2(.din(n1684),.dout(w_dff_B_4iEGNX4k6_2),.clk(gclk));
	jdff dff_B_bkqm7Fyg4_2(.din(w_dff_B_4iEGNX4k6_2),.dout(w_dff_B_bkqm7Fyg4_2),.clk(gclk));
	jdff dff_B_Asz62aTZ5_2(.din(w_dff_B_bkqm7Fyg4_2),.dout(w_dff_B_Asz62aTZ5_2),.clk(gclk));
	jdff dff_B_KWL87JfM9_2(.din(w_dff_B_Asz62aTZ5_2),.dout(w_dff_B_KWL87JfM9_2),.clk(gclk));
	jdff dff_B_g0ZBFLtY1_2(.din(w_dff_B_KWL87JfM9_2),.dout(w_dff_B_g0ZBFLtY1_2),.clk(gclk));
	jdff dff_B_oP6nXBda2_2(.din(w_dff_B_g0ZBFLtY1_2),.dout(w_dff_B_oP6nXBda2_2),.clk(gclk));
	jdff dff_B_hch7V9117_2(.din(w_dff_B_oP6nXBda2_2),.dout(w_dff_B_hch7V9117_2),.clk(gclk));
	jdff dff_B_nZY7GlY08_2(.din(w_dff_B_hch7V9117_2),.dout(w_dff_B_nZY7GlY08_2),.clk(gclk));
	jdff dff_B_VwdoIWdU2_2(.din(w_dff_B_nZY7GlY08_2),.dout(w_dff_B_VwdoIWdU2_2),.clk(gclk));
	jdff dff_B_yz6C6NLB2_2(.din(w_dff_B_VwdoIWdU2_2),.dout(w_dff_B_yz6C6NLB2_2),.clk(gclk));
	jdff dff_B_XoeOYaGt0_2(.din(w_dff_B_yz6C6NLB2_2),.dout(w_dff_B_XoeOYaGt0_2),.clk(gclk));
	jdff dff_B_e87aAuAG6_2(.din(w_dff_B_XoeOYaGt0_2),.dout(w_dff_B_e87aAuAG6_2),.clk(gclk));
	jdff dff_B_WbPBm8bm5_2(.din(w_dff_B_e87aAuAG6_2),.dout(w_dff_B_WbPBm8bm5_2),.clk(gclk));
	jdff dff_B_9mvFTDlZ6_2(.din(w_dff_B_WbPBm8bm5_2),.dout(w_dff_B_9mvFTDlZ6_2),.clk(gclk));
	jdff dff_B_TnF7dwqv5_2(.din(w_dff_B_9mvFTDlZ6_2),.dout(w_dff_B_TnF7dwqv5_2),.clk(gclk));
	jdff dff_B_9vMO3mb44_2(.din(w_dff_B_TnF7dwqv5_2),.dout(w_dff_B_9vMO3mb44_2),.clk(gclk));
	jdff dff_B_xfAlWrTt6_2(.din(w_dff_B_9vMO3mb44_2),.dout(w_dff_B_xfAlWrTt6_2),.clk(gclk));
	jdff dff_B_iKcIK2D28_2(.din(w_dff_B_xfAlWrTt6_2),.dout(w_dff_B_iKcIK2D28_2),.clk(gclk));
	jdff dff_B_EtPQ2LJz7_2(.din(w_dff_B_iKcIK2D28_2),.dout(w_dff_B_EtPQ2LJz7_2),.clk(gclk));
	jdff dff_B_iedRFMJC1_2(.din(w_dff_B_EtPQ2LJz7_2),.dout(w_dff_B_iedRFMJC1_2),.clk(gclk));
	jdff dff_B_fhj2ej8M5_2(.din(w_dff_B_iedRFMJC1_2),.dout(w_dff_B_fhj2ej8M5_2),.clk(gclk));
	jdff dff_B_UNn6pOEv9_2(.din(w_dff_B_fhj2ej8M5_2),.dout(w_dff_B_UNn6pOEv9_2),.clk(gclk));
	jdff dff_B_nJQaEDV28_2(.din(w_dff_B_UNn6pOEv9_2),.dout(w_dff_B_nJQaEDV28_2),.clk(gclk));
	jdff dff_B_iL0B8Hav0_2(.din(w_dff_B_nJQaEDV28_2),.dout(w_dff_B_iL0B8Hav0_2),.clk(gclk));
	jdff dff_B_bbmwxhks0_2(.din(w_dff_B_iL0B8Hav0_2),.dout(w_dff_B_bbmwxhks0_2),.clk(gclk));
	jdff dff_B_1Yc9nh9s0_2(.din(w_dff_B_bbmwxhks0_2),.dout(w_dff_B_1Yc9nh9s0_2),.clk(gclk));
	jdff dff_B_8cqLZpNH1_2(.din(w_dff_B_1Yc9nh9s0_2),.dout(w_dff_B_8cqLZpNH1_2),.clk(gclk));
	jdff dff_B_cI5Fv32S6_2(.din(w_dff_B_8cqLZpNH1_2),.dout(w_dff_B_cI5Fv32S6_2),.clk(gclk));
	jdff dff_B_GoHKKvWu2_2(.din(w_dff_B_cI5Fv32S6_2),.dout(w_dff_B_GoHKKvWu2_2),.clk(gclk));
	jdff dff_B_tBnbRVxq3_2(.din(w_dff_B_GoHKKvWu2_2),.dout(w_dff_B_tBnbRVxq3_2),.clk(gclk));
	jdff dff_B_jYejXZNb8_2(.din(w_dff_B_tBnbRVxq3_2),.dout(w_dff_B_jYejXZNb8_2),.clk(gclk));
	jdff dff_B_WYnXZsUE5_2(.din(w_dff_B_jYejXZNb8_2),.dout(w_dff_B_WYnXZsUE5_2),.clk(gclk));
	jdff dff_B_KfJcRmMU6_2(.din(w_dff_B_WYnXZsUE5_2),.dout(w_dff_B_KfJcRmMU6_2),.clk(gclk));
	jdff dff_B_Q6oF7kVo0_2(.din(w_dff_B_KfJcRmMU6_2),.dout(w_dff_B_Q6oF7kVo0_2),.clk(gclk));
	jdff dff_B_6i1qVTkJ0_2(.din(w_dff_B_Q6oF7kVo0_2),.dout(w_dff_B_6i1qVTkJ0_2),.clk(gclk));
	jdff dff_B_lEKhbbch0_2(.din(w_dff_B_6i1qVTkJ0_2),.dout(w_dff_B_lEKhbbch0_2),.clk(gclk));
	jdff dff_B_9CUcbquI8_2(.din(w_dff_B_lEKhbbch0_2),.dout(w_dff_B_9CUcbquI8_2),.clk(gclk));
	jdff dff_B_76qYG72q0_2(.din(w_dff_B_9CUcbquI8_2),.dout(w_dff_B_76qYG72q0_2),.clk(gclk));
	jdff dff_B_8LbPNQOY7_2(.din(w_dff_B_76qYG72q0_2),.dout(w_dff_B_8LbPNQOY7_2),.clk(gclk));
	jdff dff_B_phyzLvqW6_2(.din(w_dff_B_8LbPNQOY7_2),.dout(w_dff_B_phyzLvqW6_2),.clk(gclk));
	jdff dff_B_AXkeI9wH9_2(.din(w_dff_B_phyzLvqW6_2),.dout(w_dff_B_AXkeI9wH9_2),.clk(gclk));
	jdff dff_B_wWFUPvyS6_2(.din(w_dff_B_AXkeI9wH9_2),.dout(w_dff_B_wWFUPvyS6_2),.clk(gclk));
	jdff dff_B_al3nY6R34_2(.din(w_dff_B_wWFUPvyS6_2),.dout(w_dff_B_al3nY6R34_2),.clk(gclk));
	jdff dff_B_d02Ejx0N3_2(.din(w_dff_B_al3nY6R34_2),.dout(w_dff_B_d02Ejx0N3_2),.clk(gclk));
	jdff dff_B_JqS5l66B8_2(.din(w_dff_B_d02Ejx0N3_2),.dout(w_dff_B_JqS5l66B8_2),.clk(gclk));
	jdff dff_B_MJeIncJl2_2(.din(w_dff_B_JqS5l66B8_2),.dout(w_dff_B_MJeIncJl2_2),.clk(gclk));
	jdff dff_B_3RPeXNwE6_2(.din(w_dff_B_MJeIncJl2_2),.dout(w_dff_B_3RPeXNwE6_2),.clk(gclk));
	jdff dff_B_BKXFm4qV6_2(.din(w_dff_B_3RPeXNwE6_2),.dout(w_dff_B_BKXFm4qV6_2),.clk(gclk));
	jdff dff_B_eRWRvYFs0_2(.din(w_dff_B_BKXFm4qV6_2),.dout(w_dff_B_eRWRvYFs0_2),.clk(gclk));
	jdff dff_B_vidOmM8E0_2(.din(n1687),.dout(w_dff_B_vidOmM8E0_2),.clk(gclk));
	jdff dff_B_6E1WzGAH5_1(.din(n1685),.dout(w_dff_B_6E1WzGAH5_1),.clk(gclk));
	jdff dff_B_GMXVFmo87_2(.din(n1633),.dout(w_dff_B_GMXVFmo87_2),.clk(gclk));
	jdff dff_B_VhYiU9p90_2(.din(w_dff_B_GMXVFmo87_2),.dout(w_dff_B_VhYiU9p90_2),.clk(gclk));
	jdff dff_B_7VmPgVOa7_2(.din(w_dff_B_VhYiU9p90_2),.dout(w_dff_B_7VmPgVOa7_2),.clk(gclk));
	jdff dff_B_UBk9Vfuf4_2(.din(w_dff_B_7VmPgVOa7_2),.dout(w_dff_B_UBk9Vfuf4_2),.clk(gclk));
	jdff dff_B_z95ndv0s8_2(.din(w_dff_B_UBk9Vfuf4_2),.dout(w_dff_B_z95ndv0s8_2),.clk(gclk));
	jdff dff_B_Gj9vx9kH3_2(.din(w_dff_B_z95ndv0s8_2),.dout(w_dff_B_Gj9vx9kH3_2),.clk(gclk));
	jdff dff_B_HHglZIgO7_2(.din(w_dff_B_Gj9vx9kH3_2),.dout(w_dff_B_HHglZIgO7_2),.clk(gclk));
	jdff dff_B_WmX87N4j8_2(.din(w_dff_B_HHglZIgO7_2),.dout(w_dff_B_WmX87N4j8_2),.clk(gclk));
	jdff dff_B_aCjEWD9j5_2(.din(w_dff_B_WmX87N4j8_2),.dout(w_dff_B_aCjEWD9j5_2),.clk(gclk));
	jdff dff_B_M0JZtGP57_2(.din(w_dff_B_aCjEWD9j5_2),.dout(w_dff_B_M0JZtGP57_2),.clk(gclk));
	jdff dff_B_ID2B8IpB5_2(.din(w_dff_B_M0JZtGP57_2),.dout(w_dff_B_ID2B8IpB5_2),.clk(gclk));
	jdff dff_B_X9mdq5Y74_2(.din(w_dff_B_ID2B8IpB5_2),.dout(w_dff_B_X9mdq5Y74_2),.clk(gclk));
	jdff dff_B_rVSyZLor2_2(.din(w_dff_B_X9mdq5Y74_2),.dout(w_dff_B_rVSyZLor2_2),.clk(gclk));
	jdff dff_B_WPn96d4Q4_2(.din(w_dff_B_rVSyZLor2_2),.dout(w_dff_B_WPn96d4Q4_2),.clk(gclk));
	jdff dff_B_Z71cg9912_2(.din(w_dff_B_WPn96d4Q4_2),.dout(w_dff_B_Z71cg9912_2),.clk(gclk));
	jdff dff_B_ggK1QwuK4_2(.din(w_dff_B_Z71cg9912_2),.dout(w_dff_B_ggK1QwuK4_2),.clk(gclk));
	jdff dff_B_q9RypAz71_2(.din(w_dff_B_ggK1QwuK4_2),.dout(w_dff_B_q9RypAz71_2),.clk(gclk));
	jdff dff_B_D8UPfHhv9_2(.din(w_dff_B_q9RypAz71_2),.dout(w_dff_B_D8UPfHhv9_2),.clk(gclk));
	jdff dff_B_f6zRBvxY1_2(.din(w_dff_B_D8UPfHhv9_2),.dout(w_dff_B_f6zRBvxY1_2),.clk(gclk));
	jdff dff_B_V8j1UlyI1_2(.din(w_dff_B_f6zRBvxY1_2),.dout(w_dff_B_V8j1UlyI1_2),.clk(gclk));
	jdff dff_B_2C6bwF0m4_2(.din(w_dff_B_V8j1UlyI1_2),.dout(w_dff_B_2C6bwF0m4_2),.clk(gclk));
	jdff dff_B_nmDxdhXZ6_2(.din(w_dff_B_2C6bwF0m4_2),.dout(w_dff_B_nmDxdhXZ6_2),.clk(gclk));
	jdff dff_B_n5eS17F55_2(.din(w_dff_B_nmDxdhXZ6_2),.dout(w_dff_B_n5eS17F55_2),.clk(gclk));
	jdff dff_B_LVAZMxIP2_2(.din(w_dff_B_n5eS17F55_2),.dout(w_dff_B_LVAZMxIP2_2),.clk(gclk));
	jdff dff_B_LXhgr5xo7_2(.din(w_dff_B_LVAZMxIP2_2),.dout(w_dff_B_LXhgr5xo7_2),.clk(gclk));
	jdff dff_B_kWigknG92_2(.din(w_dff_B_LXhgr5xo7_2),.dout(w_dff_B_kWigknG92_2),.clk(gclk));
	jdff dff_B_7gnDFMqR8_2(.din(w_dff_B_kWigknG92_2),.dout(w_dff_B_7gnDFMqR8_2),.clk(gclk));
	jdff dff_B_Yw4uZofs5_2(.din(w_dff_B_7gnDFMqR8_2),.dout(w_dff_B_Yw4uZofs5_2),.clk(gclk));
	jdff dff_B_qQ3UMM6B4_2(.din(w_dff_B_Yw4uZofs5_2),.dout(w_dff_B_qQ3UMM6B4_2),.clk(gclk));
	jdff dff_B_lpDWz5xn2_2(.din(w_dff_B_qQ3UMM6B4_2),.dout(w_dff_B_lpDWz5xn2_2),.clk(gclk));
	jdff dff_B_A2nZeAre6_2(.din(w_dff_B_lpDWz5xn2_2),.dout(w_dff_B_A2nZeAre6_2),.clk(gclk));
	jdff dff_B_PKbWz6PF5_2(.din(w_dff_B_A2nZeAre6_2),.dout(w_dff_B_PKbWz6PF5_2),.clk(gclk));
	jdff dff_B_DHZPbG821_2(.din(w_dff_B_PKbWz6PF5_2),.dout(w_dff_B_DHZPbG821_2),.clk(gclk));
	jdff dff_B_KSbdqQjN2_2(.din(w_dff_B_DHZPbG821_2),.dout(w_dff_B_KSbdqQjN2_2),.clk(gclk));
	jdff dff_B_beORuMVy1_2(.din(w_dff_B_KSbdqQjN2_2),.dout(w_dff_B_beORuMVy1_2),.clk(gclk));
	jdff dff_B_R7JfVrcH7_2(.din(w_dff_B_beORuMVy1_2),.dout(w_dff_B_R7JfVrcH7_2),.clk(gclk));
	jdff dff_B_GI5B6ONl5_2(.din(w_dff_B_R7JfVrcH7_2),.dout(w_dff_B_GI5B6ONl5_2),.clk(gclk));
	jdff dff_B_ntopK4Fq5_2(.din(w_dff_B_GI5B6ONl5_2),.dout(w_dff_B_ntopK4Fq5_2),.clk(gclk));
	jdff dff_B_lNBBb5Mf1_2(.din(w_dff_B_ntopK4Fq5_2),.dout(w_dff_B_lNBBb5Mf1_2),.clk(gclk));
	jdff dff_B_tkZPKKnO0_2(.din(w_dff_B_lNBBb5Mf1_2),.dout(w_dff_B_tkZPKKnO0_2),.clk(gclk));
	jdff dff_B_AGe4Ytyv9_2(.din(w_dff_B_tkZPKKnO0_2),.dout(w_dff_B_AGe4Ytyv9_2),.clk(gclk));
	jdff dff_B_7gf4WLNu5_2(.din(w_dff_B_AGe4Ytyv9_2),.dout(w_dff_B_7gf4WLNu5_2),.clk(gclk));
	jdff dff_B_N4mBQkgr0_2(.din(w_dff_B_7gf4WLNu5_2),.dout(w_dff_B_N4mBQkgr0_2),.clk(gclk));
	jdff dff_B_CzETjaGO4_2(.din(w_dff_B_N4mBQkgr0_2),.dout(w_dff_B_CzETjaGO4_2),.clk(gclk));
	jdff dff_B_oltETmjT9_2(.din(w_dff_B_CzETjaGO4_2),.dout(w_dff_B_oltETmjT9_2),.clk(gclk));
	jdff dff_B_dpZfKvVX0_2(.din(n1636),.dout(w_dff_B_dpZfKvVX0_2),.clk(gclk));
	jdff dff_B_QKibgKDa8_1(.din(n1634),.dout(w_dff_B_QKibgKDa8_1),.clk(gclk));
	jdff dff_B_1s5tCjko0_2(.din(n1576),.dout(w_dff_B_1s5tCjko0_2),.clk(gclk));
	jdff dff_B_0cI17qcD8_2(.din(w_dff_B_1s5tCjko0_2),.dout(w_dff_B_0cI17qcD8_2),.clk(gclk));
	jdff dff_B_58pf3EQF6_2(.din(w_dff_B_0cI17qcD8_2),.dout(w_dff_B_58pf3EQF6_2),.clk(gclk));
	jdff dff_B_8IaurN1Q8_2(.din(w_dff_B_58pf3EQF6_2),.dout(w_dff_B_8IaurN1Q8_2),.clk(gclk));
	jdff dff_B_km3FnPFm5_2(.din(w_dff_B_8IaurN1Q8_2),.dout(w_dff_B_km3FnPFm5_2),.clk(gclk));
	jdff dff_B_y6yZ3j9W2_2(.din(w_dff_B_km3FnPFm5_2),.dout(w_dff_B_y6yZ3j9W2_2),.clk(gclk));
	jdff dff_B_gocjZram1_2(.din(w_dff_B_y6yZ3j9W2_2),.dout(w_dff_B_gocjZram1_2),.clk(gclk));
	jdff dff_B_1IGagMmn9_2(.din(w_dff_B_gocjZram1_2),.dout(w_dff_B_1IGagMmn9_2),.clk(gclk));
	jdff dff_B_BoHTvwfo6_2(.din(w_dff_B_1IGagMmn9_2),.dout(w_dff_B_BoHTvwfo6_2),.clk(gclk));
	jdff dff_B_uqe3gkPo4_2(.din(w_dff_B_BoHTvwfo6_2),.dout(w_dff_B_uqe3gkPo4_2),.clk(gclk));
	jdff dff_B_wyfTh3fA1_2(.din(w_dff_B_uqe3gkPo4_2),.dout(w_dff_B_wyfTh3fA1_2),.clk(gclk));
	jdff dff_B_ItWn1yZr3_2(.din(w_dff_B_wyfTh3fA1_2),.dout(w_dff_B_ItWn1yZr3_2),.clk(gclk));
	jdff dff_B_rGeIIq0s7_2(.din(w_dff_B_ItWn1yZr3_2),.dout(w_dff_B_rGeIIq0s7_2),.clk(gclk));
	jdff dff_B_liAHa5p55_2(.din(w_dff_B_rGeIIq0s7_2),.dout(w_dff_B_liAHa5p55_2),.clk(gclk));
	jdff dff_B_1DOurXRH0_2(.din(w_dff_B_liAHa5p55_2),.dout(w_dff_B_1DOurXRH0_2),.clk(gclk));
	jdff dff_B_tuA5QtV19_2(.din(w_dff_B_1DOurXRH0_2),.dout(w_dff_B_tuA5QtV19_2),.clk(gclk));
	jdff dff_B_NpocvfLw3_2(.din(w_dff_B_tuA5QtV19_2),.dout(w_dff_B_NpocvfLw3_2),.clk(gclk));
	jdff dff_B_TmzCbW5E0_2(.din(w_dff_B_NpocvfLw3_2),.dout(w_dff_B_TmzCbW5E0_2),.clk(gclk));
	jdff dff_B_voIYm9O80_2(.din(w_dff_B_TmzCbW5E0_2),.dout(w_dff_B_voIYm9O80_2),.clk(gclk));
	jdff dff_B_9RW5tuQa4_2(.din(w_dff_B_voIYm9O80_2),.dout(w_dff_B_9RW5tuQa4_2),.clk(gclk));
	jdff dff_B_2qZB7d1W7_2(.din(w_dff_B_9RW5tuQa4_2),.dout(w_dff_B_2qZB7d1W7_2),.clk(gclk));
	jdff dff_B_oFQGmyHB9_2(.din(w_dff_B_2qZB7d1W7_2),.dout(w_dff_B_oFQGmyHB9_2),.clk(gclk));
	jdff dff_B_MleDO6jT0_2(.din(w_dff_B_oFQGmyHB9_2),.dout(w_dff_B_MleDO6jT0_2),.clk(gclk));
	jdff dff_B_TjcQ3fL30_2(.din(w_dff_B_MleDO6jT0_2),.dout(w_dff_B_TjcQ3fL30_2),.clk(gclk));
	jdff dff_B_iZRbspGT7_2(.din(w_dff_B_TjcQ3fL30_2),.dout(w_dff_B_iZRbspGT7_2),.clk(gclk));
	jdff dff_B_d0tsRWLF2_2(.din(w_dff_B_iZRbspGT7_2),.dout(w_dff_B_d0tsRWLF2_2),.clk(gclk));
	jdff dff_B_jUZ15Anr9_2(.din(w_dff_B_d0tsRWLF2_2),.dout(w_dff_B_jUZ15Anr9_2),.clk(gclk));
	jdff dff_B_pyT6AlUX6_2(.din(w_dff_B_jUZ15Anr9_2),.dout(w_dff_B_pyT6AlUX6_2),.clk(gclk));
	jdff dff_B_mNHUaxJS4_2(.din(w_dff_B_pyT6AlUX6_2),.dout(w_dff_B_mNHUaxJS4_2),.clk(gclk));
	jdff dff_B_NSULHQX49_2(.din(w_dff_B_mNHUaxJS4_2),.dout(w_dff_B_NSULHQX49_2),.clk(gclk));
	jdff dff_B_OJuYZUPj1_2(.din(w_dff_B_NSULHQX49_2),.dout(w_dff_B_OJuYZUPj1_2),.clk(gclk));
	jdff dff_B_2CPpwImG4_2(.din(w_dff_B_OJuYZUPj1_2),.dout(w_dff_B_2CPpwImG4_2),.clk(gclk));
	jdff dff_B_R4gpfeSf6_2(.din(w_dff_B_2CPpwImG4_2),.dout(w_dff_B_R4gpfeSf6_2),.clk(gclk));
	jdff dff_B_OE06QjU20_2(.din(w_dff_B_R4gpfeSf6_2),.dout(w_dff_B_OE06QjU20_2),.clk(gclk));
	jdff dff_B_GJgtE1tx4_2(.din(w_dff_B_OE06QjU20_2),.dout(w_dff_B_GJgtE1tx4_2),.clk(gclk));
	jdff dff_B_EQnZijLD5_2(.din(w_dff_B_GJgtE1tx4_2),.dout(w_dff_B_EQnZijLD5_2),.clk(gclk));
	jdff dff_B_grvRkOlY1_2(.din(w_dff_B_EQnZijLD5_2),.dout(w_dff_B_grvRkOlY1_2),.clk(gclk));
	jdff dff_B_FOsTG4KS8_2(.din(w_dff_B_grvRkOlY1_2),.dout(w_dff_B_FOsTG4KS8_2),.clk(gclk));
	jdff dff_B_Uu4Xc0fB8_2(.din(w_dff_B_FOsTG4KS8_2),.dout(w_dff_B_Uu4Xc0fB8_2),.clk(gclk));
	jdff dff_B_bVmSKT6a5_2(.din(w_dff_B_Uu4Xc0fB8_2),.dout(w_dff_B_bVmSKT6a5_2),.clk(gclk));
	jdff dff_B_gEEO3E7I5_2(.din(w_dff_B_bVmSKT6a5_2),.dout(w_dff_B_gEEO3E7I5_2),.clk(gclk));
	jdff dff_B_cPxo96Ll1_2(.din(n1579),.dout(w_dff_B_cPxo96Ll1_2),.clk(gclk));
	jdff dff_B_T6U1i5sD6_1(.din(n1577),.dout(w_dff_B_T6U1i5sD6_1),.clk(gclk));
	jdff dff_B_97QZtcbo8_2(.din(n1512),.dout(w_dff_B_97QZtcbo8_2),.clk(gclk));
	jdff dff_B_c8yOQlVH8_2(.din(w_dff_B_97QZtcbo8_2),.dout(w_dff_B_c8yOQlVH8_2),.clk(gclk));
	jdff dff_B_jX9lxqyI9_2(.din(w_dff_B_c8yOQlVH8_2),.dout(w_dff_B_jX9lxqyI9_2),.clk(gclk));
	jdff dff_B_r0VF3OLf9_2(.din(w_dff_B_jX9lxqyI9_2),.dout(w_dff_B_r0VF3OLf9_2),.clk(gclk));
	jdff dff_B_tFA5BSjr3_2(.din(w_dff_B_r0VF3OLf9_2),.dout(w_dff_B_tFA5BSjr3_2),.clk(gclk));
	jdff dff_B_uA5NaYnK9_2(.din(w_dff_B_tFA5BSjr3_2),.dout(w_dff_B_uA5NaYnK9_2),.clk(gclk));
	jdff dff_B_Jk9CC1OT6_2(.din(w_dff_B_uA5NaYnK9_2),.dout(w_dff_B_Jk9CC1OT6_2),.clk(gclk));
	jdff dff_B_F7eTZm5u2_2(.din(w_dff_B_Jk9CC1OT6_2),.dout(w_dff_B_F7eTZm5u2_2),.clk(gclk));
	jdff dff_B_ic8D8o6W3_2(.din(w_dff_B_F7eTZm5u2_2),.dout(w_dff_B_ic8D8o6W3_2),.clk(gclk));
	jdff dff_B_GSgUbhqP6_2(.din(w_dff_B_ic8D8o6W3_2),.dout(w_dff_B_GSgUbhqP6_2),.clk(gclk));
	jdff dff_B_BoKDD3bt7_2(.din(w_dff_B_GSgUbhqP6_2),.dout(w_dff_B_BoKDD3bt7_2),.clk(gclk));
	jdff dff_B_LWAtVUJ64_2(.din(w_dff_B_BoKDD3bt7_2),.dout(w_dff_B_LWAtVUJ64_2),.clk(gclk));
	jdff dff_B_RR532V0c8_2(.din(w_dff_B_LWAtVUJ64_2),.dout(w_dff_B_RR532V0c8_2),.clk(gclk));
	jdff dff_B_tXPXIhhT1_2(.din(w_dff_B_RR532V0c8_2),.dout(w_dff_B_tXPXIhhT1_2),.clk(gclk));
	jdff dff_B_QWD7vBpy0_2(.din(w_dff_B_tXPXIhhT1_2),.dout(w_dff_B_QWD7vBpy0_2),.clk(gclk));
	jdff dff_B_AyJpJwkY8_2(.din(w_dff_B_QWD7vBpy0_2),.dout(w_dff_B_AyJpJwkY8_2),.clk(gclk));
	jdff dff_B_Iv6ujFZS5_2(.din(w_dff_B_AyJpJwkY8_2),.dout(w_dff_B_Iv6ujFZS5_2),.clk(gclk));
	jdff dff_B_bRWMaYzq4_2(.din(w_dff_B_Iv6ujFZS5_2),.dout(w_dff_B_bRWMaYzq4_2),.clk(gclk));
	jdff dff_B_8HPVWGUP1_2(.din(w_dff_B_bRWMaYzq4_2),.dout(w_dff_B_8HPVWGUP1_2),.clk(gclk));
	jdff dff_B_3Horefdt7_2(.din(w_dff_B_8HPVWGUP1_2),.dout(w_dff_B_3Horefdt7_2),.clk(gclk));
	jdff dff_B_AOXHcnsf1_2(.din(w_dff_B_3Horefdt7_2),.dout(w_dff_B_AOXHcnsf1_2),.clk(gclk));
	jdff dff_B_Us2NEt0j0_2(.din(w_dff_B_AOXHcnsf1_2),.dout(w_dff_B_Us2NEt0j0_2),.clk(gclk));
	jdff dff_B_IKAzVBRv4_2(.din(w_dff_B_Us2NEt0j0_2),.dout(w_dff_B_IKAzVBRv4_2),.clk(gclk));
	jdff dff_B_HwS2VOr40_2(.din(w_dff_B_IKAzVBRv4_2),.dout(w_dff_B_HwS2VOr40_2),.clk(gclk));
	jdff dff_B_WSNp20hW8_2(.din(w_dff_B_HwS2VOr40_2),.dout(w_dff_B_WSNp20hW8_2),.clk(gclk));
	jdff dff_B_bYZ5SP0d3_2(.din(w_dff_B_WSNp20hW8_2),.dout(w_dff_B_bYZ5SP0d3_2),.clk(gclk));
	jdff dff_B_vLE5msUt3_2(.din(w_dff_B_bYZ5SP0d3_2),.dout(w_dff_B_vLE5msUt3_2),.clk(gclk));
	jdff dff_B_nhQYtNyl6_2(.din(w_dff_B_vLE5msUt3_2),.dout(w_dff_B_nhQYtNyl6_2),.clk(gclk));
	jdff dff_B_1W8p3sVY5_2(.din(w_dff_B_nhQYtNyl6_2),.dout(w_dff_B_1W8p3sVY5_2),.clk(gclk));
	jdff dff_B_cvQ4GP5F6_2(.din(w_dff_B_1W8p3sVY5_2),.dout(w_dff_B_cvQ4GP5F6_2),.clk(gclk));
	jdff dff_B_4I6nkLkQ3_2(.din(w_dff_B_cvQ4GP5F6_2),.dout(w_dff_B_4I6nkLkQ3_2),.clk(gclk));
	jdff dff_B_Jej9mtvo4_2(.din(w_dff_B_4I6nkLkQ3_2),.dout(w_dff_B_Jej9mtvo4_2),.clk(gclk));
	jdff dff_B_41G6egtG0_2(.din(w_dff_B_Jej9mtvo4_2),.dout(w_dff_B_41G6egtG0_2),.clk(gclk));
	jdff dff_B_b7RFWKmF2_2(.din(w_dff_B_41G6egtG0_2),.dout(w_dff_B_b7RFWKmF2_2),.clk(gclk));
	jdff dff_B_NtiGoyX29_2(.din(w_dff_B_b7RFWKmF2_2),.dout(w_dff_B_NtiGoyX29_2),.clk(gclk));
	jdff dff_B_mJ5yHz6i7_2(.din(w_dff_B_NtiGoyX29_2),.dout(w_dff_B_mJ5yHz6i7_2),.clk(gclk));
	jdff dff_B_64mFQgHf1_2(.din(w_dff_B_mJ5yHz6i7_2),.dout(w_dff_B_64mFQgHf1_2),.clk(gclk));
	jdff dff_B_a5IKWAgM2_2(.din(n1515),.dout(w_dff_B_a5IKWAgM2_2),.clk(gclk));
	jdff dff_B_yhcxjPXC0_1(.din(n1513),.dout(w_dff_B_yhcxjPXC0_1),.clk(gclk));
	jdff dff_B_pFIWHQes1_2(.din(n1441),.dout(w_dff_B_pFIWHQes1_2),.clk(gclk));
	jdff dff_B_GotnhCGT2_2(.din(w_dff_B_pFIWHQes1_2),.dout(w_dff_B_GotnhCGT2_2),.clk(gclk));
	jdff dff_B_LTlYs43I3_2(.din(w_dff_B_GotnhCGT2_2),.dout(w_dff_B_LTlYs43I3_2),.clk(gclk));
	jdff dff_B_RHS81jZB5_2(.din(w_dff_B_LTlYs43I3_2),.dout(w_dff_B_RHS81jZB5_2),.clk(gclk));
	jdff dff_B_S3RJH4Ws2_2(.din(w_dff_B_RHS81jZB5_2),.dout(w_dff_B_S3RJH4Ws2_2),.clk(gclk));
	jdff dff_B_Tm3D5mPt7_2(.din(w_dff_B_S3RJH4Ws2_2),.dout(w_dff_B_Tm3D5mPt7_2),.clk(gclk));
	jdff dff_B_WE3qqVPP9_2(.din(w_dff_B_Tm3D5mPt7_2),.dout(w_dff_B_WE3qqVPP9_2),.clk(gclk));
	jdff dff_B_uxT1D6338_2(.din(w_dff_B_WE3qqVPP9_2),.dout(w_dff_B_uxT1D6338_2),.clk(gclk));
	jdff dff_B_jMx5779a0_2(.din(w_dff_B_uxT1D6338_2),.dout(w_dff_B_jMx5779a0_2),.clk(gclk));
	jdff dff_B_v2xwKHeb4_2(.din(w_dff_B_jMx5779a0_2),.dout(w_dff_B_v2xwKHeb4_2),.clk(gclk));
	jdff dff_B_9jKtpsFI6_2(.din(w_dff_B_v2xwKHeb4_2),.dout(w_dff_B_9jKtpsFI6_2),.clk(gclk));
	jdff dff_B_htM14mEC7_2(.din(w_dff_B_9jKtpsFI6_2),.dout(w_dff_B_htM14mEC7_2),.clk(gclk));
	jdff dff_B_n9F98El57_2(.din(w_dff_B_htM14mEC7_2),.dout(w_dff_B_n9F98El57_2),.clk(gclk));
	jdff dff_B_xoMEQcR57_2(.din(w_dff_B_n9F98El57_2),.dout(w_dff_B_xoMEQcR57_2),.clk(gclk));
	jdff dff_B_WNos43pr2_2(.din(w_dff_B_xoMEQcR57_2),.dout(w_dff_B_WNos43pr2_2),.clk(gclk));
	jdff dff_B_Mh1PnJ7f7_2(.din(w_dff_B_WNos43pr2_2),.dout(w_dff_B_Mh1PnJ7f7_2),.clk(gclk));
	jdff dff_B_RpQVY65J4_2(.din(w_dff_B_Mh1PnJ7f7_2),.dout(w_dff_B_RpQVY65J4_2),.clk(gclk));
	jdff dff_B_93VvMLb58_2(.din(w_dff_B_RpQVY65J4_2),.dout(w_dff_B_93VvMLb58_2),.clk(gclk));
	jdff dff_B_ZQYaCXxO8_2(.din(w_dff_B_93VvMLb58_2),.dout(w_dff_B_ZQYaCXxO8_2),.clk(gclk));
	jdff dff_B_t3EzFkF37_2(.din(w_dff_B_ZQYaCXxO8_2),.dout(w_dff_B_t3EzFkF37_2),.clk(gclk));
	jdff dff_B_K25tA2PS5_2(.din(w_dff_B_t3EzFkF37_2),.dout(w_dff_B_K25tA2PS5_2),.clk(gclk));
	jdff dff_B_zWRsC3bq5_2(.din(w_dff_B_K25tA2PS5_2),.dout(w_dff_B_zWRsC3bq5_2),.clk(gclk));
	jdff dff_B_7cyJ4ttE1_2(.din(w_dff_B_zWRsC3bq5_2),.dout(w_dff_B_7cyJ4ttE1_2),.clk(gclk));
	jdff dff_B_d0ojW1mo2_2(.din(w_dff_B_7cyJ4ttE1_2),.dout(w_dff_B_d0ojW1mo2_2),.clk(gclk));
	jdff dff_B_w4yjCdvI7_2(.din(w_dff_B_d0ojW1mo2_2),.dout(w_dff_B_w4yjCdvI7_2),.clk(gclk));
	jdff dff_B_6c103qEE8_2(.din(w_dff_B_w4yjCdvI7_2),.dout(w_dff_B_6c103qEE8_2),.clk(gclk));
	jdff dff_B_Hmw166ZA9_2(.din(w_dff_B_6c103qEE8_2),.dout(w_dff_B_Hmw166ZA9_2),.clk(gclk));
	jdff dff_B_Q768gosW6_2(.din(w_dff_B_Hmw166ZA9_2),.dout(w_dff_B_Q768gosW6_2),.clk(gclk));
	jdff dff_B_bxhmf6Jn1_2(.din(w_dff_B_Q768gosW6_2),.dout(w_dff_B_bxhmf6Jn1_2),.clk(gclk));
	jdff dff_B_mR8i586u6_2(.din(w_dff_B_bxhmf6Jn1_2),.dout(w_dff_B_mR8i586u6_2),.clk(gclk));
	jdff dff_B_hbex8qap6_2(.din(w_dff_B_mR8i586u6_2),.dout(w_dff_B_hbex8qap6_2),.clk(gclk));
	jdff dff_B_4AVorcFG1_2(.din(w_dff_B_hbex8qap6_2),.dout(w_dff_B_4AVorcFG1_2),.clk(gclk));
	jdff dff_B_eriIFOdA8_2(.din(w_dff_B_4AVorcFG1_2),.dout(w_dff_B_eriIFOdA8_2),.clk(gclk));
	jdff dff_B_ZYR8bUcq9_1(.din(n1442),.dout(w_dff_B_ZYR8bUcq9_1),.clk(gclk));
	jdff dff_B_4ssvc3ki2_2(.din(n1363),.dout(w_dff_B_4ssvc3ki2_2),.clk(gclk));
	jdff dff_B_kDp4w20w5_2(.din(w_dff_B_4ssvc3ki2_2),.dout(w_dff_B_kDp4w20w5_2),.clk(gclk));
	jdff dff_B_rbm0nJuE1_2(.din(w_dff_B_kDp4w20w5_2),.dout(w_dff_B_rbm0nJuE1_2),.clk(gclk));
	jdff dff_B_CRhPGjLx1_2(.din(w_dff_B_rbm0nJuE1_2),.dout(w_dff_B_CRhPGjLx1_2),.clk(gclk));
	jdff dff_B_VR0TY0En9_2(.din(w_dff_B_CRhPGjLx1_2),.dout(w_dff_B_VR0TY0En9_2),.clk(gclk));
	jdff dff_B_w7067A6k8_2(.din(w_dff_B_VR0TY0En9_2),.dout(w_dff_B_w7067A6k8_2),.clk(gclk));
	jdff dff_B_ublLwUk06_2(.din(w_dff_B_w7067A6k8_2),.dout(w_dff_B_ublLwUk06_2),.clk(gclk));
	jdff dff_B_ONZshlIA3_2(.din(w_dff_B_ublLwUk06_2),.dout(w_dff_B_ONZshlIA3_2),.clk(gclk));
	jdff dff_B_vS4z9xBE7_2(.din(w_dff_B_ONZshlIA3_2),.dout(w_dff_B_vS4z9xBE7_2),.clk(gclk));
	jdff dff_B_RZGrnvTw7_2(.din(w_dff_B_vS4z9xBE7_2),.dout(w_dff_B_RZGrnvTw7_2),.clk(gclk));
	jdff dff_B_4LIAl3iU5_2(.din(w_dff_B_RZGrnvTw7_2),.dout(w_dff_B_4LIAl3iU5_2),.clk(gclk));
	jdff dff_B_iVirvHAg5_2(.din(w_dff_B_4LIAl3iU5_2),.dout(w_dff_B_iVirvHAg5_2),.clk(gclk));
	jdff dff_B_tZsvH4Io2_2(.din(w_dff_B_iVirvHAg5_2),.dout(w_dff_B_tZsvH4Io2_2),.clk(gclk));
	jdff dff_B_9ucynOSd9_2(.din(w_dff_B_tZsvH4Io2_2),.dout(w_dff_B_9ucynOSd9_2),.clk(gclk));
	jdff dff_B_N5DiDxSP7_2(.din(w_dff_B_9ucynOSd9_2),.dout(w_dff_B_N5DiDxSP7_2),.clk(gclk));
	jdff dff_B_5BWeoAYm9_2(.din(w_dff_B_N5DiDxSP7_2),.dout(w_dff_B_5BWeoAYm9_2),.clk(gclk));
	jdff dff_B_ZHtrGXRZ0_2(.din(w_dff_B_5BWeoAYm9_2),.dout(w_dff_B_ZHtrGXRZ0_2),.clk(gclk));
	jdff dff_B_hIsLXNHo6_2(.din(w_dff_B_ZHtrGXRZ0_2),.dout(w_dff_B_hIsLXNHo6_2),.clk(gclk));
	jdff dff_B_Vh3Zg9Df7_2(.din(w_dff_B_hIsLXNHo6_2),.dout(w_dff_B_Vh3Zg9Df7_2),.clk(gclk));
	jdff dff_B_CLMI8uF79_2(.din(w_dff_B_Vh3Zg9Df7_2),.dout(w_dff_B_CLMI8uF79_2),.clk(gclk));
	jdff dff_B_L1Qd1uLb3_2(.din(w_dff_B_CLMI8uF79_2),.dout(w_dff_B_L1Qd1uLb3_2),.clk(gclk));
	jdff dff_B_IQcUPQV88_2(.din(w_dff_B_L1Qd1uLb3_2),.dout(w_dff_B_IQcUPQV88_2),.clk(gclk));
	jdff dff_B_bpggpXnK0_2(.din(w_dff_B_IQcUPQV88_2),.dout(w_dff_B_bpggpXnK0_2),.clk(gclk));
	jdff dff_B_yfeROOuA0_2(.din(w_dff_B_bpggpXnK0_2),.dout(w_dff_B_yfeROOuA0_2),.clk(gclk));
	jdff dff_B_gn6fMtlZ4_2(.din(w_dff_B_yfeROOuA0_2),.dout(w_dff_B_gn6fMtlZ4_2),.clk(gclk));
	jdff dff_B_KvxMmyCb4_2(.din(w_dff_B_gn6fMtlZ4_2),.dout(w_dff_B_KvxMmyCb4_2),.clk(gclk));
	jdff dff_B_sOps9xw27_2(.din(w_dff_B_KvxMmyCb4_2),.dout(w_dff_B_sOps9xw27_2),.clk(gclk));
	jdff dff_B_q8M89MVA6_2(.din(w_dff_B_sOps9xw27_2),.dout(w_dff_B_q8M89MVA6_2),.clk(gclk));
	jdff dff_B_9btL855A4_2(.din(w_dff_B_q8M89MVA6_2),.dout(w_dff_B_9btL855A4_2),.clk(gclk));
	jdff dff_B_7yT6s86O9_2(.din(w_dff_B_9btL855A4_2),.dout(w_dff_B_7yT6s86O9_2),.clk(gclk));
	jdff dff_B_N7HFNmL51_2(.din(n1395),.dout(w_dff_B_N7HFNmL51_2),.clk(gclk));
	jdff dff_B_3PqYq3sP3_1(.din(n1364),.dout(w_dff_B_3PqYq3sP3_1),.clk(gclk));
	jdff dff_B_OtXlyWkF9_2(.din(n1278),.dout(w_dff_B_OtXlyWkF9_2),.clk(gclk));
	jdff dff_B_MZJd5AlY4_2(.din(w_dff_B_OtXlyWkF9_2),.dout(w_dff_B_MZJd5AlY4_2),.clk(gclk));
	jdff dff_B_qM1O2MMg5_2(.din(w_dff_B_MZJd5AlY4_2),.dout(w_dff_B_qM1O2MMg5_2),.clk(gclk));
	jdff dff_B_XL6K4SKI0_2(.din(w_dff_B_qM1O2MMg5_2),.dout(w_dff_B_XL6K4SKI0_2),.clk(gclk));
	jdff dff_B_nPak7Bnr0_2(.din(w_dff_B_XL6K4SKI0_2),.dout(w_dff_B_nPak7Bnr0_2),.clk(gclk));
	jdff dff_B_6CFPvWJB5_2(.din(w_dff_B_nPak7Bnr0_2),.dout(w_dff_B_6CFPvWJB5_2),.clk(gclk));
	jdff dff_B_iVhXdDKL5_2(.din(w_dff_B_6CFPvWJB5_2),.dout(w_dff_B_iVhXdDKL5_2),.clk(gclk));
	jdff dff_B_K7NKydnj0_2(.din(w_dff_B_iVhXdDKL5_2),.dout(w_dff_B_K7NKydnj0_2),.clk(gclk));
	jdff dff_B_AGFIL2cr7_2(.din(w_dff_B_K7NKydnj0_2),.dout(w_dff_B_AGFIL2cr7_2),.clk(gclk));
	jdff dff_B_WUVTxoag8_2(.din(w_dff_B_AGFIL2cr7_2),.dout(w_dff_B_WUVTxoag8_2),.clk(gclk));
	jdff dff_B_Qmh1s1rS4_2(.din(w_dff_B_WUVTxoag8_2),.dout(w_dff_B_Qmh1s1rS4_2),.clk(gclk));
	jdff dff_B_hhUp20oT9_2(.din(w_dff_B_Qmh1s1rS4_2),.dout(w_dff_B_hhUp20oT9_2),.clk(gclk));
	jdff dff_B_SjsIbhE67_2(.din(w_dff_B_hhUp20oT9_2),.dout(w_dff_B_SjsIbhE67_2),.clk(gclk));
	jdff dff_B_0RFOmsFX8_2(.din(w_dff_B_SjsIbhE67_2),.dout(w_dff_B_0RFOmsFX8_2),.clk(gclk));
	jdff dff_B_vYHVJ21a4_2(.din(w_dff_B_0RFOmsFX8_2),.dout(w_dff_B_vYHVJ21a4_2),.clk(gclk));
	jdff dff_B_iWxfl3AW9_2(.din(w_dff_B_vYHVJ21a4_2),.dout(w_dff_B_iWxfl3AW9_2),.clk(gclk));
	jdff dff_B_noptbPDu7_2(.din(w_dff_B_iWxfl3AW9_2),.dout(w_dff_B_noptbPDu7_2),.clk(gclk));
	jdff dff_B_lAevw6P08_2(.din(w_dff_B_noptbPDu7_2),.dout(w_dff_B_lAevw6P08_2),.clk(gclk));
	jdff dff_B_ERzJiIhE7_2(.din(w_dff_B_lAevw6P08_2),.dout(w_dff_B_ERzJiIhE7_2),.clk(gclk));
	jdff dff_B_b1fEkFM42_2(.din(w_dff_B_ERzJiIhE7_2),.dout(w_dff_B_b1fEkFM42_2),.clk(gclk));
	jdff dff_B_jqWeuXVU8_2(.din(w_dff_B_b1fEkFM42_2),.dout(w_dff_B_jqWeuXVU8_2),.clk(gclk));
	jdff dff_B_xNkw5Xi87_2(.din(w_dff_B_jqWeuXVU8_2),.dout(w_dff_B_xNkw5Xi87_2),.clk(gclk));
	jdff dff_B_aZQysVSF8_2(.din(w_dff_B_xNkw5Xi87_2),.dout(w_dff_B_aZQysVSF8_2),.clk(gclk));
	jdff dff_B_N9BdXA5F1_2(.din(w_dff_B_aZQysVSF8_2),.dout(w_dff_B_N9BdXA5F1_2),.clk(gclk));
	jdff dff_B_cIzcRSxX1_2(.din(w_dff_B_N9BdXA5F1_2),.dout(w_dff_B_cIzcRSxX1_2),.clk(gclk));
	jdff dff_B_qAVhMp1z9_2(.din(w_dff_B_cIzcRSxX1_2),.dout(w_dff_B_qAVhMp1z9_2),.clk(gclk));
	jdff dff_B_rCZSACc71_2(.din(w_dff_B_qAVhMp1z9_2),.dout(w_dff_B_rCZSACc71_2),.clk(gclk));
	jdff dff_B_JzaWxUPK5_2(.din(n1310),.dout(w_dff_B_JzaWxUPK5_2),.clk(gclk));
	jdff dff_B_GEWdfR901_1(.din(n1279),.dout(w_dff_B_GEWdfR901_1),.clk(gclk));
	jdff dff_B_NjmbRh5y1_2(.din(n1188),.dout(w_dff_B_NjmbRh5y1_2),.clk(gclk));
	jdff dff_B_3TUKA2cL3_2(.din(w_dff_B_NjmbRh5y1_2),.dout(w_dff_B_3TUKA2cL3_2),.clk(gclk));
	jdff dff_B_tQRABHbm6_2(.din(w_dff_B_3TUKA2cL3_2),.dout(w_dff_B_tQRABHbm6_2),.clk(gclk));
	jdff dff_B_TWULv2pj6_2(.din(w_dff_B_tQRABHbm6_2),.dout(w_dff_B_TWULv2pj6_2),.clk(gclk));
	jdff dff_B_Zlz2yOhk7_2(.din(w_dff_B_TWULv2pj6_2),.dout(w_dff_B_Zlz2yOhk7_2),.clk(gclk));
	jdff dff_B_v6HjMCBG8_2(.din(w_dff_B_Zlz2yOhk7_2),.dout(w_dff_B_v6HjMCBG8_2),.clk(gclk));
	jdff dff_B_AgvHnm2u6_2(.din(w_dff_B_v6HjMCBG8_2),.dout(w_dff_B_AgvHnm2u6_2),.clk(gclk));
	jdff dff_B_K0LGHv5S3_2(.din(w_dff_B_AgvHnm2u6_2),.dout(w_dff_B_K0LGHv5S3_2),.clk(gclk));
	jdff dff_B_tfnngBfj8_2(.din(w_dff_B_K0LGHv5S3_2),.dout(w_dff_B_tfnngBfj8_2),.clk(gclk));
	jdff dff_B_FZfGiIqE5_2(.din(w_dff_B_tfnngBfj8_2),.dout(w_dff_B_FZfGiIqE5_2),.clk(gclk));
	jdff dff_B_H9JVhHAc0_2(.din(w_dff_B_FZfGiIqE5_2),.dout(w_dff_B_H9JVhHAc0_2),.clk(gclk));
	jdff dff_B_MHKDtimG9_2(.din(w_dff_B_H9JVhHAc0_2),.dout(w_dff_B_MHKDtimG9_2),.clk(gclk));
	jdff dff_B_59xidWHp8_2(.din(w_dff_B_MHKDtimG9_2),.dout(w_dff_B_59xidWHp8_2),.clk(gclk));
	jdff dff_B_zIisVie89_2(.din(w_dff_B_59xidWHp8_2),.dout(w_dff_B_zIisVie89_2),.clk(gclk));
	jdff dff_B_WmJUN1np3_2(.din(w_dff_B_zIisVie89_2),.dout(w_dff_B_WmJUN1np3_2),.clk(gclk));
	jdff dff_B_WgULM6H93_2(.din(w_dff_B_WmJUN1np3_2),.dout(w_dff_B_WgULM6H93_2),.clk(gclk));
	jdff dff_B_fedn4pvG9_2(.din(w_dff_B_WgULM6H93_2),.dout(w_dff_B_fedn4pvG9_2),.clk(gclk));
	jdff dff_B_BOXrLKuW2_2(.din(w_dff_B_fedn4pvG9_2),.dout(w_dff_B_BOXrLKuW2_2),.clk(gclk));
	jdff dff_B_uvlFfCrR9_2(.din(w_dff_B_BOXrLKuW2_2),.dout(w_dff_B_uvlFfCrR9_2),.clk(gclk));
	jdff dff_B_gSqHp4Qn3_2(.din(w_dff_B_uvlFfCrR9_2),.dout(w_dff_B_gSqHp4Qn3_2),.clk(gclk));
	jdff dff_B_9tzzqx2D9_2(.din(w_dff_B_gSqHp4Qn3_2),.dout(w_dff_B_9tzzqx2D9_2),.clk(gclk));
	jdff dff_B_PfRVapns3_2(.din(w_dff_B_9tzzqx2D9_2),.dout(w_dff_B_PfRVapns3_2),.clk(gclk));
	jdff dff_B_QBrN1hbE8_2(.din(w_dff_B_PfRVapns3_2),.dout(w_dff_B_QBrN1hbE8_2),.clk(gclk));
	jdff dff_B_OX7pxmD05_2(.din(w_dff_B_QBrN1hbE8_2),.dout(w_dff_B_OX7pxmD05_2),.clk(gclk));
	jdff dff_B_D9ufeY0w9_2(.din(n1219),.dout(w_dff_B_D9ufeY0w9_2),.clk(gclk));
	jdff dff_B_OGayP6UF0_1(.din(n1189),.dout(w_dff_B_OGayP6UF0_1),.clk(gclk));
	jdff dff_B_pPoq0s3E5_2(.din(n1084),.dout(w_dff_B_pPoq0s3E5_2),.clk(gclk));
	jdff dff_B_7YDyOhI02_2(.din(w_dff_B_pPoq0s3E5_2),.dout(w_dff_B_7YDyOhI02_2),.clk(gclk));
	jdff dff_B_Mgyzczwn7_2(.din(w_dff_B_7YDyOhI02_2),.dout(w_dff_B_Mgyzczwn7_2),.clk(gclk));
	jdff dff_B_WptxvJo90_2(.din(w_dff_B_Mgyzczwn7_2),.dout(w_dff_B_WptxvJo90_2),.clk(gclk));
	jdff dff_B_Z5oEdZZJ9_2(.din(w_dff_B_WptxvJo90_2),.dout(w_dff_B_Z5oEdZZJ9_2),.clk(gclk));
	jdff dff_B_CiRB4mgs6_2(.din(w_dff_B_Z5oEdZZJ9_2),.dout(w_dff_B_CiRB4mgs6_2),.clk(gclk));
	jdff dff_B_UyNeCXGl9_2(.din(w_dff_B_CiRB4mgs6_2),.dout(w_dff_B_UyNeCXGl9_2),.clk(gclk));
	jdff dff_B_LQ7cMm0f9_2(.din(w_dff_B_UyNeCXGl9_2),.dout(w_dff_B_LQ7cMm0f9_2),.clk(gclk));
	jdff dff_B_CGHJPGSj3_2(.din(w_dff_B_LQ7cMm0f9_2),.dout(w_dff_B_CGHJPGSj3_2),.clk(gclk));
	jdff dff_B_mhRCrGfW5_2(.din(w_dff_B_CGHJPGSj3_2),.dout(w_dff_B_mhRCrGfW5_2),.clk(gclk));
	jdff dff_B_3nlWnsGa8_2(.din(w_dff_B_mhRCrGfW5_2),.dout(w_dff_B_3nlWnsGa8_2),.clk(gclk));
	jdff dff_B_Pkf2jpEu2_2(.din(w_dff_B_3nlWnsGa8_2),.dout(w_dff_B_Pkf2jpEu2_2),.clk(gclk));
	jdff dff_B_Y4zq1sGt3_2(.din(w_dff_B_Pkf2jpEu2_2),.dout(w_dff_B_Y4zq1sGt3_2),.clk(gclk));
	jdff dff_B_Yw5WNjbN2_2(.din(w_dff_B_Y4zq1sGt3_2),.dout(w_dff_B_Yw5WNjbN2_2),.clk(gclk));
	jdff dff_B_TtLTdCew5_2(.din(w_dff_B_Yw5WNjbN2_2),.dout(w_dff_B_TtLTdCew5_2),.clk(gclk));
	jdff dff_B_2I0LAd8o8_2(.din(w_dff_B_TtLTdCew5_2),.dout(w_dff_B_2I0LAd8o8_2),.clk(gclk));
	jdff dff_B_5wyvDAza6_2(.din(w_dff_B_2I0LAd8o8_2),.dout(w_dff_B_5wyvDAza6_2),.clk(gclk));
	jdff dff_B_CASYQ0eH7_2(.din(w_dff_B_5wyvDAza6_2),.dout(w_dff_B_CASYQ0eH7_2),.clk(gclk));
	jdff dff_B_5WBTIYFa4_2(.din(w_dff_B_CASYQ0eH7_2),.dout(w_dff_B_5WBTIYFa4_2),.clk(gclk));
	jdff dff_B_BxoRNNht1_2(.din(w_dff_B_5WBTIYFa4_2),.dout(w_dff_B_BxoRNNht1_2),.clk(gclk));
	jdff dff_B_7bZcCXZS1_2(.din(w_dff_B_BxoRNNht1_2),.dout(w_dff_B_7bZcCXZS1_2),.clk(gclk));
	jdff dff_B_GbmpGLAX9_2(.din(n1121),.dout(w_dff_B_GbmpGLAX9_2),.clk(gclk));
	jdff dff_B_gCRseKSX3_1(.din(n1085),.dout(w_dff_B_gCRseKSX3_1),.clk(gclk));
	jdff dff_B_mlDj4PGA0_2(.din(n986),.dout(w_dff_B_mlDj4PGA0_2),.clk(gclk));
	jdff dff_B_60JDDtxq8_2(.din(w_dff_B_mlDj4PGA0_2),.dout(w_dff_B_60JDDtxq8_2),.clk(gclk));
	jdff dff_B_dXKPNGaB6_2(.din(w_dff_B_60JDDtxq8_2),.dout(w_dff_B_dXKPNGaB6_2),.clk(gclk));
	jdff dff_B_BcmT4in45_2(.din(w_dff_B_dXKPNGaB6_2),.dout(w_dff_B_BcmT4in45_2),.clk(gclk));
	jdff dff_B_nXsgOr2e6_2(.din(w_dff_B_BcmT4in45_2),.dout(w_dff_B_nXsgOr2e6_2),.clk(gclk));
	jdff dff_B_b3xcDoic3_2(.din(w_dff_B_nXsgOr2e6_2),.dout(w_dff_B_b3xcDoic3_2),.clk(gclk));
	jdff dff_B_85kXD39g6_2(.din(w_dff_B_b3xcDoic3_2),.dout(w_dff_B_85kXD39g6_2),.clk(gclk));
	jdff dff_B_TDjDuefu0_2(.din(w_dff_B_85kXD39g6_2),.dout(w_dff_B_TDjDuefu0_2),.clk(gclk));
	jdff dff_B_GkPCBVRA0_2(.din(w_dff_B_TDjDuefu0_2),.dout(w_dff_B_GkPCBVRA0_2),.clk(gclk));
	jdff dff_B_k7XBf9yh1_2(.din(w_dff_B_GkPCBVRA0_2),.dout(w_dff_B_k7XBf9yh1_2),.clk(gclk));
	jdff dff_B_KLP56cjr7_2(.din(w_dff_B_k7XBf9yh1_2),.dout(w_dff_B_KLP56cjr7_2),.clk(gclk));
	jdff dff_B_QoIdJcCd5_2(.din(w_dff_B_KLP56cjr7_2),.dout(w_dff_B_QoIdJcCd5_2),.clk(gclk));
	jdff dff_B_d6bmIbUv2_2(.din(w_dff_B_QoIdJcCd5_2),.dout(w_dff_B_d6bmIbUv2_2),.clk(gclk));
	jdff dff_B_mqnz2Oec4_2(.din(w_dff_B_d6bmIbUv2_2),.dout(w_dff_B_mqnz2Oec4_2),.clk(gclk));
	jdff dff_B_NczUmfie4_2(.din(w_dff_B_mqnz2Oec4_2),.dout(w_dff_B_NczUmfie4_2),.clk(gclk));
	jdff dff_B_ScNqzfOL9_2(.din(w_dff_B_NczUmfie4_2),.dout(w_dff_B_ScNqzfOL9_2),.clk(gclk));
	jdff dff_B_4mkaHuoa0_2(.din(w_dff_B_ScNqzfOL9_2),.dout(w_dff_B_4mkaHuoa0_2),.clk(gclk));
	jdff dff_B_SYNboMum6_2(.din(w_dff_B_4mkaHuoa0_2),.dout(w_dff_B_SYNboMum6_2),.clk(gclk));
	jdff dff_B_xixEthtw6_2(.din(n1016),.dout(w_dff_B_xixEthtw6_2),.clk(gclk));
	jdff dff_B_qeu9lj3P5_1(.din(n987),.dout(w_dff_B_qeu9lj3P5_1),.clk(gclk));
	jdff dff_B_HmnumnpZ7_2(.din(n881),.dout(w_dff_B_HmnumnpZ7_2),.clk(gclk));
	jdff dff_B_sOrVGgvY5_2(.din(w_dff_B_HmnumnpZ7_2),.dout(w_dff_B_sOrVGgvY5_2),.clk(gclk));
	jdff dff_B_iEXFjpRo6_2(.din(w_dff_B_sOrVGgvY5_2),.dout(w_dff_B_iEXFjpRo6_2),.clk(gclk));
	jdff dff_B_2GYSVV2G5_2(.din(w_dff_B_iEXFjpRo6_2),.dout(w_dff_B_2GYSVV2G5_2),.clk(gclk));
	jdff dff_B_eojb1KFr7_2(.din(w_dff_B_2GYSVV2G5_2),.dout(w_dff_B_eojb1KFr7_2),.clk(gclk));
	jdff dff_B_w2CaxaxL6_2(.din(w_dff_B_eojb1KFr7_2),.dout(w_dff_B_w2CaxaxL6_2),.clk(gclk));
	jdff dff_B_fvZqbBQc7_2(.din(w_dff_B_w2CaxaxL6_2),.dout(w_dff_B_fvZqbBQc7_2),.clk(gclk));
	jdff dff_B_4pObe9bz1_2(.din(w_dff_B_fvZqbBQc7_2),.dout(w_dff_B_4pObe9bz1_2),.clk(gclk));
	jdff dff_B_yyPU1AZ42_2(.din(w_dff_B_4pObe9bz1_2),.dout(w_dff_B_yyPU1AZ42_2),.clk(gclk));
	jdff dff_B_rDT0YzAj1_2(.din(w_dff_B_yyPU1AZ42_2),.dout(w_dff_B_rDT0YzAj1_2),.clk(gclk));
	jdff dff_B_3nyNm6ik4_2(.din(w_dff_B_rDT0YzAj1_2),.dout(w_dff_B_3nyNm6ik4_2),.clk(gclk));
	jdff dff_B_4VG4T8j56_2(.din(w_dff_B_3nyNm6ik4_2),.dout(w_dff_B_4VG4T8j56_2),.clk(gclk));
	jdff dff_B_oDQCTvP72_2(.din(w_dff_B_4VG4T8j56_2),.dout(w_dff_B_oDQCTvP72_2),.clk(gclk));
	jdff dff_B_jN30JHwD0_2(.din(w_dff_B_oDQCTvP72_2),.dout(w_dff_B_jN30JHwD0_2),.clk(gclk));
	jdff dff_B_hZonOQGc3_2(.din(w_dff_B_jN30JHwD0_2),.dout(w_dff_B_hZonOQGc3_2),.clk(gclk));
	jdff dff_B_VPqAJya48_2(.din(n911),.dout(w_dff_B_VPqAJya48_2),.clk(gclk));
	jdff dff_B_mzUSu3Sl6_1(.din(n882),.dout(w_dff_B_mzUSu3Sl6_1),.clk(gclk));
	jdff dff_B_U2zLMTSV7_2(.din(n782),.dout(w_dff_B_U2zLMTSV7_2),.clk(gclk));
	jdff dff_B_FKFziUga8_2(.din(w_dff_B_U2zLMTSV7_2),.dout(w_dff_B_FKFziUga8_2),.clk(gclk));
	jdff dff_B_VB0madkY1_2(.din(w_dff_B_FKFziUga8_2),.dout(w_dff_B_VB0madkY1_2),.clk(gclk));
	jdff dff_B_ndr0xpYE1_2(.din(w_dff_B_VB0madkY1_2),.dout(w_dff_B_ndr0xpYE1_2),.clk(gclk));
	jdff dff_B_esdRrUru9_2(.din(w_dff_B_ndr0xpYE1_2),.dout(w_dff_B_esdRrUru9_2),.clk(gclk));
	jdff dff_B_LaW8pPi32_2(.din(w_dff_B_esdRrUru9_2),.dout(w_dff_B_LaW8pPi32_2),.clk(gclk));
	jdff dff_B_R5w4YP2I5_2(.din(w_dff_B_LaW8pPi32_2),.dout(w_dff_B_R5w4YP2I5_2),.clk(gclk));
	jdff dff_B_cbGvOLHq5_2(.din(w_dff_B_R5w4YP2I5_2),.dout(w_dff_B_cbGvOLHq5_2),.clk(gclk));
	jdff dff_B_NcjOMpo80_2(.din(w_dff_B_cbGvOLHq5_2),.dout(w_dff_B_NcjOMpo80_2),.clk(gclk));
	jdff dff_B_rJhexsno1_2(.din(w_dff_B_NcjOMpo80_2),.dout(w_dff_B_rJhexsno1_2),.clk(gclk));
	jdff dff_B_lFlZ85i59_2(.din(w_dff_B_rJhexsno1_2),.dout(w_dff_B_lFlZ85i59_2),.clk(gclk));
	jdff dff_B_qZbZfeDP3_2(.din(w_dff_B_lFlZ85i59_2),.dout(w_dff_B_qZbZfeDP3_2),.clk(gclk));
	jdff dff_B_fwDr6czM6_2(.din(n805),.dout(w_dff_B_fwDr6czM6_2),.clk(gclk));
	jdff dff_B_5vWzdcRT7_1(.din(n783),.dout(w_dff_B_5vWzdcRT7_1),.clk(gclk));
	jdff dff_B_8LTdD9Av0_2(.din(n689),.dout(w_dff_B_8LTdD9Av0_2),.clk(gclk));
	jdff dff_B_az2n5Dvx8_2(.din(w_dff_B_8LTdD9Av0_2),.dout(w_dff_B_az2n5Dvx8_2),.clk(gclk));
	jdff dff_B_hLCyo4IY1_2(.din(w_dff_B_az2n5Dvx8_2),.dout(w_dff_B_hLCyo4IY1_2),.clk(gclk));
	jdff dff_B_KTHieP3o9_2(.din(w_dff_B_hLCyo4IY1_2),.dout(w_dff_B_KTHieP3o9_2),.clk(gclk));
	jdff dff_B_QJRV6pjR8_2(.din(w_dff_B_KTHieP3o9_2),.dout(w_dff_B_QJRV6pjR8_2),.clk(gclk));
	jdff dff_B_vYcwUBYG0_2(.din(w_dff_B_QJRV6pjR8_2),.dout(w_dff_B_vYcwUBYG0_2),.clk(gclk));
	jdff dff_B_zp5mS1ME4_2(.din(w_dff_B_vYcwUBYG0_2),.dout(w_dff_B_zp5mS1ME4_2),.clk(gclk));
	jdff dff_B_dVTQh3y36_2(.din(w_dff_B_zp5mS1ME4_2),.dout(w_dff_B_dVTQh3y36_2),.clk(gclk));
	jdff dff_B_kW0xO70A7_2(.din(w_dff_B_dVTQh3y36_2),.dout(w_dff_B_kW0xO70A7_2),.clk(gclk));
	jdff dff_B_Yft6KHAR0_2(.din(n705),.dout(w_dff_B_Yft6KHAR0_2),.clk(gclk));
	jdff dff_B_Q9usjkEE9_2(.din(w_dff_B_Yft6KHAR0_2),.dout(w_dff_B_Q9usjkEE9_2),.clk(gclk));
	jdff dff_B_uDBHMAkV3_1(.din(n690),.dout(w_dff_B_uDBHMAkV3_1),.clk(gclk));
	jdff dff_B_hw5kRXTC8_1(.din(w_dff_B_uDBHMAkV3_1),.dout(w_dff_B_hw5kRXTC8_1),.clk(gclk));
	jdff dff_B_xZ9luDGZ0_1(.din(w_dff_B_hw5kRXTC8_1),.dout(w_dff_B_xZ9luDGZ0_1),.clk(gclk));
	jdff dff_B_p6Xw8KO09_1(.din(w_dff_B_xZ9luDGZ0_1),.dout(w_dff_B_p6Xw8KO09_1),.clk(gclk));
	jdff dff_B_iU6lThHJ5_1(.din(w_dff_B_p6Xw8KO09_1),.dout(w_dff_B_iU6lThHJ5_1),.clk(gclk));
	jdff dff_B_zSBRfi7M7_1(.din(w_dff_B_iU6lThHJ5_1),.dout(w_dff_B_zSBRfi7M7_1),.clk(gclk));
	jdff dff_B_HDVF1MKI9_0(.din(n612),.dout(w_dff_B_HDVF1MKI9_0),.clk(gclk));
	jdff dff_B_EekNaYkb0_0(.din(w_dff_B_HDVF1MKI9_0),.dout(w_dff_B_EekNaYkb0_0),.clk(gclk));
	jdff dff_A_N1glNa8a6_0(.dout(w_n611_0[0]),.din(w_dff_A_N1glNa8a6_0),.clk(gclk));
	jdff dff_A_XdFrbmsi7_0(.dout(w_dff_A_N1glNa8a6_0),.din(w_dff_A_XdFrbmsi7_0),.clk(gclk));
	jdff dff_A_uWveNDfc0_0(.dout(w_dff_A_XdFrbmsi7_0),.din(w_dff_A_uWveNDfc0_0),.clk(gclk));
	jdff dff_B_8Jm3I2aR8_1(.din(n605),.dout(w_dff_B_8Jm3I2aR8_1),.clk(gclk));
	jdff dff_A_dGQ0nULC2_0(.dout(w_n523_0[0]),.din(w_dff_A_dGQ0nULC2_0),.clk(gclk));
	jdff dff_A_KSL9U9ae5_1(.dout(w_n523_0[1]),.din(w_dff_A_KSL9U9ae5_1),.clk(gclk));
	jdff dff_A_KSo3umKP5_1(.dout(w_dff_A_KSL9U9ae5_1),.din(w_dff_A_KSo3umKP5_1),.clk(gclk));
	jdff dff_A_Kw2ZnM0o7_1(.dout(w_n603_0[1]),.din(w_dff_A_Kw2ZnM0o7_1),.clk(gclk));
	jdff dff_A_dpJ3ydDa4_1(.dout(w_dff_A_Kw2ZnM0o7_1),.din(w_dff_A_dpJ3ydDa4_1),.clk(gclk));
	jdff dff_A_u14aLw1x1_1(.dout(w_dff_A_dpJ3ydDa4_1),.din(w_dff_A_u14aLw1x1_1),.clk(gclk));
	jdff dff_A_8HGtWYyN0_1(.dout(w_dff_A_u14aLw1x1_1),.din(w_dff_A_8HGtWYyN0_1),.clk(gclk));
	jdff dff_A_XiL1B0KF5_1(.dout(w_dff_A_8HGtWYyN0_1),.din(w_dff_A_XiL1B0KF5_1),.clk(gclk));
	jdff dff_A_zum0rnsQ5_1(.dout(w_dff_A_XiL1B0KF5_1),.din(w_dff_A_zum0rnsQ5_1),.clk(gclk));
	jdff dff_B_r5DeWLnr2_1(.din(n1793),.dout(w_dff_B_r5DeWLnr2_1),.clk(gclk));
	jdff dff_A_NXdfcoJP4_1(.dout(w_n1768_0[1]),.din(w_dff_A_NXdfcoJP4_1),.clk(gclk));
	jdff dff_B_GY0AmhZ59_1(.din(n1766),.dout(w_dff_B_GY0AmhZ59_1),.clk(gclk));
	jdff dff_B_ePK80bvI7_2(.din(n1730),.dout(w_dff_B_ePK80bvI7_2),.clk(gclk));
	jdff dff_B_cCfugXea4_2(.din(w_dff_B_ePK80bvI7_2),.dout(w_dff_B_cCfugXea4_2),.clk(gclk));
	jdff dff_B_HNzP4zuC9_2(.din(w_dff_B_cCfugXea4_2),.dout(w_dff_B_HNzP4zuC9_2),.clk(gclk));
	jdff dff_B_xLjwrGpg1_2(.din(w_dff_B_HNzP4zuC9_2),.dout(w_dff_B_xLjwrGpg1_2),.clk(gclk));
	jdff dff_B_nlfY0wlw1_2(.din(w_dff_B_xLjwrGpg1_2),.dout(w_dff_B_nlfY0wlw1_2),.clk(gclk));
	jdff dff_B_Pzt54vDd6_2(.din(w_dff_B_nlfY0wlw1_2),.dout(w_dff_B_Pzt54vDd6_2),.clk(gclk));
	jdff dff_B_x1sVaed98_2(.din(w_dff_B_Pzt54vDd6_2),.dout(w_dff_B_x1sVaed98_2),.clk(gclk));
	jdff dff_B_Ke4Ut6Fp8_2(.din(w_dff_B_x1sVaed98_2),.dout(w_dff_B_Ke4Ut6Fp8_2),.clk(gclk));
	jdff dff_B_qfNMeWtP7_2(.din(w_dff_B_Ke4Ut6Fp8_2),.dout(w_dff_B_qfNMeWtP7_2),.clk(gclk));
	jdff dff_B_fqWe8lct2_2(.din(w_dff_B_qfNMeWtP7_2),.dout(w_dff_B_fqWe8lct2_2),.clk(gclk));
	jdff dff_B_CuW57XJU7_2(.din(w_dff_B_fqWe8lct2_2),.dout(w_dff_B_CuW57XJU7_2),.clk(gclk));
	jdff dff_B_o0dZ6yOj0_2(.din(w_dff_B_CuW57XJU7_2),.dout(w_dff_B_o0dZ6yOj0_2),.clk(gclk));
	jdff dff_B_Nay2pum26_2(.din(w_dff_B_o0dZ6yOj0_2),.dout(w_dff_B_Nay2pum26_2),.clk(gclk));
	jdff dff_B_ANHQpEA33_2(.din(w_dff_B_Nay2pum26_2),.dout(w_dff_B_ANHQpEA33_2),.clk(gclk));
	jdff dff_B_IbVan7kt7_2(.din(w_dff_B_ANHQpEA33_2),.dout(w_dff_B_IbVan7kt7_2),.clk(gclk));
	jdff dff_B_HDABYoca9_2(.din(w_dff_B_IbVan7kt7_2),.dout(w_dff_B_HDABYoca9_2),.clk(gclk));
	jdff dff_B_I2vE2NPk8_2(.din(w_dff_B_HDABYoca9_2),.dout(w_dff_B_I2vE2NPk8_2),.clk(gclk));
	jdff dff_B_fZjbahRI0_2(.din(w_dff_B_I2vE2NPk8_2),.dout(w_dff_B_fZjbahRI0_2),.clk(gclk));
	jdff dff_B_6EEMmO5J1_2(.din(w_dff_B_fZjbahRI0_2),.dout(w_dff_B_6EEMmO5J1_2),.clk(gclk));
	jdff dff_B_NqDLBXqy3_2(.din(w_dff_B_6EEMmO5J1_2),.dout(w_dff_B_NqDLBXqy3_2),.clk(gclk));
	jdff dff_B_5iYD0Zbd8_2(.din(w_dff_B_NqDLBXqy3_2),.dout(w_dff_B_5iYD0Zbd8_2),.clk(gclk));
	jdff dff_B_u0fiProG1_2(.din(w_dff_B_5iYD0Zbd8_2),.dout(w_dff_B_u0fiProG1_2),.clk(gclk));
	jdff dff_B_i1p3lPvA3_2(.din(w_dff_B_u0fiProG1_2),.dout(w_dff_B_i1p3lPvA3_2),.clk(gclk));
	jdff dff_B_JxbbM03X2_2(.din(w_dff_B_i1p3lPvA3_2),.dout(w_dff_B_JxbbM03X2_2),.clk(gclk));
	jdff dff_B_jjbOOJty0_2(.din(w_dff_B_JxbbM03X2_2),.dout(w_dff_B_jjbOOJty0_2),.clk(gclk));
	jdff dff_B_LLxWuUlF7_2(.din(w_dff_B_jjbOOJty0_2),.dout(w_dff_B_LLxWuUlF7_2),.clk(gclk));
	jdff dff_B_DwzoH0JF1_2(.din(w_dff_B_LLxWuUlF7_2),.dout(w_dff_B_DwzoH0JF1_2),.clk(gclk));
	jdff dff_B_Ca5xTHUO0_2(.din(w_dff_B_DwzoH0JF1_2),.dout(w_dff_B_Ca5xTHUO0_2),.clk(gclk));
	jdff dff_B_m5J8wfJ60_2(.din(w_dff_B_Ca5xTHUO0_2),.dout(w_dff_B_m5J8wfJ60_2),.clk(gclk));
	jdff dff_B_iZnl4Rt58_2(.din(w_dff_B_m5J8wfJ60_2),.dout(w_dff_B_iZnl4Rt58_2),.clk(gclk));
	jdff dff_B_DGDq6EMk9_2(.din(w_dff_B_iZnl4Rt58_2),.dout(w_dff_B_DGDq6EMk9_2),.clk(gclk));
	jdff dff_B_hNRTvzt02_2(.din(w_dff_B_DGDq6EMk9_2),.dout(w_dff_B_hNRTvzt02_2),.clk(gclk));
	jdff dff_B_31xG7Nmt6_2(.din(w_dff_B_hNRTvzt02_2),.dout(w_dff_B_31xG7Nmt6_2),.clk(gclk));
	jdff dff_B_TQKvFGPy5_2(.din(w_dff_B_31xG7Nmt6_2),.dout(w_dff_B_TQKvFGPy5_2),.clk(gclk));
	jdff dff_B_KdSJ1KoX0_2(.din(w_dff_B_TQKvFGPy5_2),.dout(w_dff_B_KdSJ1KoX0_2),.clk(gclk));
	jdff dff_B_PzXFJFzi7_2(.din(w_dff_B_KdSJ1KoX0_2),.dout(w_dff_B_PzXFJFzi7_2),.clk(gclk));
	jdff dff_B_aGujVf8T0_2(.din(w_dff_B_PzXFJFzi7_2),.dout(w_dff_B_aGujVf8T0_2),.clk(gclk));
	jdff dff_B_VoPYT5206_2(.din(w_dff_B_aGujVf8T0_2),.dout(w_dff_B_VoPYT5206_2),.clk(gclk));
	jdff dff_B_ILRjO57R8_2(.din(w_dff_B_VoPYT5206_2),.dout(w_dff_B_ILRjO57R8_2),.clk(gclk));
	jdff dff_B_pw6AlegW4_2(.din(w_dff_B_ILRjO57R8_2),.dout(w_dff_B_pw6AlegW4_2),.clk(gclk));
	jdff dff_B_tbcR3mhi0_2(.din(w_dff_B_pw6AlegW4_2),.dout(w_dff_B_tbcR3mhi0_2),.clk(gclk));
	jdff dff_B_ocZ4SEGP9_2(.din(w_dff_B_tbcR3mhi0_2),.dout(w_dff_B_ocZ4SEGP9_2),.clk(gclk));
	jdff dff_B_TKwQSZXY8_2(.din(w_dff_B_ocZ4SEGP9_2),.dout(w_dff_B_TKwQSZXY8_2),.clk(gclk));
	jdff dff_B_MU1aIrer5_2(.din(w_dff_B_TKwQSZXY8_2),.dout(w_dff_B_MU1aIrer5_2),.clk(gclk));
	jdff dff_B_d2o0mNql3_2(.din(w_dff_B_MU1aIrer5_2),.dout(w_dff_B_d2o0mNql3_2),.clk(gclk));
	jdff dff_B_NOHnhdVs3_2(.din(w_dff_B_d2o0mNql3_2),.dout(w_dff_B_NOHnhdVs3_2),.clk(gclk));
	jdff dff_B_8q2A1Z6i4_2(.din(w_dff_B_NOHnhdVs3_2),.dout(w_dff_B_8q2A1Z6i4_2),.clk(gclk));
	jdff dff_B_4ZrVkaSV6_2(.din(w_dff_B_8q2A1Z6i4_2),.dout(w_dff_B_4ZrVkaSV6_2),.clk(gclk));
	jdff dff_B_lJgWZslt3_2(.din(w_dff_B_4ZrVkaSV6_2),.dout(w_dff_B_lJgWZslt3_2),.clk(gclk));
	jdff dff_B_DUsgVNnI2_2(.din(w_dff_B_lJgWZslt3_2),.dout(w_dff_B_DUsgVNnI2_2),.clk(gclk));
	jdff dff_B_9RcW6zgb1_2(.din(w_dff_B_DUsgVNnI2_2),.dout(w_dff_B_9RcW6zgb1_2),.clk(gclk));
	jdff dff_B_xqDSkUBz5_2(.din(n1733),.dout(w_dff_B_xqDSkUBz5_2),.clk(gclk));
	jdff dff_B_gNgsEzPQ0_1(.din(n1731),.dout(w_dff_B_gNgsEzPQ0_1),.clk(gclk));
	jdff dff_B_UeJy3oBG9_2(.din(n1689),.dout(w_dff_B_UeJy3oBG9_2),.clk(gclk));
	jdff dff_B_7S71IYYJ9_2(.din(w_dff_B_UeJy3oBG9_2),.dout(w_dff_B_7S71IYYJ9_2),.clk(gclk));
	jdff dff_B_RXNEyLjz0_2(.din(w_dff_B_7S71IYYJ9_2),.dout(w_dff_B_RXNEyLjz0_2),.clk(gclk));
	jdff dff_B_dvGNkrd43_2(.din(w_dff_B_RXNEyLjz0_2),.dout(w_dff_B_dvGNkrd43_2),.clk(gclk));
	jdff dff_B_dIE8lYaJ6_2(.din(w_dff_B_dvGNkrd43_2),.dout(w_dff_B_dIE8lYaJ6_2),.clk(gclk));
	jdff dff_B_7zSgs2rL9_2(.din(w_dff_B_dIE8lYaJ6_2),.dout(w_dff_B_7zSgs2rL9_2),.clk(gclk));
	jdff dff_B_AOYRtnH48_2(.din(w_dff_B_7zSgs2rL9_2),.dout(w_dff_B_AOYRtnH48_2),.clk(gclk));
	jdff dff_B_xVlfDaRu6_2(.din(w_dff_B_AOYRtnH48_2),.dout(w_dff_B_xVlfDaRu6_2),.clk(gclk));
	jdff dff_B_Q5Q2WDhV2_2(.din(w_dff_B_xVlfDaRu6_2),.dout(w_dff_B_Q5Q2WDhV2_2),.clk(gclk));
	jdff dff_B_IB18Sr8k6_2(.din(w_dff_B_Q5Q2WDhV2_2),.dout(w_dff_B_IB18Sr8k6_2),.clk(gclk));
	jdff dff_B_RofjhBv10_2(.din(w_dff_B_IB18Sr8k6_2),.dout(w_dff_B_RofjhBv10_2),.clk(gclk));
	jdff dff_B_Ejvc9xEw2_2(.din(w_dff_B_RofjhBv10_2),.dout(w_dff_B_Ejvc9xEw2_2),.clk(gclk));
	jdff dff_B_mWE9sFZR3_2(.din(w_dff_B_Ejvc9xEw2_2),.dout(w_dff_B_mWE9sFZR3_2),.clk(gclk));
	jdff dff_B_cYLcsKcj5_2(.din(w_dff_B_mWE9sFZR3_2),.dout(w_dff_B_cYLcsKcj5_2),.clk(gclk));
	jdff dff_B_6s16I7Nh2_2(.din(w_dff_B_cYLcsKcj5_2),.dout(w_dff_B_6s16I7Nh2_2),.clk(gclk));
	jdff dff_B_wLve7vrG2_2(.din(w_dff_B_6s16I7Nh2_2),.dout(w_dff_B_wLve7vrG2_2),.clk(gclk));
	jdff dff_B_QpVrswoV0_2(.din(w_dff_B_wLve7vrG2_2),.dout(w_dff_B_QpVrswoV0_2),.clk(gclk));
	jdff dff_B_FvWZoqPa6_2(.din(w_dff_B_QpVrswoV0_2),.dout(w_dff_B_FvWZoqPa6_2),.clk(gclk));
	jdff dff_B_PTLvPhbQ4_2(.din(w_dff_B_FvWZoqPa6_2),.dout(w_dff_B_PTLvPhbQ4_2),.clk(gclk));
	jdff dff_B_6h3tks1C3_2(.din(w_dff_B_PTLvPhbQ4_2),.dout(w_dff_B_6h3tks1C3_2),.clk(gclk));
	jdff dff_B_6MDofNqx3_2(.din(w_dff_B_6h3tks1C3_2),.dout(w_dff_B_6MDofNqx3_2),.clk(gclk));
	jdff dff_B_lvbNRr7F0_2(.din(w_dff_B_6MDofNqx3_2),.dout(w_dff_B_lvbNRr7F0_2),.clk(gclk));
	jdff dff_B_KhifAR572_2(.din(w_dff_B_lvbNRr7F0_2),.dout(w_dff_B_KhifAR572_2),.clk(gclk));
	jdff dff_B_pKmY9tj21_2(.din(w_dff_B_KhifAR572_2),.dout(w_dff_B_pKmY9tj21_2),.clk(gclk));
	jdff dff_B_HDS0TLWb8_2(.din(w_dff_B_pKmY9tj21_2),.dout(w_dff_B_HDS0TLWb8_2),.clk(gclk));
	jdff dff_B_SGCr3OSu3_2(.din(w_dff_B_HDS0TLWb8_2),.dout(w_dff_B_SGCr3OSu3_2),.clk(gclk));
	jdff dff_B_kZSg5kYB2_2(.din(w_dff_B_SGCr3OSu3_2),.dout(w_dff_B_kZSg5kYB2_2),.clk(gclk));
	jdff dff_B_bDech5iz6_2(.din(w_dff_B_kZSg5kYB2_2),.dout(w_dff_B_bDech5iz6_2),.clk(gclk));
	jdff dff_B_flcFECST9_2(.din(w_dff_B_bDech5iz6_2),.dout(w_dff_B_flcFECST9_2),.clk(gclk));
	jdff dff_B_F7zz0rJa6_2(.din(w_dff_B_flcFECST9_2),.dout(w_dff_B_F7zz0rJa6_2),.clk(gclk));
	jdff dff_B_oHMzqdI25_2(.din(w_dff_B_F7zz0rJa6_2),.dout(w_dff_B_oHMzqdI25_2),.clk(gclk));
	jdff dff_B_zEyIqyRd9_2(.din(w_dff_B_oHMzqdI25_2),.dout(w_dff_B_zEyIqyRd9_2),.clk(gclk));
	jdff dff_B_1LFhMdCH5_2(.din(w_dff_B_zEyIqyRd9_2),.dout(w_dff_B_1LFhMdCH5_2),.clk(gclk));
	jdff dff_B_udmTubbg5_2(.din(w_dff_B_1LFhMdCH5_2),.dout(w_dff_B_udmTubbg5_2),.clk(gclk));
	jdff dff_B_YLrErCGP1_2(.din(w_dff_B_udmTubbg5_2),.dout(w_dff_B_YLrErCGP1_2),.clk(gclk));
	jdff dff_B_XJFTwsvg8_2(.din(w_dff_B_YLrErCGP1_2),.dout(w_dff_B_XJFTwsvg8_2),.clk(gclk));
	jdff dff_B_qzN7AVFu1_2(.din(w_dff_B_XJFTwsvg8_2),.dout(w_dff_B_qzN7AVFu1_2),.clk(gclk));
	jdff dff_B_RHCQOPhW4_2(.din(w_dff_B_qzN7AVFu1_2),.dout(w_dff_B_RHCQOPhW4_2),.clk(gclk));
	jdff dff_B_4yo4dVHH8_2(.din(w_dff_B_RHCQOPhW4_2),.dout(w_dff_B_4yo4dVHH8_2),.clk(gclk));
	jdff dff_B_vSoP8dTC1_2(.din(w_dff_B_4yo4dVHH8_2),.dout(w_dff_B_vSoP8dTC1_2),.clk(gclk));
	jdff dff_B_3mftr2mb9_2(.din(w_dff_B_vSoP8dTC1_2),.dout(w_dff_B_3mftr2mb9_2),.clk(gclk));
	jdff dff_B_uV4YDR5P6_2(.din(w_dff_B_3mftr2mb9_2),.dout(w_dff_B_uV4YDR5P6_2),.clk(gclk));
	jdff dff_B_35pUyFmV2_2(.din(w_dff_B_uV4YDR5P6_2),.dout(w_dff_B_35pUyFmV2_2),.clk(gclk));
	jdff dff_B_oE49qvc90_2(.din(w_dff_B_35pUyFmV2_2),.dout(w_dff_B_oE49qvc90_2),.clk(gclk));
	jdff dff_B_HtFINoEQ4_2(.din(w_dff_B_oE49qvc90_2),.dout(w_dff_B_HtFINoEQ4_2),.clk(gclk));
	jdff dff_B_UJncnEO08_2(.din(w_dff_B_HtFINoEQ4_2),.dout(w_dff_B_UJncnEO08_2),.clk(gclk));
	jdff dff_B_r7iq2aZb3_2(.din(w_dff_B_UJncnEO08_2),.dout(w_dff_B_r7iq2aZb3_2),.clk(gclk));
	jdff dff_B_2HkC6nbC5_2(.din(n1692),.dout(w_dff_B_2HkC6nbC5_2),.clk(gclk));
	jdff dff_B_1mu5OWs52_1(.din(n1690),.dout(w_dff_B_1mu5OWs52_1),.clk(gclk));
	jdff dff_B_fx9haq3O3_2(.din(n1638),.dout(w_dff_B_fx9haq3O3_2),.clk(gclk));
	jdff dff_B_YfMA7yYg6_2(.din(w_dff_B_fx9haq3O3_2),.dout(w_dff_B_YfMA7yYg6_2),.clk(gclk));
	jdff dff_B_jztVFGoW9_2(.din(w_dff_B_YfMA7yYg6_2),.dout(w_dff_B_jztVFGoW9_2),.clk(gclk));
	jdff dff_B_UtV1uj8u9_2(.din(w_dff_B_jztVFGoW9_2),.dout(w_dff_B_UtV1uj8u9_2),.clk(gclk));
	jdff dff_B_ZebFH1Ax8_2(.din(w_dff_B_UtV1uj8u9_2),.dout(w_dff_B_ZebFH1Ax8_2),.clk(gclk));
	jdff dff_B_G50801TZ8_2(.din(w_dff_B_ZebFH1Ax8_2),.dout(w_dff_B_G50801TZ8_2),.clk(gclk));
	jdff dff_B_94tuSiRp4_2(.din(w_dff_B_G50801TZ8_2),.dout(w_dff_B_94tuSiRp4_2),.clk(gclk));
	jdff dff_B_TIMERHmp5_2(.din(w_dff_B_94tuSiRp4_2),.dout(w_dff_B_TIMERHmp5_2),.clk(gclk));
	jdff dff_B_Echx574a5_2(.din(w_dff_B_TIMERHmp5_2),.dout(w_dff_B_Echx574a5_2),.clk(gclk));
	jdff dff_B_tRKm64bN8_2(.din(w_dff_B_Echx574a5_2),.dout(w_dff_B_tRKm64bN8_2),.clk(gclk));
	jdff dff_B_ajetV92m8_2(.din(w_dff_B_tRKm64bN8_2),.dout(w_dff_B_ajetV92m8_2),.clk(gclk));
	jdff dff_B_5r6tFA737_2(.din(w_dff_B_ajetV92m8_2),.dout(w_dff_B_5r6tFA737_2),.clk(gclk));
	jdff dff_B_37MzKY7l3_2(.din(w_dff_B_5r6tFA737_2),.dout(w_dff_B_37MzKY7l3_2),.clk(gclk));
	jdff dff_B_V51WLoZA6_2(.din(w_dff_B_37MzKY7l3_2),.dout(w_dff_B_V51WLoZA6_2),.clk(gclk));
	jdff dff_B_Bk0ZjsuH0_2(.din(w_dff_B_V51WLoZA6_2),.dout(w_dff_B_Bk0ZjsuH0_2),.clk(gclk));
	jdff dff_B_vggDPlZB8_2(.din(w_dff_B_Bk0ZjsuH0_2),.dout(w_dff_B_vggDPlZB8_2),.clk(gclk));
	jdff dff_B_jrMZqvoa6_2(.din(w_dff_B_vggDPlZB8_2),.dout(w_dff_B_jrMZqvoa6_2),.clk(gclk));
	jdff dff_B_oZRJ3UTB2_2(.din(w_dff_B_jrMZqvoa6_2),.dout(w_dff_B_oZRJ3UTB2_2),.clk(gclk));
	jdff dff_B_8n0VR7Yz7_2(.din(w_dff_B_oZRJ3UTB2_2),.dout(w_dff_B_8n0VR7Yz7_2),.clk(gclk));
	jdff dff_B_mLwm33GN1_2(.din(w_dff_B_8n0VR7Yz7_2),.dout(w_dff_B_mLwm33GN1_2),.clk(gclk));
	jdff dff_B_EN0qF3oE4_2(.din(w_dff_B_mLwm33GN1_2),.dout(w_dff_B_EN0qF3oE4_2),.clk(gclk));
	jdff dff_B_rMNk3DzX1_2(.din(w_dff_B_EN0qF3oE4_2),.dout(w_dff_B_rMNk3DzX1_2),.clk(gclk));
	jdff dff_B_AF4cXdQd9_2(.din(w_dff_B_rMNk3DzX1_2),.dout(w_dff_B_AF4cXdQd9_2),.clk(gclk));
	jdff dff_B_XMVHqsc73_2(.din(w_dff_B_AF4cXdQd9_2),.dout(w_dff_B_XMVHqsc73_2),.clk(gclk));
	jdff dff_B_z1VVwp4Y0_2(.din(w_dff_B_XMVHqsc73_2),.dout(w_dff_B_z1VVwp4Y0_2),.clk(gclk));
	jdff dff_B_IIYiEoRg0_2(.din(w_dff_B_z1VVwp4Y0_2),.dout(w_dff_B_IIYiEoRg0_2),.clk(gclk));
	jdff dff_B_wb5hKJfC2_2(.din(w_dff_B_IIYiEoRg0_2),.dout(w_dff_B_wb5hKJfC2_2),.clk(gclk));
	jdff dff_B_3KyRdlSd7_2(.din(w_dff_B_wb5hKJfC2_2),.dout(w_dff_B_3KyRdlSd7_2),.clk(gclk));
	jdff dff_B_cEzJSqq35_2(.din(w_dff_B_3KyRdlSd7_2),.dout(w_dff_B_cEzJSqq35_2),.clk(gclk));
	jdff dff_B_tiFV97GI2_2(.din(w_dff_B_cEzJSqq35_2),.dout(w_dff_B_tiFV97GI2_2),.clk(gclk));
	jdff dff_B_59BGuEmy0_2(.din(w_dff_B_tiFV97GI2_2),.dout(w_dff_B_59BGuEmy0_2),.clk(gclk));
	jdff dff_B_tWUDG0Vs2_2(.din(w_dff_B_59BGuEmy0_2),.dout(w_dff_B_tWUDG0Vs2_2),.clk(gclk));
	jdff dff_B_UiR0cI807_2(.din(w_dff_B_tWUDG0Vs2_2),.dout(w_dff_B_UiR0cI807_2),.clk(gclk));
	jdff dff_B_08ESIBcq8_2(.din(w_dff_B_UiR0cI807_2),.dout(w_dff_B_08ESIBcq8_2),.clk(gclk));
	jdff dff_B_vAIYuKNk3_2(.din(w_dff_B_08ESIBcq8_2),.dout(w_dff_B_vAIYuKNk3_2),.clk(gclk));
	jdff dff_B_6AUDhgD76_2(.din(w_dff_B_vAIYuKNk3_2),.dout(w_dff_B_6AUDhgD76_2),.clk(gclk));
	jdff dff_B_4vd5f4yR0_2(.din(w_dff_B_6AUDhgD76_2),.dout(w_dff_B_4vd5f4yR0_2),.clk(gclk));
	jdff dff_B_oHs6fx5U7_2(.din(w_dff_B_4vd5f4yR0_2),.dout(w_dff_B_oHs6fx5U7_2),.clk(gclk));
	jdff dff_B_q7UVgjRl9_2(.din(w_dff_B_oHs6fx5U7_2),.dout(w_dff_B_q7UVgjRl9_2),.clk(gclk));
	jdff dff_B_aP3utOCb8_2(.din(w_dff_B_q7UVgjRl9_2),.dout(w_dff_B_aP3utOCb8_2),.clk(gclk));
	jdff dff_B_IzhBC1Of2_2(.din(w_dff_B_aP3utOCb8_2),.dout(w_dff_B_IzhBC1Of2_2),.clk(gclk));
	jdff dff_B_crzB92Gp2_2(.din(w_dff_B_IzhBC1Of2_2),.dout(w_dff_B_crzB92Gp2_2),.clk(gclk));
	jdff dff_B_TbklrleN4_2(.din(w_dff_B_crzB92Gp2_2),.dout(w_dff_B_TbklrleN4_2),.clk(gclk));
	jdff dff_B_wvGEp2xp2_2(.din(n1641),.dout(w_dff_B_wvGEp2xp2_2),.clk(gclk));
	jdff dff_B_A4pjQGCK7_1(.din(n1639),.dout(w_dff_B_A4pjQGCK7_1),.clk(gclk));
	jdff dff_B_FnXJUlif7_2(.din(n1581),.dout(w_dff_B_FnXJUlif7_2),.clk(gclk));
	jdff dff_B_u0Jv3aqi7_2(.din(w_dff_B_FnXJUlif7_2),.dout(w_dff_B_u0Jv3aqi7_2),.clk(gclk));
	jdff dff_B_b6lgS73J8_2(.din(w_dff_B_u0Jv3aqi7_2),.dout(w_dff_B_b6lgS73J8_2),.clk(gclk));
	jdff dff_B_AbhwuB7d4_2(.din(w_dff_B_b6lgS73J8_2),.dout(w_dff_B_AbhwuB7d4_2),.clk(gclk));
	jdff dff_B_W11WnIzr4_2(.din(w_dff_B_AbhwuB7d4_2),.dout(w_dff_B_W11WnIzr4_2),.clk(gclk));
	jdff dff_B_veHGK0tW9_2(.din(w_dff_B_W11WnIzr4_2),.dout(w_dff_B_veHGK0tW9_2),.clk(gclk));
	jdff dff_B_LCDF74L72_2(.din(w_dff_B_veHGK0tW9_2),.dout(w_dff_B_LCDF74L72_2),.clk(gclk));
	jdff dff_B_dWltNYjq9_2(.din(w_dff_B_LCDF74L72_2),.dout(w_dff_B_dWltNYjq9_2),.clk(gclk));
	jdff dff_B_3yihavyc2_2(.din(w_dff_B_dWltNYjq9_2),.dout(w_dff_B_3yihavyc2_2),.clk(gclk));
	jdff dff_B_f7VucrrQ7_2(.din(w_dff_B_3yihavyc2_2),.dout(w_dff_B_f7VucrrQ7_2),.clk(gclk));
	jdff dff_B_dPb9Go098_2(.din(w_dff_B_f7VucrrQ7_2),.dout(w_dff_B_dPb9Go098_2),.clk(gclk));
	jdff dff_B_xsBvHCo94_2(.din(w_dff_B_dPb9Go098_2),.dout(w_dff_B_xsBvHCo94_2),.clk(gclk));
	jdff dff_B_h0cos4mL5_2(.din(w_dff_B_xsBvHCo94_2),.dout(w_dff_B_h0cos4mL5_2),.clk(gclk));
	jdff dff_B_xIJW41TO3_2(.din(w_dff_B_h0cos4mL5_2),.dout(w_dff_B_xIJW41TO3_2),.clk(gclk));
	jdff dff_B_9rXEMFgp1_2(.din(w_dff_B_xIJW41TO3_2),.dout(w_dff_B_9rXEMFgp1_2),.clk(gclk));
	jdff dff_B_ZxEWPVTO8_2(.din(w_dff_B_9rXEMFgp1_2),.dout(w_dff_B_ZxEWPVTO8_2),.clk(gclk));
	jdff dff_B_46TE9PDf6_2(.din(w_dff_B_ZxEWPVTO8_2),.dout(w_dff_B_46TE9PDf6_2),.clk(gclk));
	jdff dff_B_kCQksZOY7_2(.din(w_dff_B_46TE9PDf6_2),.dout(w_dff_B_kCQksZOY7_2),.clk(gclk));
	jdff dff_B_yp6xNKAH8_2(.din(w_dff_B_kCQksZOY7_2),.dout(w_dff_B_yp6xNKAH8_2),.clk(gclk));
	jdff dff_B_Iz8mMGtd4_2(.din(w_dff_B_yp6xNKAH8_2),.dout(w_dff_B_Iz8mMGtd4_2),.clk(gclk));
	jdff dff_B_5CXB30p35_2(.din(w_dff_B_Iz8mMGtd4_2),.dout(w_dff_B_5CXB30p35_2),.clk(gclk));
	jdff dff_B_WFpXvUFk3_2(.din(w_dff_B_5CXB30p35_2),.dout(w_dff_B_WFpXvUFk3_2),.clk(gclk));
	jdff dff_B_LsTKBciX4_2(.din(w_dff_B_WFpXvUFk3_2),.dout(w_dff_B_LsTKBciX4_2),.clk(gclk));
	jdff dff_B_lxdCiglv5_2(.din(w_dff_B_LsTKBciX4_2),.dout(w_dff_B_lxdCiglv5_2),.clk(gclk));
	jdff dff_B_tUBomGYf4_2(.din(w_dff_B_lxdCiglv5_2),.dout(w_dff_B_tUBomGYf4_2),.clk(gclk));
	jdff dff_B_CDUf4V7V9_2(.din(w_dff_B_tUBomGYf4_2),.dout(w_dff_B_CDUf4V7V9_2),.clk(gclk));
	jdff dff_B_xObiIz8G8_2(.din(w_dff_B_CDUf4V7V9_2),.dout(w_dff_B_xObiIz8G8_2),.clk(gclk));
	jdff dff_B_xVzciGid0_2(.din(w_dff_B_xObiIz8G8_2),.dout(w_dff_B_xVzciGid0_2),.clk(gclk));
	jdff dff_B_MU6FulMD7_2(.din(w_dff_B_xVzciGid0_2),.dout(w_dff_B_MU6FulMD7_2),.clk(gclk));
	jdff dff_B_JNPVonrv8_2(.din(w_dff_B_MU6FulMD7_2),.dout(w_dff_B_JNPVonrv8_2),.clk(gclk));
	jdff dff_B_2bmkkxQE5_2(.din(w_dff_B_JNPVonrv8_2),.dout(w_dff_B_2bmkkxQE5_2),.clk(gclk));
	jdff dff_B_oXNII3Wb9_2(.din(w_dff_B_2bmkkxQE5_2),.dout(w_dff_B_oXNII3Wb9_2),.clk(gclk));
	jdff dff_B_783TQtc27_2(.din(w_dff_B_oXNII3Wb9_2),.dout(w_dff_B_783TQtc27_2),.clk(gclk));
	jdff dff_B_9fTZuK665_2(.din(w_dff_B_783TQtc27_2),.dout(w_dff_B_9fTZuK665_2),.clk(gclk));
	jdff dff_B_CB8uP2Fw9_2(.din(w_dff_B_9fTZuK665_2),.dout(w_dff_B_CB8uP2Fw9_2),.clk(gclk));
	jdff dff_B_1ldaiBDb7_2(.din(w_dff_B_CB8uP2Fw9_2),.dout(w_dff_B_1ldaiBDb7_2),.clk(gclk));
	jdff dff_B_PkKDIW489_2(.din(w_dff_B_1ldaiBDb7_2),.dout(w_dff_B_PkKDIW489_2),.clk(gclk));
	jdff dff_B_02l0st186_2(.din(w_dff_B_PkKDIW489_2),.dout(w_dff_B_02l0st186_2),.clk(gclk));
	jdff dff_B_Vw0RU65l8_2(.din(w_dff_B_02l0st186_2),.dout(w_dff_B_Vw0RU65l8_2),.clk(gclk));
	jdff dff_B_V4twCLF92_2(.din(n1584),.dout(w_dff_B_V4twCLF92_2),.clk(gclk));
	jdff dff_B_Z7ZDwvJ80_1(.din(n1582),.dout(w_dff_B_Z7ZDwvJ80_1),.clk(gclk));
	jdff dff_B_woEOB4hB1_2(.din(n1517),.dout(w_dff_B_woEOB4hB1_2),.clk(gclk));
	jdff dff_B_mDLFQIFL5_2(.din(w_dff_B_woEOB4hB1_2),.dout(w_dff_B_mDLFQIFL5_2),.clk(gclk));
	jdff dff_B_dJ6203jA6_2(.din(w_dff_B_mDLFQIFL5_2),.dout(w_dff_B_dJ6203jA6_2),.clk(gclk));
	jdff dff_B_lKymu9Lv4_2(.din(w_dff_B_dJ6203jA6_2),.dout(w_dff_B_lKymu9Lv4_2),.clk(gclk));
	jdff dff_B_JPkCIFal8_2(.din(w_dff_B_lKymu9Lv4_2),.dout(w_dff_B_JPkCIFal8_2),.clk(gclk));
	jdff dff_B_DbfqoEeI1_2(.din(w_dff_B_JPkCIFal8_2),.dout(w_dff_B_DbfqoEeI1_2),.clk(gclk));
	jdff dff_B_U91YbclF1_2(.din(w_dff_B_DbfqoEeI1_2),.dout(w_dff_B_U91YbclF1_2),.clk(gclk));
	jdff dff_B_fXLij1Mx7_2(.din(w_dff_B_U91YbclF1_2),.dout(w_dff_B_fXLij1Mx7_2),.clk(gclk));
	jdff dff_B_qOOmlspL1_2(.din(w_dff_B_fXLij1Mx7_2),.dout(w_dff_B_qOOmlspL1_2),.clk(gclk));
	jdff dff_B_VlyAqOLq8_2(.din(w_dff_B_qOOmlspL1_2),.dout(w_dff_B_VlyAqOLq8_2),.clk(gclk));
	jdff dff_B_rE80ocvs4_2(.din(w_dff_B_VlyAqOLq8_2),.dout(w_dff_B_rE80ocvs4_2),.clk(gclk));
	jdff dff_B_RyLxkEpr5_2(.din(w_dff_B_rE80ocvs4_2),.dout(w_dff_B_RyLxkEpr5_2),.clk(gclk));
	jdff dff_B_xfO8Phnw0_2(.din(w_dff_B_RyLxkEpr5_2),.dout(w_dff_B_xfO8Phnw0_2),.clk(gclk));
	jdff dff_B_tm6IjM5W7_2(.din(w_dff_B_xfO8Phnw0_2),.dout(w_dff_B_tm6IjM5W7_2),.clk(gclk));
	jdff dff_B_joA427e71_2(.din(w_dff_B_tm6IjM5W7_2),.dout(w_dff_B_joA427e71_2),.clk(gclk));
	jdff dff_B_jtNb9Dqs1_2(.din(w_dff_B_joA427e71_2),.dout(w_dff_B_jtNb9Dqs1_2),.clk(gclk));
	jdff dff_B_d2Bicvdq8_2(.din(w_dff_B_jtNb9Dqs1_2),.dout(w_dff_B_d2Bicvdq8_2),.clk(gclk));
	jdff dff_B_Xy2KueEx5_2(.din(w_dff_B_d2Bicvdq8_2),.dout(w_dff_B_Xy2KueEx5_2),.clk(gclk));
	jdff dff_B_p5eCBVpM5_2(.din(w_dff_B_Xy2KueEx5_2),.dout(w_dff_B_p5eCBVpM5_2),.clk(gclk));
	jdff dff_B_8r2l9ORy4_2(.din(w_dff_B_p5eCBVpM5_2),.dout(w_dff_B_8r2l9ORy4_2),.clk(gclk));
	jdff dff_B_899Nl0u35_2(.din(w_dff_B_8r2l9ORy4_2),.dout(w_dff_B_899Nl0u35_2),.clk(gclk));
	jdff dff_B_Xskf7ANf0_2(.din(w_dff_B_899Nl0u35_2),.dout(w_dff_B_Xskf7ANf0_2),.clk(gclk));
	jdff dff_B_srHJoi8r6_2(.din(w_dff_B_Xskf7ANf0_2),.dout(w_dff_B_srHJoi8r6_2),.clk(gclk));
	jdff dff_B_XrxUk0ap3_2(.din(w_dff_B_srHJoi8r6_2),.dout(w_dff_B_XrxUk0ap3_2),.clk(gclk));
	jdff dff_B_8tBkrL922_2(.din(w_dff_B_XrxUk0ap3_2),.dout(w_dff_B_8tBkrL922_2),.clk(gclk));
	jdff dff_B_bNnqb7Ur8_2(.din(w_dff_B_8tBkrL922_2),.dout(w_dff_B_bNnqb7Ur8_2),.clk(gclk));
	jdff dff_B_dOpIcEEJ1_2(.din(w_dff_B_bNnqb7Ur8_2),.dout(w_dff_B_dOpIcEEJ1_2),.clk(gclk));
	jdff dff_B_3TquZD4L8_2(.din(w_dff_B_dOpIcEEJ1_2),.dout(w_dff_B_3TquZD4L8_2),.clk(gclk));
	jdff dff_B_uzVvRaG98_2(.din(w_dff_B_3TquZD4L8_2),.dout(w_dff_B_uzVvRaG98_2),.clk(gclk));
	jdff dff_B_I5PyVKJE5_2(.din(w_dff_B_uzVvRaG98_2),.dout(w_dff_B_I5PyVKJE5_2),.clk(gclk));
	jdff dff_B_V4WBCfy56_2(.din(w_dff_B_I5PyVKJE5_2),.dout(w_dff_B_V4WBCfy56_2),.clk(gclk));
	jdff dff_B_0PjtLUVy8_2(.din(w_dff_B_V4WBCfy56_2),.dout(w_dff_B_0PjtLUVy8_2),.clk(gclk));
	jdff dff_B_ddjO5ckY1_2(.din(w_dff_B_0PjtLUVy8_2),.dout(w_dff_B_ddjO5ckY1_2),.clk(gclk));
	jdff dff_B_ULlziK0B4_2(.din(w_dff_B_ddjO5ckY1_2),.dout(w_dff_B_ULlziK0B4_2),.clk(gclk));
	jdff dff_B_fKPvmQG84_2(.din(w_dff_B_ULlziK0B4_2),.dout(w_dff_B_fKPvmQG84_2),.clk(gclk));
	jdff dff_B_bkzLefRO7_2(.din(n1520),.dout(w_dff_B_bkzLefRO7_2),.clk(gclk));
	jdff dff_B_tB5h44mQ6_1(.din(n1518),.dout(w_dff_B_tB5h44mQ6_1),.clk(gclk));
	jdff dff_B_Y6Lt9qFR1_2(.din(n1446),.dout(w_dff_B_Y6Lt9qFR1_2),.clk(gclk));
	jdff dff_B_sdmIJJiy6_2(.din(w_dff_B_Y6Lt9qFR1_2),.dout(w_dff_B_sdmIJJiy6_2),.clk(gclk));
	jdff dff_B_e0JaXbkX8_2(.din(w_dff_B_sdmIJJiy6_2),.dout(w_dff_B_e0JaXbkX8_2),.clk(gclk));
	jdff dff_B_Z5IoM4KV9_2(.din(w_dff_B_e0JaXbkX8_2),.dout(w_dff_B_Z5IoM4KV9_2),.clk(gclk));
	jdff dff_B_l7b6rMQt2_2(.din(w_dff_B_Z5IoM4KV9_2),.dout(w_dff_B_l7b6rMQt2_2),.clk(gclk));
	jdff dff_B_VIi6iYqQ0_2(.din(w_dff_B_l7b6rMQt2_2),.dout(w_dff_B_VIi6iYqQ0_2),.clk(gclk));
	jdff dff_B_eQM7WvpS7_2(.din(w_dff_B_VIi6iYqQ0_2),.dout(w_dff_B_eQM7WvpS7_2),.clk(gclk));
	jdff dff_B_yFjIxuYn2_2(.din(w_dff_B_eQM7WvpS7_2),.dout(w_dff_B_yFjIxuYn2_2),.clk(gclk));
	jdff dff_B_uLFsrxjJ0_2(.din(w_dff_B_yFjIxuYn2_2),.dout(w_dff_B_uLFsrxjJ0_2),.clk(gclk));
	jdff dff_B_Nzz2xrKI9_2(.din(w_dff_B_uLFsrxjJ0_2),.dout(w_dff_B_Nzz2xrKI9_2),.clk(gclk));
	jdff dff_B_rto4OUmf2_2(.din(w_dff_B_Nzz2xrKI9_2),.dout(w_dff_B_rto4OUmf2_2),.clk(gclk));
	jdff dff_B_LB06HmON2_2(.din(w_dff_B_rto4OUmf2_2),.dout(w_dff_B_LB06HmON2_2),.clk(gclk));
	jdff dff_B_Ns69LjTy3_2(.din(w_dff_B_LB06HmON2_2),.dout(w_dff_B_Ns69LjTy3_2),.clk(gclk));
	jdff dff_B_g8BCCC211_2(.din(w_dff_B_Ns69LjTy3_2),.dout(w_dff_B_g8BCCC211_2),.clk(gclk));
	jdff dff_B_wbnkx0T13_2(.din(w_dff_B_g8BCCC211_2),.dout(w_dff_B_wbnkx0T13_2),.clk(gclk));
	jdff dff_B_id3uFHpD0_2(.din(w_dff_B_wbnkx0T13_2),.dout(w_dff_B_id3uFHpD0_2),.clk(gclk));
	jdff dff_B_usQTZ7oR4_2(.din(w_dff_B_id3uFHpD0_2),.dout(w_dff_B_usQTZ7oR4_2),.clk(gclk));
	jdff dff_B_c6cJmcVJ2_2(.din(w_dff_B_usQTZ7oR4_2),.dout(w_dff_B_c6cJmcVJ2_2),.clk(gclk));
	jdff dff_B_EvwR6gro0_2(.din(w_dff_B_c6cJmcVJ2_2),.dout(w_dff_B_EvwR6gro0_2),.clk(gclk));
	jdff dff_B_HoIrTVtM7_2(.din(w_dff_B_EvwR6gro0_2),.dout(w_dff_B_HoIrTVtM7_2),.clk(gclk));
	jdff dff_B_DKo8EdJc7_2(.din(w_dff_B_HoIrTVtM7_2),.dout(w_dff_B_DKo8EdJc7_2),.clk(gclk));
	jdff dff_B_7mOIfWiO7_2(.din(w_dff_B_DKo8EdJc7_2),.dout(w_dff_B_7mOIfWiO7_2),.clk(gclk));
	jdff dff_B_h6fDJDHS9_2(.din(w_dff_B_7mOIfWiO7_2),.dout(w_dff_B_h6fDJDHS9_2),.clk(gclk));
	jdff dff_B_m92kKJL86_2(.din(w_dff_B_h6fDJDHS9_2),.dout(w_dff_B_m92kKJL86_2),.clk(gclk));
	jdff dff_B_XgZGUoUN4_2(.din(w_dff_B_m92kKJL86_2),.dout(w_dff_B_XgZGUoUN4_2),.clk(gclk));
	jdff dff_B_OHfZSjCa0_2(.din(w_dff_B_XgZGUoUN4_2),.dout(w_dff_B_OHfZSjCa0_2),.clk(gclk));
	jdff dff_B_X5Dacjfa3_2(.din(w_dff_B_OHfZSjCa0_2),.dout(w_dff_B_X5Dacjfa3_2),.clk(gclk));
	jdff dff_B_DllvmJjb1_2(.din(w_dff_B_X5Dacjfa3_2),.dout(w_dff_B_DllvmJjb1_2),.clk(gclk));
	jdff dff_B_GRzYs9UU0_2(.din(w_dff_B_DllvmJjb1_2),.dout(w_dff_B_GRzYs9UU0_2),.clk(gclk));
	jdff dff_B_f0pfmsU71_2(.din(w_dff_B_GRzYs9UU0_2),.dout(w_dff_B_f0pfmsU71_2),.clk(gclk));
	jdff dff_B_OaNem0ST0_2(.din(w_dff_B_f0pfmsU71_2),.dout(w_dff_B_OaNem0ST0_2),.clk(gclk));
	jdff dff_B_72E2VBGY8_2(.din(n1449),.dout(w_dff_B_72E2VBGY8_2),.clk(gclk));
	jdff dff_B_JqiJPZgx9_1(.din(n1447),.dout(w_dff_B_JqiJPZgx9_1),.clk(gclk));
	jdff dff_B_wz2j3OsE3_2(.din(n1368),.dout(w_dff_B_wz2j3OsE3_2),.clk(gclk));
	jdff dff_B_x6OCiYCV3_2(.din(w_dff_B_wz2j3OsE3_2),.dout(w_dff_B_x6OCiYCV3_2),.clk(gclk));
	jdff dff_B_XizDq3wQ9_2(.din(w_dff_B_x6OCiYCV3_2),.dout(w_dff_B_XizDq3wQ9_2),.clk(gclk));
	jdff dff_B_l7w4yQkK1_2(.din(w_dff_B_XizDq3wQ9_2),.dout(w_dff_B_l7w4yQkK1_2),.clk(gclk));
	jdff dff_B_7zhnYyxv2_2(.din(w_dff_B_l7w4yQkK1_2),.dout(w_dff_B_7zhnYyxv2_2),.clk(gclk));
	jdff dff_B_aF4DWmiM4_2(.din(w_dff_B_7zhnYyxv2_2),.dout(w_dff_B_aF4DWmiM4_2),.clk(gclk));
	jdff dff_B_N5k7GIlI5_2(.din(w_dff_B_aF4DWmiM4_2),.dout(w_dff_B_N5k7GIlI5_2),.clk(gclk));
	jdff dff_B_9cIQunZl8_2(.din(w_dff_B_N5k7GIlI5_2),.dout(w_dff_B_9cIQunZl8_2),.clk(gclk));
	jdff dff_B_rB0COoHL2_2(.din(w_dff_B_9cIQunZl8_2),.dout(w_dff_B_rB0COoHL2_2),.clk(gclk));
	jdff dff_B_8Z5bNeUv2_2(.din(w_dff_B_rB0COoHL2_2),.dout(w_dff_B_8Z5bNeUv2_2),.clk(gclk));
	jdff dff_B_I2nQITPJ1_2(.din(w_dff_B_8Z5bNeUv2_2),.dout(w_dff_B_I2nQITPJ1_2),.clk(gclk));
	jdff dff_B_62UScHEs7_2(.din(w_dff_B_I2nQITPJ1_2),.dout(w_dff_B_62UScHEs7_2),.clk(gclk));
	jdff dff_B_nC8ZqM5K7_2(.din(w_dff_B_62UScHEs7_2),.dout(w_dff_B_nC8ZqM5K7_2),.clk(gclk));
	jdff dff_B_ZoLICgUo6_2(.din(w_dff_B_nC8ZqM5K7_2),.dout(w_dff_B_ZoLICgUo6_2),.clk(gclk));
	jdff dff_B_YLU3kOcs8_2(.din(w_dff_B_ZoLICgUo6_2),.dout(w_dff_B_YLU3kOcs8_2),.clk(gclk));
	jdff dff_B_baOsjY5c2_2(.din(w_dff_B_YLU3kOcs8_2),.dout(w_dff_B_baOsjY5c2_2),.clk(gclk));
	jdff dff_B_mxpmkjTt4_2(.din(w_dff_B_baOsjY5c2_2),.dout(w_dff_B_mxpmkjTt4_2),.clk(gclk));
	jdff dff_B_ciZMMJGM1_2(.din(w_dff_B_mxpmkjTt4_2),.dout(w_dff_B_ciZMMJGM1_2),.clk(gclk));
	jdff dff_B_Q2LiyG181_2(.din(w_dff_B_ciZMMJGM1_2),.dout(w_dff_B_Q2LiyG181_2),.clk(gclk));
	jdff dff_B_rOQXuXeo8_2(.din(w_dff_B_Q2LiyG181_2),.dout(w_dff_B_rOQXuXeo8_2),.clk(gclk));
	jdff dff_B_9Bg31B148_2(.din(w_dff_B_rOQXuXeo8_2),.dout(w_dff_B_9Bg31B148_2),.clk(gclk));
	jdff dff_B_I2zr3lj56_2(.din(w_dff_B_9Bg31B148_2),.dout(w_dff_B_I2zr3lj56_2),.clk(gclk));
	jdff dff_B_vskFeLij2_2(.din(w_dff_B_I2zr3lj56_2),.dout(w_dff_B_vskFeLij2_2),.clk(gclk));
	jdff dff_B_Aq76FbGq0_2(.din(w_dff_B_vskFeLij2_2),.dout(w_dff_B_Aq76FbGq0_2),.clk(gclk));
	jdff dff_B_Eb4qjR1P0_2(.din(w_dff_B_Aq76FbGq0_2),.dout(w_dff_B_Eb4qjR1P0_2),.clk(gclk));
	jdff dff_B_nRKGAYik5_2(.din(w_dff_B_Eb4qjR1P0_2),.dout(w_dff_B_nRKGAYik5_2),.clk(gclk));
	jdff dff_B_NOQOgkWw8_2(.din(w_dff_B_nRKGAYik5_2),.dout(w_dff_B_NOQOgkWw8_2),.clk(gclk));
	jdff dff_B_PNvyRkvI3_1(.din(n1369),.dout(w_dff_B_PNvyRkvI3_1),.clk(gclk));
	jdff dff_B_94zjszsN3_2(.din(n1283),.dout(w_dff_B_94zjszsN3_2),.clk(gclk));
	jdff dff_B_Ah8ScVZB7_2(.din(w_dff_B_94zjszsN3_2),.dout(w_dff_B_Ah8ScVZB7_2),.clk(gclk));
	jdff dff_B_WqqXRcvh2_2(.din(w_dff_B_Ah8ScVZB7_2),.dout(w_dff_B_WqqXRcvh2_2),.clk(gclk));
	jdff dff_B_mRZXVqgv4_2(.din(w_dff_B_WqqXRcvh2_2),.dout(w_dff_B_mRZXVqgv4_2),.clk(gclk));
	jdff dff_B_Pwa2BY1K2_2(.din(w_dff_B_mRZXVqgv4_2),.dout(w_dff_B_Pwa2BY1K2_2),.clk(gclk));
	jdff dff_B_eCPEyWZa9_2(.din(w_dff_B_Pwa2BY1K2_2),.dout(w_dff_B_eCPEyWZa9_2),.clk(gclk));
	jdff dff_B_mE27JYPy5_2(.din(w_dff_B_eCPEyWZa9_2),.dout(w_dff_B_mE27JYPy5_2),.clk(gclk));
	jdff dff_B_BWCfL8cj3_2(.din(w_dff_B_mE27JYPy5_2),.dout(w_dff_B_BWCfL8cj3_2),.clk(gclk));
	jdff dff_B_W6MVfBXk8_2(.din(w_dff_B_BWCfL8cj3_2),.dout(w_dff_B_W6MVfBXk8_2),.clk(gclk));
	jdff dff_B_LPcYtsBO0_2(.din(w_dff_B_W6MVfBXk8_2),.dout(w_dff_B_LPcYtsBO0_2),.clk(gclk));
	jdff dff_B_77y0nqge2_2(.din(w_dff_B_LPcYtsBO0_2),.dout(w_dff_B_77y0nqge2_2),.clk(gclk));
	jdff dff_B_ZHHbx8e05_2(.din(w_dff_B_77y0nqge2_2),.dout(w_dff_B_ZHHbx8e05_2),.clk(gclk));
	jdff dff_B_YF3wRVRy4_2(.din(w_dff_B_ZHHbx8e05_2),.dout(w_dff_B_YF3wRVRy4_2),.clk(gclk));
	jdff dff_B_yOVIrUnP1_2(.din(w_dff_B_YF3wRVRy4_2),.dout(w_dff_B_yOVIrUnP1_2),.clk(gclk));
	jdff dff_B_VWrr8tZA1_2(.din(w_dff_B_yOVIrUnP1_2),.dout(w_dff_B_VWrr8tZA1_2),.clk(gclk));
	jdff dff_B_TDPBBekm7_2(.din(w_dff_B_VWrr8tZA1_2),.dout(w_dff_B_TDPBBekm7_2),.clk(gclk));
	jdff dff_B_Kx6zWY4F7_2(.din(w_dff_B_TDPBBekm7_2),.dout(w_dff_B_Kx6zWY4F7_2),.clk(gclk));
	jdff dff_B_EdVhn0Ov9_2(.din(w_dff_B_Kx6zWY4F7_2),.dout(w_dff_B_EdVhn0Ov9_2),.clk(gclk));
	jdff dff_B_0PwMVtqr8_2(.din(w_dff_B_EdVhn0Ov9_2),.dout(w_dff_B_0PwMVtqr8_2),.clk(gclk));
	jdff dff_B_oyyZiBef2_2(.din(w_dff_B_0PwMVtqr8_2),.dout(w_dff_B_oyyZiBef2_2),.clk(gclk));
	jdff dff_B_i6g2mmxq3_2(.din(w_dff_B_oyyZiBef2_2),.dout(w_dff_B_i6g2mmxq3_2),.clk(gclk));
	jdff dff_B_t4pLYhXH6_2(.din(w_dff_B_i6g2mmxq3_2),.dout(w_dff_B_t4pLYhXH6_2),.clk(gclk));
	jdff dff_B_b0JCdIFC3_2(.din(w_dff_B_t4pLYhXH6_2),.dout(w_dff_B_b0JCdIFC3_2),.clk(gclk));
	jdff dff_B_rYzcXI5W9_2(.din(w_dff_B_b0JCdIFC3_2),.dout(w_dff_B_rYzcXI5W9_2),.clk(gclk));
	jdff dff_B_4LcJR0th3_2(.din(n1308),.dout(w_dff_B_4LcJR0th3_2),.clk(gclk));
	jdff dff_B_sMQcSNB69_1(.din(n1284),.dout(w_dff_B_sMQcSNB69_1),.clk(gclk));
	jdff dff_B_qiWnmlq81_2(.din(n1193),.dout(w_dff_B_qiWnmlq81_2),.clk(gclk));
	jdff dff_B_h0j2oLgh8_2(.din(w_dff_B_qiWnmlq81_2),.dout(w_dff_B_h0j2oLgh8_2),.clk(gclk));
	jdff dff_B_ZDT7n5Hv1_2(.din(w_dff_B_h0j2oLgh8_2),.dout(w_dff_B_ZDT7n5Hv1_2),.clk(gclk));
	jdff dff_B_RlYLjQvk9_2(.din(w_dff_B_ZDT7n5Hv1_2),.dout(w_dff_B_RlYLjQvk9_2),.clk(gclk));
	jdff dff_B_jJrQumHY0_2(.din(w_dff_B_RlYLjQvk9_2),.dout(w_dff_B_jJrQumHY0_2),.clk(gclk));
	jdff dff_B_nZoprrbN3_2(.din(w_dff_B_jJrQumHY0_2),.dout(w_dff_B_nZoprrbN3_2),.clk(gclk));
	jdff dff_B_l2NmkNVe2_2(.din(w_dff_B_nZoprrbN3_2),.dout(w_dff_B_l2NmkNVe2_2),.clk(gclk));
	jdff dff_B_rtNthS4D2_2(.din(w_dff_B_l2NmkNVe2_2),.dout(w_dff_B_rtNthS4D2_2),.clk(gclk));
	jdff dff_B_SXe0O2YX3_2(.din(w_dff_B_rtNthS4D2_2),.dout(w_dff_B_SXe0O2YX3_2),.clk(gclk));
	jdff dff_B_LIFYLMSx8_2(.din(w_dff_B_SXe0O2YX3_2),.dout(w_dff_B_LIFYLMSx8_2),.clk(gclk));
	jdff dff_B_BY7AOyL14_2(.din(w_dff_B_LIFYLMSx8_2),.dout(w_dff_B_BY7AOyL14_2),.clk(gclk));
	jdff dff_B_nhyMnMBl7_2(.din(w_dff_B_BY7AOyL14_2),.dout(w_dff_B_nhyMnMBl7_2),.clk(gclk));
	jdff dff_B_YSv1apY30_2(.din(w_dff_B_nhyMnMBl7_2),.dout(w_dff_B_YSv1apY30_2),.clk(gclk));
	jdff dff_B_h4kWvDaG6_2(.din(w_dff_B_YSv1apY30_2),.dout(w_dff_B_h4kWvDaG6_2),.clk(gclk));
	jdff dff_B_KORiv8Ni3_2(.din(w_dff_B_h4kWvDaG6_2),.dout(w_dff_B_KORiv8Ni3_2),.clk(gclk));
	jdff dff_B_ZO7wDaH22_2(.din(w_dff_B_KORiv8Ni3_2),.dout(w_dff_B_ZO7wDaH22_2),.clk(gclk));
	jdff dff_B_IwsFy9vA6_2(.din(w_dff_B_ZO7wDaH22_2),.dout(w_dff_B_IwsFy9vA6_2),.clk(gclk));
	jdff dff_B_3hAzUktV8_2(.din(w_dff_B_IwsFy9vA6_2),.dout(w_dff_B_3hAzUktV8_2),.clk(gclk));
	jdff dff_B_BMwuPzhD5_2(.din(w_dff_B_3hAzUktV8_2),.dout(w_dff_B_BMwuPzhD5_2),.clk(gclk));
	jdff dff_B_Veom8jI67_2(.din(w_dff_B_BMwuPzhD5_2),.dout(w_dff_B_Veom8jI67_2),.clk(gclk));
	jdff dff_B_m6wpOOTX3_2(.din(w_dff_B_Veom8jI67_2),.dout(w_dff_B_m6wpOOTX3_2),.clk(gclk));
	jdff dff_B_9cKVxRGY2_2(.din(n1217),.dout(w_dff_B_9cKVxRGY2_2),.clk(gclk));
	jdff dff_B_pdx9xkB96_1(.din(n1194),.dout(w_dff_B_pdx9xkB96_1),.clk(gclk));
	jdff dff_B_VxD0nNwJ2_2(.din(n1089),.dout(w_dff_B_VxD0nNwJ2_2),.clk(gclk));
	jdff dff_B_BXTyLVDb1_2(.din(w_dff_B_VxD0nNwJ2_2),.dout(w_dff_B_BXTyLVDb1_2),.clk(gclk));
	jdff dff_B_haLYPqUp7_2(.din(w_dff_B_BXTyLVDb1_2),.dout(w_dff_B_haLYPqUp7_2),.clk(gclk));
	jdff dff_B_ebf72IZ39_2(.din(w_dff_B_haLYPqUp7_2),.dout(w_dff_B_ebf72IZ39_2),.clk(gclk));
	jdff dff_B_nJzcCgIt2_2(.din(w_dff_B_ebf72IZ39_2),.dout(w_dff_B_nJzcCgIt2_2),.clk(gclk));
	jdff dff_B_2l3WI0sp5_2(.din(w_dff_B_nJzcCgIt2_2),.dout(w_dff_B_2l3WI0sp5_2),.clk(gclk));
	jdff dff_B_Y4OTmPUh0_2(.din(w_dff_B_2l3WI0sp5_2),.dout(w_dff_B_Y4OTmPUh0_2),.clk(gclk));
	jdff dff_B_xKW4vRda4_2(.din(w_dff_B_Y4OTmPUh0_2),.dout(w_dff_B_xKW4vRda4_2),.clk(gclk));
	jdff dff_B_CR9zV5al8_2(.din(w_dff_B_xKW4vRda4_2),.dout(w_dff_B_CR9zV5al8_2),.clk(gclk));
	jdff dff_B_s7EP1w689_2(.din(w_dff_B_CR9zV5al8_2),.dout(w_dff_B_s7EP1w689_2),.clk(gclk));
	jdff dff_B_M51abpuQ7_2(.din(w_dff_B_s7EP1w689_2),.dout(w_dff_B_M51abpuQ7_2),.clk(gclk));
	jdff dff_B_eIwrQVmt6_2(.din(w_dff_B_M51abpuQ7_2),.dout(w_dff_B_eIwrQVmt6_2),.clk(gclk));
	jdff dff_B_NGhfny2I7_2(.din(w_dff_B_eIwrQVmt6_2),.dout(w_dff_B_NGhfny2I7_2),.clk(gclk));
	jdff dff_B_bx12cM4l8_2(.din(w_dff_B_NGhfny2I7_2),.dout(w_dff_B_bx12cM4l8_2),.clk(gclk));
	jdff dff_B_w7SSzkEF1_2(.din(w_dff_B_bx12cM4l8_2),.dout(w_dff_B_w7SSzkEF1_2),.clk(gclk));
	jdff dff_B_ylhBoDkU3_2(.din(w_dff_B_w7SSzkEF1_2),.dout(w_dff_B_ylhBoDkU3_2),.clk(gclk));
	jdff dff_B_XUlRkKmS3_2(.din(w_dff_B_ylhBoDkU3_2),.dout(w_dff_B_XUlRkKmS3_2),.clk(gclk));
	jdff dff_B_79Wcx5u26_2(.din(w_dff_B_XUlRkKmS3_2),.dout(w_dff_B_79Wcx5u26_2),.clk(gclk));
	jdff dff_B_MqZfHPqe4_2(.din(n1119),.dout(w_dff_B_MqZfHPqe4_2),.clk(gclk));
	jdff dff_B_qDrVah190_1(.din(n1090),.dout(w_dff_B_qDrVah190_1),.clk(gclk));
	jdff dff_B_bBHxkFfT2_2(.din(n991),.dout(w_dff_B_bBHxkFfT2_2),.clk(gclk));
	jdff dff_B_wqTWrfma3_2(.din(w_dff_B_bBHxkFfT2_2),.dout(w_dff_B_wqTWrfma3_2),.clk(gclk));
	jdff dff_B_SJt05p5r3_2(.din(w_dff_B_wqTWrfma3_2),.dout(w_dff_B_SJt05p5r3_2),.clk(gclk));
	jdff dff_B_NumCiepD9_2(.din(w_dff_B_SJt05p5r3_2),.dout(w_dff_B_NumCiepD9_2),.clk(gclk));
	jdff dff_B_Ig6YHL9A9_2(.din(w_dff_B_NumCiepD9_2),.dout(w_dff_B_Ig6YHL9A9_2),.clk(gclk));
	jdff dff_B_iUJjc4pH5_2(.din(w_dff_B_Ig6YHL9A9_2),.dout(w_dff_B_iUJjc4pH5_2),.clk(gclk));
	jdff dff_B_lmYmd38Z4_2(.din(w_dff_B_iUJjc4pH5_2),.dout(w_dff_B_lmYmd38Z4_2),.clk(gclk));
	jdff dff_B_Jjln5ErG9_2(.din(w_dff_B_lmYmd38Z4_2),.dout(w_dff_B_Jjln5ErG9_2),.clk(gclk));
	jdff dff_B_1OhHQiec1_2(.din(w_dff_B_Jjln5ErG9_2),.dout(w_dff_B_1OhHQiec1_2),.clk(gclk));
	jdff dff_B_UldrICCv1_2(.din(w_dff_B_1OhHQiec1_2),.dout(w_dff_B_UldrICCv1_2),.clk(gclk));
	jdff dff_B_RXC2QJlE3_2(.din(w_dff_B_UldrICCv1_2),.dout(w_dff_B_RXC2QJlE3_2),.clk(gclk));
	jdff dff_B_MBKh6QIq4_2(.din(w_dff_B_RXC2QJlE3_2),.dout(w_dff_B_MBKh6QIq4_2),.clk(gclk));
	jdff dff_B_Yz8IP7JI9_2(.din(w_dff_B_MBKh6QIq4_2),.dout(w_dff_B_Yz8IP7JI9_2),.clk(gclk));
	jdff dff_B_bEmJq9Q26_2(.din(w_dff_B_Yz8IP7JI9_2),.dout(w_dff_B_bEmJq9Q26_2),.clk(gclk));
	jdff dff_B_8iNnw4fd3_2(.din(w_dff_B_bEmJq9Q26_2),.dout(w_dff_B_8iNnw4fd3_2),.clk(gclk));
	jdff dff_B_dUlgKmam6_2(.din(n1014),.dout(w_dff_B_dUlgKmam6_2),.clk(gclk));
	jdff dff_B_OuzEvqxX7_1(.din(n992),.dout(w_dff_B_OuzEvqxX7_1),.clk(gclk));
	jdff dff_B_p575ndzE0_2(.din(n886),.dout(w_dff_B_p575ndzE0_2),.clk(gclk));
	jdff dff_B_4tIrRp6y3_2(.din(w_dff_B_p575ndzE0_2),.dout(w_dff_B_4tIrRp6y3_2),.clk(gclk));
	jdff dff_B_aJrelXs39_2(.din(w_dff_B_4tIrRp6y3_2),.dout(w_dff_B_aJrelXs39_2),.clk(gclk));
	jdff dff_B_yX0hV0zB7_2(.din(w_dff_B_aJrelXs39_2),.dout(w_dff_B_yX0hV0zB7_2),.clk(gclk));
	jdff dff_B_LLoECp1X8_2(.din(w_dff_B_yX0hV0zB7_2),.dout(w_dff_B_LLoECp1X8_2),.clk(gclk));
	jdff dff_B_0TpDOiCf3_2(.din(w_dff_B_LLoECp1X8_2),.dout(w_dff_B_0TpDOiCf3_2),.clk(gclk));
	jdff dff_B_8IhBZRR65_2(.din(w_dff_B_0TpDOiCf3_2),.dout(w_dff_B_8IhBZRR65_2),.clk(gclk));
	jdff dff_B_blKFOxBF6_2(.din(w_dff_B_8IhBZRR65_2),.dout(w_dff_B_blKFOxBF6_2),.clk(gclk));
	jdff dff_B_QEGnW7u19_2(.din(w_dff_B_blKFOxBF6_2),.dout(w_dff_B_QEGnW7u19_2),.clk(gclk));
	jdff dff_B_L4wEvSvt2_2(.din(w_dff_B_QEGnW7u19_2),.dout(w_dff_B_L4wEvSvt2_2),.clk(gclk));
	jdff dff_B_kweSgKqg4_2(.din(w_dff_B_L4wEvSvt2_2),.dout(w_dff_B_kweSgKqg4_2),.clk(gclk));
	jdff dff_B_0l63gjYM2_2(.din(w_dff_B_kweSgKqg4_2),.dout(w_dff_B_0l63gjYM2_2),.clk(gclk));
	jdff dff_B_FMIx6HkA4_2(.din(n909),.dout(w_dff_B_FMIx6HkA4_2),.clk(gclk));
	jdff dff_B_Th5MwW257_1(.din(n887),.dout(w_dff_B_Th5MwW257_1),.clk(gclk));
	jdff dff_B_NcUp0Ci72_2(.din(n787),.dout(w_dff_B_NcUp0Ci72_2),.clk(gclk));
	jdff dff_B_c3TfShXe5_2(.din(w_dff_B_NcUp0Ci72_2),.dout(w_dff_B_c3TfShXe5_2),.clk(gclk));
	jdff dff_B_fTBGaos44_2(.din(w_dff_B_c3TfShXe5_2),.dout(w_dff_B_fTBGaos44_2),.clk(gclk));
	jdff dff_B_g2SpbvpB2_2(.din(w_dff_B_fTBGaos44_2),.dout(w_dff_B_g2SpbvpB2_2),.clk(gclk));
	jdff dff_B_OxVT2tcz6_2(.din(w_dff_B_g2SpbvpB2_2),.dout(w_dff_B_OxVT2tcz6_2),.clk(gclk));
	jdff dff_B_Rlhd1RZ53_2(.din(w_dff_B_OxVT2tcz6_2),.dout(w_dff_B_Rlhd1RZ53_2),.clk(gclk));
	jdff dff_B_XFxrXvdU6_2(.din(w_dff_B_Rlhd1RZ53_2),.dout(w_dff_B_XFxrXvdU6_2),.clk(gclk));
	jdff dff_B_0hucysWl5_2(.din(w_dff_B_XFxrXvdU6_2),.dout(w_dff_B_0hucysWl5_2),.clk(gclk));
	jdff dff_B_eylds8PW2_2(.din(w_dff_B_0hucysWl5_2),.dout(w_dff_B_eylds8PW2_2),.clk(gclk));
	jdff dff_B_r2tZCzxO0_2(.din(n803),.dout(w_dff_B_r2tZCzxO0_2),.clk(gclk));
	jdff dff_B_yseD4T131_2(.din(w_dff_B_r2tZCzxO0_2),.dout(w_dff_B_yseD4T131_2),.clk(gclk));
	jdff dff_B_8UsONRXs4_1(.din(n788),.dout(w_dff_B_8UsONRXs4_1),.clk(gclk));
	jdff dff_B_i5s3NL2W3_1(.din(w_dff_B_8UsONRXs4_1),.dout(w_dff_B_i5s3NL2W3_1),.clk(gclk));
	jdff dff_B_UXBtV24U6_1(.din(w_dff_B_i5s3NL2W3_1),.dout(w_dff_B_UXBtV24U6_1),.clk(gclk));
	jdff dff_B_yhLU7zb81_1(.din(w_dff_B_UXBtV24U6_1),.dout(w_dff_B_yhLU7zb81_1),.clk(gclk));
	jdff dff_B_z1IWhVkG5_1(.din(w_dff_B_yhLU7zb81_1),.dout(w_dff_B_z1IWhVkG5_1),.clk(gclk));
	jdff dff_B_Z6o9Hakd3_1(.din(w_dff_B_z1IWhVkG5_1),.dout(w_dff_B_Z6o9Hakd3_1),.clk(gclk));
	jdff dff_B_SJeyUxvo2_0(.din(n703),.dout(w_dff_B_SJeyUxvo2_0),.clk(gclk));
	jdff dff_B_wrk2j1G20_0(.din(w_dff_B_SJeyUxvo2_0),.dout(w_dff_B_wrk2j1G20_0),.clk(gclk));
	jdff dff_A_MrsLvblf1_0(.dout(w_n702_0[0]),.din(w_dff_A_MrsLvblf1_0),.clk(gclk));
	jdff dff_A_R9Z5k56G0_0(.dout(w_dff_A_MrsLvblf1_0),.din(w_dff_A_R9Z5k56G0_0),.clk(gclk));
	jdff dff_A_sw2PtKtX2_0(.dout(w_dff_A_R9Z5k56G0_0),.din(w_dff_A_sw2PtKtX2_0),.clk(gclk));
	jdff dff_B_2psNJ8Fq6_1(.din(n696),.dout(w_dff_B_2psNJ8Fq6_1),.clk(gclk));
	jdff dff_A_vN8Ty6XF4_0(.dout(w_n607_0[0]),.din(w_dff_A_vN8Ty6XF4_0),.clk(gclk));
	jdff dff_A_Tru88F5E9_1(.dout(w_n607_0[1]),.din(w_dff_A_Tru88F5E9_1),.clk(gclk));
	jdff dff_A_srnRvMnm4_1(.dout(w_dff_A_Tru88F5E9_1),.din(w_dff_A_srnRvMnm4_1),.clk(gclk));
	jdff dff_A_z36lHbXL5_1(.dout(w_n694_0[1]),.din(w_dff_A_z36lHbXL5_1),.clk(gclk));
	jdff dff_A_Ib01DOzk8_1(.dout(w_dff_A_z36lHbXL5_1),.din(w_dff_A_Ib01DOzk8_1),.clk(gclk));
	jdff dff_A_Ou5AVYtg3_1(.dout(w_dff_A_Ib01DOzk8_1),.din(w_dff_A_Ou5AVYtg3_1),.clk(gclk));
	jdff dff_A_yDHm8PpD2_1(.dout(w_dff_A_Ou5AVYtg3_1),.din(w_dff_A_yDHm8PpD2_1),.clk(gclk));
	jdff dff_A_F1pYYuP78_1(.dout(w_dff_A_yDHm8PpD2_1),.din(w_dff_A_F1pYYuP78_1),.clk(gclk));
	jdff dff_A_04uEiypF3_1(.dout(w_dff_A_F1pYYuP78_1),.din(w_dff_A_04uEiypF3_1),.clk(gclk));
	jdff dff_B_LOyfXsth5_1(.din(n1819),.dout(w_dff_B_LOyfXsth5_1),.clk(gclk));
	jdff dff_A_Hvb89mYh3_1(.dout(w_n1801_0[1]),.din(w_dff_A_Hvb89mYh3_1),.clk(gclk));
	jdff dff_B_mSbZR5nX4_1(.din(n1799),.dout(w_dff_B_mSbZR5nX4_1),.clk(gclk));
	jdff dff_B_Ejj13FDg1_2(.din(n1770),.dout(w_dff_B_Ejj13FDg1_2),.clk(gclk));
	jdff dff_B_umvEI9Vo6_2(.din(w_dff_B_Ejj13FDg1_2),.dout(w_dff_B_umvEI9Vo6_2),.clk(gclk));
	jdff dff_B_FUzfAqvL8_2(.din(w_dff_B_umvEI9Vo6_2),.dout(w_dff_B_FUzfAqvL8_2),.clk(gclk));
	jdff dff_B_ITm47nRE0_2(.din(w_dff_B_FUzfAqvL8_2),.dout(w_dff_B_ITm47nRE0_2),.clk(gclk));
	jdff dff_B_IvY5Cxcl5_2(.din(w_dff_B_ITm47nRE0_2),.dout(w_dff_B_IvY5Cxcl5_2),.clk(gclk));
	jdff dff_B_xrEQa0iw9_2(.din(w_dff_B_IvY5Cxcl5_2),.dout(w_dff_B_xrEQa0iw9_2),.clk(gclk));
	jdff dff_B_iB3dktwx3_2(.din(w_dff_B_xrEQa0iw9_2),.dout(w_dff_B_iB3dktwx3_2),.clk(gclk));
	jdff dff_B_IcjrXihW5_2(.din(w_dff_B_iB3dktwx3_2),.dout(w_dff_B_IcjrXihW5_2),.clk(gclk));
	jdff dff_B_oCmQpDPh9_2(.din(w_dff_B_IcjrXihW5_2),.dout(w_dff_B_oCmQpDPh9_2),.clk(gclk));
	jdff dff_B_j0oG0F0G4_2(.din(w_dff_B_oCmQpDPh9_2),.dout(w_dff_B_j0oG0F0G4_2),.clk(gclk));
	jdff dff_B_z8J6ruUG0_2(.din(w_dff_B_j0oG0F0G4_2),.dout(w_dff_B_z8J6ruUG0_2),.clk(gclk));
	jdff dff_B_pGJKsymL9_2(.din(w_dff_B_z8J6ruUG0_2),.dout(w_dff_B_pGJKsymL9_2),.clk(gclk));
	jdff dff_B_L8IgM5Zy6_2(.din(w_dff_B_pGJKsymL9_2),.dout(w_dff_B_L8IgM5Zy6_2),.clk(gclk));
	jdff dff_B_8m2k3oyM8_2(.din(w_dff_B_L8IgM5Zy6_2),.dout(w_dff_B_8m2k3oyM8_2),.clk(gclk));
	jdff dff_B_YwRopqfB3_2(.din(w_dff_B_8m2k3oyM8_2),.dout(w_dff_B_YwRopqfB3_2),.clk(gclk));
	jdff dff_B_GEsXNV6y5_2(.din(w_dff_B_YwRopqfB3_2),.dout(w_dff_B_GEsXNV6y5_2),.clk(gclk));
	jdff dff_B_p0xbA5Ai8_2(.din(w_dff_B_GEsXNV6y5_2),.dout(w_dff_B_p0xbA5Ai8_2),.clk(gclk));
	jdff dff_B_q6XIlSm58_2(.din(w_dff_B_p0xbA5Ai8_2),.dout(w_dff_B_q6XIlSm58_2),.clk(gclk));
	jdff dff_B_Q5qOZsg61_2(.din(w_dff_B_q6XIlSm58_2),.dout(w_dff_B_Q5qOZsg61_2),.clk(gclk));
	jdff dff_B_qh1sDJVQ2_2(.din(w_dff_B_Q5qOZsg61_2),.dout(w_dff_B_qh1sDJVQ2_2),.clk(gclk));
	jdff dff_B_VuvW6dgs2_2(.din(w_dff_B_qh1sDJVQ2_2),.dout(w_dff_B_VuvW6dgs2_2),.clk(gclk));
	jdff dff_B_IGKpHItS6_2(.din(w_dff_B_VuvW6dgs2_2),.dout(w_dff_B_IGKpHItS6_2),.clk(gclk));
	jdff dff_B_cHEDTrUP0_2(.din(w_dff_B_IGKpHItS6_2),.dout(w_dff_B_cHEDTrUP0_2),.clk(gclk));
	jdff dff_B_0YQkRkXF8_2(.din(w_dff_B_cHEDTrUP0_2),.dout(w_dff_B_0YQkRkXF8_2),.clk(gclk));
	jdff dff_B_Kj2OZhRL7_2(.din(w_dff_B_0YQkRkXF8_2),.dout(w_dff_B_Kj2OZhRL7_2),.clk(gclk));
	jdff dff_B_OYx71PWU9_2(.din(w_dff_B_Kj2OZhRL7_2),.dout(w_dff_B_OYx71PWU9_2),.clk(gclk));
	jdff dff_B_V6KxGlsT4_2(.din(w_dff_B_OYx71PWU9_2),.dout(w_dff_B_V6KxGlsT4_2),.clk(gclk));
	jdff dff_B_g9hd9jit8_2(.din(w_dff_B_V6KxGlsT4_2),.dout(w_dff_B_g9hd9jit8_2),.clk(gclk));
	jdff dff_B_vXpvzYHM7_2(.din(w_dff_B_g9hd9jit8_2),.dout(w_dff_B_vXpvzYHM7_2),.clk(gclk));
	jdff dff_B_UjGuASmA9_2(.din(w_dff_B_vXpvzYHM7_2),.dout(w_dff_B_UjGuASmA9_2),.clk(gclk));
	jdff dff_B_WGXuEf7o3_2(.din(w_dff_B_UjGuASmA9_2),.dout(w_dff_B_WGXuEf7o3_2),.clk(gclk));
	jdff dff_B_5nc5dami1_2(.din(w_dff_B_WGXuEf7o3_2),.dout(w_dff_B_5nc5dami1_2),.clk(gclk));
	jdff dff_B_lvsYMnRp1_2(.din(w_dff_B_5nc5dami1_2),.dout(w_dff_B_lvsYMnRp1_2),.clk(gclk));
	jdff dff_B_qWuLwY080_2(.din(w_dff_B_lvsYMnRp1_2),.dout(w_dff_B_qWuLwY080_2),.clk(gclk));
	jdff dff_B_oiOybrMn6_2(.din(w_dff_B_qWuLwY080_2),.dout(w_dff_B_oiOybrMn6_2),.clk(gclk));
	jdff dff_B_r6KyqbrR0_2(.din(w_dff_B_oiOybrMn6_2),.dout(w_dff_B_r6KyqbrR0_2),.clk(gclk));
	jdff dff_B_XnZgAs7f9_2(.din(w_dff_B_r6KyqbrR0_2),.dout(w_dff_B_XnZgAs7f9_2),.clk(gclk));
	jdff dff_B_NODFih3y9_2(.din(w_dff_B_XnZgAs7f9_2),.dout(w_dff_B_NODFih3y9_2),.clk(gclk));
	jdff dff_B_fLzc46Ce3_2(.din(w_dff_B_NODFih3y9_2),.dout(w_dff_B_fLzc46Ce3_2),.clk(gclk));
	jdff dff_B_42jNCee70_2(.din(w_dff_B_fLzc46Ce3_2),.dout(w_dff_B_42jNCee70_2),.clk(gclk));
	jdff dff_B_yeWMj1072_2(.din(w_dff_B_42jNCee70_2),.dout(w_dff_B_yeWMj1072_2),.clk(gclk));
	jdff dff_B_Aojw71c43_2(.din(w_dff_B_yeWMj1072_2),.dout(w_dff_B_Aojw71c43_2),.clk(gclk));
	jdff dff_B_mU5xv5Ij6_2(.din(w_dff_B_Aojw71c43_2),.dout(w_dff_B_mU5xv5Ij6_2),.clk(gclk));
	jdff dff_B_srGj8NzH7_2(.din(w_dff_B_mU5xv5Ij6_2),.dout(w_dff_B_srGj8NzH7_2),.clk(gclk));
	jdff dff_B_4PXeIdUz4_2(.din(w_dff_B_srGj8NzH7_2),.dout(w_dff_B_4PXeIdUz4_2),.clk(gclk));
	jdff dff_B_Ko9Gsvxi5_2(.din(w_dff_B_4PXeIdUz4_2),.dout(w_dff_B_Ko9Gsvxi5_2),.clk(gclk));
	jdff dff_B_wHB96kvt5_2(.din(w_dff_B_Ko9Gsvxi5_2),.dout(w_dff_B_wHB96kvt5_2),.clk(gclk));
	jdff dff_B_ACndFeqS3_2(.din(w_dff_B_wHB96kvt5_2),.dout(w_dff_B_ACndFeqS3_2),.clk(gclk));
	jdff dff_B_ykurAHmU2_2(.din(w_dff_B_ACndFeqS3_2),.dout(w_dff_B_ykurAHmU2_2),.clk(gclk));
	jdff dff_B_fQEvWDZd2_2(.din(w_dff_B_ykurAHmU2_2),.dout(w_dff_B_fQEvWDZd2_2),.clk(gclk));
	jdff dff_B_iwbOJypr8_2(.din(w_dff_B_fQEvWDZd2_2),.dout(w_dff_B_iwbOJypr8_2),.clk(gclk));
	jdff dff_B_rXXBjKT04_2(.din(w_dff_B_iwbOJypr8_2),.dout(w_dff_B_rXXBjKT04_2),.clk(gclk));
	jdff dff_B_ZmG8bPWg0_2(.din(w_dff_B_rXXBjKT04_2),.dout(w_dff_B_ZmG8bPWg0_2),.clk(gclk));
	jdff dff_B_75PHjK6M9_2(.din(n1773),.dout(w_dff_B_75PHjK6M9_2),.clk(gclk));
	jdff dff_B_41ptGfqe8_1(.din(n1771),.dout(w_dff_B_41ptGfqe8_1),.clk(gclk));
	jdff dff_B_geUBvjFh7_2(.din(n1735),.dout(w_dff_B_geUBvjFh7_2),.clk(gclk));
	jdff dff_B_RZKNY6CS2_2(.din(w_dff_B_geUBvjFh7_2),.dout(w_dff_B_RZKNY6CS2_2),.clk(gclk));
	jdff dff_B_pf1BbJ5J8_2(.din(w_dff_B_RZKNY6CS2_2),.dout(w_dff_B_pf1BbJ5J8_2),.clk(gclk));
	jdff dff_B_EWnqIpaA8_2(.din(w_dff_B_pf1BbJ5J8_2),.dout(w_dff_B_EWnqIpaA8_2),.clk(gclk));
	jdff dff_B_Li1A4bY65_2(.din(w_dff_B_EWnqIpaA8_2),.dout(w_dff_B_Li1A4bY65_2),.clk(gclk));
	jdff dff_B_f6PjTMbV3_2(.din(w_dff_B_Li1A4bY65_2),.dout(w_dff_B_f6PjTMbV3_2),.clk(gclk));
	jdff dff_B_0H3tDfsL7_2(.din(w_dff_B_f6PjTMbV3_2),.dout(w_dff_B_0H3tDfsL7_2),.clk(gclk));
	jdff dff_B_lwAyrWz72_2(.din(w_dff_B_0H3tDfsL7_2),.dout(w_dff_B_lwAyrWz72_2),.clk(gclk));
	jdff dff_B_7HTn104q4_2(.din(w_dff_B_lwAyrWz72_2),.dout(w_dff_B_7HTn104q4_2),.clk(gclk));
	jdff dff_B_z1vOFJ5q5_2(.din(w_dff_B_7HTn104q4_2),.dout(w_dff_B_z1vOFJ5q5_2),.clk(gclk));
	jdff dff_B_WkGOZLW77_2(.din(w_dff_B_z1vOFJ5q5_2),.dout(w_dff_B_WkGOZLW77_2),.clk(gclk));
	jdff dff_B_BU0WOKZz5_2(.din(w_dff_B_WkGOZLW77_2),.dout(w_dff_B_BU0WOKZz5_2),.clk(gclk));
	jdff dff_B_cyCdttq31_2(.din(w_dff_B_BU0WOKZz5_2),.dout(w_dff_B_cyCdttq31_2),.clk(gclk));
	jdff dff_B_m9MlvMKq4_2(.din(w_dff_B_cyCdttq31_2),.dout(w_dff_B_m9MlvMKq4_2),.clk(gclk));
	jdff dff_B_60oNfWN27_2(.din(w_dff_B_m9MlvMKq4_2),.dout(w_dff_B_60oNfWN27_2),.clk(gclk));
	jdff dff_B_XQV099jo4_2(.din(w_dff_B_60oNfWN27_2),.dout(w_dff_B_XQV099jo4_2),.clk(gclk));
	jdff dff_B_MHVfk0DL6_2(.din(w_dff_B_XQV099jo4_2),.dout(w_dff_B_MHVfk0DL6_2),.clk(gclk));
	jdff dff_B_Jnz2xk1V0_2(.din(w_dff_B_MHVfk0DL6_2),.dout(w_dff_B_Jnz2xk1V0_2),.clk(gclk));
	jdff dff_B_41HSxumI2_2(.din(w_dff_B_Jnz2xk1V0_2),.dout(w_dff_B_41HSxumI2_2),.clk(gclk));
	jdff dff_B_QhLlWjY38_2(.din(w_dff_B_41HSxumI2_2),.dout(w_dff_B_QhLlWjY38_2),.clk(gclk));
	jdff dff_B_MqyGJm1L5_2(.din(w_dff_B_QhLlWjY38_2),.dout(w_dff_B_MqyGJm1L5_2),.clk(gclk));
	jdff dff_B_r41UVl7Y9_2(.din(w_dff_B_MqyGJm1L5_2),.dout(w_dff_B_r41UVl7Y9_2),.clk(gclk));
	jdff dff_B_ELVGJrJk8_2(.din(w_dff_B_r41UVl7Y9_2),.dout(w_dff_B_ELVGJrJk8_2),.clk(gclk));
	jdff dff_B_e4tBWFxm6_2(.din(w_dff_B_ELVGJrJk8_2),.dout(w_dff_B_e4tBWFxm6_2),.clk(gclk));
	jdff dff_B_vPXOdMit6_2(.din(w_dff_B_e4tBWFxm6_2),.dout(w_dff_B_vPXOdMit6_2),.clk(gclk));
	jdff dff_B_56FuqRwM2_2(.din(w_dff_B_vPXOdMit6_2),.dout(w_dff_B_56FuqRwM2_2),.clk(gclk));
	jdff dff_B_nIL7XCRY7_2(.din(w_dff_B_56FuqRwM2_2),.dout(w_dff_B_nIL7XCRY7_2),.clk(gclk));
	jdff dff_B_SIZ9O1VG9_2(.din(w_dff_B_nIL7XCRY7_2),.dout(w_dff_B_SIZ9O1VG9_2),.clk(gclk));
	jdff dff_B_k3WNy3345_2(.din(w_dff_B_SIZ9O1VG9_2),.dout(w_dff_B_k3WNy3345_2),.clk(gclk));
	jdff dff_B_c75UBdPK7_2(.din(w_dff_B_k3WNy3345_2),.dout(w_dff_B_c75UBdPK7_2),.clk(gclk));
	jdff dff_B_xmVdhNrQ0_2(.din(w_dff_B_c75UBdPK7_2),.dout(w_dff_B_xmVdhNrQ0_2),.clk(gclk));
	jdff dff_B_903JaLxB3_2(.din(w_dff_B_xmVdhNrQ0_2),.dout(w_dff_B_903JaLxB3_2),.clk(gclk));
	jdff dff_B_0mrL5mLA8_2(.din(w_dff_B_903JaLxB3_2),.dout(w_dff_B_0mrL5mLA8_2),.clk(gclk));
	jdff dff_B_jYjJuIVq3_2(.din(w_dff_B_0mrL5mLA8_2),.dout(w_dff_B_jYjJuIVq3_2),.clk(gclk));
	jdff dff_B_g0jwsfyE0_2(.din(w_dff_B_jYjJuIVq3_2),.dout(w_dff_B_g0jwsfyE0_2),.clk(gclk));
	jdff dff_B_QFvel9269_2(.din(w_dff_B_g0jwsfyE0_2),.dout(w_dff_B_QFvel9269_2),.clk(gclk));
	jdff dff_B_qogUaso08_2(.din(w_dff_B_QFvel9269_2),.dout(w_dff_B_qogUaso08_2),.clk(gclk));
	jdff dff_B_l8fT2krH8_2(.din(w_dff_B_qogUaso08_2),.dout(w_dff_B_l8fT2krH8_2),.clk(gclk));
	jdff dff_B_C7tR32BQ0_2(.din(w_dff_B_l8fT2krH8_2),.dout(w_dff_B_C7tR32BQ0_2),.clk(gclk));
	jdff dff_B_76XomXZs9_2(.din(w_dff_B_C7tR32BQ0_2),.dout(w_dff_B_76XomXZs9_2),.clk(gclk));
	jdff dff_B_J0Ufhwpm7_2(.din(w_dff_B_76XomXZs9_2),.dout(w_dff_B_J0Ufhwpm7_2),.clk(gclk));
	jdff dff_B_fTyxRqd77_2(.din(w_dff_B_J0Ufhwpm7_2),.dout(w_dff_B_fTyxRqd77_2),.clk(gclk));
	jdff dff_B_pj1VU2v43_2(.din(w_dff_B_fTyxRqd77_2),.dout(w_dff_B_pj1VU2v43_2),.clk(gclk));
	jdff dff_B_uHePrxfz2_2(.din(w_dff_B_pj1VU2v43_2),.dout(w_dff_B_uHePrxfz2_2),.clk(gclk));
	jdff dff_B_4r5AkvxC9_2(.din(w_dff_B_uHePrxfz2_2),.dout(w_dff_B_4r5AkvxC9_2),.clk(gclk));
	jdff dff_B_U7wureC74_2(.din(w_dff_B_4r5AkvxC9_2),.dout(w_dff_B_U7wureC74_2),.clk(gclk));
	jdff dff_B_gqDYvhZe3_2(.din(w_dff_B_U7wureC74_2),.dout(w_dff_B_gqDYvhZe3_2),.clk(gclk));
	jdff dff_B_uF3q11ah9_2(.din(w_dff_B_gqDYvhZe3_2),.dout(w_dff_B_uF3q11ah9_2),.clk(gclk));
	jdff dff_B_5oksoLxC0_2(.din(w_dff_B_uF3q11ah9_2),.dout(w_dff_B_5oksoLxC0_2),.clk(gclk));
	jdff dff_B_kfVdW4aC6_2(.din(n1738),.dout(w_dff_B_kfVdW4aC6_2),.clk(gclk));
	jdff dff_B_gC3Rv0z41_1(.din(n1736),.dout(w_dff_B_gC3Rv0z41_1),.clk(gclk));
	jdff dff_B_jT8LzB527_2(.din(n1694),.dout(w_dff_B_jT8LzB527_2),.clk(gclk));
	jdff dff_B_W0ZmB8Ho4_2(.din(w_dff_B_jT8LzB527_2),.dout(w_dff_B_W0ZmB8Ho4_2),.clk(gclk));
	jdff dff_B_AmiSepg94_2(.din(w_dff_B_W0ZmB8Ho4_2),.dout(w_dff_B_AmiSepg94_2),.clk(gclk));
	jdff dff_B_3fgl0hCo3_2(.din(w_dff_B_AmiSepg94_2),.dout(w_dff_B_3fgl0hCo3_2),.clk(gclk));
	jdff dff_B_Qc5DzA5Q8_2(.din(w_dff_B_3fgl0hCo3_2),.dout(w_dff_B_Qc5DzA5Q8_2),.clk(gclk));
	jdff dff_B_sW3pWa7H3_2(.din(w_dff_B_Qc5DzA5Q8_2),.dout(w_dff_B_sW3pWa7H3_2),.clk(gclk));
	jdff dff_B_FJblDYcg0_2(.din(w_dff_B_sW3pWa7H3_2),.dout(w_dff_B_FJblDYcg0_2),.clk(gclk));
	jdff dff_B_bIPXvJRG1_2(.din(w_dff_B_FJblDYcg0_2),.dout(w_dff_B_bIPXvJRG1_2),.clk(gclk));
	jdff dff_B_gsznbvZ46_2(.din(w_dff_B_bIPXvJRG1_2),.dout(w_dff_B_gsznbvZ46_2),.clk(gclk));
	jdff dff_B_5Fihdx7n4_2(.din(w_dff_B_gsznbvZ46_2),.dout(w_dff_B_5Fihdx7n4_2),.clk(gclk));
	jdff dff_B_i0yZvowo8_2(.din(w_dff_B_5Fihdx7n4_2),.dout(w_dff_B_i0yZvowo8_2),.clk(gclk));
	jdff dff_B_eWz0jVWp9_2(.din(w_dff_B_i0yZvowo8_2),.dout(w_dff_B_eWz0jVWp9_2),.clk(gclk));
	jdff dff_B_ntf0nUQE3_2(.din(w_dff_B_eWz0jVWp9_2),.dout(w_dff_B_ntf0nUQE3_2),.clk(gclk));
	jdff dff_B_doikCE2z5_2(.din(w_dff_B_ntf0nUQE3_2),.dout(w_dff_B_doikCE2z5_2),.clk(gclk));
	jdff dff_B_ipaRpm2w1_2(.din(w_dff_B_doikCE2z5_2),.dout(w_dff_B_ipaRpm2w1_2),.clk(gclk));
	jdff dff_B_yyjjj4Qy8_2(.din(w_dff_B_ipaRpm2w1_2),.dout(w_dff_B_yyjjj4Qy8_2),.clk(gclk));
	jdff dff_B_swsjroU35_2(.din(w_dff_B_yyjjj4Qy8_2),.dout(w_dff_B_swsjroU35_2),.clk(gclk));
	jdff dff_B_XQVhgTYB8_2(.din(w_dff_B_swsjroU35_2),.dout(w_dff_B_XQVhgTYB8_2),.clk(gclk));
	jdff dff_B_XMIeaaOw0_2(.din(w_dff_B_XQVhgTYB8_2),.dout(w_dff_B_XMIeaaOw0_2),.clk(gclk));
	jdff dff_B_c8b6EEaw5_2(.din(w_dff_B_XMIeaaOw0_2),.dout(w_dff_B_c8b6EEaw5_2),.clk(gclk));
	jdff dff_B_4WMR2ZzK2_2(.din(w_dff_B_c8b6EEaw5_2),.dout(w_dff_B_4WMR2ZzK2_2),.clk(gclk));
	jdff dff_B_YvCy8vvI3_2(.din(w_dff_B_4WMR2ZzK2_2),.dout(w_dff_B_YvCy8vvI3_2),.clk(gclk));
	jdff dff_B_NtPpTp807_2(.din(w_dff_B_YvCy8vvI3_2),.dout(w_dff_B_NtPpTp807_2),.clk(gclk));
	jdff dff_B_ulFXfwZm0_2(.din(w_dff_B_NtPpTp807_2),.dout(w_dff_B_ulFXfwZm0_2),.clk(gclk));
	jdff dff_B_HtplOrIW4_2(.din(w_dff_B_ulFXfwZm0_2),.dout(w_dff_B_HtplOrIW4_2),.clk(gclk));
	jdff dff_B_l1DokOau1_2(.din(w_dff_B_HtplOrIW4_2),.dout(w_dff_B_l1DokOau1_2),.clk(gclk));
	jdff dff_B_E4SZPomJ6_2(.din(w_dff_B_l1DokOau1_2),.dout(w_dff_B_E4SZPomJ6_2),.clk(gclk));
	jdff dff_B_s6U3UHmG4_2(.din(w_dff_B_E4SZPomJ6_2),.dout(w_dff_B_s6U3UHmG4_2),.clk(gclk));
	jdff dff_B_cGHYqfnb2_2(.din(w_dff_B_s6U3UHmG4_2),.dout(w_dff_B_cGHYqfnb2_2),.clk(gclk));
	jdff dff_B_TnAnl9QO9_2(.din(w_dff_B_cGHYqfnb2_2),.dout(w_dff_B_TnAnl9QO9_2),.clk(gclk));
	jdff dff_B_3gfV9m352_2(.din(w_dff_B_TnAnl9QO9_2),.dout(w_dff_B_3gfV9m352_2),.clk(gclk));
	jdff dff_B_s1tnnurs4_2(.din(w_dff_B_3gfV9m352_2),.dout(w_dff_B_s1tnnurs4_2),.clk(gclk));
	jdff dff_B_7PwPP5Cm1_2(.din(w_dff_B_s1tnnurs4_2),.dout(w_dff_B_7PwPP5Cm1_2),.clk(gclk));
	jdff dff_B_2tQ9lGuU8_2(.din(w_dff_B_7PwPP5Cm1_2),.dout(w_dff_B_2tQ9lGuU8_2),.clk(gclk));
	jdff dff_B_QmzEqv8E2_2(.din(w_dff_B_2tQ9lGuU8_2),.dout(w_dff_B_QmzEqv8E2_2),.clk(gclk));
	jdff dff_B_AS7lg4Kf4_2(.din(w_dff_B_QmzEqv8E2_2),.dout(w_dff_B_AS7lg4Kf4_2),.clk(gclk));
	jdff dff_B_whwD1eTk2_2(.din(w_dff_B_AS7lg4Kf4_2),.dout(w_dff_B_whwD1eTk2_2),.clk(gclk));
	jdff dff_B_LDEa0inY4_2(.din(w_dff_B_whwD1eTk2_2),.dout(w_dff_B_LDEa0inY4_2),.clk(gclk));
	jdff dff_B_4VzBaOai2_2(.din(w_dff_B_LDEa0inY4_2),.dout(w_dff_B_4VzBaOai2_2),.clk(gclk));
	jdff dff_B_hd3L1nA42_2(.din(w_dff_B_4VzBaOai2_2),.dout(w_dff_B_hd3L1nA42_2),.clk(gclk));
	jdff dff_B_ijvmdrRa9_2(.din(w_dff_B_hd3L1nA42_2),.dout(w_dff_B_ijvmdrRa9_2),.clk(gclk));
	jdff dff_B_xu4GHzgO6_2(.din(w_dff_B_ijvmdrRa9_2),.dout(w_dff_B_xu4GHzgO6_2),.clk(gclk));
	jdff dff_B_Ibm9RoZ63_2(.din(w_dff_B_xu4GHzgO6_2),.dout(w_dff_B_Ibm9RoZ63_2),.clk(gclk));
	jdff dff_B_NXJungvK4_2(.din(w_dff_B_Ibm9RoZ63_2),.dout(w_dff_B_NXJungvK4_2),.clk(gclk));
	jdff dff_B_BGuYp3u05_2(.din(w_dff_B_NXJungvK4_2),.dout(w_dff_B_BGuYp3u05_2),.clk(gclk));
	jdff dff_B_7bx0Xb2Q0_2(.din(n1697),.dout(w_dff_B_7bx0Xb2Q0_2),.clk(gclk));
	jdff dff_B_bCY77S658_1(.din(n1695),.dout(w_dff_B_bCY77S658_1),.clk(gclk));
	jdff dff_B_V6RJLTFs0_2(.din(n1643),.dout(w_dff_B_V6RJLTFs0_2),.clk(gclk));
	jdff dff_B_h2jtc9p91_2(.din(w_dff_B_V6RJLTFs0_2),.dout(w_dff_B_h2jtc9p91_2),.clk(gclk));
	jdff dff_B_3ltZOvc64_2(.din(w_dff_B_h2jtc9p91_2),.dout(w_dff_B_3ltZOvc64_2),.clk(gclk));
	jdff dff_B_7S3PMFjP1_2(.din(w_dff_B_3ltZOvc64_2),.dout(w_dff_B_7S3PMFjP1_2),.clk(gclk));
	jdff dff_B_88fwvHQb1_2(.din(w_dff_B_7S3PMFjP1_2),.dout(w_dff_B_88fwvHQb1_2),.clk(gclk));
	jdff dff_B_sbClGWUO8_2(.din(w_dff_B_88fwvHQb1_2),.dout(w_dff_B_sbClGWUO8_2),.clk(gclk));
	jdff dff_B_SISSsBgx5_2(.din(w_dff_B_sbClGWUO8_2),.dout(w_dff_B_SISSsBgx5_2),.clk(gclk));
	jdff dff_B_FMlXwUqq6_2(.din(w_dff_B_SISSsBgx5_2),.dout(w_dff_B_FMlXwUqq6_2),.clk(gclk));
	jdff dff_B_Cj8FaT1T8_2(.din(w_dff_B_FMlXwUqq6_2),.dout(w_dff_B_Cj8FaT1T8_2),.clk(gclk));
	jdff dff_B_92FFWy2l9_2(.din(w_dff_B_Cj8FaT1T8_2),.dout(w_dff_B_92FFWy2l9_2),.clk(gclk));
	jdff dff_B_ylJbDdbT2_2(.din(w_dff_B_92FFWy2l9_2),.dout(w_dff_B_ylJbDdbT2_2),.clk(gclk));
	jdff dff_B_TFaJemOH3_2(.din(w_dff_B_ylJbDdbT2_2),.dout(w_dff_B_TFaJemOH3_2),.clk(gclk));
	jdff dff_B_O6SJOrJG9_2(.din(w_dff_B_TFaJemOH3_2),.dout(w_dff_B_O6SJOrJG9_2),.clk(gclk));
	jdff dff_B_vOmZ0eok6_2(.din(w_dff_B_O6SJOrJG9_2),.dout(w_dff_B_vOmZ0eok6_2),.clk(gclk));
	jdff dff_B_IscFfvsp6_2(.din(w_dff_B_vOmZ0eok6_2),.dout(w_dff_B_IscFfvsp6_2),.clk(gclk));
	jdff dff_B_r8LAgrPk4_2(.din(w_dff_B_IscFfvsp6_2),.dout(w_dff_B_r8LAgrPk4_2),.clk(gclk));
	jdff dff_B_qoeSUkIe6_2(.din(w_dff_B_r8LAgrPk4_2),.dout(w_dff_B_qoeSUkIe6_2),.clk(gclk));
	jdff dff_B_mfI2KR4f3_2(.din(w_dff_B_qoeSUkIe6_2),.dout(w_dff_B_mfI2KR4f3_2),.clk(gclk));
	jdff dff_B_VGU6obil9_2(.din(w_dff_B_mfI2KR4f3_2),.dout(w_dff_B_VGU6obil9_2),.clk(gclk));
	jdff dff_B_foXoIVQb9_2(.din(w_dff_B_VGU6obil9_2),.dout(w_dff_B_foXoIVQb9_2),.clk(gclk));
	jdff dff_B_OEHadiIT7_2(.din(w_dff_B_foXoIVQb9_2),.dout(w_dff_B_OEHadiIT7_2),.clk(gclk));
	jdff dff_B_uv7ME0AH9_2(.din(w_dff_B_OEHadiIT7_2),.dout(w_dff_B_uv7ME0AH9_2),.clk(gclk));
	jdff dff_B_gbScNmri3_2(.din(w_dff_B_uv7ME0AH9_2),.dout(w_dff_B_gbScNmri3_2),.clk(gclk));
	jdff dff_B_fGgc8efR3_2(.din(w_dff_B_gbScNmri3_2),.dout(w_dff_B_fGgc8efR3_2),.clk(gclk));
	jdff dff_B_7wAcj6WB8_2(.din(w_dff_B_fGgc8efR3_2),.dout(w_dff_B_7wAcj6WB8_2),.clk(gclk));
	jdff dff_B_0cocnuP30_2(.din(w_dff_B_7wAcj6WB8_2),.dout(w_dff_B_0cocnuP30_2),.clk(gclk));
	jdff dff_B_ZJQ4THPG5_2(.din(w_dff_B_0cocnuP30_2),.dout(w_dff_B_ZJQ4THPG5_2),.clk(gclk));
	jdff dff_B_ZBK0Ce3x0_2(.din(w_dff_B_ZJQ4THPG5_2),.dout(w_dff_B_ZBK0Ce3x0_2),.clk(gclk));
	jdff dff_B_V08ECaFc4_2(.din(w_dff_B_ZBK0Ce3x0_2),.dout(w_dff_B_V08ECaFc4_2),.clk(gclk));
	jdff dff_B_rMaAlsfY6_2(.din(w_dff_B_V08ECaFc4_2),.dout(w_dff_B_rMaAlsfY6_2),.clk(gclk));
	jdff dff_B_2bGgQ2qh5_2(.din(w_dff_B_rMaAlsfY6_2),.dout(w_dff_B_2bGgQ2qh5_2),.clk(gclk));
	jdff dff_B_Xdt4naIX0_2(.din(w_dff_B_2bGgQ2qh5_2),.dout(w_dff_B_Xdt4naIX0_2),.clk(gclk));
	jdff dff_B_p5vZOwmM8_2(.din(w_dff_B_Xdt4naIX0_2),.dout(w_dff_B_p5vZOwmM8_2),.clk(gclk));
	jdff dff_B_QCKbahQL3_2(.din(w_dff_B_p5vZOwmM8_2),.dout(w_dff_B_QCKbahQL3_2),.clk(gclk));
	jdff dff_B_MGN1ipDK0_2(.din(w_dff_B_QCKbahQL3_2),.dout(w_dff_B_MGN1ipDK0_2),.clk(gclk));
	jdff dff_B_H4YxNmQo7_2(.din(w_dff_B_MGN1ipDK0_2),.dout(w_dff_B_H4YxNmQo7_2),.clk(gclk));
	jdff dff_B_XkRIf8Hz2_2(.din(w_dff_B_H4YxNmQo7_2),.dout(w_dff_B_XkRIf8Hz2_2),.clk(gclk));
	jdff dff_B_Mp2ifXT79_2(.din(w_dff_B_XkRIf8Hz2_2),.dout(w_dff_B_Mp2ifXT79_2),.clk(gclk));
	jdff dff_B_MquMrvv39_2(.din(w_dff_B_Mp2ifXT79_2),.dout(w_dff_B_MquMrvv39_2),.clk(gclk));
	jdff dff_B_U0h6fLI23_2(.din(w_dff_B_MquMrvv39_2),.dout(w_dff_B_U0h6fLI23_2),.clk(gclk));
	jdff dff_B_3rVbqRBO3_2(.din(w_dff_B_U0h6fLI23_2),.dout(w_dff_B_3rVbqRBO3_2),.clk(gclk));
	jdff dff_B_hHfKE0vn2_2(.din(n1646),.dout(w_dff_B_hHfKE0vn2_2),.clk(gclk));
	jdff dff_B_8uuf1NPF9_1(.din(n1644),.dout(w_dff_B_8uuf1NPF9_1),.clk(gclk));
	jdff dff_B_8W0a4QFq5_2(.din(n1586),.dout(w_dff_B_8W0a4QFq5_2),.clk(gclk));
	jdff dff_B_Zzr90bZu7_2(.din(w_dff_B_8W0a4QFq5_2),.dout(w_dff_B_Zzr90bZu7_2),.clk(gclk));
	jdff dff_B_oCpmkZgS4_2(.din(w_dff_B_Zzr90bZu7_2),.dout(w_dff_B_oCpmkZgS4_2),.clk(gclk));
	jdff dff_B_cSpuQyeN8_2(.din(w_dff_B_oCpmkZgS4_2),.dout(w_dff_B_cSpuQyeN8_2),.clk(gclk));
	jdff dff_B_czLHytWY8_2(.din(w_dff_B_cSpuQyeN8_2),.dout(w_dff_B_czLHytWY8_2),.clk(gclk));
	jdff dff_B_Od2bjCmf6_2(.din(w_dff_B_czLHytWY8_2),.dout(w_dff_B_Od2bjCmf6_2),.clk(gclk));
	jdff dff_B_y7pZWHVO9_2(.din(w_dff_B_Od2bjCmf6_2),.dout(w_dff_B_y7pZWHVO9_2),.clk(gclk));
	jdff dff_B_upvZbSKu0_2(.din(w_dff_B_y7pZWHVO9_2),.dout(w_dff_B_upvZbSKu0_2),.clk(gclk));
	jdff dff_B_ajmSSkjV0_2(.din(w_dff_B_upvZbSKu0_2),.dout(w_dff_B_ajmSSkjV0_2),.clk(gclk));
	jdff dff_B_G1OcHUp34_2(.din(w_dff_B_ajmSSkjV0_2),.dout(w_dff_B_G1OcHUp34_2),.clk(gclk));
	jdff dff_B_8jcfrtjq0_2(.din(w_dff_B_G1OcHUp34_2),.dout(w_dff_B_8jcfrtjq0_2),.clk(gclk));
	jdff dff_B_FdIi7iov8_2(.din(w_dff_B_8jcfrtjq0_2),.dout(w_dff_B_FdIi7iov8_2),.clk(gclk));
	jdff dff_B_8dYf9r8b4_2(.din(w_dff_B_FdIi7iov8_2),.dout(w_dff_B_8dYf9r8b4_2),.clk(gclk));
	jdff dff_B_kSqZamUx9_2(.din(w_dff_B_8dYf9r8b4_2),.dout(w_dff_B_kSqZamUx9_2),.clk(gclk));
	jdff dff_B_a6ufy1Un4_2(.din(w_dff_B_kSqZamUx9_2),.dout(w_dff_B_a6ufy1Un4_2),.clk(gclk));
	jdff dff_B_XmwejyP26_2(.din(w_dff_B_a6ufy1Un4_2),.dout(w_dff_B_XmwejyP26_2),.clk(gclk));
	jdff dff_B_rllJl9KP3_2(.din(w_dff_B_XmwejyP26_2),.dout(w_dff_B_rllJl9KP3_2),.clk(gclk));
	jdff dff_B_G2fqfeIo8_2(.din(w_dff_B_rllJl9KP3_2),.dout(w_dff_B_G2fqfeIo8_2),.clk(gclk));
	jdff dff_B_jKMgF7Qh3_2(.din(w_dff_B_G2fqfeIo8_2),.dout(w_dff_B_jKMgF7Qh3_2),.clk(gclk));
	jdff dff_B_o1VfcBMx8_2(.din(w_dff_B_jKMgF7Qh3_2),.dout(w_dff_B_o1VfcBMx8_2),.clk(gclk));
	jdff dff_B_gMCmfg1B0_2(.din(w_dff_B_o1VfcBMx8_2),.dout(w_dff_B_gMCmfg1B0_2),.clk(gclk));
	jdff dff_B_xlvvTZfE2_2(.din(w_dff_B_gMCmfg1B0_2),.dout(w_dff_B_xlvvTZfE2_2),.clk(gclk));
	jdff dff_B_BWvDlSpP4_2(.din(w_dff_B_xlvvTZfE2_2),.dout(w_dff_B_BWvDlSpP4_2),.clk(gclk));
	jdff dff_B_vVK2PL6q3_2(.din(w_dff_B_BWvDlSpP4_2),.dout(w_dff_B_vVK2PL6q3_2),.clk(gclk));
	jdff dff_B_TV50pzx35_2(.din(w_dff_B_vVK2PL6q3_2),.dout(w_dff_B_TV50pzx35_2),.clk(gclk));
	jdff dff_B_vhoxp4Az4_2(.din(w_dff_B_TV50pzx35_2),.dout(w_dff_B_vhoxp4Az4_2),.clk(gclk));
	jdff dff_B_wayJIXNz8_2(.din(w_dff_B_vhoxp4Az4_2),.dout(w_dff_B_wayJIXNz8_2),.clk(gclk));
	jdff dff_B_K2Xhf19H5_2(.din(w_dff_B_wayJIXNz8_2),.dout(w_dff_B_K2Xhf19H5_2),.clk(gclk));
	jdff dff_B_25U39w9H4_2(.din(w_dff_B_K2Xhf19H5_2),.dout(w_dff_B_25U39w9H4_2),.clk(gclk));
	jdff dff_B_Cus5OcBd0_2(.din(w_dff_B_25U39w9H4_2),.dout(w_dff_B_Cus5OcBd0_2),.clk(gclk));
	jdff dff_B_Q9jgfP202_2(.din(w_dff_B_Cus5OcBd0_2),.dout(w_dff_B_Q9jgfP202_2),.clk(gclk));
	jdff dff_B_Dccwno3t9_2(.din(w_dff_B_Q9jgfP202_2),.dout(w_dff_B_Dccwno3t9_2),.clk(gclk));
	jdff dff_B_7Nhz5uH56_2(.din(w_dff_B_Dccwno3t9_2),.dout(w_dff_B_7Nhz5uH56_2),.clk(gclk));
	jdff dff_B_UOCWkoL34_2(.din(w_dff_B_7Nhz5uH56_2),.dout(w_dff_B_UOCWkoL34_2),.clk(gclk));
	jdff dff_B_aWQQDVVC9_2(.din(w_dff_B_UOCWkoL34_2),.dout(w_dff_B_aWQQDVVC9_2),.clk(gclk));
	jdff dff_B_OGKro7M29_2(.din(w_dff_B_aWQQDVVC9_2),.dout(w_dff_B_OGKro7M29_2),.clk(gclk));
	jdff dff_B_uxlbT8043_2(.din(w_dff_B_OGKro7M29_2),.dout(w_dff_B_uxlbT8043_2),.clk(gclk));
	jdff dff_B_niD869Mu6_2(.din(n1589),.dout(w_dff_B_niD869Mu6_2),.clk(gclk));
	jdff dff_B_AjoZInzR4_1(.din(n1587),.dout(w_dff_B_AjoZInzR4_1),.clk(gclk));
	jdff dff_B_pIjbyzw96_2(.din(n1522),.dout(w_dff_B_pIjbyzw96_2),.clk(gclk));
	jdff dff_B_n5eLjJz29_2(.din(w_dff_B_pIjbyzw96_2),.dout(w_dff_B_n5eLjJz29_2),.clk(gclk));
	jdff dff_B_tZuXqGTK5_2(.din(w_dff_B_n5eLjJz29_2),.dout(w_dff_B_tZuXqGTK5_2),.clk(gclk));
	jdff dff_B_Ibq5R8j12_2(.din(w_dff_B_tZuXqGTK5_2),.dout(w_dff_B_Ibq5R8j12_2),.clk(gclk));
	jdff dff_B_Jvq2UC8s7_2(.din(w_dff_B_Ibq5R8j12_2),.dout(w_dff_B_Jvq2UC8s7_2),.clk(gclk));
	jdff dff_B_Rt1K60Na5_2(.din(w_dff_B_Jvq2UC8s7_2),.dout(w_dff_B_Rt1K60Na5_2),.clk(gclk));
	jdff dff_B_BkDZH8WR6_2(.din(w_dff_B_Rt1K60Na5_2),.dout(w_dff_B_BkDZH8WR6_2),.clk(gclk));
	jdff dff_B_tWaOV1KK1_2(.din(w_dff_B_BkDZH8WR6_2),.dout(w_dff_B_tWaOV1KK1_2),.clk(gclk));
	jdff dff_B_CJMzdSok6_2(.din(w_dff_B_tWaOV1KK1_2),.dout(w_dff_B_CJMzdSok6_2),.clk(gclk));
	jdff dff_B_ztQmL6nz0_2(.din(w_dff_B_CJMzdSok6_2),.dout(w_dff_B_ztQmL6nz0_2),.clk(gclk));
	jdff dff_B_9mqc3Ao92_2(.din(w_dff_B_ztQmL6nz0_2),.dout(w_dff_B_9mqc3Ao92_2),.clk(gclk));
	jdff dff_B_O3W17pQ15_2(.din(w_dff_B_9mqc3Ao92_2),.dout(w_dff_B_O3W17pQ15_2),.clk(gclk));
	jdff dff_B_J4Zz7LsP4_2(.din(w_dff_B_O3W17pQ15_2),.dout(w_dff_B_J4Zz7LsP4_2),.clk(gclk));
	jdff dff_B_2KWcHWup0_2(.din(w_dff_B_J4Zz7LsP4_2),.dout(w_dff_B_2KWcHWup0_2),.clk(gclk));
	jdff dff_B_QUmbG9yf1_2(.din(w_dff_B_2KWcHWup0_2),.dout(w_dff_B_QUmbG9yf1_2),.clk(gclk));
	jdff dff_B_hla1cY9Y8_2(.din(w_dff_B_QUmbG9yf1_2),.dout(w_dff_B_hla1cY9Y8_2),.clk(gclk));
	jdff dff_B_GEzHCmKz5_2(.din(w_dff_B_hla1cY9Y8_2),.dout(w_dff_B_GEzHCmKz5_2),.clk(gclk));
	jdff dff_B_auESlpph5_2(.din(w_dff_B_GEzHCmKz5_2),.dout(w_dff_B_auESlpph5_2),.clk(gclk));
	jdff dff_B_4f3I6soJ2_2(.din(w_dff_B_auESlpph5_2),.dout(w_dff_B_4f3I6soJ2_2),.clk(gclk));
	jdff dff_B_95CPVkjc1_2(.din(w_dff_B_4f3I6soJ2_2),.dout(w_dff_B_95CPVkjc1_2),.clk(gclk));
	jdff dff_B_Lvfo8yf86_2(.din(w_dff_B_95CPVkjc1_2),.dout(w_dff_B_Lvfo8yf86_2),.clk(gclk));
	jdff dff_B_GzjYyes91_2(.din(w_dff_B_Lvfo8yf86_2),.dout(w_dff_B_GzjYyes91_2),.clk(gclk));
	jdff dff_B_FEuV478o9_2(.din(w_dff_B_GzjYyes91_2),.dout(w_dff_B_FEuV478o9_2),.clk(gclk));
	jdff dff_B_0YoGJYha3_2(.din(w_dff_B_FEuV478o9_2),.dout(w_dff_B_0YoGJYha3_2),.clk(gclk));
	jdff dff_B_a09rMzAG5_2(.din(w_dff_B_0YoGJYha3_2),.dout(w_dff_B_a09rMzAG5_2),.clk(gclk));
	jdff dff_B_EzDJem7c1_2(.din(w_dff_B_a09rMzAG5_2),.dout(w_dff_B_EzDJem7c1_2),.clk(gclk));
	jdff dff_B_wCBlYzyR4_2(.din(w_dff_B_EzDJem7c1_2),.dout(w_dff_B_wCBlYzyR4_2),.clk(gclk));
	jdff dff_B_IzqOz8po1_2(.din(w_dff_B_wCBlYzyR4_2),.dout(w_dff_B_IzqOz8po1_2),.clk(gclk));
	jdff dff_B_u9zubPfy8_2(.din(w_dff_B_IzqOz8po1_2),.dout(w_dff_B_u9zubPfy8_2),.clk(gclk));
	jdff dff_B_UtBZzhJt2_2(.din(w_dff_B_u9zubPfy8_2),.dout(w_dff_B_UtBZzhJt2_2),.clk(gclk));
	jdff dff_B_n0ikSsPP2_2(.din(w_dff_B_UtBZzhJt2_2),.dout(w_dff_B_n0ikSsPP2_2),.clk(gclk));
	jdff dff_B_4GVukgXr0_2(.din(w_dff_B_n0ikSsPP2_2),.dout(w_dff_B_4GVukgXr0_2),.clk(gclk));
	jdff dff_B_8pMa8pGJ1_2(.din(w_dff_B_4GVukgXr0_2),.dout(w_dff_B_8pMa8pGJ1_2),.clk(gclk));
	jdff dff_B_wZRVoe8d1_2(.din(n1525),.dout(w_dff_B_wZRVoe8d1_2),.clk(gclk));
	jdff dff_B_CPSDcxeo0_1(.din(n1523),.dout(w_dff_B_CPSDcxeo0_1),.clk(gclk));
	jdff dff_B_pkIXgoCW0_2(.din(n1451),.dout(w_dff_B_pkIXgoCW0_2),.clk(gclk));
	jdff dff_B_qL122ReC9_2(.din(w_dff_B_pkIXgoCW0_2),.dout(w_dff_B_qL122ReC9_2),.clk(gclk));
	jdff dff_B_CEfFlcDu0_2(.din(w_dff_B_qL122ReC9_2),.dout(w_dff_B_CEfFlcDu0_2),.clk(gclk));
	jdff dff_B_OaUVFtHj8_2(.din(w_dff_B_CEfFlcDu0_2),.dout(w_dff_B_OaUVFtHj8_2),.clk(gclk));
	jdff dff_B_m5Xpi6ss2_2(.din(w_dff_B_OaUVFtHj8_2),.dout(w_dff_B_m5Xpi6ss2_2),.clk(gclk));
	jdff dff_B_Gu7VTcKj0_2(.din(w_dff_B_m5Xpi6ss2_2),.dout(w_dff_B_Gu7VTcKj0_2),.clk(gclk));
	jdff dff_B_MmVG5Zm49_2(.din(w_dff_B_Gu7VTcKj0_2),.dout(w_dff_B_MmVG5Zm49_2),.clk(gclk));
	jdff dff_B_SY2MVKr11_2(.din(w_dff_B_MmVG5Zm49_2),.dout(w_dff_B_SY2MVKr11_2),.clk(gclk));
	jdff dff_B_SvmLfalu9_2(.din(w_dff_B_SY2MVKr11_2),.dout(w_dff_B_SvmLfalu9_2),.clk(gclk));
	jdff dff_B_DPx3AT5T9_2(.din(w_dff_B_SvmLfalu9_2),.dout(w_dff_B_DPx3AT5T9_2),.clk(gclk));
	jdff dff_B_FhunLZ0A9_2(.din(w_dff_B_DPx3AT5T9_2),.dout(w_dff_B_FhunLZ0A9_2),.clk(gclk));
	jdff dff_B_D7zCsoZQ5_2(.din(w_dff_B_FhunLZ0A9_2),.dout(w_dff_B_D7zCsoZQ5_2),.clk(gclk));
	jdff dff_B_6YSeV2Bq1_2(.din(w_dff_B_D7zCsoZQ5_2),.dout(w_dff_B_6YSeV2Bq1_2),.clk(gclk));
	jdff dff_B_WSKAjr3g2_2(.din(w_dff_B_6YSeV2Bq1_2),.dout(w_dff_B_WSKAjr3g2_2),.clk(gclk));
	jdff dff_B_R7UFBQkP5_2(.din(w_dff_B_WSKAjr3g2_2),.dout(w_dff_B_R7UFBQkP5_2),.clk(gclk));
	jdff dff_B_r2PpmB2L5_2(.din(w_dff_B_R7UFBQkP5_2),.dout(w_dff_B_r2PpmB2L5_2),.clk(gclk));
	jdff dff_B_D4DvMUMe3_2(.din(w_dff_B_r2PpmB2L5_2),.dout(w_dff_B_D4DvMUMe3_2),.clk(gclk));
	jdff dff_B_bThkq4ZT6_2(.din(w_dff_B_D4DvMUMe3_2),.dout(w_dff_B_bThkq4ZT6_2),.clk(gclk));
	jdff dff_B_7giKRh5M5_2(.din(w_dff_B_bThkq4ZT6_2),.dout(w_dff_B_7giKRh5M5_2),.clk(gclk));
	jdff dff_B_YVUhQyBk8_2(.din(w_dff_B_7giKRh5M5_2),.dout(w_dff_B_YVUhQyBk8_2),.clk(gclk));
	jdff dff_B_JOFnZy7U4_2(.din(w_dff_B_YVUhQyBk8_2),.dout(w_dff_B_JOFnZy7U4_2),.clk(gclk));
	jdff dff_B_yjMxemBL2_2(.din(w_dff_B_JOFnZy7U4_2),.dout(w_dff_B_yjMxemBL2_2),.clk(gclk));
	jdff dff_B_YQvke0zO7_2(.din(w_dff_B_yjMxemBL2_2),.dout(w_dff_B_YQvke0zO7_2),.clk(gclk));
	jdff dff_B_5iujL0oo1_2(.din(w_dff_B_YQvke0zO7_2),.dout(w_dff_B_5iujL0oo1_2),.clk(gclk));
	jdff dff_B_eE3jrWdx9_2(.din(w_dff_B_5iujL0oo1_2),.dout(w_dff_B_eE3jrWdx9_2),.clk(gclk));
	jdff dff_B_J1uBbdG53_2(.din(w_dff_B_eE3jrWdx9_2),.dout(w_dff_B_J1uBbdG53_2),.clk(gclk));
	jdff dff_B_kUxMpTmz3_2(.din(w_dff_B_J1uBbdG53_2),.dout(w_dff_B_kUxMpTmz3_2),.clk(gclk));
	jdff dff_B_zzFGn0zt8_2(.din(w_dff_B_kUxMpTmz3_2),.dout(w_dff_B_zzFGn0zt8_2),.clk(gclk));
	jdff dff_B_PgDjnd6z1_2(.din(w_dff_B_zzFGn0zt8_2),.dout(w_dff_B_PgDjnd6z1_2),.clk(gclk));
	jdff dff_B_L7rgudxM0_2(.din(n1454),.dout(w_dff_B_L7rgudxM0_2),.clk(gclk));
	jdff dff_B_2eWKUzzW9_1(.din(n1452),.dout(w_dff_B_2eWKUzzW9_1),.clk(gclk));
	jdff dff_B_91JATJxl9_2(.din(n1373),.dout(w_dff_B_91JATJxl9_2),.clk(gclk));
	jdff dff_B_AQSNkDys5_2(.din(w_dff_B_91JATJxl9_2),.dout(w_dff_B_AQSNkDys5_2),.clk(gclk));
	jdff dff_B_J3129anV8_2(.din(w_dff_B_AQSNkDys5_2),.dout(w_dff_B_J3129anV8_2),.clk(gclk));
	jdff dff_B_YYa7I4iS4_2(.din(w_dff_B_J3129anV8_2),.dout(w_dff_B_YYa7I4iS4_2),.clk(gclk));
	jdff dff_B_RqZR2cBd7_2(.din(w_dff_B_YYa7I4iS4_2),.dout(w_dff_B_RqZR2cBd7_2),.clk(gclk));
	jdff dff_B_anPhin0E3_2(.din(w_dff_B_RqZR2cBd7_2),.dout(w_dff_B_anPhin0E3_2),.clk(gclk));
	jdff dff_B_Fi8zziLH7_2(.din(w_dff_B_anPhin0E3_2),.dout(w_dff_B_Fi8zziLH7_2),.clk(gclk));
	jdff dff_B_7YMmdHuy7_2(.din(w_dff_B_Fi8zziLH7_2),.dout(w_dff_B_7YMmdHuy7_2),.clk(gclk));
	jdff dff_B_oH0vbbef6_2(.din(w_dff_B_7YMmdHuy7_2),.dout(w_dff_B_oH0vbbef6_2),.clk(gclk));
	jdff dff_B_XkDJSfbK4_2(.din(w_dff_B_oH0vbbef6_2),.dout(w_dff_B_XkDJSfbK4_2),.clk(gclk));
	jdff dff_B_MlgJ31f45_2(.din(w_dff_B_XkDJSfbK4_2),.dout(w_dff_B_MlgJ31f45_2),.clk(gclk));
	jdff dff_B_EUG5hBs56_2(.din(w_dff_B_MlgJ31f45_2),.dout(w_dff_B_EUG5hBs56_2),.clk(gclk));
	jdff dff_B_HjeZR5zt2_2(.din(w_dff_B_EUG5hBs56_2),.dout(w_dff_B_HjeZR5zt2_2),.clk(gclk));
	jdff dff_B_tob1Cp0L5_2(.din(w_dff_B_HjeZR5zt2_2),.dout(w_dff_B_tob1Cp0L5_2),.clk(gclk));
	jdff dff_B_SSKae8cT4_2(.din(w_dff_B_tob1Cp0L5_2),.dout(w_dff_B_SSKae8cT4_2),.clk(gclk));
	jdff dff_B_oKdZxUj41_2(.din(w_dff_B_SSKae8cT4_2),.dout(w_dff_B_oKdZxUj41_2),.clk(gclk));
	jdff dff_B_DjMOWeJy8_2(.din(w_dff_B_oKdZxUj41_2),.dout(w_dff_B_DjMOWeJy8_2),.clk(gclk));
	jdff dff_B_XstjE5572_2(.din(w_dff_B_DjMOWeJy8_2),.dout(w_dff_B_XstjE5572_2),.clk(gclk));
	jdff dff_B_SdX8df405_2(.din(w_dff_B_XstjE5572_2),.dout(w_dff_B_SdX8df405_2),.clk(gclk));
	jdff dff_B_d6OQDYRy6_2(.din(w_dff_B_SdX8df405_2),.dout(w_dff_B_d6OQDYRy6_2),.clk(gclk));
	jdff dff_B_p0SDXEes4_2(.din(w_dff_B_d6OQDYRy6_2),.dout(w_dff_B_p0SDXEes4_2),.clk(gclk));
	jdff dff_B_3rnfloFZ3_2(.din(w_dff_B_p0SDXEes4_2),.dout(w_dff_B_3rnfloFZ3_2),.clk(gclk));
	jdff dff_B_FH9w0fmJ4_2(.din(w_dff_B_3rnfloFZ3_2),.dout(w_dff_B_FH9w0fmJ4_2),.clk(gclk));
	jdff dff_B_Wx7Efk4F4_2(.din(w_dff_B_FH9w0fmJ4_2),.dout(w_dff_B_Wx7Efk4F4_2),.clk(gclk));
	jdff dff_B_XlOikqK90_2(.din(w_dff_B_Wx7Efk4F4_2),.dout(w_dff_B_XlOikqK90_2),.clk(gclk));
	jdff dff_B_TmNOlf9n0_2(.din(n1376),.dout(w_dff_B_TmNOlf9n0_2),.clk(gclk));
	jdff dff_B_RtdkC2mD4_1(.din(n1374),.dout(w_dff_B_RtdkC2mD4_1),.clk(gclk));
	jdff dff_B_6PfcSkGz6_2(.din(n1288),.dout(w_dff_B_6PfcSkGz6_2),.clk(gclk));
	jdff dff_B_oBviVAW80_2(.din(w_dff_B_6PfcSkGz6_2),.dout(w_dff_B_oBviVAW80_2),.clk(gclk));
	jdff dff_B_PQN2gM129_2(.din(w_dff_B_oBviVAW80_2),.dout(w_dff_B_PQN2gM129_2),.clk(gclk));
	jdff dff_B_NHsx9DbZ8_2(.din(w_dff_B_PQN2gM129_2),.dout(w_dff_B_NHsx9DbZ8_2),.clk(gclk));
	jdff dff_B_Hu68tsAF5_2(.din(w_dff_B_NHsx9DbZ8_2),.dout(w_dff_B_Hu68tsAF5_2),.clk(gclk));
	jdff dff_B_fz7Cus5n0_2(.din(w_dff_B_Hu68tsAF5_2),.dout(w_dff_B_fz7Cus5n0_2),.clk(gclk));
	jdff dff_B_x06G9Chp7_2(.din(w_dff_B_fz7Cus5n0_2),.dout(w_dff_B_x06G9Chp7_2),.clk(gclk));
	jdff dff_B_swhybO3A6_2(.din(w_dff_B_x06G9Chp7_2),.dout(w_dff_B_swhybO3A6_2),.clk(gclk));
	jdff dff_B_fy4x7IpU2_2(.din(w_dff_B_swhybO3A6_2),.dout(w_dff_B_fy4x7IpU2_2),.clk(gclk));
	jdff dff_B_GT8MMnUN9_2(.din(w_dff_B_fy4x7IpU2_2),.dout(w_dff_B_GT8MMnUN9_2),.clk(gclk));
	jdff dff_B_R8GnHqlY7_2(.din(w_dff_B_GT8MMnUN9_2),.dout(w_dff_B_R8GnHqlY7_2),.clk(gclk));
	jdff dff_B_BmKcjgLl8_2(.din(w_dff_B_R8GnHqlY7_2),.dout(w_dff_B_BmKcjgLl8_2),.clk(gclk));
	jdff dff_B_KvB2Wl8E0_2(.din(w_dff_B_BmKcjgLl8_2),.dout(w_dff_B_KvB2Wl8E0_2),.clk(gclk));
	jdff dff_B_n0CsZ01L3_2(.din(w_dff_B_KvB2Wl8E0_2),.dout(w_dff_B_n0CsZ01L3_2),.clk(gclk));
	jdff dff_B_KK4ApRKM8_2(.din(w_dff_B_n0CsZ01L3_2),.dout(w_dff_B_KK4ApRKM8_2),.clk(gclk));
	jdff dff_B_7gxUUBDR9_2(.din(w_dff_B_KK4ApRKM8_2),.dout(w_dff_B_7gxUUBDR9_2),.clk(gclk));
	jdff dff_B_4f0ajlLY9_2(.din(w_dff_B_7gxUUBDR9_2),.dout(w_dff_B_4f0ajlLY9_2),.clk(gclk));
	jdff dff_B_ILKuVmAd9_2(.din(w_dff_B_4f0ajlLY9_2),.dout(w_dff_B_ILKuVmAd9_2),.clk(gclk));
	jdff dff_B_QRIHWUsw8_2(.din(w_dff_B_ILKuVmAd9_2),.dout(w_dff_B_QRIHWUsw8_2),.clk(gclk));
	jdff dff_B_HnGLTB9O7_2(.din(w_dff_B_QRIHWUsw8_2),.dout(w_dff_B_HnGLTB9O7_2),.clk(gclk));
	jdff dff_B_GP9JAZhC8_2(.din(w_dff_B_HnGLTB9O7_2),.dout(w_dff_B_GP9JAZhC8_2),.clk(gclk));
	jdff dff_B_Fo72BbEF4_1(.din(n1289),.dout(w_dff_B_Fo72BbEF4_1),.clk(gclk));
	jdff dff_B_LVlIYL3C2_2(.din(n1198),.dout(w_dff_B_LVlIYL3C2_2),.clk(gclk));
	jdff dff_B_ZWCw7MDQ5_2(.din(w_dff_B_LVlIYL3C2_2),.dout(w_dff_B_ZWCw7MDQ5_2),.clk(gclk));
	jdff dff_B_faN7JA1a0_2(.din(w_dff_B_ZWCw7MDQ5_2),.dout(w_dff_B_faN7JA1a0_2),.clk(gclk));
	jdff dff_B_zjF7C7RV7_2(.din(w_dff_B_faN7JA1a0_2),.dout(w_dff_B_zjF7C7RV7_2),.clk(gclk));
	jdff dff_B_rfzX121o4_2(.din(w_dff_B_zjF7C7RV7_2),.dout(w_dff_B_rfzX121o4_2),.clk(gclk));
	jdff dff_B_Kxrdym9R8_2(.din(w_dff_B_rfzX121o4_2),.dout(w_dff_B_Kxrdym9R8_2),.clk(gclk));
	jdff dff_B_HIpDGStJ0_2(.din(w_dff_B_Kxrdym9R8_2),.dout(w_dff_B_HIpDGStJ0_2),.clk(gclk));
	jdff dff_B_8366iCDu3_2(.din(w_dff_B_HIpDGStJ0_2),.dout(w_dff_B_8366iCDu3_2),.clk(gclk));
	jdff dff_B_8YZY78lu5_2(.din(w_dff_B_8366iCDu3_2),.dout(w_dff_B_8YZY78lu5_2),.clk(gclk));
	jdff dff_B_9NA4N8Lp3_2(.din(w_dff_B_8YZY78lu5_2),.dout(w_dff_B_9NA4N8Lp3_2),.clk(gclk));
	jdff dff_B_aLLSB5Lk2_2(.din(w_dff_B_9NA4N8Lp3_2),.dout(w_dff_B_aLLSB5Lk2_2),.clk(gclk));
	jdff dff_B_4hhFZWI41_2(.din(w_dff_B_aLLSB5Lk2_2),.dout(w_dff_B_4hhFZWI41_2),.clk(gclk));
	jdff dff_B_0fFqT3866_2(.din(w_dff_B_4hhFZWI41_2),.dout(w_dff_B_0fFqT3866_2),.clk(gclk));
	jdff dff_B_6kwJyHEd0_2(.din(w_dff_B_0fFqT3866_2),.dout(w_dff_B_6kwJyHEd0_2),.clk(gclk));
	jdff dff_B_c4BHIpOz5_2(.din(w_dff_B_6kwJyHEd0_2),.dout(w_dff_B_c4BHIpOz5_2),.clk(gclk));
	jdff dff_B_vcEkbXEZ7_2(.din(w_dff_B_c4BHIpOz5_2),.dout(w_dff_B_vcEkbXEZ7_2),.clk(gclk));
	jdff dff_B_LMs7POFQ8_2(.din(w_dff_B_vcEkbXEZ7_2),.dout(w_dff_B_LMs7POFQ8_2),.clk(gclk));
	jdff dff_B_5p8CRa7h9_2(.din(w_dff_B_LMs7POFQ8_2),.dout(w_dff_B_5p8CRa7h9_2),.clk(gclk));
	jdff dff_B_vZPtaRWA8_2(.din(n1215),.dout(w_dff_B_vZPtaRWA8_2),.clk(gclk));
	jdff dff_B_VX0TK40R4_1(.din(n1199),.dout(w_dff_B_VX0TK40R4_1),.clk(gclk));
	jdff dff_B_cz58degP2_2(.din(n1094),.dout(w_dff_B_cz58degP2_2),.clk(gclk));
	jdff dff_B_vrSXT5b96_2(.din(w_dff_B_cz58degP2_2),.dout(w_dff_B_vrSXT5b96_2),.clk(gclk));
	jdff dff_B_sHe4B7qA3_2(.din(w_dff_B_vrSXT5b96_2),.dout(w_dff_B_sHe4B7qA3_2),.clk(gclk));
	jdff dff_B_aIdpIA1u1_2(.din(w_dff_B_sHe4B7qA3_2),.dout(w_dff_B_aIdpIA1u1_2),.clk(gclk));
	jdff dff_B_I0EmQrU52_2(.din(w_dff_B_aIdpIA1u1_2),.dout(w_dff_B_I0EmQrU52_2),.clk(gclk));
	jdff dff_B_tLuahK4X4_2(.din(w_dff_B_I0EmQrU52_2),.dout(w_dff_B_tLuahK4X4_2),.clk(gclk));
	jdff dff_B_0BatgX1U8_2(.din(w_dff_B_tLuahK4X4_2),.dout(w_dff_B_0BatgX1U8_2),.clk(gclk));
	jdff dff_B_5TX5zvkd6_2(.din(w_dff_B_0BatgX1U8_2),.dout(w_dff_B_5TX5zvkd6_2),.clk(gclk));
	jdff dff_B_poBBREZb0_2(.din(w_dff_B_5TX5zvkd6_2),.dout(w_dff_B_poBBREZb0_2),.clk(gclk));
	jdff dff_B_bsSzjpNN0_2(.din(w_dff_B_poBBREZb0_2),.dout(w_dff_B_bsSzjpNN0_2),.clk(gclk));
	jdff dff_B_EXJcq01N7_2(.din(w_dff_B_bsSzjpNN0_2),.dout(w_dff_B_EXJcq01N7_2),.clk(gclk));
	jdff dff_B_kctEHTof3_2(.din(w_dff_B_EXJcq01N7_2),.dout(w_dff_B_kctEHTof3_2),.clk(gclk));
	jdff dff_B_TqhesGzM8_2(.din(w_dff_B_kctEHTof3_2),.dout(w_dff_B_TqhesGzM8_2),.clk(gclk));
	jdff dff_B_Q8XWme3d4_2(.din(w_dff_B_TqhesGzM8_2),.dout(w_dff_B_Q8XWme3d4_2),.clk(gclk));
	jdff dff_B_Y8OjuYp30_2(.din(w_dff_B_Q8XWme3d4_2),.dout(w_dff_B_Y8OjuYp30_2),.clk(gclk));
	jdff dff_B_0cS1Hx3N3_2(.din(n1117),.dout(w_dff_B_0cS1Hx3N3_2),.clk(gclk));
	jdff dff_B_bu33HQNV7_2(.din(w_dff_B_0cS1Hx3N3_2),.dout(w_dff_B_bu33HQNV7_2),.clk(gclk));
	jdff dff_B_fD5g9lbL1_1(.din(n1095),.dout(w_dff_B_fD5g9lbL1_1),.clk(gclk));
	jdff dff_B_MTQAPdOR2_2(.din(n996),.dout(w_dff_B_MTQAPdOR2_2),.clk(gclk));
	jdff dff_B_jtQ8Y7GX4_2(.din(w_dff_B_MTQAPdOR2_2),.dout(w_dff_B_jtQ8Y7GX4_2),.clk(gclk));
	jdff dff_B_10TE86aF9_2(.din(w_dff_B_jtQ8Y7GX4_2),.dout(w_dff_B_10TE86aF9_2),.clk(gclk));
	jdff dff_B_ncnuwJ2E3_2(.din(w_dff_B_10TE86aF9_2),.dout(w_dff_B_ncnuwJ2E3_2),.clk(gclk));
	jdff dff_B_bzuIbQoh6_2(.din(w_dff_B_ncnuwJ2E3_2),.dout(w_dff_B_bzuIbQoh6_2),.clk(gclk));
	jdff dff_B_21e51WDS9_2(.din(w_dff_B_bzuIbQoh6_2),.dout(w_dff_B_21e51WDS9_2),.clk(gclk));
	jdff dff_B_ERTz4txs2_2(.din(w_dff_B_21e51WDS9_2),.dout(w_dff_B_ERTz4txs2_2),.clk(gclk));
	jdff dff_B_VxRWLuUO7_2(.din(w_dff_B_ERTz4txs2_2),.dout(w_dff_B_VxRWLuUO7_2),.clk(gclk));
	jdff dff_B_O1ZusvBL0_2(.din(w_dff_B_VxRWLuUO7_2),.dout(w_dff_B_O1ZusvBL0_2),.clk(gclk));
	jdff dff_B_TDCgQw3H6_2(.din(w_dff_B_O1ZusvBL0_2),.dout(w_dff_B_TDCgQw3H6_2),.clk(gclk));
	jdff dff_B_9XHbzvvr1_2(.din(w_dff_B_TDCgQw3H6_2),.dout(w_dff_B_9XHbzvvr1_2),.clk(gclk));
	jdff dff_B_chRGbMx43_2(.din(w_dff_B_9XHbzvvr1_2),.dout(w_dff_B_chRGbMx43_2),.clk(gclk));
	jdff dff_B_a4v49fP78_2(.din(n1012),.dout(w_dff_B_a4v49fP78_2),.clk(gclk));
	jdff dff_B_wXiLleDA8_2(.din(w_dff_B_a4v49fP78_2),.dout(w_dff_B_wXiLleDA8_2),.clk(gclk));
	jdff dff_B_UFwAyNCv0_1(.din(n997),.dout(w_dff_B_UFwAyNCv0_1),.clk(gclk));
	jdff dff_B_MEHfKbew9_2(.din(n891),.dout(w_dff_B_MEHfKbew9_2),.clk(gclk));
	jdff dff_B_LrNxf9oc7_2(.din(w_dff_B_MEHfKbew9_2),.dout(w_dff_B_LrNxf9oc7_2),.clk(gclk));
	jdff dff_B_EGze31uY3_2(.din(w_dff_B_LrNxf9oc7_2),.dout(w_dff_B_EGze31uY3_2),.clk(gclk));
	jdff dff_B_X647aHxM6_2(.din(w_dff_B_EGze31uY3_2),.dout(w_dff_B_X647aHxM6_2),.clk(gclk));
	jdff dff_B_MSQ59Pwh8_2(.din(w_dff_B_X647aHxM6_2),.dout(w_dff_B_MSQ59Pwh8_2),.clk(gclk));
	jdff dff_B_RuXvByrj7_2(.din(w_dff_B_MSQ59Pwh8_2),.dout(w_dff_B_RuXvByrj7_2),.clk(gclk));
	jdff dff_B_Ps3ZqFUD9_2(.din(w_dff_B_RuXvByrj7_2),.dout(w_dff_B_Ps3ZqFUD9_2),.clk(gclk));
	jdff dff_B_f3mfKWtz7_2(.din(w_dff_B_Ps3ZqFUD9_2),.dout(w_dff_B_f3mfKWtz7_2),.clk(gclk));
	jdff dff_B_l1f4Eccm7_2(.din(w_dff_B_f3mfKWtz7_2),.dout(w_dff_B_l1f4Eccm7_2),.clk(gclk));
	jdff dff_B_XzPR8iDa5_2(.din(n907),.dout(w_dff_B_XzPR8iDa5_2),.clk(gclk));
	jdff dff_B_AJXfXcpy5_2(.din(w_dff_B_XzPR8iDa5_2),.dout(w_dff_B_AJXfXcpy5_2),.clk(gclk));
	jdff dff_B_RKXxBQcS6_2(.din(w_dff_B_AJXfXcpy5_2),.dout(w_dff_B_RKXxBQcS6_2),.clk(gclk));
	jdff dff_B_VCOEMQuA2_1(.din(n892),.dout(w_dff_B_VCOEMQuA2_1),.clk(gclk));
	jdff dff_B_yqtwYyqE3_1(.din(w_dff_B_VCOEMQuA2_1),.dout(w_dff_B_yqtwYyqE3_1),.clk(gclk));
	jdff dff_B_oh5YNsE37_1(.din(w_dff_B_yqtwYyqE3_1),.dout(w_dff_B_oh5YNsE37_1),.clk(gclk));
	jdff dff_B_Fnn0jdrm6_1(.din(w_dff_B_oh5YNsE37_1),.dout(w_dff_B_Fnn0jdrm6_1),.clk(gclk));
	jdff dff_B_A27aPuPb3_1(.din(w_dff_B_Fnn0jdrm6_1),.dout(w_dff_B_A27aPuPb3_1),.clk(gclk));
	jdff dff_B_t0DlR4tB3_1(.din(w_dff_B_A27aPuPb3_1),.dout(w_dff_B_t0DlR4tB3_1),.clk(gclk));
	jdff dff_B_wIvBc2Ns2_0(.din(n801),.dout(w_dff_B_wIvBc2Ns2_0),.clk(gclk));
	jdff dff_B_zSHMYozx7_0(.din(w_dff_B_wIvBc2Ns2_0),.dout(w_dff_B_zSHMYozx7_0),.clk(gclk));
	jdff dff_A_p4yOhTTZ4_0(.dout(w_n800_0[0]),.din(w_dff_A_p4yOhTTZ4_0),.clk(gclk));
	jdff dff_A_MqQUNCDP0_0(.dout(w_dff_A_p4yOhTTZ4_0),.din(w_dff_A_MqQUNCDP0_0),.clk(gclk));
	jdff dff_A_gsSunOMy6_0(.dout(w_dff_A_MqQUNCDP0_0),.din(w_dff_A_gsSunOMy6_0),.clk(gclk));
	jdff dff_B_mzYTa5E69_1(.din(n794),.dout(w_dff_B_mzYTa5E69_1),.clk(gclk));
	jdff dff_A_xi5AQlVt6_0(.dout(w_n698_0[0]),.din(w_dff_A_xi5AQlVt6_0),.clk(gclk));
	jdff dff_A_MZXWqFtS9_1(.dout(w_n698_0[1]),.din(w_dff_A_MZXWqFtS9_1),.clk(gclk));
	jdff dff_A_UfhNzngE2_1(.dout(w_dff_A_MZXWqFtS9_1),.din(w_dff_A_UfhNzngE2_1),.clk(gclk));
	jdff dff_A_my0qZSVl3_1(.dout(w_n792_0[1]),.din(w_dff_A_my0qZSVl3_1),.clk(gclk));
	jdff dff_A_hE7lVLGO5_1(.dout(w_dff_A_my0qZSVl3_1),.din(w_dff_A_hE7lVLGO5_1),.clk(gclk));
	jdff dff_A_71TKbdsM7_1(.dout(w_dff_A_hE7lVLGO5_1),.din(w_dff_A_71TKbdsM7_1),.clk(gclk));
	jdff dff_A_DKvQaQ6L6_1(.dout(w_dff_A_71TKbdsM7_1),.din(w_dff_A_DKvQaQ6L6_1),.clk(gclk));
	jdff dff_A_LauM8jeY5_1(.dout(w_dff_A_DKvQaQ6L6_1),.din(w_dff_A_LauM8jeY5_1),.clk(gclk));
	jdff dff_A_AW1PADH56_1(.dout(w_dff_A_LauM8jeY5_1),.din(w_dff_A_AW1PADH56_1),.clk(gclk));
	jdff dff_B_081Xrddf4_1(.din(n1843),.dout(w_dff_B_081Xrddf4_1),.clk(gclk));
	jdff dff_B_PELpkZGR6_1(.din(n1830),.dout(w_dff_B_PELpkZGR6_1),.clk(gclk));
	jdff dff_B_UPlWjVfl7_1(.din(w_dff_B_PELpkZGR6_1),.dout(w_dff_B_UPlWjVfl7_1),.clk(gclk));
	jdff dff_B_5v7Cwybu6_2(.din(n1829),.dout(w_dff_B_5v7Cwybu6_2),.clk(gclk));
	jdff dff_B_f1OG74Oz3_2(.din(w_dff_B_5v7Cwybu6_2),.dout(w_dff_B_f1OG74Oz3_2),.clk(gclk));
	jdff dff_B_qdN04MBe9_2(.din(w_dff_B_f1OG74Oz3_2),.dout(w_dff_B_qdN04MBe9_2),.clk(gclk));
	jdff dff_B_3dV18AZc7_2(.din(w_dff_B_qdN04MBe9_2),.dout(w_dff_B_3dV18AZc7_2),.clk(gclk));
	jdff dff_B_J0pmaD6N1_2(.din(w_dff_B_3dV18AZc7_2),.dout(w_dff_B_J0pmaD6N1_2),.clk(gclk));
	jdff dff_B_ZMIiXKNE4_2(.din(w_dff_B_J0pmaD6N1_2),.dout(w_dff_B_ZMIiXKNE4_2),.clk(gclk));
	jdff dff_B_r5Zq5X2H7_2(.din(w_dff_B_ZMIiXKNE4_2),.dout(w_dff_B_r5Zq5X2H7_2),.clk(gclk));
	jdff dff_B_frcr2BQ58_2(.din(w_dff_B_r5Zq5X2H7_2),.dout(w_dff_B_frcr2BQ58_2),.clk(gclk));
	jdff dff_B_6VN7LgEd2_2(.din(w_dff_B_frcr2BQ58_2),.dout(w_dff_B_6VN7LgEd2_2),.clk(gclk));
	jdff dff_B_mPJKC1FO5_2(.din(w_dff_B_6VN7LgEd2_2),.dout(w_dff_B_mPJKC1FO5_2),.clk(gclk));
	jdff dff_B_3ufNL6YE1_2(.din(w_dff_B_mPJKC1FO5_2),.dout(w_dff_B_3ufNL6YE1_2),.clk(gclk));
	jdff dff_B_G0gLPMY86_2(.din(w_dff_B_3ufNL6YE1_2),.dout(w_dff_B_G0gLPMY86_2),.clk(gclk));
	jdff dff_B_CMuiVO743_2(.din(w_dff_B_G0gLPMY86_2),.dout(w_dff_B_CMuiVO743_2),.clk(gclk));
	jdff dff_B_jbWSueBK0_2(.din(w_dff_B_CMuiVO743_2),.dout(w_dff_B_jbWSueBK0_2),.clk(gclk));
	jdff dff_B_rnx8ihFa0_2(.din(w_dff_B_jbWSueBK0_2),.dout(w_dff_B_rnx8ihFa0_2),.clk(gclk));
	jdff dff_B_lkEdDCNd5_2(.din(w_dff_B_rnx8ihFa0_2),.dout(w_dff_B_lkEdDCNd5_2),.clk(gclk));
	jdff dff_B_5Kqjs0H78_2(.din(w_dff_B_lkEdDCNd5_2),.dout(w_dff_B_5Kqjs0H78_2),.clk(gclk));
	jdff dff_B_yTlv3t160_2(.din(w_dff_B_5Kqjs0H78_2),.dout(w_dff_B_yTlv3t160_2),.clk(gclk));
	jdff dff_B_eP7KzkAU1_2(.din(w_dff_B_yTlv3t160_2),.dout(w_dff_B_eP7KzkAU1_2),.clk(gclk));
	jdff dff_B_zHfpANWv3_2(.din(w_dff_B_eP7KzkAU1_2),.dout(w_dff_B_zHfpANWv3_2),.clk(gclk));
	jdff dff_B_2VKmsVJD1_2(.din(w_dff_B_zHfpANWv3_2),.dout(w_dff_B_2VKmsVJD1_2),.clk(gclk));
	jdff dff_B_pDgrJjwb8_2(.din(w_dff_B_2VKmsVJD1_2),.dout(w_dff_B_pDgrJjwb8_2),.clk(gclk));
	jdff dff_B_NCEZoyRg9_2(.din(w_dff_B_pDgrJjwb8_2),.dout(w_dff_B_NCEZoyRg9_2),.clk(gclk));
	jdff dff_B_hpRTIMEf5_2(.din(w_dff_B_NCEZoyRg9_2),.dout(w_dff_B_hpRTIMEf5_2),.clk(gclk));
	jdff dff_B_uw15CJv09_2(.din(w_dff_B_hpRTIMEf5_2),.dout(w_dff_B_uw15CJv09_2),.clk(gclk));
	jdff dff_B_7SqJUegL5_2(.din(w_dff_B_uw15CJv09_2),.dout(w_dff_B_7SqJUegL5_2),.clk(gclk));
	jdff dff_B_fsTo1ptP8_2(.din(w_dff_B_7SqJUegL5_2),.dout(w_dff_B_fsTo1ptP8_2),.clk(gclk));
	jdff dff_B_pFdLz4Cc4_2(.din(w_dff_B_fsTo1ptP8_2),.dout(w_dff_B_pFdLz4Cc4_2),.clk(gclk));
	jdff dff_B_nGEyyGEa8_2(.din(w_dff_B_pFdLz4Cc4_2),.dout(w_dff_B_nGEyyGEa8_2),.clk(gclk));
	jdff dff_B_kkk8bx8y7_2(.din(w_dff_B_nGEyyGEa8_2),.dout(w_dff_B_kkk8bx8y7_2),.clk(gclk));
	jdff dff_B_oXHz3RBJ8_2(.din(w_dff_B_kkk8bx8y7_2),.dout(w_dff_B_oXHz3RBJ8_2),.clk(gclk));
	jdff dff_B_4cTCC7kT1_2(.din(w_dff_B_oXHz3RBJ8_2),.dout(w_dff_B_4cTCC7kT1_2),.clk(gclk));
	jdff dff_B_pSZ7TYnB4_2(.din(w_dff_B_4cTCC7kT1_2),.dout(w_dff_B_pSZ7TYnB4_2),.clk(gclk));
	jdff dff_B_pB83XQWe5_2(.din(w_dff_B_pSZ7TYnB4_2),.dout(w_dff_B_pB83XQWe5_2),.clk(gclk));
	jdff dff_B_d64f9uoR8_2(.din(w_dff_B_pB83XQWe5_2),.dout(w_dff_B_d64f9uoR8_2),.clk(gclk));
	jdff dff_B_U1DOPePd6_2(.din(w_dff_B_d64f9uoR8_2),.dout(w_dff_B_U1DOPePd6_2),.clk(gclk));
	jdff dff_B_LMq2bu8i3_2(.din(w_dff_B_U1DOPePd6_2),.dout(w_dff_B_LMq2bu8i3_2),.clk(gclk));
	jdff dff_B_TcZANVD60_2(.din(w_dff_B_LMq2bu8i3_2),.dout(w_dff_B_TcZANVD60_2),.clk(gclk));
	jdff dff_B_tcfZoO6z3_2(.din(w_dff_B_TcZANVD60_2),.dout(w_dff_B_tcfZoO6z3_2),.clk(gclk));
	jdff dff_B_S2lf0fWp3_2(.din(w_dff_B_tcfZoO6z3_2),.dout(w_dff_B_S2lf0fWp3_2),.clk(gclk));
	jdff dff_B_3CAGL5ax6_2(.din(w_dff_B_S2lf0fWp3_2),.dout(w_dff_B_3CAGL5ax6_2),.clk(gclk));
	jdff dff_B_ljXJ2ynj2_2(.din(w_dff_B_3CAGL5ax6_2),.dout(w_dff_B_ljXJ2ynj2_2),.clk(gclk));
	jdff dff_B_665JCJru3_2(.din(w_dff_B_ljXJ2ynj2_2),.dout(w_dff_B_665JCJru3_2),.clk(gclk));
	jdff dff_B_zOTBCFUP3_2(.din(w_dff_B_665JCJru3_2),.dout(w_dff_B_zOTBCFUP3_2),.clk(gclk));
	jdff dff_B_CVk7hsi26_2(.din(w_dff_B_zOTBCFUP3_2),.dout(w_dff_B_CVk7hsi26_2),.clk(gclk));
	jdff dff_B_pddNHisA9_2(.din(w_dff_B_CVk7hsi26_2),.dout(w_dff_B_pddNHisA9_2),.clk(gclk));
	jdff dff_B_OsphWy6H8_2(.din(w_dff_B_pddNHisA9_2),.dout(w_dff_B_OsphWy6H8_2),.clk(gclk));
	jdff dff_B_lhckDvac9_2(.din(w_dff_B_OsphWy6H8_2),.dout(w_dff_B_lhckDvac9_2),.clk(gclk));
	jdff dff_B_mWv5pILD7_2(.din(w_dff_B_lhckDvac9_2),.dout(w_dff_B_mWv5pILD7_2),.clk(gclk));
	jdff dff_B_nBofrBcW4_2(.din(w_dff_B_mWv5pILD7_2),.dout(w_dff_B_nBofrBcW4_2),.clk(gclk));
	jdff dff_B_bSDy59976_2(.din(w_dff_B_nBofrBcW4_2),.dout(w_dff_B_bSDy59976_2),.clk(gclk));
	jdff dff_B_JLr79cM30_2(.din(w_dff_B_bSDy59976_2),.dout(w_dff_B_JLr79cM30_2),.clk(gclk));
	jdff dff_B_T26zHkVu5_2(.din(w_dff_B_JLr79cM30_2),.dout(w_dff_B_T26zHkVu5_2),.clk(gclk));
	jdff dff_B_r62pziid6_2(.din(w_dff_B_T26zHkVu5_2),.dout(w_dff_B_r62pziid6_2),.clk(gclk));
	jdff dff_B_dLkIvAW73_2(.din(w_dff_B_r62pziid6_2),.dout(w_dff_B_dLkIvAW73_2),.clk(gclk));
	jdff dff_B_DWU7mLRu5_2(.din(w_dff_B_dLkIvAW73_2),.dout(w_dff_B_DWU7mLRu5_2),.clk(gclk));
	jdff dff_B_v6oMuJO42_2(.din(n1828),.dout(w_dff_B_v6oMuJO42_2),.clk(gclk));
	jdff dff_B_Rm6MhEQf4_2(.din(w_dff_B_v6oMuJO42_2),.dout(w_dff_B_Rm6MhEQf4_2),.clk(gclk));
	jdff dff_B_HtVBoJV96_2(.din(w_dff_B_Rm6MhEQf4_2),.dout(w_dff_B_HtVBoJV96_2),.clk(gclk));
	jdff dff_B_PVvCbUy14_2(.din(w_dff_B_HtVBoJV96_2),.dout(w_dff_B_PVvCbUy14_2),.clk(gclk));
	jdff dff_B_KmfJV7hs9_2(.din(w_dff_B_PVvCbUy14_2),.dout(w_dff_B_KmfJV7hs9_2),.clk(gclk));
	jdff dff_B_kXzCZgBD6_2(.din(w_dff_B_KmfJV7hs9_2),.dout(w_dff_B_kXzCZgBD6_2),.clk(gclk));
	jdff dff_B_fwUUWTIM0_2(.din(w_dff_B_kXzCZgBD6_2),.dout(w_dff_B_fwUUWTIM0_2),.clk(gclk));
	jdff dff_B_OHFUtWk27_2(.din(w_dff_B_fwUUWTIM0_2),.dout(w_dff_B_OHFUtWk27_2),.clk(gclk));
	jdff dff_B_Of0j8XoX2_2(.din(w_dff_B_OHFUtWk27_2),.dout(w_dff_B_Of0j8XoX2_2),.clk(gclk));
	jdff dff_B_JORh3Z2K5_2(.din(w_dff_B_Of0j8XoX2_2),.dout(w_dff_B_JORh3Z2K5_2),.clk(gclk));
	jdff dff_B_kKn3i41J6_2(.din(w_dff_B_JORh3Z2K5_2),.dout(w_dff_B_kKn3i41J6_2),.clk(gclk));
	jdff dff_B_NkkRH9ZQ8_2(.din(w_dff_B_kKn3i41J6_2),.dout(w_dff_B_NkkRH9ZQ8_2),.clk(gclk));
	jdff dff_B_2GkZ8hpD9_2(.din(w_dff_B_NkkRH9ZQ8_2),.dout(w_dff_B_2GkZ8hpD9_2),.clk(gclk));
	jdff dff_B_eujWYkjA4_2(.din(w_dff_B_2GkZ8hpD9_2),.dout(w_dff_B_eujWYkjA4_2),.clk(gclk));
	jdff dff_B_KRbT3pt91_2(.din(w_dff_B_eujWYkjA4_2),.dout(w_dff_B_KRbT3pt91_2),.clk(gclk));
	jdff dff_B_JhzzV94S2_2(.din(w_dff_B_KRbT3pt91_2),.dout(w_dff_B_JhzzV94S2_2),.clk(gclk));
	jdff dff_B_hz98RGvz8_2(.din(w_dff_B_JhzzV94S2_2),.dout(w_dff_B_hz98RGvz8_2),.clk(gclk));
	jdff dff_B_08fJ1fTh5_2(.din(w_dff_B_hz98RGvz8_2),.dout(w_dff_B_08fJ1fTh5_2),.clk(gclk));
	jdff dff_B_d6Hgq5M18_2(.din(w_dff_B_08fJ1fTh5_2),.dout(w_dff_B_d6Hgq5M18_2),.clk(gclk));
	jdff dff_B_f0vzKlBO2_2(.din(w_dff_B_d6Hgq5M18_2),.dout(w_dff_B_f0vzKlBO2_2),.clk(gclk));
	jdff dff_B_cZyrIjHG1_2(.din(w_dff_B_f0vzKlBO2_2),.dout(w_dff_B_cZyrIjHG1_2),.clk(gclk));
	jdff dff_B_KbZiRDfg4_2(.din(w_dff_B_cZyrIjHG1_2),.dout(w_dff_B_KbZiRDfg4_2),.clk(gclk));
	jdff dff_B_NSWvBMA29_2(.din(w_dff_B_KbZiRDfg4_2),.dout(w_dff_B_NSWvBMA29_2),.clk(gclk));
	jdff dff_B_1oX7jY9N5_2(.din(w_dff_B_NSWvBMA29_2),.dout(w_dff_B_1oX7jY9N5_2),.clk(gclk));
	jdff dff_B_ajKvOeor9_2(.din(w_dff_B_1oX7jY9N5_2),.dout(w_dff_B_ajKvOeor9_2),.clk(gclk));
	jdff dff_B_hRclBnZW3_2(.din(w_dff_B_ajKvOeor9_2),.dout(w_dff_B_hRclBnZW3_2),.clk(gclk));
	jdff dff_B_vlt6mRqO8_2(.din(w_dff_B_hRclBnZW3_2),.dout(w_dff_B_vlt6mRqO8_2),.clk(gclk));
	jdff dff_B_CQ4DIJ6n0_2(.din(w_dff_B_vlt6mRqO8_2),.dout(w_dff_B_CQ4DIJ6n0_2),.clk(gclk));
	jdff dff_B_O0ZoKvlz7_2(.din(w_dff_B_CQ4DIJ6n0_2),.dout(w_dff_B_O0ZoKvlz7_2),.clk(gclk));
	jdff dff_B_xMIDyI3U4_2(.din(w_dff_B_O0ZoKvlz7_2),.dout(w_dff_B_xMIDyI3U4_2),.clk(gclk));
	jdff dff_B_qLMiArfw7_2(.din(w_dff_B_xMIDyI3U4_2),.dout(w_dff_B_qLMiArfw7_2),.clk(gclk));
	jdff dff_B_zwtG02J54_2(.din(w_dff_B_qLMiArfw7_2),.dout(w_dff_B_zwtG02J54_2),.clk(gclk));
	jdff dff_B_YaN0fOWd5_2(.din(w_dff_B_zwtG02J54_2),.dout(w_dff_B_YaN0fOWd5_2),.clk(gclk));
	jdff dff_B_lysFEHkd7_2(.din(w_dff_B_YaN0fOWd5_2),.dout(w_dff_B_lysFEHkd7_2),.clk(gclk));
	jdff dff_B_VMaSCxnd1_2(.din(w_dff_B_lysFEHkd7_2),.dout(w_dff_B_VMaSCxnd1_2),.clk(gclk));
	jdff dff_B_pVXkeNhE4_2(.din(w_dff_B_VMaSCxnd1_2),.dout(w_dff_B_pVXkeNhE4_2),.clk(gclk));
	jdff dff_B_IuMVvph68_2(.din(w_dff_B_pVXkeNhE4_2),.dout(w_dff_B_IuMVvph68_2),.clk(gclk));
	jdff dff_B_GekZBews5_2(.din(w_dff_B_IuMVvph68_2),.dout(w_dff_B_GekZBews5_2),.clk(gclk));
	jdff dff_B_fEGvgOtp1_2(.din(w_dff_B_GekZBews5_2),.dout(w_dff_B_fEGvgOtp1_2),.clk(gclk));
	jdff dff_B_UapzPCYt3_2(.din(w_dff_B_fEGvgOtp1_2),.dout(w_dff_B_UapzPCYt3_2),.clk(gclk));
	jdff dff_B_0DBgrgZV6_2(.din(w_dff_B_UapzPCYt3_2),.dout(w_dff_B_0DBgrgZV6_2),.clk(gclk));
	jdff dff_B_Ui2zdgbZ5_2(.din(w_dff_B_0DBgrgZV6_2),.dout(w_dff_B_Ui2zdgbZ5_2),.clk(gclk));
	jdff dff_B_robcFZAe6_2(.din(w_dff_B_Ui2zdgbZ5_2),.dout(w_dff_B_robcFZAe6_2),.clk(gclk));
	jdff dff_B_3ITGfKaW9_2(.din(w_dff_B_robcFZAe6_2),.dout(w_dff_B_3ITGfKaW9_2),.clk(gclk));
	jdff dff_B_BDOogQE10_2(.din(w_dff_B_3ITGfKaW9_2),.dout(w_dff_B_BDOogQE10_2),.clk(gclk));
	jdff dff_B_6B4Ao2BR9_2(.din(w_dff_B_BDOogQE10_2),.dout(w_dff_B_6B4Ao2BR9_2),.clk(gclk));
	jdff dff_B_H35qfwNg9_2(.din(w_dff_B_6B4Ao2BR9_2),.dout(w_dff_B_H35qfwNg9_2),.clk(gclk));
	jdff dff_B_FyEso6WK7_2(.din(w_dff_B_H35qfwNg9_2),.dout(w_dff_B_FyEso6WK7_2),.clk(gclk));
	jdff dff_B_yBtzNJ2J0_2(.din(w_dff_B_FyEso6WK7_2),.dout(w_dff_B_yBtzNJ2J0_2),.clk(gclk));
	jdff dff_B_S0RrCZ7l0_2(.din(w_dff_B_yBtzNJ2J0_2),.dout(w_dff_B_S0RrCZ7l0_2),.clk(gclk));
	jdff dff_B_ylm2zTC42_2(.din(w_dff_B_S0RrCZ7l0_2),.dout(w_dff_B_ylm2zTC42_2),.clk(gclk));
	jdff dff_B_jTuo7NQI0_2(.din(w_dff_B_ylm2zTC42_2),.dout(w_dff_B_jTuo7NQI0_2),.clk(gclk));
	jdff dff_B_he1rIc3I5_2(.din(w_dff_B_jTuo7NQI0_2),.dout(w_dff_B_he1rIc3I5_2),.clk(gclk));
	jdff dff_B_836wzKpd8_2(.din(w_dff_B_he1rIc3I5_2),.dout(w_dff_B_836wzKpd8_2),.clk(gclk));
	jdff dff_B_7dGqTvEF8_2(.din(w_dff_B_836wzKpd8_2),.dout(w_dff_B_7dGqTvEF8_2),.clk(gclk));
	jdff dff_B_3QhjI9FW5_2(.din(w_dff_B_7dGqTvEF8_2),.dout(w_dff_B_3QhjI9FW5_2),.clk(gclk));
	jdff dff_B_KwmOwAnj1_2(.din(w_dff_B_3QhjI9FW5_2),.dout(w_dff_B_KwmOwAnj1_2),.clk(gclk));
	jdff dff_B_fosja2Hu4_2(.din(w_dff_B_KwmOwAnj1_2),.dout(w_dff_B_fosja2Hu4_2),.clk(gclk));
	jdff dff_A_aQrQ35x31_1(.dout(w_n1827_0[1]),.din(w_dff_A_aQrQ35x31_1),.clk(gclk));
	jdff dff_B_C92hqvgL8_1(.din(n1825),.dout(w_dff_B_C92hqvgL8_1),.clk(gclk));
	jdff dff_B_grHPxLff2_2(.din(n1803),.dout(w_dff_B_grHPxLff2_2),.clk(gclk));
	jdff dff_B_2t0uBdcP6_2(.din(w_dff_B_grHPxLff2_2),.dout(w_dff_B_2t0uBdcP6_2),.clk(gclk));
	jdff dff_B_Agovedgy2_2(.din(w_dff_B_2t0uBdcP6_2),.dout(w_dff_B_Agovedgy2_2),.clk(gclk));
	jdff dff_B_XnFqnkd55_2(.din(w_dff_B_Agovedgy2_2),.dout(w_dff_B_XnFqnkd55_2),.clk(gclk));
	jdff dff_B_nRECSmre3_2(.din(w_dff_B_XnFqnkd55_2),.dout(w_dff_B_nRECSmre3_2),.clk(gclk));
	jdff dff_B_Gbg1xO0r7_2(.din(w_dff_B_nRECSmre3_2),.dout(w_dff_B_Gbg1xO0r7_2),.clk(gclk));
	jdff dff_B_dLnvZYU03_2(.din(w_dff_B_Gbg1xO0r7_2),.dout(w_dff_B_dLnvZYU03_2),.clk(gclk));
	jdff dff_B_mGjCruk43_2(.din(w_dff_B_dLnvZYU03_2),.dout(w_dff_B_mGjCruk43_2),.clk(gclk));
	jdff dff_B_Ds66a7Zk9_2(.din(w_dff_B_mGjCruk43_2),.dout(w_dff_B_Ds66a7Zk9_2),.clk(gclk));
	jdff dff_B_4NHEN7pu4_2(.din(w_dff_B_Ds66a7Zk9_2),.dout(w_dff_B_4NHEN7pu4_2),.clk(gclk));
	jdff dff_B_pzRuHHUT5_2(.din(w_dff_B_4NHEN7pu4_2),.dout(w_dff_B_pzRuHHUT5_2),.clk(gclk));
	jdff dff_B_dIIfp8xh6_2(.din(w_dff_B_pzRuHHUT5_2),.dout(w_dff_B_dIIfp8xh6_2),.clk(gclk));
	jdff dff_B_jWvrj71G7_2(.din(w_dff_B_dIIfp8xh6_2),.dout(w_dff_B_jWvrj71G7_2),.clk(gclk));
	jdff dff_B_Ja1ABzjF7_2(.din(w_dff_B_jWvrj71G7_2),.dout(w_dff_B_Ja1ABzjF7_2),.clk(gclk));
	jdff dff_B_5CoJBZyy4_2(.din(w_dff_B_Ja1ABzjF7_2),.dout(w_dff_B_5CoJBZyy4_2),.clk(gclk));
	jdff dff_B_S15C6HcH4_2(.din(w_dff_B_5CoJBZyy4_2),.dout(w_dff_B_S15C6HcH4_2),.clk(gclk));
	jdff dff_B_lyuZzVzM8_2(.din(w_dff_B_S15C6HcH4_2),.dout(w_dff_B_lyuZzVzM8_2),.clk(gclk));
	jdff dff_B_yPAyk9lF2_2(.din(w_dff_B_lyuZzVzM8_2),.dout(w_dff_B_yPAyk9lF2_2),.clk(gclk));
	jdff dff_B_lk2w28Fo1_2(.din(w_dff_B_yPAyk9lF2_2),.dout(w_dff_B_lk2w28Fo1_2),.clk(gclk));
	jdff dff_B_sV5fIFD98_2(.din(w_dff_B_lk2w28Fo1_2),.dout(w_dff_B_sV5fIFD98_2),.clk(gclk));
	jdff dff_B_6zrt42610_2(.din(w_dff_B_sV5fIFD98_2),.dout(w_dff_B_6zrt42610_2),.clk(gclk));
	jdff dff_B_jtnQ4U8k3_2(.din(w_dff_B_6zrt42610_2),.dout(w_dff_B_jtnQ4U8k3_2),.clk(gclk));
	jdff dff_B_SZvDbafQ3_2(.din(w_dff_B_jtnQ4U8k3_2),.dout(w_dff_B_SZvDbafQ3_2),.clk(gclk));
	jdff dff_B_SDNxZN1g3_2(.din(w_dff_B_SZvDbafQ3_2),.dout(w_dff_B_SDNxZN1g3_2),.clk(gclk));
	jdff dff_B_dhSrtEEv9_2(.din(w_dff_B_SDNxZN1g3_2),.dout(w_dff_B_dhSrtEEv9_2),.clk(gclk));
	jdff dff_B_IBTHqlCX4_2(.din(w_dff_B_dhSrtEEv9_2),.dout(w_dff_B_IBTHqlCX4_2),.clk(gclk));
	jdff dff_B_FYvFNWhv6_2(.din(w_dff_B_IBTHqlCX4_2),.dout(w_dff_B_FYvFNWhv6_2),.clk(gclk));
	jdff dff_B_NPGUVlxb0_2(.din(w_dff_B_FYvFNWhv6_2),.dout(w_dff_B_NPGUVlxb0_2),.clk(gclk));
	jdff dff_B_MWl8q4I98_2(.din(w_dff_B_NPGUVlxb0_2),.dout(w_dff_B_MWl8q4I98_2),.clk(gclk));
	jdff dff_B_kMgM8Tg71_2(.din(w_dff_B_MWl8q4I98_2),.dout(w_dff_B_kMgM8Tg71_2),.clk(gclk));
	jdff dff_B_LSOUMlfv1_2(.din(w_dff_B_kMgM8Tg71_2),.dout(w_dff_B_LSOUMlfv1_2),.clk(gclk));
	jdff dff_B_G4BYq1t22_2(.din(w_dff_B_LSOUMlfv1_2),.dout(w_dff_B_G4BYq1t22_2),.clk(gclk));
	jdff dff_B_StOvbnaR9_2(.din(w_dff_B_G4BYq1t22_2),.dout(w_dff_B_StOvbnaR9_2),.clk(gclk));
	jdff dff_B_or6V7SCe8_2(.din(w_dff_B_StOvbnaR9_2),.dout(w_dff_B_or6V7SCe8_2),.clk(gclk));
	jdff dff_B_5XqyY2eQ6_2(.din(w_dff_B_or6V7SCe8_2),.dout(w_dff_B_5XqyY2eQ6_2),.clk(gclk));
	jdff dff_B_1dDZwQAr9_2(.din(w_dff_B_5XqyY2eQ6_2),.dout(w_dff_B_1dDZwQAr9_2),.clk(gclk));
	jdff dff_B_sD0CfKGj3_2(.din(w_dff_B_1dDZwQAr9_2),.dout(w_dff_B_sD0CfKGj3_2),.clk(gclk));
	jdff dff_B_YjL7x2uR4_2(.din(w_dff_B_sD0CfKGj3_2),.dout(w_dff_B_YjL7x2uR4_2),.clk(gclk));
	jdff dff_B_uAUcWnL02_2(.din(w_dff_B_YjL7x2uR4_2),.dout(w_dff_B_uAUcWnL02_2),.clk(gclk));
	jdff dff_B_vRsIJSpv7_2(.din(w_dff_B_uAUcWnL02_2),.dout(w_dff_B_vRsIJSpv7_2),.clk(gclk));
	jdff dff_B_42mpVIHe2_2(.din(w_dff_B_vRsIJSpv7_2),.dout(w_dff_B_42mpVIHe2_2),.clk(gclk));
	jdff dff_B_yl0REqCP3_2(.din(w_dff_B_42mpVIHe2_2),.dout(w_dff_B_yl0REqCP3_2),.clk(gclk));
	jdff dff_B_CvoZ9Ung1_2(.din(w_dff_B_yl0REqCP3_2),.dout(w_dff_B_CvoZ9Ung1_2),.clk(gclk));
	jdff dff_B_ml8z6I3A4_2(.din(w_dff_B_CvoZ9Ung1_2),.dout(w_dff_B_ml8z6I3A4_2),.clk(gclk));
	jdff dff_B_4blErXlR5_2(.din(w_dff_B_ml8z6I3A4_2),.dout(w_dff_B_4blErXlR5_2),.clk(gclk));
	jdff dff_B_7EkaFK5e0_2(.din(w_dff_B_4blErXlR5_2),.dout(w_dff_B_7EkaFK5e0_2),.clk(gclk));
	jdff dff_B_A1ZfeXeZ0_2(.din(w_dff_B_7EkaFK5e0_2),.dout(w_dff_B_A1ZfeXeZ0_2),.clk(gclk));
	jdff dff_B_U8JkEi1S5_2(.din(w_dff_B_A1ZfeXeZ0_2),.dout(w_dff_B_U8JkEi1S5_2),.clk(gclk));
	jdff dff_B_J7GcF8Kw5_2(.din(w_dff_B_U8JkEi1S5_2),.dout(w_dff_B_J7GcF8Kw5_2),.clk(gclk));
	jdff dff_B_woChbYS79_2(.din(w_dff_B_J7GcF8Kw5_2),.dout(w_dff_B_woChbYS79_2),.clk(gclk));
	jdff dff_B_EjCfjk3d5_2(.din(w_dff_B_woChbYS79_2),.dout(w_dff_B_EjCfjk3d5_2),.clk(gclk));
	jdff dff_B_kb8mRVRf4_2(.din(w_dff_B_EjCfjk3d5_2),.dout(w_dff_B_kb8mRVRf4_2),.clk(gclk));
	jdff dff_B_66jx00kP9_2(.din(w_dff_B_kb8mRVRf4_2),.dout(w_dff_B_66jx00kP9_2),.clk(gclk));
	jdff dff_B_p3eyB6Cd5_2(.din(w_dff_B_66jx00kP9_2),.dout(w_dff_B_p3eyB6Cd5_2),.clk(gclk));
	jdff dff_B_eIaXRKAC9_2(.din(w_dff_B_p3eyB6Cd5_2),.dout(w_dff_B_eIaXRKAC9_2),.clk(gclk));
	jdff dff_B_3ETeiOUN6_1(.din(n1809),.dout(w_dff_B_3ETeiOUN6_1),.clk(gclk));
	jdff dff_B_4p6E7E1O0_1(.din(w_dff_B_3ETeiOUN6_1),.dout(w_dff_B_4p6E7E1O0_1),.clk(gclk));
	jdff dff_B_r5DEL3wF3_2(.din(n1808),.dout(w_dff_B_r5DEL3wF3_2),.clk(gclk));
	jdff dff_B_41nrji832_2(.din(w_dff_B_r5DEL3wF3_2),.dout(w_dff_B_41nrji832_2),.clk(gclk));
	jdff dff_B_8F8cbYSV3_2(.din(w_dff_B_41nrji832_2),.dout(w_dff_B_8F8cbYSV3_2),.clk(gclk));
	jdff dff_B_BsFOJEvq2_2(.din(w_dff_B_8F8cbYSV3_2),.dout(w_dff_B_BsFOJEvq2_2),.clk(gclk));
	jdff dff_B_RMjv8qhD2_2(.din(w_dff_B_BsFOJEvq2_2),.dout(w_dff_B_RMjv8qhD2_2),.clk(gclk));
	jdff dff_B_Xefi5GXi6_2(.din(w_dff_B_RMjv8qhD2_2),.dout(w_dff_B_Xefi5GXi6_2),.clk(gclk));
	jdff dff_B_ZiS5HXpC5_2(.din(w_dff_B_Xefi5GXi6_2),.dout(w_dff_B_ZiS5HXpC5_2),.clk(gclk));
	jdff dff_B_UcpOn7Jw3_2(.din(w_dff_B_ZiS5HXpC5_2),.dout(w_dff_B_UcpOn7Jw3_2),.clk(gclk));
	jdff dff_B_GRDGAL5z3_2(.din(w_dff_B_UcpOn7Jw3_2),.dout(w_dff_B_GRDGAL5z3_2),.clk(gclk));
	jdff dff_B_DkiRuxjS4_2(.din(w_dff_B_GRDGAL5z3_2),.dout(w_dff_B_DkiRuxjS4_2),.clk(gclk));
	jdff dff_B_JmQDMNcD6_2(.din(w_dff_B_DkiRuxjS4_2),.dout(w_dff_B_JmQDMNcD6_2),.clk(gclk));
	jdff dff_B_40TCthHB3_2(.din(w_dff_B_JmQDMNcD6_2),.dout(w_dff_B_40TCthHB3_2),.clk(gclk));
	jdff dff_B_HLiXnyRE4_2(.din(w_dff_B_40TCthHB3_2),.dout(w_dff_B_HLiXnyRE4_2),.clk(gclk));
	jdff dff_B_J4o6ukSd5_2(.din(w_dff_B_HLiXnyRE4_2),.dout(w_dff_B_J4o6ukSd5_2),.clk(gclk));
	jdff dff_B_5NfzmMAL4_2(.din(w_dff_B_J4o6ukSd5_2),.dout(w_dff_B_5NfzmMAL4_2),.clk(gclk));
	jdff dff_B_bT8o41Ha4_2(.din(w_dff_B_5NfzmMAL4_2),.dout(w_dff_B_bT8o41Ha4_2),.clk(gclk));
	jdff dff_B_hCVkK3CI6_2(.din(w_dff_B_bT8o41Ha4_2),.dout(w_dff_B_hCVkK3CI6_2),.clk(gclk));
	jdff dff_B_Nn5HNoY04_2(.din(w_dff_B_hCVkK3CI6_2),.dout(w_dff_B_Nn5HNoY04_2),.clk(gclk));
	jdff dff_B_jGjPlxOJ2_2(.din(w_dff_B_Nn5HNoY04_2),.dout(w_dff_B_jGjPlxOJ2_2),.clk(gclk));
	jdff dff_B_sioFT1Gn2_2(.din(w_dff_B_jGjPlxOJ2_2),.dout(w_dff_B_sioFT1Gn2_2),.clk(gclk));
	jdff dff_B_s7w2bqc97_2(.din(w_dff_B_sioFT1Gn2_2),.dout(w_dff_B_s7w2bqc97_2),.clk(gclk));
	jdff dff_B_m5vN53pR8_2(.din(w_dff_B_s7w2bqc97_2),.dout(w_dff_B_m5vN53pR8_2),.clk(gclk));
	jdff dff_B_1ajmfdsi1_2(.din(w_dff_B_m5vN53pR8_2),.dout(w_dff_B_1ajmfdsi1_2),.clk(gclk));
	jdff dff_B_ZVb7hnVn9_2(.din(w_dff_B_1ajmfdsi1_2),.dout(w_dff_B_ZVb7hnVn9_2),.clk(gclk));
	jdff dff_B_kTg5F5Uw8_2(.din(w_dff_B_ZVb7hnVn9_2),.dout(w_dff_B_kTg5F5Uw8_2),.clk(gclk));
	jdff dff_B_BfAL3iO21_2(.din(w_dff_B_kTg5F5Uw8_2),.dout(w_dff_B_BfAL3iO21_2),.clk(gclk));
	jdff dff_B_vlYk47kL3_2(.din(w_dff_B_BfAL3iO21_2),.dout(w_dff_B_vlYk47kL3_2),.clk(gclk));
	jdff dff_B_m8yavwcg5_2(.din(w_dff_B_vlYk47kL3_2),.dout(w_dff_B_m8yavwcg5_2),.clk(gclk));
	jdff dff_B_HvUKYcwq5_2(.din(w_dff_B_m8yavwcg5_2),.dout(w_dff_B_HvUKYcwq5_2),.clk(gclk));
	jdff dff_B_mnqqvzLX5_2(.din(w_dff_B_HvUKYcwq5_2),.dout(w_dff_B_mnqqvzLX5_2),.clk(gclk));
	jdff dff_B_XJOE9A6E5_2(.din(w_dff_B_mnqqvzLX5_2),.dout(w_dff_B_XJOE9A6E5_2),.clk(gclk));
	jdff dff_B_PVsj90Kj4_2(.din(w_dff_B_XJOE9A6E5_2),.dout(w_dff_B_PVsj90Kj4_2),.clk(gclk));
	jdff dff_B_6B4ijnv61_2(.din(w_dff_B_PVsj90Kj4_2),.dout(w_dff_B_6B4ijnv61_2),.clk(gclk));
	jdff dff_B_JJ7eaP0L2_2(.din(w_dff_B_6B4ijnv61_2),.dout(w_dff_B_JJ7eaP0L2_2),.clk(gclk));
	jdff dff_B_OaljYqE97_2(.din(w_dff_B_JJ7eaP0L2_2),.dout(w_dff_B_OaljYqE97_2),.clk(gclk));
	jdff dff_B_Ydaoss7M1_2(.din(w_dff_B_OaljYqE97_2),.dout(w_dff_B_Ydaoss7M1_2),.clk(gclk));
	jdff dff_B_h6yxs8or0_2(.din(w_dff_B_Ydaoss7M1_2),.dout(w_dff_B_h6yxs8or0_2),.clk(gclk));
	jdff dff_B_KjWYSJ7N2_2(.din(w_dff_B_h6yxs8or0_2),.dout(w_dff_B_KjWYSJ7N2_2),.clk(gclk));
	jdff dff_B_HqwWS43L9_2(.din(w_dff_B_KjWYSJ7N2_2),.dout(w_dff_B_HqwWS43L9_2),.clk(gclk));
	jdff dff_B_YyNfbTiP0_2(.din(w_dff_B_HqwWS43L9_2),.dout(w_dff_B_YyNfbTiP0_2),.clk(gclk));
	jdff dff_B_N9BA0jPQ2_2(.din(w_dff_B_YyNfbTiP0_2),.dout(w_dff_B_N9BA0jPQ2_2),.clk(gclk));
	jdff dff_B_noWhhSHy3_2(.din(w_dff_B_N9BA0jPQ2_2),.dout(w_dff_B_noWhhSHy3_2),.clk(gclk));
	jdff dff_B_BCpTLhAm0_2(.din(w_dff_B_noWhhSHy3_2),.dout(w_dff_B_BCpTLhAm0_2),.clk(gclk));
	jdff dff_B_zRJPFy7l0_2(.din(w_dff_B_BCpTLhAm0_2),.dout(w_dff_B_zRJPFy7l0_2),.clk(gclk));
	jdff dff_B_1DRiESHt5_2(.din(w_dff_B_zRJPFy7l0_2),.dout(w_dff_B_1DRiESHt5_2),.clk(gclk));
	jdff dff_B_PgG3sjmQ2_2(.din(w_dff_B_1DRiESHt5_2),.dout(w_dff_B_PgG3sjmQ2_2),.clk(gclk));
	jdff dff_B_gZWKAKOx8_2(.din(w_dff_B_PgG3sjmQ2_2),.dout(w_dff_B_gZWKAKOx8_2),.clk(gclk));
	jdff dff_B_Lh3Q3shL4_2(.din(w_dff_B_gZWKAKOx8_2),.dout(w_dff_B_Lh3Q3shL4_2),.clk(gclk));
	jdff dff_B_lUCdtiE86_2(.din(w_dff_B_Lh3Q3shL4_2),.dout(w_dff_B_lUCdtiE86_2),.clk(gclk));
	jdff dff_B_Nozv5TuX6_2(.din(w_dff_B_lUCdtiE86_2),.dout(w_dff_B_Nozv5TuX6_2),.clk(gclk));
	jdff dff_B_AmTbGDv35_2(.din(w_dff_B_Nozv5TuX6_2),.dout(w_dff_B_AmTbGDv35_2),.clk(gclk));
	jdff dff_B_ow1ACzzW2_2(.din(w_dff_B_AmTbGDv35_2),.dout(w_dff_B_ow1ACzzW2_2),.clk(gclk));
	jdff dff_B_HFGdEqMT4_2(.din(n1807),.dout(w_dff_B_HFGdEqMT4_2),.clk(gclk));
	jdff dff_B_FNKI545q1_2(.din(w_dff_B_HFGdEqMT4_2),.dout(w_dff_B_FNKI545q1_2),.clk(gclk));
	jdff dff_B_KrnCxEr38_2(.din(w_dff_B_FNKI545q1_2),.dout(w_dff_B_KrnCxEr38_2),.clk(gclk));
	jdff dff_B_DauTOFYo8_2(.din(w_dff_B_KrnCxEr38_2),.dout(w_dff_B_DauTOFYo8_2),.clk(gclk));
	jdff dff_B_IV5fNUIQ2_2(.din(w_dff_B_DauTOFYo8_2),.dout(w_dff_B_IV5fNUIQ2_2),.clk(gclk));
	jdff dff_B_ho4FAEGm2_2(.din(w_dff_B_IV5fNUIQ2_2),.dout(w_dff_B_ho4FAEGm2_2),.clk(gclk));
	jdff dff_B_cY8mQqxw9_2(.din(w_dff_B_ho4FAEGm2_2),.dout(w_dff_B_cY8mQqxw9_2),.clk(gclk));
	jdff dff_B_D1La8O7d4_2(.din(w_dff_B_cY8mQqxw9_2),.dout(w_dff_B_D1La8O7d4_2),.clk(gclk));
	jdff dff_B_mSswtA1x9_2(.din(w_dff_B_D1La8O7d4_2),.dout(w_dff_B_mSswtA1x9_2),.clk(gclk));
	jdff dff_B_owMSigKX4_2(.din(w_dff_B_mSswtA1x9_2),.dout(w_dff_B_owMSigKX4_2),.clk(gclk));
	jdff dff_B_4QbQ19Db6_2(.din(w_dff_B_owMSigKX4_2),.dout(w_dff_B_4QbQ19Db6_2),.clk(gclk));
	jdff dff_B_8XDFSGgI4_2(.din(w_dff_B_4QbQ19Db6_2),.dout(w_dff_B_8XDFSGgI4_2),.clk(gclk));
	jdff dff_B_ViWPzmuD8_2(.din(w_dff_B_8XDFSGgI4_2),.dout(w_dff_B_ViWPzmuD8_2),.clk(gclk));
	jdff dff_B_5y5s0Fwa5_2(.din(w_dff_B_ViWPzmuD8_2),.dout(w_dff_B_5y5s0Fwa5_2),.clk(gclk));
	jdff dff_B_AROnbn3k2_2(.din(w_dff_B_5y5s0Fwa5_2),.dout(w_dff_B_AROnbn3k2_2),.clk(gclk));
	jdff dff_B_Mg6T2Yox1_2(.din(w_dff_B_AROnbn3k2_2),.dout(w_dff_B_Mg6T2Yox1_2),.clk(gclk));
	jdff dff_B_AFIxo8Gk2_2(.din(w_dff_B_Mg6T2Yox1_2),.dout(w_dff_B_AFIxo8Gk2_2),.clk(gclk));
	jdff dff_B_rylRi0Fa8_2(.din(w_dff_B_AFIxo8Gk2_2),.dout(w_dff_B_rylRi0Fa8_2),.clk(gclk));
	jdff dff_B_wbsNyRlg3_2(.din(w_dff_B_rylRi0Fa8_2),.dout(w_dff_B_wbsNyRlg3_2),.clk(gclk));
	jdff dff_B_VIYIXzl65_2(.din(w_dff_B_wbsNyRlg3_2),.dout(w_dff_B_VIYIXzl65_2),.clk(gclk));
	jdff dff_B_H0yJlRON3_2(.din(w_dff_B_VIYIXzl65_2),.dout(w_dff_B_H0yJlRON3_2),.clk(gclk));
	jdff dff_B_JmeE15He0_2(.din(w_dff_B_H0yJlRON3_2),.dout(w_dff_B_JmeE15He0_2),.clk(gclk));
	jdff dff_B_N4uAV5mt4_2(.din(w_dff_B_JmeE15He0_2),.dout(w_dff_B_N4uAV5mt4_2),.clk(gclk));
	jdff dff_B_hFx8PE626_2(.din(w_dff_B_N4uAV5mt4_2),.dout(w_dff_B_hFx8PE626_2),.clk(gclk));
	jdff dff_B_R9P3XLvI8_2(.din(w_dff_B_hFx8PE626_2),.dout(w_dff_B_R9P3XLvI8_2),.clk(gclk));
	jdff dff_B_GcIMSQIs1_2(.din(w_dff_B_R9P3XLvI8_2),.dout(w_dff_B_GcIMSQIs1_2),.clk(gclk));
	jdff dff_B_RSrqNa6d8_2(.din(w_dff_B_GcIMSQIs1_2),.dout(w_dff_B_RSrqNa6d8_2),.clk(gclk));
	jdff dff_B_I3e2HnSc6_2(.din(w_dff_B_RSrqNa6d8_2),.dout(w_dff_B_I3e2HnSc6_2),.clk(gclk));
	jdff dff_B_6v8dgnx22_2(.din(w_dff_B_I3e2HnSc6_2),.dout(w_dff_B_6v8dgnx22_2),.clk(gclk));
	jdff dff_B_VhYtEGdF0_2(.din(w_dff_B_6v8dgnx22_2),.dout(w_dff_B_VhYtEGdF0_2),.clk(gclk));
	jdff dff_B_Zk5GAJos8_2(.din(w_dff_B_VhYtEGdF0_2),.dout(w_dff_B_Zk5GAJos8_2),.clk(gclk));
	jdff dff_B_TQuqQPn63_2(.din(w_dff_B_Zk5GAJos8_2),.dout(w_dff_B_TQuqQPn63_2),.clk(gclk));
	jdff dff_B_GItCAx1e5_2(.din(w_dff_B_TQuqQPn63_2),.dout(w_dff_B_GItCAx1e5_2),.clk(gclk));
	jdff dff_B_Q7WRgSCv3_2(.din(w_dff_B_GItCAx1e5_2),.dout(w_dff_B_Q7WRgSCv3_2),.clk(gclk));
	jdff dff_B_mqDfCepF3_2(.din(w_dff_B_Q7WRgSCv3_2),.dout(w_dff_B_mqDfCepF3_2),.clk(gclk));
	jdff dff_B_w5f0Zlpc7_2(.din(w_dff_B_mqDfCepF3_2),.dout(w_dff_B_w5f0Zlpc7_2),.clk(gclk));
	jdff dff_B_M4Scfoab0_2(.din(w_dff_B_w5f0Zlpc7_2),.dout(w_dff_B_M4Scfoab0_2),.clk(gclk));
	jdff dff_B_YzKK4ROU9_2(.din(w_dff_B_M4Scfoab0_2),.dout(w_dff_B_YzKK4ROU9_2),.clk(gclk));
	jdff dff_B_8p4IIfyw3_2(.din(w_dff_B_YzKK4ROU9_2),.dout(w_dff_B_8p4IIfyw3_2),.clk(gclk));
	jdff dff_B_JVjmycqe6_2(.din(w_dff_B_8p4IIfyw3_2),.dout(w_dff_B_JVjmycqe6_2),.clk(gclk));
	jdff dff_B_h8pzWNGf7_2(.din(w_dff_B_JVjmycqe6_2),.dout(w_dff_B_h8pzWNGf7_2),.clk(gclk));
	jdff dff_B_Xdq2iI6f7_2(.din(w_dff_B_h8pzWNGf7_2),.dout(w_dff_B_Xdq2iI6f7_2),.clk(gclk));
	jdff dff_B_M0uDOyqm7_2(.din(w_dff_B_Xdq2iI6f7_2),.dout(w_dff_B_M0uDOyqm7_2),.clk(gclk));
	jdff dff_B_wYU0PGcR7_2(.din(w_dff_B_M0uDOyqm7_2),.dout(w_dff_B_wYU0PGcR7_2),.clk(gclk));
	jdff dff_B_wn0HOENM2_2(.din(w_dff_B_wYU0PGcR7_2),.dout(w_dff_B_wn0HOENM2_2),.clk(gclk));
	jdff dff_B_pG2N7egd5_2(.din(w_dff_B_wn0HOENM2_2),.dout(w_dff_B_pG2N7egd5_2),.clk(gclk));
	jdff dff_B_UsXC6kDV5_2(.din(w_dff_B_pG2N7egd5_2),.dout(w_dff_B_UsXC6kDV5_2),.clk(gclk));
	jdff dff_B_8DaWnkuS7_2(.din(w_dff_B_UsXC6kDV5_2),.dout(w_dff_B_8DaWnkuS7_2),.clk(gclk));
	jdff dff_B_yBGWBQQ73_2(.din(w_dff_B_8DaWnkuS7_2),.dout(w_dff_B_yBGWBQQ73_2),.clk(gclk));
	jdff dff_B_HMAyniji3_2(.din(w_dff_B_yBGWBQQ73_2),.dout(w_dff_B_HMAyniji3_2),.clk(gclk));
	jdff dff_B_qj2Sy5ei5_2(.din(w_dff_B_HMAyniji3_2),.dout(w_dff_B_qj2Sy5ei5_2),.clk(gclk));
	jdff dff_B_kHRFU87x7_2(.din(w_dff_B_qj2Sy5ei5_2),.dout(w_dff_B_kHRFU87x7_2),.clk(gclk));
	jdff dff_B_TSuX6jo15_2(.din(w_dff_B_kHRFU87x7_2),.dout(w_dff_B_TSuX6jo15_2),.clk(gclk));
	jdff dff_B_NjmfjCyy8_2(.din(w_dff_B_TSuX6jo15_2),.dout(w_dff_B_NjmfjCyy8_2),.clk(gclk));
	jdff dff_B_hqG9jUJl5_2(.din(n1806),.dout(w_dff_B_hqG9jUJl5_2),.clk(gclk));
	jdff dff_B_HZcRA8yf1_1(.din(n1804),.dout(w_dff_B_HZcRA8yf1_1),.clk(gclk));
	jdff dff_B_DBvI3FUx2_2(.din(n1775),.dout(w_dff_B_DBvI3FUx2_2),.clk(gclk));
	jdff dff_B_0bcAbLjy1_2(.din(w_dff_B_DBvI3FUx2_2),.dout(w_dff_B_0bcAbLjy1_2),.clk(gclk));
	jdff dff_B_pLM2oyV69_2(.din(w_dff_B_0bcAbLjy1_2),.dout(w_dff_B_pLM2oyV69_2),.clk(gclk));
	jdff dff_B_QyA5ih9P2_2(.din(w_dff_B_pLM2oyV69_2),.dout(w_dff_B_QyA5ih9P2_2),.clk(gclk));
	jdff dff_B_tlYb8Ct29_2(.din(w_dff_B_QyA5ih9P2_2),.dout(w_dff_B_tlYb8Ct29_2),.clk(gclk));
	jdff dff_B_GUWN96WQ5_2(.din(w_dff_B_tlYb8Ct29_2),.dout(w_dff_B_GUWN96WQ5_2),.clk(gclk));
	jdff dff_B_XE9YeepA2_2(.din(w_dff_B_GUWN96WQ5_2),.dout(w_dff_B_XE9YeepA2_2),.clk(gclk));
	jdff dff_B_QeLZ2IJi2_2(.din(w_dff_B_XE9YeepA2_2),.dout(w_dff_B_QeLZ2IJi2_2),.clk(gclk));
	jdff dff_B_FBoJmY6D3_2(.din(w_dff_B_QeLZ2IJi2_2),.dout(w_dff_B_FBoJmY6D3_2),.clk(gclk));
	jdff dff_B_cNUbaqCd4_2(.din(w_dff_B_FBoJmY6D3_2),.dout(w_dff_B_cNUbaqCd4_2),.clk(gclk));
	jdff dff_B_BzgW8faj8_2(.din(w_dff_B_cNUbaqCd4_2),.dout(w_dff_B_BzgW8faj8_2),.clk(gclk));
	jdff dff_B_cGdMyVA66_2(.din(w_dff_B_BzgW8faj8_2),.dout(w_dff_B_cGdMyVA66_2),.clk(gclk));
	jdff dff_B_A7Xjo4ef8_2(.din(w_dff_B_cGdMyVA66_2),.dout(w_dff_B_A7Xjo4ef8_2),.clk(gclk));
	jdff dff_B_0tvM4rOw1_2(.din(w_dff_B_A7Xjo4ef8_2),.dout(w_dff_B_0tvM4rOw1_2),.clk(gclk));
	jdff dff_B_0MFJM3tm7_2(.din(w_dff_B_0tvM4rOw1_2),.dout(w_dff_B_0MFJM3tm7_2),.clk(gclk));
	jdff dff_B_9QnjixyN7_2(.din(w_dff_B_0MFJM3tm7_2),.dout(w_dff_B_9QnjixyN7_2),.clk(gclk));
	jdff dff_B_u6xCdFJu4_2(.din(w_dff_B_9QnjixyN7_2),.dout(w_dff_B_u6xCdFJu4_2),.clk(gclk));
	jdff dff_B_zmE3oj9M0_2(.din(w_dff_B_u6xCdFJu4_2),.dout(w_dff_B_zmE3oj9M0_2),.clk(gclk));
	jdff dff_B_WtUrwfds3_2(.din(w_dff_B_zmE3oj9M0_2),.dout(w_dff_B_WtUrwfds3_2),.clk(gclk));
	jdff dff_B_4wu9n1Mw6_2(.din(w_dff_B_WtUrwfds3_2),.dout(w_dff_B_4wu9n1Mw6_2),.clk(gclk));
	jdff dff_B_nDrme8X40_2(.din(w_dff_B_4wu9n1Mw6_2),.dout(w_dff_B_nDrme8X40_2),.clk(gclk));
	jdff dff_B_6YbSQnxc5_2(.din(w_dff_B_nDrme8X40_2),.dout(w_dff_B_6YbSQnxc5_2),.clk(gclk));
	jdff dff_B_j9s88Kr50_2(.din(w_dff_B_6YbSQnxc5_2),.dout(w_dff_B_j9s88Kr50_2),.clk(gclk));
	jdff dff_B_n5MbotQ47_2(.din(w_dff_B_j9s88Kr50_2),.dout(w_dff_B_n5MbotQ47_2),.clk(gclk));
	jdff dff_B_QdihqDre8_2(.din(w_dff_B_n5MbotQ47_2),.dout(w_dff_B_QdihqDre8_2),.clk(gclk));
	jdff dff_B_VrAU1dhq1_2(.din(w_dff_B_QdihqDre8_2),.dout(w_dff_B_VrAU1dhq1_2),.clk(gclk));
	jdff dff_B_fixnhraI4_2(.din(w_dff_B_VrAU1dhq1_2),.dout(w_dff_B_fixnhraI4_2),.clk(gclk));
	jdff dff_B_XJFtRB5M8_2(.din(w_dff_B_fixnhraI4_2),.dout(w_dff_B_XJFtRB5M8_2),.clk(gclk));
	jdff dff_B_qOCNdoRj7_2(.din(w_dff_B_XJFtRB5M8_2),.dout(w_dff_B_qOCNdoRj7_2),.clk(gclk));
	jdff dff_B_AnMfmTVn5_2(.din(w_dff_B_qOCNdoRj7_2),.dout(w_dff_B_AnMfmTVn5_2),.clk(gclk));
	jdff dff_B_cznM22t16_2(.din(w_dff_B_AnMfmTVn5_2),.dout(w_dff_B_cznM22t16_2),.clk(gclk));
	jdff dff_B_bynwQf8f8_2(.din(w_dff_B_cznM22t16_2),.dout(w_dff_B_bynwQf8f8_2),.clk(gclk));
	jdff dff_B_PoecEloe9_2(.din(w_dff_B_bynwQf8f8_2),.dout(w_dff_B_PoecEloe9_2),.clk(gclk));
	jdff dff_B_YEvfCuoy8_2(.din(w_dff_B_PoecEloe9_2),.dout(w_dff_B_YEvfCuoy8_2),.clk(gclk));
	jdff dff_B_rnrDXxx41_2(.din(w_dff_B_YEvfCuoy8_2),.dout(w_dff_B_rnrDXxx41_2),.clk(gclk));
	jdff dff_B_OECkqqyE4_2(.din(w_dff_B_rnrDXxx41_2),.dout(w_dff_B_OECkqqyE4_2),.clk(gclk));
	jdff dff_B_1b1BGJsA9_2(.din(w_dff_B_OECkqqyE4_2),.dout(w_dff_B_1b1BGJsA9_2),.clk(gclk));
	jdff dff_B_TvnV2T2i9_2(.din(w_dff_B_1b1BGJsA9_2),.dout(w_dff_B_TvnV2T2i9_2),.clk(gclk));
	jdff dff_B_wiJHOoZ48_2(.din(w_dff_B_TvnV2T2i9_2),.dout(w_dff_B_wiJHOoZ48_2),.clk(gclk));
	jdff dff_B_SzOkO6av7_2(.din(w_dff_B_wiJHOoZ48_2),.dout(w_dff_B_SzOkO6av7_2),.clk(gclk));
	jdff dff_B_Uxw2Ipnu7_2(.din(w_dff_B_SzOkO6av7_2),.dout(w_dff_B_Uxw2Ipnu7_2),.clk(gclk));
	jdff dff_B_blLPoyJI9_2(.din(w_dff_B_Uxw2Ipnu7_2),.dout(w_dff_B_blLPoyJI9_2),.clk(gclk));
	jdff dff_B_yE1wnOeW0_2(.din(w_dff_B_blLPoyJI9_2),.dout(w_dff_B_yE1wnOeW0_2),.clk(gclk));
	jdff dff_B_FtgpU8QG4_2(.din(w_dff_B_yE1wnOeW0_2),.dout(w_dff_B_FtgpU8QG4_2),.clk(gclk));
	jdff dff_B_OoBrKVxl6_2(.din(w_dff_B_FtgpU8QG4_2),.dout(w_dff_B_OoBrKVxl6_2),.clk(gclk));
	jdff dff_B_b5X33vDF0_2(.din(w_dff_B_OoBrKVxl6_2),.dout(w_dff_B_b5X33vDF0_2),.clk(gclk));
	jdff dff_B_mS5tJWfv6_2(.din(w_dff_B_b5X33vDF0_2),.dout(w_dff_B_mS5tJWfv6_2),.clk(gclk));
	jdff dff_B_lk55Bam87_2(.din(w_dff_B_mS5tJWfv6_2),.dout(w_dff_B_lk55Bam87_2),.clk(gclk));
	jdff dff_B_KS0wfYEv8_2(.din(w_dff_B_lk55Bam87_2),.dout(w_dff_B_KS0wfYEv8_2),.clk(gclk));
	jdff dff_B_Dvayqm2X9_2(.din(w_dff_B_KS0wfYEv8_2),.dout(w_dff_B_Dvayqm2X9_2),.clk(gclk));
	jdff dff_B_fpdTFUYa8_2(.din(w_dff_B_Dvayqm2X9_2),.dout(w_dff_B_fpdTFUYa8_2),.clk(gclk));
	jdff dff_B_IRqDxaMe2_1(.din(n1781),.dout(w_dff_B_IRqDxaMe2_1),.clk(gclk));
	jdff dff_B_hxknXZrK4_1(.din(w_dff_B_IRqDxaMe2_1),.dout(w_dff_B_hxknXZrK4_1),.clk(gclk));
	jdff dff_B_5KS1wJEA4_2(.din(n1780),.dout(w_dff_B_5KS1wJEA4_2),.clk(gclk));
	jdff dff_B_kywnD8D52_2(.din(w_dff_B_5KS1wJEA4_2),.dout(w_dff_B_kywnD8D52_2),.clk(gclk));
	jdff dff_B_JA8KGkvM4_2(.din(w_dff_B_kywnD8D52_2),.dout(w_dff_B_JA8KGkvM4_2),.clk(gclk));
	jdff dff_B_HbnxkMWh2_2(.din(w_dff_B_JA8KGkvM4_2),.dout(w_dff_B_HbnxkMWh2_2),.clk(gclk));
	jdff dff_B_P0esF45n4_2(.din(w_dff_B_HbnxkMWh2_2),.dout(w_dff_B_P0esF45n4_2),.clk(gclk));
	jdff dff_B_XCEmDejO7_2(.din(w_dff_B_P0esF45n4_2),.dout(w_dff_B_XCEmDejO7_2),.clk(gclk));
	jdff dff_B_YEiDr6lP2_2(.din(w_dff_B_XCEmDejO7_2),.dout(w_dff_B_YEiDr6lP2_2),.clk(gclk));
	jdff dff_B_1AgA72WP7_2(.din(w_dff_B_YEiDr6lP2_2),.dout(w_dff_B_1AgA72WP7_2),.clk(gclk));
	jdff dff_B_BgpCTGJ53_2(.din(w_dff_B_1AgA72WP7_2),.dout(w_dff_B_BgpCTGJ53_2),.clk(gclk));
	jdff dff_B_WfNCh4uI6_2(.din(w_dff_B_BgpCTGJ53_2),.dout(w_dff_B_WfNCh4uI6_2),.clk(gclk));
	jdff dff_B_gH4EAu6N1_2(.din(w_dff_B_WfNCh4uI6_2),.dout(w_dff_B_gH4EAu6N1_2),.clk(gclk));
	jdff dff_B_YvK5si3a3_2(.din(w_dff_B_gH4EAu6N1_2),.dout(w_dff_B_YvK5si3a3_2),.clk(gclk));
	jdff dff_B_pGSOdx9c0_2(.din(w_dff_B_YvK5si3a3_2),.dout(w_dff_B_pGSOdx9c0_2),.clk(gclk));
	jdff dff_B_YVHKVAro5_2(.din(w_dff_B_pGSOdx9c0_2),.dout(w_dff_B_YVHKVAro5_2),.clk(gclk));
	jdff dff_B_ybRAsPRh1_2(.din(w_dff_B_YVHKVAro5_2),.dout(w_dff_B_ybRAsPRh1_2),.clk(gclk));
	jdff dff_B_dpliggGD8_2(.din(w_dff_B_ybRAsPRh1_2),.dout(w_dff_B_dpliggGD8_2),.clk(gclk));
	jdff dff_B_SYalu5ew7_2(.din(w_dff_B_dpliggGD8_2),.dout(w_dff_B_SYalu5ew7_2),.clk(gclk));
	jdff dff_B_JPK31wup3_2(.din(w_dff_B_SYalu5ew7_2),.dout(w_dff_B_JPK31wup3_2),.clk(gclk));
	jdff dff_B_2pjFRDFr0_2(.din(w_dff_B_JPK31wup3_2),.dout(w_dff_B_2pjFRDFr0_2),.clk(gclk));
	jdff dff_B_b2UZ6BZj7_2(.din(w_dff_B_2pjFRDFr0_2),.dout(w_dff_B_b2UZ6BZj7_2),.clk(gclk));
	jdff dff_B_W8ek7kr86_2(.din(w_dff_B_b2UZ6BZj7_2),.dout(w_dff_B_W8ek7kr86_2),.clk(gclk));
	jdff dff_B_aUo1xKZw6_2(.din(w_dff_B_W8ek7kr86_2),.dout(w_dff_B_aUo1xKZw6_2),.clk(gclk));
	jdff dff_B_ZqZfp8yf8_2(.din(w_dff_B_aUo1xKZw6_2),.dout(w_dff_B_ZqZfp8yf8_2),.clk(gclk));
	jdff dff_B_ZfTsfHxK5_2(.din(w_dff_B_ZqZfp8yf8_2),.dout(w_dff_B_ZfTsfHxK5_2),.clk(gclk));
	jdff dff_B_Jxaxbwb33_2(.din(w_dff_B_ZfTsfHxK5_2),.dout(w_dff_B_Jxaxbwb33_2),.clk(gclk));
	jdff dff_B_pyyKvmwy2_2(.din(w_dff_B_Jxaxbwb33_2),.dout(w_dff_B_pyyKvmwy2_2),.clk(gclk));
	jdff dff_B_L7Fcjvbs8_2(.din(w_dff_B_pyyKvmwy2_2),.dout(w_dff_B_L7Fcjvbs8_2),.clk(gclk));
	jdff dff_B_PnLBA0UL6_2(.din(w_dff_B_L7Fcjvbs8_2),.dout(w_dff_B_PnLBA0UL6_2),.clk(gclk));
	jdff dff_B_pYvE194M6_2(.din(w_dff_B_PnLBA0UL6_2),.dout(w_dff_B_pYvE194M6_2),.clk(gclk));
	jdff dff_B_Ei8ldF8G1_2(.din(w_dff_B_pYvE194M6_2),.dout(w_dff_B_Ei8ldF8G1_2),.clk(gclk));
	jdff dff_B_1PeOV0S97_2(.din(w_dff_B_Ei8ldF8G1_2),.dout(w_dff_B_1PeOV0S97_2),.clk(gclk));
	jdff dff_B_1dCMWeoB6_2(.din(w_dff_B_1PeOV0S97_2),.dout(w_dff_B_1dCMWeoB6_2),.clk(gclk));
	jdff dff_B_7PZTt0Nl6_2(.din(w_dff_B_1dCMWeoB6_2),.dout(w_dff_B_7PZTt0Nl6_2),.clk(gclk));
	jdff dff_B_Nixu45cg7_2(.din(w_dff_B_7PZTt0Nl6_2),.dout(w_dff_B_Nixu45cg7_2),.clk(gclk));
	jdff dff_B_o9BeNMxs4_2(.din(w_dff_B_Nixu45cg7_2),.dout(w_dff_B_o9BeNMxs4_2),.clk(gclk));
	jdff dff_B_dPjRhudc3_2(.din(w_dff_B_o9BeNMxs4_2),.dout(w_dff_B_dPjRhudc3_2),.clk(gclk));
	jdff dff_B_I18DbIgU8_2(.din(w_dff_B_dPjRhudc3_2),.dout(w_dff_B_I18DbIgU8_2),.clk(gclk));
	jdff dff_B_fl6qs6778_2(.din(w_dff_B_I18DbIgU8_2),.dout(w_dff_B_fl6qs6778_2),.clk(gclk));
	jdff dff_B_ryPWfqGa6_2(.din(w_dff_B_fl6qs6778_2),.dout(w_dff_B_ryPWfqGa6_2),.clk(gclk));
	jdff dff_B_9pQwhCmg7_2(.din(w_dff_B_ryPWfqGa6_2),.dout(w_dff_B_9pQwhCmg7_2),.clk(gclk));
	jdff dff_B_WMqxo3Es3_2(.din(w_dff_B_9pQwhCmg7_2),.dout(w_dff_B_WMqxo3Es3_2),.clk(gclk));
	jdff dff_B_kYVTeL8l2_2(.din(w_dff_B_WMqxo3Es3_2),.dout(w_dff_B_kYVTeL8l2_2),.clk(gclk));
	jdff dff_B_ok5uJN1p7_2(.din(w_dff_B_kYVTeL8l2_2),.dout(w_dff_B_ok5uJN1p7_2),.clk(gclk));
	jdff dff_B_siBtAxSY7_2(.din(w_dff_B_ok5uJN1p7_2),.dout(w_dff_B_siBtAxSY7_2),.clk(gclk));
	jdff dff_B_qWczEMzF2_2(.din(w_dff_B_siBtAxSY7_2),.dout(w_dff_B_qWczEMzF2_2),.clk(gclk));
	jdff dff_B_TIO3sbTp7_2(.din(w_dff_B_qWczEMzF2_2),.dout(w_dff_B_TIO3sbTp7_2),.clk(gclk));
	jdff dff_B_swwn3wE48_2(.din(w_dff_B_TIO3sbTp7_2),.dout(w_dff_B_swwn3wE48_2),.clk(gclk));
	jdff dff_B_BsNym0BD6_2(.din(w_dff_B_swwn3wE48_2),.dout(w_dff_B_BsNym0BD6_2),.clk(gclk));
	jdff dff_B_ealXpbdV2_2(.din(n1779),.dout(w_dff_B_ealXpbdV2_2),.clk(gclk));
	jdff dff_B_8iza5Kt46_2(.din(w_dff_B_ealXpbdV2_2),.dout(w_dff_B_8iza5Kt46_2),.clk(gclk));
	jdff dff_B_GXbmv8rY9_2(.din(w_dff_B_8iza5Kt46_2),.dout(w_dff_B_GXbmv8rY9_2),.clk(gclk));
	jdff dff_B_XOeGf7qs7_2(.din(w_dff_B_GXbmv8rY9_2),.dout(w_dff_B_XOeGf7qs7_2),.clk(gclk));
	jdff dff_B_v6Cgo9NB8_2(.din(w_dff_B_XOeGf7qs7_2),.dout(w_dff_B_v6Cgo9NB8_2),.clk(gclk));
	jdff dff_B_wSEXmgPU0_2(.din(w_dff_B_v6Cgo9NB8_2),.dout(w_dff_B_wSEXmgPU0_2),.clk(gclk));
	jdff dff_B_hBHke2de9_2(.din(w_dff_B_wSEXmgPU0_2),.dout(w_dff_B_hBHke2de9_2),.clk(gclk));
	jdff dff_B_UNMbelaW4_2(.din(w_dff_B_hBHke2de9_2),.dout(w_dff_B_UNMbelaW4_2),.clk(gclk));
	jdff dff_B_kobvEVYX1_2(.din(w_dff_B_UNMbelaW4_2),.dout(w_dff_B_kobvEVYX1_2),.clk(gclk));
	jdff dff_B_UnQM4R7c6_2(.din(w_dff_B_kobvEVYX1_2),.dout(w_dff_B_UnQM4R7c6_2),.clk(gclk));
	jdff dff_B_LCbHCw8t7_2(.din(w_dff_B_UnQM4R7c6_2),.dout(w_dff_B_LCbHCw8t7_2),.clk(gclk));
	jdff dff_B_HzALTBaN4_2(.din(w_dff_B_LCbHCw8t7_2),.dout(w_dff_B_HzALTBaN4_2),.clk(gclk));
	jdff dff_B_tysyyMfp0_2(.din(w_dff_B_HzALTBaN4_2),.dout(w_dff_B_tysyyMfp0_2),.clk(gclk));
	jdff dff_B_m5zu1xe02_2(.din(w_dff_B_tysyyMfp0_2),.dout(w_dff_B_m5zu1xe02_2),.clk(gclk));
	jdff dff_B_qQP2INB56_2(.din(w_dff_B_m5zu1xe02_2),.dout(w_dff_B_qQP2INB56_2),.clk(gclk));
	jdff dff_B_u60CNJ896_2(.din(w_dff_B_qQP2INB56_2),.dout(w_dff_B_u60CNJ896_2),.clk(gclk));
	jdff dff_B_PHrOfp9n6_2(.din(w_dff_B_u60CNJ896_2),.dout(w_dff_B_PHrOfp9n6_2),.clk(gclk));
	jdff dff_B_QJ3luVGO8_2(.din(w_dff_B_PHrOfp9n6_2),.dout(w_dff_B_QJ3luVGO8_2),.clk(gclk));
	jdff dff_B_HAjFXVIc1_2(.din(w_dff_B_QJ3luVGO8_2),.dout(w_dff_B_HAjFXVIc1_2),.clk(gclk));
	jdff dff_B_PMh6y69q2_2(.din(w_dff_B_HAjFXVIc1_2),.dout(w_dff_B_PMh6y69q2_2),.clk(gclk));
	jdff dff_B_xmGpfmcz5_2(.din(w_dff_B_PMh6y69q2_2),.dout(w_dff_B_xmGpfmcz5_2),.clk(gclk));
	jdff dff_B_Lk5xmkvt5_2(.din(w_dff_B_xmGpfmcz5_2),.dout(w_dff_B_Lk5xmkvt5_2),.clk(gclk));
	jdff dff_B_8AoPRLl48_2(.din(w_dff_B_Lk5xmkvt5_2),.dout(w_dff_B_8AoPRLl48_2),.clk(gclk));
	jdff dff_B_VSxlUXr04_2(.din(w_dff_B_8AoPRLl48_2),.dout(w_dff_B_VSxlUXr04_2),.clk(gclk));
	jdff dff_B_yTOMP64G7_2(.din(w_dff_B_VSxlUXr04_2),.dout(w_dff_B_yTOMP64G7_2),.clk(gclk));
	jdff dff_B_Df3n2kFg9_2(.din(w_dff_B_yTOMP64G7_2),.dout(w_dff_B_Df3n2kFg9_2),.clk(gclk));
	jdff dff_B_sg3UA50U7_2(.din(w_dff_B_Df3n2kFg9_2),.dout(w_dff_B_sg3UA50U7_2),.clk(gclk));
	jdff dff_B_oq90p8J44_2(.din(w_dff_B_sg3UA50U7_2),.dout(w_dff_B_oq90p8J44_2),.clk(gclk));
	jdff dff_B_5u973HIt0_2(.din(w_dff_B_oq90p8J44_2),.dout(w_dff_B_5u973HIt0_2),.clk(gclk));
	jdff dff_B_D8vfNS1L9_2(.din(w_dff_B_5u973HIt0_2),.dout(w_dff_B_D8vfNS1L9_2),.clk(gclk));
	jdff dff_B_Lac3mYhn1_2(.din(w_dff_B_D8vfNS1L9_2),.dout(w_dff_B_Lac3mYhn1_2),.clk(gclk));
	jdff dff_B_iJYaALo58_2(.din(w_dff_B_Lac3mYhn1_2),.dout(w_dff_B_iJYaALo58_2),.clk(gclk));
	jdff dff_B_hxm3uO8t9_2(.din(w_dff_B_iJYaALo58_2),.dout(w_dff_B_hxm3uO8t9_2),.clk(gclk));
	jdff dff_B_w41tatFL0_2(.din(w_dff_B_hxm3uO8t9_2),.dout(w_dff_B_w41tatFL0_2),.clk(gclk));
	jdff dff_B_nh76Sbsk4_2(.din(w_dff_B_w41tatFL0_2),.dout(w_dff_B_nh76Sbsk4_2),.clk(gclk));
	jdff dff_B_SldmnIo06_2(.din(w_dff_B_nh76Sbsk4_2),.dout(w_dff_B_SldmnIo06_2),.clk(gclk));
	jdff dff_B_JJZvrVZY7_2(.din(w_dff_B_SldmnIo06_2),.dout(w_dff_B_JJZvrVZY7_2),.clk(gclk));
	jdff dff_B_qSktLfQv8_2(.din(w_dff_B_JJZvrVZY7_2),.dout(w_dff_B_qSktLfQv8_2),.clk(gclk));
	jdff dff_B_xROvHceJ8_2(.din(w_dff_B_qSktLfQv8_2),.dout(w_dff_B_xROvHceJ8_2),.clk(gclk));
	jdff dff_B_dRrEVYHj5_2(.din(w_dff_B_xROvHceJ8_2),.dout(w_dff_B_dRrEVYHj5_2),.clk(gclk));
	jdff dff_B_8F4mGf0c5_2(.din(w_dff_B_dRrEVYHj5_2),.dout(w_dff_B_8F4mGf0c5_2),.clk(gclk));
	jdff dff_B_rAZiex4m4_2(.din(w_dff_B_8F4mGf0c5_2),.dout(w_dff_B_rAZiex4m4_2),.clk(gclk));
	jdff dff_B_LzIUIt3x7_2(.din(w_dff_B_rAZiex4m4_2),.dout(w_dff_B_LzIUIt3x7_2),.clk(gclk));
	jdff dff_B_HfomW0Ed8_2(.din(w_dff_B_LzIUIt3x7_2),.dout(w_dff_B_HfomW0Ed8_2),.clk(gclk));
	jdff dff_B_md8JpPnn8_2(.din(w_dff_B_HfomW0Ed8_2),.dout(w_dff_B_md8JpPnn8_2),.clk(gclk));
	jdff dff_B_SOKTh8qq0_2(.din(w_dff_B_md8JpPnn8_2),.dout(w_dff_B_SOKTh8qq0_2),.clk(gclk));
	jdff dff_B_eZk0nAOL2_2(.din(w_dff_B_SOKTh8qq0_2),.dout(w_dff_B_eZk0nAOL2_2),.clk(gclk));
	jdff dff_B_7r3JzWwv3_2(.din(w_dff_B_eZk0nAOL2_2),.dout(w_dff_B_7r3JzWwv3_2),.clk(gclk));
	jdff dff_B_UyeOzMud5_2(.din(w_dff_B_7r3JzWwv3_2),.dout(w_dff_B_UyeOzMud5_2),.clk(gclk));
	jdff dff_B_ZgDUxRu08_2(.din(w_dff_B_UyeOzMud5_2),.dout(w_dff_B_ZgDUxRu08_2),.clk(gclk));
	jdff dff_B_jQz8xYvG9_2(.din(n1778),.dout(w_dff_B_jQz8xYvG9_2),.clk(gclk));
	jdff dff_B_4H58eYGh5_1(.din(n1776),.dout(w_dff_B_4H58eYGh5_1),.clk(gclk));
	jdff dff_B_iK0CLIKr8_2(.din(n1740),.dout(w_dff_B_iK0CLIKr8_2),.clk(gclk));
	jdff dff_B_gJhXQPSx6_2(.din(w_dff_B_iK0CLIKr8_2),.dout(w_dff_B_gJhXQPSx6_2),.clk(gclk));
	jdff dff_B_clkvx3ng3_2(.din(w_dff_B_gJhXQPSx6_2),.dout(w_dff_B_clkvx3ng3_2),.clk(gclk));
	jdff dff_B_HUTX4Mc65_2(.din(w_dff_B_clkvx3ng3_2),.dout(w_dff_B_HUTX4Mc65_2),.clk(gclk));
	jdff dff_B_ICUFsK3n1_2(.din(w_dff_B_HUTX4Mc65_2),.dout(w_dff_B_ICUFsK3n1_2),.clk(gclk));
	jdff dff_B_A4EuyVaJ1_2(.din(w_dff_B_ICUFsK3n1_2),.dout(w_dff_B_A4EuyVaJ1_2),.clk(gclk));
	jdff dff_B_BT39IYJk7_2(.din(w_dff_B_A4EuyVaJ1_2),.dout(w_dff_B_BT39IYJk7_2),.clk(gclk));
	jdff dff_B_iHUdGvY64_2(.din(w_dff_B_BT39IYJk7_2),.dout(w_dff_B_iHUdGvY64_2),.clk(gclk));
	jdff dff_B_Vkybx9sd6_2(.din(w_dff_B_iHUdGvY64_2),.dout(w_dff_B_Vkybx9sd6_2),.clk(gclk));
	jdff dff_B_2hR0JXpz0_2(.din(w_dff_B_Vkybx9sd6_2),.dout(w_dff_B_2hR0JXpz0_2),.clk(gclk));
	jdff dff_B_BONtfjYJ0_2(.din(w_dff_B_2hR0JXpz0_2),.dout(w_dff_B_BONtfjYJ0_2),.clk(gclk));
	jdff dff_B_S5PEcgqK1_2(.din(w_dff_B_BONtfjYJ0_2),.dout(w_dff_B_S5PEcgqK1_2),.clk(gclk));
	jdff dff_B_EIshArMQ8_2(.din(w_dff_B_S5PEcgqK1_2),.dout(w_dff_B_EIshArMQ8_2),.clk(gclk));
	jdff dff_B_oKJfnPyo3_2(.din(w_dff_B_EIshArMQ8_2),.dout(w_dff_B_oKJfnPyo3_2),.clk(gclk));
	jdff dff_B_7MRlVLlA9_2(.din(w_dff_B_oKJfnPyo3_2),.dout(w_dff_B_7MRlVLlA9_2),.clk(gclk));
	jdff dff_B_IxnnyTHG6_2(.din(w_dff_B_7MRlVLlA9_2),.dout(w_dff_B_IxnnyTHG6_2),.clk(gclk));
	jdff dff_B_qtsZK9MU1_2(.din(w_dff_B_IxnnyTHG6_2),.dout(w_dff_B_qtsZK9MU1_2),.clk(gclk));
	jdff dff_B_aNBclOXF6_2(.din(w_dff_B_qtsZK9MU1_2),.dout(w_dff_B_aNBclOXF6_2),.clk(gclk));
	jdff dff_B_Kak0d9OD3_2(.din(w_dff_B_aNBclOXF6_2),.dout(w_dff_B_Kak0d9OD3_2),.clk(gclk));
	jdff dff_B_KeMCybJm5_2(.din(w_dff_B_Kak0d9OD3_2),.dout(w_dff_B_KeMCybJm5_2),.clk(gclk));
	jdff dff_B_81SBDW203_2(.din(w_dff_B_KeMCybJm5_2),.dout(w_dff_B_81SBDW203_2),.clk(gclk));
	jdff dff_B_1V6OoTMh3_2(.din(w_dff_B_81SBDW203_2),.dout(w_dff_B_1V6OoTMh3_2),.clk(gclk));
	jdff dff_B_RaGXJgGj1_2(.din(w_dff_B_1V6OoTMh3_2),.dout(w_dff_B_RaGXJgGj1_2),.clk(gclk));
	jdff dff_B_o8GRixEZ3_2(.din(w_dff_B_RaGXJgGj1_2),.dout(w_dff_B_o8GRixEZ3_2),.clk(gclk));
	jdff dff_B_pLjPmnNs7_2(.din(w_dff_B_o8GRixEZ3_2),.dout(w_dff_B_pLjPmnNs7_2),.clk(gclk));
	jdff dff_B_5yyJ8P2h7_2(.din(w_dff_B_pLjPmnNs7_2),.dout(w_dff_B_5yyJ8P2h7_2),.clk(gclk));
	jdff dff_B_uyht0P7T4_2(.din(w_dff_B_5yyJ8P2h7_2),.dout(w_dff_B_uyht0P7T4_2),.clk(gclk));
	jdff dff_B_gOzMkHVW5_2(.din(w_dff_B_uyht0P7T4_2),.dout(w_dff_B_gOzMkHVW5_2),.clk(gclk));
	jdff dff_B_oQjzj1si8_2(.din(w_dff_B_gOzMkHVW5_2),.dout(w_dff_B_oQjzj1si8_2),.clk(gclk));
	jdff dff_B_hlNPSmZN2_2(.din(w_dff_B_oQjzj1si8_2),.dout(w_dff_B_hlNPSmZN2_2),.clk(gclk));
	jdff dff_B_hNyIm47R4_2(.din(w_dff_B_hlNPSmZN2_2),.dout(w_dff_B_hNyIm47R4_2),.clk(gclk));
	jdff dff_B_7IPpYafO4_2(.din(w_dff_B_hNyIm47R4_2),.dout(w_dff_B_7IPpYafO4_2),.clk(gclk));
	jdff dff_B_lX9rPIp45_2(.din(w_dff_B_7IPpYafO4_2),.dout(w_dff_B_lX9rPIp45_2),.clk(gclk));
	jdff dff_B_akycZ8pd1_2(.din(w_dff_B_lX9rPIp45_2),.dout(w_dff_B_akycZ8pd1_2),.clk(gclk));
	jdff dff_B_Xrqzdsys4_2(.din(w_dff_B_akycZ8pd1_2),.dout(w_dff_B_Xrqzdsys4_2),.clk(gclk));
	jdff dff_B_plqKYCF24_2(.din(w_dff_B_Xrqzdsys4_2),.dout(w_dff_B_plqKYCF24_2),.clk(gclk));
	jdff dff_B_p29naSmn1_2(.din(w_dff_B_plqKYCF24_2),.dout(w_dff_B_p29naSmn1_2),.clk(gclk));
	jdff dff_B_HP8VGHm88_2(.din(w_dff_B_p29naSmn1_2),.dout(w_dff_B_HP8VGHm88_2),.clk(gclk));
	jdff dff_B_HdqSspbk1_2(.din(w_dff_B_HP8VGHm88_2),.dout(w_dff_B_HdqSspbk1_2),.clk(gclk));
	jdff dff_B_r0mf3nj57_2(.din(w_dff_B_HdqSspbk1_2),.dout(w_dff_B_r0mf3nj57_2),.clk(gclk));
	jdff dff_B_HIEjp3Vf1_2(.din(w_dff_B_r0mf3nj57_2),.dout(w_dff_B_HIEjp3Vf1_2),.clk(gclk));
	jdff dff_B_KZMw3vOh0_2(.din(w_dff_B_HIEjp3Vf1_2),.dout(w_dff_B_KZMw3vOh0_2),.clk(gclk));
	jdff dff_B_dJDkOySD7_2(.din(w_dff_B_KZMw3vOh0_2),.dout(w_dff_B_dJDkOySD7_2),.clk(gclk));
	jdff dff_B_GgSrqpV50_2(.din(w_dff_B_dJDkOySD7_2),.dout(w_dff_B_GgSrqpV50_2),.clk(gclk));
	jdff dff_B_aoa3D9JD2_2(.din(w_dff_B_GgSrqpV50_2),.dout(w_dff_B_aoa3D9JD2_2),.clk(gclk));
	jdff dff_B_wSk8cq3o3_2(.din(w_dff_B_aoa3D9JD2_2),.dout(w_dff_B_wSk8cq3o3_2),.clk(gclk));
	jdff dff_B_DI2GWMrx8_2(.din(w_dff_B_wSk8cq3o3_2),.dout(w_dff_B_DI2GWMrx8_2),.clk(gclk));
	jdff dff_B_Ywyy6tRh3_1(.din(n1746),.dout(w_dff_B_Ywyy6tRh3_1),.clk(gclk));
	jdff dff_B_yr9DqX8w2_1(.din(w_dff_B_Ywyy6tRh3_1),.dout(w_dff_B_yr9DqX8w2_1),.clk(gclk));
	jdff dff_B_ZBHDNJzt6_2(.din(n1745),.dout(w_dff_B_ZBHDNJzt6_2),.clk(gclk));
	jdff dff_B_RmLoZWni9_2(.din(w_dff_B_ZBHDNJzt6_2),.dout(w_dff_B_RmLoZWni9_2),.clk(gclk));
	jdff dff_B_yjM5zYcU9_2(.din(w_dff_B_RmLoZWni9_2),.dout(w_dff_B_yjM5zYcU9_2),.clk(gclk));
	jdff dff_B_n3A0exga1_2(.din(w_dff_B_yjM5zYcU9_2),.dout(w_dff_B_n3A0exga1_2),.clk(gclk));
	jdff dff_B_QtAb0TbW6_2(.din(w_dff_B_n3A0exga1_2),.dout(w_dff_B_QtAb0TbW6_2),.clk(gclk));
	jdff dff_B_0dSs4GBc5_2(.din(w_dff_B_QtAb0TbW6_2),.dout(w_dff_B_0dSs4GBc5_2),.clk(gclk));
	jdff dff_B_hC7cbqva6_2(.din(w_dff_B_0dSs4GBc5_2),.dout(w_dff_B_hC7cbqva6_2),.clk(gclk));
	jdff dff_B_gUP1Vrog7_2(.din(w_dff_B_hC7cbqva6_2),.dout(w_dff_B_gUP1Vrog7_2),.clk(gclk));
	jdff dff_B_xIHU875o3_2(.din(w_dff_B_gUP1Vrog7_2),.dout(w_dff_B_xIHU875o3_2),.clk(gclk));
	jdff dff_B_BZ5gUWDc3_2(.din(w_dff_B_xIHU875o3_2),.dout(w_dff_B_BZ5gUWDc3_2),.clk(gclk));
	jdff dff_B_SduZHkGW3_2(.din(w_dff_B_BZ5gUWDc3_2),.dout(w_dff_B_SduZHkGW3_2),.clk(gclk));
	jdff dff_B_rY42VeaF9_2(.din(w_dff_B_SduZHkGW3_2),.dout(w_dff_B_rY42VeaF9_2),.clk(gclk));
	jdff dff_B_JpIlw6kJ2_2(.din(w_dff_B_rY42VeaF9_2),.dout(w_dff_B_JpIlw6kJ2_2),.clk(gclk));
	jdff dff_B_Req1KuG09_2(.din(w_dff_B_JpIlw6kJ2_2),.dout(w_dff_B_Req1KuG09_2),.clk(gclk));
	jdff dff_B_1u2LQapE3_2(.din(w_dff_B_Req1KuG09_2),.dout(w_dff_B_1u2LQapE3_2),.clk(gclk));
	jdff dff_B_Um9K5SFx7_2(.din(w_dff_B_1u2LQapE3_2),.dout(w_dff_B_Um9K5SFx7_2),.clk(gclk));
	jdff dff_B_00UchqWP0_2(.din(w_dff_B_Um9K5SFx7_2),.dout(w_dff_B_00UchqWP0_2),.clk(gclk));
	jdff dff_B_YxL4j6fr9_2(.din(w_dff_B_00UchqWP0_2),.dout(w_dff_B_YxL4j6fr9_2),.clk(gclk));
	jdff dff_B_jmYPMs3A7_2(.din(w_dff_B_YxL4j6fr9_2),.dout(w_dff_B_jmYPMs3A7_2),.clk(gclk));
	jdff dff_B_KTaYiATc4_2(.din(w_dff_B_jmYPMs3A7_2),.dout(w_dff_B_KTaYiATc4_2),.clk(gclk));
	jdff dff_B_GT5CY0NJ1_2(.din(w_dff_B_KTaYiATc4_2),.dout(w_dff_B_GT5CY0NJ1_2),.clk(gclk));
	jdff dff_B_uPnJlxGY6_2(.din(w_dff_B_GT5CY0NJ1_2),.dout(w_dff_B_uPnJlxGY6_2),.clk(gclk));
	jdff dff_B_4TfFEFmg9_2(.din(w_dff_B_uPnJlxGY6_2),.dout(w_dff_B_4TfFEFmg9_2),.clk(gclk));
	jdff dff_B_bCnXdMgz3_2(.din(w_dff_B_4TfFEFmg9_2),.dout(w_dff_B_bCnXdMgz3_2),.clk(gclk));
	jdff dff_B_HzCfA7cZ8_2(.din(w_dff_B_bCnXdMgz3_2),.dout(w_dff_B_HzCfA7cZ8_2),.clk(gclk));
	jdff dff_B_BFKUpc1U5_2(.din(w_dff_B_HzCfA7cZ8_2),.dout(w_dff_B_BFKUpc1U5_2),.clk(gclk));
	jdff dff_B_0LRMnEKd8_2(.din(w_dff_B_BFKUpc1U5_2),.dout(w_dff_B_0LRMnEKd8_2),.clk(gclk));
	jdff dff_B_uglbfiYX0_2(.din(w_dff_B_0LRMnEKd8_2),.dout(w_dff_B_uglbfiYX0_2),.clk(gclk));
	jdff dff_B_QGDZ9MTw1_2(.din(w_dff_B_uglbfiYX0_2),.dout(w_dff_B_QGDZ9MTw1_2),.clk(gclk));
	jdff dff_B_5Meo4a0n4_2(.din(w_dff_B_QGDZ9MTw1_2),.dout(w_dff_B_5Meo4a0n4_2),.clk(gclk));
	jdff dff_B_SA7uSTSo8_2(.din(w_dff_B_5Meo4a0n4_2),.dout(w_dff_B_SA7uSTSo8_2),.clk(gclk));
	jdff dff_B_azP34OCt8_2(.din(w_dff_B_SA7uSTSo8_2),.dout(w_dff_B_azP34OCt8_2),.clk(gclk));
	jdff dff_B_pX9ORayd2_2(.din(w_dff_B_azP34OCt8_2),.dout(w_dff_B_pX9ORayd2_2),.clk(gclk));
	jdff dff_B_Me2PQC3N9_2(.din(w_dff_B_pX9ORayd2_2),.dout(w_dff_B_Me2PQC3N9_2),.clk(gclk));
	jdff dff_B_OxvjDJ3p1_2(.din(w_dff_B_Me2PQC3N9_2),.dout(w_dff_B_OxvjDJ3p1_2),.clk(gclk));
	jdff dff_B_BwER6cLT9_2(.din(w_dff_B_OxvjDJ3p1_2),.dout(w_dff_B_BwER6cLT9_2),.clk(gclk));
	jdff dff_B_sXh5Bkkm4_2(.din(w_dff_B_BwER6cLT9_2),.dout(w_dff_B_sXh5Bkkm4_2),.clk(gclk));
	jdff dff_B_deZ7pzqU8_2(.din(w_dff_B_sXh5Bkkm4_2),.dout(w_dff_B_deZ7pzqU8_2),.clk(gclk));
	jdff dff_B_TvISKjQx3_2(.din(w_dff_B_deZ7pzqU8_2),.dout(w_dff_B_TvISKjQx3_2),.clk(gclk));
	jdff dff_B_lr0asqRj2_2(.din(w_dff_B_TvISKjQx3_2),.dout(w_dff_B_lr0asqRj2_2),.clk(gclk));
	jdff dff_B_WYGTdMM76_2(.din(w_dff_B_lr0asqRj2_2),.dout(w_dff_B_WYGTdMM76_2),.clk(gclk));
	jdff dff_B_U2e5r6Nl9_2(.din(w_dff_B_WYGTdMM76_2),.dout(w_dff_B_U2e5r6Nl9_2),.clk(gclk));
	jdff dff_B_JvU7r4pt9_2(.din(w_dff_B_U2e5r6Nl9_2),.dout(w_dff_B_JvU7r4pt9_2),.clk(gclk));
	jdff dff_B_DfVGyMBd9_2(.din(w_dff_B_JvU7r4pt9_2),.dout(w_dff_B_DfVGyMBd9_2),.clk(gclk));
	jdff dff_B_dmwKZURY8_2(.din(n1744),.dout(w_dff_B_dmwKZURY8_2),.clk(gclk));
	jdff dff_B_SXHO6v2R8_2(.din(w_dff_B_dmwKZURY8_2),.dout(w_dff_B_SXHO6v2R8_2),.clk(gclk));
	jdff dff_B_AXoFbq769_2(.din(w_dff_B_SXHO6v2R8_2),.dout(w_dff_B_AXoFbq769_2),.clk(gclk));
	jdff dff_B_A6m6aOKY2_2(.din(w_dff_B_AXoFbq769_2),.dout(w_dff_B_A6m6aOKY2_2),.clk(gclk));
	jdff dff_B_bgIJkmEK1_2(.din(w_dff_B_A6m6aOKY2_2),.dout(w_dff_B_bgIJkmEK1_2),.clk(gclk));
	jdff dff_B_KTE7Lz235_2(.din(w_dff_B_bgIJkmEK1_2),.dout(w_dff_B_KTE7Lz235_2),.clk(gclk));
	jdff dff_B_gmtkPaLR3_2(.din(w_dff_B_KTE7Lz235_2),.dout(w_dff_B_gmtkPaLR3_2),.clk(gclk));
	jdff dff_B_LhX2oZAg1_2(.din(w_dff_B_gmtkPaLR3_2),.dout(w_dff_B_LhX2oZAg1_2),.clk(gclk));
	jdff dff_B_rXEFJwjP6_2(.din(w_dff_B_LhX2oZAg1_2),.dout(w_dff_B_rXEFJwjP6_2),.clk(gclk));
	jdff dff_B_GJZ9DoLp6_2(.din(w_dff_B_rXEFJwjP6_2),.dout(w_dff_B_GJZ9DoLp6_2),.clk(gclk));
	jdff dff_B_VebLElUT1_2(.din(w_dff_B_GJZ9DoLp6_2),.dout(w_dff_B_VebLElUT1_2),.clk(gclk));
	jdff dff_B_J01WigQ02_2(.din(w_dff_B_VebLElUT1_2),.dout(w_dff_B_J01WigQ02_2),.clk(gclk));
	jdff dff_B_XJU5Cm8H4_2(.din(w_dff_B_J01WigQ02_2),.dout(w_dff_B_XJU5Cm8H4_2),.clk(gclk));
	jdff dff_B_UcD1Ktzn3_2(.din(w_dff_B_XJU5Cm8H4_2),.dout(w_dff_B_UcD1Ktzn3_2),.clk(gclk));
	jdff dff_B_8PvWckt09_2(.din(w_dff_B_UcD1Ktzn3_2),.dout(w_dff_B_8PvWckt09_2),.clk(gclk));
	jdff dff_B_xnWoSRgK2_2(.din(w_dff_B_8PvWckt09_2),.dout(w_dff_B_xnWoSRgK2_2),.clk(gclk));
	jdff dff_B_v3seb3v67_2(.din(w_dff_B_xnWoSRgK2_2),.dout(w_dff_B_v3seb3v67_2),.clk(gclk));
	jdff dff_B_PFm7VDJ03_2(.din(w_dff_B_v3seb3v67_2),.dout(w_dff_B_PFm7VDJ03_2),.clk(gclk));
	jdff dff_B_H8JqCsWv3_2(.din(w_dff_B_PFm7VDJ03_2),.dout(w_dff_B_H8JqCsWv3_2),.clk(gclk));
	jdff dff_B_s5hRRsaH8_2(.din(w_dff_B_H8JqCsWv3_2),.dout(w_dff_B_s5hRRsaH8_2),.clk(gclk));
	jdff dff_B_XIEIcuha0_2(.din(w_dff_B_s5hRRsaH8_2),.dout(w_dff_B_XIEIcuha0_2),.clk(gclk));
	jdff dff_B_Qx86ozSY4_2(.din(w_dff_B_XIEIcuha0_2),.dout(w_dff_B_Qx86ozSY4_2),.clk(gclk));
	jdff dff_B_YWkvLIPl9_2(.din(w_dff_B_Qx86ozSY4_2),.dout(w_dff_B_YWkvLIPl9_2),.clk(gclk));
	jdff dff_B_Qlte1brX2_2(.din(w_dff_B_YWkvLIPl9_2),.dout(w_dff_B_Qlte1brX2_2),.clk(gclk));
	jdff dff_B_qZScaye56_2(.din(w_dff_B_Qlte1brX2_2),.dout(w_dff_B_qZScaye56_2),.clk(gclk));
	jdff dff_B_PQjzMQKF6_2(.din(w_dff_B_qZScaye56_2),.dout(w_dff_B_PQjzMQKF6_2),.clk(gclk));
	jdff dff_B_IaYODAFQ0_2(.din(w_dff_B_PQjzMQKF6_2),.dout(w_dff_B_IaYODAFQ0_2),.clk(gclk));
	jdff dff_B_EB9xEaQh4_2(.din(w_dff_B_IaYODAFQ0_2),.dout(w_dff_B_EB9xEaQh4_2),.clk(gclk));
	jdff dff_B_ik7VVAML4_2(.din(w_dff_B_EB9xEaQh4_2),.dout(w_dff_B_ik7VVAML4_2),.clk(gclk));
	jdff dff_B_WFEwjM4p7_2(.din(w_dff_B_ik7VVAML4_2),.dout(w_dff_B_WFEwjM4p7_2),.clk(gclk));
	jdff dff_B_BzHw6BKf6_2(.din(w_dff_B_WFEwjM4p7_2),.dout(w_dff_B_BzHw6BKf6_2),.clk(gclk));
	jdff dff_B_c1Yp6nVe7_2(.din(w_dff_B_BzHw6BKf6_2),.dout(w_dff_B_c1Yp6nVe7_2),.clk(gclk));
	jdff dff_B_kENMhCXh5_2(.din(w_dff_B_c1Yp6nVe7_2),.dout(w_dff_B_kENMhCXh5_2),.clk(gclk));
	jdff dff_B_fw8qvMm93_2(.din(w_dff_B_kENMhCXh5_2),.dout(w_dff_B_fw8qvMm93_2),.clk(gclk));
	jdff dff_B_hQUSD2Ng3_2(.din(w_dff_B_fw8qvMm93_2),.dout(w_dff_B_hQUSD2Ng3_2),.clk(gclk));
	jdff dff_B_u5CPnxKk6_2(.din(w_dff_B_hQUSD2Ng3_2),.dout(w_dff_B_u5CPnxKk6_2),.clk(gclk));
	jdff dff_B_hO2WXrgp2_2(.din(w_dff_B_u5CPnxKk6_2),.dout(w_dff_B_hO2WXrgp2_2),.clk(gclk));
	jdff dff_B_0BPhTIYv2_2(.din(w_dff_B_hO2WXrgp2_2),.dout(w_dff_B_0BPhTIYv2_2),.clk(gclk));
	jdff dff_B_qq5oRZqx1_2(.din(w_dff_B_0BPhTIYv2_2),.dout(w_dff_B_qq5oRZqx1_2),.clk(gclk));
	jdff dff_B_n31KSzgu9_2(.din(w_dff_B_qq5oRZqx1_2),.dout(w_dff_B_n31KSzgu9_2),.clk(gclk));
	jdff dff_B_0jfTam7d6_2(.din(w_dff_B_n31KSzgu9_2),.dout(w_dff_B_0jfTam7d6_2),.clk(gclk));
	jdff dff_B_CEhtiWqJ5_2(.din(w_dff_B_0jfTam7d6_2),.dout(w_dff_B_CEhtiWqJ5_2),.clk(gclk));
	jdff dff_B_14UZf4QF2_2(.din(w_dff_B_CEhtiWqJ5_2),.dout(w_dff_B_14UZf4QF2_2),.clk(gclk));
	jdff dff_B_S55qrRp56_2(.din(w_dff_B_14UZf4QF2_2),.dout(w_dff_B_S55qrRp56_2),.clk(gclk));
	jdff dff_B_YlIqJLc14_2(.din(w_dff_B_S55qrRp56_2),.dout(w_dff_B_YlIqJLc14_2),.clk(gclk));
	jdff dff_B_o76WopWf3_2(.din(w_dff_B_YlIqJLc14_2),.dout(w_dff_B_o76WopWf3_2),.clk(gclk));
	jdff dff_B_AdJXDMSH1_2(.din(n1743),.dout(w_dff_B_AdJXDMSH1_2),.clk(gclk));
	jdff dff_B_15EDfjX83_1(.din(n1741),.dout(w_dff_B_15EDfjX83_1),.clk(gclk));
	jdff dff_B_hw018sdB4_2(.din(n1699),.dout(w_dff_B_hw018sdB4_2),.clk(gclk));
	jdff dff_B_w1GA6uHh1_2(.din(w_dff_B_hw018sdB4_2),.dout(w_dff_B_w1GA6uHh1_2),.clk(gclk));
	jdff dff_B_WUq4pdFE3_2(.din(w_dff_B_w1GA6uHh1_2),.dout(w_dff_B_WUq4pdFE3_2),.clk(gclk));
	jdff dff_B_nl0jVKUQ3_2(.din(w_dff_B_WUq4pdFE3_2),.dout(w_dff_B_nl0jVKUQ3_2),.clk(gclk));
	jdff dff_B_5qBng3mg5_2(.din(w_dff_B_nl0jVKUQ3_2),.dout(w_dff_B_5qBng3mg5_2),.clk(gclk));
	jdff dff_B_KdTJFGpu1_2(.din(w_dff_B_5qBng3mg5_2),.dout(w_dff_B_KdTJFGpu1_2),.clk(gclk));
	jdff dff_B_eAEFeRr96_2(.din(w_dff_B_KdTJFGpu1_2),.dout(w_dff_B_eAEFeRr96_2),.clk(gclk));
	jdff dff_B_UQQ4umHl8_2(.din(w_dff_B_eAEFeRr96_2),.dout(w_dff_B_UQQ4umHl8_2),.clk(gclk));
	jdff dff_B_MNn7b7Xs9_2(.din(w_dff_B_UQQ4umHl8_2),.dout(w_dff_B_MNn7b7Xs9_2),.clk(gclk));
	jdff dff_B_LqY1PsdG1_2(.din(w_dff_B_MNn7b7Xs9_2),.dout(w_dff_B_LqY1PsdG1_2),.clk(gclk));
	jdff dff_B_G9ctXz6g4_2(.din(w_dff_B_LqY1PsdG1_2),.dout(w_dff_B_G9ctXz6g4_2),.clk(gclk));
	jdff dff_B_npYuCtBM9_2(.din(w_dff_B_G9ctXz6g4_2),.dout(w_dff_B_npYuCtBM9_2),.clk(gclk));
	jdff dff_B_zvV1A57O7_2(.din(w_dff_B_npYuCtBM9_2),.dout(w_dff_B_zvV1A57O7_2),.clk(gclk));
	jdff dff_B_MRy8ADoc4_2(.din(w_dff_B_zvV1A57O7_2),.dout(w_dff_B_MRy8ADoc4_2),.clk(gclk));
	jdff dff_B_BpPjR14f1_2(.din(w_dff_B_MRy8ADoc4_2),.dout(w_dff_B_BpPjR14f1_2),.clk(gclk));
	jdff dff_B_oUISqR6o9_2(.din(w_dff_B_BpPjR14f1_2),.dout(w_dff_B_oUISqR6o9_2),.clk(gclk));
	jdff dff_B_36X7dkTJ0_2(.din(w_dff_B_oUISqR6o9_2),.dout(w_dff_B_36X7dkTJ0_2),.clk(gclk));
	jdff dff_B_cAQL9vEU0_2(.din(w_dff_B_36X7dkTJ0_2),.dout(w_dff_B_cAQL9vEU0_2),.clk(gclk));
	jdff dff_B_Jong7ev57_2(.din(w_dff_B_cAQL9vEU0_2),.dout(w_dff_B_Jong7ev57_2),.clk(gclk));
	jdff dff_B_EkqaA7YN8_2(.din(w_dff_B_Jong7ev57_2),.dout(w_dff_B_EkqaA7YN8_2),.clk(gclk));
	jdff dff_B_CEDnOjeO9_2(.din(w_dff_B_EkqaA7YN8_2),.dout(w_dff_B_CEDnOjeO9_2),.clk(gclk));
	jdff dff_B_UE83noeL6_2(.din(w_dff_B_CEDnOjeO9_2),.dout(w_dff_B_UE83noeL6_2),.clk(gclk));
	jdff dff_B_ORLXTgM02_2(.din(w_dff_B_UE83noeL6_2),.dout(w_dff_B_ORLXTgM02_2),.clk(gclk));
	jdff dff_B_NPDXFtjq4_2(.din(w_dff_B_ORLXTgM02_2),.dout(w_dff_B_NPDXFtjq4_2),.clk(gclk));
	jdff dff_B_webvFmka7_2(.din(w_dff_B_NPDXFtjq4_2),.dout(w_dff_B_webvFmka7_2),.clk(gclk));
	jdff dff_B_35URPWFz7_2(.din(w_dff_B_webvFmka7_2),.dout(w_dff_B_35URPWFz7_2),.clk(gclk));
	jdff dff_B_JeGnx6XI0_2(.din(w_dff_B_35URPWFz7_2),.dout(w_dff_B_JeGnx6XI0_2),.clk(gclk));
	jdff dff_B_IuYgknc22_2(.din(w_dff_B_JeGnx6XI0_2),.dout(w_dff_B_IuYgknc22_2),.clk(gclk));
	jdff dff_B_5bA0Ij1U2_2(.din(w_dff_B_IuYgknc22_2),.dout(w_dff_B_5bA0Ij1U2_2),.clk(gclk));
	jdff dff_B_AooL0T7V5_2(.din(w_dff_B_5bA0Ij1U2_2),.dout(w_dff_B_AooL0T7V5_2),.clk(gclk));
	jdff dff_B_4pYvItSK8_2(.din(w_dff_B_AooL0T7V5_2),.dout(w_dff_B_4pYvItSK8_2),.clk(gclk));
	jdff dff_B_f2FJ0NOx6_2(.din(w_dff_B_4pYvItSK8_2),.dout(w_dff_B_f2FJ0NOx6_2),.clk(gclk));
	jdff dff_B_uEmygJSJ5_2(.din(w_dff_B_f2FJ0NOx6_2),.dout(w_dff_B_uEmygJSJ5_2),.clk(gclk));
	jdff dff_B_JFA7JtGe1_2(.din(w_dff_B_uEmygJSJ5_2),.dout(w_dff_B_JFA7JtGe1_2),.clk(gclk));
	jdff dff_B_3rzeB9eI1_2(.din(w_dff_B_JFA7JtGe1_2),.dout(w_dff_B_3rzeB9eI1_2),.clk(gclk));
	jdff dff_B_tcYRE7Kr5_2(.din(w_dff_B_3rzeB9eI1_2),.dout(w_dff_B_tcYRE7Kr5_2),.clk(gclk));
	jdff dff_B_JJ2X8Wkx6_2(.din(w_dff_B_tcYRE7Kr5_2),.dout(w_dff_B_JJ2X8Wkx6_2),.clk(gclk));
	jdff dff_B_5O9OFVnQ4_2(.din(w_dff_B_JJ2X8Wkx6_2),.dout(w_dff_B_5O9OFVnQ4_2),.clk(gclk));
	jdff dff_B_250ee1ss1_2(.din(w_dff_B_5O9OFVnQ4_2),.dout(w_dff_B_250ee1ss1_2),.clk(gclk));
	jdff dff_B_eXC6rSt59_2(.din(w_dff_B_250ee1ss1_2),.dout(w_dff_B_eXC6rSt59_2),.clk(gclk));
	jdff dff_B_YYr8HkEN2_2(.din(w_dff_B_eXC6rSt59_2),.dout(w_dff_B_YYr8HkEN2_2),.clk(gclk));
	jdff dff_B_ELxEnowF3_2(.din(w_dff_B_YYr8HkEN2_2),.dout(w_dff_B_ELxEnowF3_2),.clk(gclk));
	jdff dff_B_Jq1IKcFg1_2(.din(w_dff_B_ELxEnowF3_2),.dout(w_dff_B_Jq1IKcFg1_2),.clk(gclk));
	jdff dff_B_fcbH6VQR2_1(.din(n1705),.dout(w_dff_B_fcbH6VQR2_1),.clk(gclk));
	jdff dff_B_bI5IHVx85_1(.din(w_dff_B_fcbH6VQR2_1),.dout(w_dff_B_bI5IHVx85_1),.clk(gclk));
	jdff dff_B_lteTwQdY1_2(.din(n1704),.dout(w_dff_B_lteTwQdY1_2),.clk(gclk));
	jdff dff_B_iLcR157s8_2(.din(w_dff_B_lteTwQdY1_2),.dout(w_dff_B_iLcR157s8_2),.clk(gclk));
	jdff dff_B_eZMmiQCN8_2(.din(w_dff_B_iLcR157s8_2),.dout(w_dff_B_eZMmiQCN8_2),.clk(gclk));
	jdff dff_B_S5naS7Vj3_2(.din(w_dff_B_eZMmiQCN8_2),.dout(w_dff_B_S5naS7Vj3_2),.clk(gclk));
	jdff dff_B_RZeVmmhQ4_2(.din(w_dff_B_S5naS7Vj3_2),.dout(w_dff_B_RZeVmmhQ4_2),.clk(gclk));
	jdff dff_B_fxRrV9pX4_2(.din(w_dff_B_RZeVmmhQ4_2),.dout(w_dff_B_fxRrV9pX4_2),.clk(gclk));
	jdff dff_B_X8NUlGL60_2(.din(w_dff_B_fxRrV9pX4_2),.dout(w_dff_B_X8NUlGL60_2),.clk(gclk));
	jdff dff_B_xgQOqUCw7_2(.din(w_dff_B_X8NUlGL60_2),.dout(w_dff_B_xgQOqUCw7_2),.clk(gclk));
	jdff dff_B_fC2WItM03_2(.din(w_dff_B_xgQOqUCw7_2),.dout(w_dff_B_fC2WItM03_2),.clk(gclk));
	jdff dff_B_EGZFkNvT4_2(.din(w_dff_B_fC2WItM03_2),.dout(w_dff_B_EGZFkNvT4_2),.clk(gclk));
	jdff dff_B_DDLyHUMJ9_2(.din(w_dff_B_EGZFkNvT4_2),.dout(w_dff_B_DDLyHUMJ9_2),.clk(gclk));
	jdff dff_B_wfJQxeM52_2(.din(w_dff_B_DDLyHUMJ9_2),.dout(w_dff_B_wfJQxeM52_2),.clk(gclk));
	jdff dff_B_dTSHe7BF0_2(.din(w_dff_B_wfJQxeM52_2),.dout(w_dff_B_dTSHe7BF0_2),.clk(gclk));
	jdff dff_B_z2yU9exO5_2(.din(w_dff_B_dTSHe7BF0_2),.dout(w_dff_B_z2yU9exO5_2),.clk(gclk));
	jdff dff_B_2sssUxLd8_2(.din(w_dff_B_z2yU9exO5_2),.dout(w_dff_B_2sssUxLd8_2),.clk(gclk));
	jdff dff_B_awshfGlE6_2(.din(w_dff_B_2sssUxLd8_2),.dout(w_dff_B_awshfGlE6_2),.clk(gclk));
	jdff dff_B_LNURQio10_2(.din(w_dff_B_awshfGlE6_2),.dout(w_dff_B_LNURQio10_2),.clk(gclk));
	jdff dff_B_ByZzTT6o7_2(.din(w_dff_B_LNURQio10_2),.dout(w_dff_B_ByZzTT6o7_2),.clk(gclk));
	jdff dff_B_XnHKelct7_2(.din(w_dff_B_ByZzTT6o7_2),.dout(w_dff_B_XnHKelct7_2),.clk(gclk));
	jdff dff_B_A3VL9cYM8_2(.din(w_dff_B_XnHKelct7_2),.dout(w_dff_B_A3VL9cYM8_2),.clk(gclk));
	jdff dff_B_gyfyoaY33_2(.din(w_dff_B_A3VL9cYM8_2),.dout(w_dff_B_gyfyoaY33_2),.clk(gclk));
	jdff dff_B_PX5SqSWe1_2(.din(w_dff_B_gyfyoaY33_2),.dout(w_dff_B_PX5SqSWe1_2),.clk(gclk));
	jdff dff_B_SmpGvvSq4_2(.din(w_dff_B_PX5SqSWe1_2),.dout(w_dff_B_SmpGvvSq4_2),.clk(gclk));
	jdff dff_B_S3tmkxzO9_2(.din(w_dff_B_SmpGvvSq4_2),.dout(w_dff_B_S3tmkxzO9_2),.clk(gclk));
	jdff dff_B_d8v3CkdT2_2(.din(w_dff_B_S3tmkxzO9_2),.dout(w_dff_B_d8v3CkdT2_2),.clk(gclk));
	jdff dff_B_jkyGrMiy0_2(.din(w_dff_B_d8v3CkdT2_2),.dout(w_dff_B_jkyGrMiy0_2),.clk(gclk));
	jdff dff_B_UmyfR7cI8_2(.din(w_dff_B_jkyGrMiy0_2),.dout(w_dff_B_UmyfR7cI8_2),.clk(gclk));
	jdff dff_B_0gsQyXWp5_2(.din(w_dff_B_UmyfR7cI8_2),.dout(w_dff_B_0gsQyXWp5_2),.clk(gclk));
	jdff dff_B_46xgBcQX6_2(.din(w_dff_B_0gsQyXWp5_2),.dout(w_dff_B_46xgBcQX6_2),.clk(gclk));
	jdff dff_B_mj1QzL3k1_2(.din(w_dff_B_46xgBcQX6_2),.dout(w_dff_B_mj1QzL3k1_2),.clk(gclk));
	jdff dff_B_bI7ElMqh7_2(.din(w_dff_B_mj1QzL3k1_2),.dout(w_dff_B_bI7ElMqh7_2),.clk(gclk));
	jdff dff_B_g6H5fklB8_2(.din(w_dff_B_bI7ElMqh7_2),.dout(w_dff_B_g6H5fklB8_2),.clk(gclk));
	jdff dff_B_BGr92eYH7_2(.din(w_dff_B_g6H5fklB8_2),.dout(w_dff_B_BGr92eYH7_2),.clk(gclk));
	jdff dff_B_gT91Cokv4_2(.din(w_dff_B_BGr92eYH7_2),.dout(w_dff_B_gT91Cokv4_2),.clk(gclk));
	jdff dff_B_891SdkNe1_2(.din(w_dff_B_gT91Cokv4_2),.dout(w_dff_B_891SdkNe1_2),.clk(gclk));
	jdff dff_B_D53wKc4P8_2(.din(w_dff_B_891SdkNe1_2),.dout(w_dff_B_D53wKc4P8_2),.clk(gclk));
	jdff dff_B_9zP7aAPd5_2(.din(w_dff_B_D53wKc4P8_2),.dout(w_dff_B_9zP7aAPd5_2),.clk(gclk));
	jdff dff_B_BpSotqvJ2_2(.din(w_dff_B_9zP7aAPd5_2),.dout(w_dff_B_BpSotqvJ2_2),.clk(gclk));
	jdff dff_B_MwHRYxnq2_2(.din(w_dff_B_BpSotqvJ2_2),.dout(w_dff_B_MwHRYxnq2_2),.clk(gclk));
	jdff dff_B_io3x0prC6_2(.din(w_dff_B_MwHRYxnq2_2),.dout(w_dff_B_io3x0prC6_2),.clk(gclk));
	jdff dff_B_Hbpoq7ZI9_2(.din(n1703),.dout(w_dff_B_Hbpoq7ZI9_2),.clk(gclk));
	jdff dff_B_4K9zM5Yz5_2(.din(w_dff_B_Hbpoq7ZI9_2),.dout(w_dff_B_4K9zM5Yz5_2),.clk(gclk));
	jdff dff_B_GFpIGppL7_2(.din(w_dff_B_4K9zM5Yz5_2),.dout(w_dff_B_GFpIGppL7_2),.clk(gclk));
	jdff dff_B_uxbj7PjQ9_2(.din(w_dff_B_GFpIGppL7_2),.dout(w_dff_B_uxbj7PjQ9_2),.clk(gclk));
	jdff dff_B_aMkKiomu6_2(.din(w_dff_B_uxbj7PjQ9_2),.dout(w_dff_B_aMkKiomu6_2),.clk(gclk));
	jdff dff_B_3LSiX3WJ0_2(.din(w_dff_B_aMkKiomu6_2),.dout(w_dff_B_3LSiX3WJ0_2),.clk(gclk));
	jdff dff_B_WRnF1dbG2_2(.din(w_dff_B_3LSiX3WJ0_2),.dout(w_dff_B_WRnF1dbG2_2),.clk(gclk));
	jdff dff_B_YpoexdLl1_2(.din(w_dff_B_WRnF1dbG2_2),.dout(w_dff_B_YpoexdLl1_2),.clk(gclk));
	jdff dff_B_ONCPzIwO2_2(.din(w_dff_B_YpoexdLl1_2),.dout(w_dff_B_ONCPzIwO2_2),.clk(gclk));
	jdff dff_B_fAufSgq51_2(.din(w_dff_B_ONCPzIwO2_2),.dout(w_dff_B_fAufSgq51_2),.clk(gclk));
	jdff dff_B_l0RKTsTW7_2(.din(w_dff_B_fAufSgq51_2),.dout(w_dff_B_l0RKTsTW7_2),.clk(gclk));
	jdff dff_B_Z1c9yUfT4_2(.din(w_dff_B_l0RKTsTW7_2),.dout(w_dff_B_Z1c9yUfT4_2),.clk(gclk));
	jdff dff_B_uhLlVpYw7_2(.din(w_dff_B_Z1c9yUfT4_2),.dout(w_dff_B_uhLlVpYw7_2),.clk(gclk));
	jdff dff_B_PqVieLC61_2(.din(w_dff_B_uhLlVpYw7_2),.dout(w_dff_B_PqVieLC61_2),.clk(gclk));
	jdff dff_B_XDL8dbcl6_2(.din(w_dff_B_PqVieLC61_2),.dout(w_dff_B_XDL8dbcl6_2),.clk(gclk));
	jdff dff_B_INqlzx837_2(.din(w_dff_B_XDL8dbcl6_2),.dout(w_dff_B_INqlzx837_2),.clk(gclk));
	jdff dff_B_Hb9zzTJE2_2(.din(w_dff_B_INqlzx837_2),.dout(w_dff_B_Hb9zzTJE2_2),.clk(gclk));
	jdff dff_B_56KtMsJx4_2(.din(w_dff_B_Hb9zzTJE2_2),.dout(w_dff_B_56KtMsJx4_2),.clk(gclk));
	jdff dff_B_cvKGoKbM4_2(.din(w_dff_B_56KtMsJx4_2),.dout(w_dff_B_cvKGoKbM4_2),.clk(gclk));
	jdff dff_B_ZZCrM4em0_2(.din(w_dff_B_cvKGoKbM4_2),.dout(w_dff_B_ZZCrM4em0_2),.clk(gclk));
	jdff dff_B_YaQLFveC0_2(.din(w_dff_B_ZZCrM4em0_2),.dout(w_dff_B_YaQLFveC0_2),.clk(gclk));
	jdff dff_B_8UFTCT2L5_2(.din(w_dff_B_YaQLFveC0_2),.dout(w_dff_B_8UFTCT2L5_2),.clk(gclk));
	jdff dff_B_GICkqN6N8_2(.din(w_dff_B_8UFTCT2L5_2),.dout(w_dff_B_GICkqN6N8_2),.clk(gclk));
	jdff dff_B_6mlta9xD4_2(.din(w_dff_B_GICkqN6N8_2),.dout(w_dff_B_6mlta9xD4_2),.clk(gclk));
	jdff dff_B_d9rEHVlX3_2(.din(w_dff_B_6mlta9xD4_2),.dout(w_dff_B_d9rEHVlX3_2),.clk(gclk));
	jdff dff_B_NrsRAcI75_2(.din(w_dff_B_d9rEHVlX3_2),.dout(w_dff_B_NrsRAcI75_2),.clk(gclk));
	jdff dff_B_azmRlFvL6_2(.din(w_dff_B_NrsRAcI75_2),.dout(w_dff_B_azmRlFvL6_2),.clk(gclk));
	jdff dff_B_K0NkzhIB2_2(.din(w_dff_B_azmRlFvL6_2),.dout(w_dff_B_K0NkzhIB2_2),.clk(gclk));
	jdff dff_B_l6rcGCcK6_2(.din(w_dff_B_K0NkzhIB2_2),.dout(w_dff_B_l6rcGCcK6_2),.clk(gclk));
	jdff dff_B_8NaDjJ7R7_2(.din(w_dff_B_l6rcGCcK6_2),.dout(w_dff_B_8NaDjJ7R7_2),.clk(gclk));
	jdff dff_B_LEyHWSU28_2(.din(w_dff_B_8NaDjJ7R7_2),.dout(w_dff_B_LEyHWSU28_2),.clk(gclk));
	jdff dff_B_kwg80eUZ5_2(.din(w_dff_B_LEyHWSU28_2),.dout(w_dff_B_kwg80eUZ5_2),.clk(gclk));
	jdff dff_B_1raf0HVA7_2(.din(w_dff_B_kwg80eUZ5_2),.dout(w_dff_B_1raf0HVA7_2),.clk(gclk));
	jdff dff_B_290cngb96_2(.din(w_dff_B_1raf0HVA7_2),.dout(w_dff_B_290cngb96_2),.clk(gclk));
	jdff dff_B_UrUNSdwe0_2(.din(w_dff_B_290cngb96_2),.dout(w_dff_B_UrUNSdwe0_2),.clk(gclk));
	jdff dff_B_qX66UXMo7_2(.din(w_dff_B_UrUNSdwe0_2),.dout(w_dff_B_qX66UXMo7_2),.clk(gclk));
	jdff dff_B_tPxFV14z8_2(.din(w_dff_B_qX66UXMo7_2),.dout(w_dff_B_tPxFV14z8_2),.clk(gclk));
	jdff dff_B_Qd9CJMmI7_2(.din(w_dff_B_tPxFV14z8_2),.dout(w_dff_B_Qd9CJMmI7_2),.clk(gclk));
	jdff dff_B_1BzwHCJs7_2(.din(w_dff_B_Qd9CJMmI7_2),.dout(w_dff_B_1BzwHCJs7_2),.clk(gclk));
	jdff dff_B_x4Wou5S19_2(.din(w_dff_B_1BzwHCJs7_2),.dout(w_dff_B_x4Wou5S19_2),.clk(gclk));
	jdff dff_B_XXPJS6kv8_2(.din(w_dff_B_x4Wou5S19_2),.dout(w_dff_B_XXPJS6kv8_2),.clk(gclk));
	jdff dff_B_PBFYhsH57_2(.din(w_dff_B_XXPJS6kv8_2),.dout(w_dff_B_PBFYhsH57_2),.clk(gclk));
	jdff dff_B_vpqxp1Kb7_2(.din(n1702),.dout(w_dff_B_vpqxp1Kb7_2),.clk(gclk));
	jdff dff_B_9ydfEmg55_1(.din(n1700),.dout(w_dff_B_9ydfEmg55_1),.clk(gclk));
	jdff dff_B_ZMS2Vlgh3_2(.din(n1648),.dout(w_dff_B_ZMS2Vlgh3_2),.clk(gclk));
	jdff dff_B_SqCleVKN9_2(.din(w_dff_B_ZMS2Vlgh3_2),.dout(w_dff_B_SqCleVKN9_2),.clk(gclk));
	jdff dff_B_vK3Zz64v9_2(.din(w_dff_B_SqCleVKN9_2),.dout(w_dff_B_vK3Zz64v9_2),.clk(gclk));
	jdff dff_B_fXarcyMf0_2(.din(w_dff_B_vK3Zz64v9_2),.dout(w_dff_B_fXarcyMf0_2),.clk(gclk));
	jdff dff_B_Se9J04Kq3_2(.din(w_dff_B_fXarcyMf0_2),.dout(w_dff_B_Se9J04Kq3_2),.clk(gclk));
	jdff dff_B_zFJDWkud6_2(.din(w_dff_B_Se9J04Kq3_2),.dout(w_dff_B_zFJDWkud6_2),.clk(gclk));
	jdff dff_B_jJShNd7i2_2(.din(w_dff_B_zFJDWkud6_2),.dout(w_dff_B_jJShNd7i2_2),.clk(gclk));
	jdff dff_B_toKTsgxP8_2(.din(w_dff_B_jJShNd7i2_2),.dout(w_dff_B_toKTsgxP8_2),.clk(gclk));
	jdff dff_B_d9j0DKPJ6_2(.din(w_dff_B_toKTsgxP8_2),.dout(w_dff_B_d9j0DKPJ6_2),.clk(gclk));
	jdff dff_B_Nl3ZX58E8_2(.din(w_dff_B_d9j0DKPJ6_2),.dout(w_dff_B_Nl3ZX58E8_2),.clk(gclk));
	jdff dff_B_gIEUCPnm6_2(.din(w_dff_B_Nl3ZX58E8_2),.dout(w_dff_B_gIEUCPnm6_2),.clk(gclk));
	jdff dff_B_DRaPI8Wl7_2(.din(w_dff_B_gIEUCPnm6_2),.dout(w_dff_B_DRaPI8Wl7_2),.clk(gclk));
	jdff dff_B_kwuV2xiU5_2(.din(w_dff_B_DRaPI8Wl7_2),.dout(w_dff_B_kwuV2xiU5_2),.clk(gclk));
	jdff dff_B_Xk6vgI0U5_2(.din(w_dff_B_kwuV2xiU5_2),.dout(w_dff_B_Xk6vgI0U5_2),.clk(gclk));
	jdff dff_B_hq6ZSFrN0_2(.din(w_dff_B_Xk6vgI0U5_2),.dout(w_dff_B_hq6ZSFrN0_2),.clk(gclk));
	jdff dff_B_F3EP3AeZ4_2(.din(w_dff_B_hq6ZSFrN0_2),.dout(w_dff_B_F3EP3AeZ4_2),.clk(gclk));
	jdff dff_B_LAizMQ1M0_2(.din(w_dff_B_F3EP3AeZ4_2),.dout(w_dff_B_LAizMQ1M0_2),.clk(gclk));
	jdff dff_B_9F0VmLuT0_2(.din(w_dff_B_LAizMQ1M0_2),.dout(w_dff_B_9F0VmLuT0_2),.clk(gclk));
	jdff dff_B_njGHyIku0_2(.din(w_dff_B_9F0VmLuT0_2),.dout(w_dff_B_njGHyIku0_2),.clk(gclk));
	jdff dff_B_2xhwFLI90_2(.din(w_dff_B_njGHyIku0_2),.dout(w_dff_B_2xhwFLI90_2),.clk(gclk));
	jdff dff_B_s1obosXv1_2(.din(w_dff_B_2xhwFLI90_2),.dout(w_dff_B_s1obosXv1_2),.clk(gclk));
	jdff dff_B_E3TtFOE52_2(.din(w_dff_B_s1obosXv1_2),.dout(w_dff_B_E3TtFOE52_2),.clk(gclk));
	jdff dff_B_mGGnLoVQ7_2(.din(w_dff_B_E3TtFOE52_2),.dout(w_dff_B_mGGnLoVQ7_2),.clk(gclk));
	jdff dff_B_lJggEX4b9_2(.din(w_dff_B_mGGnLoVQ7_2),.dout(w_dff_B_lJggEX4b9_2),.clk(gclk));
	jdff dff_B_OaSbouYj8_2(.din(w_dff_B_lJggEX4b9_2),.dout(w_dff_B_OaSbouYj8_2),.clk(gclk));
	jdff dff_B_HLrOsYkm2_2(.din(w_dff_B_OaSbouYj8_2),.dout(w_dff_B_HLrOsYkm2_2),.clk(gclk));
	jdff dff_B_lTtlyRh95_2(.din(w_dff_B_HLrOsYkm2_2),.dout(w_dff_B_lTtlyRh95_2),.clk(gclk));
	jdff dff_B_crmkhb9j1_2(.din(w_dff_B_lTtlyRh95_2),.dout(w_dff_B_crmkhb9j1_2),.clk(gclk));
	jdff dff_B_AmQhiB013_2(.din(w_dff_B_crmkhb9j1_2),.dout(w_dff_B_AmQhiB013_2),.clk(gclk));
	jdff dff_B_iZLbhxoo7_2(.din(w_dff_B_AmQhiB013_2),.dout(w_dff_B_iZLbhxoo7_2),.clk(gclk));
	jdff dff_B_qwtc29Jh7_2(.din(w_dff_B_iZLbhxoo7_2),.dout(w_dff_B_qwtc29Jh7_2),.clk(gclk));
	jdff dff_B_nC1IgaNQ6_2(.din(w_dff_B_qwtc29Jh7_2),.dout(w_dff_B_nC1IgaNQ6_2),.clk(gclk));
	jdff dff_B_OpapyPtB9_2(.din(w_dff_B_nC1IgaNQ6_2),.dout(w_dff_B_OpapyPtB9_2),.clk(gclk));
	jdff dff_B_tILYIIsp6_2(.din(w_dff_B_OpapyPtB9_2),.dout(w_dff_B_tILYIIsp6_2),.clk(gclk));
	jdff dff_B_sQjQBrpf0_2(.din(w_dff_B_tILYIIsp6_2),.dout(w_dff_B_sQjQBrpf0_2),.clk(gclk));
	jdff dff_B_OG30zOvl3_2(.din(w_dff_B_sQjQBrpf0_2),.dout(w_dff_B_OG30zOvl3_2),.clk(gclk));
	jdff dff_B_2NPYnQza8_2(.din(w_dff_B_OG30zOvl3_2),.dout(w_dff_B_2NPYnQza8_2),.clk(gclk));
	jdff dff_B_qEOmvMIj2_2(.din(w_dff_B_2NPYnQza8_2),.dout(w_dff_B_qEOmvMIj2_2),.clk(gclk));
	jdff dff_B_ICMzF6Jr6_2(.din(w_dff_B_qEOmvMIj2_2),.dout(w_dff_B_ICMzF6Jr6_2),.clk(gclk));
	jdff dff_B_X7xodnwm1_1(.din(n1654),.dout(w_dff_B_X7xodnwm1_1),.clk(gclk));
	jdff dff_B_nlXGNjIF6_1(.din(w_dff_B_X7xodnwm1_1),.dout(w_dff_B_nlXGNjIF6_1),.clk(gclk));
	jdff dff_B_0NPQCha60_2(.din(n1653),.dout(w_dff_B_0NPQCha60_2),.clk(gclk));
	jdff dff_B_n18SuO5a3_2(.din(w_dff_B_0NPQCha60_2),.dout(w_dff_B_n18SuO5a3_2),.clk(gclk));
	jdff dff_B_t43B5j8c5_2(.din(w_dff_B_n18SuO5a3_2),.dout(w_dff_B_t43B5j8c5_2),.clk(gclk));
	jdff dff_B_F84NreC82_2(.din(w_dff_B_t43B5j8c5_2),.dout(w_dff_B_F84NreC82_2),.clk(gclk));
	jdff dff_B_AOkS4PYT5_2(.din(w_dff_B_F84NreC82_2),.dout(w_dff_B_AOkS4PYT5_2),.clk(gclk));
	jdff dff_B_SmYUXrUs2_2(.din(w_dff_B_AOkS4PYT5_2),.dout(w_dff_B_SmYUXrUs2_2),.clk(gclk));
	jdff dff_B_AnSy7udP7_2(.din(w_dff_B_SmYUXrUs2_2),.dout(w_dff_B_AnSy7udP7_2),.clk(gclk));
	jdff dff_B_S0RfVLwC6_2(.din(w_dff_B_AnSy7udP7_2),.dout(w_dff_B_S0RfVLwC6_2),.clk(gclk));
	jdff dff_B_BDYfIA1O9_2(.din(w_dff_B_S0RfVLwC6_2),.dout(w_dff_B_BDYfIA1O9_2),.clk(gclk));
	jdff dff_B_haaLgri37_2(.din(w_dff_B_BDYfIA1O9_2),.dout(w_dff_B_haaLgri37_2),.clk(gclk));
	jdff dff_B_cL3Pn4GH0_2(.din(w_dff_B_haaLgri37_2),.dout(w_dff_B_cL3Pn4GH0_2),.clk(gclk));
	jdff dff_B_J0Z3k1ML2_2(.din(w_dff_B_cL3Pn4GH0_2),.dout(w_dff_B_J0Z3k1ML2_2),.clk(gclk));
	jdff dff_B_EJoyquFC8_2(.din(w_dff_B_J0Z3k1ML2_2),.dout(w_dff_B_EJoyquFC8_2),.clk(gclk));
	jdff dff_B_ZDL4Brfd7_2(.din(w_dff_B_EJoyquFC8_2),.dout(w_dff_B_ZDL4Brfd7_2),.clk(gclk));
	jdff dff_B_TETDjt7T8_2(.din(w_dff_B_ZDL4Brfd7_2),.dout(w_dff_B_TETDjt7T8_2),.clk(gclk));
	jdff dff_B_knKaKNxA8_2(.din(w_dff_B_TETDjt7T8_2),.dout(w_dff_B_knKaKNxA8_2),.clk(gclk));
	jdff dff_B_9roTWaUf2_2(.din(w_dff_B_knKaKNxA8_2),.dout(w_dff_B_9roTWaUf2_2),.clk(gclk));
	jdff dff_B_EKtsm1xm8_2(.din(w_dff_B_9roTWaUf2_2),.dout(w_dff_B_EKtsm1xm8_2),.clk(gclk));
	jdff dff_B_Z3xbjfB47_2(.din(w_dff_B_EKtsm1xm8_2),.dout(w_dff_B_Z3xbjfB47_2),.clk(gclk));
	jdff dff_B_8xkb2ZLw7_2(.din(w_dff_B_Z3xbjfB47_2),.dout(w_dff_B_8xkb2ZLw7_2),.clk(gclk));
	jdff dff_B_29d2u9qo9_2(.din(w_dff_B_8xkb2ZLw7_2),.dout(w_dff_B_29d2u9qo9_2),.clk(gclk));
	jdff dff_B_irvvmkuX2_2(.din(w_dff_B_29d2u9qo9_2),.dout(w_dff_B_irvvmkuX2_2),.clk(gclk));
	jdff dff_B_oX2YHHF74_2(.din(w_dff_B_irvvmkuX2_2),.dout(w_dff_B_oX2YHHF74_2),.clk(gclk));
	jdff dff_B_uHYM0hIk7_2(.din(w_dff_B_oX2YHHF74_2),.dout(w_dff_B_uHYM0hIk7_2),.clk(gclk));
	jdff dff_B_swMWQBmI5_2(.din(w_dff_B_uHYM0hIk7_2),.dout(w_dff_B_swMWQBmI5_2),.clk(gclk));
	jdff dff_B_bogDKblD1_2(.din(w_dff_B_swMWQBmI5_2),.dout(w_dff_B_bogDKblD1_2),.clk(gclk));
	jdff dff_B_WnXDne0P8_2(.din(w_dff_B_bogDKblD1_2),.dout(w_dff_B_WnXDne0P8_2),.clk(gclk));
	jdff dff_B_gT2D0SUk3_2(.din(w_dff_B_WnXDne0P8_2),.dout(w_dff_B_gT2D0SUk3_2),.clk(gclk));
	jdff dff_B_TgMPwA4Q2_2(.din(w_dff_B_gT2D0SUk3_2),.dout(w_dff_B_TgMPwA4Q2_2),.clk(gclk));
	jdff dff_B_2yjlCh1N1_2(.din(w_dff_B_TgMPwA4Q2_2),.dout(w_dff_B_2yjlCh1N1_2),.clk(gclk));
	jdff dff_B_rbD5szq79_2(.din(w_dff_B_2yjlCh1N1_2),.dout(w_dff_B_rbD5szq79_2),.clk(gclk));
	jdff dff_B_15H3kabV2_2(.din(w_dff_B_rbD5szq79_2),.dout(w_dff_B_15H3kabV2_2),.clk(gclk));
	jdff dff_B_fIMasrvF3_2(.din(w_dff_B_15H3kabV2_2),.dout(w_dff_B_fIMasrvF3_2),.clk(gclk));
	jdff dff_B_0hxaG8rN4_2(.din(w_dff_B_fIMasrvF3_2),.dout(w_dff_B_0hxaG8rN4_2),.clk(gclk));
	jdff dff_B_pwCNOjhA3_2(.din(w_dff_B_0hxaG8rN4_2),.dout(w_dff_B_pwCNOjhA3_2),.clk(gclk));
	jdff dff_B_ef7mrUa07_2(.din(w_dff_B_pwCNOjhA3_2),.dout(w_dff_B_ef7mrUa07_2),.clk(gclk));
	jdff dff_B_D0bcy96T8_2(.din(n1652),.dout(w_dff_B_D0bcy96T8_2),.clk(gclk));
	jdff dff_B_7eP7DN1Y4_2(.din(w_dff_B_D0bcy96T8_2),.dout(w_dff_B_7eP7DN1Y4_2),.clk(gclk));
	jdff dff_B_rCVC8Nrv3_2(.din(w_dff_B_7eP7DN1Y4_2),.dout(w_dff_B_rCVC8Nrv3_2),.clk(gclk));
	jdff dff_B_SMQlLS9G7_2(.din(w_dff_B_rCVC8Nrv3_2),.dout(w_dff_B_SMQlLS9G7_2),.clk(gclk));
	jdff dff_B_KwZlrEUg5_2(.din(w_dff_B_SMQlLS9G7_2),.dout(w_dff_B_KwZlrEUg5_2),.clk(gclk));
	jdff dff_B_8sU7tmQn6_2(.din(w_dff_B_KwZlrEUg5_2),.dout(w_dff_B_8sU7tmQn6_2),.clk(gclk));
	jdff dff_B_bUJCqNGF9_2(.din(w_dff_B_8sU7tmQn6_2),.dout(w_dff_B_bUJCqNGF9_2),.clk(gclk));
	jdff dff_B_wTpbPT1U3_2(.din(w_dff_B_bUJCqNGF9_2),.dout(w_dff_B_wTpbPT1U3_2),.clk(gclk));
	jdff dff_B_hvL0KFLo6_2(.din(w_dff_B_wTpbPT1U3_2),.dout(w_dff_B_hvL0KFLo6_2),.clk(gclk));
	jdff dff_B_tYBrYaQC0_2(.din(w_dff_B_hvL0KFLo6_2),.dout(w_dff_B_tYBrYaQC0_2),.clk(gclk));
	jdff dff_B_Q6sD4Qeb5_2(.din(w_dff_B_tYBrYaQC0_2),.dout(w_dff_B_Q6sD4Qeb5_2),.clk(gclk));
	jdff dff_B_wff3Dzjk0_2(.din(w_dff_B_Q6sD4Qeb5_2),.dout(w_dff_B_wff3Dzjk0_2),.clk(gclk));
	jdff dff_B_al9gX4Yh0_2(.din(w_dff_B_wff3Dzjk0_2),.dout(w_dff_B_al9gX4Yh0_2),.clk(gclk));
	jdff dff_B_0asvR0wp9_2(.din(w_dff_B_al9gX4Yh0_2),.dout(w_dff_B_0asvR0wp9_2),.clk(gclk));
	jdff dff_B_D7XTMrYT5_2(.din(w_dff_B_0asvR0wp9_2),.dout(w_dff_B_D7XTMrYT5_2),.clk(gclk));
	jdff dff_B_4zdIWGLF7_2(.din(w_dff_B_D7XTMrYT5_2),.dout(w_dff_B_4zdIWGLF7_2),.clk(gclk));
	jdff dff_B_mV09WgCd9_2(.din(w_dff_B_4zdIWGLF7_2),.dout(w_dff_B_mV09WgCd9_2),.clk(gclk));
	jdff dff_B_OZxWyJjY5_2(.din(w_dff_B_mV09WgCd9_2),.dout(w_dff_B_OZxWyJjY5_2),.clk(gclk));
	jdff dff_B_ExYSN7yU2_2(.din(w_dff_B_OZxWyJjY5_2),.dout(w_dff_B_ExYSN7yU2_2),.clk(gclk));
	jdff dff_B_OGkyOXb97_2(.din(w_dff_B_ExYSN7yU2_2),.dout(w_dff_B_OGkyOXb97_2),.clk(gclk));
	jdff dff_B_bCIaheV48_2(.din(w_dff_B_OGkyOXb97_2),.dout(w_dff_B_bCIaheV48_2),.clk(gclk));
	jdff dff_B_cAWOpRNm5_2(.din(w_dff_B_bCIaheV48_2),.dout(w_dff_B_cAWOpRNm5_2),.clk(gclk));
	jdff dff_B_ZtgcNjdf2_2(.din(w_dff_B_cAWOpRNm5_2),.dout(w_dff_B_ZtgcNjdf2_2),.clk(gclk));
	jdff dff_B_PK76ddSN5_2(.din(w_dff_B_ZtgcNjdf2_2),.dout(w_dff_B_PK76ddSN5_2),.clk(gclk));
	jdff dff_B_rl7TjIv99_2(.din(w_dff_B_PK76ddSN5_2),.dout(w_dff_B_rl7TjIv99_2),.clk(gclk));
	jdff dff_B_lR7Wf5kq2_2(.din(w_dff_B_rl7TjIv99_2),.dout(w_dff_B_lR7Wf5kq2_2),.clk(gclk));
	jdff dff_B_EkuLaFIM1_2(.din(w_dff_B_lR7Wf5kq2_2),.dout(w_dff_B_EkuLaFIM1_2),.clk(gclk));
	jdff dff_B_GLbYpbuX3_2(.din(w_dff_B_EkuLaFIM1_2),.dout(w_dff_B_GLbYpbuX3_2),.clk(gclk));
	jdff dff_B_QuGF6xXi6_2(.din(w_dff_B_GLbYpbuX3_2),.dout(w_dff_B_QuGF6xXi6_2),.clk(gclk));
	jdff dff_B_BR0o74Rc7_2(.din(w_dff_B_QuGF6xXi6_2),.dout(w_dff_B_BR0o74Rc7_2),.clk(gclk));
	jdff dff_B_Ktywyk4b1_2(.din(w_dff_B_BR0o74Rc7_2),.dout(w_dff_B_Ktywyk4b1_2),.clk(gclk));
	jdff dff_B_yK91rIF66_2(.din(w_dff_B_Ktywyk4b1_2),.dout(w_dff_B_yK91rIF66_2),.clk(gclk));
	jdff dff_B_Q9QehKZ13_2(.din(w_dff_B_yK91rIF66_2),.dout(w_dff_B_Q9QehKZ13_2),.clk(gclk));
	jdff dff_B_QohVCJko7_2(.din(w_dff_B_Q9QehKZ13_2),.dout(w_dff_B_QohVCJko7_2),.clk(gclk));
	jdff dff_B_bHbVmv3S5_2(.din(w_dff_B_QohVCJko7_2),.dout(w_dff_B_bHbVmv3S5_2),.clk(gclk));
	jdff dff_B_pPjyttP71_2(.din(w_dff_B_bHbVmv3S5_2),.dout(w_dff_B_pPjyttP71_2),.clk(gclk));
	jdff dff_B_UBiOOzAm4_2(.din(w_dff_B_pPjyttP71_2),.dout(w_dff_B_UBiOOzAm4_2),.clk(gclk));
	jdff dff_B_O76LVzGe3_2(.din(w_dff_B_UBiOOzAm4_2),.dout(w_dff_B_O76LVzGe3_2),.clk(gclk));
	jdff dff_B_7ewJLvDw1_2(.din(n1651),.dout(w_dff_B_7ewJLvDw1_2),.clk(gclk));
	jdff dff_B_ZKC0WEWM3_1(.din(n1649),.dout(w_dff_B_ZKC0WEWM3_1),.clk(gclk));
	jdff dff_B_BNC8kMfX0_2(.din(n1591),.dout(w_dff_B_BNC8kMfX0_2),.clk(gclk));
	jdff dff_B_2AFvZx8t7_2(.din(w_dff_B_BNC8kMfX0_2),.dout(w_dff_B_2AFvZx8t7_2),.clk(gclk));
	jdff dff_B_vdvEouQM7_2(.din(w_dff_B_2AFvZx8t7_2),.dout(w_dff_B_vdvEouQM7_2),.clk(gclk));
	jdff dff_B_hoio2uhr0_2(.din(w_dff_B_vdvEouQM7_2),.dout(w_dff_B_hoio2uhr0_2),.clk(gclk));
	jdff dff_B_iOV2Hjtg3_2(.din(w_dff_B_hoio2uhr0_2),.dout(w_dff_B_iOV2Hjtg3_2),.clk(gclk));
	jdff dff_B_IXm6Ny388_2(.din(w_dff_B_iOV2Hjtg3_2),.dout(w_dff_B_IXm6Ny388_2),.clk(gclk));
	jdff dff_B_2ukPKuky7_2(.din(w_dff_B_IXm6Ny388_2),.dout(w_dff_B_2ukPKuky7_2),.clk(gclk));
	jdff dff_B_tSSubhgk2_2(.din(w_dff_B_2ukPKuky7_2),.dout(w_dff_B_tSSubhgk2_2),.clk(gclk));
	jdff dff_B_Rc69CJUn5_2(.din(w_dff_B_tSSubhgk2_2),.dout(w_dff_B_Rc69CJUn5_2),.clk(gclk));
	jdff dff_B_Xu3So4dr6_2(.din(w_dff_B_Rc69CJUn5_2),.dout(w_dff_B_Xu3So4dr6_2),.clk(gclk));
	jdff dff_B_DItVifN45_2(.din(w_dff_B_Xu3So4dr6_2),.dout(w_dff_B_DItVifN45_2),.clk(gclk));
	jdff dff_B_eyvana3L5_2(.din(w_dff_B_DItVifN45_2),.dout(w_dff_B_eyvana3L5_2),.clk(gclk));
	jdff dff_B_HLyMGbqo1_2(.din(w_dff_B_eyvana3L5_2),.dout(w_dff_B_HLyMGbqo1_2),.clk(gclk));
	jdff dff_B_O1tkoqEf2_2(.din(w_dff_B_HLyMGbqo1_2),.dout(w_dff_B_O1tkoqEf2_2),.clk(gclk));
	jdff dff_B_EfE2ysZA5_2(.din(w_dff_B_O1tkoqEf2_2),.dout(w_dff_B_EfE2ysZA5_2),.clk(gclk));
	jdff dff_B_0dS5CT4o2_2(.din(w_dff_B_EfE2ysZA5_2),.dout(w_dff_B_0dS5CT4o2_2),.clk(gclk));
	jdff dff_B_wXc8zhX84_2(.din(w_dff_B_0dS5CT4o2_2),.dout(w_dff_B_wXc8zhX84_2),.clk(gclk));
	jdff dff_B_clctTt8x1_2(.din(w_dff_B_wXc8zhX84_2),.dout(w_dff_B_clctTt8x1_2),.clk(gclk));
	jdff dff_B_WWG48nvQ1_2(.din(w_dff_B_clctTt8x1_2),.dout(w_dff_B_WWG48nvQ1_2),.clk(gclk));
	jdff dff_B_ez0DO1L38_2(.din(w_dff_B_WWG48nvQ1_2),.dout(w_dff_B_ez0DO1L38_2),.clk(gclk));
	jdff dff_B_2CWKtBYO2_2(.din(w_dff_B_ez0DO1L38_2),.dout(w_dff_B_2CWKtBYO2_2),.clk(gclk));
	jdff dff_B_oCquieuX0_2(.din(w_dff_B_2CWKtBYO2_2),.dout(w_dff_B_oCquieuX0_2),.clk(gclk));
	jdff dff_B_6yu15raF8_2(.din(w_dff_B_oCquieuX0_2),.dout(w_dff_B_6yu15raF8_2),.clk(gclk));
	jdff dff_B_nsPbGACH3_2(.din(w_dff_B_6yu15raF8_2),.dout(w_dff_B_nsPbGACH3_2),.clk(gclk));
	jdff dff_B_4HnGiibP4_2(.din(w_dff_B_nsPbGACH3_2),.dout(w_dff_B_4HnGiibP4_2),.clk(gclk));
	jdff dff_B_B62lF1dI8_2(.din(w_dff_B_4HnGiibP4_2),.dout(w_dff_B_B62lF1dI8_2),.clk(gclk));
	jdff dff_B_cGkTm7iv7_2(.din(w_dff_B_B62lF1dI8_2),.dout(w_dff_B_cGkTm7iv7_2),.clk(gclk));
	jdff dff_B_I1xc5ct55_2(.din(w_dff_B_cGkTm7iv7_2),.dout(w_dff_B_I1xc5ct55_2),.clk(gclk));
	jdff dff_B_2h7iqjcF0_2(.din(w_dff_B_I1xc5ct55_2),.dout(w_dff_B_2h7iqjcF0_2),.clk(gclk));
	jdff dff_B_0ZHmcmaX0_2(.din(w_dff_B_2h7iqjcF0_2),.dout(w_dff_B_0ZHmcmaX0_2),.clk(gclk));
	jdff dff_B_FmNj1nCT7_2(.din(w_dff_B_0ZHmcmaX0_2),.dout(w_dff_B_FmNj1nCT7_2),.clk(gclk));
	jdff dff_B_nGKmKZuY9_2(.din(w_dff_B_FmNj1nCT7_2),.dout(w_dff_B_nGKmKZuY9_2),.clk(gclk));
	jdff dff_B_2JtS07gc5_2(.din(w_dff_B_nGKmKZuY9_2),.dout(w_dff_B_2JtS07gc5_2),.clk(gclk));
	jdff dff_B_pzdKgBdT1_2(.din(w_dff_B_2JtS07gc5_2),.dout(w_dff_B_pzdKgBdT1_2),.clk(gclk));
	jdff dff_B_rdWGEVfD7_2(.din(w_dff_B_pzdKgBdT1_2),.dout(w_dff_B_rdWGEVfD7_2),.clk(gclk));
	jdff dff_B_4zw2Wckk3_1(.din(n1597),.dout(w_dff_B_4zw2Wckk3_1),.clk(gclk));
	jdff dff_B_jpgEFxr40_1(.din(w_dff_B_4zw2Wckk3_1),.dout(w_dff_B_jpgEFxr40_1),.clk(gclk));
	jdff dff_B_7FcKe92B1_2(.din(n1596),.dout(w_dff_B_7FcKe92B1_2),.clk(gclk));
	jdff dff_B_gt0Mjkak6_2(.din(w_dff_B_7FcKe92B1_2),.dout(w_dff_B_gt0Mjkak6_2),.clk(gclk));
	jdff dff_B_6T9qt8P13_2(.din(w_dff_B_gt0Mjkak6_2),.dout(w_dff_B_6T9qt8P13_2),.clk(gclk));
	jdff dff_B_NcJYkPxn7_2(.din(w_dff_B_6T9qt8P13_2),.dout(w_dff_B_NcJYkPxn7_2),.clk(gclk));
	jdff dff_B_VDJSfolT0_2(.din(w_dff_B_NcJYkPxn7_2),.dout(w_dff_B_VDJSfolT0_2),.clk(gclk));
	jdff dff_B_s9LaQPmQ2_2(.din(w_dff_B_VDJSfolT0_2),.dout(w_dff_B_s9LaQPmQ2_2),.clk(gclk));
	jdff dff_B_8tIsUzxP2_2(.din(w_dff_B_s9LaQPmQ2_2),.dout(w_dff_B_8tIsUzxP2_2),.clk(gclk));
	jdff dff_B_7tuKtVzO5_2(.din(w_dff_B_8tIsUzxP2_2),.dout(w_dff_B_7tuKtVzO5_2),.clk(gclk));
	jdff dff_B_r6x1NBrr6_2(.din(w_dff_B_7tuKtVzO5_2),.dout(w_dff_B_r6x1NBrr6_2),.clk(gclk));
	jdff dff_B_08WEnwmU5_2(.din(w_dff_B_r6x1NBrr6_2),.dout(w_dff_B_08WEnwmU5_2),.clk(gclk));
	jdff dff_B_Gcelk3Ma2_2(.din(w_dff_B_08WEnwmU5_2),.dout(w_dff_B_Gcelk3Ma2_2),.clk(gclk));
	jdff dff_B_UDEQTZPQ9_2(.din(w_dff_B_Gcelk3Ma2_2),.dout(w_dff_B_UDEQTZPQ9_2),.clk(gclk));
	jdff dff_B_S9xv1bjO3_2(.din(w_dff_B_UDEQTZPQ9_2),.dout(w_dff_B_S9xv1bjO3_2),.clk(gclk));
	jdff dff_B_NFUzX4r40_2(.din(w_dff_B_S9xv1bjO3_2),.dout(w_dff_B_NFUzX4r40_2),.clk(gclk));
	jdff dff_B_RC8upy0Y3_2(.din(w_dff_B_NFUzX4r40_2),.dout(w_dff_B_RC8upy0Y3_2),.clk(gclk));
	jdff dff_B_UH0dkvVo6_2(.din(w_dff_B_RC8upy0Y3_2),.dout(w_dff_B_UH0dkvVo6_2),.clk(gclk));
	jdff dff_B_2dZ8ulhM2_2(.din(w_dff_B_UH0dkvVo6_2),.dout(w_dff_B_2dZ8ulhM2_2),.clk(gclk));
	jdff dff_B_KyfxT94a6_2(.din(w_dff_B_2dZ8ulhM2_2),.dout(w_dff_B_KyfxT94a6_2),.clk(gclk));
	jdff dff_B_vVeQjTaB7_2(.din(w_dff_B_KyfxT94a6_2),.dout(w_dff_B_vVeQjTaB7_2),.clk(gclk));
	jdff dff_B_fHdOZAZR9_2(.din(w_dff_B_vVeQjTaB7_2),.dout(w_dff_B_fHdOZAZR9_2),.clk(gclk));
	jdff dff_B_aQQlbn8U9_2(.din(w_dff_B_fHdOZAZR9_2),.dout(w_dff_B_aQQlbn8U9_2),.clk(gclk));
	jdff dff_B_Pemg0udW0_2(.din(w_dff_B_aQQlbn8U9_2),.dout(w_dff_B_Pemg0udW0_2),.clk(gclk));
	jdff dff_B_gQLaWQFL5_2(.din(w_dff_B_Pemg0udW0_2),.dout(w_dff_B_gQLaWQFL5_2),.clk(gclk));
	jdff dff_B_CUdGUCs62_2(.din(w_dff_B_gQLaWQFL5_2),.dout(w_dff_B_CUdGUCs62_2),.clk(gclk));
	jdff dff_B_6RuOt6mp1_2(.din(w_dff_B_CUdGUCs62_2),.dout(w_dff_B_6RuOt6mp1_2),.clk(gclk));
	jdff dff_B_AmNTbTcf3_2(.din(w_dff_B_6RuOt6mp1_2),.dout(w_dff_B_AmNTbTcf3_2),.clk(gclk));
	jdff dff_B_G0a8hd3Z7_2(.din(w_dff_B_AmNTbTcf3_2),.dout(w_dff_B_G0a8hd3Z7_2),.clk(gclk));
	jdff dff_B_hYWoXIzD2_2(.din(w_dff_B_G0a8hd3Z7_2),.dout(w_dff_B_hYWoXIzD2_2),.clk(gclk));
	jdff dff_B_tCIblQOO6_2(.din(w_dff_B_hYWoXIzD2_2),.dout(w_dff_B_tCIblQOO6_2),.clk(gclk));
	jdff dff_B_zxD86mAu4_2(.din(w_dff_B_tCIblQOO6_2),.dout(w_dff_B_zxD86mAu4_2),.clk(gclk));
	jdff dff_B_5k0XQMr77_2(.din(w_dff_B_zxD86mAu4_2),.dout(w_dff_B_5k0XQMr77_2),.clk(gclk));
	jdff dff_B_j3hSLS2j5_2(.din(w_dff_B_5k0XQMr77_2),.dout(w_dff_B_j3hSLS2j5_2),.clk(gclk));
	jdff dff_B_bvtdjLpj9_2(.din(n1595),.dout(w_dff_B_bvtdjLpj9_2),.clk(gclk));
	jdff dff_B_hCIdtIQp0_2(.din(w_dff_B_bvtdjLpj9_2),.dout(w_dff_B_hCIdtIQp0_2),.clk(gclk));
	jdff dff_B_c9LG3Gxg3_2(.din(w_dff_B_hCIdtIQp0_2),.dout(w_dff_B_c9LG3Gxg3_2),.clk(gclk));
	jdff dff_B_TBEWTNIU2_2(.din(w_dff_B_c9LG3Gxg3_2),.dout(w_dff_B_TBEWTNIU2_2),.clk(gclk));
	jdff dff_B_9mjOgcBi6_2(.din(w_dff_B_TBEWTNIU2_2),.dout(w_dff_B_9mjOgcBi6_2),.clk(gclk));
	jdff dff_B_b8GU8LQn6_2(.din(w_dff_B_9mjOgcBi6_2),.dout(w_dff_B_b8GU8LQn6_2),.clk(gclk));
	jdff dff_B_055S17Mu4_2(.din(w_dff_B_b8GU8LQn6_2),.dout(w_dff_B_055S17Mu4_2),.clk(gclk));
	jdff dff_B_nglLsSAt2_2(.din(w_dff_B_055S17Mu4_2),.dout(w_dff_B_nglLsSAt2_2),.clk(gclk));
	jdff dff_B_hs6kqYo93_2(.din(w_dff_B_nglLsSAt2_2),.dout(w_dff_B_hs6kqYo93_2),.clk(gclk));
	jdff dff_B_hcVUC0IR4_2(.din(w_dff_B_hs6kqYo93_2),.dout(w_dff_B_hcVUC0IR4_2),.clk(gclk));
	jdff dff_B_1PL7pokc7_2(.din(w_dff_B_hcVUC0IR4_2),.dout(w_dff_B_1PL7pokc7_2),.clk(gclk));
	jdff dff_B_Qf8KEaym9_2(.din(w_dff_B_1PL7pokc7_2),.dout(w_dff_B_Qf8KEaym9_2),.clk(gclk));
	jdff dff_B_2jSFyZfJ7_2(.din(w_dff_B_Qf8KEaym9_2),.dout(w_dff_B_2jSFyZfJ7_2),.clk(gclk));
	jdff dff_B_gZOxMbrp7_2(.din(w_dff_B_2jSFyZfJ7_2),.dout(w_dff_B_gZOxMbrp7_2),.clk(gclk));
	jdff dff_B_v0vdtG773_2(.din(w_dff_B_gZOxMbrp7_2),.dout(w_dff_B_v0vdtG773_2),.clk(gclk));
	jdff dff_B_tvge0oW91_2(.din(w_dff_B_v0vdtG773_2),.dout(w_dff_B_tvge0oW91_2),.clk(gclk));
	jdff dff_B_sFk0Ya3X5_2(.din(w_dff_B_tvge0oW91_2),.dout(w_dff_B_sFk0Ya3X5_2),.clk(gclk));
	jdff dff_B_rZVCU9z56_2(.din(w_dff_B_sFk0Ya3X5_2),.dout(w_dff_B_rZVCU9z56_2),.clk(gclk));
	jdff dff_B_YOGAjIAm8_2(.din(w_dff_B_rZVCU9z56_2),.dout(w_dff_B_YOGAjIAm8_2),.clk(gclk));
	jdff dff_B_qwYDQuNE9_2(.din(w_dff_B_YOGAjIAm8_2),.dout(w_dff_B_qwYDQuNE9_2),.clk(gclk));
	jdff dff_B_3JTkb7hs3_2(.din(w_dff_B_qwYDQuNE9_2),.dout(w_dff_B_3JTkb7hs3_2),.clk(gclk));
	jdff dff_B_V4sVBbUs0_2(.din(w_dff_B_3JTkb7hs3_2),.dout(w_dff_B_V4sVBbUs0_2),.clk(gclk));
	jdff dff_B_iKiZRmR45_2(.din(w_dff_B_V4sVBbUs0_2),.dout(w_dff_B_iKiZRmR45_2),.clk(gclk));
	jdff dff_B_7bkktzIr1_2(.din(w_dff_B_iKiZRmR45_2),.dout(w_dff_B_7bkktzIr1_2),.clk(gclk));
	jdff dff_B_5rD8c5gv0_2(.din(w_dff_B_7bkktzIr1_2),.dout(w_dff_B_5rD8c5gv0_2),.clk(gclk));
	jdff dff_B_11dv5sD72_2(.din(w_dff_B_5rD8c5gv0_2),.dout(w_dff_B_11dv5sD72_2),.clk(gclk));
	jdff dff_B_4CrBkHdb8_2(.din(w_dff_B_11dv5sD72_2),.dout(w_dff_B_4CrBkHdb8_2),.clk(gclk));
	jdff dff_B_OMidsCf33_2(.din(w_dff_B_4CrBkHdb8_2),.dout(w_dff_B_OMidsCf33_2),.clk(gclk));
	jdff dff_B_BDBFFa2H9_2(.din(w_dff_B_OMidsCf33_2),.dout(w_dff_B_BDBFFa2H9_2),.clk(gclk));
	jdff dff_B_9wfcP7qg3_2(.din(w_dff_B_BDBFFa2H9_2),.dout(w_dff_B_9wfcP7qg3_2),.clk(gclk));
	jdff dff_B_9DcX31kt0_2(.din(w_dff_B_9wfcP7qg3_2),.dout(w_dff_B_9DcX31kt0_2),.clk(gclk));
	jdff dff_B_SrBj10tN2_2(.din(w_dff_B_9DcX31kt0_2),.dout(w_dff_B_SrBj10tN2_2),.clk(gclk));
	jdff dff_B_M25pG8lK2_2(.din(w_dff_B_SrBj10tN2_2),.dout(w_dff_B_M25pG8lK2_2),.clk(gclk));
	jdff dff_B_kHchIEaa6_2(.din(w_dff_B_M25pG8lK2_2),.dout(w_dff_B_kHchIEaa6_2),.clk(gclk));
	jdff dff_B_UnfEEObK3_2(.din(n1594),.dout(w_dff_B_UnfEEObK3_2),.clk(gclk));
	jdff dff_B_5Ib0KJ6z6_1(.din(n1592),.dout(w_dff_B_5Ib0KJ6z6_1),.clk(gclk));
	jdff dff_B_6mDeWR194_2(.din(n1527),.dout(w_dff_B_6mDeWR194_2),.clk(gclk));
	jdff dff_B_e6VEtXIN7_2(.din(w_dff_B_6mDeWR194_2),.dout(w_dff_B_e6VEtXIN7_2),.clk(gclk));
	jdff dff_B_UCsQuMDI3_2(.din(w_dff_B_e6VEtXIN7_2),.dout(w_dff_B_UCsQuMDI3_2),.clk(gclk));
	jdff dff_B_JRcnFvYy4_2(.din(w_dff_B_UCsQuMDI3_2),.dout(w_dff_B_JRcnFvYy4_2),.clk(gclk));
	jdff dff_B_MFX8Wkw83_2(.din(w_dff_B_JRcnFvYy4_2),.dout(w_dff_B_MFX8Wkw83_2),.clk(gclk));
	jdff dff_B_mzGL6Rjl6_2(.din(w_dff_B_MFX8Wkw83_2),.dout(w_dff_B_mzGL6Rjl6_2),.clk(gclk));
	jdff dff_B_WFH46CMZ3_2(.din(w_dff_B_mzGL6Rjl6_2),.dout(w_dff_B_WFH46CMZ3_2),.clk(gclk));
	jdff dff_B_ge74TO3H0_2(.din(w_dff_B_WFH46CMZ3_2),.dout(w_dff_B_ge74TO3H0_2),.clk(gclk));
	jdff dff_B_9nAkBgvF4_2(.din(w_dff_B_ge74TO3H0_2),.dout(w_dff_B_9nAkBgvF4_2),.clk(gclk));
	jdff dff_B_tEkRrEQx5_2(.din(w_dff_B_9nAkBgvF4_2),.dout(w_dff_B_tEkRrEQx5_2),.clk(gclk));
	jdff dff_B_eYeKBaxX4_2(.din(w_dff_B_tEkRrEQx5_2),.dout(w_dff_B_eYeKBaxX4_2),.clk(gclk));
	jdff dff_B_shl8RVuo8_2(.din(w_dff_B_eYeKBaxX4_2),.dout(w_dff_B_shl8RVuo8_2),.clk(gclk));
	jdff dff_B_vW9Omg9Y5_2(.din(w_dff_B_shl8RVuo8_2),.dout(w_dff_B_vW9Omg9Y5_2),.clk(gclk));
	jdff dff_B_mZFqtfPm4_2(.din(w_dff_B_vW9Omg9Y5_2),.dout(w_dff_B_mZFqtfPm4_2),.clk(gclk));
	jdff dff_B_khDeRDKf5_2(.din(w_dff_B_mZFqtfPm4_2),.dout(w_dff_B_khDeRDKf5_2),.clk(gclk));
	jdff dff_B_lLYUcJ0l3_2(.din(w_dff_B_khDeRDKf5_2),.dout(w_dff_B_lLYUcJ0l3_2),.clk(gclk));
	jdff dff_B_nDEpZeTr1_2(.din(w_dff_B_lLYUcJ0l3_2),.dout(w_dff_B_nDEpZeTr1_2),.clk(gclk));
	jdff dff_B_oRanvpB28_2(.din(w_dff_B_nDEpZeTr1_2),.dout(w_dff_B_oRanvpB28_2),.clk(gclk));
	jdff dff_B_Xg6cKKdn8_2(.din(w_dff_B_oRanvpB28_2),.dout(w_dff_B_Xg6cKKdn8_2),.clk(gclk));
	jdff dff_B_rUxF75Gh1_2(.din(w_dff_B_Xg6cKKdn8_2),.dout(w_dff_B_rUxF75Gh1_2),.clk(gclk));
	jdff dff_B_lATFeJ7o8_2(.din(w_dff_B_rUxF75Gh1_2),.dout(w_dff_B_lATFeJ7o8_2),.clk(gclk));
	jdff dff_B_n1s3b0gx8_2(.din(w_dff_B_lATFeJ7o8_2),.dout(w_dff_B_n1s3b0gx8_2),.clk(gclk));
	jdff dff_B_xyvqGlYi3_2(.din(w_dff_B_n1s3b0gx8_2),.dout(w_dff_B_xyvqGlYi3_2),.clk(gclk));
	jdff dff_B_ZViB0PM44_2(.din(w_dff_B_xyvqGlYi3_2),.dout(w_dff_B_ZViB0PM44_2),.clk(gclk));
	jdff dff_B_mzIA7bHb1_2(.din(w_dff_B_ZViB0PM44_2),.dout(w_dff_B_mzIA7bHb1_2),.clk(gclk));
	jdff dff_B_LMxFCVxi2_2(.din(w_dff_B_mzIA7bHb1_2),.dout(w_dff_B_LMxFCVxi2_2),.clk(gclk));
	jdff dff_B_lKy1rCvA4_2(.din(w_dff_B_LMxFCVxi2_2),.dout(w_dff_B_lKy1rCvA4_2),.clk(gclk));
	jdff dff_B_MA7Um7Op1_2(.din(w_dff_B_lKy1rCvA4_2),.dout(w_dff_B_MA7Um7Op1_2),.clk(gclk));
	jdff dff_B_onbLRaAG6_2(.din(w_dff_B_MA7Um7Op1_2),.dout(w_dff_B_onbLRaAG6_2),.clk(gclk));
	jdff dff_B_N7kavOKX5_2(.din(w_dff_B_onbLRaAG6_2),.dout(w_dff_B_N7kavOKX5_2),.clk(gclk));
	jdff dff_B_jdG9VyKO9_2(.din(w_dff_B_N7kavOKX5_2),.dout(w_dff_B_jdG9VyKO9_2),.clk(gclk));
	jdff dff_B_LSNcCxB14_1(.din(n1533),.dout(w_dff_B_LSNcCxB14_1),.clk(gclk));
	jdff dff_B_vQjzTvuR7_1(.din(w_dff_B_LSNcCxB14_1),.dout(w_dff_B_vQjzTvuR7_1),.clk(gclk));
	jdff dff_B_ibLykyi51_2(.din(n1532),.dout(w_dff_B_ibLykyi51_2),.clk(gclk));
	jdff dff_B_s9QbUPPy4_2(.din(w_dff_B_ibLykyi51_2),.dout(w_dff_B_s9QbUPPy4_2),.clk(gclk));
	jdff dff_B_JkBdRdHn1_2(.din(w_dff_B_s9QbUPPy4_2),.dout(w_dff_B_JkBdRdHn1_2),.clk(gclk));
	jdff dff_B_4Jorb95c9_2(.din(w_dff_B_JkBdRdHn1_2),.dout(w_dff_B_4Jorb95c9_2),.clk(gclk));
	jdff dff_B_1TCjGsp41_2(.din(w_dff_B_4Jorb95c9_2),.dout(w_dff_B_1TCjGsp41_2),.clk(gclk));
	jdff dff_B_mRbUQ3g31_2(.din(w_dff_B_1TCjGsp41_2),.dout(w_dff_B_mRbUQ3g31_2),.clk(gclk));
	jdff dff_B_azAAQTRp2_2(.din(w_dff_B_mRbUQ3g31_2),.dout(w_dff_B_azAAQTRp2_2),.clk(gclk));
	jdff dff_B_rzrCC7gD0_2(.din(w_dff_B_azAAQTRp2_2),.dout(w_dff_B_rzrCC7gD0_2),.clk(gclk));
	jdff dff_B_Ruytk1vZ0_2(.din(w_dff_B_rzrCC7gD0_2),.dout(w_dff_B_Ruytk1vZ0_2),.clk(gclk));
	jdff dff_B_XUH9uMB30_2(.din(w_dff_B_Ruytk1vZ0_2),.dout(w_dff_B_XUH9uMB30_2),.clk(gclk));
	jdff dff_B_MroiVKSx5_2(.din(w_dff_B_XUH9uMB30_2),.dout(w_dff_B_MroiVKSx5_2),.clk(gclk));
	jdff dff_B_Ta7dHKfX4_2(.din(w_dff_B_MroiVKSx5_2),.dout(w_dff_B_Ta7dHKfX4_2),.clk(gclk));
	jdff dff_B_pTwgOsb36_2(.din(w_dff_B_Ta7dHKfX4_2),.dout(w_dff_B_pTwgOsb36_2),.clk(gclk));
	jdff dff_B_DNcvXVLo1_2(.din(w_dff_B_pTwgOsb36_2),.dout(w_dff_B_DNcvXVLo1_2),.clk(gclk));
	jdff dff_B_EYpDFgBa6_2(.din(w_dff_B_DNcvXVLo1_2),.dout(w_dff_B_EYpDFgBa6_2),.clk(gclk));
	jdff dff_B_do05VpS64_2(.din(w_dff_B_EYpDFgBa6_2),.dout(w_dff_B_do05VpS64_2),.clk(gclk));
	jdff dff_B_VRyluxtt1_2(.din(w_dff_B_do05VpS64_2),.dout(w_dff_B_VRyluxtt1_2),.clk(gclk));
	jdff dff_B_TlAaYFG82_2(.din(w_dff_B_VRyluxtt1_2),.dout(w_dff_B_TlAaYFG82_2),.clk(gclk));
	jdff dff_B_Str4OJXp6_2(.din(w_dff_B_TlAaYFG82_2),.dout(w_dff_B_Str4OJXp6_2),.clk(gclk));
	jdff dff_B_JtTlxIsj9_2(.din(w_dff_B_Str4OJXp6_2),.dout(w_dff_B_JtTlxIsj9_2),.clk(gclk));
	jdff dff_B_Pp8lzc4Y1_2(.din(w_dff_B_JtTlxIsj9_2),.dout(w_dff_B_Pp8lzc4Y1_2),.clk(gclk));
	jdff dff_B_RVJo6Cox1_2(.din(w_dff_B_Pp8lzc4Y1_2),.dout(w_dff_B_RVJo6Cox1_2),.clk(gclk));
	jdff dff_B_O5zsZdx58_2(.din(w_dff_B_RVJo6Cox1_2),.dout(w_dff_B_O5zsZdx58_2),.clk(gclk));
	jdff dff_B_on58kIbA4_2(.din(w_dff_B_O5zsZdx58_2),.dout(w_dff_B_on58kIbA4_2),.clk(gclk));
	jdff dff_B_mdLUZads8_2(.din(w_dff_B_on58kIbA4_2),.dout(w_dff_B_mdLUZads8_2),.clk(gclk));
	jdff dff_B_Y63PJbbi7_2(.din(w_dff_B_mdLUZads8_2),.dout(w_dff_B_Y63PJbbi7_2),.clk(gclk));
	jdff dff_B_dwipn1rX2_2(.din(w_dff_B_Y63PJbbi7_2),.dout(w_dff_B_dwipn1rX2_2),.clk(gclk));
	jdff dff_B_GkoW1heP5_2(.din(w_dff_B_dwipn1rX2_2),.dout(w_dff_B_GkoW1heP5_2),.clk(gclk));
	jdff dff_B_3a0ws0L71_2(.din(n1531),.dout(w_dff_B_3a0ws0L71_2),.clk(gclk));
	jdff dff_B_6GyjjIVl4_2(.din(w_dff_B_3a0ws0L71_2),.dout(w_dff_B_6GyjjIVl4_2),.clk(gclk));
	jdff dff_B_IGZpL0219_2(.din(w_dff_B_6GyjjIVl4_2),.dout(w_dff_B_IGZpL0219_2),.clk(gclk));
	jdff dff_B_XEpzRJvB0_2(.din(w_dff_B_IGZpL0219_2),.dout(w_dff_B_XEpzRJvB0_2),.clk(gclk));
	jdff dff_B_6sXv0xHP5_2(.din(w_dff_B_XEpzRJvB0_2),.dout(w_dff_B_6sXv0xHP5_2),.clk(gclk));
	jdff dff_B_A9yybFE71_2(.din(w_dff_B_6sXv0xHP5_2),.dout(w_dff_B_A9yybFE71_2),.clk(gclk));
	jdff dff_B_8k5jswkw5_2(.din(w_dff_B_A9yybFE71_2),.dout(w_dff_B_8k5jswkw5_2),.clk(gclk));
	jdff dff_B_J8DRx8WX8_2(.din(w_dff_B_8k5jswkw5_2),.dout(w_dff_B_J8DRx8WX8_2),.clk(gclk));
	jdff dff_B_eyLxlTuN3_2(.din(w_dff_B_J8DRx8WX8_2),.dout(w_dff_B_eyLxlTuN3_2),.clk(gclk));
	jdff dff_B_IF5onHPo3_2(.din(w_dff_B_eyLxlTuN3_2),.dout(w_dff_B_IF5onHPo3_2),.clk(gclk));
	jdff dff_B_ULKHogEp3_2(.din(w_dff_B_IF5onHPo3_2),.dout(w_dff_B_ULKHogEp3_2),.clk(gclk));
	jdff dff_B_o5MC7lmz3_2(.din(w_dff_B_ULKHogEp3_2),.dout(w_dff_B_o5MC7lmz3_2),.clk(gclk));
	jdff dff_B_Egf9GCyA2_2(.din(w_dff_B_o5MC7lmz3_2),.dout(w_dff_B_Egf9GCyA2_2),.clk(gclk));
	jdff dff_B_Wp0eq3h40_2(.din(w_dff_B_Egf9GCyA2_2),.dout(w_dff_B_Wp0eq3h40_2),.clk(gclk));
	jdff dff_B_UTino0ZK6_2(.din(w_dff_B_Wp0eq3h40_2),.dout(w_dff_B_UTino0ZK6_2),.clk(gclk));
	jdff dff_B_xNTmY2ne4_2(.din(w_dff_B_UTino0ZK6_2),.dout(w_dff_B_xNTmY2ne4_2),.clk(gclk));
	jdff dff_B_mt0QN3742_2(.din(w_dff_B_xNTmY2ne4_2),.dout(w_dff_B_mt0QN3742_2),.clk(gclk));
	jdff dff_B_RU52QQuH0_2(.din(w_dff_B_mt0QN3742_2),.dout(w_dff_B_RU52QQuH0_2),.clk(gclk));
	jdff dff_B_6Ccp02qV8_2(.din(w_dff_B_RU52QQuH0_2),.dout(w_dff_B_6Ccp02qV8_2),.clk(gclk));
	jdff dff_B_zVrLvjrx1_2(.din(w_dff_B_6Ccp02qV8_2),.dout(w_dff_B_zVrLvjrx1_2),.clk(gclk));
	jdff dff_B_hPaFveAv8_2(.din(w_dff_B_zVrLvjrx1_2),.dout(w_dff_B_hPaFveAv8_2),.clk(gclk));
	jdff dff_B_lTKs7F450_2(.din(w_dff_B_hPaFveAv8_2),.dout(w_dff_B_lTKs7F450_2),.clk(gclk));
	jdff dff_B_4fYwJyMx9_2(.din(w_dff_B_lTKs7F450_2),.dout(w_dff_B_4fYwJyMx9_2),.clk(gclk));
	jdff dff_B_cVcvy8Hg7_2(.din(w_dff_B_4fYwJyMx9_2),.dout(w_dff_B_cVcvy8Hg7_2),.clk(gclk));
	jdff dff_B_KIGlNau69_2(.din(w_dff_B_cVcvy8Hg7_2),.dout(w_dff_B_KIGlNau69_2),.clk(gclk));
	jdff dff_B_1PfSOphx1_2(.din(w_dff_B_KIGlNau69_2),.dout(w_dff_B_1PfSOphx1_2),.clk(gclk));
	jdff dff_B_g8nA3w162_2(.din(w_dff_B_1PfSOphx1_2),.dout(w_dff_B_g8nA3w162_2),.clk(gclk));
	jdff dff_B_QT5HnJV77_2(.din(w_dff_B_g8nA3w162_2),.dout(w_dff_B_QT5HnJV77_2),.clk(gclk));
	jdff dff_B_ounjcS661_2(.din(w_dff_B_QT5HnJV77_2),.dout(w_dff_B_ounjcS661_2),.clk(gclk));
	jdff dff_B_irSCcU5R7_2(.din(w_dff_B_ounjcS661_2),.dout(w_dff_B_irSCcU5R7_2),.clk(gclk));
	jdff dff_B_24k6eYsp4_2(.din(n1530),.dout(w_dff_B_24k6eYsp4_2),.clk(gclk));
	jdff dff_B_eVn4YkX40_1(.din(n1528),.dout(w_dff_B_eVn4YkX40_1),.clk(gclk));
	jdff dff_B_bcA32Be96_2(.din(n1456),.dout(w_dff_B_bcA32Be96_2),.clk(gclk));
	jdff dff_B_12jGT5iy4_2(.din(w_dff_B_bcA32Be96_2),.dout(w_dff_B_12jGT5iy4_2),.clk(gclk));
	jdff dff_B_mXjMtn4r1_2(.din(w_dff_B_12jGT5iy4_2),.dout(w_dff_B_mXjMtn4r1_2),.clk(gclk));
	jdff dff_B_zEStQkLn0_2(.din(w_dff_B_mXjMtn4r1_2),.dout(w_dff_B_zEStQkLn0_2),.clk(gclk));
	jdff dff_B_Oju0jybA7_2(.din(w_dff_B_zEStQkLn0_2),.dout(w_dff_B_Oju0jybA7_2),.clk(gclk));
	jdff dff_B_kZEymnYy2_2(.din(w_dff_B_Oju0jybA7_2),.dout(w_dff_B_kZEymnYy2_2),.clk(gclk));
	jdff dff_B_9Kv2D6ss0_2(.din(w_dff_B_kZEymnYy2_2),.dout(w_dff_B_9Kv2D6ss0_2),.clk(gclk));
	jdff dff_B_To2LDRTW2_2(.din(w_dff_B_9Kv2D6ss0_2),.dout(w_dff_B_To2LDRTW2_2),.clk(gclk));
	jdff dff_B_DRh7zhKd8_2(.din(w_dff_B_To2LDRTW2_2),.dout(w_dff_B_DRh7zhKd8_2),.clk(gclk));
	jdff dff_B_ZrLYkahn4_2(.din(w_dff_B_DRh7zhKd8_2),.dout(w_dff_B_ZrLYkahn4_2),.clk(gclk));
	jdff dff_B_7om8xK6W1_2(.din(w_dff_B_ZrLYkahn4_2),.dout(w_dff_B_7om8xK6W1_2),.clk(gclk));
	jdff dff_B_juQnec570_2(.din(w_dff_B_7om8xK6W1_2),.dout(w_dff_B_juQnec570_2),.clk(gclk));
	jdff dff_B_llXl76rH8_2(.din(w_dff_B_juQnec570_2),.dout(w_dff_B_llXl76rH8_2),.clk(gclk));
	jdff dff_B_nczVXYaZ6_2(.din(w_dff_B_llXl76rH8_2),.dout(w_dff_B_nczVXYaZ6_2),.clk(gclk));
	jdff dff_B_CgQ9lM237_2(.din(w_dff_B_nczVXYaZ6_2),.dout(w_dff_B_CgQ9lM237_2),.clk(gclk));
	jdff dff_B_H4rYk0z34_2(.din(w_dff_B_CgQ9lM237_2),.dout(w_dff_B_H4rYk0z34_2),.clk(gclk));
	jdff dff_B_MtpIjnst4_2(.din(w_dff_B_H4rYk0z34_2),.dout(w_dff_B_MtpIjnst4_2),.clk(gclk));
	jdff dff_B_d2bQqD3o7_2(.din(w_dff_B_MtpIjnst4_2),.dout(w_dff_B_d2bQqD3o7_2),.clk(gclk));
	jdff dff_B_c0lx2f367_2(.din(w_dff_B_d2bQqD3o7_2),.dout(w_dff_B_c0lx2f367_2),.clk(gclk));
	jdff dff_B_VnXblzEc8_2(.din(w_dff_B_c0lx2f367_2),.dout(w_dff_B_VnXblzEc8_2),.clk(gclk));
	jdff dff_B_acjOKS6m0_2(.din(w_dff_B_VnXblzEc8_2),.dout(w_dff_B_acjOKS6m0_2),.clk(gclk));
	jdff dff_B_OKCdYD7p1_2(.din(w_dff_B_acjOKS6m0_2),.dout(w_dff_B_OKCdYD7p1_2),.clk(gclk));
	jdff dff_B_6pmO231M2_2(.din(w_dff_B_OKCdYD7p1_2),.dout(w_dff_B_6pmO231M2_2),.clk(gclk));
	jdff dff_B_11lJgs1H3_2(.din(w_dff_B_6pmO231M2_2),.dout(w_dff_B_11lJgs1H3_2),.clk(gclk));
	jdff dff_B_7htPfhn37_2(.din(w_dff_B_11lJgs1H3_2),.dout(w_dff_B_7htPfhn37_2),.clk(gclk));
	jdff dff_B_MEA4sZFM7_2(.din(w_dff_B_7htPfhn37_2),.dout(w_dff_B_MEA4sZFM7_2),.clk(gclk));
	jdff dff_B_cqr3P2Ay4_2(.din(w_dff_B_MEA4sZFM7_2),.dout(w_dff_B_cqr3P2Ay4_2),.clk(gclk));
	jdff dff_B_mGTa7ymT7_1(.din(n1462),.dout(w_dff_B_mGTa7ymT7_1),.clk(gclk));
	jdff dff_B_meQsglwa0_1(.din(w_dff_B_mGTa7ymT7_1),.dout(w_dff_B_meQsglwa0_1),.clk(gclk));
	jdff dff_B_WyQdZu1G7_2(.din(n1461),.dout(w_dff_B_WyQdZu1G7_2),.clk(gclk));
	jdff dff_B_oBi0Ul3v7_2(.din(w_dff_B_WyQdZu1G7_2),.dout(w_dff_B_oBi0Ul3v7_2),.clk(gclk));
	jdff dff_B_10I6NcpG1_2(.din(w_dff_B_oBi0Ul3v7_2),.dout(w_dff_B_10I6NcpG1_2),.clk(gclk));
	jdff dff_B_dAoGwnK16_2(.din(w_dff_B_10I6NcpG1_2),.dout(w_dff_B_dAoGwnK16_2),.clk(gclk));
	jdff dff_B_llaNNY9k5_2(.din(w_dff_B_dAoGwnK16_2),.dout(w_dff_B_llaNNY9k5_2),.clk(gclk));
	jdff dff_B_0yrPQEYH1_2(.din(w_dff_B_llaNNY9k5_2),.dout(w_dff_B_0yrPQEYH1_2),.clk(gclk));
	jdff dff_B_S8UkZmQP4_2(.din(w_dff_B_0yrPQEYH1_2),.dout(w_dff_B_S8UkZmQP4_2),.clk(gclk));
	jdff dff_B_yCnypHLG3_2(.din(w_dff_B_S8UkZmQP4_2),.dout(w_dff_B_yCnypHLG3_2),.clk(gclk));
	jdff dff_B_zAvpxqvI1_2(.din(w_dff_B_yCnypHLG3_2),.dout(w_dff_B_zAvpxqvI1_2),.clk(gclk));
	jdff dff_B_q98XcGyK4_2(.din(w_dff_B_zAvpxqvI1_2),.dout(w_dff_B_q98XcGyK4_2),.clk(gclk));
	jdff dff_B_swfoPuTx3_2(.din(w_dff_B_q98XcGyK4_2),.dout(w_dff_B_swfoPuTx3_2),.clk(gclk));
	jdff dff_B_eAFofZcY0_2(.din(w_dff_B_swfoPuTx3_2),.dout(w_dff_B_eAFofZcY0_2),.clk(gclk));
	jdff dff_B_n1LLCpb47_2(.din(w_dff_B_eAFofZcY0_2),.dout(w_dff_B_n1LLCpb47_2),.clk(gclk));
	jdff dff_B_swi9ghk14_2(.din(w_dff_B_n1LLCpb47_2),.dout(w_dff_B_swi9ghk14_2),.clk(gclk));
	jdff dff_B_Rs0wV5UK9_2(.din(w_dff_B_swi9ghk14_2),.dout(w_dff_B_Rs0wV5UK9_2),.clk(gclk));
	jdff dff_B_99iUJNDd3_2(.din(w_dff_B_Rs0wV5UK9_2),.dout(w_dff_B_99iUJNDd3_2),.clk(gclk));
	jdff dff_B_3fH8X0Og1_2(.din(w_dff_B_99iUJNDd3_2),.dout(w_dff_B_3fH8X0Og1_2),.clk(gclk));
	jdff dff_B_I6TdlgN36_2(.din(w_dff_B_3fH8X0Og1_2),.dout(w_dff_B_I6TdlgN36_2),.clk(gclk));
	jdff dff_B_hmCv5Pzt1_2(.din(w_dff_B_I6TdlgN36_2),.dout(w_dff_B_hmCv5Pzt1_2),.clk(gclk));
	jdff dff_B_Dq9MvurV8_2(.din(w_dff_B_hmCv5Pzt1_2),.dout(w_dff_B_Dq9MvurV8_2),.clk(gclk));
	jdff dff_B_3xe1moFK4_2(.din(w_dff_B_Dq9MvurV8_2),.dout(w_dff_B_3xe1moFK4_2),.clk(gclk));
	jdff dff_B_zKPuNROK4_2(.din(w_dff_B_3xe1moFK4_2),.dout(w_dff_B_zKPuNROK4_2),.clk(gclk));
	jdff dff_B_OQdcmkcf5_2(.din(w_dff_B_zKPuNROK4_2),.dout(w_dff_B_OQdcmkcf5_2),.clk(gclk));
	jdff dff_B_x0NmA8Gt4_2(.din(w_dff_B_OQdcmkcf5_2),.dout(w_dff_B_x0NmA8Gt4_2),.clk(gclk));
	jdff dff_B_1yjvzkdL5_2(.din(n1460),.dout(w_dff_B_1yjvzkdL5_2),.clk(gclk));
	jdff dff_B_Ijjsn1bS6_2(.din(w_dff_B_1yjvzkdL5_2),.dout(w_dff_B_Ijjsn1bS6_2),.clk(gclk));
	jdff dff_B_p0bRLz0k3_2(.din(w_dff_B_Ijjsn1bS6_2),.dout(w_dff_B_p0bRLz0k3_2),.clk(gclk));
	jdff dff_B_wrgEB7nz3_2(.din(w_dff_B_p0bRLz0k3_2),.dout(w_dff_B_wrgEB7nz3_2),.clk(gclk));
	jdff dff_B_8VbBVnmX6_2(.din(w_dff_B_wrgEB7nz3_2),.dout(w_dff_B_8VbBVnmX6_2),.clk(gclk));
	jdff dff_B_6kBtE20E3_2(.din(w_dff_B_8VbBVnmX6_2),.dout(w_dff_B_6kBtE20E3_2),.clk(gclk));
	jdff dff_B_CW53KMFZ8_2(.din(w_dff_B_6kBtE20E3_2),.dout(w_dff_B_CW53KMFZ8_2),.clk(gclk));
	jdff dff_B_UsQPoqyH9_2(.din(w_dff_B_CW53KMFZ8_2),.dout(w_dff_B_UsQPoqyH9_2),.clk(gclk));
	jdff dff_B_XO43nQfU9_2(.din(w_dff_B_UsQPoqyH9_2),.dout(w_dff_B_XO43nQfU9_2),.clk(gclk));
	jdff dff_B_Y4MTR1hm7_2(.din(w_dff_B_XO43nQfU9_2),.dout(w_dff_B_Y4MTR1hm7_2),.clk(gclk));
	jdff dff_B_nu9ZHmxk8_2(.din(w_dff_B_Y4MTR1hm7_2),.dout(w_dff_B_nu9ZHmxk8_2),.clk(gclk));
	jdff dff_B_Xg0YCQo83_2(.din(w_dff_B_nu9ZHmxk8_2),.dout(w_dff_B_Xg0YCQo83_2),.clk(gclk));
	jdff dff_B_JFMTEVnT9_2(.din(w_dff_B_Xg0YCQo83_2),.dout(w_dff_B_JFMTEVnT9_2),.clk(gclk));
	jdff dff_B_MZkzplGT3_2(.din(w_dff_B_JFMTEVnT9_2),.dout(w_dff_B_MZkzplGT3_2),.clk(gclk));
	jdff dff_B_tMWkEoQz2_2(.din(w_dff_B_MZkzplGT3_2),.dout(w_dff_B_tMWkEoQz2_2),.clk(gclk));
	jdff dff_B_JOlqMAD76_2(.din(w_dff_B_tMWkEoQz2_2),.dout(w_dff_B_JOlqMAD76_2),.clk(gclk));
	jdff dff_B_TW2E4hbb8_2(.din(w_dff_B_JOlqMAD76_2),.dout(w_dff_B_TW2E4hbb8_2),.clk(gclk));
	jdff dff_B_7r5Qeh8O9_2(.din(w_dff_B_TW2E4hbb8_2),.dout(w_dff_B_7r5Qeh8O9_2),.clk(gclk));
	jdff dff_B_ZXZrfq8x5_2(.din(w_dff_B_7r5Qeh8O9_2),.dout(w_dff_B_ZXZrfq8x5_2),.clk(gclk));
	jdff dff_B_f18JwbVl1_2(.din(w_dff_B_ZXZrfq8x5_2),.dout(w_dff_B_f18JwbVl1_2),.clk(gclk));
	jdff dff_B_XNgtLl0o0_2(.din(w_dff_B_f18JwbVl1_2),.dout(w_dff_B_XNgtLl0o0_2),.clk(gclk));
	jdff dff_B_erCkOw5d8_2(.din(w_dff_B_XNgtLl0o0_2),.dout(w_dff_B_erCkOw5d8_2),.clk(gclk));
	jdff dff_B_VVeSMAgY2_2(.din(w_dff_B_erCkOw5d8_2),.dout(w_dff_B_VVeSMAgY2_2),.clk(gclk));
	jdff dff_B_0XNddVoS8_2(.din(w_dff_B_VVeSMAgY2_2),.dout(w_dff_B_0XNddVoS8_2),.clk(gclk));
	jdff dff_B_6N6dtyd68_2(.din(w_dff_B_0XNddVoS8_2),.dout(w_dff_B_6N6dtyd68_2),.clk(gclk));
	jdff dff_B_zZeO24ZO9_2(.din(w_dff_B_6N6dtyd68_2),.dout(w_dff_B_zZeO24ZO9_2),.clk(gclk));
	jdff dff_B_mAl5mvvM9_2(.din(n1459),.dout(w_dff_B_mAl5mvvM9_2),.clk(gclk));
	jdff dff_B_MiHFayT22_1(.din(n1457),.dout(w_dff_B_MiHFayT22_1),.clk(gclk));
	jdff dff_B_6zRCsN5I2_2(.din(n1378),.dout(w_dff_B_6zRCsN5I2_2),.clk(gclk));
	jdff dff_B_hmc8dgcw6_2(.din(w_dff_B_6zRCsN5I2_2),.dout(w_dff_B_hmc8dgcw6_2),.clk(gclk));
	jdff dff_B_siPT53r59_2(.din(w_dff_B_hmc8dgcw6_2),.dout(w_dff_B_siPT53r59_2),.clk(gclk));
	jdff dff_B_M5VmMrFx9_2(.din(w_dff_B_siPT53r59_2),.dout(w_dff_B_M5VmMrFx9_2),.clk(gclk));
	jdff dff_B_MSfkfmxL6_2(.din(w_dff_B_M5VmMrFx9_2),.dout(w_dff_B_MSfkfmxL6_2),.clk(gclk));
	jdff dff_B_AqV1lGGE3_2(.din(w_dff_B_MSfkfmxL6_2),.dout(w_dff_B_AqV1lGGE3_2),.clk(gclk));
	jdff dff_B_IwUBOxKk4_2(.din(w_dff_B_AqV1lGGE3_2),.dout(w_dff_B_IwUBOxKk4_2),.clk(gclk));
	jdff dff_B_QxY2O6uL2_2(.din(w_dff_B_IwUBOxKk4_2),.dout(w_dff_B_QxY2O6uL2_2),.clk(gclk));
	jdff dff_B_pnjtYi0U3_2(.din(w_dff_B_QxY2O6uL2_2),.dout(w_dff_B_pnjtYi0U3_2),.clk(gclk));
	jdff dff_B_GQwWV3tM8_2(.din(w_dff_B_pnjtYi0U3_2),.dout(w_dff_B_GQwWV3tM8_2),.clk(gclk));
	jdff dff_B_2FJrH1991_2(.din(w_dff_B_GQwWV3tM8_2),.dout(w_dff_B_2FJrH1991_2),.clk(gclk));
	jdff dff_B_53qjY3DZ7_2(.din(w_dff_B_2FJrH1991_2),.dout(w_dff_B_53qjY3DZ7_2),.clk(gclk));
	jdff dff_B_tWS8GqNM7_2(.din(w_dff_B_53qjY3DZ7_2),.dout(w_dff_B_tWS8GqNM7_2),.clk(gclk));
	jdff dff_B_Ncememkz1_2(.din(w_dff_B_tWS8GqNM7_2),.dout(w_dff_B_Ncememkz1_2),.clk(gclk));
	jdff dff_B_H27Ncgy10_2(.din(w_dff_B_Ncememkz1_2),.dout(w_dff_B_H27Ncgy10_2),.clk(gclk));
	jdff dff_B_Zu0aLVpB7_2(.din(w_dff_B_H27Ncgy10_2),.dout(w_dff_B_Zu0aLVpB7_2),.clk(gclk));
	jdff dff_B_cBJZNKeD1_2(.din(w_dff_B_Zu0aLVpB7_2),.dout(w_dff_B_cBJZNKeD1_2),.clk(gclk));
	jdff dff_B_R0xnnk9L3_2(.din(w_dff_B_cBJZNKeD1_2),.dout(w_dff_B_R0xnnk9L3_2),.clk(gclk));
	jdff dff_B_QYyFxlef0_2(.din(w_dff_B_R0xnnk9L3_2),.dout(w_dff_B_QYyFxlef0_2),.clk(gclk));
	jdff dff_B_AFaUlWWF0_2(.din(w_dff_B_QYyFxlef0_2),.dout(w_dff_B_AFaUlWWF0_2),.clk(gclk));
	jdff dff_B_NeAUwhoJ1_2(.din(w_dff_B_AFaUlWWF0_2),.dout(w_dff_B_NeAUwhoJ1_2),.clk(gclk));
	jdff dff_B_YBQHYPJ85_2(.din(w_dff_B_NeAUwhoJ1_2),.dout(w_dff_B_YBQHYPJ85_2),.clk(gclk));
	jdff dff_B_N0Tsv9Tp0_2(.din(w_dff_B_YBQHYPJ85_2),.dout(w_dff_B_N0Tsv9Tp0_2),.clk(gclk));
	jdff dff_B_5LwBCvTA9_1(.din(n1384),.dout(w_dff_B_5LwBCvTA9_1),.clk(gclk));
	jdff dff_B_2UYJmSWs0_1(.din(w_dff_B_5LwBCvTA9_1),.dout(w_dff_B_2UYJmSWs0_1),.clk(gclk));
	jdff dff_B_yBjCL9c09_2(.din(n1383),.dout(w_dff_B_yBjCL9c09_2),.clk(gclk));
	jdff dff_B_WiLuKK9K3_2(.din(w_dff_B_yBjCL9c09_2),.dout(w_dff_B_WiLuKK9K3_2),.clk(gclk));
	jdff dff_B_QAyQGM3A2_2(.din(w_dff_B_WiLuKK9K3_2),.dout(w_dff_B_QAyQGM3A2_2),.clk(gclk));
	jdff dff_B_wqT00hx83_2(.din(w_dff_B_QAyQGM3A2_2),.dout(w_dff_B_wqT00hx83_2),.clk(gclk));
	jdff dff_B_fBfICTYq0_2(.din(w_dff_B_wqT00hx83_2),.dout(w_dff_B_fBfICTYq0_2),.clk(gclk));
	jdff dff_B_6HAJBTrF0_2(.din(w_dff_B_fBfICTYq0_2),.dout(w_dff_B_6HAJBTrF0_2),.clk(gclk));
	jdff dff_B_FBM7TZ6n2_2(.din(w_dff_B_6HAJBTrF0_2),.dout(w_dff_B_FBM7TZ6n2_2),.clk(gclk));
	jdff dff_B_3kmW9Kiy3_2(.din(w_dff_B_FBM7TZ6n2_2),.dout(w_dff_B_3kmW9Kiy3_2),.clk(gclk));
	jdff dff_B_4ikPSIaQ3_2(.din(w_dff_B_3kmW9Kiy3_2),.dout(w_dff_B_4ikPSIaQ3_2),.clk(gclk));
	jdff dff_B_udyCn42C1_2(.din(w_dff_B_4ikPSIaQ3_2),.dout(w_dff_B_udyCn42C1_2),.clk(gclk));
	jdff dff_B_ocRjkFt70_2(.din(w_dff_B_udyCn42C1_2),.dout(w_dff_B_ocRjkFt70_2),.clk(gclk));
	jdff dff_B_bPEcba2J5_2(.din(w_dff_B_ocRjkFt70_2),.dout(w_dff_B_bPEcba2J5_2),.clk(gclk));
	jdff dff_B_CTYdPjno3_2(.din(w_dff_B_bPEcba2J5_2),.dout(w_dff_B_CTYdPjno3_2),.clk(gclk));
	jdff dff_B_tMLHx8p98_2(.din(w_dff_B_CTYdPjno3_2),.dout(w_dff_B_tMLHx8p98_2),.clk(gclk));
	jdff dff_B_A0wU6i6D4_2(.din(w_dff_B_tMLHx8p98_2),.dout(w_dff_B_A0wU6i6D4_2),.clk(gclk));
	jdff dff_B_mHjUDGzn5_2(.din(w_dff_B_A0wU6i6D4_2),.dout(w_dff_B_mHjUDGzn5_2),.clk(gclk));
	jdff dff_B_1nUWKe6m7_2(.din(w_dff_B_mHjUDGzn5_2),.dout(w_dff_B_1nUWKe6m7_2),.clk(gclk));
	jdff dff_B_6Li8uaB89_2(.din(w_dff_B_1nUWKe6m7_2),.dout(w_dff_B_6Li8uaB89_2),.clk(gclk));
	jdff dff_B_AGZPkQLo8_2(.din(w_dff_B_6Li8uaB89_2),.dout(w_dff_B_AGZPkQLo8_2),.clk(gclk));
	jdff dff_B_Lwcvv2XE9_2(.din(w_dff_B_AGZPkQLo8_2),.dout(w_dff_B_Lwcvv2XE9_2),.clk(gclk));
	jdff dff_B_Y5Gh3Yym8_2(.din(n1382),.dout(w_dff_B_Y5Gh3Yym8_2),.clk(gclk));
	jdff dff_B_zXbVV5OP3_2(.din(w_dff_B_Y5Gh3Yym8_2),.dout(w_dff_B_zXbVV5OP3_2),.clk(gclk));
	jdff dff_B_ls6NnuRX6_2(.din(w_dff_B_zXbVV5OP3_2),.dout(w_dff_B_ls6NnuRX6_2),.clk(gclk));
	jdff dff_B_wVoB6uRS9_2(.din(w_dff_B_ls6NnuRX6_2),.dout(w_dff_B_wVoB6uRS9_2),.clk(gclk));
	jdff dff_B_iirIfLG89_2(.din(w_dff_B_wVoB6uRS9_2),.dout(w_dff_B_iirIfLG89_2),.clk(gclk));
	jdff dff_B_IXb9wSKN3_2(.din(w_dff_B_iirIfLG89_2),.dout(w_dff_B_IXb9wSKN3_2),.clk(gclk));
	jdff dff_B_Igk4Mib62_2(.din(w_dff_B_IXb9wSKN3_2),.dout(w_dff_B_Igk4Mib62_2),.clk(gclk));
	jdff dff_B_ZjaErCCv8_2(.din(w_dff_B_Igk4Mib62_2),.dout(w_dff_B_ZjaErCCv8_2),.clk(gclk));
	jdff dff_B_bcPIvtUJ4_2(.din(w_dff_B_ZjaErCCv8_2),.dout(w_dff_B_bcPIvtUJ4_2),.clk(gclk));
	jdff dff_B_hvdYaCEX5_2(.din(w_dff_B_bcPIvtUJ4_2),.dout(w_dff_B_hvdYaCEX5_2),.clk(gclk));
	jdff dff_B_gW63nihM1_2(.din(w_dff_B_hvdYaCEX5_2),.dout(w_dff_B_gW63nihM1_2),.clk(gclk));
	jdff dff_B_fpEvUovD7_2(.din(w_dff_B_gW63nihM1_2),.dout(w_dff_B_fpEvUovD7_2),.clk(gclk));
	jdff dff_B_SksLlSMZ9_2(.din(w_dff_B_fpEvUovD7_2),.dout(w_dff_B_SksLlSMZ9_2),.clk(gclk));
	jdff dff_B_SSuJn0qK5_2(.din(w_dff_B_SksLlSMZ9_2),.dout(w_dff_B_SSuJn0qK5_2),.clk(gclk));
	jdff dff_B_aV4EAW3S3_2(.din(w_dff_B_SSuJn0qK5_2),.dout(w_dff_B_aV4EAW3S3_2),.clk(gclk));
	jdff dff_B_uM4aMKp82_2(.din(w_dff_B_aV4EAW3S3_2),.dout(w_dff_B_uM4aMKp82_2),.clk(gclk));
	jdff dff_B_hAc2qsIN2_2(.din(w_dff_B_uM4aMKp82_2),.dout(w_dff_B_hAc2qsIN2_2),.clk(gclk));
	jdff dff_B_Hy3qaCsF0_2(.din(w_dff_B_hAc2qsIN2_2),.dout(w_dff_B_Hy3qaCsF0_2),.clk(gclk));
	jdff dff_B_IEPpiw0e2_2(.din(w_dff_B_Hy3qaCsF0_2),.dout(w_dff_B_IEPpiw0e2_2),.clk(gclk));
	jdff dff_B_CMeRreZc7_2(.din(w_dff_B_IEPpiw0e2_2),.dout(w_dff_B_CMeRreZc7_2),.clk(gclk));
	jdff dff_B_H42GKPi99_2(.din(w_dff_B_CMeRreZc7_2),.dout(w_dff_B_H42GKPi99_2),.clk(gclk));
	jdff dff_B_lQleofwo6_2(.din(w_dff_B_H42GKPi99_2),.dout(w_dff_B_lQleofwo6_2),.clk(gclk));
	jdff dff_B_mB60qQA78_2(.din(n1381),.dout(w_dff_B_mB60qQA78_2),.clk(gclk));
	jdff dff_B_7k9iJ5tT6_1(.din(n1379),.dout(w_dff_B_7k9iJ5tT6_1),.clk(gclk));
	jdff dff_B_SK7ixJDL3_2(.din(n1293),.dout(w_dff_B_SK7ixJDL3_2),.clk(gclk));
	jdff dff_B_sR0uFpe75_2(.din(w_dff_B_SK7ixJDL3_2),.dout(w_dff_B_sR0uFpe75_2),.clk(gclk));
	jdff dff_B_WGOTq29G5_2(.din(w_dff_B_sR0uFpe75_2),.dout(w_dff_B_WGOTq29G5_2),.clk(gclk));
	jdff dff_B_iDHRGbm33_2(.din(w_dff_B_WGOTq29G5_2),.dout(w_dff_B_iDHRGbm33_2),.clk(gclk));
	jdff dff_B_c6Mhr2Ba4_2(.din(w_dff_B_iDHRGbm33_2),.dout(w_dff_B_c6Mhr2Ba4_2),.clk(gclk));
	jdff dff_B_zAsTsVJR7_2(.din(w_dff_B_c6Mhr2Ba4_2),.dout(w_dff_B_zAsTsVJR7_2),.clk(gclk));
	jdff dff_B_rp6kxHkv3_2(.din(w_dff_B_zAsTsVJR7_2),.dout(w_dff_B_rp6kxHkv3_2),.clk(gclk));
	jdff dff_B_mzWakkxk3_2(.din(w_dff_B_rp6kxHkv3_2),.dout(w_dff_B_mzWakkxk3_2),.clk(gclk));
	jdff dff_B_azXYWqpz2_2(.din(w_dff_B_mzWakkxk3_2),.dout(w_dff_B_azXYWqpz2_2),.clk(gclk));
	jdff dff_B_nb8owcxN6_2(.din(w_dff_B_azXYWqpz2_2),.dout(w_dff_B_nb8owcxN6_2),.clk(gclk));
	jdff dff_B_PHbfqBnV0_2(.din(w_dff_B_nb8owcxN6_2),.dout(w_dff_B_PHbfqBnV0_2),.clk(gclk));
	jdff dff_B_Cn08fwCC5_2(.din(w_dff_B_PHbfqBnV0_2),.dout(w_dff_B_Cn08fwCC5_2),.clk(gclk));
	jdff dff_B_IiyBCTar5_2(.din(w_dff_B_Cn08fwCC5_2),.dout(w_dff_B_IiyBCTar5_2),.clk(gclk));
	jdff dff_B_ne1Iznhr2_2(.din(w_dff_B_IiyBCTar5_2),.dout(w_dff_B_ne1Iznhr2_2),.clk(gclk));
	jdff dff_B_BFgKVyXo3_2(.din(w_dff_B_ne1Iznhr2_2),.dout(w_dff_B_BFgKVyXo3_2),.clk(gclk));
	jdff dff_B_U0JDzBCI0_2(.din(w_dff_B_BFgKVyXo3_2),.dout(w_dff_B_U0JDzBCI0_2),.clk(gclk));
	jdff dff_B_HPMWVqFw8_2(.din(w_dff_B_U0JDzBCI0_2),.dout(w_dff_B_HPMWVqFw8_2),.clk(gclk));
	jdff dff_B_gZGtd2Gi4_2(.din(w_dff_B_HPMWVqFw8_2),.dout(w_dff_B_gZGtd2Gi4_2),.clk(gclk));
	jdff dff_B_rOjuu2xq3_2(.din(w_dff_B_gZGtd2Gi4_2),.dout(w_dff_B_rOjuu2xq3_2),.clk(gclk));
	jdff dff_B_YPFpbhph5_1(.din(n1299),.dout(w_dff_B_YPFpbhph5_1),.clk(gclk));
	jdff dff_B_DCPQC2Kw1_1(.din(w_dff_B_YPFpbhph5_1),.dout(w_dff_B_DCPQC2Kw1_1),.clk(gclk));
	jdff dff_B_WEHEShuh7_2(.din(n1298),.dout(w_dff_B_WEHEShuh7_2),.clk(gclk));
	jdff dff_B_t7WOkIAn1_2(.din(w_dff_B_WEHEShuh7_2),.dout(w_dff_B_t7WOkIAn1_2),.clk(gclk));
	jdff dff_B_TBKjdZve0_2(.din(w_dff_B_t7WOkIAn1_2),.dout(w_dff_B_TBKjdZve0_2),.clk(gclk));
	jdff dff_B_mZJxy1Tw7_2(.din(w_dff_B_TBKjdZve0_2),.dout(w_dff_B_mZJxy1Tw7_2),.clk(gclk));
	jdff dff_B_7GGeUX2V7_2(.din(w_dff_B_mZJxy1Tw7_2),.dout(w_dff_B_7GGeUX2V7_2),.clk(gclk));
	jdff dff_B_itFfMoP16_2(.din(w_dff_B_7GGeUX2V7_2),.dout(w_dff_B_itFfMoP16_2),.clk(gclk));
	jdff dff_B_N6cZe30a7_2(.din(w_dff_B_itFfMoP16_2),.dout(w_dff_B_N6cZe30a7_2),.clk(gclk));
	jdff dff_B_8RBPbisT3_2(.din(w_dff_B_N6cZe30a7_2),.dout(w_dff_B_8RBPbisT3_2),.clk(gclk));
	jdff dff_B_tqzRjAZo4_2(.din(w_dff_B_8RBPbisT3_2),.dout(w_dff_B_tqzRjAZo4_2),.clk(gclk));
	jdff dff_B_0h8o1GjY6_2(.din(w_dff_B_tqzRjAZo4_2),.dout(w_dff_B_0h8o1GjY6_2),.clk(gclk));
	jdff dff_B_puAnTaMN9_2(.din(w_dff_B_0h8o1GjY6_2),.dout(w_dff_B_puAnTaMN9_2),.clk(gclk));
	jdff dff_B_nJi0isK64_2(.din(w_dff_B_puAnTaMN9_2),.dout(w_dff_B_nJi0isK64_2),.clk(gclk));
	jdff dff_B_iMRQ4lTU9_2(.din(w_dff_B_nJi0isK64_2),.dout(w_dff_B_iMRQ4lTU9_2),.clk(gclk));
	jdff dff_B_gM7jwQeG7_2(.din(w_dff_B_iMRQ4lTU9_2),.dout(w_dff_B_gM7jwQeG7_2),.clk(gclk));
	jdff dff_B_eIEwx81R7_2(.din(w_dff_B_gM7jwQeG7_2),.dout(w_dff_B_eIEwx81R7_2),.clk(gclk));
	jdff dff_B_WTdmoGjV0_2(.din(w_dff_B_eIEwx81R7_2),.dout(w_dff_B_WTdmoGjV0_2),.clk(gclk));
	jdff dff_B_Hhmpk3g62_2(.din(n1297),.dout(w_dff_B_Hhmpk3g62_2),.clk(gclk));
	jdff dff_B_AKrMBL1h4_2(.din(w_dff_B_Hhmpk3g62_2),.dout(w_dff_B_AKrMBL1h4_2),.clk(gclk));
	jdff dff_B_fBgfm8bz8_2(.din(w_dff_B_AKrMBL1h4_2),.dout(w_dff_B_fBgfm8bz8_2),.clk(gclk));
	jdff dff_B_AdgTnOUt5_2(.din(w_dff_B_fBgfm8bz8_2),.dout(w_dff_B_AdgTnOUt5_2),.clk(gclk));
	jdff dff_B_dFoGbecY3_2(.din(w_dff_B_AdgTnOUt5_2),.dout(w_dff_B_dFoGbecY3_2),.clk(gclk));
	jdff dff_B_qX1pOQzH7_2(.din(w_dff_B_dFoGbecY3_2),.dout(w_dff_B_qX1pOQzH7_2),.clk(gclk));
	jdff dff_B_ZMKitu0y7_2(.din(w_dff_B_qX1pOQzH7_2),.dout(w_dff_B_ZMKitu0y7_2),.clk(gclk));
	jdff dff_B_9iVniqH93_2(.din(w_dff_B_ZMKitu0y7_2),.dout(w_dff_B_9iVniqH93_2),.clk(gclk));
	jdff dff_B_s7Y9Kv6W2_2(.din(w_dff_B_9iVniqH93_2),.dout(w_dff_B_s7Y9Kv6W2_2),.clk(gclk));
	jdff dff_B_fxrp6rHV6_2(.din(w_dff_B_s7Y9Kv6W2_2),.dout(w_dff_B_fxrp6rHV6_2),.clk(gclk));
	jdff dff_B_6soAIcis3_2(.din(w_dff_B_fxrp6rHV6_2),.dout(w_dff_B_6soAIcis3_2),.clk(gclk));
	jdff dff_B_EFZBgCdr0_2(.din(w_dff_B_6soAIcis3_2),.dout(w_dff_B_EFZBgCdr0_2),.clk(gclk));
	jdff dff_B_MK3I8beV8_2(.din(w_dff_B_EFZBgCdr0_2),.dout(w_dff_B_MK3I8beV8_2),.clk(gclk));
	jdff dff_B_EBLi6mFi8_2(.din(w_dff_B_MK3I8beV8_2),.dout(w_dff_B_EBLi6mFi8_2),.clk(gclk));
	jdff dff_B_UIuPmVgr4_2(.din(w_dff_B_EBLi6mFi8_2),.dout(w_dff_B_UIuPmVgr4_2),.clk(gclk));
	jdff dff_B_osNrJkuP9_2(.din(w_dff_B_UIuPmVgr4_2),.dout(w_dff_B_osNrJkuP9_2),.clk(gclk));
	jdff dff_B_Uptxipqr6_2(.din(w_dff_B_osNrJkuP9_2),.dout(w_dff_B_Uptxipqr6_2),.clk(gclk));
	jdff dff_B_aWfsZ3VJ7_2(.din(w_dff_B_Uptxipqr6_2),.dout(w_dff_B_aWfsZ3VJ7_2),.clk(gclk));
	jdff dff_B_RvqdFM2d3_2(.din(n1296),.dout(w_dff_B_RvqdFM2d3_2),.clk(gclk));
	jdff dff_B_0Gb9Fong5_1(.din(n1294),.dout(w_dff_B_0Gb9Fong5_1),.clk(gclk));
	jdff dff_B_g3Irwatn0_2(.din(n1203),.dout(w_dff_B_g3Irwatn0_2),.clk(gclk));
	jdff dff_B_S0Gbhlc82_2(.din(w_dff_B_g3Irwatn0_2),.dout(w_dff_B_S0Gbhlc82_2),.clk(gclk));
	jdff dff_B_gU5NsR8t5_2(.din(w_dff_B_S0Gbhlc82_2),.dout(w_dff_B_gU5NsR8t5_2),.clk(gclk));
	jdff dff_B_b35qg5Y62_2(.din(w_dff_B_gU5NsR8t5_2),.dout(w_dff_B_b35qg5Y62_2),.clk(gclk));
	jdff dff_B_aEIJ8oQw6_2(.din(w_dff_B_b35qg5Y62_2),.dout(w_dff_B_aEIJ8oQw6_2),.clk(gclk));
	jdff dff_B_yzTLXsOn9_2(.din(w_dff_B_aEIJ8oQw6_2),.dout(w_dff_B_yzTLXsOn9_2),.clk(gclk));
	jdff dff_B_lMm3TnGF6_2(.din(w_dff_B_yzTLXsOn9_2),.dout(w_dff_B_lMm3TnGF6_2),.clk(gclk));
	jdff dff_B_saLKSXE94_2(.din(w_dff_B_lMm3TnGF6_2),.dout(w_dff_B_saLKSXE94_2),.clk(gclk));
	jdff dff_B_G6WDknzh2_2(.din(w_dff_B_saLKSXE94_2),.dout(w_dff_B_G6WDknzh2_2),.clk(gclk));
	jdff dff_B_PQySZ21H7_2(.din(w_dff_B_G6WDknzh2_2),.dout(w_dff_B_PQySZ21H7_2),.clk(gclk));
	jdff dff_B_ud3fYL8c4_2(.din(w_dff_B_PQySZ21H7_2),.dout(w_dff_B_ud3fYL8c4_2),.clk(gclk));
	jdff dff_B_iaSJi1CZ6_2(.din(w_dff_B_ud3fYL8c4_2),.dout(w_dff_B_iaSJi1CZ6_2),.clk(gclk));
	jdff dff_B_6asxB7TE8_2(.din(w_dff_B_iaSJi1CZ6_2),.dout(w_dff_B_6asxB7TE8_2),.clk(gclk));
	jdff dff_B_y7WuCpIE4_2(.din(w_dff_B_6asxB7TE8_2),.dout(w_dff_B_y7WuCpIE4_2),.clk(gclk));
	jdff dff_B_FD98udlP0_2(.din(w_dff_B_y7WuCpIE4_2),.dout(w_dff_B_FD98udlP0_2),.clk(gclk));
	jdff dff_B_d372Oo5A1_2(.din(n1208),.dout(w_dff_B_d372Oo5A1_2),.clk(gclk));
	jdff dff_B_hyelq2598_2(.din(w_dff_B_d372Oo5A1_2),.dout(w_dff_B_hyelq2598_2),.clk(gclk));
	jdff dff_B_JYpE4nrd8_2(.din(w_dff_B_hyelq2598_2),.dout(w_dff_B_JYpE4nrd8_2),.clk(gclk));
	jdff dff_B_jjdl1HXT5_2(.din(w_dff_B_JYpE4nrd8_2),.dout(w_dff_B_jjdl1HXT5_2),.clk(gclk));
	jdff dff_B_1JzSWLQv2_2(.din(w_dff_B_jjdl1HXT5_2),.dout(w_dff_B_1JzSWLQv2_2),.clk(gclk));
	jdff dff_B_JtxHj3i14_2(.din(w_dff_B_1JzSWLQv2_2),.dout(w_dff_B_JtxHj3i14_2),.clk(gclk));
	jdff dff_B_AahmCqvJ0_2(.din(w_dff_B_JtxHj3i14_2),.dout(w_dff_B_AahmCqvJ0_2),.clk(gclk));
	jdff dff_B_igypnapb5_2(.din(w_dff_B_AahmCqvJ0_2),.dout(w_dff_B_igypnapb5_2),.clk(gclk));
	jdff dff_B_w3A1wWQ14_2(.din(w_dff_B_igypnapb5_2),.dout(w_dff_B_w3A1wWQ14_2),.clk(gclk));
	jdff dff_B_tweRq4vJ5_2(.din(w_dff_B_w3A1wWQ14_2),.dout(w_dff_B_tweRq4vJ5_2),.clk(gclk));
	jdff dff_B_Mi5d83Fo4_2(.din(w_dff_B_tweRq4vJ5_2),.dout(w_dff_B_Mi5d83Fo4_2),.clk(gclk));
	jdff dff_B_0sA4WOD92_2(.din(w_dff_B_Mi5d83Fo4_2),.dout(w_dff_B_0sA4WOD92_2),.clk(gclk));
	jdff dff_B_XVO8klnG6_2(.din(n1207),.dout(w_dff_B_XVO8klnG6_2),.clk(gclk));
	jdff dff_B_T5A98wyQ2_2(.din(w_dff_B_XVO8klnG6_2),.dout(w_dff_B_T5A98wyQ2_2),.clk(gclk));
	jdff dff_B_95UCo4TK0_2(.din(w_dff_B_T5A98wyQ2_2),.dout(w_dff_B_95UCo4TK0_2),.clk(gclk));
	jdff dff_B_KQWddzh79_2(.din(w_dff_B_95UCo4TK0_2),.dout(w_dff_B_KQWddzh79_2),.clk(gclk));
	jdff dff_B_sjtr7rUO1_2(.din(w_dff_B_KQWddzh79_2),.dout(w_dff_B_sjtr7rUO1_2),.clk(gclk));
	jdff dff_B_L7oXhL0G3_2(.din(w_dff_B_sjtr7rUO1_2),.dout(w_dff_B_L7oXhL0G3_2),.clk(gclk));
	jdff dff_B_38xMc8u08_2(.din(w_dff_B_L7oXhL0G3_2),.dout(w_dff_B_38xMc8u08_2),.clk(gclk));
	jdff dff_B_26EDGsq77_2(.din(w_dff_B_38xMc8u08_2),.dout(w_dff_B_26EDGsq77_2),.clk(gclk));
	jdff dff_B_xYulOIww0_2(.din(w_dff_B_26EDGsq77_2),.dout(w_dff_B_xYulOIww0_2),.clk(gclk));
	jdff dff_B_TV9oSqo39_2(.din(w_dff_B_xYulOIww0_2),.dout(w_dff_B_TV9oSqo39_2),.clk(gclk));
	jdff dff_B_lnBUZir81_2(.din(w_dff_B_TV9oSqo39_2),.dout(w_dff_B_lnBUZir81_2),.clk(gclk));
	jdff dff_B_f4sHwQoT5_2(.din(w_dff_B_lnBUZir81_2),.dout(w_dff_B_f4sHwQoT5_2),.clk(gclk));
	jdff dff_B_rHvJMzyq5_2(.din(w_dff_B_f4sHwQoT5_2),.dout(w_dff_B_rHvJMzyq5_2),.clk(gclk));
	jdff dff_B_fr1DhGc09_2(.din(w_dff_B_rHvJMzyq5_2),.dout(w_dff_B_fr1DhGc09_2),.clk(gclk));
	jdff dff_B_lu06mhQM1_2(.din(n1206),.dout(w_dff_B_lu06mhQM1_2),.clk(gclk));
	jdff dff_B_eYIqDh9G5_1(.din(n1204),.dout(w_dff_B_eYIqDh9G5_1),.clk(gclk));
	jdff dff_B_lPV6Fhfl4_2(.din(n1099),.dout(w_dff_B_lPV6Fhfl4_2),.clk(gclk));
	jdff dff_B_ixrbUdjT3_2(.din(w_dff_B_lPV6Fhfl4_2),.dout(w_dff_B_ixrbUdjT3_2),.clk(gclk));
	jdff dff_B_HtZglrRJ8_2(.din(w_dff_B_ixrbUdjT3_2),.dout(w_dff_B_HtZglrRJ8_2),.clk(gclk));
	jdff dff_B_ZSq65Qju7_2(.din(w_dff_B_HtZglrRJ8_2),.dout(w_dff_B_ZSq65Qju7_2),.clk(gclk));
	jdff dff_B_CbjeNfc21_2(.din(w_dff_B_ZSq65Qju7_2),.dout(w_dff_B_CbjeNfc21_2),.clk(gclk));
	jdff dff_B_dl6SEOlw9_2(.din(w_dff_B_CbjeNfc21_2),.dout(w_dff_B_dl6SEOlw9_2),.clk(gclk));
	jdff dff_B_thHIcPAa4_2(.din(w_dff_B_dl6SEOlw9_2),.dout(w_dff_B_thHIcPAa4_2),.clk(gclk));
	jdff dff_B_7vDaRG5I2_2(.din(w_dff_B_thHIcPAa4_2),.dout(w_dff_B_7vDaRG5I2_2),.clk(gclk));
	jdff dff_B_Wg7xHT2A3_2(.din(w_dff_B_7vDaRG5I2_2),.dout(w_dff_B_Wg7xHT2A3_2),.clk(gclk));
	jdff dff_B_f3hvHBZV4_2(.din(w_dff_B_Wg7xHT2A3_2),.dout(w_dff_B_f3hvHBZV4_2),.clk(gclk));
	jdff dff_B_fsycHxs66_2(.din(w_dff_B_f3hvHBZV4_2),.dout(w_dff_B_fsycHxs66_2),.clk(gclk));
	jdff dff_A_RhDR8iYU1_0(.dout(w_n1110_0[0]),.din(w_dff_A_RhDR8iYU1_0),.clk(gclk));
	jdff dff_A_MC7RPwqJ2_0(.dout(w_dff_A_RhDR8iYU1_0),.din(w_dff_A_MC7RPwqJ2_0),.clk(gclk));
	jdff dff_A_WmXhKVT75_0(.dout(w_dff_A_MC7RPwqJ2_0),.din(w_dff_A_WmXhKVT75_0),.clk(gclk));
	jdff dff_B_qHewBVZt4_2(.din(n1110),.dout(w_dff_B_qHewBVZt4_2),.clk(gclk));
	jdff dff_B_V60rxirR2_1(.din(n1104),.dout(w_dff_B_V60rxirR2_1),.clk(gclk));
	jdff dff_B_kbzGUNAt3_1(.din(w_dff_B_V60rxirR2_1),.dout(w_dff_B_kbzGUNAt3_1),.clk(gclk));
	jdff dff_B_suLSGBXS0_1(.din(w_dff_B_kbzGUNAt3_1),.dout(w_dff_B_suLSGBXS0_1),.clk(gclk));
	jdff dff_B_ML2YcFrR7_1(.din(w_dff_B_suLSGBXS0_1),.dout(w_dff_B_ML2YcFrR7_1),.clk(gclk));
	jdff dff_B_wgj4zyG66_1(.din(w_dff_B_ML2YcFrR7_1),.dout(w_dff_B_wgj4zyG66_1),.clk(gclk));
	jdff dff_B_rP85qQ8J0_1(.din(w_dff_B_wgj4zyG66_1),.dout(w_dff_B_rP85qQ8J0_1),.clk(gclk));
	jdff dff_B_NVAwxQ8j6_1(.din(n1105),.dout(w_dff_B_NVAwxQ8j6_1),.clk(gclk));
	jdff dff_B_hodFMUDZ4_1(.din(w_dff_B_NVAwxQ8j6_1),.dout(w_dff_B_hodFMUDZ4_1),.clk(gclk));
	jdff dff_A_WKPsJg287_1(.dout(w_G307gat_2[1]),.din(w_dff_A_WKPsJg287_1),.clk(gclk));
	jdff dff_A_tI8ZURF34_1(.dout(w_dff_A_WKPsJg287_1),.din(w_dff_A_tI8ZURF34_1),.clk(gclk));
	jdff dff_A_xPZGakul1_1(.dout(w_dff_A_tI8ZURF34_1),.din(w_dff_A_xPZGakul1_1),.clk(gclk));
	jdff dff_A_MEwpgw3j7_1(.dout(w_dff_A_xPZGakul1_1),.din(w_dff_A_MEwpgw3j7_1),.clk(gclk));
	jdff dff_A_d5cPW0z26_1(.dout(w_dff_A_MEwpgw3j7_1),.din(w_dff_A_d5cPW0z26_1),.clk(gclk));
	jdff dff_A_uPuFJxVi0_1(.dout(w_dff_A_d5cPW0z26_1),.din(w_dff_A_uPuFJxVi0_1),.clk(gclk));
	jdff dff_A_RSjd2ENx5_1(.dout(w_dff_A_uPuFJxVi0_1),.din(w_dff_A_RSjd2ENx5_1),.clk(gclk));
	jdff dff_B_VdZF60TW4_2(.din(n1103),.dout(w_dff_B_VdZF60TW4_2),.clk(gclk));
	jdff dff_B_k1MB6W6t7_2(.din(w_dff_B_VdZF60TW4_2),.dout(w_dff_B_k1MB6W6t7_2),.clk(gclk));
	jdff dff_B_gRaz6dBT7_2(.din(w_dff_B_k1MB6W6t7_2),.dout(w_dff_B_gRaz6dBT7_2),.clk(gclk));
	jdff dff_B_H79v9Uq58_2(.din(w_dff_B_gRaz6dBT7_2),.dout(w_dff_B_H79v9Uq58_2),.clk(gclk));
	jdff dff_B_Imlk7Eki1_2(.din(w_dff_B_H79v9Uq58_2),.dout(w_dff_B_Imlk7Eki1_2),.clk(gclk));
	jdff dff_B_hxtgEtn99_2(.din(w_dff_B_Imlk7Eki1_2),.dout(w_dff_B_hxtgEtn99_2),.clk(gclk));
	jdff dff_B_S1QBbm186_2(.din(w_dff_B_hxtgEtn99_2),.dout(w_dff_B_S1QBbm186_2),.clk(gclk));
	jdff dff_B_pkHOALHt4_2(.din(w_dff_B_S1QBbm186_2),.dout(w_dff_B_pkHOALHt4_2),.clk(gclk));
	jdff dff_B_hlGenjoK5_2(.din(w_dff_B_pkHOALHt4_2),.dout(w_dff_B_hlGenjoK5_2),.clk(gclk));
	jdff dff_B_jaHXtSYv4_2(.din(w_dff_B_hlGenjoK5_2),.dout(w_dff_B_jaHXtSYv4_2),.clk(gclk));
	jdff dff_B_BFY5D3Vg9_1(.din(n1100),.dout(w_dff_B_BFY5D3Vg9_1),.clk(gclk));
	jdff dff_B_m910XB5j8_2(.din(n1001),.dout(w_dff_B_m910XB5j8_2),.clk(gclk));
	jdff dff_B_vzdzVgz41_2(.din(w_dff_B_m910XB5j8_2),.dout(w_dff_B_vzdzVgz41_2),.clk(gclk));
	jdff dff_B_20BlkzZ02_2(.din(w_dff_B_vzdzVgz41_2),.dout(w_dff_B_20BlkzZ02_2),.clk(gclk));
	jdff dff_B_z58mmzRV5_2(.din(w_dff_B_20BlkzZ02_2),.dout(w_dff_B_z58mmzRV5_2),.clk(gclk));
	jdff dff_B_KocCuaqj5_2(.din(w_dff_B_z58mmzRV5_2),.dout(w_dff_B_KocCuaqj5_2),.clk(gclk));
	jdff dff_B_Y3yudIDv2_2(.din(w_dff_B_KocCuaqj5_2),.dout(w_dff_B_Y3yudIDv2_2),.clk(gclk));
	jdff dff_B_hgcUEBts6_2(.din(w_dff_B_Y3yudIDv2_2),.dout(w_dff_B_hgcUEBts6_2),.clk(gclk));
	jdff dff_B_N8ucdRpL4_2(.din(w_dff_B_hgcUEBts6_2),.dout(w_dff_B_N8ucdRpL4_2),.clk(gclk));
	jdff dff_B_rjpJ8Lqi1_2(.din(n1010),.dout(w_dff_B_rjpJ8Lqi1_2),.clk(gclk));
	jdff dff_B_S3wHjT2K0_2(.din(w_dff_B_rjpJ8Lqi1_2),.dout(w_dff_B_S3wHjT2K0_2),.clk(gclk));
	jdff dff_B_7hsdjXtW4_2(.din(w_dff_B_S3wHjT2K0_2),.dout(w_dff_B_7hsdjXtW4_2),.clk(gclk));
	jdff dff_B_9vzWDEwn2_2(.din(w_dff_B_7hsdjXtW4_2),.dout(w_dff_B_9vzWDEwn2_2),.clk(gclk));
	jdff dff_B_l45lPUQS4_2(.din(w_dff_B_9vzWDEwn2_2),.dout(w_dff_B_l45lPUQS4_2),.clk(gclk));
	jdff dff_A_08zg0qyi5_0(.dout(w_n1008_0[0]),.din(w_dff_A_08zg0qyi5_0),.clk(gclk));
	jdff dff_A_pMFqqMNj9_0(.dout(w_dff_A_08zg0qyi5_0),.din(w_dff_A_pMFqqMNj9_0),.clk(gclk));
	jdff dff_A_8xMT58BS1_0(.dout(w_dff_A_pMFqqMNj9_0),.din(w_dff_A_8xMT58BS1_0),.clk(gclk));
	jdff dff_A_SZgnYqYp9_0(.dout(w_n793_0[0]),.din(w_dff_A_SZgnYqYp9_0),.clk(gclk));
	jdff dff_A_tkYEQ15O7_1(.dout(w_n1006_0[1]),.din(w_dff_A_tkYEQ15O7_1),.clk(gclk));
	jdff dff_A_RxpTO1Zh9_1(.dout(w_dff_A_tkYEQ15O7_1),.din(w_dff_A_RxpTO1Zh9_1),.clk(gclk));
	jdff dff_B_0mee9hQv7_1(.din(n1002),.dout(w_dff_B_0mee9hQv7_1),.clk(gclk));
	jdff dff_B_l0KD2s4z2_1(.din(w_dff_B_0mee9hQv7_1),.dout(w_dff_B_l0KD2s4z2_1),.clk(gclk));
	jdff dff_B_oZbFmwUg7_1(.din(w_dff_B_l0KD2s4z2_1),.dout(w_dff_B_oZbFmwUg7_1),.clk(gclk));
	jdff dff_B_DCx1VC6Y7_1(.din(w_dff_B_oZbFmwUg7_1),.dout(w_dff_B_DCx1VC6Y7_1),.clk(gclk));
	jdff dff_B_rf367TDu7_1(.din(w_dff_B_DCx1VC6Y7_1),.dout(w_dff_B_rf367TDu7_1),.clk(gclk));
	jdff dff_A_mlAWXDW60_0(.dout(w_n903_0[0]),.din(w_dff_A_mlAWXDW60_0),.clk(gclk));
	jdff dff_A_rfFuhg8h4_0(.dout(w_dff_A_mlAWXDW60_0),.din(w_dff_A_rfFuhg8h4_0),.clk(gclk));
	jdff dff_A_YjJMEe3C2_0(.dout(w_dff_A_rfFuhg8h4_0),.din(w_dff_A_YjJMEe3C2_0),.clk(gclk));
	jdff dff_A_a9Fc5BLn6_0(.dout(w_n695_0[0]),.din(w_dff_A_a9Fc5BLn6_0),.clk(gclk));
	jdff dff_A_bmzQ5Z6I6_0(.dout(w_dff_A_a9Fc5BLn6_0),.din(w_dff_A_bmzQ5Z6I6_0),.clk(gclk));
	jdff dff_A_reLcFVwy2_0(.dout(w_dff_A_bmzQ5Z6I6_0),.din(w_dff_A_reLcFVwy2_0),.clk(gclk));
	jdff dff_B_9nAcROIB4_2(.din(n898),.dout(w_dff_B_9nAcROIB4_2),.clk(gclk));
	jdff dff_A_465exy0V6_1(.dout(w_n896_0[1]),.din(w_dff_A_465exy0V6_1),.clk(gclk));
	jdff dff_A_lZyKX5BD7_1(.dout(w_dff_A_465exy0V6_1),.din(w_dff_A_lZyKX5BD7_1),.clk(gclk));
	jdff dff_A_Tg2TvWQO4_1(.dout(w_dff_A_lZyKX5BD7_1),.din(w_dff_A_Tg2TvWQO4_1),.clk(gclk));
	jdff dff_A_TuVbJBvl8_1(.dout(w_dff_A_Tg2TvWQO4_1),.din(w_dff_A_TuVbJBvl8_1),.clk(gclk));
	jdff dff_A_8hSQ65zN0_1(.dout(w_dff_A_TuVbJBvl8_1),.din(w_dff_A_8hSQ65zN0_1),.clk(gclk));
	jdff dff_A_OnSTmqyq1_1(.dout(w_dff_A_u8sRXF6f7_0),.din(w_dff_A_OnSTmqyq1_1),.clk(gclk));
	jdff dff_A_u8sRXF6f7_0(.dout(w_dff_A_O7IBO4CG5_0),.din(w_dff_A_u8sRXF6f7_0),.clk(gclk));
	jdff dff_A_O7IBO4CG5_0(.dout(w_dff_A_uBqUbjxD5_0),.din(w_dff_A_O7IBO4CG5_0),.clk(gclk));
	jdff dff_A_uBqUbjxD5_0(.dout(w_dff_A_QnjCtdwm1_0),.din(w_dff_A_uBqUbjxD5_0),.clk(gclk));
	jdff dff_A_QnjCtdwm1_0(.dout(w_dff_A_aRGGjZYo6_0),.din(w_dff_A_QnjCtdwm1_0),.clk(gclk));
	jdff dff_A_aRGGjZYo6_0(.dout(w_dff_A_RjIseovg1_0),.din(w_dff_A_aRGGjZYo6_0),.clk(gclk));
	jdff dff_A_RjIseovg1_0(.dout(w_dff_A_wERotExv1_0),.din(w_dff_A_RjIseovg1_0),.clk(gclk));
	jdff dff_A_wERotExv1_0(.dout(w_dff_A_0gYpOujG3_0),.din(w_dff_A_wERotExv1_0),.clk(gclk));
	jdff dff_A_0gYpOujG3_0(.dout(w_dff_A_dyyIoITs1_0),.din(w_dff_A_0gYpOujG3_0),.clk(gclk));
	jdff dff_A_dyyIoITs1_0(.dout(w_dff_A_IRObgaE56_0),.din(w_dff_A_dyyIoITs1_0),.clk(gclk));
	jdff dff_A_IRObgaE56_0(.dout(w_dff_A_nQZ1IWK35_0),.din(w_dff_A_IRObgaE56_0),.clk(gclk));
	jdff dff_A_nQZ1IWK35_0(.dout(w_dff_A_TZ2Sz1g82_0),.din(w_dff_A_nQZ1IWK35_0),.clk(gclk));
	jdff dff_A_TZ2Sz1g82_0(.dout(w_dff_A_IjEeqSlc8_0),.din(w_dff_A_TZ2Sz1g82_0),.clk(gclk));
	jdff dff_A_IjEeqSlc8_0(.dout(w_dff_A_a5zOXXRW9_0),.din(w_dff_A_IjEeqSlc8_0),.clk(gclk));
	jdff dff_A_a5zOXXRW9_0(.dout(w_dff_A_UgOeq3E74_0),.din(w_dff_A_a5zOXXRW9_0),.clk(gclk));
	jdff dff_A_UgOeq3E74_0(.dout(w_dff_A_YhIT9Jj34_0),.din(w_dff_A_UgOeq3E74_0),.clk(gclk));
	jdff dff_A_YhIT9Jj34_0(.dout(w_dff_A_vpMQtO4F4_0),.din(w_dff_A_YhIT9Jj34_0),.clk(gclk));
	jdff dff_A_vpMQtO4F4_0(.dout(w_dff_A_ipGv5gIj3_0),.din(w_dff_A_vpMQtO4F4_0),.clk(gclk));
	jdff dff_A_ipGv5gIj3_0(.dout(w_dff_A_FbGLY1V18_0),.din(w_dff_A_ipGv5gIj3_0),.clk(gclk));
	jdff dff_A_FbGLY1V18_0(.dout(w_dff_A_7DRm5FfY8_0),.din(w_dff_A_FbGLY1V18_0),.clk(gclk));
	jdff dff_A_7DRm5FfY8_0(.dout(w_dff_A_kbvrLwRX2_0),.din(w_dff_A_7DRm5FfY8_0),.clk(gclk));
	jdff dff_A_kbvrLwRX2_0(.dout(w_dff_A_Wkw9DGp21_0),.din(w_dff_A_kbvrLwRX2_0),.clk(gclk));
	jdff dff_A_Wkw9DGp21_0(.dout(w_dff_A_UvEGBe7f5_0),.din(w_dff_A_Wkw9DGp21_0),.clk(gclk));
	jdff dff_A_UvEGBe7f5_0(.dout(w_dff_A_nRvBmrCg1_0),.din(w_dff_A_UvEGBe7f5_0),.clk(gclk));
	jdff dff_A_nRvBmrCg1_0(.dout(w_dff_A_SPsbKPKH1_0),.din(w_dff_A_nRvBmrCg1_0),.clk(gclk));
	jdff dff_A_SPsbKPKH1_0(.dout(w_dff_A_eVTDbam93_0),.din(w_dff_A_SPsbKPKH1_0),.clk(gclk));
	jdff dff_A_eVTDbam93_0(.dout(w_dff_A_Wt9gVfJI8_0),.din(w_dff_A_eVTDbam93_0),.clk(gclk));
	jdff dff_A_Wt9gVfJI8_0(.dout(w_dff_A_Eiz2eeZs1_0),.din(w_dff_A_Wt9gVfJI8_0),.clk(gclk));
	jdff dff_A_Eiz2eeZs1_0(.dout(w_dff_A_R3afGlWJ6_0),.din(w_dff_A_Eiz2eeZs1_0),.clk(gclk));
	jdff dff_A_R3afGlWJ6_0(.dout(w_dff_A_CdI7CRYe4_0),.din(w_dff_A_R3afGlWJ6_0),.clk(gclk));
	jdff dff_A_CdI7CRYe4_0(.dout(w_dff_A_KkAMD7Cx9_0),.din(w_dff_A_CdI7CRYe4_0),.clk(gclk));
	jdff dff_A_KkAMD7Cx9_0(.dout(w_dff_A_li4NKrln5_0),.din(w_dff_A_KkAMD7Cx9_0),.clk(gclk));
	jdff dff_A_li4NKrln5_0(.dout(w_dff_A_oqjCF0In6_0),.din(w_dff_A_li4NKrln5_0),.clk(gclk));
	jdff dff_A_oqjCF0In6_0(.dout(w_dff_A_FE5wqB124_0),.din(w_dff_A_oqjCF0In6_0),.clk(gclk));
	jdff dff_A_FE5wqB124_0(.dout(w_dff_A_4R16xZrH7_0),.din(w_dff_A_FE5wqB124_0),.clk(gclk));
	jdff dff_A_4R16xZrH7_0(.dout(w_dff_A_LJOV3Lxx9_0),.din(w_dff_A_4R16xZrH7_0),.clk(gclk));
	jdff dff_A_LJOV3Lxx9_0(.dout(w_dff_A_MGOwzsVF3_0),.din(w_dff_A_LJOV3Lxx9_0),.clk(gclk));
	jdff dff_A_MGOwzsVF3_0(.dout(w_dff_A_lyksgwbU2_0),.din(w_dff_A_MGOwzsVF3_0),.clk(gclk));
	jdff dff_A_lyksgwbU2_0(.dout(w_dff_A_86477Pek7_0),.din(w_dff_A_lyksgwbU2_0),.clk(gclk));
	jdff dff_A_86477Pek7_0(.dout(w_dff_A_c54GyUP38_0),.din(w_dff_A_86477Pek7_0),.clk(gclk));
	jdff dff_A_c54GyUP38_0(.dout(w_dff_A_mASEeWWt9_0),.din(w_dff_A_c54GyUP38_0),.clk(gclk));
	jdff dff_A_mASEeWWt9_0(.dout(w_dff_A_mj9Fs4110_0),.din(w_dff_A_mASEeWWt9_0),.clk(gclk));
	jdff dff_A_mj9Fs4110_0(.dout(w_dff_A_0Jazty1V2_0),.din(w_dff_A_mj9Fs4110_0),.clk(gclk));
	jdff dff_A_0Jazty1V2_0(.dout(w_dff_A_WHN79rNy5_0),.din(w_dff_A_0Jazty1V2_0),.clk(gclk));
	jdff dff_A_WHN79rNy5_0(.dout(w_dff_A_4lCsJIWU6_0),.din(w_dff_A_WHN79rNy5_0),.clk(gclk));
	jdff dff_A_4lCsJIWU6_0(.dout(w_dff_A_dE0hqBcc4_0),.din(w_dff_A_4lCsJIWU6_0),.clk(gclk));
	jdff dff_A_dE0hqBcc4_0(.dout(w_dff_A_Ls5lsSD16_0),.din(w_dff_A_dE0hqBcc4_0),.clk(gclk));
	jdff dff_A_Ls5lsSD16_0(.dout(w_dff_A_vwyglYq09_0),.din(w_dff_A_Ls5lsSD16_0),.clk(gclk));
	jdff dff_A_vwyglYq09_0(.dout(w_dff_A_kFViTijJ7_0),.din(w_dff_A_vwyglYq09_0),.clk(gclk));
	jdff dff_A_kFViTijJ7_0(.dout(w_dff_A_vPsWXsLZ0_0),.din(w_dff_A_kFViTijJ7_0),.clk(gclk));
	jdff dff_A_vPsWXsLZ0_0(.dout(w_dff_A_is7H95T40_0),.din(w_dff_A_vPsWXsLZ0_0),.clk(gclk));
	jdff dff_A_is7H95T40_0(.dout(w_dff_A_mXrHs79t9_0),.din(w_dff_A_is7H95T40_0),.clk(gclk));
	jdff dff_A_mXrHs79t9_0(.dout(w_dff_A_hKa7peHF0_0),.din(w_dff_A_mXrHs79t9_0),.clk(gclk));
	jdff dff_A_hKa7peHF0_0(.dout(w_dff_A_8dxI3AM84_0),.din(w_dff_A_hKa7peHF0_0),.clk(gclk));
	jdff dff_A_8dxI3AM84_0(.dout(w_dff_A_iuYQRbip0_0),.din(w_dff_A_8dxI3AM84_0),.clk(gclk));
	jdff dff_A_iuYQRbip0_0(.dout(w_dff_A_KnGhanup8_0),.din(w_dff_A_iuYQRbip0_0),.clk(gclk));
	jdff dff_A_KnGhanup8_0(.dout(w_dff_A_qEq9LsPR5_0),.din(w_dff_A_KnGhanup8_0),.clk(gclk));
	jdff dff_A_qEq9LsPR5_0(.dout(w_dff_A_hIjfV8Al0_0),.din(w_dff_A_qEq9LsPR5_0),.clk(gclk));
	jdff dff_A_hIjfV8Al0_0(.dout(w_dff_A_I3bJZEvu1_0),.din(w_dff_A_hIjfV8Al0_0),.clk(gclk));
	jdff dff_A_I3bJZEvu1_0(.dout(w_dff_A_VJfYeyLo8_0),.din(w_dff_A_I3bJZEvu1_0),.clk(gclk));
	jdff dff_A_VJfYeyLo8_0(.dout(w_dff_A_rR5XOtlX0_0),.din(w_dff_A_VJfYeyLo8_0),.clk(gclk));
	jdff dff_A_rR5XOtlX0_0(.dout(w_dff_A_P7RDMqrv4_0),.din(w_dff_A_rR5XOtlX0_0),.clk(gclk));
	jdff dff_A_P7RDMqrv4_0(.dout(w_dff_A_Yw1rUEkr6_0),.din(w_dff_A_P7RDMqrv4_0),.clk(gclk));
	jdff dff_A_Yw1rUEkr6_0(.dout(w_dff_A_8pWPZ5so7_0),.din(w_dff_A_Yw1rUEkr6_0),.clk(gclk));
	jdff dff_A_8pWPZ5so7_0(.dout(w_dff_A_TCKFPob91_0),.din(w_dff_A_8pWPZ5so7_0),.clk(gclk));
	jdff dff_A_TCKFPob91_0(.dout(w_dff_A_iXOKyWzx4_0),.din(w_dff_A_TCKFPob91_0),.clk(gclk));
	jdff dff_A_iXOKyWzx4_0(.dout(w_dff_A_y4qfZ9Im3_0),.din(w_dff_A_iXOKyWzx4_0),.clk(gclk));
	jdff dff_A_y4qfZ9Im3_0(.dout(w_dff_A_ZaDG8Mq34_0),.din(w_dff_A_y4qfZ9Im3_0),.clk(gclk));
	jdff dff_A_ZaDG8Mq34_0(.dout(w_dff_A_W1qK3Myh1_0),.din(w_dff_A_ZaDG8Mq34_0),.clk(gclk));
	jdff dff_A_W1qK3Myh1_0(.dout(w_dff_A_MbeK9Jcu1_0),.din(w_dff_A_W1qK3Myh1_0),.clk(gclk));
	jdff dff_A_MbeK9Jcu1_0(.dout(w_dff_A_54b37qpb1_0),.din(w_dff_A_MbeK9Jcu1_0),.clk(gclk));
	jdff dff_A_54b37qpb1_0(.dout(w_dff_A_2Efcu3yJ9_0),.din(w_dff_A_54b37qpb1_0),.clk(gclk));
	jdff dff_A_2Efcu3yJ9_0(.dout(w_dff_A_JQbFPgSh8_0),.din(w_dff_A_2Efcu3yJ9_0),.clk(gclk));
	jdff dff_A_JQbFPgSh8_0(.dout(w_dff_A_nW1ypwyI6_0),.din(w_dff_A_JQbFPgSh8_0),.clk(gclk));
	jdff dff_A_nW1ypwyI6_0(.dout(G545gat),.din(w_dff_A_nW1ypwyI6_0),.clk(gclk));
	jdff dff_A_7d1LhOvD7_2(.dout(w_dff_A_rvczDX1L2_0),.din(w_dff_A_7d1LhOvD7_2),.clk(gclk));
	jdff dff_A_rvczDX1L2_0(.dout(w_dff_A_sLsmbTZ66_0),.din(w_dff_A_rvczDX1L2_0),.clk(gclk));
	jdff dff_A_sLsmbTZ66_0(.dout(w_dff_A_Wg7qmMMc2_0),.din(w_dff_A_sLsmbTZ66_0),.clk(gclk));
	jdff dff_A_Wg7qmMMc2_0(.dout(w_dff_A_QWAcJONC2_0),.din(w_dff_A_Wg7qmMMc2_0),.clk(gclk));
	jdff dff_A_QWAcJONC2_0(.dout(w_dff_A_NXbXGzJ11_0),.din(w_dff_A_QWAcJONC2_0),.clk(gclk));
	jdff dff_A_NXbXGzJ11_0(.dout(w_dff_A_LNGtkm7A0_0),.din(w_dff_A_NXbXGzJ11_0),.clk(gclk));
	jdff dff_A_LNGtkm7A0_0(.dout(w_dff_A_v03aTqCa8_0),.din(w_dff_A_LNGtkm7A0_0),.clk(gclk));
	jdff dff_A_v03aTqCa8_0(.dout(w_dff_A_PvXQ8A7N6_0),.din(w_dff_A_v03aTqCa8_0),.clk(gclk));
	jdff dff_A_PvXQ8A7N6_0(.dout(w_dff_A_Rg34ntno7_0),.din(w_dff_A_PvXQ8A7N6_0),.clk(gclk));
	jdff dff_A_Rg34ntno7_0(.dout(w_dff_A_tJHxOajH5_0),.din(w_dff_A_Rg34ntno7_0),.clk(gclk));
	jdff dff_A_tJHxOajH5_0(.dout(w_dff_A_b9E0guGl5_0),.din(w_dff_A_tJHxOajH5_0),.clk(gclk));
	jdff dff_A_b9E0guGl5_0(.dout(w_dff_A_lw1IlMQZ0_0),.din(w_dff_A_b9E0guGl5_0),.clk(gclk));
	jdff dff_A_lw1IlMQZ0_0(.dout(w_dff_A_mYcqDf071_0),.din(w_dff_A_lw1IlMQZ0_0),.clk(gclk));
	jdff dff_A_mYcqDf071_0(.dout(w_dff_A_RiVu5ex30_0),.din(w_dff_A_mYcqDf071_0),.clk(gclk));
	jdff dff_A_RiVu5ex30_0(.dout(w_dff_A_IL7RVIdG0_0),.din(w_dff_A_RiVu5ex30_0),.clk(gclk));
	jdff dff_A_IL7RVIdG0_0(.dout(w_dff_A_Goycacxx8_0),.din(w_dff_A_IL7RVIdG0_0),.clk(gclk));
	jdff dff_A_Goycacxx8_0(.dout(w_dff_A_opmy3WvA4_0),.din(w_dff_A_Goycacxx8_0),.clk(gclk));
	jdff dff_A_opmy3WvA4_0(.dout(w_dff_A_jVbglBum3_0),.din(w_dff_A_opmy3WvA4_0),.clk(gclk));
	jdff dff_A_jVbglBum3_0(.dout(w_dff_A_Ac8D5KiO0_0),.din(w_dff_A_jVbglBum3_0),.clk(gclk));
	jdff dff_A_Ac8D5KiO0_0(.dout(w_dff_A_RZowy2XY7_0),.din(w_dff_A_Ac8D5KiO0_0),.clk(gclk));
	jdff dff_A_RZowy2XY7_0(.dout(w_dff_A_KqatYKAM2_0),.din(w_dff_A_RZowy2XY7_0),.clk(gclk));
	jdff dff_A_KqatYKAM2_0(.dout(w_dff_A_iI9MGEWT4_0),.din(w_dff_A_KqatYKAM2_0),.clk(gclk));
	jdff dff_A_iI9MGEWT4_0(.dout(w_dff_A_wHGDIevi8_0),.din(w_dff_A_iI9MGEWT4_0),.clk(gclk));
	jdff dff_A_wHGDIevi8_0(.dout(w_dff_A_wKkHWfzP7_0),.din(w_dff_A_wHGDIevi8_0),.clk(gclk));
	jdff dff_A_wKkHWfzP7_0(.dout(w_dff_A_kUIoZqy33_0),.din(w_dff_A_wKkHWfzP7_0),.clk(gclk));
	jdff dff_A_kUIoZqy33_0(.dout(w_dff_A_A78dhmsf1_0),.din(w_dff_A_kUIoZqy33_0),.clk(gclk));
	jdff dff_A_A78dhmsf1_0(.dout(w_dff_A_gIJTDeFf4_0),.din(w_dff_A_A78dhmsf1_0),.clk(gclk));
	jdff dff_A_gIJTDeFf4_0(.dout(w_dff_A_RiCB1H3h2_0),.din(w_dff_A_gIJTDeFf4_0),.clk(gclk));
	jdff dff_A_RiCB1H3h2_0(.dout(w_dff_A_lOI8om2V0_0),.din(w_dff_A_RiCB1H3h2_0),.clk(gclk));
	jdff dff_A_lOI8om2V0_0(.dout(w_dff_A_bNW4aXBV0_0),.din(w_dff_A_lOI8om2V0_0),.clk(gclk));
	jdff dff_A_bNW4aXBV0_0(.dout(w_dff_A_K3xSEreo1_0),.din(w_dff_A_bNW4aXBV0_0),.clk(gclk));
	jdff dff_A_K3xSEreo1_0(.dout(w_dff_A_dVCcKt8d7_0),.din(w_dff_A_K3xSEreo1_0),.clk(gclk));
	jdff dff_A_dVCcKt8d7_0(.dout(w_dff_A_3C7lMoD16_0),.din(w_dff_A_dVCcKt8d7_0),.clk(gclk));
	jdff dff_A_3C7lMoD16_0(.dout(w_dff_A_8iyDK62l3_0),.din(w_dff_A_3C7lMoD16_0),.clk(gclk));
	jdff dff_A_8iyDK62l3_0(.dout(w_dff_A_TB05FPcS2_0),.din(w_dff_A_8iyDK62l3_0),.clk(gclk));
	jdff dff_A_TB05FPcS2_0(.dout(w_dff_A_YY1ktvQR6_0),.din(w_dff_A_TB05FPcS2_0),.clk(gclk));
	jdff dff_A_YY1ktvQR6_0(.dout(w_dff_A_8xwuFCjV3_0),.din(w_dff_A_YY1ktvQR6_0),.clk(gclk));
	jdff dff_A_8xwuFCjV3_0(.dout(w_dff_A_8TjjNzAq3_0),.din(w_dff_A_8xwuFCjV3_0),.clk(gclk));
	jdff dff_A_8TjjNzAq3_0(.dout(w_dff_A_H1WrmOOh5_0),.din(w_dff_A_8TjjNzAq3_0),.clk(gclk));
	jdff dff_A_H1WrmOOh5_0(.dout(w_dff_A_F1bXCwum3_0),.din(w_dff_A_H1WrmOOh5_0),.clk(gclk));
	jdff dff_A_F1bXCwum3_0(.dout(w_dff_A_czNI0Agy8_0),.din(w_dff_A_F1bXCwum3_0),.clk(gclk));
	jdff dff_A_czNI0Agy8_0(.dout(w_dff_A_SE8FeqzN4_0),.din(w_dff_A_czNI0Agy8_0),.clk(gclk));
	jdff dff_A_SE8FeqzN4_0(.dout(w_dff_A_CWiZwwt58_0),.din(w_dff_A_SE8FeqzN4_0),.clk(gclk));
	jdff dff_A_CWiZwwt58_0(.dout(w_dff_A_i7kBb1Zc1_0),.din(w_dff_A_CWiZwwt58_0),.clk(gclk));
	jdff dff_A_i7kBb1Zc1_0(.dout(w_dff_A_3OHjbTN80_0),.din(w_dff_A_i7kBb1Zc1_0),.clk(gclk));
	jdff dff_A_3OHjbTN80_0(.dout(w_dff_A_nhDOU8Jb7_0),.din(w_dff_A_3OHjbTN80_0),.clk(gclk));
	jdff dff_A_nhDOU8Jb7_0(.dout(w_dff_A_80FsTp2J1_0),.din(w_dff_A_nhDOU8Jb7_0),.clk(gclk));
	jdff dff_A_80FsTp2J1_0(.dout(w_dff_A_bu4DrZPu4_0),.din(w_dff_A_80FsTp2J1_0),.clk(gclk));
	jdff dff_A_bu4DrZPu4_0(.dout(w_dff_A_AyJjQC3H0_0),.din(w_dff_A_bu4DrZPu4_0),.clk(gclk));
	jdff dff_A_AyJjQC3H0_0(.dout(w_dff_A_8EacnzDo2_0),.din(w_dff_A_AyJjQC3H0_0),.clk(gclk));
	jdff dff_A_8EacnzDo2_0(.dout(w_dff_A_wB3jjJIo3_0),.din(w_dff_A_8EacnzDo2_0),.clk(gclk));
	jdff dff_A_wB3jjJIo3_0(.dout(w_dff_A_oR9lj3Cj3_0),.din(w_dff_A_wB3jjJIo3_0),.clk(gclk));
	jdff dff_A_oR9lj3Cj3_0(.dout(w_dff_A_NjBX5f7n4_0),.din(w_dff_A_oR9lj3Cj3_0),.clk(gclk));
	jdff dff_A_NjBX5f7n4_0(.dout(w_dff_A_6d6rJqBF1_0),.din(w_dff_A_NjBX5f7n4_0),.clk(gclk));
	jdff dff_A_6d6rJqBF1_0(.dout(w_dff_A_NrdAXYeZ4_0),.din(w_dff_A_6d6rJqBF1_0),.clk(gclk));
	jdff dff_A_NrdAXYeZ4_0(.dout(w_dff_A_8bGzGdwd0_0),.din(w_dff_A_NrdAXYeZ4_0),.clk(gclk));
	jdff dff_A_8bGzGdwd0_0(.dout(w_dff_A_o2tMKMkp2_0),.din(w_dff_A_8bGzGdwd0_0),.clk(gclk));
	jdff dff_A_o2tMKMkp2_0(.dout(w_dff_A_8jEqjpPQ3_0),.din(w_dff_A_o2tMKMkp2_0),.clk(gclk));
	jdff dff_A_8jEqjpPQ3_0(.dout(w_dff_A_w3gmyqSr3_0),.din(w_dff_A_8jEqjpPQ3_0),.clk(gclk));
	jdff dff_A_w3gmyqSr3_0(.dout(w_dff_A_NFynntpd8_0),.din(w_dff_A_w3gmyqSr3_0),.clk(gclk));
	jdff dff_A_NFynntpd8_0(.dout(w_dff_A_1lAAMchZ3_0),.din(w_dff_A_NFynntpd8_0),.clk(gclk));
	jdff dff_A_1lAAMchZ3_0(.dout(w_dff_A_Ne5boROJ6_0),.din(w_dff_A_1lAAMchZ3_0),.clk(gclk));
	jdff dff_A_Ne5boROJ6_0(.dout(w_dff_A_dGOd6PBg2_0),.din(w_dff_A_Ne5boROJ6_0),.clk(gclk));
	jdff dff_A_dGOd6PBg2_0(.dout(w_dff_A_S0SUIxPg2_0),.din(w_dff_A_dGOd6PBg2_0),.clk(gclk));
	jdff dff_A_S0SUIxPg2_0(.dout(w_dff_A_jRb1ubOH0_0),.din(w_dff_A_S0SUIxPg2_0),.clk(gclk));
	jdff dff_A_jRb1ubOH0_0(.dout(w_dff_A_IInP2Buv4_0),.din(w_dff_A_jRb1ubOH0_0),.clk(gclk));
	jdff dff_A_IInP2Buv4_0(.dout(w_dff_A_eOqaNz979_0),.din(w_dff_A_IInP2Buv4_0),.clk(gclk));
	jdff dff_A_eOqaNz979_0(.dout(w_dff_A_p7U3kNJM0_0),.din(w_dff_A_eOqaNz979_0),.clk(gclk));
	jdff dff_A_p7U3kNJM0_0(.dout(w_dff_A_jtKUE8BM5_0),.din(w_dff_A_p7U3kNJM0_0),.clk(gclk));
	jdff dff_A_jtKUE8BM5_0(.dout(w_dff_A_BkkyqPNt8_0),.din(w_dff_A_jtKUE8BM5_0),.clk(gclk));
	jdff dff_A_BkkyqPNt8_0(.dout(w_dff_A_bZQbIqBj5_0),.din(w_dff_A_BkkyqPNt8_0),.clk(gclk));
	jdff dff_A_bZQbIqBj5_0(.dout(G1581gat),.din(w_dff_A_bZQbIqBj5_0),.clk(gclk));
	jdff dff_A_e8HaFF4D6_2(.dout(w_dff_A_ZZg83iRK9_0),.din(w_dff_A_e8HaFF4D6_2),.clk(gclk));
	jdff dff_A_ZZg83iRK9_0(.dout(w_dff_A_1ELkWDTe3_0),.din(w_dff_A_ZZg83iRK9_0),.clk(gclk));
	jdff dff_A_1ELkWDTe3_0(.dout(w_dff_A_vnFrLtHI5_0),.din(w_dff_A_1ELkWDTe3_0),.clk(gclk));
	jdff dff_A_vnFrLtHI5_0(.dout(w_dff_A_oDQXVNpp3_0),.din(w_dff_A_vnFrLtHI5_0),.clk(gclk));
	jdff dff_A_oDQXVNpp3_0(.dout(w_dff_A_mdfKnGhh8_0),.din(w_dff_A_oDQXVNpp3_0),.clk(gclk));
	jdff dff_A_mdfKnGhh8_0(.dout(w_dff_A_O3K9QHJD2_0),.din(w_dff_A_mdfKnGhh8_0),.clk(gclk));
	jdff dff_A_O3K9QHJD2_0(.dout(w_dff_A_2BX4wbWT0_0),.din(w_dff_A_O3K9QHJD2_0),.clk(gclk));
	jdff dff_A_2BX4wbWT0_0(.dout(w_dff_A_ixwumU436_0),.din(w_dff_A_2BX4wbWT0_0),.clk(gclk));
	jdff dff_A_ixwumU436_0(.dout(w_dff_A_tR5rl26t7_0),.din(w_dff_A_ixwumU436_0),.clk(gclk));
	jdff dff_A_tR5rl26t7_0(.dout(w_dff_A_AH08WWq24_0),.din(w_dff_A_tR5rl26t7_0),.clk(gclk));
	jdff dff_A_AH08WWq24_0(.dout(w_dff_A_dX3eqge23_0),.din(w_dff_A_AH08WWq24_0),.clk(gclk));
	jdff dff_A_dX3eqge23_0(.dout(w_dff_A_zVugR1mv3_0),.din(w_dff_A_dX3eqge23_0),.clk(gclk));
	jdff dff_A_zVugR1mv3_0(.dout(w_dff_A_JiBEC2kq1_0),.din(w_dff_A_zVugR1mv3_0),.clk(gclk));
	jdff dff_A_JiBEC2kq1_0(.dout(w_dff_A_DSkflptN6_0),.din(w_dff_A_JiBEC2kq1_0),.clk(gclk));
	jdff dff_A_DSkflptN6_0(.dout(w_dff_A_1cydg5nh3_0),.din(w_dff_A_DSkflptN6_0),.clk(gclk));
	jdff dff_A_1cydg5nh3_0(.dout(w_dff_A_KD3R02fk3_0),.din(w_dff_A_1cydg5nh3_0),.clk(gclk));
	jdff dff_A_KD3R02fk3_0(.dout(w_dff_A_Ntnv9MjG3_0),.din(w_dff_A_KD3R02fk3_0),.clk(gclk));
	jdff dff_A_Ntnv9MjG3_0(.dout(w_dff_A_NWqy4acc9_0),.din(w_dff_A_Ntnv9MjG3_0),.clk(gclk));
	jdff dff_A_NWqy4acc9_0(.dout(w_dff_A_i4GF1qP82_0),.din(w_dff_A_NWqy4acc9_0),.clk(gclk));
	jdff dff_A_i4GF1qP82_0(.dout(w_dff_A_lIzvw1CS9_0),.din(w_dff_A_i4GF1qP82_0),.clk(gclk));
	jdff dff_A_lIzvw1CS9_0(.dout(w_dff_A_JwLov5Xj2_0),.din(w_dff_A_lIzvw1CS9_0),.clk(gclk));
	jdff dff_A_JwLov5Xj2_0(.dout(w_dff_A_zL6EUY6B3_0),.din(w_dff_A_JwLov5Xj2_0),.clk(gclk));
	jdff dff_A_zL6EUY6B3_0(.dout(w_dff_A_sACBSGvS2_0),.din(w_dff_A_zL6EUY6B3_0),.clk(gclk));
	jdff dff_A_sACBSGvS2_0(.dout(w_dff_A_rObrAbyh5_0),.din(w_dff_A_sACBSGvS2_0),.clk(gclk));
	jdff dff_A_rObrAbyh5_0(.dout(w_dff_A_F8mBgC9n2_0),.din(w_dff_A_rObrAbyh5_0),.clk(gclk));
	jdff dff_A_F8mBgC9n2_0(.dout(w_dff_A_Pzjv24El2_0),.din(w_dff_A_F8mBgC9n2_0),.clk(gclk));
	jdff dff_A_Pzjv24El2_0(.dout(w_dff_A_Aif2BL8Q7_0),.din(w_dff_A_Pzjv24El2_0),.clk(gclk));
	jdff dff_A_Aif2BL8Q7_0(.dout(w_dff_A_WDTI2AWs7_0),.din(w_dff_A_Aif2BL8Q7_0),.clk(gclk));
	jdff dff_A_WDTI2AWs7_0(.dout(w_dff_A_QMehkqT62_0),.din(w_dff_A_WDTI2AWs7_0),.clk(gclk));
	jdff dff_A_QMehkqT62_0(.dout(w_dff_A_Y8lwrufa9_0),.din(w_dff_A_QMehkqT62_0),.clk(gclk));
	jdff dff_A_Y8lwrufa9_0(.dout(w_dff_A_2nP9Ufdi4_0),.din(w_dff_A_Y8lwrufa9_0),.clk(gclk));
	jdff dff_A_2nP9Ufdi4_0(.dout(w_dff_A_9ftYyt6u2_0),.din(w_dff_A_2nP9Ufdi4_0),.clk(gclk));
	jdff dff_A_9ftYyt6u2_0(.dout(w_dff_A_kWSAGsnT8_0),.din(w_dff_A_9ftYyt6u2_0),.clk(gclk));
	jdff dff_A_kWSAGsnT8_0(.dout(w_dff_A_32jPwhUT7_0),.din(w_dff_A_kWSAGsnT8_0),.clk(gclk));
	jdff dff_A_32jPwhUT7_0(.dout(w_dff_A_fkZe9YOD5_0),.din(w_dff_A_32jPwhUT7_0),.clk(gclk));
	jdff dff_A_fkZe9YOD5_0(.dout(w_dff_A_dimGw5UX6_0),.din(w_dff_A_fkZe9YOD5_0),.clk(gclk));
	jdff dff_A_dimGw5UX6_0(.dout(w_dff_A_kW56nKPb5_0),.din(w_dff_A_dimGw5UX6_0),.clk(gclk));
	jdff dff_A_kW56nKPb5_0(.dout(w_dff_A_lyDQ4kJU5_0),.din(w_dff_A_kW56nKPb5_0),.clk(gclk));
	jdff dff_A_lyDQ4kJU5_0(.dout(w_dff_A_eh7A5qZo0_0),.din(w_dff_A_lyDQ4kJU5_0),.clk(gclk));
	jdff dff_A_eh7A5qZo0_0(.dout(w_dff_A_c3Pnpf1J1_0),.din(w_dff_A_eh7A5qZo0_0),.clk(gclk));
	jdff dff_A_c3Pnpf1J1_0(.dout(w_dff_A_VDThfbob4_0),.din(w_dff_A_c3Pnpf1J1_0),.clk(gclk));
	jdff dff_A_VDThfbob4_0(.dout(w_dff_A_3GIsObAc5_0),.din(w_dff_A_VDThfbob4_0),.clk(gclk));
	jdff dff_A_3GIsObAc5_0(.dout(w_dff_A_9YWWJm5T3_0),.din(w_dff_A_3GIsObAc5_0),.clk(gclk));
	jdff dff_A_9YWWJm5T3_0(.dout(w_dff_A_ZXVFgdLK3_0),.din(w_dff_A_9YWWJm5T3_0),.clk(gclk));
	jdff dff_A_ZXVFgdLK3_0(.dout(w_dff_A_o4gPJLkS2_0),.din(w_dff_A_ZXVFgdLK3_0),.clk(gclk));
	jdff dff_A_o4gPJLkS2_0(.dout(w_dff_A_FNTkhPLx7_0),.din(w_dff_A_o4gPJLkS2_0),.clk(gclk));
	jdff dff_A_FNTkhPLx7_0(.dout(w_dff_A_1dfbKyYl6_0),.din(w_dff_A_FNTkhPLx7_0),.clk(gclk));
	jdff dff_A_1dfbKyYl6_0(.dout(w_dff_A_NkXw6eyl4_0),.din(w_dff_A_1dfbKyYl6_0),.clk(gclk));
	jdff dff_A_NkXw6eyl4_0(.dout(w_dff_A_LhDLpsCR0_0),.din(w_dff_A_NkXw6eyl4_0),.clk(gclk));
	jdff dff_A_LhDLpsCR0_0(.dout(w_dff_A_kR2dOtYY0_0),.din(w_dff_A_LhDLpsCR0_0),.clk(gclk));
	jdff dff_A_kR2dOtYY0_0(.dout(w_dff_A_NmTd3ng58_0),.din(w_dff_A_kR2dOtYY0_0),.clk(gclk));
	jdff dff_A_NmTd3ng58_0(.dout(w_dff_A_ApbI0e9z0_0),.din(w_dff_A_NmTd3ng58_0),.clk(gclk));
	jdff dff_A_ApbI0e9z0_0(.dout(w_dff_A_nj1SBpVm6_0),.din(w_dff_A_ApbI0e9z0_0),.clk(gclk));
	jdff dff_A_nj1SBpVm6_0(.dout(w_dff_A_7OoIpG8y9_0),.din(w_dff_A_nj1SBpVm6_0),.clk(gclk));
	jdff dff_A_7OoIpG8y9_0(.dout(w_dff_A_pXZbzZkY2_0),.din(w_dff_A_7OoIpG8y9_0),.clk(gclk));
	jdff dff_A_pXZbzZkY2_0(.dout(w_dff_A_fNoTmXkC1_0),.din(w_dff_A_pXZbzZkY2_0),.clk(gclk));
	jdff dff_A_fNoTmXkC1_0(.dout(w_dff_A_vnDR5rbC2_0),.din(w_dff_A_fNoTmXkC1_0),.clk(gclk));
	jdff dff_A_vnDR5rbC2_0(.dout(w_dff_A_SbuqzeQm8_0),.din(w_dff_A_vnDR5rbC2_0),.clk(gclk));
	jdff dff_A_SbuqzeQm8_0(.dout(w_dff_A_gVE3prvY1_0),.din(w_dff_A_SbuqzeQm8_0),.clk(gclk));
	jdff dff_A_gVE3prvY1_0(.dout(w_dff_A_fVXq8srf3_0),.din(w_dff_A_gVE3prvY1_0),.clk(gclk));
	jdff dff_A_fVXq8srf3_0(.dout(w_dff_A_6ZPVnYmI2_0),.din(w_dff_A_fVXq8srf3_0),.clk(gclk));
	jdff dff_A_6ZPVnYmI2_0(.dout(w_dff_A_wpIIYxmW6_0),.din(w_dff_A_6ZPVnYmI2_0),.clk(gclk));
	jdff dff_A_wpIIYxmW6_0(.dout(w_dff_A_IJVHL4aj9_0),.din(w_dff_A_wpIIYxmW6_0),.clk(gclk));
	jdff dff_A_IJVHL4aj9_0(.dout(w_dff_A_2xVWeuRV3_0),.din(w_dff_A_IJVHL4aj9_0),.clk(gclk));
	jdff dff_A_2xVWeuRV3_0(.dout(w_dff_A_W3WCDQQi3_0),.din(w_dff_A_2xVWeuRV3_0),.clk(gclk));
	jdff dff_A_W3WCDQQi3_0(.dout(w_dff_A_A7eHw9W44_0),.din(w_dff_A_W3WCDQQi3_0),.clk(gclk));
	jdff dff_A_A7eHw9W44_0(.dout(w_dff_A_pgrOyBBg0_0),.din(w_dff_A_A7eHw9W44_0),.clk(gclk));
	jdff dff_A_pgrOyBBg0_0(.dout(w_dff_A_DmqY5Xux5_0),.din(w_dff_A_pgrOyBBg0_0),.clk(gclk));
	jdff dff_A_DmqY5Xux5_0(.dout(G1901gat),.din(w_dff_A_DmqY5Xux5_0),.clk(gclk));
	jdff dff_A_Q4wViHZO3_2(.dout(w_dff_A_UKGyNndE4_0),.din(w_dff_A_Q4wViHZO3_2),.clk(gclk));
	jdff dff_A_UKGyNndE4_0(.dout(w_dff_A_qUeEvSGB0_0),.din(w_dff_A_UKGyNndE4_0),.clk(gclk));
	jdff dff_A_qUeEvSGB0_0(.dout(w_dff_A_uUFbC5Eb7_0),.din(w_dff_A_qUeEvSGB0_0),.clk(gclk));
	jdff dff_A_uUFbC5Eb7_0(.dout(w_dff_A_ABV271t69_0),.din(w_dff_A_uUFbC5Eb7_0),.clk(gclk));
	jdff dff_A_ABV271t69_0(.dout(w_dff_A_LhK1w2Fz8_0),.din(w_dff_A_ABV271t69_0),.clk(gclk));
	jdff dff_A_LhK1w2Fz8_0(.dout(w_dff_A_0xGoPeYp4_0),.din(w_dff_A_LhK1w2Fz8_0),.clk(gclk));
	jdff dff_A_0xGoPeYp4_0(.dout(w_dff_A_LbJY9ZJz3_0),.din(w_dff_A_0xGoPeYp4_0),.clk(gclk));
	jdff dff_A_LbJY9ZJz3_0(.dout(w_dff_A_rO1PLAT97_0),.din(w_dff_A_LbJY9ZJz3_0),.clk(gclk));
	jdff dff_A_rO1PLAT97_0(.dout(w_dff_A_Rn1PcijY6_0),.din(w_dff_A_rO1PLAT97_0),.clk(gclk));
	jdff dff_A_Rn1PcijY6_0(.dout(w_dff_A_VbOZqn9n0_0),.din(w_dff_A_Rn1PcijY6_0),.clk(gclk));
	jdff dff_A_VbOZqn9n0_0(.dout(w_dff_A_Kqcb5LSI4_0),.din(w_dff_A_VbOZqn9n0_0),.clk(gclk));
	jdff dff_A_Kqcb5LSI4_0(.dout(w_dff_A_IE7xaUEc8_0),.din(w_dff_A_Kqcb5LSI4_0),.clk(gclk));
	jdff dff_A_IE7xaUEc8_0(.dout(w_dff_A_QsSa10gD7_0),.din(w_dff_A_IE7xaUEc8_0),.clk(gclk));
	jdff dff_A_QsSa10gD7_0(.dout(w_dff_A_CemuLbpo5_0),.din(w_dff_A_QsSa10gD7_0),.clk(gclk));
	jdff dff_A_CemuLbpo5_0(.dout(w_dff_A_cYpjudqf8_0),.din(w_dff_A_CemuLbpo5_0),.clk(gclk));
	jdff dff_A_cYpjudqf8_0(.dout(w_dff_A_uS62HLbT8_0),.din(w_dff_A_cYpjudqf8_0),.clk(gclk));
	jdff dff_A_uS62HLbT8_0(.dout(w_dff_A_aAITNGHM8_0),.din(w_dff_A_uS62HLbT8_0),.clk(gclk));
	jdff dff_A_aAITNGHM8_0(.dout(w_dff_A_c7WM03iH2_0),.din(w_dff_A_aAITNGHM8_0),.clk(gclk));
	jdff dff_A_c7WM03iH2_0(.dout(w_dff_A_VMVN8ZTE0_0),.din(w_dff_A_c7WM03iH2_0),.clk(gclk));
	jdff dff_A_VMVN8ZTE0_0(.dout(w_dff_A_edAnMSk69_0),.din(w_dff_A_VMVN8ZTE0_0),.clk(gclk));
	jdff dff_A_edAnMSk69_0(.dout(w_dff_A_5bGqQTTI1_0),.din(w_dff_A_edAnMSk69_0),.clk(gclk));
	jdff dff_A_5bGqQTTI1_0(.dout(w_dff_A_qxJQYNKX9_0),.din(w_dff_A_5bGqQTTI1_0),.clk(gclk));
	jdff dff_A_qxJQYNKX9_0(.dout(w_dff_A_zqH6VjWv6_0),.din(w_dff_A_qxJQYNKX9_0),.clk(gclk));
	jdff dff_A_zqH6VjWv6_0(.dout(w_dff_A_fFlxY9z75_0),.din(w_dff_A_zqH6VjWv6_0),.clk(gclk));
	jdff dff_A_fFlxY9z75_0(.dout(w_dff_A_lVbwfm9p1_0),.din(w_dff_A_fFlxY9z75_0),.clk(gclk));
	jdff dff_A_lVbwfm9p1_0(.dout(w_dff_A_wIgw8zl50_0),.din(w_dff_A_lVbwfm9p1_0),.clk(gclk));
	jdff dff_A_wIgw8zl50_0(.dout(w_dff_A_VyzX67HB0_0),.din(w_dff_A_wIgw8zl50_0),.clk(gclk));
	jdff dff_A_VyzX67HB0_0(.dout(w_dff_A_YZXJXWSo8_0),.din(w_dff_A_VyzX67HB0_0),.clk(gclk));
	jdff dff_A_YZXJXWSo8_0(.dout(w_dff_A_oPgPigwE1_0),.din(w_dff_A_YZXJXWSo8_0),.clk(gclk));
	jdff dff_A_oPgPigwE1_0(.dout(w_dff_A_l47orzlV2_0),.din(w_dff_A_oPgPigwE1_0),.clk(gclk));
	jdff dff_A_l47orzlV2_0(.dout(w_dff_A_CTRyvGVw5_0),.din(w_dff_A_l47orzlV2_0),.clk(gclk));
	jdff dff_A_CTRyvGVw5_0(.dout(w_dff_A_wy5wa6GW2_0),.din(w_dff_A_CTRyvGVw5_0),.clk(gclk));
	jdff dff_A_wy5wa6GW2_0(.dout(w_dff_A_FJ4FBgg43_0),.din(w_dff_A_wy5wa6GW2_0),.clk(gclk));
	jdff dff_A_FJ4FBgg43_0(.dout(w_dff_A_wWjU7aGC3_0),.din(w_dff_A_FJ4FBgg43_0),.clk(gclk));
	jdff dff_A_wWjU7aGC3_0(.dout(w_dff_A_pnMt5kN98_0),.din(w_dff_A_wWjU7aGC3_0),.clk(gclk));
	jdff dff_A_pnMt5kN98_0(.dout(w_dff_A_Z0KSpMFG3_0),.din(w_dff_A_pnMt5kN98_0),.clk(gclk));
	jdff dff_A_Z0KSpMFG3_0(.dout(w_dff_A_k9nttZJ53_0),.din(w_dff_A_Z0KSpMFG3_0),.clk(gclk));
	jdff dff_A_k9nttZJ53_0(.dout(w_dff_A_8oN7L5TL1_0),.din(w_dff_A_k9nttZJ53_0),.clk(gclk));
	jdff dff_A_8oN7L5TL1_0(.dout(w_dff_A_KQvu6Vn18_0),.din(w_dff_A_8oN7L5TL1_0),.clk(gclk));
	jdff dff_A_KQvu6Vn18_0(.dout(w_dff_A_mO4b9Xv36_0),.din(w_dff_A_KQvu6Vn18_0),.clk(gclk));
	jdff dff_A_mO4b9Xv36_0(.dout(w_dff_A_Gqpo25ko8_0),.din(w_dff_A_mO4b9Xv36_0),.clk(gclk));
	jdff dff_A_Gqpo25ko8_0(.dout(w_dff_A_OiJChVz76_0),.din(w_dff_A_Gqpo25ko8_0),.clk(gclk));
	jdff dff_A_OiJChVz76_0(.dout(w_dff_A_0oUw4awM1_0),.din(w_dff_A_OiJChVz76_0),.clk(gclk));
	jdff dff_A_0oUw4awM1_0(.dout(w_dff_A_BUIBv3MN7_0),.din(w_dff_A_0oUw4awM1_0),.clk(gclk));
	jdff dff_A_BUIBv3MN7_0(.dout(w_dff_A_510i0Ffj1_0),.din(w_dff_A_BUIBv3MN7_0),.clk(gclk));
	jdff dff_A_510i0Ffj1_0(.dout(w_dff_A_63jS389e1_0),.din(w_dff_A_510i0Ffj1_0),.clk(gclk));
	jdff dff_A_63jS389e1_0(.dout(w_dff_A_jK0spGO02_0),.din(w_dff_A_63jS389e1_0),.clk(gclk));
	jdff dff_A_jK0spGO02_0(.dout(w_dff_A_PylGZhxj8_0),.din(w_dff_A_jK0spGO02_0),.clk(gclk));
	jdff dff_A_PylGZhxj8_0(.dout(w_dff_A_OLtjmGcU0_0),.din(w_dff_A_PylGZhxj8_0),.clk(gclk));
	jdff dff_A_OLtjmGcU0_0(.dout(w_dff_A_wCqrIRxR5_0),.din(w_dff_A_OLtjmGcU0_0),.clk(gclk));
	jdff dff_A_wCqrIRxR5_0(.dout(w_dff_A_ByPe0qEa0_0),.din(w_dff_A_wCqrIRxR5_0),.clk(gclk));
	jdff dff_A_ByPe0qEa0_0(.dout(w_dff_A_NzPsVdYV3_0),.din(w_dff_A_ByPe0qEa0_0),.clk(gclk));
	jdff dff_A_NzPsVdYV3_0(.dout(w_dff_A_Ld4GxZ712_0),.din(w_dff_A_NzPsVdYV3_0),.clk(gclk));
	jdff dff_A_Ld4GxZ712_0(.dout(w_dff_A_Jio3chGL5_0),.din(w_dff_A_Ld4GxZ712_0),.clk(gclk));
	jdff dff_A_Jio3chGL5_0(.dout(w_dff_A_Evu8NZnU2_0),.din(w_dff_A_Jio3chGL5_0),.clk(gclk));
	jdff dff_A_Evu8NZnU2_0(.dout(w_dff_A_FnrptbQf6_0),.din(w_dff_A_Evu8NZnU2_0),.clk(gclk));
	jdff dff_A_FnrptbQf6_0(.dout(w_dff_A_GcCGrIZl5_0),.din(w_dff_A_FnrptbQf6_0),.clk(gclk));
	jdff dff_A_GcCGrIZl5_0(.dout(w_dff_A_jZ55oJcH8_0),.din(w_dff_A_GcCGrIZl5_0),.clk(gclk));
	jdff dff_A_jZ55oJcH8_0(.dout(w_dff_A_PyPE5ikt1_0),.din(w_dff_A_jZ55oJcH8_0),.clk(gclk));
	jdff dff_A_PyPE5ikt1_0(.dout(w_dff_A_E5PSy3W04_0),.din(w_dff_A_PyPE5ikt1_0),.clk(gclk));
	jdff dff_A_E5PSy3W04_0(.dout(w_dff_A_bm2wDxTQ4_0),.din(w_dff_A_E5PSy3W04_0),.clk(gclk));
	jdff dff_A_bm2wDxTQ4_0(.dout(w_dff_A_BK8ocyvE5_0),.din(w_dff_A_bm2wDxTQ4_0),.clk(gclk));
	jdff dff_A_BK8ocyvE5_0(.dout(w_dff_A_gJzrV2Jq6_0),.din(w_dff_A_BK8ocyvE5_0),.clk(gclk));
	jdff dff_A_gJzrV2Jq6_0(.dout(w_dff_A_2eqOwn7e3_0),.din(w_dff_A_gJzrV2Jq6_0),.clk(gclk));
	jdff dff_A_2eqOwn7e3_0(.dout(w_dff_A_0zBuhWTA2_0),.din(w_dff_A_2eqOwn7e3_0),.clk(gclk));
	jdff dff_A_0zBuhWTA2_0(.dout(G2223gat),.din(w_dff_A_0zBuhWTA2_0),.clk(gclk));
	jdff dff_A_b8H84EUd8_2(.dout(w_dff_A_TfOUa18I0_0),.din(w_dff_A_b8H84EUd8_2),.clk(gclk));
	jdff dff_A_TfOUa18I0_0(.dout(w_dff_A_kOYBWUmp5_0),.din(w_dff_A_TfOUa18I0_0),.clk(gclk));
	jdff dff_A_kOYBWUmp5_0(.dout(w_dff_A_OsZUU0qz7_0),.din(w_dff_A_kOYBWUmp5_0),.clk(gclk));
	jdff dff_A_OsZUU0qz7_0(.dout(w_dff_A_EnPSnzTH3_0),.din(w_dff_A_OsZUU0qz7_0),.clk(gclk));
	jdff dff_A_EnPSnzTH3_0(.dout(w_dff_A_p5HfxFzY9_0),.din(w_dff_A_EnPSnzTH3_0),.clk(gclk));
	jdff dff_A_p5HfxFzY9_0(.dout(w_dff_A_R6DcDzhx9_0),.din(w_dff_A_p5HfxFzY9_0),.clk(gclk));
	jdff dff_A_R6DcDzhx9_0(.dout(w_dff_A_TBEkWVCz0_0),.din(w_dff_A_R6DcDzhx9_0),.clk(gclk));
	jdff dff_A_TBEkWVCz0_0(.dout(w_dff_A_mjo7B4Fa6_0),.din(w_dff_A_TBEkWVCz0_0),.clk(gclk));
	jdff dff_A_mjo7B4Fa6_0(.dout(w_dff_A_DOHeVL7p1_0),.din(w_dff_A_mjo7B4Fa6_0),.clk(gclk));
	jdff dff_A_DOHeVL7p1_0(.dout(w_dff_A_jTxufXdv3_0),.din(w_dff_A_DOHeVL7p1_0),.clk(gclk));
	jdff dff_A_jTxufXdv3_0(.dout(w_dff_A_PrAnHZNC9_0),.din(w_dff_A_jTxufXdv3_0),.clk(gclk));
	jdff dff_A_PrAnHZNC9_0(.dout(w_dff_A_hgyb57m38_0),.din(w_dff_A_PrAnHZNC9_0),.clk(gclk));
	jdff dff_A_hgyb57m38_0(.dout(w_dff_A_1yimvYdx1_0),.din(w_dff_A_hgyb57m38_0),.clk(gclk));
	jdff dff_A_1yimvYdx1_0(.dout(w_dff_A_pq0AN4Bz7_0),.din(w_dff_A_1yimvYdx1_0),.clk(gclk));
	jdff dff_A_pq0AN4Bz7_0(.dout(w_dff_A_S5TbOQHk3_0),.din(w_dff_A_pq0AN4Bz7_0),.clk(gclk));
	jdff dff_A_S5TbOQHk3_0(.dout(w_dff_A_tE7M3Alx8_0),.din(w_dff_A_S5TbOQHk3_0),.clk(gclk));
	jdff dff_A_tE7M3Alx8_0(.dout(w_dff_A_a9cnZ2ms4_0),.din(w_dff_A_tE7M3Alx8_0),.clk(gclk));
	jdff dff_A_a9cnZ2ms4_0(.dout(w_dff_A_H1HuJkNV0_0),.din(w_dff_A_a9cnZ2ms4_0),.clk(gclk));
	jdff dff_A_H1HuJkNV0_0(.dout(w_dff_A_cmwQA2G10_0),.din(w_dff_A_H1HuJkNV0_0),.clk(gclk));
	jdff dff_A_cmwQA2G10_0(.dout(w_dff_A_AjzvMHCx6_0),.din(w_dff_A_cmwQA2G10_0),.clk(gclk));
	jdff dff_A_AjzvMHCx6_0(.dout(w_dff_A_EbAumOFk7_0),.din(w_dff_A_AjzvMHCx6_0),.clk(gclk));
	jdff dff_A_EbAumOFk7_0(.dout(w_dff_A_ysdZlWv88_0),.din(w_dff_A_EbAumOFk7_0),.clk(gclk));
	jdff dff_A_ysdZlWv88_0(.dout(w_dff_A_Bbez2tlE5_0),.din(w_dff_A_ysdZlWv88_0),.clk(gclk));
	jdff dff_A_Bbez2tlE5_0(.dout(w_dff_A_6XLO7Fw82_0),.din(w_dff_A_Bbez2tlE5_0),.clk(gclk));
	jdff dff_A_6XLO7Fw82_0(.dout(w_dff_A_hKh6lD7L9_0),.din(w_dff_A_6XLO7Fw82_0),.clk(gclk));
	jdff dff_A_hKh6lD7L9_0(.dout(w_dff_A_cGkyTB5W4_0),.din(w_dff_A_hKh6lD7L9_0),.clk(gclk));
	jdff dff_A_cGkyTB5W4_0(.dout(w_dff_A_fMIrfBBI8_0),.din(w_dff_A_cGkyTB5W4_0),.clk(gclk));
	jdff dff_A_fMIrfBBI8_0(.dout(w_dff_A_JYUNmNKE9_0),.din(w_dff_A_fMIrfBBI8_0),.clk(gclk));
	jdff dff_A_JYUNmNKE9_0(.dout(w_dff_A_CvHAEX0k4_0),.din(w_dff_A_JYUNmNKE9_0),.clk(gclk));
	jdff dff_A_CvHAEX0k4_0(.dout(w_dff_A_Gv4SL5FF2_0),.din(w_dff_A_CvHAEX0k4_0),.clk(gclk));
	jdff dff_A_Gv4SL5FF2_0(.dout(w_dff_A_zfun9FGi9_0),.din(w_dff_A_Gv4SL5FF2_0),.clk(gclk));
	jdff dff_A_zfun9FGi9_0(.dout(w_dff_A_9NU0YyFk1_0),.din(w_dff_A_zfun9FGi9_0),.clk(gclk));
	jdff dff_A_9NU0YyFk1_0(.dout(w_dff_A_G2j0uwhU0_0),.din(w_dff_A_9NU0YyFk1_0),.clk(gclk));
	jdff dff_A_G2j0uwhU0_0(.dout(w_dff_A_PdFBEcAu9_0),.din(w_dff_A_G2j0uwhU0_0),.clk(gclk));
	jdff dff_A_PdFBEcAu9_0(.dout(w_dff_A_0WdiCdjO4_0),.din(w_dff_A_PdFBEcAu9_0),.clk(gclk));
	jdff dff_A_0WdiCdjO4_0(.dout(w_dff_A_HCUgIoKA0_0),.din(w_dff_A_0WdiCdjO4_0),.clk(gclk));
	jdff dff_A_HCUgIoKA0_0(.dout(w_dff_A_rfFoVhDr4_0),.din(w_dff_A_HCUgIoKA0_0),.clk(gclk));
	jdff dff_A_rfFoVhDr4_0(.dout(w_dff_A_hyB6LONs5_0),.din(w_dff_A_rfFoVhDr4_0),.clk(gclk));
	jdff dff_A_hyB6LONs5_0(.dout(w_dff_A_ltjay0QD0_0),.din(w_dff_A_hyB6LONs5_0),.clk(gclk));
	jdff dff_A_ltjay0QD0_0(.dout(w_dff_A_LvphP0BZ5_0),.din(w_dff_A_ltjay0QD0_0),.clk(gclk));
	jdff dff_A_LvphP0BZ5_0(.dout(w_dff_A_J2kPCyek1_0),.din(w_dff_A_LvphP0BZ5_0),.clk(gclk));
	jdff dff_A_J2kPCyek1_0(.dout(w_dff_A_yTJRrLgV9_0),.din(w_dff_A_J2kPCyek1_0),.clk(gclk));
	jdff dff_A_yTJRrLgV9_0(.dout(w_dff_A_qu3U2GnF7_0),.din(w_dff_A_yTJRrLgV9_0),.clk(gclk));
	jdff dff_A_qu3U2GnF7_0(.dout(w_dff_A_G2UL7Bd80_0),.din(w_dff_A_qu3U2GnF7_0),.clk(gclk));
	jdff dff_A_G2UL7Bd80_0(.dout(w_dff_A_wNcBxNYb8_0),.din(w_dff_A_G2UL7Bd80_0),.clk(gclk));
	jdff dff_A_wNcBxNYb8_0(.dout(w_dff_A_bDySrMfT6_0),.din(w_dff_A_wNcBxNYb8_0),.clk(gclk));
	jdff dff_A_bDySrMfT6_0(.dout(w_dff_A_d8Rc8Dj91_0),.din(w_dff_A_bDySrMfT6_0),.clk(gclk));
	jdff dff_A_d8Rc8Dj91_0(.dout(w_dff_A_PP7L8aRr7_0),.din(w_dff_A_d8Rc8Dj91_0),.clk(gclk));
	jdff dff_A_PP7L8aRr7_0(.dout(w_dff_A_RHkARyY51_0),.din(w_dff_A_PP7L8aRr7_0),.clk(gclk));
	jdff dff_A_RHkARyY51_0(.dout(w_dff_A_oh4qkzh30_0),.din(w_dff_A_RHkARyY51_0),.clk(gclk));
	jdff dff_A_oh4qkzh30_0(.dout(w_dff_A_vb6UVT9T2_0),.din(w_dff_A_oh4qkzh30_0),.clk(gclk));
	jdff dff_A_vb6UVT9T2_0(.dout(w_dff_A_a6ahhC4d8_0),.din(w_dff_A_vb6UVT9T2_0),.clk(gclk));
	jdff dff_A_a6ahhC4d8_0(.dout(w_dff_A_LgnjWNqr0_0),.din(w_dff_A_a6ahhC4d8_0),.clk(gclk));
	jdff dff_A_LgnjWNqr0_0(.dout(w_dff_A_b9I6DdCh8_0),.din(w_dff_A_LgnjWNqr0_0),.clk(gclk));
	jdff dff_A_b9I6DdCh8_0(.dout(w_dff_A_v8BwIdj35_0),.din(w_dff_A_b9I6DdCh8_0),.clk(gclk));
	jdff dff_A_v8BwIdj35_0(.dout(w_dff_A_tGAEwy2j6_0),.din(w_dff_A_v8BwIdj35_0),.clk(gclk));
	jdff dff_A_tGAEwy2j6_0(.dout(w_dff_A_NUWJri9V5_0),.din(w_dff_A_tGAEwy2j6_0),.clk(gclk));
	jdff dff_A_NUWJri9V5_0(.dout(w_dff_A_zIXL6pBc1_0),.din(w_dff_A_NUWJri9V5_0),.clk(gclk));
	jdff dff_A_zIXL6pBc1_0(.dout(w_dff_A_204SQmAl0_0),.din(w_dff_A_zIXL6pBc1_0),.clk(gclk));
	jdff dff_A_204SQmAl0_0(.dout(w_dff_A_P1U7JFDu8_0),.din(w_dff_A_204SQmAl0_0),.clk(gclk));
	jdff dff_A_P1U7JFDu8_0(.dout(w_dff_A_GOGGinFG4_0),.din(w_dff_A_P1U7JFDu8_0),.clk(gclk));
	jdff dff_A_GOGGinFG4_0(.dout(w_dff_A_sWpZw6D99_0),.din(w_dff_A_GOGGinFG4_0),.clk(gclk));
	jdff dff_A_sWpZw6D99_0(.dout(G2548gat),.din(w_dff_A_sWpZw6D99_0),.clk(gclk));
	jdff dff_A_8Uk1cOcq0_2(.dout(w_dff_A_ZNdjjxTJ1_0),.din(w_dff_A_8Uk1cOcq0_2),.clk(gclk));
	jdff dff_A_ZNdjjxTJ1_0(.dout(w_dff_A_GtvGFjjC7_0),.din(w_dff_A_ZNdjjxTJ1_0),.clk(gclk));
	jdff dff_A_GtvGFjjC7_0(.dout(w_dff_A_ghWEGvCc2_0),.din(w_dff_A_GtvGFjjC7_0),.clk(gclk));
	jdff dff_A_ghWEGvCc2_0(.dout(w_dff_A_FLSV3KvY3_0),.din(w_dff_A_ghWEGvCc2_0),.clk(gclk));
	jdff dff_A_FLSV3KvY3_0(.dout(w_dff_A_Bb4iMqSI9_0),.din(w_dff_A_FLSV3KvY3_0),.clk(gclk));
	jdff dff_A_Bb4iMqSI9_0(.dout(w_dff_A_5BoyWzza5_0),.din(w_dff_A_Bb4iMqSI9_0),.clk(gclk));
	jdff dff_A_5BoyWzza5_0(.dout(w_dff_A_Hu7weckT3_0),.din(w_dff_A_5BoyWzza5_0),.clk(gclk));
	jdff dff_A_Hu7weckT3_0(.dout(w_dff_A_nPGEJE8D5_0),.din(w_dff_A_Hu7weckT3_0),.clk(gclk));
	jdff dff_A_nPGEJE8D5_0(.dout(w_dff_A_2lmtdOzz6_0),.din(w_dff_A_nPGEJE8D5_0),.clk(gclk));
	jdff dff_A_2lmtdOzz6_0(.dout(w_dff_A_1xOC7Avq8_0),.din(w_dff_A_2lmtdOzz6_0),.clk(gclk));
	jdff dff_A_1xOC7Avq8_0(.dout(w_dff_A_i7Sdlbpb2_0),.din(w_dff_A_1xOC7Avq8_0),.clk(gclk));
	jdff dff_A_i7Sdlbpb2_0(.dout(w_dff_A_HSvDHkDo9_0),.din(w_dff_A_i7Sdlbpb2_0),.clk(gclk));
	jdff dff_A_HSvDHkDo9_0(.dout(w_dff_A_k7SyHhOQ6_0),.din(w_dff_A_HSvDHkDo9_0),.clk(gclk));
	jdff dff_A_k7SyHhOQ6_0(.dout(w_dff_A_kJpWwXy29_0),.din(w_dff_A_k7SyHhOQ6_0),.clk(gclk));
	jdff dff_A_kJpWwXy29_0(.dout(w_dff_A_UWTEAV8C2_0),.din(w_dff_A_kJpWwXy29_0),.clk(gclk));
	jdff dff_A_UWTEAV8C2_0(.dout(w_dff_A_6gvOMjes6_0),.din(w_dff_A_UWTEAV8C2_0),.clk(gclk));
	jdff dff_A_6gvOMjes6_0(.dout(w_dff_A_de6d6Jpu2_0),.din(w_dff_A_6gvOMjes6_0),.clk(gclk));
	jdff dff_A_de6d6Jpu2_0(.dout(w_dff_A_d7DrD2qF3_0),.din(w_dff_A_de6d6Jpu2_0),.clk(gclk));
	jdff dff_A_d7DrD2qF3_0(.dout(w_dff_A_VpcXFAxc1_0),.din(w_dff_A_d7DrD2qF3_0),.clk(gclk));
	jdff dff_A_VpcXFAxc1_0(.dout(w_dff_A_lzvGUfaV5_0),.din(w_dff_A_VpcXFAxc1_0),.clk(gclk));
	jdff dff_A_lzvGUfaV5_0(.dout(w_dff_A_0DNugwJW1_0),.din(w_dff_A_lzvGUfaV5_0),.clk(gclk));
	jdff dff_A_0DNugwJW1_0(.dout(w_dff_A_LAuOrVh08_0),.din(w_dff_A_0DNugwJW1_0),.clk(gclk));
	jdff dff_A_LAuOrVh08_0(.dout(w_dff_A_of0dPu3C3_0),.din(w_dff_A_LAuOrVh08_0),.clk(gclk));
	jdff dff_A_of0dPu3C3_0(.dout(w_dff_A_tJKfD2rm2_0),.din(w_dff_A_of0dPu3C3_0),.clk(gclk));
	jdff dff_A_tJKfD2rm2_0(.dout(w_dff_A_V36l25ax3_0),.din(w_dff_A_tJKfD2rm2_0),.clk(gclk));
	jdff dff_A_V36l25ax3_0(.dout(w_dff_A_anlxOSS95_0),.din(w_dff_A_V36l25ax3_0),.clk(gclk));
	jdff dff_A_anlxOSS95_0(.dout(w_dff_A_fF1kcHot1_0),.din(w_dff_A_anlxOSS95_0),.clk(gclk));
	jdff dff_A_fF1kcHot1_0(.dout(w_dff_A_CzeJ0s053_0),.din(w_dff_A_fF1kcHot1_0),.clk(gclk));
	jdff dff_A_CzeJ0s053_0(.dout(w_dff_A_31htIorp6_0),.din(w_dff_A_CzeJ0s053_0),.clk(gclk));
	jdff dff_A_31htIorp6_0(.dout(w_dff_A_Ie903EKS2_0),.din(w_dff_A_31htIorp6_0),.clk(gclk));
	jdff dff_A_Ie903EKS2_0(.dout(w_dff_A_vyUY25xC3_0),.din(w_dff_A_Ie903EKS2_0),.clk(gclk));
	jdff dff_A_vyUY25xC3_0(.dout(w_dff_A_JwsDxDiU1_0),.din(w_dff_A_vyUY25xC3_0),.clk(gclk));
	jdff dff_A_JwsDxDiU1_0(.dout(w_dff_A_xUjGRNrk5_0),.din(w_dff_A_JwsDxDiU1_0),.clk(gclk));
	jdff dff_A_xUjGRNrk5_0(.dout(w_dff_A_FjjpXrAd0_0),.din(w_dff_A_xUjGRNrk5_0),.clk(gclk));
	jdff dff_A_FjjpXrAd0_0(.dout(w_dff_A_zS849JfP3_0),.din(w_dff_A_FjjpXrAd0_0),.clk(gclk));
	jdff dff_A_zS849JfP3_0(.dout(w_dff_A_2A6zkH867_0),.din(w_dff_A_zS849JfP3_0),.clk(gclk));
	jdff dff_A_2A6zkH867_0(.dout(w_dff_A_m2Xk6hNZ6_0),.din(w_dff_A_2A6zkH867_0),.clk(gclk));
	jdff dff_A_m2Xk6hNZ6_0(.dout(w_dff_A_FRFGGGmw2_0),.din(w_dff_A_m2Xk6hNZ6_0),.clk(gclk));
	jdff dff_A_FRFGGGmw2_0(.dout(w_dff_A_t040DJOD7_0),.din(w_dff_A_FRFGGGmw2_0),.clk(gclk));
	jdff dff_A_t040DJOD7_0(.dout(w_dff_A_luahPP6e8_0),.din(w_dff_A_t040DJOD7_0),.clk(gclk));
	jdff dff_A_luahPP6e8_0(.dout(w_dff_A_jT8CVY1H6_0),.din(w_dff_A_luahPP6e8_0),.clk(gclk));
	jdff dff_A_jT8CVY1H6_0(.dout(w_dff_A_hDcxsap11_0),.din(w_dff_A_jT8CVY1H6_0),.clk(gclk));
	jdff dff_A_hDcxsap11_0(.dout(w_dff_A_TdIJKXMH6_0),.din(w_dff_A_hDcxsap11_0),.clk(gclk));
	jdff dff_A_TdIJKXMH6_0(.dout(w_dff_A_CEm9jKnO4_0),.din(w_dff_A_TdIJKXMH6_0),.clk(gclk));
	jdff dff_A_CEm9jKnO4_0(.dout(w_dff_A_2zrtAXyg6_0),.din(w_dff_A_CEm9jKnO4_0),.clk(gclk));
	jdff dff_A_2zrtAXyg6_0(.dout(w_dff_A_If2MmPWx1_0),.din(w_dff_A_2zrtAXyg6_0),.clk(gclk));
	jdff dff_A_If2MmPWx1_0(.dout(w_dff_A_DKdcllYN9_0),.din(w_dff_A_If2MmPWx1_0),.clk(gclk));
	jdff dff_A_DKdcllYN9_0(.dout(w_dff_A_Ikoz8JaA7_0),.din(w_dff_A_DKdcllYN9_0),.clk(gclk));
	jdff dff_A_Ikoz8JaA7_0(.dout(w_dff_A_Qh5t4D9u8_0),.din(w_dff_A_Ikoz8JaA7_0),.clk(gclk));
	jdff dff_A_Qh5t4D9u8_0(.dout(w_dff_A_ICyzaWu23_0),.din(w_dff_A_Qh5t4D9u8_0),.clk(gclk));
	jdff dff_A_ICyzaWu23_0(.dout(w_dff_A_F0fqGvBY9_0),.din(w_dff_A_ICyzaWu23_0),.clk(gclk));
	jdff dff_A_F0fqGvBY9_0(.dout(w_dff_A_rS0FBamH3_0),.din(w_dff_A_F0fqGvBY9_0),.clk(gclk));
	jdff dff_A_rS0FBamH3_0(.dout(w_dff_A_JGJ9vYXy5_0),.din(w_dff_A_rS0FBamH3_0),.clk(gclk));
	jdff dff_A_JGJ9vYXy5_0(.dout(w_dff_A_uIBqQaBQ8_0),.din(w_dff_A_JGJ9vYXy5_0),.clk(gclk));
	jdff dff_A_uIBqQaBQ8_0(.dout(w_dff_A_Uqvkm0sU2_0),.din(w_dff_A_uIBqQaBQ8_0),.clk(gclk));
	jdff dff_A_Uqvkm0sU2_0(.dout(w_dff_A_kKTB73Rd6_0),.din(w_dff_A_Uqvkm0sU2_0),.clk(gclk));
	jdff dff_A_kKTB73Rd6_0(.dout(w_dff_A_wFRSiLAG9_0),.din(w_dff_A_kKTB73Rd6_0),.clk(gclk));
	jdff dff_A_wFRSiLAG9_0(.dout(w_dff_A_DBujhYrI0_0),.din(w_dff_A_wFRSiLAG9_0),.clk(gclk));
	jdff dff_A_DBujhYrI0_0(.dout(w_dff_A_8D78vdMV3_0),.din(w_dff_A_DBujhYrI0_0),.clk(gclk));
	jdff dff_A_8D78vdMV3_0(.dout(G2877gat),.din(w_dff_A_8D78vdMV3_0),.clk(gclk));
	jdff dff_A_5EPJFSK63_2(.dout(w_dff_A_DOExoYER6_0),.din(w_dff_A_5EPJFSK63_2),.clk(gclk));
	jdff dff_A_DOExoYER6_0(.dout(w_dff_A_tFuCoYJZ8_0),.din(w_dff_A_DOExoYER6_0),.clk(gclk));
	jdff dff_A_tFuCoYJZ8_0(.dout(w_dff_A_znDc7feD8_0),.din(w_dff_A_tFuCoYJZ8_0),.clk(gclk));
	jdff dff_A_znDc7feD8_0(.dout(w_dff_A_hf6uyi5n3_0),.din(w_dff_A_znDc7feD8_0),.clk(gclk));
	jdff dff_A_hf6uyi5n3_0(.dout(w_dff_A_EhYx15uM5_0),.din(w_dff_A_hf6uyi5n3_0),.clk(gclk));
	jdff dff_A_EhYx15uM5_0(.dout(w_dff_A_yctUxyfm9_0),.din(w_dff_A_EhYx15uM5_0),.clk(gclk));
	jdff dff_A_yctUxyfm9_0(.dout(w_dff_A_qAeChpos2_0),.din(w_dff_A_yctUxyfm9_0),.clk(gclk));
	jdff dff_A_qAeChpos2_0(.dout(w_dff_A_7G5BdfF69_0),.din(w_dff_A_qAeChpos2_0),.clk(gclk));
	jdff dff_A_7G5BdfF69_0(.dout(w_dff_A_hkBNqklD3_0),.din(w_dff_A_7G5BdfF69_0),.clk(gclk));
	jdff dff_A_hkBNqklD3_0(.dout(w_dff_A_Ca6reP3d4_0),.din(w_dff_A_hkBNqklD3_0),.clk(gclk));
	jdff dff_A_Ca6reP3d4_0(.dout(w_dff_A_ujVpV9dA3_0),.din(w_dff_A_Ca6reP3d4_0),.clk(gclk));
	jdff dff_A_ujVpV9dA3_0(.dout(w_dff_A_PODTHDFB5_0),.din(w_dff_A_ujVpV9dA3_0),.clk(gclk));
	jdff dff_A_PODTHDFB5_0(.dout(w_dff_A_maef2V9b2_0),.din(w_dff_A_PODTHDFB5_0),.clk(gclk));
	jdff dff_A_maef2V9b2_0(.dout(w_dff_A_5RtaVRdA0_0),.din(w_dff_A_maef2V9b2_0),.clk(gclk));
	jdff dff_A_5RtaVRdA0_0(.dout(w_dff_A_GP2sS9ak0_0),.din(w_dff_A_5RtaVRdA0_0),.clk(gclk));
	jdff dff_A_GP2sS9ak0_0(.dout(w_dff_A_htKBQqzB2_0),.din(w_dff_A_GP2sS9ak0_0),.clk(gclk));
	jdff dff_A_htKBQqzB2_0(.dout(w_dff_A_NPTNKuUW0_0),.din(w_dff_A_htKBQqzB2_0),.clk(gclk));
	jdff dff_A_NPTNKuUW0_0(.dout(w_dff_A_bDOonGCq8_0),.din(w_dff_A_NPTNKuUW0_0),.clk(gclk));
	jdff dff_A_bDOonGCq8_0(.dout(w_dff_A_TJbWIYZT1_0),.din(w_dff_A_bDOonGCq8_0),.clk(gclk));
	jdff dff_A_TJbWIYZT1_0(.dout(w_dff_A_CvGGnXvv3_0),.din(w_dff_A_TJbWIYZT1_0),.clk(gclk));
	jdff dff_A_CvGGnXvv3_0(.dout(w_dff_A_cplFvibM7_0),.din(w_dff_A_CvGGnXvv3_0),.clk(gclk));
	jdff dff_A_cplFvibM7_0(.dout(w_dff_A_mUEyJ9456_0),.din(w_dff_A_cplFvibM7_0),.clk(gclk));
	jdff dff_A_mUEyJ9456_0(.dout(w_dff_A_Ntkvz3F21_0),.din(w_dff_A_mUEyJ9456_0),.clk(gclk));
	jdff dff_A_Ntkvz3F21_0(.dout(w_dff_A_XuGkLMtx1_0),.din(w_dff_A_Ntkvz3F21_0),.clk(gclk));
	jdff dff_A_XuGkLMtx1_0(.dout(w_dff_A_c8kEqfk06_0),.din(w_dff_A_XuGkLMtx1_0),.clk(gclk));
	jdff dff_A_c8kEqfk06_0(.dout(w_dff_A_gtTQ0BmB3_0),.din(w_dff_A_c8kEqfk06_0),.clk(gclk));
	jdff dff_A_gtTQ0BmB3_0(.dout(w_dff_A_yud3cl7S4_0),.din(w_dff_A_gtTQ0BmB3_0),.clk(gclk));
	jdff dff_A_yud3cl7S4_0(.dout(w_dff_A_OXLZpy2o2_0),.din(w_dff_A_yud3cl7S4_0),.clk(gclk));
	jdff dff_A_OXLZpy2o2_0(.dout(w_dff_A_XaMmCvE16_0),.din(w_dff_A_OXLZpy2o2_0),.clk(gclk));
	jdff dff_A_XaMmCvE16_0(.dout(w_dff_A_zjPs8UHG2_0),.din(w_dff_A_XaMmCvE16_0),.clk(gclk));
	jdff dff_A_zjPs8UHG2_0(.dout(w_dff_A_9YE8RIk48_0),.din(w_dff_A_zjPs8UHG2_0),.clk(gclk));
	jdff dff_A_9YE8RIk48_0(.dout(w_dff_A_OucV5Ba50_0),.din(w_dff_A_9YE8RIk48_0),.clk(gclk));
	jdff dff_A_OucV5Ba50_0(.dout(w_dff_A_wXqAISRH6_0),.din(w_dff_A_OucV5Ba50_0),.clk(gclk));
	jdff dff_A_wXqAISRH6_0(.dout(w_dff_A_BE9GZZZM2_0),.din(w_dff_A_wXqAISRH6_0),.clk(gclk));
	jdff dff_A_BE9GZZZM2_0(.dout(w_dff_A_MgWkUPIG2_0),.din(w_dff_A_BE9GZZZM2_0),.clk(gclk));
	jdff dff_A_MgWkUPIG2_0(.dout(w_dff_A_BfX6LqHl6_0),.din(w_dff_A_MgWkUPIG2_0),.clk(gclk));
	jdff dff_A_BfX6LqHl6_0(.dout(w_dff_A_XWMywfCp9_0),.din(w_dff_A_BfX6LqHl6_0),.clk(gclk));
	jdff dff_A_XWMywfCp9_0(.dout(w_dff_A_VDjwOVe88_0),.din(w_dff_A_XWMywfCp9_0),.clk(gclk));
	jdff dff_A_VDjwOVe88_0(.dout(w_dff_A_z9SvHDb44_0),.din(w_dff_A_VDjwOVe88_0),.clk(gclk));
	jdff dff_A_z9SvHDb44_0(.dout(w_dff_A_Ivyi9z878_0),.din(w_dff_A_z9SvHDb44_0),.clk(gclk));
	jdff dff_A_Ivyi9z878_0(.dout(w_dff_A_XACCBGIh2_0),.din(w_dff_A_Ivyi9z878_0),.clk(gclk));
	jdff dff_A_XACCBGIh2_0(.dout(w_dff_A_C8moW3nw2_0),.din(w_dff_A_XACCBGIh2_0),.clk(gclk));
	jdff dff_A_C8moW3nw2_0(.dout(w_dff_A_OmSf8ubk7_0),.din(w_dff_A_C8moW3nw2_0),.clk(gclk));
	jdff dff_A_OmSf8ubk7_0(.dout(w_dff_A_0kAqH5D97_0),.din(w_dff_A_OmSf8ubk7_0),.clk(gclk));
	jdff dff_A_0kAqH5D97_0(.dout(w_dff_A_3CnDak9C2_0),.din(w_dff_A_0kAqH5D97_0),.clk(gclk));
	jdff dff_A_3CnDak9C2_0(.dout(w_dff_A_ER9dLIIt3_0),.din(w_dff_A_3CnDak9C2_0),.clk(gclk));
	jdff dff_A_ER9dLIIt3_0(.dout(w_dff_A_BHu30DB33_0),.din(w_dff_A_ER9dLIIt3_0),.clk(gclk));
	jdff dff_A_BHu30DB33_0(.dout(w_dff_A_d3pgP1Ip1_0),.din(w_dff_A_BHu30DB33_0),.clk(gclk));
	jdff dff_A_d3pgP1Ip1_0(.dout(w_dff_A_BWQHLhiv4_0),.din(w_dff_A_d3pgP1Ip1_0),.clk(gclk));
	jdff dff_A_BWQHLhiv4_0(.dout(w_dff_A_FKtdbGcd0_0),.din(w_dff_A_BWQHLhiv4_0),.clk(gclk));
	jdff dff_A_FKtdbGcd0_0(.dout(w_dff_A_R0HwiVEl2_0),.din(w_dff_A_FKtdbGcd0_0),.clk(gclk));
	jdff dff_A_R0HwiVEl2_0(.dout(w_dff_A_lQAtHQA38_0),.din(w_dff_A_R0HwiVEl2_0),.clk(gclk));
	jdff dff_A_lQAtHQA38_0(.dout(w_dff_A_706FWQ9x8_0),.din(w_dff_A_lQAtHQA38_0),.clk(gclk));
	jdff dff_A_706FWQ9x8_0(.dout(w_dff_A_lB78BTCY6_0),.din(w_dff_A_706FWQ9x8_0),.clk(gclk));
	jdff dff_A_lB78BTCY6_0(.dout(w_dff_A_R3LZrqqa6_0),.din(w_dff_A_lB78BTCY6_0),.clk(gclk));
	jdff dff_A_R3LZrqqa6_0(.dout(w_dff_A_HxYS5P9r5_0),.din(w_dff_A_R3LZrqqa6_0),.clk(gclk));
	jdff dff_A_HxYS5P9r5_0(.dout(G3211gat),.din(w_dff_A_HxYS5P9r5_0),.clk(gclk));
	jdff dff_A_zuCOQdnm3_2(.dout(w_dff_A_qOywLTmq5_0),.din(w_dff_A_zuCOQdnm3_2),.clk(gclk));
	jdff dff_A_qOywLTmq5_0(.dout(w_dff_A_obdsjDGW8_0),.din(w_dff_A_qOywLTmq5_0),.clk(gclk));
	jdff dff_A_obdsjDGW8_0(.dout(w_dff_A_xlJxa8Vb2_0),.din(w_dff_A_obdsjDGW8_0),.clk(gclk));
	jdff dff_A_xlJxa8Vb2_0(.dout(w_dff_A_0bgbmw1u7_0),.din(w_dff_A_xlJxa8Vb2_0),.clk(gclk));
	jdff dff_A_0bgbmw1u7_0(.dout(w_dff_A_ILkNZUoq5_0),.din(w_dff_A_0bgbmw1u7_0),.clk(gclk));
	jdff dff_A_ILkNZUoq5_0(.dout(w_dff_A_6eI363v60_0),.din(w_dff_A_ILkNZUoq5_0),.clk(gclk));
	jdff dff_A_6eI363v60_0(.dout(w_dff_A_uA1SrmJJ7_0),.din(w_dff_A_6eI363v60_0),.clk(gclk));
	jdff dff_A_uA1SrmJJ7_0(.dout(w_dff_A_WNXOlrTT4_0),.din(w_dff_A_uA1SrmJJ7_0),.clk(gclk));
	jdff dff_A_WNXOlrTT4_0(.dout(w_dff_A_YSD7njIx0_0),.din(w_dff_A_WNXOlrTT4_0),.clk(gclk));
	jdff dff_A_YSD7njIx0_0(.dout(w_dff_A_Zqxssgrr2_0),.din(w_dff_A_YSD7njIx0_0),.clk(gclk));
	jdff dff_A_Zqxssgrr2_0(.dout(w_dff_A_Akfrz6Km5_0),.din(w_dff_A_Zqxssgrr2_0),.clk(gclk));
	jdff dff_A_Akfrz6Km5_0(.dout(w_dff_A_fKmMWVFy6_0),.din(w_dff_A_Akfrz6Km5_0),.clk(gclk));
	jdff dff_A_fKmMWVFy6_0(.dout(w_dff_A_IweDFsLr9_0),.din(w_dff_A_fKmMWVFy6_0),.clk(gclk));
	jdff dff_A_IweDFsLr9_0(.dout(w_dff_A_zQP5IMQI2_0),.din(w_dff_A_IweDFsLr9_0),.clk(gclk));
	jdff dff_A_zQP5IMQI2_0(.dout(w_dff_A_2lCCdQtA1_0),.din(w_dff_A_zQP5IMQI2_0),.clk(gclk));
	jdff dff_A_2lCCdQtA1_0(.dout(w_dff_A_I5Rk9tDT0_0),.din(w_dff_A_2lCCdQtA1_0),.clk(gclk));
	jdff dff_A_I5Rk9tDT0_0(.dout(w_dff_A_IRbZlG1X4_0),.din(w_dff_A_I5Rk9tDT0_0),.clk(gclk));
	jdff dff_A_IRbZlG1X4_0(.dout(w_dff_A_unJmHk0G7_0),.din(w_dff_A_IRbZlG1X4_0),.clk(gclk));
	jdff dff_A_unJmHk0G7_0(.dout(w_dff_A_1jJQ6CmA6_0),.din(w_dff_A_unJmHk0G7_0),.clk(gclk));
	jdff dff_A_1jJQ6CmA6_0(.dout(w_dff_A_xYVOu8Jh1_0),.din(w_dff_A_1jJQ6CmA6_0),.clk(gclk));
	jdff dff_A_xYVOu8Jh1_0(.dout(w_dff_A_WDrDF0rk5_0),.din(w_dff_A_xYVOu8Jh1_0),.clk(gclk));
	jdff dff_A_WDrDF0rk5_0(.dout(w_dff_A_Edd5FS4Z2_0),.din(w_dff_A_WDrDF0rk5_0),.clk(gclk));
	jdff dff_A_Edd5FS4Z2_0(.dout(w_dff_A_lZxAB5FU0_0),.din(w_dff_A_Edd5FS4Z2_0),.clk(gclk));
	jdff dff_A_lZxAB5FU0_0(.dout(w_dff_A_k8jVv6X26_0),.din(w_dff_A_lZxAB5FU0_0),.clk(gclk));
	jdff dff_A_k8jVv6X26_0(.dout(w_dff_A_8SPu4LWF3_0),.din(w_dff_A_k8jVv6X26_0),.clk(gclk));
	jdff dff_A_8SPu4LWF3_0(.dout(w_dff_A_7K4dkvlQ1_0),.din(w_dff_A_8SPu4LWF3_0),.clk(gclk));
	jdff dff_A_7K4dkvlQ1_0(.dout(w_dff_A_PrJMawVA5_0),.din(w_dff_A_7K4dkvlQ1_0),.clk(gclk));
	jdff dff_A_PrJMawVA5_0(.dout(w_dff_A_FC40UmaC4_0),.din(w_dff_A_PrJMawVA5_0),.clk(gclk));
	jdff dff_A_FC40UmaC4_0(.dout(w_dff_A_RmGkp7WL1_0),.din(w_dff_A_FC40UmaC4_0),.clk(gclk));
	jdff dff_A_RmGkp7WL1_0(.dout(w_dff_A_rEhQd5jb2_0),.din(w_dff_A_RmGkp7WL1_0),.clk(gclk));
	jdff dff_A_rEhQd5jb2_0(.dout(w_dff_A_80r88e0W0_0),.din(w_dff_A_rEhQd5jb2_0),.clk(gclk));
	jdff dff_A_80r88e0W0_0(.dout(w_dff_A_h4QrjZNp1_0),.din(w_dff_A_80r88e0W0_0),.clk(gclk));
	jdff dff_A_h4QrjZNp1_0(.dout(w_dff_A_121wZNT26_0),.din(w_dff_A_h4QrjZNp1_0),.clk(gclk));
	jdff dff_A_121wZNT26_0(.dout(w_dff_A_uU3aGcZC1_0),.din(w_dff_A_121wZNT26_0),.clk(gclk));
	jdff dff_A_uU3aGcZC1_0(.dout(w_dff_A_aGe0Gktb9_0),.din(w_dff_A_uU3aGcZC1_0),.clk(gclk));
	jdff dff_A_aGe0Gktb9_0(.dout(w_dff_A_WzXfX8em9_0),.din(w_dff_A_aGe0Gktb9_0),.clk(gclk));
	jdff dff_A_WzXfX8em9_0(.dout(w_dff_A_8f80AzCn1_0),.din(w_dff_A_WzXfX8em9_0),.clk(gclk));
	jdff dff_A_8f80AzCn1_0(.dout(w_dff_A_wmo9AFjC0_0),.din(w_dff_A_8f80AzCn1_0),.clk(gclk));
	jdff dff_A_wmo9AFjC0_0(.dout(w_dff_A_pYmXnEHf3_0),.din(w_dff_A_wmo9AFjC0_0),.clk(gclk));
	jdff dff_A_pYmXnEHf3_0(.dout(w_dff_A_0NJjoHbh9_0),.din(w_dff_A_pYmXnEHf3_0),.clk(gclk));
	jdff dff_A_0NJjoHbh9_0(.dout(w_dff_A_3a2wgAyG2_0),.din(w_dff_A_0NJjoHbh9_0),.clk(gclk));
	jdff dff_A_3a2wgAyG2_0(.dout(w_dff_A_P8qjI5I76_0),.din(w_dff_A_3a2wgAyG2_0),.clk(gclk));
	jdff dff_A_P8qjI5I76_0(.dout(w_dff_A_JgVGlE3Y2_0),.din(w_dff_A_P8qjI5I76_0),.clk(gclk));
	jdff dff_A_JgVGlE3Y2_0(.dout(w_dff_A_IbaDT5Bz6_0),.din(w_dff_A_JgVGlE3Y2_0),.clk(gclk));
	jdff dff_A_IbaDT5Bz6_0(.dout(w_dff_A_xVbIfwN30_0),.din(w_dff_A_IbaDT5Bz6_0),.clk(gclk));
	jdff dff_A_xVbIfwN30_0(.dout(w_dff_A_bw9XVCDf6_0),.din(w_dff_A_xVbIfwN30_0),.clk(gclk));
	jdff dff_A_bw9XVCDf6_0(.dout(w_dff_A_9LKUqm8Z1_0),.din(w_dff_A_bw9XVCDf6_0),.clk(gclk));
	jdff dff_A_9LKUqm8Z1_0(.dout(w_dff_A_3z8tURqP9_0),.din(w_dff_A_9LKUqm8Z1_0),.clk(gclk));
	jdff dff_A_3z8tURqP9_0(.dout(w_dff_A_l3by0rJL6_0),.din(w_dff_A_3z8tURqP9_0),.clk(gclk));
	jdff dff_A_l3by0rJL6_0(.dout(w_dff_A_AAdKUJSg5_0),.din(w_dff_A_l3by0rJL6_0),.clk(gclk));
	jdff dff_A_AAdKUJSg5_0(.dout(w_dff_A_pt1GigVO4_0),.din(w_dff_A_AAdKUJSg5_0),.clk(gclk));
	jdff dff_A_pt1GigVO4_0(.dout(w_dff_A_NS9ytCAQ5_0),.din(w_dff_A_pt1GigVO4_0),.clk(gclk));
	jdff dff_A_NS9ytCAQ5_0(.dout(w_dff_A_nT6kWBI53_0),.din(w_dff_A_NS9ytCAQ5_0),.clk(gclk));
	jdff dff_A_nT6kWBI53_0(.dout(G3552gat),.din(w_dff_A_nT6kWBI53_0),.clk(gclk));
	jdff dff_A_uq7HrGud8_2(.dout(w_dff_A_TMxT9gq27_0),.din(w_dff_A_uq7HrGud8_2),.clk(gclk));
	jdff dff_A_TMxT9gq27_0(.dout(w_dff_A_PsjvmN2d9_0),.din(w_dff_A_TMxT9gq27_0),.clk(gclk));
	jdff dff_A_PsjvmN2d9_0(.dout(w_dff_A_vXdKlroq6_0),.din(w_dff_A_PsjvmN2d9_0),.clk(gclk));
	jdff dff_A_vXdKlroq6_0(.dout(w_dff_A_qfwb87hp9_0),.din(w_dff_A_vXdKlroq6_0),.clk(gclk));
	jdff dff_A_qfwb87hp9_0(.dout(w_dff_A_L07fzR2f8_0),.din(w_dff_A_qfwb87hp9_0),.clk(gclk));
	jdff dff_A_L07fzR2f8_0(.dout(w_dff_A_971nGRUg1_0),.din(w_dff_A_L07fzR2f8_0),.clk(gclk));
	jdff dff_A_971nGRUg1_0(.dout(w_dff_A_SxVku1ct4_0),.din(w_dff_A_971nGRUg1_0),.clk(gclk));
	jdff dff_A_SxVku1ct4_0(.dout(w_dff_A_V3tVN4Im0_0),.din(w_dff_A_SxVku1ct4_0),.clk(gclk));
	jdff dff_A_V3tVN4Im0_0(.dout(w_dff_A_73MxvM4L4_0),.din(w_dff_A_V3tVN4Im0_0),.clk(gclk));
	jdff dff_A_73MxvM4L4_0(.dout(w_dff_A_Qr2dQSRe8_0),.din(w_dff_A_73MxvM4L4_0),.clk(gclk));
	jdff dff_A_Qr2dQSRe8_0(.dout(w_dff_A_6AuDajus5_0),.din(w_dff_A_Qr2dQSRe8_0),.clk(gclk));
	jdff dff_A_6AuDajus5_0(.dout(w_dff_A_KBSfT7WF8_0),.din(w_dff_A_6AuDajus5_0),.clk(gclk));
	jdff dff_A_KBSfT7WF8_0(.dout(w_dff_A_rN9DevVI5_0),.din(w_dff_A_KBSfT7WF8_0),.clk(gclk));
	jdff dff_A_rN9DevVI5_0(.dout(w_dff_A_rDKvsiUw2_0),.din(w_dff_A_rN9DevVI5_0),.clk(gclk));
	jdff dff_A_rDKvsiUw2_0(.dout(w_dff_A_db6qlW7L2_0),.din(w_dff_A_rDKvsiUw2_0),.clk(gclk));
	jdff dff_A_db6qlW7L2_0(.dout(w_dff_A_AjWnCn5s5_0),.din(w_dff_A_db6qlW7L2_0),.clk(gclk));
	jdff dff_A_AjWnCn5s5_0(.dout(w_dff_A_v6P0995l6_0),.din(w_dff_A_AjWnCn5s5_0),.clk(gclk));
	jdff dff_A_v6P0995l6_0(.dout(w_dff_A_HleEHpDh9_0),.din(w_dff_A_v6P0995l6_0),.clk(gclk));
	jdff dff_A_HleEHpDh9_0(.dout(w_dff_A_WVxaPR7a4_0),.din(w_dff_A_HleEHpDh9_0),.clk(gclk));
	jdff dff_A_WVxaPR7a4_0(.dout(w_dff_A_rsIb9tsD8_0),.din(w_dff_A_WVxaPR7a4_0),.clk(gclk));
	jdff dff_A_rsIb9tsD8_0(.dout(w_dff_A_MHvAQU5z9_0),.din(w_dff_A_rsIb9tsD8_0),.clk(gclk));
	jdff dff_A_MHvAQU5z9_0(.dout(w_dff_A_9XflZ5wp0_0),.din(w_dff_A_MHvAQU5z9_0),.clk(gclk));
	jdff dff_A_9XflZ5wp0_0(.dout(w_dff_A_UEueVxvp1_0),.din(w_dff_A_9XflZ5wp0_0),.clk(gclk));
	jdff dff_A_UEueVxvp1_0(.dout(w_dff_A_OIPmpoyZ1_0),.din(w_dff_A_UEueVxvp1_0),.clk(gclk));
	jdff dff_A_OIPmpoyZ1_0(.dout(w_dff_A_vImvgJRu9_0),.din(w_dff_A_OIPmpoyZ1_0),.clk(gclk));
	jdff dff_A_vImvgJRu9_0(.dout(w_dff_A_8h1GZ9yV9_0),.din(w_dff_A_vImvgJRu9_0),.clk(gclk));
	jdff dff_A_8h1GZ9yV9_0(.dout(w_dff_A_JHZmJGuN9_0),.din(w_dff_A_8h1GZ9yV9_0),.clk(gclk));
	jdff dff_A_JHZmJGuN9_0(.dout(w_dff_A_e3anqOcU8_0),.din(w_dff_A_JHZmJGuN9_0),.clk(gclk));
	jdff dff_A_e3anqOcU8_0(.dout(w_dff_A_NUDoO1gp9_0),.din(w_dff_A_e3anqOcU8_0),.clk(gclk));
	jdff dff_A_NUDoO1gp9_0(.dout(w_dff_A_BdB3dXRQ4_0),.din(w_dff_A_NUDoO1gp9_0),.clk(gclk));
	jdff dff_A_BdB3dXRQ4_0(.dout(w_dff_A_Y72CWuER7_0),.din(w_dff_A_BdB3dXRQ4_0),.clk(gclk));
	jdff dff_A_Y72CWuER7_0(.dout(w_dff_A_4KZaRmfv3_0),.din(w_dff_A_Y72CWuER7_0),.clk(gclk));
	jdff dff_A_4KZaRmfv3_0(.dout(w_dff_A_vAhxgl6A1_0),.din(w_dff_A_4KZaRmfv3_0),.clk(gclk));
	jdff dff_A_vAhxgl6A1_0(.dout(w_dff_A_tgqErB8D2_0),.din(w_dff_A_vAhxgl6A1_0),.clk(gclk));
	jdff dff_A_tgqErB8D2_0(.dout(w_dff_A_w1tZIuUt0_0),.din(w_dff_A_tgqErB8D2_0),.clk(gclk));
	jdff dff_A_w1tZIuUt0_0(.dout(w_dff_A_bXXoCxit5_0),.din(w_dff_A_w1tZIuUt0_0),.clk(gclk));
	jdff dff_A_bXXoCxit5_0(.dout(w_dff_A_RIUOzydE8_0),.din(w_dff_A_bXXoCxit5_0),.clk(gclk));
	jdff dff_A_RIUOzydE8_0(.dout(w_dff_A_uZT6NxH66_0),.din(w_dff_A_RIUOzydE8_0),.clk(gclk));
	jdff dff_A_uZT6NxH66_0(.dout(w_dff_A_6PVFqrjo6_0),.din(w_dff_A_uZT6NxH66_0),.clk(gclk));
	jdff dff_A_6PVFqrjo6_0(.dout(w_dff_A_mVpMqK286_0),.din(w_dff_A_6PVFqrjo6_0),.clk(gclk));
	jdff dff_A_mVpMqK286_0(.dout(w_dff_A_5ooabH5y0_0),.din(w_dff_A_mVpMqK286_0),.clk(gclk));
	jdff dff_A_5ooabH5y0_0(.dout(w_dff_A_LFHCtNum7_0),.din(w_dff_A_5ooabH5y0_0),.clk(gclk));
	jdff dff_A_LFHCtNum7_0(.dout(w_dff_A_mIL0jEPn8_0),.din(w_dff_A_LFHCtNum7_0),.clk(gclk));
	jdff dff_A_mIL0jEPn8_0(.dout(w_dff_A_srqtGN0P2_0),.din(w_dff_A_mIL0jEPn8_0),.clk(gclk));
	jdff dff_A_srqtGN0P2_0(.dout(w_dff_A_TAGBjDXW2_0),.din(w_dff_A_srqtGN0P2_0),.clk(gclk));
	jdff dff_A_TAGBjDXW2_0(.dout(w_dff_A_DY96cPWi0_0),.din(w_dff_A_TAGBjDXW2_0),.clk(gclk));
	jdff dff_A_DY96cPWi0_0(.dout(w_dff_A_vnoVe3jP8_0),.din(w_dff_A_DY96cPWi0_0),.clk(gclk));
	jdff dff_A_vnoVe3jP8_0(.dout(w_dff_A_VVtpKOgZ7_0),.din(w_dff_A_vnoVe3jP8_0),.clk(gclk));
	jdff dff_A_VVtpKOgZ7_0(.dout(w_dff_A_pw87yFbv8_0),.din(w_dff_A_VVtpKOgZ7_0),.clk(gclk));
	jdff dff_A_pw87yFbv8_0(.dout(w_dff_A_OubrqH7L0_0),.din(w_dff_A_pw87yFbv8_0),.clk(gclk));
	jdff dff_A_OubrqH7L0_0(.dout(G3895gat),.din(w_dff_A_OubrqH7L0_0),.clk(gclk));
	jdff dff_A_tHOt4IdH3_2(.dout(w_dff_A_7MZ2mz0k9_0),.din(w_dff_A_tHOt4IdH3_2),.clk(gclk));
	jdff dff_A_7MZ2mz0k9_0(.dout(w_dff_A_b53s00F83_0),.din(w_dff_A_7MZ2mz0k9_0),.clk(gclk));
	jdff dff_A_b53s00F83_0(.dout(w_dff_A_ON4f8Xev3_0),.din(w_dff_A_b53s00F83_0),.clk(gclk));
	jdff dff_A_ON4f8Xev3_0(.dout(w_dff_A_rcV7KJvx1_0),.din(w_dff_A_ON4f8Xev3_0),.clk(gclk));
	jdff dff_A_rcV7KJvx1_0(.dout(w_dff_A_jiCQ3TVQ2_0),.din(w_dff_A_rcV7KJvx1_0),.clk(gclk));
	jdff dff_A_jiCQ3TVQ2_0(.dout(w_dff_A_YYc3vBDR8_0),.din(w_dff_A_jiCQ3TVQ2_0),.clk(gclk));
	jdff dff_A_YYc3vBDR8_0(.dout(w_dff_A_jxbKZIqH0_0),.din(w_dff_A_YYc3vBDR8_0),.clk(gclk));
	jdff dff_A_jxbKZIqH0_0(.dout(w_dff_A_L1AwM1XF7_0),.din(w_dff_A_jxbKZIqH0_0),.clk(gclk));
	jdff dff_A_L1AwM1XF7_0(.dout(w_dff_A_dW5p6cFb7_0),.din(w_dff_A_L1AwM1XF7_0),.clk(gclk));
	jdff dff_A_dW5p6cFb7_0(.dout(w_dff_A_mCOWp0Dz3_0),.din(w_dff_A_dW5p6cFb7_0),.clk(gclk));
	jdff dff_A_mCOWp0Dz3_0(.dout(w_dff_A_BpcZKrht8_0),.din(w_dff_A_mCOWp0Dz3_0),.clk(gclk));
	jdff dff_A_BpcZKrht8_0(.dout(w_dff_A_UVpQz22G2_0),.din(w_dff_A_BpcZKrht8_0),.clk(gclk));
	jdff dff_A_UVpQz22G2_0(.dout(w_dff_A_ez836HoA6_0),.din(w_dff_A_UVpQz22G2_0),.clk(gclk));
	jdff dff_A_ez836HoA6_0(.dout(w_dff_A_RXF2V9y21_0),.din(w_dff_A_ez836HoA6_0),.clk(gclk));
	jdff dff_A_RXF2V9y21_0(.dout(w_dff_A_esYAQnNT3_0),.din(w_dff_A_RXF2V9y21_0),.clk(gclk));
	jdff dff_A_esYAQnNT3_0(.dout(w_dff_A_E7bdT8Qd7_0),.din(w_dff_A_esYAQnNT3_0),.clk(gclk));
	jdff dff_A_E7bdT8Qd7_0(.dout(w_dff_A_tWqpCV4W5_0),.din(w_dff_A_E7bdT8Qd7_0),.clk(gclk));
	jdff dff_A_tWqpCV4W5_0(.dout(w_dff_A_Bt6CXAh35_0),.din(w_dff_A_tWqpCV4W5_0),.clk(gclk));
	jdff dff_A_Bt6CXAh35_0(.dout(w_dff_A_KMM8obS68_0),.din(w_dff_A_Bt6CXAh35_0),.clk(gclk));
	jdff dff_A_KMM8obS68_0(.dout(w_dff_A_Er8mGpZx7_0),.din(w_dff_A_KMM8obS68_0),.clk(gclk));
	jdff dff_A_Er8mGpZx7_0(.dout(w_dff_A_GUNE9TJG3_0),.din(w_dff_A_Er8mGpZx7_0),.clk(gclk));
	jdff dff_A_GUNE9TJG3_0(.dout(w_dff_A_Hy7srK5u6_0),.din(w_dff_A_GUNE9TJG3_0),.clk(gclk));
	jdff dff_A_Hy7srK5u6_0(.dout(w_dff_A_ooQDCWvY6_0),.din(w_dff_A_Hy7srK5u6_0),.clk(gclk));
	jdff dff_A_ooQDCWvY6_0(.dout(w_dff_A_PjHqxL2c7_0),.din(w_dff_A_ooQDCWvY6_0),.clk(gclk));
	jdff dff_A_PjHqxL2c7_0(.dout(w_dff_A_Nm06FgkS6_0),.din(w_dff_A_PjHqxL2c7_0),.clk(gclk));
	jdff dff_A_Nm06FgkS6_0(.dout(w_dff_A_ukDWKzIP0_0),.din(w_dff_A_Nm06FgkS6_0),.clk(gclk));
	jdff dff_A_ukDWKzIP0_0(.dout(w_dff_A_psb2gkeg9_0),.din(w_dff_A_ukDWKzIP0_0),.clk(gclk));
	jdff dff_A_psb2gkeg9_0(.dout(w_dff_A_oqhmc8u12_0),.din(w_dff_A_psb2gkeg9_0),.clk(gclk));
	jdff dff_A_oqhmc8u12_0(.dout(w_dff_A_WhpULsPz1_0),.din(w_dff_A_oqhmc8u12_0),.clk(gclk));
	jdff dff_A_WhpULsPz1_0(.dout(w_dff_A_FFeUrgin0_0),.din(w_dff_A_WhpULsPz1_0),.clk(gclk));
	jdff dff_A_FFeUrgin0_0(.dout(w_dff_A_KtR2M6lK4_0),.din(w_dff_A_FFeUrgin0_0),.clk(gclk));
	jdff dff_A_KtR2M6lK4_0(.dout(w_dff_A_3GKXB7wb8_0),.din(w_dff_A_KtR2M6lK4_0),.clk(gclk));
	jdff dff_A_3GKXB7wb8_0(.dout(w_dff_A_OwuJQKDl3_0),.din(w_dff_A_3GKXB7wb8_0),.clk(gclk));
	jdff dff_A_OwuJQKDl3_0(.dout(w_dff_A_XSDVcXWM2_0),.din(w_dff_A_OwuJQKDl3_0),.clk(gclk));
	jdff dff_A_XSDVcXWM2_0(.dout(w_dff_A_LGv7DrxZ3_0),.din(w_dff_A_XSDVcXWM2_0),.clk(gclk));
	jdff dff_A_LGv7DrxZ3_0(.dout(w_dff_A_1RQp3Hw82_0),.din(w_dff_A_LGv7DrxZ3_0),.clk(gclk));
	jdff dff_A_1RQp3Hw82_0(.dout(w_dff_A_k7OETGIC4_0),.din(w_dff_A_1RQp3Hw82_0),.clk(gclk));
	jdff dff_A_k7OETGIC4_0(.dout(w_dff_A_jmvKePer1_0),.din(w_dff_A_k7OETGIC4_0),.clk(gclk));
	jdff dff_A_jmvKePer1_0(.dout(w_dff_A_CoEy92EC6_0),.din(w_dff_A_jmvKePer1_0),.clk(gclk));
	jdff dff_A_CoEy92EC6_0(.dout(w_dff_A_wfgYk0t26_0),.din(w_dff_A_CoEy92EC6_0),.clk(gclk));
	jdff dff_A_wfgYk0t26_0(.dout(w_dff_A_v0I5MAlB2_0),.din(w_dff_A_wfgYk0t26_0),.clk(gclk));
	jdff dff_A_v0I5MAlB2_0(.dout(w_dff_A_pud9JJYd8_0),.din(w_dff_A_v0I5MAlB2_0),.clk(gclk));
	jdff dff_A_pud9JJYd8_0(.dout(w_dff_A_thm4pJLX7_0),.din(w_dff_A_pud9JJYd8_0),.clk(gclk));
	jdff dff_A_thm4pJLX7_0(.dout(w_dff_A_o77bWtWN7_0),.din(w_dff_A_thm4pJLX7_0),.clk(gclk));
	jdff dff_A_o77bWtWN7_0(.dout(w_dff_A_tQlpkEYN5_0),.din(w_dff_A_o77bWtWN7_0),.clk(gclk));
	jdff dff_A_tQlpkEYN5_0(.dout(w_dff_A_DIG3mYDe4_0),.din(w_dff_A_tQlpkEYN5_0),.clk(gclk));
	jdff dff_A_DIG3mYDe4_0(.dout(w_dff_A_H5p053tj6_0),.din(w_dff_A_DIG3mYDe4_0),.clk(gclk));
	jdff dff_A_H5p053tj6_0(.dout(G4241gat),.din(w_dff_A_H5p053tj6_0),.clk(gclk));
	jdff dff_A_c2Mb5ZJa8_2(.dout(w_dff_A_2QtLixsD2_0),.din(w_dff_A_c2Mb5ZJa8_2),.clk(gclk));
	jdff dff_A_2QtLixsD2_0(.dout(w_dff_A_uuvaZpmj0_0),.din(w_dff_A_2QtLixsD2_0),.clk(gclk));
	jdff dff_A_uuvaZpmj0_0(.dout(w_dff_A_mYaJyjgA8_0),.din(w_dff_A_uuvaZpmj0_0),.clk(gclk));
	jdff dff_A_mYaJyjgA8_0(.dout(w_dff_A_mufysFVm3_0),.din(w_dff_A_mYaJyjgA8_0),.clk(gclk));
	jdff dff_A_mufysFVm3_0(.dout(w_dff_A_2OdettXL0_0),.din(w_dff_A_mufysFVm3_0),.clk(gclk));
	jdff dff_A_2OdettXL0_0(.dout(w_dff_A_a7kqf7gA5_0),.din(w_dff_A_2OdettXL0_0),.clk(gclk));
	jdff dff_A_a7kqf7gA5_0(.dout(w_dff_A_SHPEgKHV2_0),.din(w_dff_A_a7kqf7gA5_0),.clk(gclk));
	jdff dff_A_SHPEgKHV2_0(.dout(w_dff_A_FF0HUAtC9_0),.din(w_dff_A_SHPEgKHV2_0),.clk(gclk));
	jdff dff_A_FF0HUAtC9_0(.dout(w_dff_A_AIuHiakr5_0),.din(w_dff_A_FF0HUAtC9_0),.clk(gclk));
	jdff dff_A_AIuHiakr5_0(.dout(w_dff_A_XmEka2YI7_0),.din(w_dff_A_AIuHiakr5_0),.clk(gclk));
	jdff dff_A_XmEka2YI7_0(.dout(w_dff_A_NLUI8hMV8_0),.din(w_dff_A_XmEka2YI7_0),.clk(gclk));
	jdff dff_A_NLUI8hMV8_0(.dout(w_dff_A_Bml7fNx51_0),.din(w_dff_A_NLUI8hMV8_0),.clk(gclk));
	jdff dff_A_Bml7fNx51_0(.dout(w_dff_A_OmdLPao80_0),.din(w_dff_A_Bml7fNx51_0),.clk(gclk));
	jdff dff_A_OmdLPao80_0(.dout(w_dff_A_wOHgARtJ1_0),.din(w_dff_A_OmdLPao80_0),.clk(gclk));
	jdff dff_A_wOHgARtJ1_0(.dout(w_dff_A_1uVmMeJY5_0),.din(w_dff_A_wOHgARtJ1_0),.clk(gclk));
	jdff dff_A_1uVmMeJY5_0(.dout(w_dff_A_MCQdHX6S4_0),.din(w_dff_A_1uVmMeJY5_0),.clk(gclk));
	jdff dff_A_MCQdHX6S4_0(.dout(w_dff_A_e6nGIGsS4_0),.din(w_dff_A_MCQdHX6S4_0),.clk(gclk));
	jdff dff_A_e6nGIGsS4_0(.dout(w_dff_A_GvN2DDQe0_0),.din(w_dff_A_e6nGIGsS4_0),.clk(gclk));
	jdff dff_A_GvN2DDQe0_0(.dout(w_dff_A_6cqk7zSv7_0),.din(w_dff_A_GvN2DDQe0_0),.clk(gclk));
	jdff dff_A_6cqk7zSv7_0(.dout(w_dff_A_IG0gKjKu3_0),.din(w_dff_A_6cqk7zSv7_0),.clk(gclk));
	jdff dff_A_IG0gKjKu3_0(.dout(w_dff_A_fVajJqO53_0),.din(w_dff_A_IG0gKjKu3_0),.clk(gclk));
	jdff dff_A_fVajJqO53_0(.dout(w_dff_A_VX9jnV2g5_0),.din(w_dff_A_fVajJqO53_0),.clk(gclk));
	jdff dff_A_VX9jnV2g5_0(.dout(w_dff_A_T05j5q9S7_0),.din(w_dff_A_VX9jnV2g5_0),.clk(gclk));
	jdff dff_A_T05j5q9S7_0(.dout(w_dff_A_O8KAUTFA7_0),.din(w_dff_A_T05j5q9S7_0),.clk(gclk));
	jdff dff_A_O8KAUTFA7_0(.dout(w_dff_A_30WMGuhX5_0),.din(w_dff_A_O8KAUTFA7_0),.clk(gclk));
	jdff dff_A_30WMGuhX5_0(.dout(w_dff_A_qTIIqKoI4_0),.din(w_dff_A_30WMGuhX5_0),.clk(gclk));
	jdff dff_A_qTIIqKoI4_0(.dout(w_dff_A_C2fTUw5T8_0),.din(w_dff_A_qTIIqKoI4_0),.clk(gclk));
	jdff dff_A_C2fTUw5T8_0(.dout(w_dff_A_ZGz6OgcM6_0),.din(w_dff_A_C2fTUw5T8_0),.clk(gclk));
	jdff dff_A_ZGz6OgcM6_0(.dout(w_dff_A_Adb92XRc7_0),.din(w_dff_A_ZGz6OgcM6_0),.clk(gclk));
	jdff dff_A_Adb92XRc7_0(.dout(w_dff_A_VkDvRo3x6_0),.din(w_dff_A_Adb92XRc7_0),.clk(gclk));
	jdff dff_A_VkDvRo3x6_0(.dout(w_dff_A_edGDrP0i1_0),.din(w_dff_A_VkDvRo3x6_0),.clk(gclk));
	jdff dff_A_edGDrP0i1_0(.dout(w_dff_A_LyBLZUL77_0),.din(w_dff_A_edGDrP0i1_0),.clk(gclk));
	jdff dff_A_LyBLZUL77_0(.dout(w_dff_A_KSp9iXih7_0),.din(w_dff_A_LyBLZUL77_0),.clk(gclk));
	jdff dff_A_KSp9iXih7_0(.dout(w_dff_A_CqboO7gP9_0),.din(w_dff_A_KSp9iXih7_0),.clk(gclk));
	jdff dff_A_CqboO7gP9_0(.dout(w_dff_A_wTqkJNrg5_0),.din(w_dff_A_CqboO7gP9_0),.clk(gclk));
	jdff dff_A_wTqkJNrg5_0(.dout(w_dff_A_SUDamReS7_0),.din(w_dff_A_wTqkJNrg5_0),.clk(gclk));
	jdff dff_A_SUDamReS7_0(.dout(w_dff_A_xMWb35Nh5_0),.din(w_dff_A_SUDamReS7_0),.clk(gclk));
	jdff dff_A_xMWb35Nh5_0(.dout(w_dff_A_FX2pFjiI5_0),.din(w_dff_A_xMWb35Nh5_0),.clk(gclk));
	jdff dff_A_FX2pFjiI5_0(.dout(w_dff_A_YgLFpDns5_0),.din(w_dff_A_FX2pFjiI5_0),.clk(gclk));
	jdff dff_A_YgLFpDns5_0(.dout(w_dff_A_OBDpYuvZ6_0),.din(w_dff_A_YgLFpDns5_0),.clk(gclk));
	jdff dff_A_OBDpYuvZ6_0(.dout(w_dff_A_4fkCDQ9o1_0),.din(w_dff_A_OBDpYuvZ6_0),.clk(gclk));
	jdff dff_A_4fkCDQ9o1_0(.dout(w_dff_A_FxMM6J437_0),.din(w_dff_A_4fkCDQ9o1_0),.clk(gclk));
	jdff dff_A_FxMM6J437_0(.dout(w_dff_A_kqZzRckG2_0),.din(w_dff_A_FxMM6J437_0),.clk(gclk));
	jdff dff_A_kqZzRckG2_0(.dout(w_dff_A_VKpCHKDA0_0),.din(w_dff_A_kqZzRckG2_0),.clk(gclk));
	jdff dff_A_VKpCHKDA0_0(.dout(G4591gat),.din(w_dff_A_VKpCHKDA0_0),.clk(gclk));
	jdff dff_A_BoBfaVd45_2(.dout(w_dff_A_HUwlSYhX6_0),.din(w_dff_A_BoBfaVd45_2),.clk(gclk));
	jdff dff_A_HUwlSYhX6_0(.dout(w_dff_A_oIUR6dqM9_0),.din(w_dff_A_HUwlSYhX6_0),.clk(gclk));
	jdff dff_A_oIUR6dqM9_0(.dout(w_dff_A_CzJaNVTa4_0),.din(w_dff_A_oIUR6dqM9_0),.clk(gclk));
	jdff dff_A_CzJaNVTa4_0(.dout(w_dff_A_9sacLv096_0),.din(w_dff_A_CzJaNVTa4_0),.clk(gclk));
	jdff dff_A_9sacLv096_0(.dout(w_dff_A_0ZElR9Dc1_0),.din(w_dff_A_9sacLv096_0),.clk(gclk));
	jdff dff_A_0ZElR9Dc1_0(.dout(w_dff_A_HIkn0sTv5_0),.din(w_dff_A_0ZElR9Dc1_0),.clk(gclk));
	jdff dff_A_HIkn0sTv5_0(.dout(w_dff_A_wbvpgRiS7_0),.din(w_dff_A_HIkn0sTv5_0),.clk(gclk));
	jdff dff_A_wbvpgRiS7_0(.dout(w_dff_A_xAdwfQ3B9_0),.din(w_dff_A_wbvpgRiS7_0),.clk(gclk));
	jdff dff_A_xAdwfQ3B9_0(.dout(w_dff_A_deja45NH0_0),.din(w_dff_A_xAdwfQ3B9_0),.clk(gclk));
	jdff dff_A_deja45NH0_0(.dout(w_dff_A_BwkW8nvS9_0),.din(w_dff_A_deja45NH0_0),.clk(gclk));
	jdff dff_A_BwkW8nvS9_0(.dout(w_dff_A_x2m5ql8I9_0),.din(w_dff_A_BwkW8nvS9_0),.clk(gclk));
	jdff dff_A_x2m5ql8I9_0(.dout(w_dff_A_mKLxjuKN6_0),.din(w_dff_A_x2m5ql8I9_0),.clk(gclk));
	jdff dff_A_mKLxjuKN6_0(.dout(w_dff_A_MFDQ4FUW7_0),.din(w_dff_A_mKLxjuKN6_0),.clk(gclk));
	jdff dff_A_MFDQ4FUW7_0(.dout(w_dff_A_gz2DMb8F5_0),.din(w_dff_A_MFDQ4FUW7_0),.clk(gclk));
	jdff dff_A_gz2DMb8F5_0(.dout(w_dff_A_JXtw0OmZ1_0),.din(w_dff_A_gz2DMb8F5_0),.clk(gclk));
	jdff dff_A_JXtw0OmZ1_0(.dout(w_dff_A_nrJ9HFnl9_0),.din(w_dff_A_JXtw0OmZ1_0),.clk(gclk));
	jdff dff_A_nrJ9HFnl9_0(.dout(w_dff_A_1m26w6zd1_0),.din(w_dff_A_nrJ9HFnl9_0),.clk(gclk));
	jdff dff_A_1m26w6zd1_0(.dout(w_dff_A_1r3QkQAT1_0),.din(w_dff_A_1m26w6zd1_0),.clk(gclk));
	jdff dff_A_1r3QkQAT1_0(.dout(w_dff_A_uC2UPu4F6_0),.din(w_dff_A_1r3QkQAT1_0),.clk(gclk));
	jdff dff_A_uC2UPu4F6_0(.dout(w_dff_A_oxskycKV2_0),.din(w_dff_A_uC2UPu4F6_0),.clk(gclk));
	jdff dff_A_oxskycKV2_0(.dout(w_dff_A_p6BT5YFx8_0),.din(w_dff_A_oxskycKV2_0),.clk(gclk));
	jdff dff_A_p6BT5YFx8_0(.dout(w_dff_A_6JPh4bs26_0),.din(w_dff_A_p6BT5YFx8_0),.clk(gclk));
	jdff dff_A_6JPh4bs26_0(.dout(w_dff_A_wnTXVRLI8_0),.din(w_dff_A_6JPh4bs26_0),.clk(gclk));
	jdff dff_A_wnTXVRLI8_0(.dout(w_dff_A_v6j4jcbP7_0),.din(w_dff_A_wnTXVRLI8_0),.clk(gclk));
	jdff dff_A_v6j4jcbP7_0(.dout(w_dff_A_jOoIs8z15_0),.din(w_dff_A_v6j4jcbP7_0),.clk(gclk));
	jdff dff_A_jOoIs8z15_0(.dout(w_dff_A_kS8S7GOY8_0),.din(w_dff_A_jOoIs8z15_0),.clk(gclk));
	jdff dff_A_kS8S7GOY8_0(.dout(w_dff_A_EztnLaan4_0),.din(w_dff_A_kS8S7GOY8_0),.clk(gclk));
	jdff dff_A_EztnLaan4_0(.dout(w_dff_A_qgEKCMsP4_0),.din(w_dff_A_EztnLaan4_0),.clk(gclk));
	jdff dff_A_qgEKCMsP4_0(.dout(w_dff_A_daTCcLCA0_0),.din(w_dff_A_qgEKCMsP4_0),.clk(gclk));
	jdff dff_A_daTCcLCA0_0(.dout(w_dff_A_UTAKWyje5_0),.din(w_dff_A_daTCcLCA0_0),.clk(gclk));
	jdff dff_A_UTAKWyje5_0(.dout(w_dff_A_hT4eIrcv5_0),.din(w_dff_A_UTAKWyje5_0),.clk(gclk));
	jdff dff_A_hT4eIrcv5_0(.dout(w_dff_A_wIV3bZsk2_0),.din(w_dff_A_hT4eIrcv5_0),.clk(gclk));
	jdff dff_A_wIV3bZsk2_0(.dout(w_dff_A_1Vw0DgM69_0),.din(w_dff_A_wIV3bZsk2_0),.clk(gclk));
	jdff dff_A_1Vw0DgM69_0(.dout(w_dff_A_dFckzMtr4_0),.din(w_dff_A_1Vw0DgM69_0),.clk(gclk));
	jdff dff_A_dFckzMtr4_0(.dout(w_dff_A_5BEBlbZ29_0),.din(w_dff_A_dFckzMtr4_0),.clk(gclk));
	jdff dff_A_5BEBlbZ29_0(.dout(w_dff_A_PN0c7vH34_0),.din(w_dff_A_5BEBlbZ29_0),.clk(gclk));
	jdff dff_A_PN0c7vH34_0(.dout(w_dff_A_DhitR4bT0_0),.din(w_dff_A_PN0c7vH34_0),.clk(gclk));
	jdff dff_A_DhitR4bT0_0(.dout(w_dff_A_PbYHS0fY7_0),.din(w_dff_A_DhitR4bT0_0),.clk(gclk));
	jdff dff_A_PbYHS0fY7_0(.dout(w_dff_A_x8gxo9aW4_0),.din(w_dff_A_PbYHS0fY7_0),.clk(gclk));
	jdff dff_A_x8gxo9aW4_0(.dout(w_dff_A_y0Hedgor8_0),.din(w_dff_A_x8gxo9aW4_0),.clk(gclk));
	jdff dff_A_y0Hedgor8_0(.dout(w_dff_A_4FbZpWqa9_0),.din(w_dff_A_y0Hedgor8_0),.clk(gclk));
	jdff dff_A_4FbZpWqa9_0(.dout(G4946gat),.din(w_dff_A_4FbZpWqa9_0),.clk(gclk));
	jdff dff_A_KgRkqf0R7_2(.dout(w_dff_A_57TOYDhe0_0),.din(w_dff_A_KgRkqf0R7_2),.clk(gclk));
	jdff dff_A_57TOYDhe0_0(.dout(w_dff_A_fQwaJS1I2_0),.din(w_dff_A_57TOYDhe0_0),.clk(gclk));
	jdff dff_A_fQwaJS1I2_0(.dout(w_dff_A_eMsrY0Yu1_0),.din(w_dff_A_fQwaJS1I2_0),.clk(gclk));
	jdff dff_A_eMsrY0Yu1_0(.dout(w_dff_A_tahyBwYu3_0),.din(w_dff_A_eMsrY0Yu1_0),.clk(gclk));
	jdff dff_A_tahyBwYu3_0(.dout(w_dff_A_VMzGH1sg5_0),.din(w_dff_A_tahyBwYu3_0),.clk(gclk));
	jdff dff_A_VMzGH1sg5_0(.dout(w_dff_A_QaHnpNmE9_0),.din(w_dff_A_VMzGH1sg5_0),.clk(gclk));
	jdff dff_A_QaHnpNmE9_0(.dout(w_dff_A_eoRusGuQ0_0),.din(w_dff_A_QaHnpNmE9_0),.clk(gclk));
	jdff dff_A_eoRusGuQ0_0(.dout(w_dff_A_E2a54sDe0_0),.din(w_dff_A_eoRusGuQ0_0),.clk(gclk));
	jdff dff_A_E2a54sDe0_0(.dout(w_dff_A_sQMCH4ZL4_0),.din(w_dff_A_E2a54sDe0_0),.clk(gclk));
	jdff dff_A_sQMCH4ZL4_0(.dout(w_dff_A_yCGMJXXz7_0),.din(w_dff_A_sQMCH4ZL4_0),.clk(gclk));
	jdff dff_A_yCGMJXXz7_0(.dout(w_dff_A_7o0AS5ii1_0),.din(w_dff_A_yCGMJXXz7_0),.clk(gclk));
	jdff dff_A_7o0AS5ii1_0(.dout(w_dff_A_0xDEqeb50_0),.din(w_dff_A_7o0AS5ii1_0),.clk(gclk));
	jdff dff_A_0xDEqeb50_0(.dout(w_dff_A_wwATG9FF7_0),.din(w_dff_A_0xDEqeb50_0),.clk(gclk));
	jdff dff_A_wwATG9FF7_0(.dout(w_dff_A_HnjsgwUJ7_0),.din(w_dff_A_wwATG9FF7_0),.clk(gclk));
	jdff dff_A_HnjsgwUJ7_0(.dout(w_dff_A_TONDlJX68_0),.din(w_dff_A_HnjsgwUJ7_0),.clk(gclk));
	jdff dff_A_TONDlJX68_0(.dout(w_dff_A_4EGW1fdJ4_0),.din(w_dff_A_TONDlJX68_0),.clk(gclk));
	jdff dff_A_4EGW1fdJ4_0(.dout(w_dff_A_wnSFTbd79_0),.din(w_dff_A_4EGW1fdJ4_0),.clk(gclk));
	jdff dff_A_wnSFTbd79_0(.dout(w_dff_A_gMyykVh03_0),.din(w_dff_A_wnSFTbd79_0),.clk(gclk));
	jdff dff_A_gMyykVh03_0(.dout(w_dff_A_wenZNzJ06_0),.din(w_dff_A_gMyykVh03_0),.clk(gclk));
	jdff dff_A_wenZNzJ06_0(.dout(w_dff_A_VzdA0mXs9_0),.din(w_dff_A_wenZNzJ06_0),.clk(gclk));
	jdff dff_A_VzdA0mXs9_0(.dout(w_dff_A_F4832aG50_0),.din(w_dff_A_VzdA0mXs9_0),.clk(gclk));
	jdff dff_A_F4832aG50_0(.dout(w_dff_A_RbuTCF7e5_0),.din(w_dff_A_F4832aG50_0),.clk(gclk));
	jdff dff_A_RbuTCF7e5_0(.dout(w_dff_A_Bgt5IYUY9_0),.din(w_dff_A_RbuTCF7e5_0),.clk(gclk));
	jdff dff_A_Bgt5IYUY9_0(.dout(w_dff_A_Ssko7M8N9_0),.din(w_dff_A_Bgt5IYUY9_0),.clk(gclk));
	jdff dff_A_Ssko7M8N9_0(.dout(w_dff_A_lXMPsd2B7_0),.din(w_dff_A_Ssko7M8N9_0),.clk(gclk));
	jdff dff_A_lXMPsd2B7_0(.dout(w_dff_A_at9SIGRH3_0),.din(w_dff_A_lXMPsd2B7_0),.clk(gclk));
	jdff dff_A_at9SIGRH3_0(.dout(w_dff_A_MxziXfO06_0),.din(w_dff_A_at9SIGRH3_0),.clk(gclk));
	jdff dff_A_MxziXfO06_0(.dout(w_dff_A_E9eGopf17_0),.din(w_dff_A_MxziXfO06_0),.clk(gclk));
	jdff dff_A_E9eGopf17_0(.dout(w_dff_A_T8eY0KiG9_0),.din(w_dff_A_E9eGopf17_0),.clk(gclk));
	jdff dff_A_T8eY0KiG9_0(.dout(w_dff_A_5mKPFMY43_0),.din(w_dff_A_T8eY0KiG9_0),.clk(gclk));
	jdff dff_A_5mKPFMY43_0(.dout(w_dff_A_bCXUs6fO8_0),.din(w_dff_A_5mKPFMY43_0),.clk(gclk));
	jdff dff_A_bCXUs6fO8_0(.dout(w_dff_A_5gQRNCgM9_0),.din(w_dff_A_bCXUs6fO8_0),.clk(gclk));
	jdff dff_A_5gQRNCgM9_0(.dout(w_dff_A_qk7Gvbf94_0),.din(w_dff_A_5gQRNCgM9_0),.clk(gclk));
	jdff dff_A_qk7Gvbf94_0(.dout(w_dff_A_lrigsKGL7_0),.din(w_dff_A_qk7Gvbf94_0),.clk(gclk));
	jdff dff_A_lrigsKGL7_0(.dout(w_dff_A_i8B0Knw88_0),.din(w_dff_A_lrigsKGL7_0),.clk(gclk));
	jdff dff_A_i8B0Knw88_0(.dout(w_dff_A_yGXwLH0h1_0),.din(w_dff_A_i8B0Knw88_0),.clk(gclk));
	jdff dff_A_yGXwLH0h1_0(.dout(w_dff_A_liBpevxS9_0),.din(w_dff_A_yGXwLH0h1_0),.clk(gclk));
	jdff dff_A_liBpevxS9_0(.dout(w_dff_A_LGhsnsmq0_0),.din(w_dff_A_liBpevxS9_0),.clk(gclk));
	jdff dff_A_LGhsnsmq0_0(.dout(G5308gat),.din(w_dff_A_LGhsnsmq0_0),.clk(gclk));
	jdff dff_A_WOK9KqFE4_2(.dout(w_dff_A_ndBKPnsb5_0),.din(w_dff_A_WOK9KqFE4_2),.clk(gclk));
	jdff dff_A_ndBKPnsb5_0(.dout(w_dff_A_9FPoiyZj3_0),.din(w_dff_A_ndBKPnsb5_0),.clk(gclk));
	jdff dff_A_9FPoiyZj3_0(.dout(w_dff_A_MWTCJmFJ4_0),.din(w_dff_A_9FPoiyZj3_0),.clk(gclk));
	jdff dff_A_MWTCJmFJ4_0(.dout(w_dff_A_1ZDy1A874_0),.din(w_dff_A_MWTCJmFJ4_0),.clk(gclk));
	jdff dff_A_1ZDy1A874_0(.dout(w_dff_A_ZZO9IYEu9_0),.din(w_dff_A_1ZDy1A874_0),.clk(gclk));
	jdff dff_A_ZZO9IYEu9_0(.dout(w_dff_A_qduycNea2_0),.din(w_dff_A_ZZO9IYEu9_0),.clk(gclk));
	jdff dff_A_qduycNea2_0(.dout(w_dff_A_2spqaFr38_0),.din(w_dff_A_qduycNea2_0),.clk(gclk));
	jdff dff_A_2spqaFr38_0(.dout(w_dff_A_ole6pWoS9_0),.din(w_dff_A_2spqaFr38_0),.clk(gclk));
	jdff dff_A_ole6pWoS9_0(.dout(w_dff_A_KBiPeFWu1_0),.din(w_dff_A_ole6pWoS9_0),.clk(gclk));
	jdff dff_A_KBiPeFWu1_0(.dout(w_dff_A_ijdeybMF7_0),.din(w_dff_A_KBiPeFWu1_0),.clk(gclk));
	jdff dff_A_ijdeybMF7_0(.dout(w_dff_A_d622vyQJ8_0),.din(w_dff_A_ijdeybMF7_0),.clk(gclk));
	jdff dff_A_d622vyQJ8_0(.dout(w_dff_A_gCXp2lHf5_0),.din(w_dff_A_d622vyQJ8_0),.clk(gclk));
	jdff dff_A_gCXp2lHf5_0(.dout(w_dff_A_j0ID7f9B8_0),.din(w_dff_A_gCXp2lHf5_0),.clk(gclk));
	jdff dff_A_j0ID7f9B8_0(.dout(w_dff_A_ueqchTOU7_0),.din(w_dff_A_j0ID7f9B8_0),.clk(gclk));
	jdff dff_A_ueqchTOU7_0(.dout(w_dff_A_MBwDEREv2_0),.din(w_dff_A_ueqchTOU7_0),.clk(gclk));
	jdff dff_A_MBwDEREv2_0(.dout(w_dff_A_74Iev9hV4_0),.din(w_dff_A_MBwDEREv2_0),.clk(gclk));
	jdff dff_A_74Iev9hV4_0(.dout(w_dff_A_OWYvHwqG4_0),.din(w_dff_A_74Iev9hV4_0),.clk(gclk));
	jdff dff_A_OWYvHwqG4_0(.dout(w_dff_A_v62q8RnP2_0),.din(w_dff_A_OWYvHwqG4_0),.clk(gclk));
	jdff dff_A_v62q8RnP2_0(.dout(w_dff_A_Dw4O4psQ2_0),.din(w_dff_A_v62q8RnP2_0),.clk(gclk));
	jdff dff_A_Dw4O4psQ2_0(.dout(w_dff_A_xrq29jW81_0),.din(w_dff_A_Dw4O4psQ2_0),.clk(gclk));
	jdff dff_A_xrq29jW81_0(.dout(w_dff_A_GCfYRd367_0),.din(w_dff_A_xrq29jW81_0),.clk(gclk));
	jdff dff_A_GCfYRd367_0(.dout(w_dff_A_5R800uff2_0),.din(w_dff_A_GCfYRd367_0),.clk(gclk));
	jdff dff_A_5R800uff2_0(.dout(w_dff_A_iGcAk4P08_0),.din(w_dff_A_5R800uff2_0),.clk(gclk));
	jdff dff_A_iGcAk4P08_0(.dout(w_dff_A_TN8vkqXp6_0),.din(w_dff_A_iGcAk4P08_0),.clk(gclk));
	jdff dff_A_TN8vkqXp6_0(.dout(w_dff_A_CwtW7hEU5_0),.din(w_dff_A_TN8vkqXp6_0),.clk(gclk));
	jdff dff_A_CwtW7hEU5_0(.dout(w_dff_A_zRjZBrFB2_0),.din(w_dff_A_CwtW7hEU5_0),.clk(gclk));
	jdff dff_A_zRjZBrFB2_0(.dout(w_dff_A_tnAyMi1B7_0),.din(w_dff_A_zRjZBrFB2_0),.clk(gclk));
	jdff dff_A_tnAyMi1B7_0(.dout(w_dff_A_yi6Rjdes2_0),.din(w_dff_A_tnAyMi1B7_0),.clk(gclk));
	jdff dff_A_yi6Rjdes2_0(.dout(w_dff_A_fnskD6jX3_0),.din(w_dff_A_yi6Rjdes2_0),.clk(gclk));
	jdff dff_A_fnskD6jX3_0(.dout(w_dff_A_sgerVUJA3_0),.din(w_dff_A_fnskD6jX3_0),.clk(gclk));
	jdff dff_A_sgerVUJA3_0(.dout(w_dff_A_p9kkbE3G7_0),.din(w_dff_A_sgerVUJA3_0),.clk(gclk));
	jdff dff_A_p9kkbE3G7_0(.dout(w_dff_A_Ms9amRbX0_0),.din(w_dff_A_p9kkbE3G7_0),.clk(gclk));
	jdff dff_A_Ms9amRbX0_0(.dout(w_dff_A_X6YQEXw06_0),.din(w_dff_A_Ms9amRbX0_0),.clk(gclk));
	jdff dff_A_X6YQEXw06_0(.dout(w_dff_A_XJaLv4NV8_0),.din(w_dff_A_X6YQEXw06_0),.clk(gclk));
	jdff dff_A_XJaLv4NV8_0(.dout(w_dff_A_lH8qR5tA7_0),.din(w_dff_A_XJaLv4NV8_0),.clk(gclk));
	jdff dff_A_lH8qR5tA7_0(.dout(G5672gat),.din(w_dff_A_lH8qR5tA7_0),.clk(gclk));
	jdff dff_A_Mc6r1u771_2(.dout(w_dff_A_dX7JRheo4_0),.din(w_dff_A_Mc6r1u771_2),.clk(gclk));
	jdff dff_A_dX7JRheo4_0(.dout(w_dff_A_OUzDuztl7_0),.din(w_dff_A_dX7JRheo4_0),.clk(gclk));
	jdff dff_A_OUzDuztl7_0(.dout(w_dff_A_iJoGHwXF7_0),.din(w_dff_A_OUzDuztl7_0),.clk(gclk));
	jdff dff_A_iJoGHwXF7_0(.dout(w_dff_A_x3YpxVtV3_0),.din(w_dff_A_iJoGHwXF7_0),.clk(gclk));
	jdff dff_A_x3YpxVtV3_0(.dout(w_dff_A_ee2Zi4Ac3_0),.din(w_dff_A_x3YpxVtV3_0),.clk(gclk));
	jdff dff_A_ee2Zi4Ac3_0(.dout(w_dff_A_xlpeibEP4_0),.din(w_dff_A_ee2Zi4Ac3_0),.clk(gclk));
	jdff dff_A_xlpeibEP4_0(.dout(w_dff_A_j8VdFpOx2_0),.din(w_dff_A_xlpeibEP4_0),.clk(gclk));
	jdff dff_A_j8VdFpOx2_0(.dout(w_dff_A_6WjwWCuz3_0),.din(w_dff_A_j8VdFpOx2_0),.clk(gclk));
	jdff dff_A_6WjwWCuz3_0(.dout(w_dff_A_GJ3arNn35_0),.din(w_dff_A_6WjwWCuz3_0),.clk(gclk));
	jdff dff_A_GJ3arNn35_0(.dout(w_dff_A_w8sfpaRZ1_0),.din(w_dff_A_GJ3arNn35_0),.clk(gclk));
	jdff dff_A_w8sfpaRZ1_0(.dout(w_dff_A_cZz6kNqm6_0),.din(w_dff_A_w8sfpaRZ1_0),.clk(gclk));
	jdff dff_A_cZz6kNqm6_0(.dout(w_dff_A_QmjvM2kS7_0),.din(w_dff_A_cZz6kNqm6_0),.clk(gclk));
	jdff dff_A_QmjvM2kS7_0(.dout(w_dff_A_7gsmhxh15_0),.din(w_dff_A_QmjvM2kS7_0),.clk(gclk));
	jdff dff_A_7gsmhxh15_0(.dout(w_dff_A_5ENBYldk3_0),.din(w_dff_A_7gsmhxh15_0),.clk(gclk));
	jdff dff_A_5ENBYldk3_0(.dout(w_dff_A_q4x1fN763_0),.din(w_dff_A_5ENBYldk3_0),.clk(gclk));
	jdff dff_A_q4x1fN763_0(.dout(w_dff_A_tpSB7hXw1_0),.din(w_dff_A_q4x1fN763_0),.clk(gclk));
	jdff dff_A_tpSB7hXw1_0(.dout(w_dff_A_sZ23K3yj8_0),.din(w_dff_A_tpSB7hXw1_0),.clk(gclk));
	jdff dff_A_sZ23K3yj8_0(.dout(w_dff_A_HA3tr5Lf5_0),.din(w_dff_A_sZ23K3yj8_0),.clk(gclk));
	jdff dff_A_HA3tr5Lf5_0(.dout(w_dff_A_CFnht59b9_0),.din(w_dff_A_HA3tr5Lf5_0),.clk(gclk));
	jdff dff_A_CFnht59b9_0(.dout(w_dff_A_afBxeI4K3_0),.din(w_dff_A_CFnht59b9_0),.clk(gclk));
	jdff dff_A_afBxeI4K3_0(.dout(w_dff_A_Fu7jvWCu8_0),.din(w_dff_A_afBxeI4K3_0),.clk(gclk));
	jdff dff_A_Fu7jvWCu8_0(.dout(w_dff_A_XOdfpkN27_0),.din(w_dff_A_Fu7jvWCu8_0),.clk(gclk));
	jdff dff_A_XOdfpkN27_0(.dout(w_dff_A_q744yOYU7_0),.din(w_dff_A_XOdfpkN27_0),.clk(gclk));
	jdff dff_A_q744yOYU7_0(.dout(w_dff_A_fopuVnDL1_0),.din(w_dff_A_q744yOYU7_0),.clk(gclk));
	jdff dff_A_fopuVnDL1_0(.dout(w_dff_A_BUCk9ajE2_0),.din(w_dff_A_fopuVnDL1_0),.clk(gclk));
	jdff dff_A_BUCk9ajE2_0(.dout(w_dff_A_eccZzo577_0),.din(w_dff_A_BUCk9ajE2_0),.clk(gclk));
	jdff dff_A_eccZzo577_0(.dout(w_dff_A_Dpn8PgxM3_0),.din(w_dff_A_eccZzo577_0),.clk(gclk));
	jdff dff_A_Dpn8PgxM3_0(.dout(w_dff_A_IIoy88BV9_0),.din(w_dff_A_Dpn8PgxM3_0),.clk(gclk));
	jdff dff_A_IIoy88BV9_0(.dout(w_dff_A_fm2Dkq923_0),.din(w_dff_A_IIoy88BV9_0),.clk(gclk));
	jdff dff_A_fm2Dkq923_0(.dout(w_dff_A_9lpUHn895_0),.din(w_dff_A_fm2Dkq923_0),.clk(gclk));
	jdff dff_A_9lpUHn895_0(.dout(w_dff_A_yESDubGW9_0),.din(w_dff_A_9lpUHn895_0),.clk(gclk));
	jdff dff_A_yESDubGW9_0(.dout(w_dff_A_moQNCgH28_0),.din(w_dff_A_yESDubGW9_0),.clk(gclk));
	jdff dff_A_moQNCgH28_0(.dout(G5971gat),.din(w_dff_A_moQNCgH28_0),.clk(gclk));
	jdff dff_A_jiWzWt4L4_2(.dout(w_dff_A_dIDqiBOl1_0),.din(w_dff_A_jiWzWt4L4_2),.clk(gclk));
	jdff dff_A_dIDqiBOl1_0(.dout(w_dff_A_rSzBirvM6_0),.din(w_dff_A_dIDqiBOl1_0),.clk(gclk));
	jdff dff_A_rSzBirvM6_0(.dout(w_dff_A_O4pnc5ZF8_0),.din(w_dff_A_rSzBirvM6_0),.clk(gclk));
	jdff dff_A_O4pnc5ZF8_0(.dout(w_dff_A_yOzwVeDO3_0),.din(w_dff_A_O4pnc5ZF8_0),.clk(gclk));
	jdff dff_A_yOzwVeDO3_0(.dout(w_dff_A_BvvWRKY71_0),.din(w_dff_A_yOzwVeDO3_0),.clk(gclk));
	jdff dff_A_BvvWRKY71_0(.dout(w_dff_A_gZca098h3_0),.din(w_dff_A_BvvWRKY71_0),.clk(gclk));
	jdff dff_A_gZca098h3_0(.dout(w_dff_A_6QztLE7t8_0),.din(w_dff_A_gZca098h3_0),.clk(gclk));
	jdff dff_A_6QztLE7t8_0(.dout(w_dff_A_i4VIAhdq7_0),.din(w_dff_A_6QztLE7t8_0),.clk(gclk));
	jdff dff_A_i4VIAhdq7_0(.dout(w_dff_A_L3JheTda3_0),.din(w_dff_A_i4VIAhdq7_0),.clk(gclk));
	jdff dff_A_L3JheTda3_0(.dout(w_dff_A_xh6BYOtE9_0),.din(w_dff_A_L3JheTda3_0),.clk(gclk));
	jdff dff_A_xh6BYOtE9_0(.dout(w_dff_A_Djx1k5t62_0),.din(w_dff_A_xh6BYOtE9_0),.clk(gclk));
	jdff dff_A_Djx1k5t62_0(.dout(w_dff_A_lslRqdRj0_0),.din(w_dff_A_Djx1k5t62_0),.clk(gclk));
	jdff dff_A_lslRqdRj0_0(.dout(w_dff_A_0fggVyqM5_0),.din(w_dff_A_lslRqdRj0_0),.clk(gclk));
	jdff dff_A_0fggVyqM5_0(.dout(w_dff_A_ysXlWTMC6_0),.din(w_dff_A_0fggVyqM5_0),.clk(gclk));
	jdff dff_A_ysXlWTMC6_0(.dout(w_dff_A_jWZOckRJ8_0),.din(w_dff_A_ysXlWTMC6_0),.clk(gclk));
	jdff dff_A_jWZOckRJ8_0(.dout(w_dff_A_1429AVg40_0),.din(w_dff_A_jWZOckRJ8_0),.clk(gclk));
	jdff dff_A_1429AVg40_0(.dout(w_dff_A_v59ynbEa8_0),.din(w_dff_A_1429AVg40_0),.clk(gclk));
	jdff dff_A_v59ynbEa8_0(.dout(w_dff_A_i2nvBmoI1_0),.din(w_dff_A_v59ynbEa8_0),.clk(gclk));
	jdff dff_A_i2nvBmoI1_0(.dout(w_dff_A_CPDVvugB0_0),.din(w_dff_A_i2nvBmoI1_0),.clk(gclk));
	jdff dff_A_CPDVvugB0_0(.dout(w_dff_A_ib6BZRE60_0),.din(w_dff_A_CPDVvugB0_0),.clk(gclk));
	jdff dff_A_ib6BZRE60_0(.dout(w_dff_A_99663i0F7_0),.din(w_dff_A_ib6BZRE60_0),.clk(gclk));
	jdff dff_A_99663i0F7_0(.dout(w_dff_A_wVoIObD59_0),.din(w_dff_A_99663i0F7_0),.clk(gclk));
	jdff dff_A_wVoIObD59_0(.dout(w_dff_A_dQtWPCFS9_0),.din(w_dff_A_wVoIObD59_0),.clk(gclk));
	jdff dff_A_dQtWPCFS9_0(.dout(w_dff_A_Vo73PJKF6_0),.din(w_dff_A_dQtWPCFS9_0),.clk(gclk));
	jdff dff_A_Vo73PJKF6_0(.dout(w_dff_A_m75zSvps6_0),.din(w_dff_A_Vo73PJKF6_0),.clk(gclk));
	jdff dff_A_m75zSvps6_0(.dout(w_dff_A_iMMfIQ1a0_0),.din(w_dff_A_m75zSvps6_0),.clk(gclk));
	jdff dff_A_iMMfIQ1a0_0(.dout(w_dff_A_iNE2THiY9_0),.din(w_dff_A_iMMfIQ1a0_0),.clk(gclk));
	jdff dff_A_iNE2THiY9_0(.dout(w_dff_A_MukCaABT9_0),.din(w_dff_A_iNE2THiY9_0),.clk(gclk));
	jdff dff_A_MukCaABT9_0(.dout(w_dff_A_tBYGjeYF6_0),.din(w_dff_A_MukCaABT9_0),.clk(gclk));
	jdff dff_A_tBYGjeYF6_0(.dout(G6123gat),.din(w_dff_A_tBYGjeYF6_0),.clk(gclk));
	jdff dff_A_9rj7sGa51_2(.dout(w_dff_A_2rGyWqxD3_0),.din(w_dff_A_9rj7sGa51_2),.clk(gclk));
	jdff dff_A_2rGyWqxD3_0(.dout(w_dff_A_khaU6VDl5_0),.din(w_dff_A_2rGyWqxD3_0),.clk(gclk));
	jdff dff_A_khaU6VDl5_0(.dout(w_dff_A_Oh9wJ5Ih3_0),.din(w_dff_A_khaU6VDl5_0),.clk(gclk));
	jdff dff_A_Oh9wJ5Ih3_0(.dout(w_dff_A_tjVsJESb1_0),.din(w_dff_A_Oh9wJ5Ih3_0),.clk(gclk));
	jdff dff_A_tjVsJESb1_0(.dout(w_dff_A_6pAtnv5w4_0),.din(w_dff_A_tjVsJESb1_0),.clk(gclk));
	jdff dff_A_6pAtnv5w4_0(.dout(w_dff_A_5UoN3ttN7_0),.din(w_dff_A_6pAtnv5w4_0),.clk(gclk));
	jdff dff_A_5UoN3ttN7_0(.dout(w_dff_A_NuwQXmk26_0),.din(w_dff_A_5UoN3ttN7_0),.clk(gclk));
	jdff dff_A_NuwQXmk26_0(.dout(w_dff_A_3s7FdnUw9_0),.din(w_dff_A_NuwQXmk26_0),.clk(gclk));
	jdff dff_A_3s7FdnUw9_0(.dout(w_dff_A_i4t0viAy5_0),.din(w_dff_A_3s7FdnUw9_0),.clk(gclk));
	jdff dff_A_i4t0viAy5_0(.dout(w_dff_A_ir5fzIHe6_0),.din(w_dff_A_i4t0viAy5_0),.clk(gclk));
	jdff dff_A_ir5fzIHe6_0(.dout(w_dff_A_5qOx8dTl2_0),.din(w_dff_A_ir5fzIHe6_0),.clk(gclk));
	jdff dff_A_5qOx8dTl2_0(.dout(w_dff_A_rshkanSd1_0),.din(w_dff_A_5qOx8dTl2_0),.clk(gclk));
	jdff dff_A_rshkanSd1_0(.dout(w_dff_A_ORGcrKS00_0),.din(w_dff_A_rshkanSd1_0),.clk(gclk));
	jdff dff_A_ORGcrKS00_0(.dout(w_dff_A_sfQRTK811_0),.din(w_dff_A_ORGcrKS00_0),.clk(gclk));
	jdff dff_A_sfQRTK811_0(.dout(w_dff_A_X6zOP7RR0_0),.din(w_dff_A_sfQRTK811_0),.clk(gclk));
	jdff dff_A_X6zOP7RR0_0(.dout(w_dff_A_DOx1sjIz1_0),.din(w_dff_A_X6zOP7RR0_0),.clk(gclk));
	jdff dff_A_DOx1sjIz1_0(.dout(w_dff_A_Ibzrda5f4_0),.din(w_dff_A_DOx1sjIz1_0),.clk(gclk));
	jdff dff_A_Ibzrda5f4_0(.dout(w_dff_A_VOZsTIRo4_0),.din(w_dff_A_Ibzrda5f4_0),.clk(gclk));
	jdff dff_A_VOZsTIRo4_0(.dout(w_dff_A_RPMMjNOU7_0),.din(w_dff_A_VOZsTIRo4_0),.clk(gclk));
	jdff dff_A_RPMMjNOU7_0(.dout(w_dff_A_fQGSJnZe1_0),.din(w_dff_A_RPMMjNOU7_0),.clk(gclk));
	jdff dff_A_fQGSJnZe1_0(.dout(w_dff_A_cZDEOagL6_0),.din(w_dff_A_fQGSJnZe1_0),.clk(gclk));
	jdff dff_A_cZDEOagL6_0(.dout(w_dff_A_2RcTKpIL0_0),.din(w_dff_A_cZDEOagL6_0),.clk(gclk));
	jdff dff_A_2RcTKpIL0_0(.dout(w_dff_A_cxaeQwDO2_0),.din(w_dff_A_2RcTKpIL0_0),.clk(gclk));
	jdff dff_A_cxaeQwDO2_0(.dout(w_dff_A_54QgSaxP3_0),.din(w_dff_A_cxaeQwDO2_0),.clk(gclk));
	jdff dff_A_54QgSaxP3_0(.dout(w_dff_A_nLkAw5aV9_0),.din(w_dff_A_54QgSaxP3_0),.clk(gclk));
	jdff dff_A_nLkAw5aV9_0(.dout(w_dff_A_QGqAXeGI1_0),.din(w_dff_A_nLkAw5aV9_0),.clk(gclk));
	jdff dff_A_QGqAXeGI1_0(.dout(w_dff_A_uL2v6ct47_0),.din(w_dff_A_QGqAXeGI1_0),.clk(gclk));
	jdff dff_A_uL2v6ct47_0(.dout(G6150gat),.din(w_dff_A_uL2v6ct47_0),.clk(gclk));
	jdff dff_A_BV07xd3i5_2(.dout(w_dff_A_Xje03yDQ2_0),.din(w_dff_A_BV07xd3i5_2),.clk(gclk));
	jdff dff_A_Xje03yDQ2_0(.dout(w_dff_A_h3zk6Jrn3_0),.din(w_dff_A_Xje03yDQ2_0),.clk(gclk));
	jdff dff_A_h3zk6Jrn3_0(.dout(w_dff_A_E7uRVTQs3_0),.din(w_dff_A_h3zk6Jrn3_0),.clk(gclk));
	jdff dff_A_E7uRVTQs3_0(.dout(w_dff_A_78bz6EeU3_0),.din(w_dff_A_E7uRVTQs3_0),.clk(gclk));
	jdff dff_A_78bz6EeU3_0(.dout(w_dff_A_rk42nJcK8_0),.din(w_dff_A_78bz6EeU3_0),.clk(gclk));
	jdff dff_A_rk42nJcK8_0(.dout(w_dff_A_AuAcb4qo2_0),.din(w_dff_A_rk42nJcK8_0),.clk(gclk));
	jdff dff_A_AuAcb4qo2_0(.dout(w_dff_A_yCzpgHmG8_0),.din(w_dff_A_AuAcb4qo2_0),.clk(gclk));
	jdff dff_A_yCzpgHmG8_0(.dout(w_dff_A_PzbMTrsG7_0),.din(w_dff_A_yCzpgHmG8_0),.clk(gclk));
	jdff dff_A_PzbMTrsG7_0(.dout(w_dff_A_6ilraf8U8_0),.din(w_dff_A_PzbMTrsG7_0),.clk(gclk));
	jdff dff_A_6ilraf8U8_0(.dout(w_dff_A_ERJQ2PEi7_0),.din(w_dff_A_6ilraf8U8_0),.clk(gclk));
	jdff dff_A_ERJQ2PEi7_0(.dout(w_dff_A_Xglk7kj67_0),.din(w_dff_A_ERJQ2PEi7_0),.clk(gclk));
	jdff dff_A_Xglk7kj67_0(.dout(w_dff_A_0VlsmHk84_0),.din(w_dff_A_Xglk7kj67_0),.clk(gclk));
	jdff dff_A_0VlsmHk84_0(.dout(w_dff_A_XQCPMD2T6_0),.din(w_dff_A_0VlsmHk84_0),.clk(gclk));
	jdff dff_A_XQCPMD2T6_0(.dout(w_dff_A_WvWgsSb78_0),.din(w_dff_A_XQCPMD2T6_0),.clk(gclk));
	jdff dff_A_WvWgsSb78_0(.dout(w_dff_A_tiDfvPNe3_0),.din(w_dff_A_WvWgsSb78_0),.clk(gclk));
	jdff dff_A_tiDfvPNe3_0(.dout(w_dff_A_jAU90iYK9_0),.din(w_dff_A_tiDfvPNe3_0),.clk(gclk));
	jdff dff_A_jAU90iYK9_0(.dout(w_dff_A_bhup45yS8_0),.din(w_dff_A_jAU90iYK9_0),.clk(gclk));
	jdff dff_A_bhup45yS8_0(.dout(w_dff_A_TON4qgDI1_0),.din(w_dff_A_bhup45yS8_0),.clk(gclk));
	jdff dff_A_TON4qgDI1_0(.dout(w_dff_A_ALIL2MM26_0),.din(w_dff_A_TON4qgDI1_0),.clk(gclk));
	jdff dff_A_ALIL2MM26_0(.dout(w_dff_A_tpE6xbK47_0),.din(w_dff_A_ALIL2MM26_0),.clk(gclk));
	jdff dff_A_tpE6xbK47_0(.dout(w_dff_A_lQsRyypa8_0),.din(w_dff_A_tpE6xbK47_0),.clk(gclk));
	jdff dff_A_lQsRyypa8_0(.dout(w_dff_A_345vOSOY1_0),.din(w_dff_A_lQsRyypa8_0),.clk(gclk));
	jdff dff_A_345vOSOY1_0(.dout(w_dff_A_yrkWl3Vk0_0),.din(w_dff_A_345vOSOY1_0),.clk(gclk));
	jdff dff_A_yrkWl3Vk0_0(.dout(w_dff_A_mmVyKzX16_0),.din(w_dff_A_yrkWl3Vk0_0),.clk(gclk));
	jdff dff_A_mmVyKzX16_0(.dout(w_dff_A_3h3AmvJd6_0),.din(w_dff_A_mmVyKzX16_0),.clk(gclk));
	jdff dff_A_3h3AmvJd6_0(.dout(G6160gat),.din(w_dff_A_3h3AmvJd6_0),.clk(gclk));
	jdff dff_A_9g6kPTWT1_2(.dout(w_dff_A_yYzAMPrF3_0),.din(w_dff_A_9g6kPTWT1_2),.clk(gclk));
	jdff dff_A_yYzAMPrF3_0(.dout(w_dff_A_FIQC2Vn73_0),.din(w_dff_A_yYzAMPrF3_0),.clk(gclk));
	jdff dff_A_FIQC2Vn73_0(.dout(w_dff_A_2hVNT5ue5_0),.din(w_dff_A_FIQC2Vn73_0),.clk(gclk));
	jdff dff_A_2hVNT5ue5_0(.dout(w_dff_A_IpiW9ErK0_0),.din(w_dff_A_2hVNT5ue5_0),.clk(gclk));
	jdff dff_A_IpiW9ErK0_0(.dout(w_dff_A_X7b5pT8H5_0),.din(w_dff_A_IpiW9ErK0_0),.clk(gclk));
	jdff dff_A_X7b5pT8H5_0(.dout(w_dff_A_KSLVvw7z9_0),.din(w_dff_A_X7b5pT8H5_0),.clk(gclk));
	jdff dff_A_KSLVvw7z9_0(.dout(w_dff_A_rQpk7rlt3_0),.din(w_dff_A_KSLVvw7z9_0),.clk(gclk));
	jdff dff_A_rQpk7rlt3_0(.dout(w_dff_A_PhxBhS2G7_0),.din(w_dff_A_rQpk7rlt3_0),.clk(gclk));
	jdff dff_A_PhxBhS2G7_0(.dout(w_dff_A_ywX332KF8_0),.din(w_dff_A_PhxBhS2G7_0),.clk(gclk));
	jdff dff_A_ywX332KF8_0(.dout(w_dff_A_cV7qit4H8_0),.din(w_dff_A_ywX332KF8_0),.clk(gclk));
	jdff dff_A_cV7qit4H8_0(.dout(w_dff_A_1Gzg5Pmu1_0),.din(w_dff_A_cV7qit4H8_0),.clk(gclk));
	jdff dff_A_1Gzg5Pmu1_0(.dout(w_dff_A_OrmdwKwG3_0),.din(w_dff_A_1Gzg5Pmu1_0),.clk(gclk));
	jdff dff_A_OrmdwKwG3_0(.dout(w_dff_A_kzCWQrg84_0),.din(w_dff_A_OrmdwKwG3_0),.clk(gclk));
	jdff dff_A_kzCWQrg84_0(.dout(w_dff_A_jgz46Cau5_0),.din(w_dff_A_kzCWQrg84_0),.clk(gclk));
	jdff dff_A_jgz46Cau5_0(.dout(w_dff_A_XuK0fD9s2_0),.din(w_dff_A_jgz46Cau5_0),.clk(gclk));
	jdff dff_A_XuK0fD9s2_0(.dout(w_dff_A_PioRJHem1_0),.din(w_dff_A_XuK0fD9s2_0),.clk(gclk));
	jdff dff_A_PioRJHem1_0(.dout(w_dff_A_Q8l92rz44_0),.din(w_dff_A_PioRJHem1_0),.clk(gclk));
	jdff dff_A_Q8l92rz44_0(.dout(w_dff_A_zJnz07Xw2_0),.din(w_dff_A_Q8l92rz44_0),.clk(gclk));
	jdff dff_A_zJnz07Xw2_0(.dout(w_dff_A_lmS6NKWW0_0),.din(w_dff_A_zJnz07Xw2_0),.clk(gclk));
	jdff dff_A_lmS6NKWW0_0(.dout(w_dff_A_2aZ1pcVh3_0),.din(w_dff_A_lmS6NKWW0_0),.clk(gclk));
	jdff dff_A_2aZ1pcVh3_0(.dout(w_dff_A_pCuekJw62_0),.din(w_dff_A_2aZ1pcVh3_0),.clk(gclk));
	jdff dff_A_pCuekJw62_0(.dout(w_dff_A_08N4RNqu0_0),.din(w_dff_A_pCuekJw62_0),.clk(gclk));
	jdff dff_A_08N4RNqu0_0(.dout(w_dff_A_bQNov0F77_0),.din(w_dff_A_08N4RNqu0_0),.clk(gclk));
	jdff dff_A_bQNov0F77_0(.dout(w_dff_A_ZwLS8Cc48_0),.din(w_dff_A_bQNov0F77_0),.clk(gclk));
	jdff dff_A_ZwLS8Cc48_0(.dout(G6170gat),.din(w_dff_A_ZwLS8Cc48_0),.clk(gclk));
	jdff dff_A_fM5Zpmhi3_2(.dout(w_dff_A_LW1HRYzu7_0),.din(w_dff_A_fM5Zpmhi3_2),.clk(gclk));
	jdff dff_A_LW1HRYzu7_0(.dout(w_dff_A_bML1SCrV3_0),.din(w_dff_A_LW1HRYzu7_0),.clk(gclk));
	jdff dff_A_bML1SCrV3_0(.dout(w_dff_A_KkdrC1ro0_0),.din(w_dff_A_bML1SCrV3_0),.clk(gclk));
	jdff dff_A_KkdrC1ro0_0(.dout(w_dff_A_nOBiBduh0_0),.din(w_dff_A_KkdrC1ro0_0),.clk(gclk));
	jdff dff_A_nOBiBduh0_0(.dout(w_dff_A_tff23dYW3_0),.din(w_dff_A_nOBiBduh0_0),.clk(gclk));
	jdff dff_A_tff23dYW3_0(.dout(w_dff_A_Pk9lk0Yd8_0),.din(w_dff_A_tff23dYW3_0),.clk(gclk));
	jdff dff_A_Pk9lk0Yd8_0(.dout(w_dff_A_Wxs6fsYc3_0),.din(w_dff_A_Pk9lk0Yd8_0),.clk(gclk));
	jdff dff_A_Wxs6fsYc3_0(.dout(w_dff_A_ZEZOWqKD0_0),.din(w_dff_A_Wxs6fsYc3_0),.clk(gclk));
	jdff dff_A_ZEZOWqKD0_0(.dout(w_dff_A_rKRik5gr8_0),.din(w_dff_A_ZEZOWqKD0_0),.clk(gclk));
	jdff dff_A_rKRik5gr8_0(.dout(w_dff_A_C5cdIUN94_0),.din(w_dff_A_rKRik5gr8_0),.clk(gclk));
	jdff dff_A_C5cdIUN94_0(.dout(w_dff_A_z9CzoWJW0_0),.din(w_dff_A_C5cdIUN94_0),.clk(gclk));
	jdff dff_A_z9CzoWJW0_0(.dout(w_dff_A_oOn6l4V28_0),.din(w_dff_A_z9CzoWJW0_0),.clk(gclk));
	jdff dff_A_oOn6l4V28_0(.dout(w_dff_A_Xw7WBAyt0_0),.din(w_dff_A_oOn6l4V28_0),.clk(gclk));
	jdff dff_A_Xw7WBAyt0_0(.dout(w_dff_A_wgknJs2g1_0),.din(w_dff_A_Xw7WBAyt0_0),.clk(gclk));
	jdff dff_A_wgknJs2g1_0(.dout(w_dff_A_7yNV4YqP2_0),.din(w_dff_A_wgknJs2g1_0),.clk(gclk));
	jdff dff_A_7yNV4YqP2_0(.dout(w_dff_A_fcAL6fWU0_0),.din(w_dff_A_7yNV4YqP2_0),.clk(gclk));
	jdff dff_A_fcAL6fWU0_0(.dout(w_dff_A_EDALEDbp9_0),.din(w_dff_A_fcAL6fWU0_0),.clk(gclk));
	jdff dff_A_EDALEDbp9_0(.dout(w_dff_A_xzFzyeM54_0),.din(w_dff_A_EDALEDbp9_0),.clk(gclk));
	jdff dff_A_xzFzyeM54_0(.dout(w_dff_A_sQmwGAnI9_0),.din(w_dff_A_xzFzyeM54_0),.clk(gclk));
	jdff dff_A_sQmwGAnI9_0(.dout(w_dff_A_bFpczJJL5_0),.din(w_dff_A_sQmwGAnI9_0),.clk(gclk));
	jdff dff_A_bFpczJJL5_0(.dout(w_dff_A_mLs2v7d82_0),.din(w_dff_A_bFpczJJL5_0),.clk(gclk));
	jdff dff_A_mLs2v7d82_0(.dout(w_dff_A_Aa8iMiQH0_0),.din(w_dff_A_mLs2v7d82_0),.clk(gclk));
	jdff dff_A_Aa8iMiQH0_0(.dout(G6180gat),.din(w_dff_A_Aa8iMiQH0_0),.clk(gclk));
	jdff dff_A_ErYJJyU15_2(.dout(w_dff_A_oWT8ksqJ6_0),.din(w_dff_A_ErYJJyU15_2),.clk(gclk));
	jdff dff_A_oWT8ksqJ6_0(.dout(w_dff_A_2T3mfj314_0),.din(w_dff_A_oWT8ksqJ6_0),.clk(gclk));
	jdff dff_A_2T3mfj314_0(.dout(w_dff_A_djmyjo4D4_0),.din(w_dff_A_2T3mfj314_0),.clk(gclk));
	jdff dff_A_djmyjo4D4_0(.dout(w_dff_A_lVAzPl6C8_0),.din(w_dff_A_djmyjo4D4_0),.clk(gclk));
	jdff dff_A_lVAzPl6C8_0(.dout(w_dff_A_lFx7YcLt3_0),.din(w_dff_A_lVAzPl6C8_0),.clk(gclk));
	jdff dff_A_lFx7YcLt3_0(.dout(w_dff_A_zRZgQr203_0),.din(w_dff_A_lFx7YcLt3_0),.clk(gclk));
	jdff dff_A_zRZgQr203_0(.dout(w_dff_A_1vdkRwWs1_0),.din(w_dff_A_zRZgQr203_0),.clk(gclk));
	jdff dff_A_1vdkRwWs1_0(.dout(w_dff_A_2d2Tid294_0),.din(w_dff_A_1vdkRwWs1_0),.clk(gclk));
	jdff dff_A_2d2Tid294_0(.dout(w_dff_A_PoSyKR9j0_0),.din(w_dff_A_2d2Tid294_0),.clk(gclk));
	jdff dff_A_PoSyKR9j0_0(.dout(w_dff_A_5Xz4HYIk4_0),.din(w_dff_A_PoSyKR9j0_0),.clk(gclk));
	jdff dff_A_5Xz4HYIk4_0(.dout(w_dff_A_8aKbN7V35_0),.din(w_dff_A_5Xz4HYIk4_0),.clk(gclk));
	jdff dff_A_8aKbN7V35_0(.dout(w_dff_A_MdfagJWI4_0),.din(w_dff_A_8aKbN7V35_0),.clk(gclk));
	jdff dff_A_MdfagJWI4_0(.dout(w_dff_A_LooAqoFO0_0),.din(w_dff_A_MdfagJWI4_0),.clk(gclk));
	jdff dff_A_LooAqoFO0_0(.dout(w_dff_A_lmTmNccP0_0),.din(w_dff_A_LooAqoFO0_0),.clk(gclk));
	jdff dff_A_lmTmNccP0_0(.dout(w_dff_A_Ro6I1P4M6_0),.din(w_dff_A_lmTmNccP0_0),.clk(gclk));
	jdff dff_A_Ro6I1P4M6_0(.dout(w_dff_A_0Uy8eLJh2_0),.din(w_dff_A_Ro6I1P4M6_0),.clk(gclk));
	jdff dff_A_0Uy8eLJh2_0(.dout(w_dff_A_TDBduI0B3_0),.din(w_dff_A_0Uy8eLJh2_0),.clk(gclk));
	jdff dff_A_TDBduI0B3_0(.dout(w_dff_A_GbBGdva52_0),.din(w_dff_A_TDBduI0B3_0),.clk(gclk));
	jdff dff_A_GbBGdva52_0(.dout(w_dff_A_sPKB2ABh1_0),.din(w_dff_A_GbBGdva52_0),.clk(gclk));
	jdff dff_A_sPKB2ABh1_0(.dout(w_dff_A_lkA1ZPkL1_0),.din(w_dff_A_sPKB2ABh1_0),.clk(gclk));
	jdff dff_A_lkA1ZPkL1_0(.dout(G6190gat),.din(w_dff_A_lkA1ZPkL1_0),.clk(gclk));
	jdff dff_A_AzVrOdhu4_2(.dout(w_dff_A_uWjJLX7o1_0),.din(w_dff_A_AzVrOdhu4_2),.clk(gclk));
	jdff dff_A_uWjJLX7o1_0(.dout(w_dff_A_1mrElvGu7_0),.din(w_dff_A_uWjJLX7o1_0),.clk(gclk));
	jdff dff_A_1mrElvGu7_0(.dout(w_dff_A_rCc925j66_0),.din(w_dff_A_1mrElvGu7_0),.clk(gclk));
	jdff dff_A_rCc925j66_0(.dout(w_dff_A_x6hk4h9o8_0),.din(w_dff_A_rCc925j66_0),.clk(gclk));
	jdff dff_A_x6hk4h9o8_0(.dout(w_dff_A_IlsXXzrE7_0),.din(w_dff_A_x6hk4h9o8_0),.clk(gclk));
	jdff dff_A_IlsXXzrE7_0(.dout(w_dff_A_WGstDMbS8_0),.din(w_dff_A_IlsXXzrE7_0),.clk(gclk));
	jdff dff_A_WGstDMbS8_0(.dout(w_dff_A_uKI2OQuO0_0),.din(w_dff_A_WGstDMbS8_0),.clk(gclk));
	jdff dff_A_uKI2OQuO0_0(.dout(w_dff_A_cpKHbzom4_0),.din(w_dff_A_uKI2OQuO0_0),.clk(gclk));
	jdff dff_A_cpKHbzom4_0(.dout(w_dff_A_A7fIhCAC5_0),.din(w_dff_A_cpKHbzom4_0),.clk(gclk));
	jdff dff_A_A7fIhCAC5_0(.dout(w_dff_A_ivY0gT9Z9_0),.din(w_dff_A_A7fIhCAC5_0),.clk(gclk));
	jdff dff_A_ivY0gT9Z9_0(.dout(w_dff_A_T7xeaIm81_0),.din(w_dff_A_ivY0gT9Z9_0),.clk(gclk));
	jdff dff_A_T7xeaIm81_0(.dout(w_dff_A_W3a0RCIO4_0),.din(w_dff_A_T7xeaIm81_0),.clk(gclk));
	jdff dff_A_W3a0RCIO4_0(.dout(w_dff_A_odJUDopP1_0),.din(w_dff_A_W3a0RCIO4_0),.clk(gclk));
	jdff dff_A_odJUDopP1_0(.dout(w_dff_A_Yqy7GRQy4_0),.din(w_dff_A_odJUDopP1_0),.clk(gclk));
	jdff dff_A_Yqy7GRQy4_0(.dout(w_dff_A_2YDdMQ9S2_0),.din(w_dff_A_Yqy7GRQy4_0),.clk(gclk));
	jdff dff_A_2YDdMQ9S2_0(.dout(w_dff_A_1BOzJxMq6_0),.din(w_dff_A_2YDdMQ9S2_0),.clk(gclk));
	jdff dff_A_1BOzJxMq6_0(.dout(w_dff_A_1B5UmdWk3_0),.din(w_dff_A_1BOzJxMq6_0),.clk(gclk));
	jdff dff_A_1B5UmdWk3_0(.dout(w_dff_A_jAJg68wu4_0),.din(w_dff_A_1B5UmdWk3_0),.clk(gclk));
	jdff dff_A_jAJg68wu4_0(.dout(G6200gat),.din(w_dff_A_jAJg68wu4_0),.clk(gclk));
	jdff dff_A_bjPY08b41_2(.dout(w_dff_A_2jBrYvVK0_0),.din(w_dff_A_bjPY08b41_2),.clk(gclk));
	jdff dff_A_2jBrYvVK0_0(.dout(w_dff_A_sa08IdHG5_0),.din(w_dff_A_2jBrYvVK0_0),.clk(gclk));
	jdff dff_A_sa08IdHG5_0(.dout(w_dff_A_3TWzhnyY7_0),.din(w_dff_A_sa08IdHG5_0),.clk(gclk));
	jdff dff_A_3TWzhnyY7_0(.dout(w_dff_A_tCf1CIk89_0),.din(w_dff_A_3TWzhnyY7_0),.clk(gclk));
	jdff dff_A_tCf1CIk89_0(.dout(w_dff_A_2zFm7QTR3_0),.din(w_dff_A_tCf1CIk89_0),.clk(gclk));
	jdff dff_A_2zFm7QTR3_0(.dout(w_dff_A_LkHqktZR0_0),.din(w_dff_A_2zFm7QTR3_0),.clk(gclk));
	jdff dff_A_LkHqktZR0_0(.dout(w_dff_A_nRIk1TJg3_0),.din(w_dff_A_LkHqktZR0_0),.clk(gclk));
	jdff dff_A_nRIk1TJg3_0(.dout(w_dff_A_ncE8H9nG1_0),.din(w_dff_A_nRIk1TJg3_0),.clk(gclk));
	jdff dff_A_ncE8H9nG1_0(.dout(w_dff_A_LVRb8WOa1_0),.din(w_dff_A_ncE8H9nG1_0),.clk(gclk));
	jdff dff_A_LVRb8WOa1_0(.dout(w_dff_A_XedGkZsb1_0),.din(w_dff_A_LVRb8WOa1_0),.clk(gclk));
	jdff dff_A_XedGkZsb1_0(.dout(w_dff_A_ucfMcgXy8_0),.din(w_dff_A_XedGkZsb1_0),.clk(gclk));
	jdff dff_A_ucfMcgXy8_0(.dout(w_dff_A_H3XSbEDj4_0),.din(w_dff_A_ucfMcgXy8_0),.clk(gclk));
	jdff dff_A_H3XSbEDj4_0(.dout(w_dff_A_vgVmitma8_0),.din(w_dff_A_H3XSbEDj4_0),.clk(gclk));
	jdff dff_A_vgVmitma8_0(.dout(w_dff_A_o7EufxxD1_0),.din(w_dff_A_vgVmitma8_0),.clk(gclk));
	jdff dff_A_o7EufxxD1_0(.dout(w_dff_A_0I8W9pMw5_0),.din(w_dff_A_o7EufxxD1_0),.clk(gclk));
	jdff dff_A_0I8W9pMw5_0(.dout(w_dff_A_19jiXv2I0_0),.din(w_dff_A_0I8W9pMw5_0),.clk(gclk));
	jdff dff_A_19jiXv2I0_0(.dout(G6210gat),.din(w_dff_A_19jiXv2I0_0),.clk(gclk));
	jdff dff_A_DmqhRz3o5_2(.dout(w_dff_A_DgWwyF5U2_0),.din(w_dff_A_DmqhRz3o5_2),.clk(gclk));
	jdff dff_A_DgWwyF5U2_0(.dout(w_dff_A_SAeZcok29_0),.din(w_dff_A_DgWwyF5U2_0),.clk(gclk));
	jdff dff_A_SAeZcok29_0(.dout(w_dff_A_zxbBAUMZ4_0),.din(w_dff_A_SAeZcok29_0),.clk(gclk));
	jdff dff_A_zxbBAUMZ4_0(.dout(w_dff_A_nmTVdO7T7_0),.din(w_dff_A_zxbBAUMZ4_0),.clk(gclk));
	jdff dff_A_nmTVdO7T7_0(.dout(w_dff_A_FDfXMotY6_0),.din(w_dff_A_nmTVdO7T7_0),.clk(gclk));
	jdff dff_A_FDfXMotY6_0(.dout(w_dff_A_dBCUMnWG3_0),.din(w_dff_A_FDfXMotY6_0),.clk(gclk));
	jdff dff_A_dBCUMnWG3_0(.dout(w_dff_A_m4crRSXh5_0),.din(w_dff_A_dBCUMnWG3_0),.clk(gclk));
	jdff dff_A_m4crRSXh5_0(.dout(w_dff_A_vJ6qf8iR8_0),.din(w_dff_A_m4crRSXh5_0),.clk(gclk));
	jdff dff_A_vJ6qf8iR8_0(.dout(w_dff_A_95jBNy331_0),.din(w_dff_A_vJ6qf8iR8_0),.clk(gclk));
	jdff dff_A_95jBNy331_0(.dout(w_dff_A_dcPMNw3X9_0),.din(w_dff_A_95jBNy331_0),.clk(gclk));
	jdff dff_A_dcPMNw3X9_0(.dout(w_dff_A_yFIo1lZg7_0),.din(w_dff_A_dcPMNw3X9_0),.clk(gclk));
	jdff dff_A_yFIo1lZg7_0(.dout(w_dff_A_aNlcE4804_0),.din(w_dff_A_yFIo1lZg7_0),.clk(gclk));
	jdff dff_A_aNlcE4804_0(.dout(w_dff_A_39Q1XvvA2_0),.din(w_dff_A_aNlcE4804_0),.clk(gclk));
	jdff dff_A_39Q1XvvA2_0(.dout(w_dff_A_U0Pke4dh7_0),.din(w_dff_A_39Q1XvvA2_0),.clk(gclk));
	jdff dff_A_U0Pke4dh7_0(.dout(G6220gat),.din(w_dff_A_U0Pke4dh7_0),.clk(gclk));
	jdff dff_A_Gu5QXbuJ7_2(.dout(w_dff_A_kFYN7hz33_0),.din(w_dff_A_Gu5QXbuJ7_2),.clk(gclk));
	jdff dff_A_kFYN7hz33_0(.dout(w_dff_A_emrWU3Oz4_0),.din(w_dff_A_kFYN7hz33_0),.clk(gclk));
	jdff dff_A_emrWU3Oz4_0(.dout(w_dff_A_LdM5n9v23_0),.din(w_dff_A_emrWU3Oz4_0),.clk(gclk));
	jdff dff_A_LdM5n9v23_0(.dout(w_dff_A_x07z2FN34_0),.din(w_dff_A_LdM5n9v23_0),.clk(gclk));
	jdff dff_A_x07z2FN34_0(.dout(w_dff_A_BzDGGaaP5_0),.din(w_dff_A_x07z2FN34_0),.clk(gclk));
	jdff dff_A_BzDGGaaP5_0(.dout(w_dff_A_WoQ0EsWS5_0),.din(w_dff_A_BzDGGaaP5_0),.clk(gclk));
	jdff dff_A_WoQ0EsWS5_0(.dout(w_dff_A_9KzTNYGp0_0),.din(w_dff_A_WoQ0EsWS5_0),.clk(gclk));
	jdff dff_A_9KzTNYGp0_0(.dout(w_dff_A_WiLPlZry6_0),.din(w_dff_A_9KzTNYGp0_0),.clk(gclk));
	jdff dff_A_WiLPlZry6_0(.dout(w_dff_A_9g4tYXBj5_0),.din(w_dff_A_WiLPlZry6_0),.clk(gclk));
	jdff dff_A_9g4tYXBj5_0(.dout(w_dff_A_aqwKUeEP2_0),.din(w_dff_A_9g4tYXBj5_0),.clk(gclk));
	jdff dff_A_aqwKUeEP2_0(.dout(w_dff_A_37BxLqwc4_0),.din(w_dff_A_aqwKUeEP2_0),.clk(gclk));
	jdff dff_A_37BxLqwc4_0(.dout(w_dff_A_TkdbBbfy6_0),.din(w_dff_A_37BxLqwc4_0),.clk(gclk));
	jdff dff_A_TkdbBbfy6_0(.dout(G6230gat),.din(w_dff_A_TkdbBbfy6_0),.clk(gclk));
	jdff dff_A_TOoGb41g9_2(.dout(w_dff_A_OeQAHLUb8_0),.din(w_dff_A_TOoGb41g9_2),.clk(gclk));
	jdff dff_A_OeQAHLUb8_0(.dout(w_dff_A_IGYDdBTf8_0),.din(w_dff_A_OeQAHLUb8_0),.clk(gclk));
	jdff dff_A_IGYDdBTf8_0(.dout(w_dff_A_qc1UiXSs2_0),.din(w_dff_A_IGYDdBTf8_0),.clk(gclk));
	jdff dff_A_qc1UiXSs2_0(.dout(w_dff_A_aGtVqjBI9_0),.din(w_dff_A_qc1UiXSs2_0),.clk(gclk));
	jdff dff_A_aGtVqjBI9_0(.dout(w_dff_A_cXTYmrrz6_0),.din(w_dff_A_aGtVqjBI9_0),.clk(gclk));
	jdff dff_A_cXTYmrrz6_0(.dout(w_dff_A_U4Fj0e5N2_0),.din(w_dff_A_cXTYmrrz6_0),.clk(gclk));
	jdff dff_A_U4Fj0e5N2_0(.dout(w_dff_A_KSiVsY284_0),.din(w_dff_A_U4Fj0e5N2_0),.clk(gclk));
	jdff dff_A_KSiVsY284_0(.dout(w_dff_A_M1cFi3QN5_0),.din(w_dff_A_KSiVsY284_0),.clk(gclk));
	jdff dff_A_M1cFi3QN5_0(.dout(w_dff_A_Yk6xc5Rb3_0),.din(w_dff_A_M1cFi3QN5_0),.clk(gclk));
	jdff dff_A_Yk6xc5Rb3_0(.dout(w_dff_A_2HGFNCac5_0),.din(w_dff_A_Yk6xc5Rb3_0),.clk(gclk));
	jdff dff_A_2HGFNCac5_0(.dout(G6240gat),.din(w_dff_A_2HGFNCac5_0),.clk(gclk));
	jdff dff_A_CFydfasb0_2(.dout(w_dff_A_6gjinRhx1_0),.din(w_dff_A_CFydfasb0_2),.clk(gclk));
	jdff dff_A_6gjinRhx1_0(.dout(w_dff_A_ItJXiioD4_0),.din(w_dff_A_6gjinRhx1_0),.clk(gclk));
	jdff dff_A_ItJXiioD4_0(.dout(w_dff_A_QN6EevqU0_0),.din(w_dff_A_ItJXiioD4_0),.clk(gclk));
	jdff dff_A_QN6EevqU0_0(.dout(w_dff_A_YXvjz82R3_0),.din(w_dff_A_QN6EevqU0_0),.clk(gclk));
	jdff dff_A_YXvjz82R3_0(.dout(w_dff_A_j5ZdIJbF2_0),.din(w_dff_A_YXvjz82R3_0),.clk(gclk));
	jdff dff_A_j5ZdIJbF2_0(.dout(w_dff_A_WpW4oPeJ4_0),.din(w_dff_A_j5ZdIJbF2_0),.clk(gclk));
	jdff dff_A_WpW4oPeJ4_0(.dout(w_dff_A_UteeaXOf7_0),.din(w_dff_A_WpW4oPeJ4_0),.clk(gclk));
	jdff dff_A_UteeaXOf7_0(.dout(w_dff_A_bL2kAIyG7_0),.din(w_dff_A_UteeaXOf7_0),.clk(gclk));
	jdff dff_A_bL2kAIyG7_0(.dout(G6250gat),.din(w_dff_A_bL2kAIyG7_0),.clk(gclk));
	jdff dff_A_J0Xe6gJm8_2(.dout(w_dff_A_7w5cS6BW1_0),.din(w_dff_A_J0Xe6gJm8_2),.clk(gclk));
	jdff dff_A_7w5cS6BW1_0(.dout(w_dff_A_4bAsWJVA0_0),.din(w_dff_A_7w5cS6BW1_0),.clk(gclk));
	jdff dff_A_4bAsWJVA0_0(.dout(w_dff_A_gwJiPMT72_0),.din(w_dff_A_4bAsWJVA0_0),.clk(gclk));
	jdff dff_A_gwJiPMT72_0(.dout(w_dff_A_hFKyAnbg6_0),.din(w_dff_A_gwJiPMT72_0),.clk(gclk));
	jdff dff_A_hFKyAnbg6_0(.dout(w_dff_A_KKdOJg614_0),.din(w_dff_A_hFKyAnbg6_0),.clk(gclk));
	jdff dff_A_KKdOJg614_0(.dout(w_dff_A_N4F2ehqO5_0),.din(w_dff_A_KKdOJg614_0),.clk(gclk));
	jdff dff_A_N4F2ehqO5_0(.dout(G6260gat),.din(w_dff_A_N4F2ehqO5_0),.clk(gclk));
	jdff dff_A_kkcMHLRb7_2(.dout(w_dff_A_tvTGKUOh1_0),.din(w_dff_A_kkcMHLRb7_2),.clk(gclk));
	jdff dff_A_tvTGKUOh1_0(.dout(w_dff_A_SVrbNEq45_0),.din(w_dff_A_tvTGKUOh1_0),.clk(gclk));
	jdff dff_A_SVrbNEq45_0(.dout(w_dff_A_zOepyAGb0_0),.din(w_dff_A_SVrbNEq45_0),.clk(gclk));
	jdff dff_A_zOepyAGb0_0(.dout(w_dff_A_txUfsu520_0),.din(w_dff_A_zOepyAGb0_0),.clk(gclk));
	jdff dff_A_txUfsu520_0(.dout(G6270gat),.din(w_dff_A_txUfsu520_0),.clk(gclk));
	jdff dff_A_2YEfK94H7_2(.dout(w_dff_A_XH2YOm5t7_0),.din(w_dff_A_2YEfK94H7_2),.clk(gclk));
	jdff dff_A_XH2YOm5t7_0(.dout(w_dff_A_TVk2CzHW5_0),.din(w_dff_A_XH2YOm5t7_0),.clk(gclk));
	jdff dff_A_TVk2CzHW5_0(.dout(G6280gat),.din(w_dff_A_TVk2CzHW5_0),.clk(gclk));
	jdff dff_A_rdgwxBzJ1_2(.dout(G6288gat),.din(w_dff_A_rdgwxBzJ1_2),.clk(gclk));
endmodule

