module gf_c5315(G4115, G4092, G4089, G4087, G3724, G3550, G3548, G3546, G2824, G2358, G1694, G1690, G1689, G562, G552, G545, G534, G468, G435, G4091, G479, G422, G3173, G411, G556, G400, G523, G386, G373, G369, G366, G361, G348, G254, G127, G121, G119, G167, G114, G191, G112, G164, G389, G106, G103, G152, G117, G242, G100, G161, G118, G87, G97, G88, G146, G86, G83, G549, G82, G307, G3717, G46, G245, G358, G265, G11, G27, G123, G54, G116, G374, G43, G26, G31, G1497, G332, G218, G299, G372, G1, G128, G73, G14, G3552, G122, G248, G120, G109, G4, G23, G113, G76, G145, G34, G91, G49, G225, G64, G131, G351, G126, G37, G94, G149, G81, G226, G1691, G61, G80, G79, G280, G20, G67, G308, G503, G241, G70, G130, G200, G559, G132, G135, G188, G206, G209, G335, G136, G137, G141, G140, G197, G490, G155, G185, G158, G315, G170, G129, G17, G173, G176, G179, G182, G273, G293, G194, G210, G457, G53, G233, G234, G251, G289, G257, G514, G264, G288, G2174, G292, G302, G4090, G25, G316, G4088, G272, G323, G24, G203, G40, G324, G52, G331, G446, G281, G217, G338, G115, G341, G658, G807, G843, G685, G679, G654, G651, G648, G645, G742, G727, G869, G712, G854, G782, G826, G882, G818, G702, G813, G699, G696, G824, G670, G792, G762, G752, G693, G661, G1000, G998, G877, G873, G664, G871, G859, G834, G606, G787, G921, G828, G973, G939, G867, G851, G850, G865, G715, G757, G612, G849, G623, G634, G777, G772, G861, G603, G656, G767, G848, G875, G845, G747, G298, G636, G591, G601, G887, G599, G926, G688, G810, G600, G642, G809, G836, G611, G585, G949, G604, G667, G923, G144, G602, G832, G993, G594, G889, G1004, G892, G838, G802, G575, G1002, G978, G797, G593, G704, G717, G820, G737, G639, G732, G847, G673, G863, G707, G830, G632, G690, G598, G610, G682, G676, G588, G621, G615, G629, G626, G722, G815, G618, G822);
    input G4115, G4092, G4089, G4087, G3724, G3550, G3548, G3546, G2824, G2358, G1694, G1690, G1689, G562, G552, G545, G534, G468, G435, G4091, G479, G422, G3173, G411, G556, G400, G523, G386, G373, G369, G366, G361, G348, G254, G127, G121, G119, G167, G114, G191, G112, G164, G389, G106, G103, G152, G117, G242, G100, G161, G118, G87, G97, G88, G146, G86, G83, G549, G82, G307, G3717, G46, G245, G358, G265, G11, G27, G123, G54, G116, G374, G43, G26, G31, G1497, G332, G218, G299, G372, G1, G128, G73, G14, G3552, G122, G248, G120, G109, G4, G23, G113, G76, G145, G34, G91, G49, G225, G64, G131, G351, G126, G37, G94, G149, G81, G226, G1691, G61, G80, G79, G280, G20, G67, G308, G503, G241, G70, G130, G200, G559, G132, G135, G188, G206, G209, G335, G136, G137, G141, G140, G197, G490, G155, G185, G158, G315, G170, G129, G17, G173, G176, G179, G182, G273, G293, G194, G210, G457, G53, G233, G234, G251, G289, G257, G514, G264, G288, G2174, G292, G302, G4090, G25, G316, G4088, G272, G323, G24, G203, G40, G324, G52, G331, G446, G281, G217, G338, G115, G341;
    output G658, G807, G843, G685, G679, G654, G651, G648, G645, G742, G727, G869, G712, G854, G782, G826, G882, G818, G702, G813, G699, G696, G824, G670, G792, G762, G752, G693, G661, G1000, G998, G877, G873, G664, G871, G859, G834, G606, G787, G921, G828, G973, G939, G867, G851, G850, G865, G715, G757, G612, G849, G623, G634, G777, G772, G861, G603, G656, G767, G848, G875, G845, G747, G298, G636, G591, G601, G887, G599, G926, G688, G810, G600, G642, G809, G836, G611, G585, G949, G604, G667, G923, G144, G602, G832, G993, G594, G889, G1004, G892, G838, G802, G575, G1002, G978, G797, G593, G704, G717, G820, G737, G639, G732, G847, G673, G863, G707, G830, G632, G690, G598, G610, G682, G676, G588, G621, G615, G629, G626, G722, G815, G618, G822;
    wire n303;
    wire n306;
    wire n309;
    wire n313;
    wire n316;
    wire n319;
    wire n322;
    wire n326;
    wire n329;
    wire n332;
    wire n335;
    wire n338;
    wire n342;
    wire n345;
    wire n349;
    wire n352;
    wire n356;
    wire n360;
    wire n363;
    wire n366;
    wire n369;
    wire n373;
    wire n377;
    wire n380;
    wire n383;
    wire n386;
    wire n390;
    wire n393;
    wire n397;
    wire n401;
    wire n405;
    wire n408;
    wire n412;
    wire n415;
    wire n419;
    wire n423;
    wire n427;
    wire n430;
    wire n434;
    wire n438;
    wire n442;
    wire n446;
    wire n450;
    wire n454;
    wire n458;
    wire n462;
    wire n466;
    wire n470;
    wire n474;
    wire n478;
    wire n482;
    wire n486;
    wire n490;
    wire n494;
    wire n498;
    wire n502;
    wire n506;
    wire n510;
    wire n514;
    wire n518;
    wire n521;
    wire n524;
    wire n528;
    wire n532;
    wire n535;
    wire n538;
    wire n541;
    wire n545;
    wire n548;
    wire n552;
    wire n556;
    wire n559;
    wire n563;
    wire n566;
    wire n569;
    wire n573;
    wire n576;
    wire n579;
    wire n583;
    wire n587;
    wire n591;
    wire n595;
    wire n599;
    wire n603;
    wire n607;
    wire n611;
    wire n614;
    wire n618;
    wire n621;
    wire n625;
    wire n629;
    wire n633;
    wire n637;
    wire n641;
    wire n645;
    wire n649;
    wire n653;
    wire n657;
    wire n661;
    wire n665;
    wire n668;
    wire n671;
    wire n675;
    wire n679;
    wire n683;
    wire n686;
    wire n690;
    wire n693;
    wire n697;
    wire n701;
    wire n705;
    wire n709;
    wire n713;
    wire n716;
    wire n719;
    wire n723;
    wire n727;
    wire n731;
    wire n735;
    wire n739;
    wire n743;
    wire n747;
    wire n751;
    wire n755;
    wire n758;
    wire n762;
    wire n766;
    wire n770;
    wire n773;
    wire n777;
    wire n781;
    wire n785;
    wire n788;
    wire n792;
    wire n795;
    wire n799;
    wire n802;
    wire n806;
    wire n810;
    wire n814;
    wire n818;
    wire n822;
    wire n826;
    wire n830;
    wire n834;
    wire n838;
    wire n842;
    wire n846;
    wire n849;
    wire n853;
    wire n856;
    wire n860;
    wire n864;
    wire n868;
    wire n872;
    wire n876;
    wire n880;
    wire n884;
    wire n888;
    wire n891;
    wire n895;
    wire n898;
    wire n902;
    wire n906;
    wire n910;
    wire n914;
    wire n918;
    wire n922;
    wire n926;
    wire n930;
    wire n933;
    wire n937;
    wire n940;
    wire n944;
    wire n948;
    wire n952;
    wire n956;
    wire n960;
    wire n964;
    wire n968;
    wire n972;
    wire n976;
    wire n979;
    wire n983;
    wire n986;
    wire n990;
    wire n994;
    wire n998;
    wire n1002;
    wire n1006;
    wire n1010;
    wire n1014;
    wire n1018;
    wire n1021;
    wire n1025;
    wire n1028;
    wire n1032;
    wire n1036;
    wire n1040;
    wire n1044;
    wire n1048;
    wire n1052;
    wire n1056;
    wire n1060;
    wire n1064;
    wire n1068;
    wire n1071;
    wire n1075;
    wire n1078;
    wire n1082;
    wire n1086;
    wire n1090;
    wire n1094;
    wire n1098;
    wire n1102;
    wire n1106;
    wire n1110;
    wire n1113;
    wire n1117;
    wire n1120;
    wire n1124;
    wire n1128;
    wire n1132;
    wire n1136;
    wire n1140;
    wire n1144;
    wire n1148;
    wire n1152;
    wire n1156;
    wire n1159;
    wire n1163;
    wire n1166;
    wire n1170;
    wire n1174;
    wire n1178;
    wire n1182;
    wire n1186;
    wire n1190;
    wire n1194;
    wire n1198;
    wire n1202;
    wire n1205;
    wire n1208;
    wire n1212;
    wire n1216;
    wire n1220;
    wire n1224;
    wire n1228;
    wire n1232;
    wire n1236;
    wire n1240;
    wire n1244;
    wire n1248;
    wire n1252;
    wire n1256;
    wire n1259;
    wire n1263;
    wire n1266;
    wire n1270;
    wire n1274;
    wire n1278;
    wire n1282;
    wire n1285;
    wire n1289;
    wire n1293;
    wire n1297;
    wire n1301;
    wire n1304;
    wire n1308;
    wire n1311;
    wire n1315;
    wire n1319;
    wire n1323;
    wire n1326;
    wire n1330;
    wire n1333;
    wire n1337;
    wire n1341;
    wire n1345;
    wire n1349;
    wire n1353;
    wire n1356;
    wire n1360;
    wire n1363;
    wire n1367;
    wire n1371;
    wire n1375;
    wire n1379;
    wire n1383;
    wire n1387;
    wire n1391;
    wire n1395;
    wire n1399;
    wire n1402;
    wire n1406;
    wire n1410;
    wire n1414;
    wire n1418;
    wire n1421;
    wire n1425;
    wire n1429;
    wire n1433;
    wire n1437;
    wire n1441;
    wire n1444;
    wire n1448;
    wire n1452;
    wire n1456;
    wire n1460;
    wire n1463;
    wire n1467;
    wire n1471;
    wire n1474;
    wire n1478;
    wire n1481;
    wire n1485;
    wire n1489;
    wire n1493;
    wire n1497;
    wire n1501;
    wire n1505;
    wire n1509;
    wire n1513;
    wire n1517;
    wire n1521;
    wire n1525;
    wire n1529;
    wire n1533;
    wire n1536;
    wire n1540;
    wire n1544;
    wire n1548;
    wire n1552;
    wire n1556;
    wire n1560;
    wire n1563;
    wire n1567;
    wire n1571;
    wire n1575;
    wire n1579;
    wire n1583;
    wire n1587;
    wire n1591;
    wire n1595;
    wire n1599;
    wire n1602;
    wire n1606;
    wire n1610;
    wire n1613;
    wire n1617;
    wire n1621;
    wire n1625;
    wire n1629;
    wire n1633;
    wire n1637;
    wire n1640;
    wire n1644;
    wire n1648;
    wire n1652;
    wire n1656;
    wire n1660;
    wire n1664;
    wire n1668;
    wire n1672;
    wire n1676;
    wire n1680;
    wire n1684;
    wire n1688;
    wire n1692;
    wire n1696;
    wire n1699;
    wire n1703;
    wire n1707;
    wire n1711;
    wire n1715;
    wire n1719;
    wire n1723;
    wire n1727;
    wire n1731;
    wire n1735;
    wire n1738;
    wire n1742;
    wire n1745;
    wire n1749;
    wire n1752;
    wire n1756;
    wire n1760;
    wire n1763;
    wire n1767;
    wire n1771;
    wire n1774;
    wire n1778;
    wire n1782;
    wire n1786;
    wire n1790;
    wire n1794;
    wire n1798;
    wire n1802;
    wire n1806;
    wire n1810;
    wire n1814;
    wire n1818;
    wire n1822;
    wire n1826;
    wire n1830;
    wire n1834;
    wire n1838;
    wire n1842;
    wire n1846;
    wire n1850;
    wire n1854;
    wire n1858;
    wire n1862;
    wire n1866;
    wire n1870;
    wire n1874;
    wire n1878;
    wire n1882;
    wire n1886;
    wire n1890;
    wire n1894;
    wire n1898;
    wire n1901;
    wire n1905;
    wire n1909;
    wire n1913;
    wire n1916;
    wire n1920;
    wire n1924;
    wire n1928;
    wire n1932;
    wire n1936;
    wire n1940;
    wire n1944;
    wire n1948;
    wire n1952;
    wire n1956;
    wire n1960;
    wire n1963;
    wire n1966;
    wire n1970;
    wire n1974;
    wire n1978;
    wire n1981;
    wire n1985;
    wire n1988;
    wire n1992;
    wire n1996;
    wire n1999;
    wire n2003;
    wire n2007;
    wire n2010;
    wire n2013;
    wire n2017;
    wire n2020;
    wire n2024;
    wire n2028;
    wire n2032;
    wire n2036;
    wire n2040;
    wire n2044;
    wire n2047;
    wire n2051;
    wire n2054;
    wire n2058;
    wire n2062;
    wire n2065;
    wire n2069;
    wire n2073;
    wire n2077;
    wire n2081;
    wire n2085;
    wire n2089;
    wire n2093;
    wire n2097;
    wire n2101;
    wire n2104;
    wire n2108;
    wire n2111;
    wire n2115;
    wire n2119;
    wire n2123;
    wire n2127;
    wire n2131;
    wire n2135;
    wire n2139;
    wire n2143;
    wire n2147;
    wire n2150;
    wire n2153;
    wire n2157;
    wire n2160;
    wire n2164;
    wire n2168;
    wire n2172;
    wire n2175;
    wire n2178;
    wire n2181;
    wire n2185;
    wire n2188;
    wire n2191;
    wire n2195;
    wire n2199;
    wire n2203;
    wire n2207;
    wire n2211;
    wire n2215;
    wire n2219;
    wire n2223;
    wire n2227;
    wire n2230;
    wire n2233;
    wire n2236;
    wire n2240;
    wire n2244;
    wire n2248;
    wire n2252;
    wire n2256;
    wire n2260;
    wire n2264;
    wire n2268;
    wire n2271;
    wire n2274;
    wire n2278;
    wire n2282;
    wire n2286;
    wire n2290;
    wire n2294;
    wire n2298;
    wire n2302;
    wire n2306;
    wire n2310;
    wire n2314;
    wire n2317;
    wire n2321;
    wire n2325;
    wire n2329;
    wire n2333;
    wire n2337;
    wire n2341;
    wire n2345;
    wire n2349;
    wire n2352;
    wire n2356;
    wire n2360;
    wire n2364;
    wire n2368;
    wire n2372;
    wire n2376;
    wire n2380;
    wire n2384;
    wire n2387;
    wire n2391;
    wire n2394;
    wire n2398;
    wire n2402;
    wire n2406;
    wire n2410;
    wire n2414;
    wire n2418;
    wire n2422;
    wire n2426;
    wire n2430;
    wire n2433;
    wire n2436;
    wire n2439;
    wire n2443;
    wire n2447;
    wire n2451;
    wire n2455;
    wire n2459;
    wire n2463;
    wire n2467;
    wire n2471;
    wire n2475;
    wire n2479;
    wire n2483;
    wire n2486;
    wire n2490;
    wire n2494;
    wire n2498;
    wire n2502;
    wire n2506;
    wire n2510;
    wire n2514;
    wire n2518;
    wire n2521;
    wire n2525;
    wire n2529;
    wire n2533;
    wire n2537;
    wire n2541;
    wire n2545;
    wire n2549;
    wire n2553;
    wire n2557;
    wire n2560;
    wire n2563;
    wire n2567;
    wire n2571;
    wire n2575;
    wire n2579;
    wire n2583;
    wire n2587;
    wire n2591;
    wire n2595;
    wire n2598;
    wire n2601;
    wire n2605;
    wire n2609;
    wire n2613;
    wire n2617;
    wire n2621;
    wire n2625;
    wire n2629;
    wire n2633;
    wire n2637;
    wire n2641;
    wire n2645;
    wire n2649;
    wire n2653;
    wire n2656;
    wire n2660;
    wire n2664;
    wire n2668;
    wire n2672;
    wire n2676;
    wire n2680;
    wire n2684;
    wire n2688;
    wire n2692;
    wire n2696;
    wire n2700;
    wire n2704;
    wire n2708;
    wire n2711;
    wire n2714;
    wire n2717;
    wire n2721;
    wire n2725;
    wire n2728;
    wire n2732;
    wire n2736;
    wire n2740;
    wire n2743;
    wire n2746;
    wire n2750;
    wire n2754;
    wire n2758;
    wire n2762;
    wire n2765;
    wire n2768;
    wire n2772;
    wire n2775;
    wire n2779;
    wire n2783;
    wire n2787;
    wire n2790;
    wire n2794;
    wire n2798;
    wire n2802;
    wire n2805;
    wire n2809;
    wire n2812;
    wire n2816;
    wire n2820;
    wire n2824;
    wire n2828;
    wire n2832;
    wire n2835;
    wire n2839;
    wire n2843;
    wire n2847;
    wire n2851;
    wire n2855;
    wire n2858;
    wire n2862;
    wire n2866;
    wire n2870;
    wire n2873;
    wire n2877;
    wire n2881;
    wire n2884;
    wire n2888;
    wire n2892;
    wire n2896;
    wire n2899;
    wire n2902;
    wire n2906;
    wire n2910;
    wire n2914;
    wire n2918;
    wire n2921;
    wire n2925;
    wire n2929;
    wire n2933;
    wire n2937;
    wire n2941;
    wire n2944;
    wire n2948;
    wire n2952;
    wire n2956;
    wire n2960;
    wire n2964;
    wire n2968;
    wire n2972;
    wire n2975;
    wire n2978;
    wire n2982;
    wire n2986;
    wire n2990;
    wire n2994;
    wire n2998;
    wire n3002;
    wire n3006;
    wire n3010;
    wire n3014;
    wire n3018;
    wire n3021;
    wire n3025;
    wire n3028;
    wire n3032;
    wire n3036;
    wire n3040;
    wire n3044;
    wire n3048;
    wire n3052;
    wire n3056;
    wire n3060;
    wire n3063;
    wire n3067;
    wire n3070;
    wire n3074;
    wire n3078;
    wire n3082;
    wire n3086;
    wire n3090;
    wire n3094;
    wire n3098;
    wire n3102;
    wire n3105;
    wire n3109;
    wire n3112;
    wire n3116;
    wire n3120;
    wire n3124;
    wire n3128;
    wire n3132;
    wire n3136;
    wire n3140;
    wire n3144;
    wire n3147;
    wire n3151;
    wire n3154;
    wire n3158;
    wire n3162;
    wire n3166;
    wire n3170;
    wire n3174;
    wire n3178;
    wire n3182;
    wire n3186;
    wire n3190;
    wire n3194;
    wire n3198;
    wire n3202;
    wire n3206;
    wire n3210;
    wire n3214;
    wire n3218;
    wire n3222;
    wire n3226;
    wire n3230;
    wire n3234;
    wire n3238;
    wire n3242;
    wire n3246;
    wire n3250;
    wire n3254;
    wire n3258;
    wire n3262;
    wire n3266;
    wire n3270;
    wire n3274;
    wire n3278;
    wire n3282;
    wire n3286;
    wire n3290;
    wire n3294;
    wire n3298;
    wire n3302;
    wire n3306;
    wire n3310;
    wire n3314;
    wire n3318;
    wire n3322;
    wire n3326;
    wire n3330;
    wire n3334;
    wire n3338;
    wire n3342;
    wire n3346;
    wire n3350;
    wire n3354;
    wire n3358;
    wire n3362;
    wire n3366;
    wire n3370;
    wire n3374;
    wire n3378;
    wire n3382;
    wire n3386;
    wire n3390;
    wire n3394;
    wire n3398;
    wire n3402;
    wire n3406;
    wire n3410;
    wire n3414;
    wire n3418;
    wire n3422;
    wire n3426;
    wire n3430;
    wire n3434;
    wire n3438;
    wire n3442;
    wire n3446;
    wire n3450;
    wire n3454;
    wire n3458;
    wire n3462;
    wire n3466;
    wire n3470;
    wire n3474;
    wire n3478;
    wire n3482;
    wire n3486;
    wire n3490;
    wire n3494;
    wire n3498;
    wire n3502;
    wire n3506;
    wire n3510;
    wire n3514;
    wire n3518;
    wire n3522;
    wire n3526;
    wire n3530;
    wire n3534;
    wire n3538;
    wire n3542;
    wire n3546;
    wire n3550;
    wire n3554;
    wire n3558;
    wire n3562;
    wire n3566;
    wire n3570;
    wire n3574;
    wire n3578;
    wire n3582;
    wire n3586;
    wire n3590;
    wire n3594;
    wire n3598;
    wire n3602;
    wire n3606;
    wire n3610;
    wire n3614;
    wire n3618;
    wire n3621;
    wire n3624;
    wire n3628;
    wire n3631;
    wire n3635;
    wire n3638;
    wire n3641;
    wire n3645;
    wire n3648;
    wire n3652;
    wire n3656;
    wire n3660;
    wire n3664;
    wire n3668;
    wire n3672;
    wire n3676;
    wire n3680;
    wire n3684;
    wire n3688;
    wire n3692;
    wire n3696;
    wire n3700;
    wire n3704;
    wire n3707;
    wire n3711;
    wire n3715;
    wire n3718;
    wire n3722;
    wire n3726;
    wire n3729;
    wire n3732;
    wire n3736;
    wire n3740;
    wire n3744;
    wire n3748;
    wire n3751;
    wire n3755;
    wire n3759;
    wire n3763;
    wire n3767;
    wire n3770;
    wire n3774;
    wire n3778;
    wire n3781;
    wire n3785;
    wire n3788;
    wire n3792;
    wire n3796;
    wire n3800;
    wire n3804;
    wire n3808;
    wire n3812;
    wire n3816;
    wire n3819;
    wire n3823;
    wire n3827;
    wire n3831;
    wire n3835;
    wire n3839;
    wire n3843;
    wire n3847;
    wire n3850;
    wire n3854;
    wire n3858;
    wire n3862;
    wire n3866;
    wire n3869;
    wire n3873;
    wire n3876;
    wire n3880;
    wire n3884;
    wire n3888;
    wire n3892;
    wire n3896;
    wire n3900;
    wire n3904;
    wire n3907;
    wire n3911;
    wire n3915;
    wire n3919;
    wire n3923;
    wire n3926;
    wire n3930;
    wire n3933;
    wire n3937;
    wire n3941;
    wire n3945;
    wire n3949;
    wire n3953;
    wire n3957;
    wire n3961;
    wire n3965;
    wire n3969;
    wire n3973;
    wire n3977;
    wire n3981;
    wire n3985;
    wire n3989;
    wire n3993;
    wire n3997;
    wire n4001;
    wire n4005;
    wire n4009;
    wire n4013;
    wire n4017;
    wire n4021;
    wire n4025;
    wire n4029;
    wire n4032;
    wire n4036;
    wire n4040;
    wire n4044;
    wire n4048;
    wire n4052;
    wire n4056;
    wire n4060;
    wire n4064;
    wire n4068;
    wire n4072;
    wire n4076;
    wire n4080;
    wire n4084;
    wire n4088;
    wire n4092;
    wire n4096;
    wire n4100;
    wire n4103;
    wire n4107;
    wire n4110;
    wire n4114;
    wire n4118;
    wire n4122;
    wire n4126;
    wire n4130;
    wire n4134;
    wire n4138;
    wire n4142;
    wire n4146;
    wire n4150;
    wire n4154;
    wire n4158;
    wire n4162;
    wire n4166;
    wire n4170;
    wire n4174;
    wire n4178;
    wire n4182;
    wire n4186;
    wire n4190;
    wire n4194;
    wire n4198;
    wire n4202;
    wire n4206;
    wire n4210;
    wire n4214;
    wire n4218;
    wire n4222;
    wire n4226;
    wire n4230;
    wire n4234;
    wire n4238;
    wire n4242;
    wire n4246;
    wire n4250;
    wire n4254;
    wire n4258;
    wire n4262;
    wire n4266;
    wire n4270;
    wire n4274;
    wire n4278;
    wire n4282;
    wire n4286;
    wire n4290;
    wire n4294;
    wire n4298;
    wire n4302;
    wire n4306;
    wire n4310;
    wire n4314;
    wire n4318;
    wire n4322;
    wire n4326;
    wire n4330;
    wire n4334;
    wire n4338;
    wire n4342;
    wire n4346;
    wire n4350;
    wire n4354;
    wire n4358;
    wire n4362;
    wire n4366;
    wire n4370;
    wire n4374;
    wire n4378;
    wire n4382;
    wire n4386;
    wire n4390;
    wire n4394;
    wire n4398;
    wire n4402;
    wire n4406;
    wire n4410;
    wire n4414;
    wire n4418;
    wire n4422;
    wire n4426;
    wire n4430;
    wire n4434;
    wire n4438;
    wire n4442;
    wire n4446;
    wire n4450;
    wire n4454;
    wire n4458;
    wire n4462;
    wire n4466;
    wire n4470;
    wire n4474;
    wire n4478;
    wire n4482;
    wire n4486;
    wire n4490;
    wire n4494;
    wire n4498;
    wire n4502;
    wire n4506;
    wire n4510;
    wire n4514;
    wire n4518;
    wire n4522;
    wire n4526;
    wire n4530;
    wire n4534;
    wire n4538;
    wire n4542;
    wire n4546;
    wire n4550;
    wire n4554;
    wire n4558;
    wire n4561;
    wire n4564;
    wire n4567;
    wire n4571;
    wire n4575;
    wire n4579;
    wire n4583;
    wire n4586;
    wire n4590;
    wire n4594;
    wire n4598;
    wire n4602;
    wire n4606;
    wire n4610;
    wire n4613;
    wire n4616;
    wire n4620;
    wire n4624;
    wire n4627;
    wire n4630;
    wire n4634;
    wire n4638;
    wire n4642;
    wire n4646;
    wire n4650;
    wire n4654;
    wire n4658;
    wire n4662;
    wire n4666;
    wire n4670;
    wire n4674;
    wire n4678;
    wire n4682;
    wire n4686;
    wire n4690;
    wire n4694;
    wire n4698;
    wire n4702;
    wire n4706;
    wire n4710;
    wire n4713;
    wire n4717;
    wire n4721;
    wire n4725;
    wire n4729;
    wire n4733;
    wire n4737;
    wire n4741;
    wire n4745;
    wire n4749;
    wire n4753;
    wire n4757;
    wire n4761;
    wire n4765;
    wire n4769;
    wire n4773;
    wire n4777;
    wire n4781;
    wire n4785;
    wire n4789;
    wire n4793;
    wire n4797;
    wire n4801;
    wire n4805;
    wire n4809;
    wire n4813;
    wire n4817;
    wire n4821;
    wire n4825;
    wire n4829;
    wire n4833;
    wire n4837;
    wire n4841;
    wire n4845;
    wire n4849;
    wire n4853;
    wire n4857;
    wire n4861;
    wire n4865;
    wire n4869;
    wire n4873;
    wire n4877;
    wire n4881;
    wire n4885;
    wire n4889;
    wire n4893;
    wire n4897;
    wire n4901;
    wire n4905;
    wire n4908;
    wire n4912;
    wire n4916;
    wire n4919;
    wire n4923;
    wire n4927;
    wire n4931;
    wire n4935;
    wire n4939;
    wire n4943;
    wire n4947;
    wire n4951;
    wire n4955;
    wire n4959;
    wire n4963;
    wire n4967;
    wire n4971;
    wire n4975;
    wire n4979;
    wire n4983;
    wire n4987;
    wire n4991;
    wire n4995;
    wire n4999;
    wire n5003;
    wire n5007;
    wire n5011;
    wire n5015;
    wire n5019;
    wire n5023;
    wire n5027;
    wire n5031;
    wire n5035;
    wire n5039;
    wire n5043;
    wire n5047;
    wire n5051;
    wire n5055;
    wire n5059;
    wire n5063;
    wire n5067;
    wire n5071;
    wire n5075;
    wire n5079;
    wire n5083;
    wire n5087;
    wire n5091;
    wire n5095;
    wire n5099;
    wire n5103;
    wire n5107;
    wire n5111;
    wire n5115;
    wire n5119;
    wire n5123;
    wire n5127;
    wire n5131;
    wire n5135;
    wire n5139;
    wire n5143;
    wire n5147;
    wire n5151;
    wire n5155;
    wire n5159;
    wire n5163;
    wire n5167;
    wire n5171;
    wire n5175;
    wire n5179;
    wire n5183;
    wire n5187;
    wire n5191;
    wire n5195;
    wire n5199;
    wire n5203;
    wire n5207;
    wire n5211;
    wire n5215;
    wire n5219;
    wire n5223;
    wire n5227;
    wire n5231;
    wire n5235;
    wire n5239;
    wire n5243;
    wire n5247;
    wire n5251;
    wire n5254;
    wire n5258;
    wire n5262;
    wire n5265;
    wire n5269;
    wire n5273;
    wire n5276;
    wire n5280;
    wire n5284;
    wire n5288;
    wire n5292;
    wire n5296;
    wire n5299;
    wire n5302;
    wire n5305;
    wire n5309;
    wire n5313;
    wire n5317;
    wire n5321;
    wire n5325;
    wire n5329;
    wire n5333;
    wire n5337;
    wire n5341;
    wire n5345;
    wire n5349;
    wire n5353;
    wire n5357;
    wire n5360;
    wire n5364;
    wire n5367;
    wire n5371;
    wire n5375;
    wire n5379;
    wire n5383;
    wire n5387;
    wire n5391;
    wire n5395;
    wire n5399;
    wire n5403;
    wire n5407;
    wire n5411;
    wire n5415;
    wire n5419;
    wire n5422;
    wire n5426;
    wire n5430;
    wire n5434;
    wire n5438;
    wire n5442;
    wire n5446;
    wire n5450;
    wire n5454;
    wire n5458;
    wire n5462;
    wire n5466;
    wire n5470;
    wire n5473;
    wire n5477;
    wire n5481;
    wire n5485;
    wire n5489;
    wire n5493;
    wire n5497;
    wire n5501;
    wire n5505;
    wire n5509;
    wire n5512;
    wire n5516;
    wire n5520;
    wire n5524;
    wire n5528;
    wire n5532;
    wire n5536;
    wire n5540;
    wire n5544;
    wire n5548;
    wire n5552;
    wire n5556;
    wire n5560;
    wire n5564;
    wire n5568;
    wire n5572;
    wire n5576;
    wire n5580;
    wire n5583;
    wire n5587;
    wire n5590;
    wire n5594;
    wire n5598;
    wire n5601;
    wire n5605;
    wire n5608;
    wire n5612;
    wire n5616;
    wire n5620;
    wire n5624;
    wire n5628;
    wire n5632;
    wire n5636;
    wire n5640;
    wire n5644;
    wire n5648;
    wire n5652;
    wire n5656;
    wire n5660;
    wire n5663;
    wire n5666;
    wire n5669;
    wire n5673;
    wire n5676;
    wire n5679;
    wire n5683;
    wire n5687;
    wire n5691;
    wire n5695;
    wire n5699;
    wire n5703;
    wire n5707;
    wire n5714;
    wire n5718;
    wire n5721;
    wire n5725;
    wire n5729;
    wire n5733;
    wire n5737;
    wire n5741;
    wire n5745;
    wire n5749;
    wire n5756;
    wire n5759;
    wire n5762;
    wire n5765;
    wire n5768;
    wire n5771;
    wire n5774;
    wire n5777;
    wire n5780;
    wire n5783;
    wire n5786;
    wire n5789;
    wire n5792;
    wire n5795;
    wire n5798;
    wire n5801;
    wire n5805;
    wire n5809;
    wire n5813;
    wire n5817;
    wire n5821;
    wire n8401;
    wire n8404;
    wire n8407;
    wire n8410;
    wire n8413;
    wire n8416;
    wire n8419;
    wire n8422;
    wire n8425;
    wire n8428;
    wire n8431;
    wire n8434;
    wire n8436;
    wire n8439;
    wire n8442;
    wire n8445;
    wire n8448;
    wire n8451;
    wire n8454;
    wire n8457;
    wire n8461;
    wire n8464;
    wire n8467;
    wire n8470;
    wire n8473;
    wire n8476;
    wire n8478;
    wire n8481;
    wire n8484;
    wire n8487;
    wire n8490;
    wire n8493;
    wire n8496;
    wire n8499;
    wire n8502;
    wire n8505;
    wire n8509;
    wire n8512;
    wire n8515;
    wire n8518;
    wire n8521;
    wire n8524;
    wire n8527;
    wire n8530;
    wire n8533;
    wire n8536;
    wire n8539;
    wire n8542;
    wire n8545;
    wire n8548;
    wire n8551;
    wire n8554;
    wire n8556;
    wire n8559;
    wire n8563;
    wire n8566;
    wire n8569;
    wire n8572;
    wire n8575;
    wire n8577;
    wire n8580;
    wire n8583;
    wire n8586;
    wire n8589;
    wire n8593;
    wire n8596;
    wire n8599;
    wire n8602;
    wire n8605;
    wire n8608;
    wire n8611;
    wire n8614;
    wire n8617;
    wire n8620;
    wire n8623;
    wire n8625;
    wire n8628;
    wire n8631;
    wire n8634;
    wire n8637;
    wire n8640;
    wire n8643;
    wire n8646;
    wire n8649;
    wire n8652;
    wire n8656;
    wire n8659;
    wire n8662;
    wire n8665;
    wire n8668;
    wire n8671;
    wire n8674;
    wire n8677;
    wire n8680;
    wire n8683;
    wire n8686;
    wire n8689;
    wire n8691;
    wire n8694;
    wire n8697;
    wire n8700;
    wire n8703;
    wire n8706;
    wire n8709;
    wire n8712;
    wire n8715;
    wire n8718;
    wire n8722;
    wire n8725;
    wire n8728;
    wire n8731;
    wire n8734;
    wire n8737;
    wire n8740;
    wire n8743;
    wire n8746;
    wire n8749;
    wire n8752;
    wire n8755;
    wire n8758;
    wire n8761;
    wire n8764;
    wire n8767;
    wire n8770;
    wire n8773;
    wire n8776;
    wire n8779;
    wire n8782;
    wire n8785;
    wire n8788;
    wire n8791;
    wire n8794;
    wire n8797;
    wire n8800;
    wire n8803;
    wire n8806;
    wire n8809;
    wire n8812;
    wire n8815;
    wire n8818;
    wire n8821;
    wire n8824;
    wire n8827;
    wire n8830;
    wire n8833;
    wire n8836;
    wire n8839;
    wire n8842;
    wire n8845;
    wire n8848;
    wire n8851;
    wire n8854;
    wire n8857;
    wire n8860;
    wire n8863;
    wire n8866;
    wire n8869;
    wire n8872;
    wire n8875;
    wire n8878;
    wire n8881;
    wire n8884;
    wire n8887;
    wire n8890;
    wire n8893;
    wire n8896;
    wire n8899;
    wire n8901;
    wire n8904;
    wire n8908;
    wire n8911;
    wire n8914;
    wire n8917;
    wire n8920;
    wire n8922;
    wire n8925;
    wire n8928;
    wire n8931;
    wire n8934;
    wire n8937;
    wire n8940;
    wire n8943;
    wire n8946;
    wire n8949;
    wire n8952;
    wire n8956;
    wire n8959;
    wire n8962;
    wire n8965;
    wire n8968;
    wire n8971;
    wire n8974;
    wire n8977;
    wire n8980;
    wire n8983;
    wire n8986;
    wire n8989;
    wire n8992;
    wire n8995;
    wire n8998;
    wire n9001;
    wire n9004;
    wire n9007;
    wire n9010;
    wire n9012;
    wire n9015;
    wire n9018;
    wire n9021;
    wire n9024;
    wire n9027;
    wire n9030;
    wire n9034;
    wire n9037;
    wire n9040;
    wire n9043;
    wire n9046;
    wire n9049;
    wire n9052;
    wire n9055;
    wire n9058;
    wire n9061;
    wire n9064;
    wire n9067;
    wire n9070;
    wire n9073;
    wire n9076;
    wire n9079;
    wire n9082;
    wire n9084;
    wire n9087;
    wire n9090;
    wire n9093;
    wire n9096;
    wire n9099;
    wire n9102;
    wire n9105;
    wire n9108;
    wire n9111;
    wire n9114;
    wire n9117;
    wire n9120;
    wire n9123;
    wire n9126;
    wire n9129;
    wire n9132;
    wire n9135;
    wire n9138;
    wire n9141;
    wire n9144;
    wire n9147;
    wire n9150;
    wire n9153;
    wire n9156;
    wire n9159;
    wire n9162;
    wire n9165;
    wire n9168;
    wire n9171;
    wire n9174;
    wire n9177;
    wire n9180;
    wire n9183;
    wire n9186;
    wire n9189;
    wire n9192;
    wire n9195;
    wire n9198;
    wire n9201;
    wire n9204;
    wire n9207;
    wire n9210;
    wire n9213;
    wire n9216;
    wire n9219;
    wire n9222;
    wire n9225;
    wire n9228;
    wire n9231;
    wire n9234;
    wire n9237;
    wire n9240;
    wire n9243;
    wire n9246;
    wire n9249;
    wire n9252;
    wire n9255;
    wire n9258;
    wire n9262;
    wire n9265;
    wire n9268;
    wire n9271;
    wire n9274;
    wire n9277;
    wire n9280;
    wire n9283;
    wire n9286;
    wire n9289;
    wire n9292;
    wire n9295;
    wire n9298;
    wire n9301;
    wire n9303;
    wire n9306;
    wire n9309;
    wire n9312;
    wire n9315;
    wire n9318;
    wire n9321;
    wire n9324;
    wire n9327;
    wire n9330;
    wire n9333;
    wire n9336;
    wire n9339;
    wire n9342;
    wire n9345;
    wire n9348;
    wire n9351;
    wire n9354;
    wire n9357;
    wire n9360;
    wire n9363;
    wire n9366;
    wire n9369;
    wire n9372;
    wire n9375;
    wire n9379;
    wire n9382;
    wire n9385;
    wire n9388;
    wire n9391;
    wire n9394;
    wire n9397;
    wire n9400;
    wire n9403;
    wire n9406;
    wire n9409;
    wire n9412;
    wire n9415;
    wire n9418;
    wire n9421;
    wire n9424;
    wire n9427;
    wire n9429;
    wire n9432;
    wire n9435;
    wire n9439;
    wire n9442;
    wire n9445;
    wire n9448;
    wire n9451;
    wire n9454;
    wire n9457;
    wire n9460;
    wire n9463;
    wire n9466;
    wire n9469;
    wire n9472;
    wire n9475;
    wire n9478;
    wire n9481;
    wire n9483;
    wire n9486;
    wire n9489;
    wire n9492;
    wire n9495;
    wire n9498;
    wire n9501;
    wire n9504;
    wire n9508;
    wire n9511;
    wire n9514;
    wire n9517;
    wire n9520;
    wire n9523;
    wire n9526;
    wire n9529;
    wire n9532;
    wire n9535;
    wire n9538;
    wire n9541;
    wire n9544;
    wire n9547;
    wire n9550;
    wire n9553;
    wire n9556;
    wire n9559;
    wire n9562;
    wire n9565;
    wire n9567;
    wire n9570;
    wire n9573;
    wire n9576;
    wire n9579;
    wire n9582;
    wire n9585;
    wire n9588;
    wire n9591;
    wire n9594;
    wire n9597;
    wire n9600;
    wire n9603;
    wire n9606;
    wire n9609;
    wire n9613;
    wire n9615;
    wire n9618;
    wire n9621;
    wire n9624;
    wire n9627;
    wire n9630;
    wire n9633;
    wire n9636;
    wire n9639;
    wire n9642;
    wire n9645;
    wire n9648;
    wire n9651;
    wire n9654;
    wire n9657;
    wire n9660;
    wire n9664;
    wire n9667;
    wire n9670;
    wire n9673;
    wire n9676;
    wire n9679;
    wire n9682;
    wire n9685;
    wire n9688;
    wire n9691;
    wire n9694;
    wire n9697;
    wire n9700;
    wire n9703;
    wire n9705;
    wire n9708;
    wire n9711;
    wire n9714;
    wire n9717;
    wire n9720;
    wire n9723;
    wire n9726;
    wire n9729;
    wire n9732;
    wire n9735;
    wire n9738;
    wire n9741;
    wire n9744;
    wire n9747;
    wire n9750;
    wire n9753;
    wire n9756;
    wire n9759;
    wire n9762;
    wire n9765;
    wire n9768;
    wire n9771;
    wire n9774;
    wire n9777;
    wire n9781;
    wire n9783;
    wire n9786;
    wire n9789;
    wire n9792;
    wire n9795;
    wire n9798;
    wire n9801;
    wire n9804;
    wire n9807;
    wire n9810;
    wire n9813;
    wire n9816;
    wire n9819;
    wire n9822;
    wire n9825;
    wire n9828;
    wire n9831;
    wire n9834;
    wire n9837;
    wire n9840;
    wire n9843;
    wire n9846;
    wire n9849;
    wire n9852;
    wire n9855;
    wire n9858;
    wire n9861;
    wire n9864;
    wire n9868;
    wire n9871;
    wire n9874;
    wire n9877;
    wire n9880;
    wire n9883;
    wire n9886;
    wire n9889;
    wire n9892;
    wire n9895;
    wire n9898;
    wire n9901;
    wire n9904;
    wire n9907;
    wire n9909;
    wire n9912;
    wire n9916;
    wire n9919;
    wire n9922;
    wire n9925;
    wire n9927;
    wire n9930;
    wire n9934;
    wire n9937;
    wire n9940;
    wire n9943;
    wire n9946;
    wire n9949;
    wire n9952;
    wire n9955;
    wire n9958;
    wire n9961;
    wire n9964;
    wire n9967;
    wire n9970;
    wire n9973;
    wire n9976;
    wire n9979;
    wire n9982;
    wire n9985;
    wire n9988;
    wire n9991;
    wire n9994;
    wire n9997;
    wire n10000;
    wire n10003;
    wire n10006;
    wire n10009;
    wire n10012;
    wire n10015;
    wire n10018;
    wire n10021;
    wire n10024;
    wire n10026;
    wire n10029;
    wire n10032;
    wire n10035;
    wire n10038;
    wire n10041;
    wire n10044;
    wire n10047;
    wire n10050;
    wire n10053;
    wire n10056;
    wire n10059;
    wire n10062;
    wire n10065;
    wire n10068;
    wire n10071;
    wire n10074;
    wire n10077;
    wire n10080;
    wire n10083;
    wire n10086;
    wire n10089;
    wire n10093;
    wire n10096;
    wire n10099;
    wire n10102;
    wire n10105;
    wire n10108;
    wire n10111;
    wire n10114;
    wire n10117;
    wire n10120;
    wire n10123;
    wire n10126;
    wire n10129;
    wire n10132;
    wire n10134;
    wire n10137;
    wire n10140;
    wire n10144;
    wire n10147;
    wire n10150;
    wire n10153;
    wire n10156;
    wire n10159;
    wire n10162;
    wire n10165;
    wire n10168;
    wire n10171;
    wire n10174;
    wire n10177;
    wire n10180;
    wire n10183;
    wire n10185;
    wire n10188;
    wire n10191;
    wire n10195;
    wire n10198;
    wire n10201;
    wire n10204;
    wire n10207;
    wire n10210;
    wire n10213;
    wire n10216;
    wire n10219;
    wire n10222;
    wire n10225;
    wire n10228;
    wire n10231;
    wire n10234;
    wire n10237;
    wire n10240;
    wire n10243;
    wire n10246;
    wire n10249;
    wire n10252;
    wire n10255;
    wire n10258;
    wire n10261;
    wire n10264;
    wire n10267;
    wire n10270;
    wire n10273;
    wire n10276;
    wire n10279;
    wire n10282;
    wire n10285;
    wire n10288;
    wire n10291;
    wire n10294;
    wire n10297;
    wire n10300;
    wire n10303;
    wire n10306;
    wire n10309;
    wire n10312;
    wire n10315;
    wire n10318;
    wire n10321;
    wire n10324;
    wire n10327;
    wire n10330;
    wire n10333;
    wire n10336;
    wire n10339;
    wire n10342;
    wire n10345;
    wire n10348;
    wire n10351;
    wire n10354;
    wire n10357;
    wire n10360;
    wire n10363;
    wire n10366;
    wire n10369;
    wire n10372;
    wire n10375;
    wire n10378;
    wire n10381;
    wire n10384;
    wire n10387;
    wire n10390;
    wire n10393;
    wire n10396;
    wire n10399;
    wire n10402;
    wire n10405;
    wire n10408;
    wire n10411;
    wire n10414;
    wire n10417;
    wire n10420;
    wire n10423;
    wire n10426;
    wire n10429;
    wire n10432;
    wire n10435;
    wire n10438;
    wire n10441;
    wire n10444;
    wire n10447;
    wire n10450;
    wire n10453;
    wire n10456;
    wire n10459;
    wire n10462;
    wire n10465;
    wire n10468;
    wire n10471;
    wire n10474;
    wire n10477;
    wire n10480;
    wire n10483;
    wire n10486;
    wire n10489;
    wire n10492;
    wire n10495;
    wire n10498;
    wire n10501;
    wire n10504;
    wire n10507;
    wire n10510;
    wire n10513;
    wire n10516;
    wire n10519;
    wire n10521;
    wire n10524;
    wire n10528;
    wire n10531;
    wire n10534;
    wire n10536;
    wire n10539;
    wire n10542;
    wire n10545;
    wire n10548;
    wire n10551;
    wire n10554;
    wire n10558;
    wire n10561;
    wire n10564;
    wire n10567;
    wire n10570;
    wire n10573;
    wire n10576;
    wire n10579;
    wire n10582;
    wire n10585;
    wire n10588;
    wire n10591;
    wire n10594;
    wire n10597;
    wire n10600;
    wire n10603;
    wire n10606;
    wire n10609;
    wire n10611;
    wire n10614;
    wire n10617;
    wire n10620;
    wire n10623;
    wire n10626;
    wire n10629;
    wire n10632;
    wire n10635;
    wire n10638;
    wire n10641;
    wire n10644;
    wire n10647;
    wire n10651;
    wire n10654;
    wire n10656;
    wire n10659;
    wire n10662;
    wire n10665;
    wire n10668;
    wire n10671;
    wire n10674;
    wire n10677;
    wire n10680;
    wire n10684;
    wire n10687;
    wire n10690;
    wire n10693;
    wire n10696;
    wire n10699;
    wire n10702;
    wire n10705;
    wire n10708;
    wire n10711;
    wire n10714;
    wire n10717;
    wire n10720;
    wire n10723;
    wire n10726;
    wire n10729;
    wire n10732;
    wire n10735;
    wire n10738;
    wire n10741;
    wire n10744;
    wire n10747;
    wire n10750;
    wire n10753;
    wire n10756;
    wire n10759;
    wire n10762;
    wire n10765;
    wire n10768;
    wire n10771;
    wire n10774;
    wire n10777;
    wire n10780;
    wire n10783;
    wire n10786;
    wire n10789;
    wire n10792;
    wire n10795;
    wire n10798;
    wire n10801;
    wire n10804;
    wire n10807;
    wire n10809;
    wire n10812;
    wire n10815;
    wire n10818;
    wire n10821;
    wire n10825;
    wire n10828;
    wire n10831;
    wire n10834;
    wire n10837;
    wire n10840;
    wire n10843;
    wire n10846;
    wire n10849;
    wire n10852;
    wire n10855;
    wire n10858;
    wire n10861;
    wire n10864;
    wire n10867;
    wire n10870;
    wire n10873;
    wire n10876;
    wire n10879;
    wire n10882;
    wire n10885;
    wire n10888;
    wire n10891;
    wire n10894;
    wire n10897;
    wire n10900;
    wire n10903;
    wire n10906;
    wire n10909;
    wire n10912;
    wire n10915;
    wire n10918;
    wire n10921;
    wire n10924;
    wire n10927;
    wire n10929;
    wire n10932;
    wire n10935;
    wire n10938;
    wire n10941;
    wire n10944;
    wire n10947;
    wire n10950;
    wire n10953;
    wire n10956;
    wire n10959;
    wire n10963;
    wire n10966;
    wire n10968;
    wire n10971;
    wire n10974;
    wire n10978;
    wire n10981;
    wire n10984;
    wire n10987;
    wire n10990;
    wire n10993;
    wire n10996;
    wire n10999;
    wire n11002;
    wire n11005;
    wire n11008;
    wire n11011;
    wire n11014;
    wire n11017;
    wire n11020;
    wire n11023;
    wire n11025;
    wire n11028;
    wire n11031;
    wire n11034;
    wire n11037;
    wire n11040;
    wire n11043;
    wire n11046;
    wire n11049;
    wire n11052;
    wire n11055;
    wire n11058;
    wire n11061;
    wire n11064;
    wire n11067;
    wire n11070;
    wire n11073;
    wire n11076;
    wire n11079;
    wire n11082;
    wire n11086;
    wire n11089;
    wire n11091;
    wire n11094;
    wire n11097;
    wire n11100;
    wire n11103;
    wire n11106;
    wire n11109;
    wire n11113;
    wire n11116;
    wire n11119;
    wire n11122;
    wire n11125;
    wire n11128;
    wire n11131;
    wire n11134;
    wire n11137;
    wire n11140;
    wire n11143;
    wire n11146;
    wire n11149;
    wire n11152;
    wire n11155;
    wire n11158;
    wire n11161;
    wire n11164;
    wire n11167;
    wire n11170;
    wire n11173;
    wire n11176;
    wire n11179;
    wire n11182;
    wire n11185;
    wire n11188;
    wire n11191;
    wire n11194;
    wire n11197;
    wire n11200;
    wire n11203;
    wire n11206;
    wire n11209;
    wire n11212;
    wire n11215;
    wire n11218;
    wire n11221;
    wire n11224;
    wire n11227;
    wire n11230;
    wire n11233;
    wire n11236;
    wire n11239;
    wire n11242;
    wire n11245;
    wire n11248;
    wire n11251;
    wire n11254;
    wire n11257;
    wire n11260;
    wire n11263;
    wire n11266;
    wire n11269;
    wire n11272;
    wire n11275;
    wire n11277;
    wire n11280;
    wire n11283;
    wire n11286;
    wire n11289;
    wire n11292;
    wire n11295;
    wire n11298;
    wire n11301;
    wire n11304;
    wire n11307;
    wire n11311;
    wire n11314;
    wire n11317;
    wire n11320;
    wire n11323;
    wire n11325;
    wire n11328;
    wire n11331;
    wire n11334;
    wire n11337;
    wire n11340;
    wire n11343;
    wire n11346;
    wire n11349;
    wire n11352;
    wire n11355;
    wire n11358;
    wire n11361;
    wire n11364;
    wire n11367;
    wire n11370;
    wire n11373;
    wire n11377;
    wire n11380;
    wire n11383;
    wire n11386;
    wire n11389;
    wire n11392;
    wire n11395;
    wire n11398;
    wire n11401;
    wire n11404;
    wire n11406;
    wire n11409;
    wire n11413;
    wire n11416;
    wire n11419;
    wire n11422;
    wire n11425;
    wire n11428;
    wire n11431;
    wire n11434;
    wire n11437;
    wire n11440;
    wire n11443;
    wire n11446;
    wire n11449;
    wire n11452;
    wire n11455;
    wire n11457;
    wire n11460;
    wire n11463;
    wire n11466;
    wire n11470;
    wire n11473;
    wire n11476;
    wire n11479;
    wire n11482;
    wire n11485;
    wire n11488;
    wire n11491;
    wire n11494;
    wire n11497;
    wire n11500;
    wire n11503;
    wire n11506;
    wire n11509;
    wire n11512;
    wire n11515;
    wire n11518;
    wire n11521;
    wire n11524;
    wire n11527;
    wire n11530;
    wire n11533;
    wire n11536;
    wire n11539;
    wire n11542;
    wire n11545;
    wire n11547;
    wire n11550;
    wire n11553;
    wire n11556;
    wire n11559;
    wire n11562;
    wire n11565;
    wire n11568;
    wire n11571;
    wire n11574;
    wire n11577;
    wire n11580;
    wire n11583;
    wire n11586;
    wire n11589;
    wire n11592;
    wire n11595;
    wire n11598;
    wire n11601;
    wire n11604;
    wire n11607;
    wire n11610;
    wire n11613;
    wire n11616;
    wire n11619;
    wire n11623;
    wire n11626;
    wire n11629;
    wire n11632;
    wire n11635;
    wire n11638;
    wire n11641;
    wire n11644;
    wire n11647;
    wire n11650;
    wire n11653;
    wire n11656;
    wire n11659;
    wire n11662;
    wire n11665;
    wire n11668;
    wire n11671;
    wire n11674;
    wire n11677;
    wire n11680;
    wire n11683;
    wire n11686;
    wire n11689;
    wire n11692;
    wire n11694;
    wire n11697;
    wire n11700;
    wire n11703;
    wire n11706;
    wire n11709;
    wire n11712;
    wire n11715;
    wire n11718;
    wire n11721;
    wire n11724;
    wire n11727;
    wire n11730;
    wire n11733;
    wire n11736;
    wire n11739;
    wire n11742;
    wire n11745;
    wire n11748;
    wire n11751;
    wire n11754;
    wire n11757;
    wire n11760;
    wire n11763;
    wire n11766;
    wire n11769;
    wire n11772;
    wire n11775;
    wire n11778;
    wire n11781;
    wire n11784;
    wire n11787;
    wire n11790;
    wire n11793;
    wire n11796;
    wire n11799;
    wire n11802;
    wire n11805;
    wire n11808;
    wire n11811;
    wire n11814;
    wire n11817;
    wire n11820;
    wire n11823;
    wire n11826;
    wire n11829;
    wire n11832;
    wire n11835;
    wire n11838;
    wire n11841;
    wire n11844;
    wire n11847;
    wire n11850;
    wire n11853;
    wire n11856;
    wire n11859;
    wire n11862;
    wire n11865;
    wire n11868;
    wire n11871;
    wire n11874;
    wire n11877;
    wire n11880;
    wire n11883;
    wire n11886;
    wire n11890;
    wire n11893;
    wire n11896;
    wire n11899;
    wire n11902;
    wire n11905;
    wire n11908;
    wire n11911;
    wire n11914;
    wire n11917;
    wire n11920;
    wire n11923;
    wire n11926;
    wire n11929;
    wire n11932;
    wire n11935;
    wire n11938;
    wire n11941;
    wire n11944;
    wire n11947;
    wire n11950;
    wire n11953;
    wire n11955;
    wire n11958;
    wire n11961;
    wire n11964;
    wire n11967;
    wire n11970;
    wire n11973;
    wire n11976;
    wire n11979;
    wire n11982;
    wire n11985;
    wire n11988;
    wire n11991;
    wire n11994;
    wire n11997;
    wire n12000;
    wire n12003;
    wire n12006;
    wire n12009;
    wire n12012;
    wire n12015;
    wire n12018;
    wire n12021;
    wire n12024;
    wire n12027;
    wire n12030;
    wire n12033;
    wire n12036;
    wire n12039;
    wire n12042;
    wire n12045;
    wire n12048;
    wire n12051;
    wire n12054;
    wire n12057;
    wire n12060;
    wire n12063;
    wire n12066;
    wire n12070;
    wire n12073;
    wire n12076;
    wire n12079;
    wire n12082;
    wire n12085;
    wire n12088;
    wire n12091;
    wire n12094;
    wire n12097;
    wire n12100;
    wire n12103;
    wire n12106;
    wire n12109;
    wire n12112;
    wire n12115;
    wire n12118;
    wire n12121;
    wire n12124;
    wire n12127;
    wire n12130;
    wire n12132;
    wire n12136;
    wire n12139;
    wire n12142;
    wire n12145;
    wire n12148;
    wire n12151;
    wire n12154;
    wire n12157;
    wire n12160;
    wire n12163;
    wire n12166;
    wire n12169;
    wire n12172;
    wire n12175;
    wire n12178;
    wire n12181;
    wire n12184;
    wire n12187;
    wire n12190;
    wire n12193;
    wire n12196;
    wire n12199;
    wire n12201;
    wire n12204;
    wire n12207;
    wire n12210;
    wire n12213;
    wire n12216;
    wire n12219;
    wire n12222;
    wire n12225;
    wire n12228;
    wire n12231;
    wire n12234;
    wire n12237;
    wire n12240;
    wire n12243;
    wire n12246;
    wire n12249;
    wire n12252;
    wire n12255;
    wire n12258;
    wire n12261;
    wire n12264;
    wire n12267;
    wire n12270;
    wire n12273;
    wire n12276;
    wire n12279;
    wire n12282;
    wire n12285;
    wire n12288;
    wire n12291;
    wire n12294;
    wire n12297;
    wire n12300;
    wire n12303;
    wire n12306;
    wire n12309;
    wire n12312;
    wire n12315;
    wire n12318;
    wire n12321;
    wire n12324;
    wire n12327;
    wire n12330;
    wire n12333;
    wire n12336;
    wire n12339;
    wire n12342;
    wire n12345;
    wire n12348;
    wire n12351;
    wire n12354;
    wire n12357;
    wire n12360;
    wire n12363;
    wire n12366;
    wire n12369;
    wire n12372;
    wire n12375;
    wire n12378;
    wire n12381;
    wire n12384;
    wire n12387;
    wire n12390;
    wire n12393;
    wire n12396;
    wire n12399;
    wire n12402;
    wire n12405;
    wire n12408;
    wire n12411;
    wire n12414;
    wire n12417;
    wire n12420;
    wire n12424;
    wire n12427;
    wire n12430;
    wire n12433;
    wire n12436;
    wire n12439;
    wire n12442;
    wire n12445;
    wire n12448;
    wire n12451;
    wire n12454;
    wire n12457;
    wire n12460;
    wire n12463;
    wire n12466;
    wire n12469;
    wire n12472;
    wire n12475;
    wire n12478;
    wire n12481;
    wire n12484;
    wire n12487;
    wire n12490;
    wire n12492;
    wire n12495;
    wire n12498;
    wire n12501;
    wire n12504;
    wire n12507;
    wire n12510;
    wire n12513;
    wire n12516;
    wire n12519;
    wire n12522;
    wire n12525;
    wire n12528;
    wire n12531;
    wire n12534;
    wire n12537;
    wire n12540;
    wire n12543;
    wire n12546;
    wire n12549;
    wire n12552;
    wire n12555;
    wire n12558;
    wire n12561;
    wire n12564;
    wire n12567;
    wire n12570;
    wire n12573;
    wire n12576;
    wire n12579;
    wire n12582;
    wire n12585;
    wire n12588;
    wire n12591;
    wire n12594;
    wire n12597;
    wire n12600;
    wire n12603;
    wire n12606;
    wire n12609;
    wire n12612;
    wire n12615;
    wire n12618;
    wire n12621;
    wire n12624;
    wire n12627;
    wire n12630;
    wire n12633;
    wire n12636;
    wire n12639;
    wire n12642;
    wire n12645;
    wire n12648;
    wire n12651;
    wire n12654;
    wire n12657;
    wire n12660;
    wire n12663;
    wire n12666;
    wire n12669;
    wire n12672;
    wire n12675;
    wire n12678;
    wire n12681;
    wire n12684;
    wire n12687;
    wire n12690;
    wire n12693;
    wire n12696;
    wire n12699;
    wire n12702;
    wire n12705;
    wire n12708;
    wire n12711;
    wire n12714;
    wire n12717;
    wire n12720;
    wire n12723;
    wire n12727;
    wire n12730;
    wire n12733;
    wire n12736;
    wire n12739;
    wire n12742;
    wire n12745;
    wire n12748;
    wire n12751;
    wire n12754;
    wire n12757;
    wire n12760;
    wire n12763;
    wire n12766;
    wire n12769;
    wire n12772;
    wire n12775;
    wire n12778;
    wire n12781;
    wire n12784;
    wire n12786;
    wire n12790;
    wire n12793;
    wire n12796;
    wire n12799;
    wire n12802;
    wire n12805;
    wire n12808;
    wire n12811;
    wire n12814;
    wire n12817;
    wire n12820;
    wire n12823;
    wire n12826;
    wire n12829;
    wire n12832;
    wire n12835;
    wire n12838;
    wire n12841;
    wire n12844;
    wire n12847;
    wire n12850;
    wire n12853;
    wire n12856;
    wire n12859;
    wire n12862;
    wire n12864;
    wire n12867;
    wire n12870;
    wire n12873;
    wire n12876;
    wire n12879;
    wire n12882;
    wire n12885;
    wire n12888;
    wire n12891;
    wire n12894;
    wire n12897;
    wire n12900;
    wire n12903;
    wire n12906;
    wire n12909;
    wire n12912;
    wire n12915;
    wire n12918;
    wire n12921;
    wire n12924;
    wire n12927;
    wire n12930;
    wire n12933;
    wire n12936;
    wire n12939;
    wire n12942;
    wire n12945;
    wire n12948;
    wire n12951;
    wire n12954;
    wire n12957;
    wire n12960;
    wire n12963;
    wire n12966;
    wire n12969;
    wire n12972;
    wire n12975;
    wire n12978;
    wire n12981;
    wire n12984;
    wire n12987;
    wire n12990;
    wire n12993;
    wire n12996;
    wire n12999;
    wire n13002;
    wire n13005;
    wire n13008;
    wire n13011;
    wire n13014;
    wire n13017;
    wire n13020;
    wire n13023;
    wire n13026;
    wire n13029;
    wire n13032;
    wire n13035;
    wire n13038;
    wire n13041;
    wire n13044;
    wire n13047;
    wire n13050;
    wire n13053;
    wire n13056;
    wire n13059;
    wire n13062;
    wire n13065;
    wire n13068;
    wire n13071;
    wire n13074;
    wire n13077;
    wire n13080;
    wire n13083;
    wire n13087;
    wire n13090;
    wire n13093;
    wire n13096;
    wire n13099;
    wire n13102;
    wire n13105;
    wire n13108;
    wire n13111;
    wire n13114;
    wire n13117;
    wire n13120;
    wire n13123;
    wire n13126;
    wire n13129;
    wire n13132;
    wire n13135;
    wire n13138;
    wire n13141;
    wire n13144;
    wire n13147;
    wire n13150;
    wire n13152;
    wire n13155;
    wire n13158;
    wire n13161;
    wire n13164;
    wire n13167;
    wire n13170;
    wire n13173;
    wire n13176;
    wire n13179;
    wire n13182;
    wire n13185;
    wire n13188;
    wire n13191;
    wire n13194;
    wire n13197;
    wire n13200;
    wire n13203;
    wire n13206;
    wire n13209;
    wire n13213;
    wire n13216;
    wire n13219;
    wire n13222;
    wire n13225;
    wire n13228;
    wire n13231;
    wire n13234;
    wire n13237;
    wire n13240;
    wire n13243;
    wire n13246;
    wire n13249;
    wire n13252;
    wire n13255;
    wire n13258;
    wire n13261;
    wire n13264;
    wire n13267;
    wire n13270;
    wire n13273;
    wire n13276;
    wire n13279;
    wire n13282;
    wire n13285;
    wire n13288;
    wire n13291;
    wire n13294;
    wire n13297;
    wire n13300;
    wire n13303;
    wire n13306;
    wire n13309;
    wire n13312;
    wire n13315;
    wire n13318;
    wire n13321;
    wire n13324;
    wire n13327;
    wire n13330;
    wire n13333;
    wire n13335;
    wire n13338;
    wire n13342;
    wire n13345;
    wire n13348;
    wire n13351;
    wire n13354;
    wire n13357;
    wire n13360;
    wire n13363;
    wire n13366;
    wire n13369;
    wire n13372;
    wire n13375;
    wire n13378;
    wire n13381;
    wire n13384;
    wire n13387;
    wire n13390;
    wire n13393;
    wire n13396;
    wire n13399;
    wire n13402;
    wire n13405;
    wire n13407;
    wire n13410;
    wire n13413;
    wire n13416;
    wire n13419;
    wire n13422;
    wire n13425;
    wire n13428;
    wire n13431;
    wire n13434;
    wire n13437;
    wire n13440;
    wire n13443;
    wire n13446;
    wire n13449;
    wire n13452;
    wire n13455;
    wire n13458;
    wire n13461;
    wire n13464;
    wire n13468;
    wire n13471;
    wire n13474;
    wire n13477;
    wire n13480;
    wire n13483;
    wire n13486;
    wire n13489;
    wire n13492;
    wire n13495;
    wire n13497;
    wire n13501;
    wire n13504;
    wire n13507;
    wire n13510;
    wire n13513;
    wire n13516;
    wire n13519;
    wire n13522;
    wire n13525;
    wire n13528;
    wire n13531;
    wire n13534;
    wire n13537;
    wire n13540;
    wire n13543;
    wire n13546;
    wire n13549;
    wire n13552;
    wire n13555;
    wire n13558;
    wire n13561;
    wire n13564;
    wire n13567;
    wire n13570;
    wire n13573;
    wire n13576;
    wire n13579;
    wire n13582;
    wire n13585;
    wire n13588;
    wire n13591;
    wire n13594;
    wire n13597;
    wire n13600;
    wire n13603;
    wire n13606;
    wire n13609;
    wire n13612;
    wire n13615;
    wire n13618;
    wire n13621;
    wire n13624;
    wire n13627;
    wire n13630;
    wire n13633;
    wire n13636;
    wire n13639;
    wire n13642;
    wire n13645;
    wire n13648;
    wire n13651;
    wire n13653;
    wire n13656;
    wire n13659;
    wire n13662;
    wire n13665;
    wire n13668;
    wire n13671;
    wire n13675;
    wire n13678;
    wire n13681;
    wire n13684;
    wire n13687;
    wire n13690;
    wire n13693;
    wire n13696;
    wire n13699;
    wire n13702;
    wire n13705;
    wire n13708;
    wire n13711;
    wire n13714;
    wire n13717;
    wire n13720;
    wire n13723;
    wire n13726;
    wire n13728;
    wire n13731;
    wire n13734;
    wire n13737;
    wire n13740;
    wire n13744;
    wire n13747;
    wire n13750;
    wire n13753;
    wire n13756;
    wire n13759;
    wire n13762;
    wire n13765;
    wire n13767;
    wire n13770;
    wire n13773;
    wire n13776;
    wire n13779;
    wire n13782;
    wire n13786;
    wire n13789;
    wire n13792;
    wire n13795;
    wire n13798;
    wire n13801;
    wire n13804;
    wire n13807;
    wire n13810;
    wire n13813;
    wire n13816;
    wire n13819;
    wire n13822;
    wire n13825;
    wire n13828;
    wire n13831;
    wire n13834;
    wire n13837;
    wire n13840;
    wire n13843;
    wire n13846;
    wire n13849;
    wire n13852;
    wire n13855;
    wire n13858;
    wire n13861;
    wire n13864;
    wire n13867;
    wire n13870;
    wire n13873;
    wire n13876;
    wire n13879;
    wire n13882;
    wire n13885;
    wire n13888;
    wire n13891;
    wire n13894;
    wire n13897;
    wire n13900;
    wire n13903;
    wire n13906;
    wire n13909;
    wire n13912;
    wire n13915;
    wire n13918;
    wire n13921;
    wire n13924;
    wire n13927;
    wire n13930;
    wire n13933;
    wire n13936;
    wire n13939;
    wire n13942;
    wire n13945;
    wire n13948;
    wire n13951;
    wire n13954;
    wire n13957;
    wire n13960;
    wire n13963;
    wire n13966;
    wire n13969;
    wire n13972;
    wire n13975;
    wire n13978;
    wire n13981;
    wire n13984;
    wire n13987;
    wire n13990;
    wire n13993;
    wire n13996;
    wire n13999;
    wire n14002;
    wire n14005;
    wire n14008;
    wire n14011;
    wire n14014;
    wire n14017;
    wire n14020;
    wire n14023;
    wire n14026;
    wire n14029;
    wire n14032;
    wire n14035;
    wire n14038;
    wire n14041;
    wire n14044;
    wire n14047;
    wire n14050;
    wire n14053;
    wire n14056;
    wire n14059;
    wire n14062;
    wire n14065;
    wire n14068;
    wire n14071;
    wire n14074;
    wire n14077;
    wire n14080;
    wire n14083;
    wire n14086;
    wire n14089;
    wire n14092;
    wire n14095;
    wire n14098;
    wire n14101;
    wire n14104;
    wire n14107;
    wire n14110;
    wire n14113;
    wire n14116;
    wire n14119;
    wire n14122;
    wire n14125;
    wire n14128;
    wire n14131;
    wire n14134;
    wire n14137;
    wire n14140;
    wire n14143;
    wire n14146;
    wire n14149;
    wire n14152;
    wire n14155;
    wire n14158;
    wire n14161;
    wire n14164;
    wire n14167;
    wire n14170;
    wire n14173;
    wire n14176;
    wire n14179;
    wire n14182;
    wire n14185;
    wire n14188;
    wire n14191;
    wire n14194;
    wire n14197;
    wire n14200;
    wire n14203;
    wire n14206;
    wire n14209;
    wire n14212;
    wire n14215;
    wire n14218;
    wire n14221;
    wire n14224;
    wire n14227;
    wire n14230;
    wire n14233;
    wire n14236;
    wire n14239;
    wire n14242;
    wire n14245;
    wire n14248;
    wire n14250;
    wire n14253;
    wire n14256;
    wire n14260;
    wire n14263;
    wire n14266;
    wire n14268;
    wire n14271;
    wire n14274;
    wire n14277;
    wire n14280;
    wire n14283;
    wire n14286;
    wire n14289;
    wire n14292;
    wire n14295;
    wire n14298;
    wire n14301;
    wire n14304;
    wire n14308;
    wire n14311;
    wire n14314;
    wire n14317;
    wire n14320;
    wire n14323;
    wire n14325;
    wire n14328;
    wire n14331;
    wire n14334;
    wire n14337;
    wire n14341;
    wire n14344;
    wire n14346;
    wire n14349;
    wire n14353;
    wire n14356;
    wire n14359;
    wire n14362;
    wire n14365;
    wire n14368;
    wire n14371;
    wire n14374;
    wire n14377;
    wire n14380;
    wire n14383;
    wire n14386;
    wire n14389;
    wire n14392;
    wire n14395;
    wire n14398;
    wire n14401;
    wire n14404;
    wire n14407;
    wire n14410;
    wire n14413;
    wire n14416;
    wire n14419;
    wire n14422;
    wire n14425;
    wire n14428;
    wire n14430;
    wire n14433;
    wire n14436;
    wire n14439;
    wire n14442;
    wire n14445;
    wire n14448;
    wire n14451;
    wire n14454;
    wire n14457;
    wire n14460;
    wire n14463;
    wire n14466;
    wire n14469;
    wire n14472;
    wire n14475;
    wire n14478;
    wire n14481;
    wire n14484;
    wire n14487;
    wire n14490;
    wire n14493;
    wire n14496;
    wire n14499;
    wire n14502;
    wire n14505;
    wire n14508;
    wire n14511;
    wire n14514;
    wire n14517;
    wire n14520;
    wire n14524;
    wire n14527;
    wire n14529;
    wire n14532;
    wire n14535;
    wire n14538;
    wire n14541;
    wire n14544;
    wire n14547;
    wire n14550;
    wire n14553;
    wire n14556;
    wire n14559;
    wire n14562;
    wire n14565;
    wire n14568;
    wire n14571;
    wire n14575;
    wire n14578;
    wire n14581;
    wire n14584;
    wire n14587;
    wire n14590;
    wire n14593;
    wire n14596;
    wire n14599;
    wire n14602;
    wire n14605;
    wire n14608;
    wire n14611;
    wire n14614;
    wire n14617;
    wire n14620;
    wire n14623;
    wire n14626;
    wire n14629;
    wire n14632;
    wire n14635;
    wire n14638;
    wire n14641;
    wire n14644;
    wire n14647;
    wire n14650;
    wire n14653;
    wire n14656;
    wire n14659;
    wire n14662;
    wire n14665;
    wire n14668;
    wire n14671;
    wire n14674;
    wire n14677;
    wire n14680;
    wire n14683;
    wire n14686;
    wire n14689;
    wire n14692;
    wire n14695;
    wire n14698;
    wire n14701;
    wire n14704;
    wire n14707;
    wire n14710;
    wire n14713;
    wire n14716;
    wire n14719;
    wire n14722;
    wire n14725;
    wire n14727;
    wire n14730;
    wire n14733;
    wire n14736;
    wire n14740;
    wire n14743;
    wire n14745;
    wire n14748;
    wire n14751;
    wire n14754;
    wire n14757;
    wire n14760;
    wire n14763;
    wire n14766;
    wire n14769;
    wire n14772;
    wire n14775;
    wire n14778;
    wire n14781;
    wire n14784;
    wire n14787;
    wire n14790;
    wire n14793;
    wire n14796;
    wire n14799;
    wire n14802;
    wire n14805;
    wire n14808;
    wire n14811;
    wire n14814;
    wire n14817;
    wire n14820;
    wire n14823;
    wire n14826;
    wire n14829;
    wire n14832;
    wire n14835;
    wire n14838;
    wire n14841;
    wire n14844;
    wire n14847;
    wire n14850;
    wire n14853;
    wire n14856;
    wire n14859;
    wire n14862;
    wire n14865;
    wire n14868;
    wire n14871;
    wire n14874;
    wire n14878;
    wire n14881;
    wire n14884;
    wire n14887;
    wire n14890;
    wire n14893;
    wire n14896;
    wire n14899;
    wire n14902;
    wire n14905;
    wire n14908;
    wire n14911;
    wire n14914;
    wire n14917;
    wire n14920;
    wire n14923;
    wire n14926;
    wire n14929;
    wire n14932;
    wire n14935;
    wire n14938;
    wire n14941;
    wire n14944;
    wire n14947;
    wire n14950;
    wire n14953;
    wire n14956;
    wire n14959;
    wire n14962;
    wire n14965;
    wire n14968;
    wire n14971;
    wire n14974;
    wire n14977;
    wire n14980;
    wire n14983;
    wire n14986;
    wire n14989;
    wire n14992;
    wire n14995;
    wire n14998;
    wire n15001;
    wire n15004;
    wire n15007;
    wire n15010;
    wire n15013;
    wire n15016;
    wire n15019;
    wire n15022;
    wire n15025;
    wire n15028;
    wire n15031;
    wire n15034;
    wire n15037;
    wire n15039;
    wire n15043;
    wire n15046;
    wire n15049;
    wire n15052;
    wire n15055;
    wire n15057;
    wire n15060;
    wire n15063;
    wire n15067;
    wire n15070;
    wire n15073;
    wire n15076;
    wire n15079;
    wire n15082;
    wire n15085;
    wire n15088;
    wire n15091;
    wire n15094;
    wire n15097;
    wire n15100;
    wire n15103;
    wire n15106;
    wire n15109;
    wire n15111;
    wire n15114;
    wire n15117;
    wire n15120;
    wire n15123;
    wire n15126;
    wire n15129;
    wire n15132;
    wire n15135;
    wire n15138;
    wire n15141;
    wire n15144;
    wire n15147;
    wire n15150;
    wire n15153;
    wire n15156;
    wire n15159;
    wire n15162;
    wire n15165;
    wire n15168;
    wire n15171;
    wire n15174;
    wire n15177;
    wire n15180;
    wire n15183;
    wire n15186;
    wire n15189;
    wire n15192;
    wire n15196;
    wire n15199;
    wire n15202;
    wire n15205;
    wire n15208;
    wire n15211;
    wire n15214;
    wire n15217;
    wire n15220;
    wire n15223;
    wire n15226;
    wire n15229;
    wire n15232;
    wire n15235;
    wire n15238;
    wire n15241;
    wire n15244;
    wire n15247;
    wire n15250;
    wire n15253;
    wire n15256;
    wire n15259;
    wire n15262;
    wire n15265;
    wire n15268;
    wire n15271;
    wire n15274;
    wire n15277;
    wire n15280;
    wire n15283;
    wire n15286;
    wire n15289;
    wire n15292;
    wire n15295;
    wire n15298;
    wire n15301;
    wire n15304;
    wire n15307;
    wire n15310;
    wire n15313;
    wire n15316;
    wire n15319;
    wire n15321;
    wire n15324;
    wire n15327;
    wire n15330;
    wire n15333;
    wire n15336;
    wire n15339;
    wire n15342;
    wire n15345;
    wire n15348;
    wire n15351;
    wire n15354;
    wire n15357;
    wire n15360;
    wire n15363;
    wire n15366;
    wire n15369;
    wire n15372;
    wire n15375;
    wire n15378;
    wire n15381;
    wire n15385;
    wire n15388;
    wire n15391;
    wire n15394;
    wire n15397;
    wire n15400;
    wire n15403;
    wire n15406;
    wire n15409;
    wire n15412;
    wire n15415;
    wire n15418;
    wire n15421;
    wire n15424;
    wire n15427;
    wire n15430;
    wire n15433;
    wire n15436;
    wire n15439;
    wire n15442;
    wire n15445;
    wire n15448;
    wire n15451;
    wire n15453;
    wire n15456;
    wire n15459;
    wire n15462;
    wire n15465;
    wire n15468;
    wire n15471;
    wire n15474;
    wire n15477;
    wire n15480;
    wire n15483;
    wire n15486;
    wire n15489;
    wire n15492;
    wire n15495;
    wire n15498;
    wire n15501;
    wire n15504;
    wire n15507;
    wire n15510;
    wire n15513;
    wire n15516;
    wire n15519;
    wire n15522;
    wire n15525;
    wire n15528;
    wire n15531;
    wire n15534;
    wire n15537;
    wire n15540;
    wire n15543;
    wire n15546;
    wire n15549;
    wire n15552;
    wire n15555;
    wire n15558;
    wire n15561;
    wire n15564;
    wire n15567;
    wire n15571;
    wire n15574;
    wire n15577;
    wire n15580;
    wire n15583;
    wire n15586;
    wire n15589;
    wire n15592;
    wire n15595;
    wire n15597;
    wire n15600;
    wire n15604;
    wire n15607;
    wire n15609;
    wire n15612;
    wire n15615;
    wire n15618;
    wire n15621;
    wire n15624;
    wire n15627;
    wire n15630;
    wire n15633;
    wire n15636;
    wire n15639;
    wire n15642;
    wire n15645;
    wire n15648;
    wire n15651;
    wire n15654;
    wire n15657;
    wire n15660;
    wire n15663;
    wire n15666;
    wire n15669;
    wire n15672;
    wire n15675;
    wire n15678;
    wire n15681;
    wire n15684;
    wire n15687;
    wire n15690;
    wire n15693;
    wire n15696;
    wire n15699;
    wire n15702;
    wire n15705;
    wire n15708;
    wire n15711;
    wire n15714;
    wire n15717;
    wire n15720;
    wire n15723;
    wire n15726;
    wire n15729;
    wire n15732;
    wire n15735;
    wire n15738;
    wire n15741;
    wire n15744;
    wire n15747;
    wire n15750;
    wire n15753;
    wire n15756;
    wire n15759;
    wire n15762;
    wire n15765;
    wire n15768;
    wire n15771;
    wire n15774;
    wire n15777;
    wire n15780;
    wire n15783;
    wire n15787;
    wire n15790;
    wire n15793;
    wire n15796;
    wire n15799;
    wire n15802;
    wire n15805;
    wire n15808;
    wire n15811;
    wire n15814;
    wire n15817;
    wire n15820;
    wire n15823;
    wire n15826;
    wire n15829;
    wire n15832;
    wire n15835;
    wire n15838;
    wire n15841;
    wire n15844;
    wire n15847;
    wire n15850;
    wire n15853;
    wire n15855;
    wire n15858;
    wire n15861;
    wire n15864;
    wire n15867;
    wire n15870;
    wire n15873;
    wire n15876;
    wire n15879;
    wire n15882;
    wire n15885;
    wire n15888;
    wire n15891;
    wire n15894;
    wire n15897;
    wire n15900;
    wire n15903;
    wire n15906;
    wire n15909;
    wire n15912;
    wire n15915;
    wire n15918;
    wire n15921;
    wire n15924;
    wire n15927;
    wire n15930;
    wire n15933;
    wire n15936;
    wire n15939;
    wire n15942;
    wire n15945;
    wire n15948;
    wire n15951;
    wire n15954;
    wire n15957;
    wire n15960;
    wire n15963;
    wire n15966;
    wire n15969;
    wire n15972;
    wire n15976;
    wire n15979;
    wire n15982;
    wire n15985;
    wire n15988;
    wire n15991;
    wire n15994;
    wire n15997;
    wire n16000;
    wire n16002;
    wire n16005;
    wire n16008;
    wire n16012;
    wire n16015;
    wire n16017;
    wire n16020;
    wire n16023;
    wire n16026;
    wire n16029;
    wire n16032;
    wire n16035;
    wire n16038;
    wire n16041;
    wire n16044;
    wire n16047;
    wire n16050;
    wire n16053;
    wire n16056;
    wire n16059;
    wire n16062;
    wire n16065;
    wire n16068;
    wire n16071;
    wire n16074;
    wire n16077;
    wire n16080;
    wire n16083;
    wire n16086;
    wire n16089;
    wire n16092;
    wire n16095;
    wire n16098;
    wire n16101;
    wire n16104;
    wire n16107;
    wire n16111;
    wire n16113;
    wire n16116;
    wire n16119;
    wire n16122;
    wire n16125;
    wire n16128;
    wire n16131;
    wire n16134;
    wire n16137;
    wire n16140;
    wire n16143;
    wire n16146;
    wire n16149;
    wire n16152;
    wire n16155;
    wire n16158;
    wire n16161;
    wire n16164;
    wire n16167;
    wire n16170;
    wire n16173;
    wire n16176;
    wire n16179;
    wire n16182;
    wire n16185;
    wire n16188;
    wire n16191;
    wire n16194;
    wire n16198;
    wire n16201;
    wire n16204;
    wire n16207;
    wire n16210;
    wire n16213;
    wire n16216;
    wire n16219;
    wire n16222;
    wire n16225;
    wire n16228;
    wire n16231;
    wire n16234;
    wire n16237;
    wire n16240;
    wire n16243;
    wire n16246;
    wire n16249;
    wire n16252;
    wire n16255;
    wire n16258;
    wire n16261;
    wire n16264;
    wire n16267;
    wire n16270;
    wire n16273;
    wire n16276;
    wire n16279;
    wire n16282;
    wire n16285;
    wire n16288;
    wire n16291;
    wire n16294;
    wire n16297;
    wire n16300;
    wire n16303;
    wire n16306;
    wire n16309;
    wire n16312;
    wire n16315;
    wire n16318;
    wire n16321;
    wire n16324;
    wire n16327;
    wire n16330;
    wire n16332;
    wire n16335;
    wire n16338;
    wire n16341;
    wire n16344;
    wire n16347;
    wire n16350;
    wire n16353;
    wire n16356;
    wire n16359;
    wire n16362;
    wire n16365;
    wire n16368;
    wire n16371;
    wire n16374;
    wire n16377;
    wire n16380;
    wire n16383;
    wire n16386;
    wire n16389;
    wire n16392;
    wire n16395;
    wire n16398;
    wire n16401;
    wire n16404;
    wire n16407;
    wire n16410;
    wire n16413;
    wire n16416;
    wire n16419;
    wire n16422;
    wire n16425;
    wire n16428;
    wire n16431;
    wire n16434;
    wire n16437;
    wire n16440;
    wire n16443;
    wire n16446;
    wire n16449;
    wire n16452;
    wire n16455;
    wire n16458;
    wire n16461;
    wire n16464;
    wire n16467;
    wire n16470;
    wire n16473;
    wire n16476;
    wire n16479;
    wire n16482;
    wire n16485;
    wire n16488;
    wire n16491;
    wire n16494;
    wire n16497;
    wire n16500;
    wire n16503;
    wire n16506;
    wire n16509;
    wire n16512;
    wire n16515;
    wire n16518;
    wire n16521;
    wire n16524;
    wire n16527;
    wire n16530;
    wire n16533;
    wire n16536;
    wire n16539;
    wire n16542;
    wire n16545;
    wire n16548;
    wire n16551;
    wire n16554;
    wire n16557;
    wire n16560;
    wire n16563;
    wire n16566;
    wire n16569;
    wire n16572;
    wire n16575;
    wire n16578;
    wire n16581;
    wire n16584;
    wire n16587;
    wire n16590;
    wire n16593;
    wire n16596;
    wire n16599;
    wire n16602;
    wire n16605;
    wire n16608;
    wire n16611;
    wire n16614;
    wire n16617;
    wire n16620;
    wire n16623;
    wire n16626;
    wire n16629;
    wire n16632;
    wire n16635;
    wire n16638;
    wire n16641;
    wire n16644;
    wire n16647;
    wire n16650;
    wire n16653;
    wire n16656;
    wire n16659;
    wire n16662;
    wire n16665;
    wire n16668;
    wire n16671;
    wire n16674;
    wire n16677;
    wire n16680;
    wire n16683;
    wire n16686;
    wire n16689;
    wire n16692;
    wire n16695;
    wire n16698;
    wire n16701;
    wire n16704;
    wire n16707;
    wire n16710;
    wire n16713;
    wire n16716;
    wire n16719;
    wire n16722;
    wire n16725;
    wire n16728;
    wire n16731;
    wire n16734;
    wire n16737;
    wire n16740;
    wire n16743;
    wire n16746;
    wire n16749;
    wire n16752;
    wire n16755;
    wire n16758;
    wire n16761;
    wire n16764;
    wire n16767;
    wire n16770;
    wire n16773;
    wire n16776;
    wire n16779;
    wire n16782;
    wire n16785;
    wire n16788;
    wire n16791;
    wire n16794;
    wire n16797;
    wire n16800;
    wire n16803;
    wire n16806;
    wire n16809;
    wire n16812;
    wire n16815;
    wire n16818;
    wire n16821;
    wire n16824;
    wire n16827;
    wire n16830;
    wire n16833;
    wire n16836;
    wire n16839;
    wire n16842;
    wire n16845;
    wire n16848;
    wire n16851;
    wire n16854;
    wire n16857;
    wire n16860;
    wire n16863;
    wire n16866;
    wire n16869;
    wire n16872;
    wire n16875;
    wire n16879;
    wire n16882;
    wire n16885;
    wire n16888;
    wire n16891;
    wire n16894;
    wire n16897;
    wire n16900;
    wire n16903;
    wire n16906;
    wire n16909;
    wire n16912;
    wire n16915;
    wire n16918;
    wire n16921;
    wire n16924;
    wire n16927;
    wire n16930;
    wire n16933;
    wire n16936;
    wire n16939;
    wire n16942;
    wire n16945;
    wire n16948;
    wire n16951;
    wire n16954;
    wire n16957;
    wire n16960;
    wire n16963;
    wire n16966;
    wire n16969;
    wire n16972;
    wire n16975;
    wire n16978;
    wire n16981;
    wire n16984;
    wire n16987;
    wire n16990;
    wire n16993;
    wire n16996;
    wire n16999;
    wire n17002;
    wire n17005;
    wire n17008;
    wire n17011;
    wire n17014;
    wire n17017;
    wire n17020;
    wire n17023;
    wire n17026;
    wire n17029;
    wire n17032;
    wire n17035;
    wire n17038;
    wire n17041;
    wire n17044;
    wire n17047;
    wire n17050;
    wire n17053;
    wire n17056;
    wire n17059;
    wire n17062;
    wire n17065;
    wire n17068;
    wire n17071;
    wire n17074;
    wire n17077;
    wire n17080;
    wire n17083;
    wire n17086;
    wire n17089;
    wire n17092;
    wire n17095;
    wire n17098;
    wire n17101;
    wire n17104;
    wire n17106;
    wire n17110;
    wire n17113;
    wire n17115;
    wire n17119;
    wire n17121;
    wire n17125;
    wire n17127;
    wire n17131;
    wire n17133;
    wire n17136;
    wire n17139;
    wire n17143;
    wire n17146;
    wire n17149;
    wire n17151;
    wire n17155;
    wire n17158;
    wire n17160;
    wire n17164;
    wire n17166;
    wire n17169;
    wire n17172;
    wire n17175;
    wire n17178;
    wire n17181;
    wire n17184;
    wire n17187;
    wire n17190;
    wire n17193;
    wire n17196;
    wire n17199;
    wire n17202;
    wire n17205;
    wire n17208;
    wire n17212;
    wire n17214;
    wire n17217;
    wire n17221;
    wire n17224;
    wire n17227;
    wire n17230;
    wire n17233;
    wire n17236;
    wire n17238;
    wire n17241;
    wire n17244;
    wire n17247;
    wire n17250;
    wire n17253;
    wire n17256;
    wire n17259;
    wire n17263;
    wire n17266;
    wire n17269;
    wire n17272;
    wire n17274;
    wire n17278;
    wire n17280;
    wire n17283;
    wire n17286;
    wire n17289;
    wire n17292;
    wire n17295;
    wire n17298;
    wire n17302;
    wire n17305;
    wire n17307;
    wire n17310;
    wire n17313;
    wire n17316;
    wire n17319;
    wire n17322;
    wire n17325;
    wire n17328;
    wire n17331;
    wire n17334;
    wire n17337;
    wire n17340;
    wire n17343;
    wire n17346;
    wire n17349;
    wire n17352;
    wire n17355;
    wire n17358;
    wire n17361;
    wire n17364;
    wire n17367;
    wire n17370;
    wire n17373;
    wire n17377;
    wire n17379;
    wire n17383;
    wire n17386;
    wire n17389;
    wire n17392;
    wire n17395;
    wire n17397;
    wire n17400;
    wire n17403;
    wire n17406;
    wire n17409;
    wire n17412;
    wire n17415;
    wire n17418;
    wire n17421;
    wire n17424;
    wire n17427;
    wire n17430;
    wire n17433;
    wire n17436;
    wire n17439;
    wire n17442;
    wire n17445;
    wire n17448;
    wire n17451;
    wire n17454;
    wire n17457;
    wire n17460;
    wire n17463;
    wire n17466;
    wire n17469;
    wire n17473;
    wire n17476;
    wire n17479;
    wire n17482;
    wire n17485;
    wire n17488;
    wire n17491;
    wire n17493;
    wire n17497;
    wire n17500;
    wire n17503;
    wire n17506;
    wire n17509;
    wire n17512;
    wire n17515;
    wire n17517;
    wire n17520;
    wire n17523;
    wire n17526;
    wire n17529;
    wire n17532;
    wire n17535;
    wire n17538;
    wire n17541;
    wire n17545;
    wire n17547;
    wire n17550;
    wire n17553;
    wire n17556;
    wire n17559;
    wire n17562;
    wire n17566;
    wire n17569;
    wire n17572;
    wire n17575;
    wire n17578;
    wire n17581;
    wire n17584;
    wire n17587;
    wire n17590;
    wire n17593;
    wire n17595;
    wire n17598;
    wire n17601;
    wire n17604;
    wire n17607;
    wire n17610;
    wire n17613;
    wire n17616;
    wire n17619;
    wire n17622;
    wire n17625;
    wire n17628;
    wire n17631;
    wire n17634;
    wire n17637;
    wire n17640;
    wire n17643;
    wire n17646;
    wire n17649;
    wire n17652;
    wire n17655;
    wire n17658;
    wire n17661;
    wire n17664;
    wire n17668;
    wire n17671;
    wire n17673;
    wire n17676;
    wire n17679;
    wire n17683;
    wire n17685;
    wire n17688;
    wire n17691;
    wire n17694;
    wire n17697;
    wire n17700;
    wire n17703;
    wire n17706;
    wire n17709;
    wire n17712;
    wire n17715;
    wire n17718;
    wire n17721;
    wire n17724;
    wire n17727;
    wire n17730;
    wire n17733;
    wire n17736;
    wire n17739;
    wire n17742;
    wire n17745;
    wire n17748;
    wire n17752;
    wire n17755;
    wire n17757;
    wire n17760;
    wire n17763;
    wire n17766;
    wire n17769;
    wire n17772;
    wire n17775;
    wire n17779;
    wire n17782;
    wire n17784;
    wire n17787;
    wire n17790;
    wire n17793;
    wire n17796;
    wire n17799;
    wire n17802;
    wire n17805;
    wire n17808;
    wire n17811;
    wire n17814;
    wire n17818;
    wire n17820;
    wire n17824;
    wire n17827;
    wire n17829;
    wire n17832;
    wire n17836;
    wire n17838;
    wire n17841;
    wire n17844;
    wire n17847;
    wire n17850;
    wire n17853;
    wire n17856;
    wire n17859;
    wire n17862;
    wire n17865;
    wire n17868;
    wire n17871;
    wire n17874;
    wire n17877;
    wire n17880;
    wire n17884;
    wire n17887;
    wire n17889;
    wire n17892;
    wire n17896;
    wire n17898;
    wire n17901;
    wire n17904;
    wire n17908;
    wire n17910;
    wire n17913;
    wire n17916;
    wire n17919;
    wire n17922;
    wire n17925;
    wire n17928;
    wire n17931;
    wire n17934;
    wire n17937;
    wire n17940;
    wire n17943;
    wire n17946;
    wire n17949;
    wire n17952;
    wire n17955;
    wire n17958;
    wire n17961;
    wire n17964;
    wire n17967;
    wire n17970;
    wire n17973;
    wire n17976;
    wire n17979;
    wire n17983;
    wire n17985;
    wire n17988;
    wire n17991;
    wire n17994;
    wire n17997;
    wire n18000;
    wire n18003;
    wire n18006;
    wire n18009;
    wire n18012;
    wire n18015;
    wire n18018;
    wire n18021;
    wire n18024;
    wire n18027;
    wire n18030;
    wire n18033;
    wire n18036;
    wire n18039;
    wire n18042;
    wire n18045;
    wire n18048;
    wire n18051;
    wire n18054;
    wire n18057;
    wire n18060;
    wire n18063;
    wire n18066;
    wire n18069;
    wire n18072;
    wire n18075;
    wire n18078;
    wire n18081;
    wire n18084;
    wire n18087;
    wire n18090;
    wire n18094;
    wire n18096;
    wire n18099;
    wire n18102;
    wire n18105;
    wire n18108;
    wire n18111;
    wire n18114;
    wire n18117;
    wire n18120;
    wire n18123;
    wire n18126;
    wire n18129;
    wire n18132;
    wire n18135;
    wire n18138;
    wire n18141;
    wire n18144;
    wire n18147;
    wire n18150;
    wire n18153;
    wire n18156;
    wire n18159;
    wire n18162;
    wire n18165;
    wire n18168;
    wire n18171;
    wire n18174;
    wire n18177;
    wire n18180;
    wire n18183;
    wire n18186;
    wire n18189;
    wire n18192;
    wire n18196;
    wire n18199;
    wire n18202;
    wire n18205;
    wire n18208;
    wire n18211;
    wire n18214;
    wire n18217;
    wire n18220;
    wire n18223;
    wire n18226;
    wire n18229;
    wire n18232;
    wire n18235;
    wire n18238;
    wire n18241;
    wire n18244;
    wire n18247;
    wire n18250;
    wire n18253;
    wire n18256;
    wire n18259;
    wire n18262;
    wire n18265;
    wire n18268;
    wire n18271;
    wire n18274;
    wire n18277;
    wire n18280;
    wire n18282;
    wire n18285;
    wire n18288;
    wire n18292;
    wire n18295;
    wire n18298;
    wire n18301;
    wire n18304;
    wire n18307;
    wire n18310;
    wire n18313;
    wire n18316;
    wire n18319;
    wire n18321;
    wire n18324;
    wire n18327;
    wire n18330;
    wire n18333;
    wire n18336;
    wire n18339;
    wire n18342;
    wire n18345;
    wire n18348;
    wire n18351;
    wire n18354;
    wire n18357;
    wire n18361;
    wire n18363;
    wire n18366;
    wire n18369;
    wire n18372;
    wire n18375;
    wire n18379;
    wire n18382;
    wire n18385;
    wire n18388;
    wire n18391;
    wire n18393;
    wire n18396;
    wire n18399;
    wire n18402;
    wire n18405;
    wire n18408;
    wire n18411;
    wire n18414;
    wire n18417;
    wire n18420;
    wire n18423;
    wire n18426;
    wire n18429;
    wire n18432;
    wire n18435;
    wire n18438;
    wire n18441;
    wire n18444;
    wire n18447;
    wire n18450;
    wire n18453;
    wire n18456;
    wire n18459;
    wire n18462;
    wire n18466;
    wire n18469;
    wire n18471;
    wire n18474;
    wire n18477;
    wire n18480;
    wire n18483;
    wire n18486;
    wire n18489;
    wire n18492;
    wire n18495;
    wire n18498;
    wire n18501;
    wire n18505;
    wire n18508;
    wire n18510;
    wire n18513;
    wire n18516;
    wire n18519;
    wire n18522;
    wire n18526;
    wire n18529;
    wire n18531;
    wire n18534;
    wire n18537;
    wire n18540;
    wire n18543;
    wire n18546;
    wire n18549;
    wire n18552;
    wire n18555;
    wire n18558;
    wire n18562;
    wire n18564;
    wire n18568;
    wire n18571;
    wire n18574;
    wire n18577;
    wire n18579;
    wire n18582;
    wire n18585;
    wire n18589;
    wire n18592;
    wire n18595;
    wire n18597;
    wire n18600;
    wire n18603;
    wire n18606;
    wire n18609;
    wire n18612;
    wire n18615;
    wire n18618;
    wire n18621;
    wire n18624;
    wire n18627;
    wire n18630;
    wire n18633;
    wire n18636;
    wire n18639;
    wire n18642;
    wire n18646;
    wire n18649;
    wire n18652;
    wire n18655;
    wire n18658;
    wire n18661;
    wire n18664;
    wire n18667;
    wire n18670;
    wire n18673;
    wire n18676;
    wire n18679;
    wire n18682;
    wire n18685;
    wire n18687;
    wire n18690;
    wire n18694;
    wire n18697;
    wire n18700;
    wire n18703;
    wire n18706;
    wire n18709;
    wire n18712;
    wire n18715;
    wire n18718;
    wire n18721;
    wire n18724;
    wire n18727;
    wire n18729;
    wire n18732;
    wire n18735;
    wire n18738;
    wire n18741;
    wire n18744;
    wire n18747;
    wire n18750;
    wire n18753;
    wire n18756;
    wire n18759;
    wire n18762;
    wire n18765;
    wire n18768;
    wire n18771;
    wire n18774;
    wire n18777;
    wire n18780;
    wire n18783;
    wire n18786;
    wire n18789;
    wire n18792;
    wire n18795;
    wire n18798;
    wire n18801;
    wire n18804;
    wire n18807;
    wire n18811;
    wire n18814;
    wire n18817;
    wire n18820;
    wire n18823;
    wire n18826;
    wire n18828;
    wire n18831;
    wire n18834;
    wire n18837;
    wire n18840;
    wire n18843;
    wire n18846;
    wire n18849;
    wire n18852;
    wire n18855;
    wire n18858;
    wire n18861;
    wire n18864;
    wire n18867;
    wire n18870;
    wire n18874;
    wire n18877;
    wire n18880;
    wire n18883;
    wire n18886;
    wire n18889;
    wire n18892;
    wire n18894;
    wire n18897;
    wire n18900;
    wire n18903;
    wire n18906;
    wire n18909;
    wire n18912;
    wire n18915;
    wire n18918;
    wire n18921;
    wire n18924;
    wire n18927;
    wire n18930;
    wire n18933;
    wire n18936;
    wire n18940;
    wire n18943;
    wire n18945;
    wire n18948;
    wire n18951;
    wire n18954;
    wire n18958;
    wire n18961;
    wire n18964;
    wire n18966;
    wire n18969;
    wire n18972;
    wire n18976;
    wire n18978;
    wire n18981;
    wire n18984;
    wire n18988;
    wire n18990;
    wire n18993;
    wire n18996;
    wire n19000;
    wire n19002;
    wire n19005;
    wire n19008;
    wire n19011;
    wire n19015;
    wire n19017;
    wire n19020;
    wire n19023;
    wire n19027;
    wire n19030;
    wire n19033;
    wire n19035;
    wire n19038;
    wire n19041;
    wire n19045;
    wire n19047;
    wire n19050;
    wire n19053;
    wire n19056;
    wire n19059;
    wire n19062;
    wire n19065;
    wire n19068;
    wire n19071;
    wire n19074;
    wire n19077;
    wire n19080;
    wire n19083;
    wire n19086;
    wire n19089;
    wire n19093;
    wire n19095;
    wire n19098;
    wire n19101;
    wire n19105;
    wire n19107;
    wire n19110;
    wire n19113;
    wire n19116;
    wire n19119;
    wire n19122;
    wire n19125;
    wire n19129;
    wire n19131;
    wire n19134;
    wire n19137;
    wire n19140;
    wire n19143;
    wire n19146;
    wire n19149;
    wire n19152;
    wire n19156;
    wire n19159;
    wire n19161;
    wire n19164;
    wire n19167;
    wire n19170;
    wire n19174;
    wire n19176;
    wire n19179;
    wire n19182;
    wire n19185;
    wire n19188;
    wire n19191;
    wire n19194;
    wire n19197;
    wire n19200;
    wire n19203;
    wire n19206;
    wire n19210;
    wire n19213;
    wire n19216;
    wire n19218;
    wire n19221;
    wire n19224;
    wire n19227;
    wire n19230;
    wire n19233;
    wire n19236;
    wire n19239;
    wire n19242;
    wire n19245;
    wire n19248;
    wire n19251;
    wire n19254;
    wire n19258;
    wire n19261;
    wire n19264;
    wire n19267;
    wire n19269;
    wire n19272;
    wire n19275;
    wire n19278;
    wire n19282;
    wire n19284;
    wire n19287;
    wire n19290;
    wire n19293;
    wire n19296;
    wire n19299;
    wire n19302;
    wire n19305;
    wire n19308;
    wire n19311;
    wire n19314;
    wire n19317;
    wire n19320;
    wire n19323;
    wire n19326;
    wire n19330;
    wire n19333;
    wire n19335;
    wire n19338;
    wire n19341;
    wire n19345;
    wire n19347;
    wire n19350;
    wire n19353;
    wire n19356;
    wire n19359;
    wire n19362;
    wire n19365;
    wire n19368;
    wire n19371;
    wire n19374;
    wire n19377;
    wire n19380;
    wire n19383;
    wire n19386;
    wire n19389;
    wire n19393;
    wire n19395;
    wire n19398;
    wire n19401;
    wire n19405;
    wire n19407;
    wire n19410;
    wire n19413;
    wire n19416;
    wire n19419;
    wire n19422;
    wire n19425;
    wire n19429;
    wire n19431;
    wire n19434;
    wire n19437;
    wire n19440;
    wire n19443;
    wire n19446;
    wire n19449;
    wire n19452;
    wire n19455;
    wire n19458;
    wire n19461;
    wire n19465;
    wire n19468;
    wire n19470;
    wire n19473;
    wire n19476;
    wire n19479;
    wire n19482;
    wire n19486;
    wire n19488;
    wire n19491;
    wire n19494;
    wire n19497;
    wire n19500;
    wire n19503;
    wire n19506;
    wire n19509;
    wire n19512;
    wire n19515;
    wire n19518;
    wire n19521;
    wire n19524;
    wire n19527;
    wire n19530;
    wire n19533;
    wire n19536;
    wire n19539;
    wire n19543;
    wire n19546;
    wire n19548;
    wire n19551;
    wire n19554;
    wire n19557;
    wire n19560;
    wire n19563;
    wire n19566;
    wire n19570;
    wire n19572;
    wire n19575;
    wire n19578;
    wire n19581;
    wire n19584;
    wire n19587;
    wire n19590;
    wire n19593;
    wire n19596;
    wire n19599;
    wire n19602;
    wire n19605;
    wire n19608;
    wire n19611;
    wire n19614;
    wire n19617;
    wire n19620;
    wire n19623;
    wire n19626;
    wire n19629;
    wire n19632;
    wire n19635;
    wire n19638;
    wire n19641;
    wire n19644;
    wire n19647;
    wire n19650;
    wire n19653;
    wire n19656;
    wire n19659;
    wire n19662;
    wire n19665;
    wire n19668;
    wire n19671;
    wire n19674;
    wire n19677;
    wire n19680;
    wire n19683;
    wire n19686;
    wire n19689;
    wire n19692;
    wire n19695;
    wire n19698;
    wire n19701;
    wire n19704;
    wire n19707;
    wire n19710;
    wire n19713;
    wire n19716;
    wire n19719;
    wire n19722;
    wire n19725;
    wire n19728;
    wire n19731;
    wire n19734;
    wire n19737;
    wire n19740;
    wire n19743;
    wire n19746;
    wire n19749;
    wire n19752;
    wire n19755;
    wire n19758;
    wire n19761;
    wire n19764;
    wire n19767;
    wire n19770;
    wire n19773;
    wire n19776;
    wire n19779;
    wire n19782;
    wire n19785;
    wire n19788;
    wire n19791;
    wire n19794;
    wire n19797;
    wire n19800;
    wire n19803;
    wire n19806;
    wire n19809;
    wire n19812;
    wire n19815;
    wire n19818;
    wire n19821;
    wire n19824;
    wire n19827;
    wire n19830;
    wire n19833;
    wire n19836;
    wire n19839;
    wire n19842;
    wire n19845;
    wire n19848;
    wire n19851;
    wire n19854;
    wire n19857;
    wire n19860;
    wire n19863;
    wire n19866;
    wire n19869;
    wire n19872;
    wire n19875;
    wire n19878;
    wire n19881;
    wire n19884;
    wire n19887;
    wire n19890;
    wire n19893;
    wire n19896;
    wire n19899;
    wire n19902;
    wire n19905;
    wire n19908;
    wire n19911;
    wire n19914;
    wire n19917;
    wire n19920;
    wire n19923;
    wire n19926;
    wire n19929;
    wire n19932;
    wire n19935;
    wire n19938;
    wire n19941;
    wire n19944;
    wire n19947;
    wire n19950;
    wire n19953;
    wire n19956;
    wire n19959;
    wire n19962;
    wire n19965;
    wire n19968;
    wire n19971;
    wire n19974;
    wire n19977;
    wire n19980;
    wire n19983;
    wire n19986;
    wire n19989;
    wire n19992;
    wire n19995;
    wire n19998;
    wire n20001;
    wire n20004;
    wire n20007;
    wire n20010;
    wire n20013;
    wire n20016;
    wire n20019;
    wire n20022;
    wire n20025;
    wire n20028;
    wire n20031;
    wire n20034;
    wire n20037;
    wire n20040;
    wire n20043;
    wire n20046;
    wire n20049;
    wire n20052;
    wire n20055;
    wire n20058;
    wire n20061;
    wire n20064;
    wire n20067;
    wire n20070;
    wire n20073;
    wire n20076;
    wire n20079;
    wire n20082;
    wire n20085;
    wire n20088;
    wire n20091;
    wire n20094;
    wire n20097;
    wire n20100;
    wire n20103;
    wire n20106;
    wire n20109;
    wire n20112;
    wire n20115;
    wire n20118;
    wire n20121;
    wire n20124;
    wire n20127;
    wire n20130;
    wire n20133;
    wire n20136;
    wire n20139;
    wire n20142;
    wire n20145;
    wire n20148;
    wire n20151;
    wire n20154;
    wire n20157;
    wire n20160;
    wire n20163;
    wire n20166;
    wire n20169;
    wire n20172;
    wire n20175;
    wire n20178;
    wire n20181;
    wire n20184;
    wire n20187;
    wire n20190;
    wire n20193;
    wire n20196;
    wire n20199;
    wire n20202;
    wire n20205;
    wire n20208;
    wire n20211;
    wire n20214;
    wire n20217;
    wire n20220;
    wire n20224;
    wire n20227;
    wire n20229;
    wire n20232;
    wire n20235;
    wire n20238;
    wire n20241;
    wire n20244;
    wire n20247;
    wire n20250;
    wire n20253;
    wire n20256;
    wire n20259;
    wire n20262;
    wire n20265;
    wire n20268;
    wire n20271;
    wire n20274;
    wire n20277;
    wire n20280;
    wire n20283;
    wire n20286;
    wire n20289;
    wire n20292;
    wire n20295;
    wire n20298;
    wire n20301;
    wire n20304;
    wire n20307;
    wire n20310;
    wire n20313;
    wire n20316;
    wire n20319;
    wire n20322;
    wire n20325;
    wire n20328;
    wire n20331;
    wire n20334;
    wire n20337;
    wire n20340;
    wire n20343;
    wire n20346;
    wire n20349;
    wire n20352;
    wire n20355;
    wire n20358;
    wire n20361;
    wire n20364;
    wire n20367;
    wire n20370;
    wire n20373;
    wire n20376;
    wire n20379;
    wire n20382;
    wire n20385;
    wire n20388;
    wire n20391;
    wire n20394;
    wire n20397;
    wire n20400;
    wire n20403;
    wire n20406;
    wire n20409;
    wire n20412;
    wire n20415;
    wire n20418;
    wire n20421;
    wire n20424;
    wire n20427;
    wire n20430;
    wire n20433;
    wire n20436;
    wire n20439;
    wire n20442;
    wire n20445;
    wire n20448;
    wire n20451;
    wire n20454;
    wire n20457;
    wire n20460;
    wire n20463;
    wire n20466;
    wire n20469;
    wire n20472;
    wire n20475;
    wire n20478;
    wire n20481;
    wire n20484;
    wire n20487;
    wire n20490;
    wire n20493;
    wire n20496;
    wire n20499;
    wire n20502;
    wire n20505;
    wire n20508;
    wire n20511;
    wire n20514;
    wire n20517;
    wire n20520;
    wire n20523;
    wire n20526;
    wire n20529;
    wire n20532;
    wire n20535;
    wire n20538;
    wire n20541;
    wire n20544;
    wire n20547;
    wire n20550;
    wire n20554;
    wire n20557;
    wire n20560;
    wire n20563;
    wire n20566;
    wire n20569;
    wire n20572;
    wire n20575;
    wire n20578;
    wire n20581;
    wire n20584;
    wire n20587;
    wire n20590;
    wire n20593;
    wire n20596;
    wire n20599;
    wire n20602;
    wire n20605;
    wire n20608;
    wire n20611;
    wire n20614;
    wire n20617;
    wire n20620;
    wire n20623;
    wire n20626;
    wire n20629;
    wire n20632;
    wire n20634;
    wire n20637;
    wire n20640;
    wire n20643;
    wire n20646;
    wire n20649;
    wire n20652;
    wire n20655;
    wire n20658;
    wire n20661;
    wire n20664;
    wire n20667;
    wire n20670;
    wire n20673;
    wire n20676;
    wire n20679;
    wire n20682;
    wire n20685;
    wire n20688;
    wire n20691;
    wire n20694;
    wire n20697;
    wire n20700;
    wire n20703;
    wire n20706;
    wire n20709;
    wire n20712;
    wire n20715;
    wire n20718;
    wire n20721;
    wire n20724;
    wire n20727;
    wire n20730;
    wire n20733;
    wire n20736;
    wire n20739;
    wire n20742;
    wire n20745;
    wire n20748;
    wire n20751;
    wire n20754;
    wire n20757;
    wire n20760;
    wire n20763;
    wire n20766;
    wire n20769;
    wire n20772;
    wire n20775;
    wire n20778;
    wire n20781;
    wire n20784;
    wire n20787;
    wire n20790;
    wire n20793;
    wire n20796;
    wire n20799;
    wire n20802;
    wire n20805;
    wire n20808;
    wire n20811;
    wire n20814;
    wire n20817;
    wire n20820;
    wire n20823;
    wire n20826;
    wire n20829;
    wire n20832;
    wire n20835;
    wire n20838;
    wire n20841;
    wire n20844;
    wire n20847;
    wire n20850;
    wire n20853;
    wire n20856;
    wire n20859;
    wire n20862;
    wire n20865;
    wire n20868;
    wire n20871;
    wire n20874;
    wire n20877;
    wire n20883;
    wire n20886;
    wire n20889;
    wire n20892;
    wire n20895;
    wire n20898;
    wire n20901;
    wire n20904;
    wire n20907;
    wire n20910;
    wire n20913;
    wire n20916;
    wire n20919;
    wire n20922;
    wire n20925;
    wire n20928;
    wire n20931;
    wire n20934;
    wire n20937;
    wire n20940;
    wire n20943;
    wire n20946;
    wire n20949;
    wire n20952;
    wire n20955;
    wire n20958;
    wire n20964;
    wire n20967;
    wire n20970;
    wire n20973;
    wire n20976;
    wire n20979;
    wire n20982;
    wire n20985;
    wire n20988;
    wire n20991;
    wire n20994;
    wire n20997;
    wire n21000;
    wire n21003;
    wire n21006;
    wire n21009;
    wire n21012;
    wire n21015;
    wire n21018;
    wire n21021;
    wire n21024;
    wire n21027;
    wire n21030;
    wire n21033;
    wire n21036;
    wire n21039;
    wire n21045;
    wire n21048;
    wire n21051;
    wire n21054;
    wire n21057;
    wire n21060;
    wire n21063;
    wire n21066;
    wire n21069;
    wire n21072;
    wire n21075;
    wire n21078;
    wire n21081;
    wire n21084;
    wire n21087;
    wire n21090;
    wire n21093;
    wire n21096;
    wire n21099;
    wire n21102;
    wire n21105;
    wire n21108;
    wire n21111;
    wire n21114;
    wire n21117;
    wire n21120;
    wire n21126;
    wire n21129;
    wire n21132;
    wire n21135;
    wire n21138;
    wire n21141;
    wire n21144;
    wire n21147;
    wire n21150;
    wire n21153;
    wire n21156;
    wire n21159;
    wire n21162;
    wire n21165;
    wire n21168;
    wire n21171;
    wire n21174;
    wire n21177;
    wire n21180;
    wire n21183;
    wire n21186;
    wire n21189;
    wire n21192;
    wire n21195;
    wire n21198;
    wire n21201;
    wire n21207;
    wire n21210;
    wire n21213;
    wire n21216;
    wire n21219;
    wire n21222;
    wire n21225;
    wire n21228;
    wire n21231;
    wire n21234;
    wire n21237;
    wire n21240;
    wire n21243;
    wire n21246;
    wire n21249;
    wire n21252;
    wire n21255;
    wire n21258;
    wire n21261;
    wire n21264;
    wire n21267;
    wire n21270;
    wire n21273;
    wire n21276;
    wire n21279;
    wire n21282;
    wire n21288;
    wire n21291;
    wire n21294;
    wire n21297;
    wire n21300;
    wire n21303;
    wire n21306;
    wire n21309;
    wire n21312;
    wire n21315;
    wire n21318;
    wire n21321;
    wire n21324;
    wire n21327;
    wire n21330;
    wire n21333;
    wire n21336;
    wire n21339;
    wire n21342;
    wire n21345;
    wire n21348;
    wire n21351;
    wire n21354;
    wire n21357;
    wire n21360;
    wire n21363;
    wire n21369;
    wire n21372;
    wire n21375;
    wire n21378;
    wire n21381;
    wire n21384;
    wire n21387;
    wire n21390;
    wire n21393;
    wire n21396;
    wire n21399;
    wire n21402;
    wire n21405;
    wire n21408;
    wire n21411;
    wire n21414;
    wire n21417;
    wire n21420;
    wire n21423;
    wire n21426;
    wire n21429;
    wire n21432;
    wire n21435;
    wire n21438;
    wire n21441;
    wire n21444;
    wire n21450;
    wire n21453;
    wire n21456;
    wire n21459;
    wire n21462;
    wire n21465;
    wire n21468;
    wire n21471;
    wire n21474;
    wire n21477;
    wire n21480;
    wire n21483;
    wire n21486;
    wire n21489;
    wire n21492;
    wire n21495;
    wire n21498;
    wire n21501;
    wire n21504;
    wire n21507;
    wire n21510;
    wire n21513;
    wire n21516;
    wire n21519;
    wire n21522;
    wire n21525;
    wire n21531;
    wire n21534;
    wire n21537;
    wire n21540;
    wire n21543;
    wire n21546;
    wire n21549;
    wire n21552;
    wire n21555;
    wire n21558;
    wire n21561;
    wire n21564;
    wire n21567;
    wire n21570;
    wire n21573;
    wire n21576;
    wire n21579;
    wire n21582;
    wire n21585;
    wire n21588;
    wire n21591;
    wire n21594;
    wire n21597;
    wire n21600;
    wire n21603;
    wire n21606;
    wire n21612;
    wire n21615;
    wire n21618;
    wire n21621;
    wire n21624;
    wire n21627;
    wire n21630;
    wire n21633;
    wire n21636;
    wire n21639;
    wire n21642;
    wire n21645;
    wire n21648;
    wire n21651;
    wire n21654;
    wire n21657;
    wire n21660;
    wire n21663;
    wire n21666;
    wire n21669;
    wire n21672;
    wire n21675;
    wire n21678;
    wire n21681;
    wire n21684;
    wire n21687;
    wire n21693;
    wire n21696;
    wire n21699;
    wire n21702;
    wire n21705;
    wire n21708;
    wire n21711;
    wire n21714;
    wire n21717;
    wire n21720;
    wire n21723;
    wire n21726;
    wire n21729;
    wire n21732;
    wire n21735;
    wire n21738;
    wire n21741;
    wire n21744;
    wire n21747;
    wire n21750;
    wire n21753;
    wire n21756;
    wire n21759;
    wire n21762;
    wire n21765;
    wire n21768;
    wire n21774;
    wire n21777;
    wire n21780;
    wire n21783;
    wire n21786;
    wire n21789;
    wire n21792;
    wire n21795;
    wire n21798;
    wire n21801;
    wire n21804;
    wire n21807;
    wire n21810;
    wire n21813;
    wire n21816;
    wire n21819;
    wire n21822;
    wire n21825;
    wire n21828;
    wire n21831;
    wire n21834;
    wire n21837;
    wire n21840;
    wire n21843;
    wire n21846;
    wire n21849;
    wire n21855;
    wire n21858;
    wire n21861;
    wire n21864;
    wire n21867;
    wire n21870;
    wire n21873;
    wire n21876;
    wire n21879;
    wire n21882;
    wire n21885;
    wire n21888;
    wire n21891;
    wire n21894;
    wire n21897;
    wire n21900;
    wire n21903;
    wire n21906;
    wire n21909;
    wire n21912;
    wire n21915;
    wire n21918;
    wire n21921;
    wire n21924;
    wire n21927;
    wire n21930;
    wire n21936;
    wire n21939;
    wire n21942;
    wire n21945;
    wire n21948;
    wire n21951;
    wire n21954;
    wire n21957;
    wire n21960;
    wire n21963;
    wire n21966;
    wire n21969;
    wire n21972;
    wire n21975;
    wire n21978;
    wire n21981;
    wire n21984;
    wire n21987;
    wire n21990;
    wire n21993;
    wire n21996;
    wire n21999;
    wire n22002;
    wire n22005;
    wire n22008;
    wire n22011;
    wire n22017;
    wire n22020;
    wire n22023;
    wire n22026;
    wire n22029;
    wire n22032;
    wire n22035;
    wire n22038;
    wire n22041;
    wire n22044;
    wire n22047;
    wire n22050;
    wire n22053;
    wire n22056;
    wire n22059;
    wire n22062;
    wire n22065;
    wire n22068;
    wire n22071;
    wire n22074;
    wire n22077;
    wire n22080;
    wire n22083;
    wire n22086;
    wire n22089;
    wire n22092;
    wire n22098;
    wire n22101;
    wire n22104;
    wire n22107;
    wire n22110;
    wire n22113;
    wire n22116;
    wire n22119;
    wire n22122;
    wire n22125;
    wire n22128;
    wire n22131;
    wire n22134;
    wire n22137;
    wire n22140;
    wire n22143;
    wire n22146;
    wire n22149;
    wire n22152;
    wire n22155;
    wire n22158;
    wire n22161;
    wire n22164;
    wire n22167;
    wire n22170;
    wire n22173;
    wire n22179;
    wire n22182;
    wire n22185;
    wire n22188;
    wire n22191;
    wire n22194;
    wire n22197;
    wire n22200;
    wire n22203;
    wire n22206;
    wire n22209;
    wire n22212;
    wire n22215;
    wire n22218;
    wire n22221;
    wire n22224;
    wire n22227;
    wire n22230;
    wire n22233;
    wire n22236;
    wire n22239;
    wire n22242;
    wire n22245;
    wire n22248;
    wire n22251;
    wire n22254;
    wire n22260;
    wire n22263;
    wire n22266;
    wire n22269;
    wire n22272;
    wire n22275;
    wire n22278;
    wire n22281;
    wire n22284;
    wire n22287;
    wire n22290;
    wire n22293;
    wire n22296;
    wire n22299;
    wire n22302;
    wire n22305;
    wire n22308;
    wire n22311;
    wire n22314;
    wire n22317;
    wire n22320;
    wire n22323;
    wire n22326;
    wire n22329;
    wire n22332;
    wire n22338;
    wire n22341;
    wire n22344;
    wire n22347;
    wire n22350;
    wire n22353;
    wire n22356;
    wire n22359;
    wire n22362;
    wire n22365;
    wire n22368;
    wire n22371;
    wire n22374;
    wire n22377;
    wire n22380;
    wire n22383;
    wire n22386;
    wire n22389;
    wire n22392;
    wire n22395;
    wire n22398;
    wire n22401;
    wire n22404;
    wire n22407;
    wire n22410;
    wire n22416;
    wire n22419;
    wire n22422;
    wire n22425;
    wire n22428;
    wire n22431;
    wire n22434;
    wire n22437;
    wire n22440;
    wire n22443;
    wire n22446;
    wire n22449;
    wire n22452;
    wire n22455;
    wire n22458;
    wire n22461;
    wire n22464;
    wire n22467;
    wire n22470;
    wire n22473;
    wire n22476;
    wire n22479;
    wire n22482;
    wire n22485;
    wire n22488;
    wire n22494;
    wire n22497;
    wire n22500;
    wire n22503;
    wire n22506;
    wire n22509;
    wire n22512;
    wire n22515;
    wire n22518;
    wire n22521;
    wire n22524;
    wire n22527;
    wire n22530;
    wire n22533;
    wire n22536;
    wire n22539;
    wire n22542;
    wire n22545;
    wire n22548;
    wire n22551;
    wire n22554;
    wire n22557;
    wire n22560;
    wire n22563;
    wire n22566;
    wire n22569;
    wire n22575;
    wire n22578;
    wire n22581;
    wire n22584;
    wire n22587;
    wire n22590;
    wire n22593;
    wire n22596;
    wire n22599;
    wire n22602;
    wire n22605;
    wire n22608;
    wire n22611;
    wire n22614;
    wire n22617;
    wire n22620;
    wire n22623;
    wire n22626;
    wire n22629;
    wire n22632;
    wire n22635;
    wire n22638;
    wire n22641;
    wire n22644;
    wire n22647;
    wire n22650;
    wire n22656;
    wire n22659;
    wire n22662;
    wire n22665;
    wire n22668;
    wire n22671;
    wire n22674;
    wire n22677;
    wire n22680;
    wire n22683;
    wire n22686;
    wire n22689;
    wire n22692;
    wire n22695;
    wire n22698;
    wire n22701;
    wire n22704;
    wire n22707;
    wire n22710;
    wire n22713;
    wire n22716;
    wire n22719;
    wire n22722;
    wire n22725;
    wire n22728;
    wire n22731;
    wire n22737;
    wire n22740;
    wire n22743;
    wire n22746;
    wire n22749;
    wire n22752;
    wire n22755;
    wire n22758;
    wire n22761;
    wire n22764;
    wire n22767;
    wire n22770;
    wire n22773;
    wire n22776;
    wire n22779;
    wire n22782;
    wire n22785;
    wire n22788;
    wire n22791;
    wire n22794;
    wire n22797;
    wire n22800;
    wire n22803;
    wire n22806;
    wire n22809;
    wire n22812;
    wire n22818;
    wire n22821;
    wire n22824;
    wire n22827;
    wire n22830;
    wire n22833;
    wire n22836;
    wire n22839;
    wire n22842;
    wire n22845;
    wire n22848;
    wire n22851;
    wire n22854;
    wire n22857;
    wire n22860;
    wire n22863;
    wire n22866;
    wire n22869;
    wire n22872;
    wire n22875;
    wire n22878;
    wire n22881;
    wire n22884;
    wire n22887;
    wire n22890;
    wire n22893;
    wire n22899;
    wire n22902;
    wire n22905;
    wire n22908;
    wire n22911;
    wire n22914;
    wire n22917;
    wire n22920;
    wire n22923;
    wire n22926;
    wire n22929;
    wire n22932;
    wire n22935;
    wire n22938;
    wire n22941;
    wire n22944;
    wire n22947;
    wire n22950;
    wire n22953;
    wire n22956;
    wire n22959;
    wire n22962;
    wire n22965;
    wire n22968;
    wire n22971;
    wire n22974;
    wire n22980;
    wire n22983;
    wire n22986;
    wire n22989;
    wire n22992;
    wire n22995;
    wire n22998;
    wire n23001;
    wire n23004;
    wire n23007;
    wire n23010;
    wire n23013;
    wire n23016;
    wire n23019;
    wire n23022;
    wire n23025;
    wire n23028;
    wire n23031;
    wire n23034;
    wire n23037;
    wire n23040;
    wire n23043;
    wire n23046;
    wire n23049;
    wire n23055;
    wire n23058;
    wire n23061;
    wire n23064;
    wire n23067;
    wire n23070;
    wire n23073;
    wire n23076;
    wire n23079;
    wire n23082;
    wire n23085;
    wire n23088;
    wire n23091;
    wire n23094;
    wire n23097;
    wire n23100;
    wire n23103;
    wire n23106;
    wire n23109;
    wire n23112;
    wire n23115;
    wire n23118;
    wire n23121;
    wire n23124;
    wire n23127;
    wire n23133;
    wire n23136;
    wire n23139;
    wire n23142;
    wire n23145;
    wire n23148;
    wire n23151;
    wire n23154;
    wire n23157;
    wire n23160;
    wire n23163;
    wire n23166;
    wire n23169;
    wire n23172;
    wire n23175;
    wire n23178;
    wire n23181;
    wire n23184;
    wire n23187;
    wire n23190;
    wire n23193;
    wire n23196;
    wire n23199;
    wire n23202;
    wire n23205;
    wire n23208;
    wire n23214;
    wire n23217;
    wire n23220;
    wire n23223;
    wire n23226;
    wire n23229;
    wire n23232;
    wire n23235;
    wire n23238;
    wire n23241;
    wire n23244;
    wire n23247;
    wire n23250;
    wire n23253;
    wire n23256;
    wire n23259;
    wire n23262;
    wire n23265;
    wire n23268;
    wire n23271;
    wire n23274;
    wire n23277;
    wire n23280;
    wire n23283;
    wire n23286;
    wire n23289;
    wire n23295;
    wire n23298;
    wire n23301;
    wire n23304;
    wire n23307;
    wire n23310;
    wire n23313;
    wire n23316;
    wire n23319;
    wire n23322;
    wire n23325;
    wire n23328;
    wire n23331;
    wire n23334;
    wire n23337;
    wire n23340;
    wire n23343;
    wire n23346;
    wire n23349;
    wire n23352;
    wire n23355;
    wire n23358;
    wire n23361;
    wire n23364;
    wire n23367;
    wire n23370;
    wire n23376;
    wire n23379;
    wire n23382;
    wire n23385;
    wire n23388;
    wire n23391;
    wire n23394;
    wire n23397;
    wire n23400;
    wire n23403;
    wire n23406;
    wire n23409;
    wire n23412;
    wire n23415;
    wire n23418;
    wire n23421;
    wire n23424;
    wire n23427;
    wire n23430;
    wire n23433;
    wire n23436;
    wire n23439;
    wire n23442;
    wire n23445;
    wire n23448;
    wire n23451;
    wire n23457;
    wire n23460;
    wire n23463;
    wire n23466;
    wire n23469;
    wire n23472;
    wire n23475;
    wire n23478;
    wire n23481;
    wire n23484;
    wire n23487;
    wire n23490;
    wire n23493;
    wire n23496;
    wire n23499;
    wire n23502;
    wire n23505;
    wire n23508;
    wire n23511;
    wire n23514;
    wire n23517;
    wire n23520;
    wire n23523;
    wire n23526;
    wire n23529;
    wire n23532;
    wire n23538;
    wire n23541;
    wire n23544;
    wire n23547;
    wire n23550;
    wire n23553;
    wire n23556;
    wire n23559;
    wire n23562;
    wire n23565;
    wire n23568;
    wire n23571;
    wire n23574;
    wire n23577;
    wire n23580;
    wire n23583;
    wire n23586;
    wire n23589;
    wire n23592;
    wire n23595;
    wire n23598;
    wire n23601;
    wire n23604;
    wire n23607;
    wire n23610;
    wire n23613;
    wire n23619;
    wire n23622;
    wire n23625;
    wire n23628;
    wire n23631;
    wire n23634;
    wire n23637;
    wire n23640;
    wire n23643;
    wire n23646;
    wire n23649;
    wire n23652;
    wire n23655;
    wire n23658;
    wire n23661;
    wire n23664;
    wire n23667;
    wire n23670;
    wire n23673;
    wire n23676;
    wire n23679;
    wire n23682;
    wire n23685;
    wire n23691;
    wire n23694;
    wire n23697;
    wire n23700;
    wire n23703;
    wire n23706;
    wire n23709;
    wire n23712;
    wire n23715;
    wire n23718;
    wire n23721;
    wire n23724;
    wire n23727;
    wire n23730;
    wire n23733;
    wire n23736;
    wire n23739;
    wire n23742;
    wire n23745;
    wire n23748;
    wire n23751;
    wire n23754;
    wire n23757;
    wire n23763;
    wire n23766;
    wire n23769;
    wire n23772;
    wire n23775;
    wire n23778;
    wire n23781;
    wire n23784;
    wire n23787;
    wire n23790;
    wire n23793;
    wire n23796;
    wire n23799;
    wire n23802;
    wire n23805;
    wire n23808;
    wire n23811;
    wire n23814;
    wire n23817;
    wire n23820;
    wire n23823;
    wire n23826;
    wire n23829;
    wire n23835;
    wire n23838;
    wire n23841;
    wire n23844;
    wire n23847;
    wire n23850;
    wire n23853;
    wire n23856;
    wire n23859;
    wire n23862;
    wire n23865;
    wire n23868;
    wire n23871;
    wire n23874;
    wire n23877;
    wire n23880;
    wire n23883;
    wire n23886;
    wire n23889;
    wire n23892;
    wire n23895;
    wire n23898;
    wire n23901;
    wire n23904;
    wire n23910;
    wire n23913;
    wire n23916;
    wire n23919;
    wire n23922;
    wire n23925;
    wire n23928;
    wire n23931;
    wire n23934;
    wire n23937;
    wire n23940;
    wire n23943;
    wire n23946;
    wire n23949;
    wire n23952;
    wire n23955;
    wire n23958;
    wire n23961;
    wire n23964;
    wire n23967;
    wire n23970;
    wire n23973;
    wire n23979;
    wire n23982;
    wire n23985;
    wire n23988;
    wire n23991;
    wire n23994;
    wire n23997;
    wire n24000;
    wire n24003;
    wire n24006;
    wire n24009;
    wire n24012;
    wire n24015;
    wire n24018;
    wire n24021;
    wire n24024;
    wire n24027;
    wire n24030;
    wire n24033;
    wire n24036;
    wire n24039;
    wire n24042;
    wire n24048;
    wire n24051;
    wire n24054;
    wire n24057;
    wire n24060;
    wire n24063;
    wire n24066;
    wire n24069;
    wire n24072;
    wire n24075;
    wire n24078;
    wire n24081;
    wire n24084;
    wire n24087;
    wire n24090;
    wire n24093;
    wire n24096;
    wire n24099;
    wire n24102;
    wire n24105;
    wire n24108;
    wire n24111;
    wire n24117;
    wire n24120;
    wire n24123;
    wire n24126;
    wire n24129;
    wire n24132;
    wire n24135;
    wire n24138;
    wire n24141;
    wire n24144;
    wire n24147;
    wire n24150;
    wire n24153;
    wire n24156;
    wire n24159;
    wire n24162;
    wire n24165;
    wire n24168;
    wire n24171;
    wire n24174;
    wire n24177;
    wire n24180;
    wire n24186;
    wire n24189;
    wire n24192;
    wire n24195;
    wire n24198;
    wire n24201;
    wire n24204;
    wire n24207;
    wire n24210;
    wire n24213;
    wire n24216;
    wire n24219;
    wire n24222;
    wire n24225;
    wire n24228;
    wire n24231;
    wire n24234;
    wire n24237;
    wire n24240;
    wire n24246;
    wire n24249;
    wire n24252;
    wire n24255;
    wire n24258;
    wire n24261;
    wire n24264;
    wire n24267;
    wire n24270;
    wire n24273;
    wire n24276;
    wire n24279;
    wire n24282;
    wire n24285;
    wire n24288;
    wire n24291;
    wire n24294;
    wire n24297;
    wire n24303;
    wire n24306;
    wire n24309;
    wire n24312;
    wire n24315;
    wire n24318;
    wire n24321;
    wire n24324;
    wire n24327;
    wire n24330;
    wire n24333;
    wire n24336;
    wire n24339;
    wire n24342;
    wire n24345;
    wire n24348;
    wire n24354;
    wire n24357;
    wire n24360;
    wire n24363;
    wire n24366;
    wire n24369;
    wire n24372;
    wire n24375;
    wire n24378;
    wire n24381;
    wire n24384;
    wire n24387;
    wire n24390;
    wire n24393;
    wire n24396;
    wire n24399;
    wire n24402;
    wire n24408;
    wire n24411;
    wire n24414;
    wire n24417;
    wire n24420;
    wire n24423;
    wire n24426;
    wire n24429;
    wire n24432;
    wire n24435;
    wire n24438;
    wire n24441;
    wire n24444;
    wire n24447;
    wire n24450;
    wire n24453;
    wire n24456;
    wire n24462;
    wire n24465;
    wire n24468;
    wire n24471;
    wire n24474;
    wire n24477;
    wire n24480;
    wire n24483;
    wire n24486;
    wire n24489;
    wire n24492;
    wire n24495;
    wire n24498;
    wire n24501;
    wire n24504;
    wire n24507;
    wire n24513;
    wire n24516;
    wire n24519;
    wire n24522;
    wire n24525;
    wire n24528;
    wire n24531;
    wire n24534;
    wire n24537;
    wire n24540;
    wire n24543;
    wire n24546;
    wire n24549;
    wire n24552;
    wire n24555;
    wire n24558;
    wire n24561;
    wire n24564;
    wire n24567;
    wire n24570;
    wire n24573;
    wire n24576;
    wire n24582;
    wire n24585;
    wire n24588;
    wire n24591;
    wire n24594;
    wire n24597;
    wire n24600;
    wire n24603;
    wire n24606;
    wire n24609;
    wire n24612;
    wire n24615;
    wire n24618;
    wire n24621;
    wire n24624;
    wire n24627;
    wire n24630;
    wire n24633;
    wire n24636;
    wire n24639;
    wire n24642;
    wire n24645;
    wire n24651;
    wire n24654;
    wire n24657;
    wire n24660;
    wire n24663;
    wire n24666;
    wire n24669;
    wire n24672;
    wire n24675;
    wire n24678;
    wire n24681;
    wire n24684;
    wire n24687;
    wire n24693;
    wire n24696;
    wire n24699;
    wire n24702;
    wire n24705;
    wire n24708;
    wire n24711;
    wire n24714;
    wire n24717;
    wire n24720;
    wire n24723;
    wire n24726;
    wire n24729;
    wire n24732;
    wire n24738;
    wire n24741;
    wire n24744;
    wire n24747;
    wire n24750;
    wire n24753;
    wire n24756;
    wire n24759;
    wire n24762;
    wire n24765;
    wire n24768;
    wire n24771;
    wire n24774;
    wire n24780;
    wire n24783;
    wire n24786;
    wire n24789;
    wire n24792;
    wire n24795;
    wire n24798;
    wire n24801;
    wire n24804;
    wire n24807;
    wire n24810;
    wire n24813;
    wire n24816;
    wire n24819;
    wire n24825;
    wire n24828;
    wire n24831;
    wire n24834;
    wire n24837;
    wire n24840;
    wire n24843;
    wire n24846;
    wire n24849;
    wire n24852;
    wire n24855;
    wire n24858;
    wire n24861;
    wire n24864;
    wire n24867;
    wire n24870;
    wire n24873;
    wire n24876;
    wire n24879;
    wire n24885;
    wire n24888;
    wire n24891;
    wire n24894;
    wire n24897;
    wire n24900;
    wire n24903;
    wire n24906;
    wire n24909;
    wire n24912;
    wire n24915;
    wire n24918;
    wire n24921;
    wire n24924;
    wire n24930;
    wire n24933;
    wire n24936;
    wire n24939;
    wire n24942;
    wire n24945;
    wire n24948;
    wire n24951;
    wire n24954;
    wire n24957;
    wire n24960;
    wire n24963;
    wire n24966;
    wire n24969;
    wire n24972;
    wire n24975;
    wire n24978;
    wire n24984;
    wire n24987;
    wire n24990;
    wire n24993;
    wire n24996;
    wire n24999;
    wire n25002;
    wire n25005;
    wire n25008;
    wire n25014;
    wire n25017;
    wire n25020;
    wire n25023;
    wire n25026;
    wire n25029;
    wire n25032;
    wire n25035;
    wire n25038;
    wire n25041;
    wire n25044;
    wire n25047;
    wire n25050;
    wire n25056;
    wire n25059;
    wire n25062;
    wire n25065;
    wire n25068;
    wire n25071;
    wire n25074;
    wire n25077;
    wire n25080;
    wire n25083;
    wire n25086;
    wire n25089;
    wire n25095;
    wire n25098;
    wire n25101;
    wire n25104;
    wire n25107;
    wire n25110;
    wire n25113;
    wire n25116;
    wire n25119;
    wire n25122;
    wire n25125;
    wire n25128;
    wire n25131;
    wire n25137;
    wire n25140;
    wire n25143;
    wire n25146;
    wire n25149;
    wire n25152;
    wire n25155;
    wire n25158;
    wire n25161;
    wire n25164;
    wire n25167;
    wire n25170;
    wire n25173;
    wire n25176;
    wire n25179;
    wire n25185;
    wire n25188;
    wire n25191;
    wire n25194;
    wire n25197;
    wire n25200;
    wire n25203;
    wire n25206;
    wire n25209;
    wire n25212;
    wire n25215;
    wire n25218;
    wire n25221;
    wire n25227;
    wire n25230;
    wire n25233;
    wire n25236;
    wire n25239;
    wire n25242;
    wire n25245;
    wire n25248;
    wire n25251;
    wire n25254;
    wire n25257;
    wire n25260;
    wire n25266;
    wire n25269;
    wire n25272;
    wire n25275;
    wire n25278;
    wire n25281;
    wire n25284;
    wire n25287;
    wire n25290;
    wire n25293;
    wire n25296;
    wire n25299;
    wire n25302;
    wire n25305;
    wire n25311;
    wire n25314;
    wire n25317;
    wire n25320;
    wire n25323;
    wire n25326;
    wire n25329;
    wire n25332;
    wire n25335;
    wire n25338;
    wire n25341;
    wire n25344;
    wire n25347;
    wire n25350;
    wire n25353;
    wire n25359;
    wire n25362;
    wire n25365;
    wire n25368;
    wire n25371;
    wire n25374;
    wire n25377;
    wire n25380;
    wire n25383;
    wire n25386;
    wire n25389;
    wire n25392;
    wire n25395;
    wire n25398;
    wire n25401;
    wire n25404;
    wire n25410;
    wire n25413;
    wire n25416;
    wire n25419;
    wire n25422;
    wire n25425;
    wire n25428;
    wire n25431;
    wire n25434;
    wire n25437;
    wire n25440;
    wire n25443;
    wire n25446;
    wire n25449;
    wire n25452;
    wire n25455;
    wire n25458;
    wire n25461;
    wire n25464;
    wire n25470;
    wire n25473;
    wire n25476;
    wire n25479;
    wire n25482;
    wire n25485;
    wire n25488;
    wire n25491;
    wire n25494;
    wire n25497;
    wire n25500;
    wire n25503;
    wire n25506;
    wire n25509;
    wire n25512;
    wire n25515;
    wire n25518;
    wire n25521;
    wire n25527;
    wire n25530;
    wire n25533;
    wire n25536;
    wire n25539;
    wire n25542;
    wire n25545;
    wire n25551;
    wire n25554;
    wire n25557;
    wire n25560;
    wire n25563;
    wire n25566;
    wire n25572;
    wire n25575;
    wire n25578;
    wire n25581;
    wire n25584;
    wire n25587;
    wire n25590;
    wire n25593;
    wire n25596;
    wire n25599;
    wire n25602;
    wire n25608;
    wire n25611;
    wire n25614;
    wire n25617;
    wire n25620;
    wire n25623;
    wire n25626;
    wire n25629;
    wire n25632;
    wire n25635;
    wire n25638;
    wire n25644;
    wire n25647;
    wire n25650;
    wire n25653;
    wire n25656;
    wire n25659;
    wire n25662;
    wire n25668;
    wire n25671;
    wire n25674;
    wire n25677;
    wire n25680;
    wire n25683;
    wire n25686;
    wire n25689;
    wire n25695;
    wire n25698;
    wire n25701;
    wire n25704;
    wire n25707;
    wire n25710;
    wire n25713;
    wire n25716;
    wire n25719;
    wire n25722;
    wire n25728;
    wire n25731;
    wire n25734;
    wire n25737;
    wire n25740;
    wire n25743;
    wire n25746;
    wire n25749;
    wire n25752;
    wire n25758;
    wire n25761;
    wire n25764;
    wire n25767;
    wire n25770;
    wire n25773;
    wire n25776;
    wire n25782;
    wire n25785;
    wire n25788;
    wire n25791;
    wire n25794;
    wire n25797;
    wire n25800;
    wire n25803;
    wire n25809;
    wire n25812;
    wire n25815;
    wire n25818;
    wire n25821;
    wire n25824;
    wire n25827;
    wire n25830;
    wire n25833;
    wire n25836;
    wire n25842;
    wire n25845;
    wire n25848;
    wire n25851;
    wire n25854;
    wire n25857;
    wire n25860;
    wire n25863;
    wire n25866;
    wire n25872;
    wire n25875;
    wire n25878;
    wire n25881;
    wire n25884;
    wire n25887;
    wire n25893;
    wire n25896;
    wire n25899;
    wire n25902;
    wire n25905;
    wire n25908;
    wire n25911;
    wire n25914;
    wire n25917;
    wire n25923;
    wire n25926;
    wire n25929;
    wire n25932;
    wire n25935;
    wire n25938;
    wire n25941;
    wire n25944;
    wire n25947;
    wire n25953;
    wire n25956;
    wire n25959;
    wire n25962;
    wire n25965;
    wire n25968;
    wire n25971;
    wire n25974;
    wire n25980;
    wire n25983;
    wire n25986;
    wire n25989;
    wire n25992;
    wire n25998;
    wire n26001;
    wire n26004;
    wire n26007;
    wire n26010;
    wire n26013;
    wire n26016;
    wire n26019;
    wire n26022;
    wire n26028;
    wire n26031;
    wire n26034;
    wire n26037;
    wire n26040;
    wire n26043;
    wire n26046;
    wire n26049;
    wire n26052;
    wire n26058;
    wire n26061;
    wire n26064;
    wire n26067;
    wire n26070;
    wire n26073;
    wire n26076;
    wire n26079;
    wire n26085;
    wire n26088;
    wire n26091;
    wire n26094;
    wire n26097;
    wire n26100;
    wire n26106;
    wire n26109;
    wire n26112;
    wire n26115;
    wire n26118;
    wire n26121;
    wire n26124;
    wire n26127;
    wire n26130;
    wire n26136;
    wire n26139;
    wire n26142;
    wire n26145;
    wire n26148;
    wire n26151;
    wire n26157;
    wire n26160;
    wire n26163;
    wire n26166;
    wire n26169;
    wire n26172;
    wire n26175;
    wire n26181;
    wire n26184;
    wire n26187;
    wire n26190;
    wire n26193;
    wire n26196;
    wire n26202;
    wire n26205;
    wire n26208;
    wire n26211;
    wire n26214;
    wire n26217;
    wire n26220;
    wire n26223;
    wire n26226;
    wire n26229;
    wire n26232;
    wire n26238;
    wire n26241;
    wire n26244;
    wire n26247;
    wire n26250;
    wire n26253;
    wire n26256;
    wire n26259;
    wire n26262;
    wire n26265;
    wire n26268;
    wire n26271;
    wire n26274;
    wire n26277;
    wire n26280;
    wire n26283;
    wire n26289;
    wire n26292;
    wire n26295;
    wire n26298;
    wire n26301;
    wire n26307;
    wire n26310;
    wire n26313;
    wire n26316;
    wire n26319;
    wire n26322;
    wire n26325;
    wire n26328;
    wire n26334;
    wire n26337;
    wire n26340;
    wire n26343;
    wire n26346;
    wire n26349;
    wire n26355;
    wire n26358;
    wire n26361;
    wire n26364;
    wire n26367;
    wire n26370;
    wire n26373;
    wire n26376;
    wire n26379;
    wire n26385;
    wire n26388;
    wire n26391;
    wire n26397;
    wire n26400;
    wire n26406;
    wire n26409;
    wire n26412;
    wire n26418;
    wire n26421;
    wire n26424;
    wire n26430;
    wire n26433;
    wire n26436;
    wire n26439;
    wire n26445;
    wire n26448;
    wire n26451;
    wire n26457;
    wire n26460;
    wire n26463;
    wire n26469;
    wire n26472;
    wire n26475;
    wire n26478;
    wire n26484;
    wire n26487;
    wire n26490;
    wire n26496;
    wire n26499;
    wire n26505;
    wire n26508;
    wire n26514;
    wire n26520;
    wire n26523;
    wire n26526;
    wire n26532;
    wire n26535;
    wire n26541;
    wire n26544;
    wire n26550;
    wire n26553;
    wire n26559;
    wire n26562;
    wire n26565;
    wire n26568;
    wire n26571;
    wire n26577;
    wire n26580;
    wire n26583;
    wire n26586;
    wire n26589;
    jnot g0000(.din(G545), .dout(n303));
    jnot g0001(.din(G348), .dout(n306));
    jnot g0002(.din(G366), .dout(n309));
    jand g0003(.dinb(G552), .dina(G562), .dout(n313));
    jnot g0004(.din(G549), .dout(n316));
    jnot g0005(.din(G338), .dout(n319));
    jnot g0006(.din(G358), .dout(n322));
    jand g0007(.dinb(G141), .dina(G145), .dout(n326));
    jnot g0008(.din(G245), .dout(n329));
    jnot g0009(.din(G552), .dout(n332));
    jnot g0010(.din(G562), .dout(n335));
    jnot g0011(.din(G559), .dout(n338));
    jand g0012(.dinb(G1), .dina(G373), .dout(n342));
    jnot g0013(.din(G3173), .dout(n345));
    jand g0014(.dinb(n8401), .dina(n345), .dout(n349));
    jnot g0015(.din(G27), .dout(n352));
    jor g0016(.dinb(n352), .dina(n8404), .dout(n356));
    jand g0017(.dinb(G386), .dina(G556), .dout(n360));
    jnot g0018(.din(n360), .dout(n363));
    jnot g0019(.din(G140), .dout(n366));
    jnot g0020(.din(G31), .dout(n369));
    jor g0021(.dinb(n352), .dina(n369), .dout(n373));
    jor g0022(.dinb(n8407), .dina(n373), .dout(n377));
    jnot g0023(.din(G299), .dout(n380));
    jnot g0024(.din(G86), .dout(n383));
    jnot g0025(.din(G2358), .dout(n386));
    jand g0026(.dinb(n383), .dina(n386), .dout(n390));
    jnot g0027(.din(G87), .dout(n393));
    jand g0028(.dinb(n393), .dina(n8481), .dout(n397));
    jor g0029(.dinb(n373), .dina(n397), .dout(n401));
    jor g0030(.dinb(n8410), .dina(n401), .dout(n405));
    jnot g0031(.din(G88), .dout(n408));
    jand g0032(.dinb(n408), .dina(n386), .dout(n412));
    jnot g0033(.din(G34), .dout(n415));
    jand g0034(.dinb(n415), .dina(n8478), .dout(n419));
    jor g0035(.dinb(n373), .dina(n419), .dout(n423));
    jor g0036(.dinb(n8413), .dina(n423), .dout(n427));
    jnot g0037(.din(G83), .dout(n430));
    jor g0038(.dinb(n8416), .dina(n373), .dout(n434));
    jand g0039(.dinb(n8425), .dina(n386), .dout(n438));
    jand g0040(.dinb(G25), .dina(G2358), .dout(n442));
    jor g0041(.dinb(n373), .dina(n8422), .dout(n446));
    jor g0042(.dinb(n8419), .dina(n446), .dout(n450));
    jand g0043(.dinb(n8448), .dina(n450), .dout(n454));
    jand g0044(.dinb(n8434), .dina(n386), .dout(n458));
    jand g0045(.dinb(G81), .dina(G2358), .dout(n462));
    jor g0046(.dinb(n373), .dina(n8431), .dout(n466));
    jor g0047(.dinb(n8428), .dina(n466), .dout(n470));
    jand g0048(.dinb(n8436), .dina(n470), .dout(n474));
    jand g0049(.dinb(n8467), .dina(n386), .dout(n478));
    jand g0050(.dinb(G23), .dina(G2358), .dout(n482));
    jor g0051(.dinb(n373), .dina(n8464), .dout(n486));
    jor g0052(.dinb(n8461), .dina(n486), .dout(n490));
    jand g0053(.dinb(n8496), .dina(n490), .dout(n494));
    jand g0054(.dinb(G80), .dina(G2358), .dout(n498));
    jand g0055(.dinb(n8476), .dina(n386), .dout(n502));
    jor g0056(.dinb(n373), .dina(n502), .dout(n506));
    jor g0057(.dinb(n8473), .dina(n506), .dout(n510));
    jand g0058(.dinb(n8484), .dina(n510), .dout(n514));
    jand g0059(.dinb(G514), .dina(G3552), .dout(n518));
    jnot g0060(.din(G514), .dout(n521));
    jnot g0061(.din(G3546), .dout(n524));
    jand g0062(.dinb(n521), .dina(n524), .dout(n528));
    jor g0063(.dinb(n11023), .dina(n528), .dout(n532));
    jnot g0064(.din(n532), .dout(n535));
    jnot g0065(.din(G251), .dout(n538));
    jnot g0066(.din(G361), .dout(n541));
    jand g0067(.dinb(n538), .dina(n541), .dout(n545));
    jnot g0068(.din(G248), .dout(n548));
    jand g0069(.dinb(n548), .dina(n17121), .dout(n552));
    jor g0070(.dinb(n545), .dina(n552), .dout(n556));
    jnot g0071(.din(n556), .dout(n559));
    jand g0072(.dinb(n535), .dina(n559), .dout(n563));
    jnot g0073(.din(G351), .dout(n566));
    jnot g0074(.din(G3550), .dout(n569));
    jand g0075(.dinb(n566), .dina(n569), .dout(n573));
    jnot g0076(.din(G534), .dout(n576));
    jnot g0077(.din(G3552), .dout(n579));
    jand g0078(.dinb(n17160), .dina(n579), .dout(n583));
    jor g0079(.dinb(n17545), .dina(n583), .dout(n587));
    jor g0080(.dinb(n10597), .dina(n587), .dout(n591));
    jand g0081(.dinb(G351), .dina(G3546), .dout(n595));
    jand g0082(.dinb(n566), .dina(n14263), .dout(n599));
    jor g0083(.dinb(n10594), .dina(n599), .dout(n603));
    jor g0084(.dinb(n17547), .dina(n603), .dout(n607));
    jand g0085(.dinb(n591), .dina(n607), .dout(n611));
    jnot g0086(.din(G341), .dout(n614));
    jand g0087(.dinb(n614), .dina(n569), .dout(n618));
    jnot g0088(.din(G523), .dout(n621));
    jand g0089(.dinb(n17151), .dina(n579), .dout(n625));
    jor g0090(.dinb(n17983), .dina(n625), .dout(n629));
    jor g0091(.dinb(n10828), .dina(n629), .dout(n633));
    jand g0092(.dinb(G341), .dina(G3546), .dout(n637));
    jand g0093(.dinb(n614), .dina(n14263), .dout(n641));
    jor g0094(.dinb(n10825), .dina(n641), .dout(n645));
    jor g0095(.dinb(n17994), .dina(n645), .dout(n649));
    jand g0096(.dinb(n633), .dina(n649), .dout(n653));
    jand g0097(.dinb(n611), .dina(n653), .dout(n657));
    jand g0098(.dinb(n8509), .dina(n657), .dout(n661));
    jand g0099(.dinb(G248), .dina(G316), .dout(n665));
    jnot g0100(.din(G490), .dout(n668));
    jnot g0101(.din(G316), .dout(n671));
    jand g0102(.dinb(n19431), .dina(n671), .dout(n675));
    jor g0103(.dinb(n17683), .dina(n675), .dout(n679));
    jor g0104(.dinb(n17113), .dina(n679), .dout(n683));
    jnot g0105(.din(G254), .dout(n686));
    jand g0106(.dinb(n686), .dina(n671), .dout(n690));
    jnot g0107(.din(G242), .dout(n693));
    jand g0108(.dinb(n693), .dina(n17784), .dout(n697));
    jor g0109(.dinb(n690), .dina(n697), .dout(n701));
    jor g0110(.dinb(n17685), .dina(n701), .dout(n705));
    jand g0111(.dinb(n683), .dina(n705), .dout(n709));
    jand g0112(.dinb(G248), .dina(G308), .dout(n713));
    jnot g0113(.din(G479), .dout(n716));
    jnot g0114(.din(G308), .dout(n719));
    jand g0115(.dinb(n19434), .dina(n719), .dout(n723));
    jor g0116(.dinb(n17836), .dina(n723), .dout(n727));
    jor g0117(.dinb(n17104), .dina(n727), .dout(n731));
    jand g0118(.dinb(n686), .dina(n719), .dout(n735));
    jand g0119(.dinb(n693), .dina(n17106), .dout(n739));
    jor g0120(.dinb(n735), .dina(n739), .dout(n743));
    jor g0121(.dinb(n17847), .dina(n743), .dout(n747));
    jand g0122(.dinb(n731), .dina(n747), .dout(n751));
    jand g0123(.dinb(n709), .dina(n751), .dout(n755));
    jnot g0124(.din(G293), .dout(n758));
    jand g0125(.dinb(n686), .dina(n758), .dout(n762));
    jand g0126(.dinb(n693), .dina(n17736), .dout(n766));
    jor g0127(.dinb(n762), .dina(n766), .dout(n770));
    jnot g0128(.din(G302), .dout(n773));
    jand g0129(.dinb(n538), .dina(n773), .dout(n777));
    jand g0130(.dinb(n548), .dina(n17892), .dout(n781));
    jor g0131(.dinb(n777), .dina(n781), .dout(n785));
    jnot g0132(.din(n785), .dout(n788));
    jand g0133(.dinb(n11328), .dina(n788), .dout(n792));
    jnot g0134(.din(G324), .dout(n795));
    jand g0135(.dinb(n795), .dina(n569), .dout(n799));
    jnot g0136(.din(G503), .dout(n802));
    jand g0137(.dinb(n18099), .dina(n579), .dout(n806));
    jor g0138(.dinb(n17131), .dina(n806), .dout(n810));
    jor g0139(.dinb(n10348), .dina(n810), .dout(n814));
    jand g0140(.dinb(G324), .dina(G3546), .dout(n818));
    jand g0141(.dinb(n795), .dina(n14263), .dout(n822));
    jor g0142(.dinb(n10345), .dina(n822), .dout(n826));
    jor g0143(.dinb(n17133), .dina(n826), .dout(n830));
    jand g0144(.dinb(n814), .dina(n830), .dout(n834));
    jand g0145(.dinb(n792), .dina(n834), .dout(n838));
    jand g0146(.dinb(n755), .dina(n838), .dout(n842));
    jand g0147(.dinb(n661), .dina(n842), .dout(n846));
    jnot g0148(.din(G210), .dout(n849));
    jand g0149(.dinb(n849), .dina(n569), .dout(n853));
    jnot g0150(.din(G457), .dout(n856));
    jand g0151(.dinb(n19035), .dina(n579), .dout(n860));
    jor g0152(.dinb(n19045), .dina(n860), .dout(n864));
    jor g0153(.dinb(n14266), .dina(n864), .dout(n868));
    jand g0154(.dinb(G210), .dina(G3546), .dout(n872));
    jand g0155(.dinb(n849), .dina(n14263), .dout(n876));
    jor g0156(.dinb(n14260), .dina(n876), .dout(n880));
    jor g0157(.dinb(n19059), .dina(n880), .dout(n884));
    jand g0158(.dinb(n868), .dina(n884), .dout(n888));
    jnot g0159(.din(G234), .dout(n891));
    jand g0160(.dinb(n891), .dina(n569), .dout(n895));
    jnot g0161(.din(G435), .dout(n898));
    jand g0162(.dinb(n19269), .dina(n579), .dout(n902));
    jor g0163(.dinb(n19282), .dina(n902), .dout(n906));
    jor g0164(.dinb(n10423), .dina(n906), .dout(n910));
    jand g0165(.dinb(G234), .dina(G3546), .dout(n914));
    jand g0166(.dinb(n891), .dina(n14263), .dout(n918));
    jor g0167(.dinb(n10420), .dina(n918), .dout(n922));
    jor g0168(.dinb(n19296), .dina(n922), .dout(n926));
    jand g0169(.dinb(n910), .dina(n926), .dout(n930));
    jnot g0170(.din(G273), .dout(n933));
    jand g0171(.dinb(n933), .dina(n569), .dout(n937));
    jnot g0172(.din(G411), .dout(n940));
    jand g0173(.dinb(n19548), .dina(n579), .dout(n944));
    jor g0174(.dinb(n19570), .dina(n944), .dout(n948));
    jor g0175(.dinb(n10519), .dina(n948), .dout(n952));
    jand g0176(.dinb(G273), .dina(G3546), .dout(n956));
    jand g0177(.dinb(n933), .dina(n14263), .dout(n960));
    jor g0178(.dinb(n10516), .dina(n960), .dout(n964));
    jor g0179(.dinb(n19572), .dina(n964), .dout(n968));
    jand g0180(.dinb(n952), .dina(n968), .dout(n972));
    jand g0181(.dinb(n930), .dina(n972), .dout(n976));
    jnot g0182(.din(G265), .dout(n979));
    jand g0183(.dinb(n979), .dina(n569), .dout(n983));
    jnot g0184(.din(G400), .dout(n986));
    jand g0185(.dinb(n19458), .dina(n579), .dout(n990));
    jor g0186(.dinb(n19405), .dina(n990), .dout(n994));
    jor g0187(.dinb(n10768), .dina(n994), .dout(n998));
    jand g0188(.dinb(G265), .dina(G3546), .dout(n1002));
    jand g0189(.dinb(n979), .dina(n14263), .dout(n1006));
    jor g0190(.dinb(n10765), .dina(n1006), .dout(n1010));
    jor g0191(.dinb(n19419), .dina(n1010), .dout(n1014));
    jand g0192(.dinb(n998), .dina(n1014), .dout(n1018));
    jnot g0193(.din(G226), .dout(n1021));
    jand g0194(.dinb(n1021), .dina(n569), .dout(n1025));
    jnot g0195(.din(G422), .dout(n1028));
    jand g0196(.dinb(n19161), .dina(n579), .dout(n1032));
    jor g0197(.dinb(n19174), .dina(n1032), .dout(n1036));
    jor g0198(.dinb(n13645), .dina(n1036), .dout(n1040));
    jand g0199(.dinb(G226), .dina(G3546), .dout(n1044));
    jand g0200(.dinb(n1021), .dina(n14263), .dout(n1048));
    jor g0201(.dinb(n13642), .dina(n1048), .dout(n1052));
    jor g0202(.dinb(n19176), .dina(n1052), .dout(n1056));
    jand g0203(.dinb(n1040), .dina(n1056), .dout(n1060));
    jand g0204(.dinb(n1018), .dina(n1060), .dout(n1064));
    jand g0205(.dinb(n976), .dina(n1064), .dout(n1068));
    jnot g0206(.din(G218), .dout(n1071));
    jand g0207(.dinb(n1071), .dina(n569), .dout(n1075));
    jnot g0208(.din(G468), .dout(n1078));
    jand g0209(.dinb(n19152), .dina(n579), .dout(n1082));
    jor g0210(.dinb(n19105), .dina(n1082), .dout(n1086));
    jor g0211(.dinb(n13954), .dina(n1086), .dout(n1090));
    jand g0212(.dinb(G218), .dina(G3546), .dout(n1094));
    jand g0213(.dinb(n1071), .dina(n14263), .dout(n1098));
    jor g0214(.dinb(n13951), .dina(n1098), .dout(n1102));
    jor g0215(.dinb(n19119), .dina(n1102), .dout(n1106));
    jand g0216(.dinb(n1090), .dina(n1106), .dout(n1110));
    jnot g0217(.din(G257), .dout(n1113));
    jand g0218(.dinb(n1113), .dina(n569), .dout(n1117));
    jnot g0219(.din(G389), .dout(n1120));
    jand g0220(.dinb(n19335), .dina(n579), .dout(n1124));
    jor g0221(.dinb(n19345), .dina(n1124), .dout(n1128));
    jor g0222(.dinb(n10927), .dina(n1128), .dout(n1132));
    jand g0223(.dinb(G257), .dina(G3546), .dout(n1136));
    jand g0224(.dinb(n1113), .dina(n14263), .dout(n1140));
    jor g0225(.dinb(n10924), .dina(n1140), .dout(n1144));
    jor g0226(.dinb(n19359), .dina(n1144), .dout(n1148));
    jand g0227(.dinb(n1132), .dina(n1148), .dout(n1152));
    jand g0228(.dinb(n1110), .dina(n1152), .dout(n1156));
    jnot g0229(.din(G281), .dout(n1159));
    jand g0230(.dinb(n1159), .dina(n569), .dout(n1163));
    jnot g0231(.din(G374), .dout(n1166));
    jand g0232(.dinb(n19470), .dina(n579), .dout(n1170));
    jor g0233(.dinb(n19486), .dina(n1170), .dout(n1174));
    jor g0234(.dinb(n8899), .dina(n1174), .dout(n1178));
    jand g0235(.dinb(G281), .dina(G3546), .dout(n1182));
    jand g0236(.dinb(n1159), .dina(n14263), .dout(n1186));
    jor g0237(.dinb(n8896), .dina(n1186), .dout(n1190));
    jor g0238(.dinb(n19500), .dina(n1190), .dout(n1194));
    jand g0239(.dinb(n1178), .dina(n1194), .dout(n1198));
    jand g0240(.dinb(G206), .dina(G248), .dout(n1202));
    jnot g0241(.din(G446), .dout(n1205));
    jnot g0242(.din(G206), .dout(n1208));
    jand g0243(.dinb(n1208), .dina(n19434), .dout(n1212));
    jor g0244(.dinb(n19216), .dina(n1212), .dout(n1216));
    jor g0245(.dinb(n19213), .dina(n1216), .dout(n1220));
    jand g0246(.dinb(n1208), .dina(n686), .dout(n1224));
    jand g0247(.dinb(n19254), .dina(n693), .dout(n1228));
    jor g0248(.dinb(n1224), .dina(n1228), .dout(n1232));
    jor g0249(.dinb(n19227), .dina(n1232), .dout(n1236));
    jand g0250(.dinb(n1220), .dina(n1236), .dout(n1240));
    jand g0251(.dinb(n1198), .dina(n1240), .dout(n1244));
    jand g0252(.dinb(n1156), .dina(n1244), .dout(n1248));
    jand g0253(.dinb(n1068), .dina(n1248), .dout(n1252));
    jand g0254(.dinb(n14250), .dina(n1252), .dout(n1256));
    jnot g0255(.din(G335), .dout(n1259));
    jand g0256(.dinb(n1159), .dina(n1259), .dout(n1263));
    jnot g0257(.din(n1263), .dout(n1266));
    jor g0258(.dinb(n19000), .dina(n1259), .dout(n1270));
    jand g0259(.dinb(n1266), .dina(n18996), .dout(n1274));
    jxor g0260(.dinb(n19488), .dina(n1274), .dout(n1278));
    jand g0261(.dinb(n933), .dina(n1259), .dout(n1282));
    jnot g0262(.din(n1282), .dout(n1285));
    jor g0263(.dinb(n18988), .dina(n1259), .dout(n1289));
    jand g0264(.dinb(n1285), .dina(n18984), .dout(n1293));
    jxor g0265(.dinb(n19581), .dina(n1293), .dout(n1297));
    jand g0266(.dinb(n1278), .dina(n1297), .dout(n1301));
    jnot g0267(.din(n1301), .dout(n1304));
    jand g0268(.dinb(n979), .dina(n1259), .dout(n1308));
    jnot g0269(.din(n1308), .dout(n1311));
    jor g0270(.dinb(n19015), .dina(n1259), .dout(n1315));
    jand g0271(.dinb(n1311), .dina(n19011), .dout(n1319));
    jxor g0272(.dinb(n19407), .dina(n1319), .dout(n1323));
    jnot g0273(.din(n1323), .dout(n1326));
    jand g0274(.dinb(n1113), .dina(n1259), .dout(n1330));
    jnot g0275(.din(n1330), .dout(n1333));
    jor g0276(.dinb(n18943), .dina(n1259), .dout(n1337));
    jand g0277(.dinb(n1333), .dina(n18940), .dout(n1341));
    jxor g0278(.dinb(n19338), .dina(n1341), .dout(n1345));
    jor g0279(.dinb(n1326), .dina(n18921), .dout(n1349));
    jor g0280(.dinb(n1304), .dina(n1349), .dout(n1353));
    jnot g0281(.din(n1353), .dout(n1356));
    jand g0282(.dinb(n891), .dina(n1259), .dout(n1360));
    jnot g0283(.din(n1360), .dout(n1363));
    jor g0284(.dinb(n18877), .dina(n1259), .dout(n1367));
    jand g0285(.dinb(n1363), .dina(n18874), .dout(n1371));
    jxor g0286(.dinb(n19284), .dina(n1371), .dout(n1375));
    jand g0287(.dinb(n1356), .dina(n18861), .dout(n1379));
    jor g0288(.dinb(G206), .dina(G335), .dout(n1383));
    jor g0289(.dinb(n18529), .dina(n1259), .dout(n1387));
    jand g0290(.dinb(n18526), .dina(n1387), .dout(n1391));
    jxor g0291(.dinb(n19218), .dina(n1391), .dout(n1395));
    jand g0292(.dinb(n1021), .dina(n1259), .dout(n1399));
    jnot g0293(.din(n1399), .dout(n1402));
    jor g0294(.dinb(n18577), .dina(n1259), .dout(n1406));
    jand g0295(.dinb(n1402), .dina(n18574), .dout(n1410));
    jxor g0296(.dinb(n18453), .dina(n1410), .dout(n1414));
    jand g0297(.dinb(n1071), .dina(n1259), .dout(n1418));
    jnot g0298(.din(n1418), .dout(n1421));
    jor g0299(.dinb(n18571), .dina(n1259), .dout(n1425));
    jand g0300(.dinb(n1421), .dina(n18568), .dout(n1429));
    jxor g0301(.dinb(n19098), .dina(n1429), .dout(n1433));
    jor g0302(.dinb(n1414), .dina(n1433), .dout(n1437));
    jand g0303(.dinb(n849), .dina(n1259), .dout(n1441));
    jnot g0304(.din(n1441), .dout(n1444));
    jor g0305(.dinb(n18508), .dina(n1259), .dout(n1448));
    jand g0306(.dinb(n1444), .dina(n18505), .dout(n1452));
    jxor g0307(.dinb(n19038), .dina(n1452), .dout(n1456));
    jor g0308(.dinb(n1437), .dina(n18501), .dout(n1460));
    jnot g0309(.din(n1460), .dout(n1463));
    jand g0310(.dinb(n18513), .dina(n1463), .dout(n1467));
    jand g0311(.dinb(n1379), .dina(n8563), .dout(n1471));
    jnot g0312(.din(G332), .dout(n1474));
    jand g0313(.dinb(n795), .dina(n1474), .dout(n1478));
    jnot g0314(.din(n1478), .dout(n1481));
    jor g0315(.dinb(n18096), .dina(n1474), .dout(n1485));
    jand g0316(.dinb(n1481), .dina(n18094), .dout(n1489));
    jxor g0317(.dinb(n18105), .dina(n1489), .dout(n1493));
    jor g0318(.dinb(n1474), .dina(n18054), .dout(n1497));
    jxor g0319(.dinb(n18057), .dina(n1497), .dout(n1501));
    jor g0320(.dinb(G332), .dina(G341), .dout(n1505));
    jor g0321(.dinb(n1474), .dina(n17964), .dout(n1509));
    jand g0322(.dinb(n17970), .dina(n1509), .dout(n1513));
    jxor g0323(.dinb(n17985), .dina(n1513), .dout(n1517));
    jor g0324(.dinb(G332), .dina(G351), .dout(n1521));
    jor g0325(.dinb(n1474), .dina(n17931), .dout(n1525));
    jand g0326(.dinb(n17934), .dina(n1525), .dout(n1529));
    jor g0327(.dinb(n17940), .dina(n1529), .dout(n1533));
    jnot g0328(.din(n1521), .dout(n1536));
    jand g0329(.dinb(n17916), .dina(n322), .dout(n1540));
    jor g0330(.dinb(n1536), .dina(n1540), .dout(n1544));
    jor g0331(.dinb(n17523), .dina(n1544), .dout(n1548));
    jor g0332(.dinb(G332), .dina(G361), .dout(n1552));
    jor g0333(.dinb(n1474), .dina(n17910), .dout(n1556));
    jand g0334(.dinb(n17908), .dina(n1556), .dout(n1560));
    jnot g0335(.din(n1560), .dout(n1563));
    jand g0336(.dinb(n1548), .dina(n1563), .dout(n1567));
    jand g0337(.dinb(n17928), .dina(n1567), .dout(n1571));
    jand g0338(.dinb(n17305), .dina(n1571), .dout(n1575));
    jand g0339(.dinb(n17307), .dina(n1575), .dout(n1579));
    jand g0340(.dinb(n17364), .dina(n1579), .dout(n1583));
    jand g0341(.dinb(n758), .dina(n1474), .dout(n1587));
    jand g0342(.dinb(n380), .dina(n17913), .dout(n1591));
    jor g0343(.dinb(n1587), .dina(n1591), .dout(n1595));
    jand g0344(.dinb(n773), .dina(n1474), .dout(n1599));
    jnot g0345(.din(n1599), .dout(n1602));
    jor g0346(.dinb(n17887), .dina(n1474), .dout(n1606));
    jand g0347(.dinb(n1602), .dina(n17884), .dout(n1610));
    jnot g0348(.din(n1610), .dout(n1613));
    jand g0349(.dinb(n17730), .dina(n1613), .dout(n1617));
    jor g0350(.dinb(G308), .dina(G332), .dout(n1621));
    jor g0351(.dinb(n17827), .dina(n1474), .dout(n1625));
    jand g0352(.dinb(n17824), .dina(n1625), .dout(n1629));
    jxor g0353(.dinb(n17838), .dina(n1629), .dout(n1633));
    jand g0354(.dinb(n671), .dina(n1474), .dout(n1637));
    jnot g0355(.din(n1637), .dout(n1640));
    jor g0356(.dinb(n17782), .dina(n1474), .dout(n1644));
    jand g0357(.dinb(n1640), .dina(n17779), .dout(n1648));
    jxor g0358(.dinb(n17799), .dina(n1648), .dout(n1652));
    jand g0359(.dinb(n17818), .dina(n1652), .dout(n1656));
    jand g0360(.dinb(n1617), .dina(n1656), .dout(n1660));
    jand g0361(.dinb(n1583), .dina(n8515), .dout(n1664));
    jxor g0362(.dinb(G308), .dina(G316), .dout(n1668));
    jxor g0363(.dinb(n758), .dina(n17889), .dout(n1672));
    jxor g0364(.dinb(n11416), .dina(n1672), .dout(n1676));
    jxor g0365(.dinb(G361), .dina(G369), .dout(n1680));
    jxor g0366(.dinb(n795), .dina(n1680), .dout(n1684));
    jxor g0367(.dinb(G341), .dina(G351), .dout(n1688));
    jxor g0368(.dinb(n1684), .dina(n11413), .dout(n1692));
    jxor g0369(.dinb(n1676), .dina(n1692), .dout(n1696));
    jnot g0370(.din(n1696), .dout(n1699));
    jxor g0371(.dinb(G218), .dina(G226), .dout(n1703));
    jxor g0372(.dinb(n979), .dina(n19602), .dout(n1707));
    jxor g0373(.dinb(n11455), .dina(n1707), .dout(n1711));
    jxor g0374(.dinb(G281), .dina(G289), .dout(n1715));
    jxor g0375(.dinb(G234), .dina(G257), .dout(n1719));
    jxor g0376(.dinb(n1715), .dina(n1719), .dout(n1723));
    jxor g0377(.dinb(G206), .dina(G210), .dout(n1727));
    jxor g0378(.dinb(n1723), .dina(n11452), .dout(n1731));
    jxor g0379(.dinb(n1711), .dina(n1731), .dout(n1735));
    jnot g0380(.din(n1735), .dout(n1738));
    jand g0381(.dinb(n19314), .dina(n1371), .dout(n1742));
    jnot g0382(.din(n1371), .dout(n1745));
    jand g0383(.dinb(n19272), .dina(n1745), .dout(n1749));
    jnot g0384(.din(n1749), .dout(n1752));
    jand g0385(.dinb(n19347), .dina(n1341), .dout(n1756));
    jor g0386(.dinb(n19377), .dina(n1341), .dout(n1760));
    jnot g0387(.din(n1315), .dout(n1763));
    jor g0388(.dinb(n19017), .dina(n1763), .dout(n1767));
    jand g0389(.dinb(n19020), .dina(n1767), .dout(n1771));
    jnot g0390(.din(n1771), .dout(n1774));
    jand g0391(.dinb(n19518), .dina(n1274), .dout(n1778));
    jor g0392(.dinb(n19581), .dina(n1293), .dout(n1782));
    jand g0393(.dinb(n1778), .dina(n1782), .dout(n1786));
    jand g0394(.dinb(n19581), .dina(n1293), .dout(n1790));
    jand g0395(.dinb(n19446), .dina(n1319), .dout(n1794));
    jor g0396(.dinb(n1790), .dina(n1794), .dout(n1798));
    jor g0397(.dinb(n1786), .dina(n1798), .dout(n1802));
    jand g0398(.dinb(n18976), .dina(n1802), .dout(n1806));
    jand g0399(.dinb(n18894), .dina(n1806), .dout(n1810));
    jor g0400(.dinb(n18903), .dina(n1810), .dout(n1814));
    jand g0401(.dinb(n18595), .dina(n1814), .dout(n1818));
    jor g0402(.dinb(n18627), .dina(n1818), .dout(n1822));
    jand g0403(.dinb(n8556), .dina(n1822), .dout(n1826));
    jand g0404(.dinb(n19245), .dina(n1391), .dout(n1830));
    jor g0405(.dinb(n19236), .dina(n1391), .dout(n1834));
    jand g0406(.dinb(n19047), .dina(n1452), .dout(n1838));
    jor g0407(.dinb(n19077), .dina(n1452), .dout(n1842));
    jand g0408(.dinb(n19107), .dina(n1429), .dout(n1846));
    jand g0409(.dinb(n19194), .dina(n1410), .dout(n1850));
    jor g0410(.dinb(n19140), .dina(n1429), .dout(n1854));
    jand g0411(.dinb(n1850), .dina(n1854), .dout(n1858));
    jor g0412(.dinb(n18564), .dina(n1858), .dout(n1862));
    jand g0413(.dinb(n18391), .dina(n1862), .dout(n1866));
    jor g0414(.dinb(n18385), .dina(n1866), .dout(n1870));
    jand g0415(.dinb(n8554), .dina(n1870), .dout(n1874));
    jor g0416(.dinb(n8539), .dina(n1874), .dout(n1878));
    jor g0417(.dinb(n1826), .dina(n8521), .dout(n1882));
    jand g0418(.dinb(n18105), .dina(n1489), .dout(n1886));
    jor g0419(.dinb(n18105), .dina(n1489), .dout(n1890));
    jor g0420(.dinb(n18057), .dina(n1497), .dout(n1894));
    jand g0421(.dinb(n18057), .dina(n1497), .dout(n1898));
    jnot g0422(.din(n1505), .dout(n1901));
    jand g0423(.dinb(n17967), .dina(n306), .dout(n1905));
    jor g0424(.dinb(n1901), .dina(n1905), .dout(n1909));
    jand g0425(.dinb(n17976), .dina(n1909), .dout(n1913));
    jnot g0426(.din(n1913), .dout(n1916));
    jand g0427(.dinb(n1533), .dina(n17898), .dout(n1920));
    jand g0428(.dinb(n18012), .dina(n1513), .dout(n1924));
    jand g0429(.dinb(n17940), .dina(n1529), .dout(n1928));
    jor g0430(.dinb(n1924), .dina(n1928), .dout(n1932));
    jor g0431(.dinb(n1920), .dina(n1932), .dout(n1936));
    jand g0432(.dinb(n17896), .dina(n1936), .dout(n1940));
    jor g0433(.dinb(n18021), .dina(n1940), .dout(n1944));
    jand g0434(.dinb(n18033), .dina(n1944), .dout(n1948));
    jand g0435(.dinb(n18066), .dina(n1948), .dout(n1952));
    jor g0436(.dinb(n18078), .dina(n1952), .dout(n1956));
    jand g0437(.dinb(n8577), .dina(n1956), .dout(n1960));
    jnot g0438(.din(n1617), .dout(n1963));
    jnot g0439(.din(n1629), .dout(n1966));
    jor g0440(.dinb(n17829), .dina(n1966), .dout(n1970));
    jand g0441(.dinb(n17787), .dina(n1648), .dout(n1974));
    jand g0442(.dinb(n17818), .dina(n1974), .dout(n1978));
    jnot g0443(.din(n1978), .dout(n1981));
    jand g0444(.dinb(n17755), .dina(n1981), .dout(n1985));
    jnot g0445(.din(n1985), .dout(n1988));
    jor g0446(.dinb(n8575), .dina(n1988), .dout(n1992));
    jor g0447(.dinb(n1960), .dina(n8569), .dout(n1996));
    jnot g0448(.din(G4091), .dout(n1999));
    jand g0449(.dinb(n1999), .dina(n19908), .dout(n2003));
    jand g0450(.dinb(n8959), .dina(n2003), .dout(n2007));
    jnot g0451(.din(n2007), .dout(n2010));
    jnot g0452(.din(G54), .dout(n2013));
    jxor g0453(.dinb(n11089), .dina(n1560), .dout(n2017));
    jnot g0454(.din(n2017), .dout(n2020));
    jand g0455(.dinb(n19725), .dina(n2020), .dout(n2024));
    jand g0456(.dinb(n15375), .dina(n559), .dout(n2028));
    jor g0457(.dinb(n15336), .dina(n2028), .dout(n2032));
    jor g0458(.dinb(n2024), .dina(n2032), .dout(n2036));
    jand g0459(.dinb(n8920), .dina(n2036), .dout(n2040));
    jand g0460(.dinb(n10654), .dina(n2003), .dout(n2044));
    jnot g0461(.din(n2044), .dout(n2047));
    jxor g0462(.dinb(n17940), .dina(n1529), .dout(n2051));
    jnot g0463(.din(n2051), .dout(n2054));
    jand g0464(.dinb(n17901), .dina(n2054), .dout(n2058));
    jor g0465(.dinb(n1571), .dina(n2058), .dout(n2062));
    jnot g0466(.din(n2062), .dout(n2065));
    jand g0467(.dinb(n10611), .dina(n2065), .dout(n2069));
    jand g0468(.dinb(n14772), .dina(n2051), .dout(n2073));
    jor g0469(.dinb(n2069), .dina(n10609), .dout(n2077));
    jand g0470(.dinb(n10641), .dina(n2077), .dout(n2081));
    jand g0471(.dinb(n11034), .dina(n611), .dout(n2085));
    jor g0472(.dinb(n15321), .dina(n2085), .dout(n2089));
    jor g0473(.dinb(n2081), .dina(n10591), .dout(n2093));
    jand g0474(.dinb(n10579), .dina(n2093), .dout(n2097));
    jand g0475(.dinb(n8911), .dina(n2003), .dout(n2101));
    jnot g0476(.din(n2101), .dout(n2104));
    jxor g0477(.dinb(n15055), .dina(n1278), .dout(n2108));
    jnot g0478(.din(n2108), .dout(n2111));
    jand g0479(.dinb(n19764), .dina(n2111), .dout(n2115));
    jand g0480(.dinb(n11034), .dina(n1198), .dout(n2119));
    jor g0481(.dinb(n11040), .dina(n2119), .dout(n2123));
    jor g0482(.dinb(n2115), .dina(n8893), .dout(n2127));
    jand g0483(.dinb(n8890), .dina(n2127), .dout(n2131));
    jand g0484(.dinb(n14745), .dina(n1583), .dout(n2135));
    jor g0485(.dinb(n1956), .dina(n14743), .dout(n2139));
    jand g0486(.dinb(n17397), .dina(n2139), .dout(n2143));
    jor g0487(.dinb(n17739), .dina(n2143), .dout(n2147));
    jnot g0488(.din(n2147), .dout(n2150));
    jnot g0489(.din(n1595), .dout(n2153));
    jxor g0490(.dinb(n2153), .dina(n1610), .dout(n2157));
    jnot g0491(.din(n2157), .dout(n2160));
    jand g0492(.dinb(n2150), .dina(n17415), .dout(n2164));
    jand g0493(.dinb(n17442), .dina(n2147), .dout(n2168));
    jor g0494(.dinb(n2164), .dina(n14740), .dout(n2172));
    jnot g0495(.din(n2172), .dout(n2175));
    jnot g0496(.din(G4088), .dout(n2178));
    jnot g0497(.din(n2131), .dout(n2181));
    jor g0498(.dinb(n8625), .dina(n2181), .dout(n2185));
    jnot g0499(.din(G4087), .dout(n2188));
    jnot g0500(.din(n2040), .dout(n2191));
    jor g0501(.dinb(n15675), .dina(n2191), .dout(n2195));
    jand g0502(.dinb(n15595), .dina(n2195), .dout(n2199));
    jand g0503(.dinb(n2185), .dina(n8623), .dout(n2203));
    jor g0504(.dinb(n8686), .dina(n2178), .dout(n2207));
    jor g0505(.dinb(G11), .dina(G4088), .dout(n2211));
    jand g0506(.dinb(n15600), .dina(n2211), .dout(n2215));
    jand g0507(.dinb(n2207), .dina(n2215), .dout(n2219));
    jor g0508(.dinb(n2203), .dina(n8620), .dout(n2223));
    jand g0509(.dinb(n10369), .dina(n2003), .dout(n2227));
    jnot g0510(.din(n2227), .dout(n2230));
    jnot g0511(.din(n1894), .dout(n2233));
    jnot g0512(.din(n1898), .dout(n2236));
    jand g0513(.dinb(n17541), .dina(n1544), .dout(n2240));
    jor g0514(.dinb(n2240), .dina(n1563), .dout(n2244));
    jor g0515(.dinb(n17979), .dina(n1909), .dout(n2248));
    jand g0516(.dinb(n2248), .dina(n1548), .dout(n2252));
    jand g0517(.dinb(n2244), .dina(n2252), .dout(n2256));
    jor g0518(.dinb(n17958), .dina(n2256), .dout(n2260));
    jand g0519(.dinb(n17515), .dina(n2260), .dout(n2264));
    jor g0520(.dinb(n17506), .dina(n2264), .dout(n2268));
    jnot g0521(.din(n1501), .dout(n2271));
    jnot g0522(.din(n1575), .dout(n2274));
    jor g0523(.dinb(n11070), .dina(n2274), .dout(n2278));
    jor g0524(.dinb(n10363), .dina(n2278), .dout(n2282));
    jand g0525(.dinb(n17493), .dina(n2282), .dout(n2286));
    jxor g0526(.dinb(n17346), .dina(n2286), .dout(n2290));
    jand g0527(.dinb(n10626), .dina(n2290), .dout(n2294));
    jand g0528(.dinb(n11034), .dina(n834), .dout(n2298));
    jor g0529(.dinb(n11037), .dina(n2298), .dout(n2302));
    jor g0530(.dinb(n2294), .dina(n10342), .dout(n2306));
    jand g0531(.dinb(n10324), .dina(n2306), .dout(n2310));
    jand g0532(.dinb(n11116), .dina(n2003), .dout(n2314));
    jnot g0533(.din(n2314), .dout(n2317));
    jand g0534(.dinb(n17517), .dina(n2278), .dout(n2321));
    jxor g0535(.dinb(n17325), .dina(n2321), .dout(n2325));
    jand g0536(.dinb(n11103), .dina(n2325), .dout(n2329));
    jand g0537(.dinb(n19716), .dina(n535), .dout(n2333));
    jor g0538(.dinb(n15363), .dina(n2333), .dout(n2337));
    jor g0539(.dinb(n2329), .dina(n11020), .dout(n2341));
    jand g0540(.dinb(n11002), .dina(n2341), .dout(n2345));
    jand g0541(.dinb(n10834), .dina(n2003), .dout(n2349));
    jnot g0542(.din(n2349), .dout(n2352));
    jand g0543(.dinb(n11028), .dina(n653), .dout(n2356));
    jand g0544(.dinb(n11064), .dina(n1567), .dout(n2360));
    jor g0545(.dinb(n17535), .dina(n2360), .dout(n2364));
    jxor g0546(.dinb(n17298), .dina(n2364), .dout(n2368));
    jand g0547(.dinb(n19740), .dina(n2368), .dout(n2372));
    jor g0548(.dinb(n10929), .dina(n2372), .dout(n2376));
    jor g0549(.dinb(n10807), .dina(n2376), .dout(n2380));
    jand g0550(.dinb(n10795), .dina(n2380), .dout(n2384));
    jnot g0551(.din(G4089), .dout(n2387));
    jor g0552(.dinb(n8691), .dina(n2181), .dout(n2391));
    jnot g0553(.din(G4090), .dout(n2394));
    jor g0554(.dinb(n16083), .dina(n2191), .dout(n2398));
    jand g0555(.dinb(n16000), .dina(n2398), .dout(n2402));
    jand g0556(.dinb(n2391), .dina(n8689), .dout(n2406));
    jor g0557(.dinb(n8686), .dina(n2387), .dout(n2410));
    jor g0558(.dinb(G11), .dina(G4089), .dout(n2414));
    jand g0559(.dinb(n16008), .dina(n2414), .dout(n2418));
    jand g0560(.dinb(n2410), .dina(n2418), .dout(n2422));
    jor g0561(.dinb(n2406), .dina(n8683), .dout(n2426));
    jand g0562(.dinb(n10429), .dina(n2003), .dout(n2430));
    jnot g0563(.din(n2430), .dout(n2433));
    jnot g0564(.din(n1375), .dout(n2436));
    jnot g0565(.din(n1345), .dout(n2439));
    jand g0566(.dinb(n15039), .dina(n1301), .dout(n2443));
    jand g0567(.dinb(n18969), .dina(n2443), .dout(n2447));
    jand g0568(.dinb(n15037), .dina(n2447), .dout(n2451));
    jor g0569(.dinb(n1814), .dina(n15031), .dout(n2455));
    jxor g0570(.dinb(n18846), .dina(n2455), .dout(n2459));
    jand g0571(.dinb(n11091), .dina(n2459), .dout(n2463));
    jand g0572(.dinb(n11025), .dina(n930), .dout(n2467));
    jor g0573(.dinb(n15348), .dina(n2467), .dout(n2471));
    jor g0574(.dinb(n2463), .dina(n10417), .dout(n2475));
    jand g0575(.dinb(n10399), .dina(n2475), .dout(n2479));
    jand g0576(.dinb(n10966), .dina(n2003), .dout(n2483));
    jnot g0577(.din(n2483), .dout(n2486));
    jor g0578(.dinb(n1806), .dina(n2447), .dout(n2490));
    jxor g0579(.dinb(n18927), .dina(n2490), .dout(n2494));
    jand g0580(.dinb(n10956), .dina(n2494), .dout(n2498));
    jand g0581(.dinb(n11031), .dina(n1152), .dout(n2502));
    jor g0582(.dinb(n15348), .dina(n2502), .dout(n2506));
    jor g0583(.dinb(n2498), .dina(n10921), .dout(n2510));
    jand g0584(.dinb(n10909), .dina(n2510), .dout(n2514));
    jand g0585(.dinb(n10774), .dina(n2003), .dout(n2518));
    jnot g0586(.din(n2518), .dout(n2521));
    jor g0587(.dinb(n18981), .dina(n1786), .dout(n2525));
    jor g0588(.dinb(n2443), .dina(n2525), .dout(n2529));
    jxor g0589(.dinb(n18945), .dina(n2529), .dout(n2533));
    jand g0590(.dinb(n10953), .dina(n2533), .dout(n2537));
    jand g0591(.dinb(n11031), .dina(n1018), .dout(n2541));
    jor g0592(.dinb(n14733), .dina(n2541), .dout(n2545));
    jor g0593(.dinb(n2537), .dina(n10762), .dout(n2549));
    jand g0594(.dinb(n10753), .dina(n2549), .dout(n2553));
    jand g0595(.dinb(n10534), .dina(n2003), .dout(n2557));
    jnot g0596(.din(n2557), .dout(n2560));
    jnot g0597(.din(n1297), .dout(n2563));
    jand g0598(.dinb(n15055), .dina(n1278), .dout(n2567));
    jor g0599(.dinb(n18993), .dina(n2567), .dout(n2571));
    jxor g0600(.dinb(n10528), .dina(n2571), .dout(n2575));
    jand g0601(.dinb(n19824), .dina(n2575), .dout(n2579));
    jand g0602(.dinb(n11031), .dina(n972), .dout(n2583));
    jor g0603(.dinb(n14727), .dina(n2583), .dout(n2587));
    jor g0604(.dinb(n2579), .dina(n10513), .dout(n2591));
    jand g0605(.dinb(n10507), .dina(n2591), .dout(n2595));
    jnot g0606(.din(G331), .dout(n2598));
    jnot g0607(.din(n1497), .dout(n2601));
    jand g0608(.dinb(n11440), .dina(n2601), .dout(n2605));
    jand g0609(.dinb(n1489), .dina(n18048), .dout(n2609));
    jor g0610(.dinb(n11434), .dina(n2609), .dout(n2613));
    jxor g0611(.dinb(n2160), .dina(n2613), .dout(n2617));
    jor g0612(.dinb(G332), .dina(G369), .dout(n2621));
    jor g0613(.dinb(n1474), .dina(n11431), .dout(n2625));
    jand g0614(.dinb(n11428), .dina(n2625), .dout(n2629));
    jxor g0615(.dinb(n1563), .dina(n11425), .dout(n2633));
    jxor g0616(.dinb(n1909), .dina(n1529), .dout(n2637));
    jxor g0617(.dinb(n17820), .dina(n1648), .dout(n2641));
    jxor g0618(.dinb(n11422), .dina(n2641), .dout(n2645));
    jxor g0619(.dinb(n11419), .dina(n2645), .dout(n2649));
    jxor g0620(.dinb(n2617), .dina(n2649), .dout(n2653));
    jnot g0621(.din(n1289), .dout(n2656));
    jor g0622(.dinb(n18990), .dina(n2656), .dout(n2660));
    jxor g0623(.dinb(n2660), .dina(n1341), .dout(n2664));
    jxor g0624(.dinb(n1274), .dina(n1319), .dout(n2668));
    jxor g0625(.dinb(n2664), .dina(n2668), .dout(n2672));
    jor g0626(.dinb(G289), .dina(G335), .dout(n2676));
    jor g0627(.dinb(n11482), .dina(n1259), .dout(n2680));
    jand g0628(.dinb(n11479), .dina(n2680), .dout(n2684));
    jxor g0629(.dinb(n1391), .dina(n2684), .dout(n2688));
    jxor g0630(.dinb(n1371), .dina(n1410), .dout(n2692));
    jxor g0631(.dinb(n1429), .dina(n1452), .dout(n2696));
    jxor g0632(.dinb(n2692), .dina(n2696), .dout(n2700));
    jxor g0633(.dinb(n11476), .dina(n2700), .dout(n2704));
    jxor g0634(.dinb(n11470), .dina(n2704), .dout(n2708));
    jnot g0635(.din(n2708), .dout(n2711));
    jnot g0636(.din(n1395), .dout(n2714));
    jnot g0637(.din(n1870), .dout(n2717));
    jor g0638(.dinb(n18609), .dina(n2455), .dout(n2721));
    jand g0639(.dinb(n18582), .dina(n2721), .dout(n2725));
    jnot g0640(.din(n2725), .dout(n2728));
    jor g0641(.dinb(n18321), .dina(n2728), .dout(n2732));
    jand g0642(.dinb(n18363), .dina(n2732), .dout(n2736));
    jxor g0643(.dinb(n15028), .dina(n2736), .dout(n2740));
    jnot g0644(.din(n2740), .dout(n2743));
    jnot g0645(.din(n1437), .dout(n2746));
    jand g0646(.dinb(n14323), .dina(n2725), .dout(n2750));
    jor g0647(.dinb(n18393), .dina(n2750), .dout(n2754));
    jxor g0648(.dinb(n18471), .dina(n2754), .dout(n2758));
    jand g0649(.dinb(n2743), .dina(n14301), .dout(n2762));
    jnot g0650(.din(n1433), .dout(n2765));
    jnot g0651(.din(n1410), .dout(n2768));
    jand g0652(.dinb(n19164), .dina(n2768), .dout(n2772));
    jnot g0653(.din(n2772), .dout(n2775));
    jor g0654(.dinb(n18414), .dina(n2725), .dout(n2779));
    jand g0655(.dinb(n18540), .dina(n2779), .dout(n2783));
    jxor g0656(.dinb(n13948), .dina(n2783), .dout(n2787));
    jnot g0657(.din(n2787), .dout(n2790));
    jand g0658(.dinb(n8901), .dina(n2533), .dout(n2794));
    jand g0659(.dinb(n10521), .dina(n2794), .dout(n2798));
    jand g0660(.dinb(n2459), .dina(n8734), .dout(n2802));
    jnot g0661(.din(n1414), .dout(n2805));
    jxor g0662(.dinb(n18342), .dina(n2725), .dout(n2809));
    jnot g0663(.din(n2809), .dout(n2812));
    jand g0664(.dinb(n10938), .dina(n2812), .dout(n2816));
    jand g0665(.dinb(n8731), .dina(n2816), .dout(n2820));
    jand g0666(.dinb(n2790), .dina(n2820), .dout(n2824));
    jand g0667(.dinb(n2762), .dina(n8722), .dout(n2828));
    jxor g0668(.dinb(n14430), .dina(n2147), .dout(n2832));
    jnot g0669(.din(n2832), .dout(n2835));
    jand g0670(.dinb(n8922), .dina(n2835), .dout(n2839));
    jand g0671(.dinb(n2175), .dina(n11043), .dout(n2843));
    jand g0672(.dinb(n8755), .dina(n2843), .dout(n2847));
    jand g0673(.dinb(n17238), .dina(n2290), .dout(n2851));
    jand g0674(.dinb(n10809), .dina(n2851), .dout(n2855));
    jnot g0675(.din(n1648), .dout(n2858));
    jand g0676(.dinb(n17673), .dina(n2858), .dout(n2862));
    jand g0677(.dinb(n17811), .dina(n2862), .dout(n2866));
    jor g0678(.dinb(n17814), .dina(n2862), .dout(n2870));
    jnot g0679(.din(n2870), .dout(n2873));
    jor g0680(.dinb(n17757), .dina(n2139), .dout(n2877));
    jand g0681(.dinb(n14083), .dina(n2877), .dout(n2881));
    jnot g0682(.din(n2877), .dout(n2884));
    jand g0683(.dinb(n17694), .dina(n2884), .dout(n2888));
    jor g0684(.dinb(n14068), .dina(n2888), .dout(n2892));
    jor g0685(.dinb(n14065), .dina(n2892), .dout(n2896));
    jnot g0686(.din(n2896), .dout(n2899));
    jnot g0687(.din(n1652), .dout(n2902));
    jxor g0688(.dinb(n13759), .dina(n2139), .dout(n2906));
    jand g0689(.dinb(n2899), .dina(n13728), .dout(n2910));
    jand g0690(.dinb(n8749), .dina(n2910), .dout(n2914));
    jand g0691(.dinb(n2847), .dina(n2914), .dout(n2918));
    jnot g0692(.din(G1689), .dout(n2921));
    jand g0693(.dinb(n2921), .dina(n16617), .dout(n2925));
    jand g0694(.dinb(n8863), .dina(n2925), .dout(n2929));
    jand g0695(.dinb(G1689), .dina(G1690), .dout(n2933));
    jand g0696(.dinb(n8866), .dina(n2933), .dout(n2937));
    jor g0697(.dinb(n16377), .dina(n2181), .dout(n2941));
    jnot g0698(.din(G1690), .dout(n2944));
    jor g0699(.dinb(n16689), .dina(n2191), .dout(n2948));
    jand g0700(.dinb(n13492), .dina(n2948), .dout(n2952));
    jand g0701(.dinb(n2941), .dina(n8824), .dout(n2956));
    jor g0702(.dinb(n8821), .dina(n2956), .dout(n2960));
    jor g0703(.dinb(n8788), .dina(n2960), .dout(n2964));
    jand g0704(.dinb(n20757), .dina(n2964), .dout(n2968));
    jor g0705(.dinb(n20196), .dina(n2191), .dout(n2972));
    jnot g0706(.din(G1694), .dout(n2975));
    jnot g0707(.din(G1691), .dout(n2978));
    jor g0708(.dinb(n19956), .dina(n2181), .dout(n2982));
    jand g0709(.dinb(n14908), .dina(n2982), .dout(n2986));
    jand g0710(.dinb(n8875), .dina(n2986), .dout(n2990));
    jand g0711(.dinb(G1691), .dina(G1694), .dout(n2994));
    jand g0712(.dinb(n8866), .dina(n2994), .dout(n2998));
    jand g0713(.dinb(n2978), .dina(n20298), .dout(n3002));
    jand g0714(.dinb(n8863), .dina(n3002), .dout(n3006));
    jor g0715(.dinb(n8857), .dina(n3006), .dout(n3010));
    jor g0716(.dinb(n2990), .dina(n8854), .dout(n3014));
    jand g0717(.dinb(n20757), .dina(n3014), .dout(n3018));
    jnot g0718(.din(n2479), .dout(n3021));
    jor g0719(.dinb(n9216), .dina(n3021), .dout(n3025));
    jnot g0720(.din(n2310), .dout(n3028));
    jor g0721(.dinb(n9129), .dina(n3028), .dout(n3032));
    jand g0722(.dinb(n9012), .dina(n3032), .dout(n3036));
    jand g0723(.dinb(n9010), .dina(n3036), .dout(n3040));
    jor g0724(.dinb(n9514), .dina(n2178), .dout(n3044));
    jor g0725(.dinb(G43), .dina(G4088), .dout(n3048));
    jand g0726(.dinb(n15597), .dina(n3048), .dout(n3052));
    jand g0727(.dinb(n3044), .dina(n3052), .dout(n3056));
    jor g0728(.dinb(n3040), .dina(n9007), .dout(n3060));
    jnot g0729(.din(n2514), .dout(n3063));
    jor g0730(.dinb(n9177), .dina(n3063), .dout(n3067));
    jnot g0731(.din(n2345), .dout(n3070));
    jor g0732(.dinb(n9084), .dina(n3070), .dout(n3074));
    jand g0733(.dinb(n9432), .dina(n3074), .dout(n3078));
    jand g0734(.dinb(n9082), .dina(n3078), .dout(n3082));
    jor g0735(.dinb(n9613), .dina(n2178), .dout(n3086));
    jor g0736(.dinb(G76), .dina(G4088), .dout(n3090));
    jand g0737(.dinb(n15714), .dina(n3090), .dout(n3094));
    jand g0738(.dinb(n3086), .dina(n3094), .dout(n3098));
    jor g0739(.dinb(n3082), .dina(n9076), .dout(n3102));
    jnot g0740(.din(n2384), .dout(n3105));
    jor g0741(.dinb(n9339), .dina(n3105), .dout(n3109));
    jnot g0742(.din(n2553), .dout(n3112));
    jor g0743(.dinb(n9303), .dina(n3112), .dout(n3116));
    jand g0744(.dinb(n15558), .dina(n3116), .dout(n3120));
    jand g0745(.dinb(n9301), .dina(n3120), .dout(n3124));
    jor g0746(.dinb(n9781), .dina(n2178), .dout(n3128));
    jor g0747(.dinb(G73), .dina(G4088), .dout(n3132));
    jand g0748(.dinb(n15714), .dina(n3132), .dout(n3136));
    jand g0749(.dinb(n3128), .dina(n3136), .dout(n3140));
    jor g0750(.dinb(n3124), .dina(n9298), .dout(n3144));
    jnot g0751(.din(n2595), .dout(n3147));
    jor g0752(.dinb(n11754), .dina(n3147), .dout(n3151));
    jnot g0753(.din(n2097), .dout(n3154));
    jor g0754(.dinb(n11847), .dina(n3154), .dout(n3158));
    jand g0755(.dinb(n9429), .dina(n3158), .dout(n3162));
    jand g0756(.dinb(n9427), .dina(n3162), .dout(n3166));
    jor g0757(.dinb(n9916), .dina(n2178), .dout(n3170));
    jor g0758(.dinb(G67), .dina(G4088), .dout(n3174));
    jand g0759(.dinb(n15714), .dina(n3174), .dout(n3178));
    jand g0760(.dinb(n3170), .dina(n3178), .dout(n3182));
    jor g0761(.dinb(n3166), .dina(n9418), .dout(n3186));
    jor g0762(.dinb(G43), .dina(G4089), .dout(n3190));
    jor g0763(.dinb(n9514), .dina(n2387), .dout(n3194));
    jand g0764(.dinb(n16002), .dina(n3194), .dout(n3198));
    jand g0765(.dinb(n9511), .dina(n3198), .dout(n3202));
    jor g0766(.dinb(n9615), .dina(n3028), .dout(n3206));
    jor g0767(.dinb(n9567), .dina(n3021), .dout(n3210));
    jand g0768(.dinb(n3206), .dina(n3210), .dout(n3214));
    jand g0769(.dinb(n9483), .dina(n3214), .dout(n3218));
    jor g0770(.dinb(n9481), .dina(n3218), .dout(n3222));
    jor g0771(.dinb(G76), .dina(G4089), .dout(n3226));
    jor g0772(.dinb(n9613), .dina(n2387), .dout(n3230));
    jand g0773(.dinb(n9912), .dina(n3230), .dout(n3234));
    jand g0774(.dinb(n9565), .dina(n3234), .dout(n3238));
    jor g0775(.dinb(n9822), .dina(n3070), .dout(n3242));
    jor g0776(.dinb(n9741), .dina(n3063), .dout(n3246));
    jand g0777(.dinb(n3242), .dina(n9559), .dout(n3250));
    jand g0778(.dinb(n9927), .dina(n3250), .dout(n3254));
    jor g0779(.dinb(n9556), .dina(n3254), .dout(n3258));
    jor g0780(.dinb(G73), .dina(G4089), .dout(n3262));
    jor g0781(.dinb(n9781), .dina(n2387), .dout(n3266));
    jand g0782(.dinb(n9909), .dina(n3266), .dout(n3270));
    jand g0783(.dinb(n9703), .dina(n3270), .dout(n3274));
    jor g0784(.dinb(n9705), .dina(n3112), .dout(n3278));
    jor g0785(.dinb(n9783), .dina(n3105), .dout(n3282));
    jand g0786(.dinb(n3278), .dina(n3282), .dout(n3286));
    jand g0787(.dinb(n15960), .dina(n3286), .dout(n3290));
    jor g0788(.dinb(n9697), .dina(n3290), .dout(n3294));
    jor g0789(.dinb(n11547), .dina(n3147), .dout(n3298));
    jor g0790(.dinb(n11580), .dina(n3154), .dout(n3302));
    jand g0791(.dinb(n15960), .dina(n3302), .dout(n3306));
    jand g0792(.dinb(n9925), .dina(n3306), .dout(n3310));
    jor g0793(.dinb(n9916), .dina(n2387), .dout(n3314));
    jor g0794(.dinb(G67), .dina(G4089), .dout(n3318));
    jand g0795(.dinb(n16125), .dina(n3318), .dout(n3322));
    jand g0796(.dinb(n3314), .dina(n3322), .dout(n3326));
    jor g0797(.dinb(n3310), .dina(n9907), .dout(n3330));
    jor g0798(.dinb(n10071), .dina(n3028), .dout(n3334));
    jor g0799(.dinb(n16332), .dina(n3021), .dout(n3338));
    jand g0800(.dinb(n10035), .dina(n3338), .dout(n3342));
    jand g0801(.dinb(n9982), .dina(n3342), .dout(n3346));
    jand g0802(.dinb(n10438), .dina(n2925), .dout(n3350));
    jand g0803(.dinb(n10432), .dina(n2933), .dout(n3354));
    jor g0804(.dinb(n3350), .dina(n9979), .dout(n3358));
    jor g0805(.dinb(n3346), .dina(n9976), .dout(n3362));
    jand g0806(.dinb(n10134), .dina(n3362), .dout(n3366));
    jor g0807(.dinb(n10056), .dina(n3154), .dout(n3370));
    jor g0808(.dinb(n16584), .dina(n3147), .dout(n3374));
    jand g0809(.dinb(n10026), .dina(n3374), .dout(n3378));
    jand g0810(.dinb(n3370), .dina(n10024), .dout(n3382));
    jand g0811(.dinb(n10486), .dina(n2925), .dout(n3386));
    jand g0812(.dinb(n10480), .dina(n2933), .dout(n3390));
    jor g0813(.dinb(n3386), .dina(n10021), .dout(n3394));
    jor g0814(.dinb(n3382), .dina(n10018), .dout(n3398));
    jand g0815(.dinb(n10677), .dina(n3398), .dout(n3402));
    jor g0816(.dinb(n16839), .dina(n3105), .dout(n3406));
    jor g0817(.dinb(n10191), .dina(n3112), .dout(n3410));
    jand g0818(.dinb(n13455), .dina(n3410), .dout(n3414));
    jand g0819(.dinb(n10132), .dina(n3414), .dout(n3418));
    jand g0820(.dinb(n10729), .dina(n2925), .dout(n3422));
    jand g0821(.dinb(n10723), .dina(n2933), .dout(n3426));
    jor g0822(.dinb(n3422), .dina(n10129), .dout(n3430));
    jor g0823(.dinb(n3418), .dina(n10126), .dout(n3434));
    jand g0824(.dinb(n10677), .dina(n3434), .dout(n3438));
    jor g0825(.dinb(n13185), .dina(n3070), .dout(n3442));
    jor g0826(.dinb(n10185), .dina(n3063), .dout(n3446));
    jand g0827(.dinb(n13170), .dina(n3446), .dout(n3450));
    jand g0828(.dinb(n3442), .dina(n3450), .dout(n3454));
    jand g0829(.dinb(n10885), .dina(n2925), .dout(n3458));
    jand g0830(.dinb(n10879), .dina(n2933), .dout(n3462));
    jor g0831(.dinb(n3458), .dina(n10183), .dout(n3466));
    jor g0832(.dinb(n3454), .dina(n10180), .dout(n3470));
    jand g0833(.dinb(n10668), .dina(n3470), .dout(n3474));
    jand g0834(.dinb(n10438), .dina(n3002), .dout(n3478));
    jand g0835(.dinb(n10432), .dina(n2994), .dout(n3482));
    jor g0836(.dinb(n19911), .dina(n3021), .dout(n3486));
    jor g0837(.dinb(n20343), .dina(n3028), .dout(n3490));
    jand g0838(.dinb(n3486), .dina(n3490), .dout(n3494));
    jand g0839(.dinb(n10539), .dina(n3494), .dout(n3498));
    jor g0840(.dinb(n10294), .dina(n3498), .dout(n3502));
    jor g0841(.dinb(n10243), .dina(n3502), .dout(n3506));
    jand g0842(.dinb(n10656), .dina(n3506), .dout(n3510));
    jor g0843(.dinb(n20301), .dina(n3154), .dout(n3514));
    jor g0844(.dinb(n20163), .dina(n3147), .dout(n3518));
    jand g0845(.dinb(n10536), .dina(n3518), .dout(n3522));
    jand g0846(.dinb(n3514), .dina(n10489), .dout(n3526));
    jand g0847(.dinb(n10486), .dina(n3002), .dout(n3530));
    jand g0848(.dinb(n10480), .dina(n2994), .dout(n3534));
    jor g0849(.dinb(n3530), .dina(n10477), .dout(n3538));
    jor g0850(.dinb(n3526), .dina(n10474), .dout(n3542));
    jand g0851(.dinb(n10671), .dina(n3542), .dout(n3546));
    jor g0852(.dinb(n20514), .dina(n3105), .dout(n3550));
    jor g0853(.dinb(n10974), .dina(n3112), .dout(n3554));
    jand g0854(.dinb(n14871), .dina(n3554), .dout(n3558));
    jand g0855(.dinb(n10732), .dina(n3558), .dout(n3562));
    jand g0856(.dinb(n10729), .dina(n3002), .dout(n3566));
    jand g0857(.dinb(n10723), .dina(n2994), .dout(n3570));
    jor g0858(.dinb(n3566), .dina(n10720), .dout(n3574));
    jor g0859(.dinb(n3562), .dina(n10717), .dout(n3578));
    jand g0860(.dinb(n20706), .dina(n3578), .dout(n3582));
    jor g0861(.dinb(n13779), .dina(n3070), .dout(n3586));
    jor g0862(.dinb(n10968), .dina(n3063), .dout(n3590));
    jand g0863(.dinb(n13671), .dina(n3590), .dout(n3594));
    jand g0864(.dinb(n3586), .dina(n3594), .dout(n3598));
    jand g0865(.dinb(n10885), .dina(n3002), .dout(n3602));
    jand g0866(.dinb(n10879), .dina(n2994), .dout(n3606));
    jor g0867(.dinb(n3602), .dina(n10876), .dout(n3610));
    jor g0868(.dinb(n3598), .dina(n10873), .dout(n3614));
    jand g0869(.dinb(n13209), .dina(n3614), .dout(n3618));
    jnot g0870(.din(G135), .dout(n3621));
    jnot g0871(.din(G4115), .dout(n3624));
    jor g0872(.dinb(n3621), .dina(n3624), .dout(n3628));
    jnot g0873(.din(n770), .dout(n3631));
    jor g0874(.dinb(n11331), .dina(n3631), .dout(n3635));
    jnot g0875(.din(G3717), .dout(n3638));
    jnot g0876(.din(G3724), .dout(n3641));
    jxor g0877(.dinb(n11386), .dina(n2153), .dout(n3645));
    jnot g0878(.din(n3645), .dout(n3648));
    jor g0879(.dinb(n11323), .dina(n3648), .dout(n3652));
    jand g0880(.dinb(n11275), .dina(n3652), .dout(n3656));
    jand g0881(.dinb(n11257), .dina(n3656), .dout(n3660));
    jor g0882(.dinb(n11277), .dina(n2172), .dout(n3664));
    jor g0883(.dinb(G123), .dina(G3724), .dout(n3668));
    jand g0884(.dinb(n11325), .dina(n3668), .dout(n3672));
    jand g0885(.dinb(n3664), .dina(n11248), .dout(n3676));
    jor g0886(.dinb(n11200), .dina(n3676), .dout(n3680));
    jand g0887(.dinb(n11170), .dina(n3680), .dout(n3684));
    jxor g0888(.dinb(n2172), .dina(n11343), .dout(n3688));
    jand g0889(.dinb(n14829), .dina(n2003), .dout(n3692));
    jor g0890(.dinb(n14787), .dina(n2172), .dout(n3696));
    jand g0891(.dinb(n19710), .dina(n770), .dout(n3700));
    jor g0892(.dinb(n18183), .dina(n3700), .dout(n3704));
    jnot g0893(.din(n3704), .dout(n3707));
    jand g0894(.dinb(n3696), .dina(n14725), .dout(n3711));
    jor g0895(.dinb(n14689), .dina(n3711), .dout(n3715));
    jnot g0896(.din(n3715), .dout(n3718));
    jand g0897(.dinb(n14527), .dina(n2003), .dout(n3722));
    jand g0898(.dinb(n14784), .dina(n788), .dout(n3726));
    jnot g0899(.din(n3726), .dout(n3729));
    jnot g0900(.din(G4092), .dout(n3732));
    jor g0901(.dinb(n14493), .dina(n2832), .dout(n3736));
    jand g0902(.dinb(n15109), .dina(n3736), .dout(n3740));
    jand g0903(.dinb(n14428), .dina(n3740), .dout(n3744));
    jor g0904(.dinb(n14395), .dina(n3744), .dout(n3748));
    jnot g0905(.din(n3748), .dout(n3751));
    jand g0906(.dinb(n14089), .dina(n2003), .dout(n3755));
    jor g0907(.dinb(n14457), .dina(n2896), .dout(n3759));
    jand g0908(.dinb(n15189), .dina(n751), .dout(n3763));
    jor g0909(.dinb(n15129), .dina(n3763), .dout(n3767));
    jnot g0910(.din(n3767), .dout(n3770));
    jand g0911(.dinb(n3759), .dina(n14038), .dout(n3774));
    jor g0912(.dinb(n14008), .dina(n3774), .dout(n3778));
    jnot g0913(.din(n3778), .dout(n3781));
    jand g0914(.dinb(n13765), .dina(n2003), .dout(n3785));
    jnot g0915(.din(n3785), .dout(n3788));
    jand g0916(.dinb(n19785), .dina(n2906), .dout(n3792));
    jand g0917(.dinb(n15183), .dina(n709), .dout(n3796));
    jor g0918(.dinb(n15111), .dina(n3796), .dout(n3800));
    jor g0919(.dinb(n3792), .dina(n13726), .dout(n3804));
    jand g0920(.dinb(n13705), .dina(n3804), .dout(n3808));
    jand g0921(.dinb(n11457), .dina(n1735), .dout(n3812));
    jand g0922(.dinb(n2708), .dina(n11449), .dout(n3816));
    jnot g0923(.din(n2653), .dout(n3819));
    jand g0924(.dinb(n313), .dina(n360), .dout(n3823));
    jand g0925(.dinb(n11406), .dina(n3823), .dout(n3827));
    jand g0926(.dinb(n1696), .dina(n11404), .dout(n3831));
    jand g0927(.dinb(n3819), .dina(n11401), .dout(n3835));
    jand g0928(.dinb(n11389), .dina(n3835), .dout(n3839));
    jand g0929(.dinb(n15199), .dina(n2003), .dout(n3843));
    jand g0930(.dinb(n15183), .dina(n1240), .dout(n3847));
    jnot g0931(.din(n3847), .dout(n3850));
    jor g0932(.dinb(n15147), .dina(n2740), .dout(n3854));
    jand g0933(.dinb(n15060), .dina(n3854), .dout(n3858));
    jand g0934(.dinb(n14995), .dina(n3858), .dout(n3862));
    jor g0935(.dinb(n14959), .dina(n3862), .dout(n3866));
    jnot g0936(.din(n3866), .dout(n3869));
    jand g0937(.dinb(n14344), .dina(n2003), .dout(n3873));
    jnot g0938(.din(n3873), .dout(n3876));
    jand g0939(.dinb(n14331), .dina(n2758), .dout(n3880));
    jand g0940(.dinb(n19698), .dina(n888), .dout(n3884));
    jor g0941(.dinb(n18165), .dina(n3884), .dout(n3888));
    jor g0942(.dinb(n3880), .dina(n14248), .dout(n3892));
    jand g0943(.dinb(n14218), .dina(n3892), .dout(n3896));
    jand g0944(.dinb(n13960), .dina(n2003), .dout(n3900));
    jand g0945(.dinb(n19698), .dina(n1110), .dout(n3904));
    jnot g0946(.din(n3904), .dout(n3907));
    jor g0947(.dinb(n14268), .dina(n2787), .dout(n3911));
    jand g0948(.dinb(n15057), .dina(n3911), .dout(n3915));
    jand g0949(.dinb(n13921), .dina(n3915), .dout(n3919));
    jor g0950(.dinb(n13888), .dina(n3919), .dout(n3923));
    jnot g0951(.din(n3923), .dout(n3926));
    jand g0952(.dinb(n13651), .dina(n2003), .dout(n3930));
    jnot g0953(.din(n3930), .dout(n3933));
    jand g0954(.dinb(n14325), .dina(n2812), .dout(n3937));
    jand g0955(.dinb(n19686), .dina(n1060), .dout(n3941));
    jor g0956(.dinb(n18165), .dina(n3941), .dout(n3945));
    jor g0957(.dinb(n3937), .dina(n13639), .dout(n3949));
    jand g0958(.dinb(n13612), .dina(n3949), .dout(n3953));
    jor g0959(.dinb(G109), .dina(G4089), .dout(n3957));
    jor g0960(.dinb(n11686), .dina(n2387), .dout(n3961));
    jand g0961(.dinb(n12786), .dina(n3961), .dout(n3965));
    jand g0962(.dinb(n11545), .dina(n3965), .dout(n3969));
    jor g0963(.dinb(n12549), .dina(n3866), .dout(n3973));
    jor g0964(.dinb(n12666), .dina(n3715), .dout(n3977));
    jand g0965(.dinb(n15927), .dina(n3977), .dout(n3981));
    jand g0966(.dinb(n3973), .dina(n3981), .dout(n3985));
    jor g0967(.dinb(n11539), .dina(n3985), .dout(n3989));
    jor g0968(.dinb(n11787), .dina(n3715), .dout(n3993));
    jor g0969(.dinb(n11694), .dina(n3866), .dout(n3997));
    jand g0970(.dinb(n12132), .dina(n3997), .dout(n4001));
    jand g0971(.dinb(n11692), .dina(n4001), .dout(n4005));
    jor g0972(.dinb(n11686), .dina(n2178), .dout(n4009));
    jor g0973(.dinb(G109), .dina(G4088), .dout(n4013));
    jand g0974(.dinb(n15711), .dina(n4013), .dout(n4017));
    jand g0975(.dinb(n4009), .dina(n4017), .dout(n4021));
    jor g0976(.dinb(n4005), .dina(n11683), .dout(n4025));
    jor g0977(.dinb(n12012), .dina(n3748), .dout(n4029));
    jnot g0978(.din(n3896), .dout(n4032));
    jor g0979(.dinb(n11955), .dina(n4032), .dout(n4036));
    jand g0980(.dinb(n15525), .dina(n4036), .dout(n4040));
    jand g0981(.dinb(n11953), .dina(n4040), .dout(n4044));
    jor g0982(.dinb(n12484), .dina(n2178), .dout(n4048));
    jor g0983(.dinb(G46), .dina(G4088), .dout(n4052));
    jand g0984(.dinb(n15711), .dina(n4052), .dout(n4056));
    jand g0985(.dinb(n4048), .dina(n4056), .dout(n4060));
    jor g0986(.dinb(n4044), .dina(n11947), .dout(n4064));
    jor g0987(.dinb(n12363), .dina(n3778), .dout(n4068));
    jor g0988(.dinb(n12255), .dina(n3923), .dout(n4072));
    jand g0989(.dinb(n15525), .dina(n4072), .dout(n4076));
    jand g0990(.dinb(n12130), .dina(n4076), .dout(n4080));
    jor g0991(.dinb(n12790), .dina(n2178), .dout(n4084));
    jor g0992(.dinb(G100), .dina(G4088), .dout(n4088));
    jand g0993(.dinb(n15711), .dina(n4088), .dout(n4092));
    jand g0994(.dinb(n4084), .dina(n4092), .dout(n4096));
    jor g0995(.dinb(n4080), .dina(n12127), .dout(n4100));
    jnot g0996(.din(n3808), .dout(n4103));
    jor g0997(.dinb(n12312), .dina(n4103), .dout(n4107));
    jnot g0998(.din(n3953), .dout(n4110));
    jor g0999(.dinb(n12201), .dina(n4110), .dout(n4114));
    jand g1000(.dinb(n15495), .dina(n4114), .dout(n4118));
    jand g1001(.dinb(n12199), .dina(n4118), .dout(n4122));
    jor g1002(.dinb(n12853), .dina(n2178), .dout(n4126));
    jor g1003(.dinb(G91), .dina(G4088), .dout(n4130));
    jand g1004(.dinb(n15708), .dina(n4130), .dout(n4134));
    jand g1005(.dinb(n4126), .dina(n4134), .dout(n4138));
    jor g1006(.dinb(n4122), .dina(n12190), .dout(n4142));
    jor g1007(.dinb(n12609), .dina(n3748), .dout(n4146));
    jor g1008(.dinb(n12492), .dina(n4032), .dout(n4150));
    jand g1009(.dinb(n15927), .dina(n4150), .dout(n4154));
    jand g1010(.dinb(n12490), .dina(n4154), .dout(n4158));
    jor g1011(.dinb(n12484), .dina(n2387), .dout(n4162));
    jor g1012(.dinb(G46), .dina(G4089), .dout(n4166));
    jand g1013(.dinb(n16122), .dina(n4166), .dout(n4170));
    jand g1014(.dinb(n4162), .dina(n4170), .dout(n4174));
    jor g1015(.dinb(n4158), .dina(n12481), .dout(n4178));
    jor g1016(.dinb(n13026), .dina(n3778), .dout(n4182));
    jor g1017(.dinb(n12918), .dina(n3923), .dout(n4186));
    jand g1018(.dinb(n15927), .dina(n4186), .dout(n4190));
    jand g1019(.dinb(n12793), .dina(n4190), .dout(n4194));
    jor g1020(.dinb(n12790), .dina(n2387), .dout(n4198));
    jor g1021(.dinb(G100), .dina(G4089), .dout(n4202));
    jand g1022(.dinb(n16122), .dina(n4202), .dout(n4206));
    jand g1023(.dinb(n4198), .dina(n4206), .dout(n4210));
    jor g1024(.dinb(n4194), .dina(n12784), .dout(n4214));
    jor g1025(.dinb(n12975), .dina(n4103), .dout(n4218));
    jor g1026(.dinb(n12864), .dina(n4110), .dout(n4222));
    jand g1027(.dinb(n15897), .dina(n4222), .dout(n4226));
    jand g1028(.dinb(n12862), .dina(n4226), .dout(n4230));
    jor g1029(.dinb(n12853), .dina(n2387), .dout(n4234));
    jor g1030(.dinb(G91), .dina(G4089), .dout(n4238));
    jand g1031(.dinb(n16119), .dina(n4238), .dout(n4242));
    jand g1032(.dinb(n4234), .dina(n4242), .dout(n4246));
    jor g1033(.dinb(n4230), .dina(n12850), .dout(n4250));
    jor g1034(.dinb(n13173), .dina(n4103), .dout(n4254));
    jor g1035(.dinb(n16530), .dina(n4110), .dout(n4258));
    jand g1036(.dinb(n13152), .dina(n4258), .dout(n4262));
    jand g1037(.dinb(n13150), .dina(n4262), .dout(n4266));
    jand g1038(.dinb(n13564), .dina(n2925), .dout(n4270));
    jand g1039(.dinb(n13558), .dina(n2933), .dout(n4274));
    jor g1040(.dinb(n4270), .dina(n13141), .dout(n4278));
    jor g1041(.dinb(n4266), .dina(n13138), .dout(n4282));
    jand g1042(.dinb(n13191), .dina(n4282), .dout(n4286));
    jor g1043(.dinb(n13338), .dina(n3923), .dout(n4290));
    jor g1044(.dinb(n13410), .dina(n3778), .dout(n4294));
    jand g1045(.dinb(n13422), .dina(n4294), .dout(n4298));
    jand g1046(.dinb(n13273), .dina(n4298), .dout(n4302));
    jand g1047(.dinb(n14101), .dina(n2925), .dout(n4306));
    jand g1048(.dinb(n14095), .dina(n2933), .dout(n4310));
    jor g1049(.dinb(n4306), .dina(n13270), .dout(n4314));
    jor g1050(.dinb(n4302), .dina(n13267), .dout(n4318));
    jand g1051(.dinb(n14553), .dina(n4318), .dout(n4322));
    jand g1052(.dinb(n14170), .dina(n2925), .dout(n4326));
    jand g1053(.dinb(n14164), .dina(n2933), .dout(n4330));
    jor g1054(.dinb(n4326), .dina(n13342), .dout(n4334));
    jor g1055(.dinb(n16782), .dina(n3748), .dout(n4338));
    jor g1056(.dinb(n13335), .dina(n4032), .dout(n4342));
    jand g1057(.dinb(n13333), .dina(n4342), .dout(n4346));
    jand g1058(.dinb(n13419), .dina(n4346), .dout(n4350));
    jor g1059(.dinb(n13330), .dina(n4350), .dout(n4354));
    jand g1060(.dinb(n14553), .dina(n4354), .dout(n4358));
    jand g1061(.dinb(n14641), .dina(n2925), .dout(n4362));
    jand g1062(.dinb(n14635), .dina(n2933), .dout(n4366));
    jor g1063(.dinb(n4362), .dina(n13495), .dout(n4370));
    jor g1064(.dinb(n13407), .dina(n3715), .dout(n4374));
    jor g1065(.dinb(n16470), .dina(n3866), .dout(n4378));
    jand g1066(.dinb(n13405), .dina(n4378), .dout(n4382));
    jand g1067(.dinb(n13413), .dina(n4382), .dout(n4386));
    jor g1068(.dinb(n13402), .dina(n4386), .dout(n4390));
    jand g1069(.dinb(n13497), .dina(n4390), .dout(n4394));
    jor g1070(.dinb(n13767), .dina(n4103), .dout(n4398));
    jor g1071(.dinb(n20109), .dina(n4110), .dout(n4402));
    jand g1072(.dinb(n13653), .dina(n4402), .dout(n4406));
    jand g1073(.dinb(n13573), .dina(n4406), .dout(n4410));
    jand g1074(.dinb(n13564), .dina(n3002), .dout(n4414));
    jand g1075(.dinb(n13558), .dina(n2994), .dout(n4418));
    jor g1076(.dinb(n4414), .dina(n13555), .dout(n4422));
    jor g1077(.dinb(n4410), .dina(n13552), .dout(n4426));
    jand g1078(.dinb(n14535), .dina(n4426), .dout(n4430));
    jand g1079(.dinb(n14101), .dina(n3002), .dout(n4434));
    jand g1080(.dinb(n14095), .dina(n2994), .dout(n4438));
    jor g1081(.dinb(n4434), .dina(n14092), .dout(n4442));
    jor g1082(.dinb(n14838), .dina(n3778), .dout(n4446));
    jor g1083(.dinb(n14349), .dina(n3923), .dout(n4450));
    jand g1084(.dinb(n4446), .dina(n4450), .dout(n4454));
    jand g1085(.dinb(n14841), .dina(n4454), .dout(n4458));
    jor g1086(.dinb(n13840), .dina(n4458), .dout(n4462));
    jand g1087(.dinb(n14532), .dina(n4462), .dout(n4466));
    jor g1088(.dinb(n20457), .dina(n3748), .dout(n4470));
    jor g1089(.dinb(n14346), .dina(n4032), .dout(n4474));
    jand g1090(.dinb(n14844), .dina(n4474), .dout(n4478));
    jand g1091(.dinb(n14176), .dina(n4478), .dout(n4482));
    jand g1092(.dinb(n14170), .dina(n3002), .dout(n4486));
    jand g1093(.dinb(n14164), .dina(n2994), .dout(n4490));
    jor g1094(.dinb(n4486), .dina(n14161), .dout(n4494));
    jor g1095(.dinb(n4482), .dina(n14158), .dout(n4498));
    jand g1096(.dinb(n14529), .dina(n4498), .dout(n4502));
    jor g1097(.dinb(n20049), .dina(n3866), .dout(n4506));
    jor g1098(.dinb(n14835), .dina(n3715), .dout(n4510));
    jand g1099(.dinb(n14844), .dina(n4510), .dout(n4514));
    jand g1100(.dinb(n4506), .dina(n4514), .dout(n4518));
    jand g1101(.dinb(n14641), .dina(n3002), .dout(n4522));
    jand g1102(.dinb(n14635), .dina(n2994), .dout(n4526));
    jor g1103(.dinb(n4522), .dina(n14632), .dout(n4530));
    jor g1104(.dinb(n4518), .dina(n14629), .dout(n4534));
    jand g1105(.dinb(n20634), .dina(n4534), .dout(n4538));
    jand g1106(.dinb(n17868), .dina(n1988), .dout(n4542));
    jxor g1107(.dinb(n17814), .dina(n2862), .dout(n4546));
    jxor g1108(.dinb(n17718), .dina(n4546), .dout(n4550));
    jxor g1109(.dinb(n4542), .dina(n17671), .dout(n4554));
    jor g1110(.dinb(n1956), .dina(n4554), .dout(n4558));
    jnot g1111(.din(G2174), .dout(n4561));
    jnot g1112(.din(n1886), .dout(n4564));
    jnot g1113(.din(n1890), .dout(n4567));
    jor g1114(.dinb(n17491), .dina(n2268), .dout(n4571));
    jand g1115(.dinb(n17482), .dina(n4571), .dout(n4575));
    jxor g1116(.dinb(n17818), .dina(n1974), .dout(n4579));
    jxor g1117(.dinb(n2160), .dina(n4579), .dout(n4583));
    jnot g1118(.din(n1656), .dout(n4586));
    jand g1119(.dinb(n17856), .dina(n1985), .dout(n4590));
    jand g1120(.dinb(n17395), .dina(n4590), .dout(n4594));
    jxor g1121(.dinb(n17389), .dina(n4594), .dout(n4598));
    jor g1122(.dinb(n4575), .dina(n4598), .dout(n4602));
    jand g1123(.dinb(n17562), .dina(n4602), .dout(n4606));
    jand g1124(.dinb(n17377), .dina(n4606), .dout(n4610));
    jnot g1125(.din(n4610), .dout(n4613));
    jnot g1126(.din(n1583), .dout(n4616));
    jand g1127(.dinb(n17278), .dina(n4575), .dout(n4620));
    jor g1128(.dinb(n17379), .dina(n4620), .dout(n4624));
    jnot g1129(.din(n4624), .dout(n4627));
    jnot g1130(.din(n4554), .dout(n4630));
    jand g1131(.dinb(n4630), .dina(n4620), .dout(n4634));
    jor g1132(.dinb(n17556), .dina(n4634), .dout(n4638));
    jor g1133(.dinb(n4627), .dina(n4638), .dout(n4642));
    jand g1134(.dinb(n4613), .dina(n4642), .dout(n4646));
    jor g1135(.dinb(n1567), .dina(n1920), .dout(n4650));
    jxor g1136(.dinb(n1940), .dina(n17272), .dout(n4654));
    jxor g1137(.dinb(n1948), .dina(n17269), .dout(n4658));
    jor g1138(.dinb(n17634), .dina(n4658), .dout(n4662));
    jor g1139(.dinb(n17286), .dina(n1948), .dout(n4666));
    jor g1140(.dinb(n17919), .dina(n2260), .dout(n4670));
    jor g1141(.dinb(n17526), .dina(n1940), .dout(n4674));
    jor g1142(.dinb(n17289), .dina(n4674), .dout(n4678));
    jand g1143(.dinb(n17266), .dina(n4678), .dout(n4682));
    jxor g1144(.dinb(n4666), .dina(n4682), .dout(n4686));
    jor g1145(.dinb(n17593), .dina(n4686), .dout(n4690));
    jand g1146(.dinb(n17263), .dina(n4690), .dout(n4694));
    jxor g1147(.dinb(n1493), .dina(n17319), .dout(n4698));
    jxor g1148(.dinb(n17292), .dina(n2065), .dout(n4702));
    jxor g1149(.dinb(n17236), .dina(n4702), .dout(n4706));
    jxor g1150(.dinb(n4694), .dina(n17227), .dout(n4710));
    jnot g1151(.din(n4710), .dout(n4713));
    jand g1152(.dinb(n4646), .dina(n17212), .dout(n4717));
    jor g1153(.dinb(n17280), .dina(n1956), .dout(n4721));
    jor g1154(.dinb(n17664), .dina(n4721), .dout(n4725));
    jand g1155(.dinb(n17595), .dina(n4725), .dout(n4729));
    jand g1156(.dinb(n17274), .dina(n4729), .dout(n4733));
    jor g1157(.dinb(n17373), .dina(n4733), .dout(n4737));
    jand g1158(.dinb(n4737), .dina(n17214), .dout(n4741));
    jor g1159(.dinb(n17175), .dina(n4741), .dout(n4745));
    jor g1160(.dinb(n17164), .dina(n4745), .dout(n4749));
    jand g1161(.dinb(G248), .dina(G351), .dout(n4753));
    jand g1162(.dinb(n19434), .dina(n566), .dout(n4757));
    jor g1163(.dinb(n17545), .dina(n4757), .dout(n4761));
    jor g1164(.dinb(n17158), .dina(n4761), .dout(n4765));
    jand g1165(.dinb(n686), .dina(n566), .dout(n4769));
    jand g1166(.dinb(n693), .dina(n17937), .dout(n4773));
    jor g1167(.dinb(n4769), .dina(n4773), .dout(n4777));
    jor g1168(.dinb(n17949), .dina(n4777), .dout(n4781));
    jand g1169(.dinb(n4765), .dina(n4781), .dout(n4785));
    jand g1170(.dinb(G248), .dina(G341), .dout(n4789));
    jand g1171(.dinb(n19554), .dina(n614), .dout(n4793));
    jor g1172(.dinb(n17983), .dina(n4793), .dout(n4797));
    jor g1173(.dinb(n17149), .dina(n4797), .dout(n4801));
    jand g1174(.dinb(n686), .dina(n614), .dout(n4805));
    jand g1175(.dinb(n693), .dina(n17973), .dout(n4809));
    jor g1176(.dinb(n4805), .dina(n4809), .dout(n4813));
    jor g1177(.dinb(n18003), .dina(n4813), .dout(n4817));
    jand g1178(.dinb(n4801), .dina(n4817), .dout(n4821));
    jxor g1179(.dinb(n4785), .dina(n4821), .dout(n4825));
    jor g1180(.dinb(n548), .dina(n795), .dout(n4829));
    jor g1181(.dinb(n538), .dina(n18102), .dout(n4833));
    jand g1182(.dinb(n18117), .dina(n4833), .dout(n4837));
    jand g1183(.dinb(n17143), .dina(n4837), .dout(n4841));
    jor g1184(.dinb(G254), .dina(G324), .dout(n4845));
    jor g1185(.dinb(n19533), .dina(n795), .dout(n4849));
    jand g1186(.dinb(n17125), .dina(n4849), .dout(n4853));
    jand g1187(.dinb(n17127), .dina(n4853), .dout(n4857));
    jor g1188(.dinb(n4841), .dina(n4857), .dout(n4861));
    jor g1189(.dinb(n693), .dina(n18063), .dout(n4865));
    jor g1190(.dinb(n19608), .dina(n521), .dout(n4869));
    jand g1191(.dinb(n4865), .dina(n4869), .dout(n4873));
    jxor g1192(.dinb(n556), .dina(n4873), .dout(n4877));
    jxor g1193(.dinb(n4861), .dina(n17119), .dout(n4881));
    jxor g1194(.dinb(n4825), .dina(n4881), .dout(n4885));
    jxor g1195(.dinb(n17115), .dina(n788), .dout(n4889));
    jxor g1196(.dinb(n709), .dina(n751), .dout(n4893));
    jxor g1197(.dinb(n17098), .dina(n4893), .dout(n4897));
    jxor g1198(.dinb(n4885), .dina(n4897), .dout(n4901));
    jand g1199(.dinb(n17166), .dina(n4901), .dout(n4905));
    jnot g1200(.din(n4905), .dout(n4908));
    jand g1201(.dinb(n4749), .dina(n17095), .dout(n4912));
    jor g1202(.dinb(n18123), .dina(n4912), .dout(n4916));
    jnot g1203(.din(n2003), .dout(n4919));
    jor g1204(.dinb(n15259), .dina(n4919), .dout(n4923));
    jand g1205(.dinb(n4916), .dina(n15250), .dout(n4927));
    jand g1206(.dinb(G248), .dina(G273), .dout(n4931));
    jand g1207(.dinb(n19554), .dina(n933), .dout(n4935));
    jor g1208(.dinb(n19570), .dina(n4935), .dout(n4939));
    jor g1209(.dinb(n19546), .dina(n4939), .dout(n4943));
    jand g1210(.dinb(n686), .dina(n933), .dout(n4947));
    jand g1211(.dinb(n693), .dina(n19605), .dout(n4951));
    jor g1212(.dinb(n4947), .dina(n4951), .dout(n4955));
    jor g1213(.dinb(n19593), .dina(n4955), .dout(n4959));
    jand g1214(.dinb(n4943), .dina(n4959), .dout(n4963));
    jand g1215(.dinb(G248), .dina(G281), .dout(n4967));
    jand g1216(.dinb(n19554), .dina(n1159), .dout(n4971));
    jor g1217(.dinb(n19486), .dina(n4971), .dout(n4975));
    jor g1218(.dinb(n19468), .dina(n4975), .dout(n4979));
    jand g1219(.dinb(n686), .dina(n1159), .dout(n4983));
    jand g1220(.dinb(n693), .dina(n19530), .dout(n4987));
    jor g1221(.dinb(n4983), .dina(n4987), .dout(n4991));
    jor g1222(.dinb(n19509), .dina(n4991), .dout(n4995));
    jand g1223(.dinb(n4979), .dina(n4995), .dout(n4999));
    jxor g1224(.dinb(n4963), .dina(n4999), .dout(n5003));
    jor g1225(.dinb(n548), .dina(n979), .dout(n5007));
    jor g1226(.dinb(n538), .dina(n19461), .dout(n5011));
    jand g1227(.dinb(n19440), .dina(n5011), .dout(n5015));
    jand g1228(.dinb(n19429), .dina(n5015), .dout(n5019));
    jor g1229(.dinb(G254), .dina(G265), .dout(n5023));
    jor g1230(.dinb(n19539), .dina(n979), .dout(n5027));
    jand g1231(.dinb(n19393), .dina(n5027), .dout(n5031));
    jand g1232(.dinb(n19401), .dina(n5031), .dout(n5035));
    jor g1233(.dinb(n5019), .dina(n5035), .dout(n5039));
    jand g1234(.dinb(G248), .dina(G257), .dout(n5043));
    jand g1235(.dinb(n19551), .dina(n1113), .dout(n5047));
    jor g1236(.dinb(n19345), .dina(n5047), .dout(n5051));
    jor g1237(.dinb(n19333), .dina(n5051), .dout(n5055));
    jand g1238(.dinb(n686), .dina(n1113), .dout(n5059));
    jand g1239(.dinb(n693), .dina(n19389), .dout(n5063));
    jor g1240(.dinb(n5059), .dina(n5063), .dout(n5067));
    jor g1241(.dinb(n19368), .dina(n5067), .dout(n5071));
    jand g1242(.dinb(n5055), .dina(n5071), .dout(n5075));
    jand g1243(.dinb(G234), .dina(G248), .dout(n5079));
    jand g1244(.dinb(n891), .dina(n19551), .dout(n5083));
    jor g1245(.dinb(n19282), .dina(n5083), .dout(n5087));
    jor g1246(.dinb(n19267), .dina(n5087), .dout(n5091));
    jand g1247(.dinb(n891), .dina(n686), .dout(n5095));
    jand g1248(.dinb(n19326), .dina(n693), .dout(n5099));
    jor g1249(.dinb(n5095), .dina(n5099), .dout(n5103));
    jor g1250(.dinb(n19305), .dina(n5103), .dout(n5107));
    jand g1251(.dinb(n5091), .dina(n5107), .dout(n5111));
    jxor g1252(.dinb(n5075), .dina(n5111), .dout(n5115));
    jxor g1253(.dinb(n19261), .dina(n5115), .dout(n5119));
    jxor g1254(.dinb(n19258), .dina(n5119), .dout(n5123));
    jand g1255(.dinb(G226), .dina(G248), .dout(n5127));
    jand g1256(.dinb(n1021), .dina(n19551), .dout(n5131));
    jor g1257(.dinb(n19174), .dina(n5131), .dout(n5135));
    jor g1258(.dinb(n19159), .dina(n5135), .dout(n5139));
    jand g1259(.dinb(n1021), .dina(n686), .dout(n5143));
    jand g1260(.dinb(n19206), .dina(n693), .dout(n5147));
    jor g1261(.dinb(n5143), .dina(n5147), .dout(n5151));
    jor g1262(.dinb(n19185), .dina(n5151), .dout(n5155));
    jand g1263(.dinb(n5139), .dina(n5155), .dout(n5159));
    jxor g1264(.dinb(n1240), .dina(n5159), .dout(n5163));
    jor g1265(.dinb(n1071), .dina(n548), .dout(n5167));
    jor g1266(.dinb(n19131), .dina(n538), .dout(n5171));
    jand g1267(.dinb(n19134), .dina(n5171), .dout(n5175));
    jand g1268(.dinb(n19129), .dina(n5175), .dout(n5179));
    jor g1269(.dinb(G218), .dina(G254), .dout(n5183));
    jor g1270(.dinb(n1071), .dina(n19536), .dout(n5187));
    jand g1271(.dinb(n19093), .dina(n5187), .dout(n5191));
    jand g1272(.dinb(n19095), .dina(n5191), .dout(n5195));
    jor g1273(.dinb(n5179), .dina(n5195), .dout(n5199));
    jand g1274(.dinb(G210), .dina(G248), .dout(n5203));
    jand g1275(.dinb(n849), .dina(n19437), .dout(n5207));
    jor g1276(.dinb(n19045), .dina(n5207), .dout(n5211));
    jor g1277(.dinb(n19033), .dina(n5211), .dout(n5215));
    jand g1278(.dinb(n849), .dina(n686), .dout(n5219));
    jand g1279(.dinb(n19089), .dina(n693), .dout(n5223));
    jor g1280(.dinb(n5219), .dina(n5223), .dout(n5227));
    jor g1281(.dinb(n19068), .dina(n5227), .dout(n5231));
    jand g1282(.dinb(n5215), .dina(n5231), .dout(n5235));
    jxor g1283(.dinb(n5199), .dina(n5235), .dout(n5239));
    jxor g1284(.dinb(n5163), .dina(n5239), .dout(n5243));
    jxor g1285(.dinb(n5123), .dina(n19027), .dout(n5247));
    jand g1286(.dinb(n19662), .dina(n5247), .dout(n5251));
    jnot g1287(.din(n5251), .dout(n5254));
    jand g1288(.dinb(n1301), .dina(n18966), .dout(n5258));
    jor g1289(.dinb(n1806), .dina(n18964), .dout(n5262));
    jnot g1290(.din(n1270), .dout(n5265));
    jor g1291(.dinb(n19002), .dina(n5265), .dout(n5269));
    jand g1292(.dinb(n19479), .dina(n5269), .dout(n5273));
    jnot g1293(.din(n5273), .dout(n5276));
    jor g1294(.dinb(n5276), .dina(n18978), .dout(n5280));
    jand g1295(.dinb(n19563), .dina(n2660), .dout(n5284));
    jor g1296(.dinb(n5273), .dina(n5284), .dout(n5288));
    jand g1297(.dinb(n5280), .dina(n18961), .dout(n5292));
    jxor g1298(.dinb(n5262), .dina(n18958), .dout(n5296));
    jnot g1299(.din(n5296), .dout(n5299));
    jnot g1300(.din(n1756), .dout(n5302));
    jnot g1301(.din(n1760), .dout(n5305));
    jor g1302(.dinb(n19473), .dina(n5269), .dout(n5309));
    jor g1303(.dinb(n5309), .dina(n5284), .dout(n5313));
    jor g1304(.dinb(n19557), .dina(n2660), .dout(n5317));
    jor g1305(.dinb(n19395), .dina(n1767), .dout(n5321));
    jand g1306(.dinb(n5317), .dina(n5321), .dout(n5325));
    jand g1307(.dinb(n5313), .dina(n5325), .dout(n5329));
    jor g1308(.dinb(n19005), .dina(n5329), .dout(n5333));
    jor g1309(.dinb(n18892), .dina(n5333), .dout(n5337));
    jand g1310(.dinb(n18886), .dina(n5337), .dout(n5341));
    jand g1311(.dinb(n18915), .dina(n5341), .dout(n5345));
    jxor g1312(.dinb(n1278), .dina(n1297), .dout(n5349));
    jxor g1313(.dinb(n2436), .dina(n5349), .dout(n5353));
    jxor g1314(.dinb(n5345), .dina(n18826), .dout(n5357));
    jnot g1315(.din(n5357), .dout(n5360));
    jand g1316(.dinb(n18814), .dina(n5360), .dout(n5364));
    jnot g1317(.din(G1497), .dout(n5367));
    jand g1318(.dinb(n18951), .dina(n5357), .dout(n5371));
    jor g1319(.dinb(n18727), .dina(n5371), .dout(n5375));
    jor g1320(.dinb(n5364), .dina(n5375), .dout(n5379));
    jand g1321(.dinb(n5309), .dina(n5317), .dout(n5383));
    jor g1322(.dinb(n1786), .dina(n5383), .dout(n5387));
    jxor g1323(.dinb(n5333), .dina(n18828), .dout(n5391));
    jxor g1324(.dinb(n18685), .dina(n5391), .dout(n5395));
    jxor g1325(.dinb(n18834), .dina(n5341), .dout(n5399));
    jxor g1326(.dinb(n18679), .dina(n5399), .dout(n5403));
    jor g1327(.dinb(n18774), .dina(n5403), .dout(n5407));
    jand g1328(.dinb(n5379), .dina(n18676), .dout(n5411));
    jxor g1329(.dinb(n1326), .dina(n18924), .dout(n5415));
    jxor g1330(.dinb(n5411), .dina(n18670), .dout(n5419));
    jnot g1331(.din(n1846), .dout(n5422));
    jand g1332(.dinb(n2772), .dina(n5422), .dout(n5426));
    jand g1333(.dinb(n2775), .dina(n18534), .dout(n5430));
    jor g1334(.dinb(n18562), .dina(n5430), .dout(n5434));
    jxor g1335(.dinb(n18510), .dina(n1456), .dout(n5438));
    jxor g1336(.dinb(n18531), .dina(n5438), .dout(n5442));
    jxor g1337(.dinb(n5434), .dina(n18469), .dout(n5446));
    jor g1338(.dinb(n18438), .dina(n2717), .dout(n5450));
    jand g1339(.dinb(n18361), .dina(n1460), .dout(n5454));
    jor g1340(.dinb(n1870), .dina(n18319), .dout(n5458));
    jand g1341(.dinb(n5450), .dina(n18316), .dout(n5462));
    jxor g1342(.dinb(n18313), .dina(n5462), .dout(n5466));
    jand g1343(.dinb(n18579), .dina(n5466), .dout(n5470));
    jnot g1344(.din(n1742), .dout(n5473));
    jor g1345(.dinb(n18597), .dina(n5341), .dout(n5477));
    jand g1346(.dinb(n18307), .dina(n5477), .dout(n5481));
    jand g1347(.dinb(n2775), .dina(n1862), .dout(n5485));
    jor g1348(.dinb(n18562), .dina(n5485), .dout(n5489));
    jxor g1349(.dinb(n2717), .dina(n18292), .dout(n5493));
    jxor g1350(.dinb(n18459), .dina(n5493), .dout(n5497));
    jand g1351(.dinb(n5481), .dina(n5497), .dout(n5501));
    jor g1352(.dinb(n5470), .dina(n18288), .dout(n5505));
    jor g1353(.dinb(n18729), .dina(n5505), .dout(n5509));
    jnot g1354(.din(n1379), .dout(n5512));
    jand g1355(.dinb(n18280), .dina(n5501), .dout(n5516));
    jor g1356(.dinb(n18282), .dina(n1822), .dout(n5520));
    jand g1357(.dinb(n5466), .dina(n5520), .dout(n5524));
    jor g1358(.dinb(n5516), .dina(n5524), .dout(n5528));
    jor g1359(.dinb(n18687), .dina(n5528), .dout(n5532));
    jand g1360(.dinb(n5509), .dina(n5532), .dout(n5536));
    jxor g1361(.dinb(n5419), .dina(n5536), .dout(n5540));
    jor g1362(.dinb(n19611), .dina(n5540), .dout(n5544));
    jand g1363(.dinb(n18274), .dina(n5544), .dout(n5548));
    jor g1364(.dinb(n19848), .dina(n5548), .dout(n5552));
    jor g1365(.dinb(n15319), .dina(n4919), .dout(n5556));
    jand g1366(.dinb(n5552), .dina(n15310), .dout(n5560));
    jor g1367(.dinb(G14), .dina(G4088), .dout(n5564));
    jor g1368(.dinb(n16111), .dina(n2178), .dout(n5568));
    jand g1369(.dinb(n15702), .dina(n5568), .dout(n5572));
    jand g1370(.dinb(n15607), .dina(n5572), .dout(n5576));
    jand g1371(.dinb(G97), .dina(G4092), .dout(n5580));
    jnot g1372(.din(n5580), .dout(n5583));
    jand g1373(.dinb(n5552), .dina(n18250), .dout(n5587));
    jnot g1374(.din(n5587), .dout(n5590));
    jor g1375(.dinb(n15609), .dina(n5590), .dout(n5594));
    jand g1376(.dinb(G94), .dina(G4092), .dout(n5598));
    jnot g1377(.din(n5598), .dout(n5601));
    jand g1378(.dinb(n4916), .dina(n17068), .dout(n5605));
    jnot g1379(.din(n5605), .dout(n5608));
    jor g1380(.dinb(n15717), .dina(n5608), .dout(n5612));
    jand g1381(.dinb(n15453), .dina(n5612), .dout(n5616));
    jand g1382(.dinb(n15451), .dina(n5616), .dout(n5620));
    jor g1383(.dinb(n15448), .dina(n5620), .dout(n5624));
    jor g1384(.dinb(G14), .dina(G4089), .dout(n5628));
    jor g1385(.dinb(n16111), .dina(n2387), .dout(n5632));
    jand g1386(.dinb(n16113), .dina(n5632), .dout(n5636));
    jand g1387(.dinb(n16015), .dina(n5636), .dout(n5640));
    jor g1388(.dinb(n16017), .dina(n5590), .dout(n5644));
    jor g1389(.dinb(n16128), .dina(n5608), .dout(n5648));
    jand g1390(.dinb(n15855), .dina(n5648), .dout(n5652));
    jand g1391(.dinb(n15853), .dina(n5652), .dout(n5656));
    jor g1392(.dinb(n15850), .dina(n5656), .dout(n5660));
    jnot g1393(.din(G137), .dout(n5663));
    jnot g1394(.din(G179), .dout(n5666));
    jnot g1395(.din(n2933), .dout(n5669));
    jor g1396(.dinb(n20554), .dina(n5669), .dout(n5673));
    jnot g1397(.din(G176), .dout(n5676));
    jnot g1398(.din(n2925), .dout(n5679));
    jor g1399(.dinb(n20227), .dina(n5679), .dout(n5683));
    jand g1400(.dinb(n16716), .dina(n5587), .dout(n5687));
    jand g1401(.dinb(n16407), .dina(n5605), .dout(n5691));
    jor g1402(.dinb(n16620), .dina(n5691), .dout(n5695));
    jor g1403(.dinb(n16330), .dina(n5695), .dout(n5699));
    jand g1404(.dinb(n16327), .dina(n5699), .dout(n5703));
    jand g1405(.dinb(n16264), .dina(n5703), .dout(n5707));
    jor g1406(.dinb(n20632), .dina(n5707), .dout(G658));
    jnot g1407(.din(n2994), .dout(n5714));
    jor g1408(.dinb(n20554), .dina(n5714), .dout(n5718));
    jnot g1409(.din(n3002), .dout(n5721));
    jor g1410(.dinb(n20227), .dina(n5721), .dout(n5725));
    jand g1411(.dinb(n20391), .dina(n5587), .dout(n5729));
    jand g1412(.dinb(n19986), .dina(n5605), .dout(n5733));
    jor g1413(.dinb(n20229), .dina(n5733), .dout(n5737));
    jor g1414(.dinb(n17011), .dina(n5737), .dout(n5741));
    jand g1415(.dinb(n17008), .dina(n5741), .dout(n5745));
    jand g1416(.dinb(n16945), .dina(n5745), .dout(n5749));
    jor g1417(.dinb(n20632), .dina(n5749), .dout(G690));
    jdff g1418(.din(G141), .dout(n5756));
    jdff g1419(.din(G293), .dout(n5759));
    jdff g1420(.din(G3173), .dout(n5762));
    jnot g1421(.din(G545), .dout(n5765));
    jnot g1422(.din(G545), .dout(n5768));
    jdff g1423(.din(G137), .dout(n5771));
    jdff g1424(.din(G141), .dout(n5774));
    jdff g1425(.din(G1), .dout(n5777));
    jdff g1426(.din(G549), .dout(n5780));
    jdff g1427(.din(G299), .dout(n5783));
    jnot g1428(.din(G549), .dout(n5786));
    jdff g1429(.din(G1), .dout(n5789));
    jdff g1430(.din(G1), .dout(n5792));
    jdff g1431(.din(G1), .dout(n5795));
    jdff g1432(.din(G1), .dout(n5798));
    jdff g1433(.din(G299), .dout(n5801));
    jor g1434(.dinb(n8413), .dina(n423), .dout(n5805));
    jand g1435(.dinb(n1583), .dina(n8515), .dout(n5809));
    jand g1436(.dinb(n1379), .dina(n8563), .dout(n5813));
    jor g1437(.dinb(n1826), .dina(n8521), .dout(n5817));
    jor g1438(.dinb(n1960), .dina(n8569), .dout(n5821));
    jdff dff_A_Y9j4iuZu8_2(.din(n5660), .dout(G807));
    jdff dff_A_uayLeJHg8_2(.din(n5624), .dout(G767));
    jdff dff_A_Z6lxaLEo3_0(.din(n26589), .dout(G882));
    jdff dff_A_KtDh1uLu6_0(.din(n26586), .dout(n26589));
    jdff dff_A_o0pkMQJ63_0(.din(n26583), .dout(n26586));
    jdff dff_A_z297T3Oe8_0(.din(n26580), .dout(n26583));
    jdff dff_A_0DNiYuTX8_0(.din(n26577), .dout(n26580));
    jdff dff_A_d5yH2TQb2_2(.din(n5560), .dout(n26577));
    jdff dff_A_qhYBnWPj1_0(.din(n26571), .dout(G843));
    jdff dff_A_RaE1t2gH7_0(.din(n26568), .dout(n26571));
    jdff dff_A_cmeWtwhA1_0(.din(n26565), .dout(n26568));
    jdff dff_A_sTH0gPWI1_0(.din(n26562), .dout(n26565));
    jdff dff_A_LzkmumMs1_0(.din(n26559), .dout(n26562));
    jdff dff_A_EMPb80Xy4_2(.din(n4927), .dout(n26559));
    jdff dff_A_LMlsjDrx1_0(.din(n26553), .dout(G688));
    jdff dff_A_5Kjw3Tkd6_0(.din(n26550), .dout(n26553));
    jdff dff_A_et8vM2y52_2(.din(n4538), .dout(n26550));
    jdff dff_A_Bbj03Fq73_0(.din(n26544), .dout(G685));
    jdff dff_A_Kib1mxWx5_0(.din(n26541), .dout(n26544));
    jdff dff_A_BvotNGEA0_2(.din(n4502), .dout(n26541));
    jdff dff_A_Agly4Fzj9_0(.din(n26535), .dout(G682));
    jdff dff_A_gBeoBIe98_0(.din(n26532), .dout(n26535));
    jdff dff_A_EU9AjEys6_2(.din(n4466), .dout(n26532));
    jdff dff_A_FsMUJCpF2_0(.din(n26526), .dout(G679));
    jdff dff_A_XYb04rwh0_0(.din(n26523), .dout(n26526));
    jdff dff_A_lkCp01sO9_0(.din(n26520), .dout(n26523));
    jdff dff_A_JhrkJhl39_2(.din(n4430), .dout(n26520));
    jdff dff_A_iFsWFNfO5_0(.din(n26514), .dout(G654));
    jdff dff_A_W8e3w3NF5_2(.din(n4394), .dout(n26514));
    jdff dff_A_hEQsiTAf9_0(.din(n26508), .dout(G651));
    jdff dff_A_q80xYIbs9_0(.din(n26505), .dout(n26508));
    jdff dff_A_8Et3bTWw1_2(.din(n4358), .dout(n26505));
    jdff dff_A_xk7Cz47b9_0(.din(n26499), .dout(G648));
    jdff dff_A_lCoSCkNt9_0(.din(n26496), .dout(n26499));
    jdff dff_A_2tJJd17T5_2(.din(n4322), .dout(n26496));
    jdff dff_A_qSB0BDZw9_0(.din(n26490), .dout(G645));
    jdff dff_A_44bWtlZI3_0(.din(n26487), .dout(n26490));
    jdff dff_A_lQAtOq602_0(.din(n26484), .dout(n26487));
    jdff dff_A_iUpifcdH2_2(.din(n4286), .dout(n26484));
    jdff dff_A_xSGnrJLD0_0(.din(n26478), .dout(G782));
    jdff dff_A_p0FFlBzA3_0(.din(n26475), .dout(n26478));
    jdff dff_A_tvjJ54RO0_0(.din(n26472), .dout(n26475));
    jdff dff_A_L4953zrj5_0(.din(n26469), .dout(n26472));
    jdff dff_A_8lfa568n2_2(.din(n4250), .dout(n26469));
    jdff dff_A_lnSRuheC9_0(.din(n26463), .dout(G777));
    jdff dff_A_elfhUkaj9_0(.din(n26460), .dout(n26463));
    jdff dff_A_c6sjhufo6_0(.din(n26457), .dout(n26460));
    jdff dff_A_iVlpqlh74_2(.din(n4214), .dout(n26457));
    jdff dff_A_6IPccs4l1_0(.din(n26451), .dout(G772));
    jdff dff_A_pycDjWzk1_0(.din(n26448), .dout(n26451));
    jdff dff_A_mukuAoNM5_0(.din(n26445), .dout(n26448));
    jdff dff_A_YNkz6Tgg6_2(.din(n4178), .dout(n26445));
    jdff dff_A_ur4sohGn4_0(.din(n26439), .dout(G742));
    jdff dff_A_jXQAFSfX9_0(.din(n26436), .dout(n26439));
    jdff dff_A_u4CHBI0j2_0(.din(n26433), .dout(n26436));
    jdff dff_A_6DDb7pdb3_0(.din(n26430), .dout(n26433));
    jdff dff_A_LJKa69Qm9_2(.din(n4142), .dout(n26430));
    jdff dff_A_cfobi81r2_0(.din(n26424), .dout(G737));
    jdff dff_A_UsCiql2t9_0(.din(n26421), .dout(n26424));
    jdff dff_A_nwSLAHCZ1_0(.din(n26418), .dout(n26421));
    jdff dff_A_UFCuDxvQ5_2(.din(n4100), .dout(n26418));
    jdff dff_A_ejDAC4ma8_0(.din(n26412), .dout(G732));
    jdff dff_A_oJAdkQg52_0(.din(n26409), .dout(n26412));
    jdff dff_A_wmaiJ6M16_0(.din(n26406), .dout(n26409));
    jdff dff_A_1o2NTLEO3_2(.din(n4064), .dout(n26406));
    jdff dff_A_dizJkHxB8_0(.din(n26400), .dout(G727));
    jdff dff_A_HVf0SUn03_0(.din(n26397), .dout(n26400));
    jdff dff_A_9ZseDTY54_2(.din(n4025), .dout(n26397));
    jdff dff_A_0LeTCrT14_0(.din(n26391), .dout(G712));
    jdff dff_A_WpWKO3K38_0(.din(n26388), .dout(n26391));
    jdff dff_A_8Vbysi9b2_0(.din(n26385), .dout(n26388));
    jdff dff_A_9sxuK1rx0_2(.din(n3989), .dout(n26385));
    jdff dff_A_UA3c6uSj0_0(.din(n26379), .dout(G869));
    jdff dff_A_aSH3WLwF9_0(.din(n26376), .dout(n26379));
    jdff dff_A_oERts3xA4_0(.din(n26373), .dout(n26376));
    jdff dff_A_TOixvbg22_0(.din(n26370), .dout(n26373));
    jdff dff_A_eJneS3RH0_0(.din(n26367), .dout(n26370));
    jdff dff_A_2mUDQUYi4_0(.din(n26364), .dout(n26367));
    jdff dff_A_eopy3nFu1_0(.din(n26361), .dout(n26364));
    jdff dff_A_lEjOuwSH1_0(.din(n26358), .dout(n26361));
    jdff dff_A_nr5st40n4_0(.din(n26355), .dout(n26358));
    jdff dff_A_YxXv40kT5_1(.din(n3953), .dout(n26355));
    jdff dff_A_N2KlKkZ48_0(.din(n26349), .dout(G867));
    jdff dff_A_NGxlt3pd2_0(.din(n26346), .dout(n26349));
    jdff dff_A_tNXXiEgG1_0(.din(n26343), .dout(n26346));
    jdff dff_A_g4zNuHiz0_0(.din(n26340), .dout(n26343));
    jdff dff_A_H5JPP1089_0(.din(n26337), .dout(n26340));
    jdff dff_A_pllF5Uob6_0(.din(n26334), .dout(n26337));
    jdff dff_A_ybOm80nJ7_1(.din(n3926), .dout(n26334));
    jdff dff_A_T9EiKK7U8_0(.din(n26328), .dout(G865));
    jdff dff_A_N9gBLWNS1_0(.din(n26325), .dout(n26328));
    jdff dff_A_qwXK7NWB1_0(.din(n26322), .dout(n26325));
    jdff dff_A_8y39fQ1n8_0(.din(n26319), .dout(n26322));
    jdff dff_A_JKwEgMNF6_0(.din(n26316), .dout(n26319));
    jdff dff_A_ndgumlmq8_0(.din(n26313), .dout(n26316));
    jdff dff_A_RMCiEWdP1_0(.din(n26310), .dout(n26313));
    jdff dff_A_XHwCdkcM9_0(.din(n26307), .dout(n26310));
    jdff dff_A_8HK7cpkl2_1(.din(n3896), .dout(n26307));
    jdff dff_A_XuaPGdcM1_0(.din(n26301), .dout(G863));
    jdff dff_A_TZKGaMGi8_0(.din(n26298), .dout(n26301));
    jdff dff_A_ovPhs7Em2_0(.din(n26295), .dout(n26298));
    jdff dff_A_qq8TKOja5_0(.din(n26292), .dout(n26295));
    jdff dff_A_VL4u1syn8_0(.din(n26289), .dout(n26292));
    jdff dff_A_6KcRPZEY1_1(.din(n3869), .dout(n26289));
    jdff dff_A_HT2ozZiF6_0(.din(n26283), .dout(G854));
    jdff dff_A_Pop8U8747_0(.din(n26280), .dout(n26283));
    jdff dff_A_9g95h1Z50_0(.din(n26277), .dout(n26280));
    jdff dff_A_7qxCi5Hh4_0(.din(n26274), .dout(n26277));
    jdff dff_A_0OuHfazO0_0(.din(n26271), .dout(n26274));
    jdff dff_A_JgKoGoOG6_0(.din(n26268), .dout(n26271));
    jdff dff_A_GcND7V5D3_0(.din(n26265), .dout(n26268));
    jdff dff_A_K4j0spcf0_0(.din(n26262), .dout(n26265));
    jdff dff_A_NqzCJA5O3_0(.din(n26259), .dout(n26262));
    jdff dff_A_8JSSzpdP3_0(.din(n26256), .dout(n26259));
    jdff dff_A_XJybgXKZ4_0(.din(n26253), .dout(n26256));
    jdff dff_A_64wp8i3q5_0(.din(n26250), .dout(n26253));
    jdff dff_A_ofDz5DV79_0(.din(n26247), .dout(n26250));
    jdff dff_A_onCEKMEY6_0(.din(n26244), .dout(n26247));
    jdff dff_A_wAm89jr86_0(.din(n26241), .dout(n26244));
    jdff dff_A_iYY8G84B7_0(.din(n26238), .dout(n26241));
    jdff dff_A_895FGv130_2(.din(n3839), .dout(n26238));
    jdff dff_A_bVfZZB9E3_0(.din(n26232), .dout(G830));
    jdff dff_A_ElkFPYjj3_0(.din(n26229), .dout(n26232));
    jdff dff_A_jRoTd1a24_0(.din(n26226), .dout(n26229));
    jdff dff_A_rrEDsG667_0(.din(n26223), .dout(n26226));
    jdff dff_A_3NYxN2fx2_0(.din(n26220), .dout(n26223));
    jdff dff_A_sJPm82kd9_0(.din(n26217), .dout(n26220));
    jdff dff_A_HT0lfgmT0_0(.din(n26214), .dout(n26217));
    jdff dff_A_SdQ38IQz7_0(.din(n26211), .dout(n26214));
    jdff dff_A_602QKs9Q0_0(.din(n26208), .dout(n26211));
    jdff dff_A_4oM9h1By1_0(.din(n26205), .dout(n26208));
    jdff dff_A_gSlZSXwH6_0(.din(n26202), .dout(n26205));
    jdff dff_A_lO1QpRnm5_1(.din(n3808), .dout(n26202));
    jdff dff_A_PC2vSuin3_0(.din(n26196), .dout(G828));
    jdff dff_A_MdeDkIKL4_0(.din(n26193), .dout(n26196));
    jdff dff_A_hm9aLquT5_0(.din(n26190), .dout(n26193));
    jdff dff_A_BP2h6ADM8_0(.din(n26187), .dout(n26190));
    jdff dff_A_U3tmic7N8_0(.din(n26184), .dout(n26187));
    jdff dff_A_2JoAGth54_0(.din(n26181), .dout(n26184));
    jdff dff_A_EMYGxBMS3_1(.din(n3781), .dout(n26181));
    jdff dff_A_U2IuuViG0_0(.din(n26175), .dout(G826));
    jdff dff_A_JlobzhOr4_0(.din(n26172), .dout(n26175));
    jdff dff_A_QVQFkG3y9_0(.din(n26169), .dout(n26172));
    jdff dff_A_MqXftXCi9_0(.din(n26166), .dout(n26169));
    jdff dff_A_K8ITLv3f5_0(.din(n26163), .dout(n26166));
    jdff dff_A_KFbpGayW2_0(.din(n26160), .dout(n26163));
    jdff dff_A_XBmdcbDl4_0(.din(n26157), .dout(n26160));
    jdff dff_A_BfQNuq0O6_1(.din(n3751), .dout(n26157));
    jdff dff_A_gHpjmiQs1_0(.din(n26151), .dout(G824));
    jdff dff_A_mHR4cvL27_0(.din(n26148), .dout(n26151));
    jdff dff_A_0i01aeYu0_0(.din(n26145), .dout(n26148));
    jdff dff_A_IbKSO0nV9_0(.din(n26142), .dout(n26145));
    jdff dff_A_3J3C8zlF7_0(.din(n26139), .dout(n26142));
    jdff dff_A_XteXsbNS7_0(.din(n26136), .dout(n26139));
    jdff dff_A_JP0ztOG01_1(.din(n3718), .dout(n26136));
    jdff dff_A_uaOdc2z75_0(.din(n26130), .dout(G813));
    jdff dff_A_61roVGaG6_0(.din(n26127), .dout(n26130));
    jdff dff_A_pkJbzM3e8_0(.din(n26124), .dout(n26127));
    jdff dff_A_ARy93q053_0(.din(n26121), .dout(n26124));
    jdff dff_A_rNDqtyMM3_0(.din(n26118), .dout(n26121));
    jdff dff_A_DsKGo98l7_0(.din(n26115), .dout(n26118));
    jdff dff_A_WdVzl2oX6_0(.din(n26112), .dout(n26115));
    jdff dff_A_nktSdCDh8_0(.din(n26109), .dout(n26112));
    jdff dff_A_ipkVkOPj4_0(.din(n26106), .dout(n26109));
    jdff dff_A_yfUFm8z19_2(.din(n3688), .dout(n26106));
    jdff dff_A_8ZQBge4d2_0(.din(n26100), .dout(G818));
    jdff dff_A_tsj9VRhx1_0(.din(n26097), .dout(n26100));
    jdff dff_A_VnZF5srs2_0(.din(n26094), .dout(n26097));
    jdff dff_A_d1AauKi04_0(.din(n26091), .dout(n26094));
    jdff dff_A_d0mWpsIG6_0(.din(n26088), .dout(n26091));
    jdff dff_A_go1YCpUD8_0(.din(n26085), .dout(n26088));
    jdff dff_A_6D6rviAx0_2(.din(n3684), .dout(n26085));
    jdff dff_A_ubA97bsl7_0(.din(n26079), .dout(G702));
    jdff dff_A_tuWa77KN8_0(.din(n26076), .dout(n26079));
    jdff dff_A_n5ZA8VPH5_0(.din(n26073), .dout(n26076));
    jdff dff_A_xScfjUXN6_0(.din(n26070), .dout(n26073));
    jdff dff_A_MG9fIiLi9_0(.din(n26067), .dout(n26070));
    jdff dff_A_p98PBW9Q3_0(.din(n26064), .dout(n26067));
    jdff dff_A_6gwONjtW0_0(.din(n26061), .dout(n26064));
    jdff dff_A_nUEvxDSH5_0(.din(n26058), .dout(n26061));
    jdff dff_A_gyEHSMrf9_2(.din(n3618), .dout(n26058));
    jdff dff_A_CF9Du5FX7_0(.din(n26052), .dout(G699));
    jdff dff_A_YuQ5v5OO5_0(.din(n26049), .dout(n26052));
    jdff dff_A_Pe7egUoa6_0(.din(n26046), .dout(n26049));
    jdff dff_A_aFDQzf0f6_0(.din(n26043), .dout(n26046));
    jdff dff_A_OXHogqZl0_0(.din(n26040), .dout(n26043));
    jdff dff_A_u7lIUA0f9_0(.din(n26037), .dout(n26040));
    jdff dff_A_jMVx26Eo7_0(.din(n26034), .dout(n26037));
    jdff dff_A_jRRsxoCY2_0(.din(n26031), .dout(n26034));
    jdff dff_A_DeXEoGm77_0(.din(n26028), .dout(n26031));
    jdff dff_A_2N0KkA108_2(.din(n3582), .dout(n26028));
    jdff dff_A_P5M5q3K66_0(.din(n26022), .dout(G696));
    jdff dff_A_3TeE7m7O3_0(.din(n26019), .dout(n26022));
    jdff dff_A_OjxKfTJd9_0(.din(n26016), .dout(n26019));
    jdff dff_A_Otgs3z9w2_0(.din(n26013), .dout(n26016));
    jdff dff_A_VbV0U5Qh2_0(.din(n26010), .dout(n26013));
    jdff dff_A_ZR5Hs4fi9_0(.din(n26007), .dout(n26010));
    jdff dff_A_9gxXs9RW4_0(.din(n26004), .dout(n26007));
    jdff dff_A_ABvZrmUz6_0(.din(n26001), .dout(n26004));
    jdff dff_A_z29pUF2q2_0(.din(n25998), .dout(n26001));
    jdff dff_A_8eEJ4Fst4_2(.din(n3546), .dout(n25998));
    jdff dff_A_jCghNv7G4_0(.din(n25992), .dout(G676));
    jdff dff_A_hYM606gy2_0(.din(n25989), .dout(n25992));
    jdff dff_A_JvJfqCJj5_0(.din(n25986), .dout(n25989));
    jdff dff_A_fCCOpQyt7_0(.din(n25983), .dout(n25986));
    jdff dff_A_qr71TKgs6_0(.din(n25980), .dout(n25983));
    jdff dff_A_GYTpg0iA4_2(.din(n3510), .dout(n25980));
    jdff dff_A_uS2qjpmo0_0(.din(n25974), .dout(G670));
    jdff dff_A_T75FYnvw5_0(.din(n25971), .dout(n25974));
    jdff dff_A_lEPF0NfB0_0(.din(n25968), .dout(n25971));
    jdff dff_A_J7X7YSBc0_0(.din(n25965), .dout(n25968));
    jdff dff_A_CWFexcX38_0(.din(n25962), .dout(n25965));
    jdff dff_A_MSnstR2G4_0(.din(n25959), .dout(n25962));
    jdff dff_A_StUcGH4c1_0(.din(n25956), .dout(n25959));
    jdff dff_A_4QyUmgVw0_0(.din(n25953), .dout(n25956));
    jdff dff_A_IObyZMPk5_2(.din(n3474), .dout(n25953));
    jdff dff_A_11QVwRVB7_0(.din(n25947), .dout(G667));
    jdff dff_A_TRamPBMB1_0(.din(n25944), .dout(n25947));
    jdff dff_A_ucfcjsAp5_0(.din(n25941), .dout(n25944));
    jdff dff_A_bUP0NYwP1_0(.din(n25938), .dout(n25941));
    jdff dff_A_ceJUF5kM6_0(.din(n25935), .dout(n25938));
    jdff dff_A_YHclVrpf8_0(.din(n25932), .dout(n25935));
    jdff dff_A_neo7xxPE8_0(.din(n25929), .dout(n25932));
    jdff dff_A_vejniamN9_0(.din(n25926), .dout(n25929));
    jdff dff_A_udKfIzWQ4_0(.din(n25923), .dout(n25926));
    jdff dff_A_hZ4sVGkq1_2(.din(n3438), .dout(n25923));
    jdff dff_A_cytpHSzO3_0(.din(n25917), .dout(G664));
    jdff dff_A_65IWDiCl7_0(.din(n25914), .dout(n25917));
    jdff dff_A_yyGcsfkC2_0(.din(n25911), .dout(n25914));
    jdff dff_A_LoHZeWOW8_0(.din(n25908), .dout(n25911));
    jdff dff_A_MjXwIlmF3_0(.din(n25905), .dout(n25908));
    jdff dff_A_5YXDiOFk2_0(.din(n25902), .dout(n25905));
    jdff dff_A_LYkqClVd5_0(.din(n25899), .dout(n25902));
    jdff dff_A_eKQkdrWr5_0(.din(n25896), .dout(n25899));
    jdff dff_A_8c1TUqnO7_0(.din(n25893), .dout(n25896));
    jdff dff_A_kmX7ykt16_2(.din(n3402), .dout(n25893));
    jdff dff_A_h9veY0Y49_0(.din(n25887), .dout(G642));
    jdff dff_A_zry6GCFm8_0(.din(n25884), .dout(n25887));
    jdff dff_A_9pnHBrWs3_0(.din(n25881), .dout(n25884));
    jdff dff_A_UZ72JWAY2_0(.din(n25878), .dout(n25881));
    jdff dff_A_yLTkF0KQ9_0(.din(n25875), .dout(n25878));
    jdff dff_A_AFy31fML3_0(.din(n25872), .dout(n25875));
    jdff dff_A_oXtvQCRh0_2(.din(n3366), .dout(n25872));
    jdff dff_A_QVX67lTB4_0(.din(n25866), .dout(G802));
    jdff dff_A_AoKy7gAF3_0(.din(n25863), .dout(n25866));
    jdff dff_A_atVMBKUE6_0(.din(n25860), .dout(n25863));
    jdff dff_A_CBOLz7UP0_0(.din(n25857), .dout(n25860));
    jdff dff_A_H6Wft9bg2_0(.din(n25854), .dout(n25857));
    jdff dff_A_oG3gG4hH5_0(.din(n25851), .dout(n25854));
    jdff dff_A_53MU5xUe5_0(.din(n25848), .dout(n25851));
    jdff dff_A_LlrZNhX42_0(.din(n25845), .dout(n25848));
    jdff dff_A_zfoHNcgE4_0(.din(n25842), .dout(n25845));
    jdff dff_A_Oq5Agr8v8_2(.din(n3330), .dout(n25842));
    jdff dff_A_qu9L4y1s5_0(.din(n25836), .dout(G797));
    jdff dff_A_zrmWGPMr4_0(.din(n25833), .dout(n25836));
    jdff dff_A_Zr4QqwU15_0(.din(n25830), .dout(n25833));
    jdff dff_A_eq05BWI14_0(.din(n25827), .dout(n25830));
    jdff dff_A_ylGy2fok4_0(.din(n25824), .dout(n25827));
    jdff dff_A_IS7AgNOe9_0(.din(n25821), .dout(n25824));
    jdff dff_A_5orXmOyV5_0(.din(n25818), .dout(n25821));
    jdff dff_A_uWF7OVIf0_0(.din(n25815), .dout(n25818));
    jdff dff_A_PmQtesJW5_0(.din(n25812), .dout(n25815));
    jdff dff_A_M3DLpiA72_0(.din(n25809), .dout(n25812));
    jdff dff_A_JuenzXYu0_2(.din(n3294), .dout(n25809));
    jdff dff_A_R7He8G2k5_0(.din(n25803), .dout(G792));
    jdff dff_A_XcBEXdFK7_0(.din(n25800), .dout(n25803));
    jdff dff_A_LBw97b4V0_0(.din(n25797), .dout(n25800));
    jdff dff_A_8PdqdZtj4_0(.din(n25794), .dout(n25797));
    jdff dff_A_FOVkeETD8_0(.din(n25791), .dout(n25794));
    jdff dff_A_WRvWehwM1_0(.din(n25788), .dout(n25791));
    jdff dff_A_I6U6F1X47_0(.din(n25785), .dout(n25788));
    jdff dff_A_AhJMBAbg8_0(.din(n25782), .dout(n25785));
    jdff dff_A_AdHQiQye7_2(.din(n3258), .dout(n25782));
    jdff dff_A_5kDxmMZn0_0(.din(n25776), .dout(G787));
    jdff dff_A_8AryYicP2_0(.din(n25773), .dout(n25776));
    jdff dff_A_07LDldsB9_0(.din(n25770), .dout(n25773));
    jdff dff_A_utjEpEXv7_0(.din(n25767), .dout(n25770));
    jdff dff_A_guSCZ5V70_0(.din(n25764), .dout(n25767));
    jdff dff_A_3CMRcvsG8_0(.din(n25761), .dout(n25764));
    jdff dff_A_Sz9vAu1E6_0(.din(n25758), .dout(n25761));
    jdff dff_A_Zo2KDTfC2_2(.din(n3222), .dout(n25758));
    jdff dff_A_7YUUNSrQ2_0(.din(n25752), .dout(G762));
    jdff dff_A_kXSjycLt2_0(.din(n25749), .dout(n25752));
    jdff dff_A_titBxf2B9_0(.din(n25746), .dout(n25749));
    jdff dff_A_qg0TwOd41_0(.din(n25743), .dout(n25746));
    jdff dff_A_wydLsCJt6_0(.din(n25740), .dout(n25743));
    jdff dff_A_SGB4ZzDu8_0(.din(n25737), .dout(n25740));
    jdff dff_A_TvWaKho87_0(.din(n25734), .dout(n25737));
    jdff dff_A_0vWcoYRv3_0(.din(n25731), .dout(n25734));
    jdff dff_A_5DTFfIwR9_0(.din(n25728), .dout(n25731));
    jdff dff_A_esKhrEUJ8_2(.din(n3186), .dout(n25728));
    jdff dff_A_a8Qk4bxx1_0(.din(n25722), .dout(G757));
    jdff dff_A_FePXc5eJ4_0(.din(n25719), .dout(n25722));
    jdff dff_A_2Rc8y7wi0_0(.din(n25716), .dout(n25719));
    jdff dff_A_kB58hnys1_0(.din(n25713), .dout(n25716));
    jdff dff_A_Evi6oj1V5_0(.din(n25710), .dout(n25713));
    jdff dff_A_iB2f7KVS4_0(.din(n25707), .dout(n25710));
    jdff dff_A_pxTGSbKb4_0(.din(n25704), .dout(n25707));
    jdff dff_A_IvKZmHXa9_0(.din(n25701), .dout(n25704));
    jdff dff_A_TwTHJyww3_0(.din(n25698), .dout(n25701));
    jdff dff_A_AiUgCs3j2_0(.din(n25695), .dout(n25698));
    jdff dff_A_7if5Ex0z2_2(.din(n3144), .dout(n25695));
    jdff dff_A_gvDaQNL11_0(.din(n25689), .dout(G752));
    jdff dff_A_7d2cgz226_0(.din(n25686), .dout(n25689));
    jdff dff_A_alPBq42p3_0(.din(n25683), .dout(n25686));
    jdff dff_A_oa1i2zPk6_0(.din(n25680), .dout(n25683));
    jdff dff_A_hgH6Jr8k8_0(.din(n25677), .dout(n25680));
    jdff dff_A_LN3kr5iU5_0(.din(n25674), .dout(n25677));
    jdff dff_A_gsqUxdvN0_0(.din(n25671), .dout(n25674));
    jdff dff_A_Y6zRAHiT2_0(.din(n25668), .dout(n25671));
    jdff dff_A_nBX0wvip1_2(.din(n3102), .dout(n25668));
    jdff dff_A_chlM9X4k7_0(.din(n25662), .dout(G747));
    jdff dff_A_kFWA9HyF6_0(.din(n25659), .dout(n25662));
    jdff dff_A_h1qgAggJ6_0(.din(n25656), .dout(n25659));
    jdff dff_A_ppKmVk3i2_0(.din(n25653), .dout(n25656));
    jdff dff_A_EW1wDWNf1_0(.din(n25650), .dout(n25653));
    jdff dff_A_HHLtTfzI9_0(.din(n25647), .dout(n25650));
    jdff dff_A_DWhri1bT0_0(.din(n25644), .dout(n25647));
    jdff dff_A_GBVcLEQV9_2(.din(n3060), .dout(n25644));
    jdff dff_A_iBAJdm7G7_0(.din(n25638), .dout(G693));
    jdff dff_A_9U9Fyhuk2_0(.din(n25635), .dout(n25638));
    jdff dff_A_W8lInqRb8_0(.din(n25632), .dout(n25635));
    jdff dff_A_nuMBE6R39_0(.din(n25629), .dout(n25632));
    jdff dff_A_DzCJnUyy5_0(.din(n25626), .dout(n25629));
    jdff dff_A_IdYvVSNC8_0(.din(n25623), .dout(n25626));
    jdff dff_A_Rjm9jPqe8_0(.din(n25620), .dout(n25623));
    jdff dff_A_qbl5jmXt5_0(.din(n25617), .dout(n25620));
    jdff dff_A_66JR4QGx3_0(.din(n25614), .dout(n25617));
    jdff dff_A_8kfcHEHr0_0(.din(n25611), .dout(n25614));
    jdff dff_A_xvOKcKuY6_0(.din(n25608), .dout(n25611));
    jdff dff_A_7W4GWUDP1_2(.din(n3018), .dout(n25608));
    jdff dff_A_oMrIBUE60_0(.din(n25602), .dout(G661));
    jdff dff_A_pSp5ibAu8_0(.din(n25599), .dout(n25602));
    jdff dff_A_0KlY1cIq4_0(.din(n25596), .dout(n25599));
    jdff dff_A_pekoyJtn2_0(.din(n25593), .dout(n25596));
    jdff dff_A_ioNsIhzp4_0(.din(n25590), .dout(n25593));
    jdff dff_A_NNzvW05A4_0(.din(n25587), .dout(n25590));
    jdff dff_A_JIkxsbV44_0(.din(n25584), .dout(n25587));
    jdff dff_A_y9XzhXBi3_0(.din(n25581), .dout(n25584));
    jdff dff_A_0ZF7D4nz8_0(.din(n25578), .dout(n25581));
    jdff dff_A_6ish0ona2_0(.din(n25575), .dout(n25578));
    jdff dff_A_aoyZcCuj3_0(.din(n25572), .dout(n25575));
    jdff dff_A_cgdxqHwN3_2(.din(n2968), .dout(n25572));
    jdff dff_A_pmWRA6JS0_0(.din(n25566), .dout(G585));
    jdff dff_A_csXTs7Yw4_0(.din(n25563), .dout(n25566));
    jdff dff_A_26apLcSj0_0(.din(n25560), .dout(n25563));
    jdff dff_A_pLEqq7yX9_0(.din(n25557), .dout(n25560));
    jdff dff_A_01GTjzFh5_0(.din(n25554), .dout(n25557));
    jdff dff_A_ickgKFvR1_0(.din(n25551), .dout(n25554));
    jdff dff_A_RJ18dgvy4_2(.din(n2918), .dout(n25551));
    jdff dff_A_LVK68FTZ8_0(.din(n25545), .dout(G575));
    jdff dff_A_5Wi4odPO4_0(.din(n25542), .dout(n25545));
    jdff dff_A_qm8ipQwt3_0(.din(n25539), .dout(n25542));
    jdff dff_A_mIlpv17y8_0(.din(n25536), .dout(n25539));
    jdff dff_A_N39xu8ts0_0(.din(n25533), .dout(n25536));
    jdff dff_A_wUORH9CY2_0(.din(n25530), .dout(n25533));
    jdff dff_A_qiNPFECI1_0(.din(n25527), .dout(n25530));
    jdff dff_A_WTTfnauU2_2(.din(n2828), .dout(n25527));
    jdff dff_A_micxCBgF9_0(.din(n25521), .dout(G1000));
    jdff dff_A_6WPFaNR41_0(.din(n25518), .dout(n25521));
    jdff dff_A_Qcn33iHW0_0(.din(n25515), .dout(n25518));
    jdff dff_A_mAjVlnfA4_0(.din(n25512), .dout(n25515));
    jdff dff_A_WQgKZmDb2_0(.din(n25509), .dout(n25512));
    jdff dff_A_WklZoigz0_0(.din(n25506), .dout(n25509));
    jdff dff_A_fxiYAWL33_0(.din(n25503), .dout(n25506));
    jdff dff_A_6Opw3FZL5_0(.din(n25500), .dout(n25503));
    jdff dff_A_wW4156Sl2_0(.din(n25497), .dout(n25500));
    jdff dff_A_hK9kiUZD7_0(.din(n25494), .dout(n25497));
    jdff dff_A_FSZwXZ276_0(.din(n25491), .dout(n25494));
    jdff dff_A_16vCrZbw8_0(.din(n25488), .dout(n25491));
    jdff dff_A_6ZUh4y4v1_0(.din(n25485), .dout(n25488));
    jdff dff_A_JWwDsi4h2_0(.din(n25482), .dout(n25485));
    jdff dff_A_ZERoUCzr9_0(.din(n25479), .dout(n25482));
    jdff dff_A_7yPlVLkp1_0(.din(n25476), .dout(n25479));
    jdff dff_A_ryLxFFBv7_0(.din(n25473), .dout(n25476));
    jdff dff_A_nTfjI0cF2_0(.din(n25470), .dout(n25473));
    jdff dff_A_DX0Mtc6R2_1(.din(n2711), .dout(n25470));
    jdff dff_A_cLd5Q0cP9_0(.din(n25464), .dout(G998));
    jdff dff_A_csnrMbGv0_0(.din(n25461), .dout(n25464));
    jdff dff_A_cLzWTcj00_0(.din(n25458), .dout(n25461));
    jdff dff_A_xvWGgnOV7_0(.din(n25455), .dout(n25458));
    jdff dff_A_aIQslsMW3_0(.din(n25452), .dout(n25455));
    jdff dff_A_Tz4jAXf56_0(.din(n25449), .dout(n25452));
    jdff dff_A_onUMXk6V9_0(.din(n25446), .dout(n25449));
    jdff dff_A_dpReoaM02_0(.din(n25443), .dout(n25446));
    jdff dff_A_Z7PbR7z03_0(.din(n25440), .dout(n25443));
    jdff dff_A_ES9gYQ6i5_0(.din(n25437), .dout(n25440));
    jdff dff_A_ESCMdPsy2_0(.din(n25434), .dout(n25437));
    jdff dff_A_f70mi43T6_0(.din(n25431), .dout(n25434));
    jdff dff_A_S3U6ijvB5_0(.din(n25428), .dout(n25431));
    jdff dff_A_9695fvsc5_0(.din(n25425), .dout(n25428));
    jdff dff_A_lW3A9Ekv9_0(.din(n25422), .dout(n25425));
    jdff dff_A_aFRatdU13_0(.din(n25419), .dout(n25422));
    jdff dff_A_nD75eIp11_0(.din(n25416), .dout(n25419));
    jdff dff_A_OoJRoECC9_0(.din(n25413), .dout(n25416));
    jdff dff_A_XddnKyiD5_0(.din(n25410), .dout(n25413));
    jdff dff_A_32pOtW9D1_1(.din(n2653), .dout(n25410));
    jdff dff_A_dCiS2op41_0(.din(n25404), .dout(G877));
    jdff dff_A_mR46Ugkq4_0(.din(n25401), .dout(n25404));
    jdff dff_A_eEBuOLFI7_0(.din(n25398), .dout(n25401));
    jdff dff_A_pqSbxMkD1_0(.din(n25395), .dout(n25398));
    jdff dff_A_5KMMxAwb2_0(.din(n25392), .dout(n25395));
    jdff dff_A_o2a6b3xQ4_0(.din(n25389), .dout(n25392));
    jdff dff_A_7hpTfjw56_0(.din(n25386), .dout(n25389));
    jdff dff_A_Nhj46LBa6_0(.din(n25383), .dout(n25386));
    jdff dff_A_SWEKU9a34_0(.din(n25380), .dout(n25383));
    jdff dff_A_4EIEZhWY3_0(.din(n25377), .dout(n25380));
    jdff dff_A_CFAsKBJq7_0(.din(n25374), .dout(n25377));
    jdff dff_A_kvuU1oFX2_0(.din(n25371), .dout(n25374));
    jdff dff_A_moeM5zwB5_0(.din(n25368), .dout(n25371));
    jdff dff_A_eSKIkpYy0_0(.din(n25365), .dout(n25368));
    jdff dff_A_T9WIBBTr5_0(.din(n25362), .dout(n25365));
    jdff dff_A_g1MK8hkL5_0(.din(n25359), .dout(n25362));
    jdff dff_A_y5o85UER5_1(.din(n2595), .dout(n25359));
    jdff dff_A_LYLIQECz2_0(.din(n25353), .dout(G875));
    jdff dff_A_83uEDLpM4_0(.din(n25350), .dout(n25353));
    jdff dff_A_WVPwuZV38_0(.din(n25347), .dout(n25350));
    jdff dff_A_A9GE2VRZ3_0(.din(n25344), .dout(n25347));
    jdff dff_A_iAyjbgUq2_0(.din(n25341), .dout(n25344));
    jdff dff_A_fio9PFVt0_0(.din(n25338), .dout(n25341));
    jdff dff_A_MkKoFrcX8_0(.din(n25335), .dout(n25338));
    jdff dff_A_deqvx5Zb0_0(.din(n25332), .dout(n25335));
    jdff dff_A_qlFVpBF09_0(.din(n25329), .dout(n25332));
    jdff dff_A_eIEMQ4sF1_0(.din(n25326), .dout(n25329));
    jdff dff_A_3AnIbj842_0(.din(n25323), .dout(n25326));
    jdff dff_A_dBjPSm9l5_0(.din(n25320), .dout(n25323));
    jdff dff_A_nX7Q4mEr4_0(.din(n25317), .dout(n25320));
    jdff dff_A_iBqs50su2_0(.din(n25314), .dout(n25317));
    jdff dff_A_hI1Tcukw9_0(.din(n25311), .dout(n25314));
    jdff dff_A_lkGGGKZR7_1(.din(n2553), .dout(n25311));
    jdff dff_A_4MmVsxrl7_0(.din(n25305), .dout(G873));
    jdff dff_A_jYA1aPvp5_0(.din(n25302), .dout(n25305));
    jdff dff_A_EPsyu48S8_0(.din(n25299), .dout(n25302));
    jdff dff_A_tPCvkRa59_0(.din(n25296), .dout(n25299));
    jdff dff_A_O6Qpz3XO9_0(.din(n25293), .dout(n25296));
    jdff dff_A_Q1CVm3Fv4_0(.din(n25290), .dout(n25293));
    jdff dff_A_52Dt3Y2q1_0(.din(n25287), .dout(n25290));
    jdff dff_A_VjyYokhV5_0(.din(n25284), .dout(n25287));
    jdff dff_A_Qo4FkX5p5_0(.din(n25281), .dout(n25284));
    jdff dff_A_RcngK7Hr4_0(.din(n25278), .dout(n25281));
    jdff dff_A_2tKugoVb1_0(.din(n25275), .dout(n25278));
    jdff dff_A_bMXasXir8_0(.din(n25272), .dout(n25275));
    jdff dff_A_OyKzx4fv1_0(.din(n25269), .dout(n25272));
    jdff dff_A_NTttsbUL7_0(.din(n25266), .dout(n25269));
    jdff dff_A_ORWvyfmF9_1(.din(n2514), .dout(n25266));
    jdff dff_A_xk218FQj0_0(.din(n25260), .dout(G871));
    jdff dff_A_OidMD6HS4_0(.din(n25257), .dout(n25260));
    jdff dff_A_rZhRhsc42_0(.din(n25254), .dout(n25257));
    jdff dff_A_N75vCvc63_0(.din(n25251), .dout(n25254));
    jdff dff_A_h8qWiK589_0(.din(n25248), .dout(n25251));
    jdff dff_A_GQn8F1U73_0(.din(n25245), .dout(n25248));
    jdff dff_A_7o2950PG1_0(.din(n25242), .dout(n25245));
    jdff dff_A_xgoXUh0e2_0(.din(n25239), .dout(n25242));
    jdff dff_A_3rMJ9UZe3_0(.din(n25236), .dout(n25239));
    jdff dff_A_l8GjwcZV4_0(.din(n25233), .dout(n25236));
    jdff dff_A_D7X7ut397_0(.din(n25230), .dout(n25233));
    jdff dff_A_vvDe9zXd5_0(.din(n25227), .dout(n25230));
    jdff dff_A_PwVeE3Jp6_1(.din(n2479), .dout(n25227));
    jdff dff_A_SkCjaWIe4_0(.din(n25221), .dout(G859));
    jdff dff_A_xMM7kB9L9_0(.din(n25218), .dout(n25221));
    jdff dff_A_8HJp41DM4_0(.din(n25215), .dout(n25218));
    jdff dff_A_hPvTzWf08_0(.din(n25212), .dout(n25215));
    jdff dff_A_1ewGm17r1_0(.din(n25209), .dout(n25212));
    jdff dff_A_W9HPife25_0(.din(n25206), .dout(n25209));
    jdff dff_A_wPEG65Sn7_0(.din(n25203), .dout(n25206));
    jdff dff_A_tloivukf8_0(.din(n25200), .dout(n25203));
    jdff dff_A_CwDC2akM7_0(.din(n25197), .dout(n25200));
    jdff dff_A_62uB0t0e8_0(.din(n25194), .dout(n25197));
    jdff dff_A_wlbXbTYG4_0(.din(n25191), .dout(n25194));
    jdff dff_A_XrzYRPur9_0(.din(n25188), .dout(n25191));
    jdff dff_A_v0jJKr6S3_0(.din(n25185), .dout(n25188));
    jdff dff_A_uCgvuOjA0_2(.din(n2426), .dout(n25185));
    jdff dff_A_XbWshpzL5_0(.din(n25179), .dout(G836));
    jdff dff_A_gfl235sD6_0(.din(n25176), .dout(n25179));
    jdff dff_A_7j605oDE4_0(.din(n25173), .dout(n25176));
    jdff dff_A_WbPvDGwR3_0(.din(n25170), .dout(n25173));
    jdff dff_A_z73FdqE16_0(.din(n25167), .dout(n25170));
    jdff dff_A_TVBGNKJm3_0(.din(n25164), .dout(n25167));
    jdff dff_A_GoJv94Cg9_0(.din(n25161), .dout(n25164));
    jdff dff_A_iIueJcY23_0(.din(n25158), .dout(n25161));
    jdff dff_A_uZTXq8lc1_0(.din(n25155), .dout(n25158));
    jdff dff_A_J0I4b43A6_0(.din(n25152), .dout(n25155));
    jdff dff_A_9Aen7PEI7_0(.din(n25149), .dout(n25152));
    jdff dff_A_anHhA3nr4_0(.din(n25146), .dout(n25149));
    jdff dff_A_HR1U3KUx8_0(.din(n25143), .dout(n25146));
    jdff dff_A_I4BcIiKF5_0(.din(n25140), .dout(n25143));
    jdff dff_A_Qv8LXOZe8_0(.din(n25137), .dout(n25140));
    jdff dff_A_4PavxOpF1_1(.din(n2384), .dout(n25137));
    jdff dff_A_DKQ6jBI75_0(.din(n25131), .dout(G834));
    jdff dff_A_NzvvGosU3_0(.din(n25128), .dout(n25131));
    jdff dff_A_zOelNpH78_0(.din(n25125), .dout(n25128));
    jdff dff_A_KTLNCtdL9_0(.din(n25122), .dout(n25125));
    jdff dff_A_p4evVdpo6_0(.din(n25119), .dout(n25122));
    jdff dff_A_3LcXvDW19_0(.din(n25116), .dout(n25119));
    jdff dff_A_SiWz9tmd0_0(.din(n25113), .dout(n25116));
    jdff dff_A_gTNtLMVa8_0(.din(n25110), .dout(n25113));
    jdff dff_A_0Lj3NiCX0_0(.din(n25107), .dout(n25110));
    jdff dff_A_C1xp1yR35_0(.din(n25104), .dout(n25107));
    jdff dff_A_quJ1lWA34_0(.din(n25101), .dout(n25104));
    jdff dff_A_eFblj2Xf9_0(.din(n25098), .dout(n25101));
    jdff dff_A_p0u4xb6B4_0(.din(n25095), .dout(n25098));
    jdff dff_A_D28W5EYA0_1(.din(n2345), .dout(n25095));
    jdff dff_A_3qqKZWbw7_0(.din(n25089), .dout(G832));
    jdff dff_A_UUzW6DcE1_0(.din(n25086), .dout(n25089));
    jdff dff_A_jI2swj6e0_0(.din(n25083), .dout(n25086));
    jdff dff_A_uChanSAJ6_0(.din(n25080), .dout(n25083));
    jdff dff_A_6i2p1qVP1_0(.din(n25077), .dout(n25080));
    jdff dff_A_v6oYvakf3_0(.din(n25074), .dout(n25077));
    jdff dff_A_brNZPAFR7_0(.din(n25071), .dout(n25074));
    jdff dff_A_gMPz0CsY7_0(.din(n25068), .dout(n25071));
    jdff dff_A_zMQESlBm2_0(.din(n25065), .dout(n25068));
    jdff dff_A_Hq1NbPsd3_0(.din(n25062), .dout(n25065));
    jdff dff_A_nmGTiiY77_0(.din(n25059), .dout(n25062));
    jdff dff_A_sCQVAFv34_0(.din(n25056), .dout(n25059));
    jdff dff_A_lbSS0iQn2_1(.din(n2310), .dout(n25056));
    jdff dff_A_9n7I7ANS1_0(.din(n25050), .dout(G722));
    jdff dff_A_HVknhIRf2_0(.din(n25047), .dout(n25050));
    jdff dff_A_IxD0SVC77_0(.din(n25044), .dout(n25047));
    jdff dff_A_nZEMvpum1_0(.din(n25041), .dout(n25044));
    jdff dff_A_iKvcm3a23_0(.din(n25038), .dout(n25041));
    jdff dff_A_oSiMinqj7_0(.din(n25035), .dout(n25038));
    jdff dff_A_RtUT9neU7_0(.din(n25032), .dout(n25035));
    jdff dff_A_eifgiYac8_0(.din(n25029), .dout(n25032));
    jdff dff_A_22YHxR059_0(.din(n25026), .dout(n25029));
    jdff dff_A_RGKrigig4_0(.din(n25023), .dout(n25026));
    jdff dff_A_GvaxARSZ6_0(.din(n25020), .dout(n25023));
    jdff dff_A_1LBFoYk27_0(.din(n25017), .dout(n25020));
    jdff dff_A_AZvzbllH8_0(.din(n25014), .dout(n25017));
    jdff dff_A_PsMfZTAJ4_2(.din(n2223), .dout(n25014));
    jdff dff_A_TatpMFv50_0(.din(n25008), .dout(G623));
    jdff dff_A_rNfutp1c7_0(.din(n25005), .dout(n25008));
    jdff dff_A_WhBfwYZv5_0(.din(n25002), .dout(n25005));
    jdff dff_A_oK2HLNsr3_0(.din(n24999), .dout(n25002));
    jdff dff_A_xxznfzh42_0(.din(n24996), .dout(n24999));
    jdff dff_A_Vbzm2oFo6_0(.din(n24993), .dout(n24996));
    jdff dff_A_GOSnef3m9_0(.din(n24990), .dout(n24993));
    jdff dff_A_ESVnY7PM7_0(.din(n24987), .dout(n24990));
    jdff dff_A_095S7ZBa5_0(.din(n24984), .dout(n24987));
    jdff dff_A_J3A90Aak2_1(.din(n2175), .dout(n24984));
    jdff dff_A_6hXiobxC6_0(.din(n24978), .dout(G861));
    jdff dff_A_rbsSBUxY7_0(.din(n24975), .dout(n24978));
    jdff dff_A_MVi9QUKQ4_0(.din(n24972), .dout(n24975));
    jdff dff_A_wSJYx65l6_0(.din(n24969), .dout(n24972));
    jdff dff_A_2XRKEYz92_0(.din(n24966), .dout(n24969));
    jdff dff_A_kfqdzEDL3_0(.din(n24963), .dout(n24966));
    jdff dff_A_QL9xJwti7_0(.din(n24960), .dout(n24963));
    jdff dff_A_0a0JOHZa0_0(.din(n24957), .dout(n24960));
    jdff dff_A_CX8VlSlG2_0(.din(n24954), .dout(n24957));
    jdff dff_A_TKvq1jPF5_0(.din(n24951), .dout(n24954));
    jdff dff_A_JzpEgPu87_0(.din(n24948), .dout(n24951));
    jdff dff_A_pAAohuZF1_0(.din(n24945), .dout(n24948));
    jdff dff_A_jufIAScu7_0(.din(n24942), .dout(n24945));
    jdff dff_A_7m5xpbTN7_0(.din(n24939), .dout(n24942));
    jdff dff_A_hqKisNM08_0(.din(n24936), .dout(n24939));
    jdff dff_A_EG4FM7dn2_0(.din(n24933), .dout(n24936));
    jdff dff_A_gUBJuViZ4_0(.din(n24930), .dout(n24933));
    jdff dff_A_an0UBJ8I1_1(.din(n2131), .dout(n24930));
    jdff dff_A_dv6LnonX7_0(.din(n24924), .dout(G838));
    jdff dff_A_KQ3X0ZOR6_0(.din(n24921), .dout(n24924));
    jdff dff_A_QEwFEsPo3_0(.din(n24918), .dout(n24921));
    jdff dff_A_CPYOVB9c5_0(.din(n24915), .dout(n24918));
    jdff dff_A_rwGFPfjV1_0(.din(n24912), .dout(n24915));
    jdff dff_A_tDp8novG2_0(.din(n24909), .dout(n24912));
    jdff dff_A_7CfHCbMw1_0(.din(n24906), .dout(n24909));
    jdff dff_A_KQP8SEZB1_0(.din(n24903), .dout(n24906));
    jdff dff_A_pdWw09zv8_0(.din(n24900), .dout(n24903));
    jdff dff_A_wxpy3BVI8_0(.din(n24897), .dout(n24900));
    jdff dff_A_AOIUlj3i0_0(.din(n24894), .dout(n24897));
    jdff dff_A_LOuHhHfj4_0(.din(n24891), .dout(n24894));
    jdff dff_A_5WNC0i9U5_0(.din(n24888), .dout(n24891));
    jdff dff_A_eULcMGbE2_0(.din(n24885), .dout(n24888));
    jdff dff_A_9ExCEcXI6_1(.din(n2097), .dout(n24885));
    jdff dff_A_kKS3FP4J0_0(.din(n24879), .dout(G822));
    jdff dff_A_FwMUFPoV6_0(.din(n24876), .dout(n24879));
    jdff dff_A_8TAhpgxJ2_0(.din(n24873), .dout(n24876));
    jdff dff_A_0H6mhUGq6_0(.din(n24870), .dout(n24873));
    jdff dff_A_Wd7ai7VE9_0(.din(n24867), .dout(n24870));
    jdff dff_A_rGc7iKsR2_0(.din(n24864), .dout(n24867));
    jdff dff_A_XjWylWI51_0(.din(n24861), .dout(n24864));
    jdff dff_A_J3fltsUP7_0(.din(n24858), .dout(n24861));
    jdff dff_A_o7Y8otNz4_0(.din(n24855), .dout(n24858));
    jdff dff_A_YX4Gu2rD1_0(.din(n24852), .dout(n24855));
    jdff dff_A_Q196gJ983_0(.din(n24849), .dout(n24852));
    jdff dff_A_6TMyAyPJ9_0(.din(n24846), .dout(n24849));
    jdff dff_A_5o9JObNK3_0(.din(n24843), .dout(n24846));
    jdff dff_A_3KS7syv66_0(.din(n24840), .dout(n24843));
    jdff dff_A_njN7BIqv7_0(.din(n24837), .dout(n24840));
    jdff dff_A_UWlpq2183_0(.din(n24834), .dout(n24837));
    jdff dff_A_6HeZkhuj6_0(.din(n24831), .dout(n24834));
    jdff dff_A_8EZQGkaj3_0(.din(n24828), .dout(n24831));
    jdff dff_A_wAgdn2DK8_0(.din(n24825), .dout(n24828));
    jdff dff_A_hgFfuhYA3_1(.din(n2040), .dout(n24825));
    jdff dff_A_QHnbNUT07_0(.din(n24819), .dout(G629));
    jdff dff_A_JDnLuERo5_0(.din(n24816), .dout(n24819));
    jdff dff_A_hxVwygIH9_0(.din(n24813), .dout(n24816));
    jdff dff_A_sqN5JeLQ7_0(.din(n24810), .dout(n24813));
    jdff dff_A_Gf2jRHr16_0(.din(n24807), .dout(n24810));
    jdff dff_A_wHMlGAhe1_0(.din(n24804), .dout(n24807));
    jdff dff_A_TfHZUdBq6_0(.din(n24801), .dout(n24804));
    jdff dff_A_hBPpjwvc4_0(.din(n24798), .dout(n24801));
    jdff dff_A_1XTfuPD71_0(.din(n24795), .dout(n24798));
    jdff dff_A_sh5jV3hW6_0(.din(n24792), .dout(n24795));
    jdff dff_A_hz8SHt0D4_0(.din(n24789), .dout(n24792));
    jdff dff_A_c3eQQTJu4_0(.din(n24786), .dout(n24789));
    jdff dff_A_QhGHobqZ0_0(.din(n24783), .dout(n24786));
    jdff dff_A_HUDI3Dhr7_0(.din(n24780), .dout(n24783));
    jdff dff_A_Znsu090U2_2(.din(n5821), .dout(n24780));
    jdff dff_A_PCsd5L9P9_0(.din(n24774), .dout(G621));
    jdff dff_A_tjDiisG77_0(.din(n24771), .dout(n24774));
    jdff dff_A_UZitD0P75_0(.din(n24768), .dout(n24771));
    jdff dff_A_iksfG1dY1_0(.din(n24765), .dout(n24768));
    jdff dff_A_TAC9M9JF0_0(.din(n24762), .dout(n24765));
    jdff dff_A_thk2pDGw4_0(.din(n24759), .dout(n24762));
    jdff dff_A_VMqkaL9U6_0(.din(n24756), .dout(n24759));
    jdff dff_A_NrzH5RsR3_0(.din(n24753), .dout(n24756));
    jdff dff_A_Tqmo8nN45_0(.din(n24750), .dout(n24753));
    jdff dff_A_BB1WxiYa9_0(.din(n24747), .dout(n24750));
    jdff dff_A_U7OSUIat9_0(.din(n24744), .dout(n24747));
    jdff dff_A_Rt79gU1P5_0(.din(n24741), .dout(n24744));
    jdff dff_A_qvv5I8vh5_0(.din(n24738), .dout(n24741));
    jdff dff_A_B0akqYdF7_2(.din(n5817), .dout(n24738));
    jdff dff_A_BxyG4Isx5_0(.din(n24732), .dout(G618));
    jdff dff_A_GqrtkXJw6_0(.din(n24729), .dout(n24732));
    jdff dff_A_SgNjeYdC0_0(.din(n24726), .dout(n24729));
    jdff dff_A_3Svn1WWl9_0(.din(n24723), .dout(n24726));
    jdff dff_A_2tJdZ4Iw1_0(.din(n24720), .dout(n24723));
    jdff dff_A_2S9IQ4Vn5_0(.din(n24717), .dout(n24720));
    jdff dff_A_ZTqyAL0G6_0(.din(n24714), .dout(n24717));
    jdff dff_A_lo68ThQf3_0(.din(n24711), .dout(n24714));
    jdff dff_A_wHyvzA8D8_0(.din(n24708), .dout(n24711));
    jdff dff_A_f1PNTAgp5_0(.din(n24705), .dout(n24708));
    jdff dff_A_PV3IfrPl2_0(.din(n24702), .dout(n24705));
    jdff dff_A_lA1EDnP07_0(.din(n24699), .dout(n24702));
    jdff dff_A_5Ce3RTXV1_0(.din(n24696), .dout(n24699));
    jdff dff_A_oGdPn1nK8_0(.din(n24693), .dout(n24696));
    jdff dff_A_XZnSM4Bv2_2(.din(n1996), .dout(n24693));
    jdff dff_A_vaK6s1wt0_0(.din(n24687), .dout(G591));
    jdff dff_A_MFYl9Z271_0(.din(n24684), .dout(n24687));
    jdff dff_A_T0qagvLT7_0(.din(n24681), .dout(n24684));
    jdff dff_A_ylvXNnnE9_0(.din(n24678), .dout(n24681));
    jdff dff_A_imkArTzf6_0(.din(n24675), .dout(n24678));
    jdff dff_A_KQ0wm0q25_0(.din(n24672), .dout(n24675));
    jdff dff_A_74FdOBZp5_0(.din(n24669), .dout(n24672));
    jdff dff_A_GTUDroBe6_0(.din(n24666), .dout(n24669));
    jdff dff_A_agM5eRlM2_0(.din(n24663), .dout(n24666));
    jdff dff_A_KZ6E29cY1_0(.din(n24660), .dout(n24663));
    jdff dff_A_q48AADeD4_0(.din(n24657), .dout(n24660));
    jdff dff_A_hZpNyaxf5_0(.din(n24654), .dout(n24657));
    jdff dff_A_l2Yh8SJN9_0(.din(n24651), .dout(n24654));
    jdff dff_A_vKR5DkTS6_2(.din(n1882), .dout(n24651));
    jdff dff_A_DAIpVBCT2_0(.din(n24645), .dout(G1004));
    jdff dff_A_x4WjN8389_0(.din(n24642), .dout(n24645));
    jdff dff_A_3eEVLCv52_0(.din(n24639), .dout(n24642));
    jdff dff_A_vnD58Lnw5_0(.din(n24636), .dout(n24639));
    jdff dff_A_Oo3iQI7s2_0(.din(n24633), .dout(n24636));
    jdff dff_A_A3B0aA2U6_0(.din(n24630), .dout(n24633));
    jdff dff_A_ZOroC7IB1_0(.din(n24627), .dout(n24630));
    jdff dff_A_rASdqLYY9_0(.din(n24624), .dout(n24627));
    jdff dff_A_fvr5Y7cP2_0(.din(n24621), .dout(n24624));
    jdff dff_A_GQzo0G338_0(.din(n24618), .dout(n24621));
    jdff dff_A_NVQh7i3k5_0(.din(n24615), .dout(n24618));
    jdff dff_A_FTsbSBtP3_0(.din(n24612), .dout(n24615));
    jdff dff_A_rQy1K00S9_0(.din(n24609), .dout(n24612));
    jdff dff_A_w04x8hvn5_0(.din(n24606), .dout(n24609));
    jdff dff_A_3SyNmhWU4_0(.din(n24603), .dout(n24606));
    jdff dff_A_jHLZZbYD8_0(.din(n24600), .dout(n24603));
    jdff dff_A_6PKRrom93_0(.din(n24597), .dout(n24600));
    jdff dff_A_XBD0ESze7_0(.din(n24594), .dout(n24597));
    jdff dff_A_u35H4Nyf2_0(.din(n24591), .dout(n24594));
    jdff dff_A_moFeEk9L8_0(.din(n24588), .dout(n24591));
    jdff dff_A_NBBiu6xp2_0(.din(n24585), .dout(n24588));
    jdff dff_A_7s0FSjaT0_0(.din(n24582), .dout(n24585));
    jdff dff_A_tW43U9KN1_1(.din(n1738), .dout(n24582));
    jdff dff_A_GVvo75fl8_0(.din(n24576), .dout(G1002));
    jdff dff_A_DGGQpU6e9_0(.din(n24573), .dout(n24576));
    jdff dff_A_aHLi1u3A8_0(.din(n24570), .dout(n24573));
    jdff dff_A_hOU7wK100_0(.din(n24567), .dout(n24570));
    jdff dff_A_KcNSmz6o9_0(.din(n24564), .dout(n24567));
    jdff dff_A_mQ3bit1g5_0(.din(n24561), .dout(n24564));
    jdff dff_A_sV3M7dZY7_0(.din(n24558), .dout(n24561));
    jdff dff_A_rAk1AOeY4_0(.din(n24555), .dout(n24558));
    jdff dff_A_wjOrQWWf2_0(.din(n24552), .dout(n24555));
    jdff dff_A_AZEwqLtC2_0(.din(n24549), .dout(n24552));
    jdff dff_A_UYjP4O1j9_0(.din(n24546), .dout(n24549));
    jdff dff_A_TBPKl1lf1_0(.din(n24543), .dout(n24546));
    jdff dff_A_FUU9QeKu5_0(.din(n24540), .dout(n24543));
    jdff dff_A_QRrpYB9c1_0(.din(n24537), .dout(n24540));
    jdff dff_A_w6kU9sVE5_0(.din(n24534), .dout(n24537));
    jdff dff_A_jz0cGITH3_0(.din(n24531), .dout(n24534));
    jdff dff_A_Too8TLhh7_0(.din(n24528), .dout(n24531));
    jdff dff_A_BxAN3miV1_0(.din(n24525), .dout(n24528));
    jdff dff_A_QyN45Ac36_0(.din(n24522), .dout(n24525));
    jdff dff_A_BvnYNZOB3_0(.din(n24519), .dout(n24522));
    jdff dff_A_8gTHU8iS2_0(.din(n24516), .dout(n24519));
    jdff dff_A_bwbB4dfk5_0(.din(n24513), .dout(n24516));
    jdff dff_A_lYUtd87F9_1(.din(n1699), .dout(n24513));
    jdff dff_A_BlRKl12i8_0(.din(n24507), .dout(G632));
    jdff dff_A_yoJGiT3X1_0(.din(n24504), .dout(n24507));
    jdff dff_A_K6d8Q3cU9_0(.din(n24501), .dout(n24504));
    jdff dff_A_JTr66KAw8_0(.din(n24498), .dout(n24501));
    jdff dff_A_kZduCUAf2_0(.din(n24495), .dout(n24498));
    jdff dff_A_y24CL9Za1_0(.din(n24492), .dout(n24495));
    jdff dff_A_iGAv61P90_0(.din(n24489), .dout(n24492));
    jdff dff_A_4IB0tKDg2_0(.din(n24486), .dout(n24489));
    jdff dff_A_O1jl03pm7_0(.din(n24483), .dout(n24486));
    jdff dff_A_BVDzHZaB2_0(.din(n24480), .dout(n24483));
    jdff dff_A_xgaQshQA7_0(.din(n24477), .dout(n24480));
    jdff dff_A_WSB7tngo1_0(.din(n24474), .dout(n24477));
    jdff dff_A_mWkPQRQa3_0(.din(n24471), .dout(n24474));
    jdff dff_A_iJ58sCCY4_0(.din(n24468), .dout(n24471));
    jdff dff_A_fn7ZApTB9_0(.din(n24465), .dout(n24468));
    jdff dff_A_txr7Wh484_0(.din(n24462), .dout(n24465));
    jdff dff_A_RZ4RQ0L23_2(.din(n5813), .dout(n24462));
    jdff dff_A_LwtLdMpv7_0(.din(n24456), .dout(G626));
    jdff dff_B_xJVd7vh19_1(.din(G136), .dout(n8401));
    jdff dff_B_NeekBaFp4_0(.din(G2824), .dout(n8404));
    jdff dff_B_H5ICgJDO2_1(.din(n366), .dout(n8407));
    jdff dff_B_T4h4UUWo7_1(.din(n390), .dout(n8410));
    jdff dff_B_m9fN94CJ9_2(.din(n412), .dout(n8413));
    jdff dff_B_FiSJvVee4_1(.din(n430), .dout(n8416));
    jdff dff_B_V1WkeonP1_1(.din(n438), .dout(n8419));
    jdff dff_B_dFPnBT7I9_0(.din(n442), .dout(n8422));
    jdff dff_B_AUPL4UiY9_1(.din(G24), .dout(n8425));
    jdff dff_B_ELkE3jRs4_1(.din(n458), .dout(n8428));
    jdff dff_B_PDYKQJxI2_0(.din(n462), .dout(n8431));
    jdff dff_B_u5UjHSah1_1(.din(G26), .dout(n8434));
    jdff dff_A_EyYMh1gb3_0(.din(n8439), .dout(n8436));
    jdff dff_A_hBgOeFl60_0(.din(n8442), .dout(n8439));
    jdff dff_A_naU6d0v53_0(.din(n8445), .dout(n8442));
    jdff dff_A_G139qUXC6_0(.din(G141), .dout(n8445));
    jdff dff_A_isseKvlO1_1(.din(n8451), .dout(n8448));
    jdff dff_A_V6aJmz8T1_1(.din(n8454), .dout(n8451));
    jdff dff_A_z4bRBYaS8_1(.din(n8457), .dout(n8454));
    jdff dff_A_9pMjfsWj9_1(.din(G141), .dout(n8457));
    jdff dff_B_7UYQIOoi0_1(.din(n478), .dout(n8461));
    jdff dff_B_Mo4niKpk5_0(.din(n482), .dout(n8464));
    jdff dff_B_9OtLNadY3_1(.din(G79), .dout(n8467));
    jdff dff_B_KSukqhV45_1(.din(n498), .dout(n8470));
    jdff dff_B_kBiuCscR6_1(.din(n8470), .dout(n8473));
    jdff dff_B_OnyUwNWl5_1(.din(G82), .dout(n8476));
    jdff dff_A_5H7xdybX2_0(.din(G2358), .dout(n8478));
    jdff dff_A_tmZmnfvl0_1(.din(G2358), .dout(n8481));
    jdff dff_A_2bn3N6YZ7_1(.din(n8487), .dout(n8484));
    jdff dff_A_3GYoWiuU0_1(.din(n8490), .dout(n8487));
    jdff dff_A_6YSjiHj03_1(.din(n8493), .dout(n8490));
    jdff dff_A_TU9gGnzH5_1(.din(G141), .dout(n8493));
    jdff dff_A_kMWxVDrh2_2(.din(n8499), .dout(n8496));
    jdff dff_A_jZ6qwYt01_2(.din(n8502), .dout(n8499));
    jdff dff_A_bRtp74It2_2(.din(n8505), .dout(n8502));
    jdff dff_A_edFeGmke8_2(.din(G141), .dout(n8505));
    jdff dff_B_ppgzI1QW4_1(.din(n563), .dout(n8509));
    jdff dff_B_WslEtSt70_2(.din(n1660), .dout(n8512));
    jdff dff_B_tLzJNkdT5_2(.din(n8512), .dout(n8515));
    jdff dff_B_Tm0nih7h7_2(.din(n1878), .dout(n8518));
    jdff dff_B_QAeNhS517_2(.din(n8518), .dout(n8521));
    jdff dff_B_HxvTgeKW1_1(.din(n1830), .dout(n8524));
    jdff dff_B_MCOzTeU11_1(.din(n8524), .dout(n8527));
    jdff dff_B_LM8uvOAs5_1(.din(n8527), .dout(n8530));
    jdff dff_B_Wl4ntgBJ8_1(.din(n8530), .dout(n8533));
    jdff dff_B_EUhZeJeu1_1(.din(n8533), .dout(n8536));
    jdff dff_B_QUdYuxkV7_1(.din(n8536), .dout(n8539));
    jdff dff_B_0mqaafZo4_1(.din(n1834), .dout(n8542));
    jdff dff_B_wDUsRAim3_1(.din(n8542), .dout(n8545));
    jdff dff_B_0oPw1zAC4_1(.din(n8545), .dout(n8548));
    jdff dff_B_SWBiYy6v8_1(.din(n8548), .dout(n8551));
    jdff dff_B_V8QbOeQJ2_1(.din(n8551), .dout(n8554));
    jdff dff_A_qgprgtJz4_1(.din(n8559), .dout(n8556));
    jdff dff_A_27kRFvmS5_1(.din(n8563), .dout(n8559));
    jdff dff_B_Gk7CQZEh4_3(.din(n1467), .dout(n8563));
    jdff dff_B_rVPAffzR7_2(.din(n1992), .dout(n8566));
    jdff dff_B_pKIMdEps8_2(.din(n8566), .dout(n8569));
    jdff dff_B_Ug8Ns8L68_1(.din(n1963), .dout(n8572));
    jdff dff_B_faKqSggN7_1(.din(n8572), .dout(n8575));
    jdff dff_A_TUQM28mg7_0(.din(n8580), .dout(n8577));
    jdff dff_A_LqDBCJup0_0(.din(n8583), .dout(n8580));
    jdff dff_A_hOsm0uFm5_0(.din(n8586), .dout(n8583));
    jdff dff_A_33gZIik94_0(.din(n8589), .dout(n8586));
    jdff dff_A_38Pjr5fa8_0(.din(n1656), .dout(n8589));
    jdff dff_B_8A802oyh5_0(.din(n2219), .dout(n8593));
    jdff dff_B_OPIUQjYO2_0(.din(n8593), .dout(n8596));
    jdff dff_B_VKWfFFBw6_0(.din(n8596), .dout(n8599));
    jdff dff_B_3alZRvZ45_0(.din(n8599), .dout(n8602));
    jdff dff_B_ZsBQnEA47_0(.din(n8602), .dout(n8605));
    jdff dff_B_NPYzj9ey3_0(.din(n8605), .dout(n8608));
    jdff dff_B_SESaneVA4_0(.din(n8608), .dout(n8611));
    jdff dff_B_GIU1vtYK0_0(.din(n8611), .dout(n8614));
    jdff dff_B_5IETn2KG4_0(.din(n8614), .dout(n8617));
    jdff dff_B_oplNXEDL6_0(.din(n8617), .dout(n8620));
    jdff dff_B_1PScmEgp4_0(.din(n2199), .dout(n8623));
    jdff dff_A_c8nKUhZi0_1(.din(n8628), .dout(n8625));
    jdff dff_A_seo738dG0_1(.din(n8631), .dout(n8628));
    jdff dff_A_HOayV5bp4_1(.din(n8634), .dout(n8631));
    jdff dff_A_AjbdDBgO6_1(.din(n8637), .dout(n8634));
    jdff dff_A_0T4J5fkg1_1(.din(n8640), .dout(n8637));
    jdff dff_A_dmjpzGTR8_1(.din(n8643), .dout(n8640));
    jdff dff_A_EKuwZTdH8_1(.din(n8646), .dout(n8643));
    jdff dff_A_iOrnd5Pj3_1(.din(n8649), .dout(n8646));
    jdff dff_A_zISZqvFC3_1(.din(n8652), .dout(n8649));
    jdff dff_A_losgSMuX1_1(.din(n2178), .dout(n8652));
    jdff dff_B_t0Lv9bLg5_0(.din(n2422), .dout(n8656));
    jdff dff_B_IY6zNTzk1_0(.din(n8656), .dout(n8659));
    jdff dff_B_Y1Crni0n0_0(.din(n8659), .dout(n8662));
    jdff dff_B_2lQCkvPH6_0(.din(n8662), .dout(n8665));
    jdff dff_B_DwmqAbxu1_0(.din(n8665), .dout(n8668));
    jdff dff_B_yO2Ld9hd1_0(.din(n8668), .dout(n8671));
    jdff dff_B_Wm19bM8k6_0(.din(n8671), .dout(n8674));
    jdff dff_B_CCcAZDDj1_0(.din(n8674), .dout(n8677));
    jdff dff_B_IdQgVWDq7_0(.din(n8677), .dout(n8680));
    jdff dff_B_ka2cL7cq3_0(.din(n8680), .dout(n8683));
    jdff dff_B_5Pi8sLZf6_2(.din(G61), .dout(n8686));
    jdff dff_B_Zj1aWoW30_0(.din(n2402), .dout(n8689));
    jdff dff_A_aRXDzq5t5_1(.din(n8694), .dout(n8691));
    jdff dff_A_54vCDj965_1(.din(n8697), .dout(n8694));
    jdff dff_A_Tjsbs8C07_1(.din(n8700), .dout(n8697));
    jdff dff_A_DjrPyRvT1_1(.din(n8703), .dout(n8700));
    jdff dff_A_RFF4a3Id4_1(.din(n8706), .dout(n8703));
    jdff dff_A_MGMIOyFU5_1(.din(n8709), .dout(n8706));
    jdff dff_A_SmllZ8dT6_1(.din(n8712), .dout(n8709));
    jdff dff_A_R7B2ihJO3_1(.din(n8715), .dout(n8712));
    jdff dff_A_Q5mkiUxB4_1(.din(n8718), .dout(n8715));
    jdff dff_A_GStFKiis3_1(.din(n2387), .dout(n8718));
    jdff dff_B_ifnOJc1U1_0(.din(n2824), .dout(n8722));
    jdff dff_B_ynuAR34F0_1(.din(n2802), .dout(n8725));
    jdff dff_B_bZ4GVU5u1_1(.din(n8725), .dout(n8728));
    jdff dff_B_nTaXBT9q0_1(.din(n8728), .dout(n8731));
    jdff dff_B_iqLddp8R8_0(.din(n2798), .dout(n8734));
    jdff dff_B_a6qgBGCl0_1(.din(n2855), .dout(n8737));
    jdff dff_B_cm89qgb02_1(.din(n8737), .dout(n8740));
    jdff dff_B_Y4rYfPA96_1(.din(n8740), .dout(n8743));
    jdff dff_B_qLpZPYUP7_1(.din(n8743), .dout(n8746));
    jdff dff_B_AxD9PwDr3_1(.din(n8746), .dout(n8749));
    jdff dff_B_0mYtizdg0_1(.din(n2839), .dout(n8752));
    jdff dff_B_CpVbdhlH2_1(.din(n8752), .dout(n8755));
    jdff dff_B_rpc69Qrr7_1(.din(n2929), .dout(n8758));
    jdff dff_B_jNILjL1c7_1(.din(n8758), .dout(n8761));
    jdff dff_B_M9tgOfoG7_1(.din(n8761), .dout(n8764));
    jdff dff_B_iFErXtgI2_1(.din(n8764), .dout(n8767));
    jdff dff_B_emGytDbn3_1(.din(n8767), .dout(n8770));
    jdff dff_B_2fWqJBgV3_1(.din(n8770), .dout(n8773));
    jdff dff_B_YPTvsFTT1_1(.din(n8773), .dout(n8776));
    jdff dff_B_xOad4M3p8_1(.din(n8776), .dout(n8779));
    jdff dff_B_fHaFuXNL2_1(.din(n8779), .dout(n8782));
    jdff dff_B_WddvAmdt9_1(.din(n8782), .dout(n8785));
    jdff dff_B_bIlR0n4s5_1(.din(n8785), .dout(n8788));
    jdff dff_B_bepvfav89_1(.din(n2937), .dout(n8791));
    jdff dff_B_PmBeLX548_1(.din(n8791), .dout(n8794));
    jdff dff_B_rzfiyyni7_1(.din(n8794), .dout(n8797));
    jdff dff_B_KQ2RIcrD9_1(.din(n8797), .dout(n8800));
    jdff dff_B_wEc3UVnu1_1(.din(n8800), .dout(n8803));
    jdff dff_B_oAnQ5GPc4_1(.din(n8803), .dout(n8806));
    jdff dff_B_3BuDIKdG0_1(.din(n8806), .dout(n8809));
    jdff dff_B_GQUnHn8g1_1(.din(n8809), .dout(n8812));
    jdff dff_B_eqL0ZiLh0_1(.din(n8812), .dout(n8815));
    jdff dff_B_pBC8bezt1_1(.din(n8815), .dout(n8818));
    jdff dff_B_zadYHcFr1_1(.din(n8818), .dout(n8821));
    jdff dff_B_gGhJvAVX2_0(.din(n2952), .dout(n8824));
    jdff dff_B_YFsucXNK3_0(.din(n3010), .dout(n8827));
    jdff dff_B_NX7qa5h72_0(.din(n8827), .dout(n8830));
    jdff dff_B_yX0JgzqU5_0(.din(n8830), .dout(n8833));
    jdff dff_B_P8VxAMFw6_0(.din(n8833), .dout(n8836));
    jdff dff_B_hu4syHSm8_0(.din(n8836), .dout(n8839));
    jdff dff_B_JB8MMbPs8_0(.din(n8839), .dout(n8842));
    jdff dff_B_LsuiAY8o2_0(.din(n8842), .dout(n8845));
    jdff dff_B_6zHzrdVX2_0(.din(n8845), .dout(n8848));
    jdff dff_B_V17nTjdJ3_0(.din(n8848), .dout(n8851));
    jdff dff_B_Ma1gKVog9_0(.din(n8851), .dout(n8854));
    jdff dff_B_s0XwuCNn0_1(.din(n2998), .dout(n8857));
    jdff dff_B_TEwl3wgg6_2(.din(G182), .dout(n8860));
    jdff dff_B_UXYvnfD98_2(.din(n8860), .dout(n8863));
    jdff dff_B_cX4vbk7M7_2(.din(G185), .dout(n8866));
    jdff dff_B_TH3AsybK0_1(.din(n2972), .dout(n8869));
    jdff dff_B_pJs3TDkA4_1(.din(n8869), .dout(n8872));
    jdff dff_B_PSJp4qRu8_1(.din(n8872), .dout(n8875));
    jdff dff_B_llc5HBxt6_1(.din(n2104), .dout(n8878));
    jdff dff_B_tPDLTsEY6_1(.din(n8878), .dout(n8881));
    jdff dff_B_X4NEc9x47_1(.din(n8881), .dout(n8884));
    jdff dff_B_7H31U1To0_1(.din(n8884), .dout(n8887));
    jdff dff_B_0fwNjf782_1(.din(n8887), .dout(n8890));
    jdff dff_B_kwHGDFZX7_0(.din(n2123), .dout(n8893));
    jdff dff_B_u9pdidx38_1(.din(n1182), .dout(n8896));
    jdff dff_B_3XLwB3kW2_1(.din(n1163), .dout(n8899));
    jdff dff_A_0kNBMird8_0(.din(n8904), .dout(n8901));
    jdff dff_A_qnGRR56D9_0(.din(n2111), .dout(n8904));
    jdff dff_B_llH03iJn7_1(.din(G117), .dout(n8908));
    jdff dff_B_uWQdhYHv7_1(.din(n8908), .dout(n8911));
    jdff dff_B_OT9KcLqn4_1(.din(n2010), .dout(n8914));
    jdff dff_B_GrmjhGxS4_1(.din(n8914), .dout(n8917));
    jdff dff_B_Wr6GDBT12_1(.din(n8917), .dout(n8920));
    jdff dff_A_3ZG8IpOA9_0(.din(n8925), .dout(n8922));
    jdff dff_A_68n6HSoo1_0(.din(n8928), .dout(n8925));
    jdff dff_A_ATfgVxmz3_0(.din(n8931), .dout(n8928));
    jdff dff_A_pJggtBVe3_0(.din(n8934), .dout(n8931));
    jdff dff_A_FkQn2sEm6_0(.din(n8937), .dout(n8934));
    jdff dff_A_MJ8r3R6z6_0(.din(n8940), .dout(n8937));
    jdff dff_A_DDxqCbB22_0(.din(n8943), .dout(n8940));
    jdff dff_A_9lKhqlHn3_0(.din(n8946), .dout(n8943));
    jdff dff_A_biLyGV7G6_0(.din(n8949), .dout(n8946));
    jdff dff_A_HR22AKG65_0(.din(n8952), .dout(n8949));
    jdff dff_A_AFcJoeIn8_0(.din(n2020), .dout(n8952));
    jdff dff_B_VjocPBUU2_1(.din(G131), .dout(n8956));
    jdff dff_B_5JNCKSIB9_1(.din(n8956), .dout(n8959));
    jdff dff_B_6C7xYPwX4_0(.din(n3056), .dout(n8962));
    jdff dff_B_6usAEpL71_0(.din(n8962), .dout(n8965));
    jdff dff_B_DPoBePda6_0(.din(n8965), .dout(n8968));
    jdff dff_B_p43uRxwh4_0(.din(n8968), .dout(n8971));
    jdff dff_B_PXHs6AVa0_0(.din(n8971), .dout(n8974));
    jdff dff_B_NCJWC3Zs6_0(.din(n8974), .dout(n8977));
    jdff dff_B_C9UyJnCz3_0(.din(n8977), .dout(n8980));
    jdff dff_B_nT9GyZhR6_0(.din(n8980), .dout(n8983));
    jdff dff_B_4kE6BgE56_0(.din(n8983), .dout(n8986));
    jdff dff_B_GmDFS35I0_0(.din(n8986), .dout(n8989));
    jdff dff_B_VSsnlerl0_0(.din(n8989), .dout(n8992));
    jdff dff_B_SCP58RGa4_0(.din(n8992), .dout(n8995));
    jdff dff_B_017KG9S71_0(.din(n8995), .dout(n8998));
    jdff dff_B_9ldMJKpa4_0(.din(n8998), .dout(n9001));
    jdff dff_B_qmgLwixf3_0(.din(n9001), .dout(n9004));
    jdff dff_B_UIq314s07_0(.din(n9004), .dout(n9007));
    jdff dff_B_IsG2THwt3_1(.din(n3025), .dout(n9010));
    jdff dff_A_TZScAyTj2_0(.din(n9015), .dout(n9012));
    jdff dff_A_QNrzqIJH1_0(.din(n9018), .dout(n9015));
    jdff dff_A_9hnClhKi8_0(.din(n9021), .dout(n9018));
    jdff dff_A_L0En3HXn6_0(.din(n9024), .dout(n9021));
    jdff dff_A_3K82hbXV2_0(.din(n9027), .dout(n9024));
    jdff dff_A_OpI0ot5M8_0(.din(n9030), .dout(n9027));
    jdff dff_A_zylMXVli7_0(.din(n15595), .dout(n9030));
    jdff dff_B_Po2ISzVd5_0(.din(n3098), .dout(n9034));
    jdff dff_B_ZRmtmCjC7_0(.din(n9034), .dout(n9037));
    jdff dff_B_hTIicSsr5_0(.din(n9037), .dout(n9040));
    jdff dff_B_mTUB5HaQ7_0(.din(n9040), .dout(n9043));
    jdff dff_B_7hy4n0E68_0(.din(n9043), .dout(n9046));
    jdff dff_B_otWUI5sG6_0(.din(n9046), .dout(n9049));
    jdff dff_B_XS6BAxRR8_0(.din(n9049), .dout(n9052));
    jdff dff_B_HaHF3kcj8_0(.din(n9052), .dout(n9055));
    jdff dff_B_ZyqN2vLL3_0(.din(n9055), .dout(n9058));
    jdff dff_B_qYCT38415_0(.din(n9058), .dout(n9061));
    jdff dff_B_p8auc4tf7_0(.din(n9061), .dout(n9064));
    jdff dff_B_fqGVN7Vg8_0(.din(n9064), .dout(n9067));
    jdff dff_B_DXGhJf8M6_0(.din(n9067), .dout(n9070));
    jdff dff_B_uKusfTFG7_0(.din(n9070), .dout(n9073));
    jdff dff_B_EmJXUkSS3_0(.din(n9073), .dout(n9076));
    jdff dff_B_QvF7cfS06_1(.din(n3067), .dout(n9079));
    jdff dff_B_JNeHI5JZ0_1(.din(n9079), .dout(n9082));
    jdff dff_A_MQEkn3ZQ3_0(.din(n9087), .dout(n9084));
    jdff dff_A_8JSkwwNG0_0(.din(n9090), .dout(n9087));
    jdff dff_A_SD5aRq3n2_0(.din(n9093), .dout(n9090));
    jdff dff_A_yHlDPozQ3_0(.din(n9096), .dout(n9093));
    jdff dff_A_KIAw0P6t3_0(.din(n9099), .dout(n9096));
    jdff dff_A_tJYE0Yn30_0(.din(n9102), .dout(n9099));
    jdff dff_A_6uxWNdtr7_0(.din(n9105), .dout(n9102));
    jdff dff_A_UZllMLiM0_0(.din(n9108), .dout(n9105));
    jdff dff_A_t1A3h8wG4_0(.din(n9111), .dout(n9108));
    jdff dff_A_Vrkc4mDz8_0(.din(n9114), .dout(n9111));
    jdff dff_A_pjGbuDnr6_0(.din(n9117), .dout(n9114));
    jdff dff_A_Cp83xP6V3_0(.din(n9120), .dout(n9117));
    jdff dff_A_Cqi6r2G91_0(.din(n9123), .dout(n9120));
    jdff dff_A_PyUVJ6Sk0_0(.din(n9126), .dout(n9123));
    jdff dff_A_p986CboN5_0(.din(G4088), .dout(n9126));
    jdff dff_A_6a5PsfXW0_2(.din(n9132), .dout(n9129));
    jdff dff_A_XA8MWyHc0_2(.din(n9135), .dout(n9132));
    jdff dff_A_8kFdNVLW4_2(.din(n9138), .dout(n9135));
    jdff dff_A_5wl5X6Qu4_2(.din(n9141), .dout(n9138));
    jdff dff_A_2uSKnKuM9_2(.din(n9144), .dout(n9141));
    jdff dff_A_OXGEE86E0_2(.din(n9147), .dout(n9144));
    jdff dff_A_KFXFmrLM3_2(.din(n9150), .dout(n9147));
    jdff dff_A_DkQQXndv4_2(.din(n9153), .dout(n9150));
    jdff dff_A_yxXdYlDR6_2(.din(n9156), .dout(n9153));
    jdff dff_A_iG2oJDo61_2(.din(n9159), .dout(n9156));
    jdff dff_A_uGZtE6xb4_2(.din(n9162), .dout(n9159));
    jdff dff_A_m8qufn2Y3_2(.din(n9165), .dout(n9162));
    jdff dff_A_3jfaWwH20_2(.din(n9168), .dout(n9165));
    jdff dff_A_W5PlwJbf8_2(.din(n9171), .dout(n9168));
    jdff dff_A_qaMVEAhk2_2(.din(n9174), .dout(n9171));
    jdff dff_A_FgbyN03F3_2(.din(G4088), .dout(n9174));
    jdff dff_A_VvG59TxG9_0(.din(n9180), .dout(n9177));
    jdff dff_A_rzUZXHyG7_0(.din(n9183), .dout(n9180));
    jdff dff_A_nuSZUysl8_0(.din(n9186), .dout(n9183));
    jdff dff_A_OadZqIXw7_0(.din(n9189), .dout(n9186));
    jdff dff_A_k39D8FCz7_0(.din(n9192), .dout(n9189));
    jdff dff_A_wQb28WFR7_0(.din(n9195), .dout(n9192));
    jdff dff_A_Kpw8bXjQ3_0(.din(n9198), .dout(n9195));
    jdff dff_A_21fj1h7t2_0(.din(n9201), .dout(n9198));
    jdff dff_A_OayhSrbs8_0(.din(n9204), .dout(n9201));
    jdff dff_A_Uj7yy23O6_0(.din(n9207), .dout(n9204));
    jdff dff_A_0VW1blZh0_0(.din(n9210), .dout(n9207));
    jdff dff_A_aBn7HYKn3_0(.din(n9213), .dout(n9210));
    jdff dff_A_RMKQ9xKZ3_0(.din(n2178), .dout(n9213));
    jdff dff_A_wMSaZ8gK4_2(.din(n9219), .dout(n9216));
    jdff dff_A_W6bTy4494_2(.din(n9222), .dout(n9219));
    jdff dff_A_lKCBf1TV2_2(.din(n9225), .dout(n9222));
    jdff dff_A_CIauddfq1_2(.din(n9228), .dout(n9225));
    jdff dff_A_6YOhI7Sq3_2(.din(n9231), .dout(n9228));
    jdff dff_A_IKtUNxUx4_2(.din(n9234), .dout(n9231));
    jdff dff_A_FrqyaWoV3_2(.din(n9237), .dout(n9234));
    jdff dff_A_8v3wnTHs3_2(.din(n9240), .dout(n9237));
    jdff dff_A_zbAwwr7D1_2(.din(n9243), .dout(n9240));
    jdff dff_A_3GY1SmH09_2(.din(n9246), .dout(n9243));
    jdff dff_A_WVYYgkO42_2(.din(n9249), .dout(n9246));
    jdff dff_A_h1z21ejw0_2(.din(n9252), .dout(n9249));
    jdff dff_A_oATnb0JV4_2(.din(n9255), .dout(n9252));
    jdff dff_A_yvKF8FNS8_2(.din(n9258), .dout(n9255));
    jdff dff_A_szCXB5hr2_2(.din(n2178), .dout(n9258));
    jdff dff_B_K0taASR83_0(.din(n3140), .dout(n9262));
    jdff dff_B_fgCIVJWI4_0(.din(n9262), .dout(n9265));
    jdff dff_B_Q390yZn54_0(.din(n9265), .dout(n9268));
    jdff dff_B_yjwzU9cr8_0(.din(n9268), .dout(n9271));
    jdff dff_B_t7VcwXUB3_0(.din(n9271), .dout(n9274));
    jdff dff_B_kDLvE5YN3_0(.din(n9274), .dout(n9277));
    jdff dff_B_WDpM9Pgp1_0(.din(n9277), .dout(n9280));
    jdff dff_B_XiOc0Asl2_0(.din(n9280), .dout(n9283));
    jdff dff_B_peDalsoS3_0(.din(n9283), .dout(n9286));
    jdff dff_B_50vjEcMR2_0(.din(n9286), .dout(n9289));
    jdff dff_B_E6G42R591_0(.din(n9289), .dout(n9292));
    jdff dff_B_7gGHSTfS2_0(.din(n9292), .dout(n9295));
    jdff dff_B_5cicOMT37_0(.din(n9295), .dout(n9298));
    jdff dff_B_wp0a28OD5_1(.din(n3109), .dout(n9301));
    jdff dff_A_Jo3bcgaK9_1(.din(n9306), .dout(n9303));
    jdff dff_A_CDwIySkN4_1(.din(n9309), .dout(n9306));
    jdff dff_A_OnXB51Bp8_1(.din(n9312), .dout(n9309));
    jdff dff_A_M7YEE43P3_1(.din(n9315), .dout(n9312));
    jdff dff_A_kg6GLHO41_1(.din(n9318), .dout(n9315));
    jdff dff_A_sddRlp4C4_1(.din(n9321), .dout(n9318));
    jdff dff_A_zz3pZw4u9_1(.din(n9324), .dout(n9321));
    jdff dff_A_4ZzXPOML7_1(.din(n9327), .dout(n9324));
    jdff dff_A_b2kEv4le4_1(.din(n9330), .dout(n9327));
    jdff dff_A_PV1fhr5j4_1(.din(n9333), .dout(n9330));
    jdff dff_A_ReqLpIV65_1(.din(n9336), .dout(n9333));
    jdff dff_A_OTCTdaMt9_1(.din(n2178), .dout(n9336));
    jdff dff_A_0ZF2PpQz8_1(.din(n9342), .dout(n9339));
    jdff dff_A_dfc0ZRY10_1(.din(n9345), .dout(n9342));
    jdff dff_A_wZfI1sYx5_1(.din(n9348), .dout(n9345));
    jdff dff_A_L00xSYiA9_1(.din(n9351), .dout(n9348));
    jdff dff_A_9hH4qnTQ4_1(.din(n9354), .dout(n9351));
    jdff dff_A_lfyjIjk33_1(.din(n9357), .dout(n9354));
    jdff dff_A_KwGtuKwl6_1(.din(n9360), .dout(n9357));
    jdff dff_A_rDygWqJN8_1(.din(n9363), .dout(n9360));
    jdff dff_A_S0JEouFS1_1(.din(n9366), .dout(n9363));
    jdff dff_A_kWWrLE427_1(.din(n9369), .dout(n9366));
    jdff dff_A_mipak4EX4_1(.din(n9372), .dout(n9369));
    jdff dff_A_z1tFrmCv4_1(.din(n9375), .dout(n9372));
    jdff dff_A_J40c4J9p9_1(.din(G4088), .dout(n9375));
    jdff dff_B_WvLGDAOl0_0(.din(n3182), .dout(n9379));
    jdff dff_B_OdkadJJI6_0(.din(n9379), .dout(n9382));
    jdff dff_B_CmNxNxjB0_0(.din(n9382), .dout(n9385));
    jdff dff_B_oBXown095_0(.din(n9385), .dout(n9388));
    jdff dff_B_cCeYb6eM9_0(.din(n9388), .dout(n9391));
    jdff dff_B_JQWwtTVl8_0(.din(n9391), .dout(n9394));
    jdff dff_B_nUqsHqs90_0(.din(n9394), .dout(n9397));
    jdff dff_B_ml71n9Iu4_0(.din(n9397), .dout(n9400));
    jdff dff_B_Y1IV97me7_0(.din(n9400), .dout(n9403));
    jdff dff_B_yL46Ax4v3_0(.din(n9403), .dout(n9406));
    jdff dff_B_fh5LHN6Z9_0(.din(n9406), .dout(n9409));
    jdff dff_B_yEGekuBd7_0(.din(n9409), .dout(n9412));
    jdff dff_B_WT21Q8Wg1_0(.din(n9412), .dout(n9415));
    jdff dff_B_PrVErDRB6_0(.din(n9415), .dout(n9418));
    jdff dff_B_pOXsZQ7t5_1(.din(n3151), .dout(n9421));
    jdff dff_B_TzjUy8CR7_1(.din(n9421), .dout(n9424));
    jdff dff_B_BkBJegN79_1(.din(n9424), .dout(n9427));
    jdff dff_A_foNLMS0P2_0(.din(n15558), .dout(n9429));
    jdff dff_A_Hu32o2cR8_2(.din(n9435), .dout(n9432));
    jdff dff_A_ptkvh7EA1_2(.din(n15558), .dout(n9435));
    jdff dff_B_3CTSQPKb8_1(.din(n3202), .dout(n9439));
    jdff dff_B_fijrpWob9_1(.din(n9439), .dout(n9442));
    jdff dff_B_cH8S5oks3_1(.din(n9442), .dout(n9445));
    jdff dff_B_E5l4s9jY8_1(.din(n9445), .dout(n9448));
    jdff dff_B_zycsE9ZW7_1(.din(n9448), .dout(n9451));
    jdff dff_B_7ZP9AhMz0_1(.din(n9451), .dout(n9454));
    jdff dff_B_a5S6kHUC3_1(.din(n9454), .dout(n9457));
    jdff dff_B_0YZn9x8B0_1(.din(n9457), .dout(n9460));
    jdff dff_B_SbA090H36_1(.din(n9460), .dout(n9463));
    jdff dff_B_DRl243DJ4_1(.din(n9463), .dout(n9466));
    jdff dff_B_SsELJ9Fa7_1(.din(n9466), .dout(n9469));
    jdff dff_B_JRRzcMFs5_1(.din(n9469), .dout(n9472));
    jdff dff_B_2xTmNc0b9_1(.din(n9472), .dout(n9475));
    jdff dff_B_EitWhjPr9_1(.din(n9475), .dout(n9478));
    jdff dff_B_sw0kQIIT5_1(.din(n9478), .dout(n9481));
    jdff dff_A_ebht2U5w7_0(.din(n9486), .dout(n9483));
    jdff dff_A_hV5J1of21_0(.din(n9489), .dout(n9486));
    jdff dff_A_sy4FFc0i5_0(.din(n9492), .dout(n9489));
    jdff dff_A_EB8dtqpN0_0(.din(n9495), .dout(n9492));
    jdff dff_A_4nLjo1g16_0(.din(n9498), .dout(n9495));
    jdff dff_A_p4UPIfMP6_0(.din(n9501), .dout(n9498));
    jdff dff_A_olaywdnc3_0(.din(n9504), .dout(n9501));
    jdff dff_A_p2PiHSc06_0(.din(n16000), .dout(n9504));
    jdff dff_B_KLHKgBge4_1(.din(n3190), .dout(n9508));
    jdff dff_B_fm2x8dKD1_1(.din(n9508), .dout(n9511));
    jdff dff_B_h9kxZlyU6_2(.din(G37), .dout(n9514));
    jdff dff_B_fKlRZZMc0_1(.din(n3238), .dout(n9517));
    jdff dff_B_8ooZeVHK3_1(.din(n9517), .dout(n9520));
    jdff dff_B_X8ZmFST18_1(.din(n9520), .dout(n9523));
    jdff dff_B_krsKa70A5_1(.din(n9523), .dout(n9526));
    jdff dff_B_67anivFM8_1(.din(n9526), .dout(n9529));
    jdff dff_B_pcoQU6oO2_1(.din(n9529), .dout(n9532));
    jdff dff_B_qlaTCUvJ4_1(.din(n9532), .dout(n9535));
    jdff dff_B_iAz9VOY70_1(.din(n9535), .dout(n9538));
    jdff dff_B_4QN1Pk018_1(.din(n9538), .dout(n9541));
    jdff dff_B_eZD9rZFq6_1(.din(n9541), .dout(n9544));
    jdff dff_B_WIKI6WIU3_1(.din(n9544), .dout(n9547));
    jdff dff_B_gSEg92IP8_1(.din(n9547), .dout(n9550));
    jdff dff_B_1Ho6YZSd5_1(.din(n9550), .dout(n9553));
    jdff dff_B_R3xuKQ1A8_1(.din(n9553), .dout(n9556));
    jdff dff_B_3RUDA86W1_0(.din(n3246), .dout(n9559));
    jdff dff_B_FiZVK3de1_1(.din(n3226), .dout(n9562));
    jdff dff_B_dSaYggRw8_1(.din(n9562), .dout(n9565));
    jdff dff_A_CABZ38Nm4_1(.din(n9570), .dout(n9567));
    jdff dff_A_Mhpg5Sw66_1(.din(n9573), .dout(n9570));
    jdff dff_A_2f3ygkh53_1(.din(n9576), .dout(n9573));
    jdff dff_A_1pNpKMnn3_1(.din(n9579), .dout(n9576));
    jdff dff_A_UFtGMjOv9_1(.din(n9582), .dout(n9579));
    jdff dff_A_G7Upt35M5_1(.din(n9585), .dout(n9582));
    jdff dff_A_wHomhmqu2_1(.din(n9588), .dout(n9585));
    jdff dff_A_2evvlSFa6_1(.din(n9591), .dout(n9588));
    jdff dff_A_THPnx7fu3_1(.din(n9594), .dout(n9591));
    jdff dff_A_XpyDvBDb2_1(.din(n9597), .dout(n9594));
    jdff dff_A_svcPAzKj3_1(.din(n9600), .dout(n9597));
    jdff dff_A_otY84Bj83_1(.din(n9603), .dout(n9600));
    jdff dff_A_1xzMNccD6_1(.din(n9606), .dout(n9603));
    jdff dff_A_MIEN68w72_1(.din(n9609), .dout(n9606));
    jdff dff_A_p2KaDZoD7_1(.din(n2387), .dout(n9609));
    jdff dff_B_MZAmZeka7_2(.din(G20), .dout(n9613));
    jdff dff_A_4gwFou728_1(.din(n9618), .dout(n9615));
    jdff dff_A_nDKLfZ6A8_1(.din(n9621), .dout(n9618));
    jdff dff_A_LVXdMjz14_1(.din(n9624), .dout(n9621));
    jdff dff_A_UMAllwSa6_1(.din(n9627), .dout(n9624));
    jdff dff_A_ZbHJusbg5_1(.din(n9630), .dout(n9627));
    jdff dff_A_eeUq2Ocq7_1(.din(n9633), .dout(n9630));
    jdff dff_A_2cVaDhVt5_1(.din(n9636), .dout(n9633));
    jdff dff_A_n6PN850D5_1(.din(n9639), .dout(n9636));
    jdff dff_A_OSHVIPAF3_1(.din(n9642), .dout(n9639));
    jdff dff_A_MCF6eygg6_1(.din(n9645), .dout(n9642));
    jdff dff_A_ATIub3M57_1(.din(n9648), .dout(n9645));
    jdff dff_A_cZyCyK2P3_1(.din(n9651), .dout(n9648));
    jdff dff_A_8MendlBx5_1(.din(n9654), .dout(n9651));
    jdff dff_A_4GTmbS0q8_1(.din(n9657), .dout(n9654));
    jdff dff_A_R5t2f0y17_1(.din(n9660), .dout(n9657));
    jdff dff_A_DGMxBQG38_1(.din(G4089), .dout(n9660));
    jdff dff_B_U62sgSUC8_1(.din(n3274), .dout(n9664));
    jdff dff_B_xB9NwQL76_1(.din(n9664), .dout(n9667));
    jdff dff_B_y19k6eIt3_1(.din(n9667), .dout(n9670));
    jdff dff_B_s05LFa7k9_1(.din(n9670), .dout(n9673));
    jdff dff_B_i3CRBM249_1(.din(n9673), .dout(n9676));
    jdff dff_B_S6GmqtZn9_1(.din(n9676), .dout(n9679));
    jdff dff_B_ul5oidY57_1(.din(n9679), .dout(n9682));
    jdff dff_B_fdimDfiK2_1(.din(n9682), .dout(n9685));
    jdff dff_B_3GWiesPE3_1(.din(n9685), .dout(n9688));
    jdff dff_B_AUFu4Drc0_1(.din(n9688), .dout(n9691));
    jdff dff_B_KDCB6Twn2_1(.din(n9691), .dout(n9694));
    jdff dff_B_QtbKjWVe1_1(.din(n9694), .dout(n9697));
    jdff dff_B_2Krg9KE16_1(.din(n3262), .dout(n9700));
    jdff dff_B_wsR42LE81_1(.din(n9700), .dout(n9703));
    jdff dff_A_AdgkasZo8_0(.din(n9708), .dout(n9705));
    jdff dff_A_3wMHiP440_0(.din(n9711), .dout(n9708));
    jdff dff_A_2CVtRpox0_0(.din(n9714), .dout(n9711));
    jdff dff_A_JpFHzrtN9_0(.din(n9717), .dout(n9714));
    jdff dff_A_4lukrovC8_0(.din(n9720), .dout(n9717));
    jdff dff_A_7HUDM1Yw4_0(.din(n9723), .dout(n9720));
    jdff dff_A_Azb8ug1R9_0(.din(n9726), .dout(n9723));
    jdff dff_A_Bb8YF7Ma6_0(.din(n9729), .dout(n9726));
    jdff dff_A_cQkQ1UbB1_0(.din(n9732), .dout(n9729));
    jdff dff_A_pcWhhPNn3_0(.din(n9735), .dout(n9732));
    jdff dff_A_fVceHLmP6_0(.din(n9738), .dout(n9735));
    jdff dff_A_z4pdcwoX3_0(.din(n2387), .dout(n9738));
    jdff dff_A_33GAKJi55_2(.din(n9744), .dout(n9741));
    jdff dff_A_EgB1K0cH3_2(.din(n9747), .dout(n9744));
    jdff dff_A_RUC4aArw9_2(.din(n9750), .dout(n9747));
    jdff dff_A_DunTaVRw4_2(.din(n9753), .dout(n9750));
    jdff dff_A_2ZDS1ZtK8_2(.din(n9756), .dout(n9753));
    jdff dff_A_o4Hb3cco8_2(.din(n9759), .dout(n9756));
    jdff dff_A_7SqNkHp28_2(.din(n9762), .dout(n9759));
    jdff dff_A_B21LMjTn3_2(.din(n9765), .dout(n9762));
    jdff dff_A_nB8D89q28_2(.din(n9768), .dout(n9765));
    jdff dff_A_HIX9uVYh9_2(.din(n9771), .dout(n9768));
    jdff dff_A_RyWzwAUx5_2(.din(n9774), .dout(n9771));
    jdff dff_A_98xNmKra5_2(.din(n9777), .dout(n9774));
    jdff dff_A_js8pimOP0_2(.din(n2387), .dout(n9777));
    jdff dff_B_RPIWd08X5_2(.din(G17), .dout(n9781));
    jdff dff_A_H2jeIYjO1_0(.din(n9786), .dout(n9783));
    jdff dff_A_nrzLWmSR1_0(.din(n9789), .dout(n9786));
    jdff dff_A_44DkNbkz7_0(.din(n9792), .dout(n9789));
    jdff dff_A_m6WbrJ8L0_0(.din(n9795), .dout(n9792));
    jdff dff_A_lapcYyYX9_0(.din(n9798), .dout(n9795));
    jdff dff_A_O62LtL2A0_0(.din(n9801), .dout(n9798));
    jdff dff_A_5Gdr1D451_0(.din(n9804), .dout(n9801));
    jdff dff_A_XuHovybZ8_0(.din(n9807), .dout(n9804));
    jdff dff_A_Wc0Fc5UN9_0(.din(n9810), .dout(n9807));
    jdff dff_A_27Pe6pAY1_0(.din(n9813), .dout(n9810));
    jdff dff_A_pVhTbSdy7_0(.din(n9816), .dout(n9813));
    jdff dff_A_BUisNmyH8_0(.din(n9819), .dout(n9816));
    jdff dff_A_EGw3OCqi1_0(.din(G4089), .dout(n9819));
    jdff dff_A_oK2ZZWd80_2(.din(n9825), .dout(n9822));
    jdff dff_A_cbpnOs2t2_2(.din(n9828), .dout(n9825));
    jdff dff_A_1dQ0nBsJ4_2(.din(n9831), .dout(n9828));
    jdff dff_A_wnUlBMJS2_2(.din(n9834), .dout(n9831));
    jdff dff_A_tAIIr8Mb2_2(.din(n9837), .dout(n9834));
    jdff dff_A_U4VeFLT89_2(.din(n9840), .dout(n9837));
    jdff dff_A_0YTHVqHw1_2(.din(n9843), .dout(n9840));
    jdff dff_A_Uv1ru2fl1_2(.din(n9846), .dout(n9843));
    jdff dff_A_UYzecIFh4_2(.din(n9849), .dout(n9846));
    jdff dff_A_QgoiUmMT1_2(.din(n9852), .dout(n9849));
    jdff dff_A_TntnKZWC6_2(.din(n9855), .dout(n9852));
    jdff dff_A_P7p4HuS22_2(.din(n9858), .dout(n9855));
    jdff dff_A_6eMntC6i9_2(.din(n9861), .dout(n9858));
    jdff dff_A_i9DnFPfo7_2(.din(n9864), .dout(n9861));
    jdff dff_A_d2WmELSA3_2(.din(G4089), .dout(n9864));
    jdff dff_B_dwgKOCQT5_0(.din(n3326), .dout(n9868));
    jdff dff_B_MJXpMlSz8_0(.din(n9868), .dout(n9871));
    jdff dff_B_lVtnwA7P9_0(.din(n9871), .dout(n9874));
    jdff dff_B_q54FTbbG2_0(.din(n9874), .dout(n9877));
    jdff dff_B_LEZjdAOF2_0(.din(n9877), .dout(n9880));
    jdff dff_B_K5gxWMxw9_0(.din(n9880), .dout(n9883));
    jdff dff_B_jhGhSjXn1_0(.din(n9883), .dout(n9886));
    jdff dff_B_XXn0nBBT4_0(.din(n9886), .dout(n9889));
    jdff dff_B_8XvexMbO0_0(.din(n9889), .dout(n9892));
    jdff dff_B_k5ROGEeQ9_0(.din(n9892), .dout(n9895));
    jdff dff_B_dPS8gKbJ3_0(.din(n9895), .dout(n9898));
    jdff dff_B_Mqwo4kXx0_0(.din(n9898), .dout(n9901));
    jdff dff_B_tgwF8Qzt1_0(.din(n9901), .dout(n9904));
    jdff dff_B_fUQ7IRTy5_0(.din(n9904), .dout(n9907));
    jdff dff_A_YxLnYYPV2_1(.din(n16125), .dout(n9909));
    jdff dff_A_wZ5mTor86_2(.din(n16125), .dout(n9912));
    jdff dff_B_FIoheWbs5_2(.din(G70), .dout(n9916));
    jdff dff_B_IGq84fdi5_1(.din(n3298), .dout(n9919));
    jdff dff_B_Y32ShMuw6_1(.din(n9919), .dout(n9922));
    jdff dff_B_hPqcY2iD9_1(.din(n9922), .dout(n9925));
    jdff dff_A_3W4kvWNZ3_2(.din(n9930), .dout(n9927));
    jdff dff_A_nMHJbxjT1_2(.din(n15960), .dout(n9930));
    jdff dff_B_ZVmm8MNS6_0(.din(n3358), .dout(n9934));
    jdff dff_B_0A3Ro9nz0_0(.din(n9934), .dout(n9937));
    jdff dff_B_ep9uS0Mf1_0(.din(n9937), .dout(n9940));
    jdff dff_B_3aDHVfrs0_0(.din(n9940), .dout(n9943));
    jdff dff_B_ujgqR1BA0_0(.din(n9943), .dout(n9946));
    jdff dff_B_Lpe4bac67_0(.din(n9946), .dout(n9949));
    jdff dff_B_qqefWXnl8_0(.din(n9949), .dout(n9952));
    jdff dff_B_2YvTkKCA9_0(.din(n9952), .dout(n9955));
    jdff dff_B_kWAgN8za5_0(.din(n9955), .dout(n9958));
    jdff dff_B_h2W2eMv27_0(.din(n9958), .dout(n9961));
    jdff dff_B_eYQWpjpO9_0(.din(n9961), .dout(n9964));
    jdff dff_B_u2gv6qbn2_0(.din(n9964), .dout(n9967));
    jdff dff_B_65GFBJ5i0_0(.din(n9967), .dout(n9970));
    jdff dff_B_1S2oHxRv6_0(.din(n9970), .dout(n9973));
    jdff dff_B_n4Z3kC0B8_0(.din(n9973), .dout(n9976));
    jdff dff_B_69LkdRe29_0(.din(n3354), .dout(n9979));
    jdff dff_B_BFLz6QQE7_1(.din(n3334), .dout(n9982));
    jdff dff_B_WEtm194H6_0(.din(n3394), .dout(n9985));
    jdff dff_B_7IBwxlQT2_0(.din(n9985), .dout(n9988));
    jdff dff_B_HnBuq4GM7_0(.din(n9988), .dout(n9991));
    jdff dff_B_j0gK1YOY6_0(.din(n9991), .dout(n9994));
    jdff dff_B_817Q2Pqi5_0(.din(n9994), .dout(n9997));
    jdff dff_B_J9CF1wra9_0(.din(n9997), .dout(n10000));
    jdff dff_B_rC1cw62D8_0(.din(n10000), .dout(n10003));
    jdff dff_B_xWmwhYEu5_0(.din(n10003), .dout(n10006));
    jdff dff_B_NAUXOCim6_0(.din(n10006), .dout(n10009));
    jdff dff_B_NeoQELkz9_0(.din(n10009), .dout(n10012));
    jdff dff_B_nsN7kUO77_0(.din(n10012), .dout(n10015));
    jdff dff_B_Fo0Afh4i9_0(.din(n10015), .dout(n10018));
    jdff dff_B_44vAecWO2_0(.din(n3390), .dout(n10021));
    jdff dff_B_jYDj2gId5_0(.din(n3378), .dout(n10024));
    jdff dff_A_sc3jI8Q69_0(.din(n10029), .dout(n10026));
    jdff dff_A_ojvfwOxf9_0(.din(n10032), .dout(n10029));
    jdff dff_A_RUcvG7n60_0(.din(n13492), .dout(n10032));
    jdff dff_A_ax7OvO1A0_1(.din(n10038), .dout(n10035));
    jdff dff_A_1tEDy0cf0_1(.din(n10041), .dout(n10038));
    jdff dff_A_By1RKrdX8_1(.din(n10044), .dout(n10041));
    jdff dff_A_DC7nCXXN2_1(.din(n10047), .dout(n10044));
    jdff dff_A_sjV8SmEY9_1(.din(n10050), .dout(n10047));
    jdff dff_A_eihDuhsQ7_1(.din(n10053), .dout(n10050));
    jdff dff_A_ex2SzdNi7_1(.din(n13492), .dout(n10053));
    jdff dff_A_xXCSNQrE9_0(.din(n10059), .dout(n10056));
    jdff dff_A_NbS7Alik6_0(.din(n10062), .dout(n10059));
    jdff dff_A_FPGa4Tmv5_0(.din(n10065), .dout(n10062));
    jdff dff_A_4mEEVqk35_0(.din(n10068), .dout(n10065));
    jdff dff_A_BNuCiqWE6_0(.din(n16689), .dout(n10068));
    jdff dff_A_gyXkKqaX3_1(.din(n10074), .dout(n10071));
    jdff dff_A_0fZTBHr02_1(.din(n10077), .dout(n10074));
    jdff dff_A_If7SqYPf4_1(.din(n10080), .dout(n10077));
    jdff dff_A_9DpGzOIF8_1(.din(n10083), .dout(n10080));
    jdff dff_A_mKOuAFjK0_1(.din(n10086), .dout(n10083));
    jdff dff_A_L7SHkB7f7_1(.din(n10089), .dout(n10086));
    jdff dff_A_NmeBqJej4_1(.din(n16689), .dout(n10089));
    jdff dff_B_DqTLLdrs8_0(.din(n3430), .dout(n10093));
    jdff dff_B_Hg05mqed6_0(.din(n10093), .dout(n10096));
    jdff dff_B_4C7GlDBG1_0(.din(n10096), .dout(n10099));
    jdff dff_B_O1iGWmKO3_0(.din(n10099), .dout(n10102));
    jdff dff_B_uIzJ5YwN7_0(.din(n10102), .dout(n10105));
    jdff dff_B_DWi30R3v4_0(.din(n10105), .dout(n10108));
    jdff dff_B_DzHoF0Ho2_0(.din(n10108), .dout(n10111));
    jdff dff_B_6vc9JUTF5_0(.din(n10111), .dout(n10114));
    jdff dff_B_ipExecNx7_0(.din(n10114), .dout(n10117));
    jdff dff_B_IGY9THnU3_0(.din(n10117), .dout(n10120));
    jdff dff_B_dvbZwwhr3_0(.din(n10120), .dout(n10123));
    jdff dff_B_0gPtaQdm0_0(.din(n10123), .dout(n10126));
    jdff dff_B_u5p460Ly0_0(.din(n3426), .dout(n10129));
    jdff dff_B_vv2nfHoo5_1(.din(n3406), .dout(n10132));
    jdff dff_A_Z1lAP6kb0_2(.din(n10137), .dout(n10134));
    jdff dff_A_OZ82CCvQ3_2(.din(n10140), .dout(n10137));
    jdff dff_A_snODAuqc6_2(.din(n10677), .dout(n10140));
    jdff dff_B_q1kALwgv4_0(.din(n3466), .dout(n10144));
    jdff dff_B_Akr5dmJX1_0(.din(n10144), .dout(n10147));
    jdff dff_B_voAJ6e0B4_0(.din(n10147), .dout(n10150));
    jdff dff_B_LbmON4d04_0(.din(n10150), .dout(n10153));
    jdff dff_B_czf60rpt0_0(.din(n10153), .dout(n10156));
    jdff dff_B_OtENGNYd1_0(.din(n10156), .dout(n10159));
    jdff dff_B_6pjDQfW88_0(.din(n10159), .dout(n10162));
    jdff dff_B_nIM3frMz3_0(.din(n10162), .dout(n10165));
    jdff dff_B_sumYEOPg6_0(.din(n10165), .dout(n10168));
    jdff dff_B_wKto22uR8_0(.din(n10168), .dout(n10171));
    jdff dff_B_83oAMUNY6_0(.din(n10171), .dout(n10174));
    jdff dff_B_0ovZIQyE8_0(.din(n10174), .dout(n10177));
    jdff dff_B_DHFhcBXc5_0(.din(n10177), .dout(n10180));
    jdff dff_B_sFCOBFKZ8_0(.din(n3462), .dout(n10183));
    jdff dff_A_YrGfyymj5_0(.din(n10188), .dout(n10185));
    jdff dff_A_gamMfp6T9_0(.din(n16584), .dout(n10188));
    jdff dff_A_iXDsf0Av2_1(.din(n16584), .dout(n10191));
    jdff dff_B_d44rBEZQ4_1(.din(n3478), .dout(n10195));
    jdff dff_B_hLhYhoOa3_1(.din(n10195), .dout(n10198));
    jdff dff_B_Kq7EokUD6_1(.din(n10198), .dout(n10201));
    jdff dff_B_nSl6TPh82_1(.din(n10201), .dout(n10204));
    jdff dff_B_dWZPMxOD5_1(.din(n10204), .dout(n10207));
    jdff dff_B_vhe6go5h3_1(.din(n10207), .dout(n10210));
    jdff dff_B_VPO1xM0b1_1(.din(n10210), .dout(n10213));
    jdff dff_B_xl4fjvn14_1(.din(n10213), .dout(n10216));
    jdff dff_B_prMlvip00_1(.din(n10216), .dout(n10219));
    jdff dff_B_lB19PUY14_1(.din(n10219), .dout(n10222));
    jdff dff_B_fW7CWBUT3_1(.din(n10222), .dout(n10225));
    jdff dff_B_2bYdIWHR2_1(.din(n10225), .dout(n10228));
    jdff dff_B_QlE12RLM6_1(.din(n10228), .dout(n10231));
    jdff dff_B_lc1B8HQ97_1(.din(n10231), .dout(n10234));
    jdff dff_B_8HXiJ17M2_1(.din(n10234), .dout(n10237));
    jdff dff_B_IbNvrrdT9_1(.din(n10237), .dout(n10240));
    jdff dff_B_4rKzi5ft5_1(.din(n10240), .dout(n10243));
    jdff dff_B_hr4RBaw75_1(.din(n3482), .dout(n10246));
    jdff dff_B_JPTkieWH6_1(.din(n10246), .dout(n10249));
    jdff dff_B_JFrPKMCF7_1(.din(n10249), .dout(n10252));
    jdff dff_B_6bJ5mfPR9_1(.din(n10252), .dout(n10255));
    jdff dff_B_HLYyn1f77_1(.din(n10255), .dout(n10258));
    jdff dff_B_7YKmGSuK7_1(.din(n10258), .dout(n10261));
    jdff dff_B_7lvApMHE8_1(.din(n10261), .dout(n10264));
    jdff dff_B_ONpsITEh0_1(.din(n10264), .dout(n10267));
    jdff dff_B_9P3iOI6n7_1(.din(n10267), .dout(n10270));
    jdff dff_B_RWnyobUg6_1(.din(n10270), .dout(n10273));
    jdff dff_B_KZoARXLc0_1(.din(n10273), .dout(n10276));
    jdff dff_B_FqkfDwMg0_1(.din(n10276), .dout(n10279));
    jdff dff_B_IDc6rDxQ2_1(.din(n10279), .dout(n10282));
    jdff dff_B_URZBSOEB9_1(.din(n10282), .dout(n10285));
    jdff dff_B_mgwEUQS91_1(.din(n10285), .dout(n10288));
    jdff dff_B_sRWC0tdv5_1(.din(n10288), .dout(n10291));
    jdff dff_B_dzFlQmzL4_1(.din(n10291), .dout(n10294));
    jdff dff_B_tuaV0hrY5_1(.din(n2230), .dout(n10297));
    jdff dff_B_j17Q7vPS0_1(.din(n10297), .dout(n10300));
    jdff dff_B_Li0bAqfx2_1(.din(n10300), .dout(n10303));
    jdff dff_B_4DN8KS018_1(.din(n10303), .dout(n10306));
    jdff dff_B_T3Kapml73_1(.din(n10306), .dout(n10309));
    jdff dff_B_H7MzAnXL8_1(.din(n10309), .dout(n10312));
    jdff dff_B_erHClltW3_1(.din(n10312), .dout(n10315));
    jdff dff_B_VRr48Sni9_1(.din(n10315), .dout(n10318));
    jdff dff_B_GjJOhlnr9_1(.din(n10318), .dout(n10321));
    jdff dff_B_YaNA41sQ1_1(.din(n10321), .dout(n10324));
    jdff dff_B_cuEdzt2S1_0(.din(n2302), .dout(n10327));
    jdff dff_B_LPgtyoLW5_0(.din(n10327), .dout(n10330));
    jdff dff_B_uYNAnF3P9_0(.din(n10330), .dout(n10333));
    jdff dff_B_TTI3V0c07_0(.din(n10333), .dout(n10336));
    jdff dff_B_0LeQCjqX9_0(.din(n10336), .dout(n10339));
    jdff dff_B_hGo6aE1L4_0(.din(n10339), .dout(n10342));
    jdff dff_B_vrHzVBPs5_1(.din(n818), .dout(n10345));
    jdff dff_B_8P1YGzgQ2_1(.din(n799), .dout(n10348));
    jdff dff_B_Quo6qYtP7_1(.din(n2271), .dout(n10351));
    jdff dff_B_oUcrpXRb4_1(.din(n10351), .dout(n10354));
    jdff dff_B_vAZPEblA7_1(.din(n10354), .dout(n10357));
    jdff dff_B_iQPIcCBI1_1(.din(n10357), .dout(n10360));
    jdff dff_B_qwPBKtuU9_1(.din(n10360), .dout(n10363));
    jdff dff_B_7ursiyCr0_1(.din(G52), .dout(n10366));
    jdff dff_B_9EyVRvmn8_1(.din(n10366), .dout(n10369));
    jdff dff_B_DUiIQvWy4_1(.din(n2433), .dout(n10372));
    jdff dff_B_WTgw8wve6_1(.din(n10372), .dout(n10375));
    jdff dff_B_7O6ie4Ck9_1(.din(n10375), .dout(n10378));
    jdff dff_B_Ni0PLMRt2_1(.din(n10378), .dout(n10381));
    jdff dff_B_VfuJOKvu7_1(.din(n10381), .dout(n10384));
    jdff dff_B_ujPWr6ve6_1(.din(n10384), .dout(n10387));
    jdff dff_B_rbAuemPE9_1(.din(n10387), .dout(n10390));
    jdff dff_B_3TGk4T0w7_1(.din(n10390), .dout(n10393));
    jdff dff_B_ZBum0YOh9_1(.din(n10393), .dout(n10396));
    jdff dff_B_mRm8lSLm3_1(.din(n10396), .dout(n10399));
    jdff dff_B_FXetr5Jf8_0(.din(n2471), .dout(n10402));
    jdff dff_B_bj1sZqhK9_0(.din(n10402), .dout(n10405));
    jdff dff_B_ZzupltTq5_0(.din(n10405), .dout(n10408));
    jdff dff_B_RCQ0KC3s0_0(.din(n10408), .dout(n10411));
    jdff dff_B_PbjgCsSE0_0(.din(n10411), .dout(n10414));
    jdff dff_B_ZIzc92Bh0_0(.din(n10414), .dout(n10417));
    jdff dff_B_AKBIMfoM4_1(.din(n914), .dout(n10420));
    jdff dff_B_VkR0RJnO3_1(.din(n895), .dout(n10423));
    jdff dff_B_YoXDgICp1_1(.din(G122), .dout(n10426));
    jdff dff_B_7UNUH5rp2_1(.din(n10426), .dout(n10429));
    jdff dff_B_o2AF7ZD13_2(.din(G170), .dout(n10432));
    jdff dff_B_kgOnxlfu9_2(.din(G200), .dout(n10435));
    jdff dff_B_O2epEFNI8_2(.din(n10435), .dout(n10438));
    jdff dff_B_zdIME7Wv5_0(.din(n3538), .dout(n10441));
    jdff dff_B_0t4XAYSf0_0(.din(n10441), .dout(n10444));
    jdff dff_B_kdRm8gLu1_0(.din(n10444), .dout(n10447));
    jdff dff_B_M5D640MM2_0(.din(n10447), .dout(n10450));
    jdff dff_B_TnHaRBC44_0(.din(n10450), .dout(n10453));
    jdff dff_B_2hFp0IYO8_0(.din(n10453), .dout(n10456));
    jdff dff_B_D4dwODuW2_0(.din(n10456), .dout(n10459));
    jdff dff_B_bUX2u2H59_0(.din(n10459), .dout(n10462));
    jdff dff_B_9KqjEjrP8_0(.din(n10462), .dout(n10465));
    jdff dff_B_7o2KHG086_0(.din(n10465), .dout(n10468));
    jdff dff_B_oQ8gKiWd9_0(.din(n10468), .dout(n10471));
    jdff dff_B_9vShPgtL7_0(.din(n10471), .dout(n10474));
    jdff dff_B_iKYzvaD16_0(.din(n3534), .dout(n10477));
    jdff dff_B_SJjDmDZT6_2(.din(G158), .dout(n10480));
    jdff dff_B_bsAacwTI8_2(.din(G188), .dout(n10483));
    jdff dff_B_K9zwZyi23_2(.din(n10483), .dout(n10486));
    jdff dff_B_metFiBlD4_0(.din(n3522), .dout(n10489));
    jdff dff_B_XEBaaWNY0_1(.din(n2560), .dout(n10492));
    jdff dff_B_cWW7BqkY5_1(.din(n10492), .dout(n10495));
    jdff dff_B_FT55muRm4_1(.din(n10495), .dout(n10498));
    jdff dff_B_P2bFHe5K8_1(.din(n10498), .dout(n10501));
    jdff dff_B_4UIEkQYb6_1(.din(n10501), .dout(n10504));
    jdff dff_B_VwpLRZYF3_1(.din(n10504), .dout(n10507));
    jdff dff_B_GtsUyFiA0_0(.din(n2587), .dout(n10510));
    jdff dff_B_S49bTiMW9_0(.din(n10510), .dout(n10513));
    jdff dff_B_RLUsb3Cv4_1(.din(n956), .dout(n10516));
    jdff dff_B_z12meKbH6_1(.din(n937), .dout(n10519));
    jdff dff_A_0VM845kW6_0(.din(n10524), .dout(n10521));
    jdff dff_A_EsAjOgU65_0(.din(n2575), .dout(n10524));
    jdff dff_B_eJ69Mfy49_1(.din(n2563), .dout(n10528));
    jdff dff_B_uLwGAIUX9_1(.din(G126), .dout(n10531));
    jdff dff_B_PS2S0xBY7_1(.din(n10531), .dout(n10534));
    jdff dff_A_npS2ivQk8_0(.din(n14908), .dout(n10536));
    jdff dff_A_IqrBrl157_1(.din(n10542), .dout(n10539));
    jdff dff_A_U4fR8iQ06_1(.din(n10545), .dout(n10542));
    jdff dff_A_2xgFELTQ7_1(.din(n10548), .dout(n10545));
    jdff dff_A_tGcLAQFM9_1(.din(n10551), .dout(n10548));
    jdff dff_A_CX0tG5144_1(.din(n10554), .dout(n10551));
    jdff dff_A_6u7w5u6X9_1(.din(n14908), .dout(n10554));
    jdff dff_B_tlusE0j86_1(.din(n2047), .dout(n10558));
    jdff dff_B_sWwHpGJt0_1(.din(n10558), .dout(n10561));
    jdff dff_B_GuCnLKnr4_1(.din(n10561), .dout(n10564));
    jdff dff_B_4J9ddOpI5_1(.din(n10564), .dout(n10567));
    jdff dff_B_HlcYQuNT3_1(.din(n10567), .dout(n10570));
    jdff dff_B_c1L8sULW9_1(.din(n10570), .dout(n10573));
    jdff dff_B_p49FRbal8_1(.din(n10573), .dout(n10576));
    jdff dff_B_ZbyInzDL9_1(.din(n10576), .dout(n10579));
    jdff dff_B_iVd2sr9e1_0(.din(n2089), .dout(n10582));
    jdff dff_B_yRqSM7OQ3_0(.din(n10582), .dout(n10585));
    jdff dff_B_LoDdlt7O8_0(.din(n10585), .dout(n10588));
    jdff dff_B_HGmizWoM4_0(.din(n10588), .dout(n10591));
    jdff dff_B_oZOwAB332_1(.din(n595), .dout(n10594));
    jdff dff_B_hamSiRHx7_1(.din(n573), .dout(n10597));
    jdff dff_B_5IjkzF0r0_0(.din(n2073), .dout(n10600));
    jdff dff_B_7wNVapkp3_0(.din(n10600), .dout(n10603));
    jdff dff_B_kJmmPrrk2_0(.din(n10603), .dout(n10606));
    jdff dff_B_vFdVfgzK6_0(.din(n10606), .dout(n10609));
    jdff dff_A_B0xsdXZn9_0(.din(n10614), .dout(n10611));
    jdff dff_A_OTKIU66v7_0(.din(n10617), .dout(n10614));
    jdff dff_A_YV5OdHI91_0(.din(n10620), .dout(n10617));
    jdff dff_A_PPiBdDlg1_0(.din(n10623), .dout(n10620));
    jdff dff_A_xrLt9rQJ6_0(.din(n11089), .dout(n10623));
    jdff dff_A_TwveDcUk1_0(.din(n10629), .dout(n10626));
    jdff dff_A_YM1cTB718_0(.din(n10632), .dout(n10629));
    jdff dff_A_5cmZxVG40_0(.din(n10635), .dout(n10632));
    jdff dff_A_9W5ELkMv7_0(.din(n10638), .dout(n10635));
    jdff dff_A_xhrFUx5g6_0(.din(n19764), .dout(n10638));
    jdff dff_A_K8kkhlAe6_2(.din(n10644), .dout(n10641));
    jdff dff_A_dO3Ntust9_2(.din(n10647), .dout(n10644));
    jdff dff_A_2hM6Ucfa7_2(.din(n19764), .dout(n10647));
    jdff dff_B_tGjzBN9i0_1(.din(G129), .dout(n10651));
    jdff dff_B_NJuNj2kG9_1(.din(n10651), .dout(n10654));
    jdff dff_A_NnsPrOqX9_1(.din(n10659), .dout(n10656));
    jdff dff_A_qQP3m4jI7_1(.din(n10662), .dout(n10659));
    jdff dff_A_0NMZDrI95_1(.din(n10665), .dout(n10662));
    jdff dff_A_gGGJZbzA5_1(.din(n10671), .dout(n10665));
    jdff dff_A_GGM1gy4q7_2(.din(n10671), .dout(n10668));
    jdff dff_A_D9Wcx2QM8_0(.din(n10674), .dout(n10671));
    jdff dff_A_vfZVX75W4_0(.din(n20757), .dout(n10674));
    jdff dff_A_bdDwh1Wl4_1(.din(n10680), .dout(n10677));
    jdff dff_A_Jw5QYtyr4_1(.din(n20757), .dout(n10680));
    jdff dff_B_CUT3gRE58_0(.din(n3574), .dout(n10684));
    jdff dff_B_bWLS9a6V2_0(.din(n10684), .dout(n10687));
    jdff dff_B_vI2VsaJz9_0(.din(n10687), .dout(n10690));
    jdff dff_B_zGKyLPLR5_0(.din(n10690), .dout(n10693));
    jdff dff_B_0XECho6T1_0(.din(n10693), .dout(n10696));
    jdff dff_B_0ZMRQjxo5_0(.din(n10696), .dout(n10699));
    jdff dff_B_Ce7ze7A05_0(.din(n10699), .dout(n10702));
    jdff dff_B_04LfTljs7_0(.din(n10702), .dout(n10705));
    jdff dff_B_5FLfSNxX5_0(.din(n10705), .dout(n10708));
    jdff dff_B_E4IgnFj56_0(.din(n10708), .dout(n10711));
    jdff dff_B_0spYFI720_0(.din(n10711), .dout(n10714));
    jdff dff_B_0FbXlvoh7_0(.din(n10714), .dout(n10717));
    jdff dff_B_kwmSNrEv6_0(.din(n3570), .dout(n10720));
    jdff dff_B_8AGxI0Mu5_2(.din(G152), .dout(n10723));
    jdff dff_B_ASVoifaa9_2(.din(G155), .dout(n10726));
    jdff dff_B_Ajmd820Z0_2(.din(n10726), .dout(n10729));
    jdff dff_B_EFBbqyKg0_1(.din(n3550), .dout(n10732));
    jdff dff_B_NuMGKBgK4_1(.din(n2521), .dout(n10735));
    jdff dff_B_fIKJ2Mgp5_1(.din(n10735), .dout(n10738));
    jdff dff_B_d4z54aPe4_1(.din(n10738), .dout(n10741));
    jdff dff_B_MylFQXjh9_1(.din(n10741), .dout(n10744));
    jdff dff_B_hWOXd6XA6_1(.din(n10744), .dout(n10747));
    jdff dff_B_Periazxo7_1(.din(n10747), .dout(n10750));
    jdff dff_B_9P4ED7zy1_1(.din(n10750), .dout(n10753));
    jdff dff_B_U8M86RnQ3_0(.din(n2545), .dout(n10756));
    jdff dff_B_gBzeg0a72_0(.din(n10756), .dout(n10759));
    jdff dff_B_I1dON0uH7_0(.din(n10759), .dout(n10762));
    jdff dff_B_ugITFTmU9_1(.din(n1002), .dout(n10765));
    jdff dff_B_ybO4WRJc4_1(.din(n983), .dout(n10768));
    jdff dff_B_8U0Oim1p9_1(.din(G127), .dout(n10771));
    jdff dff_B_l6Ij8nIr3_1(.din(n10771), .dout(n10774));
    jdff dff_B_CG8aC8g90_1(.din(n2352), .dout(n10777));
    jdff dff_B_onHZEBtR5_1(.din(n10777), .dout(n10780));
    jdff dff_B_B3Sll7g45_1(.din(n10780), .dout(n10783));
    jdff dff_B_HHaPyPg73_1(.din(n10783), .dout(n10786));
    jdff dff_B_fieNrXQD7_1(.din(n10786), .dout(n10789));
    jdff dff_B_BFd0Oyoi6_1(.din(n10789), .dout(n10792));
    jdff dff_B_Pg0Xh79Q8_1(.din(n10792), .dout(n10795));
    jdff dff_B_8rQ7rliv3_1(.din(n2356), .dout(n10798));
    jdff dff_B_LxXzK1Q48_1(.din(n10798), .dout(n10801));
    jdff dff_B_OEziAhiQ8_1(.din(n10801), .dout(n10804));
    jdff dff_B_sStGSEa44_1(.din(n10804), .dout(n10807));
    jdff dff_A_SwyMxSwn5_0(.din(n10812), .dout(n10809));
    jdff dff_A_K1FPsr598_0(.din(n10815), .dout(n10812));
    jdff dff_A_FL9tvQGF9_0(.din(n10818), .dout(n10815));
    jdff dff_A_yezpWkaN3_0(.din(n10821), .dout(n10818));
    jdff dff_A_3lqhmAhK7_0(.din(n2368), .dout(n10821));
    jdff dff_B_90WGFX200_1(.din(n637), .dout(n10825));
    jdff dff_B_WTvEmP2Q3_1(.din(n618), .dout(n10828));
    jdff dff_B_gCPz57zM4_1(.din(G119), .dout(n10831));
    jdff dff_B_7640OupI3_1(.din(n10831), .dout(n10834));
    jdff dff_B_RnR6lCWr1_0(.din(n3610), .dout(n10837));
    jdff dff_B_bk9oqwj17_0(.din(n10837), .dout(n10840));
    jdff dff_B_zjR3F0PZ6_0(.din(n10840), .dout(n10843));
    jdff dff_B_uAVllWra0_0(.din(n10843), .dout(n10846));
    jdff dff_B_RU9gjels2_0(.din(n10846), .dout(n10849));
    jdff dff_B_vNbCm1wf4_0(.din(n10849), .dout(n10852));
    jdff dff_B_sczV63Oz7_0(.din(n10852), .dout(n10855));
    jdff dff_B_TU8pH5Wq5_0(.din(n10855), .dout(n10858));
    jdff dff_B_pA0nuJHF3_0(.din(n10858), .dout(n10861));
    jdff dff_B_iecZB5iN5_0(.din(n10861), .dout(n10864));
    jdff dff_B_EaveTiGR9_0(.din(n10864), .dout(n10867));
    jdff dff_B_I7cht51M1_0(.din(n10867), .dout(n10870));
    jdff dff_B_MEIhhaKH4_0(.din(n10870), .dout(n10873));
    jdff dff_B_l83lBKCX4_0(.din(n3606), .dout(n10876));
    jdff dff_B_ZI5yvDHv8_2(.din(G146), .dout(n10879));
    jdff dff_B_BiHPPjJQ1_2(.din(G149), .dout(n10882));
    jdff dff_B_t5CF08rg6_2(.din(n10882), .dout(n10885));
    jdff dff_B_UXzmJdT80_1(.din(n2486), .dout(n10888));
    jdff dff_B_gGE7O5iU9_1(.din(n10888), .dout(n10891));
    jdff dff_B_hU0SneQp0_1(.din(n10891), .dout(n10894));
    jdff dff_B_VzT1cfgR9_1(.din(n10894), .dout(n10897));
    jdff dff_B_I7I4M44f4_1(.din(n10897), .dout(n10900));
    jdff dff_B_3lXXAADx3_1(.din(n10900), .dout(n10903));
    jdff dff_B_GTMGHZwB8_1(.din(n10903), .dout(n10906));
    jdff dff_B_c9O17rgw7_1(.din(n10906), .dout(n10909));
    jdff dff_B_Ej5h7qih9_0(.din(n2506), .dout(n10912));
    jdff dff_B_KpAM97bC1_0(.din(n10912), .dout(n10915));
    jdff dff_B_h8VxbfjI7_0(.din(n10915), .dout(n10918));
    jdff dff_B_wazcHJKO4_0(.din(n10918), .dout(n10921));
    jdff dff_B_Ib7fXhQc1_1(.din(n1136), .dout(n10924));
    jdff dff_B_kZQ8zMyd6_1(.din(n1117), .dout(n10927));
    jdff dff_A_rNiPtXLH8_2(.din(n10932), .dout(n10929));
    jdff dff_A_3aedCEev1_2(.din(n10935), .dout(n10932));
    jdff dff_A_QMPVijS82_2(.din(n15348), .dout(n10935));
    jdff dff_A_GZeO6MGe9_0(.din(n10941), .dout(n10938));
    jdff dff_A_0WMH8yzG8_0(.din(n10944), .dout(n10941));
    jdff dff_A_cdAeYYAu1_0(.din(n10947), .dout(n10944));
    jdff dff_A_bIIZgxBS9_0(.din(n10950), .dout(n10947));
    jdff dff_A_Pp1HGQRd6_0(.din(n2494), .dout(n10950));
    jdff dff_A_za0xKMAC7_1(.din(n19824), .dout(n10953));
    jdff dff_A_7WVyANtA8_2(.din(n10959), .dout(n10956));
    jdff dff_A_Yv7YRBAz8_2(.din(n19824), .dout(n10959));
    jdff dff_B_u4wgZrrl9_1(.din(G128), .dout(n10963));
    jdff dff_B_e7Aq2xOM1_1(.din(n10963), .dout(n10966));
    jdff dff_A_0V2656ta9_0(.din(n10971), .dout(n10968));
    jdff dff_A_QiqEtPaT6_0(.din(n20163), .dout(n10971));
    jdff dff_A_LWUS1reT6_1(.din(n20163), .dout(n10974));
    jdff dff_B_l3iQHOaA7_1(.din(n2317), .dout(n10978));
    jdff dff_B_2JDzgvY80_1(.din(n10978), .dout(n10981));
    jdff dff_B_X9qMtqnv1_1(.din(n10981), .dout(n10984));
    jdff dff_B_Y1iIcmNt6_1(.din(n10984), .dout(n10987));
    jdff dff_B_0f47Wv3m5_1(.din(n10987), .dout(n10990));
    jdff dff_B_At1YA5Vh4_1(.din(n10990), .dout(n10993));
    jdff dff_B_lJZSXHvj7_1(.din(n10993), .dout(n10996));
    jdff dff_B_m1rdW9ar1_1(.din(n10996), .dout(n10999));
    jdff dff_B_BQ2EQVOl9_1(.din(n10999), .dout(n11002));
    jdff dff_B_1iNS7Nap6_0(.din(n2337), .dout(n11005));
    jdff dff_B_eMTh1SQH4_0(.din(n11005), .dout(n11008));
    jdff dff_B_SXzXfOxQ5_0(.din(n11008), .dout(n11011));
    jdff dff_B_LDLs90Uk8_0(.din(n11011), .dout(n11014));
    jdff dff_B_heqfmxww4_0(.din(n11014), .dout(n11017));
    jdff dff_B_G225qpP34_0(.din(n11017), .dout(n11020));
    jdff dff_B_Sq3v5Xdh4_1(.din(n518), .dout(n11023));
    jdff dff_A_9JjDmRhG0_0(.din(n19716), .dout(n11025));
    jdff dff_A_7TidQJ6G5_1(.din(n19716), .dout(n11028));
    jdff dff_A_Q62aijYp6_0(.din(n19716), .dout(n11031));
    jdff dff_A_QcqzsMkw0_2(.din(n19716), .dout(n11034));
    jdff dff_A_QegbFgMH0_1(.din(n15363), .dout(n11037));
    jdff dff_A_fI6T211y3_2(.din(n15363), .dout(n11040));
    jdff dff_A_ORZgCVlI8_0(.din(n11046), .dout(n11043));
    jdff dff_A_7suQ0XYU3_0(.din(n11049), .dout(n11046));
    jdff dff_A_hAkS5YAw9_0(.din(n11052), .dout(n11049));
    jdff dff_A_d6GDjhyS9_0(.din(n11055), .dout(n11052));
    jdff dff_A_97sd9oJa1_0(.din(n11058), .dout(n11055));
    jdff dff_A_7ThD62w13_0(.din(n11061), .dout(n11058));
    jdff dff_A_V7JhJi4I3_0(.din(n2325), .dout(n11061));
    jdff dff_A_crg4mZyX4_1(.din(n11067), .dout(n11064));
    jdff dff_A_Xx2je7Ng9_1(.din(n11089), .dout(n11067));
    jdff dff_A_segWPjME5_2(.din(n11073), .dout(n11070));
    jdff dff_A_yIPwBlnh7_2(.din(n11076), .dout(n11073));
    jdff dff_A_dJn9XU4r0_2(.din(n11079), .dout(n11076));
    jdff dff_A_J9WMtu723_2(.din(n11082), .dout(n11079));
    jdff dff_A_eCToI8218_2(.din(n11089), .dout(n11082));
    jdff dff_B_gMSfxgK16_3(.din(n2013), .dout(n11086));
    jdff dff_B_KcNeIWmv8_3(.din(n11086), .dout(n11089));
    jdff dff_A_1TDZkw5D4_0(.din(n11094), .dout(n11091));
    jdff dff_A_UmKYnHNg0_0(.din(n11097), .dout(n11094));
    jdff dff_A_AlWs86Wg8_0(.din(n11100), .dout(n11097));
    jdff dff_A_vWLEkGRQ2_0(.din(n19740), .dout(n11100));
    jdff dff_A_dzVduUWR0_2(.din(n11106), .dout(n11103));
    jdff dff_A_PWGx2d8f6_2(.din(n11109), .dout(n11106));
    jdff dff_A_a58CEpQU8_2(.din(n19740), .dout(n11109));
    jdff dff_B_mjLra52h0_1(.din(G130), .dout(n11113));
    jdff dff_B_4LVBH2It6_1(.din(n11113), .dout(n11116));
    jdff dff_B_SJTCTUpE8_1(.din(n3628), .dout(n11119));
    jdff dff_B_0pq8b4099_1(.din(n11119), .dout(n11122));
    jdff dff_B_wP0WAYa06_1(.din(n11122), .dout(n11125));
    jdff dff_B_FfW8U1v00_1(.din(n11125), .dout(n11128));
    jdff dff_B_dw0eGgNd5_1(.din(n11128), .dout(n11131));
    jdff dff_B_BDi1Z0Wg1_1(.din(n11131), .dout(n11134));
    jdff dff_B_NK9pg6376_1(.din(n11134), .dout(n11137));
    jdff dff_B_gxIe1wTu2_1(.din(n11137), .dout(n11140));
    jdff dff_B_jhc8k3IX3_1(.din(n11140), .dout(n11143));
    jdff dff_B_yS83qBjv9_1(.din(n11143), .dout(n11146));
    jdff dff_B_JIjnueRV8_1(.din(n11146), .dout(n11149));
    jdff dff_B_262O5ZM97_1(.din(n11149), .dout(n11152));
    jdff dff_B_h34gSi9m2_1(.din(n11152), .dout(n11155));
    jdff dff_B_wujcZsIp8_1(.din(n11155), .dout(n11158));
    jdff dff_B_rzkQElNl3_1(.din(n11158), .dout(n11161));
    jdff dff_B_YehUqUFZ2_1(.din(n11161), .dout(n11164));
    jdff dff_B_yPIn38pH5_1(.din(n11164), .dout(n11167));
    jdff dff_B_IR1js6PY9_1(.din(n11167), .dout(n11170));
    jdff dff_B_p01T7xu26_1(.din(n3660), .dout(n11173));
    jdff dff_B_x2B1v9ul5_1(.din(n11173), .dout(n11176));
    jdff dff_B_9XDQ9MuK2_1(.din(n11176), .dout(n11179));
    jdff dff_B_6rxE4lJ27_1(.din(n11179), .dout(n11182));
    jdff dff_B_S5HSk2m91_1(.din(n11182), .dout(n11185));
    jdff dff_B_fBrT7Hht7_1(.din(n11185), .dout(n11188));
    jdff dff_B_LbGTneuH2_1(.din(n11188), .dout(n11191));
    jdff dff_B_TSoGnU751_1(.din(n11191), .dout(n11194));
    jdff dff_B_giGWtHgu2_1(.din(n11194), .dout(n11197));
    jdff dff_B_AcWpHut54_1(.din(n11197), .dout(n11200));
    jdff dff_B_Y2q2okYk1_0(.din(n3672), .dout(n11203));
    jdff dff_B_pma8W6UL3_0(.din(n11203), .dout(n11206));
    jdff dff_B_jifYEoLa5_0(.din(n11206), .dout(n11209));
    jdff dff_B_ZEnctCti8_0(.din(n11209), .dout(n11212));
    jdff dff_B_EmH8pxP01_0(.din(n11212), .dout(n11215));
    jdff dff_B_Naal926N0_0(.din(n11215), .dout(n11218));
    jdff dff_B_q67KMKMI6_0(.din(n11218), .dout(n11221));
    jdff dff_B_Gmtzc4x55_0(.din(n11221), .dout(n11224));
    jdff dff_B_gWjX512N1_0(.din(n11224), .dout(n11227));
    jdff dff_B_9K9OXY3N2_0(.din(n11227), .dout(n11230));
    jdff dff_B_HwYRXSb17_0(.din(n11230), .dout(n11233));
    jdff dff_B_8KOJ0rAh4_0(.din(n11233), .dout(n11236));
    jdff dff_B_aGH9xiGJ4_0(.din(n11236), .dout(n11239));
    jdff dff_B_oL3F66b33_0(.din(n11239), .dout(n11242));
    jdff dff_B_FuoDS0bO8_0(.din(n11242), .dout(n11245));
    jdff dff_B_REvoa9Uk5_0(.din(n11245), .dout(n11248));
    jdff dff_B_t6pHtrQy5_1(.din(n3635), .dout(n11251));
    jdff dff_B_dDzzxKxE0_1(.din(n11251), .dout(n11254));
    jdff dff_B_eTcQlCR77_1(.din(n11254), .dout(n11257));
    jdff dff_B_Txjh1bF79_1(.din(n3638), .dout(n11260));
    jdff dff_B_EEK85wo98_1(.din(n11260), .dout(n11263));
    jdff dff_B_e6rApPUh7_1(.din(n11263), .dout(n11266));
    jdff dff_B_0OOP1XMK4_1(.din(n11266), .dout(n11269));
    jdff dff_B_utxupP6v0_1(.din(n11269), .dout(n11272));
    jdff dff_B_fkywhnmy6_1(.din(n11272), .dout(n11275));
    jdff dff_A_qAfsH6ps1_0(.din(n11280), .dout(n11277));
    jdff dff_A_ka0Af7gB1_0(.din(n11283), .dout(n11280));
    jdff dff_A_Y7VtoUEM8_0(.din(n11286), .dout(n11283));
    jdff dff_A_vXaZmONx2_0(.din(n11289), .dout(n11286));
    jdff dff_A_3u8AhDZ50_0(.din(n11292), .dout(n11289));
    jdff dff_A_CBmTJGOR5_0(.din(n11295), .dout(n11292));
    jdff dff_A_2n1SrRKC7_0(.din(n11298), .dout(n11295));
    jdff dff_A_FdbRZcal4_0(.din(n11301), .dout(n11298));
    jdff dff_A_XpKbW4934_0(.din(n11304), .dout(n11301));
    jdff dff_A_WAbi9woj3_0(.din(n11307), .dout(n11304));
    jdff dff_A_q0KUU9WO9_0(.din(n11323), .dout(n11307));
    jdff dff_B_1JrkY8Dv8_2(.din(n3641), .dout(n11311));
    jdff dff_B_Ozu4KnEC0_2(.din(n11311), .dout(n11314));
    jdff dff_B_llg6wm2I2_2(.din(n11314), .dout(n11317));
    jdff dff_B_nGukN8y83_2(.din(n11317), .dout(n11320));
    jdff dff_B_eBuerXZk9_2(.din(n11320), .dout(n11323));
    jdff dff_A_yY3htEE00_0(.din(G3717), .dout(n11325));
    jdff dff_A_Spe8grpu6_1(.din(n770), .dout(n11328));
    jdff dff_A_ce82iF9C0_2(.din(n11334), .dout(n11331));
    jdff dff_A_bqmsRlfN6_2(.din(n11337), .dout(n11334));
    jdff dff_A_iymLysLC7_2(.din(n11340), .dout(n11337));
    jdff dff_A_nRGnI5Q08_2(.din(G3724), .dout(n11340));
    jdff dff_A_faYPsANX9_0(.din(n11346), .dout(n11343));
    jdff dff_A_IL6xpjDa7_0(.din(n11349), .dout(n11346));
    jdff dff_A_Q6I6sg426_0(.din(n11352), .dout(n11349));
    jdff dff_A_2ESL2CEo6_0(.din(n11355), .dout(n11352));
    jdff dff_A_ZDO7B8j88_0(.din(n11358), .dout(n11355));
    jdff dff_A_zyAtjveW0_0(.din(n11361), .dout(n11358));
    jdff dff_A_VihzxTqh9_0(.din(n11364), .dout(n11361));
    jdff dff_A_l1TPZ3Kj2_0(.din(n11367), .dout(n11364));
    jdff dff_A_zOHvRT210_0(.din(n11370), .dout(n11367));
    jdff dff_A_kjwlrNqP9_0(.din(n11373), .dout(n11370));
    jdff dff_A_HFFMZKXC4_0(.din(n3648), .dout(n11373));
    jdff dff_B_2ODW0byy4_1(.din(G132), .dout(n11377));
    jdff dff_B_bR5wdcvE0_1(.din(n11377), .dout(n11380));
    jdff dff_B_YCh1T0KM1_1(.din(n11380), .dout(n11383));
    jdff dff_B_WLeseU1z1_1(.din(n11383), .dout(n11386));
    jdff dff_B_GBcMuDia6_1(.din(n3816), .dout(n11389));
    jdff dff_B_9WsjWPI97_0(.din(n3831), .dout(n11392));
    jdff dff_B_PoXP9G9H8_0(.din(n11392), .dout(n11395));
    jdff dff_B_LH6zC8nH4_0(.din(n11395), .dout(n11398));
    jdff dff_B_N5kgZ4q98_0(.din(n11398), .dout(n11401));
    jdff dff_B_tam88bC02_0(.din(n3827), .dout(n11404));
    jdff dff_A_JmBuoIrZ9_0(.din(n11409), .dout(n11406));
    jdff dff_A_FtQ5RHRX1_0(.din(G559), .dout(n11409));
    jdff dff_B_lwgdiKd39_0(.din(n1688), .dout(n11413));
    jdff dff_B_Qa0kXc944_1(.din(n1668), .dout(n11416));
    jdff dff_B_gv7JNX2u5_1(.din(n2633), .dout(n11419));
    jdff dff_B_ArBKaFRb0_1(.din(n2637), .dout(n11422));
    jdff dff_B_GgwDVmIk2_0(.din(n2629), .dout(n11425));
    jdff dff_B_xLQe94xi2_1(.din(n2621), .dout(n11428));
    jdff dff_B_Y91lCFsy5_0(.din(G372), .dout(n11431));
    jdff dff_B_UpMQVbjd6_1(.din(n2605), .dout(n11434));
    jdff dff_B_jaZ47cMA7_1(.din(n2598), .dout(n11437));
    jdff dff_B_7xINs6mG3_1(.din(n11437), .dout(n11440));
    jdff dff_B_Y2yoSY4w4_0(.din(n3812), .dout(n11443));
    jdff dff_B_jOxmupOZ6_0(.din(n11443), .dout(n11446));
    jdff dff_B_yrPwA8uG8_0(.din(n11446), .dout(n11449));
    jdff dff_B_kSKAt8eF0_0(.din(n1727), .dout(n11452));
    jdff dff_B_HIzuN37p7_1(.din(n1703), .dout(n11455));
    jdff dff_A_J483ghBZ3_0(.din(n11460), .dout(n11457));
    jdff dff_A_R1I8Dhts8_0(.din(n11463), .dout(n11460));
    jdff dff_A_bXDUOtni8_0(.din(n11466), .dout(n11463));
    jdff dff_A_lTOzkCx56_0(.din(G245), .dout(n11466));
    jdff dff_B_Lkz0kzL29_1(.din(n2672), .dout(n11470));
    jdff dff_B_FTZIdq6L0_1(.din(n2688), .dout(n11473));
    jdff dff_B_WMbiIHUO3_1(.din(n11473), .dout(n11476));
    jdff dff_B_1GSiAlF65_1(.din(n2676), .dout(n11479));
    jdff dff_B_KzVdmX5f1_1(.din(G292), .dout(n11482));
    jdff dff_B_Eh8xcU5w1_1(.din(n3969), .dout(n11485));
    jdff dff_B_R6OPvu1m6_1(.din(n11485), .dout(n11488));
    jdff dff_B_tO5YvwMX9_1(.din(n11488), .dout(n11491));
    jdff dff_B_xTqVdMq19_1(.din(n11491), .dout(n11494));
    jdff dff_B_Yn23Ap934_1(.din(n11494), .dout(n11497));
    jdff dff_B_OUA70wuN8_1(.din(n11497), .dout(n11500));
    jdff dff_B_CHoghGGr2_1(.din(n11500), .dout(n11503));
    jdff dff_B_sRwG79PK9_1(.din(n11503), .dout(n11506));
    jdff dff_B_d0vPN1jU2_1(.din(n11506), .dout(n11509));
    jdff dff_B_XgTP2XRT7_1(.din(n11509), .dout(n11512));
    jdff dff_B_xF71wDdE2_1(.din(n11512), .dout(n11515));
    jdff dff_B_vUmjxWLO5_1(.din(n11515), .dout(n11518));
    jdff dff_B_Qv13RY871_1(.din(n11518), .dout(n11521));
    jdff dff_B_WLoJdSsh8_1(.din(n11521), .dout(n11524));
    jdff dff_B_blNbS6wX1_1(.din(n11524), .dout(n11527));
    jdff dff_B_Rh31UQkH5_1(.din(n11527), .dout(n11530));
    jdff dff_B_TT1moR132_1(.din(n11530), .dout(n11533));
    jdff dff_B_Ah0S6DeG2_1(.din(n11533), .dout(n11536));
    jdff dff_B_awItk95I5_1(.din(n11536), .dout(n11539));
    jdff dff_B_LVHBRYbN7_1(.din(n3957), .dout(n11542));
    jdff dff_B_RL3xREXt5_1(.din(n11542), .dout(n11545));
    jdff dff_A_bRwySmv44_2(.din(n11550), .dout(n11547));
    jdff dff_A_hIMjxelj8_2(.din(n11553), .dout(n11550));
    jdff dff_A_0YCsWJI95_2(.din(n11556), .dout(n11553));
    jdff dff_A_NdvFqruk6_2(.din(n11559), .dout(n11556));
    jdff dff_A_vBqxePfa1_2(.din(n11562), .dout(n11559));
    jdff dff_A_klTK2TIY7_2(.din(n11565), .dout(n11562));
    jdff dff_A_8gqaPvZ35_2(.din(n11568), .dout(n11565));
    jdff dff_A_T2fUFLh32_2(.din(n11571), .dout(n11568));
    jdff dff_A_eIaYIMDb1_2(.din(n11574), .dout(n11571));
    jdff dff_A_R2KmGRb39_2(.din(n11577), .dout(n11574));
    jdff dff_A_GbTFOAwC9_2(.din(n2387), .dout(n11577));
    jdff dff_A_Jn6agjht7_2(.din(n11583), .dout(n11580));
    jdff dff_A_zK74rVjF6_2(.din(n11586), .dout(n11583));
    jdff dff_A_WoT2ruqa0_2(.din(n11589), .dout(n11586));
    jdff dff_A_fgX5Exue9_2(.din(n11592), .dout(n11589));
    jdff dff_A_QtfeuDtX3_2(.din(n11595), .dout(n11592));
    jdff dff_A_NunGVhI32_2(.din(n11598), .dout(n11595));
    jdff dff_A_ZPlxwMdM3_2(.din(n11601), .dout(n11598));
    jdff dff_A_IMnj1xPy9_2(.din(n11604), .dout(n11601));
    jdff dff_A_5zXiPppJ4_2(.din(n11607), .dout(n11604));
    jdff dff_A_5VTLUQNs7_2(.din(n11610), .dout(n11607));
    jdff dff_A_6zJ0XKoK5_2(.din(n11613), .dout(n11610));
    jdff dff_A_NWM5yy8d4_2(.din(n11616), .dout(n11613));
    jdff dff_A_BePHHIG12_2(.din(n11619), .dout(n11616));
    jdff dff_A_SuyHfsP33_2(.din(G4089), .dout(n11619));
    jdff dff_B_WRpIyDKr5_0(.din(n4021), .dout(n11623));
    jdff dff_B_G6NOgQou0_0(.din(n11623), .dout(n11626));
    jdff dff_B_AsRt94t66_0(.din(n11626), .dout(n11629));
    jdff dff_B_xa0r5KoB9_0(.din(n11629), .dout(n11632));
    jdff dff_B_VOw4BDys5_0(.din(n11632), .dout(n11635));
    jdff dff_B_9tOouuU77_0(.din(n11635), .dout(n11638));
    jdff dff_B_GIuNXjbb3_0(.din(n11638), .dout(n11641));
    jdff dff_B_xoYDG25r2_0(.din(n11641), .dout(n11644));
    jdff dff_B_3MNhwztg4_0(.din(n11644), .dout(n11647));
    jdff dff_B_tooZ1f2L3_0(.din(n11647), .dout(n11650));
    jdff dff_B_97cH0skD7_0(.din(n11650), .dout(n11653));
    jdff dff_B_VZ8CXkyb1_0(.din(n11653), .dout(n11656));
    jdff dff_B_VFOFqvPb3_0(.din(n11656), .dout(n11659));
    jdff dff_B_yYWLHLHx1_0(.din(n11659), .dout(n11662));
    jdff dff_B_BXeoeUfm2_0(.din(n11662), .dout(n11665));
    jdff dff_B_G9lWqzGc2_0(.din(n11665), .dout(n11668));
    jdff dff_B_3VyOr7uT0_0(.din(n11668), .dout(n11671));
    jdff dff_B_Pdrz4BLb9_0(.din(n11671), .dout(n11674));
    jdff dff_B_oiuRAOfW1_0(.din(n11674), .dout(n11677));
    jdff dff_B_oDyragN69_0(.din(n11677), .dout(n11680));
    jdff dff_B_VNDVWmfp6_0(.din(n11680), .dout(n11683));
    jdff dff_B_ysMN1GsA7_2(.din(G106), .dout(n11686));
    jdff dff_B_kPe973K11_1(.din(n3993), .dout(n11689));
    jdff dff_B_gFIIPHp96_1(.din(n11689), .dout(n11692));
    jdff dff_A_lNU0yOKL0_0(.din(n11697), .dout(n11694));
    jdff dff_A_5oygKVDc0_0(.din(n11700), .dout(n11697));
    jdff dff_A_Oj3gjdpi9_0(.din(n11703), .dout(n11700));
    jdff dff_A_9heJPZ8k6_0(.din(n11706), .dout(n11703));
    jdff dff_A_fGTiVtRK4_0(.din(n11709), .dout(n11706));
    jdff dff_A_nQQgaYQw0_0(.din(n11712), .dout(n11709));
    jdff dff_A_YLZyl7P60_0(.din(n11715), .dout(n11712));
    jdff dff_A_Moh6W1In2_0(.din(n11718), .dout(n11715));
    jdff dff_A_PMi9rjUu8_0(.din(n11721), .dout(n11718));
    jdff dff_A_ZKnW40b80_0(.din(n11724), .dout(n11721));
    jdff dff_A_Z8AzZGpY8_0(.din(n11727), .dout(n11724));
    jdff dff_A_gSJ0gdUE4_0(.din(n11730), .dout(n11727));
    jdff dff_A_YvUVRR3i0_0(.din(n11733), .dout(n11730));
    jdff dff_A_W1rNttzp8_0(.din(n11736), .dout(n11733));
    jdff dff_A_U71Wqot97_0(.din(n11739), .dout(n11736));
    jdff dff_A_THkQBd0N4_0(.din(n11742), .dout(n11739));
    jdff dff_A_sQllPZOP3_0(.din(n11745), .dout(n11742));
    jdff dff_A_M3Jx9hsM7_0(.din(n11748), .dout(n11745));
    jdff dff_A_m3CNYkjw4_0(.din(n11751), .dout(n11748));
    jdff dff_A_tb1vKi2D2_0(.din(n2178), .dout(n11751));
    jdff dff_A_ZBIkZu7l7_2(.din(n11757), .dout(n11754));
    jdff dff_A_6Wjp8grj5_2(.din(n11760), .dout(n11757));
    jdff dff_A_T3SAIYIW2_2(.din(n11763), .dout(n11760));
    jdff dff_A_kw7EHbiv4_2(.din(n11766), .dout(n11763));
    jdff dff_A_NtF6MYvO1_2(.din(n11769), .dout(n11766));
    jdff dff_A_6tCwbCYX8_2(.din(n11772), .dout(n11769));
    jdff dff_A_apcfSdi74_2(.din(n11775), .dout(n11772));
    jdff dff_A_ATFi6iuZ7_2(.din(n11778), .dout(n11775));
    jdff dff_A_xAlNmWun0_2(.din(n11781), .dout(n11778));
    jdff dff_A_j40pknwC0_2(.din(n11784), .dout(n11781));
    jdff dff_A_Ll5Z3cAM9_2(.din(n2178), .dout(n11784));
    jdff dff_A_xYaKMUou5_0(.din(n11790), .dout(n11787));
    jdff dff_A_aVDGvTBl0_0(.din(n11793), .dout(n11790));
    jdff dff_A_RxSHQLeR8_0(.din(n11796), .dout(n11793));
    jdff dff_A_Nnpg2m7N6_0(.din(n11799), .dout(n11796));
    jdff dff_A_Ir6YNkOk1_0(.din(n11802), .dout(n11799));
    jdff dff_A_bz7cpQx72_0(.din(n11805), .dout(n11802));
    jdff dff_A_4tC039Cp9_0(.din(n11808), .dout(n11805));
    jdff dff_A_3vRFSR4i9_0(.din(n11811), .dout(n11808));
    jdff dff_A_5vdkZwtE7_0(.din(n11814), .dout(n11811));
    jdff dff_A_a4OH2zoE8_0(.din(n11817), .dout(n11814));
    jdff dff_A_w2IaFdIS4_0(.din(n11820), .dout(n11817));
    jdff dff_A_XhCivb6b2_0(.din(n11823), .dout(n11820));
    jdff dff_A_TjHKLjft5_0(.din(n11826), .dout(n11823));
    jdff dff_A_CPCe5i563_0(.din(n11829), .dout(n11826));
    jdff dff_A_0owSNGe31_0(.din(n11832), .dout(n11829));
    jdff dff_A_mCWSBeBZ3_0(.din(n11835), .dout(n11832));
    jdff dff_A_Gop5yYRW1_0(.din(n11838), .dout(n11835));
    jdff dff_A_ANmvAQjt5_0(.din(n11841), .dout(n11838));
    jdff dff_A_EpucYBj75_0(.din(n11844), .dout(n11841));
    jdff dff_A_UAnolVtf5_0(.din(G4088), .dout(n11844));
    jdff dff_A_UL2OIh3Q1_2(.din(n11850), .dout(n11847));
    jdff dff_A_bHQMXbCU3_2(.din(n11853), .dout(n11850));
    jdff dff_A_wkO4e9Mb7_2(.din(n11856), .dout(n11853));
    jdff dff_A_X2obzv4Q0_2(.din(n11859), .dout(n11856));
    jdff dff_A_5nRUB4HX9_2(.din(n11862), .dout(n11859));
    jdff dff_A_OYYFGldD6_2(.din(n11865), .dout(n11862));
    jdff dff_A_5CJESW8C2_2(.din(n11868), .dout(n11865));
    jdff dff_A_Z56cqX7z9_2(.din(n11871), .dout(n11868));
    jdff dff_A_4nEIVHXF1_2(.din(n11874), .dout(n11871));
    jdff dff_A_6X6eDHsP7_2(.din(n11877), .dout(n11874));
    jdff dff_A_NJJxwybQ5_2(.din(n11880), .dout(n11877));
    jdff dff_A_HPTCquTi3_2(.din(n11883), .dout(n11880));
    jdff dff_A_xCSFowHo3_2(.din(n11886), .dout(n11883));
    jdff dff_A_ycHHp8f25_2(.din(G4088), .dout(n11886));
    jdff dff_B_ib0tolKH8_0(.din(n4060), .dout(n11890));
    jdff dff_B_ZHJTGL6T5_0(.din(n11890), .dout(n11893));
    jdff dff_B_rrzrgDyO1_0(.din(n11893), .dout(n11896));
    jdff dff_B_rZKLo1xI4_0(.din(n11896), .dout(n11899));
    jdff dff_B_HgiEKKdQ0_0(.din(n11899), .dout(n11902));
    jdff dff_B_ze0IZd1g9_0(.din(n11902), .dout(n11905));
    jdff dff_B_nr8ZFi4z4_0(.din(n11905), .dout(n11908));
    jdff dff_B_f3FXnLPP7_0(.din(n11908), .dout(n11911));
    jdff dff_B_UEjY8Sqi8_0(.din(n11911), .dout(n11914));
    jdff dff_B_CZsidcyL3_0(.din(n11914), .dout(n11917));
    jdff dff_B_KwH0vJ9X5_0(.din(n11917), .dout(n11920));
    jdff dff_B_jK4BFWzy9_0(.din(n11920), .dout(n11923));
    jdff dff_B_xRRWSQSy0_0(.din(n11923), .dout(n11926));
    jdff dff_B_zDEEEJlf7_0(.din(n11926), .dout(n11929));
    jdff dff_B_xj7QYRbn9_0(.din(n11929), .dout(n11932));
    jdff dff_B_sE56QogI2_0(.din(n11932), .dout(n11935));
    jdff dff_B_iMDAzPsU1_0(.din(n11935), .dout(n11938));
    jdff dff_B_2tifSvW78_0(.din(n11938), .dout(n11941));
    jdff dff_B_ydx6ld577_0(.din(n11941), .dout(n11944));
    jdff dff_B_EGaddTYu8_0(.din(n11944), .dout(n11947));
    jdff dff_B_L6RmGUHe6_1(.din(n4029), .dout(n11950));
    jdff dff_B_humdkuXK2_1(.din(n11950), .dout(n11953));
    jdff dff_A_BU7ua3pb8_1(.din(n11958), .dout(n11955));
    jdff dff_A_NzWahemj5_1(.din(n11961), .dout(n11958));
    jdff dff_A_5hpZymzW3_1(.din(n11964), .dout(n11961));
    jdff dff_A_50tdOzGC6_1(.din(n11967), .dout(n11964));
    jdff dff_A_NCM9XFF52_1(.din(n11970), .dout(n11967));
    jdff dff_A_jOjA4B3G5_1(.din(n11973), .dout(n11970));
    jdff dff_A_t6JmLTNz6_1(.din(n11976), .dout(n11973));
    jdff dff_A_CL7LuoBa3_1(.din(n11979), .dout(n11976));
    jdff dff_A_E07EwdgE8_1(.din(n11982), .dout(n11979));
    jdff dff_A_l26b1K5J8_1(.din(n11985), .dout(n11982));
    jdff dff_A_X8EoCYOa1_1(.din(n11988), .dout(n11985));
    jdff dff_A_Bfwzorlg8_1(.din(n11991), .dout(n11988));
    jdff dff_A_7dZYS9B62_1(.din(n11994), .dout(n11991));
    jdff dff_A_eJL18UmO4_1(.din(n11997), .dout(n11994));
    jdff dff_A_i4rtBFi63_1(.din(n12000), .dout(n11997));
    jdff dff_A_x9mLeMmb5_1(.din(n12003), .dout(n12000));
    jdff dff_A_AprcE3Le9_1(.din(n12006), .dout(n12003));
    jdff dff_A_vENDE7u71_1(.din(n12009), .dout(n12006));
    jdff dff_A_a30Dc9h31_1(.din(n2178), .dout(n12009));
    jdff dff_A_nERkjmNx0_1(.din(n12015), .dout(n12012));
    jdff dff_A_2B9x6Pbt1_1(.din(n12018), .dout(n12015));
    jdff dff_A_E1ohL8k44_1(.din(n12021), .dout(n12018));
    jdff dff_A_CDMp4Ikt7_1(.din(n12024), .dout(n12021));
    jdff dff_A_QRTRrZUQ5_1(.din(n12027), .dout(n12024));
    jdff dff_A_1TQ1Sbgq5_1(.din(n12030), .dout(n12027));
    jdff dff_A_0yJBJbhp4_1(.din(n12033), .dout(n12030));
    jdff dff_A_RpM7D0SV8_1(.din(n12036), .dout(n12033));
    jdff dff_A_fpNWQqcX6_1(.din(n12039), .dout(n12036));
    jdff dff_A_DnYYmT1e8_1(.din(n12042), .dout(n12039));
    jdff dff_A_9fTUwbFM1_1(.din(n12045), .dout(n12042));
    jdff dff_A_NkOUE4QV9_1(.din(n12048), .dout(n12045));
    jdff dff_A_KCDM5riV0_1(.din(n12051), .dout(n12048));
    jdff dff_A_iveCsrqg5_1(.din(n12054), .dout(n12051));
    jdff dff_A_enNOYNb38_1(.din(n12057), .dout(n12054));
    jdff dff_A_MW1Bc9OL0_1(.din(n12060), .dout(n12057));
    jdff dff_A_0cPIuAtG6_1(.din(n12063), .dout(n12060));
    jdff dff_A_qmWfOSdh2_1(.din(n12066), .dout(n12063));
    jdff dff_A_cevV5e9A0_1(.din(G4088), .dout(n12066));
    jdff dff_B_Kgrl6t8O0_0(.din(n4096), .dout(n12070));
    jdff dff_B_DLZeU8Xl6_0(.din(n12070), .dout(n12073));
    jdff dff_B_sMp9HhWS2_0(.din(n12073), .dout(n12076));
    jdff dff_B_g9U9IYyX3_0(.din(n12076), .dout(n12079));
    jdff dff_B_YwCy8oZN3_0(.din(n12079), .dout(n12082));
    jdff dff_B_wMXNHpyY5_0(.din(n12082), .dout(n12085));
    jdff dff_B_Sx8LJqTa0_0(.din(n12085), .dout(n12088));
    jdff dff_B_Ffcd17VR9_0(.din(n12088), .dout(n12091));
    jdff dff_B_IH7fL4Nm9_0(.din(n12091), .dout(n12094));
    jdff dff_B_IpeAaenE6_0(.din(n12094), .dout(n12097));
    jdff dff_B_7BFlbH6r1_0(.din(n12097), .dout(n12100));
    jdff dff_B_kBY2X3PQ8_0(.din(n12100), .dout(n12103));
    jdff dff_B_dZxcuT3S9_0(.din(n12103), .dout(n12106));
    jdff dff_B_pjaLm7MK4_0(.din(n12106), .dout(n12109));
    jdff dff_B_42xHG2kJ5_0(.din(n12109), .dout(n12112));
    jdff dff_B_UydGTAgU1_0(.din(n12112), .dout(n12115));
    jdff dff_B_c9vALxBW9_0(.din(n12115), .dout(n12118));
    jdff dff_B_JhodgRi09_0(.din(n12118), .dout(n12121));
    jdff dff_B_MLLz04vA7_0(.din(n12121), .dout(n12124));
    jdff dff_B_TSdQhI3G0_0(.din(n12124), .dout(n12127));
    jdff dff_B_IzLWxCMd6_1(.din(n4068), .dout(n12130));
    jdff dff_A_4tE30Vwy7_2(.din(n15525), .dout(n12132));
    jdff dff_B_vSewMB1y0_0(.din(n4138), .dout(n12136));
    jdff dff_B_K9I4zaTN6_0(.din(n12136), .dout(n12139));
    jdff dff_B_o2NWN9GO7_0(.din(n12139), .dout(n12142));
    jdff dff_B_vmfxdA4W9_0(.din(n12142), .dout(n12145));
    jdff dff_B_cbtK9TAa6_0(.din(n12145), .dout(n12148));
    jdff dff_B_7hdcCF510_0(.din(n12148), .dout(n12151));
    jdff dff_B_MnZpJsH21_0(.din(n12151), .dout(n12154));
    jdff dff_B_GLoHxRd08_0(.din(n12154), .dout(n12157));
    jdff dff_B_o5P7f0169_0(.din(n12157), .dout(n12160));
    jdff dff_B_A2ZDyqOk5_0(.din(n12160), .dout(n12163));
    jdff dff_B_hmoUdjim9_0(.din(n12163), .dout(n12166));
    jdff dff_B_H7AUu1EA1_0(.din(n12166), .dout(n12169));
    jdff dff_B_O1AictfI4_0(.din(n12169), .dout(n12172));
    jdff dff_B_HoPAZZOw6_0(.din(n12172), .dout(n12175));
    jdff dff_B_EcNXww7o1_0(.din(n12175), .dout(n12178));
    jdff dff_B_q3PBkS4d2_0(.din(n12178), .dout(n12181));
    jdff dff_B_Fbl7Xien0_0(.din(n12181), .dout(n12184));
    jdff dff_B_qn5bWogX8_0(.din(n12184), .dout(n12187));
    jdff dff_B_aZcDLtDG6_0(.din(n12187), .dout(n12190));
    jdff dff_B_Jq7OWrXU8_1(.din(n4107), .dout(n12193));
    jdff dff_B_ovKHhbdz1_1(.din(n12193), .dout(n12196));
    jdff dff_B_Q8ABeuZd7_1(.din(n12196), .dout(n12199));
    jdff dff_A_ki0ASF4M8_0(.din(n12204), .dout(n12201));
    jdff dff_A_lFomooOb5_0(.din(n12207), .dout(n12204));
    jdff dff_A_ZrhT11cM2_0(.din(n12210), .dout(n12207));
    jdff dff_A_3gcMCGJO1_0(.din(n12213), .dout(n12210));
    jdff dff_A_WwunhunA1_0(.din(n12216), .dout(n12213));
    jdff dff_A_NbYHYZhP2_0(.din(n12219), .dout(n12216));
    jdff dff_A_Ubr6QMM37_0(.din(n12222), .dout(n12219));
    jdff dff_A_KlvC5Bed3_0(.din(n12225), .dout(n12222));
    jdff dff_A_bpKVYhvG2_0(.din(n12228), .dout(n12225));
    jdff dff_A_14KvqGfs6_0(.din(n12231), .dout(n12228));
    jdff dff_A_dugp3Xvq2_0(.din(n12234), .dout(n12231));
    jdff dff_A_EfMp3gX20_0(.din(n12237), .dout(n12234));
    jdff dff_A_GSPtApM15_0(.din(n12240), .dout(n12237));
    jdff dff_A_sxe1NpZs7_0(.din(n12243), .dout(n12240));
    jdff dff_A_pw6QaPsH7_0(.din(n12246), .dout(n12243));
    jdff dff_A_QLx6BECE6_0(.din(n12249), .dout(n12246));
    jdff dff_A_jMObl2In7_0(.din(n12252), .dout(n12249));
    jdff dff_A_58dpKpKG9_0(.din(n2178), .dout(n12252));
    jdff dff_A_7j2i70Da2_2(.din(n12258), .dout(n12255));
    jdff dff_A_5saTnAlU9_2(.din(n12261), .dout(n12258));
    jdff dff_A_wOJZlyW08_2(.din(n12264), .dout(n12261));
    jdff dff_A_rW2uadle0_2(.din(n12267), .dout(n12264));
    jdff dff_A_QeePR53M7_2(.din(n12270), .dout(n12267));
    jdff dff_A_tXPiKJdB2_2(.din(n12273), .dout(n12270));
    jdff dff_A_HUASIeDg1_2(.din(n12276), .dout(n12273));
    jdff dff_A_3iIQOlkU6_2(.din(n12279), .dout(n12276));
    jdff dff_A_FKKUxtHb1_2(.din(n12282), .dout(n12279));
    jdff dff_A_BeAran7r8_2(.din(n12285), .dout(n12282));
    jdff dff_A_mnwn4CYJ5_2(.din(n12288), .dout(n12285));
    jdff dff_A_wmHjxtnJ2_2(.din(n12291), .dout(n12288));
    jdff dff_A_tTGgUwVC5_2(.din(n12294), .dout(n12291));
    jdff dff_A_0k1q2xTD9_2(.din(n12297), .dout(n12294));
    jdff dff_A_778z624G2_2(.din(n12300), .dout(n12297));
    jdff dff_A_HUKVj8fA4_2(.din(n12303), .dout(n12300));
    jdff dff_A_K6Iq2SXH5_2(.din(n12306), .dout(n12303));
    jdff dff_A_rh61vUaI2_2(.din(n12309), .dout(n12306));
    jdff dff_A_vwgUazEv3_2(.din(n2178), .dout(n12309));
    jdff dff_A_q0V7oPRS2_0(.din(n12315), .dout(n12312));
    jdff dff_A_JTX3UDzV4_0(.din(n12318), .dout(n12315));
    jdff dff_A_Iyijq3FQ7_0(.din(n12321), .dout(n12318));
    jdff dff_A_1kc3LsSs4_0(.din(n12324), .dout(n12321));
    jdff dff_A_itu51oVY4_0(.din(n12327), .dout(n12324));
    jdff dff_A_s6sk633O5_0(.din(n12330), .dout(n12327));
    jdff dff_A_VOyMETQt6_0(.din(n12333), .dout(n12330));
    jdff dff_A_R8iQ81MI1_0(.din(n12336), .dout(n12333));
    jdff dff_A_nqY2Uh666_0(.din(n12339), .dout(n12336));
    jdff dff_A_Z4VBhC2g9_0(.din(n12342), .dout(n12339));
    jdff dff_A_EGko19t43_0(.din(n12345), .dout(n12342));
    jdff dff_A_iT981qWw0_0(.din(n12348), .dout(n12345));
    jdff dff_A_xPFvLJPM0_0(.din(n12351), .dout(n12348));
    jdff dff_A_RBKwFwSC2_0(.din(n12354), .dout(n12351));
    jdff dff_A_PifznpmR9_0(.din(n12357), .dout(n12354));
    jdff dff_A_THl7v3H99_0(.din(n12360), .dout(n12357));
    jdff dff_A_jVEqA2kz8_0(.din(G4088), .dout(n12360));
    jdff dff_A_Jz1nKuwT1_2(.din(n12366), .dout(n12363));
    jdff dff_A_ZKftlHUA6_2(.din(n12369), .dout(n12366));
    jdff dff_A_QpGET3A94_2(.din(n12372), .dout(n12369));
    jdff dff_A_dpVnm63O7_2(.din(n12375), .dout(n12372));
    jdff dff_A_iBsoTUgp3_2(.din(n12378), .dout(n12375));
    jdff dff_A_pwfpBjgA7_2(.din(n12381), .dout(n12378));
    jdff dff_A_2heLTJ250_2(.din(n12384), .dout(n12381));
    jdff dff_A_DwYJ2Z3T6_2(.din(n12387), .dout(n12384));
    jdff dff_A_kL3I5mTA9_2(.din(n12390), .dout(n12387));
    jdff dff_A_On1pbqBq8_2(.din(n12393), .dout(n12390));
    jdff dff_A_4MEsVlrA7_2(.din(n12396), .dout(n12393));
    jdff dff_A_034kpSf43_2(.din(n12399), .dout(n12396));
    jdff dff_A_PVtJZn7T6_2(.din(n12402), .dout(n12399));
    jdff dff_A_44gbeMXv9_2(.din(n12405), .dout(n12402));
    jdff dff_A_u8NlSWp98_2(.din(n12408), .dout(n12405));
    jdff dff_A_pUhPiI5Q7_2(.din(n12411), .dout(n12408));
    jdff dff_A_iDITvLu20_2(.din(n12414), .dout(n12411));
    jdff dff_A_DWaEN6e94_2(.din(n12417), .dout(n12414));
    jdff dff_A_YEAViCjk5_2(.din(n12420), .dout(n12417));
    jdff dff_A_SBWxVdOH5_2(.din(G4088), .dout(n12420));
    jdff dff_B_n0JULlMa2_0(.din(n4174), .dout(n12424));
    jdff dff_B_6uClxzp97_0(.din(n12424), .dout(n12427));
    jdff dff_B_mASb81U03_0(.din(n12427), .dout(n12430));
    jdff dff_B_7u1vgKYg6_0(.din(n12430), .dout(n12433));
    jdff dff_B_6ZiCbqQd3_0(.din(n12433), .dout(n12436));
    jdff dff_B_DoasNh6g3_0(.din(n12436), .dout(n12439));
    jdff dff_B_ESwQ3rgW2_0(.din(n12439), .dout(n12442));
    jdff dff_B_LQ1ySkNK0_0(.din(n12442), .dout(n12445));
    jdff dff_B_4WIrFQMY0_0(.din(n12445), .dout(n12448));
    jdff dff_B_m5LPkm6d0_0(.din(n12448), .dout(n12451));
    jdff dff_B_nv4Y54bF1_0(.din(n12451), .dout(n12454));
    jdff dff_B_66LUithL5_0(.din(n12454), .dout(n12457));
    jdff dff_B_1Rt8GaNl3_0(.din(n12457), .dout(n12460));
    jdff dff_B_zPBW5Ady7_0(.din(n12460), .dout(n12463));
    jdff dff_B_NYOotvNJ2_0(.din(n12463), .dout(n12466));
    jdff dff_B_6hQY9w0h2_0(.din(n12466), .dout(n12469));
    jdff dff_B_ttaq4fJM2_0(.din(n12469), .dout(n12472));
    jdff dff_B_uSs6b6rw5_0(.din(n12472), .dout(n12475));
    jdff dff_B_htTGsVSt9_0(.din(n12475), .dout(n12478));
    jdff dff_B_pwxvlKCd3_0(.din(n12478), .dout(n12481));
    jdff dff_B_QHr4jZ8J4_2(.din(G49), .dout(n12484));
    jdff dff_B_7nPZ3Rre2_1(.din(n4146), .dout(n12487));
    jdff dff_B_1fOuwH6L7_1(.din(n12487), .dout(n12490));
    jdff dff_A_XYqQI4tr2_1(.din(n12495), .dout(n12492));
    jdff dff_A_oq3zXX0C7_1(.din(n12498), .dout(n12495));
    jdff dff_A_6zqY6HDs9_1(.din(n12501), .dout(n12498));
    jdff dff_A_oOvmg0VM2_1(.din(n12504), .dout(n12501));
    jdff dff_A_cWTMDDHd3_1(.din(n12507), .dout(n12504));
    jdff dff_A_KmnruPb86_1(.din(n12510), .dout(n12507));
    jdff dff_A_UVi6WQcO4_1(.din(n12513), .dout(n12510));
    jdff dff_A_L0DHTAX51_1(.din(n12516), .dout(n12513));
    jdff dff_A_8fx1SEuP8_1(.din(n12519), .dout(n12516));
    jdff dff_A_uVTEgqv23_1(.din(n12522), .dout(n12519));
    jdff dff_A_pem9On199_1(.din(n12525), .dout(n12522));
    jdff dff_A_6PSyUXSh4_1(.din(n12528), .dout(n12525));
    jdff dff_A_w6WjhYjx1_1(.din(n12531), .dout(n12528));
    jdff dff_A_buocVb7d9_1(.din(n12534), .dout(n12531));
    jdff dff_A_Ewn4RtIF1_1(.din(n12537), .dout(n12534));
    jdff dff_A_5EtBrdRd7_1(.din(n12540), .dout(n12537));
    jdff dff_A_0lFLGziL8_1(.din(n12543), .dout(n12540));
    jdff dff_A_ZCrqRcRk6_1(.din(n12546), .dout(n12543));
    jdff dff_A_WPWSIian4_1(.din(n2387), .dout(n12546));
    jdff dff_A_d1MpCJDD3_2(.din(n12552), .dout(n12549));
    jdff dff_A_3pxIiuSN9_2(.din(n12555), .dout(n12552));
    jdff dff_A_YSWYsvqi3_2(.din(n12558), .dout(n12555));
    jdff dff_A_fyPmQcVm8_2(.din(n12561), .dout(n12558));
    jdff dff_A_trAjfuju2_2(.din(n12564), .dout(n12561));
    jdff dff_A_FvB1Qr9T2_2(.din(n12567), .dout(n12564));
    jdff dff_A_d94azWjj7_2(.din(n12570), .dout(n12567));
    jdff dff_A_dghaaWEf4_2(.din(n12573), .dout(n12570));
    jdff dff_A_sKsSBgEk9_2(.din(n12576), .dout(n12573));
    jdff dff_A_Zg41apJI9_2(.din(n12579), .dout(n12576));
    jdff dff_A_nL5LldgU1_2(.din(n12582), .dout(n12579));
    jdff dff_A_pYk34Idd7_2(.din(n12585), .dout(n12582));
    jdff dff_A_p2CFUgv18_2(.din(n12588), .dout(n12585));
    jdff dff_A_2VVTXPgh1_2(.din(n12591), .dout(n12588));
    jdff dff_A_IXYfh8WW7_2(.din(n12594), .dout(n12591));
    jdff dff_A_hQSBjLl80_2(.din(n12597), .dout(n12594));
    jdff dff_A_7U4jiEVr8_2(.din(n12600), .dout(n12597));
    jdff dff_A_GGkEp1kd8_2(.din(n12603), .dout(n12600));
    jdff dff_A_i8NayOmt2_2(.din(n12606), .dout(n12603));
    jdff dff_A_NG1cNPox5_2(.din(n2387), .dout(n12606));
    jdff dff_A_2T0YjRoR8_1(.din(n12612), .dout(n12609));
    jdff dff_A_ukj2lMYs3_1(.din(n12615), .dout(n12612));
    jdff dff_A_v3sMnOfD6_1(.din(n12618), .dout(n12615));
    jdff dff_A_GqDT4R8b0_1(.din(n12621), .dout(n12618));
    jdff dff_A_yTlniVR09_1(.din(n12624), .dout(n12621));
    jdff dff_A_xVptjahG8_1(.din(n12627), .dout(n12624));
    jdff dff_A_fXwbrHrn6_1(.din(n12630), .dout(n12627));
    jdff dff_A_p6MkiGPY8_1(.din(n12633), .dout(n12630));
    jdff dff_A_gTLj0d0T3_1(.din(n12636), .dout(n12633));
    jdff dff_A_ydVYs9g36_1(.din(n12639), .dout(n12636));
    jdff dff_A_3TXZKoFM6_1(.din(n12642), .dout(n12639));
    jdff dff_A_t7MkKv054_1(.din(n12645), .dout(n12642));
    jdff dff_A_cuEbSjxY8_1(.din(n12648), .dout(n12645));
    jdff dff_A_oVjjiMYT7_1(.din(n12651), .dout(n12648));
    jdff dff_A_TkRUub3H9_1(.din(n12654), .dout(n12651));
    jdff dff_A_nx9bvsxe4_1(.din(n12657), .dout(n12654));
    jdff dff_A_9HOC5UXP4_1(.din(n12660), .dout(n12657));
    jdff dff_A_WmhOFS8T7_1(.din(n12663), .dout(n12660));
    jdff dff_A_TBX5Mh469_1(.din(G4089), .dout(n12663));
    jdff dff_A_8JXtxRY97_2(.din(n12669), .dout(n12666));
    jdff dff_A_fEPr5yPk6_2(.din(n12672), .dout(n12669));
    jdff dff_A_2EIqdY9a5_2(.din(n12675), .dout(n12672));
    jdff dff_A_G1ybo0jX4_2(.din(n12678), .dout(n12675));
    jdff dff_A_OLvqYejf3_2(.din(n12681), .dout(n12678));
    jdff dff_A_SlkMDmm30_2(.din(n12684), .dout(n12681));
    jdff dff_A_RBqN83Ax1_2(.din(n12687), .dout(n12684));
    jdff dff_A_rIpBa0Ap7_2(.din(n12690), .dout(n12687));
    jdff dff_A_cNl0c7bd9_2(.din(n12693), .dout(n12690));
    jdff dff_A_OXGOCku81_2(.din(n12696), .dout(n12693));
    jdff dff_A_he3bOx2Q8_2(.din(n12699), .dout(n12696));
    jdff dff_A_vSTRQghL4_2(.din(n12702), .dout(n12699));
    jdff dff_A_Kv3cKQwf0_2(.din(n12705), .dout(n12702));
    jdff dff_A_qKsaUKEO2_2(.din(n12708), .dout(n12705));
    jdff dff_A_eDAwHI2u4_2(.din(n12711), .dout(n12708));
    jdff dff_A_P8UycJDD8_2(.din(n12714), .dout(n12711));
    jdff dff_A_QxwvuVAj4_2(.din(n12717), .dout(n12714));
    jdff dff_A_rNFC4wfo5_2(.din(n12720), .dout(n12717));
    jdff dff_A_kcw9hboA7_2(.din(n12723), .dout(n12720));
    jdff dff_A_RJWpgXXD6_2(.din(G4089), .dout(n12723));
    jdff dff_B_Tx3nH3oS8_0(.din(n4210), .dout(n12727));
    jdff dff_B_hgGxcLaZ2_0(.din(n12727), .dout(n12730));
    jdff dff_B_mbycB4hs9_0(.din(n12730), .dout(n12733));
    jdff dff_B_idaAs0Bw9_0(.din(n12733), .dout(n12736));
    jdff dff_B_XzBlgQAC4_0(.din(n12736), .dout(n12739));
    jdff dff_B_Q6RuIBFz3_0(.din(n12739), .dout(n12742));
    jdff dff_B_Q7Atw7ZZ3_0(.din(n12742), .dout(n12745));
    jdff dff_B_da2HRq8B2_0(.din(n12745), .dout(n12748));
    jdff dff_B_Y1Z1LecR4_0(.din(n12748), .dout(n12751));
    jdff dff_B_ijvYExa02_0(.din(n12751), .dout(n12754));
    jdff dff_B_dsWROEKM4_0(.din(n12754), .dout(n12757));
    jdff dff_B_AYDWcRqT7_0(.din(n12757), .dout(n12760));
    jdff dff_B_fegGlux16_0(.din(n12760), .dout(n12763));
    jdff dff_B_bLveDmSc6_0(.din(n12763), .dout(n12766));
    jdff dff_B_F7XzmOPd8_0(.din(n12766), .dout(n12769));
    jdff dff_B_F3T0l02s7_0(.din(n12769), .dout(n12772));
    jdff dff_B_Xtb5aoXD7_0(.din(n12772), .dout(n12775));
    jdff dff_B_4VDLMkRI1_0(.din(n12775), .dout(n12778));
    jdff dff_B_ESMV3WSY4_0(.din(n12778), .dout(n12781));
    jdff dff_B_GRzCDFLx2_0(.din(n12781), .dout(n12784));
    jdff dff_A_RHULBzFo7_2(.din(n16122), .dout(n12786));
    jdff dff_B_uaO0d8MK4_2(.din(G103), .dout(n12790));
    jdff dff_B_T1W1r0Mi2_1(.din(n4182), .dout(n12793));
    jdff dff_B_hdS1Xd212_0(.din(n4246), .dout(n12796));
    jdff dff_B_qh3ZIsU17_0(.din(n12796), .dout(n12799));
    jdff dff_B_pnffsTc89_0(.din(n12799), .dout(n12802));
    jdff dff_B_Y2FFdj650_0(.din(n12802), .dout(n12805));
    jdff dff_B_PCe4hWqu0_0(.din(n12805), .dout(n12808));
    jdff dff_B_iIdX5ytB4_0(.din(n12808), .dout(n12811));
    jdff dff_B_8ru6XpIH6_0(.din(n12811), .dout(n12814));
    jdff dff_B_o7zdvJmS4_0(.din(n12814), .dout(n12817));
    jdff dff_B_jSKjCHVl7_0(.din(n12817), .dout(n12820));
    jdff dff_B_IPorO2iJ9_0(.din(n12820), .dout(n12823));
    jdff dff_B_wiAzWvOK8_0(.din(n12823), .dout(n12826));
    jdff dff_B_59pWEpqM0_0(.din(n12826), .dout(n12829));
    jdff dff_B_0NrHRDnN8_0(.din(n12829), .dout(n12832));
    jdff dff_B_z5Yeu1YP3_0(.din(n12832), .dout(n12835));
    jdff dff_B_2RxG98qb5_0(.din(n12835), .dout(n12838));
    jdff dff_B_evBNwruV0_0(.din(n12838), .dout(n12841));
    jdff dff_B_LO9JOhnI8_0(.din(n12841), .dout(n12844));
    jdff dff_B_LqHYB27G5_0(.din(n12844), .dout(n12847));
    jdff dff_B_tCYsu0WS0_0(.din(n12847), .dout(n12850));
    jdff dff_B_YnmLANBf9_2(.din(G40), .dout(n12853));
    jdff dff_B_WKybI4lD9_1(.din(n4218), .dout(n12856));
    jdff dff_B_Nt5hPK6m3_1(.din(n12856), .dout(n12859));
    jdff dff_B_C4l1m0gX6_1(.din(n12859), .dout(n12862));
    jdff dff_A_vnhR8o3d4_0(.din(n12867), .dout(n12864));
    jdff dff_A_GEU44v5Q4_0(.din(n12870), .dout(n12867));
    jdff dff_A_wfZ8ZsLa1_0(.din(n12873), .dout(n12870));
    jdff dff_A_F5aYLFnV1_0(.din(n12876), .dout(n12873));
    jdff dff_A_tmBuKDQV3_0(.din(n12879), .dout(n12876));
    jdff dff_A_vLkJbTwn0_0(.din(n12882), .dout(n12879));
    jdff dff_A_1WgpBUtp3_0(.din(n12885), .dout(n12882));
    jdff dff_A_ilK3GIH75_0(.din(n12888), .dout(n12885));
    jdff dff_A_Emgmwmvm8_0(.din(n12891), .dout(n12888));
    jdff dff_A_MfPtqWRG0_0(.din(n12894), .dout(n12891));
    jdff dff_A_R9fmyxep8_0(.din(n12897), .dout(n12894));
    jdff dff_A_7wRx7xaG3_0(.din(n12900), .dout(n12897));
    jdff dff_A_cHzaRFDO4_0(.din(n12903), .dout(n12900));
    jdff dff_A_G4Xxnea55_0(.din(n12906), .dout(n12903));
    jdff dff_A_MvsB6TA38_0(.din(n12909), .dout(n12906));
    jdff dff_A_iA2VBYc17_0(.din(n12912), .dout(n12909));
    jdff dff_A_GgQ1ID3J5_0(.din(n12915), .dout(n12912));
    jdff dff_A_bNh4M6Ep2_0(.din(n2387), .dout(n12915));
    jdff dff_A_TJygGqzl7_2(.din(n12921), .dout(n12918));
    jdff dff_A_iU15CS426_2(.din(n12924), .dout(n12921));
    jdff dff_A_dpzeTCi89_2(.din(n12927), .dout(n12924));
    jdff dff_A_yQgaYmtb1_2(.din(n12930), .dout(n12927));
    jdff dff_A_cfEQ7Qna0_2(.din(n12933), .dout(n12930));
    jdff dff_A_E56k601s3_2(.din(n12936), .dout(n12933));
    jdff dff_A_jio8YAFG7_2(.din(n12939), .dout(n12936));
    jdff dff_A_PZrhnLXL2_2(.din(n12942), .dout(n12939));
    jdff dff_A_jxw9vpws8_2(.din(n12945), .dout(n12942));
    jdff dff_A_cJft473K6_2(.din(n12948), .dout(n12945));
    jdff dff_A_7PRmW6Ip6_2(.din(n12951), .dout(n12948));
    jdff dff_A_v5VCptiH7_2(.din(n12954), .dout(n12951));
    jdff dff_A_O40I5Xo73_2(.din(n12957), .dout(n12954));
    jdff dff_A_lsbdGSYB5_2(.din(n12960), .dout(n12957));
    jdff dff_A_VAJHHmLj1_2(.din(n12963), .dout(n12960));
    jdff dff_A_KKh4rwpx4_2(.din(n12966), .dout(n12963));
    jdff dff_A_HFgvA4HM3_2(.din(n12969), .dout(n12966));
    jdff dff_A_IPJr4FrX8_2(.din(n12972), .dout(n12969));
    jdff dff_A_FHS91h1n8_2(.din(n2387), .dout(n12972));
    jdff dff_A_HSz7qNpi9_0(.din(n12978), .dout(n12975));
    jdff dff_A_viGMn3QI9_0(.din(n12981), .dout(n12978));
    jdff dff_A_5uhSE4tk9_0(.din(n12984), .dout(n12981));
    jdff dff_A_yD8WmPpv2_0(.din(n12987), .dout(n12984));
    jdff dff_A_pFbS3kbv3_0(.din(n12990), .dout(n12987));
    jdff dff_A_eSWenga86_0(.din(n12993), .dout(n12990));
    jdff dff_A_K2qJq7z68_0(.din(n12996), .dout(n12993));
    jdff dff_A_JJWtZTpV4_0(.din(n12999), .dout(n12996));
    jdff dff_A_yc4fj2JV3_0(.din(n13002), .dout(n12999));
    jdff dff_A_RRimMF1z8_0(.din(n13005), .dout(n13002));
    jdff dff_A_g6rtoMU50_0(.din(n13008), .dout(n13005));
    jdff dff_A_NM2AqfPu2_0(.din(n13011), .dout(n13008));
    jdff dff_A_IhdNb4sX1_0(.din(n13014), .dout(n13011));
    jdff dff_A_lpLbDs6F4_0(.din(n13017), .dout(n13014));
    jdff dff_A_2neD71Vj8_0(.din(n13020), .dout(n13017));
    jdff dff_A_y72R2Axt7_0(.din(n13023), .dout(n13020));
    jdff dff_A_Hzdn82JJ8_0(.din(G4089), .dout(n13023));
    jdff dff_A_a1Ck1LAN9_2(.din(n13029), .dout(n13026));
    jdff dff_A_O6xluIb36_2(.din(n13032), .dout(n13029));
    jdff dff_A_GiiiFa3n3_2(.din(n13035), .dout(n13032));
    jdff dff_A_rAuThIDR2_2(.din(n13038), .dout(n13035));
    jdff dff_A_DHgXbhto7_2(.din(n13041), .dout(n13038));
    jdff dff_A_7XYq4DsJ4_2(.din(n13044), .dout(n13041));
    jdff dff_A_K5jHEDma0_2(.din(n13047), .dout(n13044));
    jdff dff_A_496LZMLI8_2(.din(n13050), .dout(n13047));
    jdff dff_A_pYJCONra7_2(.din(n13053), .dout(n13050));
    jdff dff_A_FyPPEUMn5_2(.din(n13056), .dout(n13053));
    jdff dff_A_Qtz8xAoZ2_2(.din(n13059), .dout(n13056));
    jdff dff_A_d4lzdykj4_2(.din(n13062), .dout(n13059));
    jdff dff_A_KXSTPiPM8_2(.din(n13065), .dout(n13062));
    jdff dff_A_ncMREv2P8_2(.din(n13068), .dout(n13065));
    jdff dff_A_1dAyC3bT0_2(.din(n13071), .dout(n13068));
    jdff dff_A_woZw5Kyi8_2(.din(n13074), .dout(n13071));
    jdff dff_A_4uPCxWrf1_2(.din(n13077), .dout(n13074));
    jdff dff_A_uif6g65M9_2(.din(n13080), .dout(n13077));
    jdff dff_A_XOZcIZ1n5_2(.din(n13083), .dout(n13080));
    jdff dff_A_8Qwl9bBz2_2(.din(G4089), .dout(n13083));
    jdff dff_B_yYB6TAZo9_0(.din(n4278), .dout(n13087));
    jdff dff_B_N9rGxIIx6_0(.din(n13087), .dout(n13090));
    jdff dff_B_Arf4ptQS9_0(.din(n13090), .dout(n13093));
    jdff dff_B_LT7gTv8j4_0(.din(n13093), .dout(n13096));
    jdff dff_B_PPi1ZdXw9_0(.din(n13096), .dout(n13099));
    jdff dff_B_1zYuoSQ24_0(.din(n13099), .dout(n13102));
    jdff dff_B_9ZxP1CpH4_0(.din(n13102), .dout(n13105));
    jdff dff_B_dYNfhZ5W5_0(.din(n13105), .dout(n13108));
    jdff dff_B_8Ouoy7LE7_0(.din(n13108), .dout(n13111));
    jdff dff_B_15p2zQ3u1_0(.din(n13111), .dout(n13114));
    jdff dff_B_sPD79SSp3_0(.din(n13114), .dout(n13117));
    jdff dff_B_THVAymhP4_0(.din(n13117), .dout(n13120));
    jdff dff_B_h3nGbSLd0_0(.din(n13120), .dout(n13123));
    jdff dff_B_MLpbz2IM5_0(.din(n13123), .dout(n13126));
    jdff dff_B_e4BKR3X65_0(.din(n13126), .dout(n13129));
    jdff dff_B_YKawyxsP8_0(.din(n13129), .dout(n13132));
    jdff dff_B_ylHZqwYG2_0(.din(n13132), .dout(n13135));
    jdff dff_B_o3U269by6_0(.din(n13135), .dout(n13138));
    jdff dff_B_o2lYWXg34_0(.din(n4274), .dout(n13141));
    jdff dff_B_QTf9ErPX5_1(.din(n4254), .dout(n13144));
    jdff dff_B_oWAW81qD6_1(.din(n13144), .dout(n13147));
    jdff dff_B_oMESUjmC8_1(.din(n13147), .dout(n13150));
    jdff dff_A_3K5qGB1N1_0(.din(n13155), .dout(n13152));
    jdff dff_A_95xPttmD4_0(.din(n13158), .dout(n13155));
    jdff dff_A_Di47PCmo2_0(.din(n13161), .dout(n13158));
    jdff dff_A_GB3lom5E6_0(.din(n13164), .dout(n13161));
    jdff dff_A_PKL4Ihwc6_0(.din(n13167), .dout(n13164));
    jdff dff_A_VOAFHszn5_0(.din(n13455), .dout(n13167));
    jdff dff_A_APFbucbk9_1(.din(n13455), .dout(n13170));
    jdff dff_A_tXUoP4lF0_0(.din(n13176), .dout(n13173));
    jdff dff_A_Aw6lNMMU4_0(.din(n13179), .dout(n13176));
    jdff dff_A_z9ivnzQ28_0(.din(n13182), .dout(n13179));
    jdff dff_A_wAZAh3OW7_0(.din(n16839), .dout(n13182));
    jdff dff_A_VYfevSgU1_1(.din(n13188), .dout(n13185));
    jdff dff_A_IdOvsTrc2_1(.din(n16839), .dout(n13188));
    jdff dff_A_2k6ktBTe1_0(.din(n13194), .dout(n13191));
    jdff dff_A_zT7UaD024_0(.din(n13197), .dout(n13194));
    jdff dff_A_hra1La5V3_0(.din(n13200), .dout(n13197));
    jdff dff_A_uC2OrI8W5_0(.din(n13203), .dout(n13200));
    jdff dff_A_Ho32hBRl7_0(.din(n13206), .dout(n13203));
    jdff dff_A_wEzRSUOx8_0(.din(n20706), .dout(n13206));
    jdff dff_A_9uvh0oUf1_1(.din(n20706), .dout(n13209));
    jdff dff_B_Qjq07H452_0(.din(n4314), .dout(n13213));
    jdff dff_B_Ijvwahbm8_0(.din(n13213), .dout(n13216));
    jdff dff_B_U1WfJBmg3_0(.din(n13216), .dout(n13219));
    jdff dff_B_npXesAWe5_0(.din(n13219), .dout(n13222));
    jdff dff_B_Zv8jywsV7_0(.din(n13222), .dout(n13225));
    jdff dff_B_RVc9EPDD6_0(.din(n13225), .dout(n13228));
    jdff dff_B_F2soZxR53_0(.din(n13228), .dout(n13231));
    jdff dff_B_6hvB721S8_0(.din(n13231), .dout(n13234));
    jdff dff_B_lBoNCdOZ8_0(.din(n13234), .dout(n13237));
    jdff dff_B_9lUh3Cp42_0(.din(n13237), .dout(n13240));
    jdff dff_B_WSczm8ck7_0(.din(n13240), .dout(n13243));
    jdff dff_B_xbporivq5_0(.din(n13243), .dout(n13246));
    jdff dff_B_1DElu1if2_0(.din(n13246), .dout(n13249));
    jdff dff_B_yu3bNiHn0_0(.din(n13249), .dout(n13252));
    jdff dff_B_w0Eo8hmv1_0(.din(n13252), .dout(n13255));
    jdff dff_B_eZzwnoab4_0(.din(n13255), .dout(n13258));
    jdff dff_B_myS6yNBK6_0(.din(n13258), .dout(n13261));
    jdff dff_B_v9gZSm0M9_0(.din(n13261), .dout(n13264));
    jdff dff_B_k8e4oTpX8_0(.din(n13264), .dout(n13267));
    jdff dff_B_YFV8slcf0_0(.din(n4310), .dout(n13270));
    jdff dff_B_WtmtCWCJ1_1(.din(n4290), .dout(n13273));
    jdff dff_B_lXMbRhuD4_1(.din(n4334), .dout(n13276));
    jdff dff_B_HY13YXOs5_1(.din(n13276), .dout(n13279));
    jdff dff_B_FonaWKoP9_1(.din(n13279), .dout(n13282));
    jdff dff_B_i6hooBBx6_1(.din(n13282), .dout(n13285));
    jdff dff_B_pPnBGupb1_1(.din(n13285), .dout(n13288));
    jdff dff_B_r4f2I6v88_1(.din(n13288), .dout(n13291));
    jdff dff_B_o77agAi46_1(.din(n13291), .dout(n13294));
    jdff dff_B_5ZIGr0MD4_1(.din(n13294), .dout(n13297));
    jdff dff_B_fug5m2Uz6_1(.din(n13297), .dout(n13300));
    jdff dff_B_PMrZCyXN4_1(.din(n13300), .dout(n13303));
    jdff dff_B_h1rIcDDy2_1(.din(n13303), .dout(n13306));
    jdff dff_B_cUS0QtHJ5_1(.din(n13306), .dout(n13309));
    jdff dff_B_vT0DQTLX3_1(.din(n13309), .dout(n13312));
    jdff dff_B_4RuFdNRT6_1(.din(n13312), .dout(n13315));
    jdff dff_B_OX8ualn71_1(.din(n13315), .dout(n13318));
    jdff dff_B_fKIVnX7K4_1(.din(n13318), .dout(n13321));
    jdff dff_B_m6W3wUY36_1(.din(n13321), .dout(n13324));
    jdff dff_B_7enCrB7h2_1(.din(n13324), .dout(n13327));
    jdff dff_B_m5sqUrVV8_1(.din(n13327), .dout(n13330));
    jdff dff_B_ObQwgJC15_1(.din(n4338), .dout(n13333));
    jdff dff_A_5xdz7XYU7_0(.din(n16530), .dout(n13335));
    jdff dff_A_Hpy5MfOc2_1(.din(n16530), .dout(n13338));
    jdff dff_B_Ym1YPgLI8_0(.din(n4330), .dout(n13342));
    jdff dff_B_AtolZT8F9_1(.din(n4370), .dout(n13345));
    jdff dff_B_pwRJUksx3_1(.din(n13345), .dout(n13348));
    jdff dff_B_8woNUihl2_1(.din(n13348), .dout(n13351));
    jdff dff_B_skGCBfp53_1(.din(n13351), .dout(n13354));
    jdff dff_B_ZRgVQ4vv1_1(.din(n13354), .dout(n13357));
    jdff dff_B_JL4i2ARc7_1(.din(n13357), .dout(n13360));
    jdff dff_B_zbAMYEjV6_1(.din(n13360), .dout(n13363));
    jdff dff_B_aHWdyLhU9_1(.din(n13363), .dout(n13366));
    jdff dff_B_LWqd3uZb3_1(.din(n13366), .dout(n13369));
    jdff dff_B_V6K2BZu84_1(.din(n13369), .dout(n13372));
    jdff dff_B_16LEHejr9_1(.din(n13372), .dout(n13375));
    jdff dff_B_0660sNOs6_1(.din(n13375), .dout(n13378));
    jdff dff_B_daWiL30p6_1(.din(n13378), .dout(n13381));
    jdff dff_B_LD59wa0H4_1(.din(n13381), .dout(n13384));
    jdff dff_B_RkSYgIEO4_1(.din(n13384), .dout(n13387));
    jdff dff_B_xxMAb5BD6_1(.din(n13387), .dout(n13390));
    jdff dff_B_LBvUITzk2_1(.din(n13390), .dout(n13393));
    jdff dff_B_gbqBUwIl1_1(.din(n13393), .dout(n13396));
    jdff dff_B_5ibtmSeG1_1(.din(n13396), .dout(n13399));
    jdff dff_B_AZuUwZqn7_1(.din(n13399), .dout(n13402));
    jdff dff_B_EWcgwott5_1(.din(n4374), .dout(n13405));
    jdff dff_A_HFPQpTJG5_0(.din(n16782), .dout(n13407));
    jdff dff_A_ppmNuYTf8_2(.din(n16782), .dout(n13410));
    jdff dff_A_eTspS4q13_0(.din(n13416), .dout(n13413));
    jdff dff_A_yDlvjHw96_0(.din(n13422), .dout(n13416));
    jdff dff_A_1hELk9MS9_1(.din(n13422), .dout(n13419));
    jdff dff_A_4nj4cidn5_0(.din(n13425), .dout(n13422));
    jdff dff_A_76uPv6W69_0(.din(n13428), .dout(n13425));
    jdff dff_A_OEPIWn4Y0_0(.din(n13431), .dout(n13428));
    jdff dff_A_rwowK5U84_0(.din(n13434), .dout(n13431));
    jdff dff_A_luLEJHA67_0(.din(n13437), .dout(n13434));
    jdff dff_A_NTrox4ME1_0(.din(n13440), .dout(n13437));
    jdff dff_A_oTeowHYw0_0(.din(n13443), .dout(n13440));
    jdff dff_A_XzEB0ILD7_0(.din(n13446), .dout(n13443));
    jdff dff_A_DL87QF4n7_0(.din(n13449), .dout(n13446));
    jdff dff_A_c9J82Jq75_0(.din(n13452), .dout(n13449));
    jdff dff_A_VMh60d2x4_0(.din(n13492), .dout(n13452));
    jdff dff_A_yBwxPKn73_1(.din(n13458), .dout(n13455));
    jdff dff_A_DRZzqlun9_1(.din(n13461), .dout(n13458));
    jdff dff_A_pFQl3gRB8_1(.din(n13464), .dout(n13461));
    jdff dff_A_eZp5P86f6_1(.din(n13492), .dout(n13464));
    jdff dff_B_FXNeghKD8_3(.din(n2944), .dout(n13468));
    jdff dff_B_KHVOwOSr1_3(.din(n13468), .dout(n13471));
    jdff dff_B_B8UBqGIR9_3(.din(n13471), .dout(n13474));
    jdff dff_B_6qKQzCyJ9_3(.din(n13474), .dout(n13477));
    jdff dff_B_3aabpeHx6_3(.din(n13477), .dout(n13480));
    jdff dff_B_68lGMx9Z2_3(.din(n13480), .dout(n13483));
    jdff dff_B_7zwlRWqY0_3(.din(n13483), .dout(n13486));
    jdff dff_B_VhKtsMnV0_3(.din(n13486), .dout(n13489));
    jdff dff_B_XHslf9w03_3(.din(n13489), .dout(n13492));
    jdff dff_B_KcfGaCcD5_0(.din(n4366), .dout(n13495));
    jdff dff_A_0vW8M7pl8_0(.din(n14553), .dout(n13497));
    jdff dff_B_CRtjkcmB5_0(.din(n4422), .dout(n13501));
    jdff dff_B_XD00l3zH0_0(.din(n13501), .dout(n13504));
    jdff dff_B_qQ5xfVII6_0(.din(n13504), .dout(n13507));
    jdff dff_B_MOeP6t8y4_0(.din(n13507), .dout(n13510));
    jdff dff_B_pN7XJb359_0(.din(n13510), .dout(n13513));
    jdff dff_B_EZtPf5V10_0(.din(n13513), .dout(n13516));
    jdff dff_B_6nFsEehQ2_0(.din(n13516), .dout(n13519));
    jdff dff_B_qsbTU6aX5_0(.din(n13519), .dout(n13522));
    jdff dff_B_ZRSVymbL6_0(.din(n13522), .dout(n13525));
    jdff dff_B_xFuDborj1_0(.din(n13525), .dout(n13528));
    jdff dff_B_ZP3Ou09r3_0(.din(n13528), .dout(n13531));
    jdff dff_B_t1GA4otx5_0(.din(n13531), .dout(n13534));
    jdff dff_B_TYfR1S6V5_0(.din(n13534), .dout(n13537));
    jdff dff_B_nOX7kZNc2_0(.din(n13537), .dout(n13540));
    jdff dff_B_Lwbztwl10_0(.din(n13540), .dout(n13543));
    jdff dff_B_F7ipmCq31_0(.din(n13543), .dout(n13546));
    jdff dff_B_bZvC7fT64_0(.din(n13546), .dout(n13549));
    jdff dff_B_XKntAtJb8_0(.din(n13549), .dout(n13552));
    jdff dff_B_ihjrzGeK4_0(.din(n4418), .dout(n13555));
    jdff dff_B_hv1i2ayl9_2(.din(G173), .dout(n13558));
    jdff dff_B_r4QAimLG6_2(.din(G203), .dout(n13561));
    jdff dff_B_PZmhi2Ux9_2(.din(n13561), .dout(n13564));
    jdff dff_B_tiUFcGwx2_1(.din(n4398), .dout(n13567));
    jdff dff_B_5TN3qEZ67_1(.din(n13567), .dout(n13570));
    jdff dff_B_6BA4nhSw3_1(.din(n13570), .dout(n13573));
    jdff dff_B_BtdO2gts0_1(.din(n3933), .dout(n13576));
    jdff dff_B_ePHP2b9y8_1(.din(n13576), .dout(n13579));
    jdff dff_B_fcLVQSPd9_1(.din(n13579), .dout(n13582));
    jdff dff_B_EB1jyn2G3_1(.din(n13582), .dout(n13585));
    jdff dff_B_SwwdMu4Y8_1(.din(n13585), .dout(n13588));
    jdff dff_B_Y0z90IVy1_1(.din(n13588), .dout(n13591));
    jdff dff_B_6X7uMZkU6_1(.din(n13591), .dout(n13594));
    jdff dff_B_Q2EHH6wW5_1(.din(n13594), .dout(n13597));
    jdff dff_B_GyAtbnbc1_1(.din(n13597), .dout(n13600));
    jdff dff_B_uBwPSrnu7_1(.din(n13600), .dout(n13603));
    jdff dff_B_nszbMZii6_1(.din(n13603), .dout(n13606));
    jdff dff_B_kOvO2zm75_1(.din(n13606), .dout(n13609));
    jdff dff_B_7ZKBsrZl6_1(.din(n13609), .dout(n13612));
    jdff dff_B_lMTC9uL96_0(.din(n3945), .dout(n13615));
    jdff dff_B_NaHG9NqN9_0(.din(n13615), .dout(n13618));
    jdff dff_B_ePknq90s6_0(.din(n13618), .dout(n13621));
    jdff dff_B_9zm5aosW8_0(.din(n13621), .dout(n13624));
    jdff dff_B_K9NaHNCa3_0(.din(n13624), .dout(n13627));
    jdff dff_B_xDbWoImo4_0(.din(n13627), .dout(n13630));
    jdff dff_B_q0elnQ2I0_0(.din(n13630), .dout(n13633));
    jdff dff_B_Li3oPenu2_0(.din(n13633), .dout(n13636));
    jdff dff_B_75NlZSdJ8_0(.din(n13636), .dout(n13639));
    jdff dff_B_ZXo0Ajip9_1(.din(n1044), .dout(n13642));
    jdff dff_B_GWbKGlHL4_1(.din(n1025), .dout(n13645));
    jdff dff_B_UdMAZiz87_1(.din(G113), .dout(n13648));
    jdff dff_B_aljd1Jnr4_1(.din(n13648), .dout(n13651));
    jdff dff_A_vrU2TEnj8_0(.din(n13656), .dout(n13653));
    jdff dff_A_c63SQAcV4_0(.din(n13659), .dout(n13656));
    jdff dff_A_IhPVHmS03_0(.din(n13662), .dout(n13659));
    jdff dff_A_ppsnujPY6_0(.din(n13665), .dout(n13662));
    jdff dff_A_L3tuD2tc0_0(.din(n13668), .dout(n13665));
    jdff dff_A_eY1SVWxl9_0(.din(n14871), .dout(n13668));
    jdff dff_A_A9qC9FTc9_1(.din(n14871), .dout(n13671));
    jdff dff_B_wd3WBX613_1(.din(n3788), .dout(n13675));
    jdff dff_B_6TtA3TpS8_1(.din(n13675), .dout(n13678));
    jdff dff_B_5xvRDIY67_1(.din(n13678), .dout(n13681));
    jdff dff_B_8dNRyRnD0_1(.din(n13681), .dout(n13684));
    jdff dff_B_bPLbmZ3P5_1(.din(n13684), .dout(n13687));
    jdff dff_B_5aPzewHF4_1(.din(n13687), .dout(n13690));
    jdff dff_B_mUOTr4No8_1(.din(n13690), .dout(n13693));
    jdff dff_B_tCN1YVT29_1(.din(n13693), .dout(n13696));
    jdff dff_B_EHvUj70j2_1(.din(n13696), .dout(n13699));
    jdff dff_B_yJWGdK1H6_1(.din(n13699), .dout(n13702));
    jdff dff_B_J8o4nnxb3_1(.din(n13702), .dout(n13705));
    jdff dff_B_nhj6bx8W5_0(.din(n3800), .dout(n13708));
    jdff dff_B_QAm637499_0(.din(n13708), .dout(n13711));
    jdff dff_B_iyvZikVc5_0(.din(n13711), .dout(n13714));
    jdff dff_B_qxjqu7PP5_0(.din(n13714), .dout(n13717));
    jdff dff_B_sltbgdBD4_0(.din(n13717), .dout(n13720));
    jdff dff_B_Ghv57Xo84_0(.din(n13720), .dout(n13723));
    jdff dff_B_fx5k9FZY9_0(.din(n13723), .dout(n13726));
    jdff dff_A_2Oqkcr7F2_1(.din(n13731), .dout(n13728));
    jdff dff_A_qO258kTB7_1(.din(n13734), .dout(n13731));
    jdff dff_A_WqYq0zA37_1(.din(n13737), .dout(n13734));
    jdff dff_A_GxTLhJZx7_1(.din(n13740), .dout(n13737));
    jdff dff_A_wfN3sNeB6_1(.din(n2906), .dout(n13740));
    jdff dff_B_WcBNWtOU8_1(.din(n2902), .dout(n13744));
    jdff dff_B_bapi0k3s0_1(.din(n13744), .dout(n13747));
    jdff dff_B_e1ncb7Vw9_1(.din(n13747), .dout(n13750));
    jdff dff_B_ymZyGPr64_1(.din(n13750), .dout(n13753));
    jdff dff_B_ndtNxg8A0_1(.din(n13753), .dout(n13756));
    jdff dff_B_SyvHB0u91_1(.din(n13756), .dout(n13759));
    jdff dff_B_0RGx7qUb3_1(.din(G112), .dout(n13762));
    jdff dff_B_F7iw6GAC2_1(.din(n13762), .dout(n13765));
    jdff dff_A_ewr4SXXH1_0(.din(n13770), .dout(n13767));
    jdff dff_A_atevLuvj3_0(.din(n13773), .dout(n13770));
    jdff dff_A_31nNRVPo0_0(.din(n13776), .dout(n13773));
    jdff dff_A_PTfTAvJb1_0(.din(n20514), .dout(n13776));
    jdff dff_A_hdUzfdID3_1(.din(n13782), .dout(n13779));
    jdff dff_A_vpSkG3G47_1(.din(n20514), .dout(n13782));
    jdff dff_B_3gObBvtq6_1(.din(n4442), .dout(n13786));
    jdff dff_B_7BNYNatJ7_1(.din(n13786), .dout(n13789));
    jdff dff_B_vWtlvFBq7_1(.din(n13789), .dout(n13792));
    jdff dff_B_pal9sUyi5_1(.din(n13792), .dout(n13795));
    jdff dff_B_sxWPdZfA4_1(.din(n13795), .dout(n13798));
    jdff dff_B_pd2DNL1X3_1(.din(n13798), .dout(n13801));
    jdff dff_B_QU100WUX8_1(.din(n13801), .dout(n13804));
    jdff dff_B_27yDHJjp1_1(.din(n13804), .dout(n13807));
    jdff dff_B_tUL6pXNC2_1(.din(n13807), .dout(n13810));
    jdff dff_B_quc5fPgB3_1(.din(n13810), .dout(n13813));
    jdff dff_B_JY4lHCv44_1(.din(n13813), .dout(n13816));
    jdff dff_B_uGKSFA9M9_1(.din(n13816), .dout(n13819));
    jdff dff_B_qZageBzx2_1(.din(n13819), .dout(n13822));
    jdff dff_B_Kqho8I655_1(.din(n13822), .dout(n13825));
    jdff dff_B_zzhyHL5h9_1(.din(n13825), .dout(n13828));
    jdff dff_B_xYUlCryM1_1(.din(n13828), .dout(n13831));
    jdff dff_B_kAxv4aJy7_1(.din(n13831), .dout(n13834));
    jdff dff_B_T6D8dj7o7_1(.din(n13834), .dout(n13837));
    jdff dff_B_jthn2JR95_1(.din(n13837), .dout(n13840));
    jdff dff_B_FMdVkkiS9_1(.din(n3900), .dout(n13843));
    jdff dff_B_RlXyN75Z2_1(.din(n13843), .dout(n13846));
    jdff dff_B_HffqlGeD3_1(.din(n13846), .dout(n13849));
    jdff dff_B_BrRlp7DK5_1(.din(n13849), .dout(n13852));
    jdff dff_B_HtTzx4SS0_1(.din(n13852), .dout(n13855));
    jdff dff_B_g4pXpyvD2_1(.din(n13855), .dout(n13858));
    jdff dff_B_qMC45aoi3_1(.din(n13858), .dout(n13861));
    jdff dff_B_Ryg6WJ9s5_1(.din(n13861), .dout(n13864));
    jdff dff_B_mYKFUuBt2_1(.din(n13864), .dout(n13867));
    jdff dff_B_ODHRcNGn0_1(.din(n13867), .dout(n13870));
    jdff dff_B_WB9zdLi83_1(.din(n13870), .dout(n13873));
    jdff dff_B_VSfgctiF3_1(.din(n13873), .dout(n13876));
    jdff dff_B_h15wSets3_1(.din(n13876), .dout(n13879));
    jdff dff_B_nA4l5icK4_1(.din(n13879), .dout(n13882));
    jdff dff_B_FO7cTvde1_1(.din(n13882), .dout(n13885));
    jdff dff_B_IQtoGsNT7_1(.din(n13885), .dout(n13888));
    jdff dff_B_qgl7C1FO8_1(.din(n3907), .dout(n13891));
    jdff dff_B_BQmwYZ0S5_1(.din(n13891), .dout(n13894));
    jdff dff_B_wmaGa7Tq4_1(.din(n13894), .dout(n13897));
    jdff dff_B_3GEBUdvs2_1(.din(n13897), .dout(n13900));
    jdff dff_B_txWFpU7O5_1(.din(n13900), .dout(n13903));
    jdff dff_B_LLRgr22f0_1(.din(n13903), .dout(n13906));
    jdff dff_B_8WiDnjDU1_1(.din(n13906), .dout(n13909));
    jdff dff_B_4zoGhQZS1_1(.din(n13909), .dout(n13912));
    jdff dff_B_A6XYkeE92_1(.din(n13912), .dout(n13915));
    jdff dff_B_poQmnGEx7_1(.din(n13915), .dout(n13918));
    jdff dff_B_Cp2TkbYB7_1(.din(n13918), .dout(n13921));
    jdff dff_B_rM69akLu3_1(.din(n2765), .dout(n13924));
    jdff dff_B_hhR8mnqz5_1(.din(n13924), .dout(n13927));
    jdff dff_B_M8GRt5Zw8_1(.din(n13927), .dout(n13930));
    jdff dff_B_73a9uzZc8_1(.din(n13930), .dout(n13933));
    jdff dff_B_GNB9tcu21_1(.din(n13933), .dout(n13936));
    jdff dff_B_EzmdNFix3_1(.din(n13936), .dout(n13939));
    jdff dff_B_eInc3zi74_1(.din(n13939), .dout(n13942));
    jdff dff_B_gwymAcpq4_1(.din(n13942), .dout(n13945));
    jdff dff_B_6atzRXp50_1(.din(n13945), .dout(n13948));
    jdff dff_B_0c6LfmK61_1(.din(n1094), .dout(n13951));
    jdff dff_B_yOGDY6he7_1(.din(n1075), .dout(n13954));
    jdff dff_B_DevnYb509_1(.din(G53), .dout(n13957));
    jdff dff_B_3LTRgAEm6_1(.din(n13957), .dout(n13960));
    jdff dff_B_5P3q6PZK0_1(.din(n3755), .dout(n13963));
    jdff dff_B_pKYzJm8L7_1(.din(n13963), .dout(n13966));
    jdff dff_B_gh8tn6QU6_1(.din(n13966), .dout(n13969));
    jdff dff_B_pIKEtVug2_1(.din(n13969), .dout(n13972));
    jdff dff_B_YBUokWUn1_1(.din(n13972), .dout(n13975));
    jdff dff_B_UQh2oZzD2_1(.din(n13975), .dout(n13978));
    jdff dff_B_mLOE9ARC1_1(.din(n13978), .dout(n13981));
    jdff dff_B_7C5wYFeg3_1(.din(n13981), .dout(n13984));
    jdff dff_B_tCXuAXLT7_1(.din(n13984), .dout(n13987));
    jdff dff_B_D6QwLJ9m6_1(.din(n13987), .dout(n13990));
    jdff dff_B_VqM9cSes9_1(.din(n13990), .dout(n13993));
    jdff dff_B_5XZ1CRXX8_1(.din(n13993), .dout(n13996));
    jdff dff_B_GXFxBcp05_1(.din(n13996), .dout(n13999));
    jdff dff_B_QMHplCug2_1(.din(n13999), .dout(n14002));
    jdff dff_B_WPIHHPTY2_1(.din(n14002), .dout(n14005));
    jdff dff_B_kWb1quw83_1(.din(n14005), .dout(n14008));
    jdff dff_B_rEvkE60D6_0(.din(n3770), .dout(n14011));
    jdff dff_B_zINwDq7O3_0(.din(n14011), .dout(n14014));
    jdff dff_B_zQ9aCCvk7_0(.din(n14014), .dout(n14017));
    jdff dff_B_lqbikiFs9_0(.din(n14017), .dout(n14020));
    jdff dff_B_ikIkOiEX1_0(.din(n14020), .dout(n14023));
    jdff dff_B_g8HhNVks3_0(.din(n14023), .dout(n14026));
    jdff dff_B_hZfhGPNm0_0(.din(n14026), .dout(n14029));
    jdff dff_B_JHIZx4mV9_0(.din(n14029), .dout(n14032));
    jdff dff_B_OaAbXU2z9_0(.din(n14032), .dout(n14035));
    jdff dff_B_0wWjNpv39_0(.din(n14035), .dout(n14038));
    jdff dff_B_4kuolSpY5_1(.din(n2866), .dout(n14041));
    jdff dff_B_jz1Kwpoq7_1(.din(n14041), .dout(n14044));
    jdff dff_B_uH0ugx2r4_1(.din(n14044), .dout(n14047));
    jdff dff_B_YLf6kt0O4_1(.din(n14047), .dout(n14050));
    jdff dff_B_ygeRtY650_1(.din(n14050), .dout(n14053));
    jdff dff_B_RSAys7RH0_1(.din(n14053), .dout(n14056));
    jdff dff_B_PGwbWVVH2_1(.din(n14056), .dout(n14059));
    jdff dff_B_FebDitlu7_1(.din(n14059), .dout(n14062));
    jdff dff_B_ICYdCDT54_1(.din(n14062), .dout(n14065));
    jdff dff_B_pyHhzsWM4_1(.din(n2881), .dout(n14068));
    jdff dff_B_MyokzfJG6_1(.din(n2873), .dout(n14071));
    jdff dff_B_qatXc8VV6_1(.din(n14071), .dout(n14074));
    jdff dff_B_5f5v76gk3_1(.din(n14074), .dout(n14077));
    jdff dff_B_9T0J95il7_1(.din(n14077), .dout(n14080));
    jdff dff_B_0D9ogn6Y8_1(.din(n14080), .dout(n14083));
    jdff dff_B_MF9Owc8L0_1(.din(G116), .dout(n14086));
    jdff dff_B_kYjK86vv1_1(.din(n14086), .dout(n14089));
    jdff dff_B_QCQEHJBJ9_0(.din(n4438), .dout(n14092));
    jdff dff_B_NwUqWdPU1_2(.din(G167), .dout(n14095));
    jdff dff_B_KUr6AdJf3_2(.din(G197), .dout(n14098));
    jdff dff_B_6Z1okz4h3_2(.din(n14098), .dout(n14101));
    jdff dff_B_yroClNli2_0(.din(n4494), .dout(n14104));
    jdff dff_B_zdAzHRRF8_0(.din(n14104), .dout(n14107));
    jdff dff_B_6UYEQL2x2_0(.din(n14107), .dout(n14110));
    jdff dff_B_mfpd21pw8_0(.din(n14110), .dout(n14113));
    jdff dff_B_udkTUowa9_0(.din(n14113), .dout(n14116));
    jdff dff_B_hs6jSJjl1_0(.din(n14116), .dout(n14119));
    jdff dff_B_AWSvcsWE1_0(.din(n14119), .dout(n14122));
    jdff dff_B_rz8kvVKx4_0(.din(n14122), .dout(n14125));
    jdff dff_B_m0Oq0xMV3_0(.din(n14125), .dout(n14128));
    jdff dff_B_yYVWrSDQ9_0(.din(n14128), .dout(n14131));
    jdff dff_B_oNLfMOBy9_0(.din(n14131), .dout(n14134));
    jdff dff_B_zHKFq20D8_0(.din(n14134), .dout(n14137));
    jdff dff_B_4W0Uptyo6_0(.din(n14137), .dout(n14140));
    jdff dff_B_7Iq5rWsd2_0(.din(n14140), .dout(n14143));
    jdff dff_B_pMCEaWye6_0(.din(n14143), .dout(n14146));
    jdff dff_B_RssjXhAQ3_0(.din(n14146), .dout(n14149));
    jdff dff_B_8hCC8MqE5_0(.din(n14149), .dout(n14152));
    jdff dff_B_cRRZ9vyq5_0(.din(n14152), .dout(n14155));
    jdff dff_B_aECCcNub3_0(.din(n14155), .dout(n14158));
    jdff dff_B_j1n3kkOT6_0(.din(n4490), .dout(n14161));
    jdff dff_B_shkYsADX0_2(.din(G164), .dout(n14164));
    jdff dff_B_ForsF7Gk3_2(.din(G194), .dout(n14167));
    jdff dff_B_GHXBL6V70_2(.din(n14167), .dout(n14170));
    jdff dff_B_SATYeYta6_1(.din(n4470), .dout(n14173));
    jdff dff_B_IRc6Jqif2_1(.din(n14173), .dout(n14176));
    jdff dff_B_SuASEOwW9_1(.din(n3876), .dout(n14179));
    jdff dff_B_khujN4kz9_1(.din(n14179), .dout(n14182));
    jdff dff_B_F3Kxm83X1_1(.din(n14182), .dout(n14185));
    jdff dff_B_8dQBZvQ76_1(.din(n14185), .dout(n14188));
    jdff dff_B_aQaHBYYT8_1(.din(n14188), .dout(n14191));
    jdff dff_B_tlWiEksU1_1(.din(n14191), .dout(n14194));
    jdff dff_B_V4g9B0Bc1_1(.din(n14194), .dout(n14197));
    jdff dff_B_4IMke6an4_1(.din(n14197), .dout(n14200));
    jdff dff_B_is8T0Zvx8_1(.din(n14200), .dout(n14203));
    jdff dff_B_uY0k4gIV8_1(.din(n14203), .dout(n14206));
    jdff dff_B_p4AXBXKC0_1(.din(n14206), .dout(n14209));
    jdff dff_B_NTB3WyIr9_1(.din(n14209), .dout(n14212));
    jdff dff_B_KGmhtZ5V7_1(.din(n14212), .dout(n14215));
    jdff dff_B_jXg2uAaj1_1(.din(n14215), .dout(n14218));
    jdff dff_B_gDMHa5dD1_0(.din(n3888), .dout(n14221));
    jdff dff_B_hnlt39in2_0(.din(n14221), .dout(n14224));
    jdff dff_B_CzjmnqsG2_0(.din(n14224), .dout(n14227));
    jdff dff_B_Uk6SWWo31_0(.din(n14227), .dout(n14230));
    jdff dff_B_amk12isJ4_0(.din(n14230), .dout(n14233));
    jdff dff_B_aqHn981c9_0(.din(n14233), .dout(n14236));
    jdff dff_B_TOhZOnpB9_0(.din(n14236), .dout(n14239));
    jdff dff_B_Y2HgL4gd1_0(.din(n14239), .dout(n14242));
    jdff dff_B_JAOvdGPG3_0(.din(n14242), .dout(n14245));
    jdff dff_B_Vhmy5KCT8_0(.din(n14245), .dout(n14248));
    jdff dff_A_HArAgng82_1(.din(n14253), .dout(n14250));
    jdff dff_A_M0jMOAI95_1(.din(n14256), .dout(n14253));
    jdff dff_A_9OEWihJg9_1(.din(n888), .dout(n14256));
    jdff dff_B_2TSL03jK6_1(.din(n872), .dout(n14260));
    jdff dff_B_q9Ly9YM44_3(.din(G3548), .dout(n14263));
    jdff dff_B_cRRncVaF6_1(.din(n853), .dout(n14266));
    jdff dff_A_VoJQY4mK5_0(.din(n14271), .dout(n14268));
    jdff dff_A_zOK6Sc6G1_0(.din(n14274), .dout(n14271));
    jdff dff_A_W72xPigz0_0(.din(n14277), .dout(n14274));
    jdff dff_A_XUWvpTXo5_0(.din(n14280), .dout(n14277));
    jdff dff_A_7EGXfocg3_0(.din(n14283), .dout(n14280));
    jdff dff_A_jj5mAno66_0(.din(n14286), .dout(n14283));
    jdff dff_A_aKgZac1K6_0(.din(n14289), .dout(n14286));
    jdff dff_A_mDIJjcnI8_0(.din(n14292), .dout(n14289));
    jdff dff_A_moObGmSF6_0(.din(n14295), .dout(n14292));
    jdff dff_A_2m1qgmXz6_0(.din(n14298), .dout(n14295));
    jdff dff_A_O9OK7o6x9_0(.din(n19698), .dout(n14298));
    jdff dff_A_09PEiPU34_1(.din(n14304), .dout(n14301));
    jdff dff_A_uXdx9I4O0_1(.din(n2758), .dout(n14304));
    jdff dff_B_9fTv7oJp4_1(.din(n2746), .dout(n14308));
    jdff dff_B_c0RnFSPh6_1(.din(n14308), .dout(n14311));
    jdff dff_B_Wu4ANowT3_1(.din(n14311), .dout(n14314));
    jdff dff_B_Eq7yUAjh0_1(.din(n14314), .dout(n14317));
    jdff dff_B_zqJrC4xK2_1(.din(n14317), .dout(n14320));
    jdff dff_B_YgrLRGQT5_1(.din(n14320), .dout(n14323));
    jdff dff_A_yPdgnVZq1_0(.din(n14328), .dout(n14325));
    jdff dff_A_EQO7aPUZ7_0(.din(n19785), .dout(n14328));
    jdff dff_A_Sdgvmiav8_1(.din(n14334), .dout(n14331));
    jdff dff_A_IFemFwP97_1(.din(n14337), .dout(n14334));
    jdff dff_A_DB8a6sF52_1(.din(n19785), .dout(n14337));
    jdff dff_B_babhDdva3_1(.din(G114), .dout(n14341));
    jdff dff_B_Or80r8Bu4_1(.din(n14341), .dout(n14344));
    jdff dff_A_bDAjTJQY5_0(.din(n20109), .dout(n14346));
    jdff dff_A_5i6QK7o84_1(.din(n20109), .dout(n14349));
    jdff dff_B_50hXFk5M3_1(.din(n3722), .dout(n14353));
    jdff dff_B_FFfn2ho82_1(.din(n14353), .dout(n14356));
    jdff dff_B_SIN1FyzY3_1(.din(n14356), .dout(n14359));
    jdff dff_B_Yu8UBpLi6_1(.din(n14359), .dout(n14362));
    jdff dff_B_xWGtZ0OT7_1(.din(n14362), .dout(n14365));
    jdff dff_B_Kmxdsp1M9_1(.din(n14365), .dout(n14368));
    jdff dff_B_R9w9evNC0_1(.din(n14368), .dout(n14371));
    jdff dff_B_6JhyAsAc9_1(.din(n14371), .dout(n14374));
    jdff dff_B_AGGg2M6Z2_1(.din(n14374), .dout(n14377));
    jdff dff_B_cFioTv9R6_1(.din(n14377), .dout(n14380));
    jdff dff_B_wFZP9U8Z9_1(.din(n14380), .dout(n14383));
    jdff dff_B_oMLOhkRf6_1(.din(n14383), .dout(n14386));
    jdff dff_B_e3JhcnfG7_1(.din(n14386), .dout(n14389));
    jdff dff_B_ot4T40aM7_1(.din(n14389), .dout(n14392));
    jdff dff_B_UZUkPoFP0_1(.din(n14392), .dout(n14395));
    jdff dff_B_dmjTBYiW3_1(.din(n3729), .dout(n14398));
    jdff dff_B_zaz4tCVY8_1(.din(n14398), .dout(n14401));
    jdff dff_B_neIGb0Nn7_1(.din(n14401), .dout(n14404));
    jdff dff_B_w0ha3GHo1_1(.din(n14404), .dout(n14407));
    jdff dff_B_iyvx0Osu3_1(.din(n14407), .dout(n14410));
    jdff dff_B_ypEKkKHu1_1(.din(n14410), .dout(n14413));
    jdff dff_B_1HBEN5Er7_1(.din(n14413), .dout(n14416));
    jdff dff_B_9orisDh76_1(.din(n14416), .dout(n14419));
    jdff dff_B_NwbyyCxe4_1(.din(n14419), .dout(n14422));
    jdff dff_B_ovtLENyn1_1(.din(n14422), .dout(n14425));
    jdff dff_B_TA9c7iQR3_1(.din(n14425), .dout(n14428));
    jdff dff_A_KpkyMcK08_0(.din(n14433), .dout(n14430));
    jdff dff_A_AIMvmSNJ1_0(.din(n14436), .dout(n14433));
    jdff dff_A_uAYq9qwW0_0(.din(n14439), .dout(n14436));
    jdff dff_A_sXdHsCJz1_0(.din(n14442), .dout(n14439));
    jdff dff_A_Sp5I7ldP9_0(.din(n14445), .dout(n14442));
    jdff dff_A_vqtaKSFB4_0(.din(n14448), .dout(n14445));
    jdff dff_A_mlYvGYp88_0(.din(n14451), .dout(n14448));
    jdff dff_A_BDO4lIXq1_0(.din(n14454), .dout(n14451));
    jdff dff_A_M55HYp4e6_0(.din(n1613), .dout(n14454));
    jdff dff_A_5CRQ0zB80_1(.din(n14460), .dout(n14457));
    jdff dff_A_jES8ImbP5_1(.din(n14463), .dout(n14460));
    jdff dff_A_g6TZUcjN9_1(.din(n14466), .dout(n14463));
    jdff dff_A_rH4vGzSu7_1(.din(n14469), .dout(n14466));
    jdff dff_A_l22ymRVk8_1(.din(n14472), .dout(n14469));
    jdff dff_A_r41c0YZ74_1(.din(n14475), .dout(n14472));
    jdff dff_A_tsD94GUS7_1(.din(n14478), .dout(n14475));
    jdff dff_A_usWIVe4r6_1(.din(n14481), .dout(n14478));
    jdff dff_A_VbB6nsO87_1(.din(n14484), .dout(n14481));
    jdff dff_A_Gm075tNU0_1(.din(n14487), .dout(n14484));
    jdff dff_A_8x7QodEG0_1(.din(n14490), .dout(n14487));
    jdff dff_A_GPQp5Te57_1(.din(n15189), .dout(n14490));
    jdff dff_A_MpLo72ts6_2(.din(n14496), .dout(n14493));
    jdff dff_A_3E1I7apd9_2(.din(n14499), .dout(n14496));
    jdff dff_A_gY5xpIeV8_2(.din(n14502), .dout(n14499));
    jdff dff_A_DFk1rNYC3_2(.din(n14505), .dout(n14502));
    jdff dff_A_9YSRrLIq5_2(.din(n14508), .dout(n14505));
    jdff dff_A_ceGm2RIz5_2(.din(n14511), .dout(n14508));
    jdff dff_A_khqusC305_2(.din(n14514), .dout(n14511));
    jdff dff_A_ZIh2Izqh5_2(.din(n14517), .dout(n14514));
    jdff dff_A_oOh3FEj50_2(.din(n14520), .dout(n14517));
    jdff dff_A_kRe9C1FU2_2(.din(n15189), .dout(n14520));
    jdff dff_B_2Ko6HozK1_1(.din(G121), .dout(n14524));
    jdff dff_B_4nhfmZyy7_1(.din(n14524), .dout(n14527));
    jdff dff_A_kCA1roIz8_0(.din(n14535), .dout(n14529));
    jdff dff_A_Ii9nEp3G4_1(.din(n14535), .dout(n14532));
    jdff dff_A_Uantm8hy6_0(.din(n14538), .dout(n14535));
    jdff dff_A_EvlWgjHm5_0(.din(n14541), .dout(n14538));
    jdff dff_A_zFhXjUh34_0(.din(n14544), .dout(n14541));
    jdff dff_A_5SjB4z280_0(.din(n14547), .dout(n14544));
    jdff dff_A_GTGvGoaV3_0(.din(n14550), .dout(n14547));
    jdff dff_A_9SF0wWVx1_0(.din(n20706), .dout(n14550));
    jdff dff_A_5UICh8js7_1(.din(n14556), .dout(n14553));
    jdff dff_A_fvgm4vOr9_1(.din(n14559), .dout(n14556));
    jdff dff_A_jFoquQJb9_1(.din(n14562), .dout(n14559));
    jdff dff_A_rm8v5iUM7_1(.din(n14565), .dout(n14562));
    jdff dff_A_rqTSfhJM6_1(.din(n14568), .dout(n14565));
    jdff dff_A_ViVAQnti7_1(.din(n14571), .dout(n14568));
    jdff dff_A_z3v7vRp71_1(.din(n20706), .dout(n14571));
    jdff dff_B_IaT2PVUl3_0(.din(n4530), .dout(n14575));
    jdff dff_B_OPohOdCj5_0(.din(n14575), .dout(n14578));
    jdff dff_B_Sz85MPJU5_0(.din(n14578), .dout(n14581));
    jdff dff_B_aKXskUcH3_0(.din(n14581), .dout(n14584));
    jdff dff_B_9uX8harz7_0(.din(n14584), .dout(n14587));
    jdff dff_B_9QUziSNQ6_0(.din(n14587), .dout(n14590));
    jdff dff_B_dhOeJycN7_0(.din(n14590), .dout(n14593));
    jdff dff_B_jBhjZjjS2_0(.din(n14593), .dout(n14596));
    jdff dff_B_57gpdxxg8_0(.din(n14596), .dout(n14599));
    jdff dff_B_0MA2VM3V0_0(.din(n14599), .dout(n14602));
    jdff dff_B_9qarWJfO7_0(.din(n14602), .dout(n14605));
    jdff dff_B_ijD61zwB8_0(.din(n14605), .dout(n14608));
    jdff dff_B_bkfVty1l4_0(.din(n14608), .dout(n14611));
    jdff dff_B_5qIDoWML4_0(.din(n14611), .dout(n14614));
    jdff dff_B_w3f5EaIq8_0(.din(n14614), .dout(n14617));
    jdff dff_B_NRyAP7tH3_0(.din(n14617), .dout(n14620));
    jdff dff_B_fzndBmR54_0(.din(n14620), .dout(n14623));
    jdff dff_B_l1DuayOK1_0(.din(n14623), .dout(n14626));
    jdff dff_B_80SRCvM26_0(.din(n14626), .dout(n14629));
    jdff dff_B_E3wrtXIv4_0(.din(n4526), .dout(n14632));
    jdff dff_B_ZoSLA8cb9_2(.din(G161), .dout(n14635));
    jdff dff_B_7uLmyHdV4_2(.din(G191), .dout(n14638));
    jdff dff_B_fGuvLndO3_2(.din(n14638), .dout(n14641));
    jdff dff_B_V0qgLHDs2_1(.din(n3692), .dout(n14644));
    jdff dff_B_9KWmcCOm7_1(.din(n14644), .dout(n14647));
    jdff dff_B_f1VurmMl8_1(.din(n14647), .dout(n14650));
    jdff dff_B_N78XHgTI0_1(.din(n14650), .dout(n14653));
    jdff dff_B_TihVkcu21_1(.din(n14653), .dout(n14656));
    jdff dff_B_8gj5Y2tG9_1(.din(n14656), .dout(n14659));
    jdff dff_B_YJDpsx4H3_1(.din(n14659), .dout(n14662));
    jdff dff_B_HCH1NubT5_1(.din(n14662), .dout(n14665));
    jdff dff_B_XW4WyXIR5_1(.din(n14665), .dout(n14668));
    jdff dff_B_CelSJfSW6_1(.din(n14668), .dout(n14671));
    jdff dff_B_fAe2TAn28_1(.din(n14671), .dout(n14674));
    jdff dff_B_8qwtpWrV4_1(.din(n14674), .dout(n14677));
    jdff dff_B_V4Ppvtsg0_1(.din(n14677), .dout(n14680));
    jdff dff_B_34MWWBSD3_1(.din(n14680), .dout(n14683));
    jdff dff_B_G67N6VPI7_1(.din(n14683), .dout(n14686));
    jdff dff_B_BGM5W6S45_1(.din(n14686), .dout(n14689));
    jdff dff_B_GKfzRS3d7_0(.din(n3707), .dout(n14692));
    jdff dff_B_VzNzpOiO9_0(.din(n14692), .dout(n14695));
    jdff dff_B_lJ3dHqQx5_0(.din(n14695), .dout(n14698));
    jdff dff_B_QVsNxBfM1_0(.din(n14698), .dout(n14701));
    jdff dff_B_Tzipyeb02_0(.din(n14701), .dout(n14704));
    jdff dff_B_eD5iR0z97_0(.din(n14704), .dout(n14707));
    jdff dff_B_jZNhevm24_0(.din(n14707), .dout(n14710));
    jdff dff_B_yv72Z9yD3_0(.din(n14710), .dout(n14713));
    jdff dff_B_aXOr8GyN4_0(.din(n14713), .dout(n14716));
    jdff dff_B_VmEIurYj1_0(.din(n14716), .dout(n14719));
    jdff dff_B_WLwvlIPA5_0(.din(n14719), .dout(n14722));
    jdff dff_B_s4WOZmBm6_0(.din(n14722), .dout(n14725));
    jdff dff_A_BH3rsD105_1(.din(n14730), .dout(n14727));
    jdff dff_A_rLeApYgQ2_1(.din(n18183), .dout(n14730));
    jdff dff_A_nymskFp84_2(.din(n14736), .dout(n14733));
    jdff dff_A_Zoy8pnXB4_2(.din(n18183), .dout(n14736));
    jdff dff_B_7CzP2E2L3_0(.din(n2168), .dout(n14740));
    jdff dff_B_m8lrl0n79_0(.din(n2135), .dout(n14743));
    jdff dff_A_BmOSzjts1_0(.din(n14748), .dout(n14745));
    jdff dff_A_sGehzmu81_0(.din(n14751), .dout(n14748));
    jdff dff_A_Rni5PH7f7_0(.din(n14754), .dout(n14751));
    jdff dff_A_u0eNrmBu4_0(.din(n14757), .dout(n14754));
    jdff dff_A_GbWrzrA04_0(.din(n14760), .dout(n14757));
    jdff dff_A_dgYS5rF39_0(.din(n14763), .dout(n14760));
    jdff dff_A_HKIO64mQ1_0(.din(n14766), .dout(n14763));
    jdff dff_A_6WBjMV9a8_0(.din(n14769), .dout(n14766));
    jdff dff_A_IjOfffxg2_0(.din(G54), .dout(n14769));
    jdff dff_A_5zH7QhnH9_1(.din(n14775), .dout(n14772));
    jdff dff_A_wJ3Ouuzb5_1(.din(n14778), .dout(n14775));
    jdff dff_A_WbcQvHDP1_1(.din(n14781), .dout(n14778));
    jdff dff_A_w3gOLomI2_1(.din(G54), .dout(n14781));
    jdff dff_A_NxClbYBH0_0(.din(n19710), .dout(n14784));
    jdff dff_A_1Dx4HAHp7_2(.din(n14790), .dout(n14787));
    jdff dff_A_qso3eQg61_2(.din(n14793), .dout(n14790));
    jdff dff_A_xQg7Be0V8_2(.din(n14796), .dout(n14793));
    jdff dff_A_UcqKxuSJ8_2(.din(n14799), .dout(n14796));
    jdff dff_A_oZwZOjGH5_2(.din(n14802), .dout(n14799));
    jdff dff_A_xj9gEQvJ1_2(.din(n14805), .dout(n14802));
    jdff dff_A_eLxW5qXp5_2(.din(n14808), .dout(n14805));
    jdff dff_A_1CdI0S0G6_2(.din(n14811), .dout(n14808));
    jdff dff_A_rdRbeQpz7_2(.din(n14814), .dout(n14811));
    jdff dff_A_DKIsNxmh3_2(.din(n14817), .dout(n14814));
    jdff dff_A_tFqvLuoQ2_2(.din(n14820), .dout(n14817));
    jdff dff_A_nnfxkria6_2(.din(n14823), .dout(n14820));
    jdff dff_A_LFp7k7aZ3_2(.din(n14826), .dout(n14823));
    jdff dff_A_aOqhSAk29_2(.din(n19710), .dout(n14826));
    jdff dff_A_u5tFlz3S7_0(.din(n14832), .dout(n14829));
    jdff dff_A_bJ19DS6e9_0(.din(G123), .dout(n14832));
    jdff dff_A_phMaxgek3_0(.din(n20457), .dout(n14835));
    jdff dff_A_4i0Tqhj48_2(.din(n20457), .dout(n14838));
    jdff dff_A_0YtcJIVr1_2(.din(n14844), .dout(n14841));
    jdff dff_A_5ZHG9g6R5_0(.din(n14847), .dout(n14844));
    jdff dff_A_wfRDHPzP8_0(.din(n14850), .dout(n14847));
    jdff dff_A_hD979AwS9_0(.din(n14853), .dout(n14850));
    jdff dff_A_9HBBF0OZ2_0(.din(n14856), .dout(n14853));
    jdff dff_A_kNJtKEVH1_0(.din(n14859), .dout(n14856));
    jdff dff_A_A93dWc351_0(.din(n14862), .dout(n14859));
    jdff dff_A_1fpD5eUO1_0(.din(n14865), .dout(n14862));
    jdff dff_A_1UH77wLh7_0(.din(n14868), .dout(n14865));
    jdff dff_A_H4V82B3V1_0(.din(n14908), .dout(n14868));
    jdff dff_A_DKLNwFK66_1(.din(n14874), .dout(n14871));
    jdff dff_A_u2T2DKa28_1(.din(n14908), .dout(n14874));
    jdff dff_B_7eAZoxY13_3(.din(n2975), .dout(n14878));
    jdff dff_B_CWRxvdPn2_3(.din(n14878), .dout(n14881));
    jdff dff_B_4g4Q6Rvf1_3(.din(n14881), .dout(n14884));
    jdff dff_B_7pfkPapK2_3(.din(n14884), .dout(n14887));
    jdff dff_B_IGDUEajs0_3(.din(n14887), .dout(n14890));
    jdff dff_B_wcC1iBGy8_3(.din(n14890), .dout(n14893));
    jdff dff_B_ylLpoCZ65_3(.din(n14893), .dout(n14896));
    jdff dff_B_dQiEg0El9_3(.din(n14896), .dout(n14899));
    jdff dff_B_sJ1C3hQo8_3(.din(n14899), .dout(n14902));
    jdff dff_B_gaPX4nAc7_3(.din(n14902), .dout(n14905));
    jdff dff_B_djOsCc3g3_3(.din(n14905), .dout(n14908));
    jdff dff_B_FHX8TLny0_1(.din(n3843), .dout(n14911));
    jdff dff_B_P19qavdH1_1(.din(n14911), .dout(n14914));
    jdff dff_B_ycbutOvK2_1(.din(n14914), .dout(n14917));
    jdff dff_B_Soo3w26k1_1(.din(n14917), .dout(n14920));
    jdff dff_B_7pt7jynQ8_1(.din(n14920), .dout(n14923));
    jdff dff_B_mZSUNb9g1_1(.din(n14923), .dout(n14926));
    jdff dff_B_NBxSAoRi8_1(.din(n14926), .dout(n14929));
    jdff dff_B_n9wQfuIa9_1(.din(n14929), .dout(n14932));
    jdff dff_B_njhLuD006_1(.din(n14932), .dout(n14935));
    jdff dff_B_SohIp7eS4_1(.din(n14935), .dout(n14938));
    jdff dff_B_VEGbVZ7T5_1(.din(n14938), .dout(n14941));
    jdff dff_B_hel2dOG81_1(.din(n14941), .dout(n14944));
    jdff dff_B_tX8kMrfL6_1(.din(n14944), .dout(n14947));
    jdff dff_B_mlc6LtcC8_1(.din(n14947), .dout(n14950));
    jdff dff_B_5faaRwDs5_1(.din(n14950), .dout(n14953));
    jdff dff_B_HTpe1VCg2_1(.din(n14953), .dout(n14956));
    jdff dff_B_0Z5IiwPq7_1(.din(n14956), .dout(n14959));
    jdff dff_B_BjCTQoto0_1(.din(n3850), .dout(n14962));
    jdff dff_B_VckX4ovK6_1(.din(n14962), .dout(n14965));
    jdff dff_B_MbvjTpVM5_1(.din(n14965), .dout(n14968));
    jdff dff_B_LA1x1T553_1(.din(n14968), .dout(n14971));
    jdff dff_B_DEk286bu7_1(.din(n14971), .dout(n14974));
    jdff dff_B_9V0H138A9_1(.din(n14974), .dout(n14977));
    jdff dff_B_Ghu6kiR09_1(.din(n14977), .dout(n14980));
    jdff dff_B_L9lWMhdF2_1(.din(n14980), .dout(n14983));
    jdff dff_B_o8GKBQRI7_1(.din(n14983), .dout(n14986));
    jdff dff_B_iWhCo6B03_1(.din(n14986), .dout(n14989));
    jdff dff_B_i48UCTAL8_1(.din(n14989), .dout(n14992));
    jdff dff_B_E104wsN56_1(.din(n14992), .dout(n14995));
    jdff dff_B_GCUTKeC38_1(.din(n2714), .dout(n14998));
    jdff dff_B_pdUuINJl0_1(.din(n14998), .dout(n15001));
    jdff dff_B_UpfYWGsR2_1(.din(n15001), .dout(n15004));
    jdff dff_B_K3RuSd0b4_1(.din(n15004), .dout(n15007));
    jdff dff_B_4gLCdTGb0_1(.din(n15007), .dout(n15010));
    jdff dff_B_pOTZXhRw8_1(.din(n15010), .dout(n15013));
    jdff dff_B_TULGqpbe4_1(.din(n15013), .dout(n15016));
    jdff dff_B_r2KtQKQg4_1(.din(n15016), .dout(n15019));
    jdff dff_B_rLWnffD82_1(.din(n15019), .dout(n15022));
    jdff dff_B_pJBymsxM6_1(.din(n15022), .dout(n15025));
    jdff dff_B_ulWuoMYT0_1(.din(n15025), .dout(n15028));
    jdff dff_B_1etY6Mwd5_0(.din(n2451), .dout(n15031));
    jdff dff_B_GEUE8hrs9_1(.din(n2439), .dout(n15034));
    jdff dff_B_9UXiCv0m5_1(.din(n15034), .dout(n15037));
    jdff dff_A_zhbpJqqR3_1(.din(n15055), .dout(n15039));
    jdff dff_B_Djb85jzw6_3(.din(G4), .dout(n15043));
    jdff dff_B_XbMfPNC78_3(.din(n15043), .dout(n15046));
    jdff dff_B_kXpySNY15_3(.din(n15046), .dout(n15049));
    jdff dff_B_7lgsNG6L1_3(.din(n15049), .dout(n15052));
    jdff dff_B_3BFNaT9z0_3(.din(n15052), .dout(n15055));
    jdff dff_A_nshC9MZh4_0(.din(n15109), .dout(n15057));
    jdff dff_A_ZLrIieCK1_1(.din(n15063), .dout(n15060));
    jdff dff_A_Tjcoy3949_1(.din(n15109), .dout(n15063));
    jdff dff_B_6soiylNA4_3(.din(n3732), .dout(n15067));
    jdff dff_B_gaxXnFkz7_3(.din(n15067), .dout(n15070));
    jdff dff_B_D6GWk81n4_3(.din(n15070), .dout(n15073));
    jdff dff_B_hKojJ9Rp0_3(.din(n15073), .dout(n15076));
    jdff dff_B_KLBHPtCb3_3(.din(n15076), .dout(n15079));
    jdff dff_B_boVhpqj27_3(.din(n15079), .dout(n15082));
    jdff dff_B_x6UQqVXX7_3(.din(n15082), .dout(n15085));
    jdff dff_B_7XORGzGK5_3(.din(n15085), .dout(n15088));
    jdff dff_B_nu7RB4Nl2_3(.din(n15088), .dout(n15091));
    jdff dff_B_XZuJ79wq8_3(.din(n15091), .dout(n15094));
    jdff dff_B_TJkDqrhs3_3(.din(n15094), .dout(n15097));
    jdff dff_B_3PiQHyt39_3(.din(n15097), .dout(n15100));
    jdff dff_B_oqp7mgxB8_3(.din(n15100), .dout(n15103));
    jdff dff_B_G1XF9B541_3(.din(n15103), .dout(n15106));
    jdff dff_B_Vg4hOFcp5_3(.din(n15106), .dout(n15109));
    jdff dff_A_LypQKKcW0_0(.din(n15114), .dout(n15111));
    jdff dff_A_yXRHn23c6_0(.din(n15117), .dout(n15114));
    jdff dff_A_kAPst4rG7_0(.din(n15120), .dout(n15117));
    jdff dff_A_olHE7vfl9_0(.din(n15123), .dout(n15120));
    jdff dff_A_LWuJLPGe4_0(.din(n15126), .dout(n15123));
    jdff dff_A_93243qg33_0(.din(G4092), .dout(n15126));
    jdff dff_A_L9n2n8oJ8_1(.din(n15132), .dout(n15129));
    jdff dff_A_edaGDRxl6_1(.din(n15135), .dout(n15132));
    jdff dff_A_Z4Y8e3Fm2_1(.din(n15138), .dout(n15135));
    jdff dff_A_2jivuVoV2_1(.din(n15141), .dout(n15138));
    jdff dff_A_vYseTm2Q7_1(.din(n15144), .dout(n15141));
    jdff dff_A_N2iAANj73_1(.din(G4092), .dout(n15144));
    jdff dff_A_tdTttx1A4_0(.din(n15150), .dout(n15147));
    jdff dff_A_6TS6vlq43_0(.din(n15153), .dout(n15150));
    jdff dff_A_UnODfP1e7_0(.din(n15156), .dout(n15153));
    jdff dff_A_AA0Aec4E5_0(.din(n15159), .dout(n15156));
    jdff dff_A_pg1yx1tx3_0(.din(n15162), .dout(n15159));
    jdff dff_A_vqeYpe6u4_0(.din(n15165), .dout(n15162));
    jdff dff_A_T1XhDIww2_0(.din(n15168), .dout(n15165));
    jdff dff_A_riKcW56x8_0(.din(n15171), .dout(n15168));
    jdff dff_A_nmRawhVX0_0(.din(n15174), .dout(n15171));
    jdff dff_A_orhdBHcl5_0(.din(n15177), .dout(n15174));
    jdff dff_A_KUKgTNlP7_0(.din(n15180), .dout(n15177));
    jdff dff_A_jhT5jWgK2_0(.din(n15183), .dout(n15180));
    jdff dff_A_fZvtdc804_0(.din(n15186), .dout(n15183));
    jdff dff_A_UGEY9o3W6_0(.din(n19710), .dout(n15186));
    jdff dff_A_2WSEciTN5_1(.din(n15192), .dout(n15189));
    jdff dff_A_r6mjsyH68_1(.din(n19710), .dout(n15192));
    jdff dff_B_Ehju4Z324_1(.din(G115), .dout(n15196));
    jdff dff_B_uKlhyMAY6_1(.din(n15196), .dout(n15199));
    jdff dff_B_wDrfRkwT3_0(.din(n4923), .dout(n15202));
    jdff dff_B_Cwc16hRW5_0(.din(n15202), .dout(n15205));
    jdff dff_B_vWWfOqqQ9_0(.din(n15205), .dout(n15208));
    jdff dff_B_D5UDEj6N8_0(.din(n15208), .dout(n15211));
    jdff dff_B_bzNCjmpl3_0(.din(n15211), .dout(n15214));
    jdff dff_B_dLbIVf7M8_0(.din(n15214), .dout(n15217));
    jdff dff_B_3o1tM25u3_0(.din(n15217), .dout(n15220));
    jdff dff_B_SOWLTAqs1_0(.din(n15220), .dout(n15223));
    jdff dff_B_L4TOTHkU6_0(.din(n15223), .dout(n15226));
    jdff dff_B_AvUsMNqQ5_0(.din(n15226), .dout(n15229));
    jdff dff_B_qosWfwVb2_0(.din(n15229), .dout(n15232));
    jdff dff_B_0EAHIAn80_0(.din(n15232), .dout(n15235));
    jdff dff_B_4saqOU3Y3_0(.din(n15235), .dout(n15238));
    jdff dff_B_Ec75XCn20_0(.din(n15238), .dout(n15241));
    jdff dff_B_HvZxSwsH1_0(.din(n15241), .dout(n15244));
    jdff dff_B_1Y5pUuUD6_0(.din(n15244), .dout(n15247));
    jdff dff_B_ow9X3H7R6_0(.din(n15247), .dout(n15250));
    jdff dff_B_us0caNch4_1(.din(G120), .dout(n15253));
    jdff dff_B_OIAyBtWZ3_1(.din(n15253), .dout(n15256));
    jdff dff_B_qS653Y2i8_1(.din(n15256), .dout(n15259));
    jdff dff_B_o2XB3q0z2_0(.din(n5556), .dout(n15262));
    jdff dff_B_N02CtFAU5_0(.din(n15262), .dout(n15265));
    jdff dff_B_y3ymCFBe5_0(.din(n15265), .dout(n15268));
    jdff dff_B_N5YZXX2n3_0(.din(n15268), .dout(n15271));
    jdff dff_B_GVlPamiQ3_0(.din(n15271), .dout(n15274));
    jdff dff_B_BIpqgLrW3_0(.din(n15274), .dout(n15277));
    jdff dff_B_gFIt59JH6_0(.din(n15277), .dout(n15280));
    jdff dff_B_cNBuyqeU3_0(.din(n15280), .dout(n15283));
    jdff dff_B_t8gWkXLY8_0(.din(n15283), .dout(n15286));
    jdff dff_B_SPPxYmft4_0(.din(n15286), .dout(n15289));
    jdff dff_B_JMA2Ojso9_0(.din(n15289), .dout(n15292));
    jdff dff_B_bdhzgnpS6_0(.din(n15292), .dout(n15295));
    jdff dff_B_5yvKG2eJ0_0(.din(n15295), .dout(n15298));
    jdff dff_B_I2IkDyHH9_0(.din(n15298), .dout(n15301));
    jdff dff_B_61X5ZuyU4_0(.din(n15301), .dout(n15304));
    jdff dff_B_NaYOdTpP1_0(.din(n15304), .dout(n15307));
    jdff dff_B_9NRyjmDE9_0(.din(n15307), .dout(n15310));
    jdff dff_B_PBRsEGmR6_1(.din(G118), .dout(n15313));
    jdff dff_B_1u8wWBmn5_1(.din(n15313), .dout(n15316));
    jdff dff_B_E0dWacZS0_1(.din(n15316), .dout(n15319));
    jdff dff_A_YlAgmg6T7_0(.din(n15324), .dout(n15321));
    jdff dff_A_rcfcSIjf5_0(.din(n15327), .dout(n15324));
    jdff dff_A_Jn97mrZK5_0(.din(n15330), .dout(n15327));
    jdff dff_A_C4NNP8Xo9_0(.din(n15333), .dout(n15330));
    jdff dff_A_5lvsBwnu3_0(.din(n19908), .dout(n15333));
    jdff dff_A_xfi47aKt6_1(.din(n15339), .dout(n15336));
    jdff dff_A_XX8s0kTl5_1(.din(n15342), .dout(n15339));
    jdff dff_A_wcH6QTuZ3_1(.din(n15345), .dout(n15342));
    jdff dff_A_R2cCntsR9_1(.din(n19908), .dout(n15345));
    jdff dff_A_2ThLU8My3_0(.din(n15351), .dout(n15348));
    jdff dff_A_PUvMD4Qh7_0(.din(n15354), .dout(n15351));
    jdff dff_A_0T5gnU6g4_0(.din(n15357), .dout(n15354));
    jdff dff_A_RIoXXCcc6_0(.din(n15360), .dout(n15357));
    jdff dff_A_Rcqv1pnE6_0(.din(n19908), .dout(n15360));
    jdff dff_A_mFeMHTtF2_1(.din(n15366), .dout(n15363));
    jdff dff_A_v7kFF0zp0_1(.din(n15369), .dout(n15366));
    jdff dff_A_KkthLwDo4_1(.din(n15372), .dout(n15369));
    jdff dff_A_u4fEX5Gh2_1(.din(n19908), .dout(n15372));
    jdff dff_A_6vxKppbj8_0(.din(n15378), .dout(n15375));
    jdff dff_A_Q1y0rw1J0_0(.din(n15381), .dout(n15378));
    jdff dff_A_MYjoLYpB8_0(.din(n1999), .dout(n15381));
    jdff dff_B_zEo4q6Xh3_1(.din(n5576), .dout(n15385));
    jdff dff_B_BJBS0wp33_1(.din(n15385), .dout(n15388));
    jdff dff_B_nsg6w8Jg1_1(.din(n15388), .dout(n15391));
    jdff dff_B_9DeTDEkl1_1(.din(n15391), .dout(n15394));
    jdff dff_B_eqHr8K7Z4_1(.din(n15394), .dout(n15397));
    jdff dff_B_m6uGQahr0_1(.din(n15397), .dout(n15400));
    jdff dff_B_w4OiuBEM4_1(.din(n15400), .dout(n15403));
    jdff dff_B_uGzj4GnF2_1(.din(n15403), .dout(n15406));
    jdff dff_B_Cu8AVbP31_1(.din(n15406), .dout(n15409));
    jdff dff_B_3T8p3AbB2_1(.din(n15409), .dout(n15412));
    jdff dff_B_bSBCFu0d3_1(.din(n15412), .dout(n15415));
    jdff dff_B_cMV8N3sX5_1(.din(n15415), .dout(n15418));
    jdff dff_B_8oSCkhnx1_1(.din(n15418), .dout(n15421));
    jdff dff_B_pvphTkoP5_1(.din(n15421), .dout(n15424));
    jdff dff_B_P2UAXcJf8_1(.din(n15424), .dout(n15427));
    jdff dff_B_d6bv0RBw7_1(.din(n15427), .dout(n15430));
    jdff dff_B_YPFyJM4S1_1(.din(n15430), .dout(n15433));
    jdff dff_B_eiqe9rVO8_1(.din(n15433), .dout(n15436));
    jdff dff_B_u3QlNxvx7_1(.din(n15436), .dout(n15439));
    jdff dff_B_tirUx62I2_1(.din(n15439), .dout(n15442));
    jdff dff_B_rxo2Dayk1_1(.din(n15442), .dout(n15445));
    jdff dff_B_DQdEZMtx8_1(.din(n15445), .dout(n15448));
    jdff dff_B_Xab86eH79_1(.din(n5594), .dout(n15451));
    jdff dff_A_hdXM7sbV1_1(.din(n15456), .dout(n15453));
    jdff dff_A_Z0m7DK4o2_1(.din(n15459), .dout(n15456));
    jdff dff_A_Q03PM3lt4_1(.din(n15462), .dout(n15459));
    jdff dff_A_YmGFXRcK2_1(.din(n15465), .dout(n15462));
    jdff dff_A_v0v4KUoW6_1(.din(n15468), .dout(n15465));
    jdff dff_A_lEOxaR872_1(.din(n15471), .dout(n15468));
    jdff dff_A_uFJdQoKg6_1(.din(n15474), .dout(n15471));
    jdff dff_A_hWrlshFl1_1(.din(n15477), .dout(n15474));
    jdff dff_A_7UY9nmdC8_1(.din(n15480), .dout(n15477));
    jdff dff_A_niaUuaPX1_1(.din(n15483), .dout(n15480));
    jdff dff_A_sKnW5gSz2_1(.din(n15486), .dout(n15483));
    jdff dff_A_qh4CeztD9_1(.din(n15489), .dout(n15486));
    jdff dff_A_ygC8iK3D9_1(.din(n15492), .dout(n15489));
    jdff dff_A_29YK8VA16_1(.din(n15595), .dout(n15492));
    jdff dff_A_FM70XG8Q0_2(.din(n15498), .dout(n15495));
    jdff dff_A_5HkoReu22_2(.din(n15501), .dout(n15498));
    jdff dff_A_8YKp4dCs0_2(.din(n15504), .dout(n15501));
    jdff dff_A_PdafN9kM7_2(.din(n15507), .dout(n15504));
    jdff dff_A_tSoASTp51_2(.din(n15510), .dout(n15507));
    jdff dff_A_l3SVPDTu0_2(.din(n15513), .dout(n15510));
    jdff dff_A_NCeIZyn30_2(.din(n15516), .dout(n15513));
    jdff dff_A_c33zlPMx0_2(.din(n15519), .dout(n15516));
    jdff dff_A_CKntm3vl8_2(.din(n15522), .dout(n15519));
    jdff dff_A_Pbl6qVni4_2(.din(n15595), .dout(n15522));
    jdff dff_A_4ukLVA8O8_1(.din(n15528), .dout(n15525));
    jdff dff_A_8FvYFgJ17_1(.din(n15531), .dout(n15528));
    jdff dff_A_cymLraMl8_1(.din(n15534), .dout(n15531));
    jdff dff_A_APp8NyV30_1(.din(n15537), .dout(n15534));
    jdff dff_A_vADtSfHk0_1(.din(n15540), .dout(n15537));
    jdff dff_A_iB6LAnTI1_1(.din(n15543), .dout(n15540));
    jdff dff_A_C60DUzXr7_1(.din(n15546), .dout(n15543));
    jdff dff_A_CP8EoBFH8_1(.din(n15549), .dout(n15546));
    jdff dff_A_L2OZaSFY0_1(.din(n15552), .dout(n15549));
    jdff dff_A_yp4yISs39_1(.din(n15555), .dout(n15552));
    jdff dff_A_ChpFXZM95_1(.din(n15595), .dout(n15555));
    jdff dff_A_cLxXia6N4_2(.din(n15561), .dout(n15558));
    jdff dff_A_BlkVTWEQ9_2(.din(n15564), .dout(n15561));
    jdff dff_A_WIcn31uy0_2(.din(n15567), .dout(n15564));
    jdff dff_A_6zlKOZOd4_2(.din(n15595), .dout(n15567));
    jdff dff_B_ScrxC0ex8_3(.din(n2188), .dout(n15571));
    jdff dff_B_bF9HSW5h6_3(.din(n15571), .dout(n15574));
    jdff dff_B_iV8XZhOK8_3(.din(n15574), .dout(n15577));
    jdff dff_B_IgwPsuVZ1_3(.din(n15577), .dout(n15580));
    jdff dff_B_pAHPjq7V4_3(.din(n15580), .dout(n15583));
    jdff dff_B_7mfdTIcv8_3(.din(n15583), .dout(n15586));
    jdff dff_B_bDR0fVtB4_3(.din(n15586), .dout(n15589));
    jdff dff_B_3WtelaWZ0_3(.din(n15589), .dout(n15592));
    jdff dff_B_1YMFOaP55_3(.din(n15592), .dout(n15595));
    jdff dff_A_uKSr5MXa6_0(.din(G4087), .dout(n15597));
    jdff dff_A_pPMSWfET9_1(.din(G4087), .dout(n15600));
    jdff dff_B_wjVMUX9z6_1(.din(n5564), .dout(n15604));
    jdff dff_B_F1BdJIRn7_1(.din(n15604), .dout(n15607));
    jdff dff_A_J7RpXy9j0_0(.din(n15612), .dout(n15609));
    jdff dff_A_B2b2QXRq5_0(.din(n15615), .dout(n15612));
    jdff dff_A_U73T2Cer5_0(.din(n15618), .dout(n15615));
    jdff dff_A_w39mU8Y99_0(.din(n15621), .dout(n15618));
    jdff dff_A_m15o0S1P9_0(.din(n15624), .dout(n15621));
    jdff dff_A_mcMP1zUM8_0(.din(n15627), .dout(n15624));
    jdff dff_A_zjECLO450_0(.din(n15630), .dout(n15627));
    jdff dff_A_aM0peksZ5_0(.din(n15633), .dout(n15630));
    jdff dff_A_FQZO09FO5_0(.din(n15636), .dout(n15633));
    jdff dff_A_Spd7vZn46_0(.din(n15639), .dout(n15636));
    jdff dff_A_bQitdwoY1_0(.din(n15642), .dout(n15639));
    jdff dff_A_oThGbyep6_0(.din(n15645), .dout(n15642));
    jdff dff_A_BZXl5qNo8_0(.din(n15648), .dout(n15645));
    jdff dff_A_DR3dhzZL6_0(.din(n15651), .dout(n15648));
    jdff dff_A_0X6f479c5_0(.din(n15654), .dout(n15651));
    jdff dff_A_AN4zE28N9_0(.din(n15657), .dout(n15654));
    jdff dff_A_M3BwlCt59_0(.din(n15660), .dout(n15657));
    jdff dff_A_RaZXe41y5_0(.din(n15663), .dout(n15660));
    jdff dff_A_ZTLypPDO1_0(.din(n15666), .dout(n15663));
    jdff dff_A_557w5x5b3_0(.din(n15669), .dout(n15666));
    jdff dff_A_70LyU2fl4_0(.din(n15672), .dout(n15669));
    jdff dff_A_ExNRHowj8_0(.din(n2178), .dout(n15672));
    jdff dff_A_9CG4UPxr9_1(.din(n15678), .dout(n15675));
    jdff dff_A_V1YRyjog0_1(.din(n15681), .dout(n15678));
    jdff dff_A_NCDTHPr95_1(.din(n15684), .dout(n15681));
    jdff dff_A_wIyHRV9x1_1(.din(n15687), .dout(n15684));
    jdff dff_A_zYyz2T3b6_1(.din(n15690), .dout(n15687));
    jdff dff_A_Jq3nLSms4_1(.din(n15693), .dout(n15690));
    jdff dff_A_SfRM7CcV4_1(.din(n15696), .dout(n15693));
    jdff dff_A_ouvJbN4a0_1(.din(n15699), .dout(n15696));
    jdff dff_A_F4a1JVaO5_1(.din(G4088), .dout(n15699));
    jdff dff_A_FjZ8h4rR6_1(.din(n15705), .dout(n15702));
    jdff dff_A_qxidpLW09_1(.din(G4087), .dout(n15705));
    jdff dff_A_EXoqS4CX2_2(.din(G4087), .dout(n15708));
    jdff dff_A_ZtjjC1cr6_1(.din(G4087), .dout(n15711));
    jdff dff_A_yQpYbEpp5_2(.din(G4087), .dout(n15714));
    jdff dff_A_stD9tdsP3_0(.din(n15720), .dout(n15717));
    jdff dff_A_GzQHRemz8_0(.din(n15723), .dout(n15720));
    jdff dff_A_q2xxL2809_0(.din(n15726), .dout(n15723));
    jdff dff_A_wjn5NGJL4_0(.din(n15729), .dout(n15726));
    jdff dff_A_3vHb5jwq0_0(.din(n15732), .dout(n15729));
    jdff dff_A_BxOZloTC5_0(.din(n15735), .dout(n15732));
    jdff dff_A_d2LAGOai2_0(.din(n15738), .dout(n15735));
    jdff dff_A_gKJA16UU5_0(.din(n15741), .dout(n15738));
    jdff dff_A_4c45Rt3G2_0(.din(n15744), .dout(n15741));
    jdff dff_A_7f1V6vuB5_0(.din(n15747), .dout(n15744));
    jdff dff_A_IdcioEF45_0(.din(n15750), .dout(n15747));
    jdff dff_A_NXCW0Peo0_0(.din(n15753), .dout(n15750));
    jdff dff_A_cKVgP91G6_0(.din(n15756), .dout(n15753));
    jdff dff_A_Rr3erOfF6_0(.din(n15759), .dout(n15756));
    jdff dff_A_I5pOKBT10_0(.din(n15762), .dout(n15759));
    jdff dff_A_rKht7d1D0_0(.din(n15765), .dout(n15762));
    jdff dff_A_EOyZ921T3_0(.din(n15768), .dout(n15765));
    jdff dff_A_eP5pG42G3_0(.din(n15771), .dout(n15768));
    jdff dff_A_m5UgHlOP8_0(.din(n15774), .dout(n15771));
    jdff dff_A_BIn5dbuA0_0(.din(n15777), .dout(n15774));
    jdff dff_A_ZrCBTGC77_0(.din(n15780), .dout(n15777));
    jdff dff_A_xo76DDLe0_0(.din(n15783), .dout(n15780));
    jdff dff_A_e2DMmeF93_0(.din(G4088), .dout(n15783));
    jdff dff_B_5VWJlEk10_1(.din(n5640), .dout(n15787));
    jdff dff_B_FKUbdl895_1(.din(n15787), .dout(n15790));
    jdff dff_B_GhtElLy78_1(.din(n15790), .dout(n15793));
    jdff dff_B_N1ppBTzP7_1(.din(n15793), .dout(n15796));
    jdff dff_B_qaJaVZEb7_1(.din(n15796), .dout(n15799));
    jdff dff_B_DPx4D44O9_1(.din(n15799), .dout(n15802));
    jdff dff_B_MIPrLEAQ4_1(.din(n15802), .dout(n15805));
    jdff dff_B_2p7NKM7G4_1(.din(n15805), .dout(n15808));
    jdff dff_B_W4eb44Fa9_1(.din(n15808), .dout(n15811));
    jdff dff_B_WueJfSvG9_1(.din(n15811), .dout(n15814));
    jdff dff_B_i02qVWdV5_1(.din(n15814), .dout(n15817));
    jdff dff_B_tz9ImYf91_1(.din(n15817), .dout(n15820));
    jdff dff_B_kFRza5023_1(.din(n15820), .dout(n15823));
    jdff dff_B_Jw1xMxJU9_1(.din(n15823), .dout(n15826));
    jdff dff_B_rGCXZjog7_1(.din(n15826), .dout(n15829));
    jdff dff_B_A6VkFRSM6_1(.din(n15829), .dout(n15832));
    jdff dff_B_7zLHV44n1_1(.din(n15832), .dout(n15835));
    jdff dff_B_vVmKJpte0_1(.din(n15835), .dout(n15838));
    jdff dff_B_JxXsnwWw9_1(.din(n15838), .dout(n15841));
    jdff dff_B_AvTLxa0U9_1(.din(n15841), .dout(n15844));
    jdff dff_B_0COEn1EF5_1(.din(n15844), .dout(n15847));
    jdff dff_B_JZhC67786_1(.din(n15847), .dout(n15850));
    jdff dff_B_4w8ijg4L1_1(.din(n5644), .dout(n15853));
    jdff dff_A_XHd2QwV55_1(.din(n15858), .dout(n15855));
    jdff dff_A_Ap4mMjKA8_1(.din(n15861), .dout(n15858));
    jdff dff_A_v0A9eA911_1(.din(n15864), .dout(n15861));
    jdff dff_A_ysOOM7QB4_1(.din(n15867), .dout(n15864));
    jdff dff_A_Ka0TaOuV2_1(.din(n15870), .dout(n15867));
    jdff dff_A_mmrxd1oL7_1(.din(n15873), .dout(n15870));
    jdff dff_A_6bNMblGB6_1(.din(n15876), .dout(n15873));
    jdff dff_A_xji6pgNy8_1(.din(n15879), .dout(n15876));
    jdff dff_A_ToTuOMhx6_1(.din(n15882), .dout(n15879));
    jdff dff_A_6ZjksA0e1_1(.din(n15885), .dout(n15882));
    jdff dff_A_bPTvEwAl5_1(.din(n15888), .dout(n15885));
    jdff dff_A_tUZ1kFg80_1(.din(n15891), .dout(n15888));
    jdff dff_A_AzxWRYBH5_1(.din(n15894), .dout(n15891));
    jdff dff_A_MADeFKk91_1(.din(n16000), .dout(n15894));
    jdff dff_A_HSeYYdKz2_2(.din(n15900), .dout(n15897));
    jdff dff_A_vIcfKhgF2_2(.din(n15903), .dout(n15900));
    jdff dff_A_lQAzILS92_2(.din(n15906), .dout(n15903));
    jdff dff_A_vcWsDHm01_2(.din(n15909), .dout(n15906));
    jdff dff_A_N3rKhFR06_2(.din(n15912), .dout(n15909));
    jdff dff_A_kkjVur1N4_2(.din(n15915), .dout(n15912));
    jdff dff_A_vpbSd4Xr2_2(.din(n15918), .dout(n15915));
    jdff dff_A_UbJhJIwu0_2(.din(n15921), .dout(n15918));
    jdff dff_A_5Lr90UL94_2(.din(n15924), .dout(n15921));
    jdff dff_A_cFnCmMlb6_2(.din(n16000), .dout(n15924));
    jdff dff_A_duCczTxM6_1(.din(n15930), .dout(n15927));
    jdff dff_A_vsdwndrL6_1(.din(n15933), .dout(n15930));
    jdff dff_A_DnrT2OXK6_1(.din(n15936), .dout(n15933));
    jdff dff_A_oUqq3q7g6_1(.din(n15939), .dout(n15936));
    jdff dff_A_BPJPEmzi0_1(.din(n15942), .dout(n15939));
    jdff dff_A_Ej2ttc3v6_1(.din(n15945), .dout(n15942));
    jdff dff_A_o4OMuCUz2_1(.din(n15948), .dout(n15945));
    jdff dff_A_YB9OgIea1_1(.din(n15951), .dout(n15948));
    jdff dff_A_3VItfUrT1_1(.din(n15954), .dout(n15951));
    jdff dff_A_A304rUl82_1(.din(n15957), .dout(n15954));
    jdff dff_A_DhjotKiY6_1(.din(n16000), .dout(n15957));
    jdff dff_A_BhU2XX7h7_2(.din(n15963), .dout(n15960));
    jdff dff_A_2niEqCLp7_2(.din(n15966), .dout(n15963));
    jdff dff_A_YhQiCBCf8_2(.din(n15969), .dout(n15966));
    jdff dff_A_8CdQoD6j4_2(.din(n15972), .dout(n15969));
    jdff dff_A_GJS3iESA2_2(.din(n16000), .dout(n15972));
    jdff dff_B_YU5aFbwY8_3(.din(n2394), .dout(n15976));
    jdff dff_B_mASZFfYi0_3(.din(n15976), .dout(n15979));
    jdff dff_B_X7VLNaWq3_3(.din(n15979), .dout(n15982));
    jdff dff_B_QCV7Orfh1_3(.din(n15982), .dout(n15985));
    jdff dff_B_v84117wn9_3(.din(n15985), .dout(n15988));
    jdff dff_B_KIsqCmnf9_3(.din(n15988), .dout(n15991));
    jdff dff_B_YNEIxzyE8_3(.din(n15991), .dout(n15994));
    jdff dff_B_QnYnZjV90_3(.din(n15994), .dout(n15997));
    jdff dff_B_LKKyFNdM0_3(.din(n15997), .dout(n16000));
    jdff dff_A_rTzxTR3f9_0(.din(n16005), .dout(n16002));
    jdff dff_A_ghHCOaPZ1_0(.din(G4090), .dout(n16005));
    jdff dff_A_y0stXhZv5_1(.din(G4090), .dout(n16008));
    jdff dff_B_6890W6Pk6_1(.din(n5628), .dout(n16012));
    jdff dff_B_zD5UW9OE9_1(.din(n16012), .dout(n16015));
    jdff dff_A_Md6L4ZLk1_0(.din(n16020), .dout(n16017));
    jdff dff_A_L1rL8Lnv3_0(.din(n16023), .dout(n16020));
    jdff dff_A_qRNKc1yt7_0(.din(n16026), .dout(n16023));
    jdff dff_A_ePbmOZq23_0(.din(n16029), .dout(n16026));
    jdff dff_A_h4WNevPM8_0(.din(n16032), .dout(n16029));
    jdff dff_A_4BdJor4m2_0(.din(n16035), .dout(n16032));
    jdff dff_A_AiDyksuY8_0(.din(n16038), .dout(n16035));
    jdff dff_A_LiFeRp1E3_0(.din(n16041), .dout(n16038));
    jdff dff_A_MccVLTGR2_0(.din(n16044), .dout(n16041));
    jdff dff_A_FOVAUchP1_0(.din(n16047), .dout(n16044));
    jdff dff_A_AMohUKfL5_0(.din(n16050), .dout(n16047));
    jdff dff_A_xy8G4voT8_0(.din(n16053), .dout(n16050));
    jdff dff_A_EOr0CDKt2_0(.din(n16056), .dout(n16053));
    jdff dff_A_cDeiVApS6_0(.din(n16059), .dout(n16056));
    jdff dff_A_7OK8rxKQ2_0(.din(n16062), .dout(n16059));
    jdff dff_A_8K67Gti73_0(.din(n16065), .dout(n16062));
    jdff dff_A_w9dg7Net7_0(.din(n16068), .dout(n16065));
    jdff dff_A_TEtlqzdT3_0(.din(n16071), .dout(n16068));
    jdff dff_A_8HZgfnTa5_0(.din(n16074), .dout(n16071));
    jdff dff_A_mwdF4tvc7_0(.din(n16077), .dout(n16074));
    jdff dff_A_hthhEKpR5_0(.din(n16080), .dout(n16077));
    jdff dff_A_gPRdKgN45_0(.din(n2387), .dout(n16080));
    jdff dff_A_wt8bNgyy7_1(.din(n16086), .dout(n16083));
    jdff dff_A_A6De25d65_1(.din(n16089), .dout(n16086));
    jdff dff_A_OdmbJE6u6_1(.din(n16092), .dout(n16089));
    jdff dff_A_2W0nE7DX9_1(.din(n16095), .dout(n16092));
    jdff dff_A_HwNHOzNl1_1(.din(n16098), .dout(n16095));
    jdff dff_A_VBKp2dHu3_1(.din(n16101), .dout(n16098));
    jdff dff_A_txW4Kzme7_1(.din(n16104), .dout(n16101));
    jdff dff_A_1xkcgrRy6_1(.din(n16107), .dout(n16104));
    jdff dff_A_y6gLe14R0_1(.din(G4089), .dout(n16107));
    jdff dff_B_YuQ5o83W9_2(.din(G64), .dout(n16111));
    jdff dff_A_rrKM09fd4_1(.din(n16116), .dout(n16113));
    jdff dff_A_a1NFrYxL3_1(.din(G4090), .dout(n16116));
    jdff dff_A_oHlGz0YR3_2(.din(G4090), .dout(n16119));
    jdff dff_A_98uwd9An2_1(.din(G4090), .dout(n16122));
    jdff dff_A_N5K4KyUj0_2(.din(G4090), .dout(n16125));
    jdff dff_A_rdeyPKAs0_0(.din(n16131), .dout(n16128));
    jdff dff_A_rJ4BELuO9_0(.din(n16134), .dout(n16131));
    jdff dff_A_QsjLx9Ce7_0(.din(n16137), .dout(n16134));
    jdff dff_A_C9GsvAJa7_0(.din(n16140), .dout(n16137));
    jdff dff_A_y1xvDWAF2_0(.din(n16143), .dout(n16140));
    jdff dff_A_tO0Qrx1f1_0(.din(n16146), .dout(n16143));
    jdff dff_A_IEu0Uf5u3_0(.din(n16149), .dout(n16146));
    jdff dff_A_oBHPoYYs8_0(.din(n16152), .dout(n16149));
    jdff dff_A_k35eJEDi1_0(.din(n16155), .dout(n16152));
    jdff dff_A_MsesAbzI5_0(.din(n16158), .dout(n16155));
    jdff dff_A_TAEROzuT5_0(.din(n16161), .dout(n16158));
    jdff dff_A_ATy3qVdy1_0(.din(n16164), .dout(n16161));
    jdff dff_A_oHE4udjl1_0(.din(n16167), .dout(n16164));
    jdff dff_A_tAkLuTeL3_0(.din(n16170), .dout(n16167));
    jdff dff_A_MFrG6Vnt9_0(.din(n16173), .dout(n16170));
    jdff dff_A_j6HF3K6N8_0(.din(n16176), .dout(n16173));
    jdff dff_A_bPPJTE1Z3_0(.din(n16179), .dout(n16176));
    jdff dff_A_jyR1jeXn2_0(.din(n16182), .dout(n16179));
    jdff dff_A_rfIPd6nx3_0(.din(n16185), .dout(n16182));
    jdff dff_A_RSZ9pChh2_0(.din(n16188), .dout(n16185));
    jdff dff_A_ie7Z40Gz9_0(.din(n16191), .dout(n16188));
    jdff dff_A_ZPALRbNc1_0(.din(n16194), .dout(n16191));
    jdff dff_A_M6dwhNZe0_0(.din(G4089), .dout(n16194));
    jdff dff_B_bMIbFn0F5_1(.din(n5673), .dout(n16198));
    jdff dff_B_Oa9qd6IH4_1(.din(n16198), .dout(n16201));
    jdff dff_B_wGu4CYYp9_1(.din(n16201), .dout(n16204));
    jdff dff_B_Ue4dzxzn0_1(.din(n16204), .dout(n16207));
    jdff dff_B_ELSlJ2Fh7_1(.din(n16207), .dout(n16210));
    jdff dff_B_TnFwnLhE0_1(.din(n16210), .dout(n16213));
    jdff dff_B_0Mqoad4x4_1(.din(n16213), .dout(n16216));
    jdff dff_B_ltrxup4S5_1(.din(n16216), .dout(n16219));
    jdff dff_B_5LAFverN7_1(.din(n16219), .dout(n16222));
    jdff dff_B_JCr0poLX2_1(.din(n16222), .dout(n16225));
    jdff dff_B_5G8zQwIv0_1(.din(n16225), .dout(n16228));
    jdff dff_B_fP0jmasL8_1(.din(n16228), .dout(n16231));
    jdff dff_B_AB3Z6gZY9_1(.din(n16231), .dout(n16234));
    jdff dff_B_N9p2ONu75_1(.din(n16234), .dout(n16237));
    jdff dff_B_6uQeOPUq7_1(.din(n16237), .dout(n16240));
    jdff dff_B_uW0c6eat7_1(.din(n16240), .dout(n16243));
    jdff dff_B_K7gGYNGh6_1(.din(n16243), .dout(n16246));
    jdff dff_B_e9N9hQB34_1(.din(n16246), .dout(n16249));
    jdff dff_B_yBPMgex56_1(.din(n16249), .dout(n16252));
    jdff dff_B_EJ1vIkfj9_1(.din(n16252), .dout(n16255));
    jdff dff_B_3Pnvo5Wy4_1(.din(n16255), .dout(n16258));
    jdff dff_B_yxl5bIgC1_1(.din(n16258), .dout(n16261));
    jdff dff_B_OFoLb81D1_1(.din(n16261), .dout(n16264));
    jdff dff_B_BtjNFnQ62_1(.din(n5683), .dout(n16267));
    jdff dff_B_7zbOjT482_1(.din(n16267), .dout(n16270));
    jdff dff_B_X3Q2TPw86_1(.din(n16270), .dout(n16273));
    jdff dff_B_VBQ2ByaR2_1(.din(n16273), .dout(n16276));
    jdff dff_B_HP4pVqIo7_1(.din(n16276), .dout(n16279));
    jdff dff_B_szQD7lG23_1(.din(n16279), .dout(n16282));
    jdff dff_B_Wk9oLYPq2_1(.din(n16282), .dout(n16285));
    jdff dff_B_J4crlOi21_1(.din(n16285), .dout(n16288));
    jdff dff_B_d289MB6R7_1(.din(n16288), .dout(n16291));
    jdff dff_B_9qFjxQSI4_1(.din(n16291), .dout(n16294));
    jdff dff_B_lFXW8lHy0_1(.din(n16294), .dout(n16297));
    jdff dff_B_3aozawya1_1(.din(n16297), .dout(n16300));
    jdff dff_B_35hDRlGt3_1(.din(n16300), .dout(n16303));
    jdff dff_B_g8DzMmqT5_1(.din(n16303), .dout(n16306));
    jdff dff_B_1V2d6Ptw3_1(.din(n16306), .dout(n16309));
    jdff dff_B_VaCCbFQW1_1(.din(n16309), .dout(n16312));
    jdff dff_B_3lYlaJqe7_1(.din(n16312), .dout(n16315));
    jdff dff_B_vErUsyA04_1(.din(n16315), .dout(n16318));
    jdff dff_B_v4T5gsVC4_1(.din(n16318), .dout(n16321));
    jdff dff_B_0kJnOtNr6_1(.din(n16321), .dout(n16324));
    jdff dff_B_2cHRsFbU8_1(.din(n16324), .dout(n16327));
    jdff dff_B_yScOK9ru2_1(.din(n5687), .dout(n16330));
    jdff dff_A_SlYv8LDR1_0(.din(n16335), .dout(n16332));
    jdff dff_A_ItebSVhY6_0(.din(n16338), .dout(n16335));
    jdff dff_A_MdmZpCRp5_0(.din(n16341), .dout(n16338));
    jdff dff_A_F3uKWVcV2_0(.din(n16344), .dout(n16341));
    jdff dff_A_qhnKv03l0_0(.din(n16347), .dout(n16344));
    jdff dff_A_jyFXtZNu1_0(.din(n16350), .dout(n16347));
    jdff dff_A_a3kbefkD9_0(.din(n16353), .dout(n16350));
    jdff dff_A_wDfwGPd80_0(.din(n16356), .dout(n16353));
    jdff dff_A_jqIEugti6_0(.din(n16359), .dout(n16356));
    jdff dff_A_Ioz0d5Nt4_0(.din(n16362), .dout(n16359));
    jdff dff_A_wYl1bAxT8_0(.din(n16365), .dout(n16362));
    jdff dff_A_yo3MvZQ20_0(.din(n16368), .dout(n16365));
    jdff dff_A_CA7cmmFD8_0(.din(n16371), .dout(n16368));
    jdff dff_A_jAKgpXcQ3_0(.din(n16374), .dout(n16371));
    jdff dff_A_GY8z1wY53_0(.din(n2921), .dout(n16374));
    jdff dff_A_hBs0JYMO5_1(.din(n16380), .dout(n16377));
    jdff dff_A_E00msF9S8_1(.din(n16383), .dout(n16380));
    jdff dff_A_KBrCNoyH2_1(.din(n16386), .dout(n16383));
    jdff dff_A_hQt0O5c47_1(.din(n16389), .dout(n16386));
    jdff dff_A_s4HPvbzB5_1(.din(n16392), .dout(n16389));
    jdff dff_A_9XR28cZQ0_1(.din(n16395), .dout(n16392));
    jdff dff_A_SaluuUvc8_1(.din(n16398), .dout(n16395));
    jdff dff_A_IBgY35Ba8_1(.din(n16401), .dout(n16398));
    jdff dff_A_LcIc8VQ40_1(.din(n16404), .dout(n16401));
    jdff dff_A_0fxBTHVS6_1(.din(n2921), .dout(n16404));
    jdff dff_A_Sx4BI8977_1(.din(n16410), .dout(n16407));
    jdff dff_A_BgW4wWCA1_1(.din(n16413), .dout(n16410));
    jdff dff_A_zbtyXcT68_1(.din(n16416), .dout(n16413));
    jdff dff_A_RXC5pQLZ0_1(.din(n16419), .dout(n16416));
    jdff dff_A_6q7gu6kZ5_1(.din(n16422), .dout(n16419));
    jdff dff_A_PvgqQlK40_1(.din(n16425), .dout(n16422));
    jdff dff_A_krANA6Z87_1(.din(n16428), .dout(n16425));
    jdff dff_A_1naFaLhF2_1(.din(n16431), .dout(n16428));
    jdff dff_A_Ojn0kkYc3_1(.din(n16434), .dout(n16431));
    jdff dff_A_LJnRnScN6_1(.din(n16437), .dout(n16434));
    jdff dff_A_oMXIdcBD7_1(.din(n16440), .dout(n16437));
    jdff dff_A_DRrznnA01_1(.din(n16443), .dout(n16440));
    jdff dff_A_X0KzkqqW8_1(.din(n16446), .dout(n16443));
    jdff dff_A_q488RTdU3_1(.din(n16449), .dout(n16446));
    jdff dff_A_pC6vtcTT4_1(.din(n16452), .dout(n16449));
    jdff dff_A_oErH0m2e9_1(.din(n16455), .dout(n16452));
    jdff dff_A_SmdYjCkC2_1(.din(n16458), .dout(n16455));
    jdff dff_A_wv8LgdWo5_1(.din(n16461), .dout(n16458));
    jdff dff_A_vfOOW9eV1_1(.din(n16464), .dout(n16461));
    jdff dff_A_OmbFbeiy7_1(.din(n16467), .dout(n16464));
    jdff dff_A_LPoxAlm50_1(.din(n2921), .dout(n16467));
    jdff dff_A_1apXy0ad4_2(.din(n16473), .dout(n16470));
    jdff dff_A_SjCjHrU97_2(.din(n16476), .dout(n16473));
    jdff dff_A_y2R6h7587_2(.din(n16479), .dout(n16476));
    jdff dff_A_Ra9P4r6X0_2(.din(n16482), .dout(n16479));
    jdff dff_A_XXSDnZKZ6_2(.din(n16485), .dout(n16482));
    jdff dff_A_7tYfKjwv0_2(.din(n16488), .dout(n16485));
    jdff dff_A_fwTHRFFT7_2(.din(n16491), .dout(n16488));
    jdff dff_A_kes8BGOy5_2(.din(n16494), .dout(n16491));
    jdff dff_A_cIKV6sB89_2(.din(n16497), .dout(n16494));
    jdff dff_A_tBOTIIWJ7_2(.din(n16500), .dout(n16497));
    jdff dff_A_uO7t2O6z3_2(.din(n16503), .dout(n16500));
    jdff dff_A_f4Zs8oBC4_2(.din(n16506), .dout(n16503));
    jdff dff_A_Whe0g9Av0_2(.din(n16509), .dout(n16506));
    jdff dff_A_2B1qupzO7_2(.din(n16512), .dout(n16509));
    jdff dff_A_jG06aDOL0_2(.din(n16515), .dout(n16512));
    jdff dff_A_NaB2w87d7_2(.din(n16518), .dout(n16515));
    jdff dff_A_Twvw7lxj4_2(.din(n16521), .dout(n16518));
    jdff dff_A_oewqjaCp0_2(.din(n16524), .dout(n16521));
    jdff dff_A_Lt74J5M05_2(.din(n16527), .dout(n16524));
    jdff dff_A_bFcptGNJ2_2(.din(n2921), .dout(n16527));
    jdff dff_A_p4nLFl8q3_1(.din(n16533), .dout(n16530));
    jdff dff_A_EYrLqPqr0_1(.din(n16536), .dout(n16533));
    jdff dff_A_mBvmh2bY5_1(.din(n16539), .dout(n16536));
    jdff dff_A_VRP4Ngk05_1(.din(n16542), .dout(n16539));
    jdff dff_A_X82o1FL83_1(.din(n16545), .dout(n16542));
    jdff dff_A_0lDIfkg95_1(.din(n16548), .dout(n16545));
    jdff dff_A_IzmYZUuV3_1(.din(n16551), .dout(n16548));
    jdff dff_A_VGJA1fJn7_1(.din(n16554), .dout(n16551));
    jdff dff_A_LMANtSHB6_1(.din(n16557), .dout(n16554));
    jdff dff_A_ahxEezkt2_1(.din(n16560), .dout(n16557));
    jdff dff_A_x6JB4o569_1(.din(n16563), .dout(n16560));
    jdff dff_A_2QQSaOSQ2_1(.din(n16566), .dout(n16563));
    jdff dff_A_AZzYQT3o6_1(.din(n16569), .dout(n16566));
    jdff dff_A_vp6kULU05_1(.din(n16572), .dout(n16569));
    jdff dff_A_MJtMi19x2_1(.din(n16575), .dout(n16572));
    jdff dff_A_67K9j7t85_1(.din(n16578), .dout(n16575));
    jdff dff_A_fFSRRVgn1_1(.din(n16581), .dout(n16578));
    jdff dff_A_KDQYG55A6_1(.din(n2921), .dout(n16581));
    jdff dff_A_oLysiJcs3_2(.din(n16587), .dout(n16584));
    jdff dff_A_ggRoZm195_2(.din(n16590), .dout(n16587));
    jdff dff_A_b0G6MoTR1_2(.din(n16593), .dout(n16590));
    jdff dff_A_HIL9ujgO0_2(.din(n16596), .dout(n16593));
    jdff dff_A_6SxZoqee7_2(.din(n16599), .dout(n16596));
    jdff dff_A_NxmArqPE9_2(.din(n16602), .dout(n16599));
    jdff dff_A_FD6LLLM71_2(.din(n16605), .dout(n16602));
    jdff dff_A_K6hrhoON0_2(.din(n16608), .dout(n16605));
    jdff dff_A_1RU6fnuX6_2(.din(n16611), .dout(n16608));
    jdff dff_A_zpurIaVN1_2(.din(n16614), .dout(n16611));
    jdff dff_A_HLISzOAQ6_2(.din(n2921), .dout(n16614));
    jdff dff_A_oQ6hWZ8K6_1(.din(G1690), .dout(n16617));
    jdff dff_A_ZqQ5dgBf9_1(.din(n16623), .dout(n16620));
    jdff dff_A_BCD8u8gK8_1(.din(n16626), .dout(n16623));
    jdff dff_A_g8SwvjE69_1(.din(n16629), .dout(n16626));
    jdff dff_A_L21lRDsT2_1(.din(n16632), .dout(n16629));
    jdff dff_A_mjSB2XIM0_1(.din(n16635), .dout(n16632));
    jdff dff_A_Z1j81ptQ7_1(.din(n16638), .dout(n16635));
    jdff dff_A_2aaxuw399_1(.din(n16641), .dout(n16638));
    jdff dff_A_jMxfTBlk9_1(.din(n16644), .dout(n16641));
    jdff dff_A_poynQU1Y6_1(.din(n16647), .dout(n16644));
    jdff dff_A_v8Bg2hU68_1(.din(n16650), .dout(n16647));
    jdff dff_A_4U0l04jV0_1(.din(n16653), .dout(n16650));
    jdff dff_A_u4DWv6Lg0_1(.din(n16656), .dout(n16653));
    jdff dff_A_eIXvyG0r8_1(.din(n16659), .dout(n16656));
    jdff dff_A_5RWirk279_1(.din(n16662), .dout(n16659));
    jdff dff_A_yECbOnJk5_1(.din(n16665), .dout(n16662));
    jdff dff_A_c2vrPWTn6_1(.din(n16668), .dout(n16665));
    jdff dff_A_odjQJDVI1_1(.din(n16671), .dout(n16668));
    jdff dff_A_otNrD9H20_1(.din(n16674), .dout(n16671));
    jdff dff_A_YA7kGA5z9_1(.din(n16677), .dout(n16674));
    jdff dff_A_AitZwGyh9_1(.din(n16680), .dout(n16677));
    jdff dff_A_2UrOsUSd1_1(.din(n16683), .dout(n16680));
    jdff dff_A_hgNgdS730_1(.din(n16686), .dout(n16683));
    jdff dff_A_8q1v2Fau8_1(.din(G1690), .dout(n16686));
    jdff dff_A_VwzzJvf65_0(.din(n16692), .dout(n16689));
    jdff dff_A_ShNaac751_0(.din(n16695), .dout(n16692));
    jdff dff_A_5Oz4lCsW3_0(.din(n16698), .dout(n16695));
    jdff dff_A_ESwHyVEX2_0(.din(n16701), .dout(n16698));
    jdff dff_A_ji7vJUdB3_0(.din(n16704), .dout(n16701));
    jdff dff_A_CS8RqFnI3_0(.din(n16707), .dout(n16704));
    jdff dff_A_pappRIuy5_0(.din(n16710), .dout(n16707));
    jdff dff_A_E009sSDJ5_0(.din(n16713), .dout(n16710));
    jdff dff_A_DjEPVuot6_0(.din(G1689), .dout(n16713));
    jdff dff_A_63qojU8U2_2(.din(n16719), .dout(n16716));
    jdff dff_A_RfNOAa5D4_2(.din(n16722), .dout(n16719));
    jdff dff_A_iZPFkH8r6_2(.din(n16725), .dout(n16722));
    jdff dff_A_S0IfHSAp0_2(.din(n16728), .dout(n16725));
    jdff dff_A_Nq2xCbnW4_2(.din(n16731), .dout(n16728));
    jdff dff_A_crbYARKb0_2(.din(n16734), .dout(n16731));
    jdff dff_A_FgkZB9Mw4_2(.din(n16737), .dout(n16734));
    jdff dff_A_vQ3mENBJ9_2(.din(n16740), .dout(n16737));
    jdff dff_A_s85UEDSu3_2(.din(n16743), .dout(n16740));
    jdff dff_A_ibqOQKJ08_2(.din(n16746), .dout(n16743));
    jdff dff_A_5jt12NCG6_2(.din(n16749), .dout(n16746));
    jdff dff_A_VOUGfFPN2_2(.din(n16752), .dout(n16749));
    jdff dff_A_KbnJfHre1_2(.din(n16755), .dout(n16752));
    jdff dff_A_kApJddP89_2(.din(n16758), .dout(n16755));
    jdff dff_A_LIRcmzzV4_2(.din(n16761), .dout(n16758));
    jdff dff_A_DCfos2bf9_2(.din(n16764), .dout(n16761));
    jdff dff_A_10iNWcyt9_2(.din(n16767), .dout(n16764));
    jdff dff_A_iWZg5kyo0_2(.din(n16770), .dout(n16767));
    jdff dff_A_DKhhC6jr6_2(.din(n16773), .dout(n16770));
    jdff dff_A_8Bhrdh8W6_2(.din(n16776), .dout(n16773));
    jdff dff_A_X8tib3Xx3_2(.din(n16779), .dout(n16776));
    jdff dff_A_V9AeNPX94_2(.din(G1689), .dout(n16779));
    jdff dff_A_773q4Ajn8_1(.din(n16785), .dout(n16782));
    jdff dff_A_c8B6M1fH1_1(.din(n16788), .dout(n16785));
    jdff dff_A_QlWRPz4U7_1(.din(n16791), .dout(n16788));
    jdff dff_A_nnpthrqL4_1(.din(n16794), .dout(n16791));
    jdff dff_A_wPmKhg8A0_1(.din(n16797), .dout(n16794));
    jdff dff_A_cwOmZkHW5_1(.din(n16800), .dout(n16797));
    jdff dff_A_M4Db9nyY5_1(.din(n16803), .dout(n16800));
    jdff dff_A_FJJYCpmb3_1(.din(n16806), .dout(n16803));
    jdff dff_A_C8UCi4yX7_1(.din(n16809), .dout(n16806));
    jdff dff_A_eH6uomXR6_1(.din(n16812), .dout(n16809));
    jdff dff_A_zfQgTGRS8_1(.din(n16815), .dout(n16812));
    jdff dff_A_GVWeV97E2_1(.din(n16818), .dout(n16815));
    jdff dff_A_OUTm0v0B0_1(.din(n16821), .dout(n16818));
    jdff dff_A_F960wYkX9_1(.din(n16824), .dout(n16821));
    jdff dff_A_JCCE42rm0_1(.din(n16827), .dout(n16824));
    jdff dff_A_fxVNohek0_1(.din(n16830), .dout(n16827));
    jdff dff_A_rrl7vplS7_1(.din(n16833), .dout(n16830));
    jdff dff_A_gawc5Su77_1(.din(n16836), .dout(n16833));
    jdff dff_A_TRFWSf9o9_1(.din(G1689), .dout(n16836));
    jdff dff_A_2UEpnK4m7_2(.din(n16842), .dout(n16839));
    jdff dff_A_acpypHIp4_2(.din(n16845), .dout(n16842));
    jdff dff_A_3ensXNEH3_2(.din(n16848), .dout(n16845));
    jdff dff_A_9GgifZZj0_2(.din(n16851), .dout(n16848));
    jdff dff_A_SLN9LdOC7_2(.din(n16854), .dout(n16851));
    jdff dff_A_EuADFi455_2(.din(n16857), .dout(n16854));
    jdff dff_A_taIc74Ms2_2(.din(n16860), .dout(n16857));
    jdff dff_A_pYmkRsUp5_2(.din(n16863), .dout(n16860));
    jdff dff_A_BJZnq2nh9_2(.din(n16866), .dout(n16863));
    jdff dff_A_GwsTqavO7_2(.din(n16869), .dout(n16866));
    jdff dff_A_wl56k2at9_2(.din(n16872), .dout(n16869));
    jdff dff_A_dqC8Jl5g8_2(.din(n16875), .dout(n16872));
    jdff dff_A_qhYXJhut8_2(.din(G1689), .dout(n16875));
    jdff dff_B_fappLODQ3_1(.din(n5718), .dout(n16879));
    jdff dff_B_K1eSItKk0_1(.din(n16879), .dout(n16882));
    jdff dff_B_f4UNuX4U5_1(.din(n16882), .dout(n16885));
    jdff dff_B_Xe6OwQUV0_1(.din(n16885), .dout(n16888));
    jdff dff_B_vltlLjBs2_1(.din(n16888), .dout(n16891));
    jdff dff_B_ZNPbb3Je8_1(.din(n16891), .dout(n16894));
    jdff dff_B_LigNWl0D7_1(.din(n16894), .dout(n16897));
    jdff dff_B_JxbLPvAR2_1(.din(n16897), .dout(n16900));
    jdff dff_B_N8ynxXMk0_1(.din(n16900), .dout(n16903));
    jdff dff_B_84PIClfp7_1(.din(n16903), .dout(n16906));
    jdff dff_B_G8uzX2zx0_1(.din(n16906), .dout(n16909));
    jdff dff_B_a1GkaZ6l0_1(.din(n16909), .dout(n16912));
    jdff dff_B_jBZI8hw18_1(.din(n16912), .dout(n16915));
    jdff dff_B_PqLUO8oi4_1(.din(n16915), .dout(n16918));
    jdff dff_B_3ubxHMpQ4_1(.din(n16918), .dout(n16921));
    jdff dff_B_lkcI4hR56_1(.din(n16921), .dout(n16924));
    jdff dff_B_OYdWE7k76_1(.din(n16924), .dout(n16927));
    jdff dff_B_A84Spr3i9_1(.din(n16927), .dout(n16930));
    jdff dff_B_dG9LJPdV7_1(.din(n16930), .dout(n16933));
    jdff dff_B_qKANdGMn4_1(.din(n16933), .dout(n16936));
    jdff dff_B_x3SmIgxL6_1(.din(n16936), .dout(n16939));
    jdff dff_B_Zp839Tqa8_1(.din(n16939), .dout(n16942));
    jdff dff_B_4pl9l5DJ3_1(.din(n16942), .dout(n16945));
    jdff dff_B_7KxXvuiq5_1(.din(n5725), .dout(n16948));
    jdff dff_B_VwMv84VU3_1(.din(n16948), .dout(n16951));
    jdff dff_B_AztD1pwj1_1(.din(n16951), .dout(n16954));
    jdff dff_B_LyzQh7MP8_1(.din(n16954), .dout(n16957));
    jdff dff_B_dJFA7P208_1(.din(n16957), .dout(n16960));
    jdff dff_B_Fq43BFwN3_1(.din(n16960), .dout(n16963));
    jdff dff_B_G0BVtXRn7_1(.din(n16963), .dout(n16966));
    jdff dff_B_kn63FJ2r7_1(.din(n16966), .dout(n16969));
    jdff dff_B_5Zutcn3n0_1(.din(n16969), .dout(n16972));
    jdff dff_B_TAinSHb54_1(.din(n16972), .dout(n16975));
    jdff dff_B_VLJu7GQG7_1(.din(n16975), .dout(n16978));
    jdff dff_B_GNgU3cM99_1(.din(n16978), .dout(n16981));
    jdff dff_B_kIOcZ6FJ0_1(.din(n16981), .dout(n16984));
    jdff dff_B_3mwH3La20_1(.din(n16984), .dout(n16987));
    jdff dff_B_pWpPGTZd5_1(.din(n16987), .dout(n16990));
    jdff dff_B_tT7GL0eE8_1(.din(n16990), .dout(n16993));
    jdff dff_B_vevqLO3x7_1(.din(n16993), .dout(n16996));
    jdff dff_B_vQ9pZ3jq7_1(.din(n16996), .dout(n16999));
    jdff dff_B_aOWQD9044_1(.din(n16999), .dout(n17002));
    jdff dff_B_r5AAnhzs6_1(.din(n17002), .dout(n17005));
    jdff dff_B_lPnA7KxI1_1(.din(n17005), .dout(n17008));
    jdff dff_B_TvwtaERu1_1(.din(n5729), .dout(n17011));
    jdff dff_B_uMayVPtM2_0(.din(n5601), .dout(n17014));
    jdff dff_B_YehyMLQ18_0(.din(n17014), .dout(n17017));
    jdff dff_B_oyrNO1rC6_0(.din(n17017), .dout(n17020));
    jdff dff_B_Pzqkmj7s0_0(.din(n17020), .dout(n17023));
    jdff dff_B_l9nXCu7R0_0(.din(n17023), .dout(n17026));
    jdff dff_B_VuH0LG3Y0_0(.din(n17026), .dout(n17029));
    jdff dff_B_7CLkLhNS4_0(.din(n17029), .dout(n17032));
    jdff dff_B_dZfUUkFQ9_0(.din(n17032), .dout(n17035));
    jdff dff_B_R0ph8LWv6_0(.din(n17035), .dout(n17038));
    jdff dff_B_ihydbqsS0_0(.din(n17038), .dout(n17041));
    jdff dff_B_1uf5h5F70_0(.din(n17041), .dout(n17044));
    jdff dff_B_d88tFYTL8_0(.din(n17044), .dout(n17047));
    jdff dff_B_t3YGfFxZ4_0(.din(n17047), .dout(n17050));
    jdff dff_B_KLvwqxyX5_0(.din(n17050), .dout(n17053));
    jdff dff_B_seZyezCh5_0(.din(n17053), .dout(n17056));
    jdff dff_B_dJcJZI5n5_0(.din(n17056), .dout(n17059));
    jdff dff_B_wpWc3Yfc5_0(.din(n17059), .dout(n17062));
    jdff dff_B_AR7NSALd2_0(.din(n17062), .dout(n17065));
    jdff dff_B_tshotWrx4_0(.din(n17065), .dout(n17068));
    jdff dff_B_SX1hBGvL9_0(.din(n4908), .dout(n17071));
    jdff dff_B_Vu0RJXKf9_0(.din(n17071), .dout(n17074));
    jdff dff_B_n5BF50uh8_0(.din(n17074), .dout(n17077));
    jdff dff_B_Az16hyfc7_0(.din(n17077), .dout(n17080));
    jdff dff_B_HzbJxaAG6_0(.din(n17080), .dout(n17083));
    jdff dff_B_wexuEVra7_0(.din(n17083), .dout(n17086));
    jdff dff_B_oCa9GmqI7_0(.din(n17086), .dout(n17089));
    jdff dff_B_Xefk6Yl04_0(.din(n17089), .dout(n17092));
    jdff dff_B_LnFfZrMQ4_0(.din(n17092), .dout(n17095));
    jdff dff_B_vCCTPlxH9_1(.din(n4889), .dout(n17098));
    jdff dff_B_KY4oClPQ5_1(.din(n713), .dout(n17101));
    jdff dff_B_HKApNhrR4_1(.din(n17101), .dout(n17104));
    jdff dff_A_ScLRp0dH0_0(.din(G308), .dout(n17106));
    jdff dff_B_IuHkOkDX2_1(.din(n665), .dout(n17110));
    jdff dff_B_yyfaiPDj6_1(.din(n17110), .dout(n17113));
    jdff dff_A_ZpN0xOKU4_1(.din(n770), .dout(n17115));
    jdff dff_B_8Xf7QnmY4_0(.din(n4877), .dout(n17119));
    jdff dff_A_S8jCp1lV4_0(.din(G361), .dout(n17121));
    jdff dff_B_4uGaUG2h6_1(.din(n4845), .dout(n17125));
    jdff dff_A_JMj54jpY1_0(.din(n17131), .dout(n17127));
    jdff dff_B_SB3eUVwo7_2(.din(n802), .dout(n17131));
    jdff dff_A_bqOqBG597_0(.din(n17136), .dout(n17133));
    jdff dff_A_0rgalY9k1_0(.din(n17139), .dout(n17136));
    jdff dff_A_PXTYXeMl1_0(.din(G503), .dout(n17139));
    jdff dff_B_EY5P9kkJ0_1(.din(n4829), .dout(n17143));
    jdff dff_B_xQ7tHhqd7_1(.din(n4789), .dout(n17146));
    jdff dff_B_3bgIAedx2_1(.din(n17146), .dout(n17149));
    jdff dff_A_F6B7u8qa1_1(.din(G341), .dout(n17151));
    jdff dff_B_TnwyGcai3_1(.din(n4753), .dout(n17155));
    jdff dff_B_Ifi5KaPP0_1(.din(n17155), .dout(n17158));
    jdff dff_A_ngYc9BaC7_1(.din(G351), .dout(n17160));
    jdff dff_B_z7gTYVop1_1(.din(n4717), .dout(n17164));
    jdff dff_A_V7FGggCU2_0(.din(n17169), .dout(n17166));
    jdff dff_A_yTmRByLd0_0(.din(n17172), .dout(n17169));
    jdff dff_A_aUEeXtDh7_0(.din(n19686), .dout(n17172));
    jdff dff_A_ZGbPL6sO7_1(.din(n17178), .dout(n17175));
    jdff dff_A_xCDea2wl3_1(.din(n17181), .dout(n17178));
    jdff dff_A_gJgdEIrO5_1(.din(n17184), .dout(n17181));
    jdff dff_A_QtdHhHKE0_1(.din(n17187), .dout(n17184));
    jdff dff_A_8mDJimVz1_1(.din(n17190), .dout(n17187));
    jdff dff_A_FCBxGdyh3_1(.din(n17193), .dout(n17190));
    jdff dff_A_h9R3Tg6B4_1(.din(n17196), .dout(n17193));
    jdff dff_A_Bn8s0z5C4_1(.din(n17199), .dout(n17196));
    jdff dff_A_qWGh3QJT3_1(.din(n17202), .dout(n17199));
    jdff dff_A_acbRl9gy2_1(.din(n17205), .dout(n17202));
    jdff dff_A_GpYsJDvJ6_1(.din(n17208), .dout(n17205));
    jdff dff_A_Y5kv7rC74_1(.din(n19686), .dout(n17208));
    jdff dff_B_99f1ywRJ4_0(.din(n4713), .dout(n17212));
    jdff dff_A_ZotBMQ0D5_0(.din(n17217), .dout(n17214));
    jdff dff_A_TmQHv6xl0_0(.din(n4710), .dout(n17217));
    jdff dff_B_KKXQIs3M6_0(.din(n4706), .dout(n17221));
    jdff dff_B_03kMr17E1_0(.din(n17221), .dout(n17224));
    jdff dff_B_c3XXmCf30_0(.din(n17224), .dout(n17227));
    jdff dff_B_pC6Oo3Vw3_1(.din(n4698), .dout(n17230));
    jdff dff_B_BwKl9oSn1_1(.din(n17230), .dout(n17233));
    jdff dff_B_HMWdFj7t1_1(.din(n17233), .dout(n17236));
    jdff dff_A_jOpFjveP9_0(.din(n17241), .dout(n17238));
    jdff dff_A_0WBcNEnh6_0(.din(n17244), .dout(n17241));
    jdff dff_A_Colzfz4w2_0(.din(n17247), .dout(n17244));
    jdff dff_A_2gaaYJ2z9_0(.din(n17250), .dout(n17247));
    jdff dff_A_pKK52SXc3_0(.din(n17253), .dout(n17250));
    jdff dff_A_zCWqs08e9_0(.din(n17256), .dout(n17253));
    jdff dff_A_ZDmExVea5_0(.din(n17259), .dout(n17256));
    jdff dff_A_Nh5iaij37_0(.din(n2051), .dout(n17259));
    jdff dff_B_gkOm9f2C8_1(.din(n4662), .dout(n17263));
    jdff dff_B_X7h3zKJR7_1(.din(n4670), .dout(n17266));
    jdff dff_B_HFXHnHTq0_0(.din(n4654), .dout(n17269));
    jdff dff_B_YmCA8NpP5_0(.din(n4650), .dout(n17272));
    jdff dff_A_fLKCUw2Z1_0(.din(n4624), .dout(n17274));
    jdff dff_B_CGHTI8A53_1(.din(n4616), .dout(n17278));
    jdff dff_A_qr3O2Jyf8_2(.din(n17283), .dout(n17280));
    jdff dff_A_3lMUSRFd5_2(.din(n1583), .dout(n17283));
    jdff dff_A_pp4HwyNl2_0(.din(n1579), .dout(n17286));
    jdff dff_A_hISlCyLZ4_0(.din(n1575), .dout(n17289));
    jdff dff_A_PUUWdHUJ7_0(.din(n17295), .dout(n17292));
    jdff dff_A_Jhn4XrRk4_0(.din(n17305), .dout(n17295));
    jdff dff_A_TizUnkPX5_1(.din(n17305), .dout(n17298));
    jdff dff_B_8fAdz1ZW7_3(.din(n1517), .dout(n17302));
    jdff dff_B_XUuxerAk5_3(.din(n17302), .dout(n17305));
    jdff dff_A_SYi6c45J6_1(.din(n17310), .dout(n17307));
    jdff dff_A_3MEM3U4V7_1(.din(n17313), .dout(n17310));
    jdff dff_A_3umru07q0_1(.din(n17316), .dout(n17313));
    jdff dff_A_NHz2SRfK7_1(.din(n1501), .dout(n17316));
    jdff dff_A_qHr140EL7_1(.din(n17322), .dout(n17319));
    jdff dff_A_GwQxQH0o0_1(.din(n1501), .dout(n17322));
    jdff dff_A_pu0aBU7w3_2(.din(n17328), .dout(n17325));
    jdff dff_A_B2AbRm9C6_2(.din(n17331), .dout(n17328));
    jdff dff_A_RzH3MoT43_2(.din(n17334), .dout(n17331));
    jdff dff_A_UnQODbXq5_2(.din(n17337), .dout(n17334));
    jdff dff_A_QAGcJSPV5_2(.din(n17340), .dout(n17337));
    jdff dff_A_fdnYTmS70_2(.din(n17343), .dout(n17340));
    jdff dff_A_ioamGLlq1_2(.din(n1501), .dout(n17343));
    jdff dff_A_4Q6uc5GK7_1(.din(n17349), .dout(n17346));
    jdff dff_A_dsFZ2h5H1_1(.din(n17352), .dout(n17349));
    jdff dff_A_JL4ZPdIW2_1(.din(n17355), .dout(n17352));
    jdff dff_A_NFvJFWBi9_1(.din(n17358), .dout(n17355));
    jdff dff_A_2ddUJsYP3_1(.din(n17361), .dout(n17358));
    jdff dff_A_zHayOKWN5_1(.din(n1493), .dout(n17361));
    jdff dff_A_3tylgieY3_2(.din(n17367), .dout(n17364));
    jdff dff_A_qBVbiEbx0_2(.din(n17370), .dout(n17367));
    jdff dff_A_XOM3sFug4_2(.din(n1493), .dout(n17370));
    jdff dff_A_5WLf0liM1_0(.din(n4610), .dout(n17373));
    jdff dff_B_T4kygeEA9_1(.din(n4558), .dout(n17377));
    jdff dff_A_O4Bg95WV8_0(.din(n4598), .dout(n17379));
    jdff dff_B_1KSxEyng2_1(.din(n4583), .dout(n17383));
    jdff dff_B_xjS2fJOz2_1(.din(n17383), .dout(n17386));
    jdff dff_B_g9698oLR9_1(.din(n17386), .dout(n17389));
    jdff dff_B_CXq2RJea6_1(.din(n4586), .dout(n17392));
    jdff dff_B_fuURMbT48_1(.din(n17392), .dout(n17395));
    jdff dff_A_8KmR0YJP9_2(.din(n17400), .dout(n17397));
    jdff dff_A_snwGPB9Z3_2(.din(n17403), .dout(n17400));
    jdff dff_A_E2gla9Im8_2(.din(n17406), .dout(n17403));
    jdff dff_A_lvIaQO0g4_2(.din(n17409), .dout(n17406));
    jdff dff_A_8dtaMtdk8_2(.din(n17412), .dout(n17409));
    jdff dff_A_L4yrxRrg8_2(.din(n1656), .dout(n17412));
    jdff dff_A_PLnNkKAR6_2(.din(n17418), .dout(n17415));
    jdff dff_A_tPGViu0P0_2(.din(n17421), .dout(n17418));
    jdff dff_A_LiZCO5hy1_2(.din(n17424), .dout(n17421));
    jdff dff_A_38fXQmRj4_2(.din(n17427), .dout(n17424));
    jdff dff_A_JJd7wOE12_2(.din(n17430), .dout(n17427));
    jdff dff_A_NSJ5nVXs1_2(.din(n17433), .dout(n17430));
    jdff dff_A_slkS1ByX2_2(.din(n17436), .dout(n17433));
    jdff dff_A_N3Gq0osR5_2(.din(n17439), .dout(n17436));
    jdff dff_A_68PoRUC35_2(.din(n2160), .dout(n17439));
    jdff dff_A_wo7kR2uM2_1(.din(n17445), .dout(n17442));
    jdff dff_A_yLioJ1nj9_1(.din(n17448), .dout(n17445));
    jdff dff_A_lBhsoe5B3_1(.din(n17451), .dout(n17448));
    jdff dff_A_QNWnC9vh2_1(.din(n17454), .dout(n17451));
    jdff dff_A_xVD02jHt7_1(.din(n17457), .dout(n17454));
    jdff dff_A_kgVQSWxH0_1(.din(n17460), .dout(n17457));
    jdff dff_A_0fIJiKcG7_1(.din(n17463), .dout(n17460));
    jdff dff_A_jtqU0hGe6_1(.din(n17466), .dout(n17463));
    jdff dff_A_54lJdxHT6_1(.din(n17469), .dout(n17466));
    jdff dff_A_4MuFKhJy2_1(.din(n2153), .dout(n17469));
    jdff dff_B_9CdaUsTE7_1(.din(n4564), .dout(n17473));
    jdff dff_B_IcLk55ca2_1(.din(n17473), .dout(n17476));
    jdff dff_B_2Y962Pvs2_1(.din(n17476), .dout(n17479));
    jdff dff_B_Qoa6Ht6s8_1(.din(n17479), .dout(n17482));
    jdff dff_B_S0q4jkJ69_1(.din(n4567), .dout(n17485));
    jdff dff_B_7ueIVrlP4_1(.din(n17485), .dout(n17488));
    jdff dff_B_mAlA7HAG8_1(.din(n17488), .dout(n17491));
    jdff dff_A_mfsUWL0M9_1(.din(n2268), .dout(n17493));
    jdff dff_B_0iqja61s8_1(.din(n2233), .dout(n17497));
    jdff dff_B_EKjZM2YP1_1(.din(n17497), .dout(n17500));
    jdff dff_B_8z1ZQthU8_1(.din(n17500), .dout(n17503));
    jdff dff_B_WzlzO9Pe6_1(.din(n17503), .dout(n17506));
    jdff dff_B_xABjFLal2_1(.din(n2236), .dout(n17509));
    jdff dff_B_X11dDHA70_1(.din(n17509), .dout(n17512));
    jdff dff_B_N0rTAIrb9_1(.din(n17512), .dout(n17515));
    jdff dff_A_ls8UL0Zm0_1(.din(n17520), .dout(n17517));
    jdff dff_A_IYJMrDp93_1(.din(n2260), .dout(n17520));
    jdff dff_A_iWDqtKCR1_0(.din(n17545), .dout(n17523));
    jdff dff_A_wS2vt67i1_0(.din(n17529), .dout(n17526));
    jdff dff_A_2ZtELZvn1_0(.din(n17532), .dout(n17529));
    jdff dff_A_12ZkINdP0_0(.din(n2240), .dout(n17532));
    jdff dff_A_z7p6YUjr6_1(.din(n17538), .dout(n17535));
    jdff dff_A_TJs1W6DT4_1(.din(n2240), .dout(n17538));
    jdff dff_A_Gva3RcoY4_2(.din(n17545), .dout(n17541));
    jdff dff_B_8YMo3sLn6_3(.din(n576), .dout(n17545));
    jdff dff_A_eNIehFkN6_0(.din(n17550), .dout(n17547));
    jdff dff_A_9sijSR7X7_0(.din(n17553), .dout(n17550));
    jdff dff_A_YeTVb28I2_0(.din(G534), .dout(n17553));
    jdff dff_A_uj2YxGOe0_1(.din(n17559), .dout(n17556));
    jdff dff_A_uacR1U299_1(.din(n17593), .dout(n17559));
    jdff dff_A_7rkIrt1C7_2(.din(n17593), .dout(n17562));
    jdff dff_B_PgG8jdQ65_3(.din(n4561), .dout(n17566));
    jdff dff_B_G1Da8Jhw2_3(.din(n17566), .dout(n17569));
    jdff dff_B_Z2ESZr7E7_3(.din(n17569), .dout(n17572));
    jdff dff_B_FP36ZvEP7_3(.din(n17572), .dout(n17575));
    jdff dff_B_H0CS5pZQ4_3(.din(n17575), .dout(n17578));
    jdff dff_B_3ffLWUqT4_3(.din(n17578), .dout(n17581));
    jdff dff_B_nUYSVcto3_3(.din(n17581), .dout(n17584));
    jdff dff_B_Fvxerrtk9_3(.din(n17584), .dout(n17587));
    jdff dff_B_sdwmjEXH9_3(.din(n17587), .dout(n17590));
    jdff dff_B_1mfQGzjy0_3(.din(n17590), .dout(n17593));
    jdff dff_A_rBMiAk2D1_0(.din(n17598), .dout(n17595));
    jdff dff_A_OCUCIsPn8_0(.din(n17601), .dout(n17598));
    jdff dff_A_Rs7jDHPV2_0(.din(n17604), .dout(n17601));
    jdff dff_A_GzMljIXB9_0(.din(n17607), .dout(n17604));
    jdff dff_A_AbNsvuMK8_0(.din(n17610), .dout(n17607));
    jdff dff_A_LcXRCDil6_0(.din(n17613), .dout(n17610));
    jdff dff_A_kBWWMt8I3_0(.din(n17616), .dout(n17613));
    jdff dff_A_5Rwlu8WZ7_0(.din(n17619), .dout(n17616));
    jdff dff_A_J0FTVxWY9_0(.din(n17622), .dout(n17619));
    jdff dff_A_mkjfvBAA2_0(.din(n17625), .dout(n17622));
    jdff dff_A_xNidbHy21_0(.din(n17628), .dout(n17625));
    jdff dff_A_HzJQC4BY7_0(.din(n17631), .dout(n17628));
    jdff dff_A_Jsb5G67L3_0(.din(G2174), .dout(n17631));
    jdff dff_A_3XgOyV4A3_1(.din(n17637), .dout(n17634));
    jdff dff_A_l5Fp4qqx5_1(.din(n17640), .dout(n17637));
    jdff dff_A_RpzViQAF7_1(.din(n17643), .dout(n17640));
    jdff dff_A_FKCEAtMd9_1(.din(n17646), .dout(n17643));
    jdff dff_A_4leJHROL5_1(.din(n17649), .dout(n17646));
    jdff dff_A_kt02p7lV7_1(.din(n17652), .dout(n17649));
    jdff dff_A_FcLCn6tK6_1(.din(n17655), .dout(n17652));
    jdff dff_A_tRzY0CQz2_1(.din(n17658), .dout(n17655));
    jdff dff_A_0oDtY7i71_1(.din(n17661), .dout(n17658));
    jdff dff_A_ibm6KBV90_1(.din(G2174), .dout(n17661));
    jdff dff_A_xGYv2QMQ1_0(.din(n4554), .dout(n17664));
    jdff dff_B_96UzNQdT7_0(.din(n4550), .dout(n17668));
    jdff dff_B_T4ChUrjp5_0(.din(n17668), .dout(n17671));
    jdff dff_A_c6y1Byqp4_0(.din(n17676), .dout(n17673));
    jdff dff_A_akJRuCx35_0(.din(n17679), .dout(n17676));
    jdff dff_A_TG9rKCVs5_0(.din(n17683), .dout(n17679));
    jdff dff_B_dxrmcj3p8_2(.din(n668), .dout(n17683));
    jdff dff_A_BCOMpbI92_0(.din(n17688), .dout(n17685));
    jdff dff_A_jIE75rIy5_0(.din(n17691), .dout(n17688));
    jdff dff_A_DlOB61Du6_0(.din(G490), .dout(n17691));
    jdff dff_A_fl2XX5NO3_1(.din(n17697), .dout(n17694));
    jdff dff_A_KzDCsPxR0_1(.din(n17700), .dout(n17697));
    jdff dff_A_CuvyOiKi4_1(.din(n17703), .dout(n17700));
    jdff dff_A_CseopRmD1_1(.din(n17706), .dout(n17703));
    jdff dff_A_DtV5yOsa7_1(.din(n17709), .dout(n17706));
    jdff dff_A_Av5iEvP98_1(.din(n17712), .dout(n17709));
    jdff dff_A_cY01WQiF5_1(.din(n17715), .dout(n17712));
    jdff dff_A_8SolGUlR1_1(.din(n17814), .dout(n17715));
    jdff dff_A_MaZmCqmi6_0(.din(n17721), .dout(n17718));
    jdff dff_A_7DuDT1AJ7_0(.din(n17724), .dout(n17721));
    jdff dff_A_y04Tg1jh5_0(.din(n17727), .dout(n17724));
    jdff dff_A_YnXvQpkT4_0(.din(n1595), .dout(n17727));
    jdff dff_A_KcQBLqEE2_2(.din(n17733), .dout(n17730));
    jdff dff_A_lxg9sKrs5_2(.din(n1595), .dout(n17733));
    jdff dff_A_ohMqcqoZ8_1(.din(G293), .dout(n17736));
    jdff dff_A_IkZ0w3dF1_1(.din(n17742), .dout(n17739));
    jdff dff_A_LIpZI4sY9_1(.din(n17745), .dout(n17742));
    jdff dff_A_h9jhfxll5_1(.din(n17748), .dout(n17745));
    jdff dff_A_1cjKdCl93_1(.din(n1988), .dout(n17748));
    jdff dff_B_L78YjEUY2_1(.din(n1970), .dout(n17752));
    jdff dff_B_6s7BJUn44_1(.din(n17752), .dout(n17755));
    jdff dff_A_bMOUi0UJ9_1(.din(n17760), .dout(n17757));
    jdff dff_A_mU1xbz8d0_1(.din(n17763), .dout(n17760));
    jdff dff_A_89hbxUXa5_1(.din(n17766), .dout(n17763));
    jdff dff_A_9WVpNVBm1_1(.din(n17769), .dout(n17766));
    jdff dff_A_sinFkYgd5_1(.din(n17772), .dout(n17769));
    jdff dff_A_Y2fP7vZz7_1(.din(n17775), .dout(n17772));
    jdff dff_A_QbkPiTFN8_1(.din(n1974), .dout(n17775));
    jdff dff_B_asLk4WND6_0(.din(n1644), .dout(n17779));
    jdff dff_B_tschl8w45_1(.din(G323), .dout(n17782));
    jdff dff_A_gRwoKJ1I1_2(.din(G316), .dout(n17784));
    jdff dff_A_9Xax7Uze0_1(.din(n17790), .dout(n17787));
    jdff dff_A_WFQWTIZ04_1(.din(n17793), .dout(n17790));
    jdff dff_A_YhHvhUHd6_1(.din(n17796), .dout(n17793));
    jdff dff_A_S77Krj036_1(.din(G490), .dout(n17796));
    jdff dff_A_ebeDXyY83_2(.din(n17802), .dout(n17799));
    jdff dff_A_D8d91TvS3_2(.din(n17805), .dout(n17802));
    jdff dff_A_UsOjqMgw6_2(.din(n17808), .dout(n17805));
    jdff dff_A_lcGgPAjg9_2(.din(G490), .dout(n17808));
    jdff dff_A_xFdiiL3z1_0(.din(n17818), .dout(n17811));
    jdff dff_A_BrKvvSPn1_0(.din(n17818), .dout(n17814));
    jdff dff_B_r3BFdL1o3_3(.din(n1633), .dout(n17818));
    jdff dff_A_qKiqqAVL5_0(.din(n1629), .dout(n17820));
    jdff dff_B_xOOQgFa32_1(.din(n1621), .dout(n17824));
    jdff dff_B_IrD5C1yu8_1(.din(G315), .dout(n17827));
    jdff dff_A_Xsngfe2U3_0(.din(n17832), .dout(n17829));
    jdff dff_A_f4tHy0gm6_0(.din(n17836), .dout(n17832));
    jdff dff_B_zrNIoY7t3_2(.din(n716), .dout(n17836));
    jdff dff_A_exMnkZjk4_0(.din(n17841), .dout(n17838));
    jdff dff_A_fwH1ofpW3_0(.din(n17844), .dout(n17841));
    jdff dff_A_U2B1WQkS2_0(.din(G479), .dout(n17844));
    jdff dff_A_ktMtPHfW7_1(.din(n17850), .dout(n17847));
    jdff dff_A_LtTTofiA0_1(.din(n17853), .dout(n17850));
    jdff dff_A_EbD5XZ6A1_1(.din(G479), .dout(n17853));
    jdff dff_A_5E871zXd0_1(.din(n17859), .dout(n17856));
    jdff dff_A_jkidX6wY6_1(.din(n17862), .dout(n17859));
    jdff dff_A_FpBvAnXV4_1(.din(n17865), .dout(n17862));
    jdff dff_A_hVwjUmak5_1(.din(n1610), .dout(n17865));
    jdff dff_A_gEJ9SdA75_2(.din(n17871), .dout(n17868));
    jdff dff_A_Uo8RRHtf5_2(.din(n17874), .dout(n17871));
    jdff dff_A_JuVocacq3_2(.din(n17877), .dout(n17874));
    jdff dff_A_GgqagvSJ3_2(.din(n17880), .dout(n17877));
    jdff dff_A_E5nnNKxj8_2(.din(n1610), .dout(n17880));
    jdff dff_B_J7QSLHkv8_0(.din(n1606), .dout(n17884));
    jdff dff_B_G0FqcR0X5_1(.din(G307), .dout(n17887));
    jdff dff_A_etQq017Q2_0(.din(G302), .dout(n17889));
    jdff dff_A_kGtQubRU4_1(.din(G302), .dout(n17892));
    jdff dff_B_h14bxRSR8_1(.din(n1916), .dout(n17896));
    jdff dff_A_UPDBQr5m9_0(.din(n1560), .dout(n17898));
    jdff dff_A_xmHMGbPn5_1(.din(n17904), .dout(n17901));
    jdff dff_A_1wofKjqD7_1(.din(n1560), .dout(n17904));
    jdff dff_B_Ye6HFRXg6_1(.din(n1552), .dout(n17908));
    jdff dff_A_MJ0ViibJ4_0(.din(G366), .dout(n17910));
    jdff dff_A_ebIdPORu4_0(.din(G332), .dout(n17913));
    jdff dff_A_5elyxUXx2_2(.din(G332), .dout(n17916));
    jdff dff_A_HMrfA5Gf4_0(.din(n17922), .dout(n17919));
    jdff dff_A_pQe7xHr40_0(.din(n17925), .dout(n17922));
    jdff dff_A_nGDxQYAn0_0(.din(n1533), .dout(n17925));
    jdff dff_A_iHYFifiN4_2(.din(n1533), .dout(n17928));
    jdff dff_A_qeIdu1Xg2_0(.din(G358), .dout(n17931));
    jdff dff_A_jmzSzmoB4_1(.din(n1521), .dout(n17934));
    jdff dff_A_SNlAwwOi8_2(.din(G351), .dout(n17937));
    jdff dff_A_5ATc7Gsn9_0(.din(n17943), .dout(n17940));
    jdff dff_A_u6gIaMjr6_0(.din(n17946), .dout(n17943));
    jdff dff_A_LAEMmbVG5_0(.din(G534), .dout(n17946));
    jdff dff_A_0Z1fpFhw9_2(.din(n17952), .dout(n17949));
    jdff dff_A_h2orIroB3_2(.din(n17955), .dout(n17952));
    jdff dff_A_uz8yns7j3_2(.din(G534), .dout(n17955));
    jdff dff_A_wogrT4di4_0(.din(n17961), .dout(n17958));
    jdff dff_A_qDepDr3V9_0(.din(n1913), .dout(n17961));
    jdff dff_A_hItFPknl1_0(.din(G348), .dout(n17964));
    jdff dff_A_FPSHAf153_1(.din(G332), .dout(n17967));
    jdff dff_A_tpYJbV0X3_1(.din(n1505), .dout(n17970));
    jdff dff_A_r9ppHhem0_2(.din(G341), .dout(n17973));
    jdff dff_A_vNWGVL5O1_0(.din(n17983), .dout(n17976));
    jdff dff_A_jcIciAi55_2(.din(n17983), .dout(n17979));
    jdff dff_B_43Qwqhk89_3(.din(n621), .dout(n17983));
    jdff dff_A_y5zcxQJw1_0(.din(n17988), .dout(n17985));
    jdff dff_A_58qlD1fI5_0(.din(n17991), .dout(n17988));
    jdff dff_A_RzdvU1OF3_0(.din(G523), .dout(n17991));
    jdff dff_A_jc1tYchS5_1(.din(n17997), .dout(n17994));
    jdff dff_A_lp7GHm1F6_1(.din(n18000), .dout(n17997));
    jdff dff_A_5oDTPYdf1_1(.din(G523), .dout(n18000));
    jdff dff_A_yoxJaAYq4_1(.din(n18006), .dout(n18003));
    jdff dff_A_nbuYs9md5_1(.din(n18009), .dout(n18006));
    jdff dff_A_w06BWhO72_1(.din(G523), .dout(n18009));
    jdff dff_A_toLwCWIm7_2(.din(n18015), .dout(n18012));
    jdff dff_A_4lpIsodn8_2(.din(n18018), .dout(n18015));
    jdff dff_A_jo6hae3s0_2(.din(G523), .dout(n18018));
    jdff dff_A_95nW45hR3_1(.din(n18024), .dout(n18021));
    jdff dff_A_Ud1hYCRi0_1(.din(n18027), .dout(n18024));
    jdff dff_A_qV2cdtfx4_1(.din(n18030), .dout(n18027));
    jdff dff_A_8hthiOcC1_1(.din(n1898), .dout(n18030));
    jdff dff_A_mwgLu1SD4_1(.din(n18036), .dout(n18033));
    jdff dff_A_lCkwKWrU1_1(.din(n18039), .dout(n18036));
    jdff dff_A_M4yv3f1H0_1(.din(n18042), .dout(n18039));
    jdff dff_A_I7cHtpOf1_1(.din(n18045), .dout(n18042));
    jdff dff_A_XKG0JAaY6_1(.din(n1894), .dout(n18045));
    jdff dff_A_pdF4pMba5_1(.din(n18051), .dout(n18048));
    jdff dff_A_ZNLjUrh03_1(.din(n1497), .dout(n18051));
    jdff dff_A_RfHlSoqf7_0(.din(G338), .dout(n18054));
    jdff dff_A_PQmDPWnJ9_0(.din(n18060), .dout(n18057));
    jdff dff_A_3n8RWLgq4_0(.din(G514), .dout(n18060));
    jdff dff_A_khKlBzin5_2(.din(G514), .dout(n18063));
    jdff dff_A_zBOEPcfw3_1(.din(n18069), .dout(n18066));
    jdff dff_A_qwX6CVHe2_1(.din(n18072), .dout(n18069));
    jdff dff_A_A6QyrXHa2_1(.din(n18075), .dout(n18072));
    jdff dff_A_p4Fayc1v9_1(.din(n1890), .dout(n18075));
    jdff dff_A_pbft6EN75_1(.din(n18081), .dout(n18078));
    jdff dff_A_v9ao2i6o1_1(.din(n18084), .dout(n18081));
    jdff dff_A_uqg8fGWl4_1(.din(n18087), .dout(n18084));
    jdff dff_A_XfTKPgdB9_1(.din(n18090), .dout(n18087));
    jdff dff_A_1awB07r12_1(.din(n1886), .dout(n18090));
    jdff dff_B_57G6NsdX4_0(.din(n1485), .dout(n18094));
    jdff dff_A_R1RIDmXh3_1(.din(G331), .dout(n18096));
    jdff dff_A_F8Uk3U9y7_1(.din(G324), .dout(n18099));
    jdff dff_A_zFfp6bVg0_2(.din(G324), .dout(n18102));
    jdff dff_A_VICh85vW4_0(.din(n18108), .dout(n18105));
    jdff dff_A_R6CvotoX6_0(.din(n18111), .dout(n18108));
    jdff dff_A_jKyAwvkP8_0(.din(n18114), .dout(n18111));
    jdff dff_A_GN83aTc42_0(.din(G503), .dout(n18114));
    jdff dff_A_10AtPci18_2(.din(n18120), .dout(n18117));
    jdff dff_A_NJpbWQ6H2_2(.din(G503), .dout(n18120));
    jdff dff_A_EIhQxOxi1_0(.din(n18126), .dout(n18123));
    jdff dff_A_qJsf05Up1_0(.din(n18129), .dout(n18126));
    jdff dff_A_wYSDX8fS2_0(.din(n18132), .dout(n18129));
    jdff dff_A_VOUIoQCP5_0(.din(n18135), .dout(n18132));
    jdff dff_A_TAJot7FE7_0(.din(n18138), .dout(n18135));
    jdff dff_A_uISgwoQ22_0(.din(n18141), .dout(n18138));
    jdff dff_A_oTkjMKGO6_0(.din(n18144), .dout(n18141));
    jdff dff_A_9LdN4vs39_0(.din(n18147), .dout(n18144));
    jdff dff_A_kh43U5pn6_0(.din(n18150), .dout(n18147));
    jdff dff_A_4bJdu3ei3_0(.din(n18153), .dout(n18150));
    jdff dff_A_UvAzVEjK0_0(.din(n18156), .dout(n18153));
    jdff dff_A_djvkdCPF3_0(.din(n18159), .dout(n18156));
    jdff dff_A_ArpKi3J15_0(.din(n18162), .dout(n18159));
    jdff dff_A_opWE1Xsm3_0(.din(n18165), .dout(n18162));
    jdff dff_A_5H3EhhXK2_0(.din(n18168), .dout(n18165));
    jdff dff_A_AwplXlA05_0(.din(n18171), .dout(n18168));
    jdff dff_A_SvU9OCQG5_0(.din(n18174), .dout(n18171));
    jdff dff_A_PfGgEJzT3_0(.din(n18177), .dout(n18174));
    jdff dff_A_r73D5zJI9_0(.din(n18180), .dout(n18177));
    jdff dff_A_xXFR20xn1_0(.din(G4092), .dout(n18180));
    jdff dff_A_kn2ty5aY0_2(.din(n18186), .dout(n18183));
    jdff dff_A_4QZMshbv7_2(.din(n18189), .dout(n18186));
    jdff dff_A_0DjVm3660_2(.din(n18192), .dout(n18189));
    jdff dff_A_8AaK8aOG1_2(.din(G4092), .dout(n18192));
    jdff dff_B_OQgniS8Z0_0(.din(n5583), .dout(n18196));
    jdff dff_B_c7wDodW81_0(.din(n18196), .dout(n18199));
    jdff dff_B_dxlYHcWx4_0(.din(n18199), .dout(n18202));
    jdff dff_B_Ukh7m1Bv2_0(.din(n18202), .dout(n18205));
    jdff dff_B_7QClgarR9_0(.din(n18205), .dout(n18208));
    jdff dff_B_H1gZ39aE4_0(.din(n18208), .dout(n18211));
    jdff dff_B_d2uBp8jE2_0(.din(n18211), .dout(n18214));
    jdff dff_B_5OCG9Rsg8_0(.din(n18214), .dout(n18217));
    jdff dff_B_9qu58Pm82_0(.din(n18217), .dout(n18220));
    jdff dff_B_qKqzwTI43_0(.din(n18220), .dout(n18223));
    jdff dff_B_FNlDNXDC1_0(.din(n18223), .dout(n18226));
    jdff dff_B_RH52Fyov0_0(.din(n18226), .dout(n18229));
    jdff dff_B_iQyb6XoS3_0(.din(n18229), .dout(n18232));
    jdff dff_B_SkypU4MT0_0(.din(n18232), .dout(n18235));
    jdff dff_B_L8xjIghs4_0(.din(n18235), .dout(n18238));
    jdff dff_B_OnK7SI3H5_0(.din(n18238), .dout(n18241));
    jdff dff_B_WPf0bgdS4_0(.din(n18241), .dout(n18244));
    jdff dff_B_8UmPLGEf0_0(.din(n18244), .dout(n18247));
    jdff dff_B_UAoLTV0I0_0(.din(n18247), .dout(n18250));
    jdff dff_B_FRDYFa6S5_1(.din(n5254), .dout(n18253));
    jdff dff_B_vce812uo3_1(.din(n18253), .dout(n18256));
    jdff dff_B_qfHGV0D74_1(.din(n18256), .dout(n18259));
    jdff dff_B_efRlcB7r5_1(.din(n18259), .dout(n18262));
    jdff dff_B_LEQP3c7v9_1(.din(n18262), .dout(n18265));
    jdff dff_B_7dmBLewq7_1(.din(n18265), .dout(n18268));
    jdff dff_B_t6fAe9au6_1(.din(n18268), .dout(n18271));
    jdff dff_B_1X3yTzcg9_1(.din(n18271), .dout(n18274));
    jdff dff_B_6iQyRD5L9_1(.din(n5512), .dout(n18277));
    jdff dff_B_Nb21UJTq6_1(.din(n18277), .dout(n18280));
    jdff dff_A_xlkFGP9J9_2(.din(n18285), .dout(n18282));
    jdff dff_A_4SjY06lH7_2(.din(n1379), .dout(n18285));
    jdff dff_A_L7QMeyn52_1(.din(n5501), .dout(n18288));
    jdff dff_B_QoTvP5CI6_0(.din(n5489), .dout(n18292));
    jdff dff_B_kEmmUmCN9_1(.din(n5473), .dout(n18295));
    jdff dff_B_U1nnP5rN5_1(.din(n18295), .dout(n18298));
    jdff dff_B_WBi1Vhx51_1(.din(n18298), .dout(n18301));
    jdff dff_B_8IX8KGr32_1(.din(n18301), .dout(n18304));
    jdff dff_B_8cdrglPg3_1(.din(n18304), .dout(n18307));
    jdff dff_B_keaKlAXc1_1(.din(n5446), .dout(n18310));
    jdff dff_B_KfVMJ9oW4_1(.din(n18310), .dout(n18313));
    jdff dff_B_u1f4EHL35_0(.din(n5458), .dout(n18316));
    jdff dff_B_T8eDJLQt1_0(.din(n5454), .dout(n18319));
    jdff dff_A_Uws9P4kF7_1(.din(n18324), .dout(n18321));
    jdff dff_A_3trX53hq8_1(.din(n18327), .dout(n18324));
    jdff dff_A_QtIGU6nu1_1(.din(n18330), .dout(n18327));
    jdff dff_A_FyMgIb5q1_1(.din(n18333), .dout(n18330));
    jdff dff_A_oMSGCTfm4_1(.din(n18336), .dout(n18333));
    jdff dff_A_1f2BLEyN8_1(.din(n18339), .dout(n18336));
    jdff dff_A_1UZuqTSm6_1(.din(n1460), .dout(n18339));
    jdff dff_A_rUws5IQk5_1(.din(n18345), .dout(n18342));
    jdff dff_A_vvzJet7l9_1(.din(n18348), .dout(n18345));
    jdff dff_A_bID7jaFa3_1(.din(n18351), .dout(n18348));
    jdff dff_A_MTSappig0_1(.din(n18354), .dout(n18351));
    jdff dff_A_5r6h0yxY4_1(.din(n18357), .dout(n18354));
    jdff dff_A_qKtk3BAZ0_1(.din(n18361), .dout(n18357));
    jdff dff_B_06dA8gXU0_2(.din(n2805), .dout(n18361));
    jdff dff_A_moXGfcut3_2(.din(n18366), .dout(n18363));
    jdff dff_A_kxwH2KKG7_2(.din(n18369), .dout(n18366));
    jdff dff_A_4VevNxZE6_2(.din(n18372), .dout(n18369));
    jdff dff_A_MBniGXJD5_2(.din(n18375), .dout(n18372));
    jdff dff_A_GBmzx6wz4_2(.din(n2717), .dout(n18375));
    jdff dff_B_z6k5rTOH2_1(.din(n1838), .dout(n18379));
    jdff dff_B_cvGlQ0044_1(.din(n18379), .dout(n18382));
    jdff dff_B_bsMZhnDY2_1(.din(n18382), .dout(n18385));
    jdff dff_B_ttpy0CZW9_1(.din(n1842), .dout(n18388));
    jdff dff_B_3VKKs2DS2_1(.din(n18388), .dout(n18391));
    jdff dff_A_fZQ7cme07_1(.din(n18396), .dout(n18393));
    jdff dff_A_Aco4Rfxw7_1(.din(n18399), .dout(n18396));
    jdff dff_A_EUgEOsnn9_1(.din(n18402), .dout(n18399));
    jdff dff_A_khJRHsrT5_1(.din(n18405), .dout(n18402));
    jdff dff_A_OY7Q8sWP2_1(.din(n18408), .dout(n18405));
    jdff dff_A_9aUQXAKb9_1(.din(n18411), .dout(n18408));
    jdff dff_A_srQ6aHx94_1(.din(n1862), .dout(n18411));
    jdff dff_A_mi9eGh4F5_0(.din(n18417), .dout(n18414));
    jdff dff_A_rLAMROX73_0(.din(n18420), .dout(n18417));
    jdff dff_A_enGQamJO4_0(.din(n18423), .dout(n18420));
    jdff dff_A_62LuOKr94_0(.din(n18426), .dout(n18423));
    jdff dff_A_ji7Ssb0i9_0(.din(n18429), .dout(n18426));
    jdff dff_A_FHuImOqd3_0(.din(n18432), .dout(n18429));
    jdff dff_A_8VYSaQLh2_0(.din(n18435), .dout(n18432));
    jdff dff_A_F7FvTbIU6_0(.din(n1850), .dout(n18435));
    jdff dff_A_xXu241s53_0(.din(n18441), .dout(n18438));
    jdff dff_A_GPjp26wa3_0(.din(n18444), .dout(n18441));
    jdff dff_A_mqHihzL63_0(.din(n18447), .dout(n18444));
    jdff dff_A_Dp3jRNxF2_0(.din(n18450), .dout(n18447));
    jdff dff_A_1T9U05Yz1_0(.din(n1414), .dout(n18450));
    jdff dff_A_dpYbe0Vd4_0(.din(n18456), .dout(n18453));
    jdff dff_A_JOATgsfg6_0(.din(n19174), .dout(n18456));
    jdff dff_A_37apWN0E4_0(.din(n18462), .dout(n18459));
    jdff dff_A_LEtQZjGE5_0(.din(n18469), .dout(n18462));
    jdff dff_B_cPd2n3vn8_2(.din(n5442), .dout(n18466));
    jdff dff_B_pJnT534a4_2(.din(n18466), .dout(n18469));
    jdff dff_A_mirKFcdb1_1(.din(n18474), .dout(n18471));
    jdff dff_A_8b2e4GZU0_1(.din(n18477), .dout(n18474));
    jdff dff_A_1dhyPwgU6_1(.din(n18480), .dout(n18477));
    jdff dff_A_xHW8LyAM9_1(.din(n18483), .dout(n18480));
    jdff dff_A_Wjj189Lq3_1(.din(n18486), .dout(n18483));
    jdff dff_A_qGF3hIIh8_1(.din(n18489), .dout(n18486));
    jdff dff_A_oNpKmeNu2_1(.din(n18492), .dout(n18489));
    jdff dff_A_L83vThpW0_1(.din(n18495), .dout(n18492));
    jdff dff_A_PhQ3LTox0_1(.din(n18498), .dout(n18495));
    jdff dff_A_enWkxjoB9_1(.din(n1456), .dout(n18498));
    jdff dff_A_EMhCsHJR1_2(.din(n1456), .dout(n18501));
    jdff dff_B_EXzRqPhv9_0(.din(n1448), .dout(n18505));
    jdff dff_B_vbotFnb24_1(.din(G217), .dout(n18508));
    jdff dff_A_Rr5OZwbN8_0(.din(n1395), .dout(n18510));
    jdff dff_A_4x3qatY19_2(.din(n18516), .dout(n18513));
    jdff dff_A_8mxpvWCz0_2(.din(n18519), .dout(n18516));
    jdff dff_A_Yv6kDql04_2(.din(n18522), .dout(n18519));
    jdff dff_A_ib9Rh1lq1_2(.din(n1395), .dout(n18522));
    jdff dff_B_qtKr0fpF5_1(.din(n1383), .dout(n18526));
    jdff dff_B_O0nRUcvV3_1(.din(G209), .dout(n18529));
    jdff dff_A_fpZxkH2L2_0(.din(n1433), .dout(n18531));
    jdff dff_A_BmdpZ4Lh4_0(.din(n18537), .dout(n18534));
    jdff dff_A_4cNbMmsO6_0(.din(n1854), .dout(n18537));
    jdff dff_A_r3NdDLcl6_2(.din(n18543), .dout(n18540));
    jdff dff_A_mLhvBfUC2_2(.din(n18546), .dout(n18543));
    jdff dff_A_weVSCX4f8_2(.din(n18549), .dout(n18546));
    jdff dff_A_g4AstPkX1_2(.din(n18552), .dout(n18549));
    jdff dff_A_cRaF1Mbl7_2(.din(n18555), .dout(n18552));
    jdff dff_A_G6qPK8wB9_2(.din(n18558), .dout(n18555));
    jdff dff_A_xgc5JR2D4_2(.din(n2775), .dout(n18558));
    jdff dff_B_K5Phutoi0_2(.din(n5426), .dout(n18562));
    jdff dff_A_7Weigvoq1_1(.din(n1846), .dout(n18564));
    jdff dff_B_G1yOpguQ2_0(.din(n1425), .dout(n18568));
    jdff dff_B_y63hCaOL7_1(.din(G225), .dout(n18571));
    jdff dff_B_Yd1FmHXW5_0(.din(n1406), .dout(n18574));
    jdff dff_B_8f4RVvMu5_1(.din(G233), .dout(n18577));
    jdff dff_A_VySiNYam7_1(.din(n1822), .dout(n18579));
    jdff dff_A_BLVgBP3s8_0(.din(n18585), .dout(n18582));
    jdff dff_A_KaP3mLZ20_0(.din(n18595), .dout(n18585));
    jdff dff_B_8quRQZr08_2(.din(n1752), .dout(n18589));
    jdff dff_B_PGJ73wt72_2(.din(n18589), .dout(n18592));
    jdff dff_B_i8QFpFER7_2(.din(n18592), .dout(n18595));
    jdff dff_A_hyklK2l55_0(.din(n18600), .dout(n18597));
    jdff dff_A_B2v12AOc4_0(.din(n18603), .dout(n18600));
    jdff dff_A_HKTgWa7w6_0(.din(n18606), .dout(n18603));
    jdff dff_A_Awaqc4aS2_0(.din(n1749), .dout(n18606));
    jdff dff_A_2QmQ8UmM1_1(.din(n18612), .dout(n18609));
    jdff dff_A_0VGBal8i6_1(.din(n18615), .dout(n18612));
    jdff dff_A_WHOrqpLf1_1(.din(n18618), .dout(n18615));
    jdff dff_A_mp2OLete7_1(.din(n18621), .dout(n18618));
    jdff dff_A_RIzCUENo3_1(.din(n18624), .dout(n18621));
    jdff dff_A_Xw0QZFdE1_1(.din(n1742), .dout(n18624));
    jdff dff_A_MXSlLSCG9_2(.din(n18630), .dout(n18627));
    jdff dff_A_UexTmkzh5_2(.din(n18633), .dout(n18630));
    jdff dff_A_2JeTvPl28_2(.din(n18636), .dout(n18633));
    jdff dff_A_obhZ1qgF7_2(.din(n18639), .dout(n18636));
    jdff dff_A_9OxIGf3C9_2(.din(n18642), .dout(n18639));
    jdff dff_A_NxH4tdPn0_2(.din(n1742), .dout(n18642));
    jdff dff_B_kghlOlOs9_0(.din(n5415), .dout(n18646));
    jdff dff_B_h6UqhT4u7_0(.din(n18646), .dout(n18649));
    jdff dff_B_ZRUgqySz6_0(.din(n18649), .dout(n18652));
    jdff dff_B_cgW0hOZr8_0(.din(n18652), .dout(n18655));
    jdff dff_B_wcYJ1TzN1_0(.din(n18655), .dout(n18658));
    jdff dff_B_BrCnk7Kw2_0(.din(n18658), .dout(n18661));
    jdff dff_B_SmgpBJxx1_0(.din(n18661), .dout(n18664));
    jdff dff_B_jFPfXCOu8_0(.din(n18664), .dout(n18667));
    jdff dff_B_kmufscFm5_0(.din(n18667), .dout(n18670));
    jdff dff_B_2j0nYXVw6_0(.din(n5407), .dout(n18673));
    jdff dff_B_6bkGyK2w7_0(.din(n18673), .dout(n18676));
    jdff dff_B_NmUcLTXn0_1(.din(n5395), .dout(n18679));
    jdff dff_B_8COAyz5T1_1(.din(n5387), .dout(n18682));
    jdff dff_B_4grUwu5F0_1(.din(n18682), .dout(n18685));
    jdff dff_A_NxE5199g4_0(.din(n18690), .dout(n18687));
    jdff dff_A_c1571MWv0_0(.din(n18727), .dout(n18690));
    jdff dff_B_1UAZNobP5_2(.din(n5367), .dout(n18694));
    jdff dff_B_VNHm9cY24_2(.din(n18694), .dout(n18697));
    jdff dff_B_918j1l7K2_2(.din(n18697), .dout(n18700));
    jdff dff_B_VjbN95og9_2(.din(n18700), .dout(n18703));
    jdff dff_B_fivtRROq9_2(.din(n18703), .dout(n18706));
    jdff dff_B_ux2iu24m6_2(.din(n18706), .dout(n18709));
    jdff dff_B_6ape9e1y0_2(.din(n18709), .dout(n18712));
    jdff dff_B_7HdnSMWM1_2(.din(n18712), .dout(n18715));
    jdff dff_B_TWfjzTAo4_2(.din(n18715), .dout(n18718));
    jdff dff_B_3apDr30h5_2(.din(n18718), .dout(n18721));
    jdff dff_B_Ujo9Syr77_2(.din(n18721), .dout(n18724));
    jdff dff_B_fCBI0eF75_2(.din(n18724), .dout(n18727));
    jdff dff_A_Kyha9QU23_0(.din(n18732), .dout(n18729));
    jdff dff_A_LpLLVyIt7_0(.din(n18735), .dout(n18732));
    jdff dff_A_b8Zi22nb3_0(.din(n18738), .dout(n18735));
    jdff dff_A_G8jV60gn7_0(.din(n18741), .dout(n18738));
    jdff dff_A_gv9hIwzM5_0(.din(n18744), .dout(n18741));
    jdff dff_A_efNm6fAq4_0(.din(n18747), .dout(n18744));
    jdff dff_A_7lweI8Tw5_0(.din(n18750), .dout(n18747));
    jdff dff_A_MwC5JsDB6_0(.din(n18753), .dout(n18750));
    jdff dff_A_WqcEn3r81_0(.din(n18756), .dout(n18753));
    jdff dff_A_XuDmv30e4_0(.din(n18759), .dout(n18756));
    jdff dff_A_AccpODWJ0_0(.din(n18762), .dout(n18759));
    jdff dff_A_MVkNx5Pp9_0(.din(n18765), .dout(n18762));
    jdff dff_A_2UiPeyF29_0(.din(n18768), .dout(n18765));
    jdff dff_A_nSdn0rlr3_0(.din(n18771), .dout(n18768));
    jdff dff_A_USsYQNdK9_0(.din(G1497), .dout(n18771));
    jdff dff_A_4ouY8qtj9_1(.din(n18777), .dout(n18774));
    jdff dff_A_F4FUDs3M5_1(.din(n18780), .dout(n18777));
    jdff dff_A_TLumZ1LD0_1(.din(n18783), .dout(n18780));
    jdff dff_A_nq8MFM1V3_1(.din(n18786), .dout(n18783));
    jdff dff_A_OpuR5ybL5_1(.din(n18789), .dout(n18786));
    jdff dff_A_Kyfo73fF2_1(.din(n18792), .dout(n18789));
    jdff dff_A_OAl2Lzxh7_1(.din(n18795), .dout(n18792));
    jdff dff_A_D5i4tLOH4_1(.din(n18798), .dout(n18795));
    jdff dff_A_1Perz2kI6_1(.din(n18801), .dout(n18798));
    jdff dff_A_qGhmJ1uq6_1(.din(n18804), .dout(n18801));
    jdff dff_A_uod133Nn2_1(.din(n18807), .dout(n18804));
    jdff dff_A_fKRahply6_1(.din(G1497), .dout(n18807));
    jdff dff_B_KmuGB4Wa4_1(.din(n5299), .dout(n18811));
    jdff dff_B_2bHVAlJb1_1(.din(n18811), .dout(n18814));
    jdff dff_B_iWpnZ9fZ2_0(.din(n5353), .dout(n18817));
    jdff dff_B_KmjT6LZ54_0(.din(n18817), .dout(n18820));
    jdff dff_B_QXQtFWVM3_0(.din(n18820), .dout(n18823));
    jdff dff_B_KEuu4M2p9_0(.din(n18823), .dout(n18826));
    jdff dff_A_jmLmb4bc5_0(.din(n18831), .dout(n18828));
    jdff dff_A_SdXrTuRN7_0(.din(n5349), .dout(n18831));
    jdff dff_A_KftsghUC4_0(.din(n18837), .dout(n18834));
    jdff dff_A_zQUxjSjB4_0(.din(n18840), .dout(n18837));
    jdff dff_A_1iPsS97d8_0(.din(n18843), .dout(n18840));
    jdff dff_A_S4J3oz055_0(.din(n2436), .dout(n18843));
    jdff dff_A_tLTauKTU4_2(.din(n18849), .dout(n18846));
    jdff dff_A_8QoqLDaH3_2(.din(n18852), .dout(n18849));
    jdff dff_A_j64Xv3qz2_2(.din(n18855), .dout(n18852));
    jdff dff_A_i3G21l3P2_2(.din(n18858), .dout(n18855));
    jdff dff_A_QqAqicj04_2(.din(n2436), .dout(n18858));
    jdff dff_A_6POUhTop1_1(.din(n18864), .dout(n18861));
    jdff dff_A_uIGeh2Lg0_1(.din(n18867), .dout(n18864));
    jdff dff_A_Nbzwjh4j8_1(.din(n18870), .dout(n18867));
    jdff dff_A_oC8bNNVc9_1(.din(n1375), .dout(n18870));
    jdff dff_B_yCM6XrYW8_0(.din(n1367), .dout(n18874));
    jdff dff_B_LGHcPilM5_1(.din(G241), .dout(n18877));
    jdff dff_B_eWV88eXH9_1(.din(n5302), .dout(n18880));
    jdff dff_B_FjYJOSeL0_1(.din(n18880), .dout(n18883));
    jdff dff_B_xDHxEj471_1(.din(n18883), .dout(n18886));
    jdff dff_B_9qF6hteK6_1(.din(n5305), .dout(n18889));
    jdff dff_B_RS5LCjhX5_1(.din(n18889), .dout(n18892));
    jdff dff_A_Z638JVzt5_1(.din(n18897), .dout(n18894));
    jdff dff_A_CvzPEdAw0_1(.din(n18900), .dout(n18897));
    jdff dff_A_5jgei4zv9_1(.din(n1760), .dout(n18900));
    jdff dff_A_thC6SE5m2_1(.din(n18906), .dout(n18903));
    jdff dff_A_v8XxsTxc9_1(.din(n18909), .dout(n18906));
    jdff dff_A_hur0nhdE9_1(.din(n18912), .dout(n18909));
    jdff dff_A_2tTVCuS14_1(.din(n1756), .dout(n18912));
    jdff dff_A_h5ww4nX32_0(.din(n18918), .dout(n18915));
    jdff dff_A_IP7kNLv53_0(.din(n1353), .dout(n18918));
    jdff dff_A_3drH5Idj8_1(.din(n1345), .dout(n18921));
    jdff dff_A_oXcb4rub9_1(.din(n1345), .dout(n18924));
    jdff dff_A_NVFluDeo3_2(.din(n18930), .dout(n18927));
    jdff dff_A_VL4FUWSr8_2(.din(n18933), .dout(n18930));
    jdff dff_A_vLl8KNLZ3_2(.din(n18936), .dout(n18933));
    jdff dff_A_apldzcTr2_2(.din(n1345), .dout(n18936));
    jdff dff_B_36jfe22f8_0(.din(n1337), .dout(n18940));
    jdff dff_B_rh2BxCzh4_1(.din(G264), .dout(n18943));
    jdff dff_A_PZqyPr7U8_1(.din(n18948), .dout(n18945));
    jdff dff_A_ZC2bstJW3_1(.din(n1326), .dout(n18948));
    jdff dff_A_oMKzX95G8_0(.din(n18954), .dout(n18951));
    jdff dff_A_DCcBNEoT4_0(.din(n5296), .dout(n18954));
    jdff dff_B_UZ0RO1iU3_0(.din(n5292), .dout(n18958));
    jdff dff_B_xzfxRi8R7_0(.din(n5288), .dout(n18961));
    jdff dff_B_NbMeyCxI1_0(.din(n5258), .dout(n18964));
    jdff dff_A_E8RvXwhG7_0(.din(n1323), .dout(n18966));
    jdff dff_A_LlCKywvu0_1(.din(n18972), .dout(n18969));
    jdff dff_A_6f9bX2tD6_1(.din(n1323), .dout(n18972));
    jdff dff_B_I6rSOM260_1(.din(n1774), .dout(n18976));
    jdff dff_A_s88eH5Y14_0(.din(n1790), .dout(n18978));
    jdff dff_A_Qe9sEAx29_1(.din(n1790), .dout(n18981));
    jdff dff_A_NHIWFKCJ9_1(.din(n1289), .dout(n18984));
    jdff dff_B_hQ7pqEYK6_1(.din(G280), .dout(n18988));
    jdff dff_A_2L149ccd6_0(.din(n1282), .dout(n18990));
    jdff dff_A_Hv98Ul3Y0_0(.din(n1778), .dout(n18993));
    jdff dff_A_s2LmmwUv5_1(.din(n1270), .dout(n18996));
    jdff dff_B_dcyVP1xp6_1(.din(G288), .dout(n19000));
    jdff dff_A_zuN3zQmS5_0(.din(n1263), .dout(n19002));
    jdff dff_A_qDxhoPsK9_0(.din(n19008), .dout(n19005));
    jdff dff_A_hl6HUjuu1_0(.din(n1771), .dout(n19008));
    jdff dff_A_b2al5vls9_1(.din(n1315), .dout(n19011));
    jdff dff_B_WxmNg9VF5_1(.din(G272), .dout(n19015));
    jdff dff_A_v4ndQapO6_0(.din(n1308), .dout(n19017));
    jdff dff_A_vm5gbBGa0_0(.din(n19023), .dout(n19020));
    jdff dff_A_K02QV1Jy0_0(.din(n19405), .dout(n19023));
    jdff dff_B_889MNSiZ3_0(.din(n5243), .dout(n19027));
    jdff dff_B_Q1twm8zD2_1(.din(n5203), .dout(n19030));
    jdff dff_B_EtmbtrLr8_1(.din(n19030), .dout(n19033));
    jdff dff_A_oLekoJB74_0(.din(G210), .dout(n19035));
    jdff dff_A_v255Axo79_1(.din(n19041), .dout(n19038));
    jdff dff_A_begpvNal4_1(.din(n19045), .dout(n19041));
    jdff dff_B_fLnXQ0Lb0_3(.din(n856), .dout(n19045));
    jdff dff_A_8eZYEhHf5_0(.din(n19050), .dout(n19047));
    jdff dff_A_j9NSDTOJ0_0(.din(n19053), .dout(n19050));
    jdff dff_A_9ln3n0g28_0(.din(n19056), .dout(n19053));
    jdff dff_A_ofFN2KXF6_0(.din(G457), .dout(n19056));
    jdff dff_A_IvhJg8688_1(.din(n19062), .dout(n19059));
    jdff dff_A_Fz4uHTIG0_1(.din(n19065), .dout(n19062));
    jdff dff_A_L5HpIfiT5_1(.din(G457), .dout(n19065));
    jdff dff_A_j1EMTddv1_1(.din(n19071), .dout(n19068));
    jdff dff_A_1KzzcdFs5_1(.din(n19074), .dout(n19071));
    jdff dff_A_y63zbw8x4_1(.din(G457), .dout(n19074));
    jdff dff_A_cKOUHrFF9_2(.din(n19080), .dout(n19077));
    jdff dff_A_rmmWmvdv0_2(.din(n19083), .dout(n19080));
    jdff dff_A_YXtTpnJ03_2(.din(n19086), .dout(n19083));
    jdff dff_A_SfgBxLJ12_2(.din(G457), .dout(n19086));
    jdff dff_A_ObGN1cyK6_2(.din(G210), .dout(n19089));
    jdff dff_B_wX4VpuQn3_1(.din(n5183), .dout(n19093));
    jdff dff_A_5zvoiHyn4_0(.din(n19105), .dout(n19095));
    jdff dff_A_qvgEtbMD4_1(.din(n19101), .dout(n19098));
    jdff dff_A_g2ibEBXg4_1(.din(n19105), .dout(n19101));
    jdff dff_B_HKAzCg7R7_3(.din(n1078), .dout(n19105));
    jdff dff_A_ZPEVKmD71_0(.din(n19110), .dout(n19107));
    jdff dff_A_FkFWjuf19_0(.din(n19113), .dout(n19110));
    jdff dff_A_MAAjVj5D3_0(.din(n19116), .dout(n19113));
    jdff dff_A_A5Y9CIJd1_0(.din(G468), .dout(n19116));
    jdff dff_A_6IczPJFg8_1(.din(n19122), .dout(n19119));
    jdff dff_A_kk6Xg4d20_1(.din(n19125), .dout(n19122));
    jdff dff_A_UmtnvGTW6_1(.din(G468), .dout(n19125));
    jdff dff_B_d0nm04rx4_1(.din(n5167), .dout(n19129));
    jdff dff_A_omqAYVWi0_0(.din(G218), .dout(n19131));
    jdff dff_A_dOKrPts53_1(.din(n19137), .dout(n19134));
    jdff dff_A_Zllgn7rC3_1(.din(G468), .dout(n19137));
    jdff dff_A_M1BjK6yz4_2(.din(n19143), .dout(n19140));
    jdff dff_A_X80VAKJu5_2(.din(n19146), .dout(n19143));
    jdff dff_A_QVEhdUTm7_2(.din(n19149), .dout(n19146));
    jdff dff_A_C4MnImA90_2(.din(G468), .dout(n19149));
    jdff dff_A_GfG3u0CN9_0(.din(G218), .dout(n19152));
    jdff dff_B_Evnm23O15_1(.din(n5127), .dout(n19156));
    jdff dff_B_2GqOtywX5_1(.din(n19156), .dout(n19159));
    jdff dff_A_jKyEDYcW2_0(.din(G226), .dout(n19161));
    jdff dff_A_EnrzktwJ9_2(.din(n19167), .dout(n19164));
    jdff dff_A_2XBEw37y9_2(.din(n19170), .dout(n19167));
    jdff dff_A_Kof4lzNX5_2(.din(n19174), .dout(n19170));
    jdff dff_B_OzpKQcnl0_3(.din(n1028), .dout(n19174));
    jdff dff_A_p5OtCipC7_0(.din(n19179), .dout(n19176));
    jdff dff_A_LtzjnPaH2_0(.din(n19182), .dout(n19179));
    jdff dff_A_byQV1EwN1_0(.din(G422), .dout(n19182));
    jdff dff_A_67X00Ndi9_1(.din(n19188), .dout(n19185));
    jdff dff_A_uxQAF81y4_1(.din(n19191), .dout(n19188));
    jdff dff_A_sS3oEy2s3_1(.din(G422), .dout(n19191));
    jdff dff_A_e1WClZRI7_2(.din(n19197), .dout(n19194));
    jdff dff_A_pbJw1qfz5_2(.din(n19200), .dout(n19197));
    jdff dff_A_U6Ikx0Vg4_2(.din(n19203), .dout(n19200));
    jdff dff_A_M0zNXlLG7_2(.din(G422), .dout(n19203));
    jdff dff_A_gT9buK4T4_2(.din(G226), .dout(n19206));
    jdff dff_B_MT3m1v0b3_1(.din(n1202), .dout(n19210));
    jdff dff_B_Iy94drE61_1(.din(n19210), .dout(n19213));
    jdff dff_B_VYw4pF030_1(.din(n1205), .dout(n19216));
    jdff dff_A_vMNUiQfu8_0(.din(n19221), .dout(n19218));
    jdff dff_A_KR7BGXZC0_0(.din(n19224), .dout(n19221));
    jdff dff_A_ofgL8hNt0_0(.din(G446), .dout(n19224));
    jdff dff_A_PoDJRc4n1_1(.din(n19230), .dout(n19227));
    jdff dff_A_1GH9ejTP0_1(.din(n19233), .dout(n19230));
    jdff dff_A_ClsEoZwW8_1(.din(G446), .dout(n19233));
    jdff dff_A_d9umcNL71_1(.din(n19239), .dout(n19236));
    jdff dff_A_m1ayBrvp4_1(.din(n19242), .dout(n19239));
    jdff dff_A_ZxaHmWHq9_1(.din(G446), .dout(n19242));
    jdff dff_A_TKLUWJgi2_2(.din(n19248), .dout(n19245));
    jdff dff_A_77SFOBKl7_2(.din(n19251), .dout(n19248));
    jdff dff_A_Mmgn51Xh7_2(.din(G446), .dout(n19251));
    jdff dff_A_5HCCnfVr4_0(.din(G206), .dout(n19254));
    jdff dff_B_UhzF9ryi3_1(.din(n5003), .dout(n19258));
    jdff dff_B_wNMw5I5N0_1(.din(n5039), .dout(n19261));
    jdff dff_B_tRZZYgo67_1(.din(n5079), .dout(n19264));
    jdff dff_B_SeD0dRPb3_1(.din(n19264), .dout(n19267));
    jdff dff_A_IAv7bVlJ3_0(.din(G234), .dout(n19269));
    jdff dff_A_k3UyB8Po6_1(.din(n19275), .dout(n19272));
    jdff dff_A_KZ8wSDaz2_1(.din(n19278), .dout(n19275));
    jdff dff_A_vrW7pce47_1(.din(n19282), .dout(n19278));
    jdff dff_B_d2dBaqaS5_3(.din(n898), .dout(n19282));
    jdff dff_A_ixjX31sh3_0(.din(n19287), .dout(n19284));
    jdff dff_A_GtMqQLe60_0(.din(n19290), .dout(n19287));
    jdff dff_A_YbWXFDCo7_0(.din(n19293), .dout(n19290));
    jdff dff_A_ZOupd35Q9_0(.din(G435), .dout(n19293));
    jdff dff_A_4nBuZFG15_1(.din(n19299), .dout(n19296));
    jdff dff_A_fZxMoYKW5_1(.din(n19302), .dout(n19299));
    jdff dff_A_lrnp6gFq2_1(.din(G435), .dout(n19302));
    jdff dff_A_Nnii9NIS3_1(.din(n19308), .dout(n19305));
    jdff dff_A_a1yMwuBY3_1(.din(n19311), .dout(n19308));
    jdff dff_A_qaPcEWrT7_1(.din(G435), .dout(n19311));
    jdff dff_A_N81RKIix8_2(.din(n19317), .dout(n19314));
    jdff dff_A_sFDtG4JR7_2(.din(n19320), .dout(n19317));
    jdff dff_A_Noi6SRXT0_2(.din(n19323), .dout(n19320));
    jdff dff_A_8lsHxblE7_2(.din(G435), .dout(n19323));
    jdff dff_A_zJ4OzjGQ4_2(.din(G234), .dout(n19326));
    jdff dff_B_m6dmyI8h8_1(.din(n5043), .dout(n19330));
    jdff dff_B_GsQmPUvU2_1(.din(n19330), .dout(n19333));
    jdff dff_A_jWHGvtCa9_0(.din(G257), .dout(n19335));
    jdff dff_A_LwEQZpPG1_1(.din(n19341), .dout(n19338));
    jdff dff_A_SsfZd5P01_1(.din(n19345), .dout(n19341));
    jdff dff_B_9BYI8BGR2_3(.din(n1120), .dout(n19345));
    jdff dff_A_jk3Igepg2_0(.din(n19350), .dout(n19347));
    jdff dff_A_A3snWA4u5_0(.din(n19353), .dout(n19350));
    jdff dff_A_8CYTgtUW9_0(.din(n19356), .dout(n19353));
    jdff dff_A_SWo3DVyA2_0(.din(G389), .dout(n19356));
    jdff dff_A_VxC4n2dU9_1(.din(n19362), .dout(n19359));
    jdff dff_A_QxBoCB4y1_1(.din(n19365), .dout(n19362));
    jdff dff_A_VgDuH2sX9_1(.din(G389), .dout(n19365));
    jdff dff_A_McdFHEj28_1(.din(n19371), .dout(n19368));
    jdff dff_A_SSYCyo4y7_1(.din(n19374), .dout(n19371));
    jdff dff_A_RU41QhYS4_1(.din(G389), .dout(n19374));
    jdff dff_A_BYPkcyG07_2(.din(n19380), .dout(n19377));
    jdff dff_A_SpExcGnA3_2(.din(n19383), .dout(n19380));
    jdff dff_A_xlgPmUFB1_2(.din(n19386), .dout(n19383));
    jdff dff_A_A8WUKmeI4_2(.din(G389), .dout(n19386));
    jdff dff_A_CID2Snx76_2(.din(G257), .dout(n19389));
    jdff dff_B_vQWbygcP6_1(.din(n5023), .dout(n19393));
    jdff dff_A_TJDdjxDN3_1(.din(n19398), .dout(n19395));
    jdff dff_A_Fq7oCxoN3_1(.din(n19405), .dout(n19398));
    jdff dff_A_pMW24VFp3_2(.din(n19405), .dout(n19401));
    jdff dff_B_5B0514A33_3(.din(n986), .dout(n19405));
    jdff dff_A_0HziCBUR3_0(.din(n19410), .dout(n19407));
    jdff dff_A_xtl1iMlQ9_0(.din(n19413), .dout(n19410));
    jdff dff_A_I4r5TiI65_0(.din(n19416), .dout(n19413));
    jdff dff_A_PRE9t4K11_0(.din(G400), .dout(n19416));
    jdff dff_A_CDgMUzjN4_1(.din(n19422), .dout(n19419));
    jdff dff_A_mGBU1vtR5_1(.din(n19425), .dout(n19422));
    jdff dff_A_BcsnzGcI1_1(.din(G400), .dout(n19425));
    jdff dff_B_ii3wpd5b0_1(.din(n5007), .dout(n19429));
    jdff dff_A_J1GBjRnw5_0(.din(G251), .dout(n19431));
    jdff dff_A_iW6HyRsz8_0(.din(G251), .dout(n19434));
    jdff dff_A_3HPeGmjr0_2(.din(G251), .dout(n19437));
    jdff dff_A_Xe8Fmw9H8_1(.din(n19443), .dout(n19440));
    jdff dff_A_poS3m5Qm4_1(.din(G400), .dout(n19443));
    jdff dff_A_AsvBBfPu7_2(.din(n19449), .dout(n19446));
    jdff dff_A_WrXyI5iu0_2(.din(n19452), .dout(n19449));
    jdff dff_A_v6NM0Qup3_2(.din(n19455), .dout(n19452));
    jdff dff_A_OVVhrC421_2(.din(G400), .dout(n19455));
    jdff dff_A_yKhhrmpy2_1(.din(G265), .dout(n19458));
    jdff dff_A_c5SsxF4r5_2(.din(G265), .dout(n19461));
    jdff dff_B_9eh08wkv9_1(.din(n4967), .dout(n19465));
    jdff dff_B_o8C3BcRH5_1(.din(n19465), .dout(n19468));
    jdff dff_A_YLF0ccXX5_0(.din(G281), .dout(n19470));
    jdff dff_A_NuzqmZ4V1_1(.din(n19476), .dout(n19473));
    jdff dff_A_zxckjhqV0_1(.din(n19486), .dout(n19476));
    jdff dff_A_vRi5HaW28_2(.din(n19482), .dout(n19479));
    jdff dff_A_oEkkQGhu1_2(.din(n19486), .dout(n19482));
    jdff dff_B_b9meJiND4_3(.din(n1166), .dout(n19486));
    jdff dff_A_3BW8hfJP5_0(.din(n19491), .dout(n19488));
    jdff dff_A_vZMHX8wm5_0(.din(n19494), .dout(n19491));
    jdff dff_A_9TpVP1lK2_0(.din(n19497), .dout(n19494));
    jdff dff_A_oxlsLqtp8_0(.din(G374), .dout(n19497));
    jdff dff_A_kYWSXtUk2_1(.din(n19503), .dout(n19500));
    jdff dff_A_MfbTLasS1_1(.din(n19506), .dout(n19503));
    jdff dff_A_pi6uTrMi7_1(.din(G374), .dout(n19506));
    jdff dff_A_8d7Ye7kU8_1(.din(n19512), .dout(n19509));
    jdff dff_A_D5okqryN3_1(.din(n19515), .dout(n19512));
    jdff dff_A_MbOpF8PG8_1(.din(G374), .dout(n19515));
    jdff dff_A_vRwjoFX78_2(.din(n19521), .dout(n19518));
    jdff dff_A_2PR6l5d35_2(.din(n19524), .dout(n19521));
    jdff dff_A_XbVAolyy7_2(.din(n19527), .dout(n19524));
    jdff dff_A_5g6MpCxj4_2(.din(G374), .dout(n19527));
    jdff dff_A_YoDwKxKM6_2(.din(G281), .dout(n19530));
    jdff dff_A_ObhXBezk2_0(.din(G242), .dout(n19533));
    jdff dff_A_vXPYLiIZ1_1(.din(G242), .dout(n19536));
    jdff dff_A_zeUXuxX64_2(.din(G242), .dout(n19539));
    jdff dff_B_J9zxAP4D0_1(.din(n4931), .dout(n19543));
    jdff dff_B_4fm55Zox3_1(.din(n19543), .dout(n19546));
    jdff dff_A_CCG8Zxt41_0(.din(G273), .dout(n19548));
    jdff dff_A_h7Jd0gJN0_1(.din(G251), .dout(n19551));
    jdff dff_A_DQGrjRHK8_2(.din(G251), .dout(n19554));
    jdff dff_A_AKrFKqE09_1(.din(n19560), .dout(n19557));
    jdff dff_A_fWW2UeFb7_1(.din(n19570), .dout(n19560));
    jdff dff_A_JRx1cu4J3_2(.din(n19566), .dout(n19563));
    jdff dff_A_r91G5d5d1_2(.din(n19570), .dout(n19566));
    jdff dff_B_2DsNOHuP7_3(.din(n940), .dout(n19570));
    jdff dff_A_ijT9kB0A1_0(.din(n19575), .dout(n19572));
    jdff dff_A_Wwvhte7V5_0(.din(n19578), .dout(n19575));
    jdff dff_A_El7HS5tF9_0(.din(G411), .dout(n19578));
    jdff dff_A_juiEJIiC2_0(.din(n19584), .dout(n19581));
    jdff dff_A_z5CTrU3b2_0(.din(n19587), .dout(n19584));
    jdff dff_A_MFdt46Gh2_0(.din(n19590), .dout(n19587));
    jdff dff_A_lge6Nse23_0(.din(G411), .dout(n19590));
    jdff dff_A_kMCUL8xc2_2(.din(n19596), .dout(n19593));
    jdff dff_A_QctWO7aU5_2(.din(n19599), .dout(n19596));
    jdff dff_A_HuQwAL7r3_2(.din(G411), .dout(n19599));
    jdff dff_A_AK5xYz0k8_1(.din(G273), .dout(n19602));
    jdff dff_A_4imqgMe79_2(.din(G273), .dout(n19605));
    jdff dff_A_OfhDr8Jr0_2(.din(G248), .dout(n19608));
    jdff dff_A_XL4AbLks6_1(.din(n19614), .dout(n19611));
    jdff dff_A_2ZuXrpe36_1(.din(n19617), .dout(n19614));
    jdff dff_A_t8w2e87r8_1(.din(n19620), .dout(n19617));
    jdff dff_A_oPNC0mPF0_1(.din(n19623), .dout(n19620));
    jdff dff_A_5yGfR4rj6_1(.din(n19626), .dout(n19623));
    jdff dff_A_MJ6Hvoij0_1(.din(n19629), .dout(n19626));
    jdff dff_A_RCJMwuVo0_1(.din(n19632), .dout(n19629));
    jdff dff_A_VBAUcQae1_1(.din(n19635), .dout(n19632));
    jdff dff_A_q49p95m61_1(.din(n19638), .dout(n19635));
    jdff dff_A_EXDpjo6W6_1(.din(n19641), .dout(n19638));
    jdff dff_A_QOcUvxSe8_1(.din(n19644), .dout(n19641));
    jdff dff_A_T1dFYe3G1_1(.din(n19647), .dout(n19644));
    jdff dff_A_rmSyudrV7_1(.din(n19650), .dout(n19647));
    jdff dff_A_sgr2C9MX6_1(.din(n19653), .dout(n19650));
    jdff dff_A_HEfhdYZv6_1(.din(n19656), .dout(n19653));
    jdff dff_A_vd0hohDx2_1(.din(n19659), .dout(n19656));
    jdff dff_A_CQbw284R5_1(.din(n1999), .dout(n19659));
    jdff dff_A_qc0WrT8J1_2(.din(n19665), .dout(n19662));
    jdff dff_A_oCgrTsBV9_2(.din(n19668), .dout(n19665));
    jdff dff_A_HIR4MtVn9_2(.din(n19671), .dout(n19668));
    jdff dff_A_KO4VY6Sp8_2(.din(n19674), .dout(n19671));
    jdff dff_A_40Z9CLjG2_2(.din(n19677), .dout(n19674));
    jdff dff_A_8QOhCgk58_2(.din(n19680), .dout(n19677));
    jdff dff_A_YfRbn58s9_2(.din(n19683), .dout(n19680));
    jdff dff_A_oRDUx95A7_2(.din(n1999), .dout(n19683));
    jdff dff_A_xo8H0iUw2_1(.din(n19689), .dout(n19686));
    jdff dff_A_pU6HVoYk6_1(.din(n19692), .dout(n19689));
    jdff dff_A_h14ZsECt1_1(.din(n19695), .dout(n19692));
    jdff dff_A_WSPSDGqZ9_1(.din(n1999), .dout(n19695));
    jdff dff_A_9q4aPqhS1_2(.din(n19701), .dout(n19698));
    jdff dff_A_yHz3fP6c9_2(.din(n19704), .dout(n19701));
    jdff dff_A_dsMB0Ji38_2(.din(n19707), .dout(n19704));
    jdff dff_A_MsncRhbx1_2(.din(n1999), .dout(n19707));
    jdff dff_A_2uW4Q9kK5_1(.din(n19713), .dout(n19710));
    jdff dff_A_lYHRuC0r7_1(.din(n1999), .dout(n19713));
    jdff dff_A_Aur4jt7Q5_2(.din(n19719), .dout(n19716));
    jdff dff_A_71ICoD9D2_2(.din(n19722), .dout(n19719));
    jdff dff_A_dbchnsP29_2(.din(n1999), .dout(n19722));
    jdff dff_A_VjbP3K595_0(.din(n19728), .dout(n19725));
    jdff dff_A_86b8CQdR3_0(.din(n19731), .dout(n19728));
    jdff dff_A_IEo8tGwN3_0(.din(n19734), .dout(n19731));
    jdff dff_A_mljz6IqM0_0(.din(n19737), .dout(n19734));
    jdff dff_A_piDFrEPc8_0(.din(G4091), .dout(n19737));
    jdff dff_A_EitXLudL1_0(.din(n19743), .dout(n19740));
    jdff dff_A_QnZl4vUa2_0(.din(n19746), .dout(n19743));
    jdff dff_A_9Xb9cIaV5_0(.din(n19749), .dout(n19746));
    jdff dff_A_0E3KASNc4_0(.din(n19752), .dout(n19749));
    jdff dff_A_ZZv3dkAw8_0(.din(n19755), .dout(n19752));
    jdff dff_A_tUwb5tTI9_0(.din(n19758), .dout(n19755));
    jdff dff_A_sQwWNgac7_0(.din(n19761), .dout(n19758));
    jdff dff_A_WS9eeEtU1_0(.din(G4091), .dout(n19761));
    jdff dff_A_9OEWljUK9_1(.din(n19767), .dout(n19764));
    jdff dff_A_Wo73ayXj5_1(.din(n19770), .dout(n19767));
    jdff dff_A_9HeyBpws5_1(.din(n19773), .dout(n19770));
    jdff dff_A_8LSCkkyj2_1(.din(n19776), .dout(n19773));
    jdff dff_A_PIJVGkZz1_1(.din(n19779), .dout(n19776));
    jdff dff_A_Ss8MEqmn8_1(.din(n19782), .dout(n19779));
    jdff dff_A_H1SsEM2h4_1(.din(G4091), .dout(n19782));
    jdff dff_A_9MtcZvZE4_1(.din(n19788), .dout(n19785));
    jdff dff_A_KKuVZUuQ7_1(.din(n19791), .dout(n19788));
    jdff dff_A_yQfGyEy12_1(.din(n19794), .dout(n19791));
    jdff dff_A_cf86T9NH3_1(.din(n19797), .dout(n19794));
    jdff dff_A_VjAtKayS5_1(.din(n19800), .dout(n19797));
    jdff dff_A_ajbuNz1y3_1(.din(n19803), .dout(n19800));
    jdff dff_A_Szs7ReQ35_1(.din(n19806), .dout(n19803));
    jdff dff_A_UGiFwJl39_1(.din(n19809), .dout(n19806));
    jdff dff_A_t3Q4ZoCk4_1(.din(n19812), .dout(n19809));
    jdff dff_A_5QgE2dt85_1(.din(n19815), .dout(n19812));
    jdff dff_A_2I9ItvmN3_1(.din(n19818), .dout(n19815));
    jdff dff_A_XdZlMQAp8_1(.din(n19821), .dout(n19818));
    jdff dff_A_ZsiNco8d4_1(.din(G4091), .dout(n19821));
    jdff dff_A_sV38P4L49_2(.din(n19827), .dout(n19824));
    jdff dff_A_o1bSZhtG4_2(.din(n19830), .dout(n19827));
    jdff dff_A_RxDwcOHl8_2(.din(n19833), .dout(n19830));
    jdff dff_A_4GsiOF2g8_2(.din(n19836), .dout(n19833));
    jdff dff_A_id7i98L30_2(.din(n19839), .dout(n19836));
    jdff dff_A_z11Eld5C5_2(.din(n19842), .dout(n19839));
    jdff dff_A_b6se461D7_2(.din(n19845), .dout(n19842));
    jdff dff_A_pFqduqXp0_2(.din(G4091), .dout(n19845));
    jdff dff_A_r7IPFdiu7_2(.din(n19851), .dout(n19848));
    jdff dff_A_ugPDC4sW7_2(.din(n19854), .dout(n19851));
    jdff dff_A_JW7ucBXq1_2(.din(n19857), .dout(n19854));
    jdff dff_A_orSiVrM64_2(.din(n19860), .dout(n19857));
    jdff dff_A_psOsMHOR2_2(.din(n19863), .dout(n19860));
    jdff dff_A_tQ5rBqIt1_2(.din(n19866), .dout(n19863));
    jdff dff_A_TQCfDaYJ3_2(.din(n19869), .dout(n19866));
    jdff dff_A_WV4ki3Zp1_2(.din(n19872), .dout(n19869));
    jdff dff_A_hNALHbFE6_2(.din(n19875), .dout(n19872));
    jdff dff_A_YnuYCGgS8_2(.din(n19878), .dout(n19875));
    jdff dff_A_tWgS3oAK1_2(.din(n19881), .dout(n19878));
    jdff dff_A_WsPtK1r61_2(.din(n19884), .dout(n19881));
    jdff dff_A_Tvm6nn3e3_2(.din(n19887), .dout(n19884));
    jdff dff_A_DnTYD3nX1_2(.din(n19890), .dout(n19887));
    jdff dff_A_fCJhd0fm9_2(.din(n19893), .dout(n19890));
    jdff dff_A_UJ2Znemh6_2(.din(n19896), .dout(n19893));
    jdff dff_A_Ws7c9QGw6_2(.din(n19899), .dout(n19896));
    jdff dff_A_r7lXwKxe0_2(.din(n19902), .dout(n19899));
    jdff dff_A_8AcuioY74_2(.din(n19905), .dout(n19902));
    jdff dff_A_4gOJRDdD0_2(.din(G4092), .dout(n19905));
    jdff dff_A_QPoL2Yr86_1(.din(G4092), .dout(n19908));
    jdff dff_A_WSqycTFI7_0(.din(n19914), .dout(n19911));
    jdff dff_A_uUSEqkrO9_0(.din(n19917), .dout(n19914));
    jdff dff_A_ON0sg6aB4_0(.din(n19920), .dout(n19917));
    jdff dff_A_4uUDOd8n9_0(.din(n19923), .dout(n19920));
    jdff dff_A_ok1mW5CE9_0(.din(n19926), .dout(n19923));
    jdff dff_A_Qx3w1VQI2_0(.din(n19929), .dout(n19926));
    jdff dff_A_8f1KVLOG8_0(.din(n19932), .dout(n19929));
    jdff dff_A_SMf7Agkr3_0(.din(n19935), .dout(n19932));
    jdff dff_A_n88UjXSt9_0(.din(n19938), .dout(n19935));
    jdff dff_A_4EMrDtKz7_0(.din(n19941), .dout(n19938));
    jdff dff_A_2ZojMmEh2_0(.din(n19944), .dout(n19941));
    jdff dff_A_OYIlsWXH8_0(.din(n19947), .dout(n19944));
    jdff dff_A_qFgT65Bj9_0(.din(n19950), .dout(n19947));
    jdff dff_A_XCvCTKxb7_0(.din(n19953), .dout(n19950));
    jdff dff_A_SKWies1N4_0(.din(n2978), .dout(n19953));
    jdff dff_A_u3Idcy3m6_2(.din(n19959), .dout(n19956));
    jdff dff_A_LA10yz5M3_2(.din(n19962), .dout(n19959));
    jdff dff_A_TlxeCcEY4_2(.din(n19965), .dout(n19962));
    jdff dff_A_QQO0Bdfn3_2(.din(n19968), .dout(n19965));
    jdff dff_A_bSPJPTBF8_2(.din(n19971), .dout(n19968));
    jdff dff_A_EGyJJntq3_2(.din(n19974), .dout(n19971));
    jdff dff_A_D5C9xmcl9_2(.din(n19977), .dout(n19974));
    jdff dff_A_OQJO4pMg6_2(.din(n19980), .dout(n19977));
    jdff dff_A_zcNQ3ys02_2(.din(n19983), .dout(n19980));
    jdff dff_A_mZ86McBp3_2(.din(n2978), .dout(n19983));
    jdff dff_A_kSfNaV7k4_1(.din(n19989), .dout(n19986));
    jdff dff_A_XCW97tO20_1(.din(n19992), .dout(n19989));
    jdff dff_A_dsynUTGi1_1(.din(n19995), .dout(n19992));
    jdff dff_A_oLJktYkX3_1(.din(n19998), .dout(n19995));
    jdff dff_A_OhuHp5ts4_1(.din(n20001), .dout(n19998));
    jdff dff_A_dnfSHvyF5_1(.din(n20004), .dout(n20001));
    jdff dff_A_Bh0PukLk2_1(.din(n20007), .dout(n20004));
    jdff dff_A_Q7GQe5kG7_1(.din(n20010), .dout(n20007));
    jdff dff_A_VJp9CNGQ7_1(.din(n20013), .dout(n20010));
    jdff dff_A_Npfoxvkr2_1(.din(n20016), .dout(n20013));
    jdff dff_A_RRf0z1JV7_1(.din(n20019), .dout(n20016));
    jdff dff_A_0LDNOHWG8_1(.din(n20022), .dout(n20019));
    jdff dff_A_pjQgGHN08_1(.din(n20025), .dout(n20022));
    jdff dff_A_XJr2CE7J8_1(.din(n20028), .dout(n20025));
    jdff dff_A_wayGqTb63_1(.din(n20031), .dout(n20028));
    jdff dff_A_DYHgFZ441_1(.din(n20034), .dout(n20031));
    jdff dff_A_52KHvoTS2_1(.din(n20037), .dout(n20034));
    jdff dff_A_WR26FZwb7_1(.din(n20040), .dout(n20037));
    jdff dff_A_xftwfBFJ9_1(.din(n20043), .dout(n20040));
    jdff dff_A_QDnQbt1F5_1(.din(n20046), .dout(n20043));
    jdff dff_A_pQ3HAkyF6_1(.din(n2978), .dout(n20046));
    jdff dff_A_SIxGBBAz0_2(.din(n20052), .dout(n20049));
    jdff dff_A_oR8Ojy7Q8_2(.din(n20055), .dout(n20052));
    jdff dff_A_Fs10dkLd6_2(.din(n20058), .dout(n20055));
    jdff dff_A_pO8CWy865_2(.din(n20061), .dout(n20058));
    jdff dff_A_mP8DDIcz7_2(.din(n20064), .dout(n20061));
    jdff dff_A_rdAFcOJ67_2(.din(n20067), .dout(n20064));
    jdff dff_A_sTvDPdlT3_2(.din(n20070), .dout(n20067));
    jdff dff_A_bHA0pX3V9_2(.din(n20073), .dout(n20070));
    jdff dff_A_ZxqKzhHM7_2(.din(n20076), .dout(n20073));
    jdff dff_A_5LGF4Llh5_2(.din(n20079), .dout(n20076));
    jdff dff_A_YuYIoP734_2(.din(n20082), .dout(n20079));
    jdff dff_A_RMrA0vc58_2(.din(n20085), .dout(n20082));
    jdff dff_A_1DDlXiSl7_2(.din(n20088), .dout(n20085));
    jdff dff_A_A0wXchy67_2(.din(n20091), .dout(n20088));
    jdff dff_A_axxn571j7_2(.din(n20094), .dout(n20091));
    jdff dff_A_fizGF83e2_2(.din(n20097), .dout(n20094));
    jdff dff_A_7exSQ6oc8_2(.din(n20100), .dout(n20097));
    jdff dff_A_Klt8O5nc0_2(.din(n20103), .dout(n20100));
    jdff dff_A_AwGANxKm8_2(.din(n20106), .dout(n20103));
    jdff dff_A_SwhyDRds8_2(.din(n2978), .dout(n20106));
    jdff dff_A_joNpa7pj5_1(.din(n20112), .dout(n20109));
    jdff dff_A_IwgFjkYh3_1(.din(n20115), .dout(n20112));
    jdff dff_A_KLZFKEtw2_1(.din(n20118), .dout(n20115));
    jdff dff_A_7FxgQzyS8_1(.din(n20121), .dout(n20118));
    jdff dff_A_mKKPOxLH8_1(.din(n20124), .dout(n20121));
    jdff dff_A_eFGPnXsz7_1(.din(n20127), .dout(n20124));
    jdff dff_A_EHMk3NIn7_1(.din(n20130), .dout(n20127));
    jdff dff_A_NklZwVqI4_1(.din(n20133), .dout(n20130));
    jdff dff_A_Sv95TVcw6_1(.din(n20136), .dout(n20133));
    jdff dff_A_PKwUAUwU8_1(.din(n20139), .dout(n20136));
    jdff dff_A_oUP31tfa2_1(.din(n20142), .dout(n20139));
    jdff dff_A_MVYqPbwh5_1(.din(n20145), .dout(n20142));
    jdff dff_A_CRBbVg4z5_1(.din(n20148), .dout(n20145));
    jdff dff_A_8BtsdIM15_1(.din(n20151), .dout(n20148));
    jdff dff_A_vH45RwE30_1(.din(n20154), .dout(n20151));
    jdff dff_A_CBJv59lI3_1(.din(n20157), .dout(n20154));
    jdff dff_A_fDL2Gcz20_1(.din(n20160), .dout(n20157));
    jdff dff_A_b1Z1GqIh7_1(.din(n2978), .dout(n20160));
    jdff dff_A_gZloFhOf3_2(.din(n20166), .dout(n20163));
    jdff dff_A_Lu9EV3RW3_2(.din(n20169), .dout(n20166));
    jdff dff_A_jNxfeHUK6_2(.din(n20172), .dout(n20169));
    jdff dff_A_CDcBIiOV7_2(.din(n20175), .dout(n20172));
    jdff dff_A_HW3Sb6ig8_2(.din(n20178), .dout(n20175));
    jdff dff_A_C9YfbesS1_2(.din(n20181), .dout(n20178));
    jdff dff_A_pyMCgMEp8_2(.din(n20184), .dout(n20181));
    jdff dff_A_da5ylVH45_2(.din(n20187), .dout(n20184));
    jdff dff_A_9BWh89Fn8_2(.din(n20190), .dout(n20187));
    jdff dff_A_PoY3Yy488_2(.din(n20193), .dout(n20190));
    jdff dff_A_wtsjZLC43_2(.din(n2978), .dout(n20193));
    jdff dff_A_lvhsygkr0_1(.din(n20199), .dout(n20196));
    jdff dff_A_nGbJspLH0_1(.din(n20202), .dout(n20199));
    jdff dff_A_zMCP0Xa69_1(.din(n20205), .dout(n20202));
    jdff dff_A_Mtb30mf10_1(.din(n20208), .dout(n20205));
    jdff dff_A_7z7cGEbk7_1(.din(n20211), .dout(n20208));
    jdff dff_A_LLipclX71_1(.din(n20214), .dout(n20211));
    jdff dff_A_sXUPwNmt9_1(.din(n20217), .dout(n20214));
    jdff dff_A_GUx2y2KX8_1(.din(n20220), .dout(n20217));
    jdff dff_A_KCA2LkGM5_1(.din(G1691), .dout(n20220));
    jdff dff_B_JFNhjRj26_2(.din(n5676), .dout(n20224));
    jdff dff_B_SHjTvCFN8_2(.din(n20224), .dout(n20227));
    jdff dff_A_NrHeVJaU2_1(.din(n20232), .dout(n20229));
    jdff dff_A_OYuBxBoI3_1(.din(n20235), .dout(n20232));
    jdff dff_A_83w313hf4_1(.din(n20238), .dout(n20235));
    jdff dff_A_uq3IpMya7_1(.din(n20241), .dout(n20238));
    jdff dff_A_PndnQEq71_1(.din(n20244), .dout(n20241));
    jdff dff_A_tt66UUE16_1(.din(n20247), .dout(n20244));
    jdff dff_A_MkNfVwnp9_1(.din(n20250), .dout(n20247));
    jdff dff_A_6CU7N1Vx3_1(.din(n20253), .dout(n20250));
    jdff dff_A_HL2V6y215_1(.din(n20256), .dout(n20253));
    jdff dff_A_MgmqeuPb5_1(.din(n20259), .dout(n20256));
    jdff dff_A_R894gWeW2_1(.din(n20262), .dout(n20259));
    jdff dff_A_xVXb5A5Y1_1(.din(n20265), .dout(n20262));
    jdff dff_A_bvIW5vGo3_1(.din(n20268), .dout(n20265));
    jdff dff_A_aHrjlshB3_1(.din(n20271), .dout(n20268));
    jdff dff_A_n8pSpgXP7_1(.din(n20274), .dout(n20271));
    jdff dff_A_WI9PiHta0_1(.din(n20277), .dout(n20274));
    jdff dff_A_K8lD1TQj4_1(.din(n20280), .dout(n20277));
    jdff dff_A_LbbRRbec4_1(.din(n20283), .dout(n20280));
    jdff dff_A_veYxSZ2n8_1(.din(n20286), .dout(n20283));
    jdff dff_A_IR6oyroZ0_1(.din(n20289), .dout(n20286));
    jdff dff_A_o6R8sHul4_1(.din(n20292), .dout(n20289));
    jdff dff_A_rm69yGQw1_1(.din(n20295), .dout(n20292));
    jdff dff_A_PuJrd79y3_1(.din(G1694), .dout(n20295));
    jdff dff_A_dgGMwTgw5_2(.din(G1694), .dout(n20298));
    jdff dff_A_jez6q3ck6_0(.din(n20304), .dout(n20301));
    jdff dff_A_Y5Htbw501_0(.din(n20307), .dout(n20304));
    jdff dff_A_y1XNu93O5_0(.din(n20310), .dout(n20307));
    jdff dff_A_nuFK7bXb4_0(.din(n20313), .dout(n20310));
    jdff dff_A_EupK70Ep0_0(.din(n20316), .dout(n20313));
    jdff dff_A_lFRbiMll2_0(.din(n20319), .dout(n20316));
    jdff dff_A_rffl1DUk7_0(.din(n20322), .dout(n20319));
    jdff dff_A_jg5l5pMu3_0(.din(n20325), .dout(n20322));
    jdff dff_A_uU8WhNG28_0(.din(n20328), .dout(n20325));
    jdff dff_A_hKfi0Hnm4_0(.din(n20331), .dout(n20328));
    jdff dff_A_lmAqRxtF5_0(.din(n20334), .dout(n20331));
    jdff dff_A_nGpldJDP8_0(.din(n20337), .dout(n20334));
    jdff dff_A_OSok7hQx6_0(.din(n20340), .dout(n20337));
    jdff dff_A_eNq6EuQo6_0(.din(G1691), .dout(n20340));
    jdff dff_A_ZJRvuEij9_1(.din(n20346), .dout(n20343));
    jdff dff_A_DPFh9Ds93_1(.din(n20349), .dout(n20346));
    jdff dff_A_cnEbxqi33_1(.din(n20352), .dout(n20349));
    jdff dff_A_wKY5CZ829_1(.din(n20355), .dout(n20352));
    jdff dff_A_tSDqsGMI2_1(.din(n20358), .dout(n20355));
    jdff dff_A_fgD7Vqk01_1(.din(n20361), .dout(n20358));
    jdff dff_A_eqb7eVTU8_1(.din(n20364), .dout(n20361));
    jdff dff_A_6WBwahvX6_1(.din(n20367), .dout(n20364));
    jdff dff_A_nDzZ8UwB1_1(.din(n20370), .dout(n20367));
    jdff dff_A_51fD4GFb3_1(.din(n20373), .dout(n20370));
    jdff dff_A_MORzu4mx0_1(.din(n20376), .dout(n20373));
    jdff dff_A_9MzmqfIV6_1(.din(n20379), .dout(n20376));
    jdff dff_A_6UCJrQ7E3_1(.din(n20382), .dout(n20379));
    jdff dff_A_c1qCztz99_1(.din(n20385), .dout(n20382));
    jdff dff_A_Al4YqERy7_1(.din(n20388), .dout(n20385));
    jdff dff_A_XLZ3R2fU3_1(.din(G1691), .dout(n20388));
    jdff dff_A_ZtOT0hLB6_2(.din(n20394), .dout(n20391));
    jdff dff_A_pel3Qd872_2(.din(n20397), .dout(n20394));
    jdff dff_A_bqdsjcwZ5_2(.din(n20400), .dout(n20397));
    jdff dff_A_RF67uqnd0_2(.din(n20403), .dout(n20400));
    jdff dff_A_sLk00SdQ3_2(.din(n20406), .dout(n20403));
    jdff dff_A_oTAhzqlh9_2(.din(n20409), .dout(n20406));
    jdff dff_A_5DeqOacz4_2(.din(n20412), .dout(n20409));
    jdff dff_A_ApLMwgYC1_2(.din(n20415), .dout(n20412));
    jdff dff_A_r9sl2ikc0_2(.din(n20418), .dout(n20415));
    jdff dff_A_tnokxD7K6_2(.din(n20421), .dout(n20418));
    jdff dff_A_PKYjso3T5_2(.din(n20424), .dout(n20421));
    jdff dff_A_aETqB8B26_2(.din(n20427), .dout(n20424));
    jdff dff_A_XFia1uVj0_2(.din(n20430), .dout(n20427));
    jdff dff_A_e2Ael8mC2_2(.din(n20433), .dout(n20430));
    jdff dff_A_WtGp5k6j4_2(.din(n20436), .dout(n20433));
    jdff dff_A_NibZ94Xm9_2(.din(n20439), .dout(n20436));
    jdff dff_A_iq4YHuwO1_2(.din(n20442), .dout(n20439));
    jdff dff_A_GcuuUpUv0_2(.din(n20445), .dout(n20442));
    jdff dff_A_lnW7Jwxq5_2(.din(n20448), .dout(n20445));
    jdff dff_A_bf8uZ9ug9_2(.din(n20451), .dout(n20448));
    jdff dff_A_nfyhVbYY1_2(.din(n20454), .dout(n20451));
    jdff dff_A_DEUdClEX8_2(.din(G1691), .dout(n20454));
    jdff dff_A_uOHIpPs64_1(.din(n20460), .dout(n20457));
    jdff dff_A_Pe0dDGyj5_1(.din(n20463), .dout(n20460));
    jdff dff_A_RAB56aaU4_1(.din(n20466), .dout(n20463));
    jdff dff_A_HUKCjav54_1(.din(n20469), .dout(n20466));
    jdff dff_A_Rb6g0GMP0_1(.din(n20472), .dout(n20469));
    jdff dff_A_UOAqTRwi0_1(.din(n20475), .dout(n20472));
    jdff dff_A_RqlN2u1v4_1(.din(n20478), .dout(n20475));
    jdff dff_A_05hehML31_1(.din(n20481), .dout(n20478));
    jdff dff_A_IjBL1HG98_1(.din(n20484), .dout(n20481));
    jdff dff_A_lboOwYLZ3_1(.din(n20487), .dout(n20484));
    jdff dff_A_qlbNgzLd4_1(.din(n20490), .dout(n20487));
    jdff dff_A_ivzypPC02_1(.din(n20493), .dout(n20490));
    jdff dff_A_glX40HsQ0_1(.din(n20496), .dout(n20493));
    jdff dff_A_MBUqYFrl2_1(.din(n20499), .dout(n20496));
    jdff dff_A_wbaxU3AM2_1(.din(n20502), .dout(n20499));
    jdff dff_A_xAhcRo9w8_1(.din(n20505), .dout(n20502));
    jdff dff_A_RX3Z8UeR4_1(.din(n20508), .dout(n20505));
    jdff dff_A_KJeWS4oe5_1(.din(n20511), .dout(n20508));
    jdff dff_A_6aehFRuv9_1(.din(G1691), .dout(n20511));
    jdff dff_A_dMd4Dplq1_2(.din(n20517), .dout(n20514));
    jdff dff_A_4GLrp35o8_2(.din(n20520), .dout(n20517));
    jdff dff_A_WuFYFDj19_2(.din(n20523), .dout(n20520));
    jdff dff_A_5zI5gduW9_2(.din(n20526), .dout(n20523));
    jdff dff_A_JcBH96rA1_2(.din(n20529), .dout(n20526));
    jdff dff_A_RwUuL03E9_2(.din(n20532), .dout(n20529));
    jdff dff_A_qSKoB0l20_2(.din(n20535), .dout(n20532));
    jdff dff_A_JzZxz98o0_2(.din(n20538), .dout(n20535));
    jdff dff_A_KFrZBu1F1_2(.din(n20541), .dout(n20538));
    jdff dff_A_0RcGyH1M4_2(.din(n20544), .dout(n20541));
    jdff dff_A_klkUp8ao9_2(.din(n20547), .dout(n20544));
    jdff dff_A_dT8Ia2OZ0_2(.din(n20550), .dout(n20547));
    jdff dff_A_vGHTfhyW9_2(.din(G1691), .dout(n20550));
    jdff dff_B_AzGMDA8y8_2(.din(n5666), .dout(n20554));
    jdff dff_B_uy03LviU8_2(.din(n5663), .dout(n20557));
    jdff dff_B_8e51ZPui5_2(.din(n20557), .dout(n20560));
    jdff dff_B_UI1HZQrx3_2(.din(n20560), .dout(n20563));
    jdff dff_B_ONbC3eCq1_2(.din(n20563), .dout(n20566));
    jdff dff_B_lfDjGvPZ0_2(.din(n20566), .dout(n20569));
    jdff dff_B_CMs9GZ1y0_2(.din(n20569), .dout(n20572));
    jdff dff_B_4fPtujk65_2(.din(n20572), .dout(n20575));
    jdff dff_B_mWon9R7R9_2(.din(n20575), .dout(n20578));
    jdff dff_B_HuA5otXH4_2(.din(n20578), .dout(n20581));
    jdff dff_B_31jyz91C5_2(.din(n20581), .dout(n20584));
    jdff dff_B_Kj3JMYLO7_2(.din(n20584), .dout(n20587));
    jdff dff_B_rt2susp59_2(.din(n20587), .dout(n20590));
    jdff dff_B_moXigPB47_2(.din(n20590), .dout(n20593));
    jdff dff_B_Ey2tPuqD6_2(.din(n20593), .dout(n20596));
    jdff dff_B_7tL7QzxS7_2(.din(n20596), .dout(n20599));
    jdff dff_B_k5cSsR3t0_2(.din(n20599), .dout(n20602));
    jdff dff_B_4755z2Hn7_2(.din(n20602), .dout(n20605));
    jdff dff_B_s9yo5N0r9_2(.din(n20605), .dout(n20608));
    jdff dff_B_OFXG6fSg7_2(.din(n20608), .dout(n20611));
    jdff dff_B_CFnvvsaX4_2(.din(n20611), .dout(n20614));
    jdff dff_B_wk8eK7oI1_2(.din(n20614), .dout(n20617));
    jdff dff_B_VoyoSs4I0_2(.din(n20617), .dout(n20620));
    jdff dff_B_NYN7OKw15_2(.din(n20620), .dout(n20623));
    jdff dff_B_4ld0KiXW7_2(.din(n20623), .dout(n20626));
    jdff dff_B_CxtvxXxF4_2(.din(n20626), .dout(n20629));
    jdff dff_B_ZhlFiBiX3_2(.din(n20629), .dout(n20632));
    jdff dff_A_PWzSKAnh2_2(.din(n20637), .dout(n20634));
    jdff dff_A_pJu6TLUw5_2(.din(n20640), .dout(n20637));
    jdff dff_A_VaawTq0Y3_2(.din(n20643), .dout(n20640));
    jdff dff_A_yOYMrknm3_2(.din(n20646), .dout(n20643));
    jdff dff_A_s6wrYOsC1_2(.din(n20649), .dout(n20646));
    jdff dff_A_LsHyNQB36_2(.din(n20652), .dout(n20649));
    jdff dff_A_48j3K6HD4_2(.din(n20655), .dout(n20652));
    jdff dff_A_eqg8PPEo6_2(.din(n20658), .dout(n20655));
    jdff dff_A_ELQkdxmX1_2(.din(n20661), .dout(n20658));
    jdff dff_A_uuq7jWJm9_2(.din(n20664), .dout(n20661));
    jdff dff_A_LBfUyJGt2_2(.din(n20667), .dout(n20664));
    jdff dff_A_vnLBMEmj1_2(.din(n20670), .dout(n20667));
    jdff dff_A_6VPhDO5v1_2(.din(n20673), .dout(n20670));
    jdff dff_A_RMshaW478_2(.din(n20676), .dout(n20673));
    jdff dff_A_ZSAPFrF88_2(.din(n20679), .dout(n20676));
    jdff dff_A_vKJ96aS84_2(.din(n20682), .dout(n20679));
    jdff dff_A_xRPTxXmC9_2(.din(n20685), .dout(n20682));
    jdff dff_A_Io6h3bx43_2(.din(n20688), .dout(n20685));
    jdff dff_A_B9ujESKV2_2(.din(n20691), .dout(n20688));
    jdff dff_A_B02DsWh05_2(.din(n20694), .dout(n20691));
    jdff dff_A_C0zyaOhS4_2(.din(n20697), .dout(n20694));
    jdff dff_A_7KLxEBCn3_2(.din(n20700), .dout(n20697));
    jdff dff_A_6QicL7n99_2(.din(n20703), .dout(n20700));
    jdff dff_A_tdkmqNYI7_2(.din(G137), .dout(n20703));
    jdff dff_A_JaX8JiOJ9_0(.din(n20709), .dout(n20706));
    jdff dff_A_DWFiqVPp2_0(.din(n20712), .dout(n20709));
    jdff dff_A_4Y8E3njp6_0(.din(n20715), .dout(n20712));
    jdff dff_A_uTKog0qp3_0(.din(n20718), .dout(n20715));
    jdff dff_A_Yl6sBJFe7_0(.din(n20721), .dout(n20718));
    jdff dff_A_vrU1h5q76_0(.din(n20724), .dout(n20721));
    jdff dff_A_6h6MoGTq4_0(.din(n20727), .dout(n20724));
    jdff dff_A_3sz47knn2_0(.din(n20730), .dout(n20727));
    jdff dff_A_5Z5PhRWw2_0(.din(n20733), .dout(n20730));
    jdff dff_A_4qQJtJNU1_0(.din(n20736), .dout(n20733));
    jdff dff_A_qxrKAmvh1_0(.din(n20739), .dout(n20736));
    jdff dff_A_8SFuhkZz4_0(.din(n20742), .dout(n20739));
    jdff dff_A_fLt2uriD4_0(.din(n20745), .dout(n20742));
    jdff dff_A_XYpH9AIa3_0(.din(n20748), .dout(n20745));
    jdff dff_A_8HvueTtx2_0(.din(n20751), .dout(n20748));
    jdff dff_A_1IJ4gebr6_0(.din(n20754), .dout(n20751));
    jdff dff_A_yOntMPx73_0(.din(G137), .dout(n20754));
    jdff dff_A_PgPS7vHF7_1(.din(n20760), .dout(n20757));
    jdff dff_A_U7LGI2NW6_1(.din(n20763), .dout(n20760));
    jdff dff_A_5H0sIIw53_1(.din(n20766), .dout(n20763));
    jdff dff_A_vR1YJq4y5_1(.din(n20769), .dout(n20766));
    jdff dff_A_E6SiKNQJ1_1(.din(n20772), .dout(n20769));
    jdff dff_A_Dnlmsim40_1(.din(n20775), .dout(n20772));
    jdff dff_A_IfxHcgWw0_1(.din(n20778), .dout(n20775));
    jdff dff_A_CS1XUDc44_1(.din(n20781), .dout(n20778));
    jdff dff_A_lgskrCNj6_1(.din(n20784), .dout(n20781));
    jdff dff_A_TaMCCUBL4_1(.din(n20787), .dout(n20784));
    jdff dff_A_cLxrOEJU8_1(.din(n20790), .dout(n20787));
    jdff dff_A_BhUrfjsT4_1(.din(n20793), .dout(n20790));
    jdff dff_A_MyMfKrmE2_1(.din(n20796), .dout(n20793));
    jdff dff_A_UikOBbBR2_1(.din(n20799), .dout(n20796));
    jdff dff_A_fEh8IIwQ7_1(.din(G137), .dout(n20799));
    jdff dff_A_3qesbko21_1(.din(n5756), .dout(n20802));
    jdff dff_A_rZMUeqtT1_0(.din(n20802), .dout(n20805));
    jdff dff_A_2xZl2LHc0_0(.din(n20805), .dout(n20808));
    jdff dff_A_o4hKRHkh8_0(.din(n20808), .dout(n20811));
    jdff dff_A_fbl2CEZY5_0(.din(n20811), .dout(n20814));
    jdff dff_A_LmrBxr9C2_0(.din(n20814), .dout(n20817));
    jdff dff_A_DOIi9s5f9_0(.din(n20817), .dout(n20820));
    jdff dff_A_9iYeXxQm9_0(.din(n20820), .dout(n20823));
    jdff dff_A_DQTCx7PV6_0(.din(n20823), .dout(n20826));
    jdff dff_A_9pd7nHgI1_0(.din(n20826), .dout(n20829));
    jdff dff_A_U7Vz4sXe9_0(.din(n20829), .dout(n20832));
    jdff dff_A_Rk1zU4oN8_0(.din(n20832), .dout(n20835));
    jdff dff_A_8EcYE1yi1_0(.din(n20835), .dout(n20838));
    jdff dff_A_kXzompdx0_0(.din(n20838), .dout(n20841));
    jdff dff_A_N1qdQRdK4_0(.din(n20841), .dout(n20844));
    jdff dff_A_UP7Tw7xo6_0(.din(n20844), .dout(n20847));
    jdff dff_A_4BObyJuZ0_0(.din(n20847), .dout(n20850));
    jdff dff_A_9IdfYSln5_0(.din(n20850), .dout(n20853));
    jdff dff_A_jdP6U8b07_0(.din(n20853), .dout(n20856));
    jdff dff_A_kZqzrERF1_0(.din(n20856), .dout(n20859));
    jdff dff_A_JS09NjOF6_0(.din(n20859), .dout(n20862));
    jdff dff_A_izbnWL9K6_0(.din(n20862), .dout(n20865));
    jdff dff_A_WgQjA4mu7_0(.din(n20865), .dout(n20868));
    jdff dff_A_5kcqco9f3_0(.din(n20868), .dout(n20871));
    jdff dff_A_PW2Da1iG2_0(.din(n20871), .dout(n20874));
    jdff dff_A_JFty1vSw1_0(.din(n20874), .dout(n20877));
    jdff dff_A_Kk4Jsm8Y5_0(.din(n20877), .dout(G144));
    jdff dff_A_k5hS1sGE3_1(.din(n5759), .dout(n20883));
    jdff dff_A_8uWlESyb2_0(.din(n20883), .dout(n20886));
    jdff dff_A_ZxbXG1ZX7_0(.din(n20886), .dout(n20889));
    jdff dff_A_XUqMXgsB7_0(.din(n20889), .dout(n20892));
    jdff dff_A_Ke4YvWgH0_0(.din(n20892), .dout(n20895));
    jdff dff_A_jyng7xC70_0(.din(n20895), .dout(n20898));
    jdff dff_A_Y917uZt44_0(.din(n20898), .dout(n20901));
    jdff dff_A_NC2HOdeJ7_0(.din(n20901), .dout(n20904));
    jdff dff_A_4a5o1oev5_0(.din(n20904), .dout(n20907));
    jdff dff_A_cYgNx4oo5_0(.din(n20907), .dout(n20910));
    jdff dff_A_b7edN0jj3_0(.din(n20910), .dout(n20913));
    jdff dff_A_XuUOAamh3_0(.din(n20913), .dout(n20916));
    jdff dff_A_mZbRYjb50_0(.din(n20916), .dout(n20919));
    jdff dff_A_PbfIIqdM0_0(.din(n20919), .dout(n20922));
    jdff dff_A_7pT2pHSk2_0(.din(n20922), .dout(n20925));
    jdff dff_A_ROW0QVMA0_0(.din(n20925), .dout(n20928));
    jdff dff_A_6WUchvPs2_0(.din(n20928), .dout(n20931));
    jdff dff_A_P1xrhZVX1_0(.din(n20931), .dout(n20934));
    jdff dff_A_q4ZuV6WA7_0(.din(n20934), .dout(n20937));
    jdff dff_A_kKeVad1S9_0(.din(n20937), .dout(n20940));
    jdff dff_A_IevzEcxt4_0(.din(n20940), .dout(n20943));
    jdff dff_A_TeifZMw32_0(.din(n20943), .dout(n20946));
    jdff dff_A_Xm0W3xgQ8_0(.din(n20946), .dout(n20949));
    jdff dff_A_vjGNUgun3_0(.din(n20949), .dout(n20952));
    jdff dff_A_xCMijMMy9_0(.din(n20952), .dout(n20955));
    jdff dff_A_6VqqoTRR5_0(.din(n20955), .dout(n20958));
    jdff dff_A_bVoxBf3X7_0(.din(n20958), .dout(G298));
    jdff dff_A_d6kwjLVZ0_1(.din(n5762), .dout(n20964));
    jdff dff_A_Zs4FhmDx9_0(.din(n20964), .dout(n20967));
    jdff dff_A_udvjerb55_0(.din(n20967), .dout(n20970));
    jdff dff_A_jHunwUCV1_0(.din(n20970), .dout(n20973));
    jdff dff_A_ojg6VGAY8_0(.din(n20973), .dout(n20976));
    jdff dff_A_twwtg2867_0(.din(n20976), .dout(n20979));
    jdff dff_A_QQUPyo6B3_0(.din(n20979), .dout(n20982));
    jdff dff_A_aKnkfTMm3_0(.din(n20982), .dout(n20985));
    jdff dff_A_griBH8TH1_0(.din(n20985), .dout(n20988));
    jdff dff_A_WkKUe34a9_0(.din(n20988), .dout(n20991));
    jdff dff_A_cUFSCdBl4_0(.din(n20991), .dout(n20994));
    jdff dff_A_jV4oyZOf2_0(.din(n20994), .dout(n20997));
    jdff dff_A_KWia5jN18_0(.din(n20997), .dout(n21000));
    jdff dff_A_FV4HJGny4_0(.din(n21000), .dout(n21003));
    jdff dff_A_NkiHE9p90_0(.din(n21003), .dout(n21006));
    jdff dff_A_hD5vSv531_0(.din(n21006), .dout(n21009));
    jdff dff_A_mLW3L2zd3_0(.din(n21009), .dout(n21012));
    jdff dff_A_gTUaK7PN3_0(.din(n21012), .dout(n21015));
    jdff dff_A_9GUhU2QS7_0(.din(n21015), .dout(n21018));
    jdff dff_A_lpMKehaN0_0(.din(n21018), .dout(n21021));
    jdff dff_A_tLHd8NGO8_0(.din(n21021), .dout(n21024));
    jdff dff_A_osog69XA8_0(.din(n21024), .dout(n21027));
    jdff dff_A_8Y1H6pcH4_0(.din(n21027), .dout(n21030));
    jdff dff_A_8MYk7QEc1_0(.din(n21030), .dout(n21033));
    jdff dff_A_THwqZlsa1_0(.din(n21033), .dout(n21036));
    jdff dff_A_fzLeF5Br9_0(.din(n21036), .dout(n21039));
    jdff dff_A_JfqOrBRk2_0(.din(n21039), .dout(G973));
    jdff dff_A_VHpW1ILW7_1(.din(n303), .dout(n21045));
    jdff dff_A_0EdNBvdh9_0(.din(n21045), .dout(n21048));
    jdff dff_A_D4OkyQ4G9_0(.din(n21048), .dout(n21051));
    jdff dff_A_QfKA9iXQ7_0(.din(n21051), .dout(n21054));
    jdff dff_A_wOhFogC16_0(.din(n21054), .dout(n21057));
    jdff dff_A_UGs0r12P4_0(.din(n21057), .dout(n21060));
    jdff dff_A_zaSpRqku1_0(.din(n21060), .dout(n21063));
    jdff dff_A_dbPsrNvz1_0(.din(n21063), .dout(n21066));
    jdff dff_A_HoAwRdxX7_0(.din(n21066), .dout(n21069));
    jdff dff_A_8QFTlGAL7_0(.din(n21069), .dout(n21072));
    jdff dff_A_9jFSz56R8_0(.din(n21072), .dout(n21075));
    jdff dff_A_urHNbyaD5_0(.din(n21075), .dout(n21078));
    jdff dff_A_smurInE44_0(.din(n21078), .dout(n21081));
    jdff dff_A_cc0bom7j3_0(.din(n21081), .dout(n21084));
    jdff dff_A_oZePYS4c6_0(.din(n21084), .dout(n21087));
    jdff dff_A_Bo94DYig0_0(.din(n21087), .dout(n21090));
    jdff dff_A_MErWuuNG0_0(.din(n21090), .dout(n21093));
    jdff dff_A_pCcJklv01_0(.din(n21093), .dout(n21096));
    jdff dff_A_JKooQMiB5_0(.din(n21096), .dout(n21099));
    jdff dff_A_KKURhmtQ4_0(.din(n21099), .dout(n21102));
    jdff dff_A_QmFJHWQj2_0(.din(n21102), .dout(n21105));
    jdff dff_A_SFC6N8698_0(.din(n21105), .dout(n21108));
    jdff dff_A_6rukfAPk6_0(.din(n21108), .dout(n21111));
    jdff dff_A_YTZ4OCzy0_0(.din(n21111), .dout(n21114));
    jdff dff_A_OZW0BpKb4_0(.din(n21114), .dout(n21117));
    jdff dff_A_Pkn8qxHJ5_0(.din(n21117), .dout(n21120));
    jdff dff_A_PCekqYEQ0_0(.din(n21120), .dout(G594));
    jdff dff_A_2GuE02g96_1(.din(n306), .dout(n21126));
    jdff dff_A_0qKeY6Yy4_0(.din(n21126), .dout(n21129));
    jdff dff_A_P27MWUUx8_0(.din(n21129), .dout(n21132));
    jdff dff_A_kllTJxuw5_0(.din(n21132), .dout(n21135));
    jdff dff_A_XIJ9hcLF3_0(.din(n21135), .dout(n21138));
    jdff dff_A_uMbhdoe53_0(.din(n21138), .dout(n21141));
    jdff dff_A_uVwGQOzg1_0(.din(n21141), .dout(n21144));
    jdff dff_A_ajn1NoHo4_0(.din(n21144), .dout(n21147));
    jdff dff_A_ZMYKSxSU9_0(.din(n21147), .dout(n21150));
    jdff dff_A_4h0mS7gB3_0(.din(n21150), .dout(n21153));
    jdff dff_A_RrypEcrR9_0(.din(n21153), .dout(n21156));
    jdff dff_A_Xjea6bvo8_0(.din(n21156), .dout(n21159));
    jdff dff_A_QKlP35xm6_0(.din(n21159), .dout(n21162));
    jdff dff_A_ce8jm6bc2_0(.din(n21162), .dout(n21165));
    jdff dff_A_fXEt5rXm9_0(.din(n21165), .dout(n21168));
    jdff dff_A_HNZ1HHDk2_0(.din(n21168), .dout(n21171));
    jdff dff_A_cm8vsMiB2_0(.din(n21171), .dout(n21174));
    jdff dff_A_mN0D8Rpu3_0(.din(n21174), .dout(n21177));
    jdff dff_A_Q8rV6Zat7_0(.din(n21177), .dout(n21180));
    jdff dff_A_t7wZdGwX1_0(.din(n21180), .dout(n21183));
    jdff dff_A_KJ8rTuVl5_0(.din(n21183), .dout(n21186));
    jdff dff_A_zlVkK4YB4_0(.din(n21186), .dout(n21189));
    jdff dff_A_Taqzk2LZ4_0(.din(n21189), .dout(n21192));
    jdff dff_A_S6zLf6W24_0(.din(n21192), .dout(n21195));
    jdff dff_A_7r8n76n82_0(.din(n21195), .dout(n21198));
    jdff dff_A_GVBvY17J3_0(.din(n21198), .dout(n21201));
    jdff dff_A_qZdKgzVe7_0(.din(n21201), .dout(G599));
    jdff dff_A_63AobLUF2_1(.din(n309), .dout(n21207));
    jdff dff_A_dAlUDEjG1_0(.din(n21207), .dout(n21210));
    jdff dff_A_tejdBBNT0_0(.din(n21210), .dout(n21213));
    jdff dff_A_xzriuna22_0(.din(n21213), .dout(n21216));
    jdff dff_A_Mf5s9S5i2_0(.din(n21216), .dout(n21219));
    jdff dff_A_phDcnlxx3_0(.din(n21219), .dout(n21222));
    jdff dff_A_Ld3TBmQB5_0(.din(n21222), .dout(n21225));
    jdff dff_A_aCUV8FGK3_0(.din(n21225), .dout(n21228));
    jdff dff_A_ylPMQHgv6_0(.din(n21228), .dout(n21231));
    jdff dff_A_18iQsGit3_0(.din(n21231), .dout(n21234));
    jdff dff_A_HQp5Isk29_0(.din(n21234), .dout(n21237));
    jdff dff_A_4pNBlFnC9_0(.din(n21237), .dout(n21240));
    jdff dff_A_cegTMNkz5_0(.din(n21240), .dout(n21243));
    jdff dff_A_LuWf17Ek6_0(.din(n21243), .dout(n21246));
    jdff dff_A_olEg0y025_0(.din(n21246), .dout(n21249));
    jdff dff_A_tmqmlhJE8_0(.din(n21249), .dout(n21252));
    jdff dff_A_LNVrH9Rq0_0(.din(n21252), .dout(n21255));
    jdff dff_A_exksNRci6_0(.din(n21255), .dout(n21258));
    jdff dff_A_KVigNA9U1_0(.din(n21258), .dout(n21261));
    jdff dff_A_dAUd8jss8_0(.din(n21261), .dout(n21264));
    jdff dff_A_d9VRJBek8_0(.din(n21264), .dout(n21267));
    jdff dff_A_n6PlnGlr2_0(.din(n21267), .dout(n21270));
    jdff dff_A_5wiTCPxQ0_0(.din(n21270), .dout(n21273));
    jdff dff_A_Ne1VqeQd2_0(.din(n21273), .dout(n21276));
    jdff dff_A_ToJmm2N25_0(.din(n21276), .dout(n21279));
    jdff dff_A_Iy23Gdq82_0(.din(n21279), .dout(n21282));
    jdff dff_A_A0RiMfTY7_0(.din(n21282), .dout(G600));
    jdff dff_A_xSrgjd2r2_1(.din(n313), .dout(n21288));
    jdff dff_A_z1MV1RVm5_0(.din(n21288), .dout(n21291));
    jdff dff_A_NCvQSvrP0_0(.din(n21291), .dout(n21294));
    jdff dff_A_31ZmXWPA6_0(.din(n21294), .dout(n21297));
    jdff dff_A_rzdzpzl07_0(.din(n21297), .dout(n21300));
    jdff dff_A_8yCoMCvI6_0(.din(n21300), .dout(n21303));
    jdff dff_A_YwJr4WJK3_0(.din(n21303), .dout(n21306));
    jdff dff_A_Ow12GLnX5_0(.din(n21306), .dout(n21309));
    jdff dff_A_BEeT3fNA1_0(.din(n21309), .dout(n21312));
    jdff dff_A_258yxaEp7_0(.din(n21312), .dout(n21315));
    jdff dff_A_Bea28Dpj7_0(.din(n21315), .dout(n21318));
    jdff dff_A_gXe7JpOF8_0(.din(n21318), .dout(n21321));
    jdff dff_A_rRlDJQLa1_0(.din(n21321), .dout(n21324));
    jdff dff_A_jyi9a2ds0_0(.din(n21324), .dout(n21327));
    jdff dff_A_AvGh5mxf9_0(.din(n21327), .dout(n21330));
    jdff dff_A_DfVOl6jg6_0(.din(n21330), .dout(n21333));
    jdff dff_A_W1Q5HWHK8_0(.din(n21333), .dout(n21336));
    jdff dff_A_9QFRuSy82_0(.din(n21336), .dout(n21339));
    jdff dff_A_Ljxk9B0y1_0(.din(n21339), .dout(n21342));
    jdff dff_A_xkJtNxKY0_0(.din(n21342), .dout(n21345));
    jdff dff_A_RZNQa8Zp0_0(.din(n21345), .dout(n21348));
    jdff dff_A_sAMT18Ip3_0(.din(n21348), .dout(n21351));
    jdff dff_A_FOkR76ml9_0(.din(n21351), .dout(n21354));
    jdff dff_A_AXurrEUk1_0(.din(n21354), .dout(n21357));
    jdff dff_A_HhopjXlZ5_0(.din(n21357), .dout(n21360));
    jdff dff_A_EnmNRsPi0_0(.din(n21360), .dout(n21363));
    jdff dff_A_dKQThvRv8_0(.din(n21363), .dout(G601));
    jdff dff_A_FJrUYRUW2_1(.din(n316), .dout(n21369));
    jdff dff_A_midEEXwi6_0(.din(n21369), .dout(n21372));
    jdff dff_A_nEvJflSm7_0(.din(n21372), .dout(n21375));
    jdff dff_A_SESSf9AI6_0(.din(n21375), .dout(n21378));
    jdff dff_A_YsZvdVsm1_0(.din(n21378), .dout(n21381));
    jdff dff_A_btPF0H3W0_0(.din(n21381), .dout(n21384));
    jdff dff_A_M0YggQ760_0(.din(n21384), .dout(n21387));
    jdff dff_A_SzLWu1io6_0(.din(n21387), .dout(n21390));
    jdff dff_A_dZB7ziFm4_0(.din(n21390), .dout(n21393));
    jdff dff_A_9XyS5e731_0(.din(n21393), .dout(n21396));
    jdff dff_A_r8lzG5NM2_0(.din(n21396), .dout(n21399));
    jdff dff_A_QPF6Efy87_0(.din(n21399), .dout(n21402));
    jdff dff_A_sZTpVlYA9_0(.din(n21402), .dout(n21405));
    jdff dff_A_BNg0veXI8_0(.din(n21405), .dout(n21408));
    jdff dff_A_FdehvAmM2_0(.din(n21408), .dout(n21411));
    jdff dff_A_fs63tjHV7_0(.din(n21411), .dout(n21414));
    jdff dff_A_nX1Dl57M2_0(.din(n21414), .dout(n21417));
    jdff dff_A_gtSoiKOo4_0(.din(n21417), .dout(n21420));
    jdff dff_A_RMXDH7rG7_0(.din(n21420), .dout(n21423));
    jdff dff_A_ymzgro2G8_0(.din(n21423), .dout(n21426));
    jdff dff_A_eCLMDY9V5_0(.din(n21426), .dout(n21429));
    jdff dff_A_JmltyGqX9_0(.din(n21429), .dout(n21432));
    jdff dff_A_zrdcGyY85_0(.din(n21432), .dout(n21435));
    jdff dff_A_LRXr5ju66_0(.din(n21435), .dout(n21438));
    jdff dff_A_VhDntoKw5_0(.din(n21438), .dout(n21441));
    jdff dff_A_oGAw2bVZ4_0(.din(n21441), .dout(n21444));
    jdff dff_A_zYPLqGsr8_0(.din(n21444), .dout(G602));
    jdff dff_A_hsW6rtkC8_1(.din(n5765), .dout(n21450));
    jdff dff_A_szKiCzJS1_0(.din(n21450), .dout(n21453));
    jdff dff_A_yJBiMRC79_0(.din(n21453), .dout(n21456));
    jdff dff_A_Z9VSso8D1_0(.din(n21456), .dout(n21459));
    jdff dff_A_gZdKDqab3_0(.din(n21459), .dout(n21462));
    jdff dff_A_9RZ0kxKC1_0(.din(n21462), .dout(n21465));
    jdff dff_A_Tf7IENfH1_0(.din(n21465), .dout(n21468));
    jdff dff_A_6c6RHEE55_0(.din(n21468), .dout(n21471));
    jdff dff_A_Cj9JVRMP3_0(.din(n21471), .dout(n21474));
    jdff dff_A_TWAnU5KB2_0(.din(n21474), .dout(n21477));
    jdff dff_A_EYi4WWD14_0(.din(n21477), .dout(n21480));
    jdff dff_A_Jv1Yxix80_0(.din(n21480), .dout(n21483));
    jdff dff_A_GezRUYTJ9_0(.din(n21483), .dout(n21486));
    jdff dff_A_IbrxoSpm7_0(.din(n21486), .dout(n21489));
    jdff dff_A_ruY906Ta4_0(.din(n21489), .dout(n21492));
    jdff dff_A_irFwQcnP4_0(.din(n21492), .dout(n21495));
    jdff dff_A_OuKPEvKB0_0(.din(n21495), .dout(n21498));
    jdff dff_A_7c4ZfVoG7_0(.din(n21498), .dout(n21501));
    jdff dff_A_N3TJd7Gp5_0(.din(n21501), .dout(n21504));
    jdff dff_A_tgloV8av7_0(.din(n21504), .dout(n21507));
    jdff dff_A_Xets2Obk2_0(.din(n21507), .dout(n21510));
    jdff dff_A_RKyVqdFx5_0(.din(n21510), .dout(n21513));
    jdff dff_A_eXir635X9_0(.din(n21513), .dout(n21516));
    jdff dff_A_KPIQcHyP7_0(.din(n21516), .dout(n21519));
    jdff dff_A_pdkIhO8J0_0(.din(n21519), .dout(n21522));
    jdff dff_A_GNYTEDO03_0(.din(n21522), .dout(n21525));
    jdff dff_A_I2luZ5AD4_0(.din(n21525), .dout(G603));
    jdff dff_A_PX3V940Q1_1(.din(n5768), .dout(n21531));
    jdff dff_A_Szlr61vU3_0(.din(n21531), .dout(n21534));
    jdff dff_A_txxwIzN43_0(.din(n21534), .dout(n21537));
    jdff dff_A_TcaYo2gG9_0(.din(n21537), .dout(n21540));
    jdff dff_A_JhxAfswL4_0(.din(n21540), .dout(n21543));
    jdff dff_A_57InIhXx1_0(.din(n21543), .dout(n21546));
    jdff dff_A_qYmlp08P4_0(.din(n21546), .dout(n21549));
    jdff dff_A_xxcY15o56_0(.din(n21549), .dout(n21552));
    jdff dff_A_SyNuU87b4_0(.din(n21552), .dout(n21555));
    jdff dff_A_3axgsdQM0_0(.din(n21555), .dout(n21558));
    jdff dff_A_CHWLo9YL9_0(.din(n21558), .dout(n21561));
    jdff dff_A_w6Npeprv7_0(.din(n21561), .dout(n21564));
    jdff dff_A_iA6SLOYw2_0(.din(n21564), .dout(n21567));
    jdff dff_A_VpihWe7C8_0(.din(n21567), .dout(n21570));
    jdff dff_A_vmXYj26E5_0(.din(n21570), .dout(n21573));
    jdff dff_A_Wj1A375y5_0(.din(n21573), .dout(n21576));
    jdff dff_A_oUPPLDIT1_0(.din(n21576), .dout(n21579));
    jdff dff_A_fFCFGCtw3_0(.din(n21579), .dout(n21582));
    jdff dff_A_gxbjnoIh6_0(.din(n21582), .dout(n21585));
    jdff dff_A_40w87G6r0_0(.din(n21585), .dout(n21588));
    jdff dff_A_7Nczw42J7_0(.din(n21588), .dout(n21591));
    jdff dff_A_bjmRyeJX8_0(.din(n21591), .dout(n21594));
    jdff dff_A_D3aERHvU1_0(.din(n21594), .dout(n21597));
    jdff dff_A_tsTZTo0n4_0(.din(n21597), .dout(n21600));
    jdff dff_A_eOrHbXe88_0(.din(n21600), .dout(n21603));
    jdff dff_A_bmPpN7js2_0(.din(n21603), .dout(n21606));
    jdff dff_A_jf8spJsC9_0(.din(n21606), .dout(G604));
    jdff dff_A_FpfbrbRf3_1(.din(n319), .dout(n21612));
    jdff dff_A_hWBhh0uA5_0(.din(n21612), .dout(n21615));
    jdff dff_A_DF2pDixM4_0(.din(n21615), .dout(n21618));
    jdff dff_A_uuuBjRoR1_0(.din(n21618), .dout(n21621));
    jdff dff_A_WohuxkYd2_0(.din(n21621), .dout(n21624));
    jdff dff_A_Ir2xvp0x1_0(.din(n21624), .dout(n21627));
    jdff dff_A_afzONmUh7_0(.din(n21627), .dout(n21630));
    jdff dff_A_jKnjhFfZ6_0(.din(n21630), .dout(n21633));
    jdff dff_A_YS4lJjbE0_0(.din(n21633), .dout(n21636));
    jdff dff_A_sV06MLaO8_0(.din(n21636), .dout(n21639));
    jdff dff_A_8K2SK2cJ2_0(.din(n21639), .dout(n21642));
    jdff dff_A_YJ15L2IW5_0(.din(n21642), .dout(n21645));
    jdff dff_A_PkL00IS48_0(.din(n21645), .dout(n21648));
    jdff dff_A_gBzSJv3r7_0(.din(n21648), .dout(n21651));
    jdff dff_A_BVzplejU9_0(.din(n21651), .dout(n21654));
    jdff dff_A_Zj3TXxVz6_0(.din(n21654), .dout(n21657));
    jdff dff_A_tsCG02bx4_0(.din(n21657), .dout(n21660));
    jdff dff_A_D1O1SYim5_0(.din(n21660), .dout(n21663));
    jdff dff_A_HGvRUoVW5_0(.din(n21663), .dout(n21666));
    jdff dff_A_cSJqokbd4_0(.din(n21666), .dout(n21669));
    jdff dff_A_nwWD9v3C3_0(.din(n21669), .dout(n21672));
    jdff dff_A_9P9q7ot19_0(.din(n21672), .dout(n21675));
    jdff dff_A_QSwPkL6k4_0(.din(n21675), .dout(n21678));
    jdff dff_A_eo6KGMVz7_0(.din(n21678), .dout(n21681));
    jdff dff_A_3prTw2Z20_0(.din(n21681), .dout(n21684));
    jdff dff_A_ZyehewfO2_0(.din(n21684), .dout(n21687));
    jdff dff_A_nCxU7v4v1_0(.din(n21687), .dout(G611));
    jdff dff_A_ngtpAtsY5_1(.din(n322), .dout(n21693));
    jdff dff_A_dI8qiuRa9_0(.din(n21693), .dout(n21696));
    jdff dff_A_XS6ojzl56_0(.din(n21696), .dout(n21699));
    jdff dff_A_pSpZeeOU2_0(.din(n21699), .dout(n21702));
    jdff dff_A_xfaVxp8y8_0(.din(n21702), .dout(n21705));
    jdff dff_A_SQJ3DB1P9_0(.din(n21705), .dout(n21708));
    jdff dff_A_uzOI3sGp8_0(.din(n21708), .dout(n21711));
    jdff dff_A_p3Xx526u7_0(.din(n21711), .dout(n21714));
    jdff dff_A_WV6L8kQ13_0(.din(n21714), .dout(n21717));
    jdff dff_A_uexmfjaw3_0(.din(n21717), .dout(n21720));
    jdff dff_A_9MXOBaWj9_0(.din(n21720), .dout(n21723));
    jdff dff_A_I8JayFcY4_0(.din(n21723), .dout(n21726));
    jdff dff_A_PAx9P8q05_0(.din(n21726), .dout(n21729));
    jdff dff_A_4DQmtHqt2_0(.din(n21729), .dout(n21732));
    jdff dff_A_88KhvHXC0_0(.din(n21732), .dout(n21735));
    jdff dff_A_50UI5PGD0_0(.din(n21735), .dout(n21738));
    jdff dff_A_GkKeEPc17_0(.din(n21738), .dout(n21741));
    jdff dff_A_vLElKZTm0_0(.din(n21741), .dout(n21744));
    jdff dff_A_HBHEkfUe2_0(.din(n21744), .dout(n21747));
    jdff dff_A_uCqDNxO10_0(.din(n21747), .dout(n21750));
    jdff dff_A_QRwZmUjI4_0(.din(n21750), .dout(n21753));
    jdff dff_A_chnGNUjU5_0(.din(n21753), .dout(n21756));
    jdff dff_A_2GV3F85s8_0(.din(n21756), .dout(n21759));
    jdff dff_A_dnBudaaR9_0(.din(n21759), .dout(n21762));
    jdff dff_A_ZQ8Rg5qF5_0(.din(n21762), .dout(n21765));
    jdff dff_A_lq9Bm5JV2_0(.din(n21765), .dout(n21768));
    jdff dff_A_9T2mPAHf9_0(.din(n21768), .dout(G612));
    jdff dff_A_5cfRan3F4_2(.din(n326), .dout(n21774));
    jdff dff_A_TNeGIopd8_0(.din(n21774), .dout(n21777));
    jdff dff_A_cliTpmkT3_0(.din(n21777), .dout(n21780));
    jdff dff_A_DcGSxjqq2_0(.din(n21780), .dout(n21783));
    jdff dff_A_FV1UWYjJ3_0(.din(n21783), .dout(n21786));
    jdff dff_A_QhuGMRpv6_0(.din(n21786), .dout(n21789));
    jdff dff_A_gvTpK0tC8_0(.din(n21789), .dout(n21792));
    jdff dff_A_fSPPQFY42_0(.din(n21792), .dout(n21795));
    jdff dff_A_C8pYUjey9_0(.din(n21795), .dout(n21798));
    jdff dff_A_Dq5SKNWG6_0(.din(n21798), .dout(n21801));
    jdff dff_A_5Qp6DBuz4_0(.din(n21801), .dout(n21804));
    jdff dff_A_IYpkiHMX6_0(.din(n21804), .dout(n21807));
    jdff dff_A_WWeMLzkC5_0(.din(n21807), .dout(n21810));
    jdff dff_A_6bTjRrRU4_0(.din(n21810), .dout(n21813));
    jdff dff_A_MYVkEitD8_0(.din(n21813), .dout(n21816));
    jdff dff_A_cSWIX6eW9_0(.din(n21816), .dout(n21819));
    jdff dff_A_KGf7Iqt45_0(.din(n21819), .dout(n21822));
    jdff dff_A_FoV0X4GM5_0(.din(n21822), .dout(n21825));
    jdff dff_A_Bty9xsM37_0(.din(n21825), .dout(n21828));
    jdff dff_A_JufoRDEz4_0(.din(n21828), .dout(n21831));
    jdff dff_A_uk2DcbNv8_0(.din(n21831), .dout(n21834));
    jdff dff_A_3RmbsgOM2_0(.din(n21834), .dout(n21837));
    jdff dff_A_soGFIDx60_0(.din(n21837), .dout(n21840));
    jdff dff_A_0Asvl05L1_0(.din(n21840), .dout(n21843));
    jdff dff_A_vG3AJPai3_0(.din(n21843), .dout(n21846));
    jdff dff_A_2VOakzUt5_0(.din(n21846), .dout(n21849));
    jdff dff_A_mJOSM8RJ0_0(.din(n21849), .dout(G810));
    jdff dff_A_5t6DzlqV5_1(.din(n329), .dout(n21855));
    jdff dff_A_AkO6TqAN1_0(.din(n21855), .dout(n21858));
    jdff dff_A_0fViiNHk7_0(.din(n21858), .dout(n21861));
    jdff dff_A_KMSQqxDl9_0(.din(n21861), .dout(n21864));
    jdff dff_A_ClQuB2hj4_0(.din(n21864), .dout(n21867));
    jdff dff_A_56vSMsC89_0(.din(n21867), .dout(n21870));
    jdff dff_A_GGQcJnL39_0(.din(n21870), .dout(n21873));
    jdff dff_A_Ek0i76k61_0(.din(n21873), .dout(n21876));
    jdff dff_A_blfsYTeX7_0(.din(n21876), .dout(n21879));
    jdff dff_A_SSTP5gav9_0(.din(n21879), .dout(n21882));
    jdff dff_A_IUJH1Rzh6_0(.din(n21882), .dout(n21885));
    jdff dff_A_UnpMCpFA6_0(.din(n21885), .dout(n21888));
    jdff dff_A_toLzv5Wz8_0(.din(n21888), .dout(n21891));
    jdff dff_A_9cBlObww6_0(.din(n21891), .dout(n21894));
    jdff dff_A_rZeDuzOa5_0(.din(n21894), .dout(n21897));
    jdff dff_A_jzQ6eMdj7_0(.din(n21897), .dout(n21900));
    jdff dff_A_DjBUioum9_0(.din(n21900), .dout(n21903));
    jdff dff_A_CxweOoky9_0(.din(n21903), .dout(n21906));
    jdff dff_A_bkcEcDCz8_0(.din(n21906), .dout(n21909));
    jdff dff_A_Cp66eVQd7_0(.din(n21909), .dout(n21912));
    jdff dff_A_eljnh0Zq4_0(.din(n21912), .dout(n21915));
    jdff dff_A_dWtolInX2_0(.din(n21915), .dout(n21918));
    jdff dff_A_J9jSSohA0_0(.din(n21918), .dout(n21921));
    jdff dff_A_AzGZECcC4_0(.din(n21921), .dout(n21924));
    jdff dff_A_s23nZGQS9_0(.din(n21924), .dout(n21927));
    jdff dff_A_TtBkZVw68_0(.din(n21927), .dout(n21930));
    jdff dff_A_oLgyeFaj7_0(.din(n21930), .dout(G848));
    jdff dff_A_WU84By202_1(.din(n332), .dout(n21936));
    jdff dff_A_ExbZdFft7_0(.din(n21936), .dout(n21939));
    jdff dff_A_LipODtBL2_0(.din(n21939), .dout(n21942));
    jdff dff_A_IP95x7VF3_0(.din(n21942), .dout(n21945));
    jdff dff_A_ohwzvEnL0_0(.din(n21945), .dout(n21948));
    jdff dff_A_wRzVTGBz1_0(.din(n21948), .dout(n21951));
    jdff dff_A_M1J9ofQx9_0(.din(n21951), .dout(n21954));
    jdff dff_A_XxZuVF487_0(.din(n21954), .dout(n21957));
    jdff dff_A_8CmjZnUN6_0(.din(n21957), .dout(n21960));
    jdff dff_A_en6iky532_0(.din(n21960), .dout(n21963));
    jdff dff_A_vdY2E7GL0_0(.din(n21963), .dout(n21966));
    jdff dff_A_8c4tUJNl4_0(.din(n21966), .dout(n21969));
    jdff dff_A_9s12XcWn3_0(.din(n21969), .dout(n21972));
    jdff dff_A_hKg7IygA9_0(.din(n21972), .dout(n21975));
    jdff dff_A_KaKR3Fko9_0(.din(n21975), .dout(n21978));
    jdff dff_A_Dr8oBaGF7_0(.din(n21978), .dout(n21981));
    jdff dff_A_SzQjdAPg7_0(.din(n21981), .dout(n21984));
    jdff dff_A_WIXvc3nZ4_0(.din(n21984), .dout(n21987));
    jdff dff_A_be6sH0uC5_0(.din(n21987), .dout(n21990));
    jdff dff_A_2dfySpkn9_0(.din(n21990), .dout(n21993));
    jdff dff_A_x9n3u7oK2_0(.din(n21993), .dout(n21996));
    jdff dff_A_y55xJ1ku5_0(.din(n21996), .dout(n21999));
    jdff dff_A_Bdq7bNDo0_0(.din(n21999), .dout(n22002));
    jdff dff_A_7M6NhEP52_0(.din(n22002), .dout(n22005));
    jdff dff_A_k2LO6yXs7_0(.din(n22005), .dout(n22008));
    jdff dff_A_M83EPBTI6_0(.din(n22008), .dout(n22011));
    jdff dff_A_ZVtp3RYb3_0(.din(n22011), .dout(G849));
    jdff dff_A_00yBnyGB8_1(.din(n335), .dout(n22017));
    jdff dff_A_UDlJXt8c6_0(.din(n22017), .dout(n22020));
    jdff dff_A_LMDyBa0b8_0(.din(n22020), .dout(n22023));
    jdff dff_A_JjWo0d4c7_0(.din(n22023), .dout(n22026));
    jdff dff_A_seqQ42bY6_0(.din(n22026), .dout(n22029));
    jdff dff_A_9PjKnYGS6_0(.din(n22029), .dout(n22032));
    jdff dff_A_6NSocSQc1_0(.din(n22032), .dout(n22035));
    jdff dff_A_VogwunOA4_0(.din(n22035), .dout(n22038));
    jdff dff_A_RWtZAbBh4_0(.din(n22038), .dout(n22041));
    jdff dff_A_3umFCYI50_0(.din(n22041), .dout(n22044));
    jdff dff_A_TnSQms2s5_0(.din(n22044), .dout(n22047));
    jdff dff_A_m0PwIy8J4_0(.din(n22047), .dout(n22050));
    jdff dff_A_zxzhDAm66_0(.din(n22050), .dout(n22053));
    jdff dff_A_h6FErAJP6_0(.din(n22053), .dout(n22056));
    jdff dff_A_Vex5MC0l7_0(.din(n22056), .dout(n22059));
    jdff dff_A_7AhQ1E7u2_0(.din(n22059), .dout(n22062));
    jdff dff_A_3zbwA3tH1_0(.din(n22062), .dout(n22065));
    jdff dff_A_ynQ30shl7_0(.din(n22065), .dout(n22068));
    jdff dff_A_NbYM2WC09_0(.din(n22068), .dout(n22071));
    jdff dff_A_yPhRucby9_0(.din(n22071), .dout(n22074));
    jdff dff_A_g9U8ADko8_0(.din(n22074), .dout(n22077));
    jdff dff_A_xFuGE22u5_0(.din(n22077), .dout(n22080));
    jdff dff_A_P4hpayBY0_0(.din(n22080), .dout(n22083));
    jdff dff_A_hCCATq3l4_0(.din(n22083), .dout(n22086));
    jdff dff_A_fIboX2j20_0(.din(n22086), .dout(n22089));
    jdff dff_A_DHO0Yl9L6_0(.din(n22089), .dout(n22092));
    jdff dff_A_W4LvPFHI2_0(.din(n22092), .dout(G850));
    jdff dff_A_9O4gAV2i7_1(.din(n338), .dout(n22098));
    jdff dff_A_VlzhPncD2_0(.din(n22098), .dout(n22101));
    jdff dff_A_mAC2MZIc1_0(.din(n22101), .dout(n22104));
    jdff dff_A_xNV2BHgZ1_0(.din(n22104), .dout(n22107));
    jdff dff_A_2yPk94W95_0(.din(n22107), .dout(n22110));
    jdff dff_A_wrbFE21X9_0(.din(n22110), .dout(n22113));
    jdff dff_A_JEXyzaBW5_0(.din(n22113), .dout(n22116));
    jdff dff_A_WMqTFTfS4_0(.din(n22116), .dout(n22119));
    jdff dff_A_L2x21T8C4_0(.din(n22119), .dout(n22122));
    jdff dff_A_eqxLe8Ly2_0(.din(n22122), .dout(n22125));
    jdff dff_A_poOSoO2I6_0(.din(n22125), .dout(n22128));
    jdff dff_A_dPQMv4Ly5_0(.din(n22128), .dout(n22131));
    jdff dff_A_UTtF3snW4_0(.din(n22131), .dout(n22134));
    jdff dff_A_4CIW0D9p0_0(.din(n22134), .dout(n22137));
    jdff dff_A_2oWqbx8g0_0(.din(n22137), .dout(n22140));
    jdff dff_A_eGUVLsiR1_0(.din(n22140), .dout(n22143));
    jdff dff_A_gFoE7tEK5_0(.din(n22143), .dout(n22146));
    jdff dff_A_qeXe7CHZ3_0(.din(n22146), .dout(n22149));
    jdff dff_A_ll7FEGeB0_0(.din(n22149), .dout(n22152));
    jdff dff_A_yqtzfzdn2_0(.din(n22152), .dout(n22155));
    jdff dff_A_cGLikj2N9_0(.din(n22155), .dout(n22158));
    jdff dff_A_IF9OC0EY6_0(.din(n22158), .dout(n22161));
    jdff dff_A_EVMxK5z23_0(.din(n22161), .dout(n22164));
    jdff dff_A_CJUHXIz74_0(.din(n22164), .dout(n22167));
    jdff dff_A_LPG7EiUM4_0(.din(n22167), .dout(n22170));
    jdff dff_A_wd7LoYRr0_0(.din(n22170), .dout(n22173));
    jdff dff_A_ed7jCAqA2_0(.din(n22173), .dout(G851));
    jdff dff_A_wElPQzTe5_2(.din(n342), .dout(n22179));
    jdff dff_A_4AOl2UH79_0(.din(n22179), .dout(n22182));
    jdff dff_A_JlKtbfur3_0(.din(n22182), .dout(n22185));
    jdff dff_A_DkNyWvK76_0(.din(n22185), .dout(n22188));
    jdff dff_A_mJmbW3Cc4_0(.din(n22188), .dout(n22191));
    jdff dff_A_UzGttZvD9_0(.din(n22191), .dout(n22194));
    jdff dff_A_YNd6SKU43_0(.din(n22194), .dout(n22197));
    jdff dff_A_Ov1Tvs7f5_0(.din(n22197), .dout(n22200));
    jdff dff_A_dA0TC0dG4_0(.din(n22200), .dout(n22203));
    jdff dff_A_ZBWY9wqZ4_0(.din(n22203), .dout(n22206));
    jdff dff_A_AR1uQiiT7_0(.din(n22206), .dout(n22209));
    jdff dff_A_FRkgn1Go4_0(.din(n22209), .dout(n22212));
    jdff dff_A_QPLO1r0R1_0(.din(n22212), .dout(n22215));
    jdff dff_A_UBbajyiL4_0(.din(n22215), .dout(n22218));
    jdff dff_A_nmLoOm7U5_0(.din(n22218), .dout(n22221));
    jdff dff_A_cOdwUzQW6_0(.din(n22221), .dout(n22224));
    jdff dff_A_QGb8wMTu9_0(.din(n22224), .dout(n22227));
    jdff dff_A_LXWUVEv72_0(.din(n22227), .dout(n22230));
    jdff dff_A_qwnZtuUh2_0(.din(n22230), .dout(n22233));
    jdff dff_A_EhaPn7jp7_0(.din(n22233), .dout(n22236));
    jdff dff_A_MuPXOk6G3_0(.din(n22236), .dout(n22239));
    jdff dff_A_eJuhSk0E3_0(.din(n22239), .dout(n22242));
    jdff dff_A_uZ8yTvPd7_0(.din(n22242), .dout(n22245));
    jdff dff_A_eEvjbcGu3_0(.din(n22245), .dout(n22248));
    jdff dff_A_hUtW2DhM9_0(.din(n22248), .dout(n22251));
    jdff dff_A_obxRtBkU9_0(.din(n22251), .dout(n22254));
    jdff dff_A_0UmWNMxX9_0(.din(n22254), .dout(G634));
    jdff dff_A_5ftdZgkS7_2(.din(n349), .dout(n22260));
    jdff dff_A_CMaaRmQY4_0(.din(n22260), .dout(n22263));
    jdff dff_A_TeZA8vRj1_0(.din(n22263), .dout(n22266));
    jdff dff_A_bYTk6TVq9_0(.din(n22266), .dout(n22269));
    jdff dff_A_JtqXfOQ52_0(.din(n22269), .dout(n22272));
    jdff dff_A_Gl0DGDjm2_0(.din(n22272), .dout(n22275));
    jdff dff_A_XBCRh5Pa5_0(.din(n22275), .dout(n22278));
    jdff dff_A_hXemu6u64_0(.din(n22278), .dout(n22281));
    jdff dff_A_7qpG2OMS7_0(.din(n22281), .dout(n22284));
    jdff dff_A_j2lCvmCJ4_0(.din(n22284), .dout(n22287));
    jdff dff_A_lTi6JReR2_0(.din(n22287), .dout(n22290));
    jdff dff_A_9NPOSaKl7_0(.din(n22290), .dout(n22293));
    jdff dff_A_BrrOSoGj3_0(.din(n22293), .dout(n22296));
    jdff dff_A_VfwoEhfr4_0(.din(n22296), .dout(n22299));
    jdff dff_A_sgMNeLux8_0(.din(n22299), .dout(n22302));
    jdff dff_A_tuU4C99N4_0(.din(n22302), .dout(n22305));
    jdff dff_A_rzzQlwH61_0(.din(n22305), .dout(n22308));
    jdff dff_A_iGuArtNh5_0(.din(n22308), .dout(n22311));
    jdff dff_A_3Qf12oSp8_0(.din(n22311), .dout(n22314));
    jdff dff_A_8w1NMvb74_0(.din(n22314), .dout(n22317));
    jdff dff_A_aDNivSHy6_0(.din(n22317), .dout(n22320));
    jdff dff_A_yj4CGCgA1_0(.din(n22320), .dout(n22323));
    jdff dff_A_WrKFg0mw8_0(.din(n22323), .dout(n22326));
    jdff dff_A_c0JWgtOE4_0(.din(n22326), .dout(n22329));
    jdff dff_A_BzV8wqwf9_0(.din(n22329), .dout(n22332));
    jdff dff_A_4CP3EiGh6_0(.din(n22332), .dout(G815));
    jdff dff_A_nNW8Oyib6_2(.din(n356), .dout(n22338));
    jdff dff_A_n2FdJ63z5_0(.din(n22338), .dout(n22341));
    jdff dff_A_3hoEDqA48_0(.din(n22341), .dout(n22344));
    jdff dff_A_sysUsWEc8_0(.din(n22344), .dout(n22347));
    jdff dff_A_CYim9ad56_0(.din(n22347), .dout(n22350));
    jdff dff_A_bbMcMkbS4_0(.din(n22350), .dout(n22353));
    jdff dff_A_usgfN2SQ1_0(.din(n22353), .dout(n22356));
    jdff dff_A_ZHwqDeh71_0(.din(n22356), .dout(n22359));
    jdff dff_A_23SLu1YI9_0(.din(n22359), .dout(n22362));
    jdff dff_A_i3VyskVW1_0(.din(n22362), .dout(n22365));
    jdff dff_A_dtyqkMfr6_0(.din(n22365), .dout(n22368));
    jdff dff_A_U7dZrVpH5_0(.din(n22368), .dout(n22371));
    jdff dff_A_1KddJRVb4_0(.din(n22371), .dout(n22374));
    jdff dff_A_9Y8SiPe14_0(.din(n22374), .dout(n22377));
    jdff dff_A_cNKUpofq4_0(.din(n22377), .dout(n22380));
    jdff dff_A_uFhzg1g85_0(.din(n22380), .dout(n22383));
    jdff dff_A_Im1meCHG2_0(.din(n22383), .dout(n22386));
    jdff dff_A_oTmKnql35_0(.din(n22386), .dout(n22389));
    jdff dff_A_UtBCzH9v6_0(.din(n22389), .dout(n22392));
    jdff dff_A_eiCgoMAU3_0(.din(n22392), .dout(n22395));
    jdff dff_A_6lobc3xM7_0(.din(n22395), .dout(n22398));
    jdff dff_A_z3VMAUdJ6_0(.din(n22398), .dout(n22401));
    jdff dff_A_1sDwaukh1_0(.din(n22401), .dout(n22404));
    jdff dff_A_jfUiw9GR5_0(.din(n22404), .dout(n22407));
    jdff dff_A_ubHt4fJJ2_0(.din(n22407), .dout(n22410));
    jdff dff_A_lshyIWXp2_0(.din(n22410), .dout(G845));
    jdff dff_A_IZSXO4y19_1(.din(n363), .dout(n22416));
    jdff dff_A_FdvWJKLi8_0(.din(n22416), .dout(n22419));
    jdff dff_A_DrzRPN2R6_0(.din(n22419), .dout(n22422));
    jdff dff_A_2lRx43hP9_0(.din(n22422), .dout(n22425));
    jdff dff_A_32fzlnBH8_0(.din(n22425), .dout(n22428));
    jdff dff_A_7DbEmEQ39_0(.din(n22428), .dout(n22431));
    jdff dff_A_n1W7Q6ga7_0(.din(n22431), .dout(n22434));
    jdff dff_A_nP5pYstd3_0(.din(n22434), .dout(n22437));
    jdff dff_A_XSXuxrB71_0(.din(n22437), .dout(n22440));
    jdff dff_A_QCC3DIq40_0(.din(n22440), .dout(n22443));
    jdff dff_A_45UY7L592_0(.din(n22443), .dout(n22446));
    jdff dff_A_M4L6E43p3_0(.din(n22446), .dout(n22449));
    jdff dff_A_vmM6rYJd2_0(.din(n22449), .dout(n22452));
    jdff dff_A_ACNoAteu2_0(.din(n22452), .dout(n22455));
    jdff dff_A_wNhRjP6A5_0(.din(n22455), .dout(n22458));
    jdff dff_A_S0oksRfg3_0(.din(n22458), .dout(n22461));
    jdff dff_A_JZIrDp5I0_0(.din(n22461), .dout(n22464));
    jdff dff_A_KicmJWUX2_0(.din(n22464), .dout(n22467));
    jdff dff_A_PgAkvC1X2_0(.din(n22467), .dout(n22470));
    jdff dff_A_8gATiKRr1_0(.din(n22470), .dout(n22473));
    jdff dff_A_pgriklao0_0(.din(n22473), .dout(n22476));
    jdff dff_A_X5LgeMM37_0(.din(n22476), .dout(n22479));
    jdff dff_A_8HS1W8TA4_0(.din(n22479), .dout(n22482));
    jdff dff_A_lEUlsqKZ1_0(.din(n22482), .dout(n22485));
    jdff dff_A_KDgHikqk8_0(.din(n22485), .dout(n22488));
    jdff dff_A_BoNDu9p83_0(.din(n22488), .dout(G847));
    jdff dff_A_tBsHYMsf0_1(.din(n5771), .dout(n22494));
    jdff dff_A_Di9tBEy93_0(.din(n22494), .dout(n22497));
    jdff dff_A_FRrNlEBd4_0(.din(n22497), .dout(n22500));
    jdff dff_A_KDHxzONX2_0(.din(n22500), .dout(n22503));
    jdff dff_A_tb6xgNvv2_0(.din(n22503), .dout(n22506));
    jdff dff_A_16iSviNr2_0(.din(n22506), .dout(n22509));
    jdff dff_A_rlu5irWz5_0(.din(n22509), .dout(n22512));
    jdff dff_A_2TB6mGr13_0(.din(n22512), .dout(n22515));
    jdff dff_A_yIYqBvIk8_0(.din(n22515), .dout(n22518));
    jdff dff_A_nL8meCCM3_0(.din(n22518), .dout(n22521));
    jdff dff_A_fqKWxqRr2_0(.din(n22521), .dout(n22524));
    jdff dff_A_NUY8XYjB8_0(.din(n22524), .dout(n22527));
    jdff dff_A_gAw9JrmO5_0(.din(n22527), .dout(n22530));
    jdff dff_A_abkL6C4w1_0(.din(n22530), .dout(n22533));
    jdff dff_A_7fPhmR1o3_0(.din(n22533), .dout(n22536));
    jdff dff_A_ieokOxlL6_0(.din(n22536), .dout(n22539));
    jdff dff_A_xmzZY5IA8_0(.din(n22539), .dout(n22542));
    jdff dff_A_lL5ppykf2_0(.din(n22542), .dout(n22545));
    jdff dff_A_1fZ3Z1300_0(.din(n22545), .dout(n22548));
    jdff dff_A_A7DEkHDH2_0(.din(n22548), .dout(n22551));
    jdff dff_A_sdzZicac3_0(.din(n22551), .dout(n22554));
    jdff dff_A_vn2J0xgn3_0(.din(n22554), .dout(n22557));
    jdff dff_A_moB7jOxG0_0(.din(n22557), .dout(n22560));
    jdff dff_A_MpMlg4gU8_0(.din(n22560), .dout(n22563));
    jdff dff_A_E8J6kf2r8_0(.din(n22563), .dout(n22566));
    jdff dff_A_hyqtacLo7_0(.din(n22566), .dout(n22569));
    jdff dff_A_fchFTvy15_0(.din(n22569), .dout(G926));
    jdff dff_A_tPCLe9f04_1(.din(n5774), .dout(n22575));
    jdff dff_A_APa8b5xU3_0(.din(n22575), .dout(n22578));
    jdff dff_A_0kTMdKbI4_0(.din(n22578), .dout(n22581));
    jdff dff_A_AUCit7yg7_0(.din(n22581), .dout(n22584));
    jdff dff_A_QZ0dxaob8_0(.din(n22584), .dout(n22587));
    jdff dff_A_t9fDaZFZ9_0(.din(n22587), .dout(n22590));
    jdff dff_A_XEpRULQ03_0(.din(n22590), .dout(n22593));
    jdff dff_A_66Gf8kif4_0(.din(n22593), .dout(n22596));
    jdff dff_A_rHx8OWQg6_0(.din(n22596), .dout(n22599));
    jdff dff_A_mcoIyVux9_0(.din(n22599), .dout(n22602));
    jdff dff_A_s69KssoD8_0(.din(n22602), .dout(n22605));
    jdff dff_A_NFtq4UzW4_0(.din(n22605), .dout(n22608));
    jdff dff_A_UHkfVC438_0(.din(n22608), .dout(n22611));
    jdff dff_A_w0cdKska7_0(.din(n22611), .dout(n22614));
    jdff dff_A_odd9nTRY5_0(.din(n22614), .dout(n22617));
    jdff dff_A_BQ1Z48kf7_0(.din(n22617), .dout(n22620));
    jdff dff_A_nvUjCZu32_0(.din(n22620), .dout(n22623));
    jdff dff_A_nLZSCQ2u2_0(.din(n22623), .dout(n22626));
    jdff dff_A_aqnbexse8_0(.din(n22626), .dout(n22629));
    jdff dff_A_sk1Spi356_0(.din(n22629), .dout(n22632));
    jdff dff_A_pb3IABQT4_0(.din(n22632), .dout(n22635));
    jdff dff_A_ouqLDWaW0_0(.din(n22635), .dout(n22638));
    jdff dff_A_01kzzUme9_0(.din(n22638), .dout(n22641));
    jdff dff_A_KXvKvncn6_0(.din(n22641), .dout(n22644));
    jdff dff_A_ClpyFt7J9_0(.din(n22644), .dout(n22647));
    jdff dff_A_aZQfPyvd9_0(.din(n22647), .dout(n22650));
    jdff dff_A_dafibjqx9_0(.din(n22650), .dout(G923));
    jdff dff_A_mnbyVjQA2_1(.din(n5777), .dout(n22656));
    jdff dff_A_Jm13IGCP0_0(.din(n22656), .dout(n22659));
    jdff dff_A_fhbz7wsS6_0(.din(n22659), .dout(n22662));
    jdff dff_A_UlAn2Kdo1_0(.din(n22662), .dout(n22665));
    jdff dff_A_J3GvyTlB8_0(.din(n22665), .dout(n22668));
    jdff dff_A_cBNDgBw72_0(.din(n22668), .dout(n22671));
    jdff dff_A_5kuH9gVS2_0(.din(n22671), .dout(n22674));
    jdff dff_A_b052TarJ5_0(.din(n22674), .dout(n22677));
    jdff dff_A_NzKOpNRB5_0(.din(n22677), .dout(n22680));
    jdff dff_A_L5yaxj4p3_0(.din(n22680), .dout(n22683));
    jdff dff_A_317FVENG8_0(.din(n22683), .dout(n22686));
    jdff dff_A_LKKJsjVo7_0(.din(n22686), .dout(n22689));
    jdff dff_A_bCx5BuDl4_0(.din(n22689), .dout(n22692));
    jdff dff_A_6DjmhvjB9_0(.din(n22692), .dout(n22695));
    jdff dff_A_DWYFI0Vn2_0(.din(n22695), .dout(n22698));
    jdff dff_A_7e0zUIbQ6_0(.din(n22698), .dout(n22701));
    jdff dff_A_lOZo7eb14_0(.din(n22701), .dout(n22704));
    jdff dff_A_wP2WmMbE2_0(.din(n22704), .dout(n22707));
    jdff dff_A_mwwNQD667_0(.din(n22707), .dout(n22710));
    jdff dff_A_f462eIbp7_0(.din(n22710), .dout(n22713));
    jdff dff_A_6gt7HUvI4_0(.din(n22713), .dout(n22716));
    jdff dff_A_wjDFJL4O0_0(.din(n22716), .dout(n22719));
    jdff dff_A_vieZz9Ka5_0(.din(n22719), .dout(n22722));
    jdff dff_A_1qpbX8co8_0(.din(n22722), .dout(n22725));
    jdff dff_A_2bmp3zIS0_0(.din(n22725), .dout(n22728));
    jdff dff_A_RcPgZUiL4_0(.din(n22728), .dout(n22731));
    jdff dff_A_knvHDWqy4_0(.din(n22731), .dout(G921));
    jdff dff_A_HsXSJqmW2_1(.din(n5780), .dout(n22737));
    jdff dff_A_OKpwcyB81_0(.din(n22737), .dout(n22740));
    jdff dff_A_3F3vAHQd6_0(.din(n22740), .dout(n22743));
    jdff dff_A_rggA0Xjo4_0(.din(n22743), .dout(n22746));
    jdff dff_A_vtwirMfd2_0(.din(n22746), .dout(n22749));
    jdff dff_A_uSiiAwV32_0(.din(n22749), .dout(n22752));
    jdff dff_A_MMk7vI6F0_0(.din(n22752), .dout(n22755));
    jdff dff_A_XJfbGET98_0(.din(n22755), .dout(n22758));
    jdff dff_A_enUVeP9G1_0(.din(n22758), .dout(n22761));
    jdff dff_A_RW2z4dJ44_0(.din(n22761), .dout(n22764));
    jdff dff_A_9Cm7KGQt9_0(.din(n22764), .dout(n22767));
    jdff dff_A_BoATiG8v7_0(.din(n22767), .dout(n22770));
    jdff dff_A_65ZGevFm9_0(.din(n22770), .dout(n22773));
    jdff dff_A_URTE9TmN8_0(.din(n22773), .dout(n22776));
    jdff dff_A_HfyHt0xL1_0(.din(n22776), .dout(n22779));
    jdff dff_A_TUWilLHJ6_0(.din(n22779), .dout(n22782));
    jdff dff_A_myPRZoEq7_0(.din(n22782), .dout(n22785));
    jdff dff_A_N51r9fdv0_0(.din(n22785), .dout(n22788));
    jdff dff_A_zunUBKVQ0_0(.din(n22788), .dout(n22791));
    jdff dff_A_NX7Px3B18_0(.din(n22791), .dout(n22794));
    jdff dff_A_0eb4s6Ac5_0(.din(n22794), .dout(n22797));
    jdff dff_A_wKPSXQ9S5_0(.din(n22797), .dout(n22800));
    jdff dff_A_WS8MKiuX9_0(.din(n22800), .dout(n22803));
    jdff dff_A_HW2uTXjD8_0(.din(n22803), .dout(n22806));
    jdff dff_A_01lhwsU58_0(.din(n22806), .dout(n22809));
    jdff dff_A_UyJWuDAO7_0(.din(n22809), .dout(n22812));
    jdff dff_A_mfr6wMuy6_0(.din(n22812), .dout(G892));
    jdff dff_A_YrcMuZjh5_1(.din(n5783), .dout(n22818));
    jdff dff_A_jhEr5zGS5_0(.din(n22818), .dout(n22821));
    jdff dff_A_vjbUvAEs7_0(.din(n22821), .dout(n22824));
    jdff dff_A_yLelHxPb9_0(.din(n22824), .dout(n22827));
    jdff dff_A_ZDCQfVVY7_0(.din(n22827), .dout(n22830));
    jdff dff_A_CXROt8NI0_0(.din(n22830), .dout(n22833));
    jdff dff_A_u0KRek7n0_0(.din(n22833), .dout(n22836));
    jdff dff_A_sB0yXDSc6_0(.din(n22836), .dout(n22839));
    jdff dff_A_fiLpjyuf1_0(.din(n22839), .dout(n22842));
    jdff dff_A_rUUSTHGH2_0(.din(n22842), .dout(n22845));
    jdff dff_A_WLXMhlYe7_0(.din(n22845), .dout(n22848));
    jdff dff_A_mN1szGLP0_0(.din(n22848), .dout(n22851));
    jdff dff_A_kulQlXRO5_0(.din(n22851), .dout(n22854));
    jdff dff_A_iiseMS9g5_0(.din(n22854), .dout(n22857));
    jdff dff_A_q4JDALdd1_0(.din(n22857), .dout(n22860));
    jdff dff_A_Ld6FerP87_0(.din(n22860), .dout(n22863));
    jdff dff_A_rlfMbOL13_0(.din(n22863), .dout(n22866));
    jdff dff_A_3pIkzwlY5_0(.din(n22866), .dout(n22869));
    jdff dff_A_CSqsZH544_0(.din(n22869), .dout(n22872));
    jdff dff_A_XX0lVAs04_0(.din(n22872), .dout(n22875));
    jdff dff_A_5ljnhUSX1_0(.din(n22875), .dout(n22878));
    jdff dff_A_9wXbLuQx4_0(.din(n22878), .dout(n22881));
    jdff dff_A_Mj3Yn2ok4_0(.din(n22881), .dout(n22884));
    jdff dff_A_gKOno9Oj4_0(.din(n22884), .dout(n22887));
    jdff dff_A_UIzerzom4_0(.din(n22887), .dout(n22890));
    jdff dff_A_mSOx0lHj4_0(.din(n22890), .dout(n22893));
    jdff dff_A_8xdMCJWG0_0(.din(n22893), .dout(G887));
    jdff dff_A_i0f25SsS5_1(.din(n5786), .dout(n22899));
    jdff dff_A_EaoC9uBY9_0(.din(n22899), .dout(n22902));
    jdff dff_A_SSYifb0q5_0(.din(n22902), .dout(n22905));
    jdff dff_A_fxEzwhkz5_0(.din(n22905), .dout(n22908));
    jdff dff_A_gImH4YvO7_0(.din(n22908), .dout(n22911));
    jdff dff_A_mx8rY8fB6_0(.din(n22911), .dout(n22914));
    jdff dff_A_BjcwPdQA4_0(.din(n22914), .dout(n22917));
    jdff dff_A_pPx2SNbI8_0(.din(n22917), .dout(n22920));
    jdff dff_A_uyXOxEBR7_0(.din(n22920), .dout(n22923));
    jdff dff_A_8rO5yTEq1_0(.din(n22923), .dout(n22926));
    jdff dff_A_w57orzIn7_0(.din(n22926), .dout(n22929));
    jdff dff_A_ob5EmfXZ0_0(.din(n22929), .dout(n22932));
    jdff dff_A_vJT2ArS15_0(.din(n22932), .dout(n22935));
    jdff dff_A_5iai8qls3_0(.din(n22935), .dout(n22938));
    jdff dff_A_UxVvbBJv4_0(.din(n22938), .dout(n22941));
    jdff dff_A_XRKPOS2V9_0(.din(n22941), .dout(n22944));
    jdff dff_A_Vcg7Vzz66_0(.din(n22944), .dout(n22947));
    jdff dff_A_z3FQ501J3_0(.din(n22947), .dout(n22950));
    jdff dff_A_wtDX4HwP1_0(.din(n22950), .dout(n22953));
    jdff dff_A_iR93SuQP7_0(.din(n22953), .dout(n22956));
    jdff dff_A_AqdjrelI3_0(.din(n22956), .dout(n22959));
    jdff dff_A_VHv4GM3C5_0(.din(n22959), .dout(n22962));
    jdff dff_A_H8DPBpjF6_0(.din(n22962), .dout(n22965));
    jdff dff_A_VJ3md6VJ3_0(.din(n22965), .dout(n22968));
    jdff dff_A_tzFXcQsT8_0(.din(n22968), .dout(n22971));
    jdff dff_A_3mgvfYY55_0(.din(n22971), .dout(n22974));
    jdff dff_A_Tt7Kreo86_0(.din(n22974), .dout(G606));
    jdff dff_A_pkH3YkUJ5_2(.din(n377), .dout(n22980));
    jdff dff_A_bVproxhZ1_0(.din(n22980), .dout(n22983));
    jdff dff_A_NnggmJRV8_0(.din(n22983), .dout(n22986));
    jdff dff_A_Dtng7xtL1_0(.din(n22986), .dout(n22989));
    jdff dff_A_VzWPLMQo1_0(.din(n22989), .dout(n22992));
    jdff dff_A_5peywzLZ3_0(.din(n22992), .dout(n22995));
    jdff dff_A_FknypKjz8_0(.din(n22995), .dout(n22998));
    jdff dff_A_zYJzvywN2_0(.din(n22998), .dout(n23001));
    jdff dff_A_8d2IWV7w7_0(.din(n23001), .dout(n23004));
    jdff dff_A_syANXWzw9_0(.din(n23004), .dout(n23007));
    jdff dff_A_mQRD1Het5_0(.din(n23007), .dout(n23010));
    jdff dff_A_oz7vJrKv5_0(.din(n23010), .dout(n23013));
    jdff dff_A_2gabycod7_0(.din(n23013), .dout(n23016));
    jdff dff_A_RLZewH0M7_0(.din(n23016), .dout(n23019));
    jdff dff_A_SQ4fMz7y7_0(.din(n23019), .dout(n23022));
    jdff dff_A_P9lMhNpW4_0(.din(n23022), .dout(n23025));
    jdff dff_A_SbWgZuYa5_0(.din(n23025), .dout(n23028));
    jdff dff_A_3p5gu8aV5_0(.din(n23028), .dout(n23031));
    jdff dff_A_XlJ7iejh3_0(.din(n23031), .dout(n23034));
    jdff dff_A_LyygyGZP6_0(.din(n23034), .dout(n23037));
    jdff dff_A_n6ByNeGz2_0(.din(n23037), .dout(n23040));
    jdff dff_A_4Uq4ytKh1_0(.din(n23040), .dout(n23043));
    jdff dff_A_C9Nwdp014_0(.din(n23043), .dout(n23046));
    jdff dff_A_EpQxD4l68_0(.din(n23046), .dout(n23049));
    jdff dff_A_LcbV2KB71_0(.din(n23049), .dout(G656));
    jdff dff_A_f2GSdHvr4_2(.din(n373), .dout(n23055));
    jdff dff_A_4GI2vdTM9_0(.din(n23055), .dout(n23058));
    jdff dff_A_9DPRFH3j1_0(.din(n23058), .dout(n23061));
    jdff dff_A_brnb3pLh2_0(.din(n23061), .dout(n23064));
    jdff dff_A_4LTPbnYX6_0(.din(n23064), .dout(n23067));
    jdff dff_A_432jsq1W8_0(.din(n23067), .dout(n23070));
    jdff dff_A_Nv5oegAo6_0(.din(n23070), .dout(n23073));
    jdff dff_A_l7UkE0E24_0(.din(n23073), .dout(n23076));
    jdff dff_A_E7QuBlZJ4_0(.din(n23076), .dout(n23079));
    jdff dff_A_TwXQ17uT1_0(.din(n23079), .dout(n23082));
    jdff dff_A_orOK3QiK0_0(.din(n23082), .dout(n23085));
    jdff dff_A_OqWgzCzh6_0(.din(n23085), .dout(n23088));
    jdff dff_A_ck27aEon9_0(.din(n23088), .dout(n23091));
    jdff dff_A_LlKry5MB5_0(.din(n23091), .dout(n23094));
    jdff dff_A_GvQS4EHy0_0(.din(n23094), .dout(n23097));
    jdff dff_A_k3ETe60u0_0(.din(n23097), .dout(n23100));
    jdff dff_A_mY05oQWp8_0(.din(n23100), .dout(n23103));
    jdff dff_A_txr2TGNJ1_0(.din(n23103), .dout(n23106));
    jdff dff_A_HhBUpIvU3_0(.din(n23106), .dout(n23109));
    jdff dff_A_RmNhbpNS3_0(.din(n23109), .dout(n23112));
    jdff dff_A_KJrxWuKz7_0(.din(n23112), .dout(n23115));
    jdff dff_A_ab98WgBp3_0(.din(n23115), .dout(n23118));
    jdff dff_A_FEs7AWUG6_0(.din(n23118), .dout(n23121));
    jdff dff_A_BmlfKb2Z0_0(.din(n23121), .dout(n23124));
    jdff dff_A_5zh3mgN75_0(.din(n23124), .dout(n23127));
    jdff dff_A_t57oU9fo7_0(.din(n23127), .dout(G809));
    jdff dff_A_jBXFRELh6_1(.din(n5789), .dout(n23133));
    jdff dff_A_O4279mhi6_0(.din(n23133), .dout(n23136));
    jdff dff_A_gkLomz2O2_0(.din(n23136), .dout(n23139));
    jdff dff_A_5IO90M1b1_0(.din(n23139), .dout(n23142));
    jdff dff_A_w25WQnhG5_0(.din(n23142), .dout(n23145));
    jdff dff_A_Al5wD0XM5_0(.din(n23145), .dout(n23148));
    jdff dff_A_WUt9Obbs2_0(.din(n23148), .dout(n23151));
    jdff dff_A_IEARGc4p8_0(.din(n23151), .dout(n23154));
    jdff dff_A_oCdrQpEF4_0(.din(n23154), .dout(n23157));
    jdff dff_A_0P59qezH7_0(.din(n23157), .dout(n23160));
    jdff dff_A_tf3dk7eV5_0(.din(n23160), .dout(n23163));
    jdff dff_A_eU0hxtQK5_0(.din(n23163), .dout(n23166));
    jdff dff_A_J8ltMfCs6_0(.din(n23166), .dout(n23169));
    jdff dff_A_qO1vkvcG9_0(.din(n23169), .dout(n23172));
    jdff dff_A_xSu0o2Jz4_0(.din(n23172), .dout(n23175));
    jdff dff_A_m7EMncmL0_0(.din(n23175), .dout(n23178));
    jdff dff_A_rbuAS3CU6_0(.din(n23178), .dout(n23181));
    jdff dff_A_7Z6O8Y0J9_0(.din(n23181), .dout(n23184));
    jdff dff_A_WX9bIBWT6_0(.din(n23184), .dout(n23187));
    jdff dff_A_cIln2rmy5_0(.din(n23187), .dout(n23190));
    jdff dff_A_Rrj2gw9F6_0(.din(n23190), .dout(n23193));
    jdff dff_A_F36pxWCQ3_0(.din(n23193), .dout(n23196));
    jdff dff_A_kEDOBLfu4_0(.din(n23196), .dout(n23199));
    jdff dff_A_loYdKfFg6_0(.din(n23199), .dout(n23202));
    jdff dff_A_nO5ramgs1_0(.din(n23202), .dout(n23205));
    jdff dff_A_xxC0s3NU1_0(.din(n23205), .dout(n23208));
    jdff dff_A_x4ak0bCm9_0(.din(n23208), .dout(G993));
    jdff dff_A_AOkWbxaA9_1(.din(n5792), .dout(n23214));
    jdff dff_A_UrKL7IBP3_0(.din(n23214), .dout(n23217));
    jdff dff_A_OCoDPrgc0_0(.din(n23217), .dout(n23220));
    jdff dff_A_ID8Ltcb10_0(.din(n23220), .dout(n23223));
    jdff dff_A_Mz87F2Wy8_0(.din(n23223), .dout(n23226));
    jdff dff_A_HspfVHHf7_0(.din(n23226), .dout(n23229));
    jdff dff_A_zX0zbdhB7_0(.din(n23229), .dout(n23232));
    jdff dff_A_DlXVKrQM3_0(.din(n23232), .dout(n23235));
    jdff dff_A_og3hDeDi0_0(.din(n23235), .dout(n23238));
    jdff dff_A_Y8uGbWbG4_0(.din(n23238), .dout(n23241));
    jdff dff_A_sTDa7OYi2_0(.din(n23241), .dout(n23244));
    jdff dff_A_eWh4NSQ39_0(.din(n23244), .dout(n23247));
    jdff dff_A_BXFX4jj31_0(.din(n23247), .dout(n23250));
    jdff dff_A_Jnkop36Y9_0(.din(n23250), .dout(n23253));
    jdff dff_A_Vmxipy6w2_0(.din(n23253), .dout(n23256));
    jdff dff_A_Ok8Y0cGv1_0(.din(n23256), .dout(n23259));
    jdff dff_A_uwv5k4xR7_0(.din(n23259), .dout(n23262));
    jdff dff_A_qADDLnHx0_0(.din(n23262), .dout(n23265));
    jdff dff_A_kgcBYuEQ4_0(.din(n23265), .dout(n23268));
    jdff dff_A_rAveruXr9_0(.din(n23268), .dout(n23271));
    jdff dff_A_uQBIO8VC7_0(.din(n23271), .dout(n23274));
    jdff dff_A_WFc12DKO2_0(.din(n23274), .dout(n23277));
    jdff dff_A_Tr9ThHPu3_0(.din(n23277), .dout(n23280));
    jdff dff_A_cMjBiDnC8_0(.din(n23280), .dout(n23283));
    jdff dff_A_e5yMkLbO6_0(.din(n23283), .dout(n23286));
    jdff dff_A_NvcJmCpU8_0(.din(n23286), .dout(n23289));
    jdff dff_A_bBfrkhR76_0(.din(n23289), .dout(G978));
    jdff dff_A_8UBzqmtz1_1(.din(n5795), .dout(n23295));
    jdff dff_A_xAMmuwKd7_0(.din(n23295), .dout(n23298));
    jdff dff_A_FCy7xAyr4_0(.din(n23298), .dout(n23301));
    jdff dff_A_hiaAwhs56_0(.din(n23301), .dout(n23304));
    jdff dff_A_9aQqzs390_0(.din(n23304), .dout(n23307));
    jdff dff_A_V4O7HvQ07_0(.din(n23307), .dout(n23310));
    jdff dff_A_6dOjmLPT6_0(.din(n23310), .dout(n23313));
    jdff dff_A_RArkxi7X6_0(.din(n23313), .dout(n23316));
    jdff dff_A_lryukamR8_0(.din(n23316), .dout(n23319));
    jdff dff_A_a6ocVgTp5_0(.din(n23319), .dout(n23322));
    jdff dff_A_HnBEWdAw3_0(.din(n23322), .dout(n23325));
    jdff dff_A_dJ5c2YAM4_0(.din(n23325), .dout(n23328));
    jdff dff_A_RZhauPO90_0(.din(n23328), .dout(n23331));
    jdff dff_A_cFFHib127_0(.din(n23331), .dout(n23334));
    jdff dff_A_7QR5pUC97_0(.din(n23334), .dout(n23337));
    jdff dff_A_YP6GqKyh1_0(.din(n23337), .dout(n23340));
    jdff dff_A_Z3yLKJJr0_0(.din(n23340), .dout(n23343));
    jdff dff_A_n8oRfgRV9_0(.din(n23343), .dout(n23346));
    jdff dff_A_0l0E9Php1_0(.din(n23346), .dout(n23349));
    jdff dff_A_JOz6Y5zA2_0(.din(n23349), .dout(n23352));
    jdff dff_A_xgNSg37t8_0(.din(n23352), .dout(n23355));
    jdff dff_A_MDeAfenL1_0(.din(n23355), .dout(n23358));
    jdff dff_A_IUkC6Joo2_0(.din(n23358), .dout(n23361));
    jdff dff_A_b3V2Ghm33_0(.din(n23361), .dout(n23364));
    jdff dff_A_yvOhH7523_0(.din(n23364), .dout(n23367));
    jdff dff_A_t2vfrKCz6_0(.din(n23367), .dout(n23370));
    jdff dff_A_BoOOBYC89_0(.din(n23370), .dout(G949));
    jdff dff_A_SKPLdeyi8_1(.din(n5798), .dout(n23376));
    jdff dff_A_2qSTzhyE9_0(.din(n23376), .dout(n23379));
    jdff dff_A_nucsXvpf2_0(.din(n23379), .dout(n23382));
    jdff dff_A_pJq5yQqh4_0(.din(n23382), .dout(n23385));
    jdff dff_A_wu97i3l88_0(.din(n23385), .dout(n23388));
    jdff dff_A_5S0JHsZ41_0(.din(n23388), .dout(n23391));
    jdff dff_A_z7kyIMWU7_0(.din(n23391), .dout(n23394));
    jdff dff_A_PDVDedOh3_0(.din(n23394), .dout(n23397));
    jdff dff_A_WVwJhwtm7_0(.din(n23397), .dout(n23400));
    jdff dff_A_YwIrpcYa1_0(.din(n23400), .dout(n23403));
    jdff dff_A_xHz7VYgs1_0(.din(n23403), .dout(n23406));
    jdff dff_A_jXAdoxY40_0(.din(n23406), .dout(n23409));
    jdff dff_A_OmOWHH8i7_0(.din(n23409), .dout(n23412));
    jdff dff_A_u15K7vWv4_0(.din(n23412), .dout(n23415));
    jdff dff_A_tLPxEEPG4_0(.din(n23415), .dout(n23418));
    jdff dff_A_SalfHBKp8_0(.din(n23418), .dout(n23421));
    jdff dff_A_X20frKLI7_0(.din(n23421), .dout(n23424));
    jdff dff_A_ZA4oBV7I1_0(.din(n23424), .dout(n23427));
    jdff dff_A_keFdkTBZ4_0(.din(n23427), .dout(n23430));
    jdff dff_A_wH64j8n76_0(.din(n23430), .dout(n23433));
    jdff dff_A_qrSLvkpL6_0(.din(n23433), .dout(n23436));
    jdff dff_A_23jIzKqa0_0(.din(n23436), .dout(n23439));
    jdff dff_A_xymuw4o74_0(.din(n23439), .dout(n23442));
    jdff dff_A_pD3W7Z586_0(.din(n23442), .dout(n23445));
    jdff dff_A_JFYKppkd0_0(.din(n23445), .dout(n23448));
    jdff dff_A_CcltRsG24_0(.din(n23448), .dout(n23451));
    jdff dff_A_B2DvfHSf5_0(.din(n23451), .dout(G939));
    jdff dff_A_Femo9NLV5_1(.din(n5801), .dout(n23457));
    jdff dff_A_NlHBCzV31_0(.din(n23457), .dout(n23460));
    jdff dff_A_wg5gnJ2k1_0(.din(n23460), .dout(n23463));
    jdff dff_A_P479h9P96_0(.din(n23463), .dout(n23466));
    jdff dff_A_HqpFnqCb7_0(.din(n23466), .dout(n23469));
    jdff dff_A_PvnhAJg39_0(.din(n23469), .dout(n23472));
    jdff dff_A_LZll5Fm78_0(.din(n23472), .dout(n23475));
    jdff dff_A_0z4SIJqg6_0(.din(n23475), .dout(n23478));
    jdff dff_A_IFWuuGx01_0(.din(n23478), .dout(n23481));
    jdff dff_A_XSxmljR30_0(.din(n23481), .dout(n23484));
    jdff dff_A_BrKoEwES3_0(.din(n23484), .dout(n23487));
    jdff dff_A_rYEawTOG9_0(.din(n23487), .dout(n23490));
    jdff dff_A_a7fR5RQd1_0(.din(n23490), .dout(n23493));
    jdff dff_A_4IOJGG5X4_0(.din(n23493), .dout(n23496));
    jdff dff_A_W9iTcZTk2_0(.din(n23496), .dout(n23499));
    jdff dff_A_65rT7D2V2_0(.din(n23499), .dout(n23502));
    jdff dff_A_FswOCQ1x5_0(.din(n23502), .dout(n23505));
    jdff dff_A_rr1mzzEm5_0(.din(n23505), .dout(n23508));
    jdff dff_A_LzvWqzG99_0(.din(n23508), .dout(n23511));
    jdff dff_A_qHF1pcbb0_0(.din(n23511), .dout(n23514));
    jdff dff_A_OUaEY0X33_0(.din(n23514), .dout(n23517));
    jdff dff_A_0iAljFpq4_0(.din(n23517), .dout(n23520));
    jdff dff_A_YPIditjM1_0(.din(n23520), .dout(n23523));
    jdff dff_A_EN3CGhBf4_0(.din(n23523), .dout(n23526));
    jdff dff_A_W6UzBvUa9_0(.din(n23526), .dout(n23529));
    jdff dff_A_0gxnXOPP4_0(.din(n23529), .dout(n23532));
    jdff dff_A_0NxvzrgN0_0(.din(n23532), .dout(G889));
    jdff dff_A_JlUsfOTy7_1(.din(n380), .dout(n23538));
    jdff dff_A_3B9HwBPe0_0(.din(n23538), .dout(n23541));
    jdff dff_A_yStGtaew4_0(.din(n23541), .dout(n23544));
    jdff dff_A_jaLX8CQ02_0(.din(n23544), .dout(n23547));
    jdff dff_A_67wNSxP11_0(.din(n23547), .dout(n23550));
    jdff dff_A_GegosreC5_0(.din(n23550), .dout(n23553));
    jdff dff_A_XHWoNeFP3_0(.din(n23553), .dout(n23556));
    jdff dff_A_bLfiJvCO4_0(.din(n23556), .dout(n23559));
    jdff dff_A_BS0uVRY25_0(.din(n23559), .dout(n23562));
    jdff dff_A_kVvwKqRh3_0(.din(n23562), .dout(n23565));
    jdff dff_A_XGBQ3QtX9_0(.din(n23565), .dout(n23568));
    jdff dff_A_MMY6qRtf4_0(.din(n23568), .dout(n23571));
    jdff dff_A_j4alQXXo8_0(.din(n23571), .dout(n23574));
    jdff dff_A_riaw58ne8_0(.din(n23574), .dout(n23577));
    jdff dff_A_MN2uMMIk9_0(.din(n23577), .dout(n23580));
    jdff dff_A_XRWpcieE0_0(.din(n23580), .dout(n23583));
    jdff dff_A_0IZ2WCww9_0(.din(n23583), .dout(n23586));
    jdff dff_A_jKIJe3Cs1_0(.din(n23586), .dout(n23589));
    jdff dff_A_Eon0llJ00_0(.din(n23589), .dout(n23592));
    jdff dff_A_I302w8E71_0(.din(n23592), .dout(n23595));
    jdff dff_A_WbLeyYaB7_0(.din(n23595), .dout(n23598));
    jdff dff_A_WkftCjGB1_0(.din(n23598), .dout(n23601));
    jdff dff_A_mPYVDaIn7_0(.din(n23601), .dout(n23604));
    jdff dff_A_rzLVcdgv7_0(.din(n23604), .dout(n23607));
    jdff dff_A_xL5DAQUP6_0(.din(n23607), .dout(n23610));
    jdff dff_A_iTB1BQ4n3_0(.din(n23610), .dout(n23613));
    jdff dff_A_lzRGMTWg1_0(.din(n23613), .dout(G593));
    jdff dff_A_ggxnG5mk7_2(.din(n405), .dout(n23619));
    jdff dff_A_soGqoBSU8_0(.din(n23619), .dout(n23622));
    jdff dff_A_a0JslDTl1_0(.din(n23622), .dout(n23625));
    jdff dff_A_zpTnZla65_0(.din(n23625), .dout(n23628));
    jdff dff_A_tTRpNvXs0_0(.din(n23628), .dout(n23631));
    jdff dff_A_bjOdwmAc2_0(.din(n23631), .dout(n23634));
    jdff dff_A_YJ9ZAu3J6_0(.din(n23634), .dout(n23637));
    jdff dff_A_PixvskVl1_0(.din(n23637), .dout(n23640));
    jdff dff_A_p3qbVq8r3_0(.din(n23640), .dout(n23643));
    jdff dff_A_aW56xJAs5_0(.din(n23643), .dout(n23646));
    jdff dff_A_3Wlp8vE85_0(.din(n23646), .dout(n23649));
    jdff dff_A_E8mM1muW5_0(.din(n23649), .dout(n23652));
    jdff dff_A_SLFWPjY44_0(.din(n23652), .dout(n23655));
    jdff dff_A_J8kL7Sgt9_0(.din(n23655), .dout(n23658));
    jdff dff_A_sw8PUaHd1_0(.din(n23658), .dout(n23661));
    jdff dff_A_KIuylHh73_0(.din(n23661), .dout(n23664));
    jdff dff_A_sHYEi02l3_0(.din(n23664), .dout(n23667));
    jdff dff_A_yUvjfvIO8_0(.din(n23667), .dout(n23670));
    jdff dff_A_px2WHpYM5_0(.din(n23670), .dout(n23673));
    jdff dff_A_zRF8JdTh0_0(.din(n23673), .dout(n23676));
    jdff dff_A_9DUo6PBV2_0(.din(n23676), .dout(n23679));
    jdff dff_A_sgrLK5Oe7_0(.din(n23679), .dout(n23682));
    jdff dff_A_8zEUF1Kx6_0(.din(n23682), .dout(n23685));
    jdff dff_A_r5BCFrqL9_0(.din(n23685), .dout(G636));
    jdff dff_A_9Fp90GiW7_2(.din(n427), .dout(n23691));
    jdff dff_A_wkmp6lrl8_0(.din(n23691), .dout(n23694));
    jdff dff_A_Om9gIXYj8_0(.din(n23694), .dout(n23697));
    jdff dff_A_J8bKEIoc2_0(.din(n23697), .dout(n23700));
    jdff dff_A_1IR9LRMQ0_0(.din(n23700), .dout(n23703));
    jdff dff_A_Q27Pe5oZ8_0(.din(n23703), .dout(n23706));
    jdff dff_A_pmrRKuYQ3_0(.din(n23706), .dout(n23709));
    jdff dff_A_HZstU9Dd0_0(.din(n23709), .dout(n23712));
    jdff dff_A_3MOpmkng3_0(.din(n23712), .dout(n23715));
    jdff dff_A_zYDO4QhQ1_0(.din(n23715), .dout(n23718));
    jdff dff_A_CgGxoC2F7_0(.din(n23718), .dout(n23721));
    jdff dff_A_qWBRdyc79_0(.din(n23721), .dout(n23724));
    jdff dff_A_D1H3cY1Z2_0(.din(n23724), .dout(n23727));
    jdff dff_A_0l9AKiTB8_0(.din(n23727), .dout(n23730));
    jdff dff_A_XEqDzIra2_0(.din(n23730), .dout(n23733));
    jdff dff_A_SWGWLOGt5_0(.din(n23733), .dout(n23736));
    jdff dff_A_g2POdUbn9_0(.din(n23736), .dout(n23739));
    jdff dff_A_n3wg9EoG8_0(.din(n23739), .dout(n23742));
    jdff dff_A_tk4VvaVL2_0(.din(n23742), .dout(n23745));
    jdff dff_A_ViiQ19Ro7_0(.din(n23745), .dout(n23748));
    jdff dff_A_snizAxlQ4_0(.din(n23748), .dout(n23751));
    jdff dff_A_gQzsw8tX0_0(.din(n23751), .dout(n23754));
    jdff dff_A_ySsGHG3o4_0(.din(n23754), .dout(n23757));
    jdff dff_A_eJEs7m0C0_0(.din(n23757), .dout(G704));
    jdff dff_A_BaD8i8TF9_2(.din(n5805), .dout(n23763));
    jdff dff_A_xjBKTD4I1_0(.din(n23763), .dout(n23766));
    jdff dff_A_6YM20goG0_0(.din(n23766), .dout(n23769));
    jdff dff_A_MElF77n31_0(.din(n23769), .dout(n23772));
    jdff dff_A_xDGqj1qa7_0(.din(n23772), .dout(n23775));
    jdff dff_A_gMJ0bC1b7_0(.din(n23775), .dout(n23778));
    jdff dff_A_OZD5cGSG7_0(.din(n23778), .dout(n23781));
    jdff dff_A_dgKvcHDk1_0(.din(n23781), .dout(n23784));
    jdff dff_A_PqCbBv3R6_0(.din(n23784), .dout(n23787));
    jdff dff_A_fAYB8dnB5_0(.din(n23787), .dout(n23790));
    jdff dff_A_JP7SyptP2_0(.din(n23790), .dout(n23793));
    jdff dff_A_KI5jhp3e5_0(.din(n23793), .dout(n23796));
    jdff dff_A_zwuUHvm75_0(.din(n23796), .dout(n23799));
    jdff dff_A_otvnUqrg0_0(.din(n23799), .dout(n23802));
    jdff dff_A_NJ3uvGoa6_0(.din(n23802), .dout(n23805));
    jdff dff_A_3mvlPVQ53_0(.din(n23805), .dout(n23808));
    jdff dff_A_DDumhluL6_0(.din(n23808), .dout(n23811));
    jdff dff_A_8IuzqLEW7_0(.din(n23811), .dout(n23814));
    jdff dff_A_boPSc9fI5_0(.din(n23814), .dout(n23817));
    jdff dff_A_ESwuOz9u6_0(.din(n23817), .dout(n23820));
    jdff dff_A_UANjooBs1_0(.din(n23820), .dout(n23823));
    jdff dff_A_ADvYnNf58_0(.din(n23823), .dout(n23826));
    jdff dff_A_1CiA6Af43_0(.din(n23826), .dout(n23829));
    jdff dff_A_tzjUCfjA9_0(.din(n23829), .dout(G717));
    jdff dff_A_7aIGYmBt8_2(.din(n434), .dout(n23835));
    jdff dff_A_fdslbe5r7_0(.din(n23835), .dout(n23838));
    jdff dff_A_bgmIoIfr6_0(.din(n23838), .dout(n23841));
    jdff dff_A_eB9DO8Xr2_0(.din(n23841), .dout(n23844));
    jdff dff_A_FztlOzVp5_0(.din(n23844), .dout(n23847));
    jdff dff_A_GKY3LsMV0_0(.din(n23847), .dout(n23850));
    jdff dff_A_iNwDsvSD2_0(.din(n23850), .dout(n23853));
    jdff dff_A_xER18dRt8_0(.din(n23853), .dout(n23856));
    jdff dff_A_Vw79pbN41_0(.din(n23856), .dout(n23859));
    jdff dff_A_eD7oyL8r7_0(.din(n23859), .dout(n23862));
    jdff dff_A_QnfkqptZ9_0(.din(n23862), .dout(n23865));
    jdff dff_A_qkJJt8qk1_0(.din(n23865), .dout(n23868));
    jdff dff_A_v32xaZdh5_0(.din(n23868), .dout(n23871));
    jdff dff_A_EpydQUZR8_0(.din(n23871), .dout(n23874));
    jdff dff_A_oIQ15tVM3_0(.din(n23874), .dout(n23877));
    jdff dff_A_FecwbBKd7_0(.din(n23877), .dout(n23880));
    jdff dff_A_DJp5nEX43_0(.din(n23880), .dout(n23883));
    jdff dff_A_fagqzMmt2_0(.din(n23883), .dout(n23886));
    jdff dff_A_t6mYyL5t3_0(.din(n23886), .dout(n23889));
    jdff dff_A_fdUuXirF3_0(.din(n23889), .dout(n23892));
    jdff dff_A_sc2fG96P1_0(.din(n23892), .dout(n23895));
    jdff dff_A_lm5H9nBY1_0(.din(n23895), .dout(n23898));
    jdff dff_A_adDaodPF2_0(.din(n23898), .dout(n23901));
    jdff dff_A_RpYPwKbW1_0(.din(n23901), .dout(n23904));
    jdff dff_A_22ycq4ex2_0(.din(n23904), .dout(G820));
    jdff dff_A_oXh5hHFP5_2(.din(n454), .dout(n23910));
    jdff dff_A_4LtYUCoT8_0(.din(n23910), .dout(n23913));
    jdff dff_A_4iVz71ut0_0(.din(n23913), .dout(n23916));
    jdff dff_A_IWIDMaw86_0(.din(n23916), .dout(n23919));
    jdff dff_A_XkkHFvoO4_0(.din(n23919), .dout(n23922));
    jdff dff_A_IaQB31nO0_0(.din(n23922), .dout(n23925));
    jdff dff_A_CfsQocWg1_0(.din(n23925), .dout(n23928));
    jdff dff_A_eHgmuEbK1_0(.din(n23928), .dout(n23931));
    jdff dff_A_pqbmqe2y1_0(.din(n23931), .dout(n23934));
    jdff dff_A_lcQfdGmx4_0(.din(n23934), .dout(n23937));
    jdff dff_A_8QrI6YU44_0(.din(n23937), .dout(n23940));
    jdff dff_A_nX2fVv7i5_0(.din(n23940), .dout(n23943));
    jdff dff_A_2lH3SzDG5_0(.din(n23943), .dout(n23946));
    jdff dff_A_JjVnmOAe2_0(.din(n23946), .dout(n23949));
    jdff dff_A_uWwO6c0V0_0(.din(n23949), .dout(n23952));
    jdff dff_A_Scr4Xdlr9_0(.din(n23952), .dout(n23955));
    jdff dff_A_MNmT17kz0_0(.din(n23955), .dout(n23958));
    jdff dff_A_4NhZrj4o5_0(.din(n23958), .dout(n23961));
    jdff dff_A_Z3M9vFrv1_0(.din(n23961), .dout(n23964));
    jdff dff_A_HweYZHgk8_0(.din(n23964), .dout(n23967));
    jdff dff_A_yykWYldi2_0(.din(n23967), .dout(n23970));
    jdff dff_A_9OoTzEzV7_0(.din(n23970), .dout(n23973));
    jdff dff_A_Zlckauki5_0(.din(n23973), .dout(G639));
    jdff dff_A_4VBlrx7w2_2(.din(n474), .dout(n23979));
    jdff dff_A_BIlgfuI73_0(.din(n23979), .dout(n23982));
    jdff dff_A_uXeSAsFX3_0(.din(n23982), .dout(n23985));
    jdff dff_A_VomWAx9P1_0(.din(n23985), .dout(n23988));
    jdff dff_A_sRlKKdnF4_0(.din(n23988), .dout(n23991));
    jdff dff_A_duknT22U1_0(.din(n23991), .dout(n23994));
    jdff dff_A_HALbsMQM1_0(.din(n23994), .dout(n23997));
    jdff dff_A_qKlXLPIF0_0(.din(n23997), .dout(n24000));
    jdff dff_A_VXSzI9iX9_0(.din(n24000), .dout(n24003));
    jdff dff_A_xcijaDCS4_0(.din(n24003), .dout(n24006));
    jdff dff_A_5X1gZXtG7_0(.din(n24006), .dout(n24009));
    jdff dff_A_lRDBTsYm8_0(.din(n24009), .dout(n24012));
    jdff dff_A_MYOlMxxt1_0(.din(n24012), .dout(n24015));
    jdff dff_A_JdmnnDJw6_0(.din(n24015), .dout(n24018));
    jdff dff_A_Dn4OQfkn4_0(.din(n24018), .dout(n24021));
    jdff dff_A_6ygsp5KJ0_0(.din(n24021), .dout(n24024));
    jdff dff_A_rh6YIwCc6_0(.din(n24024), .dout(n24027));
    jdff dff_A_S0F2NR0R8_0(.din(n24027), .dout(n24030));
    jdff dff_A_FwX7Takh2_0(.din(n24030), .dout(n24033));
    jdff dff_A_N3KcFBa32_0(.din(n24033), .dout(n24036));
    jdff dff_A_LoEkIqHu8_0(.din(n24036), .dout(n24039));
    jdff dff_A_euh4H7FH7_0(.din(n24039), .dout(n24042));
    jdff dff_A_McPKAUHR9_0(.din(n24042), .dout(G673));
    jdff dff_A_TnyExUOt6_2(.din(n494), .dout(n24048));
    jdff dff_A_m2QxoPEi7_0(.din(n24048), .dout(n24051));
    jdff dff_A_6DCS2fUy9_0(.din(n24051), .dout(n24054));
    jdff dff_A_QxOHOkW36_0(.din(n24054), .dout(n24057));
    jdff dff_A_jyRVJxNl4_0(.din(n24057), .dout(n24060));
    jdff dff_A_BUaKj3Nn2_0(.din(n24060), .dout(n24063));
    jdff dff_A_Ti9mOnCh1_0(.din(n24063), .dout(n24066));
    jdff dff_A_VuWBPtCy4_0(.din(n24066), .dout(n24069));
    jdff dff_A_NFPZ5n9V4_0(.din(n24069), .dout(n24072));
    jdff dff_A_QyhQHejV1_0(.din(n24072), .dout(n24075));
    jdff dff_A_HtsmvrZi3_0(.din(n24075), .dout(n24078));
    jdff dff_A_T4XC26Jg7_0(.din(n24078), .dout(n24081));
    jdff dff_A_nFvlLH8c1_0(.din(n24081), .dout(n24084));
    jdff dff_A_OShEDruo9_0(.din(n24084), .dout(n24087));
    jdff dff_A_GGdVLRBB7_0(.din(n24087), .dout(n24090));
    jdff dff_A_rFgGl2NK4_0(.din(n24090), .dout(n24093));
    jdff dff_A_VahjnZhW6_0(.din(n24093), .dout(n24096));
    jdff dff_A_DEaQaxxT2_0(.din(n24096), .dout(n24099));
    jdff dff_A_gUfDPPDN6_0(.din(n24099), .dout(n24102));
    jdff dff_A_8afGv2pz2_0(.din(n24102), .dout(n24105));
    jdff dff_A_3lv0jjFW6_0(.din(n24105), .dout(n24108));
    jdff dff_A_YmzDT3ym0_0(.din(n24108), .dout(n24111));
    jdff dff_A_IfE1XxdW2_0(.din(n24111), .dout(G707));
    jdff dff_A_jviPCy004_2(.din(n514), .dout(n24117));
    jdff dff_A_04uaOXrN9_0(.din(n24117), .dout(n24120));
    jdff dff_A_UdbLiJgG5_0(.din(n24120), .dout(n24123));
    jdff dff_A_MzDfdB4P0_0(.din(n24123), .dout(n24126));
    jdff dff_A_SxgIrgyv4_0(.din(n24126), .dout(n24129));
    jdff dff_A_MHWEKNgO1_0(.din(n24129), .dout(n24132));
    jdff dff_A_WGdGq7Ey9_0(.din(n24132), .dout(n24135));
    jdff dff_A_OxGqiwtK2_0(.din(n24135), .dout(n24138));
    jdff dff_A_y1IPsVse8_0(.din(n24138), .dout(n24141));
    jdff dff_A_2B6Q3m830_0(.din(n24141), .dout(n24144));
    jdff dff_A_LX8HlE9g4_0(.din(n24144), .dout(n24147));
    jdff dff_A_xk5ejCSe6_0(.din(n24147), .dout(n24150));
    jdff dff_A_BaoSDj0W1_0(.din(n24150), .dout(n24153));
    jdff dff_A_5cs0LYHE3_0(.din(n24153), .dout(n24156));
    jdff dff_A_Ex6JadYn8_0(.din(n24156), .dout(n24159));
    jdff dff_A_fTvKbmDP0_0(.din(n24159), .dout(n24162));
    jdff dff_A_4mydeKCB9_0(.din(n24162), .dout(n24165));
    jdff dff_A_0ozEw7dI5_0(.din(n24165), .dout(n24168));
    jdff dff_A_K9IfZtmH3_0(.din(n24168), .dout(n24171));
    jdff dff_A_rJ51SNR76_0(.din(n24171), .dout(n24174));
    jdff dff_A_4YzD4k2h4_0(.din(n24174), .dout(n24177));
    jdff dff_A_dYaBkdA04_0(.din(n24177), .dout(n24180));
    jdff dff_A_u6GnkU9e7_0(.din(n24180), .dout(G715));
    jdff dff_A_FCzrs7lI1_2(.din(n846), .dout(n24186));
    jdff dff_A_ahcWene33_0(.din(n24186), .dout(n24189));
    jdff dff_A_E4ut34AA3_0(.din(n24189), .dout(n24192));
    jdff dff_A_lZiDdcn39_0(.din(n24192), .dout(n24195));
    jdff dff_A_irKjk10M5_0(.din(n24195), .dout(n24198));
    jdff dff_A_7ouXLBM22_0(.din(n24198), .dout(n24201));
    jdff dff_A_GP3KJ3lY1_0(.din(n24201), .dout(n24204));
    jdff dff_A_0rpV5NER2_0(.din(n24204), .dout(n24207));
    jdff dff_A_M6Sqze256_0(.din(n24207), .dout(n24210));
    jdff dff_A_yZ8dW7Bl7_0(.din(n24210), .dout(n24213));
    jdff dff_A_Cbq7JKkt2_0(.din(n24213), .dout(n24216));
    jdff dff_A_3zy9uUce6_0(.din(n24216), .dout(n24219));
    jdff dff_A_gLx2fgw39_0(.din(n24219), .dout(n24222));
    jdff dff_A_GvvLizGC0_0(.din(n24222), .dout(n24225));
    jdff dff_A_MfhM0JDk7_0(.din(n24225), .dout(n24228));
    jdff dff_A_yLhM6FhX1_0(.din(n24228), .dout(n24231));
    jdff dff_A_Gvzo9Uf08_0(.din(n24231), .dout(n24234));
    jdff dff_A_IOssKhkH6_0(.din(n24234), .dout(n24237));
    jdff dff_A_h5pezWX06_0(.din(n24237), .dout(n24240));
    jdff dff_A_54HgQfUU5_0(.din(n24240), .dout(G598));
    jdff dff_A_w6ptbcNI1_2(.din(n1256), .dout(n24246));
    jdff dff_A_wKcYnG6L0_0(.din(n24246), .dout(n24249));
    jdff dff_A_WLfds1zs2_0(.din(n24249), .dout(n24252));
    jdff dff_A_t8op28g67_0(.din(n24252), .dout(n24255));
    jdff dff_A_JHfpfx4h0_0(.din(n24255), .dout(n24258));
    jdff dff_A_2RMLKFdb4_0(.din(n24258), .dout(n24261));
    jdff dff_A_DDD1tYNc4_0(.din(n24261), .dout(n24264));
    jdff dff_A_s0hmulKZ0_0(.din(n24264), .dout(n24267));
    jdff dff_A_A9p0smSx1_0(.din(n24267), .dout(n24270));
    jdff dff_A_Cj9sbDPR6_0(.din(n24270), .dout(n24273));
    jdff dff_A_Kod3pKDV5_0(.din(n24273), .dout(n24276));
    jdff dff_A_7xhQmYh16_0(.din(n24276), .dout(n24279));
    jdff dff_A_vG0ZTohM3_0(.din(n24279), .dout(n24282));
    jdff dff_A_QvoG1XTB6_0(.din(n24282), .dout(n24285));
    jdff dff_A_e1pzCSdJ9_0(.din(n24285), .dout(n24288));
    jdff dff_A_CzWkz3IL9_0(.din(n24288), .dout(n24291));
    jdff dff_A_bhbvxTPo5_0(.din(n24291), .dout(n24294));
    jdff dff_A_YBZbAwDs7_0(.din(n24294), .dout(n24297));
    jdff dff_A_bi0nBdus6_0(.din(n24297), .dout(G610));
    jdff dff_A_hjs3pf4K4_2(.din(n1471), .dout(n24303));
    jdff dff_A_xktMmrAI2_0(.din(n24303), .dout(n24306));
    jdff dff_A_B0XsbOgY5_0(.din(n24306), .dout(n24309));
    jdff dff_A_hSHgTJH43_0(.din(n24309), .dout(n24312));
    jdff dff_A_bhUEti0a3_0(.din(n24312), .dout(n24315));
    jdff dff_A_LFUSm4GD1_0(.din(n24315), .dout(n24318));
    jdff dff_A_uUDNsvUN0_0(.din(n24318), .dout(n24321));
    jdff dff_A_ypLymG1f1_0(.din(n24321), .dout(n24324));
    jdff dff_A_Wl3MkFn20_0(.din(n24324), .dout(n24327));
    jdff dff_A_JT2tdUVw6_0(.din(n24327), .dout(n24330));
    jdff dff_A_OHzqKTJu2_0(.din(n24330), .dout(n24333));
    jdff dff_A_Kmwsm5hn3_0(.din(n24333), .dout(n24336));
    jdff dff_A_1hSgZx2J6_0(.din(n24336), .dout(n24339));
    jdff dff_A_mtPWx4Va4_0(.din(n24339), .dout(n24342));
    jdff dff_A_DmnnXYYn4_0(.din(n24342), .dout(n24345));
    jdff dff_A_UJa8BsNY4_0(.din(n24345), .dout(n24348));
    jdff dff_A_l2uks8bl3_0(.din(n24348), .dout(G588));
    jdff dff_A_QVvvToBY8_2(.din(n1664), .dout(n24354));
    jdff dff_A_r8UDSSn76_0(.din(n24354), .dout(n24357));
    jdff dff_A_6fgyXfer9_0(.din(n24357), .dout(n24360));
    jdff dff_A_zTl1PCT15_0(.din(n24360), .dout(n24363));
    jdff dff_A_favJvT4u8_0(.din(n24363), .dout(n24366));
    jdff dff_A_udDgwovk2_0(.din(n24366), .dout(n24369));
    jdff dff_A_fikQLPbe8_0(.din(n24369), .dout(n24372));
    jdff dff_A_QRgNZbL06_0(.din(n24372), .dout(n24375));
    jdff dff_A_A1BnklJE4_0(.din(n24375), .dout(n24378));
    jdff dff_A_ZOKzsVmy0_0(.din(n24378), .dout(n24381));
    jdff dff_A_L6JCwsmY9_0(.din(n24381), .dout(n24384));
    jdff dff_A_VdTOdjVu4_0(.din(n24384), .dout(n24387));
    jdff dff_A_1haxGdVJ2_0(.din(n24387), .dout(n24390));
    jdff dff_A_wZD9eGAg9_0(.din(n24390), .dout(n24393));
    jdff dff_A_Kvt6v9Sw6_0(.din(n24393), .dout(n24396));
    jdff dff_A_6Glt6atn6_0(.din(n24396), .dout(n24399));
    jdff dff_A_bzvNBOYj0_0(.din(n24399), .dout(n24402));
    jdff dff_A_6BM5FR752_0(.din(n24402), .dout(G615));
    jdff dff_A_VyRNnbsR6_2(.din(n5809), .dout(n24408));
    jdff dff_A_8v0iwfKN0_0(.din(n24408), .dout(n24411));
    jdff dff_A_5c3an98c5_0(.din(n24411), .dout(n24414));
    jdff dff_A_eP0RgtWU9_0(.din(n24414), .dout(n24417));
    jdff dff_A_2lkPwFN80_0(.din(n24417), .dout(n24420));
    jdff dff_A_ara8B4DS4_0(.din(n24420), .dout(n24423));
    jdff dff_A_JkxiWNce1_0(.din(n24423), .dout(n24426));
    jdff dff_A_yo4P0xeu7_0(.din(n24426), .dout(n24429));
    jdff dff_A_5BWg8Psx7_0(.din(n24429), .dout(n24432));
    jdff dff_A_c08IIq7k5_0(.din(n24432), .dout(n24435));
    jdff dff_A_vjE7kXum4_0(.din(n24435), .dout(n24438));
    jdff dff_A_OACUKO5e1_0(.din(n24438), .dout(n24441));
    jdff dff_A_EIFAbSCw3_0(.din(n24441), .dout(n24444));
    jdff dff_A_Uns95WFP8_0(.din(n24444), .dout(n24447));
    jdff dff_A_ywLwuiAb9_0(.din(n24447), .dout(n24450));
    jdff dff_A_dQbOsoUn7_0(.din(n24450), .dout(n24453));
    jdff dff_A_y1Id65Fp3_0(.din(n24453), .dout(n24456));
endmodule

