module gf_c7552(G4528, G4526, G4432, G4427, G4420, G4410, G4405, G4400, G3743, G3729, G3723, G3717, G3711, G3701, G3698, G3705, G2256, G2253, G2247, G2236, G2230, G2204, G1492, G1486, G1455, G1197, G339, G240, G239, G4393, G238, G234, G231, G228, G2239, G225, G2224, G221, G220, G219, G218, G217, G214, G236, G210, G208, G207, G209, G206, G205, G204, G1496, G203, G111, G202, G152, G100, G2218, G161, G97, G88, G223, G87, G118, G233, G53, G3749, G212, G84, G4415, G5, G222, G83, G226, G81, G82, G144, G227, G79, G64, G159, G94, G211, G66, G127, G230, G15, G61, G110, G196, G26, G23, G63, G4394, G78, G12, G62, G156, G73, G18, G9, G1459, G135, G198, G188, G199, G113, G76, G57, G237, G164, G59, G224, G35, G158, G41, G80, G55, G192, G229, G85, G114, G29, G77, G160, G75, G54, G1469, G153, G232, G194, G106, G65, G109, G216, G115, G121, G167, G124, G138, G130, G186, G4437, G200, G170, G134, G1462, G141, G150, G151, G47, G174, G154, G3737, G215, G155, G133, G185, G162, G58, G163, G165, G60, G166, G1480, G147, G168, G44, G1, G56, G169, G171, G2211, G157, G172, G2208, G193, G197, G173, G86, G175, G89, G50, G189, G213, G176, G38, G178, G179, G74, G180, G181, G69, G182, G183, G177, G184, G103, G32, G187, G112, G191, G235, G190, G195, G70, G201, G399, G370, G338, G321, G368, G362, G359, G471, G422, G344, G307, G304, G301, G273, G336, G333, G419, G327, G310, G276, G252, G295, G249, G416, G412, G382, G319, G379, G376, G365, G397, G353, G347, G394, G391, G388, G281, G330, G552, G316, G534, G554, G546, G530, G438, G270, G450, G432, G540, G418, G3, G448, G350, G484, G558, G482, G480, G404, G550, G494, G469, G524, G522, G298, G538, G442, G246, G258, G492, G548, G556, G440, G486, G544, G536, G313, G490, G542, G292, G414, G560, G528, G496, G532, G279, G526, G436, G488, G478, G324, G444, G402, G453, G278, G410, G2, G284, G408, G446, G373, G406, G264, G385, G286, G289, G356, G341);
    input G4528, G4526, G4432, G4427, G4420, G4410, G4405, G4400, G3743, G3729, G3723, G3717, G3711, G3701, G3698, G3705, G2256, G2253, G2247, G2236, G2230, G2204, G1492, G1486, G1455, G1197, G339, G240, G239, G4393, G238, G234, G231, G228, G2239, G225, G2224, G221, G220, G219, G218, G217, G214, G236, G210, G208, G207, G209, G206, G205, G204, G1496, G203, G111, G202, G152, G100, G2218, G161, G97, G88, G223, G87, G118, G233, G53, G3749, G212, G84, G4415, G5, G222, G83, G226, G81, G82, G144, G227, G79, G64, G159, G94, G211, G66, G127, G230, G15, G61, G110, G196, G26, G23, G63, G4394, G78, G12, G62, G156, G73, G18, G9, G1459, G135, G198, G188, G199, G113, G76, G57, G237, G164, G59, G224, G35, G158, G41, G80, G55, G192, G229, G85, G114, G29, G77, G160, G75, G54, G1469, G153, G232, G194, G106, G65, G109, G216, G115, G121, G167, G124, G138, G130, G186, G4437, G200, G170, G134, G1462, G141, G150, G151, G47, G174, G154, G3737, G215, G155, G133, G185, G162, G58, G163, G165, G60, G166, G1480, G147, G168, G44, G1, G56, G169, G171, G2211, G157, G172, G2208, G193, G197, G173, G86, G175, G89, G50, G189, G213, G176, G38, G178, G179, G74, G180, G181, G69, G182, G183, G177, G184, G103, G32, G187, G112, G191, G235, G190, G195, G70, G201;
    output G399, G370, G338, G321, G368, G362, G359, G471, G422, G344, G307, G304, G301, G273, G336, G333, G419, G327, G310, G276, G252, G295, G249, G416, G412, G382, G319, G379, G376, G365, G397, G353, G347, G394, G391, G388, G281, G330, G552, G316, G534, G554, G546, G530, G438, G270, G450, G432, G540, G418, G3, G448, G350, G484, G558, G482, G480, G404, G550, G494, G469, G524, G522, G298, G538, G442, G246, G258, G492, G548, G556, G440, G486, G544, G536, G313, G490, G542, G292, G414, G560, G528, G496, G532, G279, G526, G436, G488, G478, G324, G444, G402, G453, G278, G410, G2, G284, G408, G446, G373, G406, G264, G385, G286, G289, G356, G341;
    wire n316;
    wire n320;
    wire n323;
    wire n326;
    wire n330;
    wire n333;
    wire n336;
    wire n340;
    wire n344;
    wire n347;
    wire n350;
    wire n354;
    wire n357;
    wire n360;
    wire n364;
    wire n368;
    wire n371;
    wire n374;
    wire n378;
    wire n381;
    wire n384;
    wire n388;
    wire n392;
    wire n395;
    wire n398;
    wire n402;
    wire n405;
    wire n408;
    wire n412;
    wire n416;
    wire n419;
    wire n423;
    wire n426;
    wire n429;
    wire n433;
    wire n437;
    wire n441;
    wire n444;
    wire n448;
    wire n452;
    wire n455;
    wire n459;
    wire n463;
    wire n466;
    wire n470;
    wire n474;
    wire n477;
    wire n481;
    wire n485;
    wire n489;
    wire n493;
    wire n496;
    wire n499;
    wire n503;
    wire n507;
    wire n511;
    wire n514;
    wire n518;
    wire n521;
    wire n525;
    wire n529;
    wire n533;
    wire n537;
    wire n541;
    wire n545;
    wire n548;
    wire n552;
    wire n555;
    wire n558;
    wire n562;
    wire n565;
    wire n569;
    wire n573;
    wire n577;
    wire n580;
    wire n584;
    wire n588;
    wire n592;
    wire n595;
    wire n599;
    wire n603;
    wire n607;
    wire n611;
    wire n615;
    wire n618;
    wire n622;
    wire n625;
    wire n628;
    wire n632;
    wire n636;
    wire n639;
    wire n643;
    wire n647;
    wire n651;
    wire n654;
    wire n658;
    wire n662;
    wire n666;
    wire n670;
    wire n674;
    wire n678;
    wire n682;
    wire n686;
    wire n690;
    wire n694;
    wire n698;
    wire n701;
    wire n705;
    wire n709;
    wire n713;
    wire n717;
    wire n720;
    wire n724;
    wire n728;
    wire n732;
    wire n735;
    wire n739;
    wire n743;
    wire n747;
    wire n750;
    wire n754;
    wire n758;
    wire n762;
    wire n766;
    wire n770;
    wire n773;
    wire n777;
    wire n780;
    wire n784;
    wire n788;
    wire n792;
    wire n796;
    wire n800;
    wire n804;
    wire n808;
    wire n812;
    wire n815;
    wire n819;
    wire n823;
    wire n827;
    wire n831;
    wire n834;
    wire n838;
    wire n842;
    wire n846;
    wire n850;
    wire n854;
    wire n858;
    wire n862;
    wire n866;
    wire n870;
    wire n873;
    wire n877;
    wire n881;
    wire n885;
    wire n889;
    wire n892;
    wire n896;
    wire n900;
    wire n904;
    wire n908;
    wire n911;
    wire n915;
    wire n919;
    wire n923;
    wire n927;
    wire n931;
    wire n935;
    wire n938;
    wire n942;
    wire n945;
    wire n949;
    wire n953;
    wire n956;
    wire n960;
    wire n964;
    wire n968;
    wire n972;
    wire n975;
    wire n979;
    wire n983;
    wire n986;
    wire n990;
    wire n994;
    wire n998;
    wire n1002;
    wire n1005;
    wire n1009;
    wire n1013;
    wire n1017;
    wire n1021;
    wire n1024;
    wire n1028;
    wire n1031;
    wire n1034;
    wire n1038;
    wire n1042;
    wire n1046;
    wire n1050;
    wire n1053;
    wire n1057;
    wire n1061;
    wire n1065;
    wire n1069;
    wire n1072;
    wire n1075;
    wire n1079;
    wire n1083;
    wire n1087;
    wire n1091;
    wire n1094;
    wire n1098;
    wire n1101;
    wire n1104;
    wire n1108;
    wire n1112;
    wire n1116;
    wire n1120;
    wire n1123;
    wire n1127;
    wire n1130;
    wire n1133;
    wire n1137;
    wire n1141;
    wire n1145;
    wire n1149;
    wire n1152;
    wire n1156;
    wire n1159;
    wire n1162;
    wire n1166;
    wire n1170;
    wire n1174;
    wire n1178;
    wire n1181;
    wire n1185;
    wire n1188;
    wire n1191;
    wire n1195;
    wire n1199;
    wire n1203;
    wire n1207;
    wire n1210;
    wire n1214;
    wire n1217;
    wire n1220;
    wire n1224;
    wire n1228;
    wire n1232;
    wire n1236;
    wire n1240;
    wire n1244;
    wire n1248;
    wire n1252;
    wire n1256;
    wire n1260;
    wire n1264;
    wire n1268;
    wire n1272;
    wire n1276;
    wire n1280;
    wire n1284;
    wire n1288;
    wire n1292;
    wire n1296;
    wire n1300;
    wire n1304;
    wire n1307;
    wire n1311;
    wire n1315;
    wire n1319;
    wire n1323;
    wire n1326;
    wire n1330;
    wire n1333;
    wire n1336;
    wire n1340;
    wire n1344;
    wire n1348;
    wire n1352;
    wire n1355;
    wire n1359;
    wire n1363;
    wire n1367;
    wire n1371;
    wire n1374;
    wire n1378;
    wire n1382;
    wire n1386;
    wire n1390;
    wire n1394;
    wire n1398;
    wire n1401;
    wire n1404;
    wire n1408;
    wire n1412;
    wire n1415;
    wire n1419;
    wire n1423;
    wire n1427;
    wire n1431;
    wire n1434;
    wire n1438;
    wire n1442;
    wire n1446;
    wire n1449;
    wire n1452;
    wire n1455;
    wire n1459;
    wire n1463;
    wire n1467;
    wire n1471;
    wire n1474;
    wire n1478;
    wire n1482;
    wire n1486;
    wire n1490;
    wire n1493;
    wire n1497;
    wire n1501;
    wire n1505;
    wire n1509;
    wire n1512;
    wire n1516;
    wire n1519;
    wire n1523;
    wire n1527;
    wire n1531;
    wire n1535;
    wire n1539;
    wire n1543;
    wire n1547;
    wire n1551;
    wire n1554;
    wire n1558;
    wire n1561;
    wire n1564;
    wire n1568;
    wire n1571;
    wire n1575;
    wire n1579;
    wire n1583;
    wire n1586;
    wire n1590;
    wire n1594;
    wire n1598;
    wire n1602;
    wire n1605;
    wire n1609;
    wire n1613;
    wire n1617;
    wire n1621;
    wire n1625;
    wire n1629;
    wire n1633;
    wire n1637;
    wire n1641;
    wire n1645;
    wire n1649;
    wire n1653;
    wire n1657;
    wire n1661;
    wire n1665;
    wire n1669;
    wire n1673;
    wire n1677;
    wire n1681;
    wire n1685;
    wire n1689;
    wire n1693;
    wire n1697;
    wire n1701;
    wire n1705;
    wire n1708;
    wire n1711;
    wire n1715;
    wire n1719;
    wire n1723;
    wire n1727;
    wire n1730;
    wire n1734;
    wire n1738;
    wire n1741;
    wire n1745;
    wire n1749;
    wire n1753;
    wire n1757;
    wire n1761;
    wire n1765;
    wire n1769;
    wire n1773;
    wire n1777;
    wire n1781;
    wire n1785;
    wire n1789;
    wire n1793;
    wire n1797;
    wire n1800;
    wire n1804;
    wire n1808;
    wire n1812;
    wire n1820;
    wire n1824;
    wire n1828;
    wire n1832;
    wire n1836;
    wire n1840;
    wire n1844;
    wire n1848;
    wire n1852;
    wire n1856;
    wire n1860;
    wire n1864;
    wire n1868;
    wire n1872;
    wire n1876;
    wire n1880;
    wire n1884;
    wire n1888;
    wire n1892;
    wire n1896;
    wire n1900;
    wire n1904;
    wire n1907;
    wire n1911;
    wire n1915;
    wire n1919;
    wire n1923;
    wire n1927;
    wire n1931;
    wire n1935;
    wire n1939;
    wire n1943;
    wire n1947;
    wire n1951;
    wire n1955;
    wire n1959;
    wire n1963;
    wire n1967;
    wire n1971;
    wire n1975;
    wire n1979;
    wire n1983;
    wire n1987;
    wire n1991;
    wire n1995;
    wire n1999;
    wire n2003;
    wire n2007;
    wire n2011;
    wire n2015;
    wire n2019;
    wire n2023;
    wire n2027;
    wire n2030;
    wire n2034;
    wire n2038;
    wire n2042;
    wire n2046;
    wire n2050;
    wire n2054;
    wire n2058;
    wire n2061;
    wire n2065;
    wire n2069;
    wire n2073;
    wire n2077;
    wire n2081;
    wire n2085;
    wire n2089;
    wire n2093;
    wire n2097;
    wire n2101;
    wire n2105;
    wire n2109;
    wire n2112;
    wire n2115;
    wire n2119;
    wire n2123;
    wire n2127;
    wire n2131;
    wire n2135;
    wire n2138;
    wire n2142;
    wire n2146;
    wire n2150;
    wire n2154;
    wire n2158;
    wire n2162;
    wire n2166;
    wire n2170;
    wire n2174;
    wire n2178;
    wire n2182;
    wire n2186;
    wire n2190;
    wire n2193;
    wire n2197;
    wire n2201;
    wire n2205;
    wire n2209;
    wire n2213;
    wire n2217;
    wire n2221;
    wire n2225;
    wire n2229;
    wire n2233;
    wire n2237;
    wire n2241;
    wire n2245;
    wire n2249;
    wire n2253;
    wire n2257;
    wire n2261;
    wire n2265;
    wire n2269;
    wire n2273;
    wire n2277;
    wire n2281;
    wire n2285;
    wire n2289;
    wire n2293;
    wire n2297;
    wire n2301;
    wire n2305;
    wire n2309;
    wire n2313;
    wire n2317;
    wire n2321;
    wire n2325;
    wire n2329;
    wire n2333;
    wire n2337;
    wire n2341;
    wire n2345;
    wire n2349;
    wire n2353;
    wire n2357;
    wire n2361;
    wire n2365;
    wire n2369;
    wire n2373;
    wire n2377;
    wire n2381;
    wire n2384;
    wire n2388;
    wire n2392;
    wire n2396;
    wire n2400;
    wire n2404;
    wire n2408;
    wire n2412;
    wire n2415;
    wire n2419;
    wire n2423;
    wire n2427;
    wire n2431;
    wire n2435;
    wire n2439;
    wire n2443;
    wire n2447;
    wire n2451;
    wire n2455;
    wire n2459;
    wire n2463;
    wire n2467;
    wire n2471;
    wire n2475;
    wire n2479;
    wire n2483;
    wire n2487;
    wire n2491;
    wire n2495;
    wire n2499;
    wire n2503;
    wire n2507;
    wire n2511;
    wire n2515;
    wire n2519;
    wire n2523;
    wire n2527;
    wire n2531;
    wire n2535;
    wire n2539;
    wire n2543;
    wire n2547;
    wire n2551;
    wire n2555;
    wire n2559;
    wire n2563;
    wire n2567;
    wire n2571;
    wire n2575;
    wire n2579;
    wire n2583;
    wire n2587;
    wire n2591;
    wire n2595;
    wire n2599;
    wire n2603;
    wire n2607;
    wire n2611;
    wire n2615;
    wire n2619;
    wire n2623;
    wire n2627;
    wire n2631;
    wire n2635;
    wire n2639;
    wire n2643;
    wire n2647;
    wire n2651;
    wire n2654;
    wire n2658;
    wire n2662;
    wire n2666;
    wire n2670;
    wire n2674;
    wire n2678;
    wire n2682;
    wire n2686;
    wire n2690;
    wire n2694;
    wire n2698;
    wire n2702;
    wire n2706;
    wire n2710;
    wire n2714;
    wire n2718;
    wire n2722;
    wire n2726;
    wire n2730;
    wire n2734;
    wire n2738;
    wire n2742;
    wire n2746;
    wire n2750;
    wire n2754;
    wire n2758;
    wire n2762;
    wire n2766;
    wire n2770;
    wire n2774;
    wire n2778;
    wire n2782;
    wire n2786;
    wire n2790;
    wire n2794;
    wire n2798;
    wire n2802;
    wire n2806;
    wire n2810;
    wire n2813;
    wire n2817;
    wire n2821;
    wire n2825;
    wire n2829;
    wire n2833;
    wire n2837;
    wire n2840;
    wire n2844;
    wire n2848;
    wire n2852;
    wire n2856;
    wire n2860;
    wire n2864;
    wire n2868;
    wire n2872;
    wire n2876;
    wire n2880;
    wire n2884;
    wire n2888;
    wire n2892;
    wire n2895;
    wire n2899;
    wire n2903;
    wire n2907;
    wire n2910;
    wire n2914;
    wire n2918;
    wire n2922;
    wire n2925;
    wire n2929;
    wire n2933;
    wire n2937;
    wire n2941;
    wire n2945;
    wire n2949;
    wire n2952;
    wire n2956;
    wire n2960;
    wire n2964;
    wire n2968;
    wire n2971;
    wire n2975;
    wire n2979;
    wire n2983;
    wire n2987;
    wire n2991;
    wire n2995;
    wire n2999;
    wire n3003;
    wire n3007;
    wire n3011;
    wire n3015;
    wire n3019;
    wire n3023;
    wire n3027;
    wire n3031;
    wire n3034;
    wire n3037;
    wire n3041;
    wire n3045;
    wire n3049;
    wire n3053;
    wire n3057;
    wire n3061;
    wire n3065;
    wire n3069;
    wire n3073;
    wire n3077;
    wire n3081;
    wire n3085;
    wire n3089;
    wire n3093;
    wire n3097;
    wire n3101;
    wire n3105;
    wire n3109;
    wire n3113;
    wire n3117;
    wire n3121;
    wire n3125;
    wire n3129;
    wire n3133;
    wire n3137;
    wire n3141;
    wire n3145;
    wire n3149;
    wire n3153;
    wire n3157;
    wire n3161;
    wire n3165;
    wire n3169;
    wire n3173;
    wire n3176;
    wire n3179;
    wire n3182;
    wire n3186;
    wire n3190;
    wire n3194;
    wire n3198;
    wire n3202;
    wire n3206;
    wire n3210;
    wire n3213;
    wire n3217;
    wire n3221;
    wire n3225;
    wire n3229;
    wire n3233;
    wire n3237;
    wire n3241;
    wire n3245;
    wire n3249;
    wire n3253;
    wire n3257;
    wire n3261;
    wire n3265;
    wire n3269;
    wire n3272;
    wire n3275;
    wire n3278;
    wire n3282;
    wire n3286;
    wire n3290;
    wire n3294;
    wire n3298;
    wire n3301;
    wire n3305;
    wire n3309;
    wire n3313;
    wire n3317;
    wire n3321;
    wire n3325;
    wire n3329;
    wire n3333;
    wire n3337;
    wire n3341;
    wire n3344;
    wire n3347;
    wire n3350;
    wire n3354;
    wire n3358;
    wire n3362;
    wire n3366;
    wire n3370;
    wire n3373;
    wire n3377;
    wire n3380;
    wire n3384;
    wire n3388;
    wire n3391;
    wire n3395;
    wire n3399;
    wire n3403;
    wire n3407;
    wire n3410;
    wire n3414;
    wire n3418;
    wire n3421;
    wire n3425;
    wire n3428;
    wire n3432;
    wire n3436;
    wire n3440;
    wire n3444;
    wire n3448;
    wire n3452;
    wire n3456;
    wire n3460;
    wire n3464;
    wire n3468;
    wire n3472;
    wire n3476;
    wire n3480;
    wire n3484;
    wire n3488;
    wire n3492;
    wire n3496;
    wire n3500;
    wire n3504;
    wire n3508;
    wire n3512;
    wire n3516;
    wire n3520;
    wire n3524;
    wire n3528;
    wire n3531;
    wire n3535;
    wire n3538;
    wire n3542;
    wire n3546;
    wire n3550;
    wire n3553;
    wire n3557;
    wire n3561;
    wire n3565;
    wire n3569;
    wire n3573;
    wire n3577;
    wire n3581;
    wire n3585;
    wire n3589;
    wire n3593;
    wire n3597;
    wire n3601;
    wire n3605;
    wire n3609;
    wire n3613;
    wire n3617;
    wire n3621;
    wire n3625;
    wire n3628;
    wire n3632;
    wire n3635;
    wire n3639;
    wire n3643;
    wire n3647;
    wire n3651;
    wire n3655;
    wire n3659;
    wire n3663;
    wire n3667;
    wire n3671;
    wire n3675;
    wire n3679;
    wire n3683;
    wire n3687;
    wire n3691;
    wire n3694;
    wire n3698;
    wire n3702;
    wire n3706;
    wire n3710;
    wire n3714;
    wire n3718;
    wire n3722;
    wire n3726;
    wire n3729;
    wire n3733;
    wire n3737;
    wire n3741;
    wire n3745;
    wire n3749;
    wire n3753;
    wire n3757;
    wire n3761;
    wire n3765;
    wire n3768;
    wire n3772;
    wire n3776;
    wire n3780;
    wire n3784;
    wire n3788;
    wire n3792;
    wire n3796;
    wire n3800;
    wire n3804;
    wire n3807;
    wire n3811;
    wire n3815;
    wire n3819;
    wire n3823;
    wire n3827;
    wire n3831;
    wire n3834;
    wire n3838;
    wire n3842;
    wire n3846;
    wire n3850;
    wire n3854;
    wire n3858;
    wire n3862;
    wire n3866;
    wire n3869;
    wire n3873;
    wire n3877;
    wire n3881;
    wire n3885;
    wire n3889;
    wire n3893;
    wire n3897;
    wire n3901;
    wire n3905;
    wire n3909;
    wire n3913;
    wire n3917;
    wire n3921;
    wire n3925;
    wire n3929;
    wire n3933;
    wire n3937;
    wire n3941;
    wire n3945;
    wire n3949;
    wire n3953;
    wire n3956;
    wire n3960;
    wire n3964;
    wire n3968;
    wire n3972;
    wire n3976;
    wire n3980;
    wire n3984;
    wire n3987;
    wire n3991;
    wire n3994;
    wire n3998;
    wire n4002;
    wire n4005;
    wire n4009;
    wire n4012;
    wire n4016;
    wire n4020;
    wire n4024;
    wire n4028;
    wire n4032;
    wire n4035;
    wire n4039;
    wire n4043;
    wire n4047;
    wire n4051;
    wire n4055;
    wire n4058;
    wire n4062;
    wire n4065;
    wire n4069;
    wire n4073;
    wire n4076;
    wire n4080;
    wire n4083;
    wire n4087;
    wire n4091;
    wire n4095;
    wire n4099;
    wire n4103;
    wire n4107;
    wire n4111;
    wire n4114;
    wire n4117;
    wire n4120;
    wire n4123;
    wire n4126;
    wire n4129;
    wire n4132;
    wire n4136;
    wire n4140;
    wire n4144;
    wire n4148;
    wire n4152;
    wire n4156;
    wire n4160;
    wire n4164;
    wire n4168;
    wire n4172;
    wire n4176;
    wire n4179;
    wire n4182;
    wire n4185;
    wire n4188;
    wire n4191;
    wire n4194;
    wire n4197;
    wire n4200;
    wire n4204;
    wire n4208;
    wire n4212;
    wire n4216;
    wire n4220;
    wire n4224;
    wire n4228;
    wire n4232;
    wire n4236;
    wire n4239;
    wire n4243;
    wire n4246;
    wire n4250;
    wire n4254;
    wire n4258;
    wire n4262;
    wire n4266;
    wire n4269;
    wire n4273;
    wire n4277;
    wire n4280;
    wire n4284;
    wire n4288;
    wire n4292;
    wire n4296;
    wire n4300;
    wire n4304;
    wire n4308;
    wire n4312;
    wire n4316;
    wire n4320;
    wire n4324;
    wire n4328;
    wire n4332;
    wire n4336;
    wire n4340;
    wire n4344;
    wire n4347;
    wire n4350;
    wire n4353;
    wire n4357;
    wire n4361;
    wire n4365;
    wire n4369;
    wire n4377;
    wire n4381;
    wire n4385;
    wire n4389;
    wire n4393;
    wire n4397;
    wire n4401;
    wire n4405;
    wire n4409;
    wire n4413;
    wire n4417;
    wire n4421;
    wire n4424;
    wire n4428;
    wire n4432;
    wire n4436;
    wire n4440;
    wire n4444;
    wire n4448;
    wire n4452;
    wire n4456;
    wire n4464;
    wire n4468;
    wire n4472;
    wire n4476;
    wire n4479;
    wire n4482;
    wire n4485;
    wire n4488;
    wire n4492;
    wire n4496;
    wire n4500;
    wire n4503;
    wire n4507;
    wire n4511;
    wire n4515;
    wire n4519;
    wire n4523;
    wire n4527;
    wire n4531;
    wire n4535;
    wire n4539;
    wire n4543;
    wire n4547;
    wire n4551;
    wire n4555;
    wire n4559;
    wire n4563;
    wire n4567;
    wire n4571;
    wire n4575;
    wire n4579;
    wire n4583;
    wire n4586;
    wire n4590;
    wire n4594;
    wire n4598;
    wire n4602;
    wire n4606;
    wire n4610;
    wire n4614;
    wire n4617;
    wire n4621;
    wire n4625;
    wire n4629;
    wire n4633;
    wire n4637;
    wire n4641;
    wire n4645;
    wire n4649;
    wire n4653;
    wire n4657;
    wire n4661;
    wire n4665;
    wire n4668;
    wire n4672;
    wire n4676;
    wire n4679;
    wire n4683;
    wire n4686;
    wire n4690;
    wire n4694;
    wire n4698;
    wire n4702;
    wire n4706;
    wire n4710;
    wire n4714;
    wire n4718;
    wire n4722;
    wire n4726;
    wire n4730;
    wire n4734;
    wire n4738;
    wire n4742;
    wire n4746;
    wire n4750;
    wire n4754;
    wire n4758;
    wire n4762;
    wire n4766;
    wire n4770;
    wire n4774;
    wire n4778;
    wire n4782;
    wire n4786;
    wire n4789;
    wire n4793;
    wire n4797;
    wire n4801;
    wire n4805;
    wire n4809;
    wire n4813;
    wire n4817;
    wire n4821;
    wire n4825;
    wire n4828;
    wire n4832;
    wire n4836;
    wire n4840;
    wire n4844;
    wire n4848;
    wire n4852;
    wire n4856;
    wire n4860;
    wire n4864;
    wire n4868;
    wire n4872;
    wire n4875;
    wire n4879;
    wire n4882;
    wire n4886;
    wire n4890;
    wire n4894;
    wire n4897;
    wire n4901;
    wire n4905;
    wire n4909;
    wire n4913;
    wire n4917;
    wire n4921;
    wire n4925;
    wire n4928;
    wire n4932;
    wire n4936;
    wire n4940;
    wire n4944;
    wire n4948;
    wire n4952;
    wire n4956;
    wire n4960;
    wire n4964;
    wire n4968;
    wire n4972;
    wire n4976;
    wire n4980;
    wire n4984;
    wire n4988;
    wire n4991;
    wire n4995;
    wire n4999;
    wire n5003;
    wire n5007;
    wire n5011;
    wire n5015;
    wire n5019;
    wire n5023;
    wire n5027;
    wire n5031;
    wire n5035;
    wire n5039;
    wire n5043;
    wire n5047;
    wire n5051;
    wire n5054;
    wire n5058;
    wire n5061;
    wire n5065;
    wire n5069;
    wire n5073;
    wire n5077;
    wire n5081;
    wire n5084;
    wire n5088;
    wire n5091;
    wire n5095;
    wire n5099;
    wire n5103;
    wire n5107;
    wire n5111;
    wire n5115;
    wire n5119;
    wire n5122;
    wire n5126;
    wire n5130;
    wire n5134;
    wire n5138;
    wire n5142;
    wire n5146;
    wire n5150;
    wire n5154;
    wire n5158;
    wire n5162;
    wire n5166;
    wire n5170;
    wire n5174;
    wire n5178;
    wire n5182;
    wire n5186;
    wire n5190;
    wire n5193;
    wire n5197;
    wire n5201;
    wire n5205;
    wire n5209;
    wire n5213;
    wire n5217;
    wire n5221;
    wire n5225;
    wire n5229;
    wire n5233;
    wire n5237;
    wire n5241;
    wire n5245;
    wire n5249;
    wire n5253;
    wire n5257;
    wire n5261;
    wire n5265;
    wire n5268;
    wire n5272;
    wire n5276;
    wire n5280;
    wire n5283;
    wire n5287;
    wire n5291;
    wire n5295;
    wire n5299;
    wire n5303;
    wire n5307;
    wire n5311;
    wire n5315;
    wire n5318;
    wire n5321;
    wire n5325;
    wire n5329;
    wire n5332;
    wire n5336;
    wire n5340;
    wire n5344;
    wire n5348;
    wire n5352;
    wire n5356;
    wire n5360;
    wire n5364;
    wire n5367;
    wire n5370;
    wire n5373;
    wire n5376;
    wire n5379;
    wire n5382;
    wire n5385;
    wire n5388;
    wire n5391;
    wire n5394;
    wire n5397;
    wire n5400;
    wire n5403;
    wire n5406;
    wire n5409;
    wire n5412;
    wire n5415;
    wire n5418;
    wire n5421;
    wire n5424;
    wire n5427;
    wire n5430;
    wire n5433;
    wire n5436;
    wire n5439;
    wire n5442;
    wire n5445;
    wire n5448;
    wire n5451;
    wire n5454;
    wire n5457;
    wire n5460;
    wire n5463;
    wire n5466;
    wire n5469;
    wire n5472;
    wire n5475;
    wire n5478;
    wire n5481;
    wire n5484;
    wire n5487;
    wire n5490;
    wire n5494;
    wire n5497;
    wire n5501;
    wire n5504;
    wire n5508;
    wire n5516;
    wire n5532;
    wire n7855;
    wire n7858;
    wire n7861;
    wire n7865;
    wire n7868;
    wire n7871;
    wire n7874;
    wire n7877;
    wire n7880;
    wire n7883;
    wire n7886;
    wire n7889;
    wire n7892;
    wire n7895;
    wire n7898;
    wire n7901;
    wire n7904;
    wire n7907;
    wire n7910;
    wire n7913;
    wire n7916;
    wire n7919;
    wire n7922;
    wire n7925;
    wire n7928;
    wire n7931;
    wire n7934;
    wire n7937;
    wire n7940;
    wire n7943;
    wire n7946;
    wire n7949;
    wire n7952;
    wire n7955;
    wire n7958;
    wire n7961;
    wire n7964;
    wire n7967;
    wire n7970;
    wire n7973;
    wire n7976;
    wire n7979;
    wire n7982;
    wire n7985;
    wire n7988;
    wire n7991;
    wire n7994;
    wire n7997;
    wire n8000;
    wire n8003;
    wire n8006;
    wire n8009;
    wire n8012;
    wire n8015;
    wire n8018;
    wire n8021;
    wire n8024;
    wire n8027;
    wire n8030;
    wire n8033;
    wire n8036;
    wire n8039;
    wire n8042;
    wire n8045;
    wire n8048;
    wire n8051;
    wire n8054;
    wire n8056;
    wire n8060;
    wire n8063;
    wire n8066;
    wire n8069;
    wire n8072;
    wire n8075;
    wire n8078;
    wire n8081;
    wire n8084;
    wire n8087;
    wire n8090;
    wire n8093;
    wire n8096;
    wire n8099;
    wire n8102;
    wire n8105;
    wire n8108;
    wire n8111;
    wire n8114;
    wire n8117;
    wire n8120;
    wire n8123;
    wire n8126;
    wire n8129;
    wire n8132;
    wire n8135;
    wire n8138;
    wire n8141;
    wire n8144;
    wire n8147;
    wire n8150;
    wire n8153;
    wire n8156;
    wire n8159;
    wire n8162;
    wire n8165;
    wire n8168;
    wire n8171;
    wire n8174;
    wire n8177;
    wire n8180;
    wire n8183;
    wire n8186;
    wire n8189;
    wire n8192;
    wire n8195;
    wire n8198;
    wire n8201;
    wire n8204;
    wire n8207;
    wire n8210;
    wire n8213;
    wire n8216;
    wire n8219;
    wire n8222;
    wire n8225;
    wire n8228;
    wire n8231;
    wire n8234;
    wire n8237;
    wire n8240;
    wire n8243;
    wire n8246;
    wire n8249;
    wire n8252;
    wire n8255;
    wire n8258;
    wire n8261;
    wire n8264;
    wire n8267;
    wire n8270;
    wire n8273;
    wire n8276;
    wire n8279;
    wire n8282;
    wire n8285;
    wire n8288;
    wire n8291;
    wire n8294;
    wire n8297;
    wire n8300;
    wire n8303;
    wire n8306;
    wire n8309;
    wire n8312;
    wire n8315;
    wire n8318;
    wire n8321;
    wire n8324;
    wire n8326;
    wire n8329;
    wire n8333;
    wire n8336;
    wire n8338;
    wire n8342;
    wire n8345;
    wire n8348;
    wire n8351;
    wire n8354;
    wire n8357;
    wire n8360;
    wire n8362;
    wire n8365;
    wire n8368;
    wire n8371;
    wire n8375;
    wire n8378;
    wire n8381;
    wire n8384;
    wire n8387;
    wire n8390;
    wire n8393;
    wire n8396;
    wire n8399;
    wire n8402;
    wire n8405;
    wire n8408;
    wire n8411;
    wire n8414;
    wire n8417;
    wire n8420;
    wire n8423;
    wire n8426;
    wire n8429;
    wire n8432;
    wire n8435;
    wire n8438;
    wire n8441;
    wire n8444;
    wire n8447;
    wire n8450;
    wire n8453;
    wire n8456;
    wire n8459;
    wire n8462;
    wire n8465;
    wire n8468;
    wire n8471;
    wire n8474;
    wire n8477;
    wire n8480;
    wire n8483;
    wire n8486;
    wire n8489;
    wire n8492;
    wire n8495;
    wire n8498;
    wire n8501;
    wire n8504;
    wire n8507;
    wire n8510;
    wire n8513;
    wire n8516;
    wire n8519;
    wire n8522;
    wire n8525;
    wire n8528;
    wire n8531;
    wire n8534;
    wire n8537;
    wire n8540;
    wire n8543;
    wire n8546;
    wire n8549;
    wire n8552;
    wire n8555;
    wire n8558;
    wire n8561;
    wire n8564;
    wire n8567;
    wire n8570;
    wire n8573;
    wire n8576;
    wire n8579;
    wire n8582;
    wire n8585;
    wire n8588;
    wire n8591;
    wire n8594;
    wire n8597;
    wire n8600;
    wire n8603;
    wire n8606;
    wire n8609;
    wire n8612;
    wire n8615;
    wire n8618;
    wire n8621;
    wire n8624;
    wire n8627;
    wire n8630;
    wire n8633;
    wire n8636;
    wire n8639;
    wire n8642;
    wire n8645;
    wire n8648;
    wire n8651;
    wire n8654;
    wire n8657;
    wire n8660;
    wire n8662;
    wire n8665;
    wire n8668;
    wire n8671;
    wire n8675;
    wire n8677;
    wire n8680;
    wire n8683;
    wire n8687;
    wire n8690;
    wire n8693;
    wire n8696;
    wire n8699;
    wire n8702;
    wire n8705;
    wire n8708;
    wire n8711;
    wire n8714;
    wire n8717;
    wire n8720;
    wire n8723;
    wire n8726;
    wire n8729;
    wire n8732;
    wire n8735;
    wire n8738;
    wire n8741;
    wire n8744;
    wire n8747;
    wire n8750;
    wire n8753;
    wire n8756;
    wire n8759;
    wire n8762;
    wire n8765;
    wire n8768;
    wire n8771;
    wire n8774;
    wire n8777;
    wire n8780;
    wire n8783;
    wire n8785;
    wire n8788;
    wire n8792;
    wire n8795;
    wire n8797;
    wire n8800;
    wire n8804;
    wire n8807;
    wire n8810;
    wire n8813;
    wire n8816;
    wire n8819;
    wire n8822;
    wire n8825;
    wire n8828;
    wire n8831;
    wire n8834;
    wire n8837;
    wire n8840;
    wire n8843;
    wire n8846;
    wire n8849;
    wire n8852;
    wire n8855;
    wire n8858;
    wire n8861;
    wire n8864;
    wire n8867;
    wire n8870;
    wire n8873;
    wire n8876;
    wire n8879;
    wire n8882;
    wire n8885;
    wire n8888;
    wire n8891;
    wire n8894;
    wire n8897;
    wire n8900;
    wire n8903;
    wire n8906;
    wire n8909;
    wire n8912;
    wire n8915;
    wire n8918;
    wire n8921;
    wire n8924;
    wire n8927;
    wire n8930;
    wire n8933;
    wire n8936;
    wire n8939;
    wire n8942;
    wire n8945;
    wire n8948;
    wire n8951;
    wire n8954;
    wire n8957;
    wire n8960;
    wire n8963;
    wire n8966;
    wire n8969;
    wire n8972;
    wire n8975;
    wire n8978;
    wire n8981;
    wire n8984;
    wire n8987;
    wire n8990;
    wire n8993;
    wire n8996;
    wire n8999;
    wire n9002;
    wire n9005;
    wire n9008;
    wire n9011;
    wire n9014;
    wire n9017;
    wire n9020;
    wire n9023;
    wire n9026;
    wire n9029;
    wire n9032;
    wire n9035;
    wire n9038;
    wire n9041;
    wire n9044;
    wire n9047;
    wire n9050;
    wire n9053;
    wire n9056;
    wire n9059;
    wire n9062;
    wire n9065;
    wire n9068;
    wire n9071;
    wire n9074;
    wire n9077;
    wire n9080;
    wire n9083;
    wire n9086;
    wire n9089;
    wire n9092;
    wire n9095;
    wire n9098;
    wire n9101;
    wire n9104;
    wire n9107;
    wire n9110;
    wire n9113;
    wire n9116;
    wire n9119;
    wire n9122;
    wire n9125;
    wire n9128;
    wire n9131;
    wire n9134;
    wire n9137;
    wire n9140;
    wire n9143;
    wire n9146;
    wire n9149;
    wire n9152;
    wire n9155;
    wire n9158;
    wire n9161;
    wire n9164;
    wire n9167;
    wire n9170;
    wire n9173;
    wire n9176;
    wire n9179;
    wire n9182;
    wire n9185;
    wire n9188;
    wire n9191;
    wire n9194;
    wire n9197;
    wire n9200;
    wire n9203;
    wire n9206;
    wire n9209;
    wire n9212;
    wire n9215;
    wire n9218;
    wire n9221;
    wire n9224;
    wire n9227;
    wire n9230;
    wire n9233;
    wire n9236;
    wire n9239;
    wire n9242;
    wire n9245;
    wire n9248;
    wire n9251;
    wire n9254;
    wire n9257;
    wire n9260;
    wire n9263;
    wire n9266;
    wire n9269;
    wire n9272;
    wire n9275;
    wire n9278;
    wire n9281;
    wire n9284;
    wire n9287;
    wire n9290;
    wire n9293;
    wire n9296;
    wire n9299;
    wire n9302;
    wire n9305;
    wire n9307;
    wire n9311;
    wire n9314;
    wire n9317;
    wire n9320;
    wire n9323;
    wire n9326;
    wire n9328;
    wire n9331;
    wire n9335;
    wire n9337;
    wire n9340;
    wire n9344;
    wire n9347;
    wire n9349;
    wire n9353;
    wire n9356;
    wire n9359;
    wire n9362;
    wire n9364;
    wire n9368;
    wire n9371;
    wire n9374;
    wire n9377;
    wire n9380;
    wire n9383;
    wire n9386;
    wire n9389;
    wire n9392;
    wire n9395;
    wire n9398;
    wire n9401;
    wire n9404;
    wire n9407;
    wire n9410;
    wire n9413;
    wire n9416;
    wire n9419;
    wire n9422;
    wire n9425;
    wire n9428;
    wire n9431;
    wire n9433;
    wire n9437;
    wire n9439;
    wire n9443;
    wire n9446;
    wire n9449;
    wire n9452;
    wire n9455;
    wire n9458;
    wire n9461;
    wire n9464;
    wire n9467;
    wire n9469;
    wire n9472;
    wire n9475;
    wire n9479;
    wire n9482;
    wire n9485;
    wire n9487;
    wire n9491;
    wire n9494;
    wire n9496;
    wire n9500;
    wire n9503;
    wire n9506;
    wire n9509;
    wire n9512;
    wire n9515;
    wire n9518;
    wire n9521;
    wire n9523;
    wire n9527;
    wire n9530;
    wire n9532;
    wire n9536;
    wire n9539;
    wire n9542;
    wire n9545;
    wire n9548;
    wire n9551;
    wire n9554;
    wire n9557;
    wire n9560;
    wire n9563;
    wire n9566;
    wire n9569;
    wire n9572;
    wire n9575;
    wire n9578;
    wire n9581;
    wire n9584;
    wire n9586;
    wire n9590;
    wire n9593;
    wire n9596;
    wire n9599;
    wire n9602;
    wire n9605;
    wire n9608;
    wire n9611;
    wire n9614;
    wire n9617;
    wire n9620;
    wire n9623;
    wire n9626;
    wire n9629;
    wire n9632;
    wire n9635;
    wire n9638;
    wire n9641;
    wire n9644;
    wire n9647;
    wire n9650;
    wire n9653;
    wire n9656;
    wire n9659;
    wire n9662;
    wire n9665;
    wire n9668;
    wire n9671;
    wire n9674;
    wire n9677;
    wire n9680;
    wire n9683;
    wire n9686;
    wire n9689;
    wire n9692;
    wire n9695;
    wire n9698;
    wire n9701;
    wire n9704;
    wire n9707;
    wire n9710;
    wire n9713;
    wire n9716;
    wire n9719;
    wire n9722;
    wire n9725;
    wire n9728;
    wire n9731;
    wire n9734;
    wire n9737;
    wire n9740;
    wire n9743;
    wire n9746;
    wire n9749;
    wire n9752;
    wire n9755;
    wire n9758;
    wire n9761;
    wire n9764;
    wire n9767;
    wire n9770;
    wire n9773;
    wire n9776;
    wire n9779;
    wire n9782;
    wire n9785;
    wire n9788;
    wire n9791;
    wire n9794;
    wire n9797;
    wire n9800;
    wire n9802;
    wire n9805;
    wire n9808;
    wire n9811;
    wire n9814;
    wire n9817;
    wire n9820;
    wire n9823;
    wire n9826;
    wire n9829;
    wire n9832;
    wire n9835;
    wire n9838;
    wire n9841;
    wire n9844;
    wire n9847;
    wire n9850;
    wire n9853;
    wire n9856;
    wire n9859;
    wire n9862;
    wire n9865;
    wire n9868;
    wire n9871;
    wire n9874;
    wire n9877;
    wire n9880;
    wire n9883;
    wire n9886;
    wire n9889;
    wire n9892;
    wire n9895;
    wire n9898;
    wire n9901;
    wire n9904;
    wire n9907;
    wire n9910;
    wire n9913;
    wire n9916;
    wire n9920;
    wire n9923;
    wire n9926;
    wire n9929;
    wire n9932;
    wire n9935;
    wire n9938;
    wire n9941;
    wire n9944;
    wire n9947;
    wire n9950;
    wire n9953;
    wire n9956;
    wire n9959;
    wire n9962;
    wire n9965;
    wire n9968;
    wire n9971;
    wire n9974;
    wire n9977;
    wire n9980;
    wire n9983;
    wire n9986;
    wire n9989;
    wire n9992;
    wire n9995;
    wire n9998;
    wire n10001;
    wire n10004;
    wire n10007;
    wire n10010;
    wire n10013;
    wire n10016;
    wire n10018;
    wire n10022;
    wire n10025;
    wire n10028;
    wire n10031;
    wire n10034;
    wire n10037;
    wire n10040;
    wire n10043;
    wire n10046;
    wire n10049;
    wire n10052;
    wire n10055;
    wire n10058;
    wire n10061;
    wire n10064;
    wire n10067;
    wire n10070;
    wire n10073;
    wire n10076;
    wire n10079;
    wire n10082;
    wire n10085;
    wire n10088;
    wire n10091;
    wire n10094;
    wire n10097;
    wire n10100;
    wire n10103;
    wire n10106;
    wire n10109;
    wire n10112;
    wire n10115;
    wire n10118;
    wire n10121;
    wire n10124;
    wire n10127;
    wire n10130;
    wire n10133;
    wire n10136;
    wire n10139;
    wire n10142;
    wire n10145;
    wire n10148;
    wire n10151;
    wire n10154;
    wire n10157;
    wire n10160;
    wire n10163;
    wire n10166;
    wire n10169;
    wire n10172;
    wire n10175;
    wire n10178;
    wire n10181;
    wire n10184;
    wire n10187;
    wire n10190;
    wire n10193;
    wire n10196;
    wire n10199;
    wire n10202;
    wire n10205;
    wire n10208;
    wire n10211;
    wire n10214;
    wire n10217;
    wire n10220;
    wire n10223;
    wire n10226;
    wire n10229;
    wire n10232;
    wire n10235;
    wire n10238;
    wire n10241;
    wire n10244;
    wire n10247;
    wire n10250;
    wire n10253;
    wire n10256;
    wire n10259;
    wire n10262;
    wire n10265;
    wire n10268;
    wire n10271;
    wire n10274;
    wire n10277;
    wire n10280;
    wire n10283;
    wire n10286;
    wire n10289;
    wire n10292;
    wire n10295;
    wire n10298;
    wire n10301;
    wire n10304;
    wire n10307;
    wire n10310;
    wire n10313;
    wire n10316;
    wire n10319;
    wire n10322;
    wire n10325;
    wire n10328;
    wire n10331;
    wire n10334;
    wire n10337;
    wire n10340;
    wire n10343;
    wire n10346;
    wire n10349;
    wire n10352;
    wire n10355;
    wire n10358;
    wire n10361;
    wire n10364;
    wire n10367;
    wire n10370;
    wire n10373;
    wire n10376;
    wire n10379;
    wire n10382;
    wire n10385;
    wire n10388;
    wire n10391;
    wire n10393;
    wire n10396;
    wire n10399;
    wire n10402;
    wire n10405;
    wire n10408;
    wire n10411;
    wire n10414;
    wire n10417;
    wire n10420;
    wire n10423;
    wire n10426;
    wire n10429;
    wire n10432;
    wire n10435;
    wire n10438;
    wire n10441;
    wire n10444;
    wire n10447;
    wire n10450;
    wire n10453;
    wire n10456;
    wire n10459;
    wire n10462;
    wire n10465;
    wire n10468;
    wire n10471;
    wire n10474;
    wire n10477;
    wire n10481;
    wire n10484;
    wire n10487;
    wire n10490;
    wire n10493;
    wire n10496;
    wire n10499;
    wire n10502;
    wire n10505;
    wire n10508;
    wire n10511;
    wire n10514;
    wire n10517;
    wire n10520;
    wire n10523;
    wire n10526;
    wire n10529;
    wire n10532;
    wire n10535;
    wire n10538;
    wire n10541;
    wire n10544;
    wire n10547;
    wire n10550;
    wire n10553;
    wire n10556;
    wire n10559;
    wire n10562;
    wire n10565;
    wire n10568;
    wire n10571;
    wire n10574;
    wire n10577;
    wire n10580;
    wire n10583;
    wire n10586;
    wire n10589;
    wire n10592;
    wire n10595;
    wire n10598;
    wire n10601;
    wire n10604;
    wire n10607;
    wire n10610;
    wire n10613;
    wire n10616;
    wire n10619;
    wire n10621;
    wire n10624;
    wire n10627;
    wire n10630;
    wire n10633;
    wire n10636;
    wire n10639;
    wire n10642;
    wire n10645;
    wire n10648;
    wire n10651;
    wire n10654;
    wire n10657;
    wire n10660;
    wire n10663;
    wire n10666;
    wire n10669;
    wire n10672;
    wire n10675;
    wire n10678;
    wire n10681;
    wire n10684;
    wire n10687;
    wire n10690;
    wire n10693;
    wire n10696;
    wire n10699;
    wire n10703;
    wire n10706;
    wire n10709;
    wire n10712;
    wire n10715;
    wire n10718;
    wire n10721;
    wire n10724;
    wire n10727;
    wire n10730;
    wire n10733;
    wire n10736;
    wire n10739;
    wire n10742;
    wire n10745;
    wire n10748;
    wire n10751;
    wire n10754;
    wire n10757;
    wire n10760;
    wire n10763;
    wire n10766;
    wire n10769;
    wire n10771;
    wire n10774;
    wire n10777;
    wire n10780;
    wire n10783;
    wire n10786;
    wire n10789;
    wire n10792;
    wire n10795;
    wire n10798;
    wire n10801;
    wire n10804;
    wire n10807;
    wire n10810;
    wire n10813;
    wire n10816;
    wire n10819;
    wire n10822;
    wire n10825;
    wire n10828;
    wire n10831;
    wire n10834;
    wire n10837;
    wire n10840;
    wire n10843;
    wire n10846;
    wire n10849;
    wire n10852;
    wire n10855;
    wire n10858;
    wire n10861;
    wire n10864;
    wire n10867;
    wire n10870;
    wire n10873;
    wire n10876;
    wire n10879;
    wire n10882;
    wire n10885;
    wire n10888;
    wire n10891;
    wire n10894;
    wire n10898;
    wire n10901;
    wire n10904;
    wire n10907;
    wire n10910;
    wire n10913;
    wire n10916;
    wire n10918;
    wire n10921;
    wire n10924;
    wire n10927;
    wire n10930;
    wire n10933;
    wire n10937;
    wire n10940;
    wire n10943;
    wire n10946;
    wire n10949;
    wire n10952;
    wire n10955;
    wire n10958;
    wire n10961;
    wire n10964;
    wire n10967;
    wire n10970;
    wire n10973;
    wire n10976;
    wire n10979;
    wire n10982;
    wire n10985;
    wire n10988;
    wire n10991;
    wire n10994;
    wire n10997;
    wire n11000;
    wire n11003;
    wire n11006;
    wire n11009;
    wire n11012;
    wire n11015;
    wire n11018;
    wire n11020;
    wire n11023;
    wire n11026;
    wire n11029;
    wire n11032;
    wire n11035;
    wire n11039;
    wire n11042;
    wire n11045;
    wire n11048;
    wire n11051;
    wire n11054;
    wire n11057;
    wire n11060;
    wire n11063;
    wire n11065;
    wire n11068;
    wire n11071;
    wire n11074;
    wire n11077;
    wire n11080;
    wire n11083;
    wire n11086;
    wire n11089;
    wire n11092;
    wire n11095;
    wire n11099;
    wire n11102;
    wire n11105;
    wire n11108;
    wire n11111;
    wire n11114;
    wire n11117;
    wire n11120;
    wire n11122;
    wire n11125;
    wire n11128;
    wire n11131;
    wire n11134;
    wire n11137;
    wire n11140;
    wire n11143;
    wire n11146;
    wire n11149;
    wire n11152;
    wire n11155;
    wire n11158;
    wire n11161;
    wire n11164;
    wire n11167;
    wire n11170;
    wire n11173;
    wire n11176;
    wire n11179;
    wire n11182;
    wire n11185;
    wire n11188;
    wire n11191;
    wire n11194;
    wire n11197;
    wire n11200;
    wire n11203;
    wire n11206;
    wire n11209;
    wire n11212;
    wire n11215;
    wire n11218;
    wire n11221;
    wire n11224;
    wire n11228;
    wire n11231;
    wire n11234;
    wire n11237;
    wire n11240;
    wire n11243;
    wire n11246;
    wire n11249;
    wire n11252;
    wire n11255;
    wire n11258;
    wire n11261;
    wire n11264;
    wire n11267;
    wire n11270;
    wire n11273;
    wire n11276;
    wire n11279;
    wire n11282;
    wire n11285;
    wire n11288;
    wire n11291;
    wire n11294;
    wire n11297;
    wire n11300;
    wire n11303;
    wire n11306;
    wire n11309;
    wire n11312;
    wire n11315;
    wire n11318;
    wire n11321;
    wire n11324;
    wire n11327;
    wire n11330;
    wire n11333;
    wire n11336;
    wire n11339;
    wire n11342;
    wire n11345;
    wire n11348;
    wire n11351;
    wire n11354;
    wire n11357;
    wire n11360;
    wire n11363;
    wire n11366;
    wire n11369;
    wire n11372;
    wire n11375;
    wire n11378;
    wire n11381;
    wire n11384;
    wire n11387;
    wire n11390;
    wire n11393;
    wire n11396;
    wire n11399;
    wire n11401;
    wire n11404;
    wire n11407;
    wire n11410;
    wire n11413;
    wire n11416;
    wire n11419;
    wire n11422;
    wire n11425;
    wire n11428;
    wire n11431;
    wire n11434;
    wire n11437;
    wire n11440;
    wire n11443;
    wire n11446;
    wire n11449;
    wire n11452;
    wire n11455;
    wire n11458;
    wire n11461;
    wire n11464;
    wire n11467;
    wire n11470;
    wire n11473;
    wire n11477;
    wire n11480;
    wire n11483;
    wire n11486;
    wire n11489;
    wire n11492;
    wire n11495;
    wire n11498;
    wire n11500;
    wire n11503;
    wire n11506;
    wire n11509;
    wire n11512;
    wire n11515;
    wire n11518;
    wire n11521;
    wire n11524;
    wire n11527;
    wire n11530;
    wire n11533;
    wire n11536;
    wire n11539;
    wire n11542;
    wire n11545;
    wire n11548;
    wire n11551;
    wire n11554;
    wire n11557;
    wire n11560;
    wire n11563;
    wire n11567;
    wire n11569;
    wire n11572;
    wire n11575;
    wire n11578;
    wire n11581;
    wire n11585;
    wire n11588;
    wire n11591;
    wire n11594;
    wire n11597;
    wire n11600;
    wire n11603;
    wire n11606;
    wire n11609;
    wire n11612;
    wire n11615;
    wire n11618;
    wire n11621;
    wire n11624;
    wire n11627;
    wire n11630;
    wire n11633;
    wire n11636;
    wire n11639;
    wire n11642;
    wire n11645;
    wire n11648;
    wire n11651;
    wire n11654;
    wire n11657;
    wire n11660;
    wire n11663;
    wire n11666;
    wire n11669;
    wire n11672;
    wire n11675;
    wire n11678;
    wire n11681;
    wire n11684;
    wire n11687;
    wire n11690;
    wire n11693;
    wire n11696;
    wire n11699;
    wire n11702;
    wire n11705;
    wire n11708;
    wire n11711;
    wire n11714;
    wire n11717;
    wire n11720;
    wire n11723;
    wire n11726;
    wire n11729;
    wire n11732;
    wire n11735;
    wire n11738;
    wire n11741;
    wire n11744;
    wire n11747;
    wire n11750;
    wire n11753;
    wire n11756;
    wire n11759;
    wire n11762;
    wire n11765;
    wire n11768;
    wire n11771;
    wire n11774;
    wire n11777;
    wire n11780;
    wire n11783;
    wire n11786;
    wire n11789;
    wire n11792;
    wire n11795;
    wire n11798;
    wire n11801;
    wire n11804;
    wire n11807;
    wire n11810;
    wire n11813;
    wire n11816;
    wire n11819;
    wire n11822;
    wire n11825;
    wire n11828;
    wire n11831;
    wire n11834;
    wire n11837;
    wire n11840;
    wire n11843;
    wire n11846;
    wire n11849;
    wire n11852;
    wire n11855;
    wire n11858;
    wire n11861;
    wire n11864;
    wire n11867;
    wire n11870;
    wire n11873;
    wire n11876;
    wire n11879;
    wire n11882;
    wire n11885;
    wire n11888;
    wire n11891;
    wire n11894;
    wire n11897;
    wire n11900;
    wire n11903;
    wire n11906;
    wire n11909;
    wire n11912;
    wire n11915;
    wire n11918;
    wire n11921;
    wire n11924;
    wire n11927;
    wire n11930;
    wire n11933;
    wire n11936;
    wire n11939;
    wire n11942;
    wire n11945;
    wire n11948;
    wire n11951;
    wire n11954;
    wire n11957;
    wire n11960;
    wire n11963;
    wire n11966;
    wire n11969;
    wire n11972;
    wire n11975;
    wire n11978;
    wire n11981;
    wire n11984;
    wire n11987;
    wire n11990;
    wire n11993;
    wire n11996;
    wire n11999;
    wire n12002;
    wire n12005;
    wire n12008;
    wire n12011;
    wire n12014;
    wire n12017;
    wire n12020;
    wire n12023;
    wire n12026;
    wire n12029;
    wire n12032;
    wire n12035;
    wire n12038;
    wire n12041;
    wire n12044;
    wire n12047;
    wire n12050;
    wire n12053;
    wire n12056;
    wire n12059;
    wire n12062;
    wire n12065;
    wire n12068;
    wire n12071;
    wire n12074;
    wire n12077;
    wire n12080;
    wire n12083;
    wire n12086;
    wire n12089;
    wire n12092;
    wire n12095;
    wire n12097;
    wire n12101;
    wire n12104;
    wire n12107;
    wire n12110;
    wire n12113;
    wire n12116;
    wire n12119;
    wire n12122;
    wire n12125;
    wire n12128;
    wire n12131;
    wire n12134;
    wire n12137;
    wire n12140;
    wire n12143;
    wire n12146;
    wire n12149;
    wire n12152;
    wire n12155;
    wire n12158;
    wire n12161;
    wire n12164;
    wire n12167;
    wire n12170;
    wire n12173;
    wire n12176;
    wire n12179;
    wire n12182;
    wire n12185;
    wire n12188;
    wire n12191;
    wire n12194;
    wire n12197;
    wire n12200;
    wire n12203;
    wire n12206;
    wire n12209;
    wire n12212;
    wire n12215;
    wire n12218;
    wire n12221;
    wire n12224;
    wire n12227;
    wire n12230;
    wire n12232;
    wire n12235;
    wire n12238;
    wire n12241;
    wire n12244;
    wire n12247;
    wire n12250;
    wire n12253;
    wire n12257;
    wire n12260;
    wire n12262;
    wire n12265;
    wire n12268;
    wire n12271;
    wire n12274;
    wire n12277;
    wire n12280;
    wire n12283;
    wire n12286;
    wire n12289;
    wire n12292;
    wire n12295;
    wire n12298;
    wire n12301;
    wire n12304;
    wire n12307;
    wire n12310;
    wire n12313;
    wire n12316;
    wire n12319;
    wire n12322;
    wire n12325;
    wire n12328;
    wire n12331;
    wire n12334;
    wire n12337;
    wire n12340;
    wire n12343;
    wire n12347;
    wire n12350;
    wire n12352;
    wire n12355;
    wire n12358;
    wire n12361;
    wire n12364;
    wire n12367;
    wire n12370;
    wire n12373;
    wire n12376;
    wire n12379;
    wire n12382;
    wire n12385;
    wire n12388;
    wire n12391;
    wire n12394;
    wire n12397;
    wire n12400;
    wire n12403;
    wire n12406;
    wire n12409;
    wire n12412;
    wire n12415;
    wire n12418;
    wire n12422;
    wire n12425;
    wire n12428;
    wire n12431;
    wire n12434;
    wire n12437;
    wire n12440;
    wire n12443;
    wire n12446;
    wire n12448;
    wire n12451;
    wire n12454;
    wire n12457;
    wire n12460;
    wire n12463;
    wire n12466;
    wire n12469;
    wire n12472;
    wire n12475;
    wire n12478;
    wire n12481;
    wire n12484;
    wire n12487;
    wire n12490;
    wire n12493;
    wire n12496;
    wire n12499;
    wire n12502;
    wire n12505;
    wire n12508;
    wire n12511;
    wire n12514;
    wire n12517;
    wire n12520;
    wire n12524;
    wire n12526;
    wire n12529;
    wire n12532;
    wire n12535;
    wire n12538;
    wire n12541;
    wire n12544;
    wire n12547;
    wire n12550;
    wire n12553;
    wire n12556;
    wire n12559;
    wire n12562;
    wire n12565;
    wire n12568;
    wire n12571;
    wire n12574;
    wire n12577;
    wire n12580;
    wire n12583;
    wire n12586;
    wire n12589;
    wire n12592;
    wire n12595;
    wire n12598;
    wire n12601;
    wire n12604;
    wire n12607;
    wire n12610;
    wire n12613;
    wire n12616;
    wire n12619;
    wire n12622;
    wire n12626;
    wire n12628;
    wire n12631;
    wire n12634;
    wire n12637;
    wire n12640;
    wire n12643;
    wire n12646;
    wire n12649;
    wire n12652;
    wire n12656;
    wire n12658;
    wire n12661;
    wire n12664;
    wire n12667;
    wire n12670;
    wire n12673;
    wire n12676;
    wire n12679;
    wire n12682;
    wire n12685;
    wire n12688;
    wire n12691;
    wire n12694;
    wire n12697;
    wire n12700;
    wire n12703;
    wire n12706;
    wire n12710;
    wire n12712;
    wire n12715;
    wire n12718;
    wire n12721;
    wire n12725;
    wire n12728;
    wire n12731;
    wire n12734;
    wire n12737;
    wire n12740;
    wire n12743;
    wire n12746;
    wire n12749;
    wire n12752;
    wire n12755;
    wire n12758;
    wire n12761;
    wire n12764;
    wire n12767;
    wire n12770;
    wire n12773;
    wire n12776;
    wire n12779;
    wire n12782;
    wire n12785;
    wire n12788;
    wire n12791;
    wire n12794;
    wire n12797;
    wire n12800;
    wire n12803;
    wire n12806;
    wire n12809;
    wire n12812;
    wire n12815;
    wire n12818;
    wire n12821;
    wire n12823;
    wire n12826;
    wire n12829;
    wire n12832;
    wire n12835;
    wire n12838;
    wire n12841;
    wire n12844;
    wire n12847;
    wire n12850;
    wire n12853;
    wire n12856;
    wire n12859;
    wire n12862;
    wire n12865;
    wire n12869;
    wire n12872;
    wire n12875;
    wire n12878;
    wire n12881;
    wire n12884;
    wire n12887;
    wire n12890;
    wire n12893;
    wire n12896;
    wire n12899;
    wire n12902;
    wire n12905;
    wire n12908;
    wire n12911;
    wire n12914;
    wire n12917;
    wire n12920;
    wire n12923;
    wire n12926;
    wire n12929;
    wire n12932;
    wire n12935;
    wire n12938;
    wire n12941;
    wire n12944;
    wire n12947;
    wire n12950;
    wire n12953;
    wire n12956;
    wire n12959;
    wire n12962;
    wire n12965;
    wire n12968;
    wire n12970;
    wire n12973;
    wire n12976;
    wire n12979;
    wire n12982;
    wire n12985;
    wire n12988;
    wire n12991;
    wire n12994;
    wire n12997;
    wire n13000;
    wire n13003;
    wire n13006;
    wire n13009;
    wire n13012;
    wire n13015;
    wire n13018;
    wire n13021;
    wire n13024;
    wire n13027;
    wire n13030;
    wire n13033;
    wire n13036;
    wire n13039;
    wire n13042;
    wire n13045;
    wire n13048;
    wire n13051;
    wire n13054;
    wire n13057;
    wire n13060;
    wire n13063;
    wire n13066;
    wire n13069;
    wire n13072;
    wire n13075;
    wire n13078;
    wire n13081;
    wire n13084;
    wire n13087;
    wire n13090;
    wire n13093;
    wire n13096;
    wire n13099;
    wire n13102;
    wire n13105;
    wire n13108;
    wire n13111;
    wire n13114;
    wire n13117;
    wire n13120;
    wire n13123;
    wire n13126;
    wire n13129;
    wire n13132;
    wire n13135;
    wire n13138;
    wire n13141;
    wire n13144;
    wire n13147;
    wire n13150;
    wire n13153;
    wire n13156;
    wire n13159;
    wire n13162;
    wire n13165;
    wire n13168;
    wire n13171;
    wire n13174;
    wire n13177;
    wire n13180;
    wire n13183;
    wire n13186;
    wire n13189;
    wire n13192;
    wire n13195;
    wire n13198;
    wire n13201;
    wire n13204;
    wire n13207;
    wire n13210;
    wire n13213;
    wire n13216;
    wire n13219;
    wire n13222;
    wire n13225;
    wire n13228;
    wire n13231;
    wire n13234;
    wire n13237;
    wire n13240;
    wire n13243;
    wire n13246;
    wire n13249;
    wire n13252;
    wire n13255;
    wire n13258;
    wire n13261;
    wire n13264;
    wire n13267;
    wire n13270;
    wire n13273;
    wire n13276;
    wire n13279;
    wire n13282;
    wire n13285;
    wire n13288;
    wire n13291;
    wire n13294;
    wire n13297;
    wire n13300;
    wire n13303;
    wire n13306;
    wire n13309;
    wire n13312;
    wire n13316;
    wire n13319;
    wire n13322;
    wire n13324;
    wire n13327;
    wire n13330;
    wire n13333;
    wire n13336;
    wire n13339;
    wire n13342;
    wire n13345;
    wire n13348;
    wire n13351;
    wire n13354;
    wire n13357;
    wire n13360;
    wire n13363;
    wire n13366;
    wire n13369;
    wire n13372;
    wire n13375;
    wire n13378;
    wire n13382;
    wire n13385;
    wire n13387;
    wire n13390;
    wire n13393;
    wire n13396;
    wire n13399;
    wire n13402;
    wire n13405;
    wire n13408;
    wire n13411;
    wire n13414;
    wire n13417;
    wire n13420;
    wire n13423;
    wire n13426;
    wire n13429;
    wire n13432;
    wire n13435;
    wire n13438;
    wire n13441;
    wire n13444;
    wire n13447;
    wire n13450;
    wire n13453;
    wire n13456;
    wire n13459;
    wire n13462;
    wire n13465;
    wire n13468;
    wire n13471;
    wire n13474;
    wire n13477;
    wire n13480;
    wire n13483;
    wire n13486;
    wire n13489;
    wire n13492;
    wire n13495;
    wire n13498;
    wire n13501;
    wire n13504;
    wire n13507;
    wire n13510;
    wire n13513;
    wire n13516;
    wire n13519;
    wire n13522;
    wire n13525;
    wire n13528;
    wire n13531;
    wire n13534;
    wire n13537;
    wire n13540;
    wire n13543;
    wire n13546;
    wire n13549;
    wire n13552;
    wire n13555;
    wire n13558;
    wire n13561;
    wire n13564;
    wire n13567;
    wire n13570;
    wire n13573;
    wire n13576;
    wire n13579;
    wire n13582;
    wire n13585;
    wire n13588;
    wire n13591;
    wire n13594;
    wire n13597;
    wire n13600;
    wire n13603;
    wire n13606;
    wire n13610;
    wire n13613;
    wire n13615;
    wire n13618;
    wire n13621;
    wire n13624;
    wire n13627;
    wire n13630;
    wire n13633;
    wire n13636;
    wire n13639;
    wire n13642;
    wire n13645;
    wire n13648;
    wire n13651;
    wire n13654;
    wire n13657;
    wire n13660;
    wire n13663;
    wire n13666;
    wire n13669;
    wire n13672;
    wire n13675;
    wire n13678;
    wire n13681;
    wire n13684;
    wire n13687;
    wire n13690;
    wire n13693;
    wire n13696;
    wire n13699;
    wire n13702;
    wire n13705;
    wire n13708;
    wire n13711;
    wire n13715;
    wire n13718;
    wire n13720;
    wire n13723;
    wire n13726;
    wire n13729;
    wire n13732;
    wire n13735;
    wire n13738;
    wire n13741;
    wire n13744;
    wire n13747;
    wire n13750;
    wire n13753;
    wire n13756;
    wire n13759;
    wire n13762;
    wire n13765;
    wire n13768;
    wire n13771;
    wire n13774;
    wire n13777;
    wire n13780;
    wire n13783;
    wire n13786;
    wire n13789;
    wire n13792;
    wire n13795;
    wire n13798;
    wire n13801;
    wire n13804;
    wire n13807;
    wire n13810;
    wire n13813;
    wire n13816;
    wire n13819;
    wire n13822;
    wire n13826;
    wire n13829;
    wire n13832;
    wire n13835;
    wire n13837;
    wire n13840;
    wire n13843;
    wire n13846;
    wire n13849;
    wire n13853;
    wire n13856;
    wire n13859;
    wire n13862;
    wire n13864;
    wire n13867;
    wire n13870;
    wire n13873;
    wire n13876;
    wire n13879;
    wire n13882;
    wire n13885;
    wire n13888;
    wire n13891;
    wire n13894;
    wire n13897;
    wire n13900;
    wire n13903;
    wire n13906;
    wire n13909;
    wire n13912;
    wire n13915;
    wire n13918;
    wire n13921;
    wire n13924;
    wire n13927;
    wire n13930;
    wire n13933;
    wire n13936;
    wire n13939;
    wire n13942;
    wire n13945;
    wire n13948;
    wire n13951;
    wire n13954;
    wire n13957;
    wire n13960;
    wire n13963;
    wire n13966;
    wire n13969;
    wire n13972;
    wire n13975;
    wire n13978;
    wire n13981;
    wire n13984;
    wire n13987;
    wire n13990;
    wire n13993;
    wire n13996;
    wire n13999;
    wire n14002;
    wire n14005;
    wire n14008;
    wire n14011;
    wire n14014;
    wire n14017;
    wire n14020;
    wire n14023;
    wire n14026;
    wire n14029;
    wire n14032;
    wire n14035;
    wire n14038;
    wire n14041;
    wire n14044;
    wire n14047;
    wire n14050;
    wire n14053;
    wire n14056;
    wire n14059;
    wire n14062;
    wire n14065;
    wire n14068;
    wire n14071;
    wire n14074;
    wire n14077;
    wire n14080;
    wire n14083;
    wire n14086;
    wire n14089;
    wire n14092;
    wire n14095;
    wire n14098;
    wire n14101;
    wire n14104;
    wire n14107;
    wire n14110;
    wire n14113;
    wire n14116;
    wire n14119;
    wire n14122;
    wire n14126;
    wire n14128;
    wire n14131;
    wire n14134;
    wire n14137;
    wire n14140;
    wire n14143;
    wire n14146;
    wire n14149;
    wire n14152;
    wire n14155;
    wire n14158;
    wire n14161;
    wire n14164;
    wire n14167;
    wire n14170;
    wire n14173;
    wire n14176;
    wire n14179;
    wire n14182;
    wire n14185;
    wire n14188;
    wire n14191;
    wire n14194;
    wire n14197;
    wire n14200;
    wire n14203;
    wire n14206;
    wire n14209;
    wire n14212;
    wire n14215;
    wire n14218;
    wire n14221;
    wire n14224;
    wire n14227;
    wire n14230;
    wire n14233;
    wire n14236;
    wire n14239;
    wire n14242;
    wire n14245;
    wire n14248;
    wire n14251;
    wire n14254;
    wire n14257;
    wire n14260;
    wire n14263;
    wire n14266;
    wire n14269;
    wire n14272;
    wire n14275;
    wire n14278;
    wire n14281;
    wire n14284;
    wire n14287;
    wire n14290;
    wire n14293;
    wire n14296;
    wire n14299;
    wire n14302;
    wire n14305;
    wire n14308;
    wire n14311;
    wire n14314;
    wire n14317;
    wire n14320;
    wire n14323;
    wire n14326;
    wire n14329;
    wire n14333;
    wire n14336;
    wire n14338;
    wire n14341;
    wire n14344;
    wire n14347;
    wire n14350;
    wire n14353;
    wire n14356;
    wire n14359;
    wire n14362;
    wire n14366;
    wire n14369;
    wire n14372;
    wire n14374;
    wire n14377;
    wire n14380;
    wire n14383;
    wire n14386;
    wire n14389;
    wire n14392;
    wire n14395;
    wire n14398;
    wire n14401;
    wire n14404;
    wire n14407;
    wire n14410;
    wire n14413;
    wire n14416;
    wire n14419;
    wire n14422;
    wire n14425;
    wire n14428;
    wire n14431;
    wire n14434;
    wire n14437;
    wire n14441;
    wire n14444;
    wire n14446;
    wire n14449;
    wire n14452;
    wire n14455;
    wire n14458;
    wire n14461;
    wire n14464;
    wire n14467;
    wire n14470;
    wire n14473;
    wire n14476;
    wire n14479;
    wire n14482;
    wire n14485;
    wire n14488;
    wire n14491;
    wire n14494;
    wire n14497;
    wire n14500;
    wire n14503;
    wire n14506;
    wire n14509;
    wire n14513;
    wire n14516;
    wire n14519;
    wire n14521;
    wire n14524;
    wire n14527;
    wire n14530;
    wire n14533;
    wire n14536;
    wire n14539;
    wire n14542;
    wire n14545;
    wire n14548;
    wire n14551;
    wire n14554;
    wire n14557;
    wire n14560;
    wire n14563;
    wire n14566;
    wire n14569;
    wire n14572;
    wire n14575;
    wire n14578;
    wire n14581;
    wire n14584;
    wire n14587;
    wire n14590;
    wire n14593;
    wire n14596;
    wire n14599;
    wire n14602;
    wire n14605;
    wire n14608;
    wire n14611;
    wire n14614;
    wire n14617;
    wire n14620;
    wire n14623;
    wire n14626;
    wire n14629;
    wire n14632;
    wire n14635;
    wire n14638;
    wire n14641;
    wire n14644;
    wire n14647;
    wire n14650;
    wire n14653;
    wire n14656;
    wire n14659;
    wire n14662;
    wire n14665;
    wire n14668;
    wire n14671;
    wire n14674;
    wire n14677;
    wire n14680;
    wire n14683;
    wire n14686;
    wire n14689;
    wire n14692;
    wire n14695;
    wire n14698;
    wire n14701;
    wire n14704;
    wire n14707;
    wire n14710;
    wire n14713;
    wire n14716;
    wire n14719;
    wire n14722;
    wire n14725;
    wire n14728;
    wire n14731;
    wire n14734;
    wire n14737;
    wire n14740;
    wire n14743;
    wire n14746;
    wire n14749;
    wire n14752;
    wire n14755;
    wire n14758;
    wire n14761;
    wire n14764;
    wire n14767;
    wire n14770;
    wire n14773;
    wire n14776;
    wire n14779;
    wire n14782;
    wire n14785;
    wire n14788;
    wire n14791;
    wire n14794;
    wire n14797;
    wire n14800;
    wire n14803;
    wire n14806;
    wire n14809;
    wire n14812;
    wire n14815;
    wire n14818;
    wire n14821;
    wire n14824;
    wire n14827;
    wire n14830;
    wire n14833;
    wire n14836;
    wire n14839;
    wire n14843;
    wire n14846;
    wire n14849;
    wire n14851;
    wire n14854;
    wire n14857;
    wire n14860;
    wire n14863;
    wire n14866;
    wire n14869;
    wire n14872;
    wire n14875;
    wire n14878;
    wire n14881;
    wire n14884;
    wire n14887;
    wire n14890;
    wire n14893;
    wire n14896;
    wire n14899;
    wire n14902;
    wire n14905;
    wire n14908;
    wire n14911;
    wire n14914;
    wire n14917;
    wire n14920;
    wire n14923;
    wire n14926;
    wire n14929;
    wire n14932;
    wire n14935;
    wire n14938;
    wire n14941;
    wire n14944;
    wire n14947;
    wire n14950;
    wire n14953;
    wire n14956;
    wire n14959;
    wire n14962;
    wire n14966;
    wire n14969;
    wire n14972;
    wire n14974;
    wire n14977;
    wire n14980;
    wire n14983;
    wire n14986;
    wire n14989;
    wire n14992;
    wire n14995;
    wire n14998;
    wire n15001;
    wire n15004;
    wire n15007;
    wire n15010;
    wire n15013;
    wire n15016;
    wire n15019;
    wire n15022;
    wire n15025;
    wire n15028;
    wire n15031;
    wire n15034;
    wire n15037;
    wire n15040;
    wire n15043;
    wire n15046;
    wire n15049;
    wire n15052;
    wire n15055;
    wire n15058;
    wire n15061;
    wire n15064;
    wire n15068;
    wire n15070;
    wire n15073;
    wire n15076;
    wire n15079;
    wire n15082;
    wire n15085;
    wire n15088;
    wire n15091;
    wire n15094;
    wire n15097;
    wire n15100;
    wire n15103;
    wire n15106;
    wire n15109;
    wire n15112;
    wire n15115;
    wire n15118;
    wire n15121;
    wire n15124;
    wire n15127;
    wire n15130;
    wire n15133;
    wire n15136;
    wire n15139;
    wire n15142;
    wire n15145;
    wire n15148;
    wire n15151;
    wire n15154;
    wire n15157;
    wire n15160;
    wire n15163;
    wire n15166;
    wire n15169;
    wire n15172;
    wire n15175;
    wire n15178;
    wire n15181;
    wire n15184;
    wire n15187;
    wire n15190;
    wire n15193;
    wire n15196;
    wire n15199;
    wire n15202;
    wire n15205;
    wire n15208;
    wire n15211;
    wire n15214;
    wire n15217;
    wire n15220;
    wire n15223;
    wire n15226;
    wire n15229;
    wire n15232;
    wire n15235;
    wire n15238;
    wire n15241;
    wire n15244;
    wire n15247;
    wire n15250;
    wire n15253;
    wire n15256;
    wire n15259;
    wire n15262;
    wire n15265;
    wire n15268;
    wire n15271;
    wire n15274;
    wire n15277;
    wire n15280;
    wire n15283;
    wire n15286;
    wire n15289;
    wire n15292;
    wire n15295;
    wire n15298;
    wire n15301;
    wire n15304;
    wire n15307;
    wire n15310;
    wire n15313;
    wire n15316;
    wire n15319;
    wire n15322;
    wire n15325;
    wire n15328;
    wire n15331;
    wire n15334;
    wire n15337;
    wire n15340;
    wire n15343;
    wire n15346;
    wire n15349;
    wire n15352;
    wire n15356;
    wire n15358;
    wire n15361;
    wire n15364;
    wire n15367;
    wire n15370;
    wire n15373;
    wire n15376;
    wire n15379;
    wire n15382;
    wire n15385;
    wire n15388;
    wire n15391;
    wire n15394;
    wire n15397;
    wire n15400;
    wire n15403;
    wire n15406;
    wire n15409;
    wire n15412;
    wire n15415;
    wire n15418;
    wire n15421;
    wire n15424;
    wire n15427;
    wire n15430;
    wire n15433;
    wire n15436;
    wire n15439;
    wire n15442;
    wire n15445;
    wire n15448;
    wire n15451;
    wire n15454;
    wire n15457;
    wire n15460;
    wire n15463;
    wire n15466;
    wire n15469;
    wire n15473;
    wire n15475;
    wire n15478;
    wire n15481;
    wire n15484;
    wire n15487;
    wire n15490;
    wire n15493;
    wire n15496;
    wire n15500;
    wire n15503;
    wire n15506;
    wire n15508;
    wire n15511;
    wire n15514;
    wire n15517;
    wire n15521;
    wire n15524;
    wire n15527;
    wire n15530;
    wire n15533;
    wire n15536;
    wire n15539;
    wire n15542;
    wire n15545;
    wire n15548;
    wire n15551;
    wire n15554;
    wire n15557;
    wire n15560;
    wire n15563;
    wire n15566;
    wire n15569;
    wire n15572;
    wire n15575;
    wire n15578;
    wire n15581;
    wire n15584;
    wire n15587;
    wire n15590;
    wire n15593;
    wire n15596;
    wire n15599;
    wire n15602;
    wire n15605;
    wire n15608;
    wire n15611;
    wire n15614;
    wire n15617;
    wire n15620;
    wire n15623;
    wire n15625;
    wire n15628;
    wire n15631;
    wire n15634;
    wire n15637;
    wire n15640;
    wire n15643;
    wire n15646;
    wire n15649;
    wire n15652;
    wire n15655;
    wire n15658;
    wire n15661;
    wire n15664;
    wire n15668;
    wire n15671;
    wire n15674;
    wire n15677;
    wire n15679;
    wire n15682;
    wire n15685;
    wire n15688;
    wire n15691;
    wire n15694;
    wire n15697;
    wire n15701;
    wire n15704;
    wire n15707;
    wire n15710;
    wire n15713;
    wire n15716;
    wire n15719;
    wire n15722;
    wire n15725;
    wire n15727;
    wire n15730;
    wire n15733;
    wire n15736;
    wire n15739;
    wire n15742;
    wire n15745;
    wire n15748;
    wire n15751;
    wire n15754;
    wire n15757;
    wire n15760;
    wire n15763;
    wire n15766;
    wire n15769;
    wire n15773;
    wire n15776;
    wire n15779;
    wire n15782;
    wire n15785;
    wire n15788;
    wire n15791;
    wire n15794;
    wire n15797;
    wire n15800;
    wire n15803;
    wire n15806;
    wire n15809;
    wire n15812;
    wire n15815;
    wire n15817;
    wire n15821;
    wire n15824;
    wire n15827;
    wire n15830;
    wire n15833;
    wire n15836;
    wire n15839;
    wire n15842;
    wire n15845;
    wire n15848;
    wire n15850;
    wire n15853;
    wire n15856;
    wire n15859;
    wire n15862;
    wire n15865;
    wire n15868;
    wire n15871;
    wire n15874;
    wire n15877;
    wire n15880;
    wire n15883;
    wire n15886;
    wire n15889;
    wire n15892;
    wire n15895;
    wire n15898;
    wire n15901;
    wire n15904;
    wire n15907;
    wire n15911;
    wire n15914;
    wire n15917;
    wire n15920;
    wire n15923;
    wire n15926;
    wire n15929;
    wire n15931;
    wire n15934;
    wire n15937;
    wire n15940;
    wire n15943;
    wire n15946;
    wire n15949;
    wire n15952;
    wire n15955;
    wire n15958;
    wire n15961;
    wire n15964;
    wire n15967;
    wire n15970;
    wire n15973;
    wire n15976;
    wire n15979;
    wire n15982;
    wire n15985;
    wire n15988;
    wire n15992;
    wire n15994;
    wire n15998;
    wire n16001;
    wire n16003;
    wire n16006;
    wire n16009;
    wire n16012;
    wire n16015;
    wire n16018;
    wire n16021;
    wire n16024;
    wire n16027;
    wire n16030;
    wire n16033;
    wire n16036;
    wire n16039;
    wire n16042;
    wire n16045;
    wire n16048;
    wire n16051;
    wire n16054;
    wire n16057;
    wire n16060;
    wire n16063;
    wire n16066;
    wire n16069;
    wire n16072;
    wire n16075;
    wire n16078;
    wire n16081;
    wire n16084;
    wire n16087;
    wire n16090;
    wire n16093;
    wire n16096;
    wire n16099;
    wire n16102;
    wire n16105;
    wire n16108;
    wire n16111;
    wire n16114;
    wire n16117;
    wire n16120;
    wire n16124;
    wire n16126;
    wire n16129;
    wire n16132;
    wire n16135;
    wire n16138;
    wire n16141;
    wire n16144;
    wire n16147;
    wire n16150;
    wire n16153;
    wire n16156;
    wire n16159;
    wire n16162;
    wire n16165;
    wire n16168;
    wire n16171;
    wire n16174;
    wire n16177;
    wire n16181;
    wire n16183;
    wire n16186;
    wire n16189;
    wire n16192;
    wire n16195;
    wire n16198;
    wire n16201;
    wire n16204;
    wire n16207;
    wire n16210;
    wire n16213;
    wire n16216;
    wire n16219;
    wire n16222;
    wire n16225;
    wire n16228;
    wire n16231;
    wire n16234;
    wire n16237;
    wire n16240;
    wire n16243;
    wire n16246;
    wire n16249;
    wire n16252;
    wire n16255;
    wire n16258;
    wire n16261;
    wire n16264;
    wire n16267;
    wire n16270;
    wire n16273;
    wire n16276;
    wire n16279;
    wire n16282;
    wire n16285;
    wire n16289;
    wire n16292;
    wire n16295;
    wire n16298;
    wire n16300;
    wire n16303;
    wire n16306;
    wire n16309;
    wire n16313;
    wire n16316;
    wire n16319;
    wire n16322;
    wire n16324;
    wire n16328;
    wire n16330;
    wire n16333;
    wire n16336;
    wire n16339;
    wire n16342;
    wire n16346;
    wire n16349;
    wire n16351;
    wire n16354;
    wire n16357;
    wire n16360;
    wire n16363;
    wire n16366;
    wire n16369;
    wire n16372;
    wire n16375;
    wire n16378;
    wire n16381;
    wire n16384;
    wire n16387;
    wire n16390;
    wire n16393;
    wire n16396;
    wire n16399;
    wire n16403;
    wire n16406;
    wire n16409;
    wire n16412;
    wire n16415;
    wire n16418;
    wire n16421;
    wire n16424;
    wire n16427;
    wire n16430;
    wire n16433;
    wire n16436;
    wire n16439;
    wire n16442;
    wire n16445;
    wire n16447;
    wire n16450;
    wire n16453;
    wire n16456;
    wire n16459;
    wire n16462;
    wire n16465;
    wire n16469;
    wire n16472;
    wire n16475;
    wire n16478;
    wire n16481;
    wire n16484;
    wire n16487;
    wire n16490;
    wire n16493;
    wire n16496;
    wire n16499;
    wire n16502;
    wire n16505;
    wire n16507;
    wire n16510;
    wire n16513;
    wire n16516;
    wire n16519;
    wire n16522;
    wire n16525;
    wire n16528;
    wire n16531;
    wire n16534;
    wire n16537;
    wire n16540;
    wire n16543;
    wire n16546;
    wire n16549;
    wire n16552;
    wire n16555;
    wire n16558;
    wire n16561;
    wire n16564;
    wire n16567;
    wire n16570;
    wire n16573;
    wire n16576;
    wire n16579;
    wire n16582;
    wire n16585;
    wire n16588;
    wire n16591;
    wire n16594;
    wire n16597;
    wire n16600;
    wire n16603;
    wire n16606;
    wire n16609;
    wire n16612;
    wire n16615;
    wire n16618;
    wire n16621;
    wire n16624;
    wire n16627;
    wire n16630;
    wire n16633;
    wire n16636;
    wire n16639;
    wire n16643;
    wire n16646;
    wire n16649;
    wire n16652;
    wire n16655;
    wire n16658;
    wire n16661;
    wire n16664;
    wire n16666;
    wire n16669;
    wire n16672;
    wire n16675;
    wire n16678;
    wire n16681;
    wire n16684;
    wire n16687;
    wire n16690;
    wire n16693;
    wire n16696;
    wire n16699;
    wire n16702;
    wire n16705;
    wire n16708;
    wire n16711;
    wire n16714;
    wire n16717;
    wire n16720;
    wire n16723;
    wire n16726;
    wire n16729;
    wire n16732;
    wire n16735;
    wire n16738;
    wire n16741;
    wire n16744;
    wire n16747;
    wire n16750;
    wire n16753;
    wire n16756;
    wire n16759;
    wire n16762;
    wire n16765;
    wire n16768;
    wire n16771;
    wire n16774;
    wire n16777;
    wire n16780;
    wire n16783;
    wire n16786;
    wire n16789;
    wire n16792;
    wire n16795;
    wire n16798;
    wire n16801;
    wire n16804;
    wire n16807;
    wire n16810;
    wire n16813;
    wire n16816;
    wire n16819;
    wire n16822;
    wire n16825;
    wire n16829;
    wire n16832;
    wire n16835;
    wire n16838;
    wire n16840;
    wire n16843;
    wire n16846;
    wire n16849;
    wire n16853;
    wire n16856;
    wire n16858;
    wire n16861;
    wire n16864;
    wire n16867;
    wire n16870;
    wire n16873;
    wire n16876;
    wire n16879;
    wire n16882;
    wire n16885;
    wire n16888;
    wire n16891;
    wire n16894;
    wire n16897;
    wire n16900;
    wire n16903;
    wire n16906;
    wire n16909;
    wire n16912;
    wire n16915;
    wire n16918;
    wire n16921;
    wire n16924;
    wire n16927;
    wire n16930;
    wire n16933;
    wire n16936;
    wire n16939;
    wire n16942;
    wire n16945;
    wire n16948;
    wire n16951;
    wire n16954;
    wire n16957;
    wire n16960;
    wire n16963;
    wire n16966;
    wire n16969;
    wire n16972;
    wire n16975;
    wire n16978;
    wire n16981;
    wire n16984;
    wire n16987;
    wire n16990;
    wire n16993;
    wire n16996;
    wire n16999;
    wire n17002;
    wire n17006;
    wire n17009;
    wire n17012;
    wire n17015;
    wire n17017;
    wire n17020;
    wire n17023;
    wire n17026;
    wire n17029;
    wire n17032;
    wire n17035;
    wire n17038;
    wire n17041;
    wire n17044;
    wire n17047;
    wire n17050;
    wire n17053;
    wire n17056;
    wire n17059;
    wire n17062;
    wire n17065;
    wire n17068;
    wire n17071;
    wire n17074;
    wire n17078;
    wire n17081;
    wire n17084;
    wire n17087;
    wire n17089;
    wire n17092;
    wire n17095;
    wire n17098;
    wire n17101;
    wire n17104;
    wire n17107;
    wire n17110;
    wire n17113;
    wire n17116;
    wire n17119;
    wire n17122;
    wire n17125;
    wire n17128;
    wire n17131;
    wire n17134;
    wire n17137;
    wire n17140;
    wire n17143;
    wire n17146;
    wire n17149;
    wire n17152;
    wire n17155;
    wire n17159;
    wire n17162;
    wire n17165;
    wire n17168;
    wire n17171;
    wire n17174;
    wire n17176;
    wire n17179;
    wire n17182;
    wire n17185;
    wire n17189;
    wire n17192;
    wire n17195;
    wire n17198;
    wire n17201;
    wire n17204;
    wire n17207;
    wire n17210;
    wire n17213;
    wire n17216;
    wire n17219;
    wire n17222;
    wire n17225;
    wire n17228;
    wire n17231;
    wire n17234;
    wire n17237;
    wire n17240;
    wire n17242;
    wire n17245;
    wire n17248;
    wire n17251;
    wire n17254;
    wire n17257;
    wire n17260;
    wire n17263;
    wire n17266;
    wire n17269;
    wire n17272;
    wire n17275;
    wire n17278;
    wire n17281;
    wire n17284;
    wire n17287;
    wire n17290;
    wire n17293;
    wire n17296;
    wire n17299;
    wire n17302;
    wire n17305;
    wire n17308;
    wire n17311;
    wire n17314;
    wire n17317;
    wire n17320;
    wire n17323;
    wire n17326;
    wire n17329;
    wire n17332;
    wire n17335;
    wire n17338;
    wire n17341;
    wire n17344;
    wire n17347;
    wire n17350;
    wire n17353;
    wire n17356;
    wire n17359;
    wire n17362;
    wire n17365;
    wire n17368;
    wire n17371;
    wire n17374;
    wire n17377;
    wire n17380;
    wire n17384;
    wire n17387;
    wire n17390;
    wire n17393;
    wire n17396;
    wire n17399;
    wire n17402;
    wire n17405;
    wire n17408;
    wire n17411;
    wire n17414;
    wire n17417;
    wire n17420;
    wire n17423;
    wire n17425;
    wire n17428;
    wire n17432;
    wire n17435;
    wire n17438;
    wire n17441;
    wire n17444;
    wire n17447;
    wire n17450;
    wire n17453;
    wire n17456;
    wire n17459;
    wire n17461;
    wire n17464;
    wire n17467;
    wire n17471;
    wire n17473;
    wire n17476;
    wire n17479;
    wire n17482;
    wire n17485;
    wire n17489;
    wire n17492;
    wire n17494;
    wire n17498;
    wire n17501;
    wire n17504;
    wire n17507;
    wire n17510;
    wire n17513;
    wire n17515;
    wire n17518;
    wire n17521;
    wire n17524;
    wire n17527;
    wire n17530;
    wire n17533;
    wire n17536;
    wire n17539;
    wire n17542;
    wire n17545;
    wire n17548;
    wire n17551;
    wire n17554;
    wire n17557;
    wire n17561;
    wire n17564;
    wire n17566;
    wire n17569;
    wire n17572;
    wire n17575;
    wire n17578;
    wire n17582;
    wire n17585;
    wire n17587;
    wire n17590;
    wire n17593;
    wire n17596;
    wire n17599;
    wire n17602;
    wire n17605;
    wire n17608;
    wire n17611;
    wire n17614;
    wire n17617;
    wire n17620;
    wire n17623;
    wire n17626;
    wire n17629;
    wire n17632;
    wire n17635;
    wire n17638;
    wire n17641;
    wire n17644;
    wire n17647;
    wire n17650;
    wire n17653;
    wire n17656;
    wire n17659;
    wire n17662;
    wire n17665;
    wire n17668;
    wire n17671;
    wire n17674;
    wire n17677;
    wire n17680;
    wire n17683;
    wire n17686;
    wire n17690;
    wire n17693;
    wire n17696;
    wire n17699;
    wire n17701;
    wire n17704;
    wire n17707;
    wire n17711;
    wire n17713;
    wire n17716;
    wire n17719;
    wire n17722;
    wire n17725;
    wire n17729;
    wire n17731;
    wire n17734;
    wire n17737;
    wire n17740;
    wire n17743;
    wire n17746;
    wire n17749;
    wire n17753;
    wire n17756;
    wire n17759;
    wire n17761;
    wire n17764;
    wire n17767;
    wire n17771;
    wire n17774;
    wire n17777;
    wire n17780;
    wire n17783;
    wire n17786;
    wire n17789;
    wire n17792;
    wire n17795;
    wire n17798;
    wire n17801;
    wire n17803;
    wire n17806;
    wire n17809;
    wire n17812;
    wire n17815;
    wire n17818;
    wire n17821;
    wire n17824;
    wire n17827;
    wire n17830;
    wire n17833;
    wire n17836;
    wire n17839;
    wire n17842;
    wire n17845;
    wire n17848;
    wire n17851;
    wire n17854;
    wire n17857;
    wire n17860;
    wire n17863;
    wire n17866;
    wire n17869;
    wire n17872;
    wire n17875;
    wire n17878;
    wire n17881;
    wire n17884;
    wire n17887;
    wire n17890;
    wire n17893;
    wire n17896;
    wire n17899;
    wire n17902;
    wire n17905;
    wire n17908;
    wire n17911;
    wire n17915;
    wire n17918;
    wire n17921;
    wire n17924;
    wire n17927;
    wire n17929;
    wire n17932;
    wire n17935;
    wire n17938;
    wire n17941;
    wire n17944;
    wire n17947;
    wire n17950;
    wire n17953;
    wire n17956;
    wire n17959;
    wire n17962;
    wire n17965;
    wire n17968;
    wire n17971;
    wire n17975;
    wire n17978;
    wire n17980;
    wire n17983;
    wire n17987;
    wire n17990;
    wire n17993;
    wire n17996;
    wire n17998;
    wire n18001;
    wire n18004;
    wire n18007;
    wire n18010;
    wire n18013;
    wire n18016;
    wire n18019;
    wire n18022;
    wire n18025;
    wire n18028;
    wire n18031;
    wire n18034;
    wire n18037;
    wire n18040;
    wire n18043;
    wire n18046;
    wire n18050;
    wire n18053;
    wire n18055;
    wire n18058;
    wire n18061;
    wire n18064;
    wire n18067;
    wire n18070;
    wire n18073;
    wire n18076;
    wire n18079;
    wire n18082;
    wire n18085;
    wire n18088;
    wire n18091;
    wire n18094;
    wire n18097;
    wire n18100;
    wire n18103;
    wire n18107;
    wire n18110;
    wire n18112;
    wire n18115;
    wire n18118;
    wire n18121;
    wire n18124;
    wire n18127;
    wire n18130;
    wire n18133;
    wire n18136;
    wire n18139;
    wire n18142;
    wire n18145;
    wire n18148;
    wire n18151;
    wire n18155;
    wire n18158;
    wire n18161;
    wire n18163;
    wire n18166;
    wire n18169;
    wire n18172;
    wire n18175;
    wire n18178;
    wire n18181;
    wire n18184;
    wire n18188;
    wire n18191;
    wire n18194;
    wire n18197;
    wire n18200;
    wire n18203;
    wire n18206;
    wire n18209;
    wire n18212;
    wire n18215;
    wire n18218;
    wire n18221;
    wire n18224;
    wire n18226;
    wire n18229;
    wire n18232;
    wire n18235;
    wire n18238;
    wire n18241;
    wire n18244;
    wire n18247;
    wire n18250;
    wire n18253;
    wire n18256;
    wire n18259;
    wire n18262;
    wire n18265;
    wire n18268;
    wire n18271;
    wire n18274;
    wire n18277;
    wire n18280;
    wire n18283;
    wire n18286;
    wire n18289;
    wire n18292;
    wire n18295;
    wire n18298;
    wire n18301;
    wire n18304;
    wire n18307;
    wire n18310;
    wire n18313;
    wire n18316;
    wire n18319;
    wire n18322;
    wire n18326;
    wire n18329;
    wire n18331;
    wire n18334;
    wire n18337;
    wire n18340;
    wire n18343;
    wire n18347;
    wire n18349;
    wire n18352;
    wire n18355;
    wire n18358;
    wire n18361;
    wire n18364;
    wire n18367;
    wire n18370;
    wire n18373;
    wire n18376;
    wire n18379;
    wire n18382;
    wire n18385;
    wire n18389;
    wire n18391;
    wire n18394;
    wire n18397;
    wire n18400;
    wire n18403;
    wire n18406;
    wire n18409;
    wire n18412;
    wire n18415;
    wire n18419;
    wire n18422;
    wire n18424;
    wire n18427;
    wire n18430;
    wire n18433;
    wire n18436;
    wire n18439;
    wire n18442;
    wire n18445;
    wire n18448;
    wire n18451;
    wire n18454;
    wire n18457;
    wire n18460;
    wire n18463;
    wire n18466;
    wire n18470;
    wire n18473;
    wire n18475;
    wire n18478;
    wire n18481;
    wire n18484;
    wire n18487;
    wire n18490;
    wire n18493;
    wire n18496;
    wire n18499;
    wire n18502;
    wire n18505;
    wire n18508;
    wire n18511;
    wire n18514;
    wire n18517;
    wire n18520;
    wire n18523;
    wire n18526;
    wire n18529;
    wire n18532;
    wire n18535;
    wire n18539;
    wire n18542;
    wire n18544;
    wire n18547;
    wire n18550;
    wire n18553;
    wire n18556;
    wire n18559;
    wire n18562;
    wire n18565;
    wire n18568;
    wire n18571;
    wire n18574;
    wire n18577;
    wire n18580;
    wire n18583;
    wire n18586;
    wire n18589;
    wire n18592;
    wire n18595;
    wire n18598;
    wire n18601;
    wire n18604;
    wire n18607;
    wire n18610;
    wire n18613;
    wire n18616;
    wire n18619;
    wire n18622;
    wire n18625;
    wire n18628;
    wire n18631;
    wire n18634;
    wire n18637;
    wire n18640;
    wire n18643;
    wire n18646;
    wire n18649;
    wire n18652;
    wire n18655;
    wire n18658;
    wire n18661;
    wire n18664;
    wire n18667;
    wire n18670;
    wire n18673;
    wire n18676;
    wire n18679;
    wire n18685;
    wire n18688;
    wire n18691;
    wire n18694;
    wire n18697;
    wire n18700;
    wire n18703;
    wire n18706;
    wire n18709;
    wire n18712;
    wire n18715;
    wire n18718;
    wire n18721;
    wire n18724;
    wire n18727;
    wire n18730;
    wire n18733;
    wire n18736;
    wire n18739;
    wire n18742;
    wire n18745;
    wire n18748;
    wire n18751;
    wire n18754;
    wire n18757;
    wire n18760;
    wire n18763;
    wire n18766;
    wire n18769;
    wire n18772;
    wire n18775;
    wire n18778;
    wire n18781;
    wire n18784;
    wire n18787;
    wire n18790;
    wire n18793;
    wire n18799;
    wire n18802;
    wire n18805;
    wire n18808;
    wire n18811;
    wire n18814;
    wire n18817;
    wire n18820;
    wire n18823;
    wire n18826;
    wire n18829;
    wire n18832;
    wire n18835;
    wire n18838;
    wire n18841;
    wire n18844;
    wire n18847;
    wire n18850;
    wire n18853;
    wire n18856;
    wire n18859;
    wire n18862;
    wire n18865;
    wire n18868;
    wire n18871;
    wire n18874;
    wire n18877;
    wire n18880;
    wire n18883;
    wire n18886;
    wire n18889;
    wire n18892;
    wire n18895;
    wire n18898;
    wire n18901;
    wire n18904;
    wire n18907;
    wire n18913;
    wire n18916;
    wire n18919;
    wire n18922;
    wire n18925;
    wire n18928;
    wire n18931;
    wire n18934;
    wire n18937;
    wire n18940;
    wire n18943;
    wire n18946;
    wire n18949;
    wire n18952;
    wire n18955;
    wire n18958;
    wire n18961;
    wire n18964;
    wire n18967;
    wire n18970;
    wire n18973;
    wire n18976;
    wire n18979;
    wire n18982;
    wire n18985;
    wire n18988;
    wire n18991;
    wire n18994;
    wire n18997;
    wire n19000;
    wire n19003;
    wire n19006;
    wire n19009;
    wire n19012;
    wire n19015;
    wire n19018;
    wire n19021;
    wire n19027;
    wire n19030;
    wire n19033;
    wire n19036;
    wire n19039;
    wire n19042;
    wire n19045;
    wire n19048;
    wire n19051;
    wire n19054;
    wire n19057;
    wire n19060;
    wire n19063;
    wire n19066;
    wire n19069;
    wire n19072;
    wire n19075;
    wire n19078;
    wire n19081;
    wire n19084;
    wire n19087;
    wire n19090;
    wire n19093;
    wire n19096;
    wire n19099;
    wire n19102;
    wire n19105;
    wire n19108;
    wire n19111;
    wire n19114;
    wire n19117;
    wire n19120;
    wire n19123;
    wire n19126;
    wire n19129;
    wire n19132;
    wire n19135;
    wire n19141;
    wire n19144;
    wire n19147;
    wire n19150;
    wire n19153;
    wire n19156;
    wire n19159;
    wire n19162;
    wire n19165;
    wire n19168;
    wire n19171;
    wire n19174;
    wire n19177;
    wire n19180;
    wire n19183;
    wire n19186;
    wire n19189;
    wire n19192;
    wire n19195;
    wire n19198;
    wire n19201;
    wire n19204;
    wire n19207;
    wire n19210;
    wire n19213;
    wire n19216;
    wire n19219;
    wire n19222;
    wire n19225;
    wire n19228;
    wire n19231;
    wire n19234;
    wire n19237;
    wire n19240;
    wire n19243;
    wire n19246;
    wire n19249;
    wire n19255;
    wire n19258;
    wire n19261;
    wire n19264;
    wire n19267;
    wire n19270;
    wire n19273;
    wire n19276;
    wire n19279;
    wire n19282;
    wire n19285;
    wire n19288;
    wire n19291;
    wire n19294;
    wire n19297;
    wire n19300;
    wire n19303;
    wire n19306;
    wire n19309;
    wire n19312;
    wire n19315;
    wire n19318;
    wire n19321;
    wire n19324;
    wire n19327;
    wire n19330;
    wire n19333;
    wire n19336;
    wire n19339;
    wire n19342;
    wire n19345;
    wire n19348;
    wire n19351;
    wire n19354;
    wire n19357;
    wire n19360;
    wire n19363;
    wire n19369;
    wire n19372;
    wire n19375;
    wire n19378;
    wire n19381;
    wire n19384;
    wire n19387;
    wire n19390;
    wire n19393;
    wire n19396;
    wire n19399;
    wire n19402;
    wire n19405;
    wire n19408;
    wire n19411;
    wire n19414;
    wire n19417;
    wire n19420;
    wire n19423;
    wire n19426;
    wire n19429;
    wire n19432;
    wire n19435;
    wire n19438;
    wire n19441;
    wire n19444;
    wire n19447;
    wire n19450;
    wire n19453;
    wire n19456;
    wire n19459;
    wire n19462;
    wire n19465;
    wire n19468;
    wire n19471;
    wire n19474;
    wire n19477;
    wire n19483;
    wire n19486;
    wire n19489;
    wire n19492;
    wire n19495;
    wire n19498;
    wire n19501;
    wire n19504;
    wire n19507;
    wire n19510;
    wire n19513;
    wire n19516;
    wire n19519;
    wire n19522;
    wire n19525;
    wire n19528;
    wire n19531;
    wire n19534;
    wire n19537;
    wire n19540;
    wire n19543;
    wire n19546;
    wire n19549;
    wire n19552;
    wire n19555;
    wire n19558;
    wire n19561;
    wire n19564;
    wire n19567;
    wire n19570;
    wire n19573;
    wire n19576;
    wire n19579;
    wire n19582;
    wire n19585;
    wire n19588;
    wire n19591;
    wire n19597;
    wire n19600;
    wire n19603;
    wire n19606;
    wire n19609;
    wire n19612;
    wire n19615;
    wire n19618;
    wire n19621;
    wire n19624;
    wire n19627;
    wire n19630;
    wire n19633;
    wire n19636;
    wire n19639;
    wire n19642;
    wire n19645;
    wire n19648;
    wire n19651;
    wire n19654;
    wire n19657;
    wire n19660;
    wire n19663;
    wire n19666;
    wire n19669;
    wire n19672;
    wire n19675;
    wire n19678;
    wire n19681;
    wire n19684;
    wire n19687;
    wire n19690;
    wire n19693;
    wire n19696;
    wire n19699;
    wire n19702;
    wire n19705;
    wire n19711;
    wire n19714;
    wire n19717;
    wire n19720;
    wire n19723;
    wire n19726;
    wire n19729;
    wire n19732;
    wire n19735;
    wire n19738;
    wire n19741;
    wire n19744;
    wire n19747;
    wire n19750;
    wire n19753;
    wire n19756;
    wire n19759;
    wire n19762;
    wire n19765;
    wire n19768;
    wire n19771;
    wire n19774;
    wire n19777;
    wire n19780;
    wire n19783;
    wire n19786;
    wire n19789;
    wire n19792;
    wire n19795;
    wire n19798;
    wire n19801;
    wire n19804;
    wire n19807;
    wire n19810;
    wire n19813;
    wire n19816;
    wire n19819;
    wire n19825;
    wire n19828;
    wire n19831;
    wire n19834;
    wire n19837;
    wire n19840;
    wire n19843;
    wire n19846;
    wire n19849;
    wire n19852;
    wire n19855;
    wire n19858;
    wire n19861;
    wire n19864;
    wire n19867;
    wire n19870;
    wire n19873;
    wire n19876;
    wire n19879;
    wire n19882;
    wire n19885;
    wire n19888;
    wire n19891;
    wire n19894;
    wire n19897;
    wire n19900;
    wire n19903;
    wire n19906;
    wire n19909;
    wire n19912;
    wire n19915;
    wire n19918;
    wire n19921;
    wire n19924;
    wire n19927;
    wire n19930;
    wire n19933;
    wire n19939;
    wire n19942;
    wire n19945;
    wire n19948;
    wire n19951;
    wire n19954;
    wire n19957;
    wire n19960;
    wire n19963;
    wire n19966;
    wire n19969;
    wire n19972;
    wire n19975;
    wire n19978;
    wire n19981;
    wire n19984;
    wire n19987;
    wire n19990;
    wire n19993;
    wire n19996;
    wire n19999;
    wire n20002;
    wire n20005;
    wire n20008;
    wire n20011;
    wire n20014;
    wire n20017;
    wire n20020;
    wire n20023;
    wire n20026;
    wire n20029;
    wire n20032;
    wire n20035;
    wire n20038;
    wire n20041;
    wire n20044;
    wire n20047;
    wire n20053;
    wire n20056;
    wire n20059;
    wire n20062;
    wire n20065;
    wire n20068;
    wire n20071;
    wire n20074;
    wire n20077;
    wire n20080;
    wire n20083;
    wire n20086;
    wire n20089;
    wire n20092;
    wire n20095;
    wire n20098;
    wire n20101;
    wire n20104;
    wire n20107;
    wire n20110;
    wire n20113;
    wire n20116;
    wire n20119;
    wire n20122;
    wire n20125;
    wire n20128;
    wire n20131;
    wire n20134;
    wire n20137;
    wire n20140;
    wire n20143;
    wire n20146;
    wire n20149;
    wire n20152;
    wire n20155;
    wire n20158;
    wire n20161;
    wire n20167;
    wire n20170;
    wire n20173;
    wire n20176;
    wire n20179;
    wire n20182;
    wire n20185;
    wire n20188;
    wire n20191;
    wire n20194;
    wire n20197;
    wire n20200;
    wire n20203;
    wire n20206;
    wire n20209;
    wire n20212;
    wire n20215;
    wire n20218;
    wire n20221;
    wire n20224;
    wire n20227;
    wire n20230;
    wire n20233;
    wire n20236;
    wire n20239;
    wire n20242;
    wire n20245;
    wire n20248;
    wire n20251;
    wire n20254;
    wire n20257;
    wire n20260;
    wire n20263;
    wire n20266;
    wire n20269;
    wire n20272;
    wire n20275;
    wire n20281;
    wire n20284;
    wire n20287;
    wire n20290;
    wire n20293;
    wire n20296;
    wire n20299;
    wire n20302;
    wire n20305;
    wire n20308;
    wire n20311;
    wire n20314;
    wire n20317;
    wire n20320;
    wire n20323;
    wire n20326;
    wire n20329;
    wire n20332;
    wire n20335;
    wire n20338;
    wire n20341;
    wire n20344;
    wire n20347;
    wire n20350;
    wire n20353;
    wire n20356;
    wire n20359;
    wire n20362;
    wire n20365;
    wire n20368;
    wire n20371;
    wire n20374;
    wire n20377;
    wire n20380;
    wire n20383;
    wire n20386;
    wire n20389;
    wire n20395;
    wire n20398;
    wire n20401;
    wire n20404;
    wire n20407;
    wire n20410;
    wire n20413;
    wire n20416;
    wire n20419;
    wire n20422;
    wire n20425;
    wire n20428;
    wire n20431;
    wire n20434;
    wire n20437;
    wire n20440;
    wire n20443;
    wire n20446;
    wire n20449;
    wire n20452;
    wire n20455;
    wire n20458;
    wire n20461;
    wire n20464;
    wire n20467;
    wire n20470;
    wire n20473;
    wire n20476;
    wire n20479;
    wire n20482;
    wire n20485;
    wire n20488;
    wire n20491;
    wire n20494;
    wire n20497;
    wire n20500;
    wire n20503;
    wire n20509;
    wire n20512;
    wire n20515;
    wire n20518;
    wire n20521;
    wire n20524;
    wire n20527;
    wire n20530;
    wire n20533;
    wire n20536;
    wire n20539;
    wire n20542;
    wire n20545;
    wire n20548;
    wire n20551;
    wire n20554;
    wire n20557;
    wire n20560;
    wire n20563;
    wire n20566;
    wire n20569;
    wire n20572;
    wire n20575;
    wire n20578;
    wire n20581;
    wire n20584;
    wire n20587;
    wire n20590;
    wire n20593;
    wire n20596;
    wire n20599;
    wire n20602;
    wire n20605;
    wire n20608;
    wire n20611;
    wire n20614;
    wire n20617;
    wire n20623;
    wire n20626;
    wire n20629;
    wire n20632;
    wire n20635;
    wire n20638;
    wire n20641;
    wire n20644;
    wire n20647;
    wire n20650;
    wire n20653;
    wire n20656;
    wire n20659;
    wire n20662;
    wire n20665;
    wire n20668;
    wire n20671;
    wire n20674;
    wire n20677;
    wire n20680;
    wire n20683;
    wire n20686;
    wire n20689;
    wire n20692;
    wire n20695;
    wire n20698;
    wire n20701;
    wire n20704;
    wire n20707;
    wire n20710;
    wire n20713;
    wire n20716;
    wire n20719;
    wire n20722;
    wire n20725;
    wire n20728;
    wire n20731;
    wire n20737;
    wire n20740;
    wire n20743;
    wire n20746;
    wire n20749;
    wire n20752;
    wire n20755;
    wire n20758;
    wire n20761;
    wire n20764;
    wire n20767;
    wire n20770;
    wire n20773;
    wire n20776;
    wire n20779;
    wire n20782;
    wire n20785;
    wire n20788;
    wire n20791;
    wire n20794;
    wire n20797;
    wire n20800;
    wire n20803;
    wire n20806;
    wire n20809;
    wire n20812;
    wire n20815;
    wire n20818;
    wire n20821;
    wire n20824;
    wire n20827;
    wire n20830;
    wire n20833;
    wire n20836;
    wire n20839;
    wire n20842;
    wire n20845;
    wire n20851;
    wire n20854;
    wire n20857;
    wire n20860;
    wire n20863;
    wire n20866;
    wire n20869;
    wire n20872;
    wire n20875;
    wire n20878;
    wire n20881;
    wire n20884;
    wire n20887;
    wire n20890;
    wire n20893;
    wire n20896;
    wire n20899;
    wire n20902;
    wire n20905;
    wire n20908;
    wire n20911;
    wire n20914;
    wire n20917;
    wire n20920;
    wire n20923;
    wire n20926;
    wire n20929;
    wire n20932;
    wire n20935;
    wire n20938;
    wire n20941;
    wire n20944;
    wire n20947;
    wire n20950;
    wire n20953;
    wire n20956;
    wire n20959;
    wire n20965;
    wire n20968;
    wire n20971;
    wire n20974;
    wire n20977;
    wire n20980;
    wire n20983;
    wire n20986;
    wire n20989;
    wire n20992;
    wire n20995;
    wire n20998;
    wire n21001;
    wire n21004;
    wire n21007;
    wire n21010;
    wire n21013;
    wire n21016;
    wire n21019;
    wire n21022;
    wire n21025;
    wire n21028;
    wire n21031;
    wire n21034;
    wire n21037;
    wire n21040;
    wire n21043;
    wire n21046;
    wire n21049;
    wire n21052;
    wire n21055;
    wire n21058;
    wire n21061;
    wire n21064;
    wire n21067;
    wire n21070;
    wire n21073;
    wire n21079;
    wire n21082;
    wire n21085;
    wire n21088;
    wire n21091;
    wire n21094;
    wire n21097;
    wire n21100;
    wire n21103;
    wire n21106;
    wire n21109;
    wire n21112;
    wire n21115;
    wire n21118;
    wire n21121;
    wire n21124;
    wire n21127;
    wire n21130;
    wire n21133;
    wire n21136;
    wire n21139;
    wire n21142;
    wire n21145;
    wire n21148;
    wire n21151;
    wire n21154;
    wire n21157;
    wire n21160;
    wire n21163;
    wire n21166;
    wire n21169;
    wire n21172;
    wire n21175;
    wire n21178;
    wire n21181;
    wire n21184;
    wire n21187;
    wire n21193;
    wire n21196;
    wire n21199;
    wire n21202;
    wire n21205;
    wire n21208;
    wire n21211;
    wire n21214;
    wire n21217;
    wire n21220;
    wire n21223;
    wire n21226;
    wire n21229;
    wire n21232;
    wire n21235;
    wire n21238;
    wire n21241;
    wire n21244;
    wire n21247;
    wire n21250;
    wire n21253;
    wire n21256;
    wire n21259;
    wire n21262;
    wire n21265;
    wire n21268;
    wire n21271;
    wire n21274;
    wire n21277;
    wire n21280;
    wire n21283;
    wire n21286;
    wire n21289;
    wire n21292;
    wire n21295;
    wire n21298;
    wire n21301;
    wire n21307;
    wire n21310;
    wire n21313;
    wire n21316;
    wire n21319;
    wire n21322;
    wire n21325;
    wire n21328;
    wire n21331;
    wire n21334;
    wire n21337;
    wire n21340;
    wire n21343;
    wire n21346;
    wire n21349;
    wire n21352;
    wire n21355;
    wire n21358;
    wire n21361;
    wire n21364;
    wire n21367;
    wire n21370;
    wire n21373;
    wire n21376;
    wire n21379;
    wire n21382;
    wire n21385;
    wire n21388;
    wire n21391;
    wire n21394;
    wire n21397;
    wire n21400;
    wire n21403;
    wire n21406;
    wire n21409;
    wire n21412;
    wire n21415;
    wire n21421;
    wire n21424;
    wire n21427;
    wire n21430;
    wire n21433;
    wire n21436;
    wire n21439;
    wire n21442;
    wire n21445;
    wire n21448;
    wire n21451;
    wire n21454;
    wire n21457;
    wire n21460;
    wire n21463;
    wire n21466;
    wire n21469;
    wire n21472;
    wire n21475;
    wire n21478;
    wire n21481;
    wire n21484;
    wire n21487;
    wire n21490;
    wire n21493;
    wire n21496;
    wire n21499;
    wire n21502;
    wire n21505;
    wire n21508;
    wire n21511;
    wire n21514;
    wire n21517;
    wire n21520;
    wire n21523;
    wire n21526;
    wire n21529;
    wire n21535;
    wire n21538;
    wire n21541;
    wire n21544;
    wire n21547;
    wire n21550;
    wire n21553;
    wire n21556;
    wire n21559;
    wire n21562;
    wire n21565;
    wire n21568;
    wire n21571;
    wire n21574;
    wire n21577;
    wire n21580;
    wire n21583;
    wire n21586;
    wire n21589;
    wire n21592;
    wire n21595;
    wire n21598;
    wire n21601;
    wire n21604;
    wire n21607;
    wire n21610;
    wire n21613;
    wire n21616;
    wire n21619;
    wire n21622;
    wire n21625;
    wire n21628;
    wire n21631;
    wire n21634;
    wire n21637;
    wire n21640;
    wire n21643;
    wire n21649;
    wire n21652;
    wire n21655;
    wire n21658;
    wire n21661;
    wire n21664;
    wire n21667;
    wire n21670;
    wire n21673;
    wire n21676;
    wire n21679;
    wire n21682;
    wire n21685;
    wire n21688;
    wire n21691;
    wire n21694;
    wire n21697;
    wire n21700;
    wire n21703;
    wire n21706;
    wire n21709;
    wire n21712;
    wire n21715;
    wire n21718;
    wire n21721;
    wire n21724;
    wire n21727;
    wire n21730;
    wire n21733;
    wire n21736;
    wire n21739;
    wire n21742;
    wire n21745;
    wire n21748;
    wire n21751;
    wire n21754;
    wire n21757;
    wire n21763;
    wire n21766;
    wire n21769;
    wire n21772;
    wire n21775;
    wire n21778;
    wire n21781;
    wire n21784;
    wire n21787;
    wire n21790;
    wire n21793;
    wire n21796;
    wire n21799;
    wire n21802;
    wire n21805;
    wire n21808;
    wire n21811;
    wire n21814;
    wire n21817;
    wire n21820;
    wire n21823;
    wire n21826;
    wire n21829;
    wire n21832;
    wire n21835;
    wire n21838;
    wire n21841;
    wire n21844;
    wire n21847;
    wire n21850;
    wire n21853;
    wire n21856;
    wire n21859;
    wire n21862;
    wire n21865;
    wire n21868;
    wire n21871;
    wire n21877;
    wire n21880;
    wire n21883;
    wire n21886;
    wire n21889;
    wire n21892;
    wire n21895;
    wire n21898;
    wire n21901;
    wire n21904;
    wire n21907;
    wire n21910;
    wire n21913;
    wire n21916;
    wire n21919;
    wire n21922;
    wire n21925;
    wire n21928;
    wire n21931;
    wire n21934;
    wire n21937;
    wire n21940;
    wire n21943;
    wire n21946;
    wire n21949;
    wire n21952;
    wire n21955;
    wire n21958;
    wire n21961;
    wire n21964;
    wire n21967;
    wire n21970;
    wire n21973;
    wire n21976;
    wire n21979;
    wire n21982;
    wire n21985;
    wire n21991;
    wire n21994;
    wire n21997;
    wire n22000;
    wire n22003;
    wire n22006;
    wire n22009;
    wire n22012;
    wire n22015;
    wire n22018;
    wire n22021;
    wire n22024;
    wire n22027;
    wire n22030;
    wire n22033;
    wire n22036;
    wire n22039;
    wire n22042;
    wire n22045;
    wire n22048;
    wire n22051;
    wire n22054;
    wire n22057;
    wire n22060;
    wire n22063;
    wire n22066;
    wire n22069;
    wire n22072;
    wire n22075;
    wire n22078;
    wire n22081;
    wire n22084;
    wire n22087;
    wire n22090;
    wire n22093;
    wire n22096;
    wire n22099;
    wire n22105;
    wire n22108;
    wire n22111;
    wire n22114;
    wire n22117;
    wire n22120;
    wire n22123;
    wire n22126;
    wire n22129;
    wire n22132;
    wire n22135;
    wire n22138;
    wire n22141;
    wire n22144;
    wire n22147;
    wire n22150;
    wire n22153;
    wire n22156;
    wire n22159;
    wire n22162;
    wire n22165;
    wire n22168;
    wire n22171;
    wire n22174;
    wire n22177;
    wire n22180;
    wire n22183;
    wire n22186;
    wire n22189;
    wire n22192;
    wire n22195;
    wire n22198;
    wire n22201;
    wire n22204;
    wire n22207;
    wire n22210;
    wire n22213;
    wire n22219;
    wire n22222;
    wire n22225;
    wire n22228;
    wire n22231;
    wire n22234;
    wire n22237;
    wire n22240;
    wire n22243;
    wire n22246;
    wire n22249;
    wire n22252;
    wire n22255;
    wire n22258;
    wire n22261;
    wire n22264;
    wire n22267;
    wire n22270;
    wire n22273;
    wire n22276;
    wire n22279;
    wire n22282;
    wire n22285;
    wire n22288;
    wire n22291;
    wire n22294;
    wire n22297;
    wire n22300;
    wire n22303;
    wire n22306;
    wire n22309;
    wire n22312;
    wire n22315;
    wire n22318;
    wire n22321;
    wire n22324;
    wire n22327;
    wire n22333;
    wire n22336;
    wire n22339;
    wire n22342;
    wire n22345;
    wire n22348;
    wire n22351;
    wire n22354;
    wire n22357;
    wire n22360;
    wire n22363;
    wire n22366;
    wire n22369;
    wire n22372;
    wire n22375;
    wire n22378;
    wire n22381;
    wire n22384;
    wire n22387;
    wire n22390;
    wire n22393;
    wire n22396;
    wire n22399;
    wire n22402;
    wire n22405;
    wire n22408;
    wire n22411;
    wire n22414;
    wire n22417;
    wire n22420;
    wire n22423;
    wire n22426;
    wire n22429;
    wire n22432;
    wire n22435;
    wire n22438;
    wire n22441;
    wire n22447;
    wire n22450;
    wire n22453;
    wire n22456;
    wire n22459;
    wire n22462;
    wire n22465;
    wire n22468;
    wire n22471;
    wire n22474;
    wire n22477;
    wire n22480;
    wire n22483;
    wire n22486;
    wire n22489;
    wire n22492;
    wire n22495;
    wire n22498;
    wire n22501;
    wire n22504;
    wire n22507;
    wire n22510;
    wire n22513;
    wire n22516;
    wire n22519;
    wire n22522;
    wire n22525;
    wire n22528;
    wire n22531;
    wire n22534;
    wire n22537;
    wire n22540;
    wire n22543;
    wire n22546;
    wire n22549;
    wire n22552;
    wire n22555;
    wire n22561;
    wire n22564;
    wire n22567;
    wire n22570;
    wire n22573;
    wire n22576;
    wire n22579;
    wire n22582;
    wire n22585;
    wire n22588;
    wire n22591;
    wire n22594;
    wire n22597;
    wire n22600;
    wire n22603;
    wire n22606;
    wire n22609;
    wire n22612;
    wire n22615;
    wire n22618;
    wire n22621;
    wire n22624;
    wire n22627;
    wire n22630;
    wire n22633;
    wire n22636;
    wire n22639;
    wire n22642;
    wire n22645;
    wire n22648;
    wire n22651;
    wire n22654;
    wire n22657;
    wire n22660;
    wire n22663;
    wire n22666;
    wire n22669;
    wire n22675;
    wire n22678;
    wire n22681;
    wire n22684;
    wire n22687;
    wire n22690;
    wire n22693;
    wire n22696;
    wire n22699;
    wire n22702;
    wire n22705;
    wire n22708;
    wire n22711;
    wire n22714;
    wire n22717;
    wire n22720;
    wire n22723;
    wire n22726;
    wire n22729;
    wire n22732;
    wire n22735;
    wire n22738;
    wire n22741;
    wire n22744;
    wire n22747;
    wire n22750;
    wire n22753;
    wire n22756;
    wire n22759;
    wire n22762;
    wire n22765;
    wire n22768;
    wire n22771;
    wire n22774;
    wire n22777;
    wire n22780;
    wire n22783;
    wire n22789;
    wire n22792;
    wire n22795;
    wire n22798;
    wire n22801;
    wire n22804;
    wire n22807;
    wire n22810;
    wire n22813;
    wire n22816;
    wire n22819;
    wire n22822;
    wire n22825;
    wire n22828;
    wire n22831;
    wire n22834;
    wire n22837;
    wire n22840;
    wire n22843;
    wire n22846;
    wire n22849;
    wire n22852;
    wire n22855;
    wire n22858;
    wire n22861;
    wire n22864;
    wire n22867;
    wire n22870;
    wire n22873;
    wire n22876;
    wire n22879;
    wire n22882;
    wire n22885;
    wire n22888;
    wire n22891;
    wire n22894;
    wire n22897;
    wire n22903;
    wire n22906;
    wire n22909;
    wire n22912;
    wire n22915;
    wire n22918;
    wire n22921;
    wire n22924;
    wire n22927;
    wire n22930;
    wire n22933;
    wire n22936;
    wire n22939;
    wire n22942;
    wire n22945;
    wire n22948;
    wire n22951;
    wire n22954;
    wire n22957;
    wire n22960;
    wire n22963;
    wire n22966;
    wire n22969;
    wire n22972;
    wire n22975;
    wire n22978;
    wire n22981;
    wire n22984;
    wire n22987;
    wire n22990;
    wire n22993;
    wire n22996;
    wire n22999;
    wire n23002;
    wire n23005;
    wire n23008;
    wire n23011;
    wire n23017;
    wire n23020;
    wire n23023;
    wire n23026;
    wire n23029;
    wire n23032;
    wire n23035;
    wire n23038;
    wire n23041;
    wire n23044;
    wire n23047;
    wire n23050;
    wire n23053;
    wire n23056;
    wire n23059;
    wire n23062;
    wire n23065;
    wire n23068;
    wire n23071;
    wire n23074;
    wire n23077;
    wire n23080;
    wire n23083;
    wire n23086;
    wire n23089;
    wire n23092;
    wire n23095;
    wire n23098;
    wire n23101;
    wire n23104;
    wire n23107;
    wire n23110;
    wire n23113;
    wire n23116;
    wire n23119;
    wire n23122;
    wire n23125;
    wire n23131;
    wire n23134;
    wire n23137;
    wire n23140;
    wire n23143;
    wire n23146;
    wire n23149;
    wire n23152;
    wire n23155;
    wire n23158;
    wire n23161;
    wire n23164;
    wire n23167;
    wire n23170;
    wire n23173;
    wire n23176;
    wire n23179;
    wire n23182;
    wire n23185;
    wire n23188;
    wire n23191;
    wire n23194;
    wire n23197;
    wire n23200;
    wire n23203;
    wire n23206;
    wire n23209;
    wire n23212;
    wire n23215;
    wire n23218;
    wire n23221;
    wire n23224;
    wire n23227;
    wire n23230;
    wire n23233;
    wire n23236;
    wire n23239;
    wire n23245;
    wire n23248;
    wire n23251;
    wire n23254;
    wire n23257;
    wire n23260;
    wire n23263;
    wire n23266;
    wire n23269;
    wire n23272;
    wire n23275;
    wire n23278;
    wire n23281;
    wire n23284;
    wire n23287;
    wire n23290;
    wire n23293;
    wire n23296;
    wire n23299;
    wire n23302;
    wire n23305;
    wire n23308;
    wire n23311;
    wire n23314;
    wire n23317;
    wire n23320;
    wire n23323;
    wire n23326;
    wire n23329;
    wire n23332;
    wire n23335;
    wire n23338;
    wire n23341;
    wire n23344;
    wire n23347;
    wire n23353;
    wire n23356;
    wire n23359;
    wire n23362;
    wire n23365;
    wire n23368;
    wire n23371;
    wire n23374;
    wire n23377;
    wire n23380;
    wire n23383;
    wire n23386;
    wire n23389;
    wire n23392;
    wire n23395;
    wire n23398;
    wire n23401;
    wire n23404;
    wire n23407;
    wire n23410;
    wire n23413;
    wire n23416;
    wire n23419;
    wire n23422;
    wire n23425;
    wire n23428;
    wire n23431;
    wire n23434;
    wire n23437;
    wire n23440;
    wire n23443;
    wire n23446;
    wire n23449;
    wire n23452;
    wire n23455;
    wire n23461;
    wire n23464;
    wire n23467;
    wire n23470;
    wire n23473;
    wire n23476;
    wire n23479;
    wire n23482;
    wire n23485;
    wire n23488;
    wire n23491;
    wire n23494;
    wire n23497;
    wire n23500;
    wire n23503;
    wire n23506;
    wire n23509;
    wire n23512;
    wire n23515;
    wire n23518;
    wire n23521;
    wire n23524;
    wire n23527;
    wire n23530;
    wire n23533;
    wire n23536;
    wire n23539;
    wire n23542;
    wire n23545;
    wire n23548;
    wire n23551;
    wire n23554;
    wire n23557;
    wire n23560;
    wire n23563;
    wire n23569;
    wire n23572;
    wire n23575;
    wire n23578;
    wire n23581;
    wire n23584;
    wire n23587;
    wire n23590;
    wire n23593;
    wire n23596;
    wire n23599;
    wire n23602;
    wire n23605;
    wire n23608;
    wire n23611;
    wire n23614;
    wire n23617;
    wire n23620;
    wire n23623;
    wire n23626;
    wire n23629;
    wire n23632;
    wire n23635;
    wire n23638;
    wire n23641;
    wire n23644;
    wire n23647;
    wire n23650;
    wire n23653;
    wire n23656;
    wire n23659;
    wire n23662;
    wire n23665;
    wire n23668;
    wire n23671;
    wire n23677;
    wire n23680;
    wire n23683;
    wire n23686;
    wire n23689;
    wire n23692;
    wire n23695;
    wire n23698;
    wire n23701;
    wire n23704;
    wire n23707;
    wire n23710;
    wire n23713;
    wire n23716;
    wire n23719;
    wire n23722;
    wire n23725;
    wire n23728;
    wire n23731;
    wire n23734;
    wire n23737;
    wire n23740;
    wire n23743;
    wire n23746;
    wire n23749;
    wire n23752;
    wire n23755;
    wire n23758;
    wire n23761;
    wire n23764;
    wire n23767;
    wire n23770;
    wire n23773;
    wire n23776;
    wire n23779;
    wire n23782;
    wire n23785;
    wire n23791;
    wire n23794;
    wire n23797;
    wire n23800;
    wire n23803;
    wire n23806;
    wire n23809;
    wire n23812;
    wire n23815;
    wire n23818;
    wire n23821;
    wire n23824;
    wire n23827;
    wire n23830;
    wire n23833;
    wire n23836;
    wire n23839;
    wire n23842;
    wire n23845;
    wire n23848;
    wire n23851;
    wire n23854;
    wire n23857;
    wire n23860;
    wire n23863;
    wire n23866;
    wire n23869;
    wire n23872;
    wire n23875;
    wire n23878;
    wire n23881;
    wire n23884;
    wire n23887;
    wire n23890;
    wire n23893;
    wire n23896;
    wire n23899;
    wire n23905;
    wire n23908;
    wire n23911;
    wire n23914;
    wire n23917;
    wire n23920;
    wire n23923;
    wire n23926;
    wire n23929;
    wire n23932;
    wire n23935;
    wire n23938;
    wire n23941;
    wire n23944;
    wire n23947;
    wire n23950;
    wire n23953;
    wire n23956;
    wire n23959;
    wire n23962;
    wire n23965;
    wire n23968;
    wire n23971;
    wire n23974;
    wire n23977;
    wire n23980;
    wire n23983;
    wire n23986;
    wire n23989;
    wire n23992;
    wire n23995;
    wire n23998;
    wire n24001;
    wire n24004;
    wire n24007;
    wire n24010;
    wire n24016;
    wire n24019;
    wire n24022;
    wire n24025;
    wire n24028;
    wire n24031;
    wire n24034;
    wire n24037;
    wire n24040;
    wire n24043;
    wire n24046;
    wire n24049;
    wire n24052;
    wire n24055;
    wire n24058;
    wire n24061;
    wire n24064;
    wire n24067;
    wire n24070;
    wire n24073;
    wire n24076;
    wire n24079;
    wire n24082;
    wire n24085;
    wire n24088;
    wire n24091;
    wire n24094;
    wire n24097;
    wire n24100;
    wire n24103;
    wire n24106;
    wire n24109;
    wire n24112;
    wire n24115;
    wire n24118;
    wire n24121;
    wire n24124;
    wire n24130;
    wire n24133;
    wire n24136;
    wire n24139;
    wire n24142;
    wire n24145;
    wire n24148;
    wire n24151;
    wire n24154;
    wire n24157;
    wire n24160;
    wire n24163;
    wire n24166;
    wire n24169;
    wire n24172;
    wire n24175;
    wire n24178;
    wire n24181;
    wire n24184;
    wire n24187;
    wire n24190;
    wire n24193;
    wire n24196;
    wire n24199;
    wire n24202;
    wire n24205;
    wire n24208;
    wire n24211;
    wire n24214;
    wire n24217;
    wire n24220;
    wire n24223;
    wire n24226;
    wire n24229;
    wire n24232;
    wire n24235;
    wire n24241;
    wire n24244;
    wire n24247;
    wire n24250;
    wire n24253;
    wire n24256;
    wire n24259;
    wire n24262;
    wire n24265;
    wire n24268;
    wire n24271;
    wire n24274;
    wire n24277;
    wire n24280;
    wire n24283;
    wire n24286;
    wire n24289;
    wire n24292;
    wire n24295;
    wire n24298;
    wire n24301;
    wire n24304;
    wire n24307;
    wire n24310;
    wire n24313;
    wire n24316;
    wire n24319;
    wire n24322;
    wire n24325;
    wire n24328;
    wire n24331;
    wire n24334;
    wire n24337;
    wire n24340;
    wire n24343;
    wire n24349;
    wire n24352;
    wire n24355;
    wire n24358;
    wire n24361;
    wire n24364;
    wire n24367;
    wire n24370;
    wire n24373;
    wire n24376;
    wire n24379;
    wire n24382;
    wire n24385;
    wire n24388;
    wire n24391;
    wire n24394;
    wire n24397;
    wire n24400;
    wire n24403;
    wire n24406;
    wire n24409;
    wire n24412;
    wire n24415;
    wire n24418;
    wire n24421;
    wire n24424;
    wire n24427;
    wire n24430;
    wire n24433;
    wire n24436;
    wire n24439;
    wire n24442;
    wire n24445;
    wire n24448;
    wire n24451;
    wire n24454;
    wire n24457;
    wire n24463;
    wire n24466;
    wire n24469;
    wire n24472;
    wire n24475;
    wire n24478;
    wire n24481;
    wire n24484;
    wire n24487;
    wire n24490;
    wire n24493;
    wire n24496;
    wire n24499;
    wire n24502;
    wire n24505;
    wire n24508;
    wire n24511;
    wire n24514;
    wire n24517;
    wire n24520;
    wire n24523;
    wire n24526;
    wire n24529;
    wire n24532;
    wire n24535;
    wire n24538;
    wire n24541;
    wire n24544;
    wire n24547;
    wire n24550;
    wire n24553;
    wire n24556;
    wire n24559;
    wire n24562;
    wire n24565;
    wire n24571;
    wire n24574;
    wire n24577;
    wire n24580;
    wire n24583;
    wire n24586;
    wire n24589;
    wire n24592;
    wire n24595;
    wire n24598;
    wire n24601;
    wire n24604;
    wire n24607;
    wire n24610;
    wire n24613;
    wire n24616;
    wire n24619;
    wire n24622;
    wire n24625;
    wire n24628;
    wire n24631;
    wire n24634;
    wire n24637;
    wire n24640;
    wire n24643;
    wire n24646;
    wire n24649;
    wire n24652;
    wire n24655;
    wire n24658;
    wire n24661;
    wire n24664;
    wire n24667;
    wire n24670;
    wire n24673;
    wire n24676;
    wire n24679;
    wire n24685;
    wire n24688;
    wire n24691;
    wire n24694;
    wire n24697;
    wire n24700;
    wire n24703;
    wire n24706;
    wire n24709;
    wire n24712;
    wire n24715;
    wire n24718;
    wire n24721;
    wire n24724;
    wire n24727;
    wire n24730;
    wire n24733;
    wire n24736;
    wire n24739;
    wire n24742;
    wire n24745;
    wire n24748;
    wire n24751;
    wire n24754;
    wire n24757;
    wire n24760;
    wire n24763;
    wire n24766;
    wire n24769;
    wire n24772;
    wire n24775;
    wire n24778;
    wire n24781;
    wire n24784;
    wire n24787;
    wire n24790;
    wire n24793;
    wire n24799;
    wire n24802;
    wire n24805;
    wire n24808;
    wire n24811;
    wire n24814;
    wire n24817;
    wire n24820;
    wire n24823;
    wire n24826;
    wire n24829;
    wire n24832;
    wire n24835;
    wire n24838;
    wire n24841;
    wire n24844;
    wire n24847;
    wire n24850;
    wire n24853;
    wire n24856;
    wire n24859;
    wire n24862;
    wire n24865;
    wire n24868;
    wire n24871;
    wire n24874;
    wire n24877;
    wire n24880;
    wire n24883;
    wire n24886;
    wire n24889;
    wire n24892;
    wire n24898;
    wire n24901;
    wire n24904;
    wire n24907;
    wire n24910;
    wire n24913;
    wire n24916;
    wire n24919;
    wire n24922;
    wire n24925;
    wire n24931;
    wire n24934;
    wire n24937;
    wire n24940;
    wire n24943;
    wire n24946;
    wire n24949;
    wire n24952;
    wire n24955;
    wire n24958;
    wire n24964;
    wire n24967;
    wire n24970;
    wire n24973;
    wire n24976;
    wire n24979;
    wire n24982;
    wire n24985;
    wire n24988;
    wire n24991;
    wire n24994;
    wire n24997;
    wire n25000;
    wire n25003;
    wire n25006;
    wire n25009;
    wire n25012;
    wire n25015;
    wire n25018;
    wire n25021;
    wire n25024;
    wire n25027;
    wire n25030;
    wire n25033;
    wire n25039;
    wire n25042;
    wire n25045;
    wire n25048;
    wire n25051;
    wire n25054;
    wire n25057;
    wire n25060;
    wire n25063;
    wire n25066;
    wire n25069;
    wire n25072;
    wire n25075;
    wire n25078;
    wire n25081;
    wire n25084;
    wire n25087;
    wire n25090;
    wire n25093;
    wire n25096;
    wire n25099;
    wire n25102;
    wire n25105;
    wire n25108;
    wire n25111;
    wire n25114;
    wire n25120;
    wire n25123;
    wire n25126;
    wire n25129;
    wire n25132;
    wire n25135;
    wire n25138;
    wire n25141;
    wire n25144;
    wire n25147;
    wire n25150;
    wire n25153;
    wire n25156;
    wire n25159;
    wire n25162;
    wire n25165;
    wire n25168;
    wire n25171;
    wire n25174;
    wire n25177;
    wire n25180;
    wire n25183;
    wire n25186;
    wire n25189;
    wire n25192;
    wire n25195;
    wire n25198;
    wire n25201;
    wire n25204;
    wire n25210;
    wire n25213;
    wire n25216;
    wire n25219;
    wire n25222;
    wire n25225;
    wire n25228;
    wire n25231;
    wire n25234;
    wire n25237;
    wire n25240;
    wire n25243;
    wire n25246;
    wire n25249;
    wire n25252;
    wire n25255;
    wire n25258;
    wire n25261;
    wire n25264;
    wire n25267;
    wire n25270;
    wire n25273;
    wire n25276;
    wire n25279;
    wire n25282;
    wire n25285;
    wire n25288;
    wire n25291;
    wire n25294;
    wire n25297;
    wire n25303;
    wire n25306;
    wire n25309;
    wire n25312;
    wire n25315;
    wire n25318;
    wire n25321;
    wire n25324;
    wire n25327;
    wire n25330;
    wire n25333;
    wire n25336;
    wire n25339;
    wire n25342;
    wire n25345;
    wire n25348;
    wire n25351;
    wire n25354;
    wire n25357;
    wire n25363;
    wire n25366;
    wire n25369;
    wire n25372;
    wire n25375;
    wire n25378;
    wire n25381;
    wire n25384;
    wire n25387;
    wire n25390;
    wire n25393;
    wire n25396;
    wire n25399;
    wire n25402;
    wire n25405;
    wire n25408;
    wire n25411;
    wire n25414;
    wire n25417;
    wire n25420;
    wire n25423;
    wire n25429;
    wire n25432;
    wire n25435;
    wire n25438;
    wire n25441;
    wire n25444;
    wire n25447;
    wire n25450;
    wire n25453;
    wire n25456;
    wire n25459;
    wire n25462;
    wire n25465;
    wire n25468;
    wire n25471;
    wire n25474;
    wire n25477;
    wire n25480;
    wire n25483;
    wire n25486;
    wire n25489;
    wire n25495;
    wire n25498;
    wire n25501;
    wire n25504;
    wire n25507;
    wire n25510;
    wire n25513;
    wire n25516;
    wire n25519;
    wire n25522;
    wire n25525;
    wire n25528;
    wire n25531;
    wire n25534;
    wire n25537;
    wire n25540;
    wire n25543;
    wire n25546;
    wire n25549;
    wire n25552;
    wire n25555;
    wire n25558;
    wire n25561;
    wire n25567;
    wire n25570;
    wire n25573;
    wire n25576;
    wire n25579;
    wire n25582;
    wire n25585;
    wire n25588;
    wire n25591;
    wire n25594;
    wire n25597;
    wire n25600;
    wire n25603;
    wire n25606;
    wire n25609;
    wire n25612;
    wire n25615;
    wire n25618;
    wire n25621;
    wire n25624;
    wire n25627;
    wire n25630;
    wire n25633;
    wire n25636;
    wire n25639;
    wire n25642;
    wire n25645;
    wire n25651;
    wire n25654;
    wire n25657;
    wire n25660;
    wire n25663;
    wire n25666;
    wire n25669;
    wire n25672;
    wire n25675;
    wire n25678;
    wire n25681;
    wire n25684;
    wire n25687;
    wire n25690;
    wire n25693;
    wire n25696;
    wire n25699;
    wire n25702;
    wire n25705;
    wire n25708;
    wire n25711;
    wire n25714;
    wire n25717;
    wire n25720;
    wire n25723;
    wire n25726;
    wire n25729;
    wire n25732;
    wire n25735;
    wire n25741;
    wire n25744;
    wire n25747;
    wire n25750;
    wire n25753;
    wire n25756;
    wire n25759;
    wire n25762;
    wire n25765;
    wire n25768;
    wire n25771;
    wire n25774;
    wire n25777;
    wire n25780;
    wire n25783;
    wire n25786;
    wire n25789;
    wire n25792;
    wire n25795;
    wire n25798;
    wire n25801;
    wire n25804;
    wire n25807;
    wire n25810;
    wire n25813;
    wire n25816;
    wire n25819;
    wire n25822;
    wire n25828;
    wire n25831;
    wire n25834;
    wire n25837;
    wire n25840;
    wire n25843;
    wire n25846;
    wire n25849;
    wire n25852;
    wire n25855;
    wire n25861;
    wire n25864;
    wire n25867;
    wire n25870;
    wire n25873;
    wire n25876;
    wire n25879;
    wire n25882;
    wire n25885;
    wire n25888;
    wire n25894;
    wire n25897;
    wire n25900;
    wire n25906;
    wire n25909;
    wire n25912;
    wire n25915;
    wire n25918;
    wire n25921;
    wire n25924;
    wire n25927;
    wire n25930;
    wire n25933;
    wire n25936;
    wire n25939;
    wire n25942;
    wire n25945;
    wire n25948;
    wire n25951;
    wire n25954;
    wire n25957;
    wire n25960;
    wire n25963;
    wire n25969;
    wire n25972;
    wire n25975;
    wire n25978;
    wire n25981;
    wire n25987;
    wire n25990;
    wire n25993;
    wire n25996;
    wire n26002;
    wire n26005;
    wire n26008;
    wire n26011;
    wire n26014;
    wire n26017;
    wire n26020;
    wire n26023;
    wire n26029;
    wire n26032;
    wire n26035;
    wire n26038;
    wire n26041;
    wire n26044;
    wire n26047;
    wire n26050;
    wire n26056;
    wire n26062;
    wire n26068;
    wire n26074;
    wire n26077;
    wire n26080;
    wire n26083;
    wire n26086;
    wire n26089;
    wire n26092;
    wire n26095;
    wire n26098;
    wire n26101;
    wire n26104;
    wire n26107;
    wire n26110;
    wire n26113;
    wire n26116;
    wire n26119;
    wire n26122;
    wire n26125;
    wire n26128;
    wire n26131;
    wire n26134;
    wire n26137;
    wire n26140;
    wire n26143;
    wire n26149;
    wire n26152;
    wire n26155;
    wire n26158;
    wire n26161;
    wire n26167;
    wire n26170;
    wire n26173;
    wire n26176;
    wire n26179;
    wire n26185;
    wire n26188;
    wire n26191;
    wire n26194;
    wire n26197;
    wire n26203;
    wire n26206;
    wire n26209;
    wire n26212;
    wire n26215;
    wire n26218;
    wire n26221;
    wire n26227;
    wire n26230;
    wire n26233;
    wire n26236;
    wire n26239;
    wire n26242;
    wire n26245;
    wire n26248;
    wire n26251;
    wire n26254;
    wire n26257;
    wire n26260;
    wire n26263;
    wire n26266;
    wire n26269;
    wire n26272;
    wire n26275;
    wire n26278;
    wire n26281;
    wire n26287;
    wire n26293;
    wire n26299;
    wire n26302;
    wire n26305;
    wire n26308;
    wire n26311;
    wire n26314;
    wire n26317;
    wire n26320;
    wire n26323;
    wire n26326;
    wire n26329;
    wire n26332;
    wire n26335;
    wire n26338;
    wire n26341;
    wire n26344;
    wire n26347;
    wire n26353;
    wire n26356;
    wire n26359;
    wire n26362;
    wire n26365;
    wire n26368;
    wire n26371;
    wire n26374;
    wire n26377;
    wire n26380;
    wire n26383;
    wire n26386;
    wire n26389;
    wire n26392;
    wire n26395;
    wire n26398;
    wire n26401;
    wire n26407;
    wire n26410;
    wire n26413;
    wire n26416;
    wire n26419;
    wire n26422;
    wire n26425;
    wire n26428;
    wire n26431;
    wire n26434;
    wire n26437;
    wire n26440;
    wire n26443;
    wire n26446;
    wire n26449;
    wire n26452;
    wire n26455;
    wire n26461;
    wire n26464;
    wire n26467;
    wire n26470;
    wire n26473;
    wire n26476;
    wire n26479;
    wire n26482;
    wire n26485;
    wire n26488;
    wire n26491;
    wire n26494;
    wire n26497;
    wire n26500;
    wire n26503;
    wire n26506;
    wire n26509;
    wire n26515;
    wire n26518;
    wire n26521;
    wire n26524;
    wire n26527;
    wire n26530;
    wire n26533;
    wire n26536;
    wire n26539;
    wire n26542;
    wire n26545;
    wire n26548;
    wire n26554;
    wire n26557;
    wire n26560;
    wire n26563;
    wire n26566;
    wire n26569;
    wire n26572;
    wire n26575;
    wire n26578;
    wire n26581;
    wire n26584;
    wire n26587;
    wire n26590;
    wire n26596;
    wire n26599;
    wire n26602;
    wire n26605;
    wire n26608;
    wire n26611;
    wire n26614;
    wire n26617;
    wire n26620;
    wire n26623;
    wire n26626;
    wire n26629;
    wire n26632;
    wire n26635;
    wire n26638;
    wire n26644;
    wire n26647;
    wire n26650;
    wire n26653;
    wire n26656;
    wire n26659;
    wire n26662;
    wire n26665;
    wire n26668;
    wire n26671;
    wire n26674;
    wire n26677;
    wire n26680;
    wire n26683;
    wire n26686;
    wire n26689;
    wire n26692;
    wire n26698;
    wire n26701;
    wire n26704;
    wire n26707;
    wire n26710;
    wire n26719;
    wire n26722;
    wire n26725;
    wire n26728;
    wire n26731;
    wire n26734;
    wire n26737;
    wire n26740;
    wire n26743;
    wire n26746;
    wire n26749;
    wire n26752;
    wire n26755;
    wire n26758;
    wire n26761;
    wire n26764;
    wire n26770;
    wire n26773;
    wire n26776;
    wire n26779;
    wire n26782;
    wire n26785;
    wire n26788;
    wire n26791;
    wire n26794;
    wire n26797;
    wire n26800;
    wire n26803;
    wire n26806;
    wire n26809;
    wire n26812;
    wire n26815;
    wire n26818;
    wire n26821;
    wire n26824;
    wire n26827;
    jnot g0000(.din(G15), .dout(n316));
    jor g0001(.dinb(G5), .dina(G57), .dout(n320));
    jnot g0002(.din(G184), .dout(n323));
    jnot g0003(.din(G228), .dout(n326));
    jor g0004(.dinb(n323), .dina(n326), .dout(n330));
    jnot g0005(.din(G150), .dout(n333));
    jnot g0006(.din(G240), .dout(n336));
    jor g0007(.dinb(n333), .dina(n336), .dout(n340));
    jor g0008(.dinb(n330), .dina(n340), .dout(n344));
    jnot g0009(.din(G210), .dout(n347));
    jnot g0010(.din(G218), .dout(n350));
    jor g0011(.dinb(n347), .dina(n350), .dout(n354));
    jnot g0012(.din(G152), .dout(n357));
    jnot g0013(.din(G230), .dout(n360));
    jor g0014(.dinb(n357), .dina(n360), .dout(n364));
    jor g0015(.dinb(n354), .dina(n364), .dout(n368));
    jnot g0016(.din(G183), .dout(n371));
    jnot g0017(.din(G185), .dout(n374));
    jor g0018(.dinb(n371), .dina(n374), .dout(n378));
    jnot g0019(.din(G182), .dout(n381));
    jnot g0020(.din(G186), .dout(n384));
    jor g0021(.dinb(n381), .dina(n384), .dout(n388));
    jor g0022(.dinb(n378), .dina(n388), .dout(n392));
    jnot g0023(.din(G172), .dout(n395));
    jnot g0024(.din(G188), .dout(n398));
    jor g0025(.dinb(n395), .dina(n398), .dout(n402));
    jnot g0026(.din(G162), .dout(n405));
    jnot g0027(.din(G199), .dout(n408));
    jor g0028(.dinb(n405), .dina(n408), .dout(n412));
    jor g0029(.dinb(n402), .dina(n412), .dout(n416));
    jnot g0030(.din(G1197), .dout(n419));
    jor g0031(.dinb(n7855), .dina(n419), .dout(n423));
    jnot g0032(.din(G134), .dout(n426));
    jnot g0033(.din(G133), .dout(n429));
    jor g0034(.dinb(n7861), .dina(n429), .dout(n433));
    jor g0035(.dinb(n7865), .dina(n433), .dout(n437));
    jand g0036(.dinb(G1), .dina(G163), .dout(n441));
    jnot g0037(.din(G41), .dout(n444));
    jor g0038(.dinb(n18544), .dina(n444), .dout(n448));
    jor g0039(.dinb(n18394), .dina(n448), .dout(n452));
    jnot g0040(.din(G18), .dout(n455));
    jand g0041(.dinb(n455), .dina(n18397), .dout(n459));
    jand g0042(.dinb(n448), .dina(n459), .dout(n463));
    jnot g0043(.din(n463), .dout(n466));
    jand g0044(.dinb(n18389), .dina(n466), .dout(n470));
    jxor g0045(.dinb(n17860), .dina(n470), .dout(n474));
    jnot g0046(.din(G38), .dout(n477));
    jand g0047(.dinb(G1492), .dina(G4528), .dout(n481));
    jxor g0048(.dinb(n477), .dina(n481), .dout(n485));
    jand g0049(.dinb(G1496), .dina(G4528), .dout(n489));
    jor g0050(.dinb(n477), .dina(n489), .dout(n493));
    jnot g0051(.din(G1496), .dout(n496));
    jnot g0052(.din(G4528), .dout(n499));
    jor g0053(.dinb(n11032), .dina(n499), .dout(n503));
    jor g0054(.dinb(n11020), .dina(n503), .dout(n507));
    jand g0055(.dinb(n10016), .dina(n507), .dout(n511));
    jnot g0056(.din(G1486), .dout(n514));
    jand g0057(.dinb(G9), .dina(G12), .dout(n518));
    jnot g0058(.din(n518), .dout(n521));
    jor g0059(.dinb(n455), .dina(n12710), .dout(n525));
    jand g0060(.dinb(n521), .dina(n525), .dout(n529));
    jand g0061(.dinb(n12718), .dina(n529), .dout(n533));
    jxor g0062(.dinb(n12712), .dina(n529), .dout(n537));
    jor g0063(.dinb(n455), .dina(n15473), .dout(n541));
    jand g0064(.dinb(n521), .dina(n541), .dout(n545));
    jnot g0065(.din(n545), .dout(n548));
    jand g0066(.dinb(n15487), .dina(n548), .dout(n552));
    jnot g0067(.din(n552), .dout(n555));
    jnot g0068(.din(G1480), .dout(n558));
    jand g0069(.dinb(n15481), .dina(n545), .dout(n562));
    jnot g0070(.din(G106), .dout(n565));
    jor g0071(.dinb(n455), .dina(n15500), .dout(n569));
    jand g0072(.dinb(n521), .dina(n569), .dout(n573));
    jxor g0073(.dinb(n15506), .dina(n573), .dout(n577));
    jnot g0074(.din(G1462), .dout(n580));
    jor g0075(.dinb(n455), .dina(n12656), .dout(n584));
    jand g0076(.dinb(n521), .dina(n584), .dout(n588));
    jand g0077(.dinb(n12658), .dina(n588), .dout(n592));
    jnot g0078(.din(G1469), .dout(n595));
    jor g0079(.dinb(n455), .dina(n12626), .dout(n599));
    jand g0080(.dinb(n521), .dina(n599), .dout(n603));
    jxor g0081(.dinb(n12628), .dina(n603), .dout(n607));
    jand g0082(.dinb(n592), .dina(n607), .dout(n611));
    jand g0083(.dinb(n12673), .dina(n611), .dout(n615));
    jnot g0084(.din(n615), .dout(n618));
    jand g0085(.dinb(n15506), .dina(n573), .dout(n622));
    jnot g0086(.din(n622), .dout(n625));
    jnot g0087(.din(n573), .dout(n628));
    jand g0088(.dinb(n15508), .dina(n628), .dout(n632));
    jand g0089(.dinb(n12628), .dina(n603), .dout(n636));
    jnot g0090(.din(n636), .dout(n639));
    jor g0091(.dinb(n632), .dina(n639), .dout(n643));
    jand g0092(.dinb(n12524), .dina(n643), .dout(n647));
    jand g0093(.dinb(n618), .dina(n647), .dout(n651));
    jnot g0094(.din(n651), .dout(n654));
    jor g0095(.dinb(n12446), .dina(n654), .dout(n658));
    jand g0096(.dinb(n12431), .dina(n658), .dout(n662));
    jand g0097(.dinb(n11212), .dina(n662), .dout(n666));
    jor g0098(.dinb(n11120), .dina(n666), .dout(n670));
    jxor g0099(.dinb(n12658), .dina(n588), .dout(n674));
    jand g0100(.dinb(n607), .dina(n674), .dout(n678));
    jxor g0101(.dinb(n15475), .dina(n545), .dout(n682));
    jand g0102(.dinb(n577), .dina(n682), .dout(n686));
    jand g0103(.dinb(n678), .dina(n686), .dout(n690));
    jand g0104(.dinb(n12676), .dina(n690), .dout(n694));
    jor g0105(.dinb(n670), .dina(n10918), .dout(n698));
    jnot g0106(.din(G2256), .dout(n701));
    jor g0107(.dinb(n455), .dina(n15356), .dout(n705));
    jand g0108(.dinb(n521), .dina(n705), .dout(n709));
    jand g0109(.dinb(n15364), .dina(n709), .dout(n713));
    jxor g0110(.dinb(n15358), .dina(n709), .dout(n717));
    jnot g0111(.din(G2253), .dout(n720));
    jor g0112(.dinb(n455), .dina(n15068), .dout(n724));
    jand g0113(.dinb(n521), .dina(n724), .dout(n728));
    jxor g0114(.dinb(n15076), .dina(n728), .dout(n732));
    jnot g0115(.din(G2247), .dout(n735));
    jor g0116(.dinb(n455), .dina(n14966), .dout(n739));
    jand g0117(.dinb(n521), .dina(n739), .dout(n743));
    jxor g0118(.dinb(n14972), .dina(n743), .dout(n747));
    jnot g0119(.din(G2239), .dout(n750));
    jor g0120(.dinb(n455), .dina(n14843), .dout(n754));
    jand g0121(.dinb(n521), .dina(n754), .dout(n758));
    jxor g0122(.dinb(n14849), .dina(n758), .dout(n762));
    jand g0123(.dinb(n747), .dina(n762), .dout(n766));
    jand g0124(.dinb(n15058), .dina(n766), .dout(n770));
    jnot g0125(.din(n728), .dout(n773));
    jand g0126(.dinb(n15082), .dina(n773), .dout(n777));
    jnot g0127(.din(n777), .dout(n780));
    jand g0128(.dinb(n15070), .dina(n728), .dout(n784));
    jand g0129(.dinb(n14972), .dina(n743), .dout(n788));
    jand g0130(.dinb(n14849), .dina(n758), .dout(n792));
    jand g0131(.dinb(n747), .dina(n792), .dout(n796));
    jor g0132(.dinb(n14680), .dina(n796), .dout(n800));
    jor g0133(.dinb(n14519), .dina(n800), .dout(n804));
    jand g0134(.dinb(n14513), .dina(n804), .dout(n808));
    jor g0135(.dinb(n14444), .dina(n808), .dout(n812));
    jnot g0136(.din(G2236), .dout(n815));
    jor g0137(.dinb(n455), .dina(n14366), .dout(n819));
    jand g0138(.dinb(n521), .dina(n819), .dout(n823));
    jand g0139(.dinb(n14372), .dina(n823), .dout(n827));
    jor g0140(.dinb(n14372), .dina(n823), .dout(n831));
    jnot g0141(.din(G2230), .dout(n834));
    jand g0142(.dinb(n455), .dina(n14336), .dout(n838));
    jand g0143(.dinb(G18), .dina(G158), .dout(n842));
    jor g0144(.dinb(n838), .dina(n14333), .dout(n846));
    jand g0145(.dinb(n14344), .dina(n846), .dout(n850));
    jand g0146(.dinb(n831), .dina(n850), .dout(n854));
    jor g0147(.dinb(n14126), .dina(n854), .dout(n858));
    jxor g0148(.dinb(n14372), .dina(n823), .dout(n862));
    jxor g0149(.dinb(n14338), .dina(n846), .dout(n866));
    jand g0150(.dinb(n862), .dina(n866), .dout(n870));
    jnot g0151(.din(G2224), .dout(n873));
    jand g0152(.dinb(n455), .dina(n13829), .dout(n877));
    jand g0153(.dinb(G18), .dina(G159), .dout(n881));
    jor g0154(.dinb(n877), .dina(n13826), .dout(n885));
    jxor g0155(.dinb(n13835), .dina(n885), .dout(n889));
    jnot g0156(.din(G2218), .dout(n892));
    jand g0157(.dinb(n455), .dina(n13718), .dout(n896));
    jand g0158(.dinb(G18), .dina(G160), .dout(n900));
    jor g0159(.dinb(n896), .dina(n13715), .dout(n904));
    jxor g0160(.dinb(n13726), .dina(n904), .dout(n908));
    jnot g0161(.din(G2211), .dout(n911));
    jand g0162(.dinb(n455), .dina(n13613), .dout(n915));
    jand g0163(.dinb(G18), .dina(G151), .dout(n919));
    jor g0164(.dinb(n915), .dina(n13610), .dout(n923));
    jxor g0165(.dinb(n13621), .dina(n923), .dout(n927));
    jand g0166(.dinb(n908), .dina(n927), .dout(n931));
    jand g0167(.dinb(n13819), .dina(n931), .dout(n935));
    jnot g0168(.din(n885), .dout(n938));
    jand g0169(.dinb(n13837), .dina(n938), .dout(n942));
    jnot g0170(.din(n904), .dout(n945));
    jand g0171(.dinb(n13732), .dina(n945), .dout(n949));
    jand g0172(.dinb(n13615), .dina(n923), .dout(n953));
    jnot g0173(.din(n953), .dout(n956));
    jor g0174(.dinb(n949), .dina(n956), .dout(n960));
    jand g0175(.dinb(n13835), .dina(n885), .dout(n964));
    jand g0176(.dinb(n13720), .dina(n904), .dout(n968));
    jor g0177(.dinb(n964), .dina(n968), .dout(n972));
    jnot g0178(.din(n972), .dout(n975));
    jand g0179(.dinb(n960), .dina(n975), .dout(n979));
    jor g0180(.dinb(n13385), .dina(n979), .dout(n983));
    jnot g0181(.din(n983), .dout(n986));
    jor g0182(.dinb(n13322), .dina(n986), .dout(n990));
    jand g0183(.dinb(n13849), .dina(n990), .dout(n994));
    jor g0184(.dinb(n14110), .dina(n994), .dout(n998));
    jand g0185(.dinb(n13862), .dina(n986), .dout(n1002));
    jnot g0186(.din(G4437), .dout(n1005));
    jand g0187(.dinb(G18), .dina(G219), .dout(n1009));
    jand g0188(.dinb(n455), .dina(n16001), .dout(n1013));
    jor g0189(.dinb(n15998), .dina(n1013), .dout(n1017));
    jand g0190(.dinb(n16009), .dina(n1017), .dout(n1021));
    jnot g0191(.din(n1017), .dout(n1024));
    jand g0192(.dinb(n16015), .dina(n1024), .dout(n1028));
    jnot g0193(.din(n1028), .dout(n1031));
    jnot g0194(.din(G4432), .dout(n1034));
    jand g0195(.dinb(G18), .dina(G220), .dout(n1038));
    jand g0196(.dinb(n455), .dina(n16349), .dout(n1042));
    jor g0197(.dinb(n16346), .dina(n1042), .dout(n1046));
    jxor g0198(.dinb(n16357), .dina(n1046), .dout(n1050));
    jnot g0199(.din(G4420), .dout(n1053));
    jand g0200(.dinb(G18), .dina(G222), .dout(n1057));
    jand g0201(.dinb(n455), .dina(n16292), .dout(n1061));
    jor g0202(.dinb(n16289), .dina(n1061), .dout(n1065));
    jand g0203(.dinb(n16298), .dina(n1065), .dout(n1069));
    jnot g0204(.din(n1069), .dout(n1072));
    jnot g0205(.din(G4427), .dout(n1075));
    jand g0206(.dinb(G18), .dina(G221), .dout(n1079));
    jand g0207(.dinb(n455), .dina(n16316), .dout(n1083));
    jor g0208(.dinb(n16313), .dina(n1083), .dout(n1087));
    jxor g0209(.dinb(n16322), .dina(n1087), .dout(n1091));
    jnot g0210(.din(n1065), .dout(n1094));
    jand g0211(.dinb(n16300), .dina(n1094), .dout(n1098));
    jnot g0212(.din(n1098), .dout(n1101));
    jnot g0213(.din(G4415), .dout(n1104));
    jand g0214(.dinb(G18), .dina(G223), .dout(n1108));
    jand g0215(.dinb(n455), .dina(n17168), .dout(n1112));
    jor g0216(.dinb(n17165), .dina(n1112), .dout(n1116));
    jand g0217(.dinb(n17174), .dina(n1116), .dout(n1120));
    jnot g0218(.din(n1116), .dout(n1123));
    jand g0219(.dinb(n17176), .dina(n1123), .dout(n1127));
    jnot g0220(.din(n1127), .dout(n1130));
    jnot g0221(.din(G4410), .dout(n1133));
    jand g0222(.dinb(G18), .dina(G224), .dout(n1137));
    jand g0223(.dinb(n455), .dina(n16856), .dout(n1141));
    jor g0224(.dinb(n16853), .dina(n1141), .dout(n1145));
    jand g0225(.dinb(n16864), .dina(n1145), .dout(n1149));
    jnot g0226(.din(n1145), .dout(n1152));
    jand g0227(.dinb(n16870), .dina(n1152), .dout(n1156));
    jnot g0228(.din(n1156), .dout(n1159));
    jnot g0229(.din(G4405), .dout(n1162));
    jand g0230(.dinb(G18), .dina(G225), .dout(n1166));
    jand g0231(.dinb(n455), .dina(n16832), .dout(n1170));
    jor g0232(.dinb(n16829), .dina(n1170), .dout(n1174));
    jand g0233(.dinb(n16838), .dina(n1174), .dout(n1178));
    jnot g0234(.din(n1174), .dout(n1181));
    jand g0235(.dinb(n16840), .dina(n1181), .dout(n1185));
    jnot g0236(.din(n1185), .dout(n1188));
    jnot g0237(.din(G4400), .dout(n1191));
    jand g0238(.dinb(G18), .dina(G226), .dout(n1195));
    jand g0239(.dinb(n455), .dina(n17081), .dout(n1199));
    jor g0240(.dinb(n17078), .dina(n1199), .dout(n1203));
    jand g0241(.dinb(n17087), .dina(n1203), .dout(n1207));
    jnot g0242(.din(n1203), .dout(n1210));
    jand g0243(.dinb(n17089), .dina(n1210), .dout(n1214));
    jnot g0244(.din(n1214), .dout(n1217));
    jnot g0245(.din(G4394), .dout(n1220));
    jand g0246(.dinb(G18), .dina(G217), .dout(n1224));
    jand g0247(.dinb(n455), .dina(n17009), .dout(n1228));
    jor g0248(.dinb(n17006), .dina(n1228), .dout(n1232));
    jand g0249(.dinb(n17015), .dina(n1232), .dout(n1236));
    jand g0250(.dinb(n1217), .dina(n16585), .dout(n1240));
    jor g0251(.dinb(n16597), .dina(n1240), .dout(n1244));
    jand g0252(.dinb(n16505), .dina(n1244), .dout(n1248));
    jor g0253(.dinb(n16621), .dina(n1248), .dout(n1252));
    jand g0254(.dinb(n16499), .dina(n1252), .dout(n1256));
    jor g0255(.dinb(n16487), .dina(n1256), .dout(n1260));
    jand g0256(.dinb(n16445), .dina(n1260), .dout(n1264));
    jor g0257(.dinb(n16427), .dina(n1264), .dout(n1268));
    jxor g0258(.dinb(n17174), .dina(n1116), .dout(n1272));
    jxor g0259(.dinb(n17087), .dina(n1203), .dout(n1276));
    jxor g0260(.dinb(n17015), .dina(n1232), .dout(n1280));
    jand g0261(.dinb(n1276), .dina(n1280), .dout(n1284));
    jxor g0262(.dinb(n16858), .dina(n1145), .dout(n1288));
    jxor g0263(.dinb(n16838), .dina(n1174), .dout(n1292));
    jand g0264(.dinb(n1288), .dina(n1292), .dout(n1296));
    jand g0265(.dinb(n1284), .dina(n1296), .dout(n1300));
    jand g0266(.dinb(n17162), .dina(n1300), .dout(n1304));
    jnot g0267(.din(G3749), .dout(n1307));
    jand g0268(.dinb(G18), .dina(G231), .dout(n1311));
    jand g0269(.dinb(n455), .dina(n18053), .dout(n1315));
    jor g0270(.dinb(n18050), .dina(n1315), .dout(n1319));
    jand g0271(.dinb(n18061), .dina(n1319), .dout(n1323));
    jnot g0272(.din(n1319), .dout(n1326));
    jand g0273(.dinb(n18067), .dina(n1326), .dout(n1330));
    jnot g0274(.din(n1330), .dout(n1333));
    jnot g0275(.din(G3743), .dout(n1336));
    jand g0276(.dinb(G18), .dina(G232), .dout(n1340));
    jand g0277(.dinb(n455), .dina(n17996), .dout(n1344));
    jor g0278(.dinb(n17993), .dina(n1344), .dout(n1348));
    jxor g0279(.dinb(n17941), .dina(n1348), .dout(n1352));
    jnot g0280(.din(G3737), .dout(n1355));
    jand g0281(.dinb(G18), .dina(G233), .dout(n1359));
    jand g0282(.dinb(n455), .dina(n18161), .dout(n1363));
    jor g0283(.dinb(n18158), .dina(n1363), .dout(n1367));
    jxor g0284(.dinb(n18169), .dina(n1367), .dout(n1371));
    jnot g0285(.din(G3729), .dout(n1374));
    jand g0286(.dinb(G18), .dina(G234), .dout(n1378));
    jand g0287(.dinb(n455), .dina(n18110), .dout(n1382));
    jor g0288(.dinb(n18107), .dina(n1382), .dout(n1386));
    jxor g0289(.dinb(n17978), .dina(n1386), .dout(n1390));
    jand g0290(.dinb(n1371), .dina(n1390), .dout(n1394));
    jand g0291(.dinb(n17686), .dina(n1394), .dout(n1398));
    jnot g0292(.din(n1398), .dout(n1401));
    jnot g0293(.din(n1348), .dout(n1404));
    jand g0294(.dinb(n17998), .dina(n1404), .dout(n1408));
    jand g0295(.dinb(n17935), .dina(n1348), .dout(n1412));
    jnot g0296(.din(n1412), .dout(n1415));
    jand g0297(.dinb(n18163), .dina(n1367), .dout(n1419));
    jand g0298(.dinb(n17978), .dina(n1386), .dout(n1423));
    jand g0299(.dinb(n1371), .dina(n1423), .dout(n1427));
    jor g0300(.dinb(n17980), .dina(n1427), .dout(n1431));
    jnot g0301(.din(n1431), .dout(n1434));
    jand g0302(.dinb(n17585), .dina(n1434), .dout(n1438));
    jor g0303(.dinb(n17983), .dina(n1438), .dout(n1442));
    jand g0304(.dinb(n17564), .dina(n1442), .dout(n1446));
    jnot g0305(.din(n1446), .dout(n1449));
    jnot g0306(.din(n1442), .dout(n1452));
    jnot g0307(.din(G3723), .dout(n1455));
    jand g0308(.dinb(G18), .dina(G235), .dout(n1459));
    jand g0309(.dinb(n455), .dina(n18542), .dout(n1463));
    jor g0310(.dinb(n18539), .dina(n1463), .dout(n1467));
    jxor g0311(.dinb(n18553), .dina(n1467), .dout(n1471));
    jnot g0312(.din(G3717), .dout(n1474));
    jand g0313(.dinb(G18), .dina(G236), .dout(n1478));
    jand g0314(.dinb(n455), .dina(n18473), .dout(n1482));
    jor g0315(.dinb(n18470), .dina(n1482), .dout(n1486));
    jxor g0316(.dinb(n18481), .dina(n1486), .dout(n1490));
    jnot g0317(.din(G3711), .dout(n1493));
    jand g0318(.dinb(G18), .dina(G237), .dout(n1497));
    jand g0319(.dinb(n455), .dina(n18422), .dout(n1501));
    jor g0320(.dinb(n18419), .dina(n1501), .dout(n1505));
    jxor g0321(.dinb(n18427), .dina(n1505), .dout(n1509));
    jnot g0322(.din(G238), .dout(n1512));
    jor g0323(.dinb(n455), .dina(n1512), .dout(n1516));
    jnot g0324(.din(G29), .dout(n1519));
    jor g0325(.dinb(n18424), .dina(n1519), .dout(n1523));
    jand g0326(.dinb(n1516), .dina(n1523), .dout(n1527));
    jxor g0327(.dinb(n18361), .dina(n1527), .dout(n1531));
    jand g0328(.dinb(n470), .dina(n18347), .dout(n1535));
    jand g0329(.dinb(n18412), .dina(n1535), .dout(n1539));
    jand g0330(.dinb(n18460), .dina(n1539), .dout(n1543));
    jand g0331(.dinb(n18514), .dina(n1543), .dout(n1547));
    jand g0332(.dinb(n18547), .dina(n1467), .dout(n1551));
    jnot g0333(.din(n1467), .dout(n1554));
    jand g0334(.dinb(n18559), .dina(n1554), .dout(n1558));
    jnot g0335(.din(n1558), .dout(n1561));
    jnot g0336(.din(n1486), .dout(n1564));
    jand g0337(.dinb(n18487), .dina(n1564), .dout(n1568));
    jnot g0338(.din(n1568), .dout(n1571));
    jand g0339(.dinb(n18475), .dina(n1486), .dout(n1575));
    jand g0340(.dinb(n18427), .dina(n1505), .dout(n1579));
    jor g0341(.dinb(n18433), .dina(n1505), .dout(n1583));
    jnot g0342(.din(G3705), .dout(n1586));
    jand g0343(.dinb(G18), .dina(G238), .dout(n1590));
    jand g0344(.dinb(n455), .dina(n18349), .dout(n1594));
    jor g0345(.dinb(n17729), .dina(n1594), .dout(n1598));
    jor g0346(.dinb(n17737), .dina(n1598), .dout(n1602));
    jnot g0347(.din(G3701), .dout(n1605));
    jand g0348(.dinb(n455), .dina(n18391), .dout(n1609));
    jand g0349(.dinb(n17713), .dina(n1609), .dout(n1613));
    jand g0350(.dinb(n17731), .dina(n1598), .dout(n1617));
    jor g0351(.dinb(n17711), .dina(n1617), .dout(n1621));
    jand g0352(.dinb(n17725), .dina(n1621), .dout(n1625));
    jand g0353(.dinb(n18226), .dina(n1625), .dout(n1629));
    jor g0354(.dinb(n18232), .dina(n1629), .dout(n1633));
    jor g0355(.dinb(n18262), .dina(n1633), .dout(n1637));
    jand g0356(.dinb(n17759), .dina(n1637), .dout(n1641));
    jand g0357(.dinb(n17699), .dina(n1641), .dout(n1645));
    jor g0358(.dinb(n18301), .dina(n1645), .dout(n1649));
    jor g0359(.dinb(n18331), .dina(n1649), .dout(n1653));
    jor g0360(.dinb(n17251), .dina(n1649), .dout(n1657));
    jand g0361(.dinb(n1653), .dina(n1657), .dout(n1661));
    jor g0362(.dinb(n17240), .dina(n1661), .dout(n1665));
    jand g0363(.dinb(n17228), .dina(n1665), .dout(n1669));
    jand g0364(.dinb(n17216), .dina(n1669), .dout(n1673));
    jor g0365(.dinb(n17344), .dina(n1673), .dout(n1677));
    jand g0366(.dinb(n16687), .dina(n1677), .dout(n1681));
    jor g0367(.dinb(n16387), .dina(n1681), .dout(n1685));
    jand g0368(.dinb(n12968), .dina(n1685), .dout(n1689));
    jand g0369(.dinb(n16183), .dina(n1689), .dout(n1693));
    jand g0370(.dinb(n12926), .dina(n1693), .dout(n1697));
    jand g0371(.dinb(n12970), .dina(n1697), .dout(n1701));
    jand g0372(.dinb(n16351), .dina(n1046), .dout(n1705));
    jnot g0373(.din(n1705), .dout(n1708));
    jnot g0374(.din(n1046), .dout(n1711));
    jand g0375(.dinb(n16363), .dina(n1711), .dout(n1715));
    jand g0376(.dinb(n16322), .dina(n1087), .dout(n1719));
    jand g0377(.dinb(n1069), .dina(n1091), .dout(n1723));
    jor g0378(.dinb(n16181), .dina(n1723), .dout(n1727));
    jnot g0379(.din(n1727), .dout(n1730));
    jor g0380(.dinb(n16324), .dina(n1730), .dout(n1734));
    jand g0381(.dinb(n12875), .dina(n1734), .dout(n1738));
    jnot g0382(.din(n1738), .dout(n1741));
    jor g0383(.dinb(n1701), .dina(n12821), .dout(n1745));
    jand g0384(.dinb(n12779), .dina(n1745), .dout(n1749));
    jor g0385(.dinb(n13087), .dina(n1749), .dout(n1753));
    jor g0386(.dinb(n14047), .dina(n1753), .dout(n1757));
    jor g0387(.dinb(n13153), .dina(n1757), .dout(n1761));
    jand g0388(.dinb(n13207), .dina(n1761), .dout(n1765));
    jor g0389(.dinb(n14446), .dina(n1765), .dout(n1769));
    jand g0390(.dinb(n14374), .dina(n1769), .dout(n1773));
    jand g0391(.dinb(n15094), .dina(n1773), .dout(n1777));
    jor g0392(.dinb(n15262), .dina(n1777), .dout(n1781));
    jor g0393(.dinb(n10834), .dina(n1781), .dout(n1785));
    jand g0394(.dinb(n10771), .dina(n1785), .dout(n1789));
    jand g0395(.dinb(n10013), .dina(n1789), .dout(n1793));
    jand g0396(.dinb(n10018), .dina(n1793), .dout(n1797));
    jnot g0397(.din(n481), .dout(n1800));
    jand g0398(.dinb(n11026), .dina(n1800), .dout(n1804));
    jand g0399(.dinb(n11092), .dina(n496), .dout(n1808));
    jor g0400(.dinb(n1804), .dina(n9698), .dout(n1812));
    jor g0401(.dinb(n1797), .dina(n9695), .dout(G246));
    jand g0402(.dinb(G1455), .dina(G2204), .dout(n1820));
    jor g0403(.dinb(n503), .dina(n8447), .dout(n1824));
    jor g0404(.dinb(n455), .dina(n9344), .dout(n1828));
    jand g0405(.dinb(n521), .dina(n1828), .dout(n1832));
    jor g0406(.dinb(n455), .dina(n514), .dout(n1836));
    jor g0407(.dinb(G18), .dina(G88), .dout(n1840));
    jand g0408(.dinb(n1836), .dina(n9467), .dout(n1844));
    jxor g0409(.dinb(n1832), .dina(n1844), .dout(n1848));
    jor g0410(.dinb(n455), .dina(n9335), .dout(n1852));
    jand g0411(.dinb(n521), .dina(n1852), .dout(n1856));
    jor g0412(.dinb(n455), .dina(n558), .dout(n1860));
    jor g0413(.dinb(G18), .dina(G112), .dout(n1864));
    jand g0414(.dinb(n1860), .dina(n9464), .dout(n1868));
    jor g0415(.dinb(n1856), .dina(n1868), .dout(n1872));
    jand g0416(.dinb(n1856), .dina(n1868), .dout(n1876));
    jor g0417(.dinb(n455), .dina(n580), .dout(n1880));
    jor g0418(.dinb(G18), .dina(G113), .dout(n1884));
    jand g0419(.dinb(n1880), .dina(n9455), .dout(n1888));
    jand g0420(.dinb(n9349), .dina(n1888), .dout(n1892));
    jor g0421(.dinb(n455), .dina(n9353), .dout(n1896));
    jand g0422(.dinb(n521), .dina(n1896), .dout(n1900));
    jand g0423(.dinb(G18), .dina(G106), .dout(n1904));
    jnot g0424(.din(n1904), .dout(n1907));
    jor g0425(.dinb(G18), .dina(G87), .dout(n1911));
    jand g0426(.dinb(n1907), .dina(n9461), .dout(n1915));
    jxor g0427(.dinb(n1900), .dina(n1915), .dout(n1919));
    jor g0428(.dinb(n455), .dina(n9347), .dout(n1923));
    jand g0429(.dinb(n521), .dina(n1923), .dout(n1927));
    jor g0430(.dinb(n455), .dina(n595), .dout(n1931));
    jor g0431(.dinb(G18), .dina(G111), .dout(n1935));
    jand g0432(.dinb(n1931), .dina(n9458), .dout(n1939));
    jxor g0433(.dinb(n1927), .dina(n1939), .dout(n1943));
    jand g0434(.dinb(n1919), .dina(n1943), .dout(n1947));
    jand g0435(.dinb(n8360), .dina(n1947), .dout(n1951));
    jor g0436(.dinb(n8357), .dina(n1951), .dout(n1955));
    jand g0437(.dinb(n8351), .dina(n1955), .dout(n1959));
    jand g0438(.dinb(n8362), .dina(n1959), .dout(n1963));
    jor g0439(.dinb(n455), .dina(n9293), .dout(n1967));
    jand g0440(.dinb(n521), .dina(n1967), .dout(n1971));
    jor g0441(.dinb(n455), .dina(n701), .dout(n1975));
    jor g0442(.dinb(G18), .dina(G110), .dout(n1979));
    jand g0443(.dinb(n1975), .dina(n9563), .dout(n1983));
    jxor g0444(.dinb(n1971), .dina(n1983), .dout(n1987));
    jor g0445(.dinb(n455), .dina(n9290), .dout(n1991));
    jand g0446(.dinb(n521), .dina(n1991), .dout(n1995));
    jor g0447(.dinb(n455), .dina(n720), .dout(n1999));
    jor g0448(.dinb(G18), .dina(G109), .dout(n2003));
    jand g0449(.dinb(n1999), .dina(n9560), .dout(n2007));
    jxor g0450(.dinb(n1995), .dina(n2007), .dout(n2011));
    jand g0451(.dinb(n1987), .dina(n2011), .dout(n2015));
    jor g0452(.dinb(n455), .dina(n9299), .dout(n2019));
    jand g0453(.dinb(n521), .dina(n2019), .dout(n2023));
    jand g0454(.dinb(G18), .dina(G2247), .dout(n2027));
    jnot g0455(.din(n2027), .dout(n2030));
    jor g0456(.dinb(G18), .dina(G86), .dout(n2034));
    jand g0457(.dinb(n2030), .dina(n9593), .dout(n2038));
    jand g0458(.dinb(n2023), .dina(n2038), .dout(n2042));
    jor g0459(.dinb(n2023), .dina(n2038), .dout(n2046));
    jor g0460(.dinb(n455), .dina(n9296), .dout(n2050));
    jand g0461(.dinb(n521), .dina(n2050), .dout(n2054));
    jand g0462(.dinb(G18), .dina(G2239), .dout(n2058));
    jnot g0463(.din(n2058), .dout(n2061));
    jor g0464(.dinb(G18), .dina(G63), .dout(n2065));
    jand g0465(.dinb(n2061), .dina(n9590), .dout(n2069));
    jand g0466(.dinb(n2054), .dina(n2069), .dout(n2073));
    jand g0467(.dinb(n2046), .dina(n2073), .dout(n2077));
    jor g0468(.dinb(n8338), .dina(n2077), .dout(n2081));
    jand g0469(.dinb(n8342), .dina(n2081), .dout(n2085));
    jand g0470(.dinb(n1971), .dina(n1983), .dout(n2089));
    jor g0471(.dinb(n1971), .dina(n1983), .dout(n2093));
    jand g0472(.dinb(n1995), .dina(n2007), .dout(n2097));
    jand g0473(.dinb(n2093), .dina(n2097), .dout(n2101));
    jor g0474(.dinb(n8336), .dina(n2101), .dout(n2105));
    jor g0475(.dinb(n2085), .dina(n8333), .dout(n2109));
    jnot g0476(.din(n2042), .dout(n2112));
    jnot g0477(.din(n2073), .dout(n2115));
    jand g0478(.dinb(n2112), .dina(n2115), .dout(n2119));
    jand g0479(.dinb(n8342), .dina(n2119), .dout(n2123));
    jor g0480(.dinb(n455), .dina(n9305), .dout(n2127));
    jand g0481(.dinb(n521), .dina(n2127), .dout(n2131));
    jand g0482(.dinb(G18), .dina(G2236), .dout(n2135));
    jnot g0483(.din(n2135), .dout(n2138));
    jor g0484(.dinb(G18), .dina(G64), .dout(n2142));
    jand g0485(.dinb(n2138), .dina(n9575), .dout(n2146));
    jxor g0486(.dinb(n2131), .dina(n2146), .dout(n2150));
    jand g0487(.dinb(G18), .dina(G178), .dout(n2154));
    jor g0488(.dinb(n838), .dina(n9302), .dout(n2158));
    jor g0489(.dinb(n455), .dina(n834), .dout(n2162));
    jor g0490(.dinb(G18), .dina(G85), .dout(n2166));
    jand g0491(.dinb(n2162), .dina(n9572), .dout(n2170));
    jxor g0492(.dinb(n2158), .dina(n2170), .dout(n2174));
    jand g0493(.dinb(n2150), .dina(n2174), .dout(n2178));
    jand g0494(.dinb(G18), .dina(G179), .dout(n2182));
    jor g0495(.dinb(n877), .dina(n9287), .dout(n2186));
    jand g0496(.dinb(G18), .dina(G2224), .dout(n2190));
    jnot g0497(.din(n2190), .dout(n2193));
    jor g0498(.dinb(G18), .dina(G84), .dout(n2197));
    jand g0499(.dinb(n2193), .dina(n9569), .dout(n2201));
    jxor g0500(.dinb(n2186), .dina(n2201), .dout(n2205));
    jand g0501(.dinb(G18), .dina(G180), .dout(n2209));
    jor g0502(.dinb(n896), .dina(n9284), .dout(n2213));
    jor g0503(.dinb(n455), .dina(n892), .dout(n2217));
    jor g0504(.dinb(G18), .dina(G83), .dout(n2221));
    jand g0505(.dinb(n2217), .dina(n9566), .dout(n2225));
    jxor g0506(.dinb(n2213), .dina(n2225), .dout(n2229));
    jand g0507(.dinb(n2205), .dina(n2229), .dout(n2233));
    jand g0508(.dinb(G18), .dina(G171), .dout(n2237));
    jor g0509(.dinb(n915), .dina(n9311), .dout(n2241));
    jor g0510(.dinb(n455), .dina(n911), .dout(n2245));
    jor g0511(.dinb(G18), .dina(G65), .dout(n2249));
    jand g0512(.dinb(n2245), .dina(n9584), .dout(n2253));
    jand g0513(.dinb(n2241), .dina(n2253), .dout(n2257));
    jand g0514(.dinb(n2233), .dina(n8324), .dout(n2261));
    jand g0515(.dinb(n2186), .dina(n2201), .dout(n2265));
    jor g0516(.dinb(n2186), .dina(n2201), .dout(n2269));
    jand g0517(.dinb(n2213), .dina(n2225), .dout(n2273));
    jand g0518(.dinb(n2269), .dina(n2273), .dout(n2277));
    jor g0519(.dinb(n8321), .dina(n2277), .dout(n2281));
    jor g0520(.dinb(n2261), .dina(n2281), .dout(n2285));
    jand g0521(.dinb(n8326), .dina(n2285), .dout(n2289));
    jand g0522(.dinb(n2131), .dina(n2146), .dout(n2293));
    jor g0523(.dinb(n2131), .dina(n2146), .dout(n2297));
    jand g0524(.dinb(n2158), .dina(n2170), .dout(n2301));
    jand g0525(.dinb(n2297), .dina(n2301), .dout(n2305));
    jor g0526(.dinb(n8318), .dina(n2305), .dout(n2309));
    jor g0527(.dinb(n2289), .dina(n8315), .dout(n2313));
    jand g0528(.dinb(n2178), .dina(n2233), .dout(n2317));
    jand g0529(.dinb(G18), .dina(G189), .dout(n2321));
    jor g0530(.dinb(n1013), .dina(n9368), .dout(n2325));
    jor g0531(.dinb(n455), .dina(n1005), .dout(n2329));
    jor g0532(.dinb(G18), .dina(G62), .dout(n2333));
    jand g0533(.dinb(n2329), .dina(n9518), .dout(n2337));
    jxor g0534(.dinb(n2325), .dina(n2337), .dout(n2341));
    jand g0535(.dinb(G18), .dina(G190), .dout(n2345));
    jor g0536(.dinb(n1042), .dina(n9362), .dout(n2349));
    jor g0537(.dinb(n455), .dina(n1034), .dout(n2353));
    jor g0538(.dinb(G18), .dina(G61), .dout(n2357));
    jand g0539(.dinb(n2353), .dina(n9515), .dout(n2361));
    jxor g0540(.dinb(n2349), .dina(n2361), .dout(n2365));
    jand g0541(.dinb(n2341), .dina(n2365), .dout(n2369));
    jand g0542(.dinb(G18), .dina(G191), .dout(n2373));
    jor g0543(.dinb(n1083), .dina(n9395), .dout(n2377));
    jand g0544(.dinb(G18), .dina(G4427), .dout(n2381));
    jnot g0545(.din(n2381), .dout(n2384));
    jor g0546(.dinb(G18), .dina(G60), .dout(n2388));
    jand g0547(.dinb(n2384), .dina(n9512), .dout(n2392));
    jand g0548(.dinb(n2377), .dina(n2392), .dout(n2396));
    jor g0549(.dinb(n2377), .dina(n2392), .dout(n2400));
    jand g0550(.dinb(G18), .dina(G192), .dout(n2404));
    jor g0551(.dinb(n1061), .dina(n9392), .dout(n2408));
    jand g0552(.dinb(G18), .dina(G4420), .dout(n2412));
    jnot g0553(.din(n2412), .dout(n2415));
    jor g0554(.dinb(G18), .dina(G79), .dout(n2419));
    jand g0555(.dinb(n2415), .dina(n9509), .dout(n2423));
    jand g0556(.dinb(n2408), .dina(n2423), .dout(n2427));
    jand g0557(.dinb(n2400), .dina(n2427), .dout(n2431));
    jor g0558(.dinb(n8797), .dina(n2431), .dout(n2435));
    jand g0559(.dinb(n8800), .dina(n2435), .dout(n2439));
    jand g0560(.dinb(n2325), .dina(n2337), .dout(n2443));
    jor g0561(.dinb(n2325), .dina(n2337), .dout(n2447));
    jand g0562(.dinb(n2349), .dina(n2361), .dout(n2451));
    jand g0563(.dinb(n2447), .dina(n2451), .dout(n2455));
    jor g0564(.dinb(n8795), .dina(n2455), .dout(n2459));
    jor g0565(.dinb(n2439), .dina(n8792), .dout(n2463));
    jor g0566(.dinb(n2408), .dina(n2423), .dout(n2467));
    jand g0567(.dinb(n2400), .dina(n2467), .dout(n2471));
    jand g0568(.dinb(n2369), .dina(n2471), .dout(n2475));
    jand g0569(.dinb(G18), .dina(G205), .dout(n2479));
    jor g0570(.dinb(n1482), .dina(n9410), .dout(n2483));
    jor g0571(.dinb(n455), .dina(n1474), .dout(n2487));
    jor g0572(.dinb(G18), .dina(G75), .dout(n2491));
    jand g0573(.dinb(n2487), .dina(n9542), .dout(n2495));
    jor g0574(.dinb(n2483), .dina(n2495), .dout(n2499));
    jand g0575(.dinb(G18), .dina(G206), .dout(n2503));
    jor g0576(.dinb(n1501), .dina(n9404), .dout(n2507));
    jor g0577(.dinb(n455), .dina(n1493), .dout(n2511));
    jor g0578(.dinb(G18), .dina(G76), .dout(n2515));
    jand g0579(.dinb(n2511), .dina(n9548), .dout(n2519));
    jand g0580(.dinb(n2507), .dina(n2519), .dout(n2523));
    jor g0581(.dinb(G70), .dina(G89), .dout(n2527));
    jand g0582(.dinb(n1609), .dina(n8783), .dout(n2531));
    jor g0583(.dinb(n2523), .dina(n8780), .dout(n2535));
    jand g0584(.dinb(G18), .dina(G207), .dout(n2539));
    jor g0585(.dinb(n1594), .dina(n9401), .dout(n2543));
    jor g0586(.dinb(n455), .dina(n1586), .dout(n2547));
    jor g0587(.dinb(G18), .dina(G74), .dout(n2551));
    jand g0588(.dinb(n2547), .dina(n9545), .dout(n2555));
    jand g0589(.dinb(n2543), .dina(n2555), .dout(n2559));
    jor g0590(.dinb(G18), .dina(G70), .dout(n2563));
    jand g0591(.dinb(n8785), .dina(n2563), .dout(n2567));
    jor g0592(.dinb(n2559), .dina(n8777), .dout(n2571));
    jor g0593(.dinb(n2535), .dina(n2571), .dout(n2575));
    jor g0594(.dinb(n2543), .dina(n2555), .dout(n2579));
    jor g0595(.dinb(n2507), .dina(n2519), .dout(n2583));
    jand g0596(.dinb(n2579), .dina(n2583), .dout(n2587));
    jor g0597(.dinb(n8788), .dina(n2587), .dout(n2591));
    jand g0598(.dinb(n2575), .dina(n2591), .dout(n2595));
    jand g0599(.dinb(n8771), .dina(n2595), .dout(n2599));
    jand g0600(.dinb(G18), .dina(G204), .dout(n2603));
    jor g0601(.dinb(n1463), .dina(n9407), .dout(n2607));
    jor g0602(.dinb(n455), .dina(n1455), .dout(n2611));
    jor g0603(.dinb(G18), .dina(G73), .dout(n2615));
    jand g0604(.dinb(n2611), .dina(n9536), .dout(n2619));
    jand g0605(.dinb(n2607), .dina(n2619), .dout(n2623));
    jand g0606(.dinb(n2483), .dina(n2495), .dout(n2627));
    jor g0607(.dinb(n2623), .dina(n2627), .dout(n2631));
    jor g0608(.dinb(n2599), .dina(n8762), .dout(n2635));
    jor g0609(.dinb(n2607), .dina(n2619), .dout(n2639));
    jand g0610(.dinb(G18), .dina(G203), .dout(n2643));
    jor g0611(.dinb(n1382), .dina(n9437), .dout(n2647));
    jand g0612(.dinb(G18), .dina(G3729), .dout(n2651));
    jnot g0613(.din(n2651), .dout(n2654));
    jor g0614(.dinb(G18), .dina(G53), .dout(n2658));
    jand g0615(.dinb(n2654), .dina(n9530), .dout(n2662));
    jor g0616(.dinb(n2647), .dina(n2662), .dout(n2666));
    jand g0617(.dinb(n2639), .dina(n2666), .dout(n2670));
    jand g0618(.dinb(n2635), .dina(n8753), .dout(n2674));
    jand g0619(.dinb(G18), .dina(G202), .dout(n2678));
    jor g0620(.dinb(n1363), .dina(n9431), .dout(n2682));
    jor g0621(.dinb(n455), .dina(n1355), .dout(n2686));
    jor g0622(.dinb(G18), .dina(G54), .dout(n2690));
    jand g0623(.dinb(n2686), .dina(n9527), .dout(n2694));
    jand g0624(.dinb(n2682), .dina(n2694), .dout(n2698));
    jand g0625(.dinb(n2647), .dina(n2662), .dout(n2702));
    jor g0626(.dinb(n2698), .dina(n2702), .dout(n2706));
    jor g0627(.dinb(n2674), .dina(n8741), .dout(n2710));
    jand g0628(.dinb(G18), .dina(G201), .dout(n2714));
    jor g0629(.dinb(n1344), .dina(n9428), .dout(n2718));
    jor g0630(.dinb(n455), .dina(n1336), .dout(n2722));
    jor g0631(.dinb(G18), .dina(G55), .dout(n2726));
    jand g0632(.dinb(n2722), .dina(n9554), .dout(n2730));
    jxor g0633(.dinb(n2718), .dina(n2730), .dout(n2734));
    jand g0634(.dinb(G18), .dina(G200), .dout(n2738));
    jor g0635(.dinb(n1315), .dina(n9425), .dout(n2742));
    jor g0636(.dinb(n455), .dina(n1307), .dout(n2746));
    jor g0637(.dinb(G18), .dina(G56), .dout(n2750));
    jand g0638(.dinb(n2746), .dina(n9551), .dout(n2754));
    jxor g0639(.dinb(n2742), .dina(n2754), .dout(n2758));
    jand g0640(.dinb(n2734), .dina(n2758), .dout(n2762));
    jor g0641(.dinb(n2682), .dina(n2694), .dout(n2766));
    jand g0642(.dinb(n2762), .dina(n8726), .dout(n2770));
    jand g0643(.dinb(n2710), .dina(n8723), .dout(n2774));
    jand g0644(.dinb(n2742), .dina(n2754), .dout(n2778));
    jand g0645(.dinb(n2718), .dina(n2730), .dout(n2782));
    jor g0646(.dinb(n2742), .dina(n2754), .dout(n2786));
    jand g0647(.dinb(n2782), .dina(n2786), .dout(n2790));
    jor g0648(.dinb(n8708), .dina(n2790), .dout(n2794));
    jor g0649(.dinb(n2774), .dina(n8705), .dout(n2798));
    jand g0650(.dinb(G18), .dina(G187), .dout(n2802));
    jor g0651(.dinb(n1228), .dina(n9377), .dout(n2806));
    jand g0652(.dinb(G18), .dina(G4394), .dout(n2810));
    jnot g0653(.din(n2810), .dout(n2813));
    jor g0654(.dinb(G18), .dina(G77), .dout(n2817));
    jand g0655(.dinb(n2813), .dina(n9500), .dout(n2821));
    jor g0656(.dinb(n2806), .dina(n2821), .dout(n2825));
    jand g0657(.dinb(G18), .dina(G193), .dout(n2829));
    jor g0658(.dinb(n1112), .dina(n9383), .dout(n2833));
    jand g0659(.dinb(G18), .dina(G4415), .dout(n2837));
    jnot g0660(.din(n2837), .dout(n2840));
    jor g0661(.dinb(G18), .dina(G80), .dout(n2844));
    jand g0662(.dinb(n2840), .dina(n9506), .dout(n2848));
    jxor g0663(.dinb(n2833), .dina(n2848), .dout(n2852));
    jand g0664(.dinb(G18), .dina(G194), .dout(n2856));
    jor g0665(.dinb(n1141), .dina(n9380), .dout(n2860));
    jor g0666(.dinb(n455), .dina(n1133), .dout(n2864));
    jor g0667(.dinb(G18), .dina(G81), .dout(n2868));
    jand g0668(.dinb(n2864), .dina(n9503), .dout(n2872));
    jxor g0669(.dinb(n2860), .dina(n2872), .dout(n2876));
    jand g0670(.dinb(n2852), .dina(n2876), .dout(n2880));
    jand g0671(.dinb(G18), .dina(G196), .dout(n2884));
    jor g0672(.dinb(n1199), .dina(n9389), .dout(n2888));
    jand g0673(.dinb(G18), .dina(G4400), .dout(n2892));
    jnot g0674(.din(n2892), .dout(n2895));
    jor g0675(.dinb(G18), .dina(G78), .dout(n2899));
    jand g0676(.dinb(n2895), .dina(n9491), .dout(n2903));
    jand g0677(.dinb(n2888), .dina(n2903), .dout(n2907));
    jnot g0678(.din(n2907), .dout(n2910));
    jand g0679(.dinb(G18), .dina(G195), .dout(n2914));
    jor g0680(.dinb(n1170), .dina(n9386), .dout(n2918));
    jand g0681(.dinb(G18), .dina(G4405), .dout(n2922));
    jnot g0682(.din(n2922), .dout(n2925));
    jor g0683(.dinb(G18), .dina(G59), .dout(n2929));
    jand g0684(.dinb(n2925), .dina(n9485), .dout(n2933));
    jor g0685(.dinb(n2918), .dina(n2933), .dout(n2937));
    jand g0686(.dinb(n2910), .dina(n8680), .dout(n2941));
    jor g0687(.dinb(n2888), .dina(n2903), .dout(n2945));
    jand g0688(.dinb(n2918), .dina(n2933), .dout(n2949));
    jnot g0689(.din(n2949), .dout(n2952));
    jand g0690(.dinb(n8675), .dina(n2952), .dout(n2956));
    jand g0691(.dinb(n2941), .dina(n2956), .dout(n2960));
    jand g0692(.dinb(n8683), .dina(n2960), .dout(n2964));
    jand g0693(.dinb(n2806), .dina(n2821), .dout(n2968));
    jnot g0694(.din(n2968), .dout(n2971));
    jand g0695(.dinb(n2964), .dina(n8660), .dout(n2975));
    jand g0696(.dinb(n8651), .dina(n2975), .dout(n2979));
    jand g0697(.dinb(n2798), .dina(n8636), .dout(n2983));
    jand g0698(.dinb(n2833), .dina(n2848), .dout(n2987));
    jor g0699(.dinb(n2833), .dina(n2848), .dout(n2991));
    jand g0700(.dinb(n2860), .dina(n2872), .dout(n2995));
    jand g0701(.dinb(n2991), .dina(n2995), .dout(n2999));
    jor g0702(.dinb(n8627), .dina(n2999), .dout(n3003));
    jand g0703(.dinb(n2964), .dina(n8662), .dout(n3007));
    jand g0704(.dinb(n2907), .dina(n2937), .dout(n3011));
    jor g0705(.dinb(n8677), .dina(n3011), .dout(n3015));
    jand g0706(.dinb(n8687), .dina(n3015), .dout(n3019));
    jor g0707(.dinb(n3007), .dina(n8624), .dout(n3023));
    jor g0708(.dinb(n8618), .dina(n3023), .dout(n3027));
    jor g0709(.dinb(n2983), .dina(n8606), .dout(n3031));
    jnot g0710(.din(n2396), .dout(n3034));
    jnot g0711(.din(n2427), .dout(n3037));
    jand g0712(.dinb(n3034), .dina(n3037), .dout(n3041));
    jand g0713(.dinb(n3031), .dina(n8597), .dout(n3045));
    jand g0714(.dinb(n8570), .dina(n3045), .dout(n3049));
    jor g0715(.dinb(n8540), .dina(n3049), .dout(n3053));
    jxor g0716(.dinb(n2241), .dina(n2253), .dout(n3057));
    jand g0717(.dinb(n3053), .dina(n8309), .dout(n3061));
    jand g0718(.dinb(n8267), .dina(n3061), .dout(n3065));
    jor g0719(.dinb(n8228), .dina(n3065), .dout(n3069));
    jor g0720(.dinb(n2054), .dina(n2069), .dout(n3073));
    jand g0721(.dinb(n2046), .dina(n3073), .dout(n3077));
    jand g0722(.dinb(n3069), .dina(n8195), .dout(n3081));
    jand g0723(.dinb(n8147), .dina(n3081), .dout(n3085));
    jor g0724(.dinb(n8102), .dina(n3085), .dout(n3089));
    jxor g0725(.dinb(n9307), .dina(n1888), .dout(n3093));
    jxor g0726(.dinb(n1856), .dina(n1868), .dout(n3097));
    jand g0727(.dinb(n1848), .dina(n3097), .dout(n3101));
    jand g0728(.dinb(n1947), .dina(n3101), .dout(n3105));
    jand g0729(.dinb(n8054), .dina(n3105), .dout(n3109));
    jand g0730(.dinb(n3089), .dina(n8048), .dout(n3113));
    jor g0731(.dinb(G1455), .dina(G2204), .dout(n3117));
    jor g0732(.dinb(n499), .dina(n3117), .dout(n3121));
    jand g0733(.dinb(n9904), .dina(n3121), .dout(n3125));
    jand g0734(.dinb(n1832), .dina(n1844), .dout(n3129));
    jand g0735(.dinb(n1900), .dina(n1915), .dout(n3133));
    jor g0736(.dinb(n1900), .dina(n1915), .dout(n3137));
    jand g0737(.dinb(n1927), .dina(n1939), .dout(n3141));
    jand g0738(.dinb(n3137), .dina(n3141), .dout(n3145));
    jor g0739(.dinb(n7997), .dina(n3145), .dout(n3149));
    jand g0740(.dinb(n8056), .dina(n3149), .dout(n3153));
    jor g0741(.dinb(n7994), .dina(n3153), .dout(n3157));
    jor g0742(.dinb(n7985), .dina(n3157), .dout(n3161));
    jor g0743(.dinb(n3113), .dina(n7970), .dout(n3165));
    jor g0744(.dinb(n7922), .dina(n3165), .dout(n3169));
    jand g0745(.dinb(n8444), .dina(n3169), .dout(n3173));
    jnot g0746(.din(n1539), .dout(n3176));
    jnot g0747(.din(n1579), .dout(n3179));
    jnot g0748(.din(n1583), .dout(n3182));
    jand g0749(.dinb(n18352), .dina(n1527), .dout(n3186));
    jor g0750(.dinb(n18370), .dina(n1527), .dout(n3190));
    jand g0751(.dinb(n18389), .dina(n3190), .dout(n3194));
    jor g0752(.dinb(n18224), .dina(n3194), .dout(n3198));
    jor g0753(.dinb(n18221), .dina(n3198), .dout(n3202));
    jand g0754(.dinb(n18218), .dina(n3202), .dout(n3206));
    jand g0755(.dinb(n3176), .dina(n3206), .dout(n3210));
    jnot g0756(.din(n3210), .dout(n3213));
    jor g0757(.dinb(n17242), .dina(n1633), .dout(n3217));
    jand g0758(.dinb(n3213), .dina(n7868), .dout(n3221));
    jor g0759(.dinb(n18241), .dina(n3221), .dout(n3225));
    jand g0760(.dinb(n17743), .dina(n3225), .dout(n3229));
    jxor g0761(.dinb(n18499), .dina(n3229), .dout(n3233));
    jxor g0762(.dinb(n18439), .dina(n3221), .dout(n3237));
    jand g0763(.dinb(n17845), .dina(n470), .dout(n3241));
    jor g0764(.dinb(n3241), .dina(n17701), .dout(n3245));
    jand g0765(.dinb(n17716), .dina(n3245), .dout(n3249));
    jxor g0766(.dinb(n18400), .dina(n3249), .dout(n3253));
    jor g0767(.dinb(n17704), .dina(n3241), .dout(n3257));
    jxor g0768(.dinb(n18340), .dina(n3257), .dout(n3261));
    jxor g0769(.dinb(n18055), .dina(n1319), .dout(n3265));
    jor g0770(.dinb(n1669), .dina(n18013), .dout(n3269));
    jnot g0771(.din(n1547), .dout(n3272));
    jnot g0772(.din(n1551), .dout(n3275));
    jnot g0773(.din(n1575), .dout(n3278));
    jand g0774(.dinb(n18212), .dina(n3206), .dout(n3282));
    jor g0775(.dinb(n18274), .dina(n3282), .dout(n3286));
    jor g0776(.dinb(n18286), .dina(n3286), .dout(n3290));
    jand g0777(.dinb(n18203), .dina(n3290), .dout(n3294));
    jand g0778(.dinb(n18329), .dina(n3294), .dout(n3298));
    jnot g0779(.din(G4526), .dout(n3301));
    jand g0780(.dinb(n17801), .dina(n3294), .dout(n3305));
    jor g0781(.dinb(n3298), .dina(n3305), .dout(n3309));
    jand g0782(.dinb(n17566), .dina(n3309), .dout(n3313));
    jor g0783(.dinb(n17545), .dina(n3313), .dout(n3317));
    jor g0784(.dinb(n17272), .dina(n3317), .dout(n3321));
    jor g0785(.dinb(n17305), .dina(n3321), .dout(n3325));
    jand g0786(.dinb(n7871), .dina(n3325), .dout(n3329));
    jand g0787(.dinb(n17593), .dina(n1661), .dout(n3333));
    jor g0788(.dinb(n17947), .dina(n3333), .dout(n3337));
    jxor g0789(.dinb(n17650), .dina(n3337), .dout(n3341));
    jnot g0790(.din(n1371), .dout(n3344));
    jnot g0791(.din(n1423), .dout(n3347));
    jnot g0792(.din(n1386), .dout(n3350));
    jand g0793(.dinb(n18112), .dina(n3350), .dout(n3354));
    jor g0794(.dinb(n18079), .dina(n3309), .dout(n3358));
    jand g0795(.dinb(n17515), .dina(n3358), .dout(n3362));
    jxor g0796(.dinb(n18124), .dina(n3362), .dout(n3366));
    jxor g0797(.dinb(n17620), .dina(n1661), .dout(n3370));
    jnot g0798(.din(n758), .dout(n3373));
    jor g0799(.dinb(n14959), .dina(n3373), .dout(n3377));
    jnot g0800(.din(n743), .dout(n3380));
    jor g0801(.dinb(n3380), .dina(n14836), .dout(n3384));
    jand g0802(.dinb(n3377), .dina(n3384), .dout(n3388));
    jnot g0803(.din(n846), .dout(n3391));
    jxor g0804(.dinb(n14362), .dina(n3391), .dout(n3395));
    jxor g0805(.dinb(n3388), .dina(n9266), .dout(n3399));
    jxor g0806(.dinb(n13822), .dina(n945), .dout(n3403));
    jor g0807(.dinb(n15349), .dina(n773), .dout(n3407));
    jnot g0808(.din(n709), .dout(n3410));
    jor g0809(.dinb(n3410), .dina(n15061), .dout(n3414));
    jand g0810(.dinb(n3407), .dina(n3414), .dout(n3418));
    jnot g0811(.din(G141), .dout(n3421));
    jor g0812(.dinb(n9487), .dina(n3421), .dout(n3425));
    jnot g0813(.din(G161), .dout(n3428));
    jor g0814(.dinb(n455), .dina(n3428), .dout(n3432));
    jand g0815(.dinb(n3425), .dina(n3432), .dout(n3436));
    jxor g0816(.dinb(n923), .dina(n3436), .dout(n3440));
    jxor g0817(.dinb(n3418), .dina(n9263), .dout(n3444));
    jxor g0818(.dinb(n9257), .dina(n3444), .dout(n3448));
    jxor g0819(.dinb(n9251), .dina(n3448), .dout(n3452));
    jxor g0820(.dinb(n1367), .dina(n1386), .dout(n3456));
    jand g0821(.dinb(G18), .dina(G239), .dout(n3460));
    jand g0822(.dinb(n455), .dina(n9419), .dout(n3464));
    jor g0823(.dinb(n9248), .dina(n3464), .dout(n3468));
    jxor g0824(.dinb(n1564), .dina(n9245), .dout(n3472));
    jxor g0825(.dinb(n9242), .dina(n3472), .dout(n3476));
    jand g0826(.dinb(G18), .dina(G229), .dout(n3480));
    jor g0827(.dinb(n1609), .dina(n9239), .dout(n3484));
    jxor g0828(.dinb(n1598), .dina(n3484), .dout(n3488));
    jxor g0829(.dinb(n1467), .dina(n1505), .dout(n3492));
    jxor g0830(.dinb(n3488), .dina(n3492), .dout(n3496));
    jxor g0831(.dinb(n1319), .dina(n1348), .dout(n3500));
    jxor g0832(.dinb(n3496), .dina(n9236), .dout(n3504));
    jxor g0833(.dinb(n3476), .dina(n3504), .dout(n3508));
    jor g0834(.dinb(n3452), .dina(n9233), .dout(n3512));
    jor g0835(.dinb(n455), .dina(n518), .dout(n3516));
    jxor g0836(.dinb(G211), .dina(G212), .dout(n3520));
    jxor g0837(.dinb(n12656), .dina(n3520), .dout(n3524));
    jor g0838(.dinb(n3516), .dina(n3524), .dout(n3528));
    jnot g0839(.din(n569), .dout(n3531));
    jand g0840(.dinb(n3531), .dina(n603), .dout(n3535));
    jnot g0841(.din(n599), .dout(n3538));
    jand g0842(.dinb(n573), .dina(n3538), .dout(n3542));
    jor g0843(.dinb(n3535), .dina(n3542), .dout(n3546));
    jor g0844(.dinb(n12703), .dina(n548), .dout(n3550));
    jnot g0845(.din(n529), .dout(n3553));
    jor g0846(.dinb(n3553), .dina(n15466), .dout(n3557));
    jand g0847(.dinb(n3550), .dina(n3557), .dout(n3561));
    jxor g0848(.dinb(n9227), .dina(n3561), .dout(n3565));
    jxor g0849(.dinb(n9224), .dina(n3565), .dout(n3569));
    jxor g0850(.dinb(n15994), .dina(n1711), .dout(n3573));
    jxor g0851(.dinb(n1065), .dina(n1087), .dout(n3577));
    jxor g0852(.dinb(n3573), .dina(n9212), .dout(n3581));
    jxor g0853(.dinb(n1145), .dina(n1203), .dout(n3585));
    jxor g0854(.dinb(n1116), .dina(n1174), .dout(n3589));
    jxor g0855(.dinb(n3585), .dina(n3589), .dout(n3593));
    jand g0856(.dinb(G18), .dina(G227), .dout(n3597));
    jand g0857(.dinb(n455), .dina(n9374), .dout(n3601));
    jor g0858(.dinb(n9209), .dina(n3601), .dout(n3605));
    jxor g0859(.dinb(n1232), .dina(n3605), .dout(n3609));
    jxor g0860(.dinb(n3593), .dina(n9206), .dout(n3613));
    jxor g0861(.dinb(n3581), .dina(n3613), .dout(n3617));
    jor g0862(.dinb(n3569), .dina(n9203), .dout(n3621));
    jor g0863(.dinb(n3512), .dina(n9200), .dout(n3625));
    jnot g0864(.din(n2038), .dout(n3628));
    jxor g0865(.dinb(n3628), .dina(n9586), .dout(n3632));
    jnot g0866(.din(G2208), .dout(n3635));
    jor g0867(.dinb(n455), .dina(n3635), .dout(n3639));
    jor g0868(.dinb(G18), .dina(G82), .dout(n3643));
    jand g0869(.dinb(n3639), .dina(n9581), .dout(n3647));
    jxor g0870(.dinb(n2253), .dina(n3647), .dout(n3651));
    jxor g0871(.dinb(n3632), .dina(n9578), .dout(n3655));
    jxor g0872(.dinb(n2146), .dina(n2170), .dout(n3659));
    jxor g0873(.dinb(n2201), .dina(n2225), .dout(n3663));
    jxor g0874(.dinb(n3659), .dina(n3663), .dout(n3667));
    jxor g0875(.dinb(n1983), .dina(n2007), .dout(n3671));
    jxor g0876(.dinb(n3667), .dina(n9557), .dout(n3675));
    jxor g0877(.dinb(n3655), .dina(n3675), .dout(n3679));
    jxor g0878(.dinb(n2730), .dina(n2754), .dout(n3683));
    jxor g0879(.dinb(n2519), .dina(n2555), .dout(n3687));
    jxor g0880(.dinb(n3683), .dina(n3687), .dout(n3691));
    jnot g0881(.din(G3698), .dout(n3694));
    jor g0882(.dinb(n455), .dina(n3694), .dout(n3698));
    jor g0883(.dinb(G18), .dina(G69), .dout(n3702));
    jand g0884(.dinb(n3698), .dina(n9539), .dout(n3706));
    jxor g0885(.dinb(n2495), .dina(n3706), .dout(n3710));
    jor g0886(.dinb(n455), .dina(n1605), .dout(n3714));
    jand g0887(.dinb(n9532), .dina(n3714), .dout(n3718));
    jxor g0888(.dinb(n2619), .dina(n3718), .dout(n3722));
    jxor g0889(.dinb(n3710), .dina(n3722), .dout(n3726));
    jnot g0890(.din(n2662), .dout(n3729));
    jxor g0891(.dinb(n3729), .dina(n9523), .dout(n3733));
    jxor g0892(.dinb(n3726), .dina(n3733), .dout(n3737));
    jxor g0893(.dinb(n9521), .dina(n3737), .dout(n3741));
    jor g0894(.dinb(n3679), .dina(n3741), .dout(n3745));
    jxor g0895(.dinb(n2337), .dina(n2361), .dout(n3749));
    jxor g0896(.dinb(n2392), .dina(n2423), .dout(n3753));
    jxor g0897(.dinb(n3749), .dina(n3753), .dout(n3757));
    jxor g0898(.dinb(n2848), .dina(n2872), .dout(n3761));
    jand g0899(.dinb(G18), .dina(G4393), .dout(n3765));
    jnot g0900(.din(G58), .dout(n3768));
    jand g0901(.dinb(n455), .dina(n3768), .dout(n3772));
    jor g0902(.dinb(n9494), .dina(n3772), .dout(n3776));
    jxor g0903(.dinb(n2821), .dina(n3776), .dout(n3780));
    jxor g0904(.dinb(n2903), .dina(n2933), .dout(n3784));
    jxor g0905(.dinb(n3780), .dina(n3784), .dout(n3788));
    jxor g0906(.dinb(n9482), .dina(n3788), .dout(n3792));
    jxor g0907(.dinb(n9479), .dina(n3792), .dout(n3796));
    jxor g0908(.dinb(n11080), .dina(n496), .dout(n3800));
    jor g0909(.dinb(n9496), .dina(n3800), .dout(n3804));
    jnot g0910(.din(G1455), .dout(n3807));
    jxor g0911(.dinb(n3807), .dina(n9469), .dout(n3811));
    jor g0912(.dinb(n9472), .dina(n3811), .dout(n3815));
    jand g0913(.dinb(n3804), .dina(n3815), .dout(n3819));
    jxor g0914(.dinb(n1844), .dina(n1868), .dout(n3823));
    jxor g0915(.dinb(n1915), .dina(n1939), .dout(n3827));
    jxor g0916(.dinb(n3823), .dina(n3827), .dout(n3831));
    jnot g0917(.din(G1459), .dout(n3834));
    jor g0918(.dinb(n455), .dina(n3834), .dout(n3838));
    jor g0919(.dinb(G18), .dina(G114), .dout(n3842));
    jand g0920(.dinb(n3838), .dina(n9452), .dout(n3846));
    jxor g0921(.dinb(n1888), .dina(n3846), .dout(n3850));
    jxor g0922(.dinb(n3831), .dina(n9449), .dout(n3854));
    jxor g0923(.dinb(n9446), .dina(n3854), .dout(n3858));
    jor g0924(.dinb(n3796), .dina(n3858), .dout(n3862));
    jor g0925(.dinb(n3745), .dina(n3862), .dout(n3866));
    jnot g0926(.din(n2682), .dout(n3869));
    jxor g0927(.dinb(n9433), .dina(n3869), .dout(n3873));
    jxor g0928(.dinb(n2718), .dina(n2742), .dout(n3877));
    jxor g0929(.dinb(n3873), .dina(n9422), .dout(n3881));
    jand g0930(.dinb(G18), .dina(G208), .dout(n3885));
    jor g0931(.dinb(n3464), .dina(n9416), .dout(n3889));
    jand g0932(.dinb(G18), .dina(G198), .dout(n3893));
    jor g0933(.dinb(n1609), .dina(n9413), .dout(n3897));
    jxor g0934(.dinb(n3889), .dina(n3897), .dout(n3901));
    jxor g0935(.dinb(n2483), .dina(n2607), .dout(n3905));
    jxor g0936(.dinb(n3901), .dina(n3905), .dout(n3909));
    jxor g0937(.dinb(n2507), .dina(n2543), .dout(n3913));
    jxor g0938(.dinb(n3909), .dina(n9398), .dout(n3917));
    jxor g0939(.dinb(n3881), .dina(n3917), .dout(n3921));
    jxor g0940(.dinb(n2377), .dina(n2408), .dout(n3925));
    jxor g0941(.dinb(n2888), .dina(n2918), .dout(n3929));
    jxor g0942(.dinb(n3925), .dina(n3929), .dout(n3933));
    jxor g0943(.dinb(n2833), .dina(n2860), .dout(n3937));
    jand g0944(.dinb(G18), .dina(G197), .dout(n3941));
    jor g0945(.dinb(n3601), .dina(n9371), .dout(n3945));
    jxor g0946(.dinb(n2806), .dina(n3945), .dout(n3949));
    jxor g0947(.dinb(n3937), .dina(n3949), .dout(n3953));
    jnot g0948(.din(n2349), .dout(n3956));
    jxor g0949(.dinb(n9364), .dina(n3956), .dout(n3960));
    jxor g0950(.dinb(n3953), .dina(n3960), .dout(n3964));
    jxor g0951(.dinb(n9359), .dina(n3964), .dout(n3968));
    jor g0952(.dinb(n3921), .dina(n3968), .dout(n3972));
    jxor g0953(.dinb(G164), .dina(G165), .dout(n3976));
    jxor g0954(.dinb(n9356), .dina(n3976), .dout(n3980));
    jor g0955(.dinb(n3516), .dina(n3980), .dout(n3984));
    jnot g0956(.din(n1896), .dout(n3987));
    jand g0957(.dinb(n3987), .dina(n1927), .dout(n3991));
    jnot g0958(.din(n1923), .dout(n3994));
    jand g0959(.dinb(n1900), .dina(n3994), .dout(n3998));
    jor g0960(.dinb(n3991), .dina(n3998), .dout(n4002));
    jnot g0961(.din(n1856), .dout(n4005));
    jor g0962(.dinb(n9337), .dina(n4005), .dout(n4009));
    jnot g0963(.din(n1832), .dout(n4012));
    jor g0964(.dinb(n4012), .dina(n9328), .dout(n4016));
    jand g0965(.dinb(n4009), .dina(n4016), .dout(n4020));
    jxor g0966(.dinb(n9326), .dina(n4020), .dout(n4024));
    jxor g0967(.dinb(n9323), .dina(n4024), .dout(n4028));
    jor g0968(.dinb(n3972), .dina(n4028), .dout(n4032));
    jnot g0969(.din(G181), .dout(n4035));
    jor g0970(.dinb(n455), .dina(n4035), .dout(n4039));
    jand g0971(.dinb(n3425), .dina(n4039), .dout(n4043));
    jxor g0972(.dinb(n2241), .dina(n4043), .dout(n4047));
    jxor g0973(.dinb(n2131), .dina(n2158), .dout(n4051));
    jxor g0974(.dinb(n4047), .dina(n4051), .dout(n4055));
    jnot g0975(.din(n2019), .dout(n4058));
    jand g0976(.dinb(n4058), .dina(n2054), .dout(n4062));
    jnot g0977(.din(n2050), .dout(n4065));
    jand g0978(.dinb(n2023), .dina(n4065), .dout(n4069));
    jor g0979(.dinb(n4062), .dina(n4069), .dout(n4073));
    jnot g0980(.din(n1967), .dout(n4076));
    jand g0981(.dinb(n4076), .dina(n1995), .dout(n4080));
    jnot g0982(.din(n1991), .dout(n4083));
    jand g0983(.dinb(n1971), .dina(n4083), .dout(n4087));
    jor g0984(.dinb(n4080), .dina(n4087), .dout(n4091));
    jxor g0985(.dinb(n4073), .dina(n4091), .dout(n4095));
    jxor g0986(.dinb(n2186), .dina(n2213), .dout(n4099));
    jxor g0987(.dinb(n4095), .dina(n9281), .dout(n4103));
    jxor g0988(.dinb(n9275), .dina(n4103), .dout(n4107));
    jor g0989(.dinb(n4032), .dina(n9269), .dout(n4111));
    jnot g0990(.din(n927), .dout(n4114));
    jnot g0991(.din(n1021), .dout(n4117));
    jnot g0992(.din(n1050), .dout(n4120));
    jnot g0993(.din(n1091), .dout(n4123));
    jnot g0994(.din(n1268), .dout(n4126));
    jnot g0995(.din(n1304), .dout(n4129));
    jnot g0996(.din(n1323), .dout(n4132));
    jand g0997(.dinb(n15812), .dina(n3321), .dout(n4136));
    jor g0998(.dinb(n16636), .dina(n4136), .dout(n4140));
    jand g0999(.dinb(n16375), .dina(n4140), .dout(n4144));
    jor g1000(.dinb(n16078), .dina(n4144), .dout(n4148));
    jor g1001(.dinb(n16027), .dina(n4148), .dout(n4152));
    jor g1002(.dinb(n16234), .dina(n4152), .dout(n4156));
    jor g1003(.dinb(n12152), .dina(n4156), .dout(n4160));
    jand g1004(.dinb(n4160), .dina(n12823), .dout(n4164));
    jor g1005(.dinb(n13027), .dina(n4164), .dout(n4168));
    jand g1006(.dinb(n12095), .dina(n4168), .dout(n4172));
    jxor g1007(.dinb(n8513), .dina(n4172), .dout(n4176));
    jnot g1008(.din(n674), .dout(n4179));
    jnot g1009(.din(n713), .dout(n4182));
    jnot g1010(.din(n717), .dout(n4185));
    jnot g1011(.din(n812), .dout(n4188));
    jnot g1012(.din(n808), .dout(n4191));
    jnot g1013(.din(n998), .dout(n4194));
    jnot g1014(.din(n1002), .dout(n4197));
    jnot g1015(.din(n858), .dout(n4200));
    jand g1016(.dinb(n12032), .dina(n4172), .dout(n4204));
    jand g1017(.dinb(n11972), .dina(n4204), .dout(n4208));
    jor g1018(.dinb(n11921), .dina(n4208), .dout(n4212));
    jand g1019(.dinb(n11873), .dina(n4212), .dout(n4216));
    jor g1020(.dinb(n11810), .dina(n4216), .dout(n4220));
    jor g1021(.dinb(n11747), .dina(n4220), .dout(n4224));
    jand g1022(.dinb(n11666), .dina(n4224), .dout(n4228));
    jxor g1023(.dinb(n9053), .dina(n4228), .dout(n4232));
    jand g1024(.dinb(n14350), .dina(n3391), .dout(n4236));
    jnot g1025(.din(n4236), .dout(n4239));
    jand g1026(.dinb(n13324), .dina(n4172), .dout(n4243));
    jnot g1027(.din(n4243), .dout(n4246));
    jand g1028(.dinb(n13258), .dina(n4246), .dout(n4250));
    jand g1029(.dinb(n10417), .dina(n4250), .dout(n4254));
    jor g1030(.dinb(n14212), .dina(n4254), .dout(n4258));
    jxor g1031(.dinb(n13942), .dina(n4258), .dout(n4262));
    jor g1032(.dinb(n13864), .dina(n4250), .dout(n4266));
    jnot g1033(.din(n4254), .dout(n4269));
    jor g1034(.dinb(n14128), .dina(n4269), .dout(n4273));
    jand g1035(.dinb(n8807), .dina(n4273), .dout(n4277));
    jnot g1036(.din(n960), .dout(n4280));
    jor g1037(.dinb(n13387), .dina(n4280), .dout(n4284));
    jand g1038(.dinb(n13474), .dina(n1753), .dout(n4288));
    jor g1039(.dinb(n8867), .dina(n4288), .dout(n4292));
    jxor g1040(.dinb(n13744), .dina(n4292), .dout(n4296));
    jand g1041(.dinb(n13540), .dina(n1753), .dout(n4300));
    jor g1042(.dinb(n13402), .dina(n4300), .dout(n4304));
    jxor g1043(.dinb(n13639), .dina(n4304), .dout(n4308));
    jor g1044(.dinb(n662), .dina(n11569), .dout(n4312));
    jor g1045(.dinb(n12352), .dina(n1781), .dout(n4316));
    jand g1046(.dinb(n11500), .dina(n4316), .dout(n4320));
    jxor g1047(.dinb(n11122), .dina(n4320), .dout(n4324));
    jand g1048(.dinb(n12670), .dina(n678), .dout(n4328));
    jor g1049(.dinb(n654), .dina(n11483), .dout(n4332));
    jor g1050(.dinb(n12448), .dina(n1781), .dout(n4336));
    jand g1051(.dinb(n11401), .dina(n4336), .dout(n4340));
    jxor g1052(.dinb(n15370), .dina(n4340), .dout(n4344));
    jnot g1053(.din(n577), .dout(n4347));
    jnot g1054(.din(n607), .dout(n4350));
    jnot g1055(.din(n592), .dout(n4353));
    jor g1056(.dinb(n9053), .dina(n4228), .dout(n4357));
    jand g1057(.dinb(n12262), .dina(n4357), .dout(n4361));
    jor g1058(.dinb(n9146), .dina(n4361), .dout(n4365));
    jand g1059(.dinb(n12529), .dina(n4365), .dout(n4369));
    jxor g1060(.dinb(n8966), .dina(n4369), .dout(G333));
    jxor g1061(.dinb(n9146), .dina(n4361), .dout(n4377));
    jor g1062(.dinb(n9439), .dina(n4111), .dout(n4381));
    jor g1063(.dinb(n344), .dina(n392), .dout(n4385));
    jor g1064(.dinb(n368), .dina(n416), .dout(n4389));
    jor g1065(.dinb(n3625), .dina(n9197), .dout(n4393));
    jor g1066(.dinb(n9176), .dina(n4393), .dout(n4397));
    jor g1067(.dinb(n9152), .dina(n4397), .dout(n4401));
    jxor g1068(.dinb(n15178), .dina(n1773), .dout(n4405));
    jand g1069(.dinb(n14683), .dina(n1765), .dout(n4409));
    jor g1070(.dinb(n14521), .dina(n4409), .dout(n4413));
    jxor g1071(.dinb(n14974), .dina(n4413), .dout(n4417));
    jand g1072(.dinb(n14851), .dina(n3373), .dout(n4421));
    jnot g1073(.din(n4421), .dout(n4424));
    jor g1074(.dinb(n14596), .dina(n1765), .dout(n4428));
    jand g1075(.dinb(n10621), .dina(n4428), .dout(n4432));
    jxor g1076(.dinb(n14863), .dina(n4432), .dout(n4436));
    jxor g1077(.dinb(n14758), .dina(n1765), .dout(n4440));
    jxor g1078(.dinb(n16921), .dina(n1677), .dout(n4444));
    jor g1079(.dinb(n9901), .dina(n1800), .dout(n4448));
    jor g1080(.dinb(n1789), .dina(n9802), .dout(n4452));
    jand g1081(.dinb(n9800), .dina(n4452), .dout(n4456));
    jxor g1082(.dinb(n9913), .dina(n4456), .dout(G422));
    jxor g1083(.dinb(n10121), .dina(n1789), .dout(n4464));
    jand g1084(.dinb(n16741), .dina(n1677), .dout(n4468));
    jor g1085(.dinb(n16447), .dina(n4468), .dout(n4472));
    jxor g1086(.dinb(n17101), .dina(n4472), .dout(n4476));
    jnot g1087(.din(n1288), .dout(n4479));
    jnot g1088(.din(n1178), .dout(n4482));
    jnot g1089(.din(n1244), .dout(n4485));
    jnot g1090(.din(n1284), .dout(n4488));
    jand g1091(.dinb(n4485), .dina(n15725), .dout(n4492));
    jor g1092(.dinb(n16606), .dina(n4492), .dout(n4496));
    jand g1093(.dinb(n15716), .dina(n4496), .dout(n4500));
    jnot g1094(.din(n1252), .dout(n4503));
    jand g1095(.dinb(n10142), .dina(n4136), .dout(n4507));
    jor g1096(.dinb(n15679), .dina(n4507), .dout(n4511));
    jxor g1097(.dinb(n15727), .dina(n4511), .dout(n4515));
    jand g1098(.dinb(n16882), .dina(n1677), .dout(n4519));
    jor g1099(.dinb(n16507), .dina(n4519), .dout(n4523));
    jxor g1100(.dinb(n16780), .dina(n4523), .dout(n4527));
    jand g1101(.dinb(n16963), .dina(n1677), .dout(n4531));
    jor g1102(.dinb(n16540), .dina(n4531), .dout(n4535));
    jxor g1103(.dinb(n17029), .dina(n4535), .dout(n4539));
    jxor g1104(.dinb(n16003), .dina(n1017), .dout(n4543));
    jxor g1105(.dinb(n1745), .dina(n15931), .dout(n4547));
    jand g1106(.dinb(n4156), .dina(n16132), .dout(n4551));
    jxor g1107(.dinb(n12097), .dina(n4551), .dout(n4555));
    jxor g1108(.dinb(n1069), .dina(n1091), .dout(n4559));
    jor g1109(.dinb(n1689), .dina(n10190), .dout(n4563));
    jand g1110(.dinb(n4152), .dina(n4563), .dout(n4567));
    jxor g1111(.dinb(n16298), .dina(n1065), .dout(n4571));
    jxor g1112(.dinb(n1685), .dina(n15862), .dout(n4575));
    jxor g1113(.dinb(n717), .dina(n732), .dout(n4579));
    jor g1114(.dinb(n14674), .dina(n4424), .dout(n4583));
    jnot g1115(.din(n800), .dout(n4586));
    jor g1116(.dinb(n10696), .dina(n4586), .dout(n4590));
    jand g1117(.dinb(n10619), .dina(n4590), .dout(n4594));
    jxor g1118(.dinb(n10712), .dina(n4594), .dout(n4598));
    jxor g1119(.dinb(n14947), .dina(n808), .dout(n4602));
    jxor g1120(.dinb(n4598), .dina(n10616), .dout(n4606));
    jand g1121(.dinb(n4212), .dina(n10613), .dout(n4610));
    jxor g1122(.dinb(n747), .dina(n792), .dout(n4614));
    jnot g1123(.din(n4614), .dout(n4617));
    jand g1124(.dinb(n4586), .dina(n10556), .dout(n4621));
    jor g1125(.dinb(n788), .dina(n762), .dout(n4625));
    jand g1126(.dinb(n4614), .dina(n4625), .dout(n4629));
    jor g1127(.dinb(n4621), .dina(n10553), .dout(n4633));
    jxor g1128(.dinb(n812), .dina(n10712), .dout(n4637));
    jxor g1129(.dinb(n10547), .dina(n4637), .dout(n4641));
    jand g1130(.dinb(n1765), .dina(n10544), .dout(n4645));
    jor g1131(.dinb(n4610), .dina(n4645), .dout(n4649));
    jand g1132(.dinb(n10414), .dina(n990), .dout(n4653));
    jor g1133(.dinb(n14311), .dina(n4653), .dout(n4657));
    jxor g1134(.dinb(n908), .dina(n927), .dout(n4661));
    jand g1135(.dinb(n983), .dina(n10405), .dout(n4665));
    jnot g1136(.din(n4661), .dout(n4668));
    jand g1137(.dinb(n990), .dina(n10391), .dout(n4672));
    jor g1138(.dinb(n10379), .dina(n4672), .dout(n4676));
    jnot g1139(.din(n923), .dout(n4679));
    jand g1140(.dinb(n13627), .dina(n4679), .dout(n4683));
    jnot g1141(.din(n4683), .dout(n4686));
    jor g1142(.dinb(n13396), .dina(n4686), .dout(n4690));
    jor g1143(.dinb(n949), .dina(n4683), .dout(n4694));
    jand g1144(.dinb(n4690), .dina(n10373), .dout(n4698));
    jxor g1145(.dinb(n14035), .dina(n4698), .dout(n4702));
    jxor g1146(.dinb(n4676), .dina(n10370), .dout(n4706));
    jxor g1147(.dinb(n10361), .dina(n4706), .dout(n4710));
    jand g1148(.dinb(n1753), .dina(n10358), .dout(n4714));
    jand g1149(.dinb(n10487), .dina(n986), .dout(n4718));
    jor g1150(.dinb(n14293), .dina(n4718), .dout(n4722));
    jor g1151(.dinb(n968), .dina(n953), .dout(n4726));
    jand g1152(.dinb(n960), .dina(n10319), .dout(n4730));
    jxor g1153(.dinb(n14026), .dina(n4730), .dout(n4734));
    jxor g1154(.dinb(n983), .dina(n4734), .dout(n4738));
    jxor g1155(.dinb(n10393), .dina(n4738), .dout(n4742));
    jxor g1156(.dinb(n4722), .dina(n10316), .dout(n4746));
    jand g1157(.dinb(n4172), .dina(n10313), .dout(n4750));
    jor g1158(.dinb(n4714), .dina(n4750), .dout(n4754));
    jxor g1159(.dinb(n866), .dina(n889), .dout(n4758));
    jxor g1160(.dinb(n4754), .dina(n10268), .dout(n4762));
    jxor g1161(.dinb(n4649), .dina(n10196), .dout(n4766));
    jxor g1162(.dinb(n577), .dina(n682), .dout(n4770));
    jxor g1163(.dinb(n12682), .dina(n662), .dout(n4774));
    jand g1164(.dinb(n12350), .dina(n647), .dout(n4778));
    jand g1165(.dinb(n12640), .dina(n654), .dout(n4782));
    jor g1166(.dinb(n12260), .dina(n4782), .dout(n4786));
    jnot g1167(.din(n611), .dout(n4789));
    jand g1168(.dinb(n12526), .dina(n4789), .dout(n4793));
    jxor g1169(.dinb(n607), .dina(n674), .dout(n4797));
    jxor g1170(.dinb(n4793), .dina(n12230), .dout(n4801));
    jxor g1171(.dinb(n4786), .dina(n12224), .dout(n4805));
    jxor g1172(.dinb(n4774), .dina(n4805), .dout(n4809));
    jor g1173(.dinb(n1781), .dina(n12215), .dout(n4813));
    jor g1174(.dinb(n12664), .dina(n588), .dout(n4817));
    jor g1175(.dinb(n12634), .dina(n603), .dout(n4821));
    jand g1176(.dinb(n4817), .dina(n4821), .dout(n4825));
    jnot g1177(.din(n4817), .dout(n4828));
    jand g1178(.dinb(n11498), .dina(n4793), .dout(n4832));
    jor g1179(.dinb(n11492), .dina(n4832), .dout(n4836));
    jxor g1180(.dinb(n537), .dina(n607), .dout(n4840));
    jxor g1181(.dinb(n4332), .dina(n11399), .dout(n4844));
    jxor g1182(.dinb(n11384), .dina(n4844), .dout(n4848));
    jxor g1183(.dinb(n12232), .dina(n4848), .dout(n4852));
    jxor g1184(.dinb(n11567), .dina(n4852), .dout(n4856));
    jor g1185(.dinb(n4228), .dina(n11378), .dout(n4860));
    jand g1186(.dinb(n4813), .dina(n4860), .dout(n4864));
    jxor g1187(.dinb(n11318), .dina(n4864), .dout(n4868));
    jand g1188(.dinb(n11095), .dina(n481), .dout(n4872));
    jnot g1189(.din(n489), .dout(n4875));
    jor g1190(.dinb(n4872), .dina(n4875), .dout(n4879));
    jnot g1191(.din(n4872), .dout(n4882));
    jor g1192(.dinb(n11071), .dina(n4882), .dout(n4886));
    jand g1193(.dinb(n11063), .dina(n4886), .dout(n4890));
    jand g1194(.dinb(n670), .dina(n11060), .dout(n4894));
    jnot g1195(.din(n670), .dout(n4897));
    jand g1196(.dinb(n11023), .dina(n1800), .dout(n4901));
    jor g1197(.dinb(n4901), .dina(n11065), .dout(n4905));
    jor g1198(.dinb(n11083), .dina(n507), .dout(n4909));
    jand g1199(.dinb(n4905), .dina(n4909), .dout(n4913));
    jand g1200(.dinb(n4897), .dina(n11018), .dout(n4917));
    jor g1201(.dinb(n10991), .dina(n4917), .dout(n4921));
    jor g1202(.dinb(n1781), .dina(n10988), .dout(n4925));
    jnot g1203(.din(n694), .dout(n4928));
    jand g1204(.dinb(n10916), .dina(n4917), .dout(n4932));
    jand g1205(.dinb(n698), .dina(n11035), .dout(n4936));
    jor g1206(.dinb(n4932), .dina(n10769), .dout(n4940));
    jor g1207(.dinb(n4228), .dina(n10766), .dout(n4944));
    jand g1208(.dinb(n4925), .dina(n4944), .dout(n4948));
    jxor g1209(.dinb(n4868), .dina(n10715), .dout(n4952));
    jor g1210(.dinb(n16126), .dina(n1727), .dout(n4956));
    jand g1211(.dinb(n1734), .dina(n16124), .dout(n4960));
    jor g1212(.dinb(n16330), .dina(n4960), .dout(n4964));
    jxor g1213(.dinb(n4123), .dina(n15992), .dout(n4968));
    jxor g1214(.dinb(n16075), .dina(n4968), .dout(n4972));
    jxor g1215(.dinb(n4964), .dina(n15929), .dout(n4976));
    jand g1216(.dinb(n4126), .dina(n15920), .dout(n4980));
    jand g1217(.dinb(n16664), .dina(n4980), .dout(n4984));
    jand g1218(.dinb(n1091), .dina(n4571), .dout(n4988));
    jnot g1219(.din(n4988), .dout(n4991));
    jor g1220(.dinb(n16328), .dina(n4991), .dout(n4995));
    jor g1221(.dinb(n4960), .dina(n15850), .dout(n4999));
    jand g1222(.dinb(n15848), .dina(n4999), .dout(n5003));
    jxor g1223(.dinb(n1050), .dina(n1069), .dout(n5007));
    jxor g1224(.dinb(n4968), .dina(n15839), .dout(n5011));
    jxor g1225(.dinb(n5003), .dina(n15836), .dout(n5015));
    jor g1226(.dinb(n1268), .dina(n16666), .dout(n5019));
    jand g1227(.dinb(n15817), .dina(n5019), .dout(n5023));
    jor g1228(.dinb(n4984), .dina(n15815), .dout(n5027));
    jand g1229(.dinb(n1677), .dina(n5027), .dout(n5031));
    jand g1230(.dinb(n1268), .dina(n15824), .dout(n5035));
    jor g1231(.dinb(n4980), .dina(n15776), .dout(n5039));
    jand g1232(.dinb(n4136), .dina(n15773), .dout(n5043));
    jor g1233(.dinb(n5031), .dina(n5043), .dout(n5047));
    jxor g1234(.dinb(n4479), .dina(n16777), .dout(n5051));
    jnot g1235(.din(n1232), .dout(n5054));
    jand g1236(.dinb(n17017), .dina(n5054), .dout(n5058));
    jnot g1237(.din(n5058), .dout(n5061));
    jand g1238(.dinb(n16591), .dina(n5061), .dout(n5065));
    jand g1239(.dinb(n16594), .dina(n5058), .dout(n5069));
    jor g1240(.dinb(n5065), .dina(n15677), .dout(n5073));
    jxor g1241(.dinb(n17152), .dina(n5073), .dout(n5077));
    jxor g1242(.dinb(n4500), .dina(n15674), .dout(n5081));
    jnot g1243(.din(n1260), .dout(n5084));
    jxor g1244(.dinb(n1276), .dina(n1280), .dout(n5088));
    jnot g1245(.din(n5088), .dout(n5091));
    jor g1246(.dinb(n5084), .dina(n15623), .dout(n5095));
    jor g1247(.dinb(n1260), .dina(n15646), .dout(n5099));
    jor g1248(.dinb(n16720), .dina(n5099), .dout(n5103));
    jand g1249(.dinb(n5095), .dina(n5103), .dout(n5107));
    jxor g1250(.dinb(n15602), .dina(n5107), .dout(n5111));
    jor g1251(.dinb(n4136), .dina(n15596), .dout(n5115));
    jxor g1252(.dinb(n1260), .dina(n15625), .dout(n5119));
    jnot g1253(.din(n1240), .dout(n5122));
    jor g1254(.dinb(n1207), .dina(n1236), .dout(n5126));
    jand g1255(.dinb(n5122), .dina(n15590), .dout(n5130));
    jxor g1256(.dinb(n17143), .dina(n5130), .dout(n5134));
    jxor g1257(.dinb(n1252), .dina(n5134), .dout(n5138));
    jxor g1258(.dinb(n5119), .dina(n15581), .dout(n5142));
    jor g1259(.dinb(n1677), .dina(n15575), .dout(n5146));
    jand g1260(.dinb(n5115), .dina(n5146), .dout(n5150));
    jxor g1261(.dinb(n15563), .dina(n5150), .dout(n5154));
    jxor g1262(.dinb(n15521), .dina(n5154), .dout(n5158));
    jxor g1263(.dinb(n3354), .dina(n18010), .dout(n5162));
    jxor g1264(.dinb(n18155), .dina(n5162), .dout(n5166));
    jand g1265(.dinb(n17990), .dina(n1434), .dout(n5170));
    jand g1266(.dinb(n17929), .dina(n1431), .dout(n5174));
    jor g1267(.dinb(n5170), .dina(n17927), .dout(n5178));
    jxor g1268(.dinb(n17924), .dina(n5178), .dout(n5182));
    jand g1269(.dinb(n3294), .dina(n17918), .dout(n5186));
    jand g1270(.dinb(n18322), .dina(n5186), .dout(n5190));
    jnot g1271(.din(n1367), .dout(n5193));
    jand g1272(.dinb(n18175), .dina(n5193), .dout(n5197));
    jand g1273(.dinb(n5197), .dina(n3347), .dout(n5201));
    jand g1274(.dinb(n1419), .dina(n1423), .dout(n5205));
    jor g1275(.dinb(n5201), .dina(n17513), .dout(n5209));
    jor g1276(.dinb(n17587), .dina(n5209), .dout(n5213));
    jxor g1277(.dinb(n1352), .dina(n3265), .dout(n5217));
    jxor g1278(.dinb(n5213), .dina(n17510), .dout(n5221));
    jxor g1279(.dinb(n1446), .dina(n17501), .dout(n5225));
    jand g1280(.dinb(n1653), .dina(n17494), .dout(n5229));
    jor g1281(.dinb(n17764), .dina(n5229), .dout(n5233));
    jor g1282(.dinb(n17492), .dina(n5233), .dout(n5237));
    jand g1283(.dinb(n1649), .dina(n17498), .dout(n5241));
    jor g1284(.dinb(n5186), .dina(n5241), .dout(n5245));
    jor g1285(.dinb(n17803), .dina(n5245), .dout(n5249));
    jand g1286(.dinb(n5237), .dina(n17489), .dout(n5253));
    jxor g1287(.dinb(n470), .dina(n18347), .dout(n5257));
    jxor g1288(.dinb(n3198), .dina(n5257), .dout(n5261));
    jxor g1289(.dinb(n3206), .dina(n17471), .dout(n5265));
    jnot g1290(.din(n5265), .dout(n5268));
    jxor g1291(.dinb(n18389), .dina(n1471), .dout(n5272));
    jxor g1292(.dinb(n1641), .dina(n17459), .dout(n5276));
    jor g1293(.dinb(n17444), .dina(n5276), .dout(n5280));
    jnot g1294(.din(n5276), .dout(n5283));
    jor g1295(.dinb(n17461), .dina(n5283), .dout(n5287));
    jand g1296(.dinb(n17761), .dina(n5287), .dout(n5291));
    jand g1297(.dinb(n17441), .dina(n5291), .dout(n5295));
    jand g1298(.dinb(n18379), .dina(n3198), .dout(n5299));
    jand g1299(.dinb(n466), .dina(n1602), .dout(n5303));
    jor g1300(.dinb(n5299), .dina(n17435), .dout(n5307));
    jxor g1301(.dinb(n18526), .dina(n5307), .dout(n5311));
    jxor g1302(.dinb(n3210), .dina(n5311), .dout(n5315));
    jnot g1303(.din(n5315), .dout(n5318));
    jnot g1304(.din(n1543), .dout(n5321));
    jand g1305(.dinb(n17423), .dina(n3286), .dout(n5325));
    jxor g1306(.dinb(n17473), .dina(n5325), .dout(n5329));
    jnot g1307(.din(n5329), .dout(n5332));
    jor g1308(.dinb(n17420), .dina(n5332), .dout(n5336));
    jor g1309(.dinb(n17425), .dina(n5329), .dout(n5340));
    jand g1310(.dinb(n17875), .dina(n5340), .dout(n5344));
    jand g1311(.dinb(n5336), .dina(n5344), .dout(n5348));
    jor g1312(.dinb(n5295), .dina(n5348), .dout(n5352));
    jxor g1313(.dinb(n1490), .dina(n1509), .dout(n5356));
    jxor g1314(.dinb(n5352), .dina(n17414), .dout(n5360));
    jxor g1315(.dinb(n5253), .dina(n5360), .dout(n5364));
    jdff g1316(.din(G1), .dout(n5367));
    jdff g1317(.din(G1), .dout(n5370));
    jdff g1318(.din(G1459), .dout(n5373));
    jdff g1319(.din(G1469), .dout(n5376));
    jdff g1320(.din(G1480), .dout(n5379));
    jdff g1321(.din(G1486), .dout(n5382));
    jdff g1322(.din(G1492), .dout(n5385));
    jdff g1323(.din(G1496), .dout(n5388));
    jdff g1324(.din(G2208), .dout(n5391));
    jdff g1325(.din(G2218), .dout(n5394));
    jdff g1326(.din(G2224), .dout(n5397));
    jdff g1327(.din(G2230), .dout(n5400));
    jdff g1328(.din(G2236), .dout(n5403));
    jdff g1329(.din(G2239), .dout(n5406));
    jdff g1330(.din(G2247), .dout(n5409));
    jdff g1331(.din(G2253), .dout(n5412));
    jdff g1332(.din(G2256), .dout(n5415));
    jdff g1333(.din(G3698), .dout(n5418));
    jdff g1334(.din(G3701), .dout(n5421));
    jdff g1335(.din(G3705), .dout(n5424));
    jdff g1336(.din(G3711), .dout(n5427));
    jdff g1337(.din(G3717), .dout(n5430));
    jdff g1338(.din(G3723), .dout(n5433));
    jdff g1339(.din(G3729), .dout(n5436));
    jdff g1340(.din(G3737), .dout(n5439));
    jdff g1341(.din(G3743), .dout(n5442));
    jdff g1342(.din(G3749), .dout(n5445));
    jdff g1343(.din(G4393), .dout(n5448));
    jdff g1344(.din(G4400), .dout(n5451));
    jdff g1345(.din(G4405), .dout(n5454));
    jdff g1346(.din(G4410), .dout(n5457));
    jdff g1347(.din(G4415), .dout(n5460));
    jdff g1348(.din(G4420), .dout(n5463));
    jdff g1349(.din(G4427), .dout(n5466));
    jdff g1350(.din(G4432), .dout(n5469));
    jdff g1351(.din(G4437), .dout(n5472));
    jdff g1352(.din(G1462), .dout(n5475));
    jdff g1353(.din(G2211), .dout(n5478));
    jdff g1354(.din(G4394), .dout(n5481));
    jdff g1355(.din(G1), .dout(n5484));
    jdff g1356(.din(G106), .dout(n5487));
    jnot g1357(.din(G15), .dout(n5490));
    jor g1358(.dinb(n7858), .dina(n419), .dout(n5494));
    jnot g1359(.din(G15), .dout(n5497));
    jor g1360(.dinb(n7865), .dina(n433), .dout(n5501));
    jdff g1361(.din(G1), .dout(n5504));
    jand g1362(.dinb(n8444), .dina(n3169), .dout(n5508));
    jor g1363(.dinb(n1797), .dina(n9695), .dout(G270));
    jand g1364(.dinb(n8444), .dina(n3169), .dout(n5516));
    jor g1365(.dinb(n1797), .dina(n9695), .dout(G276));
    jor g1366(.dinb(n1797), .dina(n9695), .dout(G273));
    jxor g1367(.dinb(n9907), .dina(n4456), .dout(G469));
    jxor g1368(.dinb(n10121), .dina(n1789), .dout(n5532));
    jdff dff_A_qp69ew1k3_0(.din(n26827), .dout(G399));
    jdff dff_A_Tm1UH8M69_0(.din(n26824), .dout(n26827));
    jdff dff_A_2MSuZMVk5_0(.din(n26821), .dout(n26824));
    jdff dff_A_9ZIm3fD33_0(.din(n26818), .dout(n26821));
    jdff dff_A_Jt6aMDQ94_0(.din(n26815), .dout(n26818));
    jdff dff_A_1vJFTEEo4_0(.din(n26812), .dout(n26815));
    jdff dff_A_EnSTdf7g6_0(.din(n26809), .dout(n26812));
    jdff dff_A_j3c1f5To7_0(.din(n26806), .dout(n26809));
    jdff dff_A_utWrhI8o3_0(.din(n26803), .dout(n26806));
    jdff dff_A_LVLxvjpj1_0(.din(n26800), .dout(n26803));
    jdff dff_A_eVXWxF4r8_0(.din(n26797), .dout(n26800));
    jdff dff_A_sNl1j9sY2_0(.din(n26794), .dout(n26797));
    jdff dff_A_UqQwMQpd0_0(.din(n26791), .dout(n26794));
    jdff dff_A_QS29gxdM5_0(.din(n26788), .dout(n26791));
    jdff dff_A_eOFAMxXJ6_0(.din(n26785), .dout(n26788));
    jdff dff_A_PSY8VEdo3_0(.din(n26782), .dout(n26785));
    jdff dff_A_iDNk4g734_0(.din(n26779), .dout(n26782));
    jdff dff_A_4ctQpcnd2_0(.din(n26776), .dout(n26779));
    jdff dff_A_faxxTd5s3_0(.din(n26773), .dout(n26776));
    jdff dff_A_xrM9NinU7_0(.din(n26770), .dout(n26773));
    jdff dff_A_SZHKifOh5_2(.din(n5364), .dout(n26770));
    jdff dff_A_iBbCuLEp4_0(.din(n26764), .dout(G370));
    jdff dff_A_04DFZzRO4_0(.din(n26761), .dout(n26764));
    jdff dff_A_5HZDyfup5_0(.din(n26758), .dout(n26761));
    jdff dff_A_caS97pzf2_0(.din(n26755), .dout(n26758));
    jdff dff_A_HCOqsXlx4_0(.din(n26752), .dout(n26755));
    jdff dff_A_patlHC8c3_0(.din(n26749), .dout(n26752));
    jdff dff_A_bi5YO1QB7_0(.din(n26746), .dout(n26749));
    jdff dff_A_eRzlU6yE5_0(.din(n26743), .dout(n26746));
    jdff dff_A_NpIy8QxP0_0(.din(n26740), .dout(n26743));
    jdff dff_A_QBrIUpQs0_0(.din(n26737), .dout(n26740));
    jdff dff_A_BgCpmlhe9_0(.din(n26734), .dout(n26737));
    jdff dff_A_OozD2UhM1_0(.din(n26731), .dout(n26734));
    jdff dff_A_pom0h5kE6_0(.din(n26728), .dout(n26731));
    jdff dff_A_Yo2qFoKU9_0(.din(n26725), .dout(n26728));
    jdff dff_A_Jqd4xWpb1_0(.din(n26722), .dout(n26725));
    jdff dff_A_o8QafsO16_0(.din(n26719), .dout(n26722));
    jdff dff_A_oM4MwWtI5_2(.din(n5158), .dout(n26719));
    jdff dff_A_3AVLPWfs6_2(.din(n4952), .dout(G338));
    jdff dff_A_ocJ5WiQt8_0(.din(n26710), .dout(G321));
    jdff dff_A_XbNGlsgT6_0(.din(n26707), .dout(n26710));
    jdff dff_A_syg62Qgg5_0(.din(n26704), .dout(n26707));
    jdff dff_A_63iv9Lgt4_0(.din(n26701), .dout(n26704));
    jdff dff_A_mIhX1E8q9_0(.din(n26698), .dout(n26701));
    jdff dff_A_kjGGFBjr5_2(.din(n4766), .dout(n26698));
    jdff dff_A_C2zreAzv5_0(.din(n26692), .dout(G356));
    jdff dff_A_G4LGUiy17_0(.din(n26689), .dout(n26692));
    jdff dff_A_CMGYIz2W0_0(.din(n26686), .dout(n26689));
    jdff dff_A_iFGbiI5M0_0(.din(n26683), .dout(n26686));
    jdff dff_A_557gcgzR0_0(.din(n26680), .dout(n26683));
    jdff dff_A_bK9inClz4_0(.din(n26677), .dout(n26680));
    jdff dff_A_UpoGRkq93_0(.din(n26674), .dout(n26677));
    jdff dff_A_zGpUNtdD2_0(.din(n26671), .dout(n26674));
    jdff dff_A_icCUAyOh3_0(.din(n26668), .dout(n26671));
    jdff dff_A_asSJdhsN3_0(.din(n26665), .dout(n26668));
    jdff dff_A_oaqnHzPb4_0(.din(n26662), .dout(n26665));
    jdff dff_A_ZTTy8cRz9_0(.din(n26659), .dout(n26662));
    jdff dff_A_LAsdIJpO2_0(.din(n26656), .dout(n26659));
    jdff dff_A_6oZDhHqT0_0(.din(n26653), .dout(n26656));
    jdff dff_A_Hwn6ljTY8_0(.din(n26650), .dout(n26653));
    jdff dff_A_hLvOlyGW9_0(.din(n26647), .dout(n26650));
    jdff dff_A_tdsQ6rES9_0(.din(n26644), .dout(n26647));
    jdff dff_A_fSEwKRmD3_2(.din(n4575), .dout(n26644));
    jdff dff_A_wX30sGNI9_0(.din(n26638), .dout(G353));
    jdff dff_A_RrFeEEwF1_0(.din(n26635), .dout(n26638));
    jdff dff_A_o2PvDGlQ1_0(.din(n26632), .dout(n26635));
    jdff dff_A_8Wg1UBbA2_0(.din(n26629), .dout(n26632));
    jdff dff_A_klBuYOAh1_0(.din(n26626), .dout(n26629));
    jdff dff_A_3WBHduyB5_0(.din(n26623), .dout(n26626));
    jdff dff_A_z4uEjMGn0_0(.din(n26620), .dout(n26623));
    jdff dff_A_HwJX9iCr2_0(.din(n26617), .dout(n26620));
    jdff dff_A_wnqCkNDS2_0(.din(n26614), .dout(n26617));
    jdff dff_A_pl2xJzib4_0(.din(n26611), .dout(n26614));
    jdff dff_A_WQGQdT9K8_0(.din(n26608), .dout(n26611));
    jdff dff_A_nB9rpTsv6_0(.din(n26605), .dout(n26608));
    jdff dff_A_xGtgUL8o3_0(.din(n26602), .dout(n26605));
    jdff dff_A_JEcEXyYJ5_0(.din(n26599), .dout(n26602));
    jdff dff_A_hFSAKiyw3_0(.din(n26596), .dout(n26599));
    jdff dff_A_lnookEJx5_2(.din(n4567), .dout(n26596));
    jdff dff_A_Dtcr2t8E9_0(.din(n26590), .dout(G350));
    jdff dff_A_ko2P7GjQ4_0(.din(n26587), .dout(n26590));
    jdff dff_A_lCZJMyYO7_0(.din(n26584), .dout(n26587));
    jdff dff_A_fYKJRhen9_0(.din(n26581), .dout(n26584));
    jdff dff_A_hvHvB2zE9_0(.din(n26578), .dout(n26581));
    jdff dff_A_eZlrCZqr9_0(.din(n26575), .dout(n26578));
    jdff dff_A_Xy2JumR71_0(.din(n26572), .dout(n26575));
    jdff dff_A_tVFX3nj97_0(.din(n26569), .dout(n26572));
    jdff dff_A_SdAU7V2Q1_0(.din(n26566), .dout(n26569));
    jdff dff_A_BiAC9qPC4_0(.din(n26563), .dout(n26566));
    jdff dff_A_cd9govl93_0(.din(n26560), .dout(n26563));
    jdff dff_A_XZea749D9_0(.din(n26557), .dout(n26560));
    jdff dff_A_Y3duYJiR3_0(.din(n26554), .dout(n26557));
    jdff dff_A_RRVhlcbP2_2(.din(n4555), .dout(n26554));
    jdff dff_A_77ssRZCb2_0(.din(n26548), .dout(G347));
    jdff dff_A_6D9PtInS1_0(.din(n26545), .dout(n26548));
    jdff dff_A_v1AWzzSo9_0(.din(n26542), .dout(n26545));
    jdff dff_A_cigL26PG5_0(.din(n26539), .dout(n26542));
    jdff dff_A_npOvNuPR5_0(.din(n26536), .dout(n26539));
    jdff dff_A_Muat5UCv8_0(.din(n26533), .dout(n26536));
    jdff dff_A_n7JEDQ8V9_0(.din(n26530), .dout(n26533));
    jdff dff_A_I58el1FW9_0(.din(n26527), .dout(n26530));
    jdff dff_A_F4x6EZGn9_0(.din(n26524), .dout(n26527));
    jdff dff_A_joX9QhWi4_0(.din(n26521), .dout(n26524));
    jdff dff_A_64PeerYV0_0(.din(n26518), .dout(n26521));
    jdff dff_A_zjSrlHje7_0(.din(n26515), .dout(n26518));
    jdff dff_A_QExPo0Wj9_2(.din(n4547), .dout(n26515));
    jdff dff_A_f6zmQDRH2_0(.din(n26509), .dout(G368));
    jdff dff_A_tggbj35D0_0(.din(n26506), .dout(n26509));
    jdff dff_A_npPxXng34_0(.din(n26503), .dout(n26506));
    jdff dff_A_FsiRgk9F2_0(.din(n26500), .dout(n26503));
    jdff dff_A_KZnSz4oG9_0(.din(n26497), .dout(n26500));
    jdff dff_A_jphJM6sA5_0(.din(n26494), .dout(n26497));
    jdff dff_A_Uk1kWr2b3_0(.din(n26491), .dout(n26494));
    jdff dff_A_06QDEm150_0(.din(n26488), .dout(n26491));
    jdff dff_A_eHYOdJuD0_0(.din(n26485), .dout(n26488));
    jdff dff_A_LgSqa9uP7_0(.din(n26482), .dout(n26485));
    jdff dff_A_adO26Uvs3_0(.din(n26479), .dout(n26482));
    jdff dff_A_eQUQsWTy3_0(.din(n26476), .dout(n26479));
    jdff dff_A_iWlaiOJf0_0(.din(n26473), .dout(n26476));
    jdff dff_A_akKupNvi7_0(.din(n26470), .dout(n26473));
    jdff dff_A_CDe5Np1a1_0(.din(n26467), .dout(n26470));
    jdff dff_A_WhsXkAvs8_0(.din(n26464), .dout(n26467));
    jdff dff_A_WBGl0WpB8_0(.din(n26461), .dout(n26464));
    jdff dff_A_7pKYbPVy4_2(.din(n4539), .dout(n26461));
    jdff dff_A_6NQCOJIc2_0(.din(n26455), .dout(G365));
    jdff dff_A_Li7dGMDe5_0(.din(n26452), .dout(n26455));
    jdff dff_A_aOSDakV86_0(.din(n26449), .dout(n26452));
    jdff dff_A_YGpfq2Jd9_0(.din(n26446), .dout(n26449));
    jdff dff_A_5VkYQ8El0_0(.din(n26443), .dout(n26446));
    jdff dff_A_fQgQo2ye7_0(.din(n26440), .dout(n26443));
    jdff dff_A_7PP1sbCB6_0(.din(n26437), .dout(n26440));
    jdff dff_A_2UzDimiZ9_0(.din(n26434), .dout(n26437));
    jdff dff_A_TCxdCZHY1_0(.din(n26431), .dout(n26434));
    jdff dff_A_YzK76lN63_0(.din(n26428), .dout(n26431));
    jdff dff_A_72h9EVtj2_0(.din(n26425), .dout(n26428));
    jdff dff_A_xWT3jQs29_0(.din(n26422), .dout(n26425));
    jdff dff_A_uCogFCmT3_0(.din(n26419), .dout(n26422));
    jdff dff_A_YOBdtfMA2_0(.din(n26416), .dout(n26419));
    jdff dff_A_o0UazIW82_0(.din(n26413), .dout(n26416));
    jdff dff_A_6YO4tzXl6_0(.din(n26410), .dout(n26413));
    jdff dff_A_AZzDua9b3_0(.din(n26407), .dout(n26410));
    jdff dff_A_aqO8jZ6A6_2(.din(n4527), .dout(n26407));
    jdff dff_A_UPZ5k5Xb9_0(.din(n26401), .dout(G362));
    jdff dff_A_OhYKUvWI1_0(.din(n26398), .dout(n26401));
    jdff dff_A_0RTInmma9_0(.din(n26395), .dout(n26398));
    jdff dff_A_8yoyiDDb7_0(.din(n26392), .dout(n26395));
    jdff dff_A_ZqUBEiYz9_0(.din(n26389), .dout(n26392));
    jdff dff_A_CpHfLnY25_0(.din(n26386), .dout(n26389));
    jdff dff_A_XyI0mOA96_0(.din(n26383), .dout(n26386));
    jdff dff_A_6L7oKnnq6_0(.din(n26380), .dout(n26383));
    jdff dff_A_zTHqLjhk6_0(.din(n26377), .dout(n26380));
    jdff dff_A_13cYZlMt2_0(.din(n26374), .dout(n26377));
    jdff dff_A_DBJGPkYD5_0(.din(n26371), .dout(n26374));
    jdff dff_A_j7MCRLo46_0(.din(n26368), .dout(n26371));
    jdff dff_A_Wp5C6Slw5_0(.din(n26365), .dout(n26368));
    jdff dff_A_LcOUrM4m3_0(.din(n26362), .dout(n26365));
    jdff dff_A_Vc4je3797_0(.din(n26359), .dout(n26362));
    jdff dff_A_GCu76aiM2_0(.din(n26356), .dout(n26359));
    jdff dff_A_gTN6iNlU9_0(.din(n26353), .dout(n26356));
    jdff dff_A_A4XOy4fh6_2(.din(n4515), .dout(n26353));
    jdff dff_A_6wJk8jyM6_0(.din(n26347), .dout(G359));
    jdff dff_A_fy6XihzP7_0(.din(n26344), .dout(n26347));
    jdff dff_A_JWsvIb9c8_0(.din(n26341), .dout(n26344));
    jdff dff_A_Bmfi1Pd85_0(.din(n26338), .dout(n26341));
    jdff dff_A_MAHEbFBd1_0(.din(n26335), .dout(n26338));
    jdff dff_A_4k3rMu2f9_0(.din(n26332), .dout(n26335));
    jdff dff_A_n9IPYTyO1_0(.din(n26329), .dout(n26332));
    jdff dff_A_zK39wwoO4_0(.din(n26326), .dout(n26329));
    jdff dff_A_SRISsozN2_0(.din(n26323), .dout(n26326));
    jdff dff_A_Ng5PWTK74_0(.din(n26320), .dout(n26323));
    jdff dff_A_nvN9YVzL6_0(.din(n26317), .dout(n26320));
    jdff dff_A_VfdZ5erP6_0(.din(n26314), .dout(n26317));
    jdff dff_A_X3BxciBC4_0(.din(n26311), .dout(n26314));
    jdff dff_A_Lca0kmFz9_0(.din(n26308), .dout(n26311));
    jdff dff_A_tPHdV3u70_0(.din(n26305), .dout(n26308));
    jdff dff_A_bEIjtywn2_0(.din(n26302), .dout(n26305));
    jdff dff_A_JXazmYKP2_0(.din(n26299), .dout(n26302));
    jdff dff_A_gjRLzgIm3_2(.din(n4476), .dout(n26299));
    jdff dff_A_kyRgxR5R7_0(.din(n26293), .dout(G471));
    jdff dff_A_TNQyhMuw3_2(.din(n5532), .dout(n26293));
    jdff dff_A_HlcRKYcW8_0(.din(n26287), .dout(G419));
    jdff dff_A_5xWKymr18_2(.din(n4464), .dout(n26287));
    jdff dff_A_Izr64Mtx0_0(.din(n26281), .dout(G344));
    jdff dff_A_zg3xNFJl1_0(.din(n26278), .dout(n26281));
    jdff dff_A_z4pndscK5_0(.din(n26275), .dout(n26278));
    jdff dff_A_kBA3nHEg5_0(.din(n26272), .dout(n26275));
    jdff dff_A_oEcxtlaH3_0(.din(n26269), .dout(n26272));
    jdff dff_A_Cn0gG3nw8_0(.din(n26266), .dout(n26269));
    jdff dff_A_RmMNSInv4_0(.din(n26263), .dout(n26266));
    jdff dff_A_H4nuQuD29_0(.din(n26260), .dout(n26263));
    jdff dff_A_QgfBEcCl0_0(.din(n26257), .dout(n26260));
    jdff dff_A_sxzLpbNr9_0(.din(n26254), .dout(n26257));
    jdff dff_A_lNXZEEmI6_0(.din(n26251), .dout(n26254));
    jdff dff_A_LNfNVx5v9_0(.din(n26248), .dout(n26251));
    jdff dff_A_xNhO77ex5_0(.din(n26245), .dout(n26248));
    jdff dff_A_7TrXXuFg1_0(.din(n26242), .dout(n26245));
    jdff dff_A_hikfPZ1u3_0(.din(n26239), .dout(n26242));
    jdff dff_A_TRwoNDg73_0(.din(n26236), .dout(n26239));
    jdff dff_A_Tx2EeQEC5_0(.din(n26233), .dout(n26236));
    jdff dff_A_KVuEHkkb2_0(.din(n26230), .dout(n26233));
    jdff dff_A_yGWClJHQ3_0(.din(n26227), .dout(n26230));
    jdff dff_A_NpO6pto17_2(.din(n4444), .dout(n26227));
    jdff dff_A_ZNa2zk2F9_0(.din(n26221), .dout(G307));
    jdff dff_A_Enrz0vw03_0(.din(n26218), .dout(n26221));
    jdff dff_A_pN6rLBLl2_0(.din(n26215), .dout(n26218));
    jdff dff_A_OPuVijkx7_0(.din(n26212), .dout(n26215));
    jdff dff_A_1mvlSIxx1_0(.din(n26209), .dout(n26212));
    jdff dff_A_t1a9Lv1z5_0(.din(n26206), .dout(n26209));
    jdff dff_A_8RsmyaiI5_0(.din(n26203), .dout(n26206));
    jdff dff_A_xlZ8L1W07_2(.din(n4440), .dout(n26203));
    jdff dff_A_UD0mHw0Y8_0(.din(n26197), .dout(G304));
    jdff dff_A_1ORmC1Rr9_0(.din(n26194), .dout(n26197));
    jdff dff_A_33B314zn1_0(.din(n26191), .dout(n26194));
    jdff dff_A_62ACiwer7_0(.din(n26188), .dout(n26191));
    jdff dff_A_B9hm0S602_0(.din(n26185), .dout(n26188));
    jdff dff_A_5ZJ7pWXu5_2(.din(n4436), .dout(n26185));
    jdff dff_A_7s1UEE4E9_0(.din(n26179), .dout(G301));
    jdff dff_A_EQdiu7Rs7_0(.din(n26176), .dout(n26179));
    jdff dff_A_wgWE2OIF4_0(.din(n26173), .dout(n26176));
    jdff dff_A_nyc2roSQ8_0(.din(n26170), .dout(n26173));
    jdff dff_A_WL258vLB9_0(.din(n26167), .dout(n26170));
    jdff dff_A_Zf5g3S756_2(.din(n4417), .dout(n26167));
    jdff dff_A_5HB4DTtw9_0(.din(n26161), .dout(G298));
    jdff dff_A_u2QOunfA3_0(.din(n26158), .dout(n26161));
    jdff dff_A_0o1hTSuY3_0(.din(n26155), .dout(n26158));
    jdff dff_A_9k1mbw330_0(.din(n26152), .dout(n26155));
    jdff dff_A_5FuhfzB66_0(.din(n26149), .dout(n26152));
    jdff dff_A_66Kxv2s37_2(.din(n4405), .dout(n26149));
    jdff dff_A_7S3hWtba7_0(.din(n26143), .dout(G418));
    jdff dff_A_EvNvKbhg4_0(.din(n26140), .dout(n26143));
    jdff dff_A_cO5F2zJo7_0(.din(n26137), .dout(n26140));
    jdff dff_A_ja4VovS83_0(.din(n26134), .dout(n26137));
    jdff dff_A_skz1TVNd4_0(.din(n26131), .dout(n26134));
    jdff dff_A_MexYlLuv6_0(.din(n26128), .dout(n26131));
    jdff dff_A_Ztvpptee8_0(.din(n26125), .dout(n26128));
    jdff dff_A_2dEyfsHJ7_0(.din(n26122), .dout(n26125));
    jdff dff_A_Yu8avxCL4_0(.din(n26119), .dout(n26122));
    jdff dff_A_vrTN3nrh9_0(.din(n26116), .dout(n26119));
    jdff dff_A_OJOU4HGP3_0(.din(n26113), .dout(n26116));
    jdff dff_A_uN8TCNXs0_0(.din(n26110), .dout(n26113));
    jdff dff_A_ZD0wqzCR0_0(.din(n26107), .dout(n26110));
    jdff dff_A_5Faf9DTs9_0(.din(n26104), .dout(n26107));
    jdff dff_A_MSlCcuJr7_0(.din(n26101), .dout(n26104));
    jdff dff_A_sPJrOy6n7_0(.din(n26098), .dout(n26101));
    jdff dff_A_tVu4vRE77_0(.din(n26095), .dout(n26098));
    jdff dff_A_fkKoHX4M6_0(.din(n26092), .dout(n26095));
    jdff dff_A_0MxlA2ET8_0(.din(n26089), .dout(n26092));
    jdff dff_A_WfdH0IHe9_0(.din(n26086), .dout(n26089));
    jdff dff_A_RwTLNT8w2_0(.din(n26083), .dout(n26086));
    jdff dff_A_4bsi1gVk1_0(.din(n26080), .dout(n26083));
    jdff dff_A_e8tpRDF93_0(.din(n26077), .dout(n26080));
    jdff dff_A_XmzPJ8Z65_0(.din(n26074), .dout(n26077));
    jdff dff_A_DpK9MJgg0_2(.din(n4401), .dout(n26074));
    jdff dff_A_8FT8dgJl5_0(.din(n26068), .dout(G336));
    jdff dff_A_LuZMZecF1_2(.din(n4377), .dout(n26068));
    jdff dff_A_WDRkfbAT3_0(.din(n26062), .dout(G330));
    jdff dff_A_4qm3SZjK2_2(.din(n4344), .dout(n26062));
    jdff dff_A_Phw1tJnA6_0(.din(n26056), .dout(G327));
    jdff dff_A_F5JBNVEW3_2(.din(n4324), .dout(n26056));
    jdff dff_A_eOEDl1WL5_0(.din(n26050), .dout(G319));
    jdff dff_A_q2DaGNrb1_0(.din(n26047), .dout(n26050));
    jdff dff_A_CdS7RY2u4_0(.din(n26044), .dout(n26047));
    jdff dff_A_xgQlfr3r4_0(.din(n26041), .dout(n26044));
    jdff dff_A_LUjSBSBl2_0(.din(n26038), .dout(n26041));
    jdff dff_A_1rPRtXIg7_0(.din(n26035), .dout(n26038));
    jdff dff_A_5Zm3OgNo7_0(.din(n26032), .dout(n26035));
    jdff dff_A_7KFerPuq5_0(.din(n26029), .dout(n26032));
    jdff dff_A_3fDqDu737_2(.din(n4308), .dout(n26029));
    jdff dff_A_eTQMF5Qy7_0(.din(n26023), .dout(G316));
    jdff dff_A_Qp3H3yc01_0(.din(n26020), .dout(n26023));
    jdff dff_A_QndRye4D9_0(.din(n26017), .dout(n26020));
    jdff dff_A_QhnLDcRO1_0(.din(n26014), .dout(n26017));
    jdff dff_A_uimQMgSQ5_0(.din(n26011), .dout(n26014));
    jdff dff_A_cNEKW8gF0_0(.din(n26008), .dout(n26011));
    jdff dff_A_sNDuGX0S8_0(.din(n26005), .dout(n26008));
    jdff dff_A_wMVTovFG7_0(.din(n26002), .dout(n26005));
    jdff dff_A_90iJhh3S3_2(.din(n4296), .dout(n26002));
    jdff dff_A_f2y4bC435_0(.din(n25996), .dout(G313));
    jdff dff_A_TiLs4IDp0_0(.din(n25993), .dout(n25996));
    jdff dff_A_MBiSDkNg6_0(.din(n25990), .dout(n25993));
    jdff dff_A_R6jWaAUu3_0(.din(n25987), .dout(n25990));
    jdff dff_A_HM3MKpQL8_2(.din(n4277), .dout(n25987));
    jdff dff_A_8lN7DabA1_0(.din(n25981), .dout(G310));
    jdff dff_A_XSrtizU08_0(.din(n25978), .dout(n25981));
    jdff dff_A_UGyAlJ6Y0_0(.din(n25975), .dout(n25978));
    jdff dff_A_HvPMqq5t9_0(.din(n25972), .dout(n25975));
    jdff dff_A_pyMSuIju5_0(.din(n25969), .dout(n25972));
    jdff dff_A_gwDlvvGS8_2(.din(n4262), .dout(n25969));
    jdff dff_A_w4VHtvYt5_0(.din(n25963), .dout(G252));
    jdff dff_A_ASJ4J5SQ2_0(.din(n25960), .dout(n25963));
    jdff dff_A_5sNSkv1N1_0(.din(n25957), .dout(n25960));
    jdff dff_A_8qXkLzQl9_0(.din(n25954), .dout(n25957));
    jdff dff_A_l5gMOBei4_0(.din(n25951), .dout(n25954));
    jdff dff_A_1tJXCDZH5_0(.din(n25948), .dout(n25951));
    jdff dff_A_FIEAXlDu9_0(.din(n25945), .dout(n25948));
    jdff dff_A_mGLUpW3V3_0(.din(n25942), .dout(n25945));
    jdff dff_A_PYLW6zl73_0(.din(n25939), .dout(n25942));
    jdff dff_A_8S4rUr0x5_0(.din(n25936), .dout(n25939));
    jdff dff_A_n5Qvx2W22_0(.din(n25933), .dout(n25936));
    jdff dff_A_KhQG3VGM0_0(.din(n25930), .dout(n25933));
    jdff dff_A_spldhYxi7_0(.din(n25927), .dout(n25930));
    jdff dff_A_VLrYmf5Z1_0(.din(n25924), .dout(n25927));
    jdff dff_A_uDtlWOCu5_0(.din(n25921), .dout(n25924));
    jdff dff_A_1XTG5deb9_0(.din(n25918), .dout(n25921));
    jdff dff_A_xPDRx4bs8_0(.din(n25915), .dout(n25918));
    jdff dff_A_pzKquxwd5_0(.din(n25912), .dout(n25915));
    jdff dff_A_KsYWvMPz2_0(.din(n25909), .dout(n25912));
    jdff dff_A_ugdaHuIq3_0(.din(n25906), .dout(n25909));
    jdff dff_A_qDtSjULd9_1(.din(n3053), .dout(n25906));
    jdff dff_A_742KAgvO1_0(.din(n25900), .dout(G324));
    jdff dff_A_YVfZ5NnC0_0(.din(n25897), .dout(n25900));
    jdff dff_A_V6rEcdFt9_0(.din(n25894), .dout(n25897));
    jdff dff_A_zrcXL1rl7_2(.din(n4232), .dout(n25894));
    jdff dff_A_X39QseWh6_0(.din(n25888), .dout(G295));
    jdff dff_A_led1xBmg1_0(.din(n25885), .dout(n25888));
    jdff dff_A_FjvKrP1L7_0(.din(n25882), .dout(n25885));
    jdff dff_A_4o1FDuoc5_0(.din(n25879), .dout(n25882));
    jdff dff_A_fycggT6y2_0(.din(n25876), .dout(n25879));
    jdff dff_A_NZNHqxuW7_0(.din(n25873), .dout(n25876));
    jdff dff_A_vfccntIk7_0(.din(n25870), .dout(n25873));
    jdff dff_A_i6rV34jg1_0(.din(n25867), .dout(n25870));
    jdff dff_A_36wbyAAn1_0(.din(n25864), .dout(n25867));
    jdff dff_A_aK0GLROY2_0(.din(n25861), .dout(n25864));
    jdff dff_A_xfiKRwPP3_2(.din(n4176), .dout(n25861));
    jdff dff_A_ediNWG1J7_0(.din(n25855), .dout(G249));
    jdff dff_A_P125zpNw4_0(.din(n25852), .dout(n25855));
    jdff dff_A_2krjyInS3_0(.din(n25849), .dout(n25852));
    jdff dff_A_QK4jZoz99_0(.din(n25846), .dout(n25849));
    jdff dff_A_SFTo6Cfo7_0(.din(n25843), .dout(n25846));
    jdff dff_A_yUIXDO435_0(.din(n25840), .dout(n25843));
    jdff dff_A_SdsYbdir9_0(.din(n25837), .dout(n25840));
    jdff dff_A_01A7bkPs6_0(.din(n25834), .dout(n25837));
    jdff dff_A_ZyDKHbNT6_0(.din(n25831), .dout(n25834));
    jdff dff_A_OVLSzOC91_0(.din(n25828), .dout(n25831));
    jdff dff_A_ILSvZBEJ4_2(.din(n5516), .dout(n25828));
    jdff dff_A_ku4bgICf8_0(.din(n25822), .dout(G416));
    jdff dff_A_IMH9stej5_0(.din(n25819), .dout(n25822));
    jdff dff_A_mG0QgLiw8_0(.din(n25816), .dout(n25819));
    jdff dff_A_kBitKUpS4_0(.din(n25813), .dout(n25816));
    jdff dff_A_y5ZnVpJd4_0(.din(n25810), .dout(n25813));
    jdff dff_A_M23WeA3w0_0(.din(n25807), .dout(n25810));
    jdff dff_A_1P1c9G1b8_0(.din(n25804), .dout(n25807));
    jdff dff_A_XtDUCDlA7_0(.din(n25801), .dout(n25804));
    jdff dff_A_BG3MG6e71_0(.din(n25798), .dout(n25801));
    jdff dff_A_u4bbuj2R2_0(.din(n25795), .dout(n25798));
    jdff dff_A_386anNwP6_0(.din(n25792), .dout(n25795));
    jdff dff_A_slxDaHWE6_0(.din(n25789), .dout(n25792));
    jdff dff_A_Sr5tra2P7_0(.din(n25786), .dout(n25789));
    jdff dff_A_6AmY8qAZ4_0(.din(n25783), .dout(n25786));
    jdff dff_A_qBBnIvzr8_0(.din(n25780), .dout(n25783));
    jdff dff_A_S74WIrSZ4_0(.din(n25777), .dout(n25780));
    jdff dff_A_2LBlAj0V3_0(.din(n25774), .dout(n25777));
    jdff dff_A_MKOz98611_0(.din(n25771), .dout(n25774));
    jdff dff_A_uhyNS0uH7_0(.din(n25768), .dout(n25771));
    jdff dff_A_GhGmbBTX1_0(.din(n25765), .dout(n25768));
    jdff dff_A_NTX6bz143_0(.din(n25762), .dout(n25765));
    jdff dff_A_zO4s8VNy2_0(.din(n25759), .dout(n25762));
    jdff dff_A_pPRppIca7_0(.din(n25756), .dout(n25759));
    jdff dff_A_R7QPpjgf2_0(.din(n25753), .dout(n25756));
    jdff dff_A_al6xBKIX6_0(.din(n25750), .dout(n25753));
    jdff dff_A_czG8FT767_0(.din(n25747), .dout(n25750));
    jdff dff_A_shnOCCR11_0(.din(n25744), .dout(n25747));
    jdff dff_A_7ljZlT9V9_0(.din(n25741), .dout(n25744));
    jdff dff_A_qkkR41lL2_1(.din(n4111), .dout(n25741));
    jdff dff_A_fl9wfYSL3_0(.din(n25735), .dout(G414));
    jdff dff_A_wwd0LvTI7_0(.din(n25732), .dout(n25735));
    jdff dff_A_3jAjF1Gz6_0(.din(n25729), .dout(n25732));
    jdff dff_A_pC563uJb1_0(.din(n25726), .dout(n25729));
    jdff dff_A_Udi0OLKP8_0(.din(n25723), .dout(n25726));
    jdff dff_A_52KrNaZP3_0(.din(n25720), .dout(n25723));
    jdff dff_A_2uwE9oa72_0(.din(n25717), .dout(n25720));
    jdff dff_A_aYNRGjsY9_0(.din(n25714), .dout(n25717));
    jdff dff_A_E7nqzzLD2_0(.din(n25711), .dout(n25714));
    jdff dff_A_A5zHOWMX2_0(.din(n25708), .dout(n25711));
    jdff dff_A_btY6XhyT9_0(.din(n25705), .dout(n25708));
    jdff dff_A_h0ewkhsh3_0(.din(n25702), .dout(n25705));
    jdff dff_A_5LoUhNRd9_0(.din(n25699), .dout(n25702));
    jdff dff_A_hT4K5FmC9_0(.din(n25696), .dout(n25699));
    jdff dff_A_5BU2K0yv5_0(.din(n25693), .dout(n25696));
    jdff dff_A_nExZUtR06_0(.din(n25690), .dout(n25693));
    jdff dff_A_gR1jdJvZ9_0(.din(n25687), .dout(n25690));
    jdff dff_A_L0UlO98V6_0(.din(n25684), .dout(n25687));
    jdff dff_A_Kz6Ru4PS6_0(.din(n25681), .dout(n25684));
    jdff dff_A_YhKGf7wL9_0(.din(n25678), .dout(n25681));
    jdff dff_A_VycTajte5_0(.din(n25675), .dout(n25678));
    jdff dff_A_WBawVD2a9_0(.din(n25672), .dout(n25675));
    jdff dff_A_hEk6ocyy6_0(.din(n25669), .dout(n25672));
    jdff dff_A_WCLfFFzk4_0(.din(n25666), .dout(n25669));
    jdff dff_A_Of6vaUcI3_0(.din(n25663), .dout(n25666));
    jdff dff_A_t4blgWWg3_0(.din(n25660), .dout(n25663));
    jdff dff_A_X2cIBIdp3_0(.din(n25657), .dout(n25660));
    jdff dff_A_quCktKZK7_0(.din(n25654), .dout(n25657));
    jdff dff_A_lvMnoDQb4_0(.din(n25651), .dout(n25654));
    jdff dff_A_I8w0B8AP8_1(.din(n3866), .dout(n25651));
    jdff dff_A_vfpGiafr1_0(.din(n25645), .dout(G412));
    jdff dff_A_KY6aIAwW6_0(.din(n25642), .dout(n25645));
    jdff dff_A_kgzbzXtT2_0(.din(n25639), .dout(n25642));
    jdff dff_A_cplgJl6L5_0(.din(n25636), .dout(n25639));
    jdff dff_A_H9WEcLuX7_0(.din(n25633), .dout(n25636));
    jdff dff_A_r2wZF0K61_0(.din(n25630), .dout(n25633));
    jdff dff_A_GfGoUerw9_0(.din(n25627), .dout(n25630));
    jdff dff_A_o6KxQzLL7_0(.din(n25624), .dout(n25627));
    jdff dff_A_UUfhRLOj5_0(.din(n25621), .dout(n25624));
    jdff dff_A_NzGWomL06_0(.din(n25618), .dout(n25621));
    jdff dff_A_Ll27CUwy3_0(.din(n25615), .dout(n25618));
    jdff dff_A_XfMIXKrl8_0(.din(n25612), .dout(n25615));
    jdff dff_A_V0skxr0F7_0(.din(n25609), .dout(n25612));
    jdff dff_A_GugBEpix2_0(.din(n25606), .dout(n25609));
    jdff dff_A_FsukPbtM5_0(.din(n25603), .dout(n25606));
    jdff dff_A_7WFgkYER7_0(.din(n25600), .dout(n25603));
    jdff dff_A_iBsDKZqG6_0(.din(n25597), .dout(n25600));
    jdff dff_A_CBiBBm4n5_0(.din(n25594), .dout(n25597));
    jdff dff_A_0YXCL5Ik2_0(.din(n25591), .dout(n25594));
    jdff dff_A_Mt9v6H714_0(.din(n25588), .dout(n25591));
    jdff dff_A_vY0xZFyl9_0(.din(n25585), .dout(n25588));
    jdff dff_A_ZTRW8m1r2_0(.din(n25582), .dout(n25585));
    jdff dff_A_nBEVTmQl0_0(.din(n25579), .dout(n25582));
    jdff dff_A_xjFsUMIC1_0(.din(n25576), .dout(n25579));
    jdff dff_A_9BdYvwWZ5_0(.din(n25573), .dout(n25576));
    jdff dff_A_H4LIQZcz0_0(.din(n25570), .dout(n25573));
    jdff dff_A_JygE6xV54_0(.din(n25567), .dout(n25570));
    jdff dff_A_bjP8Gnko9_1(.din(n3625), .dout(n25567));
    jdff dff_A_i6ELr4Gm8_0(.din(n25561), .dout(G385));
    jdff dff_A_lvIBfCit0_0(.din(n25558), .dout(n25561));
    jdff dff_A_DH8muabI7_0(.din(n25555), .dout(n25558));
    jdff dff_A_VEG1LvX42_0(.din(n25552), .dout(n25555));
    jdff dff_A_yxYhDQmB1_0(.din(n25549), .dout(n25552));
    jdff dff_A_fbVCFjhV8_0(.din(n25546), .dout(n25549));
    jdff dff_A_moKsCxe35_0(.din(n25543), .dout(n25546));
    jdff dff_A_vHHhn0rE8_0(.din(n25540), .dout(n25543));
    jdff dff_A_bQjDTPrO9_0(.din(n25537), .dout(n25540));
    jdff dff_A_qgijVHmm8_0(.din(n25534), .dout(n25537));
    jdff dff_A_lI7zYVwi0_0(.din(n25531), .dout(n25534));
    jdff dff_A_vxK1JuXe5_0(.din(n25528), .dout(n25531));
    jdff dff_A_OJvHaqSg2_0(.din(n25525), .dout(n25528));
    jdff dff_A_HGnJh86x2_0(.din(n25522), .dout(n25525));
    jdff dff_A_xVQkVIfh8_0(.din(n25519), .dout(n25522));
    jdff dff_A_GAteg4uW2_0(.din(n25516), .dout(n25519));
    jdff dff_A_wTQvmoWW0_0(.din(n25513), .dout(n25516));
    jdff dff_A_MIY5zbxi1_0(.din(n25510), .dout(n25513));
    jdff dff_A_0cWbSjBm6_0(.din(n25507), .dout(n25510));
    jdff dff_A_7kaOGsd84_0(.din(n25504), .dout(n25507));
    jdff dff_A_Dj3tBW0L8_0(.din(n25501), .dout(n25504));
    jdff dff_A_mn0c5MFP5_0(.din(n25498), .dout(n25501));
    jdff dff_A_iZEIChW01_0(.din(n25495), .dout(n25498));
    jdff dff_A_QdpmjzBx0_2(.din(n3370), .dout(n25495));
    jdff dff_A_fyaugnMa2_0(.din(n25489), .dout(G382));
    jdff dff_A_JZvHAGLw5_0(.din(n25486), .dout(n25489));
    jdff dff_A_C1hkKMUJ3_0(.din(n25483), .dout(n25486));
    jdff dff_A_3ICkKOD14_0(.din(n25480), .dout(n25483));
    jdff dff_A_5o1x4bdg3_0(.din(n25477), .dout(n25480));
    jdff dff_A_a5EPy4Eo6_0(.din(n25474), .dout(n25477));
    jdff dff_A_y2sS8QCS1_0(.din(n25471), .dout(n25474));
    jdff dff_A_JP63ReqE8_0(.din(n25468), .dout(n25471));
    jdff dff_A_QN6sim7e1_0(.din(n25465), .dout(n25468));
    jdff dff_A_mvSPDdfY6_0(.din(n25462), .dout(n25465));
    jdff dff_A_PSRTnObD1_0(.din(n25459), .dout(n25462));
    jdff dff_A_uEyHgZvI9_0(.din(n25456), .dout(n25459));
    jdff dff_A_9ipDSy589_0(.din(n25453), .dout(n25456));
    jdff dff_A_k94ta9Te0_0(.din(n25450), .dout(n25453));
    jdff dff_A_4noCiurx9_0(.din(n25447), .dout(n25450));
    jdff dff_A_rcRwI3k86_0(.din(n25444), .dout(n25447));
    jdff dff_A_gSSZ0jMX7_0(.din(n25441), .dout(n25444));
    jdff dff_A_lUNlwOxw3_0(.din(n25438), .dout(n25441));
    jdff dff_A_nIGbZKFp1_0(.din(n25435), .dout(n25438));
    jdff dff_A_akV4xtHz7_0(.din(n25432), .dout(n25435));
    jdff dff_A_81labtvY2_0(.din(n25429), .dout(n25432));
    jdff dff_A_8hS9m2Y73_2(.din(n3366), .dout(n25429));
    jdff dff_A_Pvsn6F9o5_0(.din(n25423), .dout(G379));
    jdff dff_A_CtZh37QI7_0(.din(n25420), .dout(n25423));
    jdff dff_A_TU3bReNd5_0(.din(n25417), .dout(n25420));
    jdff dff_A_DmhPxgal5_0(.din(n25414), .dout(n25417));
    jdff dff_A_cuTUdWVQ7_0(.din(n25411), .dout(n25414));
    jdff dff_A_QZu0Vnbb5_0(.din(n25408), .dout(n25411));
    jdff dff_A_xz1zoii98_0(.din(n25405), .dout(n25408));
    jdff dff_A_TttgXi3p2_0(.din(n25402), .dout(n25405));
    jdff dff_A_npwC4EFi4_0(.din(n25399), .dout(n25402));
    jdff dff_A_ASQRqqgS8_0(.din(n25396), .dout(n25399));
    jdff dff_A_g5xImQhC7_0(.din(n25393), .dout(n25396));
    jdff dff_A_Utf0xcYh7_0(.din(n25390), .dout(n25393));
    jdff dff_A_cPHzPg2Q5_0(.din(n25387), .dout(n25390));
    jdff dff_A_AdfZZQkV9_0(.din(n25384), .dout(n25387));
    jdff dff_A_3EwZXQr04_0(.din(n25381), .dout(n25384));
    jdff dff_A_oRVU4bwl0_0(.din(n25378), .dout(n25381));
    jdff dff_A_Dn1W2jZo5_0(.din(n25375), .dout(n25378));
    jdff dff_A_lvtQbmGm9_0(.din(n25372), .dout(n25375));
    jdff dff_A_DExDC5NA7_0(.din(n25369), .dout(n25372));
    jdff dff_A_ENMl7Ul43_0(.din(n25366), .dout(n25369));
    jdff dff_A_hJfgijJH7_0(.din(n25363), .dout(n25366));
    jdff dff_A_1iQksQaM0_2(.din(n3341), .dout(n25363));
    jdff dff_A_YIe0BZdp2_0(.din(n25357), .dout(G376));
    jdff dff_A_w14rmFCR8_0(.din(n25354), .dout(n25357));
    jdff dff_A_xMdH4bvC6_0(.din(n25351), .dout(n25354));
    jdff dff_A_bnz3u5M11_0(.din(n25348), .dout(n25351));
    jdff dff_A_3Rh7J9tu3_0(.din(n25345), .dout(n25348));
    jdff dff_A_5JsqUKxw8_0(.din(n25342), .dout(n25345));
    jdff dff_A_fJTZhBr26_0(.din(n25339), .dout(n25342));
    jdff dff_A_dSTkFMBC4_0(.din(n25336), .dout(n25339));
    jdff dff_A_mYyUNWY12_0(.din(n25333), .dout(n25336));
    jdff dff_A_pOGcSKCK9_0(.din(n25330), .dout(n25333));
    jdff dff_A_Iu7M7jYm4_0(.din(n25327), .dout(n25330));
    jdff dff_A_QZwkynxl6_0(.din(n25324), .dout(n25327));
    jdff dff_A_QmAp1mWZ8_0(.din(n25321), .dout(n25324));
    jdff dff_A_rov2lSPR2_0(.din(n25318), .dout(n25321));
    jdff dff_A_qzv6Kkxg3_0(.din(n25315), .dout(n25318));
    jdff dff_A_Jr2FxMJX9_0(.din(n25312), .dout(n25315));
    jdff dff_A_joi2S2HD0_0(.din(n25309), .dout(n25312));
    jdff dff_A_Jnwu2Yhf4_0(.din(n25306), .dout(n25309));
    jdff dff_A_9mPUOZh00_0(.din(n25303), .dout(n25306));
    jdff dff_A_SGZG573Y4_2(.din(n3329), .dout(n25303));
    jdff dff_A_yAlJLw6x9_0(.din(n25297), .dout(G397));
    jdff dff_A_TQEAN2BS3_0(.din(n25294), .dout(n25297));
    jdff dff_A_FFcBnvFW4_0(.din(n25291), .dout(n25294));
    jdff dff_A_nTjrgZKe8_0(.din(n25288), .dout(n25291));
    jdff dff_A_RLqxLHBO8_0(.din(n25285), .dout(n25288));
    jdff dff_A_LcmR00Rp7_0(.din(n25282), .dout(n25285));
    jdff dff_A_uVOIUjPU9_0(.din(n25279), .dout(n25282));
    jdff dff_A_hBdyxDej5_0(.din(n25276), .dout(n25279));
    jdff dff_A_hvLRLS7Y4_0(.din(n25273), .dout(n25276));
    jdff dff_A_1DEqSVSh8_0(.din(n25270), .dout(n25273));
    jdff dff_A_PmPFXRkm5_0(.din(n25267), .dout(n25270));
    jdff dff_A_TLWD8j7q8_0(.din(n25264), .dout(n25267));
    jdff dff_A_P5bnf5xA4_0(.din(n25261), .dout(n25264));
    jdff dff_A_Qa4lUHWV6_0(.din(n25258), .dout(n25261));
    jdff dff_A_ismxpB1d4_0(.din(n25255), .dout(n25258));
    jdff dff_A_LGhfym0w3_0(.din(n25252), .dout(n25255));
    jdff dff_A_P6AVwomB9_0(.din(n25249), .dout(n25252));
    jdff dff_A_sBgo36vb4_0(.din(n25246), .dout(n25249));
    jdff dff_A_fD6h7s5w5_0(.din(n25243), .dout(n25246));
    jdff dff_A_XrCT66DO4_0(.din(n25240), .dout(n25243));
    jdff dff_A_Oqd4VR4j8_0(.din(n25237), .dout(n25240));
    jdff dff_A_HaUUTyqT3_0(.din(n25234), .dout(n25237));
    jdff dff_A_Z5vwzN8A5_0(.din(n25231), .dout(n25234));
    jdff dff_A_E6RaSHGq9_0(.din(n25228), .dout(n25231));
    jdff dff_A_4vpgJdKb8_0(.din(n25225), .dout(n25228));
    jdff dff_A_GlJUvyaM9_0(.din(n25222), .dout(n25225));
    jdff dff_A_1TmbwBDk6_0(.din(n25219), .dout(n25222));
    jdff dff_A_sfGrFQKw2_0(.din(n25216), .dout(n25219));
    jdff dff_A_XKV3xiQI6_0(.din(n25213), .dout(n25216));
    jdff dff_A_prcnguFT9_0(.din(n25210), .dout(n25213));
    jdff dff_A_JmJfu1Jx3_2(.din(n3261), .dout(n25210));
    jdff dff_A_tL4B5Qt22_0(.din(n25204), .dout(G394));
    jdff dff_A_IQkVbZHN5_0(.din(n25201), .dout(n25204));
    jdff dff_A_ZVuNEt8t7_0(.din(n25198), .dout(n25201));
    jdff dff_A_CreCEGnX4_0(.din(n25195), .dout(n25198));
    jdff dff_A_2z1wE9Tr7_0(.din(n25192), .dout(n25195));
    jdff dff_A_zKOEIkDr2_0(.din(n25189), .dout(n25192));
    jdff dff_A_s3R6TkFj3_0(.din(n25186), .dout(n25189));
    jdff dff_A_0Ee2ZB4q3_0(.din(n25183), .dout(n25186));
    jdff dff_A_948eRYST5_0(.din(n25180), .dout(n25183));
    jdff dff_A_6fJC1h071_0(.din(n25177), .dout(n25180));
    jdff dff_A_Efgp4oSm6_0(.din(n25174), .dout(n25177));
    jdff dff_A_8ePTkFr49_0(.din(n25171), .dout(n25174));
    jdff dff_A_nyu2S2zC0_0(.din(n25168), .dout(n25171));
    jdff dff_A_046HKjwD5_0(.din(n25165), .dout(n25168));
    jdff dff_A_YKfG7xbx4_0(.din(n25162), .dout(n25165));
    jdff dff_A_OPysQK8j9_0(.din(n25159), .dout(n25162));
    jdff dff_A_OGfNbo279_0(.din(n25156), .dout(n25159));
    jdff dff_A_pQXfIaEc7_0(.din(n25153), .dout(n25156));
    jdff dff_A_h6KY3otM4_0(.din(n25150), .dout(n25153));
    jdff dff_A_w9WqPI5b7_0(.din(n25147), .dout(n25150));
    jdff dff_A_GeuJQvZH1_0(.din(n25144), .dout(n25147));
    jdff dff_A_KoOHLsFp7_0(.din(n25141), .dout(n25144));
    jdff dff_A_eepxyCLY5_0(.din(n25138), .dout(n25141));
    jdff dff_A_IwHeJo6u7_0(.din(n25135), .dout(n25138));
    jdff dff_A_PgLsNzlD8_0(.din(n25132), .dout(n25135));
    jdff dff_A_v6cvdGue5_0(.din(n25129), .dout(n25132));
    jdff dff_A_U29S5hfu4_0(.din(n25126), .dout(n25129));
    jdff dff_A_yKwTG61T1_0(.din(n25123), .dout(n25126));
    jdff dff_A_VEC37Kb97_0(.din(n25120), .dout(n25123));
    jdff dff_A_lPzfP2la9_2(.din(n3253), .dout(n25120));
    jdff dff_A_MLSieQRb5_0(.din(n25114), .dout(G391));
    jdff dff_A_rPh0qnnX6_0(.din(n25111), .dout(n25114));
    jdff dff_A_fjmmPZfX7_0(.din(n25108), .dout(n25111));
    jdff dff_A_I33HmPdM2_0(.din(n25105), .dout(n25108));
    jdff dff_A_rXriJFTA6_0(.din(n25102), .dout(n25105));
    jdff dff_A_ylmtbOf76_0(.din(n25099), .dout(n25102));
    jdff dff_A_F6GX7V5k7_0(.din(n25096), .dout(n25099));
    jdff dff_A_8gjEDqU79_0(.din(n25093), .dout(n25096));
    jdff dff_A_AldomAwp8_0(.din(n25090), .dout(n25093));
    jdff dff_A_UDnVxWWn3_0(.din(n25087), .dout(n25090));
    jdff dff_A_oz2mxFWJ6_0(.din(n25084), .dout(n25087));
    jdff dff_A_sdWqi4Go1_0(.din(n25081), .dout(n25084));
    jdff dff_A_l7Pn9xLV6_0(.din(n25078), .dout(n25081));
    jdff dff_A_QpadcRY80_0(.din(n25075), .dout(n25078));
    jdff dff_A_I7WGF6fh4_0(.din(n25072), .dout(n25075));
    jdff dff_A_7Pro7rEs1_0(.din(n25069), .dout(n25072));
    jdff dff_A_7vvA95Gx0_0(.din(n25066), .dout(n25069));
    jdff dff_A_D56M6mj31_0(.din(n25063), .dout(n25066));
    jdff dff_A_DV8plbpk4_0(.din(n25060), .dout(n25063));
    jdff dff_A_63ytucfX7_0(.din(n25057), .dout(n25060));
    jdff dff_A_6y2qeYlc9_0(.din(n25054), .dout(n25057));
    jdff dff_A_Ag0jBzgQ0_0(.din(n25051), .dout(n25054));
    jdff dff_A_oYmIiRKo1_0(.din(n25048), .dout(n25051));
    jdff dff_A_Ra96J6TQ9_0(.din(n25045), .dout(n25048));
    jdff dff_A_uWUq719U4_0(.din(n25042), .dout(n25045));
    jdff dff_A_x8uJ3uU14_0(.din(n25039), .dout(n25042));
    jdff dff_A_NyvscHrC9_2(.din(n3237), .dout(n25039));
    jdff dff_A_Ij8AChXO0_0(.din(n25033), .dout(G388));
    jdff dff_A_sdKYZNvW4_0(.din(n25030), .dout(n25033));
    jdff dff_A_ftUV2bVH7_0(.din(n25027), .dout(n25030));
    jdff dff_A_NXSWMPmp2_0(.din(n25024), .dout(n25027));
    jdff dff_A_cBOkQEx37_0(.din(n25021), .dout(n25024));
    jdff dff_A_KuuqqpVz0_0(.din(n25018), .dout(n25021));
    jdff dff_A_mcyC9mh01_0(.din(n25015), .dout(n25018));
    jdff dff_A_hToYVN4Y9_0(.din(n25012), .dout(n25015));
    jdff dff_A_AYdDzrQq9_0(.din(n25009), .dout(n25012));
    jdff dff_A_w1ntX4QK4_0(.din(n25006), .dout(n25009));
    jdff dff_A_Ngvebk253_0(.din(n25003), .dout(n25006));
    jdff dff_A_JERUK1X57_0(.din(n25000), .dout(n25003));
    jdff dff_A_jOZt3TJ25_0(.din(n24997), .dout(n25000));
    jdff dff_A_Y3lDAcRw4_0(.din(n24994), .dout(n24997));
    jdff dff_A_NED2kRvc1_0(.din(n24991), .dout(n24994));
    jdff dff_A_yFOsYNUg9_0(.din(n24988), .dout(n24991));
    jdff dff_A_M0lcvcBX0_0(.din(n24985), .dout(n24988));
    jdff dff_A_Wko3XSpy7_0(.din(n24982), .dout(n24985));
    jdff dff_A_wBzVYZfD6_0(.din(n24979), .dout(n24982));
    jdff dff_A_CP0LNn3C8_0(.din(n24976), .dout(n24979));
    jdff dff_A_VqUfarth3_0(.din(n24973), .dout(n24976));
    jdff dff_A_IzCSaNRG4_0(.din(n24970), .dout(n24973));
    jdff dff_A_Nt3WlxA69_0(.din(n24967), .dout(n24970));
    jdff dff_A_bB4avgpf0_0(.din(n24964), .dout(n24967));
    jdff dff_A_oa0XxNvS3_2(.din(n3233), .dout(n24964));
    jdff dff_A_pJJ0Ihlt6_0(.din(n24958), .dout(G264));
    jdff dff_A_jfYRn6PI6_0(.din(n24955), .dout(n24958));
    jdff dff_A_Q3yJPoNu6_0(.din(n24952), .dout(n24955));
    jdff dff_A_koFrxztT6_0(.din(n24949), .dout(n24952));
    jdff dff_A_jUpYjNDe8_0(.din(n24946), .dout(n24949));
    jdff dff_A_KT01SSCm0_0(.din(n24943), .dout(n24946));
    jdff dff_A_ShHN4Y151_0(.din(n24940), .dout(n24943));
    jdff dff_A_Rpdsh7GX8_0(.din(n24937), .dout(n24940));
    jdff dff_A_Iofqhzvn3_0(.din(n24934), .dout(n24937));
    jdff dff_A_9HZvrbM50_0(.din(n24931), .dout(n24934));
    jdff dff_A_6veNz4KY3_2(.din(n5508), .dout(n24931));
    jdff dff_A_xeF3ArdW7_0(.din(n24925), .dout(G258));
    jdff dff_A_9D32lsUc0_0(.din(n24922), .dout(n24925));
    jdff dff_A_ViaN4srH4_0(.din(n24919), .dout(n24922));
    jdff dff_A_5ULdjhRT0_0(.din(n24916), .dout(n24919));
    jdff dff_A_enRZMrRj2_0(.din(n24913), .dout(n24916));
    jdff dff_A_xZOhCyG66_0(.din(n24910), .dout(n24913));
    jdff dff_A_kfVPIFvh6_0(.din(n24907), .dout(n24910));
    jdff dff_A_JZLqlW553_0(.din(n24904), .dout(n24907));
    jdff dff_A_H3VhH1vY2_0(.din(n24901), .dout(n24904));
    jdff dff_A_nzl4gXeX9_0(.din(n24898), .dout(n24901));
    jdff dff_A_C7Y9DVay5_2(.din(n3173), .dout(n24898));
    jdff dff_A_0ioXxkSG6_0(.din(n24892), .dout(G373));
    jdff dff_A_T99Xbd8v0_0(.din(n24889), .dout(n24892));
    jdff dff_A_MvRVSvZU6_0(.din(n24886), .dout(n24889));
    jdff dff_A_OxPfMyx55_0(.din(n24883), .dout(n24886));
    jdff dff_A_tHYkYDFq7_0(.din(n24880), .dout(n24883));
    jdff dff_A_B5YKQYA75_0(.din(n24877), .dout(n24880));
    jdff dff_A_BBfr5o794_0(.din(n24874), .dout(n24877));
    jdff dff_A_aFXjbadQ2_0(.din(n24871), .dout(n24874));
    jdff dff_A_5a9NCTDT6_0(.din(n24868), .dout(n24871));
    jdff dff_A_n9g5SFgC7_0(.din(G5), .dout(n7855));
    jdff dff_A_7au7tv7s7_1(.din(G5), .dout(n7858));
    jdff dff_A_QQzWuTYo3_2(.din(G5), .dout(n7861));
    jdff dff_B_eVb1uE7h3_2(.din(n426), .dout(n7865));
    jdff dff_B_QW2NFVLj0_0(.din(n3217), .dout(n7868));
    jdff dff_B_iv2qALu13_1(.din(n3269), .dout(n7871));
    jdff dff_B_JL3Uxk8f4_1(.din(n1963), .dout(n7874));
    jdff dff_B_nVkUxcQh2_1(.din(n7874), .dout(n7877));
    jdff dff_B_dZFVaLSq9_1(.din(n7877), .dout(n7880));
    jdff dff_B_bxUYwUlW2_1(.din(n7880), .dout(n7883));
    jdff dff_B_rFvENq0u8_1(.din(n7883), .dout(n7886));
    jdff dff_B_hlzU7xKp9_1(.din(n7886), .dout(n7889));
    jdff dff_B_crLpbJdd3_1(.din(n7889), .dout(n7892));
    jdff dff_B_7ugGyDHY8_1(.din(n7892), .dout(n7895));
    jdff dff_B_aM0y4fTl0_1(.din(n7895), .dout(n7898));
    jdff dff_B_oKopyVDu0_1(.din(n7898), .dout(n7901));
    jdff dff_B_VzZUjfJJ3_1(.din(n7901), .dout(n7904));
    jdff dff_B_LysNLlf65_1(.din(n7904), .dout(n7907));
    jdff dff_B_ZSK9EZ2f6_1(.din(n7907), .dout(n7910));
    jdff dff_B_w359KRXJ1_1(.din(n7910), .dout(n7913));
    jdff dff_B_QDqV3Viq0_1(.din(n7913), .dout(n7916));
    jdff dff_B_izIiGylm2_1(.din(n7916), .dout(n7919));
    jdff dff_B_BQCItuAB9_1(.din(n7919), .dout(n7922));
    jdff dff_B_8HFHMBLa2_0(.din(n3161), .dout(n7925));
    jdff dff_B_Fh2BoDEf2_0(.din(n7925), .dout(n7928));
    jdff dff_B_LVM4weCC0_0(.din(n7928), .dout(n7931));
    jdff dff_B_gW8CMy1h9_0(.din(n7931), .dout(n7934));
    jdff dff_B_cxf56XXI2_0(.din(n7934), .dout(n7937));
    jdff dff_B_EALYBs6j4_0(.din(n7937), .dout(n7940));
    jdff dff_B_RfPtmtFx6_0(.din(n7940), .dout(n7943));
    jdff dff_B_HNUnMUZf5_0(.din(n7943), .dout(n7946));
    jdff dff_B_3yh1LDUD9_0(.din(n7946), .dout(n7949));
    jdff dff_B_rPsERgDg4_0(.din(n7949), .dout(n7952));
    jdff dff_B_6aWEYUU27_0(.din(n7952), .dout(n7955));
    jdff dff_B_2gyqvWcx3_0(.din(n7955), .dout(n7958));
    jdff dff_B_OJFaf4C45_0(.din(n7958), .dout(n7961));
    jdff dff_B_agc9kbSX2_0(.din(n7961), .dout(n7964));
    jdff dff_B_QhklNHYJ1_0(.din(n7964), .dout(n7967));
    jdff dff_B_4OlEFcVr6_0(.din(n7967), .dout(n7970));
    jdff dff_B_UWyCibH59_1(.din(n3125), .dout(n7973));
    jdff dff_B_8JBo7MtE0_1(.din(n7973), .dout(n7976));
    jdff dff_B_2JDqAnWF6_1(.din(n7976), .dout(n7979));
    jdff dff_B_PNmrDce39_1(.din(n7979), .dout(n7982));
    jdff dff_B_aLZtl6TB0_1(.din(n7982), .dout(n7985));
    jdff dff_B_PVYmZCkK3_1(.din(n3129), .dout(n7988));
    jdff dff_B_rhWpG1sa2_1(.din(n7988), .dout(n7991));
    jdff dff_B_LOovrd8T7_1(.din(n7991), .dout(n7994));
    jdff dff_B_gMtGkkf78_1(.din(n3133), .dout(n7997));
    jdff dff_B_Xgr1Rhsw9_0(.din(n3109), .dout(n8000));
    jdff dff_B_QB02PcLq1_0(.din(n8000), .dout(n8003));
    jdff dff_B_oatz0fpB2_0(.din(n8003), .dout(n8006));
    jdff dff_B_XQf3rFE19_0(.din(n8006), .dout(n8009));
    jdff dff_B_vxvH3OFK4_0(.din(n8009), .dout(n8012));
    jdff dff_B_GrPooNUC1_0(.din(n8012), .dout(n8015));
    jdff dff_B_OfgiU85C0_0(.din(n8015), .dout(n8018));
    jdff dff_B_qPumAjg09_0(.din(n8018), .dout(n8021));
    jdff dff_B_V0LyciSs5_0(.din(n8021), .dout(n8024));
    jdff dff_B_Ka3Cw3Gj3_0(.din(n8024), .dout(n8027));
    jdff dff_B_BJYVUQtv6_0(.din(n8027), .dout(n8030));
    jdff dff_B_GSjd4Lz08_0(.din(n8030), .dout(n8033));
    jdff dff_B_OQGKkDLd6_0(.din(n8033), .dout(n8036));
    jdff dff_B_uRaaM5jN4_0(.din(n8036), .dout(n8039));
    jdff dff_B_Q0RK8VJb7_0(.din(n8039), .dout(n8042));
    jdff dff_B_RtWilZ243_0(.din(n8042), .dout(n8045));
    jdff dff_B_g3X5V15h0_0(.din(n8045), .dout(n8048));
    jdff dff_B_nKOYJWaS6_1(.din(n3093), .dout(n8051));
    jdff dff_B_akVBs4rW7_1(.din(n8051), .dout(n8054));
    jdff dff_A_etnL63KJ2_0(.din(n3101), .dout(n8056));
    jdff dff_B_2PwnoF0C9_1(.din(n2109), .dout(n8060));
    jdff dff_B_BGoAAQot9_1(.din(n8060), .dout(n8063));
    jdff dff_B_mjwidCI77_1(.din(n8063), .dout(n8066));
    jdff dff_B_V9nMdID11_1(.din(n8066), .dout(n8069));
    jdff dff_B_tYdbC80R0_1(.din(n8069), .dout(n8072));
    jdff dff_B_TH4u9rLa8_1(.din(n8072), .dout(n8075));
    jdff dff_B_lAxSjQ1s9_1(.din(n8075), .dout(n8078));
    jdff dff_B_5FUHYWFc4_1(.din(n8078), .dout(n8081));
    jdff dff_B_En9U1VzK2_1(.din(n8081), .dout(n8084));
    jdff dff_B_N2JrJOuG9_1(.din(n8084), .dout(n8087));
    jdff dff_B_BlWityMK6_1(.din(n8087), .dout(n8090));
    jdff dff_B_jwk2BptA6_1(.din(n8090), .dout(n8093));
    jdff dff_B_zPqGfzw23_1(.din(n8093), .dout(n8096));
    jdff dff_B_RbCkI6so9_1(.din(n8096), .dout(n8099));
    jdff dff_B_q2ed6MJC2_1(.din(n8099), .dout(n8102));
    jdff dff_B_3dj0ESMk7_1(.din(n2123), .dout(n8105));
    jdff dff_B_Ly1Pwmrj8_1(.din(n8105), .dout(n8108));
    jdff dff_B_b8V7jSAR0_1(.din(n8108), .dout(n8111));
    jdff dff_B_ISYftX5M2_1(.din(n8111), .dout(n8114));
    jdff dff_B_OJlOckdU6_1(.din(n8114), .dout(n8117));
    jdff dff_B_3UocEI9x1_1(.din(n8117), .dout(n8120));
    jdff dff_B_Zltogmk66_1(.din(n8120), .dout(n8123));
    jdff dff_B_aGNbQitz5_1(.din(n8123), .dout(n8126));
    jdff dff_B_tGTEbQFu9_1(.din(n8126), .dout(n8129));
    jdff dff_B_t4PbNbjN9_1(.din(n8129), .dout(n8132));
    jdff dff_B_k4zYkSZL1_1(.din(n8132), .dout(n8135));
    jdff dff_B_pQAnTvFN7_1(.din(n8135), .dout(n8138));
    jdff dff_B_o6SHvsb31_1(.din(n8138), .dout(n8141));
    jdff dff_B_17DmmvCM8_1(.din(n8141), .dout(n8144));
    jdff dff_B_gbMbJoQG1_1(.din(n8144), .dout(n8147));
    jdff dff_B_CFcAvKLj6_0(.din(n3077), .dout(n8150));
    jdff dff_B_rQbrq56t8_0(.din(n8150), .dout(n8153));
    jdff dff_B_HmzUSUyA1_0(.din(n8153), .dout(n8156));
    jdff dff_B_QXc6b5cQ2_0(.din(n8156), .dout(n8159));
    jdff dff_B_X0FCGtHk4_0(.din(n8159), .dout(n8162));
    jdff dff_B_PRKVWczS3_0(.din(n8162), .dout(n8165));
    jdff dff_B_FDHQqxPH7_0(.din(n8165), .dout(n8168));
    jdff dff_B_CdpEen625_0(.din(n8168), .dout(n8171));
    jdff dff_B_h5sEIVQ94_0(.din(n8171), .dout(n8174));
    jdff dff_B_hIYWDFIz8_0(.din(n8174), .dout(n8177));
    jdff dff_B_JQlIRtgm7_0(.din(n8177), .dout(n8180));
    jdff dff_B_dHo87xgk2_0(.din(n8180), .dout(n8183));
    jdff dff_B_1QSc33RG0_0(.din(n8183), .dout(n8186));
    jdff dff_B_DWOeTdVH9_0(.din(n8186), .dout(n8189));
    jdff dff_B_A988JWCx6_0(.din(n8189), .dout(n8192));
    jdff dff_B_Wrw5Hqd19_0(.din(n8192), .dout(n8195));
    jdff dff_B_udaqWIxX2_1(.din(n2313), .dout(n8198));
    jdff dff_B_UtZYf41y7_1(.din(n8198), .dout(n8201));
    jdff dff_B_SnWwyTbr1_1(.din(n8201), .dout(n8204));
    jdff dff_B_DeBSnkJO1_1(.din(n8204), .dout(n8207));
    jdff dff_B_Ibq7IEn14_1(.din(n8207), .dout(n8210));
    jdff dff_B_V5letM908_1(.din(n8210), .dout(n8213));
    jdff dff_B_xZ4Xqwaj8_1(.din(n8213), .dout(n8216));
    jdff dff_B_DR71AT8P1_1(.din(n8216), .dout(n8219));
    jdff dff_B_1HW4sbfE6_1(.din(n8219), .dout(n8222));
    jdff dff_B_hqillBlo1_1(.din(n8222), .dout(n8225));
    jdff dff_B_jilyhg740_1(.din(n8225), .dout(n8228));
    jdff dff_B_kU0byQFR8_1(.din(n2317), .dout(n8231));
    jdff dff_B_Sx1uNu5a3_1(.din(n8231), .dout(n8234));
    jdff dff_B_dZGAQpab0_1(.din(n8234), .dout(n8237));
    jdff dff_B_xLdrZaIi8_1(.din(n8237), .dout(n8240));
    jdff dff_B_JqCmj6pN7_1(.din(n8240), .dout(n8243));
    jdff dff_B_4Wuzp8db7_1(.din(n8243), .dout(n8246));
    jdff dff_B_wZtY4F0h6_1(.din(n8246), .dout(n8249));
    jdff dff_B_LWD6H3D95_1(.din(n8249), .dout(n8252));
    jdff dff_B_FyyDFzm21_1(.din(n8252), .dout(n8255));
    jdff dff_B_hSbRrYUw8_1(.din(n8255), .dout(n8258));
    jdff dff_B_UAu2N2p05_1(.din(n8258), .dout(n8261));
    jdff dff_B_hDBXXTch2_1(.din(n8261), .dout(n8264));
    jdff dff_B_6ZZMi8gg9_1(.din(n8264), .dout(n8267));
    jdff dff_B_bp3JTHAO6_0(.din(n3057), .dout(n8270));
    jdff dff_B_VOa6mjkz4_0(.din(n8270), .dout(n8273));
    jdff dff_B_obl5F4as6_0(.din(n8273), .dout(n8276));
    jdff dff_B_gcpaaMQq6_0(.din(n8276), .dout(n8279));
    jdff dff_B_C5z9MrMH0_0(.din(n8279), .dout(n8282));
    jdff dff_B_F25zxsnW1_0(.din(n8282), .dout(n8285));
    jdff dff_B_xfLNtrgX0_0(.din(n8285), .dout(n8288));
    jdff dff_B_hNdKFqWY8_0(.din(n8288), .dout(n8291));
    jdff dff_B_w78BfbYk0_0(.din(n8291), .dout(n8294));
    jdff dff_B_IN28J2OI0_0(.din(n8294), .dout(n8297));
    jdff dff_B_g0IXKYU45_0(.din(n8297), .dout(n8300));
    jdff dff_B_4iCGeQns8_0(.din(n8300), .dout(n8303));
    jdff dff_B_Cz8YghvD9_0(.din(n8303), .dout(n8306));
    jdff dff_B_cuMzDEww9_0(.din(n8306), .dout(n8309));
    jdff dff_B_1fYsCXVZ7_0(.din(n2309), .dout(n8312));
    jdff dff_B_RuudyVQP2_0(.din(n8312), .dout(n8315));
    jdff dff_B_ZkmYrJx73_1(.din(n2293), .dout(n8318));
    jdff dff_B_fNbtVY718_1(.din(n2265), .dout(n8321));
    jdff dff_B_PkOzYPwq0_0(.din(n2257), .dout(n8324));
    jdff dff_A_ZGaBYqMV5_1(.din(n8329), .dout(n8326));
    jdff dff_A_K0UyC9ij2_1(.din(n2178), .dout(n8329));
    jdff dff_B_7UnKPXbe2_0(.din(n2105), .dout(n8333));
    jdff dff_B_AysCa2sL2_1(.din(n2089), .dout(n8336));
    jdff dff_A_hL4QtHdo2_1(.din(n2042), .dout(n8338));
    jdff dff_B_9uMlF7Ay0_2(.din(n2015), .dout(n8342));
    jdff dff_B_tsEoyIJd7_1(.din(n1872), .dout(n8345));
    jdff dff_B_dobygOqp2_1(.din(n8345), .dout(n8348));
    jdff dff_B_TSRR2EAS2_1(.din(n8348), .dout(n8351));
    jdff dff_B_br1cFjSc2_1(.din(n1876), .dout(n8354));
    jdff dff_B_m7N8lvTH8_1(.din(n8354), .dout(n8357));
    jdff dff_B_XLCg4Vxz6_1(.din(n1892), .dout(n8360));
    jdff dff_A_Jl51lhWb4_1(.din(n8365), .dout(n8362));
    jdff dff_A_YFJq84cV2_1(.din(n8368), .dout(n8365));
    jdff dff_A_UCuGhZcJ5_1(.din(n8371), .dout(n8368));
    jdff dff_A_lttAXzVh7_1(.din(n1848), .dout(n8371));
    jdff dff_B_wyZkRwqg1_3(.din(n1824), .dout(n8375));
    jdff dff_B_WFFcg9b19_3(.din(n8375), .dout(n8378));
    jdff dff_B_GjJNepL59_3(.din(n8378), .dout(n8381));
    jdff dff_B_3Y7CzIhi9_3(.din(n8381), .dout(n8384));
    jdff dff_B_5FjumPSY2_3(.din(n8384), .dout(n8387));
    jdff dff_B_lnJSQtNq1_3(.din(n8387), .dout(n8390));
    jdff dff_B_VYBVRL0s7_3(.din(n8390), .dout(n8393));
    jdff dff_B_cshPhwWY7_3(.din(n8393), .dout(n8396));
    jdff dff_B_fAR5PAi63_3(.din(n8396), .dout(n8399));
    jdff dff_B_Tstrbp4H5_3(.din(n8399), .dout(n8402));
    jdff dff_B_gwZrCtHh3_3(.din(n8402), .dout(n8405));
    jdff dff_B_ecySOCm87_3(.din(n8405), .dout(n8408));
    jdff dff_B_rYNRIiR07_3(.din(n8408), .dout(n8411));
    jdff dff_B_KfHtvRn50_3(.din(n8411), .dout(n8414));
    jdff dff_B_AnFO0cLV7_3(.din(n8414), .dout(n8417));
    jdff dff_B_qLiOIZ6E7_3(.din(n8417), .dout(n8420));
    jdff dff_B_36q99d5L1_3(.din(n8420), .dout(n8423));
    jdff dff_B_jN5ZtIgq2_3(.din(n8423), .dout(n8426));
    jdff dff_B_Z4txTq0q7_3(.din(n8426), .dout(n8429));
    jdff dff_B_CNLUHhKi7_3(.din(n8429), .dout(n8432));
    jdff dff_B_iTjKjlLP6_3(.din(n8432), .dout(n8435));
    jdff dff_B_NWmhIE741_3(.din(n8435), .dout(n8438));
    jdff dff_B_moekdsPF3_3(.din(n8438), .dout(n8441));
    jdff dff_B_47SaYpgW2_3(.din(n8441), .dout(n8444));
    jdff dff_B_Xp7qq0Vb4_0(.din(n1820), .dout(n8447));
    jdff dff_B_XwvYcmZv1_1(.din(n4114), .dout(n8450));
    jdff dff_B_1KBvtN5y0_1(.din(n8450), .dout(n8453));
    jdff dff_B_Z1MCnMhS5_1(.din(n8453), .dout(n8456));
    jdff dff_B_8p0wyfGX5_1(.din(n8456), .dout(n8459));
    jdff dff_B_BTItQeXr3_1(.din(n8459), .dout(n8462));
    jdff dff_B_GcJ6Qs3N9_1(.din(n8462), .dout(n8465));
    jdff dff_B_F2Ipz71k2_1(.din(n8465), .dout(n8468));
    jdff dff_B_Dnilearv7_1(.din(n8468), .dout(n8471));
    jdff dff_B_GanduZdd6_1(.din(n8471), .dout(n8474));
    jdff dff_B_OL0A4bTl4_1(.din(n8474), .dout(n8477));
    jdff dff_B_vEEIB46e3_1(.din(n8477), .dout(n8480));
    jdff dff_B_lxQHE9iJ3_1(.din(n8480), .dout(n8483));
    jdff dff_B_YGEwG3Zv8_1(.din(n8483), .dout(n8486));
    jdff dff_B_oZNzsOXp5_1(.din(n8486), .dout(n8489));
    jdff dff_B_PzZ9sjmD6_1(.din(n8489), .dout(n8492));
    jdff dff_B_jDmQfozV5_1(.din(n8492), .dout(n8495));
    jdff dff_B_OQxyPvgY5_1(.din(n8495), .dout(n8498));
    jdff dff_B_HZJ6luck2_1(.din(n8498), .dout(n8501));
    jdff dff_B_iu6b9rUm6_1(.din(n8501), .dout(n8504));
    jdff dff_B_kEcfKRZY5_1(.din(n8504), .dout(n8507));
    jdff dff_B_nnbLFFhQ7_1(.din(n8507), .dout(n8510));
    jdff dff_B_ypHWpTQ32_1(.din(n8510), .dout(n8513));
    jdff dff_B_LxQ2xTZx8_1(.din(n2463), .dout(n8516));
    jdff dff_B_6sAumDgf3_1(.din(n8516), .dout(n8519));
    jdff dff_B_kfwgKews0_1(.din(n8519), .dout(n8522));
    jdff dff_B_7Dn82H1x6_1(.din(n8522), .dout(n8525));
    jdff dff_B_jStP1M7t8_1(.din(n8525), .dout(n8528));
    jdff dff_B_tOhu7D1u7_1(.din(n8528), .dout(n8531));
    jdff dff_B_Mag9w8OI4_1(.din(n8531), .dout(n8534));
    jdff dff_B_ZdJKHoFX8_1(.din(n8534), .dout(n8537));
    jdff dff_B_lx5nZqAc0_1(.din(n8537), .dout(n8540));
    jdff dff_B_Oo0QY9Ih6_1(.din(n2475), .dout(n8543));
    jdff dff_B_QJBBCxc72_1(.din(n8543), .dout(n8546));
    jdff dff_B_ttWn3OQ39_1(.din(n8546), .dout(n8549));
    jdff dff_B_7TZ60Xwn9_1(.din(n8549), .dout(n8552));
    jdff dff_B_ZgiK9XAF4_1(.din(n8552), .dout(n8555));
    jdff dff_B_Plyq66uC2_1(.din(n8555), .dout(n8558));
    jdff dff_B_uNYCFD427_1(.din(n8558), .dout(n8561));
    jdff dff_B_P2UJUTcZ8_1(.din(n8561), .dout(n8564));
    jdff dff_B_YTkSdiyG8_1(.din(n8564), .dout(n8567));
    jdff dff_B_hoqQbiCM6_1(.din(n8567), .dout(n8570));
    jdff dff_B_8Nz34Ps88_0(.din(n3041), .dout(n8573));
    jdff dff_B_RF3upjcN2_0(.din(n8573), .dout(n8576));
    jdff dff_B_JB2wzUzL0_0(.din(n8576), .dout(n8579));
    jdff dff_B_sQ5WW1bI7_0(.din(n8579), .dout(n8582));
    jdff dff_B_Cwm1zvf69_0(.din(n8582), .dout(n8585));
    jdff dff_B_kKSLLmd88_0(.din(n8585), .dout(n8588));
    jdff dff_B_lh8VyK5u1_0(.din(n8588), .dout(n8591));
    jdff dff_B_B2omcMka9_0(.din(n8591), .dout(n8594));
    jdff dff_B_23Ep1ycX0_0(.din(n8594), .dout(n8597));
    jdff dff_B_otYfyN7k6_0(.din(n3027), .dout(n8600));
    jdff dff_B_mFzj0fnV1_0(.din(n8600), .dout(n8603));
    jdff dff_B_JQsr2JeB4_0(.din(n8603), .dout(n8606));
    jdff dff_B_QNMsegxi0_1(.din(n3003), .dout(n8609));
    jdff dff_B_PNhe6DRF0_1(.din(n8609), .dout(n8612));
    jdff dff_B_AwPlcsak5_1(.din(n8612), .dout(n8615));
    jdff dff_B_jorYkMEJ4_1(.din(n8615), .dout(n8618));
    jdff dff_B_Hhr9qj9p0_0(.din(n3019), .dout(n8621));
    jdff dff_B_fKc0yDPw9_0(.din(n8621), .dout(n8624));
    jdff dff_B_bLFA0pqD5_1(.din(n2987), .dout(n8627));
    jdff dff_B_vETxS4Ly4_0(.din(n2979), .dout(n8630));
    jdff dff_B_1vllwRkt2_0(.din(n8630), .dout(n8633));
    jdff dff_B_4bXAa7Qs8_0(.din(n8633), .dout(n8636));
    jdff dff_B_Z2MGMkkr8_1(.din(n2825), .dout(n8639));
    jdff dff_B_e3nt4qMF6_1(.din(n8639), .dout(n8642));
    jdff dff_B_34isNXdR2_1(.din(n8642), .dout(n8645));
    jdff dff_B_3JTNGUfp6_1(.din(n8645), .dout(n8648));
    jdff dff_B_iSDLFJwX9_1(.din(n8648), .dout(n8651));
    jdff dff_B_ge5PWEz40_0(.din(n2971), .dout(n8654));
    jdff dff_B_ZDcraaM70_0(.din(n8654), .dout(n8657));
    jdff dff_B_HgrYxgY77_0(.din(n8657), .dout(n8660));
    jdff dff_A_wbodIdqm6_0(.din(n8665), .dout(n8662));
    jdff dff_A_EAfLFRDE2_0(.din(n8668), .dout(n8665));
    jdff dff_A_ZZF8lVze4_0(.din(n8671), .dout(n8668));
    jdff dff_A_A4sJ5E0u2_0(.din(n2968), .dout(n8671));
    jdff dff_B_Ah2aUiDQ3_1(.din(n2945), .dout(n8675));
    jdff dff_A_ezWMIB7q9_0(.din(n2949), .dout(n8677));
    jdff dff_A_N3BsIWX12_1(.din(n2937), .dout(n8680));
    jdff dff_A_RhqxIhuS9_1(.din(n8687), .dout(n8683));
    jdff dff_B_83cBPOSs0_2(.din(n2880), .dout(n8687));
    jdff dff_B_sdDMOuXZ9_0(.din(n2794), .dout(n8690));
    jdff dff_B_LEgRd1n37_0(.din(n8690), .dout(n8693));
    jdff dff_B_P0OTCDOI4_0(.din(n8693), .dout(n8696));
    jdff dff_B_zkNYjj430_0(.din(n8696), .dout(n8699));
    jdff dff_B_tnYWgAfx1_0(.din(n8699), .dout(n8702));
    jdff dff_B_uZ9L45DT7_0(.din(n8702), .dout(n8705));
    jdff dff_B_orv1wjnb3_1(.din(n2778), .dout(n8708));
    jdff dff_B_CNN3Tmiw0_0(.din(n2770), .dout(n8711));
    jdff dff_B_4kWLMhoZ9_0(.din(n8711), .dout(n8714));
    jdff dff_B_xFBDYDCS7_0(.din(n8714), .dout(n8717));
    jdff dff_B_JdUiZGCi0_0(.din(n8717), .dout(n8720));
    jdff dff_B_3bJApQEN4_0(.din(n8720), .dout(n8723));
    jdff dff_B_estVN0us2_0(.din(n2766), .dout(n8726));
    jdff dff_B_NehKFbxp0_0(.din(n2706), .dout(n8729));
    jdff dff_B_9iZzCCub3_0(.din(n8729), .dout(n8732));
    jdff dff_B_CidzbUxa3_0(.din(n8732), .dout(n8735));
    jdff dff_B_MapM6INs9_0(.din(n8735), .dout(n8738));
    jdff dff_B_BppfZCnu1_0(.din(n8738), .dout(n8741));
    jdff dff_B_Nz54HwJD5_0(.din(n2670), .dout(n8744));
    jdff dff_B_ID7XDYqu7_0(.din(n8744), .dout(n8747));
    jdff dff_B_DwOjqOiE3_0(.din(n8747), .dout(n8750));
    jdff dff_B_k180PTCX8_0(.din(n8750), .dout(n8753));
    jdff dff_B_gxkXCOrE5_0(.din(n2631), .dout(n8756));
    jdff dff_B_zxf4LBxI1_0(.din(n8756), .dout(n8759));
    jdff dff_B_nggOTCOy9_0(.din(n8759), .dout(n8762));
    jdff dff_B_bo2wYj5S3_1(.din(n2499), .dout(n8765));
    jdff dff_B_q6EnlDxl3_1(.din(n8765), .dout(n8768));
    jdff dff_B_ZauRDTiH8_1(.din(n8768), .dout(n8771));
    jdff dff_B_wRFYCBmU5_0(.din(n2567), .dout(n8774));
    jdff dff_B_1SRk8rnZ7_0(.din(n8774), .dout(n8777));
    jdff dff_B_RnXkE3it4_0(.din(n2531), .dout(n8780));
    jdff dff_B_BNFVeHPN2_0(.din(n2527), .dout(n8783));
    jdff dff_A_ZZDYvtpd2_0(.din(G89), .dout(n8785));
    jdff dff_A_fwEvooYQ0_0(.din(n2523), .dout(n8788));
    jdff dff_B_xCGAEQP75_0(.din(n2459), .dout(n8792));
    jdff dff_B_R2ssDfRx2_1(.din(n2443), .dout(n8795));
    jdff dff_A_Ig6Jd2UU0_1(.din(n2396), .dout(n8797));
    jdff dff_A_RuXzwzZo6_1(.din(n2369), .dout(n8800));
    jdff dff_B_s5Hp0cC17_1(.din(n4266), .dout(n8804));
    jdff dff_B_y6tAviAl7_1(.din(n8804), .dout(n8807));
    jdff dff_B_eQadKVK99_1(.din(n4284), .dout(n8810));
    jdff dff_B_QOmj15Uf4_1(.din(n8810), .dout(n8813));
    jdff dff_B_c06RZygx3_1(.din(n8813), .dout(n8816));
    jdff dff_B_sjOvuJzq8_1(.din(n8816), .dout(n8819));
    jdff dff_B_OaYYyJIi8_1(.din(n8819), .dout(n8822));
    jdff dff_B_YYagu3qC3_1(.din(n8822), .dout(n8825));
    jdff dff_B_PNEekTyH5_1(.din(n8825), .dout(n8828));
    jdff dff_B_fUtICkG03_1(.din(n8828), .dout(n8831));
    jdff dff_B_NQhm448A5_1(.din(n8831), .dout(n8834));
    jdff dff_B_26CUA39Z9_1(.din(n8834), .dout(n8837));
    jdff dff_B_tnretszl7_1(.din(n8837), .dout(n8840));
    jdff dff_B_YnwHMZT42_1(.din(n8840), .dout(n8843));
    jdff dff_B_sfp0FJc35_1(.din(n8843), .dout(n8846));
    jdff dff_B_j8VXcBKN6_1(.din(n8846), .dout(n8849));
    jdff dff_B_b2IvIusC6_1(.din(n8849), .dout(n8852));
    jdff dff_B_PAWkJtJY9_1(.din(n8852), .dout(n8855));
    jdff dff_B_v8NiatIJ7_1(.din(n8855), .dout(n8858));
    jdff dff_B_j67HeSxg9_1(.din(n8858), .dout(n8861));
    jdff dff_B_rk62XQu75_1(.din(n8861), .dout(n8864));
    jdff dff_B_Yyae2c6K8_1(.din(n8864), .dout(n8867));
    jdff dff_B_PzBMoEd49_1(.din(n4347), .dout(n8870));
    jdff dff_B_IPsu51sy8_1(.din(n8870), .dout(n8873));
    jdff dff_B_YCx18kfC2_1(.din(n8873), .dout(n8876));
    jdff dff_B_EBsTKoK00_1(.din(n8876), .dout(n8879));
    jdff dff_B_Biz1UDPJ3_1(.din(n8879), .dout(n8882));
    jdff dff_B_5rz7YNcP1_1(.din(n8882), .dout(n8885));
    jdff dff_B_veDgjCRN8_1(.din(n8885), .dout(n8888));
    jdff dff_B_LlzMOLUu9_1(.din(n8888), .dout(n8891));
    jdff dff_B_jKGlioYE1_1(.din(n8891), .dout(n8894));
    jdff dff_B_r3vDdZ8X0_1(.din(n8894), .dout(n8897));
    jdff dff_B_3AZH8EsJ1_1(.din(n8897), .dout(n8900));
    jdff dff_B_TIhj8ilP0_1(.din(n8900), .dout(n8903));
    jdff dff_B_zAuZVIdH9_1(.din(n8903), .dout(n8906));
    jdff dff_B_mHSbwIWC5_1(.din(n8906), .dout(n8909));
    jdff dff_B_r0Yh98b39_1(.din(n8909), .dout(n8912));
    jdff dff_B_lEZTA7sg4_1(.din(n8912), .dout(n8915));
    jdff dff_B_Ib8tCxxr1_1(.din(n8915), .dout(n8918));
    jdff dff_B_YW26d8oN5_1(.din(n8918), .dout(n8921));
    jdff dff_B_gtvralSJ4_1(.din(n8921), .dout(n8924));
    jdff dff_B_50cW6R5h5_1(.din(n8924), .dout(n8927));
    jdff dff_B_9vv4BaAl1_1(.din(n8927), .dout(n8930));
    jdff dff_B_lT7YcpLB1_1(.din(n8930), .dout(n8933));
    jdff dff_B_RDORgMqD4_1(.din(n8933), .dout(n8936));
    jdff dff_B_ALJ4lXBz2_1(.din(n8936), .dout(n8939));
    jdff dff_B_LX7CG5Qt4_1(.din(n8939), .dout(n8942));
    jdff dff_B_LZwkqAo59_1(.din(n8942), .dout(n8945));
    jdff dff_B_1DLfnPfQ1_1(.din(n8945), .dout(n8948));
    jdff dff_B_EcLzNYaP2_1(.din(n8948), .dout(n8951));
    jdff dff_B_5DVjiJ859_1(.din(n8951), .dout(n8954));
    jdff dff_B_97LKRyJs4_1(.din(n8954), .dout(n8957));
    jdff dff_B_hy9CQt7z0_1(.din(n8957), .dout(n8960));
    jdff dff_B_JDntq90E5_1(.din(n8960), .dout(n8963));
    jdff dff_B_Vk81izGt4_1(.din(n8963), .dout(n8966));
    jdff dff_B_ahLpG0yz2_2(.din(n4179), .dout(n8969));
    jdff dff_B_A8Ubha8d9_2(.din(n8969), .dout(n8972));
    jdff dff_B_Pfp9khLw3_2(.din(n8972), .dout(n8975));
    jdff dff_B_JRXQ9fNn1_2(.din(n8975), .dout(n8978));
    jdff dff_B_IIjiu3Bv2_2(.din(n8978), .dout(n8981));
    jdff dff_B_oLXc25eD2_2(.din(n8981), .dout(n8984));
    jdff dff_B_HiNlUkE01_2(.din(n8984), .dout(n8987));
    jdff dff_B_wsUnivT46_2(.din(n8987), .dout(n8990));
    jdff dff_B_fsDYXqJj3_2(.din(n8990), .dout(n8993));
    jdff dff_B_cLBQPQYd8_2(.din(n8993), .dout(n8996));
    jdff dff_B_6NYEkpyw4_2(.din(n8996), .dout(n8999));
    jdff dff_B_Xzmf6IqD8_2(.din(n8999), .dout(n9002));
    jdff dff_B_YNLKOk187_2(.din(n9002), .dout(n9005));
    jdff dff_B_eQvRwRHh1_2(.din(n9005), .dout(n9008));
    jdff dff_B_LlkwaQ854_2(.din(n9008), .dout(n9011));
    jdff dff_B_ofEo3QIb5_2(.din(n9011), .dout(n9014));
    jdff dff_B_sOpolSFo4_2(.din(n9014), .dout(n9017));
    jdff dff_B_sqbqov2b6_2(.din(n9017), .dout(n9020));
    jdff dff_B_zQFllWNM0_2(.din(n9020), .dout(n9023));
    jdff dff_B_cRySGfZj1_2(.din(n9023), .dout(n9026));
    jdff dff_B_x3F9zCXM5_2(.din(n9026), .dout(n9029));
    jdff dff_B_Iwz6rXXn2_2(.din(n9029), .dout(n9032));
    jdff dff_B_2wAmErmz5_2(.din(n9032), .dout(n9035));
    jdff dff_B_nPlACwd95_2(.din(n9035), .dout(n9038));
    jdff dff_B_FfWgKOYy4_2(.din(n9038), .dout(n9041));
    jdff dff_B_1ul6ytrd7_2(.din(n9041), .dout(n9044));
    jdff dff_B_C7pro73t8_2(.din(n9044), .dout(n9047));
    jdff dff_B_xetpYuPs7_2(.din(n9047), .dout(n9050));
    jdff dff_B_eapPgTTJ3_2(.din(n9050), .dout(n9053));
    jdff dff_B_Nsi5X4a68_2(.din(n4350), .dout(n9056));
    jdff dff_B_Bh2we42W7_2(.din(n9056), .dout(n9059));
    jdff dff_B_ZQeZ26oA8_2(.din(n9059), .dout(n9062));
    jdff dff_B_XFy51k1n4_2(.din(n9062), .dout(n9065));
    jdff dff_B_0Ktn2SDL8_2(.din(n9065), .dout(n9068));
    jdff dff_B_V0recqrJ1_2(.din(n9068), .dout(n9071));
    jdff dff_B_3cYDWd4q5_2(.din(n9071), .dout(n9074));
    jdff dff_B_cCwouaHD3_2(.din(n9074), .dout(n9077));
    jdff dff_B_zOLsnwPo4_2(.din(n9077), .dout(n9080));
    jdff dff_B_TW8d3bdG2_2(.din(n9080), .dout(n9083));
    jdff dff_B_ZAW1SaQB6_2(.din(n9083), .dout(n9086));
    jdff dff_B_XL2DLYm64_2(.din(n9086), .dout(n9089));
    jdff dff_B_vOkVqBPd0_2(.din(n9089), .dout(n9092));
    jdff dff_B_N2PZ3a1Q0_2(.din(n9092), .dout(n9095));
    jdff dff_B_SH94kbda1_2(.din(n9095), .dout(n9098));
    jdff dff_B_4a0rIBNL6_2(.din(n9098), .dout(n9101));
    jdff dff_B_Gor3mNL25_2(.din(n9101), .dout(n9104));
    jdff dff_B_7vaA25NE1_2(.din(n9104), .dout(n9107));
    jdff dff_B_0YPyJ8Uc4_2(.din(n9107), .dout(n9110));
    jdff dff_B_aXUwLWky9_2(.din(n9110), .dout(n9113));
    jdff dff_B_2eIhZ2w12_2(.din(n9113), .dout(n9116));
    jdff dff_B_C4w7ZstR7_2(.din(n9116), .dout(n9119));
    jdff dff_B_JjtbViYg2_2(.din(n9119), .dout(n9122));
    jdff dff_B_vGWTtvqL1_2(.din(n9122), .dout(n9125));
    jdff dff_B_7ZadreeO3_2(.din(n9125), .dout(n9128));
    jdff dff_B_agoTf6pK2_2(.din(n9128), .dout(n9131));
    jdff dff_B_lCJ7p6YX6_2(.din(n9131), .dout(n9134));
    jdff dff_B_rqPDnjiC8_2(.din(n9134), .dout(n9137));
    jdff dff_B_vuxAlKJW3_2(.din(n9137), .dout(n9140));
    jdff dff_B_gm6zH1U62_2(.din(n9140), .dout(n9143));
    jdff dff_B_rYSpOFRW4_2(.din(n9143), .dout(n9146));
    jdff dff_B_nnIPsxnx3_1(.din(n4381), .dout(n9149));
    jdff dff_B_oJ3uk5Yu9_1(.din(n9149), .dout(n9152));
    jdff dff_B_5GBMW2tW7_1(.din(n4385), .dout(n9155));
    jdff dff_B_SQrA1Ldx3_1(.din(n9155), .dout(n9158));
    jdff dff_B_QfoNWJZa1_1(.din(n9158), .dout(n9161));
    jdff dff_B_jZ1VNd3j9_1(.din(n9161), .dout(n9164));
    jdff dff_B_zbpEuFZc3_1(.din(n9164), .dout(n9167));
    jdff dff_B_6neiXGcZ2_1(.din(n9167), .dout(n9170));
    jdff dff_B_WsznJuhN4_1(.din(n9170), .dout(n9173));
    jdff dff_B_D3ju29x52_1(.din(n9173), .dout(n9176));
    jdff dff_B_NRiDnaVs1_0(.din(n4389), .dout(n9179));
    jdff dff_B_xYAtRbtz9_0(.din(n9179), .dout(n9182));
    jdff dff_B_0P283q1G0_0(.din(n9182), .dout(n9185));
    jdff dff_B_DwLSuusb8_0(.din(n9185), .dout(n9188));
    jdff dff_B_e5eFDp330_0(.din(n9188), .dout(n9191));
    jdff dff_B_qNU6KT989_0(.din(n9191), .dout(n9194));
    jdff dff_B_hU40mBNJ5_0(.din(n9194), .dout(n9197));
    jdff dff_B_rfMi1FXX7_0(.din(n3621), .dout(n9200));
    jdff dff_B_nYIWO4Zh3_0(.din(n3617), .dout(n9203));
    jdff dff_B_qZ37TkEr6_0(.din(n3609), .dout(n9206));
    jdff dff_B_iO12gpId8_1(.din(n3597), .dout(n9209));
    jdff dff_B_hETOkRjX2_0(.din(n3577), .dout(n9212));
    jdff dff_B_7CjXRu199_1(.din(n3528), .dout(n9215));
    jdff dff_B_MEpDpiEk0_1(.din(n9215), .dout(n9218));
    jdff dff_B_jhQ9ZwHH8_1(.din(n9218), .dout(n9221));
    jdff dff_B_r4wVXBmI4_1(.din(n9221), .dout(n9224));
    jdff dff_B_ElLWtjbo3_1(.din(n3546), .dout(n9227));
    jdff dff_B_yxh4zwZu0_0(.din(n3508), .dout(n9230));
    jdff dff_B_DruvH7gb4_0(.din(n9230), .dout(n9233));
    jdff dff_B_VqDCOUdL7_0(.din(n3500), .dout(n9236));
    jdff dff_B_T8lypvRC0_0(.din(n3480), .dout(n9239));
    jdff dff_B_L7MDHylB8_1(.din(n3456), .dout(n9242));
    jdff dff_B_gX7dCrmQ4_0(.din(n3468), .dout(n9245));
    jdff dff_B_8KC414ka4_1(.din(n3460), .dout(n9248));
    jdff dff_B_oSRhgFo17_1(.din(n3399), .dout(n9251));
    jdff dff_B_cxn5ESvY5_1(.din(n3403), .dout(n9254));
    jdff dff_B_31ztlG9W9_1(.din(n9254), .dout(n9257));
    jdff dff_B_LCvwGGe99_0(.din(n3440), .dout(n9260));
    jdff dff_B_jXbhs1Ts2_0(.din(n9260), .dout(n9263));
    jdff dff_B_gg1Pz5RC7_0(.din(n3395), .dout(n9266));
    jdff dff_B_dxTagTcf8_0(.din(n4107), .dout(n9269));
    jdff dff_B_8NSQiVkX4_1(.din(n4055), .dout(n9272));
    jdff dff_B_pwJz712V9_1(.din(n9272), .dout(n9275));
    jdff dff_B_9OoVwt040_0(.din(n4099), .dout(n9278));
    jdff dff_B_78xqVym44_0(.din(n9278), .dout(n9281));
    jdff dff_B_VCPo7aj54_0(.din(n2209), .dout(n9284));
    jdff dff_B_HI17SWLs1_0(.din(n2182), .dout(n9287));
    jdff dff_B_xlnYYd9P9_0(.din(G174), .dout(n9290));
    jdff dff_B_rilexsIN7_0(.din(G173), .dout(n9293));
    jdff dff_B_ACptuE0V4_0(.din(G176), .dout(n9296));
    jdff dff_B_lVJBxmwj6_0(.din(G175), .dout(n9299));
    jdff dff_B_8afCptDr6_0(.din(n2154), .dout(n9302));
    jdff dff_B_neYfZjv58_0(.din(G177), .dout(n9305));
    jdff dff_A_dvAMxUoN8_0(.din(n521), .dout(n9307));
    jdff dff_B_XobirX4R6_0(.din(n2237), .dout(n9311));
    jdff dff_B_bqA7wn954_1(.din(n3984), .dout(n9314));
    jdff dff_B_wiIQHOaU6_1(.din(n9314), .dout(n9317));
    jdff dff_B_bWgIHx2K6_1(.din(n9317), .dout(n9320));
    jdff dff_B_yr36TW4i6_1(.din(n9320), .dout(n9323));
    jdff dff_B_9B07w0IG3_1(.din(n4002), .dout(n9326));
    jdff dff_A_kPtUaf2H8_0(.din(n9331), .dout(n9328));
    jdff dff_A_PpFG70SJ1_0(.din(n1852), .dout(n9331));
    jdff dff_B_X6BYXpZV8_0(.din(G167), .dout(n9335));
    jdff dff_A_kCiJr1094_0(.din(n9340), .dout(n9337));
    jdff dff_A_2hx7wOQO9_0(.din(n1828), .dout(n9340));
    jdff dff_B_LdDA1UfB9_0(.din(G166), .dout(n9344));
    jdff dff_B_q4LyJ9mr1_0(.din(G169), .dout(n9347));
    jdff dff_A_8Cb6vKBt0_2(.din(n521), .dout(n9349));
    jdff dff_B_IC7aNWb99_0(.din(G168), .dout(n9353));
    jdff dff_B_4OUwLuKY1_1(.din(G170), .dout(n9356));
    jdff dff_B_9v9MOOrH2_1(.din(n3933), .dout(n9359));
    jdff dff_B_mVGGaIz23_0(.din(n2345), .dout(n9362));
    jdff dff_A_9BgNPRCU5_1(.din(n2325), .dout(n9364));
    jdff dff_B_mTocefGd9_0(.din(n2321), .dout(n9368));
    jdff dff_B_lnZwKp530_0(.din(n3941), .dout(n9371));
    jdff dff_B_CwWHlkEl2_0(.din(G115), .dout(n9374));
    jdff dff_B_fT6cpS2r5_0(.din(n2802), .dout(n9377));
    jdff dff_B_NfZNRfxe8_0(.din(n2856), .dout(n9380));
    jdff dff_B_fFR3xlQT2_0(.din(n2829), .dout(n9383));
    jdff dff_B_XXe0m7kV4_0(.din(n2914), .dout(n9386));
    jdff dff_B_cQLPEVoP8_0(.din(n2884), .dout(n9389));
    jdff dff_B_dnkm3fBP6_0(.din(n2404), .dout(n9392));
    jdff dff_B_fV89OfNc8_0(.din(n2373), .dout(n9395));
    jdff dff_B_g6xz6nVJ6_0(.din(n3913), .dout(n9398));
    jdff dff_B_bxk0bZM88_0(.din(n2539), .dout(n9401));
    jdff dff_B_MxQHdMvy2_0(.din(n2503), .dout(n9404));
    jdff dff_B_ZKWIEJTp2_0(.din(n2603), .dout(n9407));
    jdff dff_B_9SokRwpu0_0(.din(n2479), .dout(n9410));
    jdff dff_B_9bgLBXQJ9_0(.din(n3893), .dout(n9413));
    jdff dff_B_Jrk5eOK59_0(.din(n3885), .dout(n9416));
    jdff dff_B_1rrGnPMp2_0(.din(G44), .dout(n9419));
    jdff dff_B_5YrEWmCa8_0(.din(n3877), .dout(n9422));
    jdff dff_B_4nTjbmam1_0(.din(n2738), .dout(n9425));
    jdff dff_B_tC5oChiN6_0(.din(n2714), .dout(n9428));
    jdff dff_B_q9i22s8O9_0(.din(n2678), .dout(n9431));
    jdff dff_A_ZFgUO11s5_0(.din(n2647), .dout(n9433));
    jdff dff_B_4s9IArk87_0(.din(n2643), .dout(n9437));
    jdff dff_A_ERBY7ag16_0(.din(n3866), .dout(n9439));
    jdff dff_B_gRr2QMWX6_1(.din(n3819), .dout(n9443));
    jdff dff_B_Y00uvtA76_1(.din(n9443), .dout(n9446));
    jdff dff_B_VaOgOo7R7_0(.din(n3850), .dout(n9449));
    jdff dff_B_FIx2mURg1_0(.din(n3842), .dout(n9452));
    jdff dff_B_U8wghQvY4_0(.din(n1884), .dout(n9455));
    jdff dff_B_KVIsyAul7_0(.din(n1935), .dout(n9458));
    jdff dff_B_oVCXBg7B5_0(.din(n1911), .dout(n9461));
    jdff dff_B_PknzMfj32_0(.din(n1864), .dout(n9464));
    jdff dff_B_suekqKZF4_0(.din(n1840), .dout(n9467));
    jdff dff_A_Cid0r0AO1_0(.din(G2204), .dout(n9469));
    jdff dff_A_RIAEFIVh8_2(.din(n9475), .dout(n9472));
    jdff dff_A_1ikDeAhx6_2(.din(G18), .dout(n9475));
    jdff dff_B_UT7DX8AU3_1(.din(n3757), .dout(n9479));
    jdff dff_B_mmKU2qf88_1(.din(n3761), .dout(n9482));
    jdff dff_B_hIfhACI74_0(.din(n2929), .dout(n9485));
    jdff dff_A_HQPL7rNf1_0(.din(G18), .dout(n9487));
    jdff dff_B_lmDZK8E89_0(.din(n2899), .dout(n9491));
    jdff dff_B_VAnidCBK9_1(.din(n3765), .dout(n9494));
    jdff dff_A_t7Tf8XrA0_1(.din(n455), .dout(n9496));
    jdff dff_B_8rIQAGib9_0(.din(n2817), .dout(n9500));
    jdff dff_B_UQfx4r7m6_0(.din(n2868), .dout(n9503));
    jdff dff_B_l3G4sekk1_0(.din(n2844), .dout(n9506));
    jdff dff_B_i1Wnk4No1_0(.din(n2419), .dout(n9509));
    jdff dff_B_sQF7XcW14_0(.din(n2388), .dout(n9512));
    jdff dff_B_VMN7qhTg7_0(.din(n2357), .dout(n9515));
    jdff dff_B_bTJoSfQD1_0(.din(n2333), .dout(n9518));
    jdff dff_B_LWRHO66N8_1(.din(n3691), .dout(n9521));
    jdff dff_A_6HllCUn99_0(.din(n2694), .dout(n9523));
    jdff dff_B_DjGqyaxc6_0(.din(n2690), .dout(n9527));
    jdff dff_B_GVGkWjOU8_0(.din(n2658), .dout(n9530));
    jdff dff_A_rNjZUdEz4_0(.din(n2563), .dout(n9532));
    jdff dff_B_erXJUqiE4_0(.din(n2615), .dout(n9536));
    jdff dff_B_jCyB9P0P2_0(.din(n3702), .dout(n9539));
    jdff dff_B_LTj0zE0V5_0(.din(n2491), .dout(n9542));
    jdff dff_B_6S7kVID85_0(.din(n2551), .dout(n9545));
    jdff dff_B_bEl0xenY5_0(.din(n2515), .dout(n9548));
    jdff dff_B_K8YkDxMJ7_0(.din(n2750), .dout(n9551));
    jdff dff_B_kX1qkxWd0_0(.din(n2726), .dout(n9554));
    jdff dff_B_ZDQVdoiT8_0(.din(n3671), .dout(n9557));
    jdff dff_B_6S4NPvSl2_0(.din(n2003), .dout(n9560));
    jdff dff_B_hZpeGKhD7_0(.din(n1979), .dout(n9563));
    jdff dff_B_LlYTllIS2_0(.din(n2221), .dout(n9566));
    jdff dff_B_aJMHWVVK0_0(.din(n2197), .dout(n9569));
    jdff dff_B_IHKWq1ZS2_0(.din(n2166), .dout(n9572));
    jdff dff_B_Q1fKgDge9_0(.din(n2142), .dout(n9575));
    jdff dff_B_eweljXyV3_0(.din(n3651), .dout(n9578));
    jdff dff_B_motdm5k38_0(.din(n3643), .dout(n9581));
    jdff dff_B_NXZo4Vpb7_0(.din(n2249), .dout(n9584));
    jdff dff_A_RwjGpHMx3_0(.din(n2069), .dout(n9586));
    jdff dff_B_MevoUuZj5_0(.din(n2065), .dout(n9590));
    jdff dff_B_rZiy9hkI1_0(.din(n2034), .dout(n9593));
    jdff dff_B_7harNJMF0_3(.din(n1812), .dout(n9596));
    jdff dff_B_8OB2MLuA2_3(.din(n9596), .dout(n9599));
    jdff dff_B_YnPVhjWc0_3(.din(n9599), .dout(n9602));
    jdff dff_B_eu4nILTo8_3(.din(n9602), .dout(n9605));
    jdff dff_B_Vk2AVHSq9_3(.din(n9605), .dout(n9608));
    jdff dff_B_LJJj8OGw5_3(.din(n9608), .dout(n9611));
    jdff dff_B_HIa3BgOe6_3(.din(n9611), .dout(n9614));
    jdff dff_B_JgJYS9W98_3(.din(n9614), .dout(n9617));
    jdff dff_B_ESPycNKz5_3(.din(n9617), .dout(n9620));
    jdff dff_B_yWHsUTY29_3(.din(n9620), .dout(n9623));
    jdff dff_B_0gzNXEkO3_3(.din(n9623), .dout(n9626));
    jdff dff_B_VvcJRpKe3_3(.din(n9626), .dout(n9629));
    jdff dff_B_Pf0PwEVi3_3(.din(n9629), .dout(n9632));
    jdff dff_B_WPCQJIqE3_3(.din(n9632), .dout(n9635));
    jdff dff_B_58YVGJTN1_3(.din(n9635), .dout(n9638));
    jdff dff_B_MdRPCVhl7_3(.din(n9638), .dout(n9641));
    jdff dff_B_Oew8zBW70_3(.din(n9641), .dout(n9644));
    jdff dff_B_w0Mvhv1d9_3(.din(n9644), .dout(n9647));
    jdff dff_B_c8js4H3A1_3(.din(n9647), .dout(n9650));
    jdff dff_B_MBpvApYr2_3(.din(n9650), .dout(n9653));
    jdff dff_B_6rziHhf50_3(.din(n9653), .dout(n9656));
    jdff dff_B_YeNXfyw63_3(.din(n9656), .dout(n9659));
    jdff dff_B_yOSJnDMg0_3(.din(n9659), .dout(n9662));
    jdff dff_B_U4aXV4h35_3(.din(n9662), .dout(n9665));
    jdff dff_B_qEa75UDU2_3(.din(n9665), .dout(n9668));
    jdff dff_B_GVWJ8yq63_3(.din(n9668), .dout(n9671));
    jdff dff_B_zSMpWHB00_3(.din(n9671), .dout(n9674));
    jdff dff_B_v4tQL05P7_3(.din(n9674), .dout(n9677));
    jdff dff_B_Jl9eAITO4_3(.din(n9677), .dout(n9680));
    jdff dff_B_E0sjvPnC4_3(.din(n9680), .dout(n9683));
    jdff dff_B_jz4mq0wf2_3(.din(n9683), .dout(n9686));
    jdff dff_B_htuktq9e4_3(.din(n9686), .dout(n9689));
    jdff dff_B_cHzQtCIR4_3(.din(n9689), .dout(n9692));
    jdff dff_B_jHOlOr462_3(.din(n9692), .dout(n9695));
    jdff dff_B_ZQL03hyj8_0(.din(n1808), .dout(n9698));
    jdff dff_B_twlXeJ7q4_1(.din(n4448), .dout(n9701));
    jdff dff_B_XtVTCOOT6_1(.din(n9701), .dout(n9704));
    jdff dff_B_0ajKQru93_1(.din(n9704), .dout(n9707));
    jdff dff_B_mObBsoMl9_1(.din(n9707), .dout(n9710));
    jdff dff_B_5NRuV43X0_1(.din(n9710), .dout(n9713));
    jdff dff_B_T6QZYIjE6_1(.din(n9713), .dout(n9716));
    jdff dff_B_z2e1mNPa3_1(.din(n9716), .dout(n9719));
    jdff dff_B_JDGzKElI0_1(.din(n9719), .dout(n9722));
    jdff dff_B_jZweMMIS4_1(.din(n9722), .dout(n9725));
    jdff dff_B_rmHqHeNi5_1(.din(n9725), .dout(n9728));
    jdff dff_B_tkqYSXQp0_1(.din(n9728), .dout(n9731));
    jdff dff_B_JyJLMoj38_1(.din(n9731), .dout(n9734));
    jdff dff_B_NOccPzQb0_1(.din(n9734), .dout(n9737));
    jdff dff_B_h6faLEoc9_1(.din(n9737), .dout(n9740));
    jdff dff_B_DpojqN0o5_1(.din(n9740), .dout(n9743));
    jdff dff_B_PERSpz908_1(.din(n9743), .dout(n9746));
    jdff dff_B_Lpz9wFYH3_1(.din(n9746), .dout(n9749));
    jdff dff_B_iBF0zSIX9_1(.din(n9749), .dout(n9752));
    jdff dff_B_yEufKW7X7_1(.din(n9752), .dout(n9755));
    jdff dff_B_fq0e9X9X7_1(.din(n9755), .dout(n9758));
    jdff dff_B_FJr2wMqf2_1(.din(n9758), .dout(n9761));
    jdff dff_B_03xCJqGp8_1(.din(n9761), .dout(n9764));
    jdff dff_B_sVVjQfj48_1(.din(n9764), .dout(n9767));
    jdff dff_B_BKunGsue7_1(.din(n9767), .dout(n9770));
    jdff dff_B_8R73yoEh1_1(.din(n9770), .dout(n9773));
    jdff dff_B_qjyl5HXG2_1(.din(n9773), .dout(n9776));
    jdff dff_B_7EXr7k8h9_1(.din(n9776), .dout(n9779));
    jdff dff_B_0IJlOyoJ7_1(.din(n9779), .dout(n9782));
    jdff dff_B_sUkka6jM2_1(.din(n9782), .dout(n9785));
    jdff dff_B_RSrplJz97_1(.din(n9785), .dout(n9788));
    jdff dff_B_q3iB6P8T0_1(.din(n9788), .dout(n9791));
    jdff dff_B_gBVPGCjC2_1(.din(n9791), .dout(n9794));
    jdff dff_B_PO5zx7vC7_1(.din(n9794), .dout(n9797));
    jdff dff_B_5a4TbPj14_1(.din(n9797), .dout(n9800));
    jdff dff_A_HBTyAc6I7_0(.din(n9805), .dout(n9802));
    jdff dff_A_eMHmEffM2_0(.din(n9808), .dout(n9805));
    jdff dff_A_5RNSaOsB4_0(.din(n9811), .dout(n9808));
    jdff dff_A_7QrLGILF0_0(.din(n9814), .dout(n9811));
    jdff dff_A_UqDAvpNu7_0(.din(n9817), .dout(n9814));
    jdff dff_A_08piZveL4_0(.din(n9820), .dout(n9817));
    jdff dff_A_GLjZCPGx4_0(.din(n9823), .dout(n9820));
    jdff dff_A_dGsttuS78_0(.din(n9826), .dout(n9823));
    jdff dff_A_R3LwgNdi5_0(.din(n9829), .dout(n9826));
    jdff dff_A_z2ZIgc8r4_0(.din(n9832), .dout(n9829));
    jdff dff_A_DYkcfs9h4_0(.din(n9835), .dout(n9832));
    jdff dff_A_9ULzOk1L2_0(.din(n9838), .dout(n9835));
    jdff dff_A_a9dCG73h6_0(.din(n9841), .dout(n9838));
    jdff dff_A_V3cVFiR18_0(.din(n9844), .dout(n9841));
    jdff dff_A_xwI6hixk2_0(.din(n9847), .dout(n9844));
    jdff dff_A_83rLeqmB9_0(.din(n9850), .dout(n9847));
    jdff dff_A_XXUM6CNb9_0(.din(n9853), .dout(n9850));
    jdff dff_A_5zaQv1Fu1_0(.din(n9856), .dout(n9853));
    jdff dff_A_migGWQ6K0_0(.din(n9859), .dout(n9856));
    jdff dff_A_lbXWVGxB4_0(.din(n9862), .dout(n9859));
    jdff dff_A_uo4fPLGn1_0(.din(n9865), .dout(n9862));
    jdff dff_A_9v7X2MgY2_0(.din(n9868), .dout(n9865));
    jdff dff_A_zh8uifpR5_0(.din(n9871), .dout(n9868));
    jdff dff_A_XDFsk4m49_0(.din(n9874), .dout(n9871));
    jdff dff_A_t8tGgAvN9_0(.din(n9877), .dout(n9874));
    jdff dff_A_IvULAnd04_0(.din(n9880), .dout(n9877));
    jdff dff_A_5inUDP0s4_0(.din(n9883), .dout(n9880));
    jdff dff_A_lDbIQf1M1_0(.din(n9886), .dout(n9883));
    jdff dff_A_TLi6Ey8p3_0(.din(n9889), .dout(n9886));
    jdff dff_A_C4WFfANq9_0(.din(n9892), .dout(n9889));
    jdff dff_A_UID0nzDd2_0(.din(n9895), .dout(n9892));
    jdff dff_A_brOidayp1_0(.din(n9898), .dout(n9895));
    jdff dff_A_1NxDNOAD3_0(.din(n1804), .dout(n9898));
    jdff dff_A_wVLQgSOY1_0(.din(n11092), .dout(n9901));
    jdff dff_A_ihZcVA6G5_1(.din(n11092), .dout(n9904));
    jdff dff_A_BHKCSiIk4_0(.din(n9910), .dout(n9907));
    jdff dff_A_2FSUKeD00_0(.din(n10013), .dout(n9910));
    jdff dff_A_cEOHc9J08_1(.din(n9916), .dout(n9913));
    jdff dff_A_ehSBP0Yb4_1(.din(n10013), .dout(n9916));
    jdff dff_B_q0LQ1LIh0_3(.din(n511), .dout(n9920));
    jdff dff_B_E7JCIvke2_3(.din(n9920), .dout(n9923));
    jdff dff_B_wMLwoEFJ5_3(.din(n9923), .dout(n9926));
    jdff dff_B_FFS9hwVn0_3(.din(n9926), .dout(n9929));
    jdff dff_B_Gj4y2JOc4_3(.din(n9929), .dout(n9932));
    jdff dff_B_6PjPud009_3(.din(n9932), .dout(n9935));
    jdff dff_B_0Zy8qH1L9_3(.din(n9935), .dout(n9938));
    jdff dff_B_mHJbPJ679_3(.din(n9938), .dout(n9941));
    jdff dff_B_tBka5SwJ4_3(.din(n9941), .dout(n9944));
    jdff dff_B_DdEpOIuM5_3(.din(n9944), .dout(n9947));
    jdff dff_B_RerjznoS2_3(.din(n9947), .dout(n9950));
    jdff dff_B_6iBaV3qT7_3(.din(n9950), .dout(n9953));
    jdff dff_B_y2IhB3Wx2_3(.din(n9953), .dout(n9956));
    jdff dff_B_JFyCRsdG0_3(.din(n9956), .dout(n9959));
    jdff dff_B_KuS2jGWu0_3(.din(n9959), .dout(n9962));
    jdff dff_B_xuvGn3c46_3(.din(n9962), .dout(n9965));
    jdff dff_B_pc5SgHtI1_3(.din(n9965), .dout(n9968));
    jdff dff_B_xUOIYxBN4_3(.din(n9968), .dout(n9971));
    jdff dff_B_DVHmYXEY2_3(.din(n9971), .dout(n9974));
    jdff dff_B_vEQQW6vH5_3(.din(n9974), .dout(n9977));
    jdff dff_B_0TcigI3U1_3(.din(n9977), .dout(n9980));
    jdff dff_B_AlUWaXrM6_3(.din(n9980), .dout(n9983));
    jdff dff_B_UJ55DKDV2_3(.din(n9983), .dout(n9986));
    jdff dff_B_adZOlTAc3_3(.din(n9986), .dout(n9989));
    jdff dff_B_ZtTqyoaC8_3(.din(n9989), .dout(n9992));
    jdff dff_B_IIYzzFNh4_3(.din(n9992), .dout(n9995));
    jdff dff_B_XKCGeKdu6_3(.din(n9995), .dout(n9998));
    jdff dff_B_xIIADPOF8_3(.din(n9998), .dout(n10001));
    jdff dff_B_pKKk1fqI5_3(.din(n10001), .dout(n10004));
    jdff dff_B_3UxzEWLV4_3(.din(n10004), .dout(n10007));
    jdff dff_B_otunNgPD3_3(.din(n10007), .dout(n10010));
    jdff dff_B_nxbVmBxn9_3(.din(n10010), .dout(n10013));
    jdff dff_B_gPMZX7B71_1(.din(n493), .dout(n10016));
    jdff dff_A_DpxLS1m19_2(.din(n10121), .dout(n10018));
    jdff dff_B_Uq11c23E3_3(.din(n485), .dout(n10022));
    jdff dff_B_QhcL4qzt4_3(.din(n10022), .dout(n10025));
    jdff dff_B_1mfOWhPf0_3(.din(n10025), .dout(n10028));
    jdff dff_B_Rosh9z2W5_3(.din(n10028), .dout(n10031));
    jdff dff_B_LvtAVJsN0_3(.din(n10031), .dout(n10034));
    jdff dff_B_3RjnZiL48_3(.din(n10034), .dout(n10037));
    jdff dff_B_rPE1qjcr5_3(.din(n10037), .dout(n10040));
    jdff dff_B_a8fbWRL04_3(.din(n10040), .dout(n10043));
    jdff dff_B_epQU5li38_3(.din(n10043), .dout(n10046));
    jdff dff_B_FeAzPCQL2_3(.din(n10046), .dout(n10049));
    jdff dff_B_ZLhaZyTj5_3(.din(n10049), .dout(n10052));
    jdff dff_B_UOMizGQl3_3(.din(n10052), .dout(n10055));
    jdff dff_B_Zf7VFlvj9_3(.din(n10055), .dout(n10058));
    jdff dff_B_PlUhUOXm0_3(.din(n10058), .dout(n10061));
    jdff dff_B_7fTbE3Qs0_3(.din(n10061), .dout(n10064));
    jdff dff_B_140LrTg14_3(.din(n10064), .dout(n10067));
    jdff dff_B_meu9KNNh7_3(.din(n10067), .dout(n10070));
    jdff dff_B_MlF8rQDI4_3(.din(n10070), .dout(n10073));
    jdff dff_B_p1VP9w0V4_3(.din(n10073), .dout(n10076));
    jdff dff_B_laQWJH2k2_3(.din(n10076), .dout(n10079));
    jdff dff_B_nh8BRbDh6_3(.din(n10079), .dout(n10082));
    jdff dff_B_VLp3duVg2_3(.din(n10082), .dout(n10085));
    jdff dff_B_jIgyEFNl8_3(.din(n10085), .dout(n10088));
    jdff dff_B_LO4dsblm8_3(.din(n10088), .dout(n10091));
    jdff dff_B_ofiOtxJx9_3(.din(n10091), .dout(n10094));
    jdff dff_B_12GJp60D6_3(.din(n10094), .dout(n10097));
    jdff dff_B_tCs5qjH55_3(.din(n10097), .dout(n10100));
    jdff dff_B_FlfoBxZO6_3(.din(n10100), .dout(n10103));
    jdff dff_B_et4NPvVk8_3(.din(n10103), .dout(n10106));
    jdff dff_B_85JHcCmn5_3(.din(n10106), .dout(n10109));
    jdff dff_B_8iLpfF7G6_3(.din(n10109), .dout(n10112));
    jdff dff_B_93hIVo6c5_3(.din(n10112), .dout(n10115));
    jdff dff_B_GwLzA4Vi2_3(.din(n10115), .dout(n10118));
    jdff dff_B_ICQHecuV9_3(.din(n10118), .dout(n10121));
    jdff dff_B_wWZk4Lds0_1(.din(n4503), .dout(n10124));
    jdff dff_B_wJv8Z09L0_1(.din(n10124), .dout(n10127));
    jdff dff_B_KGtdqV2A3_1(.din(n10127), .dout(n10130));
    jdff dff_B_5tREL57K7_1(.din(n10130), .dout(n10133));
    jdff dff_B_RF5t2aVj9_1(.din(n10133), .dout(n10136));
    jdff dff_B_WcJaMcar2_1(.din(n10136), .dout(n10139));
    jdff dff_B_LQia12gc9_1(.din(n10139), .dout(n10142));
    jdff dff_B_feOQWGXI5_0(.din(n4559), .dout(n10145));
    jdff dff_B_9nxREcP01_0(.din(n10145), .dout(n10148));
    jdff dff_B_GBOVEWZc9_0(.din(n10148), .dout(n10151));
    jdff dff_B_yZhpUOE74_0(.din(n10151), .dout(n10154));
    jdff dff_B_q5H8wVDo8_0(.din(n10154), .dout(n10157));
    jdff dff_B_4SapPi330_0(.din(n10157), .dout(n10160));
    jdff dff_B_qSPEZmw36_0(.din(n10160), .dout(n10163));
    jdff dff_B_PKJyVjaC7_0(.din(n10163), .dout(n10166));
    jdff dff_B_1pLUySZd3_0(.din(n10166), .dout(n10169));
    jdff dff_B_qZd0qqtg9_0(.din(n10169), .dout(n10172));
    jdff dff_B_zb3Fl8IE9_0(.din(n10172), .dout(n10175));
    jdff dff_B_nBniW0zQ0_0(.din(n10175), .dout(n10178));
    jdff dff_B_oQY7Vf4N0_0(.din(n10178), .dout(n10181));
    jdff dff_B_hvJq30dk8_0(.din(n10181), .dout(n10184));
    jdff dff_B_NDmSaG2h9_0(.din(n10184), .dout(n10187));
    jdff dff_B_9Ijh9dG00_0(.din(n10187), .dout(n10190));
    jdff dff_B_TK2VkFiS0_0(.din(n4762), .dout(n10193));
    jdff dff_B_12HAZl668_0(.din(n10193), .dout(n10196));
    jdff dff_B_oSPfDfeT1_0(.din(n4758), .dout(n10199));
    jdff dff_B_3A12Cw1k7_0(.din(n10199), .dout(n10202));
    jdff dff_B_1NZYUUDW3_0(.din(n10202), .dout(n10205));
    jdff dff_B_DxnJ7JMd7_0(.din(n10205), .dout(n10208));
    jdff dff_B_ruU84gPK4_0(.din(n10208), .dout(n10211));
    jdff dff_B_D5dEVWu88_0(.din(n10211), .dout(n10214));
    jdff dff_B_8vozDF7V2_0(.din(n10214), .dout(n10217));
    jdff dff_B_5qcoIMpU2_0(.din(n10217), .dout(n10220));
    jdff dff_B_Ca4LTnJZ4_0(.din(n10220), .dout(n10223));
    jdff dff_B_gIhRgRjM1_0(.din(n10223), .dout(n10226));
    jdff dff_B_Zt8ILZVx8_0(.din(n10226), .dout(n10229));
    jdff dff_B_gUUhPHdx0_0(.din(n10229), .dout(n10232));
    jdff dff_B_mhhPRSfj5_0(.din(n10232), .dout(n10235));
    jdff dff_B_x2Z9RvSJ7_0(.din(n10235), .dout(n10238));
    jdff dff_B_ElOjTrJk8_0(.din(n10238), .dout(n10241));
    jdff dff_B_6a3XpskK7_0(.din(n10241), .dout(n10244));
    jdff dff_B_bLwZTJWi7_0(.din(n10244), .dout(n10247));
    jdff dff_B_OUDgAJoO4_0(.din(n10247), .dout(n10250));
    jdff dff_B_rwukpntz1_0(.din(n10250), .dout(n10253));
    jdff dff_B_9FbwB4DN9_0(.din(n10253), .dout(n10256));
    jdff dff_B_4EJ33MHl7_0(.din(n10256), .dout(n10259));
    jdff dff_B_reTKQ3Mt8_0(.din(n10259), .dout(n10262));
    jdff dff_B_GQZn4cF11_0(.din(n10262), .dout(n10265));
    jdff dff_B_AXN5zYGA4_0(.din(n10265), .dout(n10268));
    jdff dff_B_2738FR838_0(.din(n4746), .dout(n10271));
    jdff dff_B_mQA7HCfO5_0(.din(n10271), .dout(n10274));
    jdff dff_B_8fkx1HXv7_0(.din(n10274), .dout(n10277));
    jdff dff_B_HGeN4flO9_0(.din(n10277), .dout(n10280));
    jdff dff_B_u2t1JI6M1_0(.din(n10280), .dout(n10283));
    jdff dff_B_Jbq6DmhX3_0(.din(n10283), .dout(n10286));
    jdff dff_B_rqNvkiyT5_0(.din(n10286), .dout(n10289));
    jdff dff_B_80hPncZ95_0(.din(n10289), .dout(n10292));
    jdff dff_B_S7F6LStF1_0(.din(n10292), .dout(n10295));
    jdff dff_B_BRMmmpfL0_0(.din(n10295), .dout(n10298));
    jdff dff_B_nRPVgKWW5_0(.din(n10298), .dout(n10301));
    jdff dff_B_8kAVW8gB0_0(.din(n10301), .dout(n10304));
    jdff dff_B_GmWRTMoa6_0(.din(n10304), .dout(n10307));
    jdff dff_B_d4kiu3Y44_0(.din(n10307), .dout(n10310));
    jdff dff_B_GfyjoT731_0(.din(n10310), .dout(n10313));
    jdff dff_B_hephm8TV5_0(.din(n4742), .dout(n10316));
    jdff dff_B_mxWw4cXU4_0(.din(n4726), .dout(n10319));
    jdff dff_B_JFGY0C2l5_0(.din(n4710), .dout(n10322));
    jdff dff_B_ACIfsFgv6_0(.din(n10322), .dout(n10325));
    jdff dff_B_oAbW667H2_0(.din(n10325), .dout(n10328));
    jdff dff_B_Rsfrln7j2_0(.din(n10328), .dout(n10331));
    jdff dff_B_8IkfZdUQ2_0(.din(n10331), .dout(n10334));
    jdff dff_B_jZ7TKH3V2_0(.din(n10334), .dout(n10337));
    jdff dff_B_ICu2GORB2_0(.din(n10337), .dout(n10340));
    jdff dff_B_dNevHoGM4_0(.din(n10340), .dout(n10343));
    jdff dff_B_W25aDOCw2_0(.din(n10343), .dout(n10346));
    jdff dff_B_uJpGYrPR3_0(.din(n10346), .dout(n10349));
    jdff dff_B_7mnuJ1KH0_0(.din(n10349), .dout(n10352));
    jdff dff_B_s4mshVr45_0(.din(n10352), .dout(n10355));
    jdff dff_B_INOpmN2v9_0(.din(n10355), .dout(n10358));
    jdff dff_B_PL1JEJ9U9_1(.din(n4657), .dout(n10361));
    jdff dff_B_1FyWNS501_0(.din(n4702), .dout(n10364));
    jdff dff_B_NozrAiAC0_0(.din(n10364), .dout(n10367));
    jdff dff_B_b9b3rXR82_0(.din(n10367), .dout(n10370));
    jdff dff_B_KYND4Y7A2_0(.din(n4694), .dout(n10373));
    jdff dff_B_ew9BjGEv2_1(.din(n4665), .dout(n10376));
    jdff dff_B_8MmWqEbC1_1(.din(n10376), .dout(n10379));
    jdff dff_B_yv0IKcgm6_0(.din(n4668), .dout(n10382));
    jdff dff_B_N2OCdIRW9_0(.din(n10382), .dout(n10385));
    jdff dff_B_xpKKAL3M3_0(.din(n10385), .dout(n10388));
    jdff dff_B_lc2rTYBf5_0(.din(n10388), .dout(n10391));
    jdff dff_A_719EER1D0_0(.din(n10396), .dout(n10393));
    jdff dff_A_OjBgAxHs3_0(.din(n10399), .dout(n10396));
    jdff dff_A_W0PFkf9e6_0(.din(n10402), .dout(n10399));
    jdff dff_A_TtsvZyKe2_0(.din(n4661), .dout(n10402));
    jdff dff_A_gbJB54ha2_2(.din(n10408), .dout(n10405));
    jdff dff_A_PzrwB98c9_2(.din(n10411), .dout(n10408));
    jdff dff_A_7oZDXmlx4_2(.din(n4661), .dout(n10411));
    jdff dff_A_krkk7XAh3_1(.din(n10487), .dout(n10414));
    jdff dff_A_aBj6fkYF0_2(.din(n10420), .dout(n10417));
    jdff dff_A_2zKwrxka1_2(.din(n10423), .dout(n10420));
    jdff dff_A_HUrhjDSj0_2(.din(n10426), .dout(n10423));
    jdff dff_A_beI3AcAP1_2(.din(n10429), .dout(n10426));
    jdff dff_A_QhrjhUhk6_2(.din(n10432), .dout(n10429));
    jdff dff_A_5r8eP85j4_2(.din(n10435), .dout(n10432));
    jdff dff_A_WEP0MKFF0_2(.din(n10438), .dout(n10435));
    jdff dff_A_YrUKhixG1_2(.din(n10441), .dout(n10438));
    jdff dff_A_eIOkxsDs3_2(.din(n10444), .dout(n10441));
    jdff dff_A_q5O3GhCj0_2(.din(n10447), .dout(n10444));
    jdff dff_A_LsF4A0HY3_2(.din(n10450), .dout(n10447));
    jdff dff_A_jtg43NQK5_2(.din(n10453), .dout(n10450));
    jdff dff_A_7yNIHFGd2_2(.din(n10456), .dout(n10453));
    jdff dff_A_QcorbPoi1_2(.din(n10459), .dout(n10456));
    jdff dff_A_ePWatc187_2(.din(n10462), .dout(n10459));
    jdff dff_A_XQE8hrzm9_2(.din(n10465), .dout(n10462));
    jdff dff_A_gUPboYWa9_2(.din(n10468), .dout(n10465));
    jdff dff_A_t7SZ7ibq3_2(.din(n10471), .dout(n10468));
    jdff dff_A_i00KGOL32_2(.din(n10474), .dout(n10471));
    jdff dff_A_HvtO3RM12_2(.din(n10477), .dout(n10474));
    jdff dff_A_jJI5G6gM5_2(.din(n10487), .dout(n10477));
    jdff dff_B_VayDGo799_3(.din(n4239), .dout(n10481));
    jdff dff_B_rDo5NBVx2_3(.din(n10481), .dout(n10484));
    jdff dff_B_tof5vAxJ8_3(.din(n10484), .dout(n10487));
    jdff dff_B_ijaMgSks0_0(.din(n4641), .dout(n10490));
    jdff dff_B_3rEMfBpF3_0(.din(n10490), .dout(n10493));
    jdff dff_B_hK5XbLPc3_0(.din(n10493), .dout(n10496));
    jdff dff_B_bzBj97qH0_0(.din(n10496), .dout(n10499));
    jdff dff_B_GAaUEI6x9_0(.din(n10499), .dout(n10502));
    jdff dff_B_Mv1xrPiQ3_0(.din(n10502), .dout(n10505));
    jdff dff_B_r8l9RA577_0(.din(n10505), .dout(n10508));
    jdff dff_B_ChH0EEBX8_0(.din(n10508), .dout(n10511));
    jdff dff_B_BSKntXx67_0(.din(n10511), .dout(n10514));
    jdff dff_B_77aDa9LM9_0(.din(n10514), .dout(n10517));
    jdff dff_B_UtGWPSW14_0(.din(n10517), .dout(n10520));
    jdff dff_B_B4SL31yq2_0(.din(n10520), .dout(n10523));
    jdff dff_B_zfRgEin34_0(.din(n10523), .dout(n10526));
    jdff dff_B_86m7VksF8_0(.din(n10526), .dout(n10529));
    jdff dff_B_5avHTFlS5_0(.din(n10529), .dout(n10532));
    jdff dff_B_UAJSjZ4p4_0(.din(n10532), .dout(n10535));
    jdff dff_B_xP21tEYM0_0(.din(n10535), .dout(n10538));
    jdff dff_B_fYPvapMd8_0(.din(n10538), .dout(n10541));
    jdff dff_B_NGsbwMpe2_0(.din(n10541), .dout(n10544));
    jdff dff_B_4HAgZNzg2_1(.din(n4633), .dout(n10547));
    jdff dff_B_nuGxlRcY6_0(.din(n4629), .dout(n10550));
    jdff dff_B_V51AO53A2_0(.din(n10550), .dout(n10553));
    jdff dff_B_pUYv3kJb8_0(.din(n4617), .dout(n10556));
    jdff dff_B_8p8f9pN02_0(.din(n4606), .dout(n10559));
    jdff dff_B_eDA1cr683_0(.din(n10559), .dout(n10562));
    jdff dff_B_2NVuRVOw5_0(.din(n10562), .dout(n10565));
    jdff dff_B_Hr4UWyl12_0(.din(n10565), .dout(n10568));
    jdff dff_B_CXgMz9647_0(.din(n10568), .dout(n10571));
    jdff dff_B_OERe5ODg6_0(.din(n10571), .dout(n10574));
    jdff dff_B_ImMSh5TZ2_0(.din(n10574), .dout(n10577));
    jdff dff_B_QaXdQIWl1_0(.din(n10577), .dout(n10580));
    jdff dff_B_1YZVfkZN3_0(.din(n10580), .dout(n10583));
    jdff dff_B_6rUDTuxD3_0(.din(n10583), .dout(n10586));
    jdff dff_B_6lcabkyl5_0(.din(n10586), .dout(n10589));
    jdff dff_B_YhVmrNL97_0(.din(n10589), .dout(n10592));
    jdff dff_B_mSlToNXx6_0(.din(n10592), .dout(n10595));
    jdff dff_B_MefwuRR94_0(.din(n10595), .dout(n10598));
    jdff dff_B_3xR3Qjsu8_0(.din(n10598), .dout(n10601));
    jdff dff_B_wgTQbKLv9_0(.din(n10601), .dout(n10604));
    jdff dff_B_MG03m1yT9_0(.din(n10604), .dout(n10607));
    jdff dff_B_hYjjC3xx1_0(.din(n10607), .dout(n10610));
    jdff dff_B_kGTsVbyO2_0(.din(n10610), .dout(n10613));
    jdff dff_B_bZewYbaQ4_0(.din(n4602), .dout(n10616));
    jdff dff_B_Jyi5VW8h0_1(.din(n4583), .dout(n10619));
    jdff dff_A_ND9Xw4v67_1(.din(n10624), .dout(n10621));
    jdff dff_A_x46G1Kg41_1(.din(n10627), .dout(n10624));
    jdff dff_A_mBJj3KzO0_1(.din(n10630), .dout(n10627));
    jdff dff_A_YbNCaeJ37_1(.din(n10633), .dout(n10630));
    jdff dff_A_oTD6dlzB2_1(.din(n10636), .dout(n10633));
    jdff dff_A_OgqFqi3b7_1(.din(n10639), .dout(n10636));
    jdff dff_A_Ou7NyWKl8_1(.din(n10642), .dout(n10639));
    jdff dff_A_Y6s8OPQO9_1(.din(n10645), .dout(n10642));
    jdff dff_A_2VYW4K1v6_1(.din(n10648), .dout(n10645));
    jdff dff_A_7fH6kUON8_1(.din(n10651), .dout(n10648));
    jdff dff_A_cevX7o0u9_1(.din(n10654), .dout(n10651));
    jdff dff_A_b4P4GOG36_1(.din(n10657), .dout(n10654));
    jdff dff_A_tEyVDrMj6_1(.din(n10660), .dout(n10657));
    jdff dff_A_zVfKWdjQ9_1(.din(n10663), .dout(n10660));
    jdff dff_A_CAAk2uRn9_1(.din(n10666), .dout(n10663));
    jdff dff_A_PIqAJi5a8_1(.din(n10669), .dout(n10666));
    jdff dff_A_3NmO94mg2_1(.din(n10672), .dout(n10669));
    jdff dff_A_3IP9oUZD1_1(.din(n10675), .dout(n10672));
    jdff dff_A_qc6uFhI29_1(.din(n10678), .dout(n10675));
    jdff dff_A_fQOs5RJI0_1(.din(n10681), .dout(n10678));
    jdff dff_A_cHkkuZrw5_1(.din(n10684), .dout(n10681));
    jdff dff_A_yBrlKAMT0_1(.din(n10687), .dout(n10684));
    jdff dff_A_L37J9nCp5_1(.din(n10690), .dout(n10687));
    jdff dff_A_Xlj8jfvv7_1(.din(n10693), .dout(n10690));
    jdff dff_A_LPFnN2Nq5_1(.din(n4424), .dout(n10693));
    jdff dff_A_UTUX7qT57_0(.din(n10699), .dout(n10696));
    jdff dff_A_aqmJyNgr3_0(.din(n4421), .dout(n10699));
    jdff dff_B_M4BynVLC9_2(.din(n4579), .dout(n10703));
    jdff dff_B_cUsg1qKh9_2(.din(n10703), .dout(n10706));
    jdff dff_B_0E7z0d090_2(.din(n10706), .dout(n10709));
    jdff dff_B_34c1KuyF5_2(.din(n10709), .dout(n10712));
    jdff dff_B_7Lz0IC683_0(.din(n4948), .dout(n10715));
    jdff dff_B_Tq42sKlL7_0(.din(n4940), .dout(n10718));
    jdff dff_B_QJJewbSj4_0(.din(n10718), .dout(n10721));
    jdff dff_B_1AgZ3Bjn8_0(.din(n10721), .dout(n10724));
    jdff dff_B_whGa9iPH5_0(.din(n10724), .dout(n10727));
    jdff dff_B_1AnSKQfI2_0(.din(n10727), .dout(n10730));
    jdff dff_B_REgLsSAk6_0(.din(n10730), .dout(n10733));
    jdff dff_B_yoFNMVqF6_0(.din(n10733), .dout(n10736));
    jdff dff_B_LO8MsGPn6_0(.din(n10736), .dout(n10739));
    jdff dff_B_MPZomksl0_0(.din(n10739), .dout(n10742));
    jdff dff_B_qPloL37m9_0(.din(n10742), .dout(n10745));
    jdff dff_B_EQRiOYtZ7_0(.din(n10745), .dout(n10748));
    jdff dff_B_5qvJ2mKi1_0(.din(n10748), .dout(n10751));
    jdff dff_B_VEzlivPG9_0(.din(n10751), .dout(n10754));
    jdff dff_B_luoQV8yu9_0(.din(n10754), .dout(n10757));
    jdff dff_B_l96kWJPL1_0(.din(n10757), .dout(n10760));
    jdff dff_B_lT3Pp4zg7_0(.din(n10760), .dout(n10763));
    jdff dff_B_JykNhceB1_0(.din(n10763), .dout(n10766));
    jdff dff_B_JwRnG0pd9_0(.din(n4936), .dout(n10769));
    jdff dff_A_8AxGSzgb4_1(.din(n10774), .dout(n10771));
    jdff dff_A_GAnxm2I85_1(.din(n10777), .dout(n10774));
    jdff dff_A_t9iASt3X5_1(.din(n10780), .dout(n10777));
    jdff dff_A_zV6UWLfI6_1(.din(n10783), .dout(n10780));
    jdff dff_A_7y77P9SC0_1(.din(n10786), .dout(n10783));
    jdff dff_A_2RVeAT833_1(.din(n10789), .dout(n10786));
    jdff dff_A_e9Go8sPr9_1(.din(n10792), .dout(n10789));
    jdff dff_A_HxTrJinE0_1(.din(n10795), .dout(n10792));
    jdff dff_A_nYkfMcrM3_1(.din(n10798), .dout(n10795));
    jdff dff_A_hbPUZvC87_1(.din(n10801), .dout(n10798));
    jdff dff_A_OZqdLF5D0_1(.din(n10804), .dout(n10801));
    jdff dff_A_dEH2fRdO4_1(.din(n10807), .dout(n10804));
    jdff dff_A_aspEWJ8J4_1(.din(n10810), .dout(n10807));
    jdff dff_A_UPBiKVTm1_1(.din(n10813), .dout(n10810));
    jdff dff_A_mxFMN0K67_1(.din(n10816), .dout(n10813));
    jdff dff_A_r997vqh18_1(.din(n10819), .dout(n10816));
    jdff dff_A_en48fLNx7_1(.din(n10822), .dout(n10819));
    jdff dff_A_eIgdf5oS8_1(.din(n10825), .dout(n10822));
    jdff dff_A_b6NpkqnL3_1(.din(n10828), .dout(n10825));
    jdff dff_A_l9fYWk477_1(.din(n10831), .dout(n10828));
    jdff dff_A_keEUnYQ00_1(.din(n698), .dout(n10831));
    jdff dff_A_M7KmyMdH9_0(.din(n10837), .dout(n10834));
    jdff dff_A_tpY9nJRG5_0(.din(n10840), .dout(n10837));
    jdff dff_A_FNA0fCSX4_0(.din(n10843), .dout(n10840));
    jdff dff_A_cnEMWUXq2_0(.din(n10846), .dout(n10843));
    jdff dff_A_JkaivZjF0_0(.din(n10849), .dout(n10846));
    jdff dff_A_OEgsPleW8_0(.din(n10852), .dout(n10849));
    jdff dff_A_l1KiWBJ80_0(.din(n10855), .dout(n10852));
    jdff dff_A_7L673EWa7_0(.din(n10858), .dout(n10855));
    jdff dff_A_QgYzijuN2_0(.din(n10861), .dout(n10858));
    jdff dff_A_Edtt8bzm2_0(.din(n10864), .dout(n10861));
    jdff dff_A_bcSouc1D2_0(.din(n10867), .dout(n10864));
    jdff dff_A_36YJjSOi8_0(.din(n10870), .dout(n10867));
    jdff dff_A_cC7PaEWc9_0(.din(n10873), .dout(n10870));
    jdff dff_A_CaRJ8C2P2_0(.din(n10876), .dout(n10873));
    jdff dff_A_AR8wxLEs0_0(.din(n10879), .dout(n10876));
    jdff dff_A_Uv5lnRWA8_0(.din(n10882), .dout(n10879));
    jdff dff_A_iMxzCyTs2_0(.din(n10885), .dout(n10882));
    jdff dff_A_xpiY8Ufd5_0(.din(n10888), .dout(n10885));
    jdff dff_A_liH9GRf56_0(.din(n10891), .dout(n10888));
    jdff dff_A_9gO6g7tX7_0(.din(n10894), .dout(n10891));
    jdff dff_A_msS3zn0b7_0(.din(n670), .dout(n10894));
    jdff dff_B_OnYKiijy7_1(.din(n4928), .dout(n10898));
    jdff dff_B_BwhpK7Re8_1(.din(n10898), .dout(n10901));
    jdff dff_B_u7raKxTd3_1(.din(n10901), .dout(n10904));
    jdff dff_B_p95jurqh9_1(.din(n10904), .dout(n10907));
    jdff dff_B_rIxcZSoR5_1(.din(n10907), .dout(n10910));
    jdff dff_B_i4G7rVJD8_1(.din(n10910), .dout(n10913));
    jdff dff_B_28qkGFQB2_1(.din(n10913), .dout(n10916));
    jdff dff_A_UHdhm1WF6_1(.din(n10921), .dout(n10918));
    jdff dff_A_ThXDYTK74_1(.din(n10924), .dout(n10921));
    jdff dff_A_wahFABi94_1(.din(n10927), .dout(n10924));
    jdff dff_A_qhGdko7W8_1(.din(n10930), .dout(n10927));
    jdff dff_A_oh1B2yho0_1(.din(n10933), .dout(n10930));
    jdff dff_A_StSoeVLD8_1(.din(n694), .dout(n10933));
    jdff dff_B_oiF3CoFo6_0(.din(n4921), .dout(n10937));
    jdff dff_B_K5OSU1ID5_0(.din(n10937), .dout(n10940));
    jdff dff_B_uYuGoqJ38_0(.din(n10940), .dout(n10943));
    jdff dff_B_5A1JMwbV0_0(.din(n10943), .dout(n10946));
    jdff dff_B_Bib73DXc3_0(.din(n10946), .dout(n10949));
    jdff dff_B_gxFZF1cC6_0(.din(n10949), .dout(n10952));
    jdff dff_B_T1a1nCr90_0(.din(n10952), .dout(n10955));
    jdff dff_B_cmmUvgXQ2_0(.din(n10955), .dout(n10958));
    jdff dff_B_VcA1N3op7_0(.din(n10958), .dout(n10961));
    jdff dff_B_DpD6zRwG4_0(.din(n10961), .dout(n10964));
    jdff dff_B_9EtzbZrf0_0(.din(n10964), .dout(n10967));
    jdff dff_B_shyeRnQy5_0(.din(n10967), .dout(n10970));
    jdff dff_B_SzAEIMD45_0(.din(n10970), .dout(n10973));
    jdff dff_B_Dkxpceow1_0(.din(n10973), .dout(n10976));
    jdff dff_B_ir71D0UF7_0(.din(n10976), .dout(n10979));
    jdff dff_B_6iJ4ZQlC5_0(.din(n10979), .dout(n10982));
    jdff dff_B_R6auYvqy2_0(.din(n10982), .dout(n10985));
    jdff dff_B_Nrh579qe2_0(.din(n10985), .dout(n10988));
    jdff dff_B_iVnIzRsb0_1(.din(n4894), .dout(n10991));
    jdff dff_B_rUCszkdl1_0(.din(n4913), .dout(n10994));
    jdff dff_B_IKQhlY9y6_0(.din(n10994), .dout(n10997));
    jdff dff_B_RGnY6viN6_0(.din(n10997), .dout(n11000));
    jdff dff_B_sJYrScQ83_0(.din(n11000), .dout(n11003));
    jdff dff_B_YpX15TpO5_0(.din(n11003), .dout(n11006));
    jdff dff_B_1MTnPnjM5_0(.din(n11006), .dout(n11009));
    jdff dff_B_9wr4v2i46_0(.din(n11009), .dout(n11012));
    jdff dff_B_7M0PEGo79_0(.din(n11012), .dout(n11015));
    jdff dff_B_myCTkUXi8_0(.din(n11015), .dout(n11018));
    jdff dff_A_QNIvOtTH5_2(.din(n496), .dout(n11020));
    jdff dff_A_4pDBzIkj8_0(.din(n477), .dout(n11023));
    jdff dff_A_AoXjLKEa2_0(.din(n11029), .dout(n11026));
    jdff dff_A_0RqgLhFE7_0(.din(G38), .dout(n11029));
    jdff dff_A_AV8fO8in9_1(.din(G38), .dout(n11032));
    jdff dff_A_GEC2RqG04_0(.din(n11060), .dout(n11035));
    jdff dff_B_k6xiZitH3_2(.din(n4890), .dout(n11039));
    jdff dff_B_h91Oegy59_2(.din(n11039), .dout(n11042));
    jdff dff_B_ceZN13d44_2(.din(n11042), .dout(n11045));
    jdff dff_B_gItFd5wj3_2(.din(n11045), .dout(n11048));
    jdff dff_B_UaCCBgEI4_2(.din(n11048), .dout(n11051));
    jdff dff_B_6cX0yVnW7_2(.din(n11051), .dout(n11054));
    jdff dff_B_yeZl5t8Z9_2(.din(n11054), .dout(n11057));
    jdff dff_B_n59tdYKQ9_2(.din(n11057), .dout(n11060));
    jdff dff_B_GB5UhtBF0_1(.din(n4879), .dout(n11063));
    jdff dff_A_JsrNYtsM8_0(.din(n11068), .dout(n11065));
    jdff dff_A_XrVfKjOm6_0(.din(n489), .dout(n11068));
    jdff dff_A_HXEhRKtJ6_2(.din(n11074), .dout(n11071));
    jdff dff_A_TygEWVQm6_2(.din(n11077), .dout(n11074));
    jdff dff_A_om8WZW3x7_2(.din(G1496), .dout(n11077));
    jdff dff_A_jj8FWGRv1_0(.din(G1492), .dout(n11080));
    jdff dff_A_5EyIJLb49_2(.din(n11086), .dout(n11083));
    jdff dff_A_z84Sivjb7_2(.din(n11089), .dout(n11086));
    jdff dff_A_0Ti9dv7b3_2(.din(G1492), .dout(n11089));
    jdff dff_A_FQOPaHzv0_0(.din(G38), .dout(n11092));
    jdff dff_A_sWXvFQX26_2(.din(G38), .dout(n11095));
    jdff dff_B_kXl7AKD53_1(.din(n533), .dout(n11099));
    jdff dff_B_gXPd4Jwn9_1(.din(n11099), .dout(n11102));
    jdff dff_B_skhcZKns8_1(.din(n11102), .dout(n11105));
    jdff dff_B_3MxGaw4F7_1(.din(n11105), .dout(n11108));
    jdff dff_B_1leuiOL64_1(.din(n11108), .dout(n11111));
    jdff dff_B_6za001C86_1(.din(n11111), .dout(n11114));
    jdff dff_B_1VpL3ITN8_1(.din(n11114), .dout(n11117));
    jdff dff_B_GP6CBlmT3_1(.din(n11117), .dout(n11120));
    jdff dff_A_2scM1JL69_0(.din(n11125), .dout(n11122));
    jdff dff_A_HT7AMlND8_0(.din(n11128), .dout(n11125));
    jdff dff_A_3ny3aAEH1_0(.din(n11131), .dout(n11128));
    jdff dff_A_Wp3jAbI40_0(.din(n11134), .dout(n11131));
    jdff dff_A_5spAxOzI6_0(.din(n11137), .dout(n11134));
    jdff dff_A_19uBMY4k7_0(.din(n11140), .dout(n11137));
    jdff dff_A_7ylir7V19_0(.din(n11143), .dout(n11140));
    jdff dff_A_clLEDIGw9_0(.din(n11146), .dout(n11143));
    jdff dff_A_ePeB584u3_0(.din(n11149), .dout(n11146));
    jdff dff_A_CT1Zwr7E6_0(.din(n11152), .dout(n11149));
    jdff dff_A_NA3emlrz5_0(.din(n11155), .dout(n11152));
    jdff dff_A_1tUvtlUT3_0(.din(n11158), .dout(n11155));
    jdff dff_A_7EcG6Nh41_0(.din(n11161), .dout(n11158));
    jdff dff_A_4n9Cq2BZ1_0(.din(n11164), .dout(n11161));
    jdff dff_A_xbcpzsOe3_0(.din(n11167), .dout(n11164));
    jdff dff_A_pWnRGosz6_0(.din(n11170), .dout(n11167));
    jdff dff_A_Nfs8BZD57_0(.din(n11173), .dout(n11170));
    jdff dff_A_fVC9dVDB5_0(.din(n11176), .dout(n11173));
    jdff dff_A_9jIclCX84_0(.din(n11179), .dout(n11176));
    jdff dff_A_G9eBYFVB8_0(.din(n11182), .dout(n11179));
    jdff dff_A_73VINfOf7_0(.din(n11185), .dout(n11182));
    jdff dff_A_q4Rcgtd79_0(.din(n11188), .dout(n11185));
    jdff dff_A_VuJDRYHz4_0(.din(n11191), .dout(n11188));
    jdff dff_A_PFxXQQEF3_0(.din(n11194), .dout(n11191));
    jdff dff_A_biG1YBpe4_0(.din(n11197), .dout(n11194));
    jdff dff_A_UOo25iMB9_0(.din(n11200), .dout(n11197));
    jdff dff_A_2DWOwWGn1_0(.din(n11203), .dout(n11200));
    jdff dff_A_otJcy7zp3_0(.din(n11206), .dout(n11203));
    jdff dff_A_P3Kbsd9q8_0(.din(n11209), .dout(n11206));
    jdff dff_A_9QatQ9tk9_0(.din(n12676), .dout(n11209));
    jdff dff_A_SiChp53D2_2(.din(n11215), .dout(n11212));
    jdff dff_A_OpQKdVDa4_2(.din(n11218), .dout(n11215));
    jdff dff_A_CsClAuT21_2(.din(n11221), .dout(n11218));
    jdff dff_A_iNggLAeh1_2(.din(n11224), .dout(n11221));
    jdff dff_A_khjwgLvX2_2(.din(n12676), .dout(n11224));
    jdff dff_B_4URZCTKT2_1(.din(n4770), .dout(n11228));
    jdff dff_B_IIRAvDTi4_1(.din(n11228), .dout(n11231));
    jdff dff_B_H9669h9Z1_1(.din(n11231), .dout(n11234));
    jdff dff_B_XCrdcWAr7_1(.din(n11234), .dout(n11237));
    jdff dff_B_MScwB68L7_1(.din(n11237), .dout(n11240));
    jdff dff_B_n5I8J8zb3_1(.din(n11240), .dout(n11243));
    jdff dff_B_VecfdJva2_1(.din(n11243), .dout(n11246));
    jdff dff_B_lmdSCRQa8_1(.din(n11246), .dout(n11249));
    jdff dff_B_dQLeCAFX5_1(.din(n11249), .dout(n11252));
    jdff dff_B_52g9Ls848_1(.din(n11252), .dout(n11255));
    jdff dff_B_NATieFFa3_1(.din(n11255), .dout(n11258));
    jdff dff_B_2ZjSOoZk1_1(.din(n11258), .dout(n11261));
    jdff dff_B_K565x8eR5_1(.din(n11261), .dout(n11264));
    jdff dff_B_jJYMotSy6_1(.din(n11264), .dout(n11267));
    jdff dff_B_DPT6iVDN3_1(.din(n11267), .dout(n11270));
    jdff dff_B_2Rq562tP6_1(.din(n11270), .dout(n11273));
    jdff dff_B_v5OaJ4Ow5_1(.din(n11273), .dout(n11276));
    jdff dff_B_1eXPyZuP0_1(.din(n11276), .dout(n11279));
    jdff dff_B_2yN8lW562_1(.din(n11279), .dout(n11282));
    jdff dff_B_4bfEc6Q59_1(.din(n11282), .dout(n11285));
    jdff dff_B_iKOJSfaE1_1(.din(n11285), .dout(n11288));
    jdff dff_B_OBsVua4Z4_1(.din(n11288), .dout(n11291));
    jdff dff_B_dUJDzBcM6_1(.din(n11291), .dout(n11294));
    jdff dff_B_YoHRC7kQ1_1(.din(n11294), .dout(n11297));
    jdff dff_B_KUJFyn363_1(.din(n11297), .dout(n11300));
    jdff dff_B_a0A0R9iS4_1(.din(n11300), .dout(n11303));
    jdff dff_B_iBqu3Y7d7_1(.din(n11303), .dout(n11306));
    jdff dff_B_57n7TXKg3_1(.din(n11306), .dout(n11309));
    jdff dff_B_EzkNbk9Z3_1(.din(n11309), .dout(n11312));
    jdff dff_B_YaANBgLp9_1(.din(n11312), .dout(n11315));
    jdff dff_B_QwCIe8H74_1(.din(n11315), .dout(n11318));
    jdff dff_B_zAPGi7sQ9_0(.din(n4856), .dout(n11321));
    jdff dff_B_kpcEDEf08_0(.din(n11321), .dout(n11324));
    jdff dff_B_cxTFnbYF4_0(.din(n11324), .dout(n11327));
    jdff dff_B_uPPHhfSG4_0(.din(n11327), .dout(n11330));
    jdff dff_B_XK8ll53l8_0(.din(n11330), .dout(n11333));
    jdff dff_B_azRK4Jwg0_0(.din(n11333), .dout(n11336));
    jdff dff_B_QVinhlI20_0(.din(n11336), .dout(n11339));
    jdff dff_B_rawBPdkp5_0(.din(n11339), .dout(n11342));
    jdff dff_B_fexPNuMS8_0(.din(n11342), .dout(n11345));
    jdff dff_B_MaMLRemh2_0(.din(n11345), .dout(n11348));
    jdff dff_B_A901igYJ6_0(.din(n11348), .dout(n11351));
    jdff dff_B_dxs6qdP81_0(.din(n11351), .dout(n11354));
    jdff dff_B_LVMcigG42_0(.din(n11354), .dout(n11357));
    jdff dff_B_EOpICpsq9_0(.din(n11357), .dout(n11360));
    jdff dff_B_sA3whaAc2_0(.din(n11360), .dout(n11363));
    jdff dff_B_gvLAsJf49_0(.din(n11363), .dout(n11366));
    jdff dff_B_vfS4H3GJ8_0(.din(n11366), .dout(n11369));
    jdff dff_B_IU8FPb0D3_0(.din(n11369), .dout(n11372));
    jdff dff_B_3IfdK66J1_0(.din(n11372), .dout(n11375));
    jdff dff_B_AHUCtzZZ4_0(.din(n11375), .dout(n11378));
    jdff dff_B_VG3jWbMU3_1(.din(n4836), .dout(n11381));
    jdff dff_B_Wz9LiyGS3_1(.din(n11381), .dout(n11384));
    jdff dff_B_xStXXyDX5_0(.din(n4840), .dout(n11387));
    jdff dff_B_8C6OP5B58_0(.din(n11387), .dout(n11390));
    jdff dff_B_EkJW2d739_0(.din(n11390), .dout(n11393));
    jdff dff_B_GfHZKRgn0_0(.din(n11393), .dout(n11396));
    jdff dff_B_7TJ07BqD6_0(.din(n11396), .dout(n11399));
    jdff dff_A_FGO3VwDe7_1(.din(n11404), .dout(n11401));
    jdff dff_A_4GxBDFuK5_1(.din(n11407), .dout(n11404));
    jdff dff_A_9Dandry36_1(.din(n11410), .dout(n11407));
    jdff dff_A_WsZgq4ld1_1(.din(n11413), .dout(n11410));
    jdff dff_A_62agWQZ76_1(.din(n11416), .dout(n11413));
    jdff dff_A_AquFdCbi3_1(.din(n11419), .dout(n11416));
    jdff dff_A_FE4fiykW8_1(.din(n11422), .dout(n11419));
    jdff dff_A_pOPNpuih6_1(.din(n11425), .dout(n11422));
    jdff dff_A_A4OjkDoC9_1(.din(n11428), .dout(n11425));
    jdff dff_A_96IQSY3P0_1(.din(n11431), .dout(n11428));
    jdff dff_A_rcEpXCLT9_1(.din(n11434), .dout(n11431));
    jdff dff_A_FueC69Vb4_1(.din(n11437), .dout(n11434));
    jdff dff_A_VZSUXcJR1_1(.din(n11440), .dout(n11437));
    jdff dff_A_XdQMZGYT8_1(.din(n11443), .dout(n11440));
    jdff dff_A_KKXS9DGc4_1(.din(n11446), .dout(n11443));
    jdff dff_A_iEOT29u52_1(.din(n11449), .dout(n11446));
    jdff dff_A_xhJreGxM4_1(.din(n11452), .dout(n11449));
    jdff dff_A_5rZqYOZF2_1(.din(n11455), .dout(n11452));
    jdff dff_A_JMGaejtI5_1(.din(n11458), .dout(n11455));
    jdff dff_A_6kHtavVd7_1(.din(n11461), .dout(n11458));
    jdff dff_A_BtTuPcIS1_1(.din(n11464), .dout(n11461));
    jdff dff_A_VTtE4p5y2_1(.din(n11467), .dout(n11464));
    jdff dff_A_aMUHQ7Iu9_1(.din(n11470), .dout(n11467));
    jdff dff_A_G14UZ7Ts8_1(.din(n11473), .dout(n11470));
    jdff dff_A_xuCJl1nq8_1(.din(n4332), .dout(n11473));
    jdff dff_B_6dr2HROu8_0(.din(n4328), .dout(n11477));
    jdff dff_B_CJN2F4J86_0(.din(n11477), .dout(n11480));
    jdff dff_B_6Xm9GNkp1_0(.din(n11480), .dout(n11483));
    jdff dff_B_jvy3VoAt6_1(.din(n4825), .dout(n11486));
    jdff dff_B_iTP5sQCM5_1(.din(n11486), .dout(n11489));
    jdff dff_B_SFXMS2uJ4_1(.din(n11489), .dout(n11492));
    jdff dff_B_qVejruuc3_1(.din(n4828), .dout(n11495));
    jdff dff_B_zpFoqYh97_1(.din(n11495), .dout(n11498));
    jdff dff_A_qQNwmH5o6_1(.din(n11503), .dout(n11500));
    jdff dff_A_nVFKisTE2_1(.din(n11506), .dout(n11503));
    jdff dff_A_ktLMMZcL7_1(.din(n11509), .dout(n11506));
    jdff dff_A_SLotKsRL8_1(.din(n11512), .dout(n11509));
    jdff dff_A_EzpjlKyO6_1(.din(n11515), .dout(n11512));
    jdff dff_A_HfGWA7UL9_1(.din(n11518), .dout(n11515));
    jdff dff_A_hKV06LHL6_1(.din(n11521), .dout(n11518));
    jdff dff_A_7nE0DL139_1(.din(n11524), .dout(n11521));
    jdff dff_A_YmS8dCMC5_1(.din(n11527), .dout(n11524));
    jdff dff_A_UbIBYy1D3_1(.din(n11530), .dout(n11527));
    jdff dff_A_k0dx8DWQ3_1(.din(n11533), .dout(n11530));
    jdff dff_A_0m2DTqYc6_1(.din(n11536), .dout(n11533));
    jdff dff_A_TCvrdDZE9_1(.din(n11539), .dout(n11536));
    jdff dff_A_7Ayixigf7_1(.din(n11542), .dout(n11539));
    jdff dff_A_Iq0hghM34_1(.din(n11545), .dout(n11542));
    jdff dff_A_nYKAr1b15_1(.din(n11548), .dout(n11545));
    jdff dff_A_ARd6ITmS7_1(.din(n11551), .dout(n11548));
    jdff dff_A_GXlCHxSq3_1(.din(n11554), .dout(n11551));
    jdff dff_A_1i44VYq57_1(.din(n11557), .dout(n11554));
    jdff dff_A_xdS4xNOl2_1(.din(n11560), .dout(n11557));
    jdff dff_A_6GealkN51_1(.din(n11563), .dout(n11560));
    jdff dff_A_OQiWABd12_1(.din(n11567), .dout(n11563));
    jdff dff_B_H8oXmmA94_2(.din(n4312), .dout(n11567));
    jdff dff_A_nfikk4AQ6_0(.din(n11572), .dout(n11569));
    jdff dff_A_lkcE2c0P4_0(.din(n11575), .dout(n11572));
    jdff dff_A_qxMPcfHI4_0(.din(n11578), .dout(n11575));
    jdff dff_A_h4etcT9V1_0(.din(n11581), .dout(n11578));
    jdff dff_A_iWAGMO7h6_0(.din(n690), .dout(n11581));
    jdff dff_B_bFGdTcFl7_1(.din(n4182), .dout(n11585));
    jdff dff_B_uktRUa4U6_1(.din(n11585), .dout(n11588));
    jdff dff_B_yPB3bYIt8_1(.din(n11588), .dout(n11591));
    jdff dff_B_SnoR0ISc2_1(.din(n11591), .dout(n11594));
    jdff dff_B_a6kOW1KS8_1(.din(n11594), .dout(n11597));
    jdff dff_B_mZtiIKQf2_1(.din(n11597), .dout(n11600));
    jdff dff_B_pZ9D4wAW0_1(.din(n11600), .dout(n11603));
    jdff dff_B_GclWk9i40_1(.din(n11603), .dout(n11606));
    jdff dff_B_NEiHFAHC2_1(.din(n11606), .dout(n11609));
    jdff dff_B_aR29EeWm8_1(.din(n11609), .dout(n11612));
    jdff dff_B_URtq9owT4_1(.din(n11612), .dout(n11615));
    jdff dff_B_4g3291wX8_1(.din(n11615), .dout(n11618));
    jdff dff_B_X2fhvDj11_1(.din(n11618), .dout(n11621));
    jdff dff_B_JJ2mHynC8_1(.din(n11621), .dout(n11624));
    jdff dff_B_gUZoFocb4_1(.din(n11624), .dout(n11627));
    jdff dff_B_GFxji9EJ8_1(.din(n11627), .dout(n11630));
    jdff dff_B_HE4ZSF592_1(.din(n11630), .dout(n11633));
    jdff dff_B_48tK7MUN0_1(.din(n11633), .dout(n11636));
    jdff dff_B_Su3kwOrT5_1(.din(n11636), .dout(n11639));
    jdff dff_B_DkS7F9ki1_1(.din(n11639), .dout(n11642));
    jdff dff_B_OiLJXAWd0_1(.din(n11642), .dout(n11645));
    jdff dff_B_jet4qFZK3_1(.din(n11645), .dout(n11648));
    jdff dff_B_0LPA7P8j1_1(.din(n11648), .dout(n11651));
    jdff dff_B_lInV46iW7_1(.din(n11651), .dout(n11654));
    jdff dff_B_8xwmUzaQ2_1(.din(n11654), .dout(n11657));
    jdff dff_B_sn5wKndL8_1(.din(n11657), .dout(n11660));
    jdff dff_B_k4OnJtg44_1(.din(n11660), .dout(n11663));
    jdff dff_B_zmbOQOvP3_1(.din(n11663), .dout(n11666));
    jdff dff_B_U3fnmt7e9_1(.din(n4185), .dout(n11669));
    jdff dff_B_PXcm5kGH7_1(.din(n11669), .dout(n11672));
    jdff dff_B_Du06je7b1_1(.din(n11672), .dout(n11675));
    jdff dff_B_4e5OsMwi1_1(.din(n11675), .dout(n11678));
    jdff dff_B_Nt7kok2D2_1(.din(n11678), .dout(n11681));
    jdff dff_B_LHcp6NtL3_1(.din(n11681), .dout(n11684));
    jdff dff_B_s0BKhxcC7_1(.din(n11684), .dout(n11687));
    jdff dff_B_uXUOpUnp0_1(.din(n11687), .dout(n11690));
    jdff dff_B_IuDRgzOw6_1(.din(n11690), .dout(n11693));
    jdff dff_B_iX6HCfrX8_1(.din(n11693), .dout(n11696));
    jdff dff_B_TkAQmy2F6_1(.din(n11696), .dout(n11699));
    jdff dff_B_HZP9cHmN3_1(.din(n11699), .dout(n11702));
    jdff dff_B_SErHn3Co3_1(.din(n11702), .dout(n11705));
    jdff dff_B_a5KWdw619_1(.din(n11705), .dout(n11708));
    jdff dff_B_6nfR4x0N9_1(.din(n11708), .dout(n11711));
    jdff dff_B_oqP1e4z64_1(.din(n11711), .dout(n11714));
    jdff dff_B_HrBH1RxL0_1(.din(n11714), .dout(n11717));
    jdff dff_B_yxSWqYma7_1(.din(n11717), .dout(n11720));
    jdff dff_B_o8Emg5SK9_1(.din(n11720), .dout(n11723));
    jdff dff_B_Rktz6AM47_1(.din(n11723), .dout(n11726));
    jdff dff_B_0QIdrxkI4_1(.din(n11726), .dout(n11729));
    jdff dff_B_Cf7HDrTi8_1(.din(n11729), .dout(n11732));
    jdff dff_B_ZsIJhXav8_1(.din(n11732), .dout(n11735));
    jdff dff_B_MpGPcPli1_1(.din(n11735), .dout(n11738));
    jdff dff_B_QxqAoEww1_1(.din(n11738), .dout(n11741));
    jdff dff_B_usKxzaUL4_1(.din(n11741), .dout(n11744));
    jdff dff_B_vp9A2Y2X7_1(.din(n11744), .dout(n11747));
    jdff dff_B_cESwo7Oj0_1(.din(n4188), .dout(n11750));
    jdff dff_B_R69Topu95_1(.din(n11750), .dout(n11753));
    jdff dff_B_67skyuQZ3_1(.din(n11753), .dout(n11756));
    jdff dff_B_AxBhauOz4_1(.din(n11756), .dout(n11759));
    jdff dff_B_KEgrpVWj1_1(.din(n11759), .dout(n11762));
    jdff dff_B_8zSm99nB1_1(.din(n11762), .dout(n11765));
    jdff dff_B_gPFETUWy8_1(.din(n11765), .dout(n11768));
    jdff dff_B_BQXFmObV5_1(.din(n11768), .dout(n11771));
    jdff dff_B_pKtYLJ7Z5_1(.din(n11771), .dout(n11774));
    jdff dff_B_wV0BdER56_1(.din(n11774), .dout(n11777));
    jdff dff_B_JPv22FWC9_1(.din(n11777), .dout(n11780));
    jdff dff_B_XnJiykrU9_1(.din(n11780), .dout(n11783));
    jdff dff_B_FL6Sb9Lk6_1(.din(n11783), .dout(n11786));
    jdff dff_B_T0wtvQYU4_1(.din(n11786), .dout(n11789));
    jdff dff_B_cCF5SyOg4_1(.din(n11789), .dout(n11792));
    jdff dff_B_KX9axuSC7_1(.din(n11792), .dout(n11795));
    jdff dff_B_NOkpmACW8_1(.din(n11795), .dout(n11798));
    jdff dff_B_Jb6RIUga0_1(.din(n11798), .dout(n11801));
    jdff dff_B_vdkrFCYN1_1(.din(n11801), .dout(n11804));
    jdff dff_B_ZsqlCYh01_1(.din(n11804), .dout(n11807));
    jdff dff_B_rnCe3Ork8_1(.din(n11807), .dout(n11810));
    jdff dff_B_k128GXOQ4_1(.din(n4191), .dout(n11813));
    jdff dff_B_8v1f5lu64_1(.din(n11813), .dout(n11816));
    jdff dff_B_qDMTBvTM4_1(.din(n11816), .dout(n11819));
    jdff dff_B_RpTJ8ne29_1(.din(n11819), .dout(n11822));
    jdff dff_B_AshLw6qE3_1(.din(n11822), .dout(n11825));
    jdff dff_B_Tc9xDrxg9_1(.din(n11825), .dout(n11828));
    jdff dff_B_5mxyAtXC7_1(.din(n11828), .dout(n11831));
    jdff dff_B_nrRkeC0n1_1(.din(n11831), .dout(n11834));
    jdff dff_B_sJ1BlAHw3_1(.din(n11834), .dout(n11837));
    jdff dff_B_NgtP7nAb7_1(.din(n11837), .dout(n11840));
    jdff dff_B_rae1xR3N7_1(.din(n11840), .dout(n11843));
    jdff dff_B_IK8yuc0C4_1(.din(n11843), .dout(n11846));
    jdff dff_B_3kuzFPr53_1(.din(n11846), .dout(n11849));
    jdff dff_B_CyWgGN208_1(.din(n11849), .dout(n11852));
    jdff dff_B_NNvIj3sz2_1(.din(n11852), .dout(n11855));
    jdff dff_B_qnAH5L7I0_1(.din(n11855), .dout(n11858));
    jdff dff_B_RgWgAMLJ0_1(.din(n11858), .dout(n11861));
    jdff dff_B_Jrt6afgO4_1(.din(n11861), .dout(n11864));
    jdff dff_B_4gExAVhN2_1(.din(n11864), .dout(n11867));
    jdff dff_B_lwVZCQWe7_1(.din(n11867), .dout(n11870));
    jdff dff_B_nd1RsLIr9_1(.din(n11870), .dout(n11873));
    jdff dff_B_HCXKnUV56_1(.din(n4194), .dout(n11876));
    jdff dff_B_44gYAvYT5_1(.din(n11876), .dout(n11879));
    jdff dff_B_ODsjwKZU9_1(.din(n11879), .dout(n11882));
    jdff dff_B_ohRFURxK8_1(.din(n11882), .dout(n11885));
    jdff dff_B_hw8qqWUl6_1(.din(n11885), .dout(n11888));
    jdff dff_B_ZFrDDfpJ6_1(.din(n11888), .dout(n11891));
    jdff dff_B_D5IQZtkR1_1(.din(n11891), .dout(n11894));
    jdff dff_B_UPCU2CmB6_1(.din(n11894), .dout(n11897));
    jdff dff_B_u6yzwprT5_1(.din(n11897), .dout(n11900));
    jdff dff_B_BonRRWPv8_1(.din(n11900), .dout(n11903));
    jdff dff_B_77XlgZEc1_1(.din(n11903), .dout(n11906));
    jdff dff_B_Akr6oeE66_1(.din(n11906), .dout(n11909));
    jdff dff_B_D03abrMJ9_1(.din(n11909), .dout(n11912));
    jdff dff_B_8lvX44m70_1(.din(n11912), .dout(n11915));
    jdff dff_B_MQlJAE9M7_1(.din(n11915), .dout(n11918));
    jdff dff_B_NAgtVxZD0_1(.din(n11918), .dout(n11921));
    jdff dff_B_Y5YldpcH8_1(.din(n4197), .dout(n11924));
    jdff dff_B_DP4CX1mM1_1(.din(n11924), .dout(n11927));
    jdff dff_B_5tklbAaM3_1(.din(n11927), .dout(n11930));
    jdff dff_B_Byl5Z62t8_1(.din(n11930), .dout(n11933));
    jdff dff_B_ytgcOuN60_1(.din(n11933), .dout(n11936));
    jdff dff_B_0kADtmeq4_1(.din(n11936), .dout(n11939));
    jdff dff_B_u6FH1tbz5_1(.din(n11939), .dout(n11942));
    jdff dff_B_jW935lNA8_1(.din(n11942), .dout(n11945));
    jdff dff_B_rLGvwbtD6_1(.din(n11945), .dout(n11948));
    jdff dff_B_nlH3rkY76_1(.din(n11948), .dout(n11951));
    jdff dff_B_i7s5kYnd1_1(.din(n11951), .dout(n11954));
    jdff dff_B_wYoPpZ6N7_1(.din(n11954), .dout(n11957));
    jdff dff_B_YTdOoUHr3_1(.din(n11957), .dout(n11960));
    jdff dff_B_e52IBdTD4_1(.din(n11960), .dout(n11963));
    jdff dff_B_j0QpTQHF5_1(.din(n11963), .dout(n11966));
    jdff dff_B_TOdfTB2l7_1(.din(n11966), .dout(n11969));
    jdff dff_B_rHabs0Ds3_1(.din(n11969), .dout(n11972));
    jdff dff_B_xlnIwjUB5_1(.din(n4200), .dout(n11975));
    jdff dff_B_epeUJmat6_1(.din(n11975), .dout(n11978));
    jdff dff_B_3bOwUSDR6_1(.din(n11978), .dout(n11981));
    jdff dff_B_7oCASZGe3_1(.din(n11981), .dout(n11984));
    jdff dff_B_4VyW49zX9_1(.din(n11984), .dout(n11987));
    jdff dff_B_pk97WiTA1_1(.din(n11987), .dout(n11990));
    jdff dff_B_xZKYKqV27_1(.din(n11990), .dout(n11993));
    jdff dff_B_Mz1q1YI47_1(.din(n11993), .dout(n11996));
    jdff dff_B_o1XJSCTh3_1(.din(n11996), .dout(n11999));
    jdff dff_B_IGC0S6jD6_1(.din(n11999), .dout(n12002));
    jdff dff_B_aTPdqReg6_1(.din(n12002), .dout(n12005));
    jdff dff_B_vxIYgitq5_1(.din(n12005), .dout(n12008));
    jdff dff_B_ZXtwGK773_1(.din(n12008), .dout(n12011));
    jdff dff_B_2iFnCUuU8_1(.din(n12011), .dout(n12014));
    jdff dff_B_RsyCdviq3_1(.din(n12014), .dout(n12017));
    jdff dff_B_nfriTmIm4_1(.din(n12017), .dout(n12020));
    jdff dff_B_oO0jZObY5_1(.din(n12020), .dout(n12023));
    jdff dff_B_BrvrR8gC2_1(.din(n12023), .dout(n12026));
    jdff dff_B_LJxHPsYZ4_1(.din(n12026), .dout(n12029));
    jdff dff_B_luDCltd93_1(.din(n12029), .dout(n12032));
    jdff dff_B_jDfHQxtX6_1(.din(n4117), .dout(n12035));
    jdff dff_B_padfVtME6_1(.din(n12035), .dout(n12038));
    jdff dff_B_YNsgfuEa4_1(.din(n12038), .dout(n12041));
    jdff dff_B_ySbCi0UA4_1(.din(n12041), .dout(n12044));
    jdff dff_B_sT2LG1VA4_1(.din(n12044), .dout(n12047));
    jdff dff_B_VkuhmvWQ4_1(.din(n12047), .dout(n12050));
    jdff dff_B_weELPwBH8_1(.din(n12050), .dout(n12053));
    jdff dff_B_MoK8K3V77_1(.din(n12053), .dout(n12056));
    jdff dff_B_aFiCM8Xa7_1(.din(n12056), .dout(n12059));
    jdff dff_B_RmXhfKrA5_1(.din(n12059), .dout(n12062));
    jdff dff_B_A9342yTM3_1(.din(n12062), .dout(n12065));
    jdff dff_B_DuUQPFvb7_1(.din(n12065), .dout(n12068));
    jdff dff_B_uo74DPz82_1(.din(n12068), .dout(n12071));
    jdff dff_B_PncgLYtv6_1(.din(n12071), .dout(n12074));
    jdff dff_B_1oMPnq7s8_1(.din(n12074), .dout(n12077));
    jdff dff_B_Y4voQsKt4_1(.din(n12077), .dout(n12080));
    jdff dff_B_6ZOy3w3J2_1(.din(n12080), .dout(n12083));
    jdff dff_B_OcKKJx5L0_1(.din(n12083), .dout(n12086));
    jdff dff_B_MLZPxglE7_1(.din(n12086), .dout(n12089));
    jdff dff_B_1H8NVeIm3_1(.din(n12089), .dout(n12092));
    jdff dff_B_ikio3lpP7_1(.din(n12092), .dout(n12095));
    jdff dff_A_IuxooMrp3_0(.din(n12152), .dout(n12097));
    jdff dff_B_g5yGYdSh2_2(.din(n4120), .dout(n12101));
    jdff dff_B_roBgkliS7_2(.din(n12101), .dout(n12104));
    jdff dff_B_5yXtPHCI4_2(.din(n12104), .dout(n12107));
    jdff dff_B_czORjX8i6_2(.din(n12107), .dout(n12110));
    jdff dff_B_vkNiYCuI6_2(.din(n12110), .dout(n12113));
    jdff dff_B_AamhJqBS7_2(.din(n12113), .dout(n12116));
    jdff dff_B_omN9lnRC1_2(.din(n12116), .dout(n12119));
    jdff dff_B_BvWSSrzu4_2(.din(n12119), .dout(n12122));
    jdff dff_B_V4gj3nKw4_2(.din(n12122), .dout(n12125));
    jdff dff_B_SMP7N7Ck0_2(.din(n12125), .dout(n12128));
    jdff dff_B_Up4m6slZ1_2(.din(n12128), .dout(n12131));
    jdff dff_B_UrTGNWhK7_2(.din(n12131), .dout(n12134));
    jdff dff_B_mBdl030i6_2(.din(n12134), .dout(n12137));
    jdff dff_B_8pQKnd758_2(.din(n12137), .dout(n12140));
    jdff dff_B_6ObSEDAw4_2(.din(n12140), .dout(n12143));
    jdff dff_B_KGY4CxUr5_2(.din(n12143), .dout(n12146));
    jdff dff_B_qXfQcp5F7_2(.din(n12146), .dout(n12149));
    jdff dff_B_Y5woxDGt8_2(.din(n12149), .dout(n12152));
    jdff dff_B_AGhvN9KA2_0(.din(n4809), .dout(n12155));
    jdff dff_B_0gJncxEk9_0(.din(n12155), .dout(n12158));
    jdff dff_B_AdBgfhpW3_0(.din(n12158), .dout(n12161));
    jdff dff_B_0TCVwuZs8_0(.din(n12161), .dout(n12164));
    jdff dff_B_rfKLOvf55_0(.din(n12164), .dout(n12167));
    jdff dff_B_05v4G4EF4_0(.din(n12167), .dout(n12170));
    jdff dff_B_FOqQI0gV0_0(.din(n12170), .dout(n12173));
    jdff dff_B_8ImvVHjO3_0(.din(n12173), .dout(n12176));
    jdff dff_B_X2YReIlf9_0(.din(n12176), .dout(n12179));
    jdff dff_B_LZXWKBZ50_0(.din(n12179), .dout(n12182));
    jdff dff_B_9xnFQAWl5_0(.din(n12182), .dout(n12185));
    jdff dff_B_98YENKx82_0(.din(n12185), .dout(n12188));
    jdff dff_B_E4vM521R1_0(.din(n12188), .dout(n12191));
    jdff dff_B_L07YgFGf5_0(.din(n12191), .dout(n12194));
    jdff dff_B_svOPQ0IX8_0(.din(n12194), .dout(n12197));
    jdff dff_B_XoqK1Qrf7_0(.din(n12197), .dout(n12200));
    jdff dff_B_mNVELAZ65_0(.din(n12200), .dout(n12203));
    jdff dff_B_wNjScP6a2_0(.din(n12203), .dout(n12206));
    jdff dff_B_F1pYMPkp7_0(.din(n12206), .dout(n12209));
    jdff dff_B_f6SH1Swa5_0(.din(n12209), .dout(n12212));
    jdff dff_B_QktJqICt2_0(.din(n12212), .dout(n12215));
    jdff dff_B_sF6oPbsM6_0(.din(n4801), .dout(n12218));
    jdff dff_B_5kIPSHbN4_0(.din(n12218), .dout(n12221));
    jdff dff_B_4T9BR8210_0(.din(n12221), .dout(n12224));
    jdff dff_B_Kzz4PDiU8_0(.din(n4797), .dout(n12227));
    jdff dff_B_nODN7bvz1_0(.din(n12227), .dout(n12230));
    jdff dff_A_gwZYhnKO5_1(.din(n12235), .dout(n12232));
    jdff dff_A_RvPdg9DA4_1(.din(n12238), .dout(n12235));
    jdff dff_A_r5vwT7TT8_1(.din(n12241), .dout(n12238));
    jdff dff_A_0EY8Gc0Y3_1(.din(n12244), .dout(n12241));
    jdff dff_A_L9KEOYBB9_1(.din(n12247), .dout(n12244));
    jdff dff_A_m5ViydYv5_1(.din(n12250), .dout(n12247));
    jdff dff_A_yoPZSWl13_1(.din(n12253), .dout(n12250));
    jdff dff_A_qWKx2dOq8_1(.din(n674), .dout(n12253));
    jdff dff_B_eFgGSVwm2_1(.din(n4778), .dout(n12257));
    jdff dff_B_0FngQeLD3_1(.din(n12257), .dout(n12260));
    jdff dff_A_eZXnlpvS8_1(.din(n12265), .dout(n12262));
    jdff dff_A_6h3bIYF37_1(.din(n12268), .dout(n12265));
    jdff dff_A_7VYmYoYr9_1(.din(n12271), .dout(n12268));
    jdff dff_A_2poalKMA2_1(.din(n12274), .dout(n12271));
    jdff dff_A_KIx2VHi19_1(.din(n12277), .dout(n12274));
    jdff dff_A_5cO6ktaw9_1(.din(n12280), .dout(n12277));
    jdff dff_A_JejYPRDo3_1(.din(n12283), .dout(n12280));
    jdff dff_A_wCJ2uaZ43_1(.din(n12286), .dout(n12283));
    jdff dff_A_6xxYKv2a0_1(.din(n12289), .dout(n12286));
    jdff dff_A_tylyX5up8_1(.din(n12292), .dout(n12289));
    jdff dff_A_EZadv2aC4_1(.din(n12295), .dout(n12292));
    jdff dff_A_K311HNM89_1(.din(n12298), .dout(n12295));
    jdff dff_A_3pwP2hv86_1(.din(n12301), .dout(n12298));
    jdff dff_A_4NJksY3z7_1(.din(n12304), .dout(n12301));
    jdff dff_A_1Mj12XJM8_1(.din(n12307), .dout(n12304));
    jdff dff_A_fEZDBPaJ9_1(.din(n12310), .dout(n12307));
    jdff dff_A_9ZwlWKzu7_1(.din(n12313), .dout(n12310));
    jdff dff_A_BZTD7tpw2_1(.din(n12316), .dout(n12313));
    jdff dff_A_qjjDobR02_1(.din(n12319), .dout(n12316));
    jdff dff_A_OjhF358c0_1(.din(n12322), .dout(n12319));
    jdff dff_A_Tz7kdlG23_1(.din(n12325), .dout(n12322));
    jdff dff_A_9McRTXCu6_1(.din(n12328), .dout(n12325));
    jdff dff_A_XBoqCcEx7_1(.din(n12331), .dout(n12328));
    jdff dff_A_fdzOriLl1_1(.din(n12334), .dout(n12331));
    jdff dff_A_vYHgwxc30_1(.din(n12337), .dout(n12334));
    jdff dff_A_PZw6Hh9P7_1(.din(n12340), .dout(n12337));
    jdff dff_A_jarPTf8q0_1(.din(n12343), .dout(n12340));
    jdff dff_A_Mo5ZWezW7_1(.din(n12350), .dout(n12343));
    jdff dff_B_AnofVKPO2_2(.din(n4353), .dout(n12347));
    jdff dff_B_lJ5QNjnV4_2(.din(n12347), .dout(n12350));
    jdff dff_A_g92e85O21_2(.din(n12355), .dout(n12352));
    jdff dff_A_aglXCVb96_2(.din(n12358), .dout(n12355));
    jdff dff_A_YWRAjuvE8_2(.din(n12361), .dout(n12358));
    jdff dff_A_i34odZJ98_2(.din(n12364), .dout(n12361));
    jdff dff_A_3uf1oS8C3_2(.din(n12367), .dout(n12364));
    jdff dff_A_fYTI9cJ48_2(.din(n12370), .dout(n12367));
    jdff dff_A_AevRGeN78_2(.din(n12373), .dout(n12370));
    jdff dff_A_3J8NWZDi6_2(.din(n12376), .dout(n12373));
    jdff dff_A_TnqrOvdt0_2(.din(n12379), .dout(n12376));
    jdff dff_A_51aRyeB72_2(.din(n12382), .dout(n12379));
    jdff dff_A_woUc07xg0_2(.din(n12385), .dout(n12382));
    jdff dff_A_IjzyheDb7_2(.din(n12388), .dout(n12385));
    jdff dff_A_CxhTikps9_2(.din(n12391), .dout(n12388));
    jdff dff_A_MQNbCX390_2(.din(n12394), .dout(n12391));
    jdff dff_A_UE8spiDH8_2(.din(n12397), .dout(n12394));
    jdff dff_A_qrthNcPY3_2(.din(n12400), .dout(n12397));
    jdff dff_A_nXS0nba76_2(.din(n12403), .dout(n12400));
    jdff dff_A_W52wLRxE4_2(.din(n12406), .dout(n12403));
    jdff dff_A_jRNRbCtR5_2(.din(n12409), .dout(n12406));
    jdff dff_A_v90dEzJ47_2(.din(n12412), .dout(n12409));
    jdff dff_A_DvqT2GfO2_2(.din(n12415), .dout(n12412));
    jdff dff_A_gAZ44v0g8_2(.din(n12418), .dout(n12415));
    jdff dff_A_C5SgrmPL0_2(.din(n662), .dout(n12418));
    jdff dff_B_Xzk5kxbQ0_1(.din(n555), .dout(n12422));
    jdff dff_B_EDueLPXN5_1(.din(n12422), .dout(n12425));
    jdff dff_B_pYGNNO9i9_1(.din(n12425), .dout(n12428));
    jdff dff_B_9j5IoNto8_1(.din(n12428), .dout(n12431));
    jdff dff_B_RWZ0nrv75_1(.din(n562), .dout(n12434));
    jdff dff_B_erbnnowH2_1(.din(n12434), .dout(n12437));
    jdff dff_B_R04qSkmn0_1(.din(n12437), .dout(n12440));
    jdff dff_B_ZQDWXIqq6_1(.din(n12440), .dout(n12443));
    jdff dff_B_Cw6wK2kq0_1(.din(n12443), .dout(n12446));
    jdff dff_A_BrJEZedj3_2(.din(n12451), .dout(n12448));
    jdff dff_A_HHPEyq3M9_2(.din(n12454), .dout(n12451));
    jdff dff_A_CJL8xyZz6_2(.din(n12457), .dout(n12454));
    jdff dff_A_dVODatoS0_2(.din(n12460), .dout(n12457));
    jdff dff_A_oU1ZM55K8_2(.din(n12463), .dout(n12460));
    jdff dff_A_sGjIIncj7_2(.din(n12466), .dout(n12463));
    jdff dff_A_6llkRCZ02_2(.din(n12469), .dout(n12466));
    jdff dff_A_SIOtIOml7_2(.din(n12472), .dout(n12469));
    jdff dff_A_glWGlEd73_2(.din(n12475), .dout(n12472));
    jdff dff_A_Cgz9fZJ48_2(.din(n12478), .dout(n12475));
    jdff dff_A_OILiBMmN9_2(.din(n12481), .dout(n12478));
    jdff dff_A_XSWRAldS2_2(.din(n12484), .dout(n12481));
    jdff dff_A_9HBIlFH77_2(.din(n12487), .dout(n12484));
    jdff dff_A_skJRAPsS0_2(.din(n12490), .dout(n12487));
    jdff dff_A_SPi4HDhp5_2(.din(n12493), .dout(n12490));
    jdff dff_A_LoqPWNol5_2(.din(n12496), .dout(n12493));
    jdff dff_A_UUzoMG4o9_2(.din(n12499), .dout(n12496));
    jdff dff_A_lhgEor1P6_2(.din(n12502), .dout(n12499));
    jdff dff_A_zMNFwiqL0_2(.din(n12505), .dout(n12502));
    jdff dff_A_jYck3y3b9_2(.din(n12508), .dout(n12505));
    jdff dff_A_2NPYQQ0K2_2(.din(n12511), .dout(n12508));
    jdff dff_A_BzExDJok8_2(.din(n12514), .dout(n12511));
    jdff dff_A_lXNnTDcK2_2(.din(n12517), .dout(n12514));
    jdff dff_A_r0jkB8Pt3_2(.din(n12520), .dout(n12517));
    jdff dff_A_Amuwpa848_2(.din(n654), .dout(n12520));
    jdff dff_B_ip9tF0zH7_1(.din(n625), .dout(n12524));
    jdff dff_A_0KsNRUZ00_0(.din(n639), .dout(n12526));
    jdff dff_A_Vzst1tsa8_1(.din(n12532), .dout(n12529));
    jdff dff_A_HW0CNNaM1_1(.din(n12535), .dout(n12532));
    jdff dff_A_LiijGa0q0_1(.din(n12538), .dout(n12535));
    jdff dff_A_Rk8SrjUc5_1(.din(n12541), .dout(n12538));
    jdff dff_A_DSp4yWnr1_1(.din(n12544), .dout(n12541));
    jdff dff_A_LmdZapYT8_1(.din(n12547), .dout(n12544));
    jdff dff_A_Q4snMDE10_1(.din(n12550), .dout(n12547));
    jdff dff_A_nczq2ASh7_1(.din(n12553), .dout(n12550));
    jdff dff_A_rqdMaNH98_1(.din(n12556), .dout(n12553));
    jdff dff_A_K1SvHrs10_1(.din(n12559), .dout(n12556));
    jdff dff_A_Z4gY4QN91_1(.din(n12562), .dout(n12559));
    jdff dff_A_v3e3znSJ6_1(.din(n12565), .dout(n12562));
    jdff dff_A_986pFOJR1_1(.din(n12568), .dout(n12565));
    jdff dff_A_5DzojULb4_1(.din(n12571), .dout(n12568));
    jdff dff_A_Wrp4ADXB5_1(.din(n12574), .dout(n12571));
    jdff dff_A_EKEE6Tlo2_1(.din(n12577), .dout(n12574));
    jdff dff_A_b7NjEgFW8_1(.din(n12580), .dout(n12577));
    jdff dff_A_A9wfmooN6_1(.din(n12583), .dout(n12580));
    jdff dff_A_mTKAX2b75_1(.din(n12586), .dout(n12583));
    jdff dff_A_Z0DGIgll9_1(.din(n12589), .dout(n12586));
    jdff dff_A_Xxub7PmQ3_1(.din(n12592), .dout(n12589));
    jdff dff_A_Pq2XUUwU2_1(.din(n12595), .dout(n12592));
    jdff dff_A_jcUCBrq45_1(.din(n12598), .dout(n12595));
    jdff dff_A_dkolpX118_1(.din(n12601), .dout(n12598));
    jdff dff_A_njsPvHKF3_1(.din(n12604), .dout(n12601));
    jdff dff_A_hbAV5I5r2_1(.din(n12607), .dout(n12604));
    jdff dff_A_RhSNtQ7o7_1(.din(n12610), .dout(n12607));
    jdff dff_A_vHpQMJM47_1(.din(n12613), .dout(n12610));
    jdff dff_A_Apmk8SeQ1_1(.din(n12616), .dout(n12613));
    jdff dff_A_BhdubKHE1_1(.din(n12619), .dout(n12616));
    jdff dff_A_5xjHTlCY6_1(.din(n12622), .dout(n12619));
    jdff dff_A_nsaHze9V0_1(.din(n639), .dout(n12622));
    jdff dff_B_bZf3Y5AV4_0(.din(G216), .dout(n12626));
    jdff dff_A_rOTyxRsQ1_0(.din(n12631), .dout(n12628));
    jdff dff_A_BBzGkKiJ5_0(.din(n595), .dout(n12631));
    jdff dff_A_ueWiOO963_1(.din(n12637), .dout(n12634));
    jdff dff_A_oj1IjktD9_1(.din(n595), .dout(n12637));
    jdff dff_A_MChL85tW9_0(.din(n12643), .dout(n12640));
    jdff dff_A_XMXSjf4L9_0(.din(n12646), .dout(n12643));
    jdff dff_A_UyLnJLpV5_0(.din(n12649), .dout(n12646));
    jdff dff_A_XvxZdTNf7_0(.din(n12652), .dout(n12649));
    jdff dff_A_wx8BE9BM7_0(.din(n592), .dout(n12652));
    jdff dff_B_SYp4AUKk5_2(.din(G209), .dout(n12656));
    jdff dff_A_5XFw2BK36_0(.din(n12661), .dout(n12658));
    jdff dff_A_qqy3ED7z2_0(.din(n580), .dout(n12661));
    jdff dff_A_GpfuqmSP6_1(.din(n12667), .dout(n12664));
    jdff dff_A_JXnlarNW9_1(.din(n580), .dout(n12667));
    jdff dff_A_j3rjMdM79_0(.din(n577), .dout(n12670));
    jdff dff_A_SRJSWJeu4_2(.din(n577), .dout(n12673));
    jdff dff_A_vKP5qq0L8_0(.din(n12679), .dout(n12676));
    jdff dff_A_t6sCCjTH2_0(.din(n537), .dout(n12679));
    jdff dff_A_p5p2AGaa0_2(.din(n12685), .dout(n12682));
    jdff dff_A_zbGCICaN3_2(.din(n12688), .dout(n12685));
    jdff dff_A_eO1qbKxK0_2(.din(n12691), .dout(n12688));
    jdff dff_A_bSvOCi7B0_2(.din(n12694), .dout(n12691));
    jdff dff_A_TP1DRJpF5_2(.din(n12697), .dout(n12694));
    jdff dff_A_zxZQCvQJ6_2(.din(n12700), .dout(n12697));
    jdff dff_A_idthlT9g4_2(.din(n537), .dout(n12700));
    jdff dff_A_kjpjMtHF4_0(.din(n12706), .dout(n12703));
    jdff dff_A_tkqNoS2v5_0(.din(n525), .dout(n12706));
    jdff dff_B_a909KlhV4_0(.din(G213), .dout(n12710));
    jdff dff_A_X1TuwsZf3_1(.din(n12715), .dout(n12712));
    jdff dff_A_nuxPCBOz4_1(.din(n514), .dout(n12715));
    jdff dff_A_FM3mH6a44_2(.din(n12721), .dout(n12718));
    jdff dff_A_fWSAdVKo6_2(.din(n514), .dout(n12721));
    jdff dff_B_dxI4Drpe8_1(.din(n1031), .dout(n12725));
    jdff dff_B_pmThCi3D0_1(.din(n12725), .dout(n12728));
    jdff dff_B_iAKDS9Hl0_1(.din(n12728), .dout(n12731));
    jdff dff_B_fLkGQpSK7_1(.din(n12731), .dout(n12734));
    jdff dff_B_ouyj905a4_1(.din(n12734), .dout(n12737));
    jdff dff_B_wsYh0W1j6_1(.din(n12737), .dout(n12740));
    jdff dff_B_s7kfYvyR7_1(.din(n12740), .dout(n12743));
    jdff dff_B_djipIL9X3_1(.din(n12743), .dout(n12746));
    jdff dff_B_HaqvBl8E4_1(.din(n12746), .dout(n12749));
    jdff dff_B_3wgKmfbH2_1(.din(n12749), .dout(n12752));
    jdff dff_B_g1HA1iMZ8_1(.din(n12752), .dout(n12755));
    jdff dff_B_hV6BjzUi4_1(.din(n12755), .dout(n12758));
    jdff dff_B_gLD3NANP0_1(.din(n12758), .dout(n12761));
    jdff dff_B_6uYLmdzp6_1(.din(n12761), .dout(n12764));
    jdff dff_B_1XOwPlP90_1(.din(n12764), .dout(n12767));
    jdff dff_B_jhN7ONri7_1(.din(n12767), .dout(n12770));
    jdff dff_B_jQqlgt9b9_1(.din(n12770), .dout(n12773));
    jdff dff_B_eOrW3sMd4_1(.din(n12773), .dout(n12776));
    jdff dff_B_ivJcWUpd4_1(.din(n12776), .dout(n12779));
    jdff dff_B_A9ljM3pL5_0(.din(n1741), .dout(n12782));
    jdff dff_B_vWTXuyzV1_0(.din(n12782), .dout(n12785));
    jdff dff_B_gFmnUpz72_0(.din(n12785), .dout(n12788));
    jdff dff_B_5hs3d9dS8_0(.din(n12788), .dout(n12791));
    jdff dff_B_glKRk3gR5_0(.din(n12791), .dout(n12794));
    jdff dff_B_9rtOB0Lq3_0(.din(n12794), .dout(n12797));
    jdff dff_B_3yjIZrto9_0(.din(n12797), .dout(n12800));
    jdff dff_B_O2veVFGl5_0(.din(n12800), .dout(n12803));
    jdff dff_B_7TVa7QrY6_0(.din(n12803), .dout(n12806));
    jdff dff_B_sagEw58q7_0(.din(n12806), .dout(n12809));
    jdff dff_B_c6HAdUaN2_0(.din(n12809), .dout(n12812));
    jdff dff_B_lAEfoLb51_0(.din(n12812), .dout(n12815));
    jdff dff_B_n6A6nBpW3_0(.din(n12815), .dout(n12818));
    jdff dff_B_pce0MwIA2_0(.din(n12818), .dout(n12821));
    jdff dff_A_I7xDzB0S6_0(.din(n12826), .dout(n12823));
    jdff dff_A_cNv0txgm3_0(.din(n12829), .dout(n12826));
    jdff dff_A_aoVUsHNH4_0(.din(n12832), .dout(n12829));
    jdff dff_A_uMMjXF7A7_0(.din(n12835), .dout(n12832));
    jdff dff_A_jRglSfii3_0(.din(n12838), .dout(n12835));
    jdff dff_A_5hsSyzRu8_0(.din(n12841), .dout(n12838));
    jdff dff_A_aXu3DKeP5_0(.din(n12844), .dout(n12841));
    jdff dff_A_nmfzxFhA3_0(.din(n12847), .dout(n12844));
    jdff dff_A_USPKJ8132_0(.din(n12850), .dout(n12847));
    jdff dff_A_X2pZoTDj5_0(.din(n12853), .dout(n12850));
    jdff dff_A_f4xdTZ1k0_0(.din(n12856), .dout(n12853));
    jdff dff_A_Rszs5hxt9_0(.din(n12859), .dout(n12856));
    jdff dff_A_0C7stwN52_0(.din(n12862), .dout(n12859));
    jdff dff_A_JicpSNRF3_0(.din(n12865), .dout(n12862));
    jdff dff_A_b1VtYyyq2_0(.din(n1738), .dout(n12865));
    jdff dff_B_4l6EjjZ92_1(.din(n1708), .dout(n12869));
    jdff dff_B_4mONRwjK5_1(.din(n12869), .dout(n12872));
    jdff dff_B_2OvdcqoQ8_1(.din(n12872), .dout(n12875));
    jdff dff_B_tWHvgilG5_1(.din(n1072), .dout(n12878));
    jdff dff_B_j3c8LBmL0_1(.din(n12878), .dout(n12881));
    jdff dff_B_NRkqAHc08_1(.din(n12881), .dout(n12884));
    jdff dff_B_UU5OWMm29_1(.din(n12884), .dout(n12887));
    jdff dff_B_FF9BiwNp5_1(.din(n12887), .dout(n12890));
    jdff dff_B_ydLvFe607_1(.din(n12890), .dout(n12893));
    jdff dff_B_OaK0ATQs6_1(.din(n12893), .dout(n12896));
    jdff dff_B_BkLkavyk7_1(.din(n12896), .dout(n12899));
    jdff dff_B_xt3rlacS3_1(.din(n12899), .dout(n12902));
    jdff dff_B_Nb90LzJ29_1(.din(n12902), .dout(n12905));
    jdff dff_B_xEI4AJRJ0_1(.din(n12905), .dout(n12908));
    jdff dff_B_BuNIFx2m3_1(.din(n12908), .dout(n12911));
    jdff dff_B_uwJGeuQo2_1(.din(n12911), .dout(n12914));
    jdff dff_B_fLrw1hNJ4_1(.din(n12914), .dout(n12917));
    jdff dff_B_KpiQnyyo5_1(.din(n12917), .dout(n12920));
    jdff dff_B_4YOywbhc6_1(.din(n12920), .dout(n12923));
    jdff dff_B_pE2wBYNa4_1(.din(n12923), .dout(n12926));
    jdff dff_B_ZCvoo7Hx9_1(.din(n1101), .dout(n12929));
    jdff dff_B_pW0r1VbN2_1(.din(n12929), .dout(n12932));
    jdff dff_B_ZnnPsRxJ0_1(.din(n12932), .dout(n12935));
    jdff dff_B_MQNi7O0W7_1(.din(n12935), .dout(n12938));
    jdff dff_B_aoeJBiiz8_1(.din(n12938), .dout(n12941));
    jdff dff_B_P0hiPupE3_1(.din(n12941), .dout(n12944));
    jdff dff_B_HR0JZQQm7_1(.din(n12944), .dout(n12947));
    jdff dff_B_BPWMRp4e6_1(.din(n12947), .dout(n12950));
    jdff dff_B_hD6mkblq0_1(.din(n12950), .dout(n12953));
    jdff dff_B_bOk8bYvH9_1(.din(n12953), .dout(n12956));
    jdff dff_B_sBFOXOMN7_1(.din(n12956), .dout(n12959));
    jdff dff_B_vvQeQ9IZ6_1(.din(n12959), .dout(n12962));
    jdff dff_B_KrkYt20q1_1(.din(n12962), .dout(n12965));
    jdff dff_B_qToOmZvf7_1(.din(n12965), .dout(n12968));
    jdff dff_A_4AY1VK1h7_1(.din(n12973), .dout(n12970));
    jdff dff_A_OiCKnY8w5_1(.din(n12976), .dout(n12973));
    jdff dff_A_e0Ejqhux7_1(.din(n12979), .dout(n12976));
    jdff dff_A_5h6Q7F6G2_1(.din(n12982), .dout(n12979));
    jdff dff_A_kBBqhWdO2_1(.din(n12985), .dout(n12982));
    jdff dff_A_A1dL6dWk5_1(.din(n12988), .dout(n12985));
    jdff dff_A_n0BAAhXE8_1(.din(n12991), .dout(n12988));
    jdff dff_A_8vjMpDMc9_1(.din(n12994), .dout(n12991));
    jdff dff_A_F3FI9HFu1_1(.din(n12997), .dout(n12994));
    jdff dff_A_bUTvmJwf9_1(.din(n13000), .dout(n12997));
    jdff dff_A_W6Q6hwAB4_1(.din(n13003), .dout(n13000));
    jdff dff_A_CcYGYwLY7_1(.din(n13006), .dout(n13003));
    jdff dff_A_UGw49bNO0_1(.din(n13009), .dout(n13006));
    jdff dff_A_elMZDeJw5_1(.din(n13012), .dout(n13009));
    jdff dff_A_IATSXNEX0_1(.din(n13015), .dout(n13012));
    jdff dff_A_7TcVFsax4_1(.din(n13018), .dout(n13015));
    jdff dff_A_YY9Wa9DR3_1(.din(n13021), .dout(n13018));
    jdff dff_A_wAQ3i3Jc9_1(.din(n13024), .dout(n13021));
    jdff dff_A_6rMMNjas3_1(.din(n1050), .dout(n13024));
    jdff dff_A_mysvAp8W3_0(.din(n13030), .dout(n13027));
    jdff dff_A_W2jLkjl70_0(.din(n13033), .dout(n13030));
    jdff dff_A_wBl7ND0M6_0(.din(n13036), .dout(n13033));
    jdff dff_A_1kHYwltR7_0(.din(n13039), .dout(n13036));
    jdff dff_A_wVENETGK6_0(.din(n13042), .dout(n13039));
    jdff dff_A_9T32hcbM6_0(.din(n13045), .dout(n13042));
    jdff dff_A_cIucq7oY5_0(.din(n13048), .dout(n13045));
    jdff dff_A_DIfLTP544_0(.din(n13051), .dout(n13048));
    jdff dff_A_FEqIZsnq9_0(.din(n13054), .dout(n13051));
    jdff dff_A_EurOJcZ53_0(.din(n13057), .dout(n13054));
    jdff dff_A_8oSIy0W82_0(.din(n13060), .dout(n13057));
    jdff dff_A_4nbLLgR66_0(.din(n13063), .dout(n13060));
    jdff dff_A_N0awK1a70_0(.din(n13066), .dout(n13063));
    jdff dff_A_hY21ZafV7_0(.din(n13069), .dout(n13066));
    jdff dff_A_4jEY70Uv7_0(.din(n13072), .dout(n13069));
    jdff dff_A_hVdWN37r8_0(.din(n13075), .dout(n13072));
    jdff dff_A_bZG6rCt02_0(.din(n13078), .dout(n13075));
    jdff dff_A_j8Yyd3C18_0(.din(n13081), .dout(n13078));
    jdff dff_A_TytrfGEn0_0(.din(n13084), .dout(n13081));
    jdff dff_A_nQGtR75U2_0(.din(n1028), .dout(n13084));
    jdff dff_A_wXmX0e7m5_1(.din(n13090), .dout(n13087));
    jdff dff_A_dhNvzuby7_1(.din(n13093), .dout(n13090));
    jdff dff_A_DJqP3u7M2_1(.din(n13096), .dout(n13093));
    jdff dff_A_7Fqir6Uc3_1(.din(n13099), .dout(n13096));
    jdff dff_A_lRaNFEFP2_1(.din(n13102), .dout(n13099));
    jdff dff_A_4lf6tUkl5_1(.din(n13105), .dout(n13102));
    jdff dff_A_xVpNistd5_1(.din(n13108), .dout(n13105));
    jdff dff_A_4Q0HkovC8_1(.din(n13111), .dout(n13108));
    jdff dff_A_05cVpLKY5_1(.din(n13114), .dout(n13111));
    jdff dff_A_I3EHgkKR5_1(.din(n13117), .dout(n13114));
    jdff dff_A_TDuqIGv35_1(.din(n13120), .dout(n13117));
    jdff dff_A_H5Du67Uf9_1(.din(n13123), .dout(n13120));
    jdff dff_A_4FXWiXsM1_1(.din(n13126), .dout(n13123));
    jdff dff_A_DavtVEpX0_1(.din(n13129), .dout(n13126));
    jdff dff_A_Cfo0Ft2p4_1(.din(n13132), .dout(n13129));
    jdff dff_A_92OGamdW0_1(.din(n13135), .dout(n13132));
    jdff dff_A_lUlKWWju8_1(.din(n13138), .dout(n13135));
    jdff dff_A_IsUwWonB5_1(.din(n13141), .dout(n13138));
    jdff dff_A_ZAjNNJfD7_1(.din(n13144), .dout(n13141));
    jdff dff_A_1VSTvnbX6_1(.din(n13147), .dout(n13144));
    jdff dff_A_gHh1LAwz8_1(.din(n13150), .dout(n13147));
    jdff dff_A_RxW72wH48_1(.din(n1021), .dout(n13150));
    jdff dff_A_pV3i2Oqw1_1(.din(n13156), .dout(n13153));
    jdff dff_A_rZ0hgTC95_1(.din(n13159), .dout(n13156));
    jdff dff_A_hQTC4fE15_1(.din(n13162), .dout(n13159));
    jdff dff_A_mslwNtHw0_1(.din(n13165), .dout(n13162));
    jdff dff_A_ijRyzMBZ9_1(.din(n13168), .dout(n13165));
    jdff dff_A_wlVkLV6h4_1(.din(n13171), .dout(n13168));
    jdff dff_A_yWUIeNXJ3_1(.din(n13174), .dout(n13171));
    jdff dff_A_pQb2xkDp4_1(.din(n13177), .dout(n13174));
    jdff dff_A_8yZtTeNR1_1(.din(n13180), .dout(n13177));
    jdff dff_A_HSRsi5bl1_1(.din(n13183), .dout(n13180));
    jdff dff_A_cFUZ2Tor7_1(.din(n13186), .dout(n13183));
    jdff dff_A_3YjeGyEk6_1(.din(n13189), .dout(n13186));
    jdff dff_A_kodrTzqj5_1(.din(n13192), .dout(n13189));
    jdff dff_A_lMCx3fHi1_1(.din(n13195), .dout(n13192));
    jdff dff_A_ySDlUllu3_1(.din(n13198), .dout(n13195));
    jdff dff_A_fNRZdPWU1_1(.din(n13201), .dout(n13198));
    jdff dff_A_wmgdaXR69_1(.din(n13204), .dout(n13201));
    jdff dff_A_AJ2RaLHq2_1(.din(n1002), .dout(n13204));
    jdff dff_A_ZHrf0Wum6_1(.din(n13210), .dout(n13207));
    jdff dff_A_tIa5nNvV2_1(.din(n13213), .dout(n13210));
    jdff dff_A_g1XOuA2k6_1(.din(n13216), .dout(n13213));
    jdff dff_A_5RRLB7Y64_1(.din(n13219), .dout(n13216));
    jdff dff_A_CpQPaSC28_1(.din(n13222), .dout(n13219));
    jdff dff_A_BTgskNrm5_1(.din(n13225), .dout(n13222));
    jdff dff_A_4IMIwSgI0_1(.din(n13228), .dout(n13225));
    jdff dff_A_8XtrJMHW8_1(.din(n13231), .dout(n13228));
    jdff dff_A_FXU8MAlH3_1(.din(n13234), .dout(n13231));
    jdff dff_A_pfxgqJCX4_1(.din(n13237), .dout(n13234));
    jdff dff_A_nNkPY3zj6_1(.din(n13240), .dout(n13237));
    jdff dff_A_2CeUZ8G02_1(.din(n13243), .dout(n13240));
    jdff dff_A_mRi2UOy46_1(.din(n13246), .dout(n13243));
    jdff dff_A_bxcvZCMb8_1(.din(n13249), .dout(n13246));
    jdff dff_A_ELfkE1sR4_1(.din(n13252), .dout(n13249));
    jdff dff_A_SzNhROO54_1(.din(n13255), .dout(n13252));
    jdff dff_A_YKcXgaSB9_1(.din(n998), .dout(n13255));
    jdff dff_A_2h3sDGq20_0(.din(n13261), .dout(n13258));
    jdff dff_A_xQp4L2oT1_0(.din(n13264), .dout(n13261));
    jdff dff_A_lP7LBitw2_0(.din(n13267), .dout(n13264));
    jdff dff_A_NeiOiegw4_0(.din(n13270), .dout(n13267));
    jdff dff_A_YCAS7qFR3_0(.din(n13273), .dout(n13270));
    jdff dff_A_aVVmcqqy9_0(.din(n13276), .dout(n13273));
    jdff dff_A_xqJnR9AY2_0(.din(n13279), .dout(n13276));
    jdff dff_A_5pBWwoNE3_0(.din(n13282), .dout(n13279));
    jdff dff_A_3Y0zYfS50_0(.din(n13285), .dout(n13282));
    jdff dff_A_QA8uoGzG6_0(.din(n13288), .dout(n13285));
    jdff dff_A_Ei0Pduxf5_0(.din(n13291), .dout(n13288));
    jdff dff_A_AzQzgRyV6_0(.din(n13294), .dout(n13291));
    jdff dff_A_tVVeXCWX9_0(.din(n13297), .dout(n13294));
    jdff dff_A_M04ERNrn8_0(.din(n13300), .dout(n13297));
    jdff dff_A_DURmX0lG4_0(.din(n13303), .dout(n13300));
    jdff dff_A_HshRxNag0_0(.din(n13306), .dout(n13303));
    jdff dff_A_qnv7e2B19_0(.din(n13309), .dout(n13306));
    jdff dff_A_M68AdHPb8_0(.din(n13312), .dout(n13309));
    jdff dff_A_IHcVICTS5_0(.din(n990), .dout(n13312));
    jdff dff_B_tus5eRkm1_1(.din(n935), .dout(n13316));
    jdff dff_B_eAXF9DqD6_1(.din(n13316), .dout(n13319));
    jdff dff_B_gyQ2zbRa9_1(.din(n13319), .dout(n13322));
    jdff dff_A_tuc5fw9a7_0(.din(n13327), .dout(n13324));
    jdff dff_A_IS805HAQ7_0(.din(n13330), .dout(n13327));
    jdff dff_A_UFxIPcbP1_0(.din(n13333), .dout(n13330));
    jdff dff_A_yetBByJb6_0(.din(n13336), .dout(n13333));
    jdff dff_A_ZQPQV9Ht5_0(.din(n13339), .dout(n13336));
    jdff dff_A_fDVTvTrs4_0(.din(n13342), .dout(n13339));
    jdff dff_A_LR0mbwcR8_0(.din(n13345), .dout(n13342));
    jdff dff_A_WnKG3TWf8_0(.din(n13348), .dout(n13345));
    jdff dff_A_x4xG804r2_0(.din(n13351), .dout(n13348));
    jdff dff_A_rXbJPyvP6_0(.din(n13354), .dout(n13351));
    jdff dff_A_YUovUFfc3_0(.din(n13357), .dout(n13354));
    jdff dff_A_oDpyawyB1_0(.din(n13360), .dout(n13357));
    jdff dff_A_J66xRmJJ2_0(.din(n13363), .dout(n13360));
    jdff dff_A_bvfMJeKd6_0(.din(n13366), .dout(n13363));
    jdff dff_A_qbs6oP5o0_0(.din(n13369), .dout(n13366));
    jdff dff_A_mMtwPRWV7_0(.din(n13372), .dout(n13369));
    jdff dff_A_9hRxczGh1_0(.din(n13375), .dout(n13372));
    jdff dff_A_2OlbOgEd7_0(.din(n13378), .dout(n13375));
    jdff dff_A_U03xe2o77_0(.din(n983), .dout(n13378));
    jdff dff_B_Yv1yDio26_1(.din(n942), .dout(n13382));
    jdff dff_B_GMRm2J0a2_1(.din(n13382), .dout(n13385));
    jdff dff_A_DgLoT3Cl6_0(.din(n13390), .dout(n13387));
    jdff dff_A_EeUnnpzw5_0(.din(n13393), .dout(n13390));
    jdff dff_A_heQPLmxD8_0(.din(n968), .dout(n13393));
    jdff dff_A_HhlvpK5i5_2(.din(n13399), .dout(n13396));
    jdff dff_A_8J2edwd05_2(.din(n968), .dout(n13399));
    jdff dff_A_wEhkXbVQ8_1(.din(n13405), .dout(n13402));
    jdff dff_A_hoEmSdRR5_1(.din(n13408), .dout(n13405));
    jdff dff_A_Yqac6JF91_1(.din(n13411), .dout(n13408));
    jdff dff_A_cQq5FWtM1_1(.din(n13414), .dout(n13411));
    jdff dff_A_kkyJwqUr4_1(.din(n13417), .dout(n13414));
    jdff dff_A_MVluvxhh8_1(.din(n13420), .dout(n13417));
    jdff dff_A_JqRgh5A39_1(.din(n13423), .dout(n13420));
    jdff dff_A_XAPlT4QL3_1(.din(n13426), .dout(n13423));
    jdff dff_A_uH5x4HXz4_1(.din(n13429), .dout(n13426));
    jdff dff_A_JDkxCPk02_1(.din(n13432), .dout(n13429));
    jdff dff_A_EU9PD6dJ6_1(.din(n13435), .dout(n13432));
    jdff dff_A_nlTJAkyk4_1(.din(n13438), .dout(n13435));
    jdff dff_A_ihrt3K1E9_1(.din(n13441), .dout(n13438));
    jdff dff_A_Xijo1cgG4_1(.din(n13444), .dout(n13441));
    jdff dff_A_dkJWDnAp9_1(.din(n13447), .dout(n13444));
    jdff dff_A_28sMcNK85_1(.din(n13450), .dout(n13447));
    jdff dff_A_OMaqpi0d6_1(.din(n13453), .dout(n13450));
    jdff dff_A_j1cVR0RX7_1(.din(n13456), .dout(n13453));
    jdff dff_A_ks5Qe54q5_1(.din(n13459), .dout(n13456));
    jdff dff_A_4dWtdapo3_1(.din(n13462), .dout(n13459));
    jdff dff_A_zpqqx4lL9_1(.din(n13465), .dout(n13462));
    jdff dff_A_xLymxBEh4_1(.din(n13468), .dout(n13465));
    jdff dff_A_FquwOoCd0_1(.din(n13471), .dout(n13468));
    jdff dff_A_JIc1SOCK2_1(.din(n953), .dout(n13471));
    jdff dff_A_GqDk9loR0_0(.din(n13477), .dout(n13474));
    jdff dff_A_4Le9nGDZ9_0(.din(n13480), .dout(n13477));
    jdff dff_A_OS89iIST8_0(.din(n13483), .dout(n13480));
    jdff dff_A_MBUxQrmc6_0(.din(n13486), .dout(n13483));
    jdff dff_A_oFywIdMs1_0(.din(n13489), .dout(n13486));
    jdff dff_A_GRSvb2ma3_0(.din(n13492), .dout(n13489));
    jdff dff_A_VLOtDGPW1_0(.din(n13495), .dout(n13492));
    jdff dff_A_5ucflLL96_0(.din(n13498), .dout(n13495));
    jdff dff_A_zZEu0zwH3_0(.din(n13501), .dout(n13498));
    jdff dff_A_s0PqEE7h4_0(.din(n13504), .dout(n13501));
    jdff dff_A_bsGkyXTe7_0(.din(n13507), .dout(n13504));
    jdff dff_A_3b34rWmF2_0(.din(n13510), .dout(n13507));
    jdff dff_A_zJq1VtZc4_0(.din(n13513), .dout(n13510));
    jdff dff_A_66Rg3Y1y9_0(.din(n13516), .dout(n13513));
    jdff dff_A_ScUGOy2X8_0(.din(n13519), .dout(n13516));
    jdff dff_A_dKUNbawA1_0(.din(n13522), .dout(n13519));
    jdff dff_A_a5IIealN0_0(.din(n13525), .dout(n13522));
    jdff dff_A_uNdcLaJw2_0(.din(n13528), .dout(n13525));
    jdff dff_A_Nm6jfFKM7_0(.din(n13531), .dout(n13528));
    jdff dff_A_ONH35l2Y7_0(.din(n13534), .dout(n13531));
    jdff dff_A_99OCfEXo9_0(.din(n13537), .dout(n13534));
    jdff dff_A_NTePZsvj2_0(.din(n931), .dout(n13537));
    jdff dff_A_7x6e1Cwz1_2(.din(n13543), .dout(n13540));
    jdff dff_A_h0mCwTHF4_2(.din(n13546), .dout(n13543));
    jdff dff_A_a2L6b9wV5_2(.din(n13549), .dout(n13546));
    jdff dff_A_RIidhpSp9_2(.din(n13552), .dout(n13549));
    jdff dff_A_FUPkHfDt6_2(.din(n13555), .dout(n13552));
    jdff dff_A_Z8wG2pGa3_2(.din(n13558), .dout(n13555));
    jdff dff_A_3nBVnkpo2_2(.din(n13561), .dout(n13558));
    jdff dff_A_y1aQQWlZ6_2(.din(n13564), .dout(n13561));
    jdff dff_A_1vWIW1Rv9_2(.din(n13567), .dout(n13564));
    jdff dff_A_UpnmtUR61_2(.din(n13570), .dout(n13567));
    jdff dff_A_99gaBX5H7_2(.din(n13573), .dout(n13570));
    jdff dff_A_SJJq44Bw8_2(.din(n13576), .dout(n13573));
    jdff dff_A_uc3cELp54_2(.din(n13579), .dout(n13576));
    jdff dff_A_s8lCTllk8_2(.din(n13582), .dout(n13579));
    jdff dff_A_17Tjddwp7_2(.din(n13585), .dout(n13582));
    jdff dff_A_tNy0GlAU6_2(.din(n13588), .dout(n13585));
    jdff dff_A_zr4HOGbH2_2(.din(n13591), .dout(n13588));
    jdff dff_A_zVRQU6PJ5_2(.din(n13594), .dout(n13591));
    jdff dff_A_t0EtXzjT4_2(.din(n13597), .dout(n13594));
    jdff dff_A_dymjYP6Y2_2(.din(n13600), .dout(n13597));
    jdff dff_A_E2nBjFEw2_2(.din(n13603), .dout(n13600));
    jdff dff_A_SKdSkvRK0_2(.din(n13606), .dout(n13603));
    jdff dff_A_oyn8YtEy2_2(.din(n927), .dout(n13606));
    jdff dff_B_tvoDF4FO0_0(.din(n919), .dout(n13610));
    jdff dff_B_0RG5tioS2_0(.din(G147), .dout(n13613));
    jdff dff_A_tpcB4Xpz7_1(.din(n13618), .dout(n13615));
    jdff dff_A_kyLWR7fF2_1(.din(n911), .dout(n13618));
    jdff dff_A_WCVFLqku1_2(.din(n13624), .dout(n13621));
    jdff dff_A_O9ZEuD0F3_2(.din(n911), .dout(n13624));
    jdff dff_A_cxp9Ss3B8_1(.din(n13630), .dout(n13627));
    jdff dff_A_M4kje5Xf9_1(.din(n13633), .dout(n13630));
    jdff dff_A_6v2Rtka73_1(.din(n13636), .dout(n13633));
    jdff dff_A_SR3YcPDr8_1(.din(G2211), .dout(n13636));
    jdff dff_A_PFQbUgFH1_1(.din(n13642), .dout(n13639));
    jdff dff_A_Th03vIP36_1(.din(n13645), .dout(n13642));
    jdff dff_A_ZKmtSBG20_1(.din(n13648), .dout(n13645));
    jdff dff_A_RkLwn8DP2_1(.din(n13651), .dout(n13648));
    jdff dff_A_TTpxHY2E4_1(.din(n13654), .dout(n13651));
    jdff dff_A_C2fZkQEP0_1(.din(n13657), .dout(n13654));
    jdff dff_A_0xmRz43N0_1(.din(n13660), .dout(n13657));
    jdff dff_A_2RU396mk8_1(.din(n13663), .dout(n13660));
    jdff dff_A_jNqaqBZC6_1(.din(n13666), .dout(n13663));
    jdff dff_A_jJlfJYnV6_1(.din(n13669), .dout(n13666));
    jdff dff_A_jN5FDuS95_1(.din(n13672), .dout(n13669));
    jdff dff_A_nyXxN85x1_1(.din(n13675), .dout(n13672));
    jdff dff_A_EZt5qb8B7_1(.din(n13678), .dout(n13675));
    jdff dff_A_7X9AVkNe8_1(.din(n13681), .dout(n13678));
    jdff dff_A_iQ8Yl5Ej1_1(.din(n13684), .dout(n13681));
    jdff dff_A_ROcfoLcr4_1(.din(n13687), .dout(n13684));
    jdff dff_A_vSmminsJ0_1(.din(n13690), .dout(n13687));
    jdff dff_A_NUDMmJ1L5_1(.din(n13693), .dout(n13690));
    jdff dff_A_a5HHw5Zd5_1(.din(n13696), .dout(n13693));
    jdff dff_A_o38x5oMh6_1(.din(n13699), .dout(n13696));
    jdff dff_A_VmET2hKb8_1(.din(n13702), .dout(n13699));
    jdff dff_A_YNAHWE8k5_1(.din(n13705), .dout(n13702));
    jdff dff_A_y5Wqknl02_1(.din(n13708), .dout(n13705));
    jdff dff_A_UgbKSko40_1(.din(n13711), .dout(n13708));
    jdff dff_A_mti1uzGy6_1(.din(n908), .dout(n13711));
    jdff dff_B_MQuA8mp51_0(.din(n900), .dout(n13715));
    jdff dff_B_i95EsnAB8_0(.din(G138), .dout(n13718));
    jdff dff_A_J2I59kpR2_1(.din(n13723), .dout(n13720));
    jdff dff_A_KfIMhN2W7_1(.din(n892), .dout(n13723));
    jdff dff_A_ZJQ3nsOw6_2(.din(n13729), .dout(n13726));
    jdff dff_A_vtutKMai1_2(.din(n892), .dout(n13729));
    jdff dff_A_sRfhcl926_1(.din(n13735), .dout(n13732));
    jdff dff_A_ihW1BRz73_1(.din(n13738), .dout(n13735));
    jdff dff_A_XHsNrMzL4_1(.din(n13741), .dout(n13738));
    jdff dff_A_MCNX1YCM4_1(.din(G2218), .dout(n13741));
    jdff dff_A_K2FeAn602_1(.din(n13747), .dout(n13744));
    jdff dff_A_lkVNIif41_1(.din(n13750), .dout(n13747));
    jdff dff_A_5OAbYRuu6_1(.din(n13753), .dout(n13750));
    jdff dff_A_m59Tvl0e4_1(.din(n13756), .dout(n13753));
    jdff dff_A_3B1BqbPB2_1(.din(n13759), .dout(n13756));
    jdff dff_A_KcalhAAw7_1(.din(n13762), .dout(n13759));
    jdff dff_A_126Nwlt32_1(.din(n13765), .dout(n13762));
    jdff dff_A_8gbLF7Hy3_1(.din(n13768), .dout(n13765));
    jdff dff_A_8R3nUI8J7_1(.din(n13771), .dout(n13768));
    jdff dff_A_XbsvL4823_1(.din(n13774), .dout(n13771));
    jdff dff_A_9xyuKzU62_1(.din(n13777), .dout(n13774));
    jdff dff_A_sqdGKtFa8_1(.din(n13780), .dout(n13777));
    jdff dff_A_1KBnA3xU1_1(.din(n13783), .dout(n13780));
    jdff dff_A_JrGpFuJX4_1(.din(n13786), .dout(n13783));
    jdff dff_A_vkXhnAcW9_1(.din(n13789), .dout(n13786));
    jdff dff_A_oxU45Yxl4_1(.din(n13792), .dout(n13789));
    jdff dff_A_XhlpIIz80_1(.din(n13795), .dout(n13792));
    jdff dff_A_EKDNYNzA3_1(.din(n13798), .dout(n13795));
    jdff dff_A_S6jx6gYA3_1(.din(n13801), .dout(n13798));
    jdff dff_A_Z31eQSZF6_1(.din(n13804), .dout(n13801));
    jdff dff_A_DZZnkvIi2_1(.din(n13807), .dout(n13804));
    jdff dff_A_9cFfsQxC2_1(.din(n13810), .dout(n13807));
    jdff dff_A_qogrGZcT3_1(.din(n13813), .dout(n13810));
    jdff dff_A_O3raPL9z5_1(.din(n13816), .dout(n13813));
    jdff dff_A_5A8AnfSW3_1(.din(n889), .dout(n13816));
    jdff dff_A_PvTO2xKm6_2(.din(n889), .dout(n13819));
    jdff dff_A_u8HoK95L0_1(.din(n885), .dout(n13822));
    jdff dff_B_s4eA4dZI1_0(.din(n881), .dout(n13826));
    jdff dff_B_FXRdcySs7_0(.din(G144), .dout(n13829));
    jdff dff_B_1p7mmdux0_2(.din(n873), .dout(n13832));
    jdff dff_B_JpelzHeC9_2(.din(n13832), .dout(n13835));
    jdff dff_A_M8I6GfXi6_0(.din(n13840), .dout(n13837));
    jdff dff_A_NQpzEZHc9_0(.din(n13843), .dout(n13840));
    jdff dff_A_ihlNcuCP0_0(.din(n13846), .dout(n13843));
    jdff dff_A_hBAC02z23_0(.din(G2224), .dout(n13846));
    jdff dff_A_cjpTw9ug5_1(.din(n13862), .dout(n13849));
    jdff dff_B_VNDBVOTU3_2(.din(n870), .dout(n13853));
    jdff dff_B_RtRPpRmP0_2(.din(n13853), .dout(n13856));
    jdff dff_B_VqLeReC87_2(.din(n13856), .dout(n13859));
    jdff dff_B_La6GKKE27_2(.din(n13859), .dout(n13862));
    jdff dff_A_HnBWU2jf4_1(.din(n13867), .dout(n13864));
    jdff dff_A_1Vt5rRGr6_1(.din(n13870), .dout(n13867));
    jdff dff_A_Dgt347V98_1(.din(n13873), .dout(n13870));
    jdff dff_A_aLjvMWy45_1(.din(n13876), .dout(n13873));
    jdff dff_A_nwifDyRU6_1(.din(n13879), .dout(n13876));
    jdff dff_A_M8CUetKr4_1(.din(n13882), .dout(n13879));
    jdff dff_A_UffxN78d5_1(.din(n13885), .dout(n13882));
    jdff dff_A_p7TklzM11_1(.din(n13888), .dout(n13885));
    jdff dff_A_lu1XPUva1_1(.din(n13891), .dout(n13888));
    jdff dff_A_xUke9Sjr9_1(.din(n13894), .dout(n13891));
    jdff dff_A_N7g21i1s1_1(.din(n13897), .dout(n13894));
    jdff dff_A_ZS28p3fN6_1(.din(n13900), .dout(n13897));
    jdff dff_A_76zefZ4f4_1(.din(n13903), .dout(n13900));
    jdff dff_A_hVXxn5s43_1(.din(n13906), .dout(n13903));
    jdff dff_A_vvj5LD029_1(.din(n13909), .dout(n13906));
    jdff dff_A_FR1jVPtN9_1(.din(n13912), .dout(n13909));
    jdff dff_A_6A0JHep92_1(.din(n13915), .dout(n13912));
    jdff dff_A_0VlJsJY14_1(.din(n13918), .dout(n13915));
    jdff dff_A_IBc3Xsp34_1(.din(n13921), .dout(n13918));
    jdff dff_A_VlQXuF739_1(.din(n13924), .dout(n13921));
    jdff dff_A_zq2jNuoz6_1(.din(n13927), .dout(n13924));
    jdff dff_A_BWZ39dDq9_1(.din(n13930), .dout(n13927));
    jdff dff_A_xPtfVNsz4_1(.din(n13933), .dout(n13930));
    jdff dff_A_Bu5drJXT4_1(.din(n13936), .dout(n13933));
    jdff dff_A_z48JbY1H5_1(.din(n13939), .dout(n13936));
    jdff dff_A_4UQNzWyN7_1(.din(n866), .dout(n13939));
    jdff dff_A_TYg8Tdpr4_0(.din(n13945), .dout(n13942));
    jdff dff_A_jMkhOUGu5_0(.din(n13948), .dout(n13945));
    jdff dff_A_9ygve7a99_0(.din(n13951), .dout(n13948));
    jdff dff_A_bDWqOgy68_0(.din(n13954), .dout(n13951));
    jdff dff_A_4wlQ1R3V9_0(.din(n13957), .dout(n13954));
    jdff dff_A_h1X0O4xv7_0(.din(n13960), .dout(n13957));
    jdff dff_A_3zzVk0uX3_0(.din(n13963), .dout(n13960));
    jdff dff_A_RI2R0slG6_0(.din(n13966), .dout(n13963));
    jdff dff_A_aZaxS6Bx2_0(.din(n13969), .dout(n13966));
    jdff dff_A_H1S0Lj2M4_0(.din(n13972), .dout(n13969));
    jdff dff_A_GRgmCoC55_0(.din(n13975), .dout(n13972));
    jdff dff_A_qQkC2sPC0_0(.din(n13978), .dout(n13975));
    jdff dff_A_hEXqIV035_0(.din(n13981), .dout(n13978));
    jdff dff_A_CAsVwaVG4_0(.din(n13984), .dout(n13981));
    jdff dff_A_ntPRJ1Yt2_0(.din(n13987), .dout(n13984));
    jdff dff_A_UfHD95A03_0(.din(n13990), .dout(n13987));
    jdff dff_A_xwjjFYpY0_0(.din(n13993), .dout(n13990));
    jdff dff_A_HY38IcR00_0(.din(n13996), .dout(n13993));
    jdff dff_A_lgy4JPt34_0(.din(n13999), .dout(n13996));
    jdff dff_A_vL5RymjX7_0(.din(n14002), .dout(n13999));
    jdff dff_A_dhVN3lCB6_0(.din(n14005), .dout(n14002));
    jdff dff_A_prACCyXJ7_0(.din(n14008), .dout(n14005));
    jdff dff_A_rz6XL2OO5_0(.din(n14011), .dout(n14008));
    jdff dff_A_u4ZDMtqK4_0(.din(n14014), .dout(n14011));
    jdff dff_A_28w2Jigz5_0(.din(n14017), .dout(n14014));
    jdff dff_A_cP91ZrdY0_0(.din(n14020), .dout(n14017));
    jdff dff_A_ADIvEDMc5_0(.din(n14023), .dout(n14020));
    jdff dff_A_NO57E4si4_0(.din(n862), .dout(n14023));
    jdff dff_A_31WWWRHU3_1(.din(n14029), .dout(n14026));
    jdff dff_A_1aLQFsMz9_1(.din(n14032), .dout(n14029));
    jdff dff_A_QVBtoqvc1_1(.din(n862), .dout(n14032));
    jdff dff_A_xC4ZM0WA6_2(.din(n14038), .dout(n14035));
    jdff dff_A_QF1WnZsW7_2(.din(n14041), .dout(n14038));
    jdff dff_A_Dujt7ChK9_2(.din(n14044), .dout(n14041));
    jdff dff_A_iJUqX09N6_2(.din(n862), .dout(n14044));
    jdff dff_A_g2m1xBFl8_1(.din(n14050), .dout(n14047));
    jdff dff_A_B0oME9l07_1(.din(n14053), .dout(n14050));
    jdff dff_A_9jqs9Xlx5_1(.din(n14056), .dout(n14053));
    jdff dff_A_uaDqfkQw2_1(.din(n14059), .dout(n14056));
    jdff dff_A_IvlrDlFz0_1(.din(n14062), .dout(n14059));
    jdff dff_A_vWMoivkc3_1(.din(n14065), .dout(n14062));
    jdff dff_A_OU0AZkxh6_1(.din(n14068), .dout(n14065));
    jdff dff_A_hOFzT9tM4_1(.din(n14071), .dout(n14068));
    jdff dff_A_kXitvI2w6_1(.din(n14074), .dout(n14071));
    jdff dff_A_kEHsHiiy8_1(.din(n14077), .dout(n14074));
    jdff dff_A_igPE98EO4_1(.din(n14080), .dout(n14077));
    jdff dff_A_MdzvNzrV6_1(.din(n14083), .dout(n14080));
    jdff dff_A_FhSiNrK38_1(.din(n14086), .dout(n14083));
    jdff dff_A_aH8OxooQ2_1(.din(n14089), .dout(n14086));
    jdff dff_A_Qu7i0AOX5_1(.din(n14092), .dout(n14089));
    jdff dff_A_KUTh1DLr8_1(.din(n14095), .dout(n14092));
    jdff dff_A_Ua2Ycfdy6_1(.din(n14098), .dout(n14095));
    jdff dff_A_gHT68AVI8_1(.din(n14101), .dout(n14098));
    jdff dff_A_qNbB8PSW1_1(.din(n14104), .dout(n14101));
    jdff dff_A_pmqbbcJL1_1(.din(n14107), .dout(n14104));
    jdff dff_A_X9cBIOx54_1(.din(n858), .dout(n14107));
    jdff dff_A_5Z81xz2U1_2(.din(n14113), .dout(n14110));
    jdff dff_A_LnyJASmM1_2(.din(n14116), .dout(n14113));
    jdff dff_A_j0ldxZUh0_2(.din(n14119), .dout(n14116));
    jdff dff_A_HIduge0I7_2(.din(n14122), .dout(n14119));
    jdff dff_A_l6iDbYvx2_2(.din(n858), .dout(n14122));
    jdff dff_B_ROfqi5sd5_1(.din(n827), .dout(n14126));
    jdff dff_A_r9uNt09E4_0(.din(n14131), .dout(n14128));
    jdff dff_A_rkdl9ovW0_0(.din(n14134), .dout(n14131));
    jdff dff_A_RK9WZi2Q1_0(.din(n14137), .dout(n14134));
    jdff dff_A_43ymp5HH0_0(.din(n14140), .dout(n14137));
    jdff dff_A_PlUjBCk18_0(.din(n14143), .dout(n14140));
    jdff dff_A_nalhsrNs8_0(.din(n14146), .dout(n14143));
    jdff dff_A_gTodIcZt1_0(.din(n14149), .dout(n14146));
    jdff dff_A_0c4x3L2H1_0(.din(n14152), .dout(n14149));
    jdff dff_A_8Wunz3Gz6_0(.din(n14155), .dout(n14152));
    jdff dff_A_F96IB2Yj5_0(.din(n14158), .dout(n14155));
    jdff dff_A_cVlb8Lai2_0(.din(n14161), .dout(n14158));
    jdff dff_A_q4kPMBVf3_0(.din(n14164), .dout(n14161));
    jdff dff_A_7ecolecs9_0(.din(n14167), .dout(n14164));
    jdff dff_A_dLJrDbS01_0(.din(n14170), .dout(n14167));
    jdff dff_A_YNLs3Fpt1_0(.din(n14173), .dout(n14170));
    jdff dff_A_nWYj38gu5_0(.din(n14176), .dout(n14173));
    jdff dff_A_fjHQlS0k7_0(.din(n14179), .dout(n14176));
    jdff dff_A_FmFN1t1E6_0(.din(n14182), .dout(n14179));
    jdff dff_A_07zxERxa6_0(.din(n14185), .dout(n14182));
    jdff dff_A_hE3TMeAi0_0(.din(n14188), .dout(n14185));
    jdff dff_A_vf7Phuzu2_0(.din(n14191), .dout(n14188));
    jdff dff_A_1k4KbDb68_0(.din(n14194), .dout(n14191));
    jdff dff_A_wAN75iSl7_0(.din(n14197), .dout(n14194));
    jdff dff_A_YRBUIWw11_0(.din(n14200), .dout(n14197));
    jdff dff_A_9lgaDUz22_0(.din(n14203), .dout(n14200));
    jdff dff_A_HkY0Ozwo5_0(.din(n14206), .dout(n14203));
    jdff dff_A_pC9SxTcg1_0(.din(n14209), .dout(n14206));
    jdff dff_A_wPtHeeCc1_0(.din(n850), .dout(n14209));
    jdff dff_A_3ZpI47qr9_1(.din(n14215), .dout(n14212));
    jdff dff_A_bFQNGcgB9_1(.din(n14218), .dout(n14215));
    jdff dff_A_MZshv5gh3_1(.din(n14221), .dout(n14218));
    jdff dff_A_TwH1swP31_1(.din(n14224), .dout(n14221));
    jdff dff_A_8HORNGw25_1(.din(n14227), .dout(n14224));
    jdff dff_A_xFMB9gpv5_1(.din(n14230), .dout(n14227));
    jdff dff_A_5NdSYsBJ7_1(.din(n14233), .dout(n14230));
    jdff dff_A_vcR82Vn03_1(.din(n14236), .dout(n14233));
    jdff dff_A_reVZ7qnZ6_1(.din(n14239), .dout(n14236));
    jdff dff_A_DrHrwRI04_1(.din(n14242), .dout(n14239));
    jdff dff_A_tbLMEGHm9_1(.din(n14245), .dout(n14242));
    jdff dff_A_0u21JPMa1_1(.din(n14248), .dout(n14245));
    jdff dff_A_9W78x3VH4_1(.din(n14251), .dout(n14248));
    jdff dff_A_oHtssPdj0_1(.din(n14254), .dout(n14251));
    jdff dff_A_C2oswGKJ7_1(.din(n14257), .dout(n14254));
    jdff dff_A_ez8dfd7Z7_1(.din(n14260), .dout(n14257));
    jdff dff_A_V8dlpBUk4_1(.din(n14263), .dout(n14260));
    jdff dff_A_y6e35GZE3_1(.din(n14266), .dout(n14263));
    jdff dff_A_YErLJ0Y63_1(.din(n14269), .dout(n14266));
    jdff dff_A_JWPlhfRX4_1(.din(n14272), .dout(n14269));
    jdff dff_A_oghk7Wwo4_1(.din(n14275), .dout(n14272));
    jdff dff_A_ZE5QrrRW7_1(.din(n14278), .dout(n14275));
    jdff dff_A_jiaZanyy9_1(.din(n14281), .dout(n14278));
    jdff dff_A_qTxX4T0S2_1(.din(n14284), .dout(n14281));
    jdff dff_A_Ni3xbxCS0_1(.din(n14287), .dout(n14284));
    jdff dff_A_D5Uy5jKu4_1(.din(n14290), .dout(n14287));
    jdff dff_A_6Hqpq9og1_1(.din(n850), .dout(n14290));
    jdff dff_A_hi7zk1CR7_1(.din(n14296), .dout(n14293));
    jdff dff_A_LF35YLmI6_1(.din(n14299), .dout(n14296));
    jdff dff_A_zcRclED08_1(.din(n14302), .dout(n14299));
    jdff dff_A_fJ6Z2Fym0_1(.din(n14305), .dout(n14302));
    jdff dff_A_H6YW1Fir0_1(.din(n14308), .dout(n14305));
    jdff dff_A_ELfZLHUX2_1(.din(n850), .dout(n14308));
    jdff dff_A_tbc2fNk24_2(.din(n14314), .dout(n14311));
    jdff dff_A_ZO8xir4g0_2(.din(n14317), .dout(n14314));
    jdff dff_A_llcSN2BG4_2(.din(n14320), .dout(n14317));
    jdff dff_A_pUa3w54x3_2(.din(n14323), .dout(n14320));
    jdff dff_A_g3dRlHVv4_2(.din(n14326), .dout(n14323));
    jdff dff_A_4iMejImJ9_2(.din(n14329), .dout(n14326));
    jdff dff_A_9WxyhcV15_2(.din(n850), .dout(n14329));
    jdff dff_B_4ktNGoya8_0(.din(n842), .dout(n14333));
    jdff dff_B_W1sljb7y0_0(.din(G135), .dout(n14336));
    jdff dff_A_K55uznzv1_1(.din(n14341), .dout(n14338));
    jdff dff_A_JnxynNQZ7_1(.din(n834), .dout(n14341));
    jdff dff_A_iSt3pmoL4_2(.din(n14347), .dout(n14344));
    jdff dff_A_fzA0RuAB8_2(.din(n834), .dout(n14347));
    jdff dff_A_62mwjYD83_1(.din(n14353), .dout(n14350));
    jdff dff_A_KHSdDUvG7_1(.din(n14356), .dout(n14353));
    jdff dff_A_WpstJHKE4_1(.din(n14359), .dout(n14356));
    jdff dff_A_cqRjat6f7_1(.din(G2230), .dout(n14359));
    jdff dff_A_tqesnuAW6_1(.din(n823), .dout(n14362));
    jdff dff_B_1NhAGwVz7_0(.din(G157), .dout(n14366));
    jdff dff_B_K5txonfB4_3(.din(n815), .dout(n14369));
    jdff dff_B_ZTy8EqPV4_3(.din(n14369), .dout(n14372));
    jdff dff_A_MbeNTaRo8_2(.din(n14377), .dout(n14374));
    jdff dff_A_VqFYbCB53_2(.din(n14380), .dout(n14377));
    jdff dff_A_tg13M2sT7_2(.din(n14383), .dout(n14380));
    jdff dff_A_6XrtcXTY6_2(.din(n14386), .dout(n14383));
    jdff dff_A_jPNMqTsu8_2(.din(n14389), .dout(n14386));
    jdff dff_A_iMez3pks7_2(.din(n14392), .dout(n14389));
    jdff dff_A_ZwyOmiDg8_2(.din(n14395), .dout(n14392));
    jdff dff_A_1pWxHSlY1_2(.din(n14398), .dout(n14395));
    jdff dff_A_JDyQ9ai18_2(.din(n14401), .dout(n14398));
    jdff dff_A_iR6B7duH2_2(.din(n14404), .dout(n14401));
    jdff dff_A_OaDpa0iQ4_2(.din(n14407), .dout(n14404));
    jdff dff_A_dyS1aMqS3_2(.din(n14410), .dout(n14407));
    jdff dff_A_6pCGcHdt6_2(.din(n14413), .dout(n14410));
    jdff dff_A_yYbDhjX34_2(.din(n14416), .dout(n14413));
    jdff dff_A_hQ8yQrNP2_2(.din(n14419), .dout(n14416));
    jdff dff_A_41mxgmIB7_2(.din(n14422), .dout(n14419));
    jdff dff_A_pYHGwCkf2_2(.din(n14425), .dout(n14422));
    jdff dff_A_2D8usgXT5_2(.din(n14428), .dout(n14425));
    jdff dff_A_hYOCOZMz8_2(.din(n14431), .dout(n14428));
    jdff dff_A_FQOKUYsv5_2(.din(n14434), .dout(n14431));
    jdff dff_A_BfJp3bsu6_2(.din(n14437), .dout(n14434));
    jdff dff_A_yOGMEFVi3_2(.din(n812), .dout(n14437));
    jdff dff_B_bEDm3zYn1_1(.din(n770), .dout(n14441));
    jdff dff_B_BiI0ZTCU1_1(.din(n14441), .dout(n14444));
    jdff dff_A_wjKWvZBb3_0(.din(n14449), .dout(n14446));
    jdff dff_A_dJgKxRIC5_0(.din(n14452), .dout(n14449));
    jdff dff_A_1ZBRyKC30_0(.din(n14455), .dout(n14452));
    jdff dff_A_cVv02Nlj1_0(.din(n14458), .dout(n14455));
    jdff dff_A_rRkeo3GP2_0(.din(n14461), .dout(n14458));
    jdff dff_A_bldm7o9G6_0(.din(n14464), .dout(n14461));
    jdff dff_A_sBerXbpX6_0(.din(n14467), .dout(n14464));
    jdff dff_A_kEVfi8W48_0(.din(n14470), .dout(n14467));
    jdff dff_A_itbCi6411_0(.din(n14473), .dout(n14470));
    jdff dff_A_ePQy4ze88_0(.din(n14476), .dout(n14473));
    jdff dff_A_gpQCK13v9_0(.din(n14479), .dout(n14476));
    jdff dff_A_VgxrRdz78_0(.din(n14482), .dout(n14479));
    jdff dff_A_2ObhRrl09_0(.din(n14485), .dout(n14482));
    jdff dff_A_2D63Mkir0_0(.din(n14488), .dout(n14485));
    jdff dff_A_ssscaKOB5_0(.din(n14491), .dout(n14488));
    jdff dff_A_YYVbMTHo0_0(.din(n14494), .dout(n14491));
    jdff dff_A_YoUP7csR4_0(.din(n14497), .dout(n14494));
    jdff dff_A_RHxQU68j4_0(.din(n14500), .dout(n14497));
    jdff dff_A_Ol441Uz21_0(.din(n14503), .dout(n14500));
    jdff dff_A_bxayRSXS9_0(.din(n14506), .dout(n14503));
    jdff dff_A_KChkSnBZ2_0(.din(n14509), .dout(n14506));
    jdff dff_A_YDSTlRFl9_0(.din(n808), .dout(n14509));
    jdff dff_B_pVUVu6oE9_1(.din(n780), .dout(n14513));
    jdff dff_B_VEsaFXyh2_1(.din(n784), .dout(n14516));
    jdff dff_B_2P3d0CEE3_1(.din(n14516), .dout(n14519));
    jdff dff_A_Yx4risHu8_1(.din(n14524), .dout(n14521));
    jdff dff_A_LPyXdJn96_1(.din(n14527), .dout(n14524));
    jdff dff_A_YRV2LOo14_1(.din(n14530), .dout(n14527));
    jdff dff_A_jPrX1cbm8_1(.din(n14533), .dout(n14530));
    jdff dff_A_BQ09mqDV6_1(.din(n14536), .dout(n14533));
    jdff dff_A_hnGbZB4c2_1(.din(n14539), .dout(n14536));
    jdff dff_A_LoWAeYgW8_1(.din(n14542), .dout(n14539));
    jdff dff_A_aga1Qr7U6_1(.din(n14545), .dout(n14542));
    jdff dff_A_E6b3rdbL2_1(.din(n14548), .dout(n14545));
    jdff dff_A_H2JKbEBc0_1(.din(n14551), .dout(n14548));
    jdff dff_A_tHGxxEfW7_1(.din(n14554), .dout(n14551));
    jdff dff_A_SV50TXc59_1(.din(n14557), .dout(n14554));
    jdff dff_A_ZCa0qgEb5_1(.din(n14560), .dout(n14557));
    jdff dff_A_seWYdYZu5_1(.din(n14563), .dout(n14560));
    jdff dff_A_esdau1Ez5_1(.din(n14566), .dout(n14563));
    jdff dff_A_88KGpDJV7_1(.din(n14569), .dout(n14566));
    jdff dff_A_sKYU1zDx5_1(.din(n14572), .dout(n14569));
    jdff dff_A_o83YnuwY8_1(.din(n14575), .dout(n14572));
    jdff dff_A_Tp2bWoNb3_1(.din(n14578), .dout(n14575));
    jdff dff_A_hXMuAwq23_1(.din(n14581), .dout(n14578));
    jdff dff_A_aNHrWs2m3_1(.din(n14584), .dout(n14581));
    jdff dff_A_DCRuM31d7_1(.din(n14587), .dout(n14584));
    jdff dff_A_cYntFtSi4_1(.din(n14590), .dout(n14587));
    jdff dff_A_kiwYSKer5_1(.din(n14593), .dout(n14590));
    jdff dff_A_DBXmQNFG7_1(.din(n800), .dout(n14593));
    jdff dff_A_7PWrwykw5_1(.din(n14599), .dout(n14596));
    jdff dff_A_tVTt4gd04_1(.din(n14602), .dout(n14599));
    jdff dff_A_gLGe0Teh8_1(.din(n14605), .dout(n14602));
    jdff dff_A_9zluSdTd1_1(.din(n14608), .dout(n14605));
    jdff dff_A_tlvcJgdQ4_1(.din(n14611), .dout(n14608));
    jdff dff_A_SJerHwCp5_1(.din(n14614), .dout(n14611));
    jdff dff_A_O0RnGL9Z6_1(.din(n14617), .dout(n14614));
    jdff dff_A_8c5mLC0Q5_1(.din(n14620), .dout(n14617));
    jdff dff_A_iUP3jbLH0_1(.din(n14623), .dout(n14620));
    jdff dff_A_iLH3P6Ny7_1(.din(n14626), .dout(n14623));
    jdff dff_A_iraFo22z3_1(.din(n14629), .dout(n14626));
    jdff dff_A_BIz3xtaL1_1(.din(n14632), .dout(n14629));
    jdff dff_A_9wo9M0UM2_1(.din(n14635), .dout(n14632));
    jdff dff_A_ZlWK9vG67_1(.din(n14638), .dout(n14635));
    jdff dff_A_mrAwvEfd2_1(.din(n14641), .dout(n14638));
    jdff dff_A_RW5hLxVc4_1(.din(n14644), .dout(n14641));
    jdff dff_A_5WviFnyq4_1(.din(n14647), .dout(n14644));
    jdff dff_A_Pmjqmfgp6_1(.din(n14650), .dout(n14647));
    jdff dff_A_cW8swT584_1(.din(n14653), .dout(n14650));
    jdff dff_A_yiEcr5Fi0_1(.din(n14656), .dout(n14653));
    jdff dff_A_7fMavj4h1_1(.din(n14659), .dout(n14656));
    jdff dff_A_kMawKvbe0_1(.din(n14662), .dout(n14659));
    jdff dff_A_Wj9KDVlV5_1(.din(n14665), .dout(n14662));
    jdff dff_A_GxaZnX183_1(.din(n14668), .dout(n14665));
    jdff dff_A_Wdxvnsr97_1(.din(n14671), .dout(n14668));
    jdff dff_A_nRvZGQid1_1(.din(n792), .dout(n14671));
    jdff dff_A_vlI9QMAP8_1(.din(n14677), .dout(n14674));
    jdff dff_A_mfUBjL8h2_1(.din(n788), .dout(n14677));
    jdff dff_A_jGvha8wF0_2(.din(n788), .dout(n14680));
    jdff dff_A_kggdpM1j0_0(.din(n14686), .dout(n14683));
    jdff dff_A_0oJUP1386_0(.din(n14689), .dout(n14686));
    jdff dff_A_k5pLKUhv3_0(.din(n14692), .dout(n14689));
    jdff dff_A_mJqz6rnL6_0(.din(n14695), .dout(n14692));
    jdff dff_A_PDW4LpkL6_0(.din(n14698), .dout(n14695));
    jdff dff_A_OmW5Xfae5_0(.din(n14701), .dout(n14698));
    jdff dff_A_EA2hOLsY0_0(.din(n14704), .dout(n14701));
    jdff dff_A_WbU7slYa3_0(.din(n14707), .dout(n14704));
    jdff dff_A_d7qouoRC9_0(.din(n14710), .dout(n14707));
    jdff dff_A_1P1smI3R2_0(.din(n14713), .dout(n14710));
    jdff dff_A_Fg6V4p2y1_0(.din(n14716), .dout(n14713));
    jdff dff_A_ydOLMp6N6_0(.din(n14719), .dout(n14716));
    jdff dff_A_EmUjLuic3_0(.din(n14722), .dout(n14719));
    jdff dff_A_LUvcrnHy4_0(.din(n14725), .dout(n14722));
    jdff dff_A_QTbTcMfe2_0(.din(n14728), .dout(n14725));
    jdff dff_A_xjM7abYy4_0(.din(n14731), .dout(n14728));
    jdff dff_A_g46lyfAZ5_0(.din(n14734), .dout(n14731));
    jdff dff_A_AiEyQROX8_0(.din(n14737), .dout(n14734));
    jdff dff_A_XEDLWGuX6_0(.din(n14740), .dout(n14737));
    jdff dff_A_S0iiNFFp4_0(.din(n14743), .dout(n14740));
    jdff dff_A_sXogL2F34_0(.din(n14746), .dout(n14743));
    jdff dff_A_Hf4XiKpk9_0(.din(n14749), .dout(n14746));
    jdff dff_A_gl02tlid9_0(.din(n14752), .dout(n14749));
    jdff dff_A_2G7fOMRi7_0(.din(n14755), .dout(n14752));
    jdff dff_A_b9i0mVPX4_0(.din(n766), .dout(n14755));
    jdff dff_A_387xNCBw7_1(.din(n14761), .dout(n14758));
    jdff dff_A_mTJizaas6_1(.din(n14764), .dout(n14761));
    jdff dff_A_eBFFZHSR0_1(.din(n14767), .dout(n14764));
    jdff dff_A_m7l1VNKy0_1(.din(n14770), .dout(n14767));
    jdff dff_A_lbqrYRH56_1(.din(n14773), .dout(n14770));
    jdff dff_A_2RPepJyl2_1(.din(n14776), .dout(n14773));
    jdff dff_A_vsDihIaw3_1(.din(n14779), .dout(n14776));
    jdff dff_A_HR0oxJQG8_1(.din(n14782), .dout(n14779));
    jdff dff_A_euFO73gY0_1(.din(n14785), .dout(n14782));
    jdff dff_A_y5wHyyBy4_1(.din(n14788), .dout(n14785));
    jdff dff_A_bTwg9hed6_1(.din(n14791), .dout(n14788));
    jdff dff_A_PUmlXlX87_1(.din(n14794), .dout(n14791));
    jdff dff_A_Tmg5YTKb6_1(.din(n14797), .dout(n14794));
    jdff dff_A_z8vE3lil5_1(.din(n14800), .dout(n14797));
    jdff dff_A_Uu017SPj2_1(.din(n14803), .dout(n14800));
    jdff dff_A_SMs7wOsT4_1(.din(n14806), .dout(n14803));
    jdff dff_A_ozyoaQiE6_1(.din(n14809), .dout(n14806));
    jdff dff_A_ItrCI28u1_1(.din(n14812), .dout(n14809));
    jdff dff_A_LY8xMpdE4_1(.din(n14815), .dout(n14812));
    jdff dff_A_w6LFbHZM6_1(.din(n14818), .dout(n14815));
    jdff dff_A_ydoMcFHd3_1(.din(n14821), .dout(n14818));
    jdff dff_A_zMW1l7rV8_1(.din(n14824), .dout(n14821));
    jdff dff_A_pWMSAPij5_1(.din(n14827), .dout(n14824));
    jdff dff_A_ERRnKHiM3_1(.din(n14830), .dout(n14827));
    jdff dff_A_GVpSceM11_1(.din(n14833), .dout(n14830));
    jdff dff_A_R1lrvgxA0_1(.din(n762), .dout(n14833));
    jdff dff_A_ixPLp55g3_0(.din(n14839), .dout(n14836));
    jdff dff_A_Dxy3LhG70_0(.din(n754), .dout(n14839));
    jdff dff_B_wEA3Mhyp8_0(.din(G156), .dout(n14843));
    jdff dff_B_q2wugx5I4_2(.din(n750), .dout(n14846));
    jdff dff_B_59IVopTg7_2(.din(n14846), .dout(n14849));
    jdff dff_A_3wBuw7q61_2(.din(n14854), .dout(n14851));
    jdff dff_A_nKOwR62T0_2(.din(n14857), .dout(n14854));
    jdff dff_A_AUMhxIV25_2(.din(n14860), .dout(n14857));
    jdff dff_A_LcmCCn9p0_2(.din(G2239), .dout(n14860));
    jdff dff_A_pAmu6KRT6_0(.din(n14866), .dout(n14863));
    jdff dff_A_BdNNkt7t5_0(.din(n14869), .dout(n14866));
    jdff dff_A_GVtHqrqw2_0(.din(n14872), .dout(n14869));
    jdff dff_A_zema3Pci6_0(.din(n14875), .dout(n14872));
    jdff dff_A_pbkPyzqZ3_0(.din(n14878), .dout(n14875));
    jdff dff_A_1snCvRQM9_0(.din(n14881), .dout(n14878));
    jdff dff_A_fvnDjC625_0(.din(n14884), .dout(n14881));
    jdff dff_A_u8A8dzar6_0(.din(n14887), .dout(n14884));
    jdff dff_A_xPZ30kMI6_0(.din(n14890), .dout(n14887));
    jdff dff_A_igY3nnvL2_0(.din(n14893), .dout(n14890));
    jdff dff_A_F5ZTxqAJ1_0(.din(n14896), .dout(n14893));
    jdff dff_A_MTgprWJy7_0(.din(n14899), .dout(n14896));
    jdff dff_A_G0bKuq5s8_0(.din(n14902), .dout(n14899));
    jdff dff_A_RYW8Liwf4_0(.din(n14905), .dout(n14902));
    jdff dff_A_NOoDreEn2_0(.din(n14908), .dout(n14905));
    jdff dff_A_jnJX9vzc5_0(.din(n14911), .dout(n14908));
    jdff dff_A_sH9JF1vV8_0(.din(n14914), .dout(n14911));
    jdff dff_A_NrXAo8iN2_0(.din(n14917), .dout(n14914));
    jdff dff_A_KCGuJm2B2_0(.din(n14920), .dout(n14917));
    jdff dff_A_kfLL1v7W8_0(.din(n14923), .dout(n14920));
    jdff dff_A_GgfWM8fP3_0(.din(n14926), .dout(n14923));
    jdff dff_A_Qqjm0Ki83_0(.din(n14929), .dout(n14926));
    jdff dff_A_2aihjCnZ1_0(.din(n14932), .dout(n14929));
    jdff dff_A_elxtFNZ21_0(.din(n14935), .dout(n14932));
    jdff dff_A_c7ZQRUbS3_0(.din(n14938), .dout(n14935));
    jdff dff_A_Ar18Dr8B6_0(.din(n14941), .dout(n14938));
    jdff dff_A_cd83q31D9_0(.din(n14944), .dout(n14941));
    jdff dff_A_OuOmfGs39_0(.din(n747), .dout(n14944));
    jdff dff_A_UYjlfQK17_2(.din(n14950), .dout(n14947));
    jdff dff_A_YLcjpomc1_2(.din(n14953), .dout(n14950));
    jdff dff_A_yvXqhH371_2(.din(n14956), .dout(n14953));
    jdff dff_A_ky3EWdLW5_2(.din(n747), .dout(n14956));
    jdff dff_A_9FBXsJ5D7_0(.din(n14962), .dout(n14959));
    jdff dff_A_rZYiXbkz5_0(.din(n739), .dout(n14962));
    jdff dff_B_F1xHy1Kr0_0(.din(G155), .dout(n14966));
    jdff dff_B_aLOuqT6y1_2(.din(n735), .dout(n14969));
    jdff dff_B_qfxNow3q4_2(.din(n14969), .dout(n14972));
    jdff dff_A_09Rzbv0n9_1(.din(n14977), .dout(n14974));
    jdff dff_A_zEQnSkvr7_1(.din(n14980), .dout(n14977));
    jdff dff_A_xGnoXxZc2_1(.din(n14983), .dout(n14980));
    jdff dff_A_sg9lbXIo8_1(.din(n14986), .dout(n14983));
    jdff dff_A_H6LTrRNq3_1(.din(n14989), .dout(n14986));
    jdff dff_A_suG4h3MQ2_1(.din(n14992), .dout(n14989));
    jdff dff_A_XwqpMb7r3_1(.din(n14995), .dout(n14992));
    jdff dff_A_gr4pZuZk5_1(.din(n14998), .dout(n14995));
    jdff dff_A_Zezn3gTG3_1(.din(n15001), .dout(n14998));
    jdff dff_A_79D3nSYZ5_1(.din(n15004), .dout(n15001));
    jdff dff_A_0m4mJ7o25_1(.din(n15007), .dout(n15004));
    jdff dff_A_RMSrkFxh6_1(.din(n15010), .dout(n15007));
    jdff dff_A_CmqjsdPN6_1(.din(n15013), .dout(n15010));
    jdff dff_A_fll1kGTT8_1(.din(n15016), .dout(n15013));
    jdff dff_A_4E0of3rE9_1(.din(n15019), .dout(n15016));
    jdff dff_A_moFGrM1t2_1(.din(n15022), .dout(n15019));
    jdff dff_A_Mjxs4LXI1_1(.din(n15025), .dout(n15022));
    jdff dff_A_36A6DOYl2_1(.din(n15028), .dout(n15025));
    jdff dff_A_zF5Nd7pD3_1(.din(n15031), .dout(n15028));
    jdff dff_A_RwvSeBfy3_1(.din(n15034), .dout(n15031));
    jdff dff_A_5gnAqyom9_1(.din(n15037), .dout(n15034));
    jdff dff_A_DhltJnR27_1(.din(n15040), .dout(n15037));
    jdff dff_A_cPYjnrig9_1(.din(n15043), .dout(n15040));
    jdff dff_A_hrEXM8FB1_1(.din(n15046), .dout(n15043));
    jdff dff_A_xddUA2Jw4_1(.din(n15049), .dout(n15046));
    jdff dff_A_cXhmlniw5_1(.din(n15052), .dout(n15049));
    jdff dff_A_1Ymh6j8A3_1(.din(n15055), .dout(n15052));
    jdff dff_A_YUTW2DAO3_1(.din(n732), .dout(n15055));
    jdff dff_A_9gVNd9nX7_2(.din(n732), .dout(n15058));
    jdff dff_A_4arLlfmD9_0(.din(n15064), .dout(n15061));
    jdff dff_A_Etqypq3F7_0(.din(n724), .dout(n15064));
    jdff dff_B_8UG59Vca7_0(.din(G154), .dout(n15068));
    jdff dff_A_QX1Bx6I01_1(.din(n15073), .dout(n15070));
    jdff dff_A_Ggj1yM443_1(.din(n720), .dout(n15073));
    jdff dff_A_HTMGDVHZ1_2(.din(n15079), .dout(n15076));
    jdff dff_A_K5ZBCKeC9_2(.din(n720), .dout(n15079));
    jdff dff_A_DY0byoKN3_1(.din(n15085), .dout(n15082));
    jdff dff_A_poaqWqFO4_1(.din(n15088), .dout(n15085));
    jdff dff_A_otUmM6eA6_1(.din(n15091), .dout(n15088));
    jdff dff_A_Pn0AJcb18_1(.din(G2253), .dout(n15091));
    jdff dff_A_baD3Q3CB8_1(.din(n15097), .dout(n15094));
    jdff dff_A_1R9bhMXu3_1(.din(n15100), .dout(n15097));
    jdff dff_A_wWKFtqNt8_1(.din(n15103), .dout(n15100));
    jdff dff_A_71pj1lpB6_1(.din(n15106), .dout(n15103));
    jdff dff_A_ryRSPHHA3_1(.din(n15109), .dout(n15106));
    jdff dff_A_KavIGZoi1_1(.din(n15112), .dout(n15109));
    jdff dff_A_OjjPaYin5_1(.din(n15115), .dout(n15112));
    jdff dff_A_49iVaXPm4_1(.din(n15118), .dout(n15115));
    jdff dff_A_uL3r89oo2_1(.din(n15121), .dout(n15118));
    jdff dff_A_K5wvCeqg4_1(.din(n15124), .dout(n15121));
    jdff dff_A_8GZUAg3f1_1(.din(n15127), .dout(n15124));
    jdff dff_A_y6Lu6vUt2_1(.din(n15130), .dout(n15127));
    jdff dff_A_yWVwfS0b3_1(.din(n15133), .dout(n15130));
    jdff dff_A_uSkAOhDH6_1(.din(n15136), .dout(n15133));
    jdff dff_A_yh9jPnZQ7_1(.din(n15139), .dout(n15136));
    jdff dff_A_CAjnkr406_1(.din(n15142), .dout(n15139));
    jdff dff_A_bZpG9w7x0_1(.din(n15145), .dout(n15142));
    jdff dff_A_3nTGLdvQ8_1(.din(n15148), .dout(n15145));
    jdff dff_A_Tqr5ye7V0_1(.din(n15151), .dout(n15148));
    jdff dff_A_MrxSu1Kd1_1(.din(n15154), .dout(n15151));
    jdff dff_A_z8TgFc517_1(.din(n15157), .dout(n15154));
    jdff dff_A_iYFIVBXd1_1(.din(n15160), .dout(n15157));
    jdff dff_A_CKmlYBeT8_1(.din(n15163), .dout(n15160));
    jdff dff_A_Lq8qeYY98_1(.din(n15166), .dout(n15163));
    jdff dff_A_AY0Ygbpn0_1(.din(n15169), .dout(n15166));
    jdff dff_A_tR2DfjdY3_1(.din(n15172), .dout(n15169));
    jdff dff_A_udk0DvfK8_1(.din(n15175), .dout(n15172));
    jdff dff_A_fHouZqGt3_1(.din(n717), .dout(n15175));
    jdff dff_A_C5gFqW8C7_2(.din(n15181), .dout(n15178));
    jdff dff_A_AzhajSGA9_2(.din(n15184), .dout(n15181));
    jdff dff_A_anWRxKrp5_2(.din(n15187), .dout(n15184));
    jdff dff_A_CEBS9loZ4_2(.din(n15190), .dout(n15187));
    jdff dff_A_zWpz9K373_2(.din(n15193), .dout(n15190));
    jdff dff_A_tS34ImiE8_2(.din(n15196), .dout(n15193));
    jdff dff_A_i9BEr20I3_2(.din(n15199), .dout(n15196));
    jdff dff_A_6BNDKbQJ5_2(.din(n15202), .dout(n15199));
    jdff dff_A_wHvaS5eP5_2(.din(n15205), .dout(n15202));
    jdff dff_A_2UJBnGw15_2(.din(n15208), .dout(n15205));
    jdff dff_A_YHYPlSnV9_2(.din(n15211), .dout(n15208));
    jdff dff_A_NmpRpQDc7_2(.din(n15214), .dout(n15211));
    jdff dff_A_IIb8Gdv16_2(.din(n15217), .dout(n15214));
    jdff dff_A_QwKkJGS42_2(.din(n15220), .dout(n15217));
    jdff dff_A_FpE1NfNw5_2(.din(n15223), .dout(n15220));
    jdff dff_A_ZAXYdkzJ8_2(.din(n15226), .dout(n15223));
    jdff dff_A_b3I5VCR79_2(.din(n15229), .dout(n15226));
    jdff dff_A_M8tnH8qC1_2(.din(n15232), .dout(n15229));
    jdff dff_A_TzFzFNrV6_2(.din(n15235), .dout(n15232));
    jdff dff_A_xkqkMJMN6_2(.din(n15238), .dout(n15235));
    jdff dff_A_jvauE3K24_2(.din(n15241), .dout(n15238));
    jdff dff_A_QQKBQqh65_2(.din(n15244), .dout(n15241));
    jdff dff_A_tUUVP2Vy9_2(.din(n15247), .dout(n15244));
    jdff dff_A_BHs6HxvU7_2(.din(n15250), .dout(n15247));
    jdff dff_A_VmcHDvd72_2(.din(n15253), .dout(n15250));
    jdff dff_A_U6iUWgwA8_2(.din(n15256), .dout(n15253));
    jdff dff_A_FNcJlQLL3_2(.din(n15259), .dout(n15256));
    jdff dff_A_wqPvJ2r96_2(.din(n717), .dout(n15259));
    jdff dff_A_JPCot2ZB7_1(.din(n15265), .dout(n15262));
    jdff dff_A_L7qavIXQ2_1(.din(n15268), .dout(n15265));
    jdff dff_A_AbUAfjVv8_1(.din(n15271), .dout(n15268));
    jdff dff_A_0vjlAh087_1(.din(n15274), .dout(n15271));
    jdff dff_A_rbzNotZQ9_1(.din(n15277), .dout(n15274));
    jdff dff_A_LIx7qTrD6_1(.din(n15280), .dout(n15277));
    jdff dff_A_TH2h2Jyo1_1(.din(n15283), .dout(n15280));
    jdff dff_A_63KIUd6P4_1(.din(n15286), .dout(n15283));
    jdff dff_A_LytSijHB7_1(.din(n15289), .dout(n15286));
    jdff dff_A_T6Pw4CQE5_1(.din(n15292), .dout(n15289));
    jdff dff_A_FecUEcXq0_1(.din(n15295), .dout(n15292));
    jdff dff_A_jfqI3rik3_1(.din(n15298), .dout(n15295));
    jdff dff_A_2VydCtZr7_1(.din(n15301), .dout(n15298));
    jdff dff_A_RwDE5Bnv0_1(.din(n15304), .dout(n15301));
    jdff dff_A_3wkFOEgy6_1(.din(n15307), .dout(n15304));
    jdff dff_A_r1jNPOol5_1(.din(n15310), .dout(n15307));
    jdff dff_A_qv6uDbQW6_1(.din(n15313), .dout(n15310));
    jdff dff_A_IxbBvkpg9_1(.din(n15316), .dout(n15313));
    jdff dff_A_nM5uXi1V4_1(.din(n15319), .dout(n15316));
    jdff dff_A_xs1WsFzi4_1(.din(n15322), .dout(n15319));
    jdff dff_A_h2OQWkcC5_1(.din(n15325), .dout(n15322));
    jdff dff_A_ZW4vS40h0_1(.din(n15328), .dout(n15325));
    jdff dff_A_BrYgqhBT2_1(.din(n15331), .dout(n15328));
    jdff dff_A_WVcPQJbm0_1(.din(n15334), .dout(n15331));
    jdff dff_A_lFLkfp0b5_1(.din(n15337), .dout(n15334));
    jdff dff_A_y8sCxpDE5_1(.din(n15340), .dout(n15337));
    jdff dff_A_vKkxQUhC6_1(.din(n15343), .dout(n15340));
    jdff dff_A_mXJSl3Zk9_1(.din(n15346), .dout(n15343));
    jdff dff_A_6GHje0Ez4_1(.din(n713), .dout(n15346));
    jdff dff_A_HvRZD6YI7_0(.din(n15352), .dout(n15349));
    jdff dff_A_3oLcbMUW2_0(.din(n705), .dout(n15352));
    jdff dff_B_KrwkUrhI8_0(.din(G153), .dout(n15356));
    jdff dff_A_GKk1bp1A7_1(.din(n15361), .dout(n15358));
    jdff dff_A_J5y6YU0r4_1(.din(n701), .dout(n15361));
    jdff dff_A_dIpyqVQs2_2(.din(n15367), .dout(n15364));
    jdff dff_A_fzPZDmtX3_2(.din(n701), .dout(n15367));
    jdff dff_A_bUrptudo5_1(.din(n15373), .dout(n15370));
    jdff dff_A_aAH0WpaF9_1(.din(n15376), .dout(n15373));
    jdff dff_A_lNPuLJKy0_1(.din(n15379), .dout(n15376));
    jdff dff_A_8RIx3fbU2_1(.din(n15382), .dout(n15379));
    jdff dff_A_40hxMOXx5_1(.din(n15385), .dout(n15382));
    jdff dff_A_Tfq0k3aS0_1(.din(n15388), .dout(n15385));
    jdff dff_A_rLdU8sJG5_1(.din(n15391), .dout(n15388));
    jdff dff_A_GsibDraX6_1(.din(n15394), .dout(n15391));
    jdff dff_A_QlKpmL7l1_1(.din(n15397), .dout(n15394));
    jdff dff_A_idxDFid54_1(.din(n15400), .dout(n15397));
    jdff dff_A_pFynIBHc3_1(.din(n15403), .dout(n15400));
    jdff dff_A_KylSvzqG0_1(.din(n15406), .dout(n15403));
    jdff dff_A_JRn941Bw9_1(.din(n15409), .dout(n15406));
    jdff dff_A_hnYhUgvT6_1(.din(n15412), .dout(n15409));
    jdff dff_A_bKtJ0jLs3_1(.din(n15415), .dout(n15412));
    jdff dff_A_Lf6bnXpT7_1(.din(n15418), .dout(n15415));
    jdff dff_A_EsfkNbea7_1(.din(n15421), .dout(n15418));
    jdff dff_A_eRFKiswX8_1(.din(n15424), .dout(n15421));
    jdff dff_A_sHTJBg2x2_1(.din(n15427), .dout(n15424));
    jdff dff_A_zBdsHkwr0_1(.din(n15430), .dout(n15427));
    jdff dff_A_24gcnJs55_1(.din(n15433), .dout(n15430));
    jdff dff_A_2yoa0Xmg3_1(.din(n15436), .dout(n15433));
    jdff dff_A_I5NxoADI0_1(.din(n15439), .dout(n15436));
    jdff dff_A_dWsgIMZl3_1(.din(n15442), .dout(n15439));
    jdff dff_A_W9XIvgWl1_1(.din(n15445), .dout(n15442));
    jdff dff_A_5avsFQRR6_1(.din(n15448), .dout(n15445));
    jdff dff_A_huoydXMQ2_1(.din(n15451), .dout(n15448));
    jdff dff_A_hYt7MMz02_1(.din(n15454), .dout(n15451));
    jdff dff_A_NlVCp1mj4_1(.din(n15457), .dout(n15454));
    jdff dff_A_O4cQ5JZr6_1(.din(n15460), .dout(n15457));
    jdff dff_A_SKbTFCZj2_1(.din(n15463), .dout(n15460));
    jdff dff_A_1zVdYsML7_1(.din(n682), .dout(n15463));
    jdff dff_A_rGde2L1r5_0(.din(n15469), .dout(n15466));
    jdff dff_A_zj7Wtcb85_0(.din(n541), .dout(n15469));
    jdff dff_B_vxvT3Qbl3_0(.din(G214), .dout(n15473));
    jdff dff_A_ZmpSsmGr0_1(.din(n15478), .dout(n15475));
    jdff dff_A_DY0VH9bL9_1(.din(n558), .dout(n15478));
    jdff dff_A_w1WJmkCq5_2(.din(n15484), .dout(n15481));
    jdff dff_A_4u7xADtA8_2(.din(n558), .dout(n15484));
    jdff dff_A_ob5eTzHp9_2(.din(n15490), .dout(n15487));
    jdff dff_A_3RoiRSzn7_2(.din(n15493), .dout(n15490));
    jdff dff_A_1guXg5S94_2(.din(n15496), .dout(n15493));
    jdff dff_A_lACnqkSy8_2(.din(G1480), .dout(n15496));
    jdff dff_B_ZagUfvbl0_0(.din(G215), .dout(n15500));
    jdff dff_B_wPxDIRJ71_2(.din(n565), .dout(n15503));
    jdff dff_B_8TkpM3NK2_2(.din(n15503), .dout(n15506));
    jdff dff_A_hV1GeVxG4_0(.din(n15511), .dout(n15508));
    jdff dff_A_B1dGCImi7_0(.din(n15514), .dout(n15511));
    jdff dff_A_jwPzA63V8_0(.din(n15517), .dout(n15514));
    jdff dff_A_Ooh0LBXd5_0(.din(G106), .dout(n15517));
    jdff dff_B_03bsOFBl3_1(.din(n5047), .dout(n15521));
    jdff dff_B_65zW7JSU8_1(.din(n5051), .dout(n15524));
    jdff dff_B_dDmxprc12_1(.din(n15524), .dout(n15527));
    jdff dff_B_3SWdjrQz8_1(.din(n15527), .dout(n15530));
    jdff dff_B_lEXq7Dmk5_1(.din(n15530), .dout(n15533));
    jdff dff_B_q2YQNKPl0_1(.din(n15533), .dout(n15536));
    jdff dff_B_84g7pzSx1_1(.din(n15536), .dout(n15539));
    jdff dff_B_UsAZKtNS6_1(.din(n15539), .dout(n15542));
    jdff dff_B_7H7EWBKK6_1(.din(n15542), .dout(n15545));
    jdff dff_B_C6KzTMwc7_1(.din(n15545), .dout(n15548));
    jdff dff_B_r0ROCC9s4_1(.din(n15548), .dout(n15551));
    jdff dff_B_IjIqbyHH4_1(.din(n15551), .dout(n15554));
    jdff dff_B_flmF78nX9_1(.din(n15554), .dout(n15557));
    jdff dff_B_aofrh8mi9_1(.din(n15557), .dout(n15560));
    jdff dff_B_c6sAlVSH7_1(.din(n15560), .dout(n15563));
    jdff dff_B_sqaBfIcu0_0(.din(n5142), .dout(n15566));
    jdff dff_B_Ao6mYGi31_0(.din(n15566), .dout(n15569));
    jdff dff_B_UuW7iBjA1_0(.din(n15569), .dout(n15572));
    jdff dff_B_zXwjkqDF0_0(.din(n15572), .dout(n15575));
    jdff dff_B_WYToY6Qz7_0(.din(n5138), .dout(n15578));
    jdff dff_B_iiTVZbst1_0(.din(n15578), .dout(n15581));
    jdff dff_B_dWg3EtNZ9_0(.din(n5126), .dout(n15584));
    jdff dff_B_2ddakiyz8_0(.din(n15584), .dout(n15587));
    jdff dff_B_23s7cY9T8_0(.din(n15587), .dout(n15590));
    jdff dff_B_v0dM5hOn8_0(.din(n5111), .dout(n15593));
    jdff dff_B_qgka1V8r4_0(.din(n15593), .dout(n15596));
    jdff dff_B_cVuH9BZP5_1(.din(n5081), .dout(n15599));
    jdff dff_B_USdYKckw6_1(.din(n15599), .dout(n15602));
    jdff dff_B_uWWG181A2_0(.din(n5091), .dout(n15605));
    jdff dff_B_rnq9dnf40_0(.din(n15605), .dout(n15608));
    jdff dff_B_aqxciPkK8_0(.din(n15608), .dout(n15611));
    jdff dff_B_zcygb30n6_0(.din(n15611), .dout(n15614));
    jdff dff_B_jjk4JYtM5_0(.din(n15614), .dout(n15617));
    jdff dff_B_mORKMFCh6_0(.din(n15617), .dout(n15620));
    jdff dff_B_zwd4YUXK8_0(.din(n15620), .dout(n15623));
    jdff dff_A_PAVCvIjB5_0(.din(n15628), .dout(n15625));
    jdff dff_A_OgBIZFUB7_0(.din(n15631), .dout(n15628));
    jdff dff_A_mN0ce6hD7_0(.din(n15634), .dout(n15631));
    jdff dff_A_jWx3Jy360_0(.din(n15637), .dout(n15634));
    jdff dff_A_sNwyBztz9_0(.din(n15640), .dout(n15637));
    jdff dff_A_mwdLIJc12_0(.din(n15643), .dout(n15640));
    jdff dff_A_uzD2hOmg0_0(.din(n5088), .dout(n15643));
    jdff dff_A_CNVqdke96_1(.din(n15649), .dout(n15646));
    jdff dff_A_XjAjlG513_1(.din(n15652), .dout(n15649));
    jdff dff_A_whqrPRhn5_1(.din(n15655), .dout(n15652));
    jdff dff_A_hZU2Twyh5_1(.din(n15658), .dout(n15655));
    jdff dff_A_4UNpTZPn2_1(.din(n15661), .dout(n15658));
    jdff dff_A_bqsqtYaC7_1(.din(n15664), .dout(n15661));
    jdff dff_A_BGKrLFec7_1(.din(n5088), .dout(n15664));
    jdff dff_B_uLmvtIRD8_0(.din(n5077), .dout(n15668));
    jdff dff_B_Rvwz1Ntt5_0(.din(n15668), .dout(n15671));
    jdff dff_B_I4GYQyWz0_0(.din(n15671), .dout(n15674));
    jdff dff_B_FFuF2WM68_0(.din(n5069), .dout(n15677));
    jdff dff_A_eZkA2yIW6_1(.din(n15682), .dout(n15679));
    jdff dff_A_IjDgqFsP6_1(.din(n15685), .dout(n15682));
    jdff dff_A_05DUFI563_1(.din(n15688), .dout(n15685));
    jdff dff_A_WPxaR21L2_1(.din(n15691), .dout(n15688));
    jdff dff_A_K8H2s6xj3_1(.din(n15694), .dout(n15691));
    jdff dff_A_MWmQHqrw8_1(.din(n15697), .dout(n15694));
    jdff dff_A_H227V6P77_1(.din(n4500), .dout(n15697));
    jdff dff_B_qwYIpRNY4_1(.din(n4482), .dout(n15701));
    jdff dff_B_oUKrvhW93_1(.din(n15701), .dout(n15704));
    jdff dff_B_yJorNVda5_1(.din(n15704), .dout(n15707));
    jdff dff_B_mp19wXpG4_1(.din(n15707), .dout(n15710));
    jdff dff_B_j7ri32Ll5_1(.din(n15710), .dout(n15713));
    jdff dff_B_rqgIY5ES8_1(.din(n15713), .dout(n15716));
    jdff dff_B_EKprS7Q16_0(.din(n4488), .dout(n15719));
    jdff dff_B_bGDSMlsM5_0(.din(n15719), .dout(n15722));
    jdff dff_B_CnVb1Lwf1_0(.din(n15722), .dout(n15725));
    jdff dff_A_TabvV23X2_1(.din(n15730), .dout(n15727));
    jdff dff_A_vswOw34m7_1(.din(n15733), .dout(n15730));
    jdff dff_A_M1TycP0p7_1(.din(n15736), .dout(n15733));
    jdff dff_A_dfIKLkOG9_1(.din(n15739), .dout(n15736));
    jdff dff_A_DdevqCW49_1(.din(n15742), .dout(n15739));
    jdff dff_A_MLEKQuC59_1(.din(n15745), .dout(n15742));
    jdff dff_A_ngUTuCte4_1(.din(n15748), .dout(n15745));
    jdff dff_A_x3DqQd8p4_1(.din(n15751), .dout(n15748));
    jdff dff_A_Sg5V6eJQ8_1(.din(n15754), .dout(n15751));
    jdff dff_A_o9f56Jhc7_1(.din(n15757), .dout(n15754));
    jdff dff_A_39Do16BY4_1(.din(n15760), .dout(n15757));
    jdff dff_A_ahBHxoSc6_1(.din(n15763), .dout(n15760));
    jdff dff_A_n6i6XZTi2_1(.din(n15766), .dout(n15763));
    jdff dff_A_oWXDgH8R3_1(.din(n15769), .dout(n15766));
    jdff dff_A_07VbPBFq4_1(.din(n4479), .dout(n15769));
    jdff dff_B_1eGYARXL9_0(.din(n5039), .dout(n15773));
    jdff dff_B_JC4Q6jwA2_0(.din(n5035), .dout(n15776));
    jdff dff_B_wwtBx1AL7_1(.din(n4132), .dout(n15779));
    jdff dff_B_Zd7shYUE7_1(.din(n15779), .dout(n15782));
    jdff dff_B_4RDfK5419_1(.din(n15782), .dout(n15785));
    jdff dff_B_cpxQha6Z2_1(.din(n15785), .dout(n15788));
    jdff dff_B_kyDp6uk88_1(.din(n15788), .dout(n15791));
    jdff dff_B_oJVVuy8x8_1(.din(n15791), .dout(n15794));
    jdff dff_B_SEwrgOtF6_1(.din(n15794), .dout(n15797));
    jdff dff_B_NudPdGMP0_1(.din(n15797), .dout(n15800));
    jdff dff_B_tVNopkYn6_1(.din(n15800), .dout(n15803));
    jdff dff_B_eDtWO0qj3_1(.din(n15803), .dout(n15806));
    jdff dff_B_hMF0gLGw1_1(.din(n15806), .dout(n15809));
    jdff dff_B_R7AEYJd50_1(.din(n15809), .dout(n15812));
    jdff dff_B_eZ81QOBf4_0(.din(n5023), .dout(n15815));
    jdff dff_A_3BncMQJW6_1(.din(n15824), .dout(n15817));
    jdff dff_B_4FNzd9Pc5_2(.din(n5015), .dout(n15821));
    jdff dff_B_24mtxUlb8_2(.din(n15821), .dout(n15824));
    jdff dff_B_kBZpwD7o1_0(.din(n5011), .dout(n15827));
    jdff dff_B_hm3K74fN6_0(.din(n15827), .dout(n15830));
    jdff dff_B_XEqBx23A8_0(.din(n15830), .dout(n15833));
    jdff dff_B_4xMheUue8_0(.din(n15833), .dout(n15836));
    jdff dff_B_FkQP94Gv6_0(.din(n5007), .dout(n15839));
    jdff dff_B_CO0nfNWu6_1(.din(n4995), .dout(n15842));
    jdff dff_B_QDA88Cd25_1(.din(n15842), .dout(n15845));
    jdff dff_B_EU2ykJhL3_1(.din(n15845), .dout(n15848));
    jdff dff_A_h2VvtMUM2_0(.din(n15853), .dout(n15850));
    jdff dff_A_WMngvtCD5_0(.din(n15856), .dout(n15853));
    jdff dff_A_mRLmi6Zn1_0(.din(n15859), .dout(n15856));
    jdff dff_A_W85UgazU7_0(.din(n4988), .dout(n15859));
    jdff dff_A_9CJyk6me6_1(.din(n15865), .dout(n15862));
    jdff dff_A_JfAr3Uyd2_1(.din(n15868), .dout(n15865));
    jdff dff_A_aTcH09wp5_1(.din(n15871), .dout(n15868));
    jdff dff_A_pHS2QGSq2_1(.din(n15874), .dout(n15871));
    jdff dff_A_ipZqOBiQ8_1(.din(n15877), .dout(n15874));
    jdff dff_A_oTx87bls5_1(.din(n15880), .dout(n15877));
    jdff dff_A_iqqYYH0K0_1(.din(n15883), .dout(n15880));
    jdff dff_A_vygkvrDe7_1(.din(n15886), .dout(n15883));
    jdff dff_A_bRsDcaSe0_1(.din(n15889), .dout(n15886));
    jdff dff_A_TF5cqGEb7_1(.din(n15892), .dout(n15889));
    jdff dff_A_8IWkgJBx5_1(.din(n15895), .dout(n15892));
    jdff dff_A_LoRLtfpl3_1(.din(n15898), .dout(n15895));
    jdff dff_A_UEjyKK6E7_1(.din(n15901), .dout(n15898));
    jdff dff_A_TR24fotw6_1(.din(n15904), .dout(n15901));
    jdff dff_A_tVeRf5z89_1(.din(n15907), .dout(n15904));
    jdff dff_A_mdctKRx36_1(.din(n4571), .dout(n15907));
    jdff dff_B_uMxn8nPI8_0(.din(n4976), .dout(n15911));
    jdff dff_B_0VGiGqZB7_0(.din(n15911), .dout(n15914));
    jdff dff_B_M3G9IcnN5_0(.din(n15914), .dout(n15917));
    jdff dff_B_mrMzToCv7_0(.din(n15917), .dout(n15920));
    jdff dff_B_bLVqyfKW6_0(.din(n4972), .dout(n15923));
    jdff dff_B_d6WT5pj18_0(.din(n15923), .dout(n15926));
    jdff dff_B_qoeLEU5k2_0(.din(n15926), .dout(n15929));
    jdff dff_A_qdiTRg3f2_1(.din(n15934), .dout(n15931));
    jdff dff_A_PVUmlWos8_1(.din(n15937), .dout(n15934));
    jdff dff_A_reUXqUeJ4_1(.din(n15940), .dout(n15937));
    jdff dff_A_5EqcL14M4_1(.din(n15943), .dout(n15940));
    jdff dff_A_HQovdrkH7_1(.din(n15946), .dout(n15943));
    jdff dff_A_5tmnPJWJ9_1(.din(n15949), .dout(n15946));
    jdff dff_A_cZzw0s9p4_1(.din(n15952), .dout(n15949));
    jdff dff_A_VqPGuDRg5_1(.din(n15955), .dout(n15952));
    jdff dff_A_mnaXM1OV5_1(.din(n15958), .dout(n15955));
    jdff dff_A_XV4JvTtJ0_1(.din(n15961), .dout(n15958));
    jdff dff_A_WknRXqOa9_1(.din(n15964), .dout(n15961));
    jdff dff_A_X0XqqPhE6_1(.din(n15967), .dout(n15964));
    jdff dff_A_EdZdUDdb8_1(.din(n15970), .dout(n15967));
    jdff dff_A_NXxsCLP79_1(.din(n15973), .dout(n15970));
    jdff dff_A_Clg8QBrH5_1(.din(n15976), .dout(n15973));
    jdff dff_A_JRCBIb8S9_1(.din(n15979), .dout(n15976));
    jdff dff_A_ML0wQCZb4_1(.din(n15982), .dout(n15979));
    jdff dff_A_9g0Gj25A9_1(.din(n15985), .dout(n15982));
    jdff dff_A_WmUiygcc7_1(.din(n15988), .dout(n15985));
    jdff dff_A_NRvr2xNV3_1(.din(n15992), .dout(n15988));
    jdff dff_B_XkcTUA521_2(.din(n4543), .dout(n15992));
    jdff dff_A_FmgsxsHO6_2(.din(n1017), .dout(n15994));
    jdff dff_B_Wb2jObOc6_1(.din(n1009), .dout(n15998));
    jdff dff_B_K91H5ioU1_0(.din(G66), .dout(n16001));
    jdff dff_A_pdW84Udt4_0(.din(n16006), .dout(n16003));
    jdff dff_A_KG5akhGz9_0(.din(n1005), .dout(n16006));
    jdff dff_A_CtKtQLz32_2(.din(n16012), .dout(n16009));
    jdff dff_A_qIxN32vE1_2(.din(n1005), .dout(n16012));
    jdff dff_A_9VwgKFyQ5_1(.din(n16018), .dout(n16015));
    jdff dff_A_Rph632JF4_1(.din(n16021), .dout(n16018));
    jdff dff_A_ruSKVlVn2_1(.din(n16024), .dout(n16021));
    jdff dff_A_bdb0wrOh4_1(.din(G4437), .dout(n16024));
    jdff dff_A_cUYEEm9U4_1(.din(n16030), .dout(n16027));
    jdff dff_A_Y9db0dxp5_1(.din(n16033), .dout(n16030));
    jdff dff_A_cAcLb03K7_1(.din(n16036), .dout(n16033));
    jdff dff_A_VKnKUEpK1_1(.din(n16039), .dout(n16036));
    jdff dff_A_MH9i3ecq1_1(.din(n16042), .dout(n16039));
    jdff dff_A_CFcnAxKv8_1(.din(n16045), .dout(n16042));
    jdff dff_A_3dSPtnlF5_1(.din(n16048), .dout(n16045));
    jdff dff_A_PlV3Rsls8_1(.din(n16051), .dout(n16048));
    jdff dff_A_rWD19SEB3_1(.din(n16054), .dout(n16051));
    jdff dff_A_0q8P4K7e5_1(.din(n16057), .dout(n16054));
    jdff dff_A_jlJRbxIg0_1(.din(n16060), .dout(n16057));
    jdff dff_A_VPXYOjKq6_1(.din(n16063), .dout(n16060));
    jdff dff_A_sLEVuBb67_1(.din(n16066), .dout(n16063));
    jdff dff_A_PzXjsi4a4_1(.din(n16069), .dout(n16066));
    jdff dff_A_KfWFhUva8_1(.din(n16072), .dout(n16069));
    jdff dff_A_sEhCQmEg5_1(.din(n4123), .dout(n16072));
    jdff dff_A_gcnzPzKn1_0(.din(n1098), .dout(n16075));
    jdff dff_A_gxjgvuVr0_1(.din(n16081), .dout(n16078));
    jdff dff_A_P1G8j8sL8_1(.din(n16084), .dout(n16081));
    jdff dff_A_OmPDAgAM1_1(.din(n16087), .dout(n16084));
    jdff dff_A_woM42a805_1(.din(n16090), .dout(n16087));
    jdff dff_A_Mz2LidRZ3_1(.din(n16093), .dout(n16090));
    jdff dff_A_QtMsrQbs7_1(.din(n16096), .dout(n16093));
    jdff dff_A_qGmwrrV43_1(.din(n16099), .dout(n16096));
    jdff dff_A_u2yqOSGB8_1(.din(n16102), .dout(n16099));
    jdff dff_A_FuSfG6mH8_1(.din(n16105), .dout(n16102));
    jdff dff_A_uEB1B4xG0_1(.din(n16108), .dout(n16105));
    jdff dff_A_qi908Ma83_1(.din(n16111), .dout(n16108));
    jdff dff_A_A9YZY4lC3_1(.din(n16114), .dout(n16111));
    jdff dff_A_vKpHolfe5_1(.din(n16117), .dout(n16114));
    jdff dff_A_ilokYAdb2_1(.din(n16120), .dout(n16117));
    jdff dff_A_xxYf9NAS1_1(.din(n1098), .dout(n16120));
    jdff dff_B_X5UPQFDB0_0(.din(n4956), .dout(n16124));
    jdff dff_A_NbdGURKy2_0(.din(n16129), .dout(n16126));
    jdff dff_A_Sv7nSz9l8_0(.din(n1705), .dout(n16129));
    jdff dff_A_FFXW9yYQ2_0(.din(n16135), .dout(n16132));
    jdff dff_A_tFkBshhu5_0(.din(n16138), .dout(n16135));
    jdff dff_A_SPOO0Qee5_0(.din(n16141), .dout(n16138));
    jdff dff_A_dLaasbX10_0(.din(n16144), .dout(n16141));
    jdff dff_A_ACfXfwOd5_0(.din(n16147), .dout(n16144));
    jdff dff_A_OKGU5iSW0_0(.din(n16150), .dout(n16147));
    jdff dff_A_HWnCfUvs6_0(.din(n16153), .dout(n16150));
    jdff dff_A_qa8Kysc94_0(.din(n16156), .dout(n16153));
    jdff dff_A_WSlPrr977_0(.din(n16159), .dout(n16156));
    jdff dff_A_AMiEeM2x1_0(.din(n16162), .dout(n16159));
    jdff dff_A_4KU2qdNu9_0(.din(n16165), .dout(n16162));
    jdff dff_A_cP1V2UuK0_0(.din(n16168), .dout(n16165));
    jdff dff_A_EgStRu3Z1_0(.din(n16171), .dout(n16168));
    jdff dff_A_fZaJ32m37_0(.din(n16174), .dout(n16171));
    jdff dff_A_DoHWcUNe7_0(.din(n16177), .dout(n16174));
    jdff dff_A_RF0FdYnX6_0(.din(n1730), .dout(n16177));
    jdff dff_B_0gubTSiJ7_1(.din(n1719), .dout(n16181));
    jdff dff_A_X3wpJNbL7_2(.din(n16186), .dout(n16183));
    jdff dff_A_xa0iUHlC0_2(.din(n16189), .dout(n16186));
    jdff dff_A_F4pBuDFz7_2(.din(n16192), .dout(n16189));
    jdff dff_A_3WTyAe7S4_2(.din(n16195), .dout(n16192));
    jdff dff_A_6C1fHsB43_2(.din(n16198), .dout(n16195));
    jdff dff_A_ndzhgdq44_2(.din(n16201), .dout(n16198));
    jdff dff_A_8oZU5jxL3_2(.din(n16204), .dout(n16201));
    jdff dff_A_YXHTOKGL7_2(.din(n16207), .dout(n16204));
    jdff dff_A_nxsvG44V5_2(.din(n16210), .dout(n16207));
    jdff dff_A_GkxlOikL3_2(.din(n16213), .dout(n16210));
    jdff dff_A_RiUiXrFZ1_2(.din(n16216), .dout(n16213));
    jdff dff_A_n5DF96ap2_2(.din(n16219), .dout(n16216));
    jdff dff_A_egbsKCSp0_2(.din(n16222), .dout(n16219));
    jdff dff_A_bGYEB6pl8_2(.din(n16225), .dout(n16222));
    jdff dff_A_0Z6mcsHj6_2(.din(n16228), .dout(n16225));
    jdff dff_A_tnuH08Or1_2(.din(n16231), .dout(n16228));
    jdff dff_A_rPeFpmjZ9_2(.din(n1091), .dout(n16231));
    jdff dff_A_WpnNlCOD7_0(.din(n16237), .dout(n16234));
    jdff dff_A_lIoSxRE81_0(.din(n16240), .dout(n16237));
    jdff dff_A_V1kp8t771_0(.din(n16243), .dout(n16240));
    jdff dff_A_7QRC78JY0_0(.din(n16246), .dout(n16243));
    jdff dff_A_Lw0NA0X93_0(.din(n16249), .dout(n16246));
    jdff dff_A_UZoUoleR8_0(.din(n16252), .dout(n16249));
    jdff dff_A_E761DXP95_0(.din(n16255), .dout(n16252));
    jdff dff_A_QaSYnA678_0(.din(n16258), .dout(n16255));
    jdff dff_A_eUgnv7qh7_0(.din(n16261), .dout(n16258));
    jdff dff_A_m9MJl1UE7_0(.din(n16264), .dout(n16261));
    jdff dff_A_5U7xi0fk0_0(.din(n16267), .dout(n16264));
    jdff dff_A_PzPvBfxc1_0(.din(n16270), .dout(n16267));
    jdff dff_A_VU7ydF1Q8_0(.din(n16273), .dout(n16270));
    jdff dff_A_eUTDHlIA4_0(.din(n16276), .dout(n16273));
    jdff dff_A_txV26H1W3_0(.din(n16279), .dout(n16276));
    jdff dff_A_zSSjrwjo9_0(.din(n16282), .dout(n16279));
    jdff dff_A_6BYmRLtj1_0(.din(n16285), .dout(n16282));
    jdff dff_A_lCny2K5N7_0(.din(n1069), .dout(n16285));
    jdff dff_B_1BBgLLMX6_1(.din(n1057), .dout(n16289));
    jdff dff_B_ZDKRkgen7_0(.din(G35), .dout(n16292));
    jdff dff_B_DR692JWO3_2(.din(n1053), .dout(n16295));
    jdff dff_B_o50higMX4_2(.din(n16295), .dout(n16298));
    jdff dff_A_GhDTW6uW7_0(.din(n16303), .dout(n16300));
    jdff dff_A_yfxtB0Mj6_0(.din(n16306), .dout(n16303));
    jdff dff_A_5gr2MZxc3_0(.din(n16309), .dout(n16306));
    jdff dff_A_QOT75w8e3_0(.din(G4420), .dout(n16309));
    jdff dff_B_hfhO92eX9_1(.din(n1079), .dout(n16313));
    jdff dff_B_Tf4sktAQ5_0(.din(G32), .dout(n16316));
    jdff dff_B_RoOexd8W5_2(.din(n1075), .dout(n16319));
    jdff dff_B_s3BtrIMB0_2(.din(n16319), .dout(n16322));
    jdff dff_A_9ccwibTO2_1(.din(n16328), .dout(n16324));
    jdff dff_B_xsOrJPyQ6_2(.din(n1715), .dout(n16328));
    jdff dff_A_OJnxlWYq1_2(.din(n16333), .dout(n16330));
    jdff dff_A_qSmO3sxM0_2(.din(n16336), .dout(n16333));
    jdff dff_A_9LQtxqQs0_2(.din(n16339), .dout(n16336));
    jdff dff_A_cyokqCZy9_2(.din(n16342), .dout(n16339));
    jdff dff_A_VgXoLfYa4_2(.din(n1050), .dout(n16342));
    jdff dff_B_S7QK8PnQ1_1(.din(n1038), .dout(n16346));
    jdff dff_B_GlAauAlX5_0(.din(G50), .dout(n16349));
    jdff dff_A_4t9OGUoO9_1(.din(n16354), .dout(n16351));
    jdff dff_A_ze2TbJmO2_1(.din(n1034), .dout(n16354));
    jdff dff_A_McacbpMI7_2(.din(n16360), .dout(n16357));
    jdff dff_A_DSMLlou83_2(.din(n1034), .dout(n16360));
    jdff dff_A_lhwAhZoi6_1(.din(n16366), .dout(n16363));
    jdff dff_A_QUdhUQBY9_1(.din(n16369), .dout(n16366));
    jdff dff_A_AzityleY0_1(.din(n16372), .dout(n16369));
    jdff dff_A_ttAswpf56_1(.din(G4432), .dout(n16372));
    jdff dff_A_TLQRb0oS4_1(.din(n16378), .dout(n16375));
    jdff dff_A_fojp8nj44_1(.din(n16381), .dout(n16378));
    jdff dff_A_TiY8jbIF4_1(.din(n16384), .dout(n16381));
    jdff dff_A_Uy6kw2GG4_1(.din(n4126), .dout(n16384));
    jdff dff_A_QAA4dzyl1_1(.din(n16390), .dout(n16387));
    jdff dff_A_icwwhiNp2_1(.din(n16393), .dout(n16390));
    jdff dff_A_BzJeaHSw9_1(.din(n16396), .dout(n16393));
    jdff dff_A_O2xbLzO42_1(.din(n16399), .dout(n16396));
    jdff dff_A_qmdxOz5k3_1(.din(n1268), .dout(n16399));
    jdff dff_B_a6OhZh6Y1_1(.din(n1120), .dout(n16403));
    jdff dff_B_f82gaWqz6_1(.din(n16403), .dout(n16406));
    jdff dff_B_tH0iE8Zk9_1(.din(n16406), .dout(n16409));
    jdff dff_B_1xEumEkB4_1(.din(n16409), .dout(n16412));
    jdff dff_B_qjwCuMP90_1(.din(n16412), .dout(n16415));
    jdff dff_B_0H8kGMJe9_1(.din(n16415), .dout(n16418));
    jdff dff_B_0osHwrEi3_1(.din(n16418), .dout(n16421));
    jdff dff_B_zL3CkYRw0_1(.din(n16421), .dout(n16424));
    jdff dff_B_w5dep8MM1_1(.din(n16424), .dout(n16427));
    jdff dff_B_14DQgkg33_1(.din(n1130), .dout(n16430));
    jdff dff_B_iS5JGtt31_1(.din(n16430), .dout(n16433));
    jdff dff_B_1LTYs2VH4_1(.din(n16433), .dout(n16436));
    jdff dff_B_CXbr2tSP6_1(.din(n16436), .dout(n16439));
    jdff dff_B_6gyHgv593_1(.din(n16439), .dout(n16442));
    jdff dff_B_o9pz9yqM5_1(.din(n16442), .dout(n16445));
    jdff dff_A_7qvt01Gw7_1(.din(n16450), .dout(n16447));
    jdff dff_A_EeAwhK9t6_1(.din(n16453), .dout(n16450));
    jdff dff_A_jVlUQMio7_1(.din(n16456), .dout(n16453));
    jdff dff_A_HybwZxUB0_1(.din(n16459), .dout(n16456));
    jdff dff_A_45QPxJd27_1(.din(n16462), .dout(n16459));
    jdff dff_A_9zizjlgD3_1(.din(n16465), .dout(n16462));
    jdff dff_A_a2DMK6Mh4_1(.din(n1260), .dout(n16465));
    jdff dff_B_yiMi5WIJ2_1(.din(n1149), .dout(n16469));
    jdff dff_B_RPzbXaBE0_1(.din(n16469), .dout(n16472));
    jdff dff_B_oicmsVBS8_1(.din(n16472), .dout(n16475));
    jdff dff_B_EEYomzKA0_1(.din(n16475), .dout(n16478));
    jdff dff_B_Z9Yjz69g1_1(.din(n16478), .dout(n16481));
    jdff dff_B_nPL5O5D18_1(.din(n16481), .dout(n16484));
    jdff dff_B_aKKKoBAO2_1(.din(n16484), .dout(n16487));
    jdff dff_B_Me8b3bQA0_1(.din(n1159), .dout(n16490));
    jdff dff_B_zoefxJOB6_1(.din(n16490), .dout(n16493));
    jdff dff_B_oRD1y27v5_1(.din(n16493), .dout(n16496));
    jdff dff_B_Hit352gK4_1(.din(n16496), .dout(n16499));
    jdff dff_B_LBb1e79w3_1(.din(n1188), .dout(n16502));
    jdff dff_B_Md0cH27z3_1(.din(n16502), .dout(n16505));
    jdff dff_A_j7Vpwvjf1_0(.din(n16510), .dout(n16507));
    jdff dff_A_nMqu4bjN2_0(.din(n16513), .dout(n16510));
    jdff dff_A_cU02PYpS4_0(.din(n16516), .dout(n16513));
    jdff dff_A_RgqDsN3a3_0(.din(n16519), .dout(n16516));
    jdff dff_A_6Lo7wcKL3_0(.din(n16522), .dout(n16519));
    jdff dff_A_2ImJFL3k4_0(.din(n16525), .dout(n16522));
    jdff dff_A_BrNc2Zwt0_0(.din(n16528), .dout(n16525));
    jdff dff_A_ZB5F9ZHS6_0(.din(n16531), .dout(n16528));
    jdff dff_A_wY4cOqzB6_0(.din(n16534), .dout(n16531));
    jdff dff_A_ujQXfP9L6_0(.din(n16537), .dout(n16534));
    jdff dff_A_TRgHmW7P3_0(.din(n1244), .dout(n16537));
    jdff dff_A_h6jXJq6t3_1(.din(n16543), .dout(n16540));
    jdff dff_A_MhbFbLx72_1(.din(n16546), .dout(n16543));
    jdff dff_A_KdPodqNV8_1(.din(n16549), .dout(n16546));
    jdff dff_A_a4AEExw83_1(.din(n16552), .dout(n16549));
    jdff dff_A_fuN38Th80_1(.din(n16555), .dout(n16552));
    jdff dff_A_XYunfvvK4_1(.din(n16558), .dout(n16555));
    jdff dff_A_CIq3GO9s4_1(.din(n16561), .dout(n16558));
    jdff dff_A_4NkmOesI3_1(.din(n16564), .dout(n16561));
    jdff dff_A_gxjmdQNJ1_1(.din(n16567), .dout(n16564));
    jdff dff_A_BfOUIvdr8_1(.din(n16570), .dout(n16567));
    jdff dff_A_nbD5zfLn8_1(.din(n16573), .dout(n16570));
    jdff dff_A_Nx1p4Kpj3_1(.din(n16576), .dout(n16573));
    jdff dff_A_DfWVp4ef4_1(.din(n16579), .dout(n16576));
    jdff dff_A_MGkzqXCE2_1(.din(n16582), .dout(n16579));
    jdff dff_A_hFM6fXmV7_1(.din(n1236), .dout(n16582));
    jdff dff_A_kkEaQzo72_2(.din(n16588), .dout(n16585));
    jdff dff_A_md8RtMPF9_2(.din(n1236), .dout(n16588));
    jdff dff_A_9H7CSzP19_0(.din(n1214), .dout(n16591));
    jdff dff_A_oQuHNRS80_1(.din(n1207), .dout(n16594));
    jdff dff_A_R95kl5eb2_2(.din(n16600), .dout(n16597));
    jdff dff_A_gKKIKIjz5_2(.din(n16603), .dout(n16600));
    jdff dff_A_dGv0HnBV7_2(.din(n1207), .dout(n16603));
    jdff dff_A_xtbKG4df1_0(.din(n16609), .dout(n16606));
    jdff dff_A_itcAS2LG7_0(.din(n16612), .dout(n16609));
    jdff dff_A_VWIuIhjw6_0(.din(n16615), .dout(n16612));
    jdff dff_A_u9hrOZe56_0(.din(n16618), .dout(n16615));
    jdff dff_A_HAQrLaVw1_0(.din(n1185), .dout(n16618));
    jdff dff_A_E4QIsxER2_1(.din(n16624), .dout(n16621));
    jdff dff_A_QisLD6h50_1(.din(n16627), .dout(n16624));
    jdff dff_A_GngKVSlr5_1(.din(n16630), .dout(n16627));
    jdff dff_A_yLqtJmZL3_1(.din(n16633), .dout(n16630));
    jdff dff_A_3WoZ6Qs11_1(.din(n1178), .dout(n16633));
    jdff dff_A_aMyWZKbS1_1(.din(n16639), .dout(n16636));
    jdff dff_A_oKs18H4K4_1(.din(n16664), .dout(n16639));
    jdff dff_B_iS4GFBys8_2(.din(n4129), .dout(n16643));
    jdff dff_B_OC3cbWcf6_2(.din(n16643), .dout(n16646));
    jdff dff_B_hsmlqB6f6_2(.din(n16646), .dout(n16649));
    jdff dff_B_7CLyjbwD3_2(.din(n16649), .dout(n16652));
    jdff dff_B_6GTJuSD64_2(.din(n16652), .dout(n16655));
    jdff dff_B_qZe0Y4ZI8_2(.din(n16655), .dout(n16658));
    jdff dff_B_yU4cyUmK7_2(.din(n16658), .dout(n16661));
    jdff dff_B_jm3SBMPv0_2(.din(n16661), .dout(n16664));
    jdff dff_A_V9Yu8TzO9_0(.din(n16669), .dout(n16666));
    jdff dff_A_QQEgXUCX7_0(.din(n16672), .dout(n16669));
    jdff dff_A_Ydu3eo0F2_0(.din(n16675), .dout(n16672));
    jdff dff_A_nVS25w047_0(.din(n16678), .dout(n16675));
    jdff dff_A_XWCBOf1L4_0(.din(n16681), .dout(n16678));
    jdff dff_A_13P1wu2X7_0(.din(n16684), .dout(n16681));
    jdff dff_A_ljIFcQ6O6_0(.din(n1304), .dout(n16684));
    jdff dff_A_fcEi5dX74_2(.din(n16690), .dout(n16687));
    jdff dff_A_pFRmMylo5_2(.din(n16693), .dout(n16690));
    jdff dff_A_Y0RvLGZH2_2(.din(n16696), .dout(n16693));
    jdff dff_A_addw5Elf2_2(.din(n16699), .dout(n16696));
    jdff dff_A_aOM5wPos3_2(.din(n16702), .dout(n16699));
    jdff dff_A_a0xwW19R2_2(.din(n16705), .dout(n16702));
    jdff dff_A_m7BPBVeD9_2(.din(n16708), .dout(n16705));
    jdff dff_A_pglbKG1h6_2(.din(n16711), .dout(n16708));
    jdff dff_A_PQfki17f3_2(.din(n16714), .dout(n16711));
    jdff dff_A_BbqT1xbR5_2(.din(n16717), .dout(n16714));
    jdff dff_A_2EevMicO9_2(.din(n1304), .dout(n16717));
    jdff dff_A_j45oVpwh7_0(.din(n16723), .dout(n16720));
    jdff dff_A_jiux9eNi8_0(.din(n16726), .dout(n16723));
    jdff dff_A_bplawuSj0_0(.din(n16729), .dout(n16726));
    jdff dff_A_y4JmTDcA8_0(.din(n16732), .dout(n16729));
    jdff dff_A_WfVSZ6Rn1_0(.din(n16735), .dout(n16732));
    jdff dff_A_amHkDlX56_0(.din(n16738), .dout(n16735));
    jdff dff_A_IYP4Qtpr2_0(.din(n1300), .dout(n16738));
    jdff dff_A_f47I2eI74_1(.din(n16744), .dout(n16741));
    jdff dff_A_9iXGh8Hf9_1(.din(n16747), .dout(n16744));
    jdff dff_A_rXPU0POp2_1(.din(n16750), .dout(n16747));
    jdff dff_A_YSOuSMyB4_1(.din(n16753), .dout(n16750));
    jdff dff_A_HwNhSJvh4_1(.din(n16756), .dout(n16753));
    jdff dff_A_eYogqwxd6_1(.din(n16759), .dout(n16756));
    jdff dff_A_VANahx7h4_1(.din(n16762), .dout(n16759));
    jdff dff_A_q7M6kJU42_1(.din(n16765), .dout(n16762));
    jdff dff_A_q4eSgDJJ1_1(.din(n16768), .dout(n16765));
    jdff dff_A_vULS35Ya7_1(.din(n16771), .dout(n16768));
    jdff dff_A_vjUkS9AR4_1(.din(n16774), .dout(n16771));
    jdff dff_A_nSimRdzg0_1(.din(n1300), .dout(n16774));
    jdff dff_A_m1xlhcAx1_0(.din(n1292), .dout(n16777));
    jdff dff_A_eWSBL3Rl6_1(.din(n16783), .dout(n16780));
    jdff dff_A_tDpN4mup8_1(.din(n16786), .dout(n16783));
    jdff dff_A_IvD4zRpv4_1(.din(n16789), .dout(n16786));
    jdff dff_A_STxpAMYJ6_1(.din(n16792), .dout(n16789));
    jdff dff_A_Zz1qrTBt0_1(.din(n16795), .dout(n16792));
    jdff dff_A_UPRVCcTd1_1(.din(n16798), .dout(n16795));
    jdff dff_A_GWv2Ifkk4_1(.din(n16801), .dout(n16798));
    jdff dff_A_3n4UuHX64_1(.din(n16804), .dout(n16801));
    jdff dff_A_eXxIkS7S1_1(.din(n16807), .dout(n16804));
    jdff dff_A_rVEXEA3D4_1(.din(n16810), .dout(n16807));
    jdff dff_A_f10blSsZ4_1(.din(n16813), .dout(n16810));
    jdff dff_A_mqsdTUsB8_1(.din(n16816), .dout(n16813));
    jdff dff_A_yJoL8IxM9_1(.din(n16819), .dout(n16816));
    jdff dff_A_pnN4e0tt2_1(.din(n16822), .dout(n16819));
    jdff dff_A_icuiq9cj9_1(.din(n16825), .dout(n16822));
    jdff dff_A_Jy21ZVUD4_1(.din(n1292), .dout(n16825));
    jdff dff_B_lncsuzpc2_1(.din(n1166), .dout(n16829));
    jdff dff_B_NdacBAVQ8_0(.din(G94), .dout(n16832));
    jdff dff_B_MCOGhzGZ9_2(.din(n1162), .dout(n16835));
    jdff dff_B_JLLYtHSi6_2(.din(n16835), .dout(n16838));
    jdff dff_A_jsUAqiQy4_0(.din(n16843), .dout(n16840));
    jdff dff_A_Nwk7wgF06_0(.din(n16846), .dout(n16843));
    jdff dff_A_5POAQ0Lp3_0(.din(n16849), .dout(n16846));
    jdff dff_A_KsBxcwTl2_0(.din(G4405), .dout(n16849));
    jdff dff_B_eBTD6XLU8_1(.din(n1137), .dout(n16853));
    jdff dff_B_VTqLAKE61_0(.din(G121), .dout(n16856));
    jdff dff_A_fD6XjZkR4_1(.din(n16861), .dout(n16858));
    jdff dff_A_hOgeOUPF7_1(.din(n1133), .dout(n16861));
    jdff dff_A_wLnxcjBH0_2(.din(n16867), .dout(n16864));
    jdff dff_A_iC5C8OjB4_2(.din(n1133), .dout(n16867));
    jdff dff_A_DeYJNhYT6_1(.din(n16873), .dout(n16870));
    jdff dff_A_YXAAON592_1(.din(n16876), .dout(n16873));
    jdff dff_A_yT4V3izG7_1(.din(n16879), .dout(n16876));
    jdff dff_A_RQNKq2ED1_1(.din(G4410), .dout(n16879));
    jdff dff_A_H1TkR1ev1_0(.din(n16885), .dout(n16882));
    jdff dff_A_w25X416A8_0(.din(n16888), .dout(n16885));
    jdff dff_A_lUCU7CAt0_0(.din(n16891), .dout(n16888));
    jdff dff_A_VOURb8ns2_0(.din(n16894), .dout(n16891));
    jdff dff_A_Q1cYFrFu1_0(.din(n16897), .dout(n16894));
    jdff dff_A_xwFz6suw3_0(.din(n16900), .dout(n16897));
    jdff dff_A_e9mg32bY4_0(.din(n16903), .dout(n16900));
    jdff dff_A_kGhswp7n5_0(.din(n16906), .dout(n16903));
    jdff dff_A_XH39Dzng4_0(.din(n16909), .dout(n16906));
    jdff dff_A_UhNbnvkD5_0(.din(n16912), .dout(n16909));
    jdff dff_A_F7SLceJQ5_0(.din(n16915), .dout(n16912));
    jdff dff_A_fviSfmSJ5_0(.din(n16918), .dout(n16915));
    jdff dff_A_LqCO2wEt1_0(.din(n1284), .dout(n16918));
    jdff dff_A_L8Jt8ksO4_0(.din(n16924), .dout(n16921));
    jdff dff_A_4y45Qwkg8_0(.din(n16927), .dout(n16924));
    jdff dff_A_yAcqsvcv1_0(.din(n16930), .dout(n16927));
    jdff dff_A_hnsfD6Wa9_0(.din(n16933), .dout(n16930));
    jdff dff_A_Ec1vrAUN4_0(.din(n16936), .dout(n16933));
    jdff dff_A_Q4gWlfxQ5_0(.din(n16939), .dout(n16936));
    jdff dff_A_tc4wjIme4_0(.din(n16942), .dout(n16939));
    jdff dff_A_WKkDVb398_0(.din(n16945), .dout(n16942));
    jdff dff_A_zWBuL2iM5_0(.din(n16948), .dout(n16945));
    jdff dff_A_7nbNurT41_0(.din(n16951), .dout(n16948));
    jdff dff_A_1UPCQan38_0(.din(n16954), .dout(n16951));
    jdff dff_A_Db3vSDXQ2_0(.din(n16957), .dout(n16954));
    jdff dff_A_fgRorDQ94_0(.din(n16960), .dout(n16957));
    jdff dff_A_834GmKxn6_0(.din(n1280), .dout(n16960));
    jdff dff_A_mr411PyE1_2(.din(n16966), .dout(n16963));
    jdff dff_A_diwNUycN8_2(.din(n16969), .dout(n16966));
    jdff dff_A_z8Of0bIP4_2(.din(n16972), .dout(n16969));
    jdff dff_A_cL81nsjY6_2(.din(n16975), .dout(n16972));
    jdff dff_A_i3EjHGms9_2(.din(n16978), .dout(n16975));
    jdff dff_A_65K3OV268_2(.din(n16981), .dout(n16978));
    jdff dff_A_eq2zt1Y13_2(.din(n16984), .dout(n16981));
    jdff dff_A_OtOJedEa0_2(.din(n16987), .dout(n16984));
    jdff dff_A_TBsNULbG4_2(.din(n16990), .dout(n16987));
    jdff dff_A_7AA5fqZw8_2(.din(n16993), .dout(n16990));
    jdff dff_A_AzHJQS0M2_2(.din(n16996), .dout(n16993));
    jdff dff_A_eg8aB7iI1_2(.din(n16999), .dout(n16996));
    jdff dff_A_rGfyodch6_2(.din(n17002), .dout(n16999));
    jdff dff_A_vgM6wKl89_2(.din(n1280), .dout(n17002));
    jdff dff_B_zfeiiKV59_1(.din(n1224), .dout(n17006));
    jdff dff_B_B9vMYkRe1_0(.din(G118), .dout(n17009));
    jdff dff_B_qmQ8RXc35_2(.din(n1220), .dout(n17012));
    jdff dff_B_mbNgPm2M9_2(.din(n17012), .dout(n17015));
    jdff dff_A_fBS8ixlD8_2(.din(n17020), .dout(n17017));
    jdff dff_A_UaorlTs97_2(.din(n17023), .dout(n17020));
    jdff dff_A_WWwU03BM3_2(.din(n17026), .dout(n17023));
    jdff dff_A_E5eUml0l6_2(.din(G4394), .dout(n17026));
    jdff dff_A_YjrnoYQ10_1(.din(n17032), .dout(n17029));
    jdff dff_A_6V5Tyu9B5_1(.din(n17035), .dout(n17032));
    jdff dff_A_IrR3M08e7_1(.din(n17038), .dout(n17035));
    jdff dff_A_CjzTuaok6_1(.din(n17041), .dout(n17038));
    jdff dff_A_Ai8doFeD4_1(.din(n17044), .dout(n17041));
    jdff dff_A_B4W2SeIN8_1(.din(n17047), .dout(n17044));
    jdff dff_A_h7He2goE9_1(.din(n17050), .dout(n17047));
    jdff dff_A_C3wFZKjy1_1(.din(n17053), .dout(n17050));
    jdff dff_A_aoA6KkSh8_1(.din(n17056), .dout(n17053));
    jdff dff_A_lwRixicT2_1(.din(n17059), .dout(n17056));
    jdff dff_A_JcXsaGgX0_1(.din(n17062), .dout(n17059));
    jdff dff_A_kkzKgLQU8_1(.din(n17065), .dout(n17062));
    jdff dff_A_ytGAotxk2_1(.din(n17068), .dout(n17065));
    jdff dff_A_UbRdQzBQ3_1(.din(n17071), .dout(n17068));
    jdff dff_A_FI0vtvFW6_1(.din(n17074), .dout(n17071));
    jdff dff_A_XafuP8tA7_1(.din(n1276), .dout(n17074));
    jdff dff_B_Ay4BhMt72_1(.din(n1195), .dout(n17078));
    jdff dff_B_d32fgfP58_0(.din(G97), .dout(n17081));
    jdff dff_B_XMHt8AVL9_2(.din(n1191), .dout(n17084));
    jdff dff_B_o3YYZP3c6_2(.din(n17084), .dout(n17087));
    jdff dff_A_psUMw5Bv8_0(.din(n17092), .dout(n17089));
    jdff dff_A_ew2MzLwk9_0(.din(n17095), .dout(n17092));
    jdff dff_A_8ek1yGCB3_0(.din(n17098), .dout(n17095));
    jdff dff_A_pTOs2fBc6_0(.din(G4400), .dout(n17098));
    jdff dff_A_6MdOfsxL0_0(.din(n17104), .dout(n17101));
    jdff dff_A_AIIYD2so7_0(.din(n17107), .dout(n17104));
    jdff dff_A_REoYckIc9_0(.din(n17110), .dout(n17107));
    jdff dff_A_KUOvir0x7_0(.din(n17113), .dout(n17110));
    jdff dff_A_d40E8XcC7_0(.din(n17116), .dout(n17113));
    jdff dff_A_ynijqlNQ3_0(.din(n17119), .dout(n17116));
    jdff dff_A_Kpdj06vu8_0(.din(n17122), .dout(n17119));
    jdff dff_A_7xQjhrrT7_0(.din(n17125), .dout(n17122));
    jdff dff_A_INjiewfE2_0(.din(n17128), .dout(n17125));
    jdff dff_A_ejd5kZHd0_0(.din(n17131), .dout(n17128));
    jdff dff_A_6p5yPW499_0(.din(n17134), .dout(n17131));
    jdff dff_A_4AXJbFjP3_0(.din(n17137), .dout(n17134));
    jdff dff_A_gvkPwK1R6_0(.din(n17140), .dout(n17137));
    jdff dff_A_hguD7QRp5_0(.din(n17162), .dout(n17140));
    jdff dff_A_tYjulFFW0_1(.din(n17146), .dout(n17143));
    jdff dff_A_txsL6BBs8_1(.din(n17149), .dout(n17146));
    jdff dff_A_zkIvd3R72_1(.din(n17162), .dout(n17149));
    jdff dff_A_iDFAnv7Y7_2(.din(n17155), .dout(n17152));
    jdff dff_A_Pvhb6ZV98_2(.din(n17162), .dout(n17155));
    jdff dff_B_S8Z1ZWjF1_3(.din(n1272), .dout(n17159));
    jdff dff_B_w0b9mGea6_3(.din(n17159), .dout(n17162));
    jdff dff_B_hpaCQnrD8_1(.din(n1108), .dout(n17165));
    jdff dff_B_zO4tm7vU4_0(.din(G47), .dout(n17168));
    jdff dff_B_TXLOIQC71_2(.din(n1104), .dout(n17171));
    jdff dff_B_6kXN9UvO1_2(.din(n17171), .dout(n17174));
    jdff dff_A_a3ffRSgg9_0(.din(n17179), .dout(n17176));
    jdff dff_A_nM7jgZub7_0(.din(n17182), .dout(n17179));
    jdff dff_A_I120n9PQ1_0(.din(n17185), .dout(n17182));
    jdff dff_A_9AKXfkfi4_0(.din(G4415), .dout(n17185));
    jdff dff_B_aV689boM3_1(.din(n1333), .dout(n17189));
    jdff dff_B_EMrRo1jj1_1(.din(n17189), .dout(n17192));
    jdff dff_B_LFNDJRb97_1(.din(n17192), .dout(n17195));
    jdff dff_B_PaXEQWEA3_1(.din(n17195), .dout(n17198));
    jdff dff_B_yKZFxwnm6_1(.din(n17198), .dout(n17201));
    jdff dff_B_8AhLXQQP6_1(.din(n17201), .dout(n17204));
    jdff dff_B_MdLgWlRM9_1(.din(n17204), .dout(n17207));
    jdff dff_B_xiawR7N49_1(.din(n17207), .dout(n17210));
    jdff dff_B_T6NLPMsr0_1(.din(n17210), .dout(n17213));
    jdff dff_B_VXnoGf3b7_1(.din(n17213), .dout(n17216));
    jdff dff_B_XvmBW3hC8_1(.din(n1449), .dout(n17219));
    jdff dff_B_skb62kuA6_1(.din(n17219), .dout(n17222));
    jdff dff_B_P7LsQFV40_1(.din(n17222), .dout(n17225));
    jdff dff_B_DN46X9li4_1(.din(n17225), .dout(n17228));
    jdff dff_B_W5HpanmD0_1(.din(n1452), .dout(n17231));
    jdff dff_B_FNWAFQOO8_1(.din(n17231), .dout(n17234));
    jdff dff_B_xZN7lzeh2_1(.din(n17234), .dout(n17237));
    jdff dff_B_arJKPxfw8_1(.din(n17237), .dout(n17240));
    jdff dff_A_2ydoM0Lz3_0(.din(n17245), .dout(n17242));
    jdff dff_A_0Q5F53ju8_0(.din(n17248), .dout(n17245));
    jdff dff_A_eGfvfQ5k5_0(.din(n17860), .dout(n17248));
    jdff dff_A_sYy0gg4E5_1(.din(n17254), .dout(n17251));
    jdff dff_A_HTS5qAX63_1(.din(n17257), .dout(n17254));
    jdff dff_A_rWmUNWKg4_1(.din(n17260), .dout(n17257));
    jdff dff_A_1qpZwEpq4_1(.din(n17263), .dout(n17260));
    jdff dff_A_fj54Z1BF9_1(.din(n17266), .dout(n17263));
    jdff dff_A_HL8nOjL58_1(.din(n17269), .dout(n17266));
    jdff dff_A_dzxADrtF4_1(.din(n17860), .dout(n17269));
    jdff dff_A_U4zVM82Y9_0(.din(n17275), .dout(n17272));
    jdff dff_A_n9LvWGKt4_0(.din(n17278), .dout(n17275));
    jdff dff_A_M2ofONVP6_0(.din(n17281), .dout(n17278));
    jdff dff_A_p6MopZZu3_0(.din(n17284), .dout(n17281));
    jdff dff_A_ahdM1dSZ2_0(.din(n17287), .dout(n17284));
    jdff dff_A_Z2ePpNmk0_0(.din(n17290), .dout(n17287));
    jdff dff_A_TutWKrlk6_0(.din(n17293), .dout(n17290));
    jdff dff_A_npGINIGV7_0(.din(n17296), .dout(n17293));
    jdff dff_A_iIlM0pb63_0(.din(n17299), .dout(n17296));
    jdff dff_A_SApXtcds4_0(.din(n17302), .dout(n17299));
    jdff dff_A_I8ZCmTMw6_0(.din(n1330), .dout(n17302));
    jdff dff_A_zL1CMt5T3_1(.din(n17308), .dout(n17305));
    jdff dff_A_zdNmMN4z5_1(.din(n17311), .dout(n17308));
    jdff dff_A_Kutyw1wQ0_1(.din(n17314), .dout(n17311));
    jdff dff_A_cVl90BdP7_1(.din(n17317), .dout(n17314));
    jdff dff_A_tWk0h5Mk6_1(.din(n17320), .dout(n17317));
    jdff dff_A_ONqJEs5t9_1(.din(n17323), .dout(n17320));
    jdff dff_A_2RymdssX3_1(.din(n17326), .dout(n17323));
    jdff dff_A_gnpfGqTm5_1(.din(n17329), .dout(n17326));
    jdff dff_A_JJmyLzV54_1(.din(n17332), .dout(n17329));
    jdff dff_A_7g1m9XmN6_1(.din(n17335), .dout(n17332));
    jdff dff_A_MTC5u9nW3_1(.din(n17338), .dout(n17335));
    jdff dff_A_Kvr04JiN4_1(.din(n17341), .dout(n17338));
    jdff dff_A_UOjkKZjf8_1(.din(n1323), .dout(n17341));
    jdff dff_A_vf1lO32r1_2(.din(n17347), .dout(n17344));
    jdff dff_A_I6NJZyvv3_2(.din(n17350), .dout(n17347));
    jdff dff_A_tpefdaWu0_2(.din(n17353), .dout(n17350));
    jdff dff_A_xg2SzjY73_2(.din(n17356), .dout(n17353));
    jdff dff_A_HtcKTuk79_2(.din(n17359), .dout(n17356));
    jdff dff_A_z767cB1A0_2(.din(n17362), .dout(n17359));
    jdff dff_A_LwSPtd0c8_2(.din(n17365), .dout(n17362));
    jdff dff_A_68v2XJIJ9_2(.din(n17368), .dout(n17365));
    jdff dff_A_uNmMGJuS4_2(.din(n17371), .dout(n17368));
    jdff dff_A_Sm5KmY0V8_2(.din(n17374), .dout(n17371));
    jdff dff_A_zAvLW0qS0_2(.din(n17377), .dout(n17374));
    jdff dff_A_3mdVLWpU8_2(.din(n17380), .dout(n17377));
    jdff dff_A_Jif3DlyP9_2(.din(n1323), .dout(n17380));
    jdff dff_B_sazdHijE6_0(.din(n5356), .dout(n17384));
    jdff dff_B_SrJEm8ST2_0(.din(n17384), .dout(n17387));
    jdff dff_B_Q71OLlIm8_0(.din(n17387), .dout(n17390));
    jdff dff_B_yLAvauhF0_0(.din(n17390), .dout(n17393));
    jdff dff_B_roJCGVcF8_0(.din(n17393), .dout(n17396));
    jdff dff_B_8LVKQobM8_0(.din(n17396), .dout(n17399));
    jdff dff_B_bzKPX9cf4_0(.din(n17399), .dout(n17402));
    jdff dff_B_d1aAI8ly4_0(.din(n17402), .dout(n17405));
    jdff dff_B_Az2yaSxJ4_0(.din(n17405), .dout(n17408));
    jdff dff_B_ozeg8SWK8_0(.din(n17408), .dout(n17411));
    jdff dff_B_dE3sVdpW8_0(.din(n17411), .dout(n17414));
    jdff dff_B_N05BqhbP3_1(.din(n5318), .dout(n17417));
    jdff dff_B_NIqczoov3_1(.din(n17417), .dout(n17420));
    jdff dff_B_qI4S16l17_1(.din(n5321), .dout(n17423));
    jdff dff_A_3xDhesA69_0(.din(n17428), .dout(n17425));
    jdff dff_A_o1ibeUd56_0(.din(n5315), .dout(n17428));
    jdff dff_B_pLSfkFdq2_0(.din(n5303), .dout(n17432));
    jdff dff_B_r2mzG9rG0_0(.din(n17432), .dout(n17435));
    jdff dff_B_6dtNDip40_1(.din(n5280), .dout(n17438));
    jdff dff_B_9hQjcZU16_1(.din(n17438), .dout(n17441));
    jdff dff_B_pGs50NTd7_1(.din(n5268), .dout(n17444));
    jdff dff_B_9fCmHICZ8_0(.din(n5272), .dout(n17447));
    jdff dff_B_2NxGL0PU0_0(.din(n17447), .dout(n17450));
    jdff dff_B_oOQZMAY02_0(.din(n17450), .dout(n17453));
    jdff dff_B_uBDpo2xi1_0(.din(n17453), .dout(n17456));
    jdff dff_B_fEle8DqW2_0(.din(n17456), .dout(n17459));
    jdff dff_A_T9LZAj526_0(.din(n17464), .dout(n17461));
    jdff dff_A_OtQD0IBF3_0(.din(n17467), .dout(n17464));
    jdff dff_A_6NPsbDMG0_0(.din(n5265), .dout(n17467));
    jdff dff_B_5Ifwxcif7_0(.din(n5261), .dout(n17471));
    jdff dff_A_UWlumCSz6_0(.din(n17476), .dout(n17473));
    jdff dff_A_r61HzQDy6_0(.din(n17479), .dout(n17476));
    jdff dff_A_tf5p52Ec4_0(.din(n17482), .dout(n17479));
    jdff dff_A_dPrAgsv13_0(.din(n17485), .dout(n17482));
    jdff dff_A_dOaRQNjy6_0(.din(n5257), .dout(n17485));
    jdff dff_B_NWmQF8Ab9_0(.din(n5249), .dout(n17489));
    jdff dff_B_YtMXNCep7_1(.din(n5190), .dout(n17492));
    jdff dff_A_cU7m0Lw71_1(.din(n17498), .dout(n17494));
    jdff dff_B_w8rOjI4n1_2(.din(n5225), .dout(n17498));
    jdff dff_B_3XopZPmy5_0(.din(n5221), .dout(n17501));
    jdff dff_B_vR2uCBVR6_0(.din(n5217), .dout(n17504));
    jdff dff_B_3KXtXQqc2_0(.din(n17504), .dout(n17507));
    jdff dff_B_ZmV7R1xK6_0(.din(n17507), .dout(n17510));
    jdff dff_B_0XqqsElB1_0(.din(n5205), .dout(n17513));
    jdff dff_A_LuCcrrTp7_1(.din(n17518), .dout(n17515));
    jdff dff_A_YmjYPiIJ5_1(.din(n17521), .dout(n17518));
    jdff dff_A_4RzCVLNv9_1(.din(n17524), .dout(n17521));
    jdff dff_A_RvvrxBSi0_1(.din(n17527), .dout(n17524));
    jdff dff_A_C86U8i2H1_1(.din(n17530), .dout(n17527));
    jdff dff_A_b9c2Mbgn9_1(.din(n17533), .dout(n17530));
    jdff dff_A_r3qnJ5C00_1(.din(n17536), .dout(n17533));
    jdff dff_A_QtZCvjht7_1(.din(n17539), .dout(n17536));
    jdff dff_A_BZUMQKgO2_1(.din(n17542), .dout(n17539));
    jdff dff_A_Da3PXiuw3_1(.din(n3347), .dout(n17542));
    jdff dff_A_GpkEY0jh0_1(.din(n17548), .dout(n17545));
    jdff dff_A_J8hwEzkF8_1(.din(n17551), .dout(n17548));
    jdff dff_A_xIQ7gbAj8_1(.din(n17554), .dout(n17551));
    jdff dff_A_HG3c8mgp8_1(.din(n17557), .dout(n17554));
    jdff dff_A_9j1YVS9y4_1(.din(n1446), .dout(n17557));
    jdff dff_B_9MsAzG8q7_1(.din(n1401), .dout(n17561));
    jdff dff_B_Q8FR69JP3_1(.din(n17561), .dout(n17564));
    jdff dff_A_SXs6JVZ94_0(.din(n17569), .dout(n17566));
    jdff dff_A_Av51p9Z88_0(.din(n17572), .dout(n17569));
    jdff dff_A_3GBMsHpT0_0(.din(n17575), .dout(n17572));
    jdff dff_A_h8BPYLPv4_0(.din(n17578), .dout(n17575));
    jdff dff_A_4HO5pGpq3_0(.din(n1442), .dout(n17578));
    jdff dff_B_R97nAaRo7_1(.din(n1415), .dout(n17582));
    jdff dff_B_1aY1013Z9_1(.din(n17582), .dout(n17585));
    jdff dff_A_Rq9lncRI9_0(.din(n17590), .dout(n17587));
    jdff dff_A_tPE7GcZP7_0(.din(n1394), .dout(n17590));
    jdff dff_A_2CcqA3Wp5_1(.din(n17596), .dout(n17593));
    jdff dff_A_A4Tkes5G2_1(.din(n17599), .dout(n17596));
    jdff dff_A_5mzia1uA7_1(.din(n17602), .dout(n17599));
    jdff dff_A_TNobmL449_1(.din(n17605), .dout(n17602));
    jdff dff_A_AZoqO2o88_1(.din(n17608), .dout(n17605));
    jdff dff_A_tYXA1acM7_1(.din(n17611), .dout(n17608));
    jdff dff_A_794GiRhN5_1(.din(n17614), .dout(n17611));
    jdff dff_A_gnJKtLYn9_1(.din(n17617), .dout(n17614));
    jdff dff_A_0KXMix2R7_1(.din(n1394), .dout(n17617));
    jdff dff_A_a6MHcINx3_0(.din(n17623), .dout(n17620));
    jdff dff_A_P0ECXsiM0_0(.din(n17626), .dout(n17623));
    jdff dff_A_K58WcmBV6_0(.din(n17629), .dout(n17626));
    jdff dff_A_f7lECtP44_0(.din(n17632), .dout(n17629));
    jdff dff_A_9nNDEB4q5_0(.din(n17635), .dout(n17632));
    jdff dff_A_tvzVDIrl0_0(.din(n17638), .dout(n17635));
    jdff dff_A_4odcy0QT3_0(.din(n17641), .dout(n17638));
    jdff dff_A_emGEHPlv5_0(.din(n17644), .dout(n17641));
    jdff dff_A_FLmQyZFF2_0(.din(n17647), .dout(n17644));
    jdff dff_A_eybIkGQx0_0(.din(n1390), .dout(n17647));
    jdff dff_A_dDpbM4O12_1(.din(n17653), .dout(n17650));
    jdff dff_A_L6t83EmZ4_1(.din(n17656), .dout(n17653));
    jdff dff_A_fzUHu6em2_1(.din(n17659), .dout(n17656));
    jdff dff_A_6BKBDSwR7_1(.din(n17662), .dout(n17659));
    jdff dff_A_S8jMWJYh0_1(.din(n17665), .dout(n17662));
    jdff dff_A_baKVXvgD7_1(.din(n17668), .dout(n17665));
    jdff dff_A_LVitKlWq9_1(.din(n17671), .dout(n17668));
    jdff dff_A_HZOXCUEY6_1(.din(n17674), .dout(n17671));
    jdff dff_A_wlaO9dSU5_1(.din(n17677), .dout(n17674));
    jdff dff_A_bykxBIGm9_1(.din(n17680), .dout(n17677));
    jdff dff_A_7SqSx9tl8_1(.din(n17683), .dout(n17680));
    jdff dff_A_kmmA1FoC8_1(.din(n1352), .dout(n17683));
    jdff dff_A_R7HIKgfX4_2(.din(n1352), .dout(n17686));
    jdff dff_B_vH4nvQFC5_1(.din(n1561), .dout(n17690));
    jdff dff_B_AjURoX3e3_1(.din(n17690), .dout(n17693));
    jdff dff_B_H3ACOtNF0_1(.din(n17693), .dout(n17696));
    jdff dff_B_KOksx7kp3_1(.din(n17696), .dout(n17699));
    jdff dff_A_Bwoqm0jQ7_0(.din(n1621), .dout(n17701));
    jdff dff_A_9oJWk3Pj8_0(.din(n17707), .dout(n17704));
    jdff dff_A_nBMtiG5B5_0(.din(n17711), .dout(n17707));
    jdff dff_B_eLWVEYyq7_2(.din(n1613), .dout(n17711));
    jdff dff_A_UqyDJu4D5_1(.din(n1605), .dout(n17713));
    jdff dff_A_Icd7JuWI5_1(.din(n17719), .dout(n17716));
    jdff dff_A_RwBj1TKk8_1(.din(n17722), .dout(n17719));
    jdff dff_A_kXj7iwpq7_1(.din(n1602), .dout(n17722));
    jdff dff_A_yUGoHWWg2_2(.din(n1602), .dout(n17725));
    jdff dff_B_pTaV3zpz2_1(.din(n1590), .dout(n17729));
    jdff dff_A_kF5LMZdN8_1(.din(n17734), .dout(n17731));
    jdff dff_A_A1OPI00p8_1(.din(n1586), .dout(n17734));
    jdff dff_A_v4wmxwJL6_2(.din(n17740), .dout(n17737));
    jdff dff_A_2GrllwjR3_2(.din(n1586), .dout(n17740));
    jdff dff_A_PZOFBsFT3_0(.din(n17746), .dout(n17743));
    jdff dff_A_kjJgJEyu9_0(.din(n17749), .dout(n17746));
    jdff dff_A_UjSvI0Ny8_0(.din(n17759), .dout(n17749));
    jdff dff_B_5lt25F7C8_2(.din(n1571), .dout(n17753));
    jdff dff_B_uoIN38tW4_2(.din(n17753), .dout(n17756));
    jdff dff_B_aEhxahxj8_2(.din(n17756), .dout(n17759));
    jdff dff_A_Rkv4QTmw4_0(.din(n17801), .dout(n17761));
    jdff dff_A_dEMNL1jD3_1(.din(n17767), .dout(n17764));
    jdff dff_A_dlGEQ5aM2_1(.din(n17801), .dout(n17767));
    jdff dff_B_uHsnKISb7_3(.din(n3301), .dout(n17771));
    jdff dff_B_HCaRfry94_3(.din(n17771), .dout(n17774));
    jdff dff_B_CHuIJ1FZ5_3(.din(n17774), .dout(n17777));
    jdff dff_B_YKTqkjlu3_3(.din(n17777), .dout(n17780));
    jdff dff_B_GBC6tgsS0_3(.din(n17780), .dout(n17783));
    jdff dff_B_fNNYFwtv6_3(.din(n17783), .dout(n17786));
    jdff dff_B_vRBwmbzP8_3(.din(n17786), .dout(n17789));
    jdff dff_B_Zzbkcf9B6_3(.din(n17789), .dout(n17792));
    jdff dff_B_jM3c1MzT9_3(.din(n17792), .dout(n17795));
    jdff dff_B_EsOLP7h00_3(.din(n17795), .dout(n17798));
    jdff dff_B_18wAMXjE5_3(.din(n17798), .dout(n17801));
    jdff dff_A_ZB8TSSX78_0(.din(n17806), .dout(n17803));
    jdff dff_A_e4bLKr3j3_0(.din(n17809), .dout(n17806));
    jdff dff_A_C5lxxWGP2_0(.din(n17812), .dout(n17809));
    jdff dff_A_SFO0hwky9_0(.din(n17815), .dout(n17812));
    jdff dff_A_NT4AtEq80_0(.din(n17818), .dout(n17815));
    jdff dff_A_fQAJd3EL8_0(.din(n17821), .dout(n17818));
    jdff dff_A_5yjwNBpz2_0(.din(n17824), .dout(n17821));
    jdff dff_A_SelS453N1_0(.din(n17827), .dout(n17824));
    jdff dff_A_qrO3UpGs9_0(.din(n17830), .dout(n17827));
    jdff dff_A_p2bKUdqv7_0(.din(n17833), .dout(n17830));
    jdff dff_A_WH1e1dBZ8_0(.din(n17836), .dout(n17833));
    jdff dff_A_4Iu5KSXc9_0(.din(n17839), .dout(n17836));
    jdff dff_A_rkpjtdP25_0(.din(n17842), .dout(n17839));
    jdff dff_A_WgW83LfH5_0(.din(G4526), .dout(n17842));
    jdff dff_A_XxhC2lv49_2(.din(n17848), .dout(n17845));
    jdff dff_A_KjHWuwaD6_2(.din(n17851), .dout(n17848));
    jdff dff_A_wROp01Cy2_2(.din(n17854), .dout(n17851));
    jdff dff_A_N2XdCU0N8_2(.din(n17857), .dout(n17854));
    jdff dff_A_vIdPQ6qN6_2(.din(G4526), .dout(n17857));
    jdff dff_A_kaQKAcE87_1(.din(n17863), .dout(n17860));
    jdff dff_A_pQu3n5bo0_1(.din(n17866), .dout(n17863));
    jdff dff_A_rof2vaeC3_1(.din(n17869), .dout(n17866));
    jdff dff_A_KzlUK4uX4_1(.din(n17872), .dout(n17869));
    jdff dff_A_AAVX09nF5_1(.din(G4526), .dout(n17872));
    jdff dff_A_WFnPfGsW1_2(.din(n17878), .dout(n17875));
    jdff dff_A_9fMpdCo01_2(.din(n17881), .dout(n17878));
    jdff dff_A_xeuuFKas7_2(.din(n17884), .dout(n17881));
    jdff dff_A_n39KGL7a6_2(.din(n17887), .dout(n17884));
    jdff dff_A_1wZzwL965_2(.din(n17890), .dout(n17887));
    jdff dff_A_GbpiApuL1_2(.din(n17893), .dout(n17890));
    jdff dff_A_iubDQSNR7_2(.din(n17896), .dout(n17893));
    jdff dff_A_zIkDMXcZ8_2(.din(n17899), .dout(n17896));
    jdff dff_A_8se1Bysi3_2(.din(n17902), .dout(n17899));
    jdff dff_A_dKJHBT0a7_2(.din(n17905), .dout(n17902));
    jdff dff_A_5gsDfRXy5_2(.din(n17908), .dout(n17905));
    jdff dff_A_CThn5KxT9_2(.din(n17911), .dout(n17908));
    jdff dff_A_M4E1PaT90_2(.din(G4526), .dout(n17911));
    jdff dff_B_B17T1vBb1_0(.din(n5182), .dout(n17915));
    jdff dff_B_ivaSIiH18_0(.din(n17915), .dout(n17918));
    jdff dff_B_x4WMh0ub5_1(.din(n5166), .dout(n17921));
    jdff dff_B_mGxIXwGq5_1(.din(n17921), .dout(n17924));
    jdff dff_B_JV2A6PtL3_0(.din(n5174), .dout(n17927));
    jdff dff_A_aUsyYBN80_0(.din(n17932), .dout(n17929));
    jdff dff_A_iag1hkad3_0(.din(n1412), .dout(n17932));
    jdff dff_A_8w9F53vG1_1(.din(n17938), .dout(n17935));
    jdff dff_A_9ZEcId8N2_1(.din(n1336), .dout(n17938));
    jdff dff_A_pQHBUbia0_2(.din(n17944), .dout(n17941));
    jdff dff_A_agWuWEKK0_2(.din(n1336), .dout(n17944));
    jdff dff_A_xCO3wEwh1_1(.din(n17950), .dout(n17947));
    jdff dff_A_X7auKSNU3_1(.din(n17953), .dout(n17950));
    jdff dff_A_LkTghKlY6_1(.din(n17956), .dout(n17953));
    jdff dff_A_VZOYcmTX5_1(.din(n17959), .dout(n17956));
    jdff dff_A_TrvEIaVe4_1(.din(n17962), .dout(n17959));
    jdff dff_A_nwt7supn4_1(.din(n17965), .dout(n17962));
    jdff dff_A_QRLz4kkM9_1(.din(n17968), .dout(n17965));
    jdff dff_A_ge2KhoMZ4_1(.din(n17971), .dout(n17968));
    jdff dff_A_6QjljWL94_1(.din(n1431), .dout(n17971));
    jdff dff_B_bDqZolpk9_2(.din(n1374), .dout(n17975));
    jdff dff_B_BXVAVGHI5_2(.din(n17975), .dout(n17978));
    jdff dff_A_NJ16sLVB1_1(.din(n1419), .dout(n17980));
    jdff dff_A_PWYghY9h1_1(.din(n17990), .dout(n17983));
    jdff dff_B_XqLl8wJC5_2(.din(n1408), .dout(n17987));
    jdff dff_B_tJHYdyLG7_2(.din(n17987), .dout(n17990));
    jdff dff_B_0Y1cWcdy6_1(.din(n1340), .dout(n17993));
    jdff dff_B_Vz2Xni5H6_0(.din(G124), .dout(n17996));
    jdff dff_A_C4MMxLEe2_1(.din(n18001), .dout(n17998));
    jdff dff_A_pDhCs61i9_1(.din(n18004), .dout(n18001));
    jdff dff_A_1GwjxuQt0_1(.din(n18007), .dout(n18004));
    jdff dff_A_ggo8CN6V0_1(.din(G3743), .dout(n18007));
    jdff dff_A_689w9I3n8_1(.din(n3265), .dout(n18010));
    jdff dff_A_K5ZrTf5f6_2(.din(n18016), .dout(n18013));
    jdff dff_A_Hn9NuiWs7_2(.din(n18019), .dout(n18016));
    jdff dff_A_oezZcvdH4_2(.din(n18022), .dout(n18019));
    jdff dff_A_rewglPAF1_2(.din(n18025), .dout(n18022));
    jdff dff_A_kvJ3T86d4_2(.din(n18028), .dout(n18025));
    jdff dff_A_fJWjDWHI5_2(.din(n18031), .dout(n18028));
    jdff dff_A_QGWFhGrH0_2(.din(n18034), .dout(n18031));
    jdff dff_A_kWpWYWT03_2(.din(n18037), .dout(n18034));
    jdff dff_A_fO1wqDCy3_2(.din(n18040), .dout(n18037));
    jdff dff_A_rXWtukPu0_2(.din(n18043), .dout(n18040));
    jdff dff_A_WRFvq4cH9_2(.din(n18046), .dout(n18043));
    jdff dff_A_zIaVZtZh8_2(.din(n3265), .dout(n18046));
    jdff dff_B_izFmWNtm7_1(.din(n1311), .dout(n18050));
    jdff dff_B_pbQHyWMd6_0(.din(G100), .dout(n18053));
    jdff dff_A_10QKI3Aw8_0(.din(n18058), .dout(n18055));
    jdff dff_A_bSEYi0OK8_0(.din(n1307), .dout(n18058));
    jdff dff_A_zKkWUVVK3_2(.din(n18064), .dout(n18061));
    jdff dff_A_ouNZOQcj1_2(.din(n1307), .dout(n18064));
    jdff dff_A_WlxqNpyP9_1(.din(n18070), .dout(n18067));
    jdff dff_A_JwtNIGmY0_1(.din(n18073), .dout(n18070));
    jdff dff_A_ysaxURk58_1(.din(n18076), .dout(n18073));
    jdff dff_A_zBnmxytd5_1(.din(G3749), .dout(n18076));
    jdff dff_A_pDtEMtL68_1(.din(n18082), .dout(n18079));
    jdff dff_A_O7Jo6SXl6_1(.din(n18085), .dout(n18082));
    jdff dff_A_3wySArqs6_1(.din(n18088), .dout(n18085));
    jdff dff_A_NYHHFhxm7_1(.din(n18091), .dout(n18088));
    jdff dff_A_KayMGbHT1_1(.din(n18094), .dout(n18091));
    jdff dff_A_lLFT9WMi5_1(.din(n18097), .dout(n18094));
    jdff dff_A_wKof2ftZ0_1(.din(n18100), .dout(n18097));
    jdff dff_A_Zpy5zA207_1(.din(n18103), .dout(n18100));
    jdff dff_A_ym1Eibhz7_1(.din(n3354), .dout(n18103));
    jdff dff_B_lULSSn2v6_1(.din(n1378), .dout(n18107));
    jdff dff_B_0p2ojq8i8_0(.din(G130), .dout(n18110));
    jdff dff_A_SsXq4vV18_2(.din(n18115), .dout(n18112));
    jdff dff_A_fzEbCmmv1_2(.din(n18118), .dout(n18115));
    jdff dff_A_Myy3nlgI8_2(.din(n18121), .dout(n18118));
    jdff dff_A_Uq2Gp1T96_2(.din(G3729), .dout(n18121));
    jdff dff_A_IcAFC0mS5_1(.din(n18127), .dout(n18124));
    jdff dff_A_EZ39tuNI9_1(.din(n18130), .dout(n18127));
    jdff dff_A_OCosiyvZ4_1(.din(n18133), .dout(n18130));
    jdff dff_A_BUTLgfjH3_1(.din(n18136), .dout(n18133));
    jdff dff_A_AP5bIcxU3_1(.din(n18139), .dout(n18136));
    jdff dff_A_FtDVlJMR1_1(.din(n18142), .dout(n18139));
    jdff dff_A_CqddQdSg5_1(.din(n18145), .dout(n18142));
    jdff dff_A_JN1pSXGJ2_1(.din(n18148), .dout(n18145));
    jdff dff_A_kCk5ZQvw1_1(.din(n18151), .dout(n18148));
    jdff dff_A_eNTiblVA7_1(.din(n18155), .dout(n18151));
    jdff dff_B_dqPP4jvQ7_2(.din(n3344), .dout(n18155));
    jdff dff_B_XueDhB7k7_1(.din(n1359), .dout(n18158));
    jdff dff_B_XAFmI2px1_0(.din(G127), .dout(n18161));
    jdff dff_A_G4DRRie31_1(.din(n18166), .dout(n18163));
    jdff dff_A_hKABPv192_1(.din(n1355), .dout(n18166));
    jdff dff_A_SqMPRcZC1_2(.din(n18172), .dout(n18169));
    jdff dff_A_OtRZhWkL0_2(.din(n1355), .dout(n18172));
    jdff dff_A_BuLXbkO42_1(.din(n18178), .dout(n18175));
    jdff dff_A_7NPCYtjt2_1(.din(n18181), .dout(n18178));
    jdff dff_A_cHu6eCAS9_1(.din(n18184), .dout(n18181));
    jdff dff_A_wq8328gB9_1(.din(G3737), .dout(n18184));
    jdff dff_B_LtWNy6fy1_1(.din(n3275), .dout(n18188));
    jdff dff_B_rO78xemd1_1(.din(n18188), .dout(n18191));
    jdff dff_B_QrSECUrD8_1(.din(n18191), .dout(n18194));
    jdff dff_B_t2W9AHbf2_1(.din(n18194), .dout(n18197));
    jdff dff_B_xEOXWKi15_1(.din(n18197), .dout(n18200));
    jdff dff_B_bqNfjuoh2_1(.din(n18200), .dout(n18203));
    jdff dff_B_iuGSE1wl9_1(.din(n3278), .dout(n18206));
    jdff dff_B_bxk3BgJ65_1(.din(n18206), .dout(n18209));
    jdff dff_B_45VyFlQB5_1(.din(n18209), .dout(n18212));
    jdff dff_B_ZdHS22Za8_1(.din(n3179), .dout(n18215));
    jdff dff_B_Tjb98FfF9_1(.din(n18215), .dout(n18218));
    jdff dff_B_8t3jpyCn9_1(.din(n3182), .dout(n18221));
    jdff dff_B_q4V9eCAW1_1(.din(n3186), .dout(n18224));
    jdff dff_A_cysCXh4O1_1(.din(n18229), .dout(n18226));
    jdff dff_A_bU3HxgH34_1(.din(n1583), .dout(n18229));
    jdff dff_A_FTVzuvmY1_1(.din(n18235), .dout(n18232));
    jdff dff_A_Ynu68b1n4_1(.din(n18238), .dout(n18235));
    jdff dff_A_PDijplF23_1(.din(n1579), .dout(n18238));
    jdff dff_A_OGbbccXe7_1(.din(n18244), .dout(n18241));
    jdff dff_A_FuBjQKpz4_1(.din(n18247), .dout(n18244));
    jdff dff_A_reYAtjlZ6_1(.din(n18250), .dout(n18247));
    jdff dff_A_6P3ypGPy3_1(.din(n18253), .dout(n18250));
    jdff dff_A_NUufaEzV0_1(.din(n18256), .dout(n18253));
    jdff dff_A_2vpKgsog9_1(.din(n18259), .dout(n18256));
    jdff dff_A_ce8Cg8FA8_1(.din(n1575), .dout(n18259));
    jdff dff_A_qPcqFAnM7_2(.din(n18265), .dout(n18262));
    jdff dff_A_b96WBDRe8_2(.din(n18268), .dout(n18265));
    jdff dff_A_JmNaSGB24_2(.din(n18271), .dout(n18268));
    jdff dff_A_zA6O4Agt9_2(.din(n1575), .dout(n18271));
    jdff dff_A_XI4CKZxJ1_0(.din(n18277), .dout(n18274));
    jdff dff_A_kG63O8gK8_0(.din(n18280), .dout(n18277));
    jdff dff_A_hkHSszR17_0(.din(n18283), .dout(n18280));
    jdff dff_A_nJFI4ewU7_0(.din(n1568), .dout(n18283));
    jdff dff_A_tgb0i89Y2_0(.din(n18289), .dout(n18286));
    jdff dff_A_0e2A0Xbb2_0(.din(n18292), .dout(n18289));
    jdff dff_A_vjFv8mU73_0(.din(n18295), .dout(n18292));
    jdff dff_A_wcqp9dnb6_0(.din(n18298), .dout(n18295));
    jdff dff_A_9aQUFTwP0_0(.din(n1558), .dout(n18298));
    jdff dff_A_9fFv3bbF7_1(.din(n18304), .dout(n18301));
    jdff dff_A_ryOVwv122_1(.din(n18307), .dout(n18304));
    jdff dff_A_uuO3hIu62_1(.din(n18310), .dout(n18307));
    jdff dff_A_lAilQdBT7_1(.din(n18313), .dout(n18310));
    jdff dff_A_igMw3oUG4_1(.din(n18316), .dout(n18313));
    jdff dff_A_LWSNA2DT0_1(.din(n18319), .dout(n18316));
    jdff dff_A_wGTAaL9u6_1(.din(n1551), .dout(n18319));
    jdff dff_A_5np9xzlW8_0(.din(n18329), .dout(n18322));
    jdff dff_B_ddE4oc3f2_2(.din(n3272), .dout(n18326));
    jdff dff_B_IrzrFxNw3_2(.din(n18326), .dout(n18329));
    jdff dff_A_I66KZtkK6_1(.din(n18334), .dout(n18331));
    jdff dff_A_vpPwzcMV9_1(.din(n18337), .dout(n18334));
    jdff dff_A_Xub83BwO5_1(.din(n1547), .dout(n18337));
    jdff dff_A_Q4gslOok1_1(.din(n18343), .dout(n18340));
    jdff dff_A_VjQZaMGs4_1(.din(n18347), .dout(n18343));
    jdff dff_B_NUMZYu669_3(.din(n1531), .dout(n18347));
    jdff dff_A_tj16hwk92_0(.din(G29), .dout(n18349));
    jdff dff_A_3SL7naHL2_0(.din(n18355), .dout(n18352));
    jdff dff_A_L4pp5dTu2_0(.din(n18358), .dout(n18355));
    jdff dff_A_4z0juuWj9_0(.din(G3705), .dout(n18358));
    jdff dff_A_eorgmWoP0_2(.din(n18364), .dout(n18361));
    jdff dff_A_EIYJuf6S6_2(.din(n18367), .dout(n18364));
    jdff dff_A_YPFFoyh43_2(.din(G3705), .dout(n18367));
    jdff dff_A_V0MKqD0R2_2(.din(n18373), .dout(n18370));
    jdff dff_A_zSq0MprW8_2(.din(n18376), .dout(n18373));
    jdff dff_A_w8ug4njh8_2(.din(G3705), .dout(n18376));
    jdff dff_A_8QWeCkZB8_0(.din(n18382), .dout(n18379));
    jdff dff_A_qoaZTQKb9_0(.din(n18385), .dout(n18382));
    jdff dff_A_8u8zz0hI7_0(.din(n463), .dout(n18385));
    jdff dff_B_bRLAOsI35_3(.din(n452), .dout(n18389));
    jdff dff_A_ox4zSsWX7_0(.din(G41), .dout(n18391));
    jdff dff_A_8S7dEa0i4_1(.din(n18397), .dout(n18394));
    jdff dff_A_Pqsjnv4v5_0(.din(G3701), .dout(n18397));
    jdff dff_A_xcezbmkX0_1(.din(n18403), .dout(n18400));
    jdff dff_A_ueHqDwNa9_1(.din(n18406), .dout(n18403));
    jdff dff_A_J7rztvn01_1(.din(n18409), .dout(n18406));
    jdff dff_A_gg61SxAS4_1(.din(n1509), .dout(n18409));
    jdff dff_A_ZKNFV40b0_2(.din(n18415), .dout(n18412));
    jdff dff_A_fEUrzPyw6_2(.din(n1509), .dout(n18415));
    jdff dff_B_C6xg2Z3Z4_1(.din(n1497), .dout(n18419));
    jdff dff_B_imc1wVcA6_0(.din(G26), .dout(n18422));
    jdff dff_A_h8yjWpDz5_1(.din(G18), .dout(n18424));
    jdff dff_A_xz0LDdqJ7_0(.din(n18430), .dout(n18427));
    jdff dff_A_oKX0JHAy5_0(.din(n1493), .dout(n18430));
    jdff dff_A_CKSZqIIO0_2(.din(n18436), .dout(n18433));
    jdff dff_A_nAx8PBdD7_2(.din(n1493), .dout(n18436));
    jdff dff_A_EtjwFWbC2_1(.din(n18442), .dout(n18439));
    jdff dff_A_xJI09LtI7_1(.din(n18445), .dout(n18442));
    jdff dff_A_DkSJbuj46_1(.din(n18448), .dout(n18445));
    jdff dff_A_J8W2vvAm2_1(.din(n18451), .dout(n18448));
    jdff dff_A_9Y44Fhkp4_1(.din(n18454), .dout(n18451));
    jdff dff_A_EXP6f9nN5_1(.din(n18457), .dout(n18454));
    jdff dff_A_tikeZxdx1_1(.din(n1490), .dout(n18457));
    jdff dff_A_WtEFTgVK8_2(.din(n18463), .dout(n18460));
    jdff dff_A_6fV3kaxC7_2(.din(n18466), .dout(n18463));
    jdff dff_A_FSv2gqVb9_2(.din(n1490), .dout(n18466));
    jdff dff_B_eSI8rUsk5_1(.din(n1478), .dout(n18470));
    jdff dff_B_qWV7iYu50_0(.din(G23), .dout(n18473));
    jdff dff_A_9I9RuQo60_1(.din(n18478), .dout(n18475));
    jdff dff_A_imEWMNjW5_1(.din(n1474), .dout(n18478));
    jdff dff_A_lZJY7RlZ8_2(.din(n18484), .dout(n18481));
    jdff dff_A_woTKomL55_2(.din(n1474), .dout(n18484));
    jdff dff_A_1G0kWD285_1(.din(n18490), .dout(n18487));
    jdff dff_A_hyOa1aWo8_1(.din(n18493), .dout(n18490));
    jdff dff_A_PNL2GcxS9_1(.din(n18496), .dout(n18493));
    jdff dff_A_x0EMkzxd8_1(.din(G3717), .dout(n18496));
    jdff dff_A_jObMJrur8_0(.din(n18502), .dout(n18499));
    jdff dff_A_mKzlczDt4_0(.din(n18505), .dout(n18502));
    jdff dff_A_KtpsS1Dp0_0(.din(n18508), .dout(n18505));
    jdff dff_A_KEHmf4lu0_0(.din(n18511), .dout(n18508));
    jdff dff_A_Gs5W5Cso5_0(.din(n18514), .dout(n18511));
    jdff dff_A_ZBMCsjP81_0(.din(n18517), .dout(n18514));
    jdff dff_A_DhWvulUT0_0(.din(n18520), .dout(n18517));
    jdff dff_A_iimobAsk6_0(.din(n18523), .dout(n18520));
    jdff dff_A_3kVY6l0E9_0(.din(n1471), .dout(n18523));
    jdff dff_A_XNShdIJK8_1(.din(n18529), .dout(n18526));
    jdff dff_A_haP4sgFU1_1(.din(n18532), .dout(n18529));
    jdff dff_A_Qcljl5nJ4_1(.din(n18535), .dout(n18532));
    jdff dff_A_wND6vBd05_1(.din(n1471), .dout(n18535));
    jdff dff_B_A084MN4E7_1(.din(n1459), .dout(n18539));
    jdff dff_B_uNyvENmp2_0(.din(G103), .dout(n18542));
    jdff dff_A_sd1wNqVa8_2(.din(G18), .dout(n18544));
    jdff dff_A_QttmMOPF5_1(.din(n18550), .dout(n18547));
    jdff dff_A_Ovq9bdPh2_1(.din(n1455), .dout(n18550));
    jdff dff_A_zoLh1nev8_2(.din(n18556), .dout(n18553));
    jdff dff_A_erNsfYQU8_2(.din(n1455), .dout(n18556));
    jdff dff_A_nAynoQZb3_1(.din(n18562), .dout(n18559));
    jdff dff_A_8rwikamZ4_1(.din(n18565), .dout(n18562));
    jdff dff_A_OQjVDZsr1_1(.din(n18568), .dout(n18565));
    jdff dff_A_RgggCuSl6_1(.din(G3723), .dout(n18568));
    jdff dff_A_StDwqhMe5_1(.din(n5367), .dout(n18571));
    jdff dff_A_SeHU1hgo8_0(.din(n18571), .dout(n18574));
    jdff dff_A_T3vqXCwM2_0(.din(n18574), .dout(n18577));
    jdff dff_A_KoxgZOEF1_0(.din(n18577), .dout(n18580));
    jdff dff_A_bWecyCwf2_0(.din(n18580), .dout(n18583));
    jdff dff_A_AzJeX3xC8_0(.din(n18583), .dout(n18586));
    jdff dff_A_sL5HqlXH6_0(.din(n18586), .dout(n18589));
    jdff dff_A_jEGO6G9f3_0(.din(n18589), .dout(n18592));
    jdff dff_A_ol50RqS85_0(.din(n18592), .dout(n18595));
    jdff dff_A_V7E4IWB67_0(.din(n18595), .dout(n18598));
    jdff dff_A_WAdk7IEB6_0(.din(n18598), .dout(n18601));
    jdff dff_A_VOrFJZH17_0(.din(n18601), .dout(n18604));
    jdff dff_A_2mO9BGRa1_0(.din(n18604), .dout(n18607));
    jdff dff_A_7MkaPO6t1_0(.din(n18607), .dout(n18610));
    jdff dff_A_yGAzjzMr3_0(.din(n18610), .dout(n18613));
    jdff dff_A_QldLZweh7_0(.din(n18613), .dout(n18616));
    jdff dff_A_LRwXOCGr6_0(.din(n18616), .dout(n18619));
    jdff dff_A_cUxzD6Z81_0(.din(n18619), .dout(n18622));
    jdff dff_A_w1EMWtID4_0(.din(n18622), .dout(n18625));
    jdff dff_A_ICd6E9qD0_0(.din(n18625), .dout(n18628));
    jdff dff_A_Iewlz38u3_0(.din(n18628), .dout(n18631));
    jdff dff_A_UpIfp7D50_0(.din(n18631), .dout(n18634));
    jdff dff_A_TTQnkFMr2_0(.din(n18634), .dout(n18637));
    jdff dff_A_u2fcHUyK2_0(.din(n18637), .dout(n18640));
    jdff dff_A_KLwZPYX23_0(.din(n18640), .dout(n18643));
    jdff dff_A_YP5NO6vp6_0(.din(n18643), .dout(n18646));
    jdff dff_A_gV3La4kk8_0(.din(n18646), .dout(n18649));
    jdff dff_A_eB55MZVj0_0(.din(n18649), .dout(n18652));
    jdff dff_A_hKEjw8si9_0(.din(n18652), .dout(n18655));
    jdff dff_A_TGt4jsAn4_0(.din(n18655), .dout(n18658));
    jdff dff_A_fe7BH65t8_0(.din(n18658), .dout(n18661));
    jdff dff_A_NxO8nnaY3_0(.din(n18661), .dout(n18664));
    jdff dff_A_zwJRnC6v8_0(.din(n18664), .dout(n18667));
    jdff dff_A_5W9wWePd1_0(.din(n18667), .dout(n18670));
    jdff dff_A_WjqOJxsZ7_0(.din(n18670), .dout(n18673));
    jdff dff_A_7qk2mgLd2_0(.din(n18673), .dout(n18676));
    jdff dff_A_KhKWKH7s8_0(.din(n18676), .dout(n18679));
    jdff dff_A_3r7eKSVv3_0(.din(n18679), .dout(G2));
    jdff dff_A_lnaQpt5X0_1(.din(n5370), .dout(n18685));
    jdff dff_A_akETpjd88_0(.din(n18685), .dout(n18688));
    jdff dff_A_BRWlUsTg0_0(.din(n18688), .dout(n18691));
    jdff dff_A_jbhnCSo23_0(.din(n18691), .dout(n18694));
    jdff dff_A_CvAgXfbh8_0(.din(n18694), .dout(n18697));
    jdff dff_A_JOO9heH96_0(.din(n18697), .dout(n18700));
    jdff dff_A_cb9wsTnb1_0(.din(n18700), .dout(n18703));
    jdff dff_A_H4a7cb6z9_0(.din(n18703), .dout(n18706));
    jdff dff_A_0h2NUQrw5_0(.din(n18706), .dout(n18709));
    jdff dff_A_Er9z4s6r0_0(.din(n18709), .dout(n18712));
    jdff dff_A_nuuhhDUB4_0(.din(n18712), .dout(n18715));
    jdff dff_A_Y0tSrl9Y2_0(.din(n18715), .dout(n18718));
    jdff dff_A_c3mtIW6s2_0(.din(n18718), .dout(n18721));
    jdff dff_A_ZAyTBcY43_0(.din(n18721), .dout(n18724));
    jdff dff_A_Jb4htPzv0_0(.din(n18724), .dout(n18727));
    jdff dff_A_Kno6wHgd8_0(.din(n18727), .dout(n18730));
    jdff dff_A_asZ4ybZH5_0(.din(n18730), .dout(n18733));
    jdff dff_A_JcMTuyK20_0(.din(n18733), .dout(n18736));
    jdff dff_A_E9klAfIO8_0(.din(n18736), .dout(n18739));
    jdff dff_A_aFhFIG2k8_0(.din(n18739), .dout(n18742));
    jdff dff_A_pC5ZSHLp6_0(.din(n18742), .dout(n18745));
    jdff dff_A_dcZZo00o8_0(.din(n18745), .dout(n18748));
    jdff dff_A_57l2aB2k0_0(.din(n18748), .dout(n18751));
    jdff dff_A_cZa7Y2LU5_0(.din(n18751), .dout(n18754));
    jdff dff_A_VtBhzFD22_0(.din(n18754), .dout(n18757));
    jdff dff_A_ZEnx1QJh6_0(.din(n18757), .dout(n18760));
    jdff dff_A_4lPC5YK68_0(.din(n18760), .dout(n18763));
    jdff dff_A_vR5xfdH05_0(.din(n18763), .dout(n18766));
    jdff dff_A_5pce0cdr3_0(.din(n18766), .dout(n18769));
    jdff dff_A_ULxU10nX0_0(.din(n18769), .dout(n18772));
    jdff dff_A_vRm0XJat8_0(.din(n18772), .dout(n18775));
    jdff dff_A_NoNuQYZl5_0(.din(n18775), .dout(n18778));
    jdff dff_A_kqJI1BYN8_0(.din(n18778), .dout(n18781));
    jdff dff_A_33yiYwlA9_0(.din(n18781), .dout(n18784));
    jdff dff_A_FetlggL45_0(.din(n18784), .dout(n18787));
    jdff dff_A_qErBFBCE0_0(.din(n18787), .dout(n18790));
    jdff dff_A_h2R4569f1_0(.din(n18790), .dout(n18793));
    jdff dff_A_Ka7CPswc2_0(.din(n18793), .dout(G3));
    jdff dff_A_nByzfYml7_1(.din(n5373), .dout(n18799));
    jdff dff_A_J2dNTYMk9_0(.din(n18799), .dout(n18802));
    jdff dff_A_JlQzPGxX6_0(.din(n18802), .dout(n18805));
    jdff dff_A_hNT8dqZ58_0(.din(n18805), .dout(n18808));
    jdff dff_A_RilbSa9c8_0(.din(n18808), .dout(n18811));
    jdff dff_A_92Y45FwU6_0(.din(n18811), .dout(n18814));
    jdff dff_A_r1OWdJB38_0(.din(n18814), .dout(n18817));
    jdff dff_A_d3Oa4mE99_0(.din(n18817), .dout(n18820));
    jdff dff_A_m8qSEMKx5_0(.din(n18820), .dout(n18823));
    jdff dff_A_Kol595Eo5_0(.din(n18823), .dout(n18826));
    jdff dff_A_JTDHGrp79_0(.din(n18826), .dout(n18829));
    jdff dff_A_uwkSKMaW8_0(.din(n18829), .dout(n18832));
    jdff dff_A_vfBdUksM7_0(.din(n18832), .dout(n18835));
    jdff dff_A_02ugSumQ8_0(.din(n18835), .dout(n18838));
    jdff dff_A_7VOvqwFU2_0(.din(n18838), .dout(n18841));
    jdff dff_A_ZBMacSA12_0(.din(n18841), .dout(n18844));
    jdff dff_A_MugumP369_0(.din(n18844), .dout(n18847));
    jdff dff_A_1giOurUF3_0(.din(n18847), .dout(n18850));
    jdff dff_A_cor92Twd7_0(.din(n18850), .dout(n18853));
    jdff dff_A_3AHtEvjq0_0(.din(n18853), .dout(n18856));
    jdff dff_A_oDe15tqa7_0(.din(n18856), .dout(n18859));
    jdff dff_A_LzM80Iw81_0(.din(n18859), .dout(n18862));
    jdff dff_A_O3R5Eqsw7_0(.din(n18862), .dout(n18865));
    jdff dff_A_ax8DhLVl6_0(.din(n18865), .dout(n18868));
    jdff dff_A_XmvNloMl0_0(.din(n18868), .dout(n18871));
    jdff dff_A_v7bhiMPO1_0(.din(n18871), .dout(n18874));
    jdff dff_A_b14A3KCN9_0(.din(n18874), .dout(n18877));
    jdff dff_A_A8Uh0u299_0(.din(n18877), .dout(n18880));
    jdff dff_A_3vw78fWU2_0(.din(n18880), .dout(n18883));
    jdff dff_A_IVFV1qeD7_0(.din(n18883), .dout(n18886));
    jdff dff_A_cDn6Vza06_0(.din(n18886), .dout(n18889));
    jdff dff_A_U3Ur1uFB9_0(.din(n18889), .dout(n18892));
    jdff dff_A_gjmkPsRA6_0(.din(n18892), .dout(n18895));
    jdff dff_A_bm8orVMl7_0(.din(n18895), .dout(n18898));
    jdff dff_A_eTtD0IZL0_0(.din(n18898), .dout(n18901));
    jdff dff_A_v33XOql27_0(.din(n18901), .dout(n18904));
    jdff dff_A_mSnL3nEr0_0(.din(n18904), .dout(n18907));
    jdff dff_A_PC9rFL5d2_0(.din(n18907), .dout(G450));
    jdff dff_A_X1gH7vPc7_1(.din(n5376), .dout(n18913));
    jdff dff_A_ydkh7xRL8_0(.din(n18913), .dout(n18916));
    jdff dff_A_FCvaEbTU9_0(.din(n18916), .dout(n18919));
    jdff dff_A_yJcuvwvd0_0(.din(n18919), .dout(n18922));
    jdff dff_A_CLlJzujA7_0(.din(n18922), .dout(n18925));
    jdff dff_A_25TzLaDL2_0(.din(n18925), .dout(n18928));
    jdff dff_A_GCGFgT1b1_0(.din(n18928), .dout(n18931));
    jdff dff_A_svYKQF5g5_0(.din(n18931), .dout(n18934));
    jdff dff_A_7bwT5q4B2_0(.din(n18934), .dout(n18937));
    jdff dff_A_cfzUSbMH7_0(.din(n18937), .dout(n18940));
    jdff dff_A_zverzQER2_0(.din(n18940), .dout(n18943));
    jdff dff_A_0N9Zz3165_0(.din(n18943), .dout(n18946));
    jdff dff_A_q3lNx0fH3_0(.din(n18946), .dout(n18949));
    jdff dff_A_S9xkrVUq0_0(.din(n18949), .dout(n18952));
    jdff dff_A_KzOr32x21_0(.din(n18952), .dout(n18955));
    jdff dff_A_cbP674Kv9_0(.din(n18955), .dout(n18958));
    jdff dff_A_atdhSgYQ0_0(.din(n18958), .dout(n18961));
    jdff dff_A_XEooD6Y84_0(.din(n18961), .dout(n18964));
    jdff dff_A_PMEDLE3F2_0(.din(n18964), .dout(n18967));
    jdff dff_A_unq1obuO9_0(.din(n18967), .dout(n18970));
    jdff dff_A_9pChAC9s5_0(.din(n18970), .dout(n18973));
    jdff dff_A_OxLpBcm77_0(.din(n18973), .dout(n18976));
    jdff dff_A_DNwDOW2w1_0(.din(n18976), .dout(n18979));
    jdff dff_A_MmIfOmpd2_0(.din(n18979), .dout(n18982));
    jdff dff_A_UhhXUQQY4_0(.din(n18982), .dout(n18985));
    jdff dff_A_xN8E6Ghb2_0(.din(n18985), .dout(n18988));
    jdff dff_A_PXYf0dZq4_0(.din(n18988), .dout(n18991));
    jdff dff_A_hfN5wi7i8_0(.din(n18991), .dout(n18994));
    jdff dff_A_oPajINVY9_0(.din(n18994), .dout(n18997));
    jdff dff_A_pnYtcv6T3_0(.din(n18997), .dout(n19000));
    jdff dff_A_YkqGDftS9_0(.din(n19000), .dout(n19003));
    jdff dff_A_RtToPjVr3_0(.din(n19003), .dout(n19006));
    jdff dff_A_ilREnJUH4_0(.din(n19006), .dout(n19009));
    jdff dff_A_FeK7bATw0_0(.din(n19009), .dout(n19012));
    jdff dff_A_lKYIe5Vw6_0(.din(n19012), .dout(n19015));
    jdff dff_A_wWOuanCo7_0(.din(n19015), .dout(n19018));
    jdff dff_A_E4l51J4X3_0(.din(n19018), .dout(n19021));
    jdff dff_A_f9ECAxSt3_0(.din(n19021), .dout(G448));
    jdff dff_A_uLsdXGj77_1(.din(n5379), .dout(n19027));
    jdff dff_A_NX1FLLKx8_0(.din(n19027), .dout(n19030));
    jdff dff_A_i1fIY9VA9_0(.din(n19030), .dout(n19033));
    jdff dff_A_vinnMVKQ3_0(.din(n19033), .dout(n19036));
    jdff dff_A_Z6MLrGcd7_0(.din(n19036), .dout(n19039));
    jdff dff_A_8HtCx68v9_0(.din(n19039), .dout(n19042));
    jdff dff_A_gZq3zVus4_0(.din(n19042), .dout(n19045));
    jdff dff_A_l7tOmevN2_0(.din(n19045), .dout(n19048));
    jdff dff_A_OgqSDkSL2_0(.din(n19048), .dout(n19051));
    jdff dff_A_lPJuA1QS4_0(.din(n19051), .dout(n19054));
    jdff dff_A_nn0FKwip9_0(.din(n19054), .dout(n19057));
    jdff dff_A_NsBrquGu9_0(.din(n19057), .dout(n19060));
    jdff dff_A_CSnJrBrw5_0(.din(n19060), .dout(n19063));
    jdff dff_A_gP7CTIag1_0(.din(n19063), .dout(n19066));
    jdff dff_A_L5iHt3dr8_0(.din(n19066), .dout(n19069));
    jdff dff_A_K6JvbFWp4_0(.din(n19069), .dout(n19072));
    jdff dff_A_9fcGjbCy8_0(.din(n19072), .dout(n19075));
    jdff dff_A_wS6cb22j4_0(.din(n19075), .dout(n19078));
    jdff dff_A_GX3cdPUI3_0(.din(n19078), .dout(n19081));
    jdff dff_A_Lkvpz61y5_0(.din(n19081), .dout(n19084));
    jdff dff_A_GQehuQGn9_0(.din(n19084), .dout(n19087));
    jdff dff_A_BMg5TUVv2_0(.din(n19087), .dout(n19090));
    jdff dff_A_wZ2f8pTL6_0(.din(n19090), .dout(n19093));
    jdff dff_A_83ZOiplb4_0(.din(n19093), .dout(n19096));
    jdff dff_A_cE5GgqAB8_0(.din(n19096), .dout(n19099));
    jdff dff_A_GgNHQkRp9_0(.din(n19099), .dout(n19102));
    jdff dff_A_vIWR0YOL4_0(.din(n19102), .dout(n19105));
    jdff dff_A_w0W6kF634_0(.din(n19105), .dout(n19108));
    jdff dff_A_8os3EzAM6_0(.din(n19108), .dout(n19111));
    jdff dff_A_7nuPcMTJ8_0(.din(n19111), .dout(n19114));
    jdff dff_A_fXIeBo3c7_0(.din(n19114), .dout(n19117));
    jdff dff_A_DTuzhzlB3_0(.din(n19117), .dout(n19120));
    jdff dff_A_vbAbtqJV7_0(.din(n19120), .dout(n19123));
    jdff dff_A_FDpsTSAO0_0(.din(n19123), .dout(n19126));
    jdff dff_A_3PMa9iHI6_0(.din(n19126), .dout(n19129));
    jdff dff_A_cPOODtLB6_0(.din(n19129), .dout(n19132));
    jdff dff_A_cH04DPs96_0(.din(n19132), .dout(n19135));
    jdff dff_A_ybJM6jXC5_0(.din(n19135), .dout(G444));
    jdff dff_A_2l1hqVy46_1(.din(n5382), .dout(n19141));
    jdff dff_A_9d3UVCu13_0(.din(n19141), .dout(n19144));
    jdff dff_A_KGfjFnLn0_0(.din(n19144), .dout(n19147));
    jdff dff_A_Z6Fss6RC9_0(.din(n19147), .dout(n19150));
    jdff dff_A_tf6WkaWM4_0(.din(n19150), .dout(n19153));
    jdff dff_A_Jau20yRE0_0(.din(n19153), .dout(n19156));
    jdff dff_A_H4CrkWjr8_0(.din(n19156), .dout(n19159));
    jdff dff_A_qMt4R6XX4_0(.din(n19159), .dout(n19162));
    jdff dff_A_tRWnFen94_0(.din(n19162), .dout(n19165));
    jdff dff_A_pPyLbdqA5_0(.din(n19165), .dout(n19168));
    jdff dff_A_aFPXLgXY1_0(.din(n19168), .dout(n19171));
    jdff dff_A_8MX3tftK2_0(.din(n19171), .dout(n19174));
    jdff dff_A_mSxr0lMG2_0(.din(n19174), .dout(n19177));
    jdff dff_A_CAYi5kPi8_0(.din(n19177), .dout(n19180));
    jdff dff_A_tk7VeiD46_0(.din(n19180), .dout(n19183));
    jdff dff_A_2YjvvqZ29_0(.din(n19183), .dout(n19186));
    jdff dff_A_oYZRwpwO7_0(.din(n19186), .dout(n19189));
    jdff dff_A_dic5qb4a4_0(.din(n19189), .dout(n19192));
    jdff dff_A_OmWpxsGv9_0(.din(n19192), .dout(n19195));
    jdff dff_A_bZp5g0I93_0(.din(n19195), .dout(n19198));
    jdff dff_A_kinliT5j2_0(.din(n19198), .dout(n19201));
    jdff dff_A_5Hc9Ldb98_0(.din(n19201), .dout(n19204));
    jdff dff_A_Dwc2Xno58_0(.din(n19204), .dout(n19207));
    jdff dff_A_rmc3rdFx6_0(.din(n19207), .dout(n19210));
    jdff dff_A_3HQ4aECa5_0(.din(n19210), .dout(n19213));
    jdff dff_A_6L5t83EB3_0(.din(n19213), .dout(n19216));
    jdff dff_A_jNTqtUKP1_0(.din(n19216), .dout(n19219));
    jdff dff_A_e5cC8NpR5_0(.din(n19219), .dout(n19222));
    jdff dff_A_vFOy2fyY4_0(.din(n19222), .dout(n19225));
    jdff dff_A_8EL24QTX0_0(.din(n19225), .dout(n19228));
    jdff dff_A_nqbQipO56_0(.din(n19228), .dout(n19231));
    jdff dff_A_5cxFsShh1_0(.din(n19231), .dout(n19234));
    jdff dff_A_nowipb605_0(.din(n19234), .dout(n19237));
    jdff dff_A_SHE8aMfO7_0(.din(n19237), .dout(n19240));
    jdff dff_A_5wO5d7hK3_0(.din(n19240), .dout(n19243));
    jdff dff_A_dfNJmO6F8_0(.din(n19243), .dout(n19246));
    jdff dff_A_q2Ks7Jvr8_0(.din(n19246), .dout(n19249));
    jdff dff_A_2rX7MfhW7_0(.din(n19249), .dout(G442));
    jdff dff_A_HiWLfWKP7_1(.din(n5385), .dout(n19255));
    jdff dff_A_0UCvrhVi4_0(.din(n19255), .dout(n19258));
    jdff dff_A_n8cv8puG5_0(.din(n19258), .dout(n19261));
    jdff dff_A_RYvqZK1l1_0(.din(n19261), .dout(n19264));
    jdff dff_A_ENzhW5jK9_0(.din(n19264), .dout(n19267));
    jdff dff_A_dVMDnWrn3_0(.din(n19267), .dout(n19270));
    jdff dff_A_8e1c2y0W5_0(.din(n19270), .dout(n19273));
    jdff dff_A_xRJmrmeE0_0(.din(n19273), .dout(n19276));
    jdff dff_A_ATMFP5mw9_0(.din(n19276), .dout(n19279));
    jdff dff_A_fNIQnVzC4_0(.din(n19279), .dout(n19282));
    jdff dff_A_C12bCA4o3_0(.din(n19282), .dout(n19285));
    jdff dff_A_8ZbMhV4i6_0(.din(n19285), .dout(n19288));
    jdff dff_A_y9pz8Om91_0(.din(n19288), .dout(n19291));
    jdff dff_A_9NF812NG2_0(.din(n19291), .dout(n19294));
    jdff dff_A_iqBQPIcQ3_0(.din(n19294), .dout(n19297));
    jdff dff_A_RCkWIBlx8_0(.din(n19297), .dout(n19300));
    jdff dff_A_bY3ubHh02_0(.din(n19300), .dout(n19303));
    jdff dff_A_QfxCFLnc7_0(.din(n19303), .dout(n19306));
    jdff dff_A_xfmKH9L01_0(.din(n19306), .dout(n19309));
    jdff dff_A_KpNIUVEs0_0(.din(n19309), .dout(n19312));
    jdff dff_A_MIrF1B9i2_0(.din(n19312), .dout(n19315));
    jdff dff_A_HzGvQglx0_0(.din(n19315), .dout(n19318));
    jdff dff_A_4twZSC3O2_0(.din(n19318), .dout(n19321));
    jdff dff_A_kSagvAEW3_0(.din(n19321), .dout(n19324));
    jdff dff_A_IolfRFdE2_0(.din(n19324), .dout(n19327));
    jdff dff_A_GriAU1Pt1_0(.din(n19327), .dout(n19330));
    jdff dff_A_667x8J2q8_0(.din(n19330), .dout(n19333));
    jdff dff_A_vLmPdVaY4_0(.din(n19333), .dout(n19336));
    jdff dff_A_9cXdnejb2_0(.din(n19336), .dout(n19339));
    jdff dff_A_c9vUUgNJ6_0(.din(n19339), .dout(n19342));
    jdff dff_A_dSk0q1FY6_0(.din(n19342), .dout(n19345));
    jdff dff_A_p8LBrKaF4_0(.din(n19345), .dout(n19348));
    jdff dff_A_LmEwFyAl4_0(.din(n19348), .dout(n19351));
    jdff dff_A_ipSodC7T5_0(.din(n19351), .dout(n19354));
    jdff dff_A_frVC1RHd9_0(.din(n19354), .dout(n19357));
    jdff dff_A_9SQwtwIr4_0(.din(n19357), .dout(n19360));
    jdff dff_A_pYiQIiIQ6_0(.din(n19360), .dout(n19363));
    jdff dff_A_S2TA1OUr4_0(.din(n19363), .dout(G440));
    jdff dff_A_kvGxlUzO4_1(.din(n5388), .dout(n19369));
    jdff dff_A_HQiO5ttM3_0(.din(n19369), .dout(n19372));
    jdff dff_A_wDMwpEe39_0(.din(n19372), .dout(n19375));
    jdff dff_A_D25LVPdq9_0(.din(n19375), .dout(n19378));
    jdff dff_A_LdqQ8GS96_0(.din(n19378), .dout(n19381));
    jdff dff_A_g5SNYsFV2_0(.din(n19381), .dout(n19384));
    jdff dff_A_7VIbVF2i0_0(.din(n19384), .dout(n19387));
    jdff dff_A_u5gsozjE8_0(.din(n19387), .dout(n19390));
    jdff dff_A_bYkPkdv60_0(.din(n19390), .dout(n19393));
    jdff dff_A_h6GV5PaT1_0(.din(n19393), .dout(n19396));
    jdff dff_A_5GOGn6aE4_0(.din(n19396), .dout(n19399));
    jdff dff_A_4RwAOoPy3_0(.din(n19399), .dout(n19402));
    jdff dff_A_PO8kIc2X7_0(.din(n19402), .dout(n19405));
    jdff dff_A_G0oO1yNn5_0(.din(n19405), .dout(n19408));
    jdff dff_A_wcG2Op2J1_0(.din(n19408), .dout(n19411));
    jdff dff_A_GH70SxUr8_0(.din(n19411), .dout(n19414));
    jdff dff_A_CcWFvBEL0_0(.din(n19414), .dout(n19417));
    jdff dff_A_sf5jpRQu8_0(.din(n19417), .dout(n19420));
    jdff dff_A_0WgsX7tT0_0(.din(n19420), .dout(n19423));
    jdff dff_A_nnPg39Tz2_0(.din(n19423), .dout(n19426));
    jdff dff_A_SHnaC6LD5_0(.din(n19426), .dout(n19429));
    jdff dff_A_WaTtFhQm2_0(.din(n19429), .dout(n19432));
    jdff dff_A_hD38IotZ8_0(.din(n19432), .dout(n19435));
    jdff dff_A_rGzf70ts7_0(.din(n19435), .dout(n19438));
    jdff dff_A_xRDBuaYF9_0(.din(n19438), .dout(n19441));
    jdff dff_A_xcQvfbi58_0(.din(n19441), .dout(n19444));
    jdff dff_A_SQGo8CdU4_0(.din(n19444), .dout(n19447));
    jdff dff_A_LWbBRtU55_0(.din(n19447), .dout(n19450));
    jdff dff_A_SvM85YHX4_0(.din(n19450), .dout(n19453));
    jdff dff_A_c7snQ1q51_0(.din(n19453), .dout(n19456));
    jdff dff_A_14omzql55_0(.din(n19456), .dout(n19459));
    jdff dff_A_uIKWQI7U1_0(.din(n19459), .dout(n19462));
    jdff dff_A_GTQTm0DE4_0(.din(n19462), .dout(n19465));
    jdff dff_A_wYryfeQU2_0(.din(n19465), .dout(n19468));
    jdff dff_A_R2ME4zqR4_0(.din(n19468), .dout(n19471));
    jdff dff_A_V5LgGH9N4_0(.din(n19471), .dout(n19474));
    jdff dff_A_wCgTN6nU2_0(.din(n19474), .dout(n19477));
    jdff dff_A_pp9IsZJP3_0(.din(n19477), .dout(G438));
    jdff dff_A_fKxVyEvG8_1(.din(n5391), .dout(n19483));
    jdff dff_A_F92hdeRJ0_0(.din(n19483), .dout(n19486));
    jdff dff_A_lh4qTxSA6_0(.din(n19486), .dout(n19489));
    jdff dff_A_Lj4aZEHl3_0(.din(n19489), .dout(n19492));
    jdff dff_A_Ch9i7imW9_0(.din(n19492), .dout(n19495));
    jdff dff_A_kCkxOE5N3_0(.din(n19495), .dout(n19498));
    jdff dff_A_dnWzRb6X7_0(.din(n19498), .dout(n19501));
    jdff dff_A_2SrkhawT5_0(.din(n19501), .dout(n19504));
    jdff dff_A_J4ggTXvG5_0(.din(n19504), .dout(n19507));
    jdff dff_A_laU8SMs35_0(.din(n19507), .dout(n19510));
    jdff dff_A_z1f7J1W22_0(.din(n19510), .dout(n19513));
    jdff dff_A_FsoH9K6T3_0(.din(n19513), .dout(n19516));
    jdff dff_A_IoUyw4J14_0(.din(n19516), .dout(n19519));
    jdff dff_A_QURQmPgQ3_0(.din(n19519), .dout(n19522));
    jdff dff_A_aLGroFPl3_0(.din(n19522), .dout(n19525));
    jdff dff_A_LfcpGE3l3_0(.din(n19525), .dout(n19528));
    jdff dff_A_EqJmcoBQ9_0(.din(n19528), .dout(n19531));
    jdff dff_A_LUMKoF214_0(.din(n19531), .dout(n19534));
    jdff dff_A_3yUQLkN69_0(.din(n19534), .dout(n19537));
    jdff dff_A_bqDVKuKK3_0(.din(n19537), .dout(n19540));
    jdff dff_A_SAUFHYGW9_0(.din(n19540), .dout(n19543));
    jdff dff_A_TAfyRZJC0_0(.din(n19543), .dout(n19546));
    jdff dff_A_LBPJll499_0(.din(n19546), .dout(n19549));
    jdff dff_A_c2nudf8R7_0(.din(n19549), .dout(n19552));
    jdff dff_A_KcmDLKqn1_0(.din(n19552), .dout(n19555));
    jdff dff_A_s16URw4I2_0(.din(n19555), .dout(n19558));
    jdff dff_A_5JPYUQsM5_0(.din(n19558), .dout(n19561));
    jdff dff_A_Idu8qWNB6_0(.din(n19561), .dout(n19564));
    jdff dff_A_1WWExI6x8_0(.din(n19564), .dout(n19567));
    jdff dff_A_0mnoZRSQ5_0(.din(n19567), .dout(n19570));
    jdff dff_A_CF2GSWek0_0(.din(n19570), .dout(n19573));
    jdff dff_A_VQpVfuAR4_0(.din(n19573), .dout(n19576));
    jdff dff_A_e170Ure11_0(.din(n19576), .dout(n19579));
    jdff dff_A_3VILppcH7_0(.din(n19579), .dout(n19582));
    jdff dff_A_l4NAm9en6_0(.din(n19582), .dout(n19585));
    jdff dff_A_fDmTOJTi1_0(.din(n19585), .dout(n19588));
    jdff dff_A_hph6m4e00_0(.din(n19588), .dout(n19591));
    jdff dff_A_PSZgYxFA9_0(.din(n19591), .dout(G496));
    jdff dff_A_AcwEvtBl8_1(.din(n5394), .dout(n19597));
    jdff dff_A_6OWjTLXC6_0(.din(n19597), .dout(n19600));
    jdff dff_A_rpdzzsy26_0(.din(n19600), .dout(n19603));
    jdff dff_A_RRnxiAJm6_0(.din(n19603), .dout(n19606));
    jdff dff_A_Prlg8BjP1_0(.din(n19606), .dout(n19609));
    jdff dff_A_3bCnMy7x4_0(.din(n19609), .dout(n19612));
    jdff dff_A_LGjH8Pn65_0(.din(n19612), .dout(n19615));
    jdff dff_A_VYde3mL26_0(.din(n19615), .dout(n19618));
    jdff dff_A_aBaFFw074_0(.din(n19618), .dout(n19621));
    jdff dff_A_YqWJ6E5b9_0(.din(n19621), .dout(n19624));
    jdff dff_A_ZRs2QVpA7_0(.din(n19624), .dout(n19627));
    jdff dff_A_9oebRl9I6_0(.din(n19627), .dout(n19630));
    jdff dff_A_hpjYXzxN6_0(.din(n19630), .dout(n19633));
    jdff dff_A_OBgwRlmI9_0(.din(n19633), .dout(n19636));
    jdff dff_A_EnWHsSSQ6_0(.din(n19636), .dout(n19639));
    jdff dff_A_ZqKAs4xj1_0(.din(n19639), .dout(n19642));
    jdff dff_A_mcCDbzoh3_0(.din(n19642), .dout(n19645));
    jdff dff_A_4APlkpIW4_0(.din(n19645), .dout(n19648));
    jdff dff_A_yGrE6SZE2_0(.din(n19648), .dout(n19651));
    jdff dff_A_ch7R156V2_0(.din(n19651), .dout(n19654));
    jdff dff_A_bbSEe4Wi5_0(.din(n19654), .dout(n19657));
    jdff dff_A_ebmEU7UJ1_0(.din(n19657), .dout(n19660));
    jdff dff_A_ww67YbTu2_0(.din(n19660), .dout(n19663));
    jdff dff_A_HNskSIVu3_0(.din(n19663), .dout(n19666));
    jdff dff_A_VKUvB8OA4_0(.din(n19666), .dout(n19669));
    jdff dff_A_XE5PC3Zx2_0(.din(n19669), .dout(n19672));
    jdff dff_A_iRRtSOHo3_0(.din(n19672), .dout(n19675));
    jdff dff_A_UhSxZrF77_0(.din(n19675), .dout(n19678));
    jdff dff_A_kTeJyuOT2_0(.din(n19678), .dout(n19681));
    jdff dff_A_vWv3fmiR5_0(.din(n19681), .dout(n19684));
    jdff dff_A_w1lbupO53_0(.din(n19684), .dout(n19687));
    jdff dff_A_nBVCXKhB1_0(.din(n19687), .dout(n19690));
    jdff dff_A_QbV8s2JN4_0(.din(n19690), .dout(n19693));
    jdff dff_A_0d02QCDj3_0(.din(n19693), .dout(n19696));
    jdff dff_A_Cy6LBfrM8_0(.din(n19696), .dout(n19699));
    jdff dff_A_K8hUt43B8_0(.din(n19699), .dout(n19702));
    jdff dff_A_JecLXnvU4_0(.din(n19702), .dout(n19705));
    jdff dff_A_NGD2okon1_0(.din(n19705), .dout(G494));
    jdff dff_A_z4lHrBEn5_1(.din(n5397), .dout(n19711));
    jdff dff_A_wMXkQfNZ7_0(.din(n19711), .dout(n19714));
    jdff dff_A_PIHhjbMF1_0(.din(n19714), .dout(n19717));
    jdff dff_A_7XwEtK6h9_0(.din(n19717), .dout(n19720));
    jdff dff_A_VeQmwW8d0_0(.din(n19720), .dout(n19723));
    jdff dff_A_1IcuaTuF8_0(.din(n19723), .dout(n19726));
    jdff dff_A_Q0bxyaBG9_0(.din(n19726), .dout(n19729));
    jdff dff_A_AC23EK8I0_0(.din(n19729), .dout(n19732));
    jdff dff_A_1YFYwp1q0_0(.din(n19732), .dout(n19735));
    jdff dff_A_0uSb1EZf5_0(.din(n19735), .dout(n19738));
    jdff dff_A_fba7M4lh6_0(.din(n19738), .dout(n19741));
    jdff dff_A_1V4bVSun7_0(.din(n19741), .dout(n19744));
    jdff dff_A_GWUFa7EB2_0(.din(n19744), .dout(n19747));
    jdff dff_A_ydN3znsn0_0(.din(n19747), .dout(n19750));
    jdff dff_A_Wwalok0z5_0(.din(n19750), .dout(n19753));
    jdff dff_A_hVfJakKe3_0(.din(n19753), .dout(n19756));
    jdff dff_A_c6vz4bpA5_0(.din(n19756), .dout(n19759));
    jdff dff_A_eAhWjZ4y4_0(.din(n19759), .dout(n19762));
    jdff dff_A_5QBs58y93_0(.din(n19762), .dout(n19765));
    jdff dff_A_QME7xHGK3_0(.din(n19765), .dout(n19768));
    jdff dff_A_KUCDi4qU8_0(.din(n19768), .dout(n19771));
    jdff dff_A_bKhBPAJF1_0(.din(n19771), .dout(n19774));
    jdff dff_A_M1Vyk1d97_0(.din(n19774), .dout(n19777));
    jdff dff_A_n9aHY8JG4_0(.din(n19777), .dout(n19780));
    jdff dff_A_jnuSaW5o8_0(.din(n19780), .dout(n19783));
    jdff dff_A_WUqwmtjw0_0(.din(n19783), .dout(n19786));
    jdff dff_A_KQt9Ye494_0(.din(n19786), .dout(n19789));
    jdff dff_A_mNYPkUIT3_0(.din(n19789), .dout(n19792));
    jdff dff_A_WPAyqyhM6_0(.din(n19792), .dout(n19795));
    jdff dff_A_sDJbfh4v8_0(.din(n19795), .dout(n19798));
    jdff dff_A_eF4yq6ZG2_0(.din(n19798), .dout(n19801));
    jdff dff_A_rRUU0rwy4_0(.din(n19801), .dout(n19804));
    jdff dff_A_SRz56pQD2_0(.din(n19804), .dout(n19807));
    jdff dff_A_U23LyN9s0_0(.din(n19807), .dout(n19810));
    jdff dff_A_houm0qa04_0(.din(n19810), .dout(n19813));
    jdff dff_A_EWxXOe9A8_0(.din(n19813), .dout(n19816));
    jdff dff_A_RA96IEze4_0(.din(n19816), .dout(n19819));
    jdff dff_A_8oeq2vBk5_0(.din(n19819), .dout(G492));
    jdff dff_A_36IIFIIA7_1(.din(n5400), .dout(n19825));
    jdff dff_A_FkmA8tq38_0(.din(n19825), .dout(n19828));
    jdff dff_A_9aGlH3DO0_0(.din(n19828), .dout(n19831));
    jdff dff_A_lMSm5W6U6_0(.din(n19831), .dout(n19834));
    jdff dff_A_prz6a1sx7_0(.din(n19834), .dout(n19837));
    jdff dff_A_3cQzEwjl6_0(.din(n19837), .dout(n19840));
    jdff dff_A_A3wrVfxj6_0(.din(n19840), .dout(n19843));
    jdff dff_A_ngJ6Fizn9_0(.din(n19843), .dout(n19846));
    jdff dff_A_ePkytt8P6_0(.din(n19846), .dout(n19849));
    jdff dff_A_nKeN6kf55_0(.din(n19849), .dout(n19852));
    jdff dff_A_ukFQpkC67_0(.din(n19852), .dout(n19855));
    jdff dff_A_9wB1IUS94_0(.din(n19855), .dout(n19858));
    jdff dff_A_0sQPsP7I3_0(.din(n19858), .dout(n19861));
    jdff dff_A_IYpIvJiJ2_0(.din(n19861), .dout(n19864));
    jdff dff_A_OvqoPMTn3_0(.din(n19864), .dout(n19867));
    jdff dff_A_9QwibUCc8_0(.din(n19867), .dout(n19870));
    jdff dff_A_R1ICejDp3_0(.din(n19870), .dout(n19873));
    jdff dff_A_oN2D5d8m5_0(.din(n19873), .dout(n19876));
    jdff dff_A_YuYOUTou0_0(.din(n19876), .dout(n19879));
    jdff dff_A_U6BGYJb88_0(.din(n19879), .dout(n19882));
    jdff dff_A_47TVOq246_0(.din(n19882), .dout(n19885));
    jdff dff_A_PbVCMIuH5_0(.din(n19885), .dout(n19888));
    jdff dff_A_ufFMvqlb0_0(.din(n19888), .dout(n19891));
    jdff dff_A_1M54oIVD0_0(.din(n19891), .dout(n19894));
    jdff dff_A_BrK1dTY31_0(.din(n19894), .dout(n19897));
    jdff dff_A_YaIfHXcC6_0(.din(n19897), .dout(n19900));
    jdff dff_A_gcwgr0Rl8_0(.din(n19900), .dout(n19903));
    jdff dff_A_ybpOetFU3_0(.din(n19903), .dout(n19906));
    jdff dff_A_6hEOK7Eq8_0(.din(n19906), .dout(n19909));
    jdff dff_A_4Yhz2anG0_0(.din(n19909), .dout(n19912));
    jdff dff_A_zRVHWq2I9_0(.din(n19912), .dout(n19915));
    jdff dff_A_32HSNbuY5_0(.din(n19915), .dout(n19918));
    jdff dff_A_xA2Dcb131_0(.din(n19918), .dout(n19921));
    jdff dff_A_cd7WkMJc1_0(.din(n19921), .dout(n19924));
    jdff dff_A_P6yfV3Ci3_0(.din(n19924), .dout(n19927));
    jdff dff_A_DKS9rln26_0(.din(n19927), .dout(n19930));
    jdff dff_A_gKtsmjWV7_0(.din(n19930), .dout(n19933));
    jdff dff_A_Kcmhynvt0_0(.din(n19933), .dout(G490));
    jdff dff_A_DXzas7OV3_1(.din(n5403), .dout(n19939));
    jdff dff_A_DitevIQt4_0(.din(n19939), .dout(n19942));
    jdff dff_A_gXqQdEKN7_0(.din(n19942), .dout(n19945));
    jdff dff_A_cqb7lCs85_0(.din(n19945), .dout(n19948));
    jdff dff_A_KZ6waLow6_0(.din(n19948), .dout(n19951));
    jdff dff_A_KeltLhp16_0(.din(n19951), .dout(n19954));
    jdff dff_A_Wt7Ebn225_0(.din(n19954), .dout(n19957));
    jdff dff_A_mlvYLxPi1_0(.din(n19957), .dout(n19960));
    jdff dff_A_M0xobwCI7_0(.din(n19960), .dout(n19963));
    jdff dff_A_D25uNUG66_0(.din(n19963), .dout(n19966));
    jdff dff_A_Cn9l1ycb3_0(.din(n19966), .dout(n19969));
    jdff dff_A_nYnI3YW30_0(.din(n19969), .dout(n19972));
    jdff dff_A_XlR2KVD69_0(.din(n19972), .dout(n19975));
    jdff dff_A_lFNeG9137_0(.din(n19975), .dout(n19978));
    jdff dff_A_7s3CsHRd6_0(.din(n19978), .dout(n19981));
    jdff dff_A_szt6NtZ92_0(.din(n19981), .dout(n19984));
    jdff dff_A_AQOP14g49_0(.din(n19984), .dout(n19987));
    jdff dff_A_aC1yb7r84_0(.din(n19987), .dout(n19990));
    jdff dff_A_0AJZRDpq0_0(.din(n19990), .dout(n19993));
    jdff dff_A_IOWH5kqj7_0(.din(n19993), .dout(n19996));
    jdff dff_A_CuRnAuZp7_0(.din(n19996), .dout(n19999));
    jdff dff_A_O6yepDJU3_0(.din(n19999), .dout(n20002));
    jdff dff_A_lkxaeDzS6_0(.din(n20002), .dout(n20005));
    jdff dff_A_oPkwPXyi7_0(.din(n20005), .dout(n20008));
    jdff dff_A_M3HGtLT02_0(.din(n20008), .dout(n20011));
    jdff dff_A_F3Ojr0sb4_0(.din(n20011), .dout(n20014));
    jdff dff_A_7Xl7WXQP8_0(.din(n20014), .dout(n20017));
    jdff dff_A_KsFnX82u9_0(.din(n20017), .dout(n20020));
    jdff dff_A_5KInHmCx2_0(.din(n20020), .dout(n20023));
    jdff dff_A_MSMhMbcC5_0(.din(n20023), .dout(n20026));
    jdff dff_A_lEu24tQd8_0(.din(n20026), .dout(n20029));
    jdff dff_A_6FfYaLH39_0(.din(n20029), .dout(n20032));
    jdff dff_A_NT84FmHo9_0(.din(n20032), .dout(n20035));
    jdff dff_A_2fnemDXS9_0(.din(n20035), .dout(n20038));
    jdff dff_A_hADZS1ol7_0(.din(n20038), .dout(n20041));
    jdff dff_A_HFGnETG61_0(.din(n20041), .dout(n20044));
    jdff dff_A_J3VE4y9D9_0(.din(n20044), .dout(n20047));
    jdff dff_A_oSWjikhs8_0(.din(n20047), .dout(G488));
    jdff dff_A_8wLrcBEf7_1(.din(n5406), .dout(n20053));
    jdff dff_A_MBtpf6nG4_0(.din(n20053), .dout(n20056));
    jdff dff_A_zTds5Dbw1_0(.din(n20056), .dout(n20059));
    jdff dff_A_dLAi06If4_0(.din(n20059), .dout(n20062));
    jdff dff_A_i9I3egDZ9_0(.din(n20062), .dout(n20065));
    jdff dff_A_5gnGIPUa4_0(.din(n20065), .dout(n20068));
    jdff dff_A_7Nvh6Vgj4_0(.din(n20068), .dout(n20071));
    jdff dff_A_erCiyXWt7_0(.din(n20071), .dout(n20074));
    jdff dff_A_TYHneHoA3_0(.din(n20074), .dout(n20077));
    jdff dff_A_FWqguuIS8_0(.din(n20077), .dout(n20080));
    jdff dff_A_Kz9cUupp4_0(.din(n20080), .dout(n20083));
    jdff dff_A_LhcF0VFA1_0(.din(n20083), .dout(n20086));
    jdff dff_A_TWLJK79o0_0(.din(n20086), .dout(n20089));
    jdff dff_A_AhAOzCav7_0(.din(n20089), .dout(n20092));
    jdff dff_A_pJDYz61E3_0(.din(n20092), .dout(n20095));
    jdff dff_A_MgswgbaL1_0(.din(n20095), .dout(n20098));
    jdff dff_A_mBbmJr9x4_0(.din(n20098), .dout(n20101));
    jdff dff_A_mwi9elKe0_0(.din(n20101), .dout(n20104));
    jdff dff_A_8h8XM6yw7_0(.din(n20104), .dout(n20107));
    jdff dff_A_0Fb1Z5739_0(.din(n20107), .dout(n20110));
    jdff dff_A_QdUUU36t8_0(.din(n20110), .dout(n20113));
    jdff dff_A_UZ1PALCw1_0(.din(n20113), .dout(n20116));
    jdff dff_A_K0ll3kxt0_0(.din(n20116), .dout(n20119));
    jdff dff_A_tdS0yNrO9_0(.din(n20119), .dout(n20122));
    jdff dff_A_fUBM5kay7_0(.din(n20122), .dout(n20125));
    jdff dff_A_1LCeM0fm7_0(.din(n20125), .dout(n20128));
    jdff dff_A_a6FGzUCU1_0(.din(n20128), .dout(n20131));
    jdff dff_A_cDyH5COV3_0(.din(n20131), .dout(n20134));
    jdff dff_A_anFDywGS0_0(.din(n20134), .dout(n20137));
    jdff dff_A_PqpMyNmQ3_0(.din(n20137), .dout(n20140));
    jdff dff_A_NJDgWsIe4_0(.din(n20140), .dout(n20143));
    jdff dff_A_A4NiK8Pt5_0(.din(n20143), .dout(n20146));
    jdff dff_A_JZ2xUKIN3_0(.din(n20146), .dout(n20149));
    jdff dff_A_wjYWRq041_0(.din(n20149), .dout(n20152));
    jdff dff_A_RCutgdgV5_0(.din(n20152), .dout(n20155));
    jdff dff_A_RuGhyXir1_0(.din(n20155), .dout(n20158));
    jdff dff_A_MySFxhTV8_0(.din(n20158), .dout(n20161));
    jdff dff_A_es4GlcNn2_0(.din(n20161), .dout(G486));
    jdff dff_A_0XQfGMjy7_1(.din(n5409), .dout(n20167));
    jdff dff_A_GmWmMbMS4_0(.din(n20167), .dout(n20170));
    jdff dff_A_xfon8w0f5_0(.din(n20170), .dout(n20173));
    jdff dff_A_dpXPvg7D6_0(.din(n20173), .dout(n20176));
    jdff dff_A_CVj0Pjvs7_0(.din(n20176), .dout(n20179));
    jdff dff_A_qAfRDUAY1_0(.din(n20179), .dout(n20182));
    jdff dff_A_QfNvzWUm6_0(.din(n20182), .dout(n20185));
    jdff dff_A_eNVXP6yO2_0(.din(n20185), .dout(n20188));
    jdff dff_A_OLvJPhHz4_0(.din(n20188), .dout(n20191));
    jdff dff_A_hcvwTh5I5_0(.din(n20191), .dout(n20194));
    jdff dff_A_bCeKO90o8_0(.din(n20194), .dout(n20197));
    jdff dff_A_s8ITB5Uc1_0(.din(n20197), .dout(n20200));
    jdff dff_A_RjgeXgxr9_0(.din(n20200), .dout(n20203));
    jdff dff_A_u3rMyb6D9_0(.din(n20203), .dout(n20206));
    jdff dff_A_Tn0hMPUG9_0(.din(n20206), .dout(n20209));
    jdff dff_A_SWymwAb43_0(.din(n20209), .dout(n20212));
    jdff dff_A_bzW8e2QY6_0(.din(n20212), .dout(n20215));
    jdff dff_A_siXEcYW97_0(.din(n20215), .dout(n20218));
    jdff dff_A_Ecx6SjWU4_0(.din(n20218), .dout(n20221));
    jdff dff_A_VwCWuPYR3_0(.din(n20221), .dout(n20224));
    jdff dff_A_eZclCqGA6_0(.din(n20224), .dout(n20227));
    jdff dff_A_jL2jo5bH9_0(.din(n20227), .dout(n20230));
    jdff dff_A_AOQ49JsI8_0(.din(n20230), .dout(n20233));
    jdff dff_A_iZMLTyxH9_0(.din(n20233), .dout(n20236));
    jdff dff_A_oKnyiuwN2_0(.din(n20236), .dout(n20239));
    jdff dff_A_9fE7aXkZ7_0(.din(n20239), .dout(n20242));
    jdff dff_A_H9OV5D8P3_0(.din(n20242), .dout(n20245));
    jdff dff_A_tS1YKY697_0(.din(n20245), .dout(n20248));
    jdff dff_A_CDkfbcBc1_0(.din(n20248), .dout(n20251));
    jdff dff_A_b8Mrjkzo9_0(.din(n20251), .dout(n20254));
    jdff dff_A_efP6I1qo1_0(.din(n20254), .dout(n20257));
    jdff dff_A_Ty0eUYJ12_0(.din(n20257), .dout(n20260));
    jdff dff_A_xDMHUktA4_0(.din(n20260), .dout(n20263));
    jdff dff_A_mDxoQrm45_0(.din(n20263), .dout(n20266));
    jdff dff_A_uCFJA9Sx9_0(.din(n20266), .dout(n20269));
    jdff dff_A_xQXYupyA1_0(.din(n20269), .dout(n20272));
    jdff dff_A_vNexCwex3_0(.din(n20272), .dout(n20275));
    jdff dff_A_gZjphLfx4_0(.din(n20275), .dout(G484));
    jdff dff_A_azIhLlon4_1(.din(n5412), .dout(n20281));
    jdff dff_A_aX7lGb0V6_0(.din(n20281), .dout(n20284));
    jdff dff_A_BVr18Mkg6_0(.din(n20284), .dout(n20287));
    jdff dff_A_7IjS7lU89_0(.din(n20287), .dout(n20290));
    jdff dff_A_f0wHBvQ86_0(.din(n20290), .dout(n20293));
    jdff dff_A_5gzUUM279_0(.din(n20293), .dout(n20296));
    jdff dff_A_nTOv59km5_0(.din(n20296), .dout(n20299));
    jdff dff_A_O0HAABJw1_0(.din(n20299), .dout(n20302));
    jdff dff_A_aOl1XXUs2_0(.din(n20302), .dout(n20305));
    jdff dff_A_fhLYO8NA7_0(.din(n20305), .dout(n20308));
    jdff dff_A_xaMWc1gD3_0(.din(n20308), .dout(n20311));
    jdff dff_A_SyVGQfqx2_0(.din(n20311), .dout(n20314));
    jdff dff_A_19Y0Xrxv7_0(.din(n20314), .dout(n20317));
    jdff dff_A_QXfnmOgn3_0(.din(n20317), .dout(n20320));
    jdff dff_A_MDxKriLN4_0(.din(n20320), .dout(n20323));
    jdff dff_A_KwSkPwEL1_0(.din(n20323), .dout(n20326));
    jdff dff_A_fGAuh8jG0_0(.din(n20326), .dout(n20329));
    jdff dff_A_Vl3eqJhC7_0(.din(n20329), .dout(n20332));
    jdff dff_A_9JF6gBlC6_0(.din(n20332), .dout(n20335));
    jdff dff_A_3wCsGf8m6_0(.din(n20335), .dout(n20338));
    jdff dff_A_E5FGXIej3_0(.din(n20338), .dout(n20341));
    jdff dff_A_vuSVhI3f8_0(.din(n20341), .dout(n20344));
    jdff dff_A_sgL9W5m90_0(.din(n20344), .dout(n20347));
    jdff dff_A_lgmrrzQR3_0(.din(n20347), .dout(n20350));
    jdff dff_A_jvqZIyvX9_0(.din(n20350), .dout(n20353));
    jdff dff_A_92QMTkZo8_0(.din(n20353), .dout(n20356));
    jdff dff_A_DhptXEy64_0(.din(n20356), .dout(n20359));
    jdff dff_A_kbsjlWvv7_0(.din(n20359), .dout(n20362));
    jdff dff_A_xMmYfnOj8_0(.din(n20362), .dout(n20365));
    jdff dff_A_GRJr3iAi0_0(.din(n20365), .dout(n20368));
    jdff dff_A_ZWEhvrVo6_0(.din(n20368), .dout(n20371));
    jdff dff_A_UP7ljwom8_0(.din(n20371), .dout(n20374));
    jdff dff_A_uvrF2HIT8_0(.din(n20374), .dout(n20377));
    jdff dff_A_lWV9yiZL0_0(.din(n20377), .dout(n20380));
    jdff dff_A_I2oZQKlL1_0(.din(n20380), .dout(n20383));
    jdff dff_A_Z2UxhWsj7_0(.din(n20383), .dout(n20386));
    jdff dff_A_IjTnKPUP4_0(.din(n20386), .dout(n20389));
    jdff dff_A_0bdAFRdb1_0(.din(n20389), .dout(G482));
    jdff dff_A_OfRm1bFs5_1(.din(n5415), .dout(n20395));
    jdff dff_A_6KmIy3PK6_0(.din(n20395), .dout(n20398));
    jdff dff_A_aYfHaKv06_0(.din(n20398), .dout(n20401));
    jdff dff_A_ZejgaIp97_0(.din(n20401), .dout(n20404));
    jdff dff_A_yzGc5Yw31_0(.din(n20404), .dout(n20407));
    jdff dff_A_xqMcAvkU1_0(.din(n20407), .dout(n20410));
    jdff dff_A_R59MYq8p2_0(.din(n20410), .dout(n20413));
    jdff dff_A_tiPOHG574_0(.din(n20413), .dout(n20416));
    jdff dff_A_zkTwiCE67_0(.din(n20416), .dout(n20419));
    jdff dff_A_2Z5sOrnG3_0(.din(n20419), .dout(n20422));
    jdff dff_A_0g1jZ2Ei2_0(.din(n20422), .dout(n20425));
    jdff dff_A_sxPu2aiE8_0(.din(n20425), .dout(n20428));
    jdff dff_A_qXHISY2e5_0(.din(n20428), .dout(n20431));
    jdff dff_A_5V6AmOpN0_0(.din(n20431), .dout(n20434));
    jdff dff_A_IeZXgIph9_0(.din(n20434), .dout(n20437));
    jdff dff_A_6HeGVw1M1_0(.din(n20437), .dout(n20440));
    jdff dff_A_bxVfAVKx8_0(.din(n20440), .dout(n20443));
    jdff dff_A_UF25iH2F4_0(.din(n20443), .dout(n20446));
    jdff dff_A_7lydPKM67_0(.din(n20446), .dout(n20449));
    jdff dff_A_12i31rrE7_0(.din(n20449), .dout(n20452));
    jdff dff_A_aZccxvds0_0(.din(n20452), .dout(n20455));
    jdff dff_A_Jg6GTRmk2_0(.din(n20455), .dout(n20458));
    jdff dff_A_uO8ThcsR6_0(.din(n20458), .dout(n20461));
    jdff dff_A_ryiJoZyX0_0(.din(n20461), .dout(n20464));
    jdff dff_A_x43oecP31_0(.din(n20464), .dout(n20467));
    jdff dff_A_LcnKBECF8_0(.din(n20467), .dout(n20470));
    jdff dff_A_askDIDOz1_0(.din(n20470), .dout(n20473));
    jdff dff_A_yp5eiI6D2_0(.din(n20473), .dout(n20476));
    jdff dff_A_0pgN7H7a9_0(.din(n20476), .dout(n20479));
    jdff dff_A_J0Cl8Llt1_0(.din(n20479), .dout(n20482));
    jdff dff_A_MsnsuOBh0_0(.din(n20482), .dout(n20485));
    jdff dff_A_JlaKHGbb1_0(.din(n20485), .dout(n20488));
    jdff dff_A_7H0JS3R56_0(.din(n20488), .dout(n20491));
    jdff dff_A_S70F4loh0_0(.din(n20491), .dout(n20494));
    jdff dff_A_L0KI4wXP4_0(.din(n20494), .dout(n20497));
    jdff dff_A_NrQNIThS3_0(.din(n20497), .dout(n20500));
    jdff dff_A_B7IuYAhl5_0(.din(n20500), .dout(n20503));
    jdff dff_A_M8AkHDF90_0(.din(n20503), .dout(G480));
    jdff dff_A_4CAs5RJf1_1(.din(n5418), .dout(n20509));
    jdff dff_A_QMx2GvSa2_0(.din(n20509), .dout(n20512));
    jdff dff_A_pSrOzuj04_0(.din(n20512), .dout(n20515));
    jdff dff_A_w6mjS1H76_0(.din(n20515), .dout(n20518));
    jdff dff_A_KIIoL9qz8_0(.din(n20518), .dout(n20521));
    jdff dff_A_geGPXntj4_0(.din(n20521), .dout(n20524));
    jdff dff_A_8ZxDRM5e6_0(.din(n20524), .dout(n20527));
    jdff dff_A_Jn6DX5Do3_0(.din(n20527), .dout(n20530));
    jdff dff_A_Q8F5g7S29_0(.din(n20530), .dout(n20533));
    jdff dff_A_UxBbbfbk4_0(.din(n20533), .dout(n20536));
    jdff dff_A_AjFpM39c8_0(.din(n20536), .dout(n20539));
    jdff dff_A_1m3PDwZa2_0(.din(n20539), .dout(n20542));
    jdff dff_A_vmH4HACf8_0(.din(n20542), .dout(n20545));
    jdff dff_A_xwXVKDmV3_0(.din(n20545), .dout(n20548));
    jdff dff_A_eAEiSS7W8_0(.din(n20548), .dout(n20551));
    jdff dff_A_YO3aOyis2_0(.din(n20551), .dout(n20554));
    jdff dff_A_8tlymgnb3_0(.din(n20554), .dout(n20557));
    jdff dff_A_kZWwcbLK3_0(.din(n20557), .dout(n20560));
    jdff dff_A_QN2zhAZ00_0(.din(n20560), .dout(n20563));
    jdff dff_A_Iw8tVeJe3_0(.din(n20563), .dout(n20566));
    jdff dff_A_A3NyS7Sa5_0(.din(n20566), .dout(n20569));
    jdff dff_A_4b5jcwNx0_0(.din(n20569), .dout(n20572));
    jdff dff_A_sch38MpP0_0(.din(n20572), .dout(n20575));
    jdff dff_A_oTwkmGe08_0(.din(n20575), .dout(n20578));
    jdff dff_A_zgtpWmSx4_0(.din(n20578), .dout(n20581));
    jdff dff_A_4x3UBLSF8_0(.din(n20581), .dout(n20584));
    jdff dff_A_yxhFuPQj5_0(.din(n20584), .dout(n20587));
    jdff dff_A_OLMT80EA4_0(.din(n20587), .dout(n20590));
    jdff dff_A_8owFwn9k2_0(.din(n20590), .dout(n20593));
    jdff dff_A_XP7bJKId0_0(.din(n20593), .dout(n20596));
    jdff dff_A_5aZy4HNv7_0(.din(n20596), .dout(n20599));
    jdff dff_A_s5UK2fwQ1_0(.din(n20599), .dout(n20602));
    jdff dff_A_dIiYmdtN4_0(.din(n20602), .dout(n20605));
    jdff dff_A_OZgHfJat0_0(.din(n20605), .dout(n20608));
    jdff dff_A_4XJbp7bv6_0(.din(n20608), .dout(n20611));
    jdff dff_A_gPxA2HPg8_0(.din(n20611), .dout(n20614));
    jdff dff_A_pGa0lBVM3_0(.din(n20614), .dout(n20617));
    jdff dff_A_L3bN9oRH5_0(.din(n20617), .dout(G560));
    jdff dff_A_C0h2PJSo2_1(.din(n5421), .dout(n20623));
    jdff dff_A_3ZlSs3ql0_0(.din(n20623), .dout(n20626));
    jdff dff_A_u4y4jl7v3_0(.din(n20626), .dout(n20629));
    jdff dff_A_s6AQ10ey3_0(.din(n20629), .dout(n20632));
    jdff dff_A_nxrKI0JN5_0(.din(n20632), .dout(n20635));
    jdff dff_A_4ln3jjCC8_0(.din(n20635), .dout(n20638));
    jdff dff_A_5Yh2akrM3_0(.din(n20638), .dout(n20641));
    jdff dff_A_yFRi18p44_0(.din(n20641), .dout(n20644));
    jdff dff_A_oYyNcA7M6_0(.din(n20644), .dout(n20647));
    jdff dff_A_oNu8gdjv7_0(.din(n20647), .dout(n20650));
    jdff dff_A_RTGOMqj45_0(.din(n20650), .dout(n20653));
    jdff dff_A_9SOpOpus0_0(.din(n20653), .dout(n20656));
    jdff dff_A_ABGEGEJA6_0(.din(n20656), .dout(n20659));
    jdff dff_A_SIe8LqtX6_0(.din(n20659), .dout(n20662));
    jdff dff_A_iVpJPaOb8_0(.din(n20662), .dout(n20665));
    jdff dff_A_6BmYJTgU8_0(.din(n20665), .dout(n20668));
    jdff dff_A_GrpZCmGt9_0(.din(n20668), .dout(n20671));
    jdff dff_A_Ij9f2J918_0(.din(n20671), .dout(n20674));
    jdff dff_A_RLU4wszg0_0(.din(n20674), .dout(n20677));
    jdff dff_A_LgTtKnGd6_0(.din(n20677), .dout(n20680));
    jdff dff_A_6anem5Lo0_0(.din(n20680), .dout(n20683));
    jdff dff_A_we5WbZM39_0(.din(n20683), .dout(n20686));
    jdff dff_A_2CQsupRd5_0(.din(n20686), .dout(n20689));
    jdff dff_A_ps2xr9Xj4_0(.din(n20689), .dout(n20692));
    jdff dff_A_O9lqSmp91_0(.din(n20692), .dout(n20695));
    jdff dff_A_WVvNACZO4_0(.din(n20695), .dout(n20698));
    jdff dff_A_Vk368qoA7_0(.din(n20698), .dout(n20701));
    jdff dff_A_7zsfv1wu5_0(.din(n20701), .dout(n20704));
    jdff dff_A_bLGWfnQL5_0(.din(n20704), .dout(n20707));
    jdff dff_A_dAcC6USf3_0(.din(n20707), .dout(n20710));
    jdff dff_A_JIUqB4bi5_0(.din(n20710), .dout(n20713));
    jdff dff_A_vEfoIVrU5_0(.din(n20713), .dout(n20716));
    jdff dff_A_4ED88eQB2_0(.din(n20716), .dout(n20719));
    jdff dff_A_fptj2er38_0(.din(n20719), .dout(n20722));
    jdff dff_A_hPEzMaVO1_0(.din(n20722), .dout(n20725));
    jdff dff_A_TttMYAGY1_0(.din(n20725), .dout(n20728));
    jdff dff_A_0ZNHaH8t7_0(.din(n20728), .dout(n20731));
    jdff dff_A_1kvOQdXn9_0(.din(n20731), .dout(G542));
    jdff dff_A_pxhHMs847_1(.din(n5424), .dout(n20737));
    jdff dff_A_VsW5jftS6_0(.din(n20737), .dout(n20740));
    jdff dff_A_JgySY6F13_0(.din(n20740), .dout(n20743));
    jdff dff_A_9sVR3Bsm9_0(.din(n20743), .dout(n20746));
    jdff dff_A_4IHpVARz4_0(.din(n20746), .dout(n20749));
    jdff dff_A_jeD6TjU52_0(.din(n20749), .dout(n20752));
    jdff dff_A_udeU1dBJ2_0(.din(n20752), .dout(n20755));
    jdff dff_A_WadM1TZy1_0(.din(n20755), .dout(n20758));
    jdff dff_A_iG0Oa1QY8_0(.din(n20758), .dout(n20761));
    jdff dff_A_yqICLXAO0_0(.din(n20761), .dout(n20764));
    jdff dff_A_XR9DT6Ab2_0(.din(n20764), .dout(n20767));
    jdff dff_A_W7zwRZey1_0(.din(n20767), .dout(n20770));
    jdff dff_A_5CeLt9wu6_0(.din(n20770), .dout(n20773));
    jdff dff_A_zCdns82z9_0(.din(n20773), .dout(n20776));
    jdff dff_A_o19kE1385_0(.din(n20776), .dout(n20779));
    jdff dff_A_CRP9tPGI1_0(.din(n20779), .dout(n20782));
    jdff dff_A_BYt7de0p9_0(.din(n20782), .dout(n20785));
    jdff dff_A_uR1WvLjb3_0(.din(n20785), .dout(n20788));
    jdff dff_A_3dSBGSdb4_0(.din(n20788), .dout(n20791));
    jdff dff_A_PYstLBrc4_0(.din(n20791), .dout(n20794));
    jdff dff_A_qS2eEVGC4_0(.din(n20794), .dout(n20797));
    jdff dff_A_rO4RnK5C1_0(.din(n20797), .dout(n20800));
    jdff dff_A_iTjdMU746_0(.din(n20800), .dout(n20803));
    jdff dff_A_iBVr8gmg1_0(.din(n20803), .dout(n20806));
    jdff dff_A_TNdRy4995_0(.din(n20806), .dout(n20809));
    jdff dff_A_bdntXmWL8_0(.din(n20809), .dout(n20812));
    jdff dff_A_C6YvucMg7_0(.din(n20812), .dout(n20815));
    jdff dff_A_5jVqDDGp3_0(.din(n20815), .dout(n20818));
    jdff dff_A_Ofw10gvI4_0(.din(n20818), .dout(n20821));
    jdff dff_A_lYmDq50Z4_0(.din(n20821), .dout(n20824));
    jdff dff_A_hsfvckSQ1_0(.din(n20824), .dout(n20827));
    jdff dff_A_LBYiaKUj8_0(.din(n20827), .dout(n20830));
    jdff dff_A_ecvZcZ1M3_0(.din(n20830), .dout(n20833));
    jdff dff_A_cK3SquUy9_0(.din(n20833), .dout(n20836));
    jdff dff_A_AO3odD4Z5_0(.din(n20836), .dout(n20839));
    jdff dff_A_pDZLOiEj7_0(.din(n20839), .dout(n20842));
    jdff dff_A_GjZBSWIH4_0(.din(n20842), .dout(n20845));
    jdff dff_A_Im9h7vRQ0_0(.din(n20845), .dout(G558));
    jdff dff_A_PaiAskYr6_1(.din(n5427), .dout(n20851));
    jdff dff_A_PEa039RS9_0(.din(n20851), .dout(n20854));
    jdff dff_A_HjVD2Ytw1_0(.din(n20854), .dout(n20857));
    jdff dff_A_yT9STdds6_0(.din(n20857), .dout(n20860));
    jdff dff_A_RFgEf2nd3_0(.din(n20860), .dout(n20863));
    jdff dff_A_NzQEx5ya8_0(.din(n20863), .dout(n20866));
    jdff dff_A_kikej6Xq9_0(.din(n20866), .dout(n20869));
    jdff dff_A_h2d6Zx2W3_0(.din(n20869), .dout(n20872));
    jdff dff_A_LCDAcrbe1_0(.din(n20872), .dout(n20875));
    jdff dff_A_fMLPRsZ55_0(.din(n20875), .dout(n20878));
    jdff dff_A_7aDMI00h7_0(.din(n20878), .dout(n20881));
    jdff dff_A_SFh5HPZa5_0(.din(n20881), .dout(n20884));
    jdff dff_A_Mm7RvVhS7_0(.din(n20884), .dout(n20887));
    jdff dff_A_Jpov4B8I8_0(.din(n20887), .dout(n20890));
    jdff dff_A_cjL4xQIG5_0(.din(n20890), .dout(n20893));
    jdff dff_A_PSSwYHHx5_0(.din(n20893), .dout(n20896));
    jdff dff_A_2oZDLeZX0_0(.din(n20896), .dout(n20899));
    jdff dff_A_4KsZuqwr2_0(.din(n20899), .dout(n20902));
    jdff dff_A_iwURB6rR4_0(.din(n20902), .dout(n20905));
    jdff dff_A_h5hsiT301_0(.din(n20905), .dout(n20908));
    jdff dff_A_EAP9Fzxq8_0(.din(n20908), .dout(n20911));
    jdff dff_A_MTzjLy4Z3_0(.din(n20911), .dout(n20914));
    jdff dff_A_QyV2OEZm1_0(.din(n20914), .dout(n20917));
    jdff dff_A_LzccGiWz1_0(.din(n20917), .dout(n20920));
    jdff dff_A_4z79Vr0M3_0(.din(n20920), .dout(n20923));
    jdff dff_A_Mq503fkA3_0(.din(n20923), .dout(n20926));
    jdff dff_A_jZeqrxm32_0(.din(n20926), .dout(n20929));
    jdff dff_A_czPnHY5l5_0(.din(n20929), .dout(n20932));
    jdff dff_A_6O0aTqTv1_0(.din(n20932), .dout(n20935));
    jdff dff_A_pjbuSGrh8_0(.din(n20935), .dout(n20938));
    jdff dff_A_hCIu31mj5_0(.din(n20938), .dout(n20941));
    jdff dff_A_L8q86LG33_0(.din(n20941), .dout(n20944));
    jdff dff_A_lBlhLQ2q3_0(.din(n20944), .dout(n20947));
    jdff dff_A_7udL8dx51_0(.din(n20947), .dout(n20950));
    jdff dff_A_UKvZ8OJJ2_0(.din(n20950), .dout(n20953));
    jdff dff_A_XrhJPh4c1_0(.din(n20953), .dout(n20956));
    jdff dff_A_SPebHgFh5_0(.din(n20956), .dout(n20959));
    jdff dff_A_FWlxy7J35_0(.din(n20959), .dout(G556));
    jdff dff_A_Nu4uyITW4_1(.din(n5430), .dout(n20965));
    jdff dff_A_KYGZMWuo6_0(.din(n20965), .dout(n20968));
    jdff dff_A_V4M1shWF4_0(.din(n20968), .dout(n20971));
    jdff dff_A_mYA8b5aI6_0(.din(n20971), .dout(n20974));
    jdff dff_A_rOxpbbnc1_0(.din(n20974), .dout(n20977));
    jdff dff_A_uIPU12619_0(.din(n20977), .dout(n20980));
    jdff dff_A_4uOo96oq0_0(.din(n20980), .dout(n20983));
    jdff dff_A_oUpgZ5rd5_0(.din(n20983), .dout(n20986));
    jdff dff_A_yN3MoL568_0(.din(n20986), .dout(n20989));
    jdff dff_A_Szwxe2ap6_0(.din(n20989), .dout(n20992));
    jdff dff_A_pMU5co2v7_0(.din(n20992), .dout(n20995));
    jdff dff_A_XbsXp4Hc6_0(.din(n20995), .dout(n20998));
    jdff dff_A_6zhj1UlZ9_0(.din(n20998), .dout(n21001));
    jdff dff_A_PYzorhCM0_0(.din(n21001), .dout(n21004));
    jdff dff_A_IpYh18977_0(.din(n21004), .dout(n21007));
    jdff dff_A_WJTv4oxh6_0(.din(n21007), .dout(n21010));
    jdff dff_A_7zD783ES2_0(.din(n21010), .dout(n21013));
    jdff dff_A_THVfvlSd4_0(.din(n21013), .dout(n21016));
    jdff dff_A_8k2dkvxx0_0(.din(n21016), .dout(n21019));
    jdff dff_A_pVcpbkyG8_0(.din(n21019), .dout(n21022));
    jdff dff_A_jcA1LeCl9_0(.din(n21022), .dout(n21025));
    jdff dff_A_ER5x3I9I6_0(.din(n21025), .dout(n21028));
    jdff dff_A_cDRioxeM9_0(.din(n21028), .dout(n21031));
    jdff dff_A_ABZ6XXaD7_0(.din(n21031), .dout(n21034));
    jdff dff_A_gZZUu6lb2_0(.din(n21034), .dout(n21037));
    jdff dff_A_sLQNeUj59_0(.din(n21037), .dout(n21040));
    jdff dff_A_ceg1PngX7_0(.din(n21040), .dout(n21043));
    jdff dff_A_w16ZXeoN1_0(.din(n21043), .dout(n21046));
    jdff dff_A_oagw8f2y1_0(.din(n21046), .dout(n21049));
    jdff dff_A_CqzgH1EY3_0(.din(n21049), .dout(n21052));
    jdff dff_A_wrhauYB39_0(.din(n21052), .dout(n21055));
    jdff dff_A_tQKxpYIC2_0(.din(n21055), .dout(n21058));
    jdff dff_A_RzdnuyV65_0(.din(n21058), .dout(n21061));
    jdff dff_A_aH1I6zrz7_0(.din(n21061), .dout(n21064));
    jdff dff_A_TRsc783g3_0(.din(n21064), .dout(n21067));
    jdff dff_A_im4eF1Z26_0(.din(n21067), .dout(n21070));
    jdff dff_A_jd4bV5Tj0_0(.din(n21070), .dout(n21073));
    jdff dff_A_JKCsMSY77_0(.din(n21073), .dout(G554));
    jdff dff_A_Ol3YBVCw1_1(.din(n5433), .dout(n21079));
    jdff dff_A_3xSYrUPJ1_0(.din(n21079), .dout(n21082));
    jdff dff_A_SUusDXpc7_0(.din(n21082), .dout(n21085));
    jdff dff_A_UOfqOoHs5_0(.din(n21085), .dout(n21088));
    jdff dff_A_qsE9DeKb3_0(.din(n21088), .dout(n21091));
    jdff dff_A_HuUsKLXL9_0(.din(n21091), .dout(n21094));
    jdff dff_A_g31GadDR8_0(.din(n21094), .dout(n21097));
    jdff dff_A_FdiocZBN3_0(.din(n21097), .dout(n21100));
    jdff dff_A_FMYTCX8M9_0(.din(n21100), .dout(n21103));
    jdff dff_A_nF5Gf2cQ6_0(.din(n21103), .dout(n21106));
    jdff dff_A_55I86xLm8_0(.din(n21106), .dout(n21109));
    jdff dff_A_mACA9E8N1_0(.din(n21109), .dout(n21112));
    jdff dff_A_V49O5pIP8_0(.din(n21112), .dout(n21115));
    jdff dff_A_9SMjUDta9_0(.din(n21115), .dout(n21118));
    jdff dff_A_a9xdFmh85_0(.din(n21118), .dout(n21121));
    jdff dff_A_9lYXErQp7_0(.din(n21121), .dout(n21124));
    jdff dff_A_C5MZFXZ75_0(.din(n21124), .dout(n21127));
    jdff dff_A_bpCqdoll5_0(.din(n21127), .dout(n21130));
    jdff dff_A_L4yJ4DLO0_0(.din(n21130), .dout(n21133));
    jdff dff_A_QPFjJrQi9_0(.din(n21133), .dout(n21136));
    jdff dff_A_fEJvXimn8_0(.din(n21136), .dout(n21139));
    jdff dff_A_5IUykv0K0_0(.din(n21139), .dout(n21142));
    jdff dff_A_VsHqff184_0(.din(n21142), .dout(n21145));
    jdff dff_A_0UGzpnuI2_0(.din(n21145), .dout(n21148));
    jdff dff_A_zjP89fBS5_0(.din(n21148), .dout(n21151));
    jdff dff_A_6QF1TzX20_0(.din(n21151), .dout(n21154));
    jdff dff_A_jZB9fzoP3_0(.din(n21154), .dout(n21157));
    jdff dff_A_57zNAon70_0(.din(n21157), .dout(n21160));
    jdff dff_A_bwdy6hBL9_0(.din(n21160), .dout(n21163));
    jdff dff_A_MAliRglB3_0(.din(n21163), .dout(n21166));
    jdff dff_A_qiO91mHu9_0(.din(n21166), .dout(n21169));
    jdff dff_A_GFjYQP9P8_0(.din(n21169), .dout(n21172));
    jdff dff_A_8oHigkgq9_0(.din(n21172), .dout(n21175));
    jdff dff_A_B7zQoqDe2_0(.din(n21175), .dout(n21178));
    jdff dff_A_wk72eYIK2_0(.din(n21178), .dout(n21181));
    jdff dff_A_C0aK5UtC3_0(.din(n21181), .dout(n21184));
    jdff dff_A_3Ntfvrp73_0(.din(n21184), .dout(n21187));
    jdff dff_A_9BShlmBg5_0(.din(n21187), .dout(G552));
    jdff dff_A_vskJrkeb7_1(.din(n5436), .dout(n21193));
    jdff dff_A_UXRGTtyt8_0(.din(n21193), .dout(n21196));
    jdff dff_A_IkSHepBD2_0(.din(n21196), .dout(n21199));
    jdff dff_A_zFEDy7cc2_0(.din(n21199), .dout(n21202));
    jdff dff_A_rA0VUDm33_0(.din(n21202), .dout(n21205));
    jdff dff_A_xiplURXD8_0(.din(n21205), .dout(n21208));
    jdff dff_A_8mkM6KpS5_0(.din(n21208), .dout(n21211));
    jdff dff_A_PR9l0QZ11_0(.din(n21211), .dout(n21214));
    jdff dff_A_SEXLDF4N1_0(.din(n21214), .dout(n21217));
    jdff dff_A_KBiiob3w8_0(.din(n21217), .dout(n21220));
    jdff dff_A_9WPEtNDk8_0(.din(n21220), .dout(n21223));
    jdff dff_A_KJ3QnQ0p9_0(.din(n21223), .dout(n21226));
    jdff dff_A_lktW1RCq9_0(.din(n21226), .dout(n21229));
    jdff dff_A_vqgQ8fcO2_0(.din(n21229), .dout(n21232));
    jdff dff_A_3gaC2I0l1_0(.din(n21232), .dout(n21235));
    jdff dff_A_u4c3Jyrf9_0(.din(n21235), .dout(n21238));
    jdff dff_A_e5XpNalE0_0(.din(n21238), .dout(n21241));
    jdff dff_A_haPEPRUE0_0(.din(n21241), .dout(n21244));
    jdff dff_A_5836id9O3_0(.din(n21244), .dout(n21247));
    jdff dff_A_DiVwlFmt9_0(.din(n21247), .dout(n21250));
    jdff dff_A_vTIAIXSj4_0(.din(n21250), .dout(n21253));
    jdff dff_A_VPgE7vpf6_0(.din(n21253), .dout(n21256));
    jdff dff_A_AXCSkW7H8_0(.din(n21256), .dout(n21259));
    jdff dff_A_GQlxiqb36_0(.din(n21259), .dout(n21262));
    jdff dff_A_fvYAw2d11_0(.din(n21262), .dout(n21265));
    jdff dff_A_fzBALfbb9_0(.din(n21265), .dout(n21268));
    jdff dff_A_z5Ba6lRk8_0(.din(n21268), .dout(n21271));
    jdff dff_A_RwwqTgD14_0(.din(n21271), .dout(n21274));
    jdff dff_A_JSUOVrrD5_0(.din(n21274), .dout(n21277));
    jdff dff_A_P6epez6C6_0(.din(n21277), .dout(n21280));
    jdff dff_A_wp7nBcW56_0(.din(n21280), .dout(n21283));
    jdff dff_A_wKKZ6bcq6_0(.din(n21283), .dout(n21286));
    jdff dff_A_orWLLVAh9_0(.din(n21286), .dout(n21289));
    jdff dff_A_oPsjac513_0(.din(n21289), .dout(n21292));
    jdff dff_A_onglniyU2_0(.din(n21292), .dout(n21295));
    jdff dff_A_eZ0JpgUC2_0(.din(n21295), .dout(n21298));
    jdff dff_A_ZIEpFpLb1_0(.din(n21298), .dout(n21301));
    jdff dff_A_JpkdzXt20_0(.din(n21301), .dout(G550));
    jdff dff_A_RaK8syet9_1(.din(n5439), .dout(n21307));
    jdff dff_A_Pb0FOVEH6_0(.din(n21307), .dout(n21310));
    jdff dff_A_cNh3RjrQ9_0(.din(n21310), .dout(n21313));
    jdff dff_A_ubaG4VGD3_0(.din(n21313), .dout(n21316));
    jdff dff_A_L3uNG30D4_0(.din(n21316), .dout(n21319));
    jdff dff_A_IBFinrlo6_0(.din(n21319), .dout(n21322));
    jdff dff_A_CXm6vD924_0(.din(n21322), .dout(n21325));
    jdff dff_A_Ko6wFLrb9_0(.din(n21325), .dout(n21328));
    jdff dff_A_O95VmH619_0(.din(n21328), .dout(n21331));
    jdff dff_A_FuicjDch4_0(.din(n21331), .dout(n21334));
    jdff dff_A_9zh2Pvub1_0(.din(n21334), .dout(n21337));
    jdff dff_A_5B7ZAKeH5_0(.din(n21337), .dout(n21340));
    jdff dff_A_kyiH4Rgi2_0(.din(n21340), .dout(n21343));
    jdff dff_A_R6e2XuF09_0(.din(n21343), .dout(n21346));
    jdff dff_A_BaCSXDmo4_0(.din(n21346), .dout(n21349));
    jdff dff_A_xk4RxYvX4_0(.din(n21349), .dout(n21352));
    jdff dff_A_LcaHG0SP1_0(.din(n21352), .dout(n21355));
    jdff dff_A_E7OIItkO5_0(.din(n21355), .dout(n21358));
    jdff dff_A_TMCGoWJI1_0(.din(n21358), .dout(n21361));
    jdff dff_A_cRBGF4Ah5_0(.din(n21361), .dout(n21364));
    jdff dff_A_wAmiWsAq9_0(.din(n21364), .dout(n21367));
    jdff dff_A_OPHZwJFJ1_0(.din(n21367), .dout(n21370));
    jdff dff_A_2HsX3HrD8_0(.din(n21370), .dout(n21373));
    jdff dff_A_y8o5wT4a7_0(.din(n21373), .dout(n21376));
    jdff dff_A_ocYDhLiT6_0(.din(n21376), .dout(n21379));
    jdff dff_A_qdlBs3d92_0(.din(n21379), .dout(n21382));
    jdff dff_A_egPTUtCl0_0(.din(n21382), .dout(n21385));
    jdff dff_A_2qERvLwG6_0(.din(n21385), .dout(n21388));
    jdff dff_A_Rfq5qPW86_0(.din(n21388), .dout(n21391));
    jdff dff_A_PbSay1IH1_0(.din(n21391), .dout(n21394));
    jdff dff_A_YJjrWvDO5_0(.din(n21394), .dout(n21397));
    jdff dff_A_ICQVzuXr5_0(.din(n21397), .dout(n21400));
    jdff dff_A_PjGBXlrt5_0(.din(n21400), .dout(n21403));
    jdff dff_A_KEQio50c4_0(.din(n21403), .dout(n21406));
    jdff dff_A_cw6n8IGT6_0(.din(n21406), .dout(n21409));
    jdff dff_A_SOWjsBFD4_0(.din(n21409), .dout(n21412));
    jdff dff_A_e5wWdgSw4_0(.din(n21412), .dout(n21415));
    jdff dff_A_kzLLaeop0_0(.din(n21415), .dout(G548));
    jdff dff_A_rcmF46MD0_1(.din(n5442), .dout(n21421));
    jdff dff_A_TIKAjhuU9_0(.din(n21421), .dout(n21424));
    jdff dff_A_ZRN1dQRs5_0(.din(n21424), .dout(n21427));
    jdff dff_A_myDFnknc2_0(.din(n21427), .dout(n21430));
    jdff dff_A_Pr60PBI84_0(.din(n21430), .dout(n21433));
    jdff dff_A_v9xMhqA74_0(.din(n21433), .dout(n21436));
    jdff dff_A_sTaudX3u8_0(.din(n21436), .dout(n21439));
    jdff dff_A_WkRKEYxj7_0(.din(n21439), .dout(n21442));
    jdff dff_A_8p3Y9tIm7_0(.din(n21442), .dout(n21445));
    jdff dff_A_63qalUZc9_0(.din(n21445), .dout(n21448));
    jdff dff_A_Y0gpKUP46_0(.din(n21448), .dout(n21451));
    jdff dff_A_Nl6H9Dbz0_0(.din(n21451), .dout(n21454));
    jdff dff_A_VBNYUmul2_0(.din(n21454), .dout(n21457));
    jdff dff_A_OZfGCYwu9_0(.din(n21457), .dout(n21460));
    jdff dff_A_cJtEl5kD8_0(.din(n21460), .dout(n21463));
    jdff dff_A_iEHPrY3h4_0(.din(n21463), .dout(n21466));
    jdff dff_A_hmaNOJpJ2_0(.din(n21466), .dout(n21469));
    jdff dff_A_UPoEbzff2_0(.din(n21469), .dout(n21472));
    jdff dff_A_JGzFKfVt4_0(.din(n21472), .dout(n21475));
    jdff dff_A_RAiL0qDq9_0(.din(n21475), .dout(n21478));
    jdff dff_A_xq0VoqIJ2_0(.din(n21478), .dout(n21481));
    jdff dff_A_OyMd5xR60_0(.din(n21481), .dout(n21484));
    jdff dff_A_JmEGPCpi9_0(.din(n21484), .dout(n21487));
    jdff dff_A_gJSuG6s35_0(.din(n21487), .dout(n21490));
    jdff dff_A_ARddEvWE7_0(.din(n21490), .dout(n21493));
    jdff dff_A_DbDzDBwI0_0(.din(n21493), .dout(n21496));
    jdff dff_A_Lupy8mqA7_0(.din(n21496), .dout(n21499));
    jdff dff_A_0VTU5TVu6_0(.din(n21499), .dout(n21502));
    jdff dff_A_SDITtrK46_0(.din(n21502), .dout(n21505));
    jdff dff_A_FVF7AGru3_0(.din(n21505), .dout(n21508));
    jdff dff_A_ICynjAzX7_0(.din(n21508), .dout(n21511));
    jdff dff_A_66klPyMA8_0(.din(n21511), .dout(n21514));
    jdff dff_A_V3PxxPoI9_0(.din(n21514), .dout(n21517));
    jdff dff_A_1cnWBF4V9_0(.din(n21517), .dout(n21520));
    jdff dff_A_ycaRZFlL9_0(.din(n21520), .dout(n21523));
    jdff dff_A_pbDOYEnG0_0(.din(n21523), .dout(n21526));
    jdff dff_A_bX0Ptm3l1_0(.din(n21526), .dout(n21529));
    jdff dff_A_ObZeEgSA1_0(.din(n21529), .dout(G546));
    jdff dff_A_dxxPtiY89_1(.din(n5445), .dout(n21535));
    jdff dff_A_G97i5TXp7_0(.din(n21535), .dout(n21538));
    jdff dff_A_VHRF8OEO2_0(.din(n21538), .dout(n21541));
    jdff dff_A_I3eEu5BT4_0(.din(n21541), .dout(n21544));
    jdff dff_A_0ANP60F64_0(.din(n21544), .dout(n21547));
    jdff dff_A_PmBYg4Oq2_0(.din(n21547), .dout(n21550));
    jdff dff_A_XfqgMaMf9_0(.din(n21550), .dout(n21553));
    jdff dff_A_QdgbZmrm1_0(.din(n21553), .dout(n21556));
    jdff dff_A_b1Dk2QaW7_0(.din(n21556), .dout(n21559));
    jdff dff_A_yuhXJrgn8_0(.din(n21559), .dout(n21562));
    jdff dff_A_wxgERnc01_0(.din(n21562), .dout(n21565));
    jdff dff_A_T692Kb5M9_0(.din(n21565), .dout(n21568));
    jdff dff_A_E21QNLKS4_0(.din(n21568), .dout(n21571));
    jdff dff_A_W4iO5Nsn4_0(.din(n21571), .dout(n21574));
    jdff dff_A_eGycNfi15_0(.din(n21574), .dout(n21577));
    jdff dff_A_nW0dzScY3_0(.din(n21577), .dout(n21580));
    jdff dff_A_Outscrxx1_0(.din(n21580), .dout(n21583));
    jdff dff_A_VMIh675L0_0(.din(n21583), .dout(n21586));
    jdff dff_A_ORckzife0_0(.din(n21586), .dout(n21589));
    jdff dff_A_uxMBtKj98_0(.din(n21589), .dout(n21592));
    jdff dff_A_EvTsR43w5_0(.din(n21592), .dout(n21595));
    jdff dff_A_POHudtj46_0(.din(n21595), .dout(n21598));
    jdff dff_A_Cn5eg88Q0_0(.din(n21598), .dout(n21601));
    jdff dff_A_kCv8v0yV1_0(.din(n21601), .dout(n21604));
    jdff dff_A_BkYbtoU89_0(.din(n21604), .dout(n21607));
    jdff dff_A_2s01hytV1_0(.din(n21607), .dout(n21610));
    jdff dff_A_x0MQOnZ92_0(.din(n21610), .dout(n21613));
    jdff dff_A_YFmCDhea8_0(.din(n21613), .dout(n21616));
    jdff dff_A_JE7Bxocw3_0(.din(n21616), .dout(n21619));
    jdff dff_A_MSq3OtVs5_0(.din(n21619), .dout(n21622));
    jdff dff_A_LVicT9iL1_0(.din(n21622), .dout(n21625));
    jdff dff_A_yykhCNPr0_0(.din(n21625), .dout(n21628));
    jdff dff_A_kbhJRXdQ6_0(.din(n21628), .dout(n21631));
    jdff dff_A_2tqiUYdu1_0(.din(n21631), .dout(n21634));
    jdff dff_A_DKAYhMC89_0(.din(n21634), .dout(n21637));
    jdff dff_A_bjHWOuXD7_0(.din(n21637), .dout(n21640));
    jdff dff_A_RDsF7P6a8_0(.din(n21640), .dout(n21643));
    jdff dff_A_QYJkjfVl0_0(.din(n21643), .dout(G544));
    jdff dff_A_k9lEreo95_1(.din(n5448), .dout(n21649));
    jdff dff_A_0nwAKcp88_0(.din(n21649), .dout(n21652));
    jdff dff_A_jGNhNoDc3_0(.din(n21652), .dout(n21655));
    jdff dff_A_ejCxPrz08_0(.din(n21655), .dout(n21658));
    jdff dff_A_w4MTPZZ84_0(.din(n21658), .dout(n21661));
    jdff dff_A_Sgf2csNq0_0(.din(n21661), .dout(n21664));
    jdff dff_A_8cjCODhm6_0(.din(n21664), .dout(n21667));
    jdff dff_A_DreVlXB93_0(.din(n21667), .dout(n21670));
    jdff dff_A_QvaNNxVW7_0(.din(n21670), .dout(n21673));
    jdff dff_A_Eae8EmhX1_0(.din(n21673), .dout(n21676));
    jdff dff_A_KDUKBNT96_0(.din(n21676), .dout(n21679));
    jdff dff_A_CJS2jRgH4_0(.din(n21679), .dout(n21682));
    jdff dff_A_0pg6gr2N2_0(.din(n21682), .dout(n21685));
    jdff dff_A_rUgAKxQk2_0(.din(n21685), .dout(n21688));
    jdff dff_A_F62ckR6d5_0(.din(n21688), .dout(n21691));
    jdff dff_A_hqze5srK4_0(.din(n21691), .dout(n21694));
    jdff dff_A_DYinpXFB0_0(.din(n21694), .dout(n21697));
    jdff dff_A_USTYARax8_0(.din(n21697), .dout(n21700));
    jdff dff_A_weaCHrdm0_0(.din(n21700), .dout(n21703));
    jdff dff_A_lIvf3hr91_0(.din(n21703), .dout(n21706));
    jdff dff_A_uy2MvhMz9_0(.din(n21706), .dout(n21709));
    jdff dff_A_4Non3de70_0(.din(n21709), .dout(n21712));
    jdff dff_A_MPeLjYBn4_0(.din(n21712), .dout(n21715));
    jdff dff_A_VpYkl1ja7_0(.din(n21715), .dout(n21718));
    jdff dff_A_uRS1m2v22_0(.din(n21718), .dout(n21721));
    jdff dff_A_dcCxrZNW1_0(.din(n21721), .dout(n21724));
    jdff dff_A_Zx2B5KrL4_0(.din(n21724), .dout(n21727));
    jdff dff_A_qJJSCMbZ0_0(.din(n21727), .dout(n21730));
    jdff dff_A_XFyMPW0X9_0(.din(n21730), .dout(n21733));
    jdff dff_A_B7epnpWG3_0(.din(n21733), .dout(n21736));
    jdff dff_A_JUZHmBjy2_0(.din(n21736), .dout(n21739));
    jdff dff_A_VXZs3TAF0_0(.din(n21739), .dout(n21742));
    jdff dff_A_MAqTSXBt9_0(.din(n21742), .dout(n21745));
    jdff dff_A_QOjK9iD20_0(.din(n21745), .dout(n21748));
    jdff dff_A_U2EDWbT94_0(.din(n21748), .dout(n21751));
    jdff dff_A_KkTw2BSX2_0(.din(n21751), .dout(n21754));
    jdff dff_A_CP1kEolh0_0(.din(n21754), .dout(n21757));
    jdff dff_A_19ElGh7A7_0(.din(n21757), .dout(G540));
    jdff dff_A_OvoAegEm6_1(.din(n5451), .dout(n21763));
    jdff dff_A_ydkyoe2X6_0(.din(n21763), .dout(n21766));
    jdff dff_A_wh0eUoIo5_0(.din(n21766), .dout(n21769));
    jdff dff_A_7d98hpyX4_0(.din(n21769), .dout(n21772));
    jdff dff_A_rgZN6Zkb7_0(.din(n21772), .dout(n21775));
    jdff dff_A_xVug889p9_0(.din(n21775), .dout(n21778));
    jdff dff_A_ZZBzL6wA1_0(.din(n21778), .dout(n21781));
    jdff dff_A_GpDI3p6U6_0(.din(n21781), .dout(n21784));
    jdff dff_A_aVuUX56V4_0(.din(n21784), .dout(n21787));
    jdff dff_A_qwj7MtCH2_0(.din(n21787), .dout(n21790));
    jdff dff_A_X6n74ntP7_0(.din(n21790), .dout(n21793));
    jdff dff_A_M2xpWZOp0_0(.din(n21793), .dout(n21796));
    jdff dff_A_KrfvbOPY0_0(.din(n21796), .dout(n21799));
    jdff dff_A_mZ4nhya30_0(.din(n21799), .dout(n21802));
    jdff dff_A_KhIoE2iT8_0(.din(n21802), .dout(n21805));
    jdff dff_A_Ujr24iPF8_0(.din(n21805), .dout(n21808));
    jdff dff_A_B8fAShn17_0(.din(n21808), .dout(n21811));
    jdff dff_A_Ih6dd4rl0_0(.din(n21811), .dout(n21814));
    jdff dff_A_raRKZkES9_0(.din(n21814), .dout(n21817));
    jdff dff_A_yIUv6Glp2_0(.din(n21817), .dout(n21820));
    jdff dff_A_NWV0efjI5_0(.din(n21820), .dout(n21823));
    jdff dff_A_5vsPEcrY6_0(.din(n21823), .dout(n21826));
    jdff dff_A_yuhaGSUP4_0(.din(n21826), .dout(n21829));
    jdff dff_A_WbIpVahl1_0(.din(n21829), .dout(n21832));
    jdff dff_A_5nQjm3KJ8_0(.din(n21832), .dout(n21835));
    jdff dff_A_mbRarS1g5_0(.din(n21835), .dout(n21838));
    jdff dff_A_N5QgfnDu5_0(.din(n21838), .dout(n21841));
    jdff dff_A_Pb2yFNHE9_0(.din(n21841), .dout(n21844));
    jdff dff_A_Czc2e6Vp5_0(.din(n21844), .dout(n21847));
    jdff dff_A_hKmT7x8c4_0(.din(n21847), .dout(n21850));
    jdff dff_A_DDidJ2n95_0(.din(n21850), .dout(n21853));
    jdff dff_A_I59aTpTO1_0(.din(n21853), .dout(n21856));
    jdff dff_A_18OEmnbb0_0(.din(n21856), .dout(n21859));
    jdff dff_A_L3RXcbDh0_0(.din(n21859), .dout(n21862));
    jdff dff_A_4I5IVXMF3_0(.din(n21862), .dout(n21865));
    jdff dff_A_EWOwMrOK0_0(.din(n21865), .dout(n21868));
    jdff dff_A_0VpkrRIy8_0(.din(n21868), .dout(n21871));
    jdff dff_A_y10T6j0N4_0(.din(n21871), .dout(G538));
    jdff dff_A_tWFx69fK7_1(.din(n5454), .dout(n21877));
    jdff dff_A_rBXTNuUt5_0(.din(n21877), .dout(n21880));
    jdff dff_A_o1iutIEO7_0(.din(n21880), .dout(n21883));
    jdff dff_A_gOWLBNeg9_0(.din(n21883), .dout(n21886));
    jdff dff_A_UGtPa2xC2_0(.din(n21886), .dout(n21889));
    jdff dff_A_nNwuuTzu5_0(.din(n21889), .dout(n21892));
    jdff dff_A_cqqhmPMK6_0(.din(n21892), .dout(n21895));
    jdff dff_A_ikMW08vh6_0(.din(n21895), .dout(n21898));
    jdff dff_A_RU6Ktixm8_0(.din(n21898), .dout(n21901));
    jdff dff_A_RlfKC6hj9_0(.din(n21901), .dout(n21904));
    jdff dff_A_fNk6dXlS5_0(.din(n21904), .dout(n21907));
    jdff dff_A_EYhkACvk6_0(.din(n21907), .dout(n21910));
    jdff dff_A_KdJX0QZ25_0(.din(n21910), .dout(n21913));
    jdff dff_A_TV58zjAa9_0(.din(n21913), .dout(n21916));
    jdff dff_A_zBTMu70L5_0(.din(n21916), .dout(n21919));
    jdff dff_A_EsETY64J9_0(.din(n21919), .dout(n21922));
    jdff dff_A_xvGjPyfh0_0(.din(n21922), .dout(n21925));
    jdff dff_A_65jCh6314_0(.din(n21925), .dout(n21928));
    jdff dff_A_yY971RDm1_0(.din(n21928), .dout(n21931));
    jdff dff_A_wcM56EJB3_0(.din(n21931), .dout(n21934));
    jdff dff_A_tFAjRxPB6_0(.din(n21934), .dout(n21937));
    jdff dff_A_QHXXRhc95_0(.din(n21937), .dout(n21940));
    jdff dff_A_FzEdkxbu0_0(.din(n21940), .dout(n21943));
    jdff dff_A_dmwX4KAX6_0(.din(n21943), .dout(n21946));
    jdff dff_A_LZUxxINK8_0(.din(n21946), .dout(n21949));
    jdff dff_A_XqCnE4RS6_0(.din(n21949), .dout(n21952));
    jdff dff_A_234JKLKH4_0(.din(n21952), .dout(n21955));
    jdff dff_A_g1iWwlxg0_0(.din(n21955), .dout(n21958));
    jdff dff_A_OyIrr8827_0(.din(n21958), .dout(n21961));
    jdff dff_A_6vm2bBBs2_0(.din(n21961), .dout(n21964));
    jdff dff_A_W5AHB6tU7_0(.din(n21964), .dout(n21967));
    jdff dff_A_dQ0E8VZA2_0(.din(n21967), .dout(n21970));
    jdff dff_A_OTO4CLrO6_0(.din(n21970), .dout(n21973));
    jdff dff_A_hBNXpWWr1_0(.din(n21973), .dout(n21976));
    jdff dff_A_k2jTy2Qw9_0(.din(n21976), .dout(n21979));
    jdff dff_A_JtbBrwXu8_0(.din(n21979), .dout(n21982));
    jdff dff_A_PxN5ufQQ4_0(.din(n21982), .dout(n21985));
    jdff dff_A_IRFD80KQ9_0(.din(n21985), .dout(G536));
    jdff dff_A_WpSOD8rp3_1(.din(n5457), .dout(n21991));
    jdff dff_A_CdT4sQSo2_0(.din(n21991), .dout(n21994));
    jdff dff_A_HMHE3DiA7_0(.din(n21994), .dout(n21997));
    jdff dff_A_x67nYRTP7_0(.din(n21997), .dout(n22000));
    jdff dff_A_mcfY7cTk4_0(.din(n22000), .dout(n22003));
    jdff dff_A_fSiYOQJI0_0(.din(n22003), .dout(n22006));
    jdff dff_A_38EpSSyU5_0(.din(n22006), .dout(n22009));
    jdff dff_A_g6CO0Dzi9_0(.din(n22009), .dout(n22012));
    jdff dff_A_00OqCLVW3_0(.din(n22012), .dout(n22015));
    jdff dff_A_TsAWrXEj4_0(.din(n22015), .dout(n22018));
    jdff dff_A_IlTOizfN3_0(.din(n22018), .dout(n22021));
    jdff dff_A_RISActYd1_0(.din(n22021), .dout(n22024));
    jdff dff_A_H5j4OuP52_0(.din(n22024), .dout(n22027));
    jdff dff_A_adGiQ2RC5_0(.din(n22027), .dout(n22030));
    jdff dff_A_FiyPuiCJ2_0(.din(n22030), .dout(n22033));
    jdff dff_A_XFCBeme97_0(.din(n22033), .dout(n22036));
    jdff dff_A_CkcwRHEs5_0(.din(n22036), .dout(n22039));
    jdff dff_A_Tv2cXZev3_0(.din(n22039), .dout(n22042));
    jdff dff_A_J507qUcA2_0(.din(n22042), .dout(n22045));
    jdff dff_A_MEHbksYP3_0(.din(n22045), .dout(n22048));
    jdff dff_A_GjJV2pwR2_0(.din(n22048), .dout(n22051));
    jdff dff_A_a93uWquw8_0(.din(n22051), .dout(n22054));
    jdff dff_A_eYCmwouk4_0(.din(n22054), .dout(n22057));
    jdff dff_A_AFiznRLh2_0(.din(n22057), .dout(n22060));
    jdff dff_A_h5VXymDw1_0(.din(n22060), .dout(n22063));
    jdff dff_A_TZ63m7H05_0(.din(n22063), .dout(n22066));
    jdff dff_A_hrfWgdWW8_0(.din(n22066), .dout(n22069));
    jdff dff_A_UgHRdBhH4_0(.din(n22069), .dout(n22072));
    jdff dff_A_B6M3UwiU8_0(.din(n22072), .dout(n22075));
    jdff dff_A_FR305U978_0(.din(n22075), .dout(n22078));
    jdff dff_A_GWB1OvPB0_0(.din(n22078), .dout(n22081));
    jdff dff_A_1KLeYKf19_0(.din(n22081), .dout(n22084));
    jdff dff_A_pA7G6NbE5_0(.din(n22084), .dout(n22087));
    jdff dff_A_FOwIA3GO4_0(.din(n22087), .dout(n22090));
    jdff dff_A_3Lcnqqwp8_0(.din(n22090), .dout(n22093));
    jdff dff_A_qi1yUlle9_0(.din(n22093), .dout(n22096));
    jdff dff_A_g93qrmQt4_0(.din(n22096), .dout(n22099));
    jdff dff_A_lMOuGJNH0_0(.din(n22099), .dout(G534));
    jdff dff_A_0Bt12MFX2_1(.din(n5460), .dout(n22105));
    jdff dff_A_rz54Zfzl8_0(.din(n22105), .dout(n22108));
    jdff dff_A_QOlJGFcz9_0(.din(n22108), .dout(n22111));
    jdff dff_A_mMDuSWno3_0(.din(n22111), .dout(n22114));
    jdff dff_A_HKdk1ZV48_0(.din(n22114), .dout(n22117));
    jdff dff_A_u2bfEMbj0_0(.din(n22117), .dout(n22120));
    jdff dff_A_wn1z2M069_0(.din(n22120), .dout(n22123));
    jdff dff_A_BQyIudlE2_0(.din(n22123), .dout(n22126));
    jdff dff_A_UuF8KJMG0_0(.din(n22126), .dout(n22129));
    jdff dff_A_vrQXckRA3_0(.din(n22129), .dout(n22132));
    jdff dff_A_htRr66EF8_0(.din(n22132), .dout(n22135));
    jdff dff_A_tPtjB26c0_0(.din(n22135), .dout(n22138));
    jdff dff_A_A0nrnv027_0(.din(n22138), .dout(n22141));
    jdff dff_A_cBlnpneQ5_0(.din(n22141), .dout(n22144));
    jdff dff_A_sGINlGaG2_0(.din(n22144), .dout(n22147));
    jdff dff_A_9ejt6TRu9_0(.din(n22147), .dout(n22150));
    jdff dff_A_FTc2yuNf2_0(.din(n22150), .dout(n22153));
    jdff dff_A_Qo0qyAeu0_0(.din(n22153), .dout(n22156));
    jdff dff_A_GYg1aoAD3_0(.din(n22156), .dout(n22159));
    jdff dff_A_oUYbyAmX5_0(.din(n22159), .dout(n22162));
    jdff dff_A_v2oLe0R57_0(.din(n22162), .dout(n22165));
    jdff dff_A_wfmD05pD2_0(.din(n22165), .dout(n22168));
    jdff dff_A_Q70oevZG8_0(.din(n22168), .dout(n22171));
    jdff dff_A_j9sDj5rm9_0(.din(n22171), .dout(n22174));
    jdff dff_A_W7AnjYws3_0(.din(n22174), .dout(n22177));
    jdff dff_A_Y0mNZce09_0(.din(n22177), .dout(n22180));
    jdff dff_A_hQAGEpKD2_0(.din(n22180), .dout(n22183));
    jdff dff_A_vQBBfBVH8_0(.din(n22183), .dout(n22186));
    jdff dff_A_LpnxXwLD7_0(.din(n22186), .dout(n22189));
    jdff dff_A_MWFhbBBb3_0(.din(n22189), .dout(n22192));
    jdff dff_A_Ns6dSFxd8_0(.din(n22192), .dout(n22195));
    jdff dff_A_A3DMHh212_0(.din(n22195), .dout(n22198));
    jdff dff_A_Gorq8wbJ5_0(.din(n22198), .dout(n22201));
    jdff dff_A_WotqE8j32_0(.din(n22201), .dout(n22204));
    jdff dff_A_wD6MLlh62_0(.din(n22204), .dout(n22207));
    jdff dff_A_IHPxW33Q6_0(.din(n22207), .dout(n22210));
    jdff dff_A_thYjKvrw5_0(.din(n22210), .dout(n22213));
    jdff dff_A_SfYhXbFh8_0(.din(n22213), .dout(G532));
    jdff dff_A_Btoykzj63_1(.din(n5463), .dout(n22219));
    jdff dff_A_DBPTFWA46_0(.din(n22219), .dout(n22222));
    jdff dff_A_1iZsiXTt0_0(.din(n22222), .dout(n22225));
    jdff dff_A_10uOhHhX1_0(.din(n22225), .dout(n22228));
    jdff dff_A_BKq4JrHR1_0(.din(n22228), .dout(n22231));
    jdff dff_A_Ptj17vIZ4_0(.din(n22231), .dout(n22234));
    jdff dff_A_7lme9fO97_0(.din(n22234), .dout(n22237));
    jdff dff_A_6QkS7RX48_0(.din(n22237), .dout(n22240));
    jdff dff_A_GO9a7j7J8_0(.din(n22240), .dout(n22243));
    jdff dff_A_93u88cEs6_0(.din(n22243), .dout(n22246));
    jdff dff_A_05SoZ6GH4_0(.din(n22246), .dout(n22249));
    jdff dff_A_MS2eqpsR2_0(.din(n22249), .dout(n22252));
    jdff dff_A_PXDy0tFB9_0(.din(n22252), .dout(n22255));
    jdff dff_A_GvDIfDeg8_0(.din(n22255), .dout(n22258));
    jdff dff_A_BvgvXHtP6_0(.din(n22258), .dout(n22261));
    jdff dff_A_tDA1uXjO3_0(.din(n22261), .dout(n22264));
    jdff dff_A_uJD1uhaZ6_0(.din(n22264), .dout(n22267));
    jdff dff_A_l6BGa1Kh6_0(.din(n22267), .dout(n22270));
    jdff dff_A_1h69Ug5y4_0(.din(n22270), .dout(n22273));
    jdff dff_A_lGcKFsVI7_0(.din(n22273), .dout(n22276));
    jdff dff_A_gP1jGYPA2_0(.din(n22276), .dout(n22279));
    jdff dff_A_9pX1HmKe5_0(.din(n22279), .dout(n22282));
    jdff dff_A_OgPKySg30_0(.din(n22282), .dout(n22285));
    jdff dff_A_WW5Y83WK3_0(.din(n22285), .dout(n22288));
    jdff dff_A_fb7eTxiX1_0(.din(n22288), .dout(n22291));
    jdff dff_A_tuH7XCB63_0(.din(n22291), .dout(n22294));
    jdff dff_A_eJFWAKch7_0(.din(n22294), .dout(n22297));
    jdff dff_A_2cYrZ14W2_0(.din(n22297), .dout(n22300));
    jdff dff_A_Gzc1oqwx2_0(.din(n22300), .dout(n22303));
    jdff dff_A_sJdCtwPd5_0(.din(n22303), .dout(n22306));
    jdff dff_A_UkTyILvP7_0(.din(n22306), .dout(n22309));
    jdff dff_A_1WsKbfvO8_0(.din(n22309), .dout(n22312));
    jdff dff_A_cSIiDGfg7_0(.din(n22312), .dout(n22315));
    jdff dff_A_uTekU42l4_0(.din(n22315), .dout(n22318));
    jdff dff_A_lxZTtf413_0(.din(n22318), .dout(n22321));
    jdff dff_A_86D7dpH85_0(.din(n22321), .dout(n22324));
    jdff dff_A_phxFdKTc5_0(.din(n22324), .dout(n22327));
    jdff dff_A_wiS1sg8g9_0(.din(n22327), .dout(G530));
    jdff dff_A_Mp0c0e9T0_1(.din(n5466), .dout(n22333));
    jdff dff_A_QAN1kA3n9_0(.din(n22333), .dout(n22336));
    jdff dff_A_ZLWJaSWH5_0(.din(n22336), .dout(n22339));
    jdff dff_A_9iINOz5i0_0(.din(n22339), .dout(n22342));
    jdff dff_A_UHSRuxXA0_0(.din(n22342), .dout(n22345));
    jdff dff_A_bobjiQpk6_0(.din(n22345), .dout(n22348));
    jdff dff_A_06zGBEtv9_0(.din(n22348), .dout(n22351));
    jdff dff_A_zawuMBcn0_0(.din(n22351), .dout(n22354));
    jdff dff_A_LHrGMtDa1_0(.din(n22354), .dout(n22357));
    jdff dff_A_YmhHv6QF0_0(.din(n22357), .dout(n22360));
    jdff dff_A_vZ6Yf7Ir1_0(.din(n22360), .dout(n22363));
    jdff dff_A_UW4jf6w40_0(.din(n22363), .dout(n22366));
    jdff dff_A_1vubCZQV2_0(.din(n22366), .dout(n22369));
    jdff dff_A_jrvG67F59_0(.din(n22369), .dout(n22372));
    jdff dff_A_gK1eM2kv2_0(.din(n22372), .dout(n22375));
    jdff dff_A_IIAWXZjE5_0(.din(n22375), .dout(n22378));
    jdff dff_A_Cwa9wFxL1_0(.din(n22378), .dout(n22381));
    jdff dff_A_nA96BF973_0(.din(n22381), .dout(n22384));
    jdff dff_A_V3UQUgxY9_0(.din(n22384), .dout(n22387));
    jdff dff_A_E4GdjO9Q8_0(.din(n22387), .dout(n22390));
    jdff dff_A_tAHhD5eq9_0(.din(n22390), .dout(n22393));
    jdff dff_A_bHB88nvE1_0(.din(n22393), .dout(n22396));
    jdff dff_A_9XwpDm3b1_0(.din(n22396), .dout(n22399));
    jdff dff_A_kCFIHhXa8_0(.din(n22399), .dout(n22402));
    jdff dff_A_tOIP03Re8_0(.din(n22402), .dout(n22405));
    jdff dff_A_dyv9nxPW5_0(.din(n22405), .dout(n22408));
    jdff dff_A_xKrQk2kV3_0(.din(n22408), .dout(n22411));
    jdff dff_A_aa9KrGIT1_0(.din(n22411), .dout(n22414));
    jdff dff_A_kbFOTB0W7_0(.din(n22414), .dout(n22417));
    jdff dff_A_69HdGNk67_0(.din(n22417), .dout(n22420));
    jdff dff_A_1YYDhmyB3_0(.din(n22420), .dout(n22423));
    jdff dff_A_lOghKWBG3_0(.din(n22423), .dout(n22426));
    jdff dff_A_CcIk14aE8_0(.din(n22426), .dout(n22429));
    jdff dff_A_qh42paZS2_0(.din(n22429), .dout(n22432));
    jdff dff_A_9kBu6i9W7_0(.din(n22432), .dout(n22435));
    jdff dff_A_RkerbP610_0(.din(n22435), .dout(n22438));
    jdff dff_A_Pzq9DuDH9_0(.din(n22438), .dout(n22441));
    jdff dff_A_qWJuqif76_0(.din(n22441), .dout(G528));
    jdff dff_A_ReeCzHam0_1(.din(n5469), .dout(n22447));
    jdff dff_A_VAtd6ojO6_0(.din(n22447), .dout(n22450));
    jdff dff_A_fgLIz7579_0(.din(n22450), .dout(n22453));
    jdff dff_A_e6psGgm19_0(.din(n22453), .dout(n22456));
    jdff dff_A_HU1Er5R40_0(.din(n22456), .dout(n22459));
    jdff dff_A_p0ejQOe19_0(.din(n22459), .dout(n22462));
    jdff dff_A_OakH9ahz8_0(.din(n22462), .dout(n22465));
    jdff dff_A_namE0PEt9_0(.din(n22465), .dout(n22468));
    jdff dff_A_bKBHiHXY7_0(.din(n22468), .dout(n22471));
    jdff dff_A_5JS1xSX60_0(.din(n22471), .dout(n22474));
    jdff dff_A_BdGG74w49_0(.din(n22474), .dout(n22477));
    jdff dff_A_LxevbDgk3_0(.din(n22477), .dout(n22480));
    jdff dff_A_dyX5QeVm6_0(.din(n22480), .dout(n22483));
    jdff dff_A_7wrVGsvS6_0(.din(n22483), .dout(n22486));
    jdff dff_A_mdvTV2M94_0(.din(n22486), .dout(n22489));
    jdff dff_A_ZOXB797B5_0(.din(n22489), .dout(n22492));
    jdff dff_A_XqDhwwTU2_0(.din(n22492), .dout(n22495));
    jdff dff_A_FN2meJcS4_0(.din(n22495), .dout(n22498));
    jdff dff_A_UWDI1rcn2_0(.din(n22498), .dout(n22501));
    jdff dff_A_nQ5FjT9j2_0(.din(n22501), .dout(n22504));
    jdff dff_A_VMdq6R6P3_0(.din(n22504), .dout(n22507));
    jdff dff_A_UcPK5xLx8_0(.din(n22507), .dout(n22510));
    jdff dff_A_VaMgQ7rf1_0(.din(n22510), .dout(n22513));
    jdff dff_A_3KRlIzmx2_0(.din(n22513), .dout(n22516));
    jdff dff_A_1iZOStDw8_0(.din(n22516), .dout(n22519));
    jdff dff_A_WlBN6Pna2_0(.din(n22519), .dout(n22522));
    jdff dff_A_wYWfktBK4_0(.din(n22522), .dout(n22525));
    jdff dff_A_c278mtd82_0(.din(n22525), .dout(n22528));
    jdff dff_A_6Kt4kC7J3_0(.din(n22528), .dout(n22531));
    jdff dff_A_JxCayiBq8_0(.din(n22531), .dout(n22534));
    jdff dff_A_2EzZnyBp1_0(.din(n22534), .dout(n22537));
    jdff dff_A_tJsHhYII5_0(.din(n22537), .dout(n22540));
    jdff dff_A_BDPAqsf18_0(.din(n22540), .dout(n22543));
    jdff dff_A_LDtMW9hx8_0(.din(n22543), .dout(n22546));
    jdff dff_A_9K7Cq7G98_0(.din(n22546), .dout(n22549));
    jdff dff_A_vSWIXsnq3_0(.din(n22549), .dout(n22552));
    jdff dff_A_JsxhfXln5_0(.din(n22552), .dout(n22555));
    jdff dff_A_R8bl4UCH7_0(.din(n22555), .dout(G526));
    jdff dff_A_wNDkqV9X6_1(.din(n5472), .dout(n22561));
    jdff dff_A_r0WQzJi04_0(.din(n22561), .dout(n22564));
    jdff dff_A_L7TZ5b2t1_0(.din(n22564), .dout(n22567));
    jdff dff_A_S8GueEaO6_0(.din(n22567), .dout(n22570));
    jdff dff_A_d2iAScxU8_0(.din(n22570), .dout(n22573));
    jdff dff_A_PeyvzLzQ4_0(.din(n22573), .dout(n22576));
    jdff dff_A_ajzfxveW1_0(.din(n22576), .dout(n22579));
    jdff dff_A_Iy9YAmz36_0(.din(n22579), .dout(n22582));
    jdff dff_A_W35tNQns1_0(.din(n22582), .dout(n22585));
    jdff dff_A_lWT33Ufv7_0(.din(n22585), .dout(n22588));
    jdff dff_A_ScI156pN7_0(.din(n22588), .dout(n22591));
    jdff dff_A_FAqIWjmC6_0(.din(n22591), .dout(n22594));
    jdff dff_A_fyOoPG2X5_0(.din(n22594), .dout(n22597));
    jdff dff_A_3OgmrwKD1_0(.din(n22597), .dout(n22600));
    jdff dff_A_Fs0ju9HF8_0(.din(n22600), .dout(n22603));
    jdff dff_A_uCWLPIYQ2_0(.din(n22603), .dout(n22606));
    jdff dff_A_LW9T8MCW7_0(.din(n22606), .dout(n22609));
    jdff dff_A_IYKKslCv1_0(.din(n22609), .dout(n22612));
    jdff dff_A_4nNAy4ns5_0(.din(n22612), .dout(n22615));
    jdff dff_A_oCRZZGWp7_0(.din(n22615), .dout(n22618));
    jdff dff_A_XsdgfgUC7_0(.din(n22618), .dout(n22621));
    jdff dff_A_xABX73f49_0(.din(n22621), .dout(n22624));
    jdff dff_A_zyGl4EHl4_0(.din(n22624), .dout(n22627));
    jdff dff_A_e3Ydfltt6_0(.din(n22627), .dout(n22630));
    jdff dff_A_Y83BffQe9_0(.din(n22630), .dout(n22633));
    jdff dff_A_sKtdNFkT7_0(.din(n22633), .dout(n22636));
    jdff dff_A_tJtXXvJM5_0(.din(n22636), .dout(n22639));
    jdff dff_A_stbY7ACb3_0(.din(n22639), .dout(n22642));
    jdff dff_A_mHiYY7PV6_0(.din(n22642), .dout(n22645));
    jdff dff_A_pxrAQ3mi1_0(.din(n22645), .dout(n22648));
    jdff dff_A_vDJsEelS6_0(.din(n22648), .dout(n22651));
    jdff dff_A_nMMYk4NR7_0(.din(n22651), .dout(n22654));
    jdff dff_A_f6L6XOUy6_0(.din(n22654), .dout(n22657));
    jdff dff_A_7l4D5zCO0_0(.din(n22657), .dout(n22660));
    jdff dff_A_TooqVmUK2_0(.din(n22660), .dout(n22663));
    jdff dff_A_fTxHXQjX8_0(.din(n22663), .dout(n22666));
    jdff dff_A_HTCSvGZZ3_0(.din(n22666), .dout(n22669));
    jdff dff_A_4hC2oC508_0(.din(n22669), .dout(G524));
    jdff dff_A_TnC3fYtR3_1(.din(n316), .dout(n22675));
    jdff dff_A_OusjvvD54_0(.din(n22675), .dout(n22678));
    jdff dff_A_X91AlhYc5_0(.din(n22678), .dout(n22681));
    jdff dff_A_MyYDfWOG7_0(.din(n22681), .dout(n22684));
    jdff dff_A_Ugd1jy1D7_0(.din(n22684), .dout(n22687));
    jdff dff_A_DkDYaxly0_0(.din(n22687), .dout(n22690));
    jdff dff_A_CUQTXiKE8_0(.din(n22690), .dout(n22693));
    jdff dff_A_7NUqq3zw5_0(.din(n22693), .dout(n22696));
    jdff dff_A_vLtl5ggm3_0(.din(n22696), .dout(n22699));
    jdff dff_A_njdB9fOO3_0(.din(n22699), .dout(n22702));
    jdff dff_A_fCkscxnd0_0(.din(n22702), .dout(n22705));
    jdff dff_A_IqkPXJAb0_0(.din(n22705), .dout(n22708));
    jdff dff_A_er7grrb98_0(.din(n22708), .dout(n22711));
    jdff dff_A_OKNEDAyD6_0(.din(n22711), .dout(n22714));
    jdff dff_A_aaO32Qjc1_0(.din(n22714), .dout(n22717));
    jdff dff_A_j6ckGRFj5_0(.din(n22717), .dout(n22720));
    jdff dff_A_j9CNGlJS8_0(.din(n22720), .dout(n22723));
    jdff dff_A_qJBXjZCB1_0(.din(n22723), .dout(n22726));
    jdff dff_A_K2dViIzc0_0(.din(n22726), .dout(n22729));
    jdff dff_A_RxcO7qo52_0(.din(n22729), .dout(n22732));
    jdff dff_A_RUL3SLqx6_0(.din(n22732), .dout(n22735));
    jdff dff_A_DlqLsbAj3_0(.din(n22735), .dout(n22738));
    jdff dff_A_VAF0i8ZA2_0(.din(n22738), .dout(n22741));
    jdff dff_A_aWDQUBIU0_0(.din(n22741), .dout(n22744));
    jdff dff_A_ojutfHwt4_0(.din(n22744), .dout(n22747));
    jdff dff_A_mPYCv19x1_0(.din(n22747), .dout(n22750));
    jdff dff_A_8hb3iYw81_0(.din(n22750), .dout(n22753));
    jdff dff_A_3zIjocPC5_0(.din(n22753), .dout(n22756));
    jdff dff_A_PypNKC9r3_0(.din(n22756), .dout(n22759));
    jdff dff_A_xW0JxjF53_0(.din(n22759), .dout(n22762));
    jdff dff_A_4VMtYlsa4_0(.din(n22762), .dout(n22765));
    jdff dff_A_ivYYIrsJ4_0(.din(n22765), .dout(n22768));
    jdff dff_A_ftxL8Nqp4_0(.din(n22768), .dout(n22771));
    jdff dff_A_q3D0uZNR4_0(.din(n22771), .dout(n22774));
    jdff dff_A_wB1HIsRx4_0(.din(n22774), .dout(n22777));
    jdff dff_A_TqJ2Mjfy5_0(.din(n22777), .dout(n22780));
    jdff dff_A_Uj2ECwpB9_0(.din(n22780), .dout(n22783));
    jdff dff_A_Xetz9aSM4_0(.din(n22783), .dout(G279));
    jdff dff_A_3rxkWg5S9_1(.din(n5475), .dout(n22789));
    jdff dff_A_LE2rjmPW1_0(.din(n22789), .dout(n22792));
    jdff dff_A_QytUHVI58_0(.din(n22792), .dout(n22795));
    jdff dff_A_KorsMJiw9_0(.din(n22795), .dout(n22798));
    jdff dff_A_pgbKMHN99_0(.din(n22798), .dout(n22801));
    jdff dff_A_BXE8Vq7z6_0(.din(n22801), .dout(n22804));
    jdff dff_A_04mTBibP3_0(.din(n22804), .dout(n22807));
    jdff dff_A_KaB9jzjV7_0(.din(n22807), .dout(n22810));
    jdff dff_A_9pC5nFss3_0(.din(n22810), .dout(n22813));
    jdff dff_A_CwEBZBp51_0(.din(n22813), .dout(n22816));
    jdff dff_A_l9Vh7Do05_0(.din(n22816), .dout(n22819));
    jdff dff_A_vOvfAFlI4_0(.din(n22819), .dout(n22822));
    jdff dff_A_YIdbzm4r7_0(.din(n22822), .dout(n22825));
    jdff dff_A_mZUaz71h5_0(.din(n22825), .dout(n22828));
    jdff dff_A_HPPW8HyZ8_0(.din(n22828), .dout(n22831));
    jdff dff_A_wR0eZlHq0_0(.din(n22831), .dout(n22834));
    jdff dff_A_rimFFKaY6_0(.din(n22834), .dout(n22837));
    jdff dff_A_RkKW1rvY3_0(.din(n22837), .dout(n22840));
    jdff dff_A_QhWst42O8_0(.din(n22840), .dout(n22843));
    jdff dff_A_PKO1MUXk5_0(.din(n22843), .dout(n22846));
    jdff dff_A_OwNzPaYB5_0(.din(n22846), .dout(n22849));
    jdff dff_A_7UITA4t27_0(.din(n22849), .dout(n22852));
    jdff dff_A_CXJqxKHW3_0(.din(n22852), .dout(n22855));
    jdff dff_A_I73LU5FT4_0(.din(n22855), .dout(n22858));
    jdff dff_A_4ltZu5ML1_0(.din(n22858), .dout(n22861));
    jdff dff_A_9Tkyn4VC7_0(.din(n22861), .dout(n22864));
    jdff dff_A_Lg4ALZlf9_0(.din(n22864), .dout(n22867));
    jdff dff_A_hKpMjOIw7_0(.din(n22867), .dout(n22870));
    jdff dff_A_nLo2os3J5_0(.din(n22870), .dout(n22873));
    jdff dff_A_KA2T3DwW2_0(.din(n22873), .dout(n22876));
    jdff dff_A_f4BbQmFp5_0(.din(n22876), .dout(n22879));
    jdff dff_A_K06CakgD0_0(.din(n22879), .dout(n22882));
    jdff dff_A_eKKYvRWU5_0(.din(n22882), .dout(n22885));
    jdff dff_A_YHgJ9OAa6_0(.din(n22885), .dout(n22888));
    jdff dff_A_qtR2F5Pr4_0(.din(n22888), .dout(n22891));
    jdff dff_A_zKxJyPZ97_0(.din(n22891), .dout(n22894));
    jdff dff_A_xK5nuJMO5_0(.din(n22894), .dout(n22897));
    jdff dff_A_NIFIvBQ92_0(.din(n22897), .dout(G436));
    jdff dff_A_VGhsnYzH9_1(.din(n5478), .dout(n22903));
    jdff dff_A_k0kxFyxg5_0(.din(n22903), .dout(n22906));
    jdff dff_A_0Kub6lVs4_0(.din(n22906), .dout(n22909));
    jdff dff_A_vpkqxgEZ9_0(.din(n22909), .dout(n22912));
    jdff dff_A_3D01UMmf6_0(.din(n22912), .dout(n22915));
    jdff dff_A_EHtETE1Z0_0(.din(n22915), .dout(n22918));
    jdff dff_A_Pv3fbyyt1_0(.din(n22918), .dout(n22921));
    jdff dff_A_4E9fniZY7_0(.din(n22921), .dout(n22924));
    jdff dff_A_MYc4JEl05_0(.din(n22924), .dout(n22927));
    jdff dff_A_oe8rHOUi9_0(.din(n22927), .dout(n22930));
    jdff dff_A_OWaAt6vZ5_0(.din(n22930), .dout(n22933));
    jdff dff_A_jkL1XRRL0_0(.din(n22933), .dout(n22936));
    jdff dff_A_pOnNXAhg8_0(.din(n22936), .dout(n22939));
    jdff dff_A_MNOt3Rpk5_0(.din(n22939), .dout(n22942));
    jdff dff_A_8bnmCgFn2_0(.din(n22942), .dout(n22945));
    jdff dff_A_GFqcIxkx0_0(.din(n22945), .dout(n22948));
    jdff dff_A_hK3okQKZ0_0(.din(n22948), .dout(n22951));
    jdff dff_A_6zYNJLny9_0(.din(n22951), .dout(n22954));
    jdff dff_A_MEoDZomE2_0(.din(n22954), .dout(n22957));
    jdff dff_A_JnNj51JT8_0(.din(n22957), .dout(n22960));
    jdff dff_A_JprOozQS7_0(.din(n22960), .dout(n22963));
    jdff dff_A_Ip0iVPii6_0(.din(n22963), .dout(n22966));
    jdff dff_A_R0sbkSL78_0(.din(n22966), .dout(n22969));
    jdff dff_A_tllcEnYY0_0(.din(n22969), .dout(n22972));
    jdff dff_A_0tEM0fhe1_0(.din(n22972), .dout(n22975));
    jdff dff_A_SMqhLXjc6_0(.din(n22975), .dout(n22978));
    jdff dff_A_qgBiWEHo1_0(.din(n22978), .dout(n22981));
    jdff dff_A_Fp9Uf06n7_0(.din(n22981), .dout(n22984));
    jdff dff_A_nSo6I93q6_0(.din(n22984), .dout(n22987));
    jdff dff_A_acXF0J0C6_0(.din(n22987), .dout(n22990));
    jdff dff_A_VCkrEa8s3_0(.din(n22990), .dout(n22993));
    jdff dff_A_dJHNVGkm4_0(.din(n22993), .dout(n22996));
    jdff dff_A_cgUuihUD0_0(.din(n22996), .dout(n22999));
    jdff dff_A_ntG72hgR0_0(.din(n22999), .dout(n23002));
    jdff dff_A_uYXQn4582_0(.din(n23002), .dout(n23005));
    jdff dff_A_28I0bMga3_0(.din(n23005), .dout(n23008));
    jdff dff_A_FIyxzINt4_0(.din(n23008), .dout(n23011));
    jdff dff_A_dMSxsxpb2_0(.din(n23011), .dout(G478));
    jdff dff_A_JFXSKKkp5_1(.din(n5481), .dout(n23017));
    jdff dff_A_KmRG8YSZ8_0(.din(n23017), .dout(n23020));
    jdff dff_A_Hmd9HzlN3_0(.din(n23020), .dout(n23023));
    jdff dff_A_cjGxqako2_0(.din(n23023), .dout(n23026));
    jdff dff_A_tyW7NXjR8_0(.din(n23026), .dout(n23029));
    jdff dff_A_aWyQiUHD4_0(.din(n23029), .dout(n23032));
    jdff dff_A_CBYYRz818_0(.din(n23032), .dout(n23035));
    jdff dff_A_Rf3WrN775_0(.din(n23035), .dout(n23038));
    jdff dff_A_tgxb4eBv7_0(.din(n23038), .dout(n23041));
    jdff dff_A_astaUZVK0_0(.din(n23041), .dout(n23044));
    jdff dff_A_EbzHxp4j0_0(.din(n23044), .dout(n23047));
    jdff dff_A_TbGuQqq25_0(.din(n23047), .dout(n23050));
    jdff dff_A_dns6CZ698_0(.din(n23050), .dout(n23053));
    jdff dff_A_5nmK8d0p2_0(.din(n23053), .dout(n23056));
    jdff dff_A_OQJ8q4XR8_0(.din(n23056), .dout(n23059));
    jdff dff_A_AWSAZYem2_0(.din(n23059), .dout(n23062));
    jdff dff_A_k3YahAFL4_0(.din(n23062), .dout(n23065));
    jdff dff_A_56F7Au5a4_0(.din(n23065), .dout(n23068));
    jdff dff_A_zlQKHLze9_0(.din(n23068), .dout(n23071));
    jdff dff_A_kxFPVAmC5_0(.din(n23071), .dout(n23074));
    jdff dff_A_cUiNiaLE9_0(.din(n23074), .dout(n23077));
    jdff dff_A_LqlnNlhh8_0(.din(n23077), .dout(n23080));
    jdff dff_A_EoJ7s8AD2_0(.din(n23080), .dout(n23083));
    jdff dff_A_XVGMf8mF1_0(.din(n23083), .dout(n23086));
    jdff dff_A_xhiXXSCI6_0(.din(n23086), .dout(n23089));
    jdff dff_A_RsnUzjIM7_0(.din(n23089), .dout(n23092));
    jdff dff_A_nubtNemo2_0(.din(n23092), .dout(n23095));
    jdff dff_A_nEZtyRX62_0(.din(n23095), .dout(n23098));
    jdff dff_A_ME7rmiYF4_0(.din(n23098), .dout(n23101));
    jdff dff_A_Z058oID48_0(.din(n23101), .dout(n23104));
    jdff dff_A_wOc3JKWb7_0(.din(n23104), .dout(n23107));
    jdff dff_A_oIxqCI0V0_0(.din(n23107), .dout(n23110));
    jdff dff_A_i0LZDUdt2_0(.din(n23110), .dout(n23113));
    jdff dff_A_WHKvjddF5_0(.din(n23113), .dout(n23116));
    jdff dff_A_m07byV5r5_0(.din(n23116), .dout(n23119));
    jdff dff_A_0Lf6114F7_0(.din(n23119), .dout(n23122));
    jdff dff_A_MEU3uGmb7_0(.din(n23122), .dout(n23125));
    jdff dff_A_Vj3nW6U86_0(.din(n23125), .dout(G522));
    jdff dff_A_158BVJfx5_2(.din(n320), .dout(n23131));
    jdff dff_A_CLL2gg4d5_0(.din(n23131), .dout(n23134));
    jdff dff_A_9oE5xXgH8_0(.din(n23134), .dout(n23137));
    jdff dff_A_5Dm0OX310_0(.din(n23137), .dout(n23140));
    jdff dff_A_xacIzu1s5_0(.din(n23140), .dout(n23143));
    jdff dff_A_pemjsvk11_0(.din(n23143), .dout(n23146));
    jdff dff_A_VZZHPRUb7_0(.din(n23146), .dout(n23149));
    jdff dff_A_CFT6vBDo3_0(.din(n23149), .dout(n23152));
    jdff dff_A_b8zK4la92_0(.din(n23152), .dout(n23155));
    jdff dff_A_3Xb9YTFB0_0(.din(n23155), .dout(n23158));
    jdff dff_A_3sKgfhgL1_0(.din(n23158), .dout(n23161));
    jdff dff_A_miJLNjiY1_0(.din(n23161), .dout(n23164));
    jdff dff_A_Ih7lLUxj2_0(.din(n23164), .dout(n23167));
    jdff dff_A_wZ1HvS8d8_0(.din(n23167), .dout(n23170));
    jdff dff_A_8D0Z7R2P1_0(.din(n23170), .dout(n23173));
    jdff dff_A_ku5aXqcm2_0(.din(n23173), .dout(n23176));
    jdff dff_A_j4LrhcMD0_0(.din(n23176), .dout(n23179));
    jdff dff_A_RCMzzZ511_0(.din(n23179), .dout(n23182));
    jdff dff_A_ZmeHSxo71_0(.din(n23182), .dout(n23185));
    jdff dff_A_MNGIbMlA0_0(.din(n23185), .dout(n23188));
    jdff dff_A_EySmUv1b4_0(.din(n23188), .dout(n23191));
    jdff dff_A_fkQkFkf26_0(.din(n23191), .dout(n23194));
    jdff dff_A_QC3yvEuU0_0(.din(n23194), .dout(n23197));
    jdff dff_A_mOYl6UFY1_0(.din(n23197), .dout(n23200));
    jdff dff_A_nh36QvYs6_0(.din(n23200), .dout(n23203));
    jdff dff_A_etqlJ6TU7_0(.din(n23203), .dout(n23206));
    jdff dff_A_NjIgqH7Q1_0(.din(n23206), .dout(n23209));
    jdff dff_A_TGmHPZnS2_0(.din(n23209), .dout(n23212));
    jdff dff_A_EEN8P03i3_0(.din(n23212), .dout(n23215));
    jdff dff_A_rl3A3UPi4_0(.din(n23215), .dout(n23218));
    jdff dff_A_bYRWAxlR4_0(.din(n23218), .dout(n23221));
    jdff dff_A_o4VX0bgv8_0(.din(n23221), .dout(n23224));
    jdff dff_A_iRGSMRKl2_0(.din(n23224), .dout(n23227));
    jdff dff_A_Md8CSjuT2_0(.din(n23227), .dout(n23230));
    jdff dff_A_sYVzjdXt8_0(.din(n23230), .dout(n23233));
    jdff dff_A_J7k3LctK6_0(.din(n23233), .dout(n23236));
    jdff dff_A_FVVC0TFo0_0(.din(n23236), .dout(n23239));
    jdff dff_A_kWgYBNDK3_0(.din(n23239), .dout(G402));
    jdff dff_A_GynMmCSi4_1(.din(n344), .dout(n23245));
    jdff dff_A_vj1i6Q4W4_0(.din(n23245), .dout(n23248));
    jdff dff_A_9iyTVvLU4_0(.din(n23248), .dout(n23251));
    jdff dff_A_BIS7cSYb4_0(.din(n23251), .dout(n23254));
    jdff dff_A_DSrrF1LD0_0(.din(n23254), .dout(n23257));
    jdff dff_A_VIcrETCE7_0(.din(n23257), .dout(n23260));
    jdff dff_A_ZWUV3q6f1_0(.din(n23260), .dout(n23263));
    jdff dff_A_TJ3rlJPR7_0(.din(n23263), .dout(n23266));
    jdff dff_A_88fEcWo73_0(.din(n23266), .dout(n23269));
    jdff dff_A_e4qr6Kim1_0(.din(n23269), .dout(n23272));
    jdff dff_A_DIRzeKGR5_0(.din(n23272), .dout(n23275));
    jdff dff_A_qqwVFXsz4_0(.din(n23275), .dout(n23278));
    jdff dff_A_xqHEpXaw2_0(.din(n23278), .dout(n23281));
    jdff dff_A_WY0X2efS1_0(.din(n23281), .dout(n23284));
    jdff dff_A_hJ3ZGWct2_0(.din(n23284), .dout(n23287));
    jdff dff_A_nawroWYY6_0(.din(n23287), .dout(n23290));
    jdff dff_A_aTs9Zv9f3_0(.din(n23290), .dout(n23293));
    jdff dff_A_q8GdOi1s4_0(.din(n23293), .dout(n23296));
    jdff dff_A_VvfLsch44_0(.din(n23296), .dout(n23299));
    jdff dff_A_XimVxw858_0(.din(n23299), .dout(n23302));
    jdff dff_A_667T2w5h1_0(.din(n23302), .dout(n23305));
    jdff dff_A_HR4KjMBJ0_0(.din(n23305), .dout(n23308));
    jdff dff_A_0RwHo2li2_0(.din(n23308), .dout(n23311));
    jdff dff_A_JcJogVNy6_0(.din(n23311), .dout(n23314));
    jdff dff_A_YAUbcyV69_0(.din(n23314), .dout(n23317));
    jdff dff_A_Gs4iSEBu7_0(.din(n23317), .dout(n23320));
    jdff dff_A_Pkj2Y5nd5_0(.din(n23320), .dout(n23323));
    jdff dff_A_WFMLinim1_0(.din(n23323), .dout(n23326));
    jdff dff_A_RcIwekHA4_0(.din(n23326), .dout(n23329));
    jdff dff_A_0xaU0Cuh0_0(.din(n23329), .dout(n23332));
    jdff dff_A_HTAEPPW28_0(.din(n23332), .dout(n23335));
    jdff dff_A_Rdlf2Vif7_0(.din(n23335), .dout(n23338));
    jdff dff_A_PXw3ExlL2_0(.din(n23338), .dout(n23341));
    jdff dff_A_aCpWcBb56_0(.din(n23341), .dout(n23344));
    jdff dff_A_CpcPe3Hn7_0(.din(n23344), .dout(n23347));
    jdff dff_A_ao8jql5i9_0(.din(n23347), .dout(G404));
    jdff dff_A_QtSapZun2_1(.din(n368), .dout(n23353));
    jdff dff_A_Ni8tMVZk0_0(.din(n23353), .dout(n23356));
    jdff dff_A_Yr13wJqq8_0(.din(n23356), .dout(n23359));
    jdff dff_A_5HzB6MDS0_0(.din(n23359), .dout(n23362));
    jdff dff_A_Mmh4FKkW1_0(.din(n23362), .dout(n23365));
    jdff dff_A_NUUm0Deu7_0(.din(n23365), .dout(n23368));
    jdff dff_A_Eg47cOYr6_0(.din(n23368), .dout(n23371));
    jdff dff_A_DHI7KS9M8_0(.din(n23371), .dout(n23374));
    jdff dff_A_vF4yevS25_0(.din(n23374), .dout(n23377));
    jdff dff_A_a2Re9Td98_0(.din(n23377), .dout(n23380));
    jdff dff_A_rtUhi4762_0(.din(n23380), .dout(n23383));
    jdff dff_A_9rU4JBHW4_0(.din(n23383), .dout(n23386));
    jdff dff_A_EbPVg9GJ5_0(.din(n23386), .dout(n23389));
    jdff dff_A_tXaxjFRS5_0(.din(n23389), .dout(n23392));
    jdff dff_A_1etpoojM9_0(.din(n23392), .dout(n23395));
    jdff dff_A_ffGf5HGF1_0(.din(n23395), .dout(n23398));
    jdff dff_A_mdA6x57w6_0(.din(n23398), .dout(n23401));
    jdff dff_A_pM1xlMzH9_0(.din(n23401), .dout(n23404));
    jdff dff_A_BQVMZrRw0_0(.din(n23404), .dout(n23407));
    jdff dff_A_qB8ix4dM5_0(.din(n23407), .dout(n23410));
    jdff dff_A_UckGQ84b8_0(.din(n23410), .dout(n23413));
    jdff dff_A_3DyiCViY7_0(.din(n23413), .dout(n23416));
    jdff dff_A_lI64x69H9_0(.din(n23416), .dout(n23419));
    jdff dff_A_xABE00sC0_0(.din(n23419), .dout(n23422));
    jdff dff_A_9ifPF6r31_0(.din(n23422), .dout(n23425));
    jdff dff_A_aUxtXqlF6_0(.din(n23425), .dout(n23428));
    jdff dff_A_rsRX30xy1_0(.din(n23428), .dout(n23431));
    jdff dff_A_FHMB4Ax24_0(.din(n23431), .dout(n23434));
    jdff dff_A_4XAdbL8E9_0(.din(n23434), .dout(n23437));
    jdff dff_A_61Kaltr52_0(.din(n23437), .dout(n23440));
    jdff dff_A_xLSKHv535_0(.din(n23440), .dout(n23443));
    jdff dff_A_QUvfsMu10_0(.din(n23443), .dout(n23446));
    jdff dff_A_k9lcU8oD2_0(.din(n23446), .dout(n23449));
    jdff dff_A_SeTd8ZPF5_0(.din(n23449), .dout(n23452));
    jdff dff_A_G0pdch835_0(.din(n23452), .dout(n23455));
    jdff dff_A_1efeAtYx5_0(.din(n23455), .dout(G406));
    jdff dff_A_iYRibRUl1_1(.din(n392), .dout(n23461));
    jdff dff_A_DtfApZ644_0(.din(n23461), .dout(n23464));
    jdff dff_A_spBeFz7Q1_0(.din(n23464), .dout(n23467));
    jdff dff_A_zggI7YUb0_0(.din(n23467), .dout(n23470));
    jdff dff_A_uqnBezBm3_0(.din(n23470), .dout(n23473));
    jdff dff_A_4M7CeSQk3_0(.din(n23473), .dout(n23476));
    jdff dff_A_DJ6AhKP72_0(.din(n23476), .dout(n23479));
    jdff dff_A_BFztI4Bh1_0(.din(n23479), .dout(n23482));
    jdff dff_A_cqJA7KfR5_0(.din(n23482), .dout(n23485));
    jdff dff_A_zsGQi5M20_0(.din(n23485), .dout(n23488));
    jdff dff_A_UlVdO9237_0(.din(n23488), .dout(n23491));
    jdff dff_A_wUk8zebQ7_0(.din(n23491), .dout(n23494));
    jdff dff_A_pmgoKI551_0(.din(n23494), .dout(n23497));
    jdff dff_A_rM84gTKC2_0(.din(n23497), .dout(n23500));
    jdff dff_A_HrFf6mQx3_0(.din(n23500), .dout(n23503));
    jdff dff_A_YfYXewFo9_0(.din(n23503), .dout(n23506));
    jdff dff_A_r2MSjyaJ9_0(.din(n23506), .dout(n23509));
    jdff dff_A_jcBqriGy5_0(.din(n23509), .dout(n23512));
    jdff dff_A_jwfMJWPO3_0(.din(n23512), .dout(n23515));
    jdff dff_A_l0XUuEHd6_0(.din(n23515), .dout(n23518));
    jdff dff_A_TLmp5ND70_0(.din(n23518), .dout(n23521));
    jdff dff_A_CQbFnLfr6_0(.din(n23521), .dout(n23524));
    jdff dff_A_SKbKcetk1_0(.din(n23524), .dout(n23527));
    jdff dff_A_L6IqURT07_0(.din(n23527), .dout(n23530));
    jdff dff_A_1RlyPywy1_0(.din(n23530), .dout(n23533));
    jdff dff_A_YM7WnGRF9_0(.din(n23533), .dout(n23536));
    jdff dff_A_EIe6eaZE5_0(.din(n23536), .dout(n23539));
    jdff dff_A_lslajPSF1_0(.din(n23539), .dout(n23542));
    jdff dff_A_e8ZfvcSP1_0(.din(n23542), .dout(n23545));
    jdff dff_A_9SlHEK3L8_0(.din(n23545), .dout(n23548));
    jdff dff_A_CIp6Cpqx5_0(.din(n23548), .dout(n23551));
    jdff dff_A_c906w5Tr0_0(.din(n23551), .dout(n23554));
    jdff dff_A_KzHKDdGE1_0(.din(n23554), .dout(n23557));
    jdff dff_A_UBBuUfUc6_0(.din(n23557), .dout(n23560));
    jdff dff_A_6wW9gcSs6_0(.din(n23560), .dout(n23563));
    jdff dff_A_kJxTHZ8z4_0(.din(n23563), .dout(G408));
    jdff dff_A_tsINoMcR6_1(.din(n416), .dout(n23569));
    jdff dff_A_XIOyU0On8_0(.din(n23569), .dout(n23572));
    jdff dff_A_DKq3e43b4_0(.din(n23572), .dout(n23575));
    jdff dff_A_czLKlFlI1_0(.din(n23575), .dout(n23578));
    jdff dff_A_kneUDeSo9_0(.din(n23578), .dout(n23581));
    jdff dff_A_asRLFjFv8_0(.din(n23581), .dout(n23584));
    jdff dff_A_dmSL62r85_0(.din(n23584), .dout(n23587));
    jdff dff_A_WGYuRayh3_0(.din(n23587), .dout(n23590));
    jdff dff_A_t6Yo5nF36_0(.din(n23590), .dout(n23593));
    jdff dff_A_ff0bDvq20_0(.din(n23593), .dout(n23596));
    jdff dff_A_YprfJ5oT0_0(.din(n23596), .dout(n23599));
    jdff dff_A_joTFkHDa9_0(.din(n23599), .dout(n23602));
    jdff dff_A_e3zsG0NN4_0(.din(n23602), .dout(n23605));
    jdff dff_A_GiAcPx413_0(.din(n23605), .dout(n23608));
    jdff dff_A_dK4zzXzr1_0(.din(n23608), .dout(n23611));
    jdff dff_A_Ht2WsStZ1_0(.din(n23611), .dout(n23614));
    jdff dff_A_cQMboIm72_0(.din(n23614), .dout(n23617));
    jdff dff_A_8ON1Eriq9_0(.din(n23617), .dout(n23620));
    jdff dff_A_v8lLApdP1_0(.din(n23620), .dout(n23623));
    jdff dff_A_zuxOMWEg1_0(.din(n23623), .dout(n23626));
    jdff dff_A_XM4UcsAw0_0(.din(n23626), .dout(n23629));
    jdff dff_A_2hzFlrvq5_0(.din(n23629), .dout(n23632));
    jdff dff_A_MfntoeHo8_0(.din(n23632), .dout(n23635));
    jdff dff_A_sNo8GWjO7_0(.din(n23635), .dout(n23638));
    jdff dff_A_gQqToHrd4_0(.din(n23638), .dout(n23641));
    jdff dff_A_dmv0xlOx5_0(.din(n23641), .dout(n23644));
    jdff dff_A_Axk2z5rC2_0(.din(n23644), .dout(n23647));
    jdff dff_A_YnNXsQSi6_0(.din(n23647), .dout(n23650));
    jdff dff_A_HYgM8sFp3_0(.din(n23650), .dout(n23653));
    jdff dff_A_4jlBtAG66_0(.din(n23653), .dout(n23656));
    jdff dff_A_qu88kCpS4_0(.din(n23656), .dout(n23659));
    jdff dff_A_vZjIRnTp8_0(.din(n23659), .dout(n23662));
    jdff dff_A_YBpAlVzF8_0(.din(n23662), .dout(n23665));
    jdff dff_A_wUcfwBcW0_0(.din(n23665), .dout(n23668));
    jdff dff_A_97LBmKt26_0(.din(n23668), .dout(n23671));
    jdff dff_A_E8Kfagdu4_0(.din(n23671), .dout(G410));
    jdff dff_A_qBosUjhi3_1(.din(n5484), .dout(n23677));
    jdff dff_A_XmgoDoCt4_0(.din(n23677), .dout(n23680));
    jdff dff_A_itObX5ox0_0(.din(n23680), .dout(n23683));
    jdff dff_A_Rpp4e2bC3_0(.din(n23683), .dout(n23686));
    jdff dff_A_lTkrdVcb8_0(.din(n23686), .dout(n23689));
    jdff dff_A_D5p6PecJ3_0(.din(n23689), .dout(n23692));
    jdff dff_A_JXSZ5SvE0_0(.din(n23692), .dout(n23695));
    jdff dff_A_3Z2f4XkW7_0(.din(n23695), .dout(n23698));
    jdff dff_A_A9OrukCD7_0(.din(n23698), .dout(n23701));
    jdff dff_A_NAYmCd8j7_0(.din(n23701), .dout(n23704));
    jdff dff_A_xupyWn3O3_0(.din(n23704), .dout(n23707));
    jdff dff_A_H4RuCvSp8_0(.din(n23707), .dout(n23710));
    jdff dff_A_zZ1EwvVA0_0(.din(n23710), .dout(n23713));
    jdff dff_A_czCWPgKP9_0(.din(n23713), .dout(n23716));
    jdff dff_A_xNdcvHzM6_0(.din(n23716), .dout(n23719));
    jdff dff_A_j87HSMIm3_0(.din(n23719), .dout(n23722));
    jdff dff_A_GmbMW3xD9_0(.din(n23722), .dout(n23725));
    jdff dff_A_C18XUQQa7_0(.din(n23725), .dout(n23728));
    jdff dff_A_naa32m2T6_0(.din(n23728), .dout(n23731));
    jdff dff_A_cOfx9NFv1_0(.din(n23731), .dout(n23734));
    jdff dff_A_4hpYc9fY4_0(.din(n23734), .dout(n23737));
    jdff dff_A_XsJpSv5p8_0(.din(n23737), .dout(n23740));
    jdff dff_A_fqUaLZyf4_0(.din(n23740), .dout(n23743));
    jdff dff_A_8RZ7vtGk9_0(.din(n23743), .dout(n23746));
    jdff dff_A_ODlXNWHL3_0(.din(n23746), .dout(n23749));
    jdff dff_A_4swP6WIa2_0(.din(n23749), .dout(n23752));
    jdff dff_A_d6Mo7nOM4_0(.din(n23752), .dout(n23755));
    jdff dff_A_KTfYlTgG4_0(.din(n23755), .dout(n23758));
    jdff dff_A_Zyw4Hh4c6_0(.din(n23758), .dout(n23761));
    jdff dff_A_n2kFEPZK1_0(.din(n23761), .dout(n23764));
    jdff dff_A_aJ1zcPEv6_0(.din(n23764), .dout(n23767));
    jdff dff_A_6irygS6R2_0(.din(n23767), .dout(n23770));
    jdff dff_A_bolcnoIS3_0(.din(n23770), .dout(n23773));
    jdff dff_A_uSEjDQWZ8_0(.din(n23773), .dout(n23776));
    jdff dff_A_KL8TYi5m6_0(.din(n23776), .dout(n23779));
    jdff dff_A_kQwDryEX1_0(.din(n23779), .dout(n23782));
    jdff dff_A_xbTcNRte5_0(.din(n23782), .dout(n23785));
    jdff dff_A_lAwUlNW61_0(.din(n23785), .dout(G432));
    jdff dff_A_7CPkUKba1_1(.din(n5487), .dout(n23791));
    jdff dff_A_hFHRnq6W9_0(.din(n23791), .dout(n23794));
    jdff dff_A_cRkVY68A8_0(.din(n23794), .dout(n23797));
    jdff dff_A_IwjzF4j26_0(.din(n23797), .dout(n23800));
    jdff dff_A_JdS5G9fi0_0(.din(n23800), .dout(n23803));
    jdff dff_A_fOQ4OWmk6_0(.din(n23803), .dout(n23806));
    jdff dff_A_mLoOTjCq3_0(.din(n23806), .dout(n23809));
    jdff dff_A_HsuMZptG0_0(.din(n23809), .dout(n23812));
    jdff dff_A_ND3CZ08G8_0(.din(n23812), .dout(n23815));
    jdff dff_A_9BvbREtT2_0(.din(n23815), .dout(n23818));
    jdff dff_A_a4PKNzHV1_0(.din(n23818), .dout(n23821));
    jdff dff_A_5NBegsxh8_0(.din(n23821), .dout(n23824));
    jdff dff_A_dF4jaW3N3_0(.din(n23824), .dout(n23827));
    jdff dff_A_99JjSqbQ1_0(.din(n23827), .dout(n23830));
    jdff dff_A_p2BmPM2V6_0(.din(n23830), .dout(n23833));
    jdff dff_A_4ZozXwag7_0(.din(n23833), .dout(n23836));
    jdff dff_A_htkz3Bcv2_0(.din(n23836), .dout(n23839));
    jdff dff_A_btiXgu8q3_0(.din(n23839), .dout(n23842));
    jdff dff_A_FnFL6dh00_0(.din(n23842), .dout(n23845));
    jdff dff_A_afGZXWsr7_0(.din(n23845), .dout(n23848));
    jdff dff_A_v2n8Ng6n3_0(.din(n23848), .dout(n23851));
    jdff dff_A_d2BlWLgO1_0(.din(n23851), .dout(n23854));
    jdff dff_A_0Q0zobza8_0(.din(n23854), .dout(n23857));
    jdff dff_A_bgYQnZzi9_0(.din(n23857), .dout(n23860));
    jdff dff_A_5H3xuNUW5_0(.din(n23860), .dout(n23863));
    jdff dff_A_S7AHO3mo4_0(.din(n23863), .dout(n23866));
    jdff dff_A_jtWoDO2h5_0(.din(n23866), .dout(n23869));
    jdff dff_A_gBOFoBxy4_0(.din(n23869), .dout(n23872));
    jdff dff_A_RhFHycWi4_0(.din(n23872), .dout(n23875));
    jdff dff_A_DT78MEPQ2_0(.din(n23875), .dout(n23878));
    jdff dff_A_Oc6JN0xg0_0(.din(n23878), .dout(n23881));
    jdff dff_A_HdxBD7nt4_0(.din(n23881), .dout(n23884));
    jdff dff_A_bInwR5Tk5_0(.din(n23884), .dout(n23887));
    jdff dff_A_JFFF6dnL9_0(.din(n23887), .dout(n23890));
    jdff dff_A_xooZ55Ga8_0(.din(n23890), .dout(n23893));
    jdff dff_A_A4jbgDlv0_0(.din(n23893), .dout(n23896));
    jdff dff_A_GgnUw7223_0(.din(n23896), .dout(n23899));
    jdff dff_A_DK5nqAm15_0(.din(n23899), .dout(G446));
    jdff dff_A_ssThCr5Y4_2(.din(n423), .dout(n23905));
    jdff dff_A_M4P5kbJ74_0(.din(n23905), .dout(n23908));
    jdff dff_A_jl8WAa2z7_0(.din(n23908), .dout(n23911));
    jdff dff_A_5NHkHYdl1_0(.din(n23911), .dout(n23914));
    jdff dff_A_p1QNopHh9_0(.din(n23914), .dout(n23917));
    jdff dff_A_CKsYa0bN9_0(.din(n23917), .dout(n23920));
    jdff dff_A_fUcmldH32_0(.din(n23920), .dout(n23923));
    jdff dff_A_YXJAhgpv8_0(.din(n23923), .dout(n23926));
    jdff dff_A_bw2fKbEw5_0(.din(n23926), .dout(n23929));
    jdff dff_A_FJJLuoSa8_0(.din(n23929), .dout(n23932));
    jdff dff_A_o7Hz3tdQ5_0(.din(n23932), .dout(n23935));
    jdff dff_A_kzHlWNOg3_0(.din(n23935), .dout(n23938));
    jdff dff_A_PUqeC5lp1_0(.din(n23938), .dout(n23941));
    jdff dff_A_P07lZhrt0_0(.din(n23941), .dout(n23944));
    jdff dff_A_totwC3zQ5_0(.din(n23944), .dout(n23947));
    jdff dff_A_cMqDTa7Z0_0(.din(n23947), .dout(n23950));
    jdff dff_A_iBdouH5S5_0(.din(n23950), .dout(n23953));
    jdff dff_A_3VKFQcpz6_0(.din(n23953), .dout(n23956));
    jdff dff_A_T9P5G9uA4_0(.din(n23956), .dout(n23959));
    jdff dff_A_5rr3c4HZ8_0(.din(n23959), .dout(n23962));
    jdff dff_A_d8ncZiCq3_0(.din(n23962), .dout(n23965));
    jdff dff_A_KYIgKngs5_0(.din(n23965), .dout(n23968));
    jdff dff_A_qTx1po8g7_0(.din(n23968), .dout(n23971));
    jdff dff_A_0tW622NM2_0(.din(n23971), .dout(n23974));
    jdff dff_A_sdiKqK4P3_0(.din(n23974), .dout(n23977));
    jdff dff_A_gzziJXjC0_0(.din(n23977), .dout(n23980));
    jdff dff_A_USJhQbOg3_0(.din(n23980), .dout(n23983));
    jdff dff_A_LBF6doIT2_0(.din(n23983), .dout(n23986));
    jdff dff_A_fBpDS66K8_0(.din(n23986), .dout(n23989));
    jdff dff_A_icL07ajY8_0(.din(n23989), .dout(n23992));
    jdff dff_A_SS5zIw232_0(.din(n23992), .dout(n23995));
    jdff dff_A_qCEiOyxe6_0(.din(n23995), .dout(n23998));
    jdff dff_A_S4fqUD1W6_0(.din(n23998), .dout(n24001));
    jdff dff_A_VMd4BWbO7_0(.din(n24001), .dout(n24004));
    jdff dff_A_72TtIEga5_0(.din(n24004), .dout(n24007));
    jdff dff_A_GRCmtOQz2_0(.din(n24007), .dout(n24010));
    jdff dff_A_bM2a9uym8_0(.din(n24010), .dout(G284));
    jdff dff_A_2CM4RefF3_1(.din(n5490), .dout(n24016));
    jdff dff_A_n5yoZDCf8_0(.din(n24016), .dout(n24019));
    jdff dff_A_bKF5IE3v5_0(.din(n24019), .dout(n24022));
    jdff dff_A_4zRKyYlP0_0(.din(n24022), .dout(n24025));
    jdff dff_A_VWD6FnwO0_0(.din(n24025), .dout(n24028));
    jdff dff_A_c7AkPyDO7_0(.din(n24028), .dout(n24031));
    jdff dff_A_NU8Yegop7_0(.din(n24031), .dout(n24034));
    jdff dff_A_FjyWPSxX2_0(.din(n24034), .dout(n24037));
    jdff dff_A_qX7D6fDA9_0(.din(n24037), .dout(n24040));
    jdff dff_A_jiIR7V6H0_0(.din(n24040), .dout(n24043));
    jdff dff_A_u69AqvrK0_0(.din(n24043), .dout(n24046));
    jdff dff_A_TSC8EBos4_0(.din(n24046), .dout(n24049));
    jdff dff_A_TMTyYm9x4_0(.din(n24049), .dout(n24052));
    jdff dff_A_iVmQubmu0_0(.din(n24052), .dout(n24055));
    jdff dff_A_4kYU3pSG2_0(.din(n24055), .dout(n24058));
    jdff dff_A_TOO6hyuv1_0(.din(n24058), .dout(n24061));
    jdff dff_A_pqZdBcaF9_0(.din(n24061), .dout(n24064));
    jdff dff_A_Fbjf0KqF1_0(.din(n24064), .dout(n24067));
    jdff dff_A_dB48OhgZ7_0(.din(n24067), .dout(n24070));
    jdff dff_A_zCkggYEu9_0(.din(n24070), .dout(n24073));
    jdff dff_A_XrWLbXV64_0(.din(n24073), .dout(n24076));
    jdff dff_A_nDeGW0gs1_0(.din(n24076), .dout(n24079));
    jdff dff_A_AWxxHpcb5_0(.din(n24079), .dout(n24082));
    jdff dff_A_KMlUbPeh0_0(.din(n24082), .dout(n24085));
    jdff dff_A_uLqjC8R84_0(.din(n24085), .dout(n24088));
    jdff dff_A_Wiwszthh8_0(.din(n24088), .dout(n24091));
    jdff dff_A_GQtNPTjH2_0(.din(n24091), .dout(n24094));
    jdff dff_A_ul6SvONu8_0(.din(n24094), .dout(n24097));
    jdff dff_A_3C3pdOhQ0_0(.din(n24097), .dout(n24100));
    jdff dff_A_gwXh8D4n5_0(.din(n24100), .dout(n24103));
    jdff dff_A_CwSzkxRm1_0(.din(n24103), .dout(n24106));
    jdff dff_A_N1pluRYG2_0(.din(n24106), .dout(n24109));
    jdff dff_A_Xa6DPwYr3_0(.din(n24109), .dout(n24112));
    jdff dff_A_GU7r6nvd5_0(.din(n24112), .dout(n24115));
    jdff dff_A_mrVNT3gD6_0(.din(n24115), .dout(n24118));
    jdff dff_A_coFlINwc6_0(.din(n24118), .dout(n24121));
    jdff dff_A_2i4GnoHT7_0(.din(n24121), .dout(n24124));
    jdff dff_A_GEUJn6gc6_0(.din(n24124), .dout(G286));
    jdff dff_A_ZwTqURVo7_2(.din(n5494), .dout(n24130));
    jdff dff_A_plbNHkHT8_0(.din(n24130), .dout(n24133));
    jdff dff_A_62v67yL61_0(.din(n24133), .dout(n24136));
    jdff dff_A_lzLj9gwB7_0(.din(n24136), .dout(n24139));
    jdff dff_A_AMqU5Q7T1_0(.din(n24139), .dout(n24142));
    jdff dff_A_rKxjZvUk8_0(.din(n24142), .dout(n24145));
    jdff dff_A_IokWATAQ4_0(.din(n24145), .dout(n24148));
    jdff dff_A_BgZ99lLa4_0(.din(n24148), .dout(n24151));
    jdff dff_A_pJnvJxP37_0(.din(n24151), .dout(n24154));
    jdff dff_A_yxQp2DIN4_0(.din(n24154), .dout(n24157));
    jdff dff_A_ocwSjP7n9_0(.din(n24157), .dout(n24160));
    jdff dff_A_tgOR6fJn0_0(.din(n24160), .dout(n24163));
    jdff dff_A_h4ApIzZf9_0(.din(n24163), .dout(n24166));
    jdff dff_A_EKQhDHtQ6_0(.din(n24166), .dout(n24169));
    jdff dff_A_rTmEYGpL2_0(.din(n24169), .dout(n24172));
    jdff dff_A_Oh1EcsKi0_0(.din(n24172), .dout(n24175));
    jdff dff_A_QbVMJAyt6_0(.din(n24175), .dout(n24178));
    jdff dff_A_x38VK13U7_0(.din(n24178), .dout(n24181));
    jdff dff_A_Lf3y1ZlA5_0(.din(n24181), .dout(n24184));
    jdff dff_A_pkU8CXXw0_0(.din(n24184), .dout(n24187));
    jdff dff_A_yUQyUETs8_0(.din(n24187), .dout(n24190));
    jdff dff_A_kq3u3yqe7_0(.din(n24190), .dout(n24193));
    jdff dff_A_v9ZiQGw37_0(.din(n24193), .dout(n24196));
    jdff dff_A_4ryWWJ1Q2_0(.din(n24196), .dout(n24199));
    jdff dff_A_wzbqZFOy7_0(.din(n24199), .dout(n24202));
    jdff dff_A_j1ezqyNl7_0(.din(n24202), .dout(n24205));
    jdff dff_A_blHQsdka1_0(.din(n24205), .dout(n24208));
    jdff dff_A_5eU4ibM80_0(.din(n24208), .dout(n24211));
    jdff dff_A_AHgRfG8G2_0(.din(n24211), .dout(n24214));
    jdff dff_A_frXSsZH08_0(.din(n24214), .dout(n24217));
    jdff dff_A_0vJJS7Pc9_0(.din(n24217), .dout(n24220));
    jdff dff_A_EqH1qAAp1_0(.din(n24220), .dout(n24223));
    jdff dff_A_uUWmgIk26_0(.din(n24223), .dout(n24226));
    jdff dff_A_Xwr63UvT2_0(.din(n24226), .dout(n24229));
    jdff dff_A_aNtfbfzQ8_0(.din(n24229), .dout(n24232));
    jdff dff_A_n5p0vNWm1_0(.din(n24232), .dout(n24235));
    jdff dff_A_16veWjrJ2_0(.din(n24235), .dout(G289));
    jdff dff_A_x6bwFvue0_2(.din(n437), .dout(n24241));
    jdff dff_A_vJTDuolT8_0(.din(n24241), .dout(n24244));
    jdff dff_A_mVRE5PBb3_0(.din(n24244), .dout(n24247));
    jdff dff_A_j4HHhwUy1_0(.din(n24247), .dout(n24250));
    jdff dff_A_8ymnaPga4_0(.din(n24250), .dout(n24253));
    jdff dff_A_gMawEEuw6_0(.din(n24253), .dout(n24256));
    jdff dff_A_kkOSS41X7_0(.din(n24256), .dout(n24259));
    jdff dff_A_FokBI5dd4_0(.din(n24259), .dout(n24262));
    jdff dff_A_eKfA5OVK9_0(.din(n24262), .dout(n24265));
    jdff dff_A_oLhL8F5V8_0(.din(n24265), .dout(n24268));
    jdff dff_A_xm5UzF4w4_0(.din(n24268), .dout(n24271));
    jdff dff_A_xirkfDEl9_0(.din(n24271), .dout(n24274));
    jdff dff_A_VSyMBy6L9_0(.din(n24274), .dout(n24277));
    jdff dff_A_hwPy5vzu4_0(.din(n24277), .dout(n24280));
    jdff dff_A_bVZYnrVS2_0(.din(n24280), .dout(n24283));
    jdff dff_A_qKLwvFUP1_0(.din(n24283), .dout(n24286));
    jdff dff_A_PWdW3zAt4_0(.din(n24286), .dout(n24289));
    jdff dff_A_xPZrV0SC3_0(.din(n24289), .dout(n24292));
    jdff dff_A_fJaFXqRS8_0(.din(n24292), .dout(n24295));
    jdff dff_A_TPgnHYr46_0(.din(n24295), .dout(n24298));
    jdff dff_A_xAKLmj6O5_0(.din(n24298), .dout(n24301));
    jdff dff_A_QWWWZ0AH4_0(.din(n24301), .dout(n24304));
    jdff dff_A_s6o5VFmK0_0(.din(n24304), .dout(n24307));
    jdff dff_A_gXKFYeAi4_0(.din(n24307), .dout(n24310));
    jdff dff_A_KfUohfH77_0(.din(n24310), .dout(n24313));
    jdff dff_A_IxFXTg752_0(.din(n24313), .dout(n24316));
    jdff dff_A_fjgkxzkq0_0(.din(n24316), .dout(n24319));
    jdff dff_A_cR61TyC04_0(.din(n24319), .dout(n24322));
    jdff dff_A_lJS3UL8m0_0(.din(n24322), .dout(n24325));
    jdff dff_A_jzmgkfkQ5_0(.din(n24325), .dout(n24328));
    jdff dff_A_T7UAfG1r1_0(.din(n24328), .dout(n24331));
    jdff dff_A_PVcoIPhT0_0(.din(n24331), .dout(n24334));
    jdff dff_A_of390Vzo3_0(.din(n24334), .dout(n24337));
    jdff dff_A_GDUSIUm76_0(.din(n24337), .dout(n24340));
    jdff dff_A_hYnJaZzd3_0(.din(n24340), .dout(n24343));
    jdff dff_A_3SV0BPMb8_0(.din(n24343), .dout(G292));
    jdff dff_A_0w6Csyvn8_1(.din(n5497), .dout(n24349));
    jdff dff_A_aJRzz02e8_0(.din(n24349), .dout(n24352));
    jdff dff_A_ySSvZSMX1_0(.din(n24352), .dout(n24355));
    jdff dff_A_817qS1Yx7_0(.din(n24355), .dout(n24358));
    jdff dff_A_vwTRdGvn7_0(.din(n24358), .dout(n24361));
    jdff dff_A_NmgrfalF8_0(.din(n24361), .dout(n24364));
    jdff dff_A_DMZsHzAL7_0(.din(n24364), .dout(n24367));
    jdff dff_A_wcMw7NWP6_0(.din(n24367), .dout(n24370));
    jdff dff_A_3gaDqzmV2_0(.din(n24370), .dout(n24373));
    jdff dff_A_WOxNUutk7_0(.din(n24373), .dout(n24376));
    jdff dff_A_Tpyuw7Lb4_0(.din(n24376), .dout(n24379));
    jdff dff_A_vGyNWZlW9_0(.din(n24379), .dout(n24382));
    jdff dff_A_vY89ozsT9_0(.din(n24382), .dout(n24385));
    jdff dff_A_W92VnVZr5_0(.din(n24385), .dout(n24388));
    jdff dff_A_1S4h1ec35_0(.din(n24388), .dout(n24391));
    jdff dff_A_nQYf6h6r3_0(.din(n24391), .dout(n24394));
    jdff dff_A_XFgQYpmq3_0(.din(n24394), .dout(n24397));
    jdff dff_A_dTAP4cXN1_0(.din(n24397), .dout(n24400));
    jdff dff_A_vCjQO0hF3_0(.din(n24400), .dout(n24403));
    jdff dff_A_32bftMGQ8_0(.din(n24403), .dout(n24406));
    jdff dff_A_T4hKSIS77_0(.din(n24406), .dout(n24409));
    jdff dff_A_REX2j62H4_0(.din(n24409), .dout(n24412));
    jdff dff_A_Gq3lznHz2_0(.din(n24412), .dout(n24415));
    jdff dff_A_QhEIEVDd9_0(.din(n24415), .dout(n24418));
    jdff dff_A_bHzDProK3_0(.din(n24418), .dout(n24421));
    jdff dff_A_ykyFEO5f6_0(.din(n24421), .dout(n24424));
    jdff dff_A_lNTfgc6s7_0(.din(n24424), .dout(n24427));
    jdff dff_A_oOdCMo2h3_0(.din(n24427), .dout(n24430));
    jdff dff_A_ZESI0Ss79_0(.din(n24430), .dout(n24433));
    jdff dff_A_EWfjLcQY6_0(.din(n24433), .dout(n24436));
    jdff dff_A_qmZVpdSi9_0(.din(n24436), .dout(n24439));
    jdff dff_A_2vQLWaaH3_0(.din(n24439), .dout(n24442));
    jdff dff_A_03PM1Ut50_0(.din(n24442), .dout(n24445));
    jdff dff_A_UhMHdjPL6_0(.din(n24445), .dout(n24448));
    jdff dff_A_uz1hkg592_0(.din(n24448), .dout(n24451));
    jdff dff_A_cCEHWIOR6_0(.din(n24451), .dout(n24454));
    jdff dff_A_9Pj9fEaC9_0(.din(n24454), .dout(n24457));
    jdff dff_A_vT7Mf1cx5_0(.din(n24457), .dout(G341));
    jdff dff_A_UKxWtnJd8_2(.din(n5501), .dout(n24463));
    jdff dff_A_RuP9411f3_0(.din(n24463), .dout(n24466));
    jdff dff_A_ALhJE6hN7_0(.din(n24466), .dout(n24469));
    jdff dff_A_GbNS7SoF3_0(.din(n24469), .dout(n24472));
    jdff dff_A_cn5ShnvJ9_0(.din(n24472), .dout(n24475));
    jdff dff_A_qwTw1RaX2_0(.din(n24475), .dout(n24478));
    jdff dff_A_PNs8KCUb1_0(.din(n24478), .dout(n24481));
    jdff dff_A_93QzkCA82_0(.din(n24481), .dout(n24484));
    jdff dff_A_xglkL6wa8_0(.din(n24484), .dout(n24487));
    jdff dff_A_LXbpOo1Z0_0(.din(n24487), .dout(n24490));
    jdff dff_A_Xvh2uMQd3_0(.din(n24490), .dout(n24493));
    jdff dff_A_LRBna6GA3_0(.din(n24493), .dout(n24496));
    jdff dff_A_AESoj9m69_0(.din(n24496), .dout(n24499));
    jdff dff_A_SXECSwnZ7_0(.din(n24499), .dout(n24502));
    jdff dff_A_DKCrPw4f9_0(.din(n24502), .dout(n24505));
    jdff dff_A_eXmqM5jx6_0(.din(n24505), .dout(n24508));
    jdff dff_A_w4oSo3Yn8_0(.din(n24508), .dout(n24511));
    jdff dff_A_91V8v4Y38_0(.din(n24511), .dout(n24514));
    jdff dff_A_nULIvwbz1_0(.din(n24514), .dout(n24517));
    jdff dff_A_2c8d4vxf3_0(.din(n24517), .dout(n24520));
    jdff dff_A_rND2kL1W5_0(.din(n24520), .dout(n24523));
    jdff dff_A_vZpAs4mw8_0(.din(n24523), .dout(n24526));
    jdff dff_A_BZ0hxsoU0_0(.din(n24526), .dout(n24529));
    jdff dff_A_BDOGNpk46_0(.din(n24529), .dout(n24532));
    jdff dff_A_TZznJtTl5_0(.din(n24532), .dout(n24535));
    jdff dff_A_ZYFuPgoN6_0(.din(n24535), .dout(n24538));
    jdff dff_A_c1vNB3sB2_0(.din(n24538), .dout(n24541));
    jdff dff_A_tmxk6DYN5_0(.din(n24541), .dout(n24544));
    jdff dff_A_Flz6wzH57_0(.din(n24544), .dout(n24547));
    jdff dff_A_WzZOrcEQ3_0(.din(n24547), .dout(n24550));
    jdff dff_A_Pd7S7EJy4_0(.din(n24550), .dout(n24553));
    jdff dff_A_fVJNAEaJ9_0(.din(n24553), .dout(n24556));
    jdff dff_A_j7TRNiBv1_0(.din(n24556), .dout(n24559));
    jdff dff_A_jWybCdhP2_0(.din(n24559), .dout(n24562));
    jdff dff_A_RWyN0RFi0_0(.din(n24562), .dout(n24565));
    jdff dff_A_jQgGwhbs3_0(.din(n24565), .dout(G281));
    jdff dff_A_M0HT7wKV8_1(.din(n5504), .dout(n24571));
    jdff dff_A_XEH1iaR35_0(.din(n24571), .dout(n24574));
    jdff dff_A_CqiTVAVZ2_0(.din(n24574), .dout(n24577));
    jdff dff_A_bsfuE8Sl1_0(.din(n24577), .dout(n24580));
    jdff dff_A_zWxyzn3l5_0(.din(n24580), .dout(n24583));
    jdff dff_A_WzuUtemE3_0(.din(n24583), .dout(n24586));
    jdff dff_A_paBSIU5t2_0(.din(n24586), .dout(n24589));
    jdff dff_A_nu7sBOC97_0(.din(n24589), .dout(n24592));
    jdff dff_A_HzvtWlB31_0(.din(n24592), .dout(n24595));
    jdff dff_A_kuGB9u1T4_0(.din(n24595), .dout(n24598));
    jdff dff_A_q0C6jZsZ7_0(.din(n24598), .dout(n24601));
    jdff dff_A_ATNOlEmw6_0(.din(n24601), .dout(n24604));
    jdff dff_A_l78yR6Lg3_0(.din(n24604), .dout(n24607));
    jdff dff_A_WeboNXlf9_0(.din(n24607), .dout(n24610));
    jdff dff_A_6Xgt1Nuk4_0(.din(n24610), .dout(n24613));
    jdff dff_A_BxZix9QQ3_0(.din(n24613), .dout(n24616));
    jdff dff_A_FwZWJJCL2_0(.din(n24616), .dout(n24619));
    jdff dff_A_lID18ov26_0(.din(n24619), .dout(n24622));
    jdff dff_A_AjzjY1pl6_0(.din(n24622), .dout(n24625));
    jdff dff_A_oNu8Qi0D7_0(.din(n24625), .dout(n24628));
    jdff dff_A_aZE4mLlt9_0(.din(n24628), .dout(n24631));
    jdff dff_A_bZMU7YKQ7_0(.din(n24631), .dout(n24634));
    jdff dff_A_RR9XyXBC3_0(.din(n24634), .dout(n24637));
    jdff dff_A_wrF4K1iO4_0(.din(n24637), .dout(n24640));
    jdff dff_A_x9NQhUqe8_0(.din(n24640), .dout(n24643));
    jdff dff_A_gOZDgZ043_0(.din(n24643), .dout(n24646));
    jdff dff_A_ZjsyHjk21_0(.din(n24646), .dout(n24649));
    jdff dff_A_S0Qy6RCn4_0(.din(n24649), .dout(n24652));
    jdff dff_A_d9rpGd3U9_0(.din(n24652), .dout(n24655));
    jdff dff_A_BUfKz0sK4_0(.din(n24655), .dout(n24658));
    jdff dff_A_xK4mRano6_0(.din(n24658), .dout(n24661));
    jdff dff_A_2RJVWX3P4_0(.din(n24661), .dout(n24664));
    jdff dff_A_KniBZR9T5_0(.din(n24664), .dout(n24667));
    jdff dff_A_sAHh03771_0(.din(n24667), .dout(n24670));
    jdff dff_A_iQckNP664_0(.din(n24670), .dout(n24673));
    jdff dff_A_v3a1Duhj4_0(.din(n24673), .dout(n24676));
    jdff dff_A_KWBqBybj2_0(.din(n24676), .dout(n24679));
    jdff dff_A_vcCgEMvk3_0(.din(n24679), .dout(G453));
    jdff dff_A_EbglPHaX6_2(.din(n441), .dout(n24685));
    jdff dff_A_swV84blL3_0(.din(n24685), .dout(n24688));
    jdff dff_A_MoTpyETq4_0(.din(n24688), .dout(n24691));
    jdff dff_A_befxaSdt5_0(.din(n24691), .dout(n24694));
    jdff dff_A_nj1S3wB41_0(.din(n24694), .dout(n24697));
    jdff dff_A_7C4MqCvJ4_0(.din(n24697), .dout(n24700));
    jdff dff_A_NJpT3PZq6_0(.din(n24700), .dout(n24703));
    jdff dff_A_rUUp3FX02_0(.din(n24703), .dout(n24706));
    jdff dff_A_fSutrgXe6_0(.din(n24706), .dout(n24709));
    jdff dff_A_VgcIlFzG8_0(.din(n24709), .dout(n24712));
    jdff dff_A_69izWaog9_0(.din(n24712), .dout(n24715));
    jdff dff_A_Cdzp4wZp7_0(.din(n24715), .dout(n24718));
    jdff dff_A_virqKLAN5_0(.din(n24718), .dout(n24721));
    jdff dff_A_5ENM3xos9_0(.din(n24721), .dout(n24724));
    jdff dff_A_V2tqs1vF0_0(.din(n24724), .dout(n24727));
    jdff dff_A_wk30Ygv81_0(.din(n24727), .dout(n24730));
    jdff dff_A_110pMlfj1_0(.din(n24730), .dout(n24733));
    jdff dff_A_hWdkipOI8_0(.din(n24733), .dout(n24736));
    jdff dff_A_GQm3qUCT1_0(.din(n24736), .dout(n24739));
    jdff dff_A_iIUXtAtb7_0(.din(n24739), .dout(n24742));
    jdff dff_A_ZsJAKTfe5_0(.din(n24742), .dout(n24745));
    jdff dff_A_qXeYCbkh8_0(.din(n24745), .dout(n24748));
    jdff dff_A_RFNpAnF93_0(.din(n24748), .dout(n24751));
    jdff dff_A_EjXHQbSF4_0(.din(n24751), .dout(n24754));
    jdff dff_A_40eeJVPZ1_0(.din(n24754), .dout(n24757));
    jdff dff_A_5QtKENZk9_0(.din(n24757), .dout(n24760));
    jdff dff_A_wkcGo9BV7_0(.din(n24760), .dout(n24763));
    jdff dff_A_Oit6hlsp3_0(.din(n24763), .dout(n24766));
    jdff dff_A_RmnDTltQ2_0(.din(n24766), .dout(n24769));
    jdff dff_A_EtNNyMz02_0(.din(n24769), .dout(n24772));
    jdff dff_A_rIrObztX0_0(.din(n24772), .dout(n24775));
    jdff dff_A_9dE3pU650_0(.din(n24775), .dout(n24778));
    jdff dff_A_6L9Z9La10_0(.din(n24778), .dout(n24781));
    jdff dff_A_rfwuTdbL8_0(.din(n24781), .dout(n24784));
    jdff dff_A_XcD2rOzf0_0(.din(n24784), .dout(n24787));
    jdff dff_A_siWTAYaz3_0(.din(n24787), .dout(n24790));
    jdff dff_A_POP02OC74_0(.din(n24790), .dout(n24793));
    jdff dff_A_rz4eBgoh6_0(.din(n24793), .dout(G278));
    jdff dff_A_S8QuRzkE0_2(.din(n474), .dout(n24799));
    jdff dff_A_dseyb2v74_0(.din(n24799), .dout(n24802));
    jdff dff_A_OUFirTFu9_0(.din(n24802), .dout(n24805));
    jdff dff_A_0TFd1sSJ4_0(.din(n24805), .dout(n24808));
    jdff dff_A_kXRCpNYU6_0(.din(n24808), .dout(n24811));
    jdff dff_A_YUdKZbFq6_0(.din(n24811), .dout(n24814));
    jdff dff_A_W5OsBaa58_0(.din(n24814), .dout(n24817));
    jdff dff_A_uu9vKEwQ8_0(.din(n24817), .dout(n24820));
    jdff dff_A_FMlwMk116_0(.din(n24820), .dout(n24823));
    jdff dff_A_XAK0UxfS4_0(.din(n24823), .dout(n24826));
    jdff dff_A_fvgllW6Q1_0(.din(n24826), .dout(n24829));
    jdff dff_A_XCi5mrWq6_0(.din(n24829), .dout(n24832));
    jdff dff_A_vMeoGz8n2_0(.din(n24832), .dout(n24835));
    jdff dff_A_0Bdpm1em9_0(.din(n24835), .dout(n24838));
    jdff dff_A_3nVUNd1z4_0(.din(n24838), .dout(n24841));
    jdff dff_A_q6yS1vd01_0(.din(n24841), .dout(n24844));
    jdff dff_A_VeUuPMa17_0(.din(n24844), .dout(n24847));
    jdff dff_A_XNT9SGAd2_0(.din(n24847), .dout(n24850));
    jdff dff_A_x7xCGkqj3_0(.din(n24850), .dout(n24853));
    jdff dff_A_T0wCi8o12_0(.din(n24853), .dout(n24856));
    jdff dff_A_Cely64dP6_0(.din(n24856), .dout(n24859));
    jdff dff_A_nrExZfeL0_0(.din(n24859), .dout(n24862));
    jdff dff_A_rQYLfaUN2_0(.din(n24862), .dout(n24865));
    jdff dff_A_12TaG0F05_0(.din(n24865), .dout(n24868));
endmodule

