/*
gf_sqrt:
	jxor: 3736
	jspl: 4699
	jspl3: 8046
	jnot: 4189
	jand: 8731
	jor: 8388

Summary:
	jxor: 3736
	jspl: 4699
	jspl3: 8046
	jnot: 4189
	jand: 8731
	jor: 8388

The maximum logic level gap of any gate:
	gf_sqrt: 2
*/

module gf_sqrt(gclk, a, asqrt);
	input gclk;
	input [127:0] a;
	output [63:0] asqrt;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n276;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n333;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n342;
	wire n343;
	wire n345;
	wire n346;
	wire n347;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1038;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1328;
	wire n1329;
	wire n1330;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1667;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1673;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1684;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1690;
	wire n1691;
	wire n1692;
	wire n1693;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1707;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire n1718;
	wire n1719;
	wire n1720;
	wire n1721;
	wire n1722;
	wire n1723;
	wire n1724;
	wire n1725;
	wire n1726;
	wire n1727;
	wire n1728;
	wire n1729;
	wire n1730;
	wire n1731;
	wire n1732;
	wire n1733;
	wire n1734;
	wire n1735;
	wire n1736;
	wire n1737;
	wire n1738;
	wire n1739;
	wire n1740;
	wire n1741;
	wire n1742;
	wire n1743;
	wire n1744;
	wire n1745;
	wire n1746;
	wire n1747;
	wire n1748;
	wire n1749;
	wire n1750;
	wire n1751;
	wire n1752;
	wire n1753;
	wire n1754;
	wire n1755;
	wire n1756;
	wire n1757;
	wire n1758;
	wire n1759;
	wire n1760;
	wire n1761;
	wire n1762;
	wire n1763;
	wire n1764;
	wire n1765;
	wire n1766;
	wire n1767;
	wire n1768;
	wire n1769;
	wire n1770;
	wire n1771;
	wire n1772;
	wire n1773;
	wire n1774;
	wire n1775;
	wire n1776;
	wire n1777;
	wire n1778;
	wire n1779;
	wire n1780;
	wire n1781;
	wire n1782;
	wire n1783;
	wire n1784;
	wire n1785;
	wire n1786;
	wire n1787;
	wire n1788;
	wire n1789;
	wire n1790;
	wire n1791;
	wire n1792;
	wire n1793;
	wire n1794;
	wire n1795;
	wire n1796;
	wire n1797;
	wire n1798;
	wire n1799;
	wire n1800;
	wire n1801;
	wire n1802;
	wire n1803;
	wire n1804;
	wire n1805;
	wire n1806;
	wire n1807;
	wire n1808;
	wire n1809;
	wire n1810;
	wire n1811;
	wire n1812;
	wire n1813;
	wire n1814;
	wire n1815;
	wire n1816;
	wire n1817;
	wire n1818;
	wire n1819;
	wire n1821;
	wire n1822;
	wire n1823;
	wire n1824;
	wire n1825;
	wire n1826;
	wire n1827;
	wire n1828;
	wire n1829;
	wire n1830;
	wire n1831;
	wire n1832;
	wire n1833;
	wire n1834;
	wire n1835;
	wire n1836;
	wire n1837;
	wire n1838;
	wire n1839;
	wire n1840;
	wire n1841;
	wire n1842;
	wire n1843;
	wire n1844;
	wire n1845;
	wire n1846;
	wire n1847;
	wire n1848;
	wire n1849;
	wire n1850;
	wire n1851;
	wire n1852;
	wire n1853;
	wire n1854;
	wire n1855;
	wire n1856;
	wire n1857;
	wire n1858;
	wire n1859;
	wire n1860;
	wire n1861;
	wire n1862;
	wire n1863;
	wire n1864;
	wire n1865;
	wire n1866;
	wire n1867;
	wire n1868;
	wire n1869;
	wire n1870;
	wire n1871;
	wire n1872;
	wire n1873;
	wire n1874;
	wire n1875;
	wire n1876;
	wire n1877;
	wire n1878;
	wire n1879;
	wire n1880;
	wire n1881;
	wire n1882;
	wire n1883;
	wire n1884;
	wire n1885;
	wire n1886;
	wire n1887;
	wire n1888;
	wire n1889;
	wire n1890;
	wire n1891;
	wire n1892;
	wire n1893;
	wire n1894;
	wire n1895;
	wire n1896;
	wire n1897;
	wire n1898;
	wire n1899;
	wire n1900;
	wire n1901;
	wire n1902;
	wire n1903;
	wire n1904;
	wire n1905;
	wire n1906;
	wire n1907;
	wire n1908;
	wire n1909;
	wire n1910;
	wire n1911;
	wire n1912;
	wire n1913;
	wire n1914;
	wire n1915;
	wire n1916;
	wire n1917;
	wire n1918;
	wire n1919;
	wire n1920;
	wire n1921;
	wire n1922;
	wire n1923;
	wire n1924;
	wire n1925;
	wire n1926;
	wire n1927;
	wire n1928;
	wire n1929;
	wire n1930;
	wire n1931;
	wire n1932;
	wire n1933;
	wire n1934;
	wire n1935;
	wire n1936;
	wire n1937;
	wire n1938;
	wire n1939;
	wire n1940;
	wire n1941;
	wire n1942;
	wire n1943;
	wire n1944;
	wire n1945;
	wire n1946;
	wire n1947;
	wire n1948;
	wire n1949;
	wire n1950;
	wire n1951;
	wire n1952;
	wire n1953;
	wire n1954;
	wire n1955;
	wire n1956;
	wire n1957;
	wire n1958;
	wire n1959;
	wire n1960;
	wire n1961;
	wire n1962;
	wire n1963;
	wire n1964;
	wire n1965;
	wire n1966;
	wire n1967;
	wire n1968;
	wire n1969;
	wire n1970;
	wire n1971;
	wire n1972;
	wire n1973;
	wire n1974;
	wire n1975;
	wire n1976;
	wire n1977;
	wire n1978;
	wire n1979;
	wire n1980;
	wire n1981;
	wire n1982;
	wire n1983;
	wire n1984;
	wire n1985;
	wire n1986;
	wire n1987;
	wire n1988;
	wire n1989;
	wire n1990;
	wire n1991;
	wire n1992;
	wire n1993;
	wire n1994;
	wire n1995;
	wire n1996;
	wire n1997;
	wire n1998;
	wire n1999;
	wire n2000;
	wire n2001;
	wire n2002;
	wire n2003;
	wire n2004;
	wire n2005;
	wire n2006;
	wire n2007;
	wire n2008;
	wire n2009;
	wire n2010;
	wire n2011;
	wire n2012;
	wire n2013;
	wire n2014;
	wire n2015;
	wire n2016;
	wire n2017;
	wire n2018;
	wire n2019;
	wire n2020;
	wire n2021;
	wire n2022;
	wire n2023;
	wire n2024;
	wire n2025;
	wire n2026;
	wire n2027;
	wire n2028;
	wire n2029;
	wire n2030;
	wire n2031;
	wire n2032;
	wire n2033;
	wire n2034;
	wire n2035;
	wire n2036;
	wire n2037;
	wire n2038;
	wire n2039;
	wire n2040;
	wire n2041;
	wire n2042;
	wire n2043;
	wire n2044;
	wire n2045;
	wire n2046;
	wire n2047;
	wire n2048;
	wire n2049;
	wire n2050;
	wire n2051;
	wire n2052;
	wire n2053;
	wire n2054;
	wire n2055;
	wire n2056;
	wire n2057;
	wire n2058;
	wire n2059;
	wire n2060;
	wire n2061;
	wire n2062;
	wire n2063;
	wire n2064;
	wire n2065;
	wire n2066;
	wire n2067;
	wire n2068;
	wire n2069;
	wire n2070;
	wire n2071;
	wire n2072;
	wire n2073;
	wire n2074;
	wire n2075;
	wire n2076;
	wire n2077;
	wire n2078;
	wire n2079;
	wire n2080;
	wire n2081;
	wire n2082;
	wire n2083;
	wire n2084;
	wire n2085;
	wire n2086;
	wire n2087;
	wire n2088;
	wire n2089;
	wire n2090;
	wire n2091;
	wire n2092;
	wire n2093;
	wire n2094;
	wire n2095;
	wire n2096;
	wire n2097;
	wire n2098;
	wire n2099;
	wire n2100;
	wire n2101;
	wire n2103;
	wire n2104;
	wire n2105;
	wire n2106;
	wire n2107;
	wire n2108;
	wire n2109;
	wire n2110;
	wire n2111;
	wire n2112;
	wire n2113;
	wire n2114;
	wire n2115;
	wire n2116;
	wire n2117;
	wire n2118;
	wire n2119;
	wire n2120;
	wire n2121;
	wire n2122;
	wire n2123;
	wire n2124;
	wire n2125;
	wire n2126;
	wire n2127;
	wire n2128;
	wire n2129;
	wire n2130;
	wire n2131;
	wire n2132;
	wire n2133;
	wire n2134;
	wire n2135;
	wire n2136;
	wire n2137;
	wire n2138;
	wire n2139;
	wire n2140;
	wire n2141;
	wire n2142;
	wire n2143;
	wire n2144;
	wire n2145;
	wire n2146;
	wire n2147;
	wire n2148;
	wire n2149;
	wire n2150;
	wire n2151;
	wire n2152;
	wire n2153;
	wire n2154;
	wire n2155;
	wire n2156;
	wire n2157;
	wire n2158;
	wire n2159;
	wire n2160;
	wire n2161;
	wire n2162;
	wire n2163;
	wire n2164;
	wire n2165;
	wire n2166;
	wire n2167;
	wire n2168;
	wire n2169;
	wire n2170;
	wire n2171;
	wire n2172;
	wire n2173;
	wire n2174;
	wire n2175;
	wire n2176;
	wire n2177;
	wire n2178;
	wire n2179;
	wire n2180;
	wire n2181;
	wire n2182;
	wire n2183;
	wire n2184;
	wire n2185;
	wire n2186;
	wire n2187;
	wire n2188;
	wire n2189;
	wire n2190;
	wire n2191;
	wire n2192;
	wire n2193;
	wire n2194;
	wire n2195;
	wire n2196;
	wire n2197;
	wire n2198;
	wire n2199;
	wire n2200;
	wire n2201;
	wire n2202;
	wire n2203;
	wire n2204;
	wire n2205;
	wire n2206;
	wire n2207;
	wire n2208;
	wire n2209;
	wire n2210;
	wire n2211;
	wire n2212;
	wire n2213;
	wire n2214;
	wire n2215;
	wire n2216;
	wire n2217;
	wire n2218;
	wire n2219;
	wire n2220;
	wire n2221;
	wire n2222;
	wire n2223;
	wire n2224;
	wire n2225;
	wire n2226;
	wire n2227;
	wire n2228;
	wire n2229;
	wire n2230;
	wire n2231;
	wire n2232;
	wire n2233;
	wire n2234;
	wire n2235;
	wire n2236;
	wire n2238;
	wire n2239;
	wire n2240;
	wire n2241;
	wire n2242;
	wire n2243;
	wire n2244;
	wire n2245;
	wire n2246;
	wire n2247;
	wire n2248;
	wire n2249;
	wire n2252;
	wire n2253;
	wire n2254;
	wire n2255;
	wire n2256;
	wire n2257;
	wire n2258;
	wire n2259;
	wire n2260;
	wire n2261;
	wire n2262;
	wire n2263;
	wire n2265;
	wire n2266;
	wire n2267;
	wire n2268;
	wire n2269;
	wire n2270;
	wire n2271;
	wire n2272;
	wire n2273;
	wire n2274;
	wire n2275;
	wire n2276;
	wire n2277;
	wire n2278;
	wire n2279;
	wire n2280;
	wire n2281;
	wire n2282;
	wire n2283;
	wire n2284;
	wire n2285;
	wire n2286;
	wire n2287;
	wire n2288;
	wire n2289;
	wire n2290;
	wire n2291;
	wire n2292;
	wire n2293;
	wire n2294;
	wire n2295;
	wire n2296;
	wire n2297;
	wire n2298;
	wire n2299;
	wire n2300;
	wire n2301;
	wire n2302;
	wire n2303;
	wire n2304;
	wire n2305;
	wire n2306;
	wire n2307;
	wire n2308;
	wire n2309;
	wire n2310;
	wire n2311;
	wire n2312;
	wire n2313;
	wire n2314;
	wire n2315;
	wire n2316;
	wire n2317;
	wire n2318;
	wire n2319;
	wire n2320;
	wire n2321;
	wire n2322;
	wire n2323;
	wire n2324;
	wire n2325;
	wire n2326;
	wire n2327;
	wire n2328;
	wire n2329;
	wire n2330;
	wire n2331;
	wire n2332;
	wire n2333;
	wire n2334;
	wire n2335;
	wire n2336;
	wire n2337;
	wire n2338;
	wire n2339;
	wire n2340;
	wire n2341;
	wire n2342;
	wire n2343;
	wire n2345;
	wire n2346;
	wire n2347;
	wire n2348;
	wire n2349;
	wire n2350;
	wire n2351;
	wire n2352;
	wire n2353;
	wire n2354;
	wire n2355;
	wire n2356;
	wire n2357;
	wire n2358;
	wire n2359;
	wire n2360;
	wire n2361;
	wire n2362;
	wire n2363;
	wire n2364;
	wire n2365;
	wire n2366;
	wire n2367;
	wire n2368;
	wire n2369;
	wire n2370;
	wire n2371;
	wire n2372;
	wire n2373;
	wire n2374;
	wire n2375;
	wire n2376;
	wire n2377;
	wire n2378;
	wire n2379;
	wire n2380;
	wire n2381;
	wire n2382;
	wire n2383;
	wire n2384;
	wire n2385;
	wire n2386;
	wire n2387;
	wire n2388;
	wire n2389;
	wire n2390;
	wire n2391;
	wire n2392;
	wire n2393;
	wire n2394;
	wire n2395;
	wire n2396;
	wire n2397;
	wire n2398;
	wire n2399;
	wire n2400;
	wire n2401;
	wire n2402;
	wire n2403;
	wire n2404;
	wire n2405;
	wire n2406;
	wire n2407;
	wire n2408;
	wire n2409;
	wire n2410;
	wire n2411;
	wire n2412;
	wire n2413;
	wire n2414;
	wire n2415;
	wire n2416;
	wire n2417;
	wire n2418;
	wire n2419;
	wire n2420;
	wire n2421;
	wire n2422;
	wire n2423;
	wire n2424;
	wire n2425;
	wire n2426;
	wire n2427;
	wire n2428;
	wire n2429;
	wire n2430;
	wire n2431;
	wire n2432;
	wire n2433;
	wire n2434;
	wire n2435;
	wire n2436;
	wire n2437;
	wire n2438;
	wire n2439;
	wire n2440;
	wire n2441;
	wire n2442;
	wire n2443;
	wire n2444;
	wire n2445;
	wire n2446;
	wire n2447;
	wire n2448;
	wire n2449;
	wire n2450;
	wire n2451;
	wire n2452;
	wire n2453;
	wire n2454;
	wire n2455;
	wire n2456;
	wire n2457;
	wire n2458;
	wire n2459;
	wire n2460;
	wire n2461;
	wire n2462;
	wire n2463;
	wire n2464;
	wire n2465;
	wire n2466;
	wire n2467;
	wire n2468;
	wire n2469;
	wire n2470;
	wire n2471;
	wire n2472;
	wire n2473;
	wire n2474;
	wire n2475;
	wire n2476;
	wire n2477;
	wire n2478;
	wire n2479;
	wire n2480;
	wire n2481;
	wire n2482;
	wire n2483;
	wire n2484;
	wire n2485;
	wire n2486;
	wire n2487;
	wire n2488;
	wire n2489;
	wire n2490;
	wire n2491;
	wire n2492;
	wire n2493;
	wire n2494;
	wire n2495;
	wire n2496;
	wire n2497;
	wire n2498;
	wire n2499;
	wire n2500;
	wire n2501;
	wire n2502;
	wire n2503;
	wire n2504;
	wire n2505;
	wire n2506;
	wire n2507;
	wire n2508;
	wire n2509;
	wire n2510;
	wire n2511;
	wire n2512;
	wire n2513;
	wire n2514;
	wire n2515;
	wire n2516;
	wire n2517;
	wire n2518;
	wire n2519;
	wire n2520;
	wire n2521;
	wire n2522;
	wire n2523;
	wire n2524;
	wire n2525;
	wire n2526;
	wire n2527;
	wire n2528;
	wire n2529;
	wire n2530;
	wire n2531;
	wire n2532;
	wire n2533;
	wire n2534;
	wire n2535;
	wire n2536;
	wire n2537;
	wire n2538;
	wire n2539;
	wire n2540;
	wire n2541;
	wire n2542;
	wire n2543;
	wire n2544;
	wire n2545;
	wire n2546;
	wire n2547;
	wire n2548;
	wire n2549;
	wire n2550;
	wire n2551;
	wire n2552;
	wire n2553;
	wire n2554;
	wire n2555;
	wire n2556;
	wire n2557;
	wire n2558;
	wire n2559;
	wire n2560;
	wire n2561;
	wire n2563;
	wire n2564;
	wire n2565;
	wire n2566;
	wire n2567;
	wire n2568;
	wire n2569;
	wire n2570;
	wire n2571;
	wire n2572;
	wire n2573;
	wire n2574;
	wire n2575;
	wire n2576;
	wire n2577;
	wire n2578;
	wire n2579;
	wire n2580;
	wire n2581;
	wire n2582;
	wire n2583;
	wire n2584;
	wire n2585;
	wire n2586;
	wire n2587;
	wire n2588;
	wire n2589;
	wire n2590;
	wire n2591;
	wire n2592;
	wire n2593;
	wire n2594;
	wire n2595;
	wire n2596;
	wire n2597;
	wire n2598;
	wire n2599;
	wire n2600;
	wire n2601;
	wire n2602;
	wire n2603;
	wire n2604;
	wire n2605;
	wire n2606;
	wire n2607;
	wire n2608;
	wire n2609;
	wire n2610;
	wire n2611;
	wire n2612;
	wire n2613;
	wire n2614;
	wire n2615;
	wire n2616;
	wire n2617;
	wire n2618;
	wire n2619;
	wire n2620;
	wire n2621;
	wire n2622;
	wire n2623;
	wire n2624;
	wire n2625;
	wire n2626;
	wire n2627;
	wire n2628;
	wire n2629;
	wire n2630;
	wire n2631;
	wire n2632;
	wire n2633;
	wire n2634;
	wire n2635;
	wire n2636;
	wire n2637;
	wire n2638;
	wire n2639;
	wire n2640;
	wire n2641;
	wire n2642;
	wire n2643;
	wire n2644;
	wire n2645;
	wire n2646;
	wire n2647;
	wire n2648;
	wire n2649;
	wire n2650;
	wire n2651;
	wire n2652;
	wire n2653;
	wire n2654;
	wire n2655;
	wire n2656;
	wire n2657;
	wire n2658;
	wire n2659;
	wire n2660;
	wire n2661;
	wire n2662;
	wire n2663;
	wire n2664;
	wire n2665;
	wire n2666;
	wire n2667;
	wire n2668;
	wire n2669;
	wire n2670;
	wire n2671;
	wire n2672;
	wire n2673;
	wire n2674;
	wire n2675;
	wire n2676;
	wire n2677;
	wire n2678;
	wire n2679;
	wire n2680;
	wire n2681;
	wire n2682;
	wire n2683;
	wire n2684;
	wire n2685;
	wire n2686;
	wire n2687;
	wire n2688;
	wire n2689;
	wire n2690;
	wire n2691;
	wire n2692;
	wire n2693;
	wire n2694;
	wire n2695;
	wire n2696;
	wire n2697;
	wire n2698;
	wire n2699;
	wire n2700;
	wire n2701;
	wire n2702;
	wire n2703;
	wire n2704;
	wire n2705;
	wire n2706;
	wire n2707;
	wire n2708;
	wire n2709;
	wire n2710;
	wire n2711;
	wire n2712;
	wire n2713;
	wire n2714;
	wire n2715;
	wire n2716;
	wire n2717;
	wire n2719;
	wire n2720;
	wire n2721;
	wire n2722;
	wire n2723;
	wire n2724;
	wire n2725;
	wire n2726;
	wire n2727;
	wire n2728;
	wire n2729;
	wire n2730;
	wire n2733;
	wire n2734;
	wire n2735;
	wire n2736;
	wire n2737;
	wire n2738;
	wire n2739;
	wire n2740;
	wire n2741;
	wire n2742;
	wire n2743;
	wire n2744;
	wire n2746;
	wire n2747;
	wire n2748;
	wire n2749;
	wire n2750;
	wire n2751;
	wire n2752;
	wire n2753;
	wire n2754;
	wire n2755;
	wire n2756;
	wire n2757;
	wire n2758;
	wire n2759;
	wire n2760;
	wire n2761;
	wire n2762;
	wire n2763;
	wire n2764;
	wire n2765;
	wire n2766;
	wire n2767;
	wire n2768;
	wire n2769;
	wire n2770;
	wire n2771;
	wire n2772;
	wire n2773;
	wire n2774;
	wire n2775;
	wire n2776;
	wire n2777;
	wire n2778;
	wire n2779;
	wire n2780;
	wire n2781;
	wire n2782;
	wire n2783;
	wire n2784;
	wire n2785;
	wire n2786;
	wire n2787;
	wire n2788;
	wire n2789;
	wire n2790;
	wire n2791;
	wire n2792;
	wire n2793;
	wire n2794;
	wire n2795;
	wire n2796;
	wire n2797;
	wire n2798;
	wire n2799;
	wire n2800;
	wire n2801;
	wire n2802;
	wire n2803;
	wire n2804;
	wire n2805;
	wire n2806;
	wire n2807;
	wire n2808;
	wire n2809;
	wire n2810;
	wire n2811;
	wire n2812;
	wire n2813;
	wire n2814;
	wire n2815;
	wire n2816;
	wire n2817;
	wire n2818;
	wire n2819;
	wire n2820;
	wire n2821;
	wire n2822;
	wire n2823;
	wire n2824;
	wire n2825;
	wire n2826;
	wire n2827;
	wire n2828;
	wire n2829;
	wire n2830;
	wire n2831;
	wire n2833;
	wire n2834;
	wire n2835;
	wire n2836;
	wire n2837;
	wire n2838;
	wire n2839;
	wire n2840;
	wire n2841;
	wire n2842;
	wire n2843;
	wire n2844;
	wire n2845;
	wire n2846;
	wire n2847;
	wire n2848;
	wire n2849;
	wire n2850;
	wire n2851;
	wire n2852;
	wire n2853;
	wire n2854;
	wire n2855;
	wire n2856;
	wire n2857;
	wire n2858;
	wire n2859;
	wire n2860;
	wire n2861;
	wire n2862;
	wire n2863;
	wire n2864;
	wire n2865;
	wire n2866;
	wire n2867;
	wire n2868;
	wire n2869;
	wire n2870;
	wire n2871;
	wire n2872;
	wire n2873;
	wire n2874;
	wire n2875;
	wire n2876;
	wire n2877;
	wire n2878;
	wire n2879;
	wire n2880;
	wire n2881;
	wire n2882;
	wire n2883;
	wire n2884;
	wire n2885;
	wire n2886;
	wire n2887;
	wire n2888;
	wire n2889;
	wire n2890;
	wire n2891;
	wire n2892;
	wire n2893;
	wire n2894;
	wire n2895;
	wire n2896;
	wire n2897;
	wire n2898;
	wire n2899;
	wire n2900;
	wire n2901;
	wire n2902;
	wire n2903;
	wire n2904;
	wire n2905;
	wire n2906;
	wire n2907;
	wire n2908;
	wire n2909;
	wire n2910;
	wire n2911;
	wire n2912;
	wire n2913;
	wire n2914;
	wire n2915;
	wire n2916;
	wire n2917;
	wire n2918;
	wire n2919;
	wire n2920;
	wire n2921;
	wire n2922;
	wire n2923;
	wire n2924;
	wire n2925;
	wire n2926;
	wire n2927;
	wire n2928;
	wire n2929;
	wire n2930;
	wire n2931;
	wire n2932;
	wire n2933;
	wire n2934;
	wire n2935;
	wire n2936;
	wire n2937;
	wire n2938;
	wire n2939;
	wire n2940;
	wire n2941;
	wire n2942;
	wire n2943;
	wire n2944;
	wire n2945;
	wire n2946;
	wire n2947;
	wire n2948;
	wire n2949;
	wire n2950;
	wire n2951;
	wire n2952;
	wire n2953;
	wire n2954;
	wire n2955;
	wire n2956;
	wire n2957;
	wire n2958;
	wire n2959;
	wire n2960;
	wire n2961;
	wire n2962;
	wire n2963;
	wire n2964;
	wire n2965;
	wire n2966;
	wire n2967;
	wire n2968;
	wire n2969;
	wire n2970;
	wire n2971;
	wire n2972;
	wire n2973;
	wire n2974;
	wire n2975;
	wire n2976;
	wire n2977;
	wire n2978;
	wire n2979;
	wire n2980;
	wire n2981;
	wire n2982;
	wire n2983;
	wire n2984;
	wire n2985;
	wire n2986;
	wire n2987;
	wire n2988;
	wire n2989;
	wire n2990;
	wire n2991;
	wire n2992;
	wire n2993;
	wire n2994;
	wire n2995;
	wire n2996;
	wire n2997;
	wire n2998;
	wire n2999;
	wire n3000;
	wire n3001;
	wire n3002;
	wire n3003;
	wire n3004;
	wire n3005;
	wire n3006;
	wire n3007;
	wire n3008;
	wire n3009;
	wire n3010;
	wire n3011;
	wire n3012;
	wire n3013;
	wire n3014;
	wire n3015;
	wire n3016;
	wire n3017;
	wire n3018;
	wire n3019;
	wire n3020;
	wire n3021;
	wire n3022;
	wire n3023;
	wire n3024;
	wire n3025;
	wire n3026;
	wire n3027;
	wire n3028;
	wire n3029;
	wire n3030;
	wire n3031;
	wire n3032;
	wire n3033;
	wire n3034;
	wire n3035;
	wire n3036;
	wire n3037;
	wire n3038;
	wire n3039;
	wire n3040;
	wire n3041;
	wire n3042;
	wire n3043;
	wire n3044;
	wire n3045;
	wire n3046;
	wire n3047;
	wire n3048;
	wire n3049;
	wire n3050;
	wire n3051;
	wire n3052;
	wire n3053;
	wire n3054;
	wire n3055;
	wire n3056;
	wire n3057;
	wire n3058;
	wire n3059;
	wire n3060;
	wire n3061;
	wire n3062;
	wire n3063;
	wire n3064;
	wire n3065;
	wire n3066;
	wire n3067;
	wire n3068;
	wire n3069;
	wire n3070;
	wire n3071;
	wire n3072;
	wire n3073;
	wire n3075;
	wire n3076;
	wire n3077;
	wire n3078;
	wire n3079;
	wire n3080;
	wire n3081;
	wire n3082;
	wire n3083;
	wire n3084;
	wire n3085;
	wire n3086;
	wire n3087;
	wire n3088;
	wire n3089;
	wire n3090;
	wire n3091;
	wire n3092;
	wire n3093;
	wire n3094;
	wire n3095;
	wire n3096;
	wire n3097;
	wire n3098;
	wire n3099;
	wire n3100;
	wire n3101;
	wire n3102;
	wire n3103;
	wire n3104;
	wire n3105;
	wire n3106;
	wire n3107;
	wire n3108;
	wire n3109;
	wire n3110;
	wire n3111;
	wire n3112;
	wire n3113;
	wire n3114;
	wire n3115;
	wire n3116;
	wire n3117;
	wire n3118;
	wire n3119;
	wire n3120;
	wire n3121;
	wire n3122;
	wire n3123;
	wire n3124;
	wire n3125;
	wire n3126;
	wire n3127;
	wire n3128;
	wire n3129;
	wire n3130;
	wire n3131;
	wire n3132;
	wire n3133;
	wire n3134;
	wire n3135;
	wire n3136;
	wire n3137;
	wire n3138;
	wire n3139;
	wire n3140;
	wire n3141;
	wire n3142;
	wire n3143;
	wire n3144;
	wire n3145;
	wire n3146;
	wire n3147;
	wire n3148;
	wire n3149;
	wire n3150;
	wire n3151;
	wire n3152;
	wire n3153;
	wire n3154;
	wire n3155;
	wire n3156;
	wire n3157;
	wire n3158;
	wire n3159;
	wire n3160;
	wire n3161;
	wire n3162;
	wire n3163;
	wire n3164;
	wire n3165;
	wire n3166;
	wire n3167;
	wire n3168;
	wire n3169;
	wire n3170;
	wire n3171;
	wire n3172;
	wire n3173;
	wire n3174;
	wire n3175;
	wire n3176;
	wire n3177;
	wire n3178;
	wire n3179;
	wire n3180;
	wire n3181;
	wire n3182;
	wire n3183;
	wire n3184;
	wire n3185;
	wire n3186;
	wire n3187;
	wire n3188;
	wire n3189;
	wire n3190;
	wire n3191;
	wire n3192;
	wire n3193;
	wire n3194;
	wire n3195;
	wire n3196;
	wire n3197;
	wire n3198;
	wire n3199;
	wire n3200;
	wire n3201;
	wire n3202;
	wire n3203;
	wire n3204;
	wire n3205;
	wire n3206;
	wire n3207;
	wire n3208;
	wire n3209;
	wire n3210;
	wire n3211;
	wire n3212;
	wire n3213;
	wire n3214;
	wire n3215;
	wire n3216;
	wire n3217;
	wire n3218;
	wire n3219;
	wire n3220;
	wire n3221;
	wire n3222;
	wire n3223;
	wire n3224;
	wire n3225;
	wire n3226;
	wire n3227;
	wire n3228;
	wire n3229;
	wire n3230;
	wire n3231;
	wire n3232;
	wire n3233;
	wire n3234;
	wire n3235;
	wire n3236;
	wire n3237;
	wire n3238;
	wire n3239;
	wire n3240;
	wire n3241;
	wire n3242;
	wire n3243;
	wire n3244;
	wire n3245;
	wire n3246;
	wire n3247;
	wire n3248;
	wire n3249;
	wire n3250;
	wire n3251;
	wire n3252;
	wire n3253;
	wire n3254;
	wire n3255;
	wire n3257;
	wire n3258;
	wire n3259;
	wire n3260;
	wire n3261;
	wire n3262;
	wire n3263;
	wire n3264;
	wire n3265;
	wire n3266;
	wire n3267;
	wire n3268;
	wire n3269;
	wire n3270;
	wire n3271;
	wire n3272;
	wire n3273;
	wire n3274;
	wire n3275;
	wire n3276;
	wire n3277;
	wire n3278;
	wire n3279;
	wire n3280;
	wire n3281;
	wire n3282;
	wire n3283;
	wire n3284;
	wire n3285;
	wire n3286;
	wire n3287;
	wire n3288;
	wire n3289;
	wire n3290;
	wire n3291;
	wire n3292;
	wire n3293;
	wire n3294;
	wire n3295;
	wire n3296;
	wire n3297;
	wire n3298;
	wire n3299;
	wire n3300;
	wire n3301;
	wire n3302;
	wire n3303;
	wire n3304;
	wire n3305;
	wire n3306;
	wire n3307;
	wire n3308;
	wire n3309;
	wire n3310;
	wire n3311;
	wire n3312;
	wire n3313;
	wire n3314;
	wire n3315;
	wire n3316;
	wire n3317;
	wire n3318;
	wire n3319;
	wire n3320;
	wire n3321;
	wire n3322;
	wire n3323;
	wire n3324;
	wire n3325;
	wire n3326;
	wire n3327;
	wire n3328;
	wire n3329;
	wire n3330;
	wire n3331;
	wire n3332;
	wire n3333;
	wire n3334;
	wire n3335;
	wire n3336;
	wire n3337;
	wire n3338;
	wire n3339;
	wire n3340;
	wire n3341;
	wire n3342;
	wire n3343;
	wire n3344;
	wire n3345;
	wire n3346;
	wire n3347;
	wire n3348;
	wire n3349;
	wire n3350;
	wire n3351;
	wire n3352;
	wire n3353;
	wire n3354;
	wire n3355;
	wire n3356;
	wire n3357;
	wire n3358;
	wire n3359;
	wire n3360;
	wire n3361;
	wire n3362;
	wire n3363;
	wire n3364;
	wire n3365;
	wire n3366;
	wire n3367;
	wire n3368;
	wire n3369;
	wire n3370;
	wire n3371;
	wire n3372;
	wire n3373;
	wire n3374;
	wire n3375;
	wire n3376;
	wire n3377;
	wire n3378;
	wire n3379;
	wire n3380;
	wire n3381;
	wire n3382;
	wire n3383;
	wire n3384;
	wire n3385;
	wire n3386;
	wire n3387;
	wire n3388;
	wire n3389;
	wire n3390;
	wire n3391;
	wire n3392;
	wire n3393;
	wire n3394;
	wire n3395;
	wire n3396;
	wire n3397;
	wire n3398;
	wire n3399;
	wire n3400;
	wire n3401;
	wire n3402;
	wire n3403;
	wire n3404;
	wire n3405;
	wire n3406;
	wire n3407;
	wire n3408;
	wire n3409;
	wire n3410;
	wire n3411;
	wire n3412;
	wire n3413;
	wire n3414;
	wire n3415;
	wire n3416;
	wire n3417;
	wire n3418;
	wire n3419;
	wire n3420;
	wire n3421;
	wire n3422;
	wire n3423;
	wire n3424;
	wire n3425;
	wire n3426;
	wire n3427;
	wire n3428;
	wire n3429;
	wire n3430;
	wire n3431;
	wire n3432;
	wire n3433;
	wire n3434;
	wire n3435;
	wire n3436;
	wire n3437;
	wire n3438;
	wire n3439;
	wire n3440;
	wire n3441;
	wire n3442;
	wire n3443;
	wire n3444;
	wire n3445;
	wire n3446;
	wire n3447;
	wire n3448;
	wire n3449;
	wire n3450;
	wire n3451;
	wire n3452;
	wire n3453;
	wire n3454;
	wire n3455;
	wire n3456;
	wire n3457;
	wire n3458;
	wire n3459;
	wire n3460;
	wire n3461;
	wire n3462;
	wire n3463;
	wire n3464;
	wire n3465;
	wire n3466;
	wire n3467;
	wire n3468;
	wire n3469;
	wire n3470;
	wire n3471;
	wire n3472;
	wire n3473;
	wire n3474;
	wire n3475;
	wire n3476;
	wire n3477;
	wire n3478;
	wire n3479;
	wire n3480;
	wire n3481;
	wire n3482;
	wire n3483;
	wire n3484;
	wire n3485;
	wire n3486;
	wire n3487;
	wire n3488;
	wire n3489;
	wire n3490;
	wire n3491;
	wire n3492;
	wire n3493;
	wire n3494;
	wire n3495;
	wire n3496;
	wire n3497;
	wire n3498;
	wire n3499;
	wire n3500;
	wire n3501;
	wire n3502;
	wire n3503;
	wire n3504;
	wire n3505;
	wire n3506;
	wire n3507;
	wire n3508;
	wire n3509;
	wire n3510;
	wire n3511;
	wire n3512;
	wire n3513;
	wire n3514;
	wire n3515;
	wire n3516;
	wire n3517;
	wire n3518;
	wire n3519;
	wire n3520;
	wire n3521;
	wire n3522;
	wire n3523;
	wire n3524;
	wire n3526;
	wire n3527;
	wire n3528;
	wire n3529;
	wire n3530;
	wire n3531;
	wire n3532;
	wire n3533;
	wire n3534;
	wire n3535;
	wire n3536;
	wire n3537;
	wire n3538;
	wire n3539;
	wire n3540;
	wire n3541;
	wire n3542;
	wire n3543;
	wire n3544;
	wire n3545;
	wire n3546;
	wire n3547;
	wire n3548;
	wire n3549;
	wire n3550;
	wire n3551;
	wire n3552;
	wire n3553;
	wire n3554;
	wire n3555;
	wire n3556;
	wire n3557;
	wire n3558;
	wire n3559;
	wire n3560;
	wire n3561;
	wire n3562;
	wire n3563;
	wire n3564;
	wire n3565;
	wire n3566;
	wire n3567;
	wire n3568;
	wire n3569;
	wire n3570;
	wire n3571;
	wire n3572;
	wire n3573;
	wire n3574;
	wire n3575;
	wire n3576;
	wire n3577;
	wire n3578;
	wire n3579;
	wire n3580;
	wire n3581;
	wire n3582;
	wire n3583;
	wire n3584;
	wire n3585;
	wire n3586;
	wire n3587;
	wire n3588;
	wire n3589;
	wire n3590;
	wire n3591;
	wire n3592;
	wire n3593;
	wire n3594;
	wire n3595;
	wire n3596;
	wire n3597;
	wire n3598;
	wire n3599;
	wire n3600;
	wire n3601;
	wire n3602;
	wire n3603;
	wire n3604;
	wire n3605;
	wire n3606;
	wire n3607;
	wire n3608;
	wire n3609;
	wire n3610;
	wire n3611;
	wire n3612;
	wire n3613;
	wire n3614;
	wire n3615;
	wire n3616;
	wire n3617;
	wire n3618;
	wire n3619;
	wire n3620;
	wire n3621;
	wire n3622;
	wire n3623;
	wire n3624;
	wire n3625;
	wire n3626;
	wire n3627;
	wire n3628;
	wire n3629;
	wire n3630;
	wire n3631;
	wire n3635;
	wire n3636;
	wire n3637;
	wire n3638;
	wire n3639;
	wire n3640;
	wire n3642;
	wire n3643;
	wire n3644;
	wire n3645;
	wire n3646;
	wire n3647;
	wire n3648;
	wire n3649;
	wire n3650;
	wire n3651;
	wire n3652;
	wire n3653;
	wire n3654;
	wire n3655;
	wire n3656;
	wire n3657;
	wire n3658;
	wire n3659;
	wire n3660;
	wire n3661;
	wire n3662;
	wire n3663;
	wire n3664;
	wire n3665;
	wire n3666;
	wire n3667;
	wire n3668;
	wire n3669;
	wire n3670;
	wire n3671;
	wire n3672;
	wire n3673;
	wire n3674;
	wire n3675;
	wire n3676;
	wire n3677;
	wire n3678;
	wire n3679;
	wire n3680;
	wire n3681;
	wire n3682;
	wire n3683;
	wire n3684;
	wire n3685;
	wire n3686;
	wire n3687;
	wire n3688;
	wire n3689;
	wire n3690;
	wire n3691;
	wire n3692;
	wire n3693;
	wire n3694;
	wire n3695;
	wire n3696;
	wire n3697;
	wire n3698;
	wire n3699;
	wire n3700;
	wire n3701;
	wire n3702;
	wire n3703;
	wire n3704;
	wire n3705;
	wire n3706;
	wire n3707;
	wire n3708;
	wire n3709;
	wire n3710;
	wire n3711;
	wire n3712;
	wire n3713;
	wire n3714;
	wire n3715;
	wire n3716;
	wire n3717;
	wire n3718;
	wire n3719;
	wire n3720;
	wire n3721;
	wire n3722;
	wire n3723;
	wire n3724;
	wire n3725;
	wire n3726;
	wire n3727;
	wire n3728;
	wire n3729;
	wire n3730;
	wire n3731;
	wire n3732;
	wire n3733;
	wire n3734;
	wire n3735;
	wire n3736;
	wire n3737;
	wire n3738;
	wire n3739;
	wire n3740;
	wire n3741;
	wire n3742;
	wire n3743;
	wire n3744;
	wire n3745;
	wire n3746;
	wire n3747;
	wire n3748;
	wire n3749;
	wire n3750;
	wire n3751;
	wire n3752;
	wire n3753;
	wire n3754;
	wire n3755;
	wire n3756;
	wire n3757;
	wire n3758;
	wire n3759;
	wire n3760;
	wire n3761;
	wire n3762;
	wire n3763;
	wire n3764;
	wire n3765;
	wire n3766;
	wire n3767;
	wire n3768;
	wire n3769;
	wire n3770;
	wire n3771;
	wire n3772;
	wire n3773;
	wire n3774;
	wire n3775;
	wire n3776;
	wire n3777;
	wire n3778;
	wire n3779;
	wire n3780;
	wire n3781;
	wire n3782;
	wire n3783;
	wire n3784;
	wire n3785;
	wire n3786;
	wire n3787;
	wire n3788;
	wire n3789;
	wire n3790;
	wire n3791;
	wire n3792;
	wire n3793;
	wire n3794;
	wire n3795;
	wire n3796;
	wire n3797;
	wire n3798;
	wire n3799;
	wire n3800;
	wire n3801;
	wire n3802;
	wire n3803;
	wire n3804;
	wire n3805;
	wire n3806;
	wire n3807;
	wire n3808;
	wire n3809;
	wire n3810;
	wire n3811;
	wire n3812;
	wire n3813;
	wire n3814;
	wire n3815;
	wire n3816;
	wire n3817;
	wire n3818;
	wire n3819;
	wire n3820;
	wire n3821;
	wire n3822;
	wire n3823;
	wire n3824;
	wire n3825;
	wire n3826;
	wire n3827;
	wire n3828;
	wire n3829;
	wire n3830;
	wire n3832;
	wire n3833;
	wire n3834;
	wire n3835;
	wire n3836;
	wire n3837;
	wire n3838;
	wire n3839;
	wire n3840;
	wire n3841;
	wire n3842;
	wire n3843;
	wire n3844;
	wire n3845;
	wire n3846;
	wire n3847;
	wire n3848;
	wire n3849;
	wire n3850;
	wire n3851;
	wire n3852;
	wire n3853;
	wire n3854;
	wire n3855;
	wire n3856;
	wire n3857;
	wire n3858;
	wire n3859;
	wire n3860;
	wire n3861;
	wire n3862;
	wire n3863;
	wire n3864;
	wire n3865;
	wire n3866;
	wire n3867;
	wire n3868;
	wire n3869;
	wire n3870;
	wire n3871;
	wire n3872;
	wire n3873;
	wire n3874;
	wire n3875;
	wire n3876;
	wire n3877;
	wire n3878;
	wire n3879;
	wire n3880;
	wire n3881;
	wire n3882;
	wire n3883;
	wire n3884;
	wire n3885;
	wire n3886;
	wire n3887;
	wire n3888;
	wire n3889;
	wire n3890;
	wire n3891;
	wire n3892;
	wire n3893;
	wire n3894;
	wire n3895;
	wire n3896;
	wire n3897;
	wire n3898;
	wire n3899;
	wire n3900;
	wire n3901;
	wire n3902;
	wire n3903;
	wire n3904;
	wire n3905;
	wire n3906;
	wire n3907;
	wire n3908;
	wire n3909;
	wire n3910;
	wire n3911;
	wire n3912;
	wire n3913;
	wire n3914;
	wire n3915;
	wire n3916;
	wire n3917;
	wire n3918;
	wire n3919;
	wire n3920;
	wire n3921;
	wire n3922;
	wire n3923;
	wire n3924;
	wire n3925;
	wire n3926;
	wire n3927;
	wire n3928;
	wire n3929;
	wire n3930;
	wire n3931;
	wire n3932;
	wire n3933;
	wire n3934;
	wire n3935;
	wire n3936;
	wire n3937;
	wire n3938;
	wire n3939;
	wire n3940;
	wire n3941;
	wire n3942;
	wire n3943;
	wire n3944;
	wire n3945;
	wire n3946;
	wire n3947;
	wire n3948;
	wire n3949;
	wire n3950;
	wire n3951;
	wire n3952;
	wire n3953;
	wire n3954;
	wire n3955;
	wire n3956;
	wire n3957;
	wire n3958;
	wire n3959;
	wire n3960;
	wire n3961;
	wire n3962;
	wire n3963;
	wire n3964;
	wire n3965;
	wire n3966;
	wire n3967;
	wire n3968;
	wire n3969;
	wire n3970;
	wire n3971;
	wire n3972;
	wire n3973;
	wire n3974;
	wire n3975;
	wire n3976;
	wire n3977;
	wire n3978;
	wire n3979;
	wire n3980;
	wire n3981;
	wire n3982;
	wire n3983;
	wire n3984;
	wire n3985;
	wire n3986;
	wire n3987;
	wire n3988;
	wire n3989;
	wire n3990;
	wire n3991;
	wire n3992;
	wire n3993;
	wire n3994;
	wire n3995;
	wire n3996;
	wire n3997;
	wire n3998;
	wire n3999;
	wire n4000;
	wire n4001;
	wire n4002;
	wire n4003;
	wire n4004;
	wire n4005;
	wire n4006;
	wire n4007;
	wire n4008;
	wire n4009;
	wire n4010;
	wire n4011;
	wire n4012;
	wire n4013;
	wire n4014;
	wire n4015;
	wire n4016;
	wire n4017;
	wire n4018;
	wire n4019;
	wire n4020;
	wire n4021;
	wire n4022;
	wire n4023;
	wire n4024;
	wire n4025;
	wire n4026;
	wire n4027;
	wire n4028;
	wire n4029;
	wire n4030;
	wire n4031;
	wire n4032;
	wire n4033;
	wire n4034;
	wire n4035;
	wire n4036;
	wire n4037;
	wire n4038;
	wire n4039;
	wire n4040;
	wire n4041;
	wire n4042;
	wire n4043;
	wire n4044;
	wire n4045;
	wire n4046;
	wire n4047;
	wire n4048;
	wire n4049;
	wire n4050;
	wire n4051;
	wire n4052;
	wire n4053;
	wire n4054;
	wire n4055;
	wire n4056;
	wire n4057;
	wire n4058;
	wire n4059;
	wire n4060;
	wire n4061;
	wire n4062;
	wire n4063;
	wire n4064;
	wire n4065;
	wire n4066;
	wire n4067;
	wire n4068;
	wire n4069;
	wire n4070;
	wire n4071;
	wire n4072;
	wire n4073;
	wire n4074;
	wire n4075;
	wire n4076;
	wire n4077;
	wire n4078;
	wire n4079;
	wire n4080;
	wire n4081;
	wire n4082;
	wire n4083;
	wire n4084;
	wire n4085;
	wire n4086;
	wire n4087;
	wire n4088;
	wire n4089;
	wire n4090;
	wire n4091;
	wire n4092;
	wire n4093;
	wire n4094;
	wire n4095;
	wire n4096;
	wire n4097;
	wire n4098;
	wire n4099;
	wire n4100;
	wire n4101;
	wire n4102;
	wire n4103;
	wire n4104;
	wire n4105;
	wire n4106;
	wire n4107;
	wire n4108;
	wire n4109;
	wire n4110;
	wire n4111;
	wire n4112;
	wire n4113;
	wire n4114;
	wire n4115;
	wire n4116;
	wire n4117;
	wire n4118;
	wire n4119;
	wire n4120;
	wire n4121;
	wire n4122;
	wire n4123;
	wire n4124;
	wire n4125;
	wire n4126;
	wire n4127;
	wire n4128;
	wire n4129;
	wire n4130;
	wire n4131;
	wire n4132;
	wire n4133;
	wire n4134;
	wire n4135;
	wire n4136;
	wire n4137;
	wire n4138;
	wire n4139;
	wire n4140;
	wire n4141;
	wire n4142;
	wire n4143;
	wire n4144;
	wire n4145;
	wire n4146;
	wire n4147;
	wire n4148;
	wire n4149;
	wire n4150;
	wire n4151;
	wire n4152;
	wire n4153;
	wire n4154;
	wire n4155;
	wire n4156;
	wire n4157;
	wire n4158;
	wire n4159;
	wire n4160;
	wire n4161;
	wire n4162;
	wire n4163;
	wire n4164;
	wire n4165;
	wire n4166;
	wire n4167;
	wire n4168;
	wire n4169;
	wire n4170;
	wire n4171;
	wire n4172;
	wire n4173;
	wire n4174;
	wire n4175;
	wire n4176;
	wire n4177;
	wire n4178;
	wire n4179;
	wire n4180;
	wire n4181;
	wire n4182;
	wire n4183;
	wire n4184;
	wire n4185;
	wire n4186;
	wire n4187;
	wire n4188;
	wire n4189;
	wire n4190;
	wire n4191;
	wire n4192;
	wire n4193;
	wire n4194;
	wire n4195;
	wire n4196;
	wire n4197;
	wire n4198;
	wire n4199;
	wire n4200;
	wire n4201;
	wire n4202;
	wire n4203;
	wire n4204;
	wire n4205;
	wire n4206;
	wire n4207;
	wire n4208;
	wire n4209;
	wire n4210;
	wire n4211;
	wire n4212;
	wire n4213;
	wire n4214;
	wire n4215;
	wire n4216;
	wire n4217;
	wire n4218;
	wire n4219;
	wire n4220;
	wire n4221;
	wire n4222;
	wire n4223;
	wire n4224;
	wire n4225;
	wire n4226;
	wire n4227;
	wire n4228;
	wire n4229;
	wire n4230;
	wire n4231;
	wire n4232;
	wire n4233;
	wire n4234;
	wire n4235;
	wire n4237;
	wire n4238;
	wire n4239;
	wire n4240;
	wire n4241;
	wire n4242;
	wire n4243;
	wire n4244;
	wire n4245;
	wire n4246;
	wire n4247;
	wire n4248;
	wire n4249;
	wire n4250;
	wire n4251;
	wire n4252;
	wire n4253;
	wire n4254;
	wire n4255;
	wire n4256;
	wire n4257;
	wire n4258;
	wire n4259;
	wire n4260;
	wire n4261;
	wire n4262;
	wire n4263;
	wire n4264;
	wire n4265;
	wire n4266;
	wire n4267;
	wire n4268;
	wire n4269;
	wire n4270;
	wire n4271;
	wire n4272;
	wire n4273;
	wire n4274;
	wire n4275;
	wire n4276;
	wire n4277;
	wire n4278;
	wire n4279;
	wire n4280;
	wire n4281;
	wire n4282;
	wire n4283;
	wire n4284;
	wire n4285;
	wire n4286;
	wire n4287;
	wire n4288;
	wire n4289;
	wire n4290;
	wire n4291;
	wire n4292;
	wire n4293;
	wire n4294;
	wire n4295;
	wire n4296;
	wire n4297;
	wire n4298;
	wire n4299;
	wire n4300;
	wire n4301;
	wire n4302;
	wire n4303;
	wire n4304;
	wire n4305;
	wire n4306;
	wire n4307;
	wire n4308;
	wire n4309;
	wire n4310;
	wire n4311;
	wire n4312;
	wire n4313;
	wire n4314;
	wire n4315;
	wire n4316;
	wire n4317;
	wire n4318;
	wire n4319;
	wire n4320;
	wire n4321;
	wire n4322;
	wire n4323;
	wire n4324;
	wire n4325;
	wire n4326;
	wire n4327;
	wire n4328;
	wire n4329;
	wire n4330;
	wire n4331;
	wire n4332;
	wire n4333;
	wire n4334;
	wire n4335;
	wire n4336;
	wire n4337;
	wire n4338;
	wire n4339;
	wire n4340;
	wire n4341;
	wire n4342;
	wire n4343;
	wire n4344;
	wire n4345;
	wire n4346;
	wire n4347;
	wire n4348;
	wire n4349;
	wire n4350;
	wire n4351;
	wire n4352;
	wire n4353;
	wire n4354;
	wire n4355;
	wire n4356;
	wire n4357;
	wire n4358;
	wire n4359;
	wire n4360;
	wire n4361;
	wire n4362;
	wire n4363;
	wire n4364;
	wire n4365;
	wire n4366;
	wire n4367;
	wire n4368;
	wire n4369;
	wire n4370;
	wire n4371;
	wire n4372;
	wire n4373;
	wire n4374;
	wire n4375;
	wire n4376;
	wire n4377;
	wire n4378;
	wire n4379;
	wire n4380;
	wire n4381;
	wire n4382;
	wire n4383;
	wire n4384;
	wire n4385;
	wire n4386;
	wire n4387;
	wire n4388;
	wire n4389;
	wire n4390;
	wire n4391;
	wire n4392;
	wire n4393;
	wire n4394;
	wire n4395;
	wire n4396;
	wire n4397;
	wire n4398;
	wire n4399;
	wire n4400;
	wire n4401;
	wire n4402;
	wire n4403;
	wire n4404;
	wire n4405;
	wire n4406;
	wire n4407;
	wire n4408;
	wire n4409;
	wire n4410;
	wire n4411;
	wire n4412;
	wire n4413;
	wire n4414;
	wire n4415;
	wire n4416;
	wire n4417;
	wire n4418;
	wire n4419;
	wire n4420;
	wire n4421;
	wire n4422;
	wire n4423;
	wire n4424;
	wire n4425;
	wire n4426;
	wire n4427;
	wire n4428;
	wire n4429;
	wire n4430;
	wire n4431;
	wire n4432;
	wire n4433;
	wire n4434;
	wire n4435;
	wire n4436;
	wire n4437;
	wire n4438;
	wire n4439;
	wire n4440;
	wire n4441;
	wire n4442;
	wire n4443;
	wire n4444;
	wire n4445;
	wire n4446;
	wire n4447;
	wire n4448;
	wire n4449;
	wire n4450;
	wire n4452;
	wire n4453;
	wire n4454;
	wire n4455;
	wire n4456;
	wire n4457;
	wire n4458;
	wire n4459;
	wire n4460;
	wire n4461;
	wire n4462;
	wire n4463;
	wire n4464;
	wire n4465;
	wire n4466;
	wire n4467;
	wire n4468;
	wire n4469;
	wire n4470;
	wire n4471;
	wire n4472;
	wire n4473;
	wire n4474;
	wire n4475;
	wire n4476;
	wire n4477;
	wire n4478;
	wire n4479;
	wire n4480;
	wire n4481;
	wire n4482;
	wire n4483;
	wire n4484;
	wire n4485;
	wire n4486;
	wire n4487;
	wire n4488;
	wire n4489;
	wire n4490;
	wire n4491;
	wire n4492;
	wire n4493;
	wire n4494;
	wire n4495;
	wire n4496;
	wire n4497;
	wire n4498;
	wire n4499;
	wire n4500;
	wire n4501;
	wire n4502;
	wire n4503;
	wire n4504;
	wire n4505;
	wire n4506;
	wire n4507;
	wire n4508;
	wire n4509;
	wire n4510;
	wire n4511;
	wire n4512;
	wire n4513;
	wire n4514;
	wire n4515;
	wire n4516;
	wire n4517;
	wire n4518;
	wire n4519;
	wire n4520;
	wire n4521;
	wire n4522;
	wire n4523;
	wire n4524;
	wire n4525;
	wire n4526;
	wire n4527;
	wire n4528;
	wire n4529;
	wire n4530;
	wire n4531;
	wire n4532;
	wire n4533;
	wire n4534;
	wire n4535;
	wire n4536;
	wire n4537;
	wire n4538;
	wire n4539;
	wire n4540;
	wire n4541;
	wire n4542;
	wire n4543;
	wire n4544;
	wire n4545;
	wire n4546;
	wire n4547;
	wire n4548;
	wire n4549;
	wire n4550;
	wire n4551;
	wire n4552;
	wire n4553;
	wire n4554;
	wire n4555;
	wire n4556;
	wire n4557;
	wire n4558;
	wire n4559;
	wire n4560;
	wire n4561;
	wire n4562;
	wire n4563;
	wire n4564;
	wire n4565;
	wire n4566;
	wire n4567;
	wire n4568;
	wire n4569;
	wire n4570;
	wire n4571;
	wire n4572;
	wire n4573;
	wire n4574;
	wire n4575;
	wire n4576;
	wire n4577;
	wire n4578;
	wire n4579;
	wire n4580;
	wire n4581;
	wire n4582;
	wire n4583;
	wire n4584;
	wire n4585;
	wire n4586;
	wire n4587;
	wire n4588;
	wire n4589;
	wire n4590;
	wire n4591;
	wire n4592;
	wire n4593;
	wire n4594;
	wire n4595;
	wire n4596;
	wire n4597;
	wire n4598;
	wire n4599;
	wire n4600;
	wire n4601;
	wire n4602;
	wire n4603;
	wire n4604;
	wire n4605;
	wire n4606;
	wire n4607;
	wire n4608;
	wire n4609;
	wire n4610;
	wire n4611;
	wire n4612;
	wire n4613;
	wire n4614;
	wire n4615;
	wire n4616;
	wire n4617;
	wire n4618;
	wire n4619;
	wire n4620;
	wire n4621;
	wire n4622;
	wire n4623;
	wire n4624;
	wire n4625;
	wire n4626;
	wire n4627;
	wire n4628;
	wire n4629;
	wire n4630;
	wire n4631;
	wire n4632;
	wire n4633;
	wire n4634;
	wire n4635;
	wire n4636;
	wire n4637;
	wire n4638;
	wire n4639;
	wire n4640;
	wire n4641;
	wire n4642;
	wire n4643;
	wire n4644;
	wire n4645;
	wire n4646;
	wire n4647;
	wire n4648;
	wire n4649;
	wire n4650;
	wire n4651;
	wire n4652;
	wire n4653;
	wire n4654;
	wire n4655;
	wire n4656;
	wire n4657;
	wire n4658;
	wire n4659;
	wire n4660;
	wire n4661;
	wire n4662;
	wire n4663;
	wire n4664;
	wire n4665;
	wire n4666;
	wire n4667;
	wire n4668;
	wire n4669;
	wire n4670;
	wire n4671;
	wire n4672;
	wire n4673;
	wire n4674;
	wire n4675;
	wire n4676;
	wire n4677;
	wire n4678;
	wire n4679;
	wire n4680;
	wire n4681;
	wire n4682;
	wire n4683;
	wire n4684;
	wire n4685;
	wire n4686;
	wire n4687;
	wire n4688;
	wire n4689;
	wire n4690;
	wire n4691;
	wire n4692;
	wire n4693;
	wire n4694;
	wire n4695;
	wire n4696;
	wire n4697;
	wire n4698;
	wire n4699;
	wire n4700;
	wire n4701;
	wire n4702;
	wire n4703;
	wire n4704;
	wire n4705;
	wire n4706;
	wire n4707;
	wire n4708;
	wire n4709;
	wire n4710;
	wire n4711;
	wire n4712;
	wire n4713;
	wire n4714;
	wire n4715;
	wire n4716;
	wire n4717;
	wire n4718;
	wire n4719;
	wire n4720;
	wire n4721;
	wire n4722;
	wire n4723;
	wire n4724;
	wire n4725;
	wire n4726;
	wire n4727;
	wire n4728;
	wire n4729;
	wire n4730;
	wire n4731;
	wire n4732;
	wire n4733;
	wire n4734;
	wire n4735;
	wire n4736;
	wire n4737;
	wire n4738;
	wire n4739;
	wire n4740;
	wire n4741;
	wire n4742;
	wire n4743;
	wire n4744;
	wire n4745;
	wire n4746;
	wire n4747;
	wire n4748;
	wire n4749;
	wire n4750;
	wire n4751;
	wire n4752;
	wire n4753;
	wire n4754;
	wire n4755;
	wire n4756;
	wire n4757;
	wire n4758;
	wire n4759;
	wire n4760;
	wire n4761;
	wire n4762;
	wire n4763;
	wire n4764;
	wire n4765;
	wire n4766;
	wire n4767;
	wire n4768;
	wire n4769;
	wire n4770;
	wire n4771;
	wire n4772;
	wire n4773;
	wire n4774;
	wire n4775;
	wire n4776;
	wire n4777;
	wire n4778;
	wire n4779;
	wire n4780;
	wire n4781;
	wire n4782;
	wire n4783;
	wire n4784;
	wire n4785;
	wire n4786;
	wire n4787;
	wire n4788;
	wire n4789;
	wire n4790;
	wire n4791;
	wire n4792;
	wire n4793;
	wire n4794;
	wire n4795;
	wire n4796;
	wire n4797;
	wire n4798;
	wire n4799;
	wire n4800;
	wire n4801;
	wire n4802;
	wire n4803;
	wire n4804;
	wire n4805;
	wire n4806;
	wire n4807;
	wire n4808;
	wire n4809;
	wire n4810;
	wire n4811;
	wire n4812;
	wire n4813;
	wire n4814;
	wire n4815;
	wire n4816;
	wire n4817;
	wire n4818;
	wire n4819;
	wire n4820;
	wire n4821;
	wire n4822;
	wire n4823;
	wire n4824;
	wire n4825;
	wire n4826;
	wire n4827;
	wire n4828;
	wire n4829;
	wire n4830;
	wire n4831;
	wire n4832;
	wire n4833;
	wire n4834;
	wire n4835;
	wire n4836;
	wire n4837;
	wire n4838;
	wire n4839;
	wire n4840;
	wire n4841;
	wire n4842;
	wire n4843;
	wire n4844;
	wire n4845;
	wire n4846;
	wire n4847;
	wire n4848;
	wire n4849;
	wire n4850;
	wire n4851;
	wire n4852;
	wire n4853;
	wire n4854;
	wire n4855;
	wire n4856;
	wire n4857;
	wire n4858;
	wire n4859;
	wire n4860;
	wire n4861;
	wire n4862;
	wire n4863;
	wire n4864;
	wire n4865;
	wire n4866;
	wire n4867;
	wire n4868;
	wire n4869;
	wire n4870;
	wire n4871;
	wire n4872;
	wire n4873;
	wire n4874;
	wire n4875;
	wire n4876;
	wire n4877;
	wire n4878;
	wire n4879;
	wire n4880;
	wire n4881;
	wire n4882;
	wire n4883;
	wire n4884;
	wire n4885;
	wire n4886;
	wire n4887;
	wire n4888;
	wire n4889;
	wire n4890;
	wire n4891;
	wire n4892;
	wire n4894;
	wire n4895;
	wire n4896;
	wire n4897;
	wire n4898;
	wire n4899;
	wire n4900;
	wire n4901;
	wire n4902;
	wire n4903;
	wire n4904;
	wire n4905;
	wire n4906;
	wire n4907;
	wire n4908;
	wire n4909;
	wire n4910;
	wire n4911;
	wire n4912;
	wire n4913;
	wire n4914;
	wire n4915;
	wire n4916;
	wire n4917;
	wire n4918;
	wire n4919;
	wire n4920;
	wire n4921;
	wire n4922;
	wire n4923;
	wire n4924;
	wire n4925;
	wire n4926;
	wire n4927;
	wire n4928;
	wire n4929;
	wire n4930;
	wire n4931;
	wire n4932;
	wire n4933;
	wire n4934;
	wire n4935;
	wire n4936;
	wire n4937;
	wire n4938;
	wire n4939;
	wire n4940;
	wire n4941;
	wire n4942;
	wire n4943;
	wire n4944;
	wire n4945;
	wire n4946;
	wire n4947;
	wire n4948;
	wire n4949;
	wire n4950;
	wire n4951;
	wire n4952;
	wire n4953;
	wire n4954;
	wire n4955;
	wire n4956;
	wire n4957;
	wire n4958;
	wire n4959;
	wire n4960;
	wire n4961;
	wire n4962;
	wire n4963;
	wire n4964;
	wire n4965;
	wire n4966;
	wire n4967;
	wire n4968;
	wire n4969;
	wire n4970;
	wire n4971;
	wire n4972;
	wire n4973;
	wire n4974;
	wire n4975;
	wire n4976;
	wire n4977;
	wire n4978;
	wire n4979;
	wire n4980;
	wire n4981;
	wire n4982;
	wire n4983;
	wire n4984;
	wire n4985;
	wire n4986;
	wire n4987;
	wire n4988;
	wire n4989;
	wire n4990;
	wire n4991;
	wire n4992;
	wire n4993;
	wire n4994;
	wire n4995;
	wire n4996;
	wire n4997;
	wire n4998;
	wire n4999;
	wire n5000;
	wire n5001;
	wire n5002;
	wire n5003;
	wire n5004;
	wire n5005;
	wire n5006;
	wire n5007;
	wire n5008;
	wire n5009;
	wire n5010;
	wire n5011;
	wire n5012;
	wire n5013;
	wire n5014;
	wire n5015;
	wire n5016;
	wire n5017;
	wire n5018;
	wire n5019;
	wire n5020;
	wire n5021;
	wire n5022;
	wire n5023;
	wire n5024;
	wire n5025;
	wire n5026;
	wire n5027;
	wire n5028;
	wire n5029;
	wire n5030;
	wire n5031;
	wire n5032;
	wire n5033;
	wire n5034;
	wire n5035;
	wire n5036;
	wire n5037;
	wire n5038;
	wire n5039;
	wire n5040;
	wire n5041;
	wire n5042;
	wire n5043;
	wire n5044;
	wire n5045;
	wire n5046;
	wire n5047;
	wire n5048;
	wire n5049;
	wire n5050;
	wire n5051;
	wire n5052;
	wire n5053;
	wire n5054;
	wire n5055;
	wire n5056;
	wire n5057;
	wire n5058;
	wire n5059;
	wire n5060;
	wire n5061;
	wire n5062;
	wire n5063;
	wire n5064;
	wire n5065;
	wire n5066;
	wire n5067;
	wire n5068;
	wire n5069;
	wire n5070;
	wire n5071;
	wire n5072;
	wire n5073;
	wire n5074;
	wire n5075;
	wire n5076;
	wire n5077;
	wire n5078;
	wire n5079;
	wire n5080;
	wire n5081;
	wire n5082;
	wire n5083;
	wire n5084;
	wire n5085;
	wire n5086;
	wire n5087;
	wire n5088;
	wire n5089;
	wire n5090;
	wire n5091;
	wire n5092;
	wire n5093;
	wire n5094;
	wire n5095;
	wire n5096;
	wire n5097;
	wire n5098;
	wire n5099;
	wire n5100;
	wire n5101;
	wire n5102;
	wire n5103;
	wire n5104;
	wire n5105;
	wire n5107;
	wire n5108;
	wire n5109;
	wire n5110;
	wire n5111;
	wire n5112;
	wire n5113;
	wire n5114;
	wire n5115;
	wire n5116;
	wire n5117;
	wire n5118;
	wire n5121;
	wire n5122;
	wire n5123;
	wire n5124;
	wire n5125;
	wire n5126;
	wire n5127;
	wire n5128;
	wire n5129;
	wire n5130;
	wire n5131;
	wire n5132;
	wire n5134;
	wire n5135;
	wire n5136;
	wire n5137;
	wire n5138;
	wire n5139;
	wire n5140;
	wire n5141;
	wire n5142;
	wire n5143;
	wire n5144;
	wire n5145;
	wire n5146;
	wire n5147;
	wire n5148;
	wire n5149;
	wire n5150;
	wire n5151;
	wire n5152;
	wire n5153;
	wire n5154;
	wire n5155;
	wire n5156;
	wire n5157;
	wire n5158;
	wire n5159;
	wire n5160;
	wire n5161;
	wire n5162;
	wire n5163;
	wire n5164;
	wire n5165;
	wire n5166;
	wire n5167;
	wire n5168;
	wire n5169;
	wire n5170;
	wire n5171;
	wire n5172;
	wire n5173;
	wire n5174;
	wire n5175;
	wire n5176;
	wire n5177;
	wire n5178;
	wire n5179;
	wire n5180;
	wire n5181;
	wire n5182;
	wire n5183;
	wire n5184;
	wire n5185;
	wire n5186;
	wire n5187;
	wire n5188;
	wire n5189;
	wire n5190;
	wire n5191;
	wire n5192;
	wire n5193;
	wire n5194;
	wire n5195;
	wire n5196;
	wire n5197;
	wire n5198;
	wire n5199;
	wire n5200;
	wire n5201;
	wire n5202;
	wire n5203;
	wire n5204;
	wire n5205;
	wire n5206;
	wire n5207;
	wire n5208;
	wire n5209;
	wire n5210;
	wire n5211;
	wire n5212;
	wire n5213;
	wire n5214;
	wire n5215;
	wire n5216;
	wire n5217;
	wire n5218;
	wire n5219;
	wire n5220;
	wire n5221;
	wire n5222;
	wire n5223;
	wire n5224;
	wire n5225;
	wire n5226;
	wire n5227;
	wire n5228;
	wire n5229;
	wire n5230;
	wire n5231;
	wire n5232;
	wire n5233;
	wire n5234;
	wire n5235;
	wire n5236;
	wire n5237;
	wire n5238;
	wire n5239;
	wire n5240;
	wire n5241;
	wire n5242;
	wire n5243;
	wire n5244;
	wire n5245;
	wire n5246;
	wire n5247;
	wire n5248;
	wire n5249;
	wire n5250;
	wire n5251;
	wire n5252;
	wire n5253;
	wire n5254;
	wire n5255;
	wire n5256;
	wire n5257;
	wire n5259;
	wire n5260;
	wire n5261;
	wire n5262;
	wire n5263;
	wire n5264;
	wire n5265;
	wire n5266;
	wire n5267;
	wire n5268;
	wire n5269;
	wire n5270;
	wire n5271;
	wire n5272;
	wire n5273;
	wire n5274;
	wire n5275;
	wire n5276;
	wire n5277;
	wire n5278;
	wire n5279;
	wire n5280;
	wire n5281;
	wire n5282;
	wire n5283;
	wire n5284;
	wire n5285;
	wire n5286;
	wire n5287;
	wire n5288;
	wire n5289;
	wire n5290;
	wire n5291;
	wire n5292;
	wire n5293;
	wire n5294;
	wire n5295;
	wire n5296;
	wire n5297;
	wire n5298;
	wire n5299;
	wire n5300;
	wire n5301;
	wire n5302;
	wire n5303;
	wire n5304;
	wire n5305;
	wire n5306;
	wire n5307;
	wire n5308;
	wire n5309;
	wire n5310;
	wire n5311;
	wire n5312;
	wire n5313;
	wire n5314;
	wire n5315;
	wire n5316;
	wire n5317;
	wire n5318;
	wire n5319;
	wire n5320;
	wire n5321;
	wire n5322;
	wire n5323;
	wire n5324;
	wire n5325;
	wire n5326;
	wire n5327;
	wire n5328;
	wire n5329;
	wire n5330;
	wire n5331;
	wire n5332;
	wire n5333;
	wire n5334;
	wire n5335;
	wire n5336;
	wire n5337;
	wire n5338;
	wire n5339;
	wire n5340;
	wire n5341;
	wire n5342;
	wire n5343;
	wire n5344;
	wire n5345;
	wire n5346;
	wire n5347;
	wire n5348;
	wire n5349;
	wire n5350;
	wire n5351;
	wire n5352;
	wire n5353;
	wire n5354;
	wire n5355;
	wire n5356;
	wire n5357;
	wire n5358;
	wire n5359;
	wire n5360;
	wire n5361;
	wire n5362;
	wire n5363;
	wire n5364;
	wire n5365;
	wire n5366;
	wire n5367;
	wire n5368;
	wire n5369;
	wire n5370;
	wire n5371;
	wire n5372;
	wire n5373;
	wire n5374;
	wire n5375;
	wire n5376;
	wire n5377;
	wire n5378;
	wire n5379;
	wire n5380;
	wire n5381;
	wire n5382;
	wire n5383;
	wire n5384;
	wire n5385;
	wire n5386;
	wire n5387;
	wire n5388;
	wire n5389;
	wire n5390;
	wire n5391;
	wire n5392;
	wire n5393;
	wire n5394;
	wire n5395;
	wire n5396;
	wire n5397;
	wire n5398;
	wire n5399;
	wire n5400;
	wire n5401;
	wire n5402;
	wire n5403;
	wire n5404;
	wire n5405;
	wire n5406;
	wire n5407;
	wire n5408;
	wire n5409;
	wire n5410;
	wire n5411;
	wire n5412;
	wire n5413;
	wire n5414;
	wire n5415;
	wire n5416;
	wire n5417;
	wire n5418;
	wire n5419;
	wire n5420;
	wire n5421;
	wire n5422;
	wire n5423;
	wire n5424;
	wire n5425;
	wire n5426;
	wire n5427;
	wire n5428;
	wire n5429;
	wire n5430;
	wire n5431;
	wire n5432;
	wire n5433;
	wire n5434;
	wire n5435;
	wire n5436;
	wire n5437;
	wire n5438;
	wire n5439;
	wire n5440;
	wire n5441;
	wire n5442;
	wire n5443;
	wire n5444;
	wire n5445;
	wire n5446;
	wire n5447;
	wire n5448;
	wire n5449;
	wire n5450;
	wire n5451;
	wire n5452;
	wire n5453;
	wire n5454;
	wire n5455;
	wire n5456;
	wire n5457;
	wire n5458;
	wire n5459;
	wire n5460;
	wire n5461;
	wire n5462;
	wire n5463;
	wire n5464;
	wire n5465;
	wire n5466;
	wire n5467;
	wire n5468;
	wire n5469;
	wire n5470;
	wire n5471;
	wire n5472;
	wire n5473;
	wire n5474;
	wire n5475;
	wire n5476;
	wire n5477;
	wire n5478;
	wire n5479;
	wire n5480;
	wire n5481;
	wire n5482;
	wire n5483;
	wire n5484;
	wire n5485;
	wire n5486;
	wire n5487;
	wire n5488;
	wire n5489;
	wire n5490;
	wire n5491;
	wire n5492;
	wire n5493;
	wire n5494;
	wire n5495;
	wire n5496;
	wire n5497;
	wire n5498;
	wire n5499;
	wire n5500;
	wire n5501;
	wire n5502;
	wire n5503;
	wire n5504;
	wire n5505;
	wire n5506;
	wire n5507;
	wire n5508;
	wire n5509;
	wire n5510;
	wire n5511;
	wire n5512;
	wire n5513;
	wire n5514;
	wire n5515;
	wire n5516;
	wire n5517;
	wire n5518;
	wire n5519;
	wire n5520;
	wire n5521;
	wire n5522;
	wire n5523;
	wire n5524;
	wire n5525;
	wire n5526;
	wire n5527;
	wire n5528;
	wire n5529;
	wire n5530;
	wire n5531;
	wire n5532;
	wire n5533;
	wire n5534;
	wire n5535;
	wire n5536;
	wire n5537;
	wire n5538;
	wire n5539;
	wire n5540;
	wire n5541;
	wire n5542;
	wire n5543;
	wire n5544;
	wire n5545;
	wire n5546;
	wire n5547;
	wire n5548;
	wire n5549;
	wire n5550;
	wire n5551;
	wire n5552;
	wire n5553;
	wire n5554;
	wire n5555;
	wire n5556;
	wire n5557;
	wire n5558;
	wire n5559;
	wire n5560;
	wire n5561;
	wire n5562;
	wire n5563;
	wire n5564;
	wire n5565;
	wire n5566;
	wire n5567;
	wire n5568;
	wire n5569;
	wire n5570;
	wire n5571;
	wire n5572;
	wire n5573;
	wire n5574;
	wire n5575;
	wire n5576;
	wire n5577;
	wire n5578;
	wire n5579;
	wire n5580;
	wire n5581;
	wire n5582;
	wire n5583;
	wire n5584;
	wire n5585;
	wire n5586;
	wire n5587;
	wire n5588;
	wire n5589;
	wire n5590;
	wire n5591;
	wire n5592;
	wire n5593;
	wire n5594;
	wire n5595;
	wire n5597;
	wire n5598;
	wire n5599;
	wire n5600;
	wire n5601;
	wire n5602;
	wire n5603;
	wire n5604;
	wire n5605;
	wire n5606;
	wire n5607;
	wire n5608;
	wire n5609;
	wire n5610;
	wire n5611;
	wire n5612;
	wire n5613;
	wire n5614;
	wire n5615;
	wire n5616;
	wire n5617;
	wire n5618;
	wire n5619;
	wire n5620;
	wire n5621;
	wire n5622;
	wire n5623;
	wire n5624;
	wire n5625;
	wire n5626;
	wire n5627;
	wire n5628;
	wire n5629;
	wire n5630;
	wire n5631;
	wire n5632;
	wire n5633;
	wire n5634;
	wire n5635;
	wire n5636;
	wire n5637;
	wire n5638;
	wire n5639;
	wire n5640;
	wire n5641;
	wire n5642;
	wire n5643;
	wire n5644;
	wire n5645;
	wire n5646;
	wire n5647;
	wire n5648;
	wire n5649;
	wire n5650;
	wire n5651;
	wire n5652;
	wire n5653;
	wire n5654;
	wire n5655;
	wire n5656;
	wire n5657;
	wire n5658;
	wire n5659;
	wire n5660;
	wire n5661;
	wire n5662;
	wire n5663;
	wire n5664;
	wire n5665;
	wire n5666;
	wire n5667;
	wire n5668;
	wire n5669;
	wire n5670;
	wire n5671;
	wire n5672;
	wire n5673;
	wire n5674;
	wire n5675;
	wire n5676;
	wire n5677;
	wire n5678;
	wire n5679;
	wire n5680;
	wire n5681;
	wire n5682;
	wire n5683;
	wire n5684;
	wire n5685;
	wire n5686;
	wire n5687;
	wire n5688;
	wire n5689;
	wire n5690;
	wire n5691;
	wire n5692;
	wire n5693;
	wire n5694;
	wire n5695;
	wire n5696;
	wire n5697;
	wire n5698;
	wire n5699;
	wire n5700;
	wire n5701;
	wire n5702;
	wire n5703;
	wire n5704;
	wire n5705;
	wire n5706;
	wire n5707;
	wire n5708;
	wire n5709;
	wire n5710;
	wire n5711;
	wire n5712;
	wire n5713;
	wire n5714;
	wire n5715;
	wire n5716;
	wire n5717;
	wire n5718;
	wire n5719;
	wire n5720;
	wire n5721;
	wire n5722;
	wire n5723;
	wire n5724;
	wire n5725;
	wire n5726;
	wire n5727;
	wire n5728;
	wire n5729;
	wire n5730;
	wire n5731;
	wire n5732;
	wire n5733;
	wire n5734;
	wire n5735;
	wire n5736;
	wire n5737;
	wire n5738;
	wire n5739;
	wire n5740;
	wire n5741;
	wire n5742;
	wire n5743;
	wire n5744;
	wire n5745;
	wire n5746;
	wire n5747;
	wire n5748;
	wire n5749;
	wire n5750;
	wire n5751;
	wire n5752;
	wire n5753;
	wire n5754;
	wire n5755;
	wire n5756;
	wire n5757;
	wire n5758;
	wire n5759;
	wire n5760;
	wire n5761;
	wire n5762;
	wire n5763;
	wire n5764;
	wire n5765;
	wire n5766;
	wire n5767;
	wire n5768;
	wire n5769;
	wire n5770;
	wire n5771;
	wire n5772;
	wire n5773;
	wire n5774;
	wire n5775;
	wire n5776;
	wire n5777;
	wire n5778;
	wire n5779;
	wire n5780;
	wire n5781;
	wire n5782;
	wire n5783;
	wire n5784;
	wire n5785;
	wire n5786;
	wire n5787;
	wire n5788;
	wire n5789;
	wire n5790;
	wire n5791;
	wire n5792;
	wire n5793;
	wire n5794;
	wire n5795;
	wire n5796;
	wire n5797;
	wire n5798;
	wire n5799;
	wire n5800;
	wire n5801;
	wire n5802;
	wire n5803;
	wire n5804;
	wire n5805;
	wire n5806;
	wire n5807;
	wire n5808;
	wire n5809;
	wire n5810;
	wire n5811;
	wire n5812;
	wire n5813;
	wire n5814;
	wire n5815;
	wire n5816;
	wire n5817;
	wire n5818;
	wire n5819;
	wire n5820;
	wire n5821;
	wire n5822;
	wire n5823;
	wire n5824;
	wire n5826;
	wire n5827;
	wire n5828;
	wire n5829;
	wire n5830;
	wire n5831;
	wire n5832;
	wire n5833;
	wire n5834;
	wire n5835;
	wire n5836;
	wire n5837;
	wire n5840;
	wire n5841;
	wire n5842;
	wire n5843;
	wire n5844;
	wire n5845;
	wire n5846;
	wire n5847;
	wire n5848;
	wire n5849;
	wire n5850;
	wire n5851;
	wire n5852;
	wire n5853;
	wire n5854;
	wire n5856;
	wire n5857;
	wire n5858;
	wire n5859;
	wire n5860;
	wire n5861;
	wire n5862;
	wire n5863;
	wire n5864;
	wire n5865;
	wire n5866;
	wire n5867;
	wire n5868;
	wire n5869;
	wire n5870;
	wire n5871;
	wire n5872;
	wire n5873;
	wire n5874;
	wire n5875;
	wire n5876;
	wire n5877;
	wire n5878;
	wire n5879;
	wire n5880;
	wire n5881;
	wire n5882;
	wire n5883;
	wire n5884;
	wire n5885;
	wire n5886;
	wire n5887;
	wire n5888;
	wire n5889;
	wire n5890;
	wire n5891;
	wire n5892;
	wire n5893;
	wire n5894;
	wire n5895;
	wire n5896;
	wire n5897;
	wire n5898;
	wire n5899;
	wire n5900;
	wire n5901;
	wire n5902;
	wire n5903;
	wire n5904;
	wire n5905;
	wire n5906;
	wire n5907;
	wire n5908;
	wire n5909;
	wire n5910;
	wire n5911;
	wire n5912;
	wire n5913;
	wire n5914;
	wire n5915;
	wire n5916;
	wire n5917;
	wire n5918;
	wire n5919;
	wire n5920;
	wire n5921;
	wire n5922;
	wire n5923;
	wire n5924;
	wire n5925;
	wire n5926;
	wire n5927;
	wire n5928;
	wire n5929;
	wire n5930;
	wire n5931;
	wire n5932;
	wire n5933;
	wire n5934;
	wire n5935;
	wire n5936;
	wire n5937;
	wire n5938;
	wire n5939;
	wire n5940;
	wire n5941;
	wire n5942;
	wire n5943;
	wire n5944;
	wire n5945;
	wire n5946;
	wire n5947;
	wire n5948;
	wire n5949;
	wire n5950;
	wire n5951;
	wire n5952;
	wire n5953;
	wire n5954;
	wire n5955;
	wire n5956;
	wire n5957;
	wire n5958;
	wire n5959;
	wire n5960;
	wire n5961;
	wire n5962;
	wire n5963;
	wire n5964;
	wire n5965;
	wire n5966;
	wire n5967;
	wire n5968;
	wire n5969;
	wire n5970;
	wire n5971;
	wire n5972;
	wire n5973;
	wire n5974;
	wire n5975;
	wire n5976;
	wire n5977;
	wire n5978;
	wire n5979;
	wire n5980;
	wire n5981;
	wire n5982;
	wire n5983;
	wire n5984;
	wire n5985;
	wire n5986;
	wire n5987;
	wire n5989;
	wire n5990;
	wire n5991;
	wire n5992;
	wire n5993;
	wire n5994;
	wire n5995;
	wire n5996;
	wire n5997;
	wire n5998;
	wire n5999;
	wire n6000;
	wire n6001;
	wire n6002;
	wire n6003;
	wire n6004;
	wire n6005;
	wire n6006;
	wire n6007;
	wire n6008;
	wire n6009;
	wire n6010;
	wire n6011;
	wire n6012;
	wire n6013;
	wire n6014;
	wire n6015;
	wire n6016;
	wire n6017;
	wire n6018;
	wire n6019;
	wire n6020;
	wire n6021;
	wire n6022;
	wire n6023;
	wire n6024;
	wire n6025;
	wire n6026;
	wire n6027;
	wire n6028;
	wire n6029;
	wire n6030;
	wire n6031;
	wire n6032;
	wire n6033;
	wire n6034;
	wire n6035;
	wire n6036;
	wire n6037;
	wire n6038;
	wire n6039;
	wire n6040;
	wire n6041;
	wire n6042;
	wire n6043;
	wire n6044;
	wire n6045;
	wire n6046;
	wire n6047;
	wire n6048;
	wire n6049;
	wire n6050;
	wire n6051;
	wire n6052;
	wire n6053;
	wire n6054;
	wire n6055;
	wire n6056;
	wire n6057;
	wire n6058;
	wire n6059;
	wire n6060;
	wire n6061;
	wire n6062;
	wire n6063;
	wire n6064;
	wire n6065;
	wire n6066;
	wire n6067;
	wire n6068;
	wire n6069;
	wire n6070;
	wire n6071;
	wire n6072;
	wire n6073;
	wire n6074;
	wire n6075;
	wire n6076;
	wire n6077;
	wire n6078;
	wire n6079;
	wire n6080;
	wire n6081;
	wire n6082;
	wire n6083;
	wire n6084;
	wire n6085;
	wire n6086;
	wire n6087;
	wire n6088;
	wire n6089;
	wire n6090;
	wire n6091;
	wire n6092;
	wire n6093;
	wire n6094;
	wire n6095;
	wire n6096;
	wire n6097;
	wire n6098;
	wire n6099;
	wire n6100;
	wire n6101;
	wire n6102;
	wire n6103;
	wire n6104;
	wire n6105;
	wire n6106;
	wire n6107;
	wire n6108;
	wire n6109;
	wire n6110;
	wire n6111;
	wire n6112;
	wire n6113;
	wire n6114;
	wire n6115;
	wire n6116;
	wire n6117;
	wire n6118;
	wire n6119;
	wire n6120;
	wire n6121;
	wire n6122;
	wire n6123;
	wire n6124;
	wire n6125;
	wire n6126;
	wire n6127;
	wire n6128;
	wire n6129;
	wire n6130;
	wire n6131;
	wire n6132;
	wire n6133;
	wire n6134;
	wire n6135;
	wire n6136;
	wire n6137;
	wire n6138;
	wire n6139;
	wire n6140;
	wire n6141;
	wire n6142;
	wire n6143;
	wire n6144;
	wire n6145;
	wire n6146;
	wire n6147;
	wire n6148;
	wire n6149;
	wire n6150;
	wire n6151;
	wire n6152;
	wire n6153;
	wire n6154;
	wire n6155;
	wire n6156;
	wire n6157;
	wire n6158;
	wire n6159;
	wire n6160;
	wire n6161;
	wire n6162;
	wire n6163;
	wire n6164;
	wire n6165;
	wire n6166;
	wire n6167;
	wire n6168;
	wire n6169;
	wire n6170;
	wire n6171;
	wire n6172;
	wire n6173;
	wire n6174;
	wire n6175;
	wire n6176;
	wire n6177;
	wire n6178;
	wire n6179;
	wire n6180;
	wire n6181;
	wire n6182;
	wire n6183;
	wire n6184;
	wire n6185;
	wire n6186;
	wire n6187;
	wire n6188;
	wire n6189;
	wire n6190;
	wire n6191;
	wire n6192;
	wire n6193;
	wire n6194;
	wire n6195;
	wire n6196;
	wire n6197;
	wire n6198;
	wire n6199;
	wire n6200;
	wire n6201;
	wire n6202;
	wire n6204;
	wire n6205;
	wire n6206;
	wire n6207;
	wire n6208;
	wire n6209;
	wire n6210;
	wire n6211;
	wire n6212;
	wire n6213;
	wire n6214;
	wire n6215;
	wire n6216;
	wire n6217;
	wire n6218;
	wire n6219;
	wire n6220;
	wire n6221;
	wire n6222;
	wire n6223;
	wire n6224;
	wire n6225;
	wire n6226;
	wire n6227;
	wire n6228;
	wire n6229;
	wire n6230;
	wire n6231;
	wire n6232;
	wire n6233;
	wire n6234;
	wire n6235;
	wire n6236;
	wire n6237;
	wire n6238;
	wire n6239;
	wire n6240;
	wire n6241;
	wire n6242;
	wire n6243;
	wire n6244;
	wire n6245;
	wire n6246;
	wire n6247;
	wire n6248;
	wire n6249;
	wire n6250;
	wire n6251;
	wire n6252;
	wire n6253;
	wire n6254;
	wire n6255;
	wire n6256;
	wire n6257;
	wire n6258;
	wire n6259;
	wire n6260;
	wire n6261;
	wire n6262;
	wire n6263;
	wire n6264;
	wire n6265;
	wire n6266;
	wire n6267;
	wire n6268;
	wire n6269;
	wire n6270;
	wire n6271;
	wire n6272;
	wire n6273;
	wire n6274;
	wire n6275;
	wire n6276;
	wire n6277;
	wire n6278;
	wire n6279;
	wire n6280;
	wire n6281;
	wire n6282;
	wire n6283;
	wire n6284;
	wire n6285;
	wire n6286;
	wire n6287;
	wire n6288;
	wire n6289;
	wire n6290;
	wire n6291;
	wire n6292;
	wire n6293;
	wire n6294;
	wire n6295;
	wire n6296;
	wire n6297;
	wire n6298;
	wire n6299;
	wire n6300;
	wire n6301;
	wire n6302;
	wire n6303;
	wire n6304;
	wire n6305;
	wire n6306;
	wire n6307;
	wire n6308;
	wire n6309;
	wire n6310;
	wire n6311;
	wire n6312;
	wire n6313;
	wire n6314;
	wire n6315;
	wire n6316;
	wire n6317;
	wire n6318;
	wire n6319;
	wire n6320;
	wire n6321;
	wire n6322;
	wire n6323;
	wire n6324;
	wire n6325;
	wire n6326;
	wire n6327;
	wire n6328;
	wire n6329;
	wire n6330;
	wire n6331;
	wire n6332;
	wire n6333;
	wire n6334;
	wire n6335;
	wire n6336;
	wire n6337;
	wire n6338;
	wire n6339;
	wire n6340;
	wire n6341;
	wire n6342;
	wire n6343;
	wire n6344;
	wire n6345;
	wire n6348;
	wire n6349;
	wire n6351;
	wire n6352;
	wire n6353;
	wire n6354;
	wire n6355;
	wire n6357;
	wire n6358;
	wire n6359;
	wire n6360;
	wire n6361;
	wire n6362;
	wire n6363;
	wire n6364;
	wire n6365;
	wire n6366;
	wire n6367;
	wire n6368;
	wire n6369;
	wire n6370;
	wire n6371;
	wire n6372;
	wire n6373;
	wire n6374;
	wire n6375;
	wire n6376;
	wire n6377;
	wire n6378;
	wire n6379;
	wire n6380;
	wire n6381;
	wire n6382;
	wire n6383;
	wire n6384;
	wire n6385;
	wire n6386;
	wire n6387;
	wire n6388;
	wire n6389;
	wire n6390;
	wire n6391;
	wire n6392;
	wire n6393;
	wire n6394;
	wire n6395;
	wire n6396;
	wire n6397;
	wire n6398;
	wire n6399;
	wire n6400;
	wire n6401;
	wire n6402;
	wire n6403;
	wire n6404;
	wire n6405;
	wire n6406;
	wire n6407;
	wire n6408;
	wire n6409;
	wire n6410;
	wire n6411;
	wire n6412;
	wire n6413;
	wire n6414;
	wire n6415;
	wire n6416;
	wire n6417;
	wire n6418;
	wire n6419;
	wire n6420;
	wire n6421;
	wire n6422;
	wire n6423;
	wire n6424;
	wire n6425;
	wire n6426;
	wire n6427;
	wire n6428;
	wire n6429;
	wire n6430;
	wire n6431;
	wire n6432;
	wire n6433;
	wire n6434;
	wire n6435;
	wire n6436;
	wire n6437;
	wire n6438;
	wire n6439;
	wire n6440;
	wire n6441;
	wire n6442;
	wire n6443;
	wire n6444;
	wire n6445;
	wire n6446;
	wire n6447;
	wire n6448;
	wire n6449;
	wire n6450;
	wire n6451;
	wire n6452;
	wire n6453;
	wire n6454;
	wire n6455;
	wire n6456;
	wire n6457;
	wire n6458;
	wire n6459;
	wire n6460;
	wire n6461;
	wire n6462;
	wire n6463;
	wire n6464;
	wire n6465;
	wire n6466;
	wire n6467;
	wire n6468;
	wire n6469;
	wire n6470;
	wire n6471;
	wire n6472;
	wire n6473;
	wire n6474;
	wire n6475;
	wire n6476;
	wire n6477;
	wire n6478;
	wire n6479;
	wire n6480;
	wire n6481;
	wire n6482;
	wire n6483;
	wire n6484;
	wire n6485;
	wire n6486;
	wire n6487;
	wire n6488;
	wire n6489;
	wire n6490;
	wire n6491;
	wire n6492;
	wire n6493;
	wire n6494;
	wire n6495;
	wire n6496;
	wire n6497;
	wire n6498;
	wire n6499;
	wire n6500;
	wire n6501;
	wire n6502;
	wire n6503;
	wire n6504;
	wire n6505;
	wire n6506;
	wire n6507;
	wire n6508;
	wire n6509;
	wire n6510;
	wire n6511;
	wire n6512;
	wire n6513;
	wire n6514;
	wire n6515;
	wire n6516;
	wire n6517;
	wire n6518;
	wire n6519;
	wire n6520;
	wire n6521;
	wire n6522;
	wire n6523;
	wire n6524;
	wire n6525;
	wire n6526;
	wire n6527;
	wire n6528;
	wire n6529;
	wire n6530;
	wire n6531;
	wire n6532;
	wire n6533;
	wire n6534;
	wire n6535;
	wire n6536;
	wire n6537;
	wire n6538;
	wire n6539;
	wire n6540;
	wire n6541;
	wire n6542;
	wire n6543;
	wire n6544;
	wire n6545;
	wire n6546;
	wire n6547;
	wire n6548;
	wire n6549;
	wire n6550;
	wire n6551;
	wire n6552;
	wire n6553;
	wire n6554;
	wire n6555;
	wire n6556;
	wire n6557;
	wire n6558;
	wire n6559;
	wire n6560;
	wire n6561;
	wire n6562;
	wire n6563;
	wire n6564;
	wire n6565;
	wire n6566;
	wire n6567;
	wire n6568;
	wire n6569;
	wire n6570;
	wire n6571;
	wire n6572;
	wire n6573;
	wire n6574;
	wire n6575;
	wire n6576;
	wire n6577;
	wire n6578;
	wire n6579;
	wire n6580;
	wire n6581;
	wire n6582;
	wire n6583;
	wire n6584;
	wire n6585;
	wire n6586;
	wire n6587;
	wire n6588;
	wire n6589;
	wire n6590;
	wire n6591;
	wire n6592;
	wire n6593;
	wire n6594;
	wire n6595;
	wire n6596;
	wire n6597;
	wire n6598;
	wire n6599;
	wire n6600;
	wire n6601;
	wire n6602;
	wire n6603;
	wire n6604;
	wire n6606;
	wire n6607;
	wire n6608;
	wire n6609;
	wire n6610;
	wire n6611;
	wire n6612;
	wire n6613;
	wire n6614;
	wire n6615;
	wire n6616;
	wire n6617;
	wire n6618;
	wire n6619;
	wire n6620;
	wire n6621;
	wire n6622;
	wire n6623;
	wire n6624;
	wire n6625;
	wire n6626;
	wire n6627;
	wire n6628;
	wire n6629;
	wire n6630;
	wire n6631;
	wire n6632;
	wire n6633;
	wire n6634;
	wire n6635;
	wire n6636;
	wire n6637;
	wire n6638;
	wire n6639;
	wire n6640;
	wire n6641;
	wire n6642;
	wire n6643;
	wire n6644;
	wire n6645;
	wire n6646;
	wire n6647;
	wire n6648;
	wire n6649;
	wire n6650;
	wire n6651;
	wire n6652;
	wire n6653;
	wire n6654;
	wire n6655;
	wire n6656;
	wire n6657;
	wire n6658;
	wire n6659;
	wire n6660;
	wire n6661;
	wire n6662;
	wire n6663;
	wire n6664;
	wire n6665;
	wire n6666;
	wire n6667;
	wire n6668;
	wire n6669;
	wire n6670;
	wire n6671;
	wire n6672;
	wire n6673;
	wire n6674;
	wire n6675;
	wire n6676;
	wire n6677;
	wire n6678;
	wire n6679;
	wire n6680;
	wire n6681;
	wire n6682;
	wire n6683;
	wire n6684;
	wire n6685;
	wire n6686;
	wire n6687;
	wire n6688;
	wire n6689;
	wire n6690;
	wire n6691;
	wire n6692;
	wire n6693;
	wire n6694;
	wire n6695;
	wire n6696;
	wire n6697;
	wire n6698;
	wire n6699;
	wire n6700;
	wire n6701;
	wire n6702;
	wire n6703;
	wire n6704;
	wire n6705;
	wire n6706;
	wire n6707;
	wire n6708;
	wire n6709;
	wire n6710;
	wire n6711;
	wire n6712;
	wire n6713;
	wire n6714;
	wire n6715;
	wire n6716;
	wire n6717;
	wire n6718;
	wire n6719;
	wire n6720;
	wire n6721;
	wire n6722;
	wire n6723;
	wire n6724;
	wire n6725;
	wire n6726;
	wire n6727;
	wire n6728;
	wire n6729;
	wire n6730;
	wire n6731;
	wire n6732;
	wire n6733;
	wire n6734;
	wire n6735;
	wire n6736;
	wire n6737;
	wire n6738;
	wire n6739;
	wire n6740;
	wire n6741;
	wire n6742;
	wire n6743;
	wire n6744;
	wire n6745;
	wire n6746;
	wire n6747;
	wire n6748;
	wire n6749;
	wire n6750;
	wire n6751;
	wire n6752;
	wire n6753;
	wire n6754;
	wire n6755;
	wire n6756;
	wire n6757;
	wire n6758;
	wire n6759;
	wire n6760;
	wire n6761;
	wire n6762;
	wire n6763;
	wire n6764;
	wire n6765;
	wire n6766;
	wire n6767;
	wire n6768;
	wire n6769;
	wire n6770;
	wire n6771;
	wire n6772;
	wire n6773;
	wire n6774;
	wire n6775;
	wire n6776;
	wire n6777;
	wire n6778;
	wire n6779;
	wire n6780;
	wire n6781;
	wire n6782;
	wire n6783;
	wire n6784;
	wire n6785;
	wire n6786;
	wire n6787;
	wire n6788;
	wire n6789;
	wire n6790;
	wire n6791;
	wire n6792;
	wire n6793;
	wire n6794;
	wire n6795;
	wire n6796;
	wire n6797;
	wire n6798;
	wire n6799;
	wire n6800;
	wire n6801;
	wire n6802;
	wire n6803;
	wire n6804;
	wire n6805;
	wire n6806;
	wire n6807;
	wire n6808;
	wire n6809;
	wire n6810;
	wire n6811;
	wire n6812;
	wire n6813;
	wire n6814;
	wire n6815;
	wire n6816;
	wire n6817;
	wire n6818;
	wire n6819;
	wire n6820;
	wire n6821;
	wire n6822;
	wire n6823;
	wire n6824;
	wire n6825;
	wire n6826;
	wire n6827;
	wire n6828;
	wire n6829;
	wire n6830;
	wire n6831;
	wire n6832;
	wire n6833;
	wire n6834;
	wire n6835;
	wire n6836;
	wire n6837;
	wire n6838;
	wire n6839;
	wire n6840;
	wire n6841;
	wire n6842;
	wire n6843;
	wire n6844;
	wire n6845;
	wire n6846;
	wire n6847;
	wire n6848;
	wire n6849;
	wire n6850;
	wire n6851;
	wire n6852;
	wire n6853;
	wire n6854;
	wire n6855;
	wire n6856;
	wire n6857;
	wire n6858;
	wire n6859;
	wire n6860;
	wire n6861;
	wire n6862;
	wire n6863;
	wire n6864;
	wire n6865;
	wire n6866;
	wire n6867;
	wire n6868;
	wire n6869;
	wire n6870;
	wire n6871;
	wire n6872;
	wire n6873;
	wire n6874;
	wire n6875;
	wire n6876;
	wire n6877;
	wire n6878;
	wire n6879;
	wire n6880;
	wire n6881;
	wire n6882;
	wire n6883;
	wire n6884;
	wire n6885;
	wire n6886;
	wire n6887;
	wire n6888;
	wire n6889;
	wire n6890;
	wire n6891;
	wire n6892;
	wire n6893;
	wire n6894;
	wire n6895;
	wire n6896;
	wire n6897;
	wire n6898;
	wire n6899;
	wire n6900;
	wire n6901;
	wire n6902;
	wire n6903;
	wire n6904;
	wire n6905;
	wire n6906;
	wire n6907;
	wire n6908;
	wire n6909;
	wire n6910;
	wire n6911;
	wire n6912;
	wire n6913;
	wire n6914;
	wire n6915;
	wire n6916;
	wire n6917;
	wire n6918;
	wire n6919;
	wire n6920;
	wire n6921;
	wire n6922;
	wire n6923;
	wire n6924;
	wire n6925;
	wire n6926;
	wire n6927;
	wire n6928;
	wire n6929;
	wire n6930;
	wire n6931;
	wire n6932;
	wire n6933;
	wire n6934;
	wire n6935;
	wire n6936;
	wire n6937;
	wire n6938;
	wire n6939;
	wire n6940;
	wire n6941;
	wire n6942;
	wire n6943;
	wire n6944;
	wire n6945;
	wire n6946;
	wire n6947;
	wire n6948;
	wire n6949;
	wire n6950;
	wire n6951;
	wire n6952;
	wire n6953;
	wire n6954;
	wire n6955;
	wire n6956;
	wire n6957;
	wire n6958;
	wire n6959;
	wire n6960;
	wire n6961;
	wire n6962;
	wire n6963;
	wire n6964;
	wire n6965;
	wire n6966;
	wire n6967;
	wire n6968;
	wire n6969;
	wire n6970;
	wire n6971;
	wire n6972;
	wire n6973;
	wire n6974;
	wire n6975;
	wire n6976;
	wire n6977;
	wire n6978;
	wire n6979;
	wire n6980;
	wire n6981;
	wire n6982;
	wire n6983;
	wire n6984;
	wire n6985;
	wire n6986;
	wire n6987;
	wire n6988;
	wire n6989;
	wire n6990;
	wire n6991;
	wire n6992;
	wire n6993;
	wire n6994;
	wire n6995;
	wire n6996;
	wire n6997;
	wire n6998;
	wire n6999;
	wire n7000;
	wire n7001;
	wire n7002;
	wire n7003;
	wire n7004;
	wire n7005;
	wire n7006;
	wire n7007;
	wire n7008;
	wire n7009;
	wire n7010;
	wire n7011;
	wire n7012;
	wire n7013;
	wire n7014;
	wire n7015;
	wire n7016;
	wire n7017;
	wire n7018;
	wire n7019;
	wire n7020;
	wire n7021;
	wire n7022;
	wire n7023;
	wire n7024;
	wire n7025;
	wire n7026;
	wire n7027;
	wire n7028;
	wire n7029;
	wire n7030;
	wire n7031;
	wire n7032;
	wire n7033;
	wire n7034;
	wire n7035;
	wire n7036;
	wire n7037;
	wire n7038;
	wire n7039;
	wire n7040;
	wire n7041;
	wire n7042;
	wire n7043;
	wire n7044;
	wire n7045;
	wire n7046;
	wire n7047;
	wire n7048;
	wire n7049;
	wire n7050;
	wire n7051;
	wire n7052;
	wire n7053;
	wire n7054;
	wire n7055;
	wire n7056;
	wire n7057;
	wire n7058;
	wire n7059;
	wire n7060;
	wire n7061;
	wire n7062;
	wire n7063;
	wire n7064;
	wire n7065;
	wire n7066;
	wire n7067;
	wire n7068;
	wire n7069;
	wire n7070;
	wire n7071;
	wire n7072;
	wire n7073;
	wire n7074;
	wire n7075;
	wire n7076;
	wire n7077;
	wire n7078;
	wire n7079;
	wire n7080;
	wire n7081;
	wire n7082;
	wire n7083;
	wire n7084;
	wire n7085;
	wire n7086;
	wire n7087;
	wire n7088;
	wire n7089;
	wire n7090;
	wire n7091;
	wire n7092;
	wire n7093;
	wire n7094;
	wire n7095;
	wire n7096;
	wire n7097;
	wire n7098;
	wire n7099;
	wire n7100;
	wire n7101;
	wire n7102;
	wire n7103;
	wire n7104;
	wire n7105;
	wire n7106;
	wire n7107;
	wire n7108;
	wire n7109;
	wire n7110;
	wire n7111;
	wire n7112;
	wire n7113;
	wire n7114;
	wire n7115;
	wire n7116;
	wire n7117;
	wire n7118;
	wire n7119;
	wire n7120;
	wire n7121;
	wire n7122;
	wire n7123;
	wire n7124;
	wire n7125;
	wire n7126;
	wire n7127;
	wire n7128;
	wire n7129;
	wire n7130;
	wire n7131;
	wire n7132;
	wire n7133;
	wire n7134;
	wire n7135;
	wire n7136;
	wire n7137;
	wire n7138;
	wire n7139;
	wire n7140;
	wire n7141;
	wire n7142;
	wire n7143;
	wire n7145;
	wire n7146;
	wire n7147;
	wire n7148;
	wire n7149;
	wire n7150;
	wire n7151;
	wire n7152;
	wire n7153;
	wire n7154;
	wire n7155;
	wire n7156;
	wire n7157;
	wire n7158;
	wire n7159;
	wire n7160;
	wire n7161;
	wire n7162;
	wire n7163;
	wire n7164;
	wire n7165;
	wire n7166;
	wire n7167;
	wire n7168;
	wire n7169;
	wire n7170;
	wire n7171;
	wire n7172;
	wire n7173;
	wire n7174;
	wire n7175;
	wire n7176;
	wire n7177;
	wire n7178;
	wire n7179;
	wire n7180;
	wire n7181;
	wire n7182;
	wire n7183;
	wire n7184;
	wire n7185;
	wire n7186;
	wire n7187;
	wire n7188;
	wire n7189;
	wire n7190;
	wire n7191;
	wire n7192;
	wire n7193;
	wire n7194;
	wire n7195;
	wire n7196;
	wire n7197;
	wire n7198;
	wire n7199;
	wire n7200;
	wire n7201;
	wire n7202;
	wire n7203;
	wire n7204;
	wire n7205;
	wire n7206;
	wire n7207;
	wire n7208;
	wire n7209;
	wire n7210;
	wire n7211;
	wire n7212;
	wire n7213;
	wire n7214;
	wire n7215;
	wire n7216;
	wire n7217;
	wire n7218;
	wire n7219;
	wire n7220;
	wire n7221;
	wire n7222;
	wire n7223;
	wire n7224;
	wire n7225;
	wire n7226;
	wire n7227;
	wire n7228;
	wire n7229;
	wire n7230;
	wire n7231;
	wire n7232;
	wire n7233;
	wire n7234;
	wire n7235;
	wire n7236;
	wire n7237;
	wire n7238;
	wire n7239;
	wire n7240;
	wire n7241;
	wire n7242;
	wire n7243;
	wire n7244;
	wire n7245;
	wire n7246;
	wire n7247;
	wire n7248;
	wire n7249;
	wire n7250;
	wire n7251;
	wire n7252;
	wire n7253;
	wire n7254;
	wire n7255;
	wire n7256;
	wire n7257;
	wire n7258;
	wire n7259;
	wire n7260;
	wire n7261;
	wire n7262;
	wire n7263;
	wire n7264;
	wire n7265;
	wire n7266;
	wire n7267;
	wire n7268;
	wire n7269;
	wire n7270;
	wire n7271;
	wire n7272;
	wire n7273;
	wire n7274;
	wire n7275;
	wire n7276;
	wire n7277;
	wire n7278;
	wire n7279;
	wire n7280;
	wire n7281;
	wire n7282;
	wire n7283;
	wire n7284;
	wire n7285;
	wire n7286;
	wire n7287;
	wire n7288;
	wire n7289;
	wire n7290;
	wire n7291;
	wire n7292;
	wire n7293;
	wire n7294;
	wire n7295;
	wire n7296;
	wire n7297;
	wire n7298;
	wire n7299;
	wire n7300;
	wire n7301;
	wire n7302;
	wire n7303;
	wire n7304;
	wire n7305;
	wire n7306;
	wire n7307;
	wire n7308;
	wire n7309;
	wire n7310;
	wire n7311;
	wire n7312;
	wire n7313;
	wire n7314;
	wire n7315;
	wire n7316;
	wire n7317;
	wire n7318;
	wire n7319;
	wire n7320;
	wire n7321;
	wire n7322;
	wire n7323;
	wire n7324;
	wire n7325;
	wire n7326;
	wire n7327;
	wire n7328;
	wire n7329;
	wire n7330;
	wire n7331;
	wire n7332;
	wire n7333;
	wire n7334;
	wire n7335;
	wire n7336;
	wire n7337;
	wire n7338;
	wire n7339;
	wire n7340;
	wire n7341;
	wire n7342;
	wire n7343;
	wire n7344;
	wire n7345;
	wire n7346;
	wire n7347;
	wire n7348;
	wire n7349;
	wire n7350;
	wire n7351;
	wire n7352;
	wire n7353;
	wire n7354;
	wire n7355;
	wire n7356;
	wire n7357;
	wire n7358;
	wire n7359;
	wire n7360;
	wire n7361;
	wire n7362;
	wire n7363;
	wire n7364;
	wire n7365;
	wire n7366;
	wire n7367;
	wire n7368;
	wire n7369;
	wire n7370;
	wire n7371;
	wire n7372;
	wire n7373;
	wire n7374;
	wire n7375;
	wire n7376;
	wire n7377;
	wire n7378;
	wire n7379;
	wire n7380;
	wire n7381;
	wire n7382;
	wire n7383;
	wire n7384;
	wire n7385;
	wire n7386;
	wire n7387;
	wire n7388;
	wire n7389;
	wire n7390;
	wire n7391;
	wire n7392;
	wire n7393;
	wire n7394;
	wire n7395;
	wire n7396;
	wire n7397;
	wire n7398;
	wire n7399;
	wire n7400;
	wire n7401;
	wire n7402;
	wire n7403;
	wire n7404;
	wire n7405;
	wire n7406;
	wire n7407;
	wire n7408;
	wire n7409;
	wire n7410;
	wire n7411;
	wire n7412;
	wire n7413;
	wire n7414;
	wire n7415;
	wire n7417;
	wire n7418;
	wire n7419;
	wire n7420;
	wire n7421;
	wire n7422;
	wire n7423;
	wire n7424;
	wire n7425;
	wire n7426;
	wire n7427;
	wire n7428;
	wire n7429;
	wire n7430;
	wire n7431;
	wire n7432;
	wire n7433;
	wire n7434;
	wire n7435;
	wire n7436;
	wire n7437;
	wire n7438;
	wire n7439;
	wire n7440;
	wire n7441;
	wire n7442;
	wire n7443;
	wire n7444;
	wire n7445;
	wire n7446;
	wire n7447;
	wire n7448;
	wire n7449;
	wire n7450;
	wire n7451;
	wire n7452;
	wire n7453;
	wire n7454;
	wire n7455;
	wire n7456;
	wire n7457;
	wire n7458;
	wire n7459;
	wire n7460;
	wire n7461;
	wire n7462;
	wire n7463;
	wire n7464;
	wire n7465;
	wire n7466;
	wire n7467;
	wire n7468;
	wire n7469;
	wire n7470;
	wire n7471;
	wire n7472;
	wire n7473;
	wire n7474;
	wire n7475;
	wire n7476;
	wire n7477;
	wire n7478;
	wire n7479;
	wire n7480;
	wire n7481;
	wire n7482;
	wire n7483;
	wire n7484;
	wire n7485;
	wire n7486;
	wire n7487;
	wire n7488;
	wire n7489;
	wire n7490;
	wire n7491;
	wire n7492;
	wire n7493;
	wire n7494;
	wire n7495;
	wire n7496;
	wire n7497;
	wire n7498;
	wire n7499;
	wire n7500;
	wire n7501;
	wire n7502;
	wire n7503;
	wire n7504;
	wire n7505;
	wire n7506;
	wire n7507;
	wire n7508;
	wire n7509;
	wire n7510;
	wire n7511;
	wire n7512;
	wire n7513;
	wire n7514;
	wire n7515;
	wire n7516;
	wire n7517;
	wire n7518;
	wire n7519;
	wire n7520;
	wire n7521;
	wire n7522;
	wire n7523;
	wire n7524;
	wire n7525;
	wire n7526;
	wire n7527;
	wire n7528;
	wire n7529;
	wire n7530;
	wire n7531;
	wire n7532;
	wire n7533;
	wire n7534;
	wire n7535;
	wire n7536;
	wire n7537;
	wire n7538;
	wire n7539;
	wire n7540;
	wire n7541;
	wire n7542;
	wire n7543;
	wire n7544;
	wire n7545;
	wire n7546;
	wire n7547;
	wire n7548;
	wire n7549;
	wire n7550;
	wire n7551;
	wire n7552;
	wire n7553;
	wire n7554;
	wire n7555;
	wire n7556;
	wire n7557;
	wire n7558;
	wire n7559;
	wire n7560;
	wire n7561;
	wire n7562;
	wire n7563;
	wire n7564;
	wire n7565;
	wire n7566;
	wire n7567;
	wire n7568;
	wire n7569;
	wire n7570;
	wire n7571;
	wire n7572;
	wire n7573;
	wire n7574;
	wire n7575;
	wire n7576;
	wire n7577;
	wire n7578;
	wire n7579;
	wire n7580;
	wire n7581;
	wire n7582;
	wire n7583;
	wire n7584;
	wire n7585;
	wire n7586;
	wire n7587;
	wire n7588;
	wire n7589;
	wire n7590;
	wire n7591;
	wire n7592;
	wire n7593;
	wire n7594;
	wire n7595;
	wire n7596;
	wire n7597;
	wire n7598;
	wire n7599;
	wire n7600;
	wire n7601;
	wire n7602;
	wire n7603;
	wire n7604;
	wire n7605;
	wire n7606;
	wire n7607;
	wire n7608;
	wire n7609;
	wire n7610;
	wire n7611;
	wire n7612;
	wire n7613;
	wire n7614;
	wire n7615;
	wire n7616;
	wire n7617;
	wire n7618;
	wire n7619;
	wire n7620;
	wire n7621;
	wire n7622;
	wire n7623;
	wire n7624;
	wire n7625;
	wire n7626;
	wire n7627;
	wire n7628;
	wire n7629;
	wire n7630;
	wire n7631;
	wire n7632;
	wire n7633;
	wire n7634;
	wire n7635;
	wire n7636;
	wire n7637;
	wire n7638;
	wire n7639;
	wire n7640;
	wire n7641;
	wire n7642;
	wire n7643;
	wire n7644;
	wire n7645;
	wire n7646;
	wire n7647;
	wire n7648;
	wire n7649;
	wire n7650;
	wire n7651;
	wire n7652;
	wire n7653;
	wire n7654;
	wire n7655;
	wire n7656;
	wire n7657;
	wire n7658;
	wire n7659;
	wire n7660;
	wire n7661;
	wire n7662;
	wire n7663;
	wire n7664;
	wire n7665;
	wire n7666;
	wire n7667;
	wire n7668;
	wire n7669;
	wire n7670;
	wire n7671;
	wire n7672;
	wire n7673;
	wire n7674;
	wire n7675;
	wire n7676;
	wire n7677;
	wire n7678;
	wire n7679;
	wire n7680;
	wire n7681;
	wire n7682;
	wire n7683;
	wire n7684;
	wire n7685;
	wire n7686;
	wire n7687;
	wire n7688;
	wire n7689;
	wire n7690;
	wire n7691;
	wire n7692;
	wire n7693;
	wire n7694;
	wire n7695;
	wire n7696;
	wire n7697;
	wire n7698;
	wire n7699;
	wire n7700;
	wire n7701;
	wire n7702;
	wire n7703;
	wire n7704;
	wire n7705;
	wire n7706;
	wire n7707;
	wire n7708;
	wire n7709;
	wire n7710;
	wire n7711;
	wire n7712;
	wire n7713;
	wire n7714;
	wire n7715;
	wire n7716;
	wire n7717;
	wire n7718;
	wire n7719;
	wire n7720;
	wire n7721;
	wire n7722;
	wire n7723;
	wire n7724;
	wire n7725;
	wire n7726;
	wire n7727;
	wire n7728;
	wire n7729;
	wire n7730;
	wire n7731;
	wire n7732;
	wire n7733;
	wire n7734;
	wire n7735;
	wire n7736;
	wire n7737;
	wire n7738;
	wire n7739;
	wire n7740;
	wire n7741;
	wire n7742;
	wire n7743;
	wire n7744;
	wire n7745;
	wire n7746;
	wire n7747;
	wire n7748;
	wire n7749;
	wire n7750;
	wire n7751;
	wire n7752;
	wire n7753;
	wire n7754;
	wire n7755;
	wire n7756;
	wire n7757;
	wire n7758;
	wire n7759;
	wire n7760;
	wire n7761;
	wire n7762;
	wire n7763;
	wire n7764;
	wire n7765;
	wire n7766;
	wire n7767;
	wire n7768;
	wire n7769;
	wire n7770;
	wire n7771;
	wire n7772;
	wire n7773;
	wire n7774;
	wire n7775;
	wire n7776;
	wire n7777;
	wire n7778;
	wire n7779;
	wire n7780;
	wire n7781;
	wire n7782;
	wire n7783;
	wire n7784;
	wire n7785;
	wire n7786;
	wire n7787;
	wire n7788;
	wire n7789;
	wire n7790;
	wire n7791;
	wire n7792;
	wire n7793;
	wire n7794;
	wire n7795;
	wire n7796;
	wire n7797;
	wire n7798;
	wire n7799;
	wire n7800;
	wire n7801;
	wire n7802;
	wire n7803;
	wire n7804;
	wire n7805;
	wire n7806;
	wire n7807;
	wire n7808;
	wire n7809;
	wire n7810;
	wire n7811;
	wire n7812;
	wire n7813;
	wire n7814;
	wire n7815;
	wire n7816;
	wire n7817;
	wire n7818;
	wire n7819;
	wire n7820;
	wire n7821;
	wire n7822;
	wire n7823;
	wire n7824;
	wire n7825;
	wire n7826;
	wire n7827;
	wire n7828;
	wire n7829;
	wire n7830;
	wire n7831;
	wire n7832;
	wire n7833;
	wire n7834;
	wire n7835;
	wire n7836;
	wire n7837;
	wire n7838;
	wire n7839;
	wire n7840;
	wire n7841;
	wire n7842;
	wire n7843;
	wire n7844;
	wire n7845;
	wire n7846;
	wire n7847;
	wire n7848;
	wire n7849;
	wire n7850;
	wire n7851;
	wire n7852;
	wire n7853;
	wire n7854;
	wire n7855;
	wire n7856;
	wire n7857;
	wire n7858;
	wire n7859;
	wire n7860;
	wire n7861;
	wire n7862;
	wire n7863;
	wire n7864;
	wire n7865;
	wire n7866;
	wire n7867;
	wire n7868;
	wire n7869;
	wire n7870;
	wire n7871;
	wire n7872;
	wire n7873;
	wire n7874;
	wire n7875;
	wire n7876;
	wire n7877;
	wire n7878;
	wire n7879;
	wire n7880;
	wire n7881;
	wire n7882;
	wire n7883;
	wire n7884;
	wire n7885;
	wire n7886;
	wire n7887;
	wire n7888;
	wire n7889;
	wire n7890;
	wire n7891;
	wire n7892;
	wire n7893;
	wire n7894;
	wire n7895;
	wire n7896;
	wire n7897;
	wire n7898;
	wire n7899;
	wire n7900;
	wire n7901;
	wire n7902;
	wire n7903;
	wire n7904;
	wire n7905;
	wire n7906;
	wire n7907;
	wire n7908;
	wire n7909;
	wire n7910;
	wire n7911;
	wire n7912;
	wire n7913;
	wire n7914;
	wire n7915;
	wire n7916;
	wire n7917;
	wire n7918;
	wire n7919;
	wire n7920;
	wire n7921;
	wire n7922;
	wire n7923;
	wire n7924;
	wire n7925;
	wire n7926;
	wire n7927;
	wire n7928;
	wire n7929;
	wire n7930;
	wire n7931;
	wire n7932;
	wire n7933;
	wire n7934;
	wire n7935;
	wire n7936;
	wire n7937;
	wire n7938;
	wire n7939;
	wire n7940;
	wire n7941;
	wire n7942;
	wire n7943;
	wire n7944;
	wire n7945;
	wire n7946;
	wire n7947;
	wire n7948;
	wire n7949;
	wire n7950;
	wire n7951;
	wire n7952;
	wire n7953;
	wire n7954;
	wire n7955;
	wire n7956;
	wire n7957;
	wire n7958;
	wire n7959;
	wire n7960;
	wire n7961;
	wire n7962;
	wire n7963;
	wire n7964;
	wire n7965;
	wire n7966;
	wire n7967;
	wire n7968;
	wire n7969;
	wire n7970;
	wire n7971;
	wire n7972;
	wire n7973;
	wire n7974;
	wire n7975;
	wire n7976;
	wire n7977;
	wire n7978;
	wire n7979;
	wire n7980;
	wire n7981;
	wire n7982;
	wire n7983;
	wire n7984;
	wire n7985;
	wire n7986;
	wire n7987;
	wire n7989;
	wire n7990;
	wire n7991;
	wire n7992;
	wire n7993;
	wire n7994;
	wire n7995;
	wire n7996;
	wire n7997;
	wire n7998;
	wire n7999;
	wire n8000;
	wire n8001;
	wire n8002;
	wire n8003;
	wire n8004;
	wire n8005;
	wire n8006;
	wire n8007;
	wire n8008;
	wire n8009;
	wire n8010;
	wire n8011;
	wire n8012;
	wire n8013;
	wire n8014;
	wire n8015;
	wire n8016;
	wire n8017;
	wire n8018;
	wire n8019;
	wire n8020;
	wire n8021;
	wire n8022;
	wire n8023;
	wire n8024;
	wire n8025;
	wire n8026;
	wire n8027;
	wire n8028;
	wire n8029;
	wire n8030;
	wire n8031;
	wire n8032;
	wire n8033;
	wire n8034;
	wire n8035;
	wire n8036;
	wire n8037;
	wire n8038;
	wire n8039;
	wire n8040;
	wire n8041;
	wire n8042;
	wire n8043;
	wire n8044;
	wire n8045;
	wire n8046;
	wire n8047;
	wire n8048;
	wire n8049;
	wire n8050;
	wire n8051;
	wire n8052;
	wire n8053;
	wire n8054;
	wire n8055;
	wire n8056;
	wire n8057;
	wire n8058;
	wire n8059;
	wire n8060;
	wire n8061;
	wire n8062;
	wire n8063;
	wire n8064;
	wire n8065;
	wire n8066;
	wire n8067;
	wire n8068;
	wire n8069;
	wire n8070;
	wire n8071;
	wire n8072;
	wire n8073;
	wire n8074;
	wire n8075;
	wire n8076;
	wire n8077;
	wire n8078;
	wire n8079;
	wire n8080;
	wire n8081;
	wire n8082;
	wire n8083;
	wire n8084;
	wire n8085;
	wire n8086;
	wire n8087;
	wire n8088;
	wire n8089;
	wire n8090;
	wire n8091;
	wire n8092;
	wire n8093;
	wire n8094;
	wire n8095;
	wire n8096;
	wire n8097;
	wire n8098;
	wire n8099;
	wire n8100;
	wire n8101;
	wire n8102;
	wire n8103;
	wire n8104;
	wire n8105;
	wire n8106;
	wire n8107;
	wire n8108;
	wire n8109;
	wire n8110;
	wire n8111;
	wire n8112;
	wire n8113;
	wire n8114;
	wire n8115;
	wire n8116;
	wire n8117;
	wire n8118;
	wire n8119;
	wire n8120;
	wire n8121;
	wire n8122;
	wire n8123;
	wire n8124;
	wire n8125;
	wire n8126;
	wire n8127;
	wire n8128;
	wire n8129;
	wire n8130;
	wire n8131;
	wire n8132;
	wire n8133;
	wire n8134;
	wire n8135;
	wire n8136;
	wire n8137;
	wire n8138;
	wire n8139;
	wire n8140;
	wire n8141;
	wire n8142;
	wire n8143;
	wire n8144;
	wire n8145;
	wire n8146;
	wire n8147;
	wire n8148;
	wire n8149;
	wire n8150;
	wire n8151;
	wire n8152;
	wire n8153;
	wire n8154;
	wire n8155;
	wire n8156;
	wire n8157;
	wire n8158;
	wire n8159;
	wire n8160;
	wire n8161;
	wire n8162;
	wire n8163;
	wire n8164;
	wire n8165;
	wire n8166;
	wire n8167;
	wire n8168;
	wire n8169;
	wire n8170;
	wire n8171;
	wire n8172;
	wire n8173;
	wire n8174;
	wire n8175;
	wire n8176;
	wire n8177;
	wire n8178;
	wire n8179;
	wire n8180;
	wire n8181;
	wire n8182;
	wire n8183;
	wire n8184;
	wire n8185;
	wire n8186;
	wire n8187;
	wire n8188;
	wire n8189;
	wire n8190;
	wire n8191;
	wire n8192;
	wire n8193;
	wire n8194;
	wire n8195;
	wire n8196;
	wire n8197;
	wire n8198;
	wire n8199;
	wire n8200;
	wire n8201;
	wire n8202;
	wire n8203;
	wire n8204;
	wire n8205;
	wire n8206;
	wire n8207;
	wire n8208;
	wire n8209;
	wire n8210;
	wire n8211;
	wire n8212;
	wire n8213;
	wire n8214;
	wire n8215;
	wire n8216;
	wire n8217;
	wire n8218;
	wire n8219;
	wire n8220;
	wire n8221;
	wire n8222;
	wire n8223;
	wire n8224;
	wire n8225;
	wire n8226;
	wire n8227;
	wire n8228;
	wire n8229;
	wire n8230;
	wire n8231;
	wire n8232;
	wire n8233;
	wire n8234;
	wire n8235;
	wire n8236;
	wire n8237;
	wire n8238;
	wire n8239;
	wire n8240;
	wire n8241;
	wire n8242;
	wire n8243;
	wire n8244;
	wire n8245;
	wire n8246;
	wire n8247;
	wire n8248;
	wire n8249;
	wire n8250;
	wire n8251;
	wire n8252;
	wire n8253;
	wire n8254;
	wire n8255;
	wire n8256;
	wire n8257;
	wire n8258;
	wire n8259;
	wire n8260;
	wire n8261;
	wire n8262;
	wire n8263;
	wire n8264;
	wire n8265;
	wire n8266;
	wire n8267;
	wire n8268;
	wire n8269;
	wire n8270;
	wire n8271;
	wire n8272;
	wire n8274;
	wire n8275;
	wire n8276;
	wire n8277;
	wire n8278;
	wire n8279;
	wire n8280;
	wire n8281;
	wire n8282;
	wire n8283;
	wire n8284;
	wire n8285;
	wire n8286;
	wire n8287;
	wire n8288;
	wire n8289;
	wire n8290;
	wire n8291;
	wire n8292;
	wire n8293;
	wire n8294;
	wire n8295;
	wire n8296;
	wire n8297;
	wire n8298;
	wire n8299;
	wire n8300;
	wire n8301;
	wire n8302;
	wire n8303;
	wire n8304;
	wire n8305;
	wire n8306;
	wire n8307;
	wire n8308;
	wire n8309;
	wire n8310;
	wire n8311;
	wire n8312;
	wire n8313;
	wire n8314;
	wire n8315;
	wire n8316;
	wire n8317;
	wire n8318;
	wire n8319;
	wire n8320;
	wire n8321;
	wire n8322;
	wire n8323;
	wire n8324;
	wire n8325;
	wire n8326;
	wire n8327;
	wire n8328;
	wire n8329;
	wire n8330;
	wire n8331;
	wire n8332;
	wire n8333;
	wire n8334;
	wire n8335;
	wire n8336;
	wire n8337;
	wire n8338;
	wire n8339;
	wire n8340;
	wire n8341;
	wire n8342;
	wire n8343;
	wire n8344;
	wire n8345;
	wire n8346;
	wire n8347;
	wire n8348;
	wire n8349;
	wire n8350;
	wire n8351;
	wire n8352;
	wire n8353;
	wire n8354;
	wire n8355;
	wire n8356;
	wire n8357;
	wire n8358;
	wire n8359;
	wire n8360;
	wire n8361;
	wire n8362;
	wire n8363;
	wire n8364;
	wire n8365;
	wire n8366;
	wire n8367;
	wire n8368;
	wire n8369;
	wire n8370;
	wire n8371;
	wire n8372;
	wire n8373;
	wire n8374;
	wire n8375;
	wire n8376;
	wire n8377;
	wire n8378;
	wire n8379;
	wire n8380;
	wire n8381;
	wire n8382;
	wire n8383;
	wire n8384;
	wire n8385;
	wire n8386;
	wire n8387;
	wire n8388;
	wire n8389;
	wire n8390;
	wire n8391;
	wire n8392;
	wire n8393;
	wire n8394;
	wire n8395;
	wire n8396;
	wire n8397;
	wire n8398;
	wire n8399;
	wire n8400;
	wire n8401;
	wire n8402;
	wire n8403;
	wire n8404;
	wire n8405;
	wire n8406;
	wire n8407;
	wire n8408;
	wire n8409;
	wire n8410;
	wire n8411;
	wire n8412;
	wire n8413;
	wire n8414;
	wire n8415;
	wire n8416;
	wire n8417;
	wire n8418;
	wire n8419;
	wire n8420;
	wire n8421;
	wire n8422;
	wire n8423;
	wire n8424;
	wire n8425;
	wire n8426;
	wire n8427;
	wire n8428;
	wire n8429;
	wire n8430;
	wire n8431;
	wire n8432;
	wire n8433;
	wire n8434;
	wire n8435;
	wire n8436;
	wire n8437;
	wire n8438;
	wire n8439;
	wire n8440;
	wire n8441;
	wire n8442;
	wire n8443;
	wire n8444;
	wire n8445;
	wire n8446;
	wire n8447;
	wire n8448;
	wire n8449;
	wire n8450;
	wire n8451;
	wire n8452;
	wire n8453;
	wire n8454;
	wire n8455;
	wire n8456;
	wire n8457;
	wire n8458;
	wire n8459;
	wire n8460;
	wire n8461;
	wire n8462;
	wire n8463;
	wire n8464;
	wire n8465;
	wire n8466;
	wire n8467;
	wire n8468;
	wire n8469;
	wire n8470;
	wire n8471;
	wire n8472;
	wire n8473;
	wire n8474;
	wire n8475;
	wire n8476;
	wire n8477;
	wire n8478;
	wire n8479;
	wire n8480;
	wire n8481;
	wire n8482;
	wire n8483;
	wire n8484;
	wire n8485;
	wire n8486;
	wire n8487;
	wire n8488;
	wire n8489;
	wire n8490;
	wire n8491;
	wire n8492;
	wire n8493;
	wire n8494;
	wire n8495;
	wire n8496;
	wire n8497;
	wire n8498;
	wire n8499;
	wire n8500;
	wire n8501;
	wire n8502;
	wire n8503;
	wire n8504;
	wire n8505;
	wire n8506;
	wire n8507;
	wire n8508;
	wire n8509;
	wire n8510;
	wire n8511;
	wire n8512;
	wire n8513;
	wire n8514;
	wire n8515;
	wire n8516;
	wire n8517;
	wire n8518;
	wire n8519;
	wire n8520;
	wire n8521;
	wire n8522;
	wire n8523;
	wire n8524;
	wire n8525;
	wire n8526;
	wire n8527;
	wire n8528;
	wire n8529;
	wire n8530;
	wire n8531;
	wire n8532;
	wire n8533;
	wire n8534;
	wire n8535;
	wire n8536;
	wire n8537;
	wire n8538;
	wire n8539;
	wire n8540;
	wire n8541;
	wire n8542;
	wire n8543;
	wire n8544;
	wire n8545;
	wire n8546;
	wire n8547;
	wire n8548;
	wire n8549;
	wire n8550;
	wire n8551;
	wire n8552;
	wire n8553;
	wire n8554;
	wire n8555;
	wire n8556;
	wire n8557;
	wire n8558;
	wire n8559;
	wire n8560;
	wire n8561;
	wire n8562;
	wire n8563;
	wire n8564;
	wire n8565;
	wire n8566;
	wire n8567;
	wire n8568;
	wire n8569;
	wire n8570;
	wire n8571;
	wire n8572;
	wire n8573;
	wire n8574;
	wire n8575;
	wire n8576;
	wire n8577;
	wire n8578;
	wire n8579;
	wire n8580;
	wire n8581;
	wire n8582;
	wire n8583;
	wire n8584;
	wire n8585;
	wire n8586;
	wire n8587;
	wire n8588;
	wire n8589;
	wire n8590;
	wire n8591;
	wire n8592;
	wire n8593;
	wire n8594;
	wire n8595;
	wire n8596;
	wire n8597;
	wire n8598;
	wire n8599;
	wire n8600;
	wire n8601;
	wire n8602;
	wire n8603;
	wire n8604;
	wire n8605;
	wire n8606;
	wire n8607;
	wire n8608;
	wire n8609;
	wire n8610;
	wire n8611;
	wire n8612;
	wire n8613;
	wire n8614;
	wire n8615;
	wire n8616;
	wire n8617;
	wire n8618;
	wire n8619;
	wire n8620;
	wire n8621;
	wire n8622;
	wire n8623;
	wire n8624;
	wire n8625;
	wire n8626;
	wire n8627;
	wire n8628;
	wire n8629;
	wire n8630;
	wire n8631;
	wire n8632;
	wire n8633;
	wire n8634;
	wire n8635;
	wire n8636;
	wire n8637;
	wire n8638;
	wire n8639;
	wire n8640;
	wire n8641;
	wire n8642;
	wire n8643;
	wire n8644;
	wire n8645;
	wire n8646;
	wire n8647;
	wire n8648;
	wire n8649;
	wire n8650;
	wire n8651;
	wire n8652;
	wire n8653;
	wire n8654;
	wire n8655;
	wire n8656;
	wire n8657;
	wire n8658;
	wire n8659;
	wire n8660;
	wire n8661;
	wire n8662;
	wire n8663;
	wire n8664;
	wire n8665;
	wire n8666;
	wire n8667;
	wire n8668;
	wire n8669;
	wire n8670;
	wire n8671;
	wire n8672;
	wire n8673;
	wire n8674;
	wire n8675;
	wire n8676;
	wire n8677;
	wire n8678;
	wire n8679;
	wire n8680;
	wire n8681;
	wire n8682;
	wire n8683;
	wire n8684;
	wire n8685;
	wire n8686;
	wire n8687;
	wire n8688;
	wire n8689;
	wire n8690;
	wire n8691;
	wire n8692;
	wire n8693;
	wire n8694;
	wire n8695;
	wire n8696;
	wire n8697;
	wire n8698;
	wire n8699;
	wire n8700;
	wire n8701;
	wire n8702;
	wire n8703;
	wire n8704;
	wire n8705;
	wire n8707;
	wire n8708;
	wire n8709;
	wire n8710;
	wire n8711;
	wire n8712;
	wire n8713;
	wire n8714;
	wire n8715;
	wire n8716;
	wire n8717;
	wire n8718;
	wire n8719;
	wire n8720;
	wire n8721;
	wire n8722;
	wire n8723;
	wire n8724;
	wire n8725;
	wire n8726;
	wire n8727;
	wire n8728;
	wire n8729;
	wire n8730;
	wire n8731;
	wire n8732;
	wire n8733;
	wire n8734;
	wire n8735;
	wire n8736;
	wire n8737;
	wire n8738;
	wire n8739;
	wire n8740;
	wire n8741;
	wire n8742;
	wire n8743;
	wire n8744;
	wire n8745;
	wire n8746;
	wire n8747;
	wire n8748;
	wire n8749;
	wire n8750;
	wire n8751;
	wire n8752;
	wire n8753;
	wire n8754;
	wire n8755;
	wire n8756;
	wire n8757;
	wire n8758;
	wire n8759;
	wire n8760;
	wire n8761;
	wire n8762;
	wire n8763;
	wire n8764;
	wire n8765;
	wire n8766;
	wire n8767;
	wire n8768;
	wire n8769;
	wire n8770;
	wire n8771;
	wire n8772;
	wire n8773;
	wire n8774;
	wire n8775;
	wire n8776;
	wire n8777;
	wire n8778;
	wire n8779;
	wire n8780;
	wire n8781;
	wire n8782;
	wire n8783;
	wire n8784;
	wire n8785;
	wire n8786;
	wire n8787;
	wire n8788;
	wire n8789;
	wire n8790;
	wire n8791;
	wire n8792;
	wire n8793;
	wire n8794;
	wire n8795;
	wire n8796;
	wire n8797;
	wire n8798;
	wire n8799;
	wire n8800;
	wire n8801;
	wire n8802;
	wire n8803;
	wire n8804;
	wire n8805;
	wire n8806;
	wire n8807;
	wire n8808;
	wire n8809;
	wire n8810;
	wire n8811;
	wire n8812;
	wire n8813;
	wire n8814;
	wire n8815;
	wire n8816;
	wire n8817;
	wire n8818;
	wire n8819;
	wire n8820;
	wire n8821;
	wire n8822;
	wire n8823;
	wire n8824;
	wire n8825;
	wire n8826;
	wire n8827;
	wire n8828;
	wire n8829;
	wire n8830;
	wire n8831;
	wire n8832;
	wire n8833;
	wire n8834;
	wire n8835;
	wire n8836;
	wire n8837;
	wire n8838;
	wire n8839;
	wire n8840;
	wire n8841;
	wire n8842;
	wire n8843;
	wire n8844;
	wire n8845;
	wire n8846;
	wire n8847;
	wire n8848;
	wire n8849;
	wire n8850;
	wire n8851;
	wire n8852;
	wire n8853;
	wire n8854;
	wire n8855;
	wire n8856;
	wire n8857;
	wire n8858;
	wire n8859;
	wire n8860;
	wire n8861;
	wire n8862;
	wire n8863;
	wire n8864;
	wire n8865;
	wire n8866;
	wire n8867;
	wire n8868;
	wire n8869;
	wire n8870;
	wire n8871;
	wire n8872;
	wire n8873;
	wire n8874;
	wire n8875;
	wire n8876;
	wire n8877;
	wire n8878;
	wire n8882;
	wire n8883;
	wire n8884;
	wire n8885;
	wire n8886;
	wire n8887;
	wire n8888;
	wire n8890;
	wire n8891;
	wire n8892;
	wire n8893;
	wire n8894;
	wire n8895;
	wire n8896;
	wire n8897;
	wire n8898;
	wire n8899;
	wire n8900;
	wire n8901;
	wire n8902;
	wire n8903;
	wire n8904;
	wire n8905;
	wire n8906;
	wire n8907;
	wire n8908;
	wire n8909;
	wire n8910;
	wire n8911;
	wire n8912;
	wire n8913;
	wire n8914;
	wire n8915;
	wire n8916;
	wire n8917;
	wire n8918;
	wire n8919;
	wire n8920;
	wire n8921;
	wire n8922;
	wire n8923;
	wire n8924;
	wire n8925;
	wire n8926;
	wire n8927;
	wire n8928;
	wire n8929;
	wire n8930;
	wire n8931;
	wire n8932;
	wire n8933;
	wire n8934;
	wire n8935;
	wire n8936;
	wire n8937;
	wire n8938;
	wire n8939;
	wire n8940;
	wire n8941;
	wire n8942;
	wire n8943;
	wire n8944;
	wire n8945;
	wire n8946;
	wire n8947;
	wire n8948;
	wire n8949;
	wire n8950;
	wire n8951;
	wire n8952;
	wire n8953;
	wire n8954;
	wire n8955;
	wire n8956;
	wire n8957;
	wire n8958;
	wire n8959;
	wire n8960;
	wire n8961;
	wire n8962;
	wire n8963;
	wire n8964;
	wire n8965;
	wire n8966;
	wire n8967;
	wire n8968;
	wire n8969;
	wire n8970;
	wire n8971;
	wire n8972;
	wire n8973;
	wire n8974;
	wire n8975;
	wire n8976;
	wire n8977;
	wire n8978;
	wire n8979;
	wire n8980;
	wire n8981;
	wire n8982;
	wire n8983;
	wire n8984;
	wire n8985;
	wire n8986;
	wire n8987;
	wire n8988;
	wire n8989;
	wire n8990;
	wire n8991;
	wire n8992;
	wire n8993;
	wire n8994;
	wire n8995;
	wire n8996;
	wire n8997;
	wire n8998;
	wire n8999;
	wire n9000;
	wire n9001;
	wire n9002;
	wire n9003;
	wire n9004;
	wire n9005;
	wire n9006;
	wire n9007;
	wire n9008;
	wire n9009;
	wire n9010;
	wire n9011;
	wire n9012;
	wire n9013;
	wire n9014;
	wire n9015;
	wire n9016;
	wire n9017;
	wire n9018;
	wire n9019;
	wire n9020;
	wire n9021;
	wire n9022;
	wire n9023;
	wire n9024;
	wire n9025;
	wire n9026;
	wire n9027;
	wire n9028;
	wire n9029;
	wire n9030;
	wire n9031;
	wire n9032;
	wire n9033;
	wire n9034;
	wire n9035;
	wire n9036;
	wire n9037;
	wire n9038;
	wire n9039;
	wire n9040;
	wire n9041;
	wire n9042;
	wire n9043;
	wire n9044;
	wire n9045;
	wire n9046;
	wire n9047;
	wire n9048;
	wire n9049;
	wire n9050;
	wire n9051;
	wire n9052;
	wire n9053;
	wire n9054;
	wire n9055;
	wire n9056;
	wire n9057;
	wire n9058;
	wire n9059;
	wire n9060;
	wire n9061;
	wire n9062;
	wire n9063;
	wire n9064;
	wire n9065;
	wire n9066;
	wire n9067;
	wire n9068;
	wire n9069;
	wire n9070;
	wire n9071;
	wire n9072;
	wire n9073;
	wire n9074;
	wire n9075;
	wire n9076;
	wire n9077;
	wire n9078;
	wire n9079;
	wire n9080;
	wire n9081;
	wire n9082;
	wire n9083;
	wire n9084;
	wire n9085;
	wire n9086;
	wire n9087;
	wire n9088;
	wire n9089;
	wire n9090;
	wire n9091;
	wire n9092;
	wire n9093;
	wire n9094;
	wire n9095;
	wire n9096;
	wire n9097;
	wire n9098;
	wire n9099;
	wire n9100;
	wire n9101;
	wire n9102;
	wire n9103;
	wire n9104;
	wire n9105;
	wire n9106;
	wire n9107;
	wire n9108;
	wire n9109;
	wire n9110;
	wire n9111;
	wire n9112;
	wire n9113;
	wire n9114;
	wire n9115;
	wire n9116;
	wire n9117;
	wire n9118;
	wire n9119;
	wire n9120;
	wire n9121;
	wire n9122;
	wire n9123;
	wire n9124;
	wire n9125;
	wire n9126;
	wire n9127;
	wire n9128;
	wire n9129;
	wire n9130;
	wire n9131;
	wire n9132;
	wire n9133;
	wire n9134;
	wire n9135;
	wire n9136;
	wire n9137;
	wire n9138;
	wire n9139;
	wire n9140;
	wire n9141;
	wire n9142;
	wire n9143;
	wire n9144;
	wire n9145;
	wire n9146;
	wire n9147;
	wire n9148;
	wire n9149;
	wire n9150;
	wire n9151;
	wire n9152;
	wire n9153;
	wire n9154;
	wire n9155;
	wire n9156;
	wire n9157;
	wire n9158;
	wire n9159;
	wire n9160;
	wire n9161;
	wire n9162;
	wire n9163;
	wire n9164;
	wire n9165;
	wire n9166;
	wire n9167;
	wire n9168;
	wire n9169;
	wire n9170;
	wire n9171;
	wire n9172;
	wire n9173;
	wire n9174;
	wire n9175;
	wire n9176;
	wire n9177;
	wire n9178;
	wire n9179;
	wire n9180;
	wire n9181;
	wire n9182;
	wire n9184;
	wire n9185;
	wire n9186;
	wire n9187;
	wire n9188;
	wire n9189;
	wire n9190;
	wire n9191;
	wire n9192;
	wire n9193;
	wire n9194;
	wire n9195;
	wire n9196;
	wire n9197;
	wire n9198;
	wire n9199;
	wire n9200;
	wire n9201;
	wire n9202;
	wire n9203;
	wire n9204;
	wire n9205;
	wire n9206;
	wire n9207;
	wire n9208;
	wire n9209;
	wire n9210;
	wire n9211;
	wire n9212;
	wire n9213;
	wire n9214;
	wire n9215;
	wire n9216;
	wire n9217;
	wire n9218;
	wire n9219;
	wire n9220;
	wire n9221;
	wire n9222;
	wire n9223;
	wire n9224;
	wire n9225;
	wire n9226;
	wire n9227;
	wire n9228;
	wire n9229;
	wire n9230;
	wire n9231;
	wire n9232;
	wire n9233;
	wire n9234;
	wire n9235;
	wire n9236;
	wire n9237;
	wire n9238;
	wire n9239;
	wire n9240;
	wire n9241;
	wire n9242;
	wire n9243;
	wire n9244;
	wire n9245;
	wire n9246;
	wire n9247;
	wire n9248;
	wire n9249;
	wire n9250;
	wire n9251;
	wire n9252;
	wire n9253;
	wire n9254;
	wire n9255;
	wire n9256;
	wire n9257;
	wire n9258;
	wire n9259;
	wire n9260;
	wire n9261;
	wire n9262;
	wire n9263;
	wire n9264;
	wire n9265;
	wire n9266;
	wire n9267;
	wire n9268;
	wire n9269;
	wire n9270;
	wire n9271;
	wire n9272;
	wire n9273;
	wire n9274;
	wire n9275;
	wire n9276;
	wire n9277;
	wire n9278;
	wire n9279;
	wire n9280;
	wire n9281;
	wire n9282;
	wire n9283;
	wire n9284;
	wire n9285;
	wire n9286;
	wire n9287;
	wire n9288;
	wire n9289;
	wire n9290;
	wire n9291;
	wire n9292;
	wire n9293;
	wire n9294;
	wire n9295;
	wire n9296;
	wire n9297;
	wire n9298;
	wire n9299;
	wire n9300;
	wire n9301;
	wire n9302;
	wire n9303;
	wire n9304;
	wire n9305;
	wire n9306;
	wire n9307;
	wire n9308;
	wire n9309;
	wire n9310;
	wire n9311;
	wire n9312;
	wire n9313;
	wire n9314;
	wire n9315;
	wire n9316;
	wire n9317;
	wire n9318;
	wire n9319;
	wire n9320;
	wire n9321;
	wire n9322;
	wire n9323;
	wire n9324;
	wire n9325;
	wire n9326;
	wire n9327;
	wire n9328;
	wire n9329;
	wire n9330;
	wire n9331;
	wire n9332;
	wire n9333;
	wire n9334;
	wire n9335;
	wire n9336;
	wire n9337;
	wire n9338;
	wire n9339;
	wire n9340;
	wire n9341;
	wire n9342;
	wire n9343;
	wire n9344;
	wire n9345;
	wire n9346;
	wire n9347;
	wire n9348;
	wire n9349;
	wire n9350;
	wire n9351;
	wire n9352;
	wire n9353;
	wire n9354;
	wire n9355;
	wire n9356;
	wire n9357;
	wire n9358;
	wire n9359;
	wire n9360;
	wire n9361;
	wire n9362;
	wire n9363;
	wire n9364;
	wire n9365;
	wire n9366;
	wire n9367;
	wire n9368;
	wire n9369;
	wire n9370;
	wire n9371;
	wire n9372;
	wire n9373;
	wire n9374;
	wire n9375;
	wire n9376;
	wire n9377;
	wire n9378;
	wire n9379;
	wire n9380;
	wire n9381;
	wire n9382;
	wire n9383;
	wire n9384;
	wire n9385;
	wire n9386;
	wire n9387;
	wire n9388;
	wire n9389;
	wire n9390;
	wire n9391;
	wire n9392;
	wire n9393;
	wire n9394;
	wire n9395;
	wire n9396;
	wire n9397;
	wire n9398;
	wire n9399;
	wire n9400;
	wire n9401;
	wire n9402;
	wire n9403;
	wire n9404;
	wire n9405;
	wire n9406;
	wire n9407;
	wire n9408;
	wire n9409;
	wire n9410;
	wire n9411;
	wire n9412;
	wire n9413;
	wire n9414;
	wire n9415;
	wire n9416;
	wire n9417;
	wire n9418;
	wire n9419;
	wire n9420;
	wire n9421;
	wire n9422;
	wire n9423;
	wire n9424;
	wire n9425;
	wire n9426;
	wire n9427;
	wire n9428;
	wire n9429;
	wire n9430;
	wire n9431;
	wire n9432;
	wire n9433;
	wire n9434;
	wire n9435;
	wire n9436;
	wire n9437;
	wire n9438;
	wire n9439;
	wire n9440;
	wire n9441;
	wire n9442;
	wire n9443;
	wire n9444;
	wire n9445;
	wire n9446;
	wire n9447;
	wire n9448;
	wire n9449;
	wire n9450;
	wire n9451;
	wire n9452;
	wire n9453;
	wire n9454;
	wire n9455;
	wire n9456;
	wire n9457;
	wire n9458;
	wire n9459;
	wire n9460;
	wire n9461;
	wire n9462;
	wire n9463;
	wire n9464;
	wire n9465;
	wire n9466;
	wire n9467;
	wire n9468;
	wire n9469;
	wire n9470;
	wire n9471;
	wire n9472;
	wire n9473;
	wire n9474;
	wire n9475;
	wire n9476;
	wire n9477;
	wire n9478;
	wire n9479;
	wire n9480;
	wire n9481;
	wire n9482;
	wire n9483;
	wire n9484;
	wire n9485;
	wire n9486;
	wire n9487;
	wire n9488;
	wire n9489;
	wire n9490;
	wire n9491;
	wire n9492;
	wire n9493;
	wire n9494;
	wire n9495;
	wire n9496;
	wire n9497;
	wire n9498;
	wire n9499;
	wire n9500;
	wire n9501;
	wire n9502;
	wire n9503;
	wire n9504;
	wire n9505;
	wire n9506;
	wire n9507;
	wire n9508;
	wire n9509;
	wire n9510;
	wire n9511;
	wire n9512;
	wire n9513;
	wire n9514;
	wire n9515;
	wire n9516;
	wire n9517;
	wire n9518;
	wire n9519;
	wire n9520;
	wire n9521;
	wire n9522;
	wire n9523;
	wire n9524;
	wire n9525;
	wire n9526;
	wire n9527;
	wire n9528;
	wire n9529;
	wire n9530;
	wire n9531;
	wire n9532;
	wire n9533;
	wire n9534;
	wire n9535;
	wire n9536;
	wire n9537;
	wire n9538;
	wire n9539;
	wire n9540;
	wire n9541;
	wire n9542;
	wire n9543;
	wire n9544;
	wire n9545;
	wire n9546;
	wire n9547;
	wire n9548;
	wire n9549;
	wire n9550;
	wire n9551;
	wire n9552;
	wire n9553;
	wire n9554;
	wire n9555;
	wire n9556;
	wire n9557;
	wire n9558;
	wire n9559;
	wire n9560;
	wire n9561;
	wire n9562;
	wire n9563;
	wire n9564;
	wire n9565;
	wire n9566;
	wire n9567;
	wire n9568;
	wire n9569;
	wire n9570;
	wire n9571;
	wire n9572;
	wire n9573;
	wire n9574;
	wire n9575;
	wire n9576;
	wire n9577;
	wire n9578;
	wire n9579;
	wire n9580;
	wire n9581;
	wire n9582;
	wire n9583;
	wire n9584;
	wire n9585;
	wire n9586;
	wire n9587;
	wire n9588;
	wire n9589;
	wire n9590;
	wire n9591;
	wire n9592;
	wire n9593;
	wire n9594;
	wire n9595;
	wire n9596;
	wire n9597;
	wire n9598;
	wire n9599;
	wire n9600;
	wire n9601;
	wire n9602;
	wire n9603;
	wire n9604;
	wire n9605;
	wire n9606;
	wire n9607;
	wire n9608;
	wire n9609;
	wire n9610;
	wire n9611;
	wire n9612;
	wire n9613;
	wire n9614;
	wire n9615;
	wire n9616;
	wire n9617;
	wire n9618;
	wire n9619;
	wire n9620;
	wire n9621;
	wire n9622;
	wire n9623;
	wire n9624;
	wire n9625;
	wire n9626;
	wire n9627;
	wire n9628;
	wire n9629;
	wire n9630;
	wire n9631;
	wire n9632;
	wire n9633;
	wire n9634;
	wire n9635;
	wire n9636;
	wire n9637;
	wire n9638;
	wire n9639;
	wire n9640;
	wire n9641;
	wire n9642;
	wire n9643;
	wire n9644;
	wire n9645;
	wire n9646;
	wire n9647;
	wire n9648;
	wire n9649;
	wire n9650;
	wire n9651;
	wire n9652;
	wire n9653;
	wire n9654;
	wire n9655;
	wire n9656;
	wire n9657;
	wire n9658;
	wire n9659;
	wire n9660;
	wire n9661;
	wire n9662;
	wire n9663;
	wire n9664;
	wire n9665;
	wire n9666;
	wire n9667;
	wire n9668;
	wire n9669;
	wire n9670;
	wire n9671;
	wire n9672;
	wire n9673;
	wire n9674;
	wire n9675;
	wire n9676;
	wire n9677;
	wire n9678;
	wire n9679;
	wire n9680;
	wire n9681;
	wire n9682;
	wire n9683;
	wire n9684;
	wire n9685;
	wire n9686;
	wire n9687;
	wire n9688;
	wire n9689;
	wire n9690;
	wire n9691;
	wire n9692;
	wire n9693;
	wire n9694;
	wire n9695;
	wire n9696;
	wire n9697;
	wire n9698;
	wire n9699;
	wire n9700;
	wire n9701;
	wire n9702;
	wire n9703;
	wire n9704;
	wire n9705;
	wire n9706;
	wire n9707;
	wire n9708;
	wire n9709;
	wire n9710;
	wire n9711;
	wire n9712;
	wire n9713;
	wire n9714;
	wire n9715;
	wire n9716;
	wire n9717;
	wire n9718;
	wire n9719;
	wire n9720;
	wire n9721;
	wire n9722;
	wire n9723;
	wire n9724;
	wire n9725;
	wire n9726;
	wire n9727;
	wire n9728;
	wire n9729;
	wire n9730;
	wire n9731;
	wire n9732;
	wire n9733;
	wire n9734;
	wire n9735;
	wire n9736;
	wire n9737;
	wire n9738;
	wire n9739;
	wire n9740;
	wire n9741;
	wire n9742;
	wire n9743;
	wire n9744;
	wire n9745;
	wire n9746;
	wire n9747;
	wire n9748;
	wire n9749;
	wire n9750;
	wire n9751;
	wire n9752;
	wire n9753;
	wire n9754;
	wire n9755;
	wire n9756;
	wire n9757;
	wire n9758;
	wire n9759;
	wire n9760;
	wire n9761;
	wire n9762;
	wire n9763;
	wire n9764;
	wire n9765;
	wire n9766;
	wire n9767;
	wire n9768;
	wire n9769;
	wire n9770;
	wire n9771;
	wire n9772;
	wire n9773;
	wire n9774;
	wire n9775;
	wire n9776;
	wire n9777;
	wire n9778;
	wire n9779;
	wire n9780;
	wire n9781;
	wire n9782;
	wire n9783;
	wire n9784;
	wire n9785;
	wire n9786;
	wire n9787;
	wire n9788;
	wire n9789;
	wire n9790;
	wire n9791;
	wire n9792;
	wire n9793;
	wire n9794;
	wire n9795;
	wire n9796;
	wire n9797;
	wire n9798;
	wire n9799;
	wire n9800;
	wire n9801;
	wire n9802;
	wire n9803;
	wire n9804;
	wire n9805;
	wire n9806;
	wire n9807;
	wire n9808;
	wire n9809;
	wire n9810;
	wire n9811;
	wire n9812;
	wire n9813;
	wire n9814;
	wire n9815;
	wire n9816;
	wire n9817;
	wire n9818;
	wire n9819;
	wire n9820;
	wire n9821;
	wire n9822;
	wire n9824;
	wire n9825;
	wire n9826;
	wire n9827;
	wire n9828;
	wire n9829;
	wire n9830;
	wire n9831;
	wire n9832;
	wire n9833;
	wire n9834;
	wire n9835;
	wire n9836;
	wire n9837;
	wire n9838;
	wire n9839;
	wire n9840;
	wire n9841;
	wire n9842;
	wire n9843;
	wire n9844;
	wire n9845;
	wire n9846;
	wire n9847;
	wire n9848;
	wire n9849;
	wire n9850;
	wire n9851;
	wire n9852;
	wire n9853;
	wire n9854;
	wire n9855;
	wire n9856;
	wire n9857;
	wire n9858;
	wire n9859;
	wire n9860;
	wire n9861;
	wire n9862;
	wire n9863;
	wire n9864;
	wire n9865;
	wire n9866;
	wire n9867;
	wire n9868;
	wire n9869;
	wire n9870;
	wire n9871;
	wire n9872;
	wire n9873;
	wire n9874;
	wire n9875;
	wire n9876;
	wire n9877;
	wire n9878;
	wire n9879;
	wire n9880;
	wire n9881;
	wire n9882;
	wire n9883;
	wire n9884;
	wire n9885;
	wire n9886;
	wire n9887;
	wire n9888;
	wire n9889;
	wire n9890;
	wire n9891;
	wire n9892;
	wire n9893;
	wire n9894;
	wire n9895;
	wire n9896;
	wire n9897;
	wire n9898;
	wire n9899;
	wire n9900;
	wire n9901;
	wire n9902;
	wire n9903;
	wire n9904;
	wire n9905;
	wire n9906;
	wire n9907;
	wire n9908;
	wire n9909;
	wire n9910;
	wire n9911;
	wire n9912;
	wire n9913;
	wire n9914;
	wire n9915;
	wire n9916;
	wire n9917;
	wire n9918;
	wire n9919;
	wire n9920;
	wire n9921;
	wire n9922;
	wire n9923;
	wire n9924;
	wire n9925;
	wire n9926;
	wire n9927;
	wire n9928;
	wire n9929;
	wire n9930;
	wire n9931;
	wire n9932;
	wire n9933;
	wire n9934;
	wire n9935;
	wire n9936;
	wire n9937;
	wire n9938;
	wire n9939;
	wire n9940;
	wire n9941;
	wire n9942;
	wire n9943;
	wire n9944;
	wire n9945;
	wire n9946;
	wire n9947;
	wire n9948;
	wire n9949;
	wire n9950;
	wire n9951;
	wire n9952;
	wire n9953;
	wire n9954;
	wire n9955;
	wire n9956;
	wire n9957;
	wire n9958;
	wire n9959;
	wire n9960;
	wire n9961;
	wire n9962;
	wire n9963;
	wire n9964;
	wire n9965;
	wire n9966;
	wire n9967;
	wire n9968;
	wire n9969;
	wire n9970;
	wire n9971;
	wire n9972;
	wire n9973;
	wire n9974;
	wire n9975;
	wire n9976;
	wire n9977;
	wire n9978;
	wire n9979;
	wire n9980;
	wire n9981;
	wire n9982;
	wire n9983;
	wire n9984;
	wire n9985;
	wire n9986;
	wire n9987;
	wire n9988;
	wire n9989;
	wire n9990;
	wire n9991;
	wire n9992;
	wire n9993;
	wire n9994;
	wire n9995;
	wire n9996;
	wire n9997;
	wire n9998;
	wire n9999;
	wire n10000;
	wire n10001;
	wire n10002;
	wire n10003;
	wire n10004;
	wire n10005;
	wire n10006;
	wire n10007;
	wire n10008;
	wire n10009;
	wire n10010;
	wire n10011;
	wire n10012;
	wire n10013;
	wire n10014;
	wire n10015;
	wire n10016;
	wire n10017;
	wire n10018;
	wire n10019;
	wire n10020;
	wire n10021;
	wire n10022;
	wire n10023;
	wire n10024;
	wire n10025;
	wire n10026;
	wire n10027;
	wire n10028;
	wire n10029;
	wire n10030;
	wire n10031;
	wire n10032;
	wire n10033;
	wire n10034;
	wire n10035;
	wire n10036;
	wire n10037;
	wire n10038;
	wire n10039;
	wire n10040;
	wire n10041;
	wire n10042;
	wire n10043;
	wire n10044;
	wire n10045;
	wire n10046;
	wire n10047;
	wire n10048;
	wire n10049;
	wire n10050;
	wire n10051;
	wire n10052;
	wire n10053;
	wire n10054;
	wire n10055;
	wire n10056;
	wire n10057;
	wire n10058;
	wire n10059;
	wire n10060;
	wire n10061;
	wire n10062;
	wire n10063;
	wire n10064;
	wire n10065;
	wire n10066;
	wire n10067;
	wire n10068;
	wire n10069;
	wire n10070;
	wire n10071;
	wire n10072;
	wire n10073;
	wire n10074;
	wire n10075;
	wire n10076;
	wire n10077;
	wire n10078;
	wire n10079;
	wire n10080;
	wire n10081;
	wire n10082;
	wire n10083;
	wire n10084;
	wire n10085;
	wire n10086;
	wire n10087;
	wire n10088;
	wire n10089;
	wire n10090;
	wire n10091;
	wire n10092;
	wire n10093;
	wire n10094;
	wire n10095;
	wire n10096;
	wire n10097;
	wire n10098;
	wire n10099;
	wire n10100;
	wire n10101;
	wire n10102;
	wire n10103;
	wire n10104;
	wire n10105;
	wire n10106;
	wire n10107;
	wire n10108;
	wire n10109;
	wire n10110;
	wire n10111;
	wire n10112;
	wire n10113;
	wire n10114;
	wire n10115;
	wire n10116;
	wire n10117;
	wire n10118;
	wire n10119;
	wire n10120;
	wire n10121;
	wire n10122;
	wire n10123;
	wire n10124;
	wire n10125;
	wire n10126;
	wire n10127;
	wire n10128;
	wire n10129;
	wire n10130;
	wire n10131;
	wire n10132;
	wire n10134;
	wire n10135;
	wire n10136;
	wire n10137;
	wire n10138;
	wire n10139;
	wire n10140;
	wire n10141;
	wire n10142;
	wire n10143;
	wire n10144;
	wire n10145;
	wire n10146;
	wire n10147;
	wire n10148;
	wire n10149;
	wire n10150;
	wire n10151;
	wire n10152;
	wire n10153;
	wire n10154;
	wire n10155;
	wire n10156;
	wire n10157;
	wire n10158;
	wire n10159;
	wire n10160;
	wire n10161;
	wire n10162;
	wire n10163;
	wire n10164;
	wire n10165;
	wire n10166;
	wire n10167;
	wire n10168;
	wire n10169;
	wire n10170;
	wire n10171;
	wire n10172;
	wire n10173;
	wire n10174;
	wire n10175;
	wire n10176;
	wire n10177;
	wire n10178;
	wire n10179;
	wire n10180;
	wire n10181;
	wire n10182;
	wire n10183;
	wire n10184;
	wire n10185;
	wire n10186;
	wire n10187;
	wire n10188;
	wire n10189;
	wire n10190;
	wire n10191;
	wire n10192;
	wire n10193;
	wire n10194;
	wire n10195;
	wire n10196;
	wire n10197;
	wire n10198;
	wire n10199;
	wire n10200;
	wire n10201;
	wire n10202;
	wire n10203;
	wire n10204;
	wire n10205;
	wire n10206;
	wire n10207;
	wire n10208;
	wire n10209;
	wire n10210;
	wire n10211;
	wire n10212;
	wire n10213;
	wire n10214;
	wire n10215;
	wire n10216;
	wire n10217;
	wire n10218;
	wire n10219;
	wire n10220;
	wire n10221;
	wire n10222;
	wire n10223;
	wire n10224;
	wire n10225;
	wire n10226;
	wire n10227;
	wire n10228;
	wire n10229;
	wire n10230;
	wire n10231;
	wire n10232;
	wire n10233;
	wire n10234;
	wire n10235;
	wire n10236;
	wire n10237;
	wire n10238;
	wire n10239;
	wire n10240;
	wire n10241;
	wire n10242;
	wire n10243;
	wire n10244;
	wire n10245;
	wire n10246;
	wire n10247;
	wire n10248;
	wire n10249;
	wire n10250;
	wire n10251;
	wire n10252;
	wire n10253;
	wire n10254;
	wire n10255;
	wire n10256;
	wire n10257;
	wire n10258;
	wire n10259;
	wire n10260;
	wire n10261;
	wire n10262;
	wire n10263;
	wire n10264;
	wire n10265;
	wire n10266;
	wire n10267;
	wire n10268;
	wire n10269;
	wire n10270;
	wire n10271;
	wire n10272;
	wire n10273;
	wire n10274;
	wire n10275;
	wire n10276;
	wire n10277;
	wire n10278;
	wire n10279;
	wire n10280;
	wire n10281;
	wire n10282;
	wire n10283;
	wire n10284;
	wire n10285;
	wire n10286;
	wire n10287;
	wire n10288;
	wire n10289;
	wire n10290;
	wire n10291;
	wire n10292;
	wire n10293;
	wire n10294;
	wire n10295;
	wire n10296;
	wire n10297;
	wire n10298;
	wire n10299;
	wire n10300;
	wire n10301;
	wire n10302;
	wire n10303;
	wire n10304;
	wire n10305;
	wire n10306;
	wire n10307;
	wire n10308;
	wire n10309;
	wire n10310;
	wire n10311;
	wire n10312;
	wire n10313;
	wire n10314;
	wire n10315;
	wire n10316;
	wire n10317;
	wire n10318;
	wire n10319;
	wire n10320;
	wire n10321;
	wire n10322;
	wire n10323;
	wire n10324;
	wire n10325;
	wire n10326;
	wire n10327;
	wire n10328;
	wire n10329;
	wire n10330;
	wire n10331;
	wire n10332;
	wire n10333;
	wire n10334;
	wire n10335;
	wire n10336;
	wire n10337;
	wire n10338;
	wire n10339;
	wire n10340;
	wire n10341;
	wire n10342;
	wire n10343;
	wire n10344;
	wire n10345;
	wire n10346;
	wire n10347;
	wire n10348;
	wire n10349;
	wire n10350;
	wire n10351;
	wire n10352;
	wire n10353;
	wire n10354;
	wire n10355;
	wire n10356;
	wire n10357;
	wire n10358;
	wire n10359;
	wire n10360;
	wire n10361;
	wire n10362;
	wire n10363;
	wire n10364;
	wire n10365;
	wire n10366;
	wire n10367;
	wire n10368;
	wire n10369;
	wire n10370;
	wire n10371;
	wire n10372;
	wire n10373;
	wire n10374;
	wire n10375;
	wire n10376;
	wire n10377;
	wire n10378;
	wire n10379;
	wire n10380;
	wire n10381;
	wire n10382;
	wire n10383;
	wire n10384;
	wire n10385;
	wire n10386;
	wire n10387;
	wire n10388;
	wire n10389;
	wire n10390;
	wire n10391;
	wire n10392;
	wire n10393;
	wire n10394;
	wire n10395;
	wire n10396;
	wire n10397;
	wire n10398;
	wire n10399;
	wire n10400;
	wire n10401;
	wire n10402;
	wire n10403;
	wire n10404;
	wire n10405;
	wire n10406;
	wire n10407;
	wire n10408;
	wire n10409;
	wire n10410;
	wire n10411;
	wire n10412;
	wire n10413;
	wire n10414;
	wire n10415;
	wire n10416;
	wire n10417;
	wire n10418;
	wire n10419;
	wire n10420;
	wire n10421;
	wire n10422;
	wire n10423;
	wire n10424;
	wire n10425;
	wire n10426;
	wire n10427;
	wire n10428;
	wire n10429;
	wire n10430;
	wire n10431;
	wire n10432;
	wire n10433;
	wire n10434;
	wire n10435;
	wire n10436;
	wire n10437;
	wire n10438;
	wire n10439;
	wire n10440;
	wire n10441;
	wire n10442;
	wire n10443;
	wire n10444;
	wire n10445;
	wire n10446;
	wire n10447;
	wire n10448;
	wire n10449;
	wire n10450;
	wire n10451;
	wire n10452;
	wire n10453;
	wire n10454;
	wire n10455;
	wire n10456;
	wire n10457;
	wire n10458;
	wire n10459;
	wire n10460;
	wire n10461;
	wire n10462;
	wire n10463;
	wire n10464;
	wire n10465;
	wire n10466;
	wire n10467;
	wire n10468;
	wire n10469;
	wire n10470;
	wire n10471;
	wire n10472;
	wire n10473;
	wire n10474;
	wire n10475;
	wire n10476;
	wire n10477;
	wire n10478;
	wire n10479;
	wire n10480;
	wire n10481;
	wire n10482;
	wire n10483;
	wire n10484;
	wire n10485;
	wire n10486;
	wire n10487;
	wire n10488;
	wire n10489;
	wire n10490;
	wire n10491;
	wire n10492;
	wire n10493;
	wire n10494;
	wire n10495;
	wire n10496;
	wire n10497;
	wire n10498;
	wire n10499;
	wire n10500;
	wire n10501;
	wire n10502;
	wire n10503;
	wire n10504;
	wire n10505;
	wire n10506;
	wire n10507;
	wire n10508;
	wire n10509;
	wire n10510;
	wire n10511;
	wire n10512;
	wire n10513;
	wire n10514;
	wire n10515;
	wire n10516;
	wire n10517;
	wire n10518;
	wire n10519;
	wire n10520;
	wire n10521;
	wire n10522;
	wire n10523;
	wire n10524;
	wire n10525;
	wire n10526;
	wire n10527;
	wire n10528;
	wire n10529;
	wire n10530;
	wire n10531;
	wire n10532;
	wire n10533;
	wire n10534;
	wire n10535;
	wire n10536;
	wire n10537;
	wire n10538;
	wire n10539;
	wire n10540;
	wire n10541;
	wire n10542;
	wire n10543;
	wire n10544;
	wire n10545;
	wire n10546;
	wire n10547;
	wire n10548;
	wire n10549;
	wire n10550;
	wire n10551;
	wire n10552;
	wire n10553;
	wire n10554;
	wire n10555;
	wire n10556;
	wire n10557;
	wire n10558;
	wire n10559;
	wire n10560;
	wire n10561;
	wire n10562;
	wire n10563;
	wire n10564;
	wire n10565;
	wire n10566;
	wire n10567;
	wire n10568;
	wire n10569;
	wire n10570;
	wire n10571;
	wire n10572;
	wire n10573;
	wire n10574;
	wire n10575;
	wire n10576;
	wire n10577;
	wire n10578;
	wire n10579;
	wire n10580;
	wire n10581;
	wire n10582;
	wire n10583;
	wire n10584;
	wire n10585;
	wire n10586;
	wire n10587;
	wire n10588;
	wire n10589;
	wire n10590;
	wire n10591;
	wire n10592;
	wire n10593;
	wire n10594;
	wire n10595;
	wire n10596;
	wire n10597;
	wire n10598;
	wire n10599;
	wire n10600;
	wire n10601;
	wire n10602;
	wire n10603;
	wire n10604;
	wire n10605;
	wire n10606;
	wire n10607;
	wire n10608;
	wire n10609;
	wire n10610;
	wire n10611;
	wire n10612;
	wire n10613;
	wire n10614;
	wire n10615;
	wire n10616;
	wire n10617;
	wire n10618;
	wire n10619;
	wire n10620;
	wire n10621;
	wire n10622;
	wire n10623;
	wire n10624;
	wire n10625;
	wire n10626;
	wire n10627;
	wire n10628;
	wire n10629;
	wire n10630;
	wire n10631;
	wire n10632;
	wire n10633;
	wire n10634;
	wire n10635;
	wire n10636;
	wire n10637;
	wire n10638;
	wire n10639;
	wire n10640;
	wire n10641;
	wire n10642;
	wire n10643;
	wire n10644;
	wire n10645;
	wire n10646;
	wire n10647;
	wire n10648;
	wire n10649;
	wire n10650;
	wire n10651;
	wire n10652;
	wire n10653;
	wire n10654;
	wire n10655;
	wire n10656;
	wire n10657;
	wire n10658;
	wire n10659;
	wire n10660;
	wire n10661;
	wire n10662;
	wire n10663;
	wire n10664;
	wire n10665;
	wire n10666;
	wire n10667;
	wire n10668;
	wire n10669;
	wire n10670;
	wire n10671;
	wire n10672;
	wire n10673;
	wire n10674;
	wire n10675;
	wire n10676;
	wire n10677;
	wire n10678;
	wire n10679;
	wire n10680;
	wire n10681;
	wire n10682;
	wire n10683;
	wire n10684;
	wire n10685;
	wire n10686;
	wire n10687;
	wire n10688;
	wire n10689;
	wire n10690;
	wire n10691;
	wire n10692;
	wire n10693;
	wire n10694;
	wire n10695;
	wire n10696;
	wire n10697;
	wire n10698;
	wire n10699;
	wire n10700;
	wire n10701;
	wire n10702;
	wire n10703;
	wire n10704;
	wire n10705;
	wire n10706;
	wire n10707;
	wire n10708;
	wire n10709;
	wire n10710;
	wire n10711;
	wire n10712;
	wire n10713;
	wire n10714;
	wire n10715;
	wire n10716;
	wire n10717;
	wire n10718;
	wire n10719;
	wire n10720;
	wire n10721;
	wire n10722;
	wire n10723;
	wire n10724;
	wire n10725;
	wire n10726;
	wire n10727;
	wire n10728;
	wire n10729;
	wire n10730;
	wire n10731;
	wire n10732;
	wire n10733;
	wire n10734;
	wire n10735;
	wire n10736;
	wire n10737;
	wire n10738;
	wire n10739;
	wire n10740;
	wire n10741;
	wire n10742;
	wire n10743;
	wire n10744;
	wire n10745;
	wire n10746;
	wire n10747;
	wire n10748;
	wire n10749;
	wire n10750;
	wire n10751;
	wire n10752;
	wire n10753;
	wire n10754;
	wire n10755;
	wire n10756;
	wire n10757;
	wire n10758;
	wire n10759;
	wire n10760;
	wire n10761;
	wire n10762;
	wire n10763;
	wire n10764;
	wire n10765;
	wire n10766;
	wire n10767;
	wire n10768;
	wire n10769;
	wire n10770;
	wire n10771;
	wire n10772;
	wire n10773;
	wire n10774;
	wire n10775;
	wire n10776;
	wire n10777;
	wire n10778;
	wire n10779;
	wire n10780;
	wire n10781;
	wire n10782;
	wire n10783;
	wire n10784;
	wire n10785;
	wire n10786;
	wire n10787;
	wire n10788;
	wire n10789;
	wire n10790;
	wire n10791;
	wire n10792;
	wire n10793;
	wire n10794;
	wire n10795;
	wire n10796;
	wire n10797;
	wire n10798;
	wire n10799;
	wire n10800;
	wire n10801;
	wire n10802;
	wire n10803;
	wire n10805;
	wire n10806;
	wire n10807;
	wire n10808;
	wire n10809;
	wire n10810;
	wire n10811;
	wire n10812;
	wire n10813;
	wire n10814;
	wire n10815;
	wire n10816;
	wire n10817;
	wire n10818;
	wire n10819;
	wire n10820;
	wire n10821;
	wire n10822;
	wire n10823;
	wire n10824;
	wire n10825;
	wire n10826;
	wire n10827;
	wire n10828;
	wire n10829;
	wire n10830;
	wire n10831;
	wire n10832;
	wire n10833;
	wire n10834;
	wire n10835;
	wire n10836;
	wire n10837;
	wire n10838;
	wire n10839;
	wire n10840;
	wire n10841;
	wire n10842;
	wire n10843;
	wire n10844;
	wire n10845;
	wire n10846;
	wire n10847;
	wire n10848;
	wire n10849;
	wire n10850;
	wire n10851;
	wire n10852;
	wire n10853;
	wire n10854;
	wire n10855;
	wire n10856;
	wire n10857;
	wire n10858;
	wire n10859;
	wire n10860;
	wire n10861;
	wire n10862;
	wire n10863;
	wire n10864;
	wire n10865;
	wire n10866;
	wire n10867;
	wire n10868;
	wire n10869;
	wire n10870;
	wire n10871;
	wire n10872;
	wire n10873;
	wire n10874;
	wire n10875;
	wire n10876;
	wire n10877;
	wire n10878;
	wire n10879;
	wire n10880;
	wire n10881;
	wire n10882;
	wire n10883;
	wire n10884;
	wire n10885;
	wire n10886;
	wire n10887;
	wire n10888;
	wire n10889;
	wire n10890;
	wire n10891;
	wire n10892;
	wire n10893;
	wire n10894;
	wire n10895;
	wire n10896;
	wire n10897;
	wire n10898;
	wire n10899;
	wire n10900;
	wire n10901;
	wire n10902;
	wire n10903;
	wire n10904;
	wire n10905;
	wire n10906;
	wire n10907;
	wire n10908;
	wire n10909;
	wire n10910;
	wire n10911;
	wire n10912;
	wire n10913;
	wire n10914;
	wire n10915;
	wire n10916;
	wire n10917;
	wire n10918;
	wire n10919;
	wire n10920;
	wire n10921;
	wire n10922;
	wire n10923;
	wire n10924;
	wire n10925;
	wire n10926;
	wire n10927;
	wire n10928;
	wire n10929;
	wire n10930;
	wire n10931;
	wire n10932;
	wire n10933;
	wire n10934;
	wire n10935;
	wire n10936;
	wire n10937;
	wire n10938;
	wire n10939;
	wire n10940;
	wire n10941;
	wire n10942;
	wire n10943;
	wire n10944;
	wire n10945;
	wire n10946;
	wire n10947;
	wire n10948;
	wire n10949;
	wire n10950;
	wire n10951;
	wire n10952;
	wire n10953;
	wire n10954;
	wire n10955;
	wire n10956;
	wire n10957;
	wire n10958;
	wire n10959;
	wire n10960;
	wire n10961;
	wire n10962;
	wire n10963;
	wire n10964;
	wire n10965;
	wire n10966;
	wire n10967;
	wire n10968;
	wire n10969;
	wire n10970;
	wire n10971;
	wire n10972;
	wire n10973;
	wire n10974;
	wire n10975;
	wire n10976;
	wire n10977;
	wire n10978;
	wire n10979;
	wire n10980;
	wire n10981;
	wire n10982;
	wire n10983;
	wire n10984;
	wire n10985;
	wire n10986;
	wire n10987;
	wire n10988;
	wire n10989;
	wire n10990;
	wire n10991;
	wire n10992;
	wire n10993;
	wire n10994;
	wire n10995;
	wire n10996;
	wire n10997;
	wire n10998;
	wire n10999;
	wire n11000;
	wire n11001;
	wire n11002;
	wire n11003;
	wire n11004;
	wire n11005;
	wire n11006;
	wire n11007;
	wire n11008;
	wire n11009;
	wire n11010;
	wire n11011;
	wire n11012;
	wire n11013;
	wire n11014;
	wire n11015;
	wire n11016;
	wire n11017;
	wire n11018;
	wire n11019;
	wire n11020;
	wire n11021;
	wire n11022;
	wire n11023;
	wire n11024;
	wire n11025;
	wire n11026;
	wire n11027;
	wire n11028;
	wire n11029;
	wire n11030;
	wire n11031;
	wire n11032;
	wire n11033;
	wire n11034;
	wire n11035;
	wire n11036;
	wire n11037;
	wire n11038;
	wire n11039;
	wire n11040;
	wire n11041;
	wire n11042;
	wire n11043;
	wire n11044;
	wire n11045;
	wire n11046;
	wire n11047;
	wire n11048;
	wire n11049;
	wire n11050;
	wire n11051;
	wire n11052;
	wire n11053;
	wire n11054;
	wire n11055;
	wire n11056;
	wire n11057;
	wire n11058;
	wire n11059;
	wire n11060;
	wire n11061;
	wire n11062;
	wire n11063;
	wire n11064;
	wire n11065;
	wire n11066;
	wire n11067;
	wire n11068;
	wire n11069;
	wire n11070;
	wire n11071;
	wire n11072;
	wire n11073;
	wire n11074;
	wire n11075;
	wire n11076;
	wire n11077;
	wire n11078;
	wire n11079;
	wire n11080;
	wire n11081;
	wire n11082;
	wire n11083;
	wire n11084;
	wire n11085;
	wire n11086;
	wire n11087;
	wire n11088;
	wire n11089;
	wire n11090;
	wire n11091;
	wire n11092;
	wire n11093;
	wire n11094;
	wire n11095;
	wire n11096;
	wire n11097;
	wire n11098;
	wire n11099;
	wire n11100;
	wire n11101;
	wire n11102;
	wire n11103;
	wire n11104;
	wire n11105;
	wire n11106;
	wire n11107;
	wire n11108;
	wire n11109;
	wire n11110;
	wire n11111;
	wire n11112;
	wire n11113;
	wire n11114;
	wire n11115;
	wire n11116;
	wire n11117;
	wire n11118;
	wire n11119;
	wire n11120;
	wire n11121;
	wire n11122;
	wire n11123;
	wire n11124;
	wire n11125;
	wire n11126;
	wire n11127;
	wire n11128;
	wire n11129;
	wire n11130;
	wire n11131;
	wire n11132;
	wire n11133;
	wire n11134;
	wire n11135;
	wire n11137;
	wire n11138;
	wire n11139;
	wire n11140;
	wire n11141;
	wire n11142;
	wire n11143;
	wire n11144;
	wire n11145;
	wire n11146;
	wire n11147;
	wire n11148;
	wire n11149;
	wire n11150;
	wire n11151;
	wire n11152;
	wire n11153;
	wire n11154;
	wire n11155;
	wire n11156;
	wire n11157;
	wire n11158;
	wire n11159;
	wire n11160;
	wire n11161;
	wire n11162;
	wire n11163;
	wire n11164;
	wire n11165;
	wire n11166;
	wire n11167;
	wire n11168;
	wire n11169;
	wire n11170;
	wire n11171;
	wire n11172;
	wire n11173;
	wire n11174;
	wire n11175;
	wire n11176;
	wire n11177;
	wire n11178;
	wire n11179;
	wire n11180;
	wire n11181;
	wire n11182;
	wire n11183;
	wire n11184;
	wire n11185;
	wire n11186;
	wire n11187;
	wire n11188;
	wire n11189;
	wire n11190;
	wire n11191;
	wire n11192;
	wire n11193;
	wire n11194;
	wire n11195;
	wire n11196;
	wire n11197;
	wire n11198;
	wire n11199;
	wire n11200;
	wire n11201;
	wire n11202;
	wire n11203;
	wire n11204;
	wire n11205;
	wire n11206;
	wire n11207;
	wire n11208;
	wire n11209;
	wire n11210;
	wire n11211;
	wire n11212;
	wire n11213;
	wire n11214;
	wire n11215;
	wire n11216;
	wire n11217;
	wire n11218;
	wire n11219;
	wire n11220;
	wire n11221;
	wire n11222;
	wire n11223;
	wire n11224;
	wire n11225;
	wire n11226;
	wire n11227;
	wire n11228;
	wire n11229;
	wire n11230;
	wire n11231;
	wire n11232;
	wire n11233;
	wire n11234;
	wire n11235;
	wire n11236;
	wire n11237;
	wire n11238;
	wire n11239;
	wire n11240;
	wire n11241;
	wire n11242;
	wire n11243;
	wire n11244;
	wire n11245;
	wire n11246;
	wire n11247;
	wire n11248;
	wire n11249;
	wire n11250;
	wire n11251;
	wire n11252;
	wire n11253;
	wire n11254;
	wire n11255;
	wire n11256;
	wire n11257;
	wire n11258;
	wire n11259;
	wire n11260;
	wire n11261;
	wire n11262;
	wire n11263;
	wire n11264;
	wire n11265;
	wire n11266;
	wire n11267;
	wire n11268;
	wire n11269;
	wire n11270;
	wire n11271;
	wire n11272;
	wire n11273;
	wire n11274;
	wire n11275;
	wire n11276;
	wire n11277;
	wire n11278;
	wire n11279;
	wire n11280;
	wire n11281;
	wire n11282;
	wire n11283;
	wire n11284;
	wire n11285;
	wire n11286;
	wire n11287;
	wire n11288;
	wire n11289;
	wire n11290;
	wire n11291;
	wire n11292;
	wire n11293;
	wire n11294;
	wire n11295;
	wire n11296;
	wire n11297;
	wire n11298;
	wire n11299;
	wire n11300;
	wire n11301;
	wire n11302;
	wire n11303;
	wire n11304;
	wire n11305;
	wire n11306;
	wire n11307;
	wire n11308;
	wire n11309;
	wire n11310;
	wire n11311;
	wire n11312;
	wire n11313;
	wire n11314;
	wire n11315;
	wire n11316;
	wire n11317;
	wire n11318;
	wire n11319;
	wire n11320;
	wire n11321;
	wire n11322;
	wire n11323;
	wire n11324;
	wire n11325;
	wire n11326;
	wire n11327;
	wire n11328;
	wire n11329;
	wire n11330;
	wire n11331;
	wire n11332;
	wire n11333;
	wire n11334;
	wire n11335;
	wire n11336;
	wire n11337;
	wire n11338;
	wire n11339;
	wire n11340;
	wire n11341;
	wire n11342;
	wire n11343;
	wire n11344;
	wire n11345;
	wire n11346;
	wire n11347;
	wire n11348;
	wire n11349;
	wire n11350;
	wire n11351;
	wire n11352;
	wire n11353;
	wire n11354;
	wire n11355;
	wire n11356;
	wire n11357;
	wire n11358;
	wire n11359;
	wire n11360;
	wire n11361;
	wire n11362;
	wire n11363;
	wire n11364;
	wire n11365;
	wire n11366;
	wire n11367;
	wire n11368;
	wire n11369;
	wire n11370;
	wire n11371;
	wire n11372;
	wire n11373;
	wire n11374;
	wire n11375;
	wire n11376;
	wire n11377;
	wire n11378;
	wire n11379;
	wire n11380;
	wire n11381;
	wire n11382;
	wire n11383;
	wire n11384;
	wire n11385;
	wire n11386;
	wire n11387;
	wire n11388;
	wire n11389;
	wire n11390;
	wire n11391;
	wire n11392;
	wire n11393;
	wire n11394;
	wire n11395;
	wire n11396;
	wire n11397;
	wire n11398;
	wire n11399;
	wire n11400;
	wire n11401;
	wire n11402;
	wire n11403;
	wire n11404;
	wire n11405;
	wire n11406;
	wire n11407;
	wire n11408;
	wire n11409;
	wire n11410;
	wire n11411;
	wire n11412;
	wire n11413;
	wire n11414;
	wire n11415;
	wire n11416;
	wire n11417;
	wire n11418;
	wire n11419;
	wire n11420;
	wire n11421;
	wire n11422;
	wire n11423;
	wire n11424;
	wire n11425;
	wire n11426;
	wire n11427;
	wire n11428;
	wire n11429;
	wire n11430;
	wire n11431;
	wire n11432;
	wire n11433;
	wire n11434;
	wire n11435;
	wire n11436;
	wire n11437;
	wire n11438;
	wire n11439;
	wire n11440;
	wire n11441;
	wire n11442;
	wire n11443;
	wire n11444;
	wire n11445;
	wire n11446;
	wire n11447;
	wire n11448;
	wire n11449;
	wire n11450;
	wire n11451;
	wire n11452;
	wire n11453;
	wire n11454;
	wire n11455;
	wire n11456;
	wire n11457;
	wire n11458;
	wire n11459;
	wire n11460;
	wire n11461;
	wire n11462;
	wire n11463;
	wire n11464;
	wire n11465;
	wire n11466;
	wire n11467;
	wire n11468;
	wire n11469;
	wire n11470;
	wire n11471;
	wire n11472;
	wire n11473;
	wire n11474;
	wire n11475;
	wire n11476;
	wire n11477;
	wire n11478;
	wire n11479;
	wire n11480;
	wire n11481;
	wire n11482;
	wire n11483;
	wire n11484;
	wire n11485;
	wire n11486;
	wire n11487;
	wire n11488;
	wire n11489;
	wire n11490;
	wire n11491;
	wire n11492;
	wire n11493;
	wire n11494;
	wire n11495;
	wire n11496;
	wire n11497;
	wire n11498;
	wire n11499;
	wire n11500;
	wire n11501;
	wire n11502;
	wire n11503;
	wire n11504;
	wire n11505;
	wire n11506;
	wire n11507;
	wire n11508;
	wire n11509;
	wire n11510;
	wire n11511;
	wire n11512;
	wire n11513;
	wire n11514;
	wire n11515;
	wire n11516;
	wire n11517;
	wire n11518;
	wire n11519;
	wire n11520;
	wire n11521;
	wire n11522;
	wire n11523;
	wire n11524;
	wire n11525;
	wire n11526;
	wire n11527;
	wire n11528;
	wire n11529;
	wire n11530;
	wire n11531;
	wire n11532;
	wire n11533;
	wire n11534;
	wire n11535;
	wire n11536;
	wire n11537;
	wire n11538;
	wire n11539;
	wire n11540;
	wire n11541;
	wire n11542;
	wire n11543;
	wire n11544;
	wire n11545;
	wire n11546;
	wire n11547;
	wire n11548;
	wire n11549;
	wire n11550;
	wire n11551;
	wire n11552;
	wire n11553;
	wire n11554;
	wire n11555;
	wire n11556;
	wire n11557;
	wire n11558;
	wire n11559;
	wire n11560;
	wire n11561;
	wire n11562;
	wire n11563;
	wire n11564;
	wire n11565;
	wire n11566;
	wire n11567;
	wire n11568;
	wire n11569;
	wire n11570;
	wire n11571;
	wire n11572;
	wire n11573;
	wire n11574;
	wire n11575;
	wire n11576;
	wire n11577;
	wire n11578;
	wire n11579;
	wire n11580;
	wire n11581;
	wire n11582;
	wire n11583;
	wire n11584;
	wire n11585;
	wire n11586;
	wire n11587;
	wire n11588;
	wire n11589;
	wire n11590;
	wire n11591;
	wire n11592;
	wire n11593;
	wire n11594;
	wire n11595;
	wire n11596;
	wire n11597;
	wire n11598;
	wire n11599;
	wire n11600;
	wire n11601;
	wire n11602;
	wire n11603;
	wire n11604;
	wire n11605;
	wire n11606;
	wire n11607;
	wire n11608;
	wire n11609;
	wire n11610;
	wire n11611;
	wire n11612;
	wire n11613;
	wire n11614;
	wire n11615;
	wire n11616;
	wire n11617;
	wire n11618;
	wire n11619;
	wire n11620;
	wire n11621;
	wire n11622;
	wire n11623;
	wire n11624;
	wire n11625;
	wire n11626;
	wire n11627;
	wire n11628;
	wire n11629;
	wire n11630;
	wire n11631;
	wire n11632;
	wire n11633;
	wire n11634;
	wire n11635;
	wire n11636;
	wire n11637;
	wire n11638;
	wire n11639;
	wire n11640;
	wire n11641;
	wire n11642;
	wire n11643;
	wire n11644;
	wire n11645;
	wire n11646;
	wire n11647;
	wire n11648;
	wire n11649;
	wire n11650;
	wire n11651;
	wire n11652;
	wire n11653;
	wire n11654;
	wire n11656;
	wire n11657;
	wire n11658;
	wire n11659;
	wire n11660;
	wire n11661;
	wire n11662;
	wire n11663;
	wire n11664;
	wire n11665;
	wire n11666;
	wire n11667;
	wire n11668;
	wire n11669;
	wire n11670;
	wire n11671;
	wire n11672;
	wire n11673;
	wire n11674;
	wire n11675;
	wire n11676;
	wire n11677;
	wire n11678;
	wire n11679;
	wire n11680;
	wire n11681;
	wire n11682;
	wire n11683;
	wire n11684;
	wire n11685;
	wire n11686;
	wire n11687;
	wire n11688;
	wire n11689;
	wire n11690;
	wire n11691;
	wire n11692;
	wire n11693;
	wire n11694;
	wire n11695;
	wire n11696;
	wire n11697;
	wire n11698;
	wire n11699;
	wire n11700;
	wire n11701;
	wire n11702;
	wire n11703;
	wire n11704;
	wire n11705;
	wire n11706;
	wire n11707;
	wire n11708;
	wire n11709;
	wire n11710;
	wire n11711;
	wire n11712;
	wire n11713;
	wire n11714;
	wire n11715;
	wire n11716;
	wire n11717;
	wire n11718;
	wire n11719;
	wire n11720;
	wire n11721;
	wire n11722;
	wire n11723;
	wire n11724;
	wire n11725;
	wire n11726;
	wire n11727;
	wire n11728;
	wire n11729;
	wire n11730;
	wire n11731;
	wire n11732;
	wire n11733;
	wire n11734;
	wire n11735;
	wire n11736;
	wire n11737;
	wire n11738;
	wire n11739;
	wire n11740;
	wire n11741;
	wire n11742;
	wire n11743;
	wire n11744;
	wire n11745;
	wire n11746;
	wire n11747;
	wire n11748;
	wire n11749;
	wire n11750;
	wire n11751;
	wire n11752;
	wire n11753;
	wire n11754;
	wire n11755;
	wire n11756;
	wire n11757;
	wire n11758;
	wire n11759;
	wire n11760;
	wire n11761;
	wire n11762;
	wire n11763;
	wire n11764;
	wire n11765;
	wire n11766;
	wire n11767;
	wire n11768;
	wire n11769;
	wire n11770;
	wire n11771;
	wire n11772;
	wire n11773;
	wire n11774;
	wire n11775;
	wire n11776;
	wire n11777;
	wire n11778;
	wire n11779;
	wire n11780;
	wire n11781;
	wire n11782;
	wire n11783;
	wire n11784;
	wire n11785;
	wire n11786;
	wire n11787;
	wire n11788;
	wire n11789;
	wire n11790;
	wire n11791;
	wire n11792;
	wire n11793;
	wire n11794;
	wire n11795;
	wire n11796;
	wire n11797;
	wire n11798;
	wire n11799;
	wire n11800;
	wire n11801;
	wire n11802;
	wire n11803;
	wire n11804;
	wire n11805;
	wire n11806;
	wire n11807;
	wire n11808;
	wire n11809;
	wire n11810;
	wire n11811;
	wire n11812;
	wire n11813;
	wire n11814;
	wire n11815;
	wire n11816;
	wire n11817;
	wire n11818;
	wire n11819;
	wire n11820;
	wire n11821;
	wire n11822;
	wire n11823;
	wire n11824;
	wire n11825;
	wire n11826;
	wire n11827;
	wire n11828;
	wire n11829;
	wire n11830;
	wire n11831;
	wire n11832;
	wire n11833;
	wire n11834;
	wire n11835;
	wire n11836;
	wire n11837;
	wire n11838;
	wire n11839;
	wire n11840;
	wire n11841;
	wire n11842;
	wire n11843;
	wire n11844;
	wire n11845;
	wire n11846;
	wire n11847;
	wire n11851;
	wire n11852;
	wire n11853;
	wire n11854;
	wire n11855;
	wire n11856;
	wire n11858;
	wire n11859;
	wire n11860;
	wire n11861;
	wire n11862;
	wire n11863;
	wire n11864;
	wire n11865;
	wire n11866;
	wire n11867;
	wire n11868;
	wire n11869;
	wire n11870;
	wire n11871;
	wire n11872;
	wire n11873;
	wire n11874;
	wire n11875;
	wire n11876;
	wire n11877;
	wire n11878;
	wire n11879;
	wire n11880;
	wire n11881;
	wire n11882;
	wire n11883;
	wire n11884;
	wire n11885;
	wire n11886;
	wire n11887;
	wire n11888;
	wire n11889;
	wire n11890;
	wire n11891;
	wire n11892;
	wire n11893;
	wire n11894;
	wire n11895;
	wire n11896;
	wire n11897;
	wire n11898;
	wire n11899;
	wire n11900;
	wire n11901;
	wire n11902;
	wire n11903;
	wire n11904;
	wire n11905;
	wire n11906;
	wire n11907;
	wire n11908;
	wire n11909;
	wire n11910;
	wire n11911;
	wire n11912;
	wire n11913;
	wire n11914;
	wire n11915;
	wire n11916;
	wire n11917;
	wire n11918;
	wire n11919;
	wire n11920;
	wire n11921;
	wire n11922;
	wire n11923;
	wire n11924;
	wire n11925;
	wire n11926;
	wire n11927;
	wire n11928;
	wire n11929;
	wire n11930;
	wire n11931;
	wire n11932;
	wire n11933;
	wire n11934;
	wire n11935;
	wire n11936;
	wire n11937;
	wire n11938;
	wire n11939;
	wire n11940;
	wire n11941;
	wire n11942;
	wire n11943;
	wire n11944;
	wire n11945;
	wire n11946;
	wire n11947;
	wire n11948;
	wire n11949;
	wire n11950;
	wire n11951;
	wire n11952;
	wire n11953;
	wire n11954;
	wire n11955;
	wire n11956;
	wire n11957;
	wire n11958;
	wire n11959;
	wire n11960;
	wire n11961;
	wire n11962;
	wire n11963;
	wire n11964;
	wire n11965;
	wire n11966;
	wire n11967;
	wire n11968;
	wire n11969;
	wire n11970;
	wire n11971;
	wire n11972;
	wire n11973;
	wire n11974;
	wire n11975;
	wire n11976;
	wire n11977;
	wire n11978;
	wire n11979;
	wire n11980;
	wire n11981;
	wire n11982;
	wire n11983;
	wire n11984;
	wire n11985;
	wire n11986;
	wire n11987;
	wire n11988;
	wire n11989;
	wire n11990;
	wire n11991;
	wire n11992;
	wire n11993;
	wire n11994;
	wire n11995;
	wire n11996;
	wire n11997;
	wire n11998;
	wire n11999;
	wire n12000;
	wire n12001;
	wire n12002;
	wire n12003;
	wire n12004;
	wire n12005;
	wire n12006;
	wire n12007;
	wire n12008;
	wire n12009;
	wire n12010;
	wire n12011;
	wire n12012;
	wire n12013;
	wire n12014;
	wire n12015;
	wire n12016;
	wire n12017;
	wire n12018;
	wire n12019;
	wire n12020;
	wire n12021;
	wire n12022;
	wire n12023;
	wire n12024;
	wire n12025;
	wire n12026;
	wire n12027;
	wire n12028;
	wire n12029;
	wire n12030;
	wire n12031;
	wire n12032;
	wire n12033;
	wire n12034;
	wire n12035;
	wire n12036;
	wire n12037;
	wire n12038;
	wire n12039;
	wire n12040;
	wire n12041;
	wire n12042;
	wire n12043;
	wire n12044;
	wire n12045;
	wire n12046;
	wire n12047;
	wire n12048;
	wire n12049;
	wire n12050;
	wire n12051;
	wire n12052;
	wire n12053;
	wire n12054;
	wire n12055;
	wire n12056;
	wire n12057;
	wire n12058;
	wire n12059;
	wire n12060;
	wire n12061;
	wire n12062;
	wire n12063;
	wire n12064;
	wire n12065;
	wire n12066;
	wire n12067;
	wire n12068;
	wire n12069;
	wire n12070;
	wire n12071;
	wire n12072;
	wire n12073;
	wire n12074;
	wire n12075;
	wire n12076;
	wire n12077;
	wire n12078;
	wire n12079;
	wire n12080;
	wire n12081;
	wire n12082;
	wire n12083;
	wire n12084;
	wire n12085;
	wire n12086;
	wire n12087;
	wire n12088;
	wire n12089;
	wire n12090;
	wire n12091;
	wire n12092;
	wire n12093;
	wire n12094;
	wire n12095;
	wire n12096;
	wire n12097;
	wire n12098;
	wire n12099;
	wire n12100;
	wire n12101;
	wire n12102;
	wire n12103;
	wire n12104;
	wire n12105;
	wire n12106;
	wire n12107;
	wire n12108;
	wire n12109;
	wire n12110;
	wire n12111;
	wire n12112;
	wire n12113;
	wire n12114;
	wire n12115;
	wire n12116;
	wire n12117;
	wire n12118;
	wire n12119;
	wire n12120;
	wire n12121;
	wire n12122;
	wire n12123;
	wire n12124;
	wire n12125;
	wire n12126;
	wire n12127;
	wire n12128;
	wire n12129;
	wire n12130;
	wire n12131;
	wire n12132;
	wire n12133;
	wire n12134;
	wire n12135;
	wire n12136;
	wire n12137;
	wire n12138;
	wire n12139;
	wire n12140;
	wire n12141;
	wire n12142;
	wire n12143;
	wire n12144;
	wire n12145;
	wire n12146;
	wire n12147;
	wire n12148;
	wire n12149;
	wire n12150;
	wire n12151;
	wire n12152;
	wire n12153;
	wire n12154;
	wire n12155;
	wire n12156;
	wire n12157;
	wire n12158;
	wire n12159;
	wire n12160;
	wire n12161;
	wire n12162;
	wire n12163;
	wire n12164;
	wire n12165;
	wire n12166;
	wire n12167;
	wire n12168;
	wire n12169;
	wire n12170;
	wire n12171;
	wire n12172;
	wire n12173;
	wire n12174;
	wire n12175;
	wire n12176;
	wire n12177;
	wire n12179;
	wire n12180;
	wire n12181;
	wire n12182;
	wire n12183;
	wire n12184;
	wire n12185;
	wire n12186;
	wire n12187;
	wire n12188;
	wire n12189;
	wire n12190;
	wire n12193;
	wire n12194;
	wire n12195;
	wire n12196;
	wire n12197;
	wire n12198;
	wire n12199;
	wire n12200;
	wire n12201;
	wire n12202;
	wire n12203;
	wire n12204;
	wire n12205;
	wire n12206;
	wire n12207;
	wire n12209;
	wire n12210;
	wire n12211;
	wire n12212;
	wire n12213;
	wire n12214;
	wire n12215;
	wire n12216;
	wire n12217;
	wire n12218;
	wire n12219;
	wire n12220;
	wire n12221;
	wire n12222;
	wire n12223;
	wire n12224;
	wire n12225;
	wire n12226;
	wire n12227;
	wire n12228;
	wire n12229;
	wire n12230;
	wire n12231;
	wire n12232;
	wire n12233;
	wire n12234;
	wire n12235;
	wire n12236;
	wire n12237;
	wire n12238;
	wire n12239;
	wire n12240;
	wire n12241;
	wire n12242;
	wire n12243;
	wire n12244;
	wire n12245;
	wire n12246;
	wire n12247;
	wire n12248;
	wire n12249;
	wire n12250;
	wire n12251;
	wire n12252;
	wire n12253;
	wire n12254;
	wire n12255;
	wire n12256;
	wire n12257;
	wire n12258;
	wire n12259;
	wire n12260;
	wire n12261;
	wire n12262;
	wire n12263;
	wire n12264;
	wire n12265;
	wire n12266;
	wire n12267;
	wire n12268;
	wire n12269;
	wire n12270;
	wire n12271;
	wire n12272;
	wire n12273;
	wire n12274;
	wire n12275;
	wire n12276;
	wire n12277;
	wire n12278;
	wire n12279;
	wire n12280;
	wire n12281;
	wire n12282;
	wire n12283;
	wire n12284;
	wire n12285;
	wire n12286;
	wire n12287;
	wire n12288;
	wire n12289;
	wire n12290;
	wire n12291;
	wire n12292;
	wire n12293;
	wire n12294;
	wire n12295;
	wire n12296;
	wire n12297;
	wire n12298;
	wire n12299;
	wire n12300;
	wire n12301;
	wire n12302;
	wire n12303;
	wire n12304;
	wire n12305;
	wire n12306;
	wire n12307;
	wire n12308;
	wire n12309;
	wire n12310;
	wire n12311;
	wire n12312;
	wire n12313;
	wire n12314;
	wire n12315;
	wire n12316;
	wire n12317;
	wire n12318;
	wire n12319;
	wire n12320;
	wire n12321;
	wire n12322;
	wire n12323;
	wire n12324;
	wire n12325;
	wire n12326;
	wire n12327;
	wire n12328;
	wire n12329;
	wire n12330;
	wire n12331;
	wire n12332;
	wire n12333;
	wire n12334;
	wire n12335;
	wire n12336;
	wire n12337;
	wire n12338;
	wire n12339;
	wire n12340;
	wire n12341;
	wire n12342;
	wire n12343;
	wire n12344;
	wire n12345;
	wire n12346;
	wire n12347;
	wire n12348;
	wire n12349;
	wire n12350;
	wire n12351;
	wire n12352;
	wire n12353;
	wire n12354;
	wire n12355;
	wire n12356;
	wire n12357;
	wire n12358;
	wire n12359;
	wire n12360;
	wire n12361;
	wire n12362;
	wire n12363;
	wire n12364;
	wire n12365;
	wire n12366;
	wire n12367;
	wire n12368;
	wire n12369;
	wire n12370;
	wire n12371;
	wire n12372;
	wire n12373;
	wire n12374;
	wire n12375;
	wire n12376;
	wire n12377;
	wire n12378;
	wire n12379;
	wire n12380;
	wire n12381;
	wire n12382;
	wire n12383;
	wire n12384;
	wire n12385;
	wire n12386;
	wire n12387;
	wire n12388;
	wire n12389;
	wire n12390;
	wire n12391;
	wire n12392;
	wire n12393;
	wire n12394;
	wire n12395;
	wire n12396;
	wire n12397;
	wire n12398;
	wire n12399;
	wire n12400;
	wire n12401;
	wire n12402;
	wire n12403;
	wire n12404;
	wire n12405;
	wire n12406;
	wire n12407;
	wire n12408;
	wire n12410;
	wire n12411;
	wire n12412;
	wire n12413;
	wire n12414;
	wire n12415;
	wire n12416;
	wire n12417;
	wire n12418;
	wire n12419;
	wire n12420;
	wire n12421;
	wire n12422;
	wire n12423;
	wire n12424;
	wire n12425;
	wire n12426;
	wire n12427;
	wire n12428;
	wire n12429;
	wire n12430;
	wire n12431;
	wire n12432;
	wire n12433;
	wire n12434;
	wire n12435;
	wire n12436;
	wire n12437;
	wire n12438;
	wire n12439;
	wire n12440;
	wire n12441;
	wire n12442;
	wire n12443;
	wire n12444;
	wire n12445;
	wire n12446;
	wire n12447;
	wire n12448;
	wire n12449;
	wire n12450;
	wire n12451;
	wire n12452;
	wire n12453;
	wire n12454;
	wire n12455;
	wire n12456;
	wire n12457;
	wire n12458;
	wire n12459;
	wire n12460;
	wire n12461;
	wire n12462;
	wire n12463;
	wire n12464;
	wire n12465;
	wire n12466;
	wire n12467;
	wire n12468;
	wire n12469;
	wire n12470;
	wire n12471;
	wire n12472;
	wire n12473;
	wire n12474;
	wire n12475;
	wire n12476;
	wire n12477;
	wire n12478;
	wire n12479;
	wire n12480;
	wire n12481;
	wire n12482;
	wire n12483;
	wire n12484;
	wire n12485;
	wire n12486;
	wire n12487;
	wire n12488;
	wire n12489;
	wire n12490;
	wire n12491;
	wire n12492;
	wire n12493;
	wire n12494;
	wire n12495;
	wire n12496;
	wire n12497;
	wire n12498;
	wire n12499;
	wire n12500;
	wire n12501;
	wire n12502;
	wire n12503;
	wire n12504;
	wire n12505;
	wire n12506;
	wire n12507;
	wire n12508;
	wire n12509;
	wire n12510;
	wire n12511;
	wire n12512;
	wire n12513;
	wire n12514;
	wire n12515;
	wire n12516;
	wire n12517;
	wire n12518;
	wire n12519;
	wire n12520;
	wire n12521;
	wire n12522;
	wire n12523;
	wire n12524;
	wire n12525;
	wire n12526;
	wire n12527;
	wire n12528;
	wire n12529;
	wire n12530;
	wire n12531;
	wire n12532;
	wire n12533;
	wire n12534;
	wire n12535;
	wire n12536;
	wire n12537;
	wire n12538;
	wire n12539;
	wire n12540;
	wire n12541;
	wire n12542;
	wire n12543;
	wire n12544;
	wire n12545;
	wire n12546;
	wire n12547;
	wire n12548;
	wire n12549;
	wire n12550;
	wire n12551;
	wire n12552;
	wire n12553;
	wire n12554;
	wire n12555;
	wire n12556;
	wire n12557;
	wire n12558;
	wire n12559;
	wire n12560;
	wire n12561;
	wire n12562;
	wire n12563;
	wire n12564;
	wire n12565;
	wire n12566;
	wire n12567;
	wire n12568;
	wire n12569;
	wire n12570;
	wire n12571;
	wire n12572;
	wire n12573;
	wire n12574;
	wire n12575;
	wire n12576;
	wire n12577;
	wire n12578;
	wire n12579;
	wire n12580;
	wire n12581;
	wire n12582;
	wire n12583;
	wire n12584;
	wire n12585;
	wire n12586;
	wire n12587;
	wire n12588;
	wire n12589;
	wire n12590;
	wire n12591;
	wire n12592;
	wire n12593;
	wire n12594;
	wire n12595;
	wire n12596;
	wire n12597;
	wire n12598;
	wire n12599;
	wire n12600;
	wire n12601;
	wire n12602;
	wire n12603;
	wire n12604;
	wire n12605;
	wire n12606;
	wire n12607;
	wire n12608;
	wire n12609;
	wire n12610;
	wire n12611;
	wire n12612;
	wire n12613;
	wire n12614;
	wire n12615;
	wire n12616;
	wire n12617;
	wire n12618;
	wire n12619;
	wire n12620;
	wire n12621;
	wire n12622;
	wire n12623;
	wire n12624;
	wire n12625;
	wire n12626;
	wire n12627;
	wire n12628;
	wire n12629;
	wire n12630;
	wire n12631;
	wire n12632;
	wire n12633;
	wire n12634;
	wire n12635;
	wire n12636;
	wire n12637;
	wire n12638;
	wire n12639;
	wire n12640;
	wire n12641;
	wire n12642;
	wire n12643;
	wire n12644;
	wire n12645;
	wire n12646;
	wire n12647;
	wire n12648;
	wire n12649;
	wire n12650;
	wire n12651;
	wire n12652;
	wire n12653;
	wire n12654;
	wire n12655;
	wire n12656;
	wire n12657;
	wire n12658;
	wire n12659;
	wire n12660;
	wire n12661;
	wire n12662;
	wire n12663;
	wire n12664;
	wire n12665;
	wire n12666;
	wire n12667;
	wire n12668;
	wire n12669;
	wire n12670;
	wire n12671;
	wire n12672;
	wire n12673;
	wire n12674;
	wire n12675;
	wire n12676;
	wire n12677;
	wire n12678;
	wire n12679;
	wire n12680;
	wire n12681;
	wire n12682;
	wire n12683;
	wire n12684;
	wire n12685;
	wire n12686;
	wire n12687;
	wire n12688;
	wire n12689;
	wire n12690;
	wire n12691;
	wire n12692;
	wire n12693;
	wire n12694;
	wire n12695;
	wire n12696;
	wire n12697;
	wire n12698;
	wire n12699;
	wire n12700;
	wire n12701;
	wire n12702;
	wire n12703;
	wire n12704;
	wire n12705;
	wire n12706;
	wire n12707;
	wire n12708;
	wire n12709;
	wire n12710;
	wire n12711;
	wire n12712;
	wire n12713;
	wire n12714;
	wire n12715;
	wire n12716;
	wire n12717;
	wire n12718;
	wire n12719;
	wire n12720;
	wire n12721;
	wire n12722;
	wire n12723;
	wire n12724;
	wire n12725;
	wire n12726;
	wire n12727;
	wire n12728;
	wire n12729;
	wire n12730;
	wire n12731;
	wire n12732;
	wire n12733;
	wire n12734;
	wire n12735;
	wire n12736;
	wire n12737;
	wire n12738;
	wire n12739;
	wire n12740;
	wire n12741;
	wire n12742;
	wire n12743;
	wire n12744;
	wire n12745;
	wire n12746;
	wire n12747;
	wire n12748;
	wire n12749;
	wire n12750;
	wire n12751;
	wire n12752;
	wire n12753;
	wire n12754;
	wire n12755;
	wire n12756;
	wire n12757;
	wire n12758;
	wire n12759;
	wire n12760;
	wire n12761;
	wire n12762;
	wire n12763;
	wire n12764;
	wire n12765;
	wire n12766;
	wire n12767;
	wire n12768;
	wire n12769;
	wire n12770;
	wire n12771;
	wire n12772;
	wire n12773;
	wire n12774;
	wire n12775;
	wire n12776;
	wire n12777;
	wire n12778;
	wire n12779;
	wire n12780;
	wire n12781;
	wire n12782;
	wire n12783;
	wire n12784;
	wire n12785;
	wire n12786;
	wire n12787;
	wire n12788;
	wire n12789;
	wire n12790;
	wire n12791;
	wire n12792;
	wire n12793;
	wire n12794;
	wire n12795;
	wire n12796;
	wire n12797;
	wire n12798;
	wire n12799;
	wire n12800;
	wire n12801;
	wire n12802;
	wire n12803;
	wire n12804;
	wire n12805;
	wire n12806;
	wire n12807;
	wire n12808;
	wire n12809;
	wire n12810;
	wire n12811;
	wire n12812;
	wire n12813;
	wire n12814;
	wire n12815;
	wire n12816;
	wire n12817;
	wire n12818;
	wire n12819;
	wire n12820;
	wire n12821;
	wire n12822;
	wire n12823;
	wire n12824;
	wire n12825;
	wire n12826;
	wire n12827;
	wire n12828;
	wire n12829;
	wire n12830;
	wire n12831;
	wire n12832;
	wire n12833;
	wire n12834;
	wire n12835;
	wire n12836;
	wire n12837;
	wire n12838;
	wire n12839;
	wire n12840;
	wire n12841;
	wire n12842;
	wire n12843;
	wire n12844;
	wire n12845;
	wire n12846;
	wire n12847;
	wire n12848;
	wire n12849;
	wire n12850;
	wire n12851;
	wire n12852;
	wire n12853;
	wire n12854;
	wire n12855;
	wire n12856;
	wire n12857;
	wire n12858;
	wire n12859;
	wire n12860;
	wire n12861;
	wire n12862;
	wire n12863;
	wire n12864;
	wire n12865;
	wire n12866;
	wire n12867;
	wire n12868;
	wire n12869;
	wire n12870;
	wire n12871;
	wire n12872;
	wire n12873;
	wire n12874;
	wire n12875;
	wire n12876;
	wire n12877;
	wire n12878;
	wire n12879;
	wire n12880;
	wire n12881;
	wire n12882;
	wire n12883;
	wire n12884;
	wire n12885;
	wire n12886;
	wire n12887;
	wire n12888;
	wire n12889;
	wire n12890;
	wire n12891;
	wire n12892;
	wire n12893;
	wire n12894;
	wire n12895;
	wire n12896;
	wire n12897;
	wire n12898;
	wire n12899;
	wire n12900;
	wire n12901;
	wire n12902;
	wire n12903;
	wire n12904;
	wire n12905;
	wire n12906;
	wire n12907;
	wire n12908;
	wire n12909;
	wire n12910;
	wire n12911;
	wire n12912;
	wire n12913;
	wire n12914;
	wire n12915;
	wire n12916;
	wire n12917;
	wire n12918;
	wire n12919;
	wire n12920;
	wire n12921;
	wire n12922;
	wire n12923;
	wire n12924;
	wire n12925;
	wire n12926;
	wire n12927;
	wire n12928;
	wire n12929;
	wire n12930;
	wire n12931;
	wire n12932;
	wire n12933;
	wire n12934;
	wire n12935;
	wire n12937;
	wire n12938;
	wire n12939;
	wire n12940;
	wire n12941;
	wire n12942;
	wire n12943;
	wire n12944;
	wire n12945;
	wire n12946;
	wire n12947;
	wire n12948;
	wire n12949;
	wire n12950;
	wire n12951;
	wire n12952;
	wire n12953;
	wire n12954;
	wire n12955;
	wire n12956;
	wire n12957;
	wire n12958;
	wire n12959;
	wire n12960;
	wire n12961;
	wire n12962;
	wire n12963;
	wire n12964;
	wire n12965;
	wire n12966;
	wire n12967;
	wire n12968;
	wire n12969;
	wire n12970;
	wire n12971;
	wire n12972;
	wire n12973;
	wire n12974;
	wire n12975;
	wire n12976;
	wire n12977;
	wire n12978;
	wire n12979;
	wire n12980;
	wire n12981;
	wire n12982;
	wire n12983;
	wire n12984;
	wire n12985;
	wire n12986;
	wire n12987;
	wire n12988;
	wire n12989;
	wire n12990;
	wire n12991;
	wire n12992;
	wire n12993;
	wire n12994;
	wire n12995;
	wire n12996;
	wire n12997;
	wire n12998;
	wire n12999;
	wire n13000;
	wire n13001;
	wire n13002;
	wire n13003;
	wire n13004;
	wire n13005;
	wire n13006;
	wire n13007;
	wire n13008;
	wire n13009;
	wire n13010;
	wire n13011;
	wire n13012;
	wire n13013;
	wire n13014;
	wire n13015;
	wire n13016;
	wire n13017;
	wire n13018;
	wire n13019;
	wire n13020;
	wire n13021;
	wire n13022;
	wire n13023;
	wire n13024;
	wire n13025;
	wire n13026;
	wire n13027;
	wire n13028;
	wire n13029;
	wire n13030;
	wire n13031;
	wire n13032;
	wire n13033;
	wire n13034;
	wire n13035;
	wire n13036;
	wire n13037;
	wire n13038;
	wire n13039;
	wire n13040;
	wire n13041;
	wire n13042;
	wire n13043;
	wire n13044;
	wire n13045;
	wire n13046;
	wire n13047;
	wire n13048;
	wire n13049;
	wire n13050;
	wire n13051;
	wire n13052;
	wire n13053;
	wire n13054;
	wire n13055;
	wire n13056;
	wire n13057;
	wire n13058;
	wire n13059;
	wire n13060;
	wire n13061;
	wire n13062;
	wire n13063;
	wire n13064;
	wire n13065;
	wire n13066;
	wire n13067;
	wire n13068;
	wire n13069;
	wire n13070;
	wire n13071;
	wire n13072;
	wire n13073;
	wire n13074;
	wire n13075;
	wire n13076;
	wire n13077;
	wire n13078;
	wire n13079;
	wire n13080;
	wire n13081;
	wire n13082;
	wire n13083;
	wire n13084;
	wire n13085;
	wire n13086;
	wire n13087;
	wire n13088;
	wire n13089;
	wire n13090;
	wire n13091;
	wire n13092;
	wire n13093;
	wire n13094;
	wire n13095;
	wire n13096;
	wire n13097;
	wire n13098;
	wire n13099;
	wire n13100;
	wire n13101;
	wire n13102;
	wire n13103;
	wire n13104;
	wire n13105;
	wire n13106;
	wire n13107;
	wire n13108;
	wire n13109;
	wire n13110;
	wire n13111;
	wire n13112;
	wire n13113;
	wire n13114;
	wire n13115;
	wire n13116;
	wire n13117;
	wire n13118;
	wire n13119;
	wire n13120;
	wire n13121;
	wire n13122;
	wire n13123;
	wire n13124;
	wire n13125;
	wire n13126;
	wire n13127;
	wire n13128;
	wire n13129;
	wire n13130;
	wire n13131;
	wire n13132;
	wire n13133;
	wire n13134;
	wire n13135;
	wire n13136;
	wire n13137;
	wire n13138;
	wire n13139;
	wire n13140;
	wire n13141;
	wire n13142;
	wire n13143;
	wire n13144;
	wire n13145;
	wire n13146;
	wire n13147;
	wire n13148;
	wire n13149;
	wire n13150;
	wire n13151;
	wire n13152;
	wire n13153;
	wire n13154;
	wire n13155;
	wire n13156;
	wire n13157;
	wire n13158;
	wire n13159;
	wire n13160;
	wire n13161;
	wire n13162;
	wire n13163;
	wire n13164;
	wire n13165;
	wire n13166;
	wire n13167;
	wire n13168;
	wire n13169;
	wire n13170;
	wire n13171;
	wire n13172;
	wire n13173;
	wire n13174;
	wire n13175;
	wire n13176;
	wire n13177;
	wire n13178;
	wire n13179;
	wire n13180;
	wire n13181;
	wire n13182;
	wire n13183;
	wire n13184;
	wire n13185;
	wire n13186;
	wire n13187;
	wire n13188;
	wire n13189;
	wire n13190;
	wire n13191;
	wire n13192;
	wire n13193;
	wire n13194;
	wire n13195;
	wire n13196;
	wire n13197;
	wire n13198;
	wire n13199;
	wire n13200;
	wire n13201;
	wire n13202;
	wire n13203;
	wire n13204;
	wire n13205;
	wire n13206;
	wire n13207;
	wire n13208;
	wire n13209;
	wire n13210;
	wire n13211;
	wire n13212;
	wire n13213;
	wire n13214;
	wire n13215;
	wire n13216;
	wire n13217;
	wire n13218;
	wire n13219;
	wire n13220;
	wire n13221;
	wire n13222;
	wire n13223;
	wire n13224;
	wire n13225;
	wire n13226;
	wire n13227;
	wire n13228;
	wire n13229;
	wire n13230;
	wire n13231;
	wire n13232;
	wire n13233;
	wire n13234;
	wire n13235;
	wire n13236;
	wire n13237;
	wire n13238;
	wire n13239;
	wire n13240;
	wire n13241;
	wire n13242;
	wire n13243;
	wire n13244;
	wire n13245;
	wire n13246;
	wire n13247;
	wire n13248;
	wire n13249;
	wire n13250;
	wire n13251;
	wire n13252;
	wire n13253;
	wire n13254;
	wire n13255;
	wire n13256;
	wire n13257;
	wire n13258;
	wire n13259;
	wire n13260;
	wire n13261;
	wire n13262;
	wire n13263;
	wire n13264;
	wire n13265;
	wire n13266;
	wire n13267;
	wire n13268;
	wire n13269;
	wire n13270;
	wire n13271;
	wire n13272;
	wire n13273;
	wire n13274;
	wire n13275;
	wire n13276;
	wire n13277;
	wire n13278;
	wire n13279;
	wire n13280;
	wire n13281;
	wire n13282;
	wire n13283;
	wire n13284;
	wire n13285;
	wire n13286;
	wire n13287;
	wire n13288;
	wire n13289;
	wire n13290;
	wire n13291;
	wire n13292;
	wire n13293;
	wire n13294;
	wire n13296;
	wire n13297;
	wire n13298;
	wire n13299;
	wire n13300;
	wire n13301;
	wire n13302;
	wire n13303;
	wire n13304;
	wire n13305;
	wire n13306;
	wire n13307;
	wire n13308;
	wire n13309;
	wire n13310;
	wire n13311;
	wire n13312;
	wire n13313;
	wire n13314;
	wire n13315;
	wire n13316;
	wire n13317;
	wire n13318;
	wire n13319;
	wire n13320;
	wire n13321;
	wire n13322;
	wire n13323;
	wire n13324;
	wire n13325;
	wire n13326;
	wire n13327;
	wire n13328;
	wire n13329;
	wire n13330;
	wire n13331;
	wire n13332;
	wire n13333;
	wire n13334;
	wire n13335;
	wire n13336;
	wire n13337;
	wire n13338;
	wire n13339;
	wire n13340;
	wire n13341;
	wire n13342;
	wire n13343;
	wire n13344;
	wire n13345;
	wire n13346;
	wire n13347;
	wire n13348;
	wire n13349;
	wire n13350;
	wire n13351;
	wire n13352;
	wire n13353;
	wire n13354;
	wire n13355;
	wire n13356;
	wire n13357;
	wire n13358;
	wire n13359;
	wire n13360;
	wire n13361;
	wire n13362;
	wire n13363;
	wire n13364;
	wire n13365;
	wire n13366;
	wire n13367;
	wire n13368;
	wire n13369;
	wire n13370;
	wire n13371;
	wire n13372;
	wire n13373;
	wire n13374;
	wire n13375;
	wire n13376;
	wire n13377;
	wire n13378;
	wire n13379;
	wire n13380;
	wire n13381;
	wire n13382;
	wire n13383;
	wire n13384;
	wire n13385;
	wire n13386;
	wire n13387;
	wire n13388;
	wire n13389;
	wire n13390;
	wire n13391;
	wire n13392;
	wire n13393;
	wire n13394;
	wire n13395;
	wire n13396;
	wire n13397;
	wire n13398;
	wire n13399;
	wire n13400;
	wire n13401;
	wire n13402;
	wire n13403;
	wire n13404;
	wire n13405;
	wire n13406;
	wire n13407;
	wire n13408;
	wire n13409;
	wire n13410;
	wire n13411;
	wire n13412;
	wire n13413;
	wire n13414;
	wire n13415;
	wire n13416;
	wire n13417;
	wire n13418;
	wire n13419;
	wire n13420;
	wire n13421;
	wire n13422;
	wire n13423;
	wire n13424;
	wire n13425;
	wire n13426;
	wire n13427;
	wire n13428;
	wire n13429;
	wire n13430;
	wire n13431;
	wire n13432;
	wire n13433;
	wire n13434;
	wire n13435;
	wire n13436;
	wire n13437;
	wire n13438;
	wire n13439;
	wire n13440;
	wire n13441;
	wire n13442;
	wire n13443;
	wire n13444;
	wire n13445;
	wire n13446;
	wire n13447;
	wire n13448;
	wire n13449;
	wire n13450;
	wire n13451;
	wire n13452;
	wire n13453;
	wire n13454;
	wire n13455;
	wire n13456;
	wire n13457;
	wire n13458;
	wire n13459;
	wire n13460;
	wire n13461;
	wire n13462;
	wire n13463;
	wire n13464;
	wire n13465;
	wire n13466;
	wire n13467;
	wire n13468;
	wire n13469;
	wire n13470;
	wire n13471;
	wire n13472;
	wire n13473;
	wire n13474;
	wire n13475;
	wire n13476;
	wire n13477;
	wire n13478;
	wire n13479;
	wire n13480;
	wire n13481;
	wire n13482;
	wire n13483;
	wire n13484;
	wire n13485;
	wire n13486;
	wire n13487;
	wire n13488;
	wire n13489;
	wire n13490;
	wire n13491;
	wire n13492;
	wire n13493;
	wire n13494;
	wire n13495;
	wire n13496;
	wire n13497;
	wire n13498;
	wire n13499;
	wire n13500;
	wire n13501;
	wire n13502;
	wire n13503;
	wire n13504;
	wire n13505;
	wire n13506;
	wire n13507;
	wire n13508;
	wire n13509;
	wire n13510;
	wire n13511;
	wire n13512;
	wire n13513;
	wire n13514;
	wire n13515;
	wire n13516;
	wire n13517;
	wire n13518;
	wire n13519;
	wire n13520;
	wire n13521;
	wire n13522;
	wire n13523;
	wire n13524;
	wire n13525;
	wire n13526;
	wire n13527;
	wire n13528;
	wire n13529;
	wire n13530;
	wire n13531;
	wire n13532;
	wire n13533;
	wire n13534;
	wire n13535;
	wire n13536;
	wire n13537;
	wire n13538;
	wire n13539;
	wire n13540;
	wire n13541;
	wire n13542;
	wire n13543;
	wire n13544;
	wire n13545;
	wire n13546;
	wire n13547;
	wire n13548;
	wire n13549;
	wire n13550;
	wire n13551;
	wire n13552;
	wire n13553;
	wire n13554;
	wire n13555;
	wire n13556;
	wire n13557;
	wire n13558;
	wire n13559;
	wire n13560;
	wire n13561;
	wire n13562;
	wire n13563;
	wire n13564;
	wire n13565;
	wire n13566;
	wire n13567;
	wire n13568;
	wire n13569;
	wire n13570;
	wire n13571;
	wire n13572;
	wire n13573;
	wire n13574;
	wire n13575;
	wire n13576;
	wire n13577;
	wire n13578;
	wire n13579;
	wire n13580;
	wire n13581;
	wire n13582;
	wire n13583;
	wire n13584;
	wire n13585;
	wire n13586;
	wire n13587;
	wire n13588;
	wire n13589;
	wire n13590;
	wire n13591;
	wire n13592;
	wire n13593;
	wire n13594;
	wire n13595;
	wire n13596;
	wire n13597;
	wire n13598;
	wire n13599;
	wire n13600;
	wire n13601;
	wire n13602;
	wire n13603;
	wire n13604;
	wire n13605;
	wire n13606;
	wire n13607;
	wire n13608;
	wire n13609;
	wire n13610;
	wire n13611;
	wire n13612;
	wire n13613;
	wire n13614;
	wire n13615;
	wire n13616;
	wire n13617;
	wire n13618;
	wire n13619;
	wire n13620;
	wire n13621;
	wire n13622;
	wire n13623;
	wire n13624;
	wire n13625;
	wire n13626;
	wire n13627;
	wire n13628;
	wire n13629;
	wire n13630;
	wire n13631;
	wire n13632;
	wire n13633;
	wire n13634;
	wire n13635;
	wire n13636;
	wire n13637;
	wire n13638;
	wire n13639;
	wire n13640;
	wire n13641;
	wire n13642;
	wire n13643;
	wire n13644;
	wire n13645;
	wire n13646;
	wire n13647;
	wire n13648;
	wire n13649;
	wire n13650;
	wire n13651;
	wire n13652;
	wire n13653;
	wire n13654;
	wire n13655;
	wire n13656;
	wire n13657;
	wire n13658;
	wire n13659;
	wire n13660;
	wire n13661;
	wire n13662;
	wire n13663;
	wire n13664;
	wire n13665;
	wire n13666;
	wire n13667;
	wire n13668;
	wire n13669;
	wire n13670;
	wire n13671;
	wire n13672;
	wire n13673;
	wire n13674;
	wire n13675;
	wire n13676;
	wire n13677;
	wire n13678;
	wire n13679;
	wire n13680;
	wire n13681;
	wire n13682;
	wire n13683;
	wire n13684;
	wire n13685;
	wire n13686;
	wire n13687;
	wire n13688;
	wire n13689;
	wire n13690;
	wire n13691;
	wire n13692;
	wire n13693;
	wire n13694;
	wire n13695;
	wire n13696;
	wire n13697;
	wire n13698;
	wire n13699;
	wire n13700;
	wire n13701;
	wire n13702;
	wire n13703;
	wire n13704;
	wire n13705;
	wire n13706;
	wire n13707;
	wire n13708;
	wire n13709;
	wire n13710;
	wire n13711;
	wire n13712;
	wire n13713;
	wire n13714;
	wire n13715;
	wire n13716;
	wire n13717;
	wire n13718;
	wire n13719;
	wire n13720;
	wire n13721;
	wire n13722;
	wire n13723;
	wire n13724;
	wire n13725;
	wire n13726;
	wire n13727;
	wire n13728;
	wire n13729;
	wire n13730;
	wire n13731;
	wire n13732;
	wire n13733;
	wire n13734;
	wire n13735;
	wire n13736;
	wire n13737;
	wire n13738;
	wire n13739;
	wire n13740;
	wire n13741;
	wire n13742;
	wire n13743;
	wire n13744;
	wire n13745;
	wire n13746;
	wire n13747;
	wire n13748;
	wire n13749;
	wire n13750;
	wire n13751;
	wire n13752;
	wire n13753;
	wire n13754;
	wire n13755;
	wire n13756;
	wire n13757;
	wire n13758;
	wire n13759;
	wire n13760;
	wire n13761;
	wire n13762;
	wire n13763;
	wire n13764;
	wire n13765;
	wire n13766;
	wire n13767;
	wire n13768;
	wire n13769;
	wire n13770;
	wire n13771;
	wire n13772;
	wire n13773;
	wire n13774;
	wire n13775;
	wire n13776;
	wire n13777;
	wire n13778;
	wire n13779;
	wire n13780;
	wire n13781;
	wire n13782;
	wire n13783;
	wire n13784;
	wire n13785;
	wire n13786;
	wire n13787;
	wire n13788;
	wire n13789;
	wire n13790;
	wire n13791;
	wire n13792;
	wire n13793;
	wire n13794;
	wire n13795;
	wire n13796;
	wire n13797;
	wire n13798;
	wire n13799;
	wire n13800;
	wire n13801;
	wire n13802;
	wire n13803;
	wire n13804;
	wire n13805;
	wire n13806;
	wire n13807;
	wire n13808;
	wire n13809;
	wire n13810;
	wire n13811;
	wire n13812;
	wire n13813;
	wire n13814;
	wire n13815;
	wire n13816;
	wire n13817;
	wire n13818;
	wire n13819;
	wire n13820;
	wire n13821;
	wire n13822;
	wire n13823;
	wire n13824;
	wire n13825;
	wire n13826;
	wire n13827;
	wire n13828;
	wire n13829;
	wire n13830;
	wire n13831;
	wire n13832;
	wire n13833;
	wire n13834;
	wire n13835;
	wire n13836;
	wire n13837;
	wire n13838;
	wire n13839;
	wire n13840;
	wire n13841;
	wire n13842;
	wire n13843;
	wire n13844;
	wire n13845;
	wire n13846;
	wire n13847;
	wire n13848;
	wire n13849;
	wire n13850;
	wire n13851;
	wire n13852;
	wire n13853;
	wire n13854;
	wire n13855;
	wire n13856;
	wire n13857;
	wire n13858;
	wire n13859;
	wire n13860;
	wire n13861;
	wire n13862;
	wire n13863;
	wire n13864;
	wire n13865;
	wire n13866;
	wire n13867;
	wire n13868;
	wire n13869;
	wire n13870;
	wire n13871;
	wire n13872;
	wire n13873;
	wire n13874;
	wire n13875;
	wire n13876;
	wire n13877;
	wire n13878;
	wire n13879;
	wire n13880;
	wire n13881;
	wire n13882;
	wire n13883;
	wire n13884;
	wire n13885;
	wire n13886;
	wire n13887;
	wire n13888;
	wire n13889;
	wire n13890;
	wire n13891;
	wire n13892;
	wire n13893;
	wire n13894;
	wire n13895;
	wire n13896;
	wire n13897;
	wire n13898;
	wire n13899;
	wire n13900;
	wire n13901;
	wire n13902;
	wire n13903;
	wire n13904;
	wire n13905;
	wire n13906;
	wire n13907;
	wire n13908;
	wire n13909;
	wire n13910;
	wire n13911;
	wire n13912;
	wire n13913;
	wire n13914;
	wire n13915;
	wire n13916;
	wire n13917;
	wire n13918;
	wire n13919;
	wire n13920;
	wire n13921;
	wire n13922;
	wire n13923;
	wire n13924;
	wire n13925;
	wire n13926;
	wire n13927;
	wire n13928;
	wire n13929;
	wire n13930;
	wire n13931;
	wire n13932;
	wire n13933;
	wire n13934;
	wire n13935;
	wire n13936;
	wire n13937;
	wire n13938;
	wire n13939;
	wire n13940;
	wire n13941;
	wire n13942;
	wire n13943;
	wire n13944;
	wire n13945;
	wire n13946;
	wire n13947;
	wire n13948;
	wire n13949;
	wire n13950;
	wire n13951;
	wire n13952;
	wire n13953;
	wire n13954;
	wire n13955;
	wire n13956;
	wire n13957;
	wire n13958;
	wire n13959;
	wire n13960;
	wire n13961;
	wire n13962;
	wire n13963;
	wire n13964;
	wire n13965;
	wire n13966;
	wire n13967;
	wire n13968;
	wire n13969;
	wire n13970;
	wire n13971;
	wire n13972;
	wire n13973;
	wire n13974;
	wire n13975;
	wire n13976;
	wire n13977;
	wire n13978;
	wire n13979;
	wire n13980;
	wire n13981;
	wire n13982;
	wire n13983;
	wire n13984;
	wire n13985;
	wire n13986;
	wire n13987;
	wire n13988;
	wire n13989;
	wire n13990;
	wire n13991;
	wire n13992;
	wire n13993;
	wire n13994;
	wire n13995;
	wire n13996;
	wire n13997;
	wire n13998;
	wire n13999;
	wire n14000;
	wire n14001;
	wire n14002;
	wire n14003;
	wire n14004;
	wire n14005;
	wire n14006;
	wire n14007;
	wire n14008;
	wire n14009;
	wire n14010;
	wire n14011;
	wire n14012;
	wire n14013;
	wire n14014;
	wire n14015;
	wire n14016;
	wire n14017;
	wire n14018;
	wire n14019;
	wire n14020;
	wire n14021;
	wire n14022;
	wire n14023;
	wire n14024;
	wire n14025;
	wire n14026;
	wire n14027;
	wire n14028;
	wire n14029;
	wire n14030;
	wire n14031;
	wire n14032;
	wire n14033;
	wire n14034;
	wire n14035;
	wire n14036;
	wire n14037;
	wire n14038;
	wire n14039;
	wire n14040;
	wire n14041;
	wire n14042;
	wire n14043;
	wire n14044;
	wire n14045;
	wire n14046;
	wire n14047;
	wire n14048;
	wire n14049;
	wire n14050;
	wire n14051;
	wire n14052;
	wire n14053;
	wire n14054;
	wire n14055;
	wire n14056;
	wire n14057;
	wire n14058;
	wire n14059;
	wire n14060;
	wire n14061;
	wire n14062;
	wire n14063;
	wire n14064;
	wire n14065;
	wire n14066;
	wire n14067;
	wire n14068;
	wire n14070;
	wire n14071;
	wire n14072;
	wire n14073;
	wire n14074;
	wire n14075;
	wire n14076;
	wire n14077;
	wire n14078;
	wire n14079;
	wire n14080;
	wire n14081;
	wire n14082;
	wire n14083;
	wire n14084;
	wire n14085;
	wire n14086;
	wire n14087;
	wire n14088;
	wire n14089;
	wire n14090;
	wire n14091;
	wire n14092;
	wire n14093;
	wire n14094;
	wire n14095;
	wire n14096;
	wire n14097;
	wire n14098;
	wire n14099;
	wire n14100;
	wire n14101;
	wire n14102;
	wire n14103;
	wire n14104;
	wire n14105;
	wire n14106;
	wire n14107;
	wire n14108;
	wire n14109;
	wire n14110;
	wire n14111;
	wire n14112;
	wire n14113;
	wire n14114;
	wire n14115;
	wire n14116;
	wire n14117;
	wire n14118;
	wire n14119;
	wire n14120;
	wire n14121;
	wire n14122;
	wire n14123;
	wire n14124;
	wire n14125;
	wire n14126;
	wire n14127;
	wire n14128;
	wire n14129;
	wire n14130;
	wire n14131;
	wire n14132;
	wire n14133;
	wire n14134;
	wire n14135;
	wire n14136;
	wire n14137;
	wire n14138;
	wire n14139;
	wire n14140;
	wire n14141;
	wire n14142;
	wire n14143;
	wire n14144;
	wire n14145;
	wire n14146;
	wire n14147;
	wire n14148;
	wire n14149;
	wire n14150;
	wire n14151;
	wire n14152;
	wire n14153;
	wire n14154;
	wire n14155;
	wire n14156;
	wire n14157;
	wire n14158;
	wire n14159;
	wire n14160;
	wire n14161;
	wire n14162;
	wire n14163;
	wire n14164;
	wire n14165;
	wire n14166;
	wire n14167;
	wire n14168;
	wire n14169;
	wire n14170;
	wire n14171;
	wire n14172;
	wire n14173;
	wire n14174;
	wire n14175;
	wire n14176;
	wire n14177;
	wire n14178;
	wire n14179;
	wire n14180;
	wire n14181;
	wire n14182;
	wire n14183;
	wire n14184;
	wire n14185;
	wire n14186;
	wire n14187;
	wire n14188;
	wire n14189;
	wire n14190;
	wire n14191;
	wire n14192;
	wire n14193;
	wire n14194;
	wire n14195;
	wire n14196;
	wire n14197;
	wire n14198;
	wire n14199;
	wire n14200;
	wire n14201;
	wire n14202;
	wire n14203;
	wire n14204;
	wire n14205;
	wire n14206;
	wire n14207;
	wire n14208;
	wire n14209;
	wire n14210;
	wire n14211;
	wire n14212;
	wire n14213;
	wire n14214;
	wire n14215;
	wire n14216;
	wire n14217;
	wire n14218;
	wire n14219;
	wire n14220;
	wire n14221;
	wire n14222;
	wire n14223;
	wire n14224;
	wire n14225;
	wire n14226;
	wire n14227;
	wire n14228;
	wire n14229;
	wire n14230;
	wire n14231;
	wire n14232;
	wire n14233;
	wire n14234;
	wire n14235;
	wire n14236;
	wire n14237;
	wire n14238;
	wire n14239;
	wire n14240;
	wire n14241;
	wire n14242;
	wire n14243;
	wire n14244;
	wire n14245;
	wire n14246;
	wire n14247;
	wire n14248;
	wire n14249;
	wire n14250;
	wire n14251;
	wire n14252;
	wire n14253;
	wire n14254;
	wire n14255;
	wire n14256;
	wire n14257;
	wire n14258;
	wire n14259;
	wire n14260;
	wire n14261;
	wire n14262;
	wire n14263;
	wire n14264;
	wire n14265;
	wire n14266;
	wire n14267;
	wire n14268;
	wire n14269;
	wire n14270;
	wire n14271;
	wire n14272;
	wire n14273;
	wire n14274;
	wire n14275;
	wire n14276;
	wire n14277;
	wire n14278;
	wire n14279;
	wire n14280;
	wire n14281;
	wire n14282;
	wire n14283;
	wire n14284;
	wire n14285;
	wire n14286;
	wire n14287;
	wire n14288;
	wire n14289;
	wire n14290;
	wire n14291;
	wire n14292;
	wire n14293;
	wire n14294;
	wire n14295;
	wire n14296;
	wire n14297;
	wire n14298;
	wire n14299;
	wire n14300;
	wire n14301;
	wire n14302;
	wire n14303;
	wire n14304;
	wire n14305;
	wire n14306;
	wire n14307;
	wire n14308;
	wire n14309;
	wire n14310;
	wire n14311;
	wire n14312;
	wire n14313;
	wire n14314;
	wire n14315;
	wire n14316;
	wire n14317;
	wire n14318;
	wire n14319;
	wire n14320;
	wire n14321;
	wire n14322;
	wire n14323;
	wire n14324;
	wire n14325;
	wire n14326;
	wire n14327;
	wire n14328;
	wire n14329;
	wire n14330;
	wire n14331;
	wire n14332;
	wire n14333;
	wire n14334;
	wire n14335;
	wire n14336;
	wire n14337;
	wire n14338;
	wire n14339;
	wire n14340;
	wire n14341;
	wire n14342;
	wire n14343;
	wire n14344;
	wire n14345;
	wire n14346;
	wire n14347;
	wire n14348;
	wire n14349;
	wire n14350;
	wire n14351;
	wire n14352;
	wire n14353;
	wire n14354;
	wire n14355;
	wire n14356;
	wire n14357;
	wire n14358;
	wire n14359;
	wire n14360;
	wire n14361;
	wire n14362;
	wire n14363;
	wire n14364;
	wire n14365;
	wire n14366;
	wire n14367;
	wire n14368;
	wire n14369;
	wire n14370;
	wire n14371;
	wire n14372;
	wire n14373;
	wire n14374;
	wire n14375;
	wire n14376;
	wire n14377;
	wire n14378;
	wire n14379;
	wire n14380;
	wire n14381;
	wire n14382;
	wire n14383;
	wire n14384;
	wire n14385;
	wire n14386;
	wire n14387;
	wire n14388;
	wire n14389;
	wire n14390;
	wire n14391;
	wire n14392;
	wire n14393;
	wire n14394;
	wire n14395;
	wire n14396;
	wire n14397;
	wire n14398;
	wire n14399;
	wire n14400;
	wire n14401;
	wire n14402;
	wire n14403;
	wire n14404;
	wire n14405;
	wire n14406;
	wire n14407;
	wire n14408;
	wire n14409;
	wire n14410;
	wire n14411;
	wire n14412;
	wire n14413;
	wire n14414;
	wire n14415;
	wire n14416;
	wire n14417;
	wire n14418;
	wire n14419;
	wire n14420;
	wire n14421;
	wire n14422;
	wire n14423;
	wire n14424;
	wire n14425;
	wire n14426;
	wire n14427;
	wire n14429;
	wire n14430;
	wire n14431;
	wire n14432;
	wire n14433;
	wire n14434;
	wire n14435;
	wire n14436;
	wire n14437;
	wire n14438;
	wire n14439;
	wire n14440;
	wire n14443;
	wire n14444;
	wire n14445;
	wire n14446;
	wire n14447;
	wire n14448;
	wire n14449;
	wire n14450;
	wire n14451;
	wire n14452;
	wire n14453;
	wire n14454;
	wire n14456;
	wire n14457;
	wire n14458;
	wire n14459;
	wire n14460;
	wire n14461;
	wire n14462;
	wire n14463;
	wire n14464;
	wire n14465;
	wire n14466;
	wire n14467;
	wire n14468;
	wire n14469;
	wire n14470;
	wire n14471;
	wire n14472;
	wire n14473;
	wire n14474;
	wire n14475;
	wire n14476;
	wire n14477;
	wire n14478;
	wire n14479;
	wire n14480;
	wire n14481;
	wire n14482;
	wire n14483;
	wire n14484;
	wire n14485;
	wire n14486;
	wire n14487;
	wire n14488;
	wire n14489;
	wire n14490;
	wire n14491;
	wire n14492;
	wire n14493;
	wire n14494;
	wire n14495;
	wire n14496;
	wire n14497;
	wire n14498;
	wire n14499;
	wire n14500;
	wire n14501;
	wire n14502;
	wire n14503;
	wire n14504;
	wire n14505;
	wire n14506;
	wire n14507;
	wire n14508;
	wire n14509;
	wire n14510;
	wire n14511;
	wire n14512;
	wire n14513;
	wire n14514;
	wire n14515;
	wire n14516;
	wire n14517;
	wire n14518;
	wire n14519;
	wire n14520;
	wire n14521;
	wire n14522;
	wire n14523;
	wire n14524;
	wire n14525;
	wire n14526;
	wire n14527;
	wire n14528;
	wire n14529;
	wire n14530;
	wire n14531;
	wire n14532;
	wire n14533;
	wire n14534;
	wire n14535;
	wire n14536;
	wire n14537;
	wire n14538;
	wire n14539;
	wire n14540;
	wire n14541;
	wire n14542;
	wire n14543;
	wire n14544;
	wire n14545;
	wire n14546;
	wire n14547;
	wire n14548;
	wire n14549;
	wire n14550;
	wire n14551;
	wire n14552;
	wire n14553;
	wire n14554;
	wire n14555;
	wire n14556;
	wire n14557;
	wire n14558;
	wire n14559;
	wire n14560;
	wire n14561;
	wire n14562;
	wire n14563;
	wire n14564;
	wire n14565;
	wire n14566;
	wire n14567;
	wire n14568;
	wire n14569;
	wire n14570;
	wire n14571;
	wire n14572;
	wire n14573;
	wire n14574;
	wire n14575;
	wire n14576;
	wire n14577;
	wire n14578;
	wire n14579;
	wire n14580;
	wire n14581;
	wire n14582;
	wire n14583;
	wire n14584;
	wire n14585;
	wire n14586;
	wire n14587;
	wire n14588;
	wire n14589;
	wire n14590;
	wire n14591;
	wire n14592;
	wire n14593;
	wire n14594;
	wire n14595;
	wire n14596;
	wire n14597;
	wire n14598;
	wire n14599;
	wire n14600;
	wire n14601;
	wire n14602;
	wire n14603;
	wire n14604;
	wire n14605;
	wire n14606;
	wire n14607;
	wire n14608;
	wire n14609;
	wire n14610;
	wire n14611;
	wire n14612;
	wire n14613;
	wire n14614;
	wire n14615;
	wire n14616;
	wire n14617;
	wire n14618;
	wire n14619;
	wire n14620;
	wire n14621;
	wire n14622;
	wire n14623;
	wire n14624;
	wire n14625;
	wire n14626;
	wire n14627;
	wire n14628;
	wire n14629;
	wire n14630;
	wire n14631;
	wire n14632;
	wire n14633;
	wire n14634;
	wire n14635;
	wire n14636;
	wire n14637;
	wire n14638;
	wire n14639;
	wire n14640;
	wire n14641;
	wire n14642;
	wire n14643;
	wire n14644;
	wire n14645;
	wire n14646;
	wire n14647;
	wire n14648;
	wire n14649;
	wire n14650;
	wire n14651;
	wire n14652;
	wire n14653;
	wire n14654;
	wire n14655;
	wire n14656;
	wire n14657;
	wire n14658;
	wire n14659;
	wire n14660;
	wire n14661;
	wire n14662;
	wire n14663;
	wire n14664;
	wire n14665;
	wire n14666;
	wire n14667;
	wire n14668;
	wire n14669;
	wire n14670;
	wire n14671;
	wire n14672;
	wire n14674;
	wire n14675;
	wire n14676;
	wire n14677;
	wire n14678;
	wire n14679;
	wire n14680;
	wire n14681;
	wire n14682;
	wire n14683;
	wire n14684;
	wire n14685;
	wire n14686;
	wire n14687;
	wire n14688;
	wire n14689;
	wire n14690;
	wire n14691;
	wire n14692;
	wire n14693;
	wire n14694;
	wire n14695;
	wire n14696;
	wire n14697;
	wire n14698;
	wire n14699;
	wire n14700;
	wire n14701;
	wire n14702;
	wire n14703;
	wire n14704;
	wire n14705;
	wire n14706;
	wire n14707;
	wire n14708;
	wire n14709;
	wire n14710;
	wire n14711;
	wire n14712;
	wire n14713;
	wire n14714;
	wire n14715;
	wire n14716;
	wire n14717;
	wire n14718;
	wire n14719;
	wire n14720;
	wire n14721;
	wire n14722;
	wire n14723;
	wire n14724;
	wire n14725;
	wire n14726;
	wire n14727;
	wire n14728;
	wire n14729;
	wire n14730;
	wire n14731;
	wire n14732;
	wire n14733;
	wire n14734;
	wire n14735;
	wire n14736;
	wire n14737;
	wire n14738;
	wire n14739;
	wire n14740;
	wire n14741;
	wire n14742;
	wire n14743;
	wire n14744;
	wire n14745;
	wire n14746;
	wire n14747;
	wire n14748;
	wire n14749;
	wire n14750;
	wire n14751;
	wire n14752;
	wire n14753;
	wire n14754;
	wire n14755;
	wire n14756;
	wire n14757;
	wire n14758;
	wire n14759;
	wire n14760;
	wire n14761;
	wire n14762;
	wire n14763;
	wire n14764;
	wire n14765;
	wire n14766;
	wire n14767;
	wire n14768;
	wire n14769;
	wire n14770;
	wire n14771;
	wire n14772;
	wire n14773;
	wire n14774;
	wire n14775;
	wire n14776;
	wire n14777;
	wire n14778;
	wire n14779;
	wire n14780;
	wire n14781;
	wire n14782;
	wire n14783;
	wire n14784;
	wire n14785;
	wire n14786;
	wire n14787;
	wire n14788;
	wire n14789;
	wire n14790;
	wire n14791;
	wire n14792;
	wire n14793;
	wire n14794;
	wire n14795;
	wire n14796;
	wire n14797;
	wire n14798;
	wire n14799;
	wire n14800;
	wire n14801;
	wire n14802;
	wire n14803;
	wire n14804;
	wire n14805;
	wire n14806;
	wire n14807;
	wire n14808;
	wire n14809;
	wire n14810;
	wire n14811;
	wire n14812;
	wire n14813;
	wire n14814;
	wire n14815;
	wire n14816;
	wire n14817;
	wire n14818;
	wire n14819;
	wire n14820;
	wire n14821;
	wire n14822;
	wire n14823;
	wire n14824;
	wire n14825;
	wire n14826;
	wire n14827;
	wire n14828;
	wire n14829;
	wire n14830;
	wire n14831;
	wire n14832;
	wire n14833;
	wire n14834;
	wire n14835;
	wire n14836;
	wire n14837;
	wire n14838;
	wire n14839;
	wire n14840;
	wire n14841;
	wire n14842;
	wire n14843;
	wire n14844;
	wire n14845;
	wire n14846;
	wire n14847;
	wire n14848;
	wire n14849;
	wire n14850;
	wire n14851;
	wire n14852;
	wire n14853;
	wire n14854;
	wire n14855;
	wire n14856;
	wire n14857;
	wire n14858;
	wire n14859;
	wire n14860;
	wire n14861;
	wire n14862;
	wire n14863;
	wire n14864;
	wire n14865;
	wire n14866;
	wire n14867;
	wire n14868;
	wire n14869;
	wire n14870;
	wire n14871;
	wire n14872;
	wire n14873;
	wire n14874;
	wire n14875;
	wire n14876;
	wire n14877;
	wire n14878;
	wire n14879;
	wire n14880;
	wire n14881;
	wire n14882;
	wire n14883;
	wire n14884;
	wire n14885;
	wire n14886;
	wire n14887;
	wire n14888;
	wire n14889;
	wire n14890;
	wire n14891;
	wire n14892;
	wire n14893;
	wire n14894;
	wire n14895;
	wire n14896;
	wire n14897;
	wire n14898;
	wire n14899;
	wire n14900;
	wire n14901;
	wire n14902;
	wire n14903;
	wire n14904;
	wire n14905;
	wire n14906;
	wire n14907;
	wire n14908;
	wire n14909;
	wire n14910;
	wire n14911;
	wire n14912;
	wire n14913;
	wire n14914;
	wire n14915;
	wire n14916;
	wire n14917;
	wire n14918;
	wire n14919;
	wire n14920;
	wire n14921;
	wire n14922;
	wire n14923;
	wire n14924;
	wire n14925;
	wire n14926;
	wire n14927;
	wire n14928;
	wire n14929;
	wire n14930;
	wire n14931;
	wire n14932;
	wire n14933;
	wire n14934;
	wire n14935;
	wire n14936;
	wire n14937;
	wire n14938;
	wire n14939;
	wire n14940;
	wire n14941;
	wire n14942;
	wire n14943;
	wire n14944;
	wire n14945;
	wire n14946;
	wire n14947;
	wire n14948;
	wire n14949;
	wire n14950;
	wire n14951;
	wire n14952;
	wire n14953;
	wire n14954;
	wire n14955;
	wire n14956;
	wire n14957;
	wire n14958;
	wire n14959;
	wire n14960;
	wire n14961;
	wire n14962;
	wire n14963;
	wire n14964;
	wire n14965;
	wire n14966;
	wire n14967;
	wire n14968;
	wire n14969;
	wire n14970;
	wire n14971;
	wire n14972;
	wire n14973;
	wire n14974;
	wire n14975;
	wire n14976;
	wire n14977;
	wire n14978;
	wire n14979;
	wire n14980;
	wire n14981;
	wire n14982;
	wire n14983;
	wire n14984;
	wire n14985;
	wire n14986;
	wire n14987;
	wire n14988;
	wire n14989;
	wire n14990;
	wire n14991;
	wire n14992;
	wire n14993;
	wire n14994;
	wire n14995;
	wire n14996;
	wire n14997;
	wire n14998;
	wire n14999;
	wire n15000;
	wire n15001;
	wire n15002;
	wire n15003;
	wire n15004;
	wire n15005;
	wire n15006;
	wire n15007;
	wire n15008;
	wire n15009;
	wire n15010;
	wire n15011;
	wire n15012;
	wire n15013;
	wire n15014;
	wire n15015;
	wire n15016;
	wire n15017;
	wire n15018;
	wire n15019;
	wire n15020;
	wire n15021;
	wire n15022;
	wire n15023;
	wire n15024;
	wire n15025;
	wire n15026;
	wire n15027;
	wire n15028;
	wire n15029;
	wire n15030;
	wire n15031;
	wire n15032;
	wire n15033;
	wire n15034;
	wire n15035;
	wire n15036;
	wire n15037;
	wire n15038;
	wire n15039;
	wire n15040;
	wire n15041;
	wire n15042;
	wire n15043;
	wire n15044;
	wire n15045;
	wire n15046;
	wire n15047;
	wire n15048;
	wire n15049;
	wire n15050;
	wire n15051;
	wire n15052;
	wire n15053;
	wire n15054;
	wire n15055;
	wire n15056;
	wire n15057;
	wire n15058;
	wire n15059;
	wire n15060;
	wire n15061;
	wire n15062;
	wire n15063;
	wire n15064;
	wire n15065;
	wire n15066;
	wire n15067;
	wire n15068;
	wire n15069;
	wire n15070;
	wire n15071;
	wire n15072;
	wire n15073;
	wire n15074;
	wire n15075;
	wire n15076;
	wire n15077;
	wire n15078;
	wire n15079;
	wire n15080;
	wire n15081;
	wire n15082;
	wire n15083;
	wire n15084;
	wire n15085;
	wire n15086;
	wire n15087;
	wire n15088;
	wire n15089;
	wire n15090;
	wire n15091;
	wire n15092;
	wire n15093;
	wire n15094;
	wire n15095;
	wire n15096;
	wire n15097;
	wire n15098;
	wire n15099;
	wire n15100;
	wire n15101;
	wire n15102;
	wire n15103;
	wire n15104;
	wire n15105;
	wire n15106;
	wire n15107;
	wire n15108;
	wire n15109;
	wire n15110;
	wire n15111;
	wire n15112;
	wire n15113;
	wire n15114;
	wire n15115;
	wire n15116;
	wire n15117;
	wire n15118;
	wire n15119;
	wire n15120;
	wire n15121;
	wire n15122;
	wire n15123;
	wire n15124;
	wire n15125;
	wire n15126;
	wire n15127;
	wire n15128;
	wire n15129;
	wire n15130;
	wire n15131;
	wire n15132;
	wire n15133;
	wire n15134;
	wire n15135;
	wire n15136;
	wire n15137;
	wire n15138;
	wire n15139;
	wire n15140;
	wire n15141;
	wire n15142;
	wire n15143;
	wire n15144;
	wire n15145;
	wire n15146;
	wire n15147;
	wire n15148;
	wire n15149;
	wire n15150;
	wire n15151;
	wire n15152;
	wire n15153;
	wire n15154;
	wire n15155;
	wire n15156;
	wire n15157;
	wire n15158;
	wire n15159;
	wire n15160;
	wire n15161;
	wire n15162;
	wire n15163;
	wire n15164;
	wire n15165;
	wire n15166;
	wire n15167;
	wire n15168;
	wire n15169;
	wire n15170;
	wire n15171;
	wire n15172;
	wire n15173;
	wire n15174;
	wire n15175;
	wire n15176;
	wire n15177;
	wire n15178;
	wire n15179;
	wire n15180;
	wire n15181;
	wire n15182;
	wire n15183;
	wire n15184;
	wire n15185;
	wire n15186;
	wire n15187;
	wire n15188;
	wire n15189;
	wire n15190;
	wire n15191;
	wire n15192;
	wire n15193;
	wire n15194;
	wire n15195;
	wire n15196;
	wire n15197;
	wire n15198;
	wire n15199;
	wire n15200;
	wire n15201;
	wire n15202;
	wire n15203;
	wire n15204;
	wire n15205;
	wire n15206;
	wire n15207;
	wire n15208;
	wire n15209;
	wire n15210;
	wire n15211;
	wire n15212;
	wire n15213;
	wire n15214;
	wire n15215;
	wire n15216;
	wire n15217;
	wire n15218;
	wire n15219;
	wire n15220;
	wire n15221;
	wire n15222;
	wire n15223;
	wire n15224;
	wire n15225;
	wire n15226;
	wire n15227;
	wire n15228;
	wire n15229;
	wire n15230;
	wire n15231;
	wire n15232;
	wire n15233;
	wire n15234;
	wire n15235;
	wire n15236;
	wire n15237;
	wire n15238;
	wire n15239;
	wire n15240;
	wire n15241;
	wire n15242;
	wire n15243;
	wire n15244;
	wire n15245;
	wire n15247;
	wire n15248;
	wire n15249;
	wire n15250;
	wire n15251;
	wire n15252;
	wire n15253;
	wire n15254;
	wire n15255;
	wire n15256;
	wire n15257;
	wire n15258;
	wire n15259;
	wire n15260;
	wire n15261;
	wire n15262;
	wire n15263;
	wire n15264;
	wire n15265;
	wire n15266;
	wire n15267;
	wire n15268;
	wire n15269;
	wire n15270;
	wire n15271;
	wire n15272;
	wire n15273;
	wire n15274;
	wire n15275;
	wire n15276;
	wire n15277;
	wire n15278;
	wire n15279;
	wire n15280;
	wire n15281;
	wire n15282;
	wire n15283;
	wire n15284;
	wire n15285;
	wire n15286;
	wire n15287;
	wire n15288;
	wire n15289;
	wire n15290;
	wire n15291;
	wire n15292;
	wire n15293;
	wire n15294;
	wire n15295;
	wire n15296;
	wire n15297;
	wire n15298;
	wire n15299;
	wire n15300;
	wire n15301;
	wire n15302;
	wire n15303;
	wire n15304;
	wire n15305;
	wire n15306;
	wire n15307;
	wire n15308;
	wire n15309;
	wire n15310;
	wire n15311;
	wire n15312;
	wire n15313;
	wire n15314;
	wire n15315;
	wire n15316;
	wire n15317;
	wire n15318;
	wire n15319;
	wire n15320;
	wire n15321;
	wire n15322;
	wire n15323;
	wire n15324;
	wire n15325;
	wire n15326;
	wire n15327;
	wire n15328;
	wire n15329;
	wire n15330;
	wire n15331;
	wire n15332;
	wire n15333;
	wire n15334;
	wire n15335;
	wire n15336;
	wire n15337;
	wire n15338;
	wire n15339;
	wire n15340;
	wire n15341;
	wire n15342;
	wire n15343;
	wire n15344;
	wire n15345;
	wire n15346;
	wire n15347;
	wire n15348;
	wire n15349;
	wire n15350;
	wire n15351;
	wire n15352;
	wire n15353;
	wire n15354;
	wire n15355;
	wire n15356;
	wire n15357;
	wire n15358;
	wire n15359;
	wire n15360;
	wire n15361;
	wire n15362;
	wire n15363;
	wire n15364;
	wire n15365;
	wire n15366;
	wire n15367;
	wire n15368;
	wire n15369;
	wire n15370;
	wire n15371;
	wire n15372;
	wire n15373;
	wire n15374;
	wire n15375;
	wire n15376;
	wire n15377;
	wire n15378;
	wire n15379;
	wire n15380;
	wire n15381;
	wire n15382;
	wire n15383;
	wire n15384;
	wire n15385;
	wire n15386;
	wire n15387;
	wire n15388;
	wire n15389;
	wire n15390;
	wire n15391;
	wire n15392;
	wire n15393;
	wire n15394;
	wire n15395;
	wire n15396;
	wire n15397;
	wire n15398;
	wire n15399;
	wire n15400;
	wire n15401;
	wire n15402;
	wire n15403;
	wire n15404;
	wire n15405;
	wire n15406;
	wire n15407;
	wire n15408;
	wire n15409;
	wire n15410;
	wire n15411;
	wire n15412;
	wire n15413;
	wire n15414;
	wire n15415;
	wire n15416;
	wire n15417;
	wire n15418;
	wire n15419;
	wire n15420;
	wire n15421;
	wire n15422;
	wire n15423;
	wire n15424;
	wire n15425;
	wire n15426;
	wire n15427;
	wire n15428;
	wire n15429;
	wire n15430;
	wire n15431;
	wire n15432;
	wire n15433;
	wire n15434;
	wire n15435;
	wire n15436;
	wire n15437;
	wire n15438;
	wire n15439;
	wire n15440;
	wire n15441;
	wire n15442;
	wire n15443;
	wire n15444;
	wire n15445;
	wire n15446;
	wire n15447;
	wire n15448;
	wire n15449;
	wire n15450;
	wire n15451;
	wire n15452;
	wire n15453;
	wire n15454;
	wire n15455;
	wire n15456;
	wire n15457;
	wire n15458;
	wire n15459;
	wire n15460;
	wire n15461;
	wire n15462;
	wire n15463;
	wire n15464;
	wire n15465;
	wire n15466;
	wire n15467;
	wire n15468;
	wire n15469;
	wire n15470;
	wire n15471;
	wire n15472;
	wire n15473;
	wire n15474;
	wire n15475;
	wire n15476;
	wire n15477;
	wire n15478;
	wire n15479;
	wire n15480;
	wire n15481;
	wire n15482;
	wire n15483;
	wire n15484;
	wire n15485;
	wire n15486;
	wire n15487;
	wire n15488;
	wire n15489;
	wire n15490;
	wire n15491;
	wire n15492;
	wire n15493;
	wire n15494;
	wire n15495;
	wire n15496;
	wire n15497;
	wire n15498;
	wire n15499;
	wire n15500;
	wire n15501;
	wire n15502;
	wire n15503;
	wire n15504;
	wire n15505;
	wire n15506;
	wire n15507;
	wire n15508;
	wire n15509;
	wire n15510;
	wire n15511;
	wire n15512;
	wire n15513;
	wire n15514;
	wire n15515;
	wire n15516;
	wire n15517;
	wire n15518;
	wire n15519;
	wire n15520;
	wire n15521;
	wire n15522;
	wire n15523;
	wire n15524;
	wire n15525;
	wire n15526;
	wire n15527;
	wire n15528;
	wire n15529;
	wire n15530;
	wire n15531;
	wire n15532;
	wire n15533;
	wire n15534;
	wire n15535;
	wire n15536;
	wire n15537;
	wire n15538;
	wire n15539;
	wire n15540;
	wire n15541;
	wire n15542;
	wire n15543;
	wire n15544;
	wire n15545;
	wire n15546;
	wire n15547;
	wire n15548;
	wire n15549;
	wire n15550;
	wire n15551;
	wire n15552;
	wire n15553;
	wire n15554;
	wire n15555;
	wire n15556;
	wire n15557;
	wire n15558;
	wire n15559;
	wire n15560;
	wire n15561;
	wire n15562;
	wire n15563;
	wire n15564;
	wire n15565;
	wire n15566;
	wire n15567;
	wire n15568;
	wire n15569;
	wire n15570;
	wire n15571;
	wire n15572;
	wire n15573;
	wire n15574;
	wire n15575;
	wire n15576;
	wire n15577;
	wire n15578;
	wire n15579;
	wire n15580;
	wire n15581;
	wire n15582;
	wire n15583;
	wire n15584;
	wire n15585;
	wire n15586;
	wire n15587;
	wire n15588;
	wire n15589;
	wire n15590;
	wire n15591;
	wire n15592;
	wire n15593;
	wire n15594;
	wire n15595;
	wire n15596;
	wire n15597;
	wire n15598;
	wire n15599;
	wire n15600;
	wire n15601;
	wire n15602;
	wire n15603;
	wire n15604;
	wire n15605;
	wire n15606;
	wire n15607;
	wire n15608;
	wire n15609;
	wire n15610;
	wire n15611;
	wire n15612;
	wire n15613;
	wire n15614;
	wire n15615;
	wire n15616;
	wire n15617;
	wire n15618;
	wire n15619;
	wire n15620;
	wire n15621;
	wire n15622;
	wire n15623;
	wire n15624;
	wire n15625;
	wire n15626;
	wire n15627;
	wire n15628;
	wire n15629;
	wire n15630;
	wire n15631;
	wire n15632;
	wire n15633;
	wire n15634;
	wire n15635;
	wire n15636;
	wire n15637;
	wire n15638;
	wire n15639;
	wire n15641;
	wire n15642;
	wire n15643;
	wire n15644;
	wire n15645;
	wire n15646;
	wire n15647;
	wire n15648;
	wire n15649;
	wire n15650;
	wire n15651;
	wire n15652;
	wire n15653;
	wire n15654;
	wire n15655;
	wire n15656;
	wire n15657;
	wire n15658;
	wire n15659;
	wire n15660;
	wire n15661;
	wire n15662;
	wire n15663;
	wire n15664;
	wire n15665;
	wire n15666;
	wire n15667;
	wire n15668;
	wire n15669;
	wire n15670;
	wire n15671;
	wire n15672;
	wire n15673;
	wire n15674;
	wire n15675;
	wire n15676;
	wire n15677;
	wire n15678;
	wire n15679;
	wire n15680;
	wire n15681;
	wire n15682;
	wire n15683;
	wire n15684;
	wire n15685;
	wire n15686;
	wire n15687;
	wire n15688;
	wire n15689;
	wire n15690;
	wire n15691;
	wire n15692;
	wire n15693;
	wire n15694;
	wire n15695;
	wire n15696;
	wire n15697;
	wire n15698;
	wire n15699;
	wire n15700;
	wire n15701;
	wire n15702;
	wire n15703;
	wire n15704;
	wire n15705;
	wire n15706;
	wire n15707;
	wire n15708;
	wire n15709;
	wire n15710;
	wire n15711;
	wire n15712;
	wire n15713;
	wire n15714;
	wire n15715;
	wire n15716;
	wire n15717;
	wire n15718;
	wire n15719;
	wire n15720;
	wire n15721;
	wire n15722;
	wire n15723;
	wire n15724;
	wire n15725;
	wire n15726;
	wire n15727;
	wire n15728;
	wire n15729;
	wire n15730;
	wire n15731;
	wire n15732;
	wire n15733;
	wire n15734;
	wire n15735;
	wire n15736;
	wire n15737;
	wire n15738;
	wire n15739;
	wire n15740;
	wire n15741;
	wire n15742;
	wire n15743;
	wire n15744;
	wire n15745;
	wire n15746;
	wire n15747;
	wire n15748;
	wire n15749;
	wire n15750;
	wire n15751;
	wire n15752;
	wire n15753;
	wire n15754;
	wire n15755;
	wire n15756;
	wire n15757;
	wire n15758;
	wire n15759;
	wire n15760;
	wire n15761;
	wire n15762;
	wire n15763;
	wire n15764;
	wire n15765;
	wire n15766;
	wire n15767;
	wire n15768;
	wire n15769;
	wire n15770;
	wire n15771;
	wire n15772;
	wire n15773;
	wire n15774;
	wire n15775;
	wire n15776;
	wire n15777;
	wire n15778;
	wire n15779;
	wire n15780;
	wire n15781;
	wire n15782;
	wire n15783;
	wire n15784;
	wire n15785;
	wire n15786;
	wire n15787;
	wire n15788;
	wire n15789;
	wire n15790;
	wire n15791;
	wire n15792;
	wire n15793;
	wire n15794;
	wire n15795;
	wire n15796;
	wire n15797;
	wire n15798;
	wire n15799;
	wire n15800;
	wire n15801;
	wire n15802;
	wire n15803;
	wire n15804;
	wire n15805;
	wire n15806;
	wire n15807;
	wire n15808;
	wire n15809;
	wire n15810;
	wire n15811;
	wire n15812;
	wire n15813;
	wire n15814;
	wire n15815;
	wire n15816;
	wire n15817;
	wire n15818;
	wire n15819;
	wire n15820;
	wire n15821;
	wire n15822;
	wire n15823;
	wire n15824;
	wire n15825;
	wire n15826;
	wire n15827;
	wire n15828;
	wire n15829;
	wire n15830;
	wire n15831;
	wire n15832;
	wire n15833;
	wire n15834;
	wire n15835;
	wire n15836;
	wire n15837;
	wire n15838;
	wire n15839;
	wire n15840;
	wire n15841;
	wire n15842;
	wire n15843;
	wire n15844;
	wire n15845;
	wire n15846;
	wire n15847;
	wire n15848;
	wire n15849;
	wire n15850;
	wire n15851;
	wire n15852;
	wire n15853;
	wire n15854;
	wire n15855;
	wire n15856;
	wire n15857;
	wire n15858;
	wire n15859;
	wire n15860;
	wire n15861;
	wire n15862;
	wire n15863;
	wire n15864;
	wire n15865;
	wire n15866;
	wire n15867;
	wire n15868;
	wire n15869;
	wire n15870;
	wire n15871;
	wire n15872;
	wire n15873;
	wire n15874;
	wire n15875;
	wire n15876;
	wire n15877;
	wire n15878;
	wire n15879;
	wire n15880;
	wire n15881;
	wire n15882;
	wire n15883;
	wire n15884;
	wire n15885;
	wire n15886;
	wire n15887;
	wire n15888;
	wire n15889;
	wire n15890;
	wire n15891;
	wire n15892;
	wire n15893;
	wire n15894;
	wire n15895;
	wire n15896;
	wire n15897;
	wire n15898;
	wire n15899;
	wire n15900;
	wire n15901;
	wire n15902;
	wire n15903;
	wire n15904;
	wire n15905;
	wire n15906;
	wire n15907;
	wire n15908;
	wire n15909;
	wire n15910;
	wire n15911;
	wire n15912;
	wire n15913;
	wire n15914;
	wire n15915;
	wire n15916;
	wire n15917;
	wire n15918;
	wire n15919;
	wire n15920;
	wire n15921;
	wire n15922;
	wire n15923;
	wire n15924;
	wire n15925;
	wire n15926;
	wire n15927;
	wire n15928;
	wire n15929;
	wire n15930;
	wire n15931;
	wire n15932;
	wire n15933;
	wire n15934;
	wire n15935;
	wire n15936;
	wire n15937;
	wire n15938;
	wire n15939;
	wire n15940;
	wire n15941;
	wire n15942;
	wire n15943;
	wire n15944;
	wire n15945;
	wire n15946;
	wire n15947;
	wire n15948;
	wire n15949;
	wire n15950;
	wire n15951;
	wire n15952;
	wire n15953;
	wire n15954;
	wire n15955;
	wire n15956;
	wire n15957;
	wire n15958;
	wire n15959;
	wire n15960;
	wire n15961;
	wire n15962;
	wire n15963;
	wire n15964;
	wire n15965;
	wire n15966;
	wire n15967;
	wire n15968;
	wire n15969;
	wire n15970;
	wire n15971;
	wire n15972;
	wire n15973;
	wire n15974;
	wire n15975;
	wire n15976;
	wire n15977;
	wire n15978;
	wire n15979;
	wire n15980;
	wire n15981;
	wire n15982;
	wire n15983;
	wire n15984;
	wire n15985;
	wire n15986;
	wire n15987;
	wire n15988;
	wire n15989;
	wire n15990;
	wire n15991;
	wire n15992;
	wire n15993;
	wire n15994;
	wire n15995;
	wire n15996;
	wire n15997;
	wire n15998;
	wire n15999;
	wire n16000;
	wire n16001;
	wire n16002;
	wire n16003;
	wire n16004;
	wire n16005;
	wire n16006;
	wire n16007;
	wire n16008;
	wire n16009;
	wire n16010;
	wire n16011;
	wire n16012;
	wire n16013;
	wire n16014;
	wire n16015;
	wire n16016;
	wire n16017;
	wire n16018;
	wire n16019;
	wire n16020;
	wire n16021;
	wire n16022;
	wire n16023;
	wire n16024;
	wire n16025;
	wire n16026;
	wire n16027;
	wire n16028;
	wire n16029;
	wire n16030;
	wire n16031;
	wire n16032;
	wire n16033;
	wire n16034;
	wire n16035;
	wire n16036;
	wire n16037;
	wire n16038;
	wire n16039;
	wire n16040;
	wire n16041;
	wire n16042;
	wire n16043;
	wire n16044;
	wire n16045;
	wire n16046;
	wire n16047;
	wire n16048;
	wire n16049;
	wire n16050;
	wire n16051;
	wire n16052;
	wire n16053;
	wire n16054;
	wire n16055;
	wire n16056;
	wire n16057;
	wire n16058;
	wire n16059;
	wire n16060;
	wire n16061;
	wire n16062;
	wire n16063;
	wire n16064;
	wire n16065;
	wire n16066;
	wire n16067;
	wire n16068;
	wire n16069;
	wire n16070;
	wire n16071;
	wire n16072;
	wire n16073;
	wire n16074;
	wire n16075;
	wire n16076;
	wire n16077;
	wire n16078;
	wire n16079;
	wire n16080;
	wire n16081;
	wire n16082;
	wire n16083;
	wire n16084;
	wire n16085;
	wire n16086;
	wire n16087;
	wire n16088;
	wire n16089;
	wire n16090;
	wire n16091;
	wire n16092;
	wire n16093;
	wire n16094;
	wire n16095;
	wire n16096;
	wire n16097;
	wire n16098;
	wire n16099;
	wire n16100;
	wire n16101;
	wire n16102;
	wire n16103;
	wire n16104;
	wire n16105;
	wire n16106;
	wire n16107;
	wire n16108;
	wire n16109;
	wire n16110;
	wire n16111;
	wire n16112;
	wire n16113;
	wire n16114;
	wire n16115;
	wire n16116;
	wire n16117;
	wire n16118;
	wire n16119;
	wire n16120;
	wire n16121;
	wire n16122;
	wire n16123;
	wire n16124;
	wire n16125;
	wire n16126;
	wire n16127;
	wire n16128;
	wire n16129;
	wire n16130;
	wire n16131;
	wire n16132;
	wire n16133;
	wire n16134;
	wire n16135;
	wire n16136;
	wire n16137;
	wire n16138;
	wire n16139;
	wire n16140;
	wire n16141;
	wire n16142;
	wire n16143;
	wire n16144;
	wire n16145;
	wire n16146;
	wire n16147;
	wire n16148;
	wire n16149;
	wire n16150;
	wire n16151;
	wire n16152;
	wire n16153;
	wire n16154;
	wire n16155;
	wire n16156;
	wire n16157;
	wire n16158;
	wire n16159;
	wire n16160;
	wire n16161;
	wire n16162;
	wire n16163;
	wire n16164;
	wire n16165;
	wire n16166;
	wire n16167;
	wire n16168;
	wire n16169;
	wire n16170;
	wire n16171;
	wire n16172;
	wire n16173;
	wire n16174;
	wire n16175;
	wire n16176;
	wire n16177;
	wire n16178;
	wire n16179;
	wire n16180;
	wire n16181;
	wire n16182;
	wire n16183;
	wire n16184;
	wire n16185;
	wire n16186;
	wire n16187;
	wire n16188;
	wire n16189;
	wire n16190;
	wire n16191;
	wire n16192;
	wire n16193;
	wire n16194;
	wire n16195;
	wire n16196;
	wire n16197;
	wire n16198;
	wire n16199;
	wire n16200;
	wire n16201;
	wire n16202;
	wire n16203;
	wire n16204;
	wire n16205;
	wire n16206;
	wire n16207;
	wire n16208;
	wire n16209;
	wire n16210;
	wire n16211;
	wire n16212;
	wire n16213;
	wire n16214;
	wire n16215;
	wire n16216;
	wire n16217;
	wire n16218;
	wire n16219;
	wire n16220;
	wire n16221;
	wire n16222;
	wire n16223;
	wire n16224;
	wire n16225;
	wire n16226;
	wire n16227;
	wire n16228;
	wire n16229;
	wire n16230;
	wire n16231;
	wire n16232;
	wire n16233;
	wire n16234;
	wire n16235;
	wire n16236;
	wire n16237;
	wire n16238;
	wire n16239;
	wire n16240;
	wire n16241;
	wire n16242;
	wire n16243;
	wire n16244;
	wire n16245;
	wire n16246;
	wire n16247;
	wire n16248;
	wire n16249;
	wire n16250;
	wire n16251;
	wire n16252;
	wire n16253;
	wire n16254;
	wire n16255;
	wire n16256;
	wire n16257;
	wire n16258;
	wire n16259;
	wire n16260;
	wire n16261;
	wire n16262;
	wire n16263;
	wire n16264;
	wire n16265;
	wire n16266;
	wire n16267;
	wire n16268;
	wire n16269;
	wire n16270;
	wire n16271;
	wire n16272;
	wire n16273;
	wire n16274;
	wire n16275;
	wire n16276;
	wire n16277;
	wire n16278;
	wire n16279;
	wire n16280;
	wire n16281;
	wire n16282;
	wire n16283;
	wire n16284;
	wire n16285;
	wire n16286;
	wire n16287;
	wire n16288;
	wire n16289;
	wire n16290;
	wire n16291;
	wire n16292;
	wire n16293;
	wire n16294;
	wire n16295;
	wire n16296;
	wire n16297;
	wire n16298;
	wire n16299;
	wire n16300;
	wire n16301;
	wire n16302;
	wire n16303;
	wire n16304;
	wire n16305;
	wire n16306;
	wire n16307;
	wire n16308;
	wire n16309;
	wire n16310;
	wire n16311;
	wire n16312;
	wire n16313;
	wire n16314;
	wire n16315;
	wire n16316;
	wire n16317;
	wire n16318;
	wire n16319;
	wire n16320;
	wire n16321;
	wire n16322;
	wire n16323;
	wire n16324;
	wire n16325;
	wire n16326;
	wire n16327;
	wire n16328;
	wire n16329;
	wire n16330;
	wire n16331;
	wire n16332;
	wire n16333;
	wire n16334;
	wire n16335;
	wire n16336;
	wire n16337;
	wire n16338;
	wire n16339;
	wire n16340;
	wire n16341;
	wire n16342;
	wire n16343;
	wire n16344;
	wire n16345;
	wire n16346;
	wire n16347;
	wire n16348;
	wire n16349;
	wire n16350;
	wire n16351;
	wire n16352;
	wire n16353;
	wire n16354;
	wire n16355;
	wire n16356;
	wire n16357;
	wire n16358;
	wire n16359;
	wire n16360;
	wire n16361;
	wire n16362;
	wire n16363;
	wire n16364;
	wire n16365;
	wire n16366;
	wire n16367;
	wire n16368;
	wire n16369;
	wire n16370;
	wire n16371;
	wire n16372;
	wire n16373;
	wire n16374;
	wire n16375;
	wire n16376;
	wire n16377;
	wire n16378;
	wire n16379;
	wire n16380;
	wire n16381;
	wire n16382;
	wire n16383;
	wire n16384;
	wire n16385;
	wire n16386;
	wire n16387;
	wire n16388;
	wire n16389;
	wire n16390;
	wire n16391;
	wire n16392;
	wire n16393;
	wire n16394;
	wire n16395;
	wire n16396;
	wire n16397;
	wire n16398;
	wire n16399;
	wire n16400;
	wire n16401;
	wire n16402;
	wire n16403;
	wire n16404;
	wire n16405;
	wire n16406;
	wire n16407;
	wire n16408;
	wire n16409;
	wire n16410;
	wire n16411;
	wire n16412;
	wire n16413;
	wire n16414;
	wire n16415;
	wire n16416;
	wire n16417;
	wire n16418;
	wire n16419;
	wire n16420;
	wire n16421;
	wire n16422;
	wire n16423;
	wire n16424;
	wire n16425;
	wire n16426;
	wire n16427;
	wire n16428;
	wire n16429;
	wire n16430;
	wire n16431;
	wire n16432;
	wire n16433;
	wire n16434;
	wire n16435;
	wire n16436;
	wire n16437;
	wire n16438;
	wire n16439;
	wire n16440;
	wire n16441;
	wire n16442;
	wire n16443;
	wire n16444;
	wire n16445;
	wire n16446;
	wire n16447;
	wire n16448;
	wire n16449;
	wire n16450;
	wire n16451;
	wire n16452;
	wire n16453;
	wire n16454;
	wire n16455;
	wire n16456;
	wire n16457;
	wire n16458;
	wire n16459;
	wire n16460;
	wire n16461;
	wire n16462;
	wire n16463;
	wire n16464;
	wire n16465;
	wire n16466;
	wire n16467;
	wire n16468;
	wire n16469;
	wire n16470;
	wire n16471;
	wire n16472;
	wire n16473;
	wire n16475;
	wire n16476;
	wire n16477;
	wire n16478;
	wire n16479;
	wire n16480;
	wire n16481;
	wire n16482;
	wire n16483;
	wire n16484;
	wire n16485;
	wire n16486;
	wire n16487;
	wire n16488;
	wire n16489;
	wire n16490;
	wire n16491;
	wire n16492;
	wire n16493;
	wire n16494;
	wire n16495;
	wire n16496;
	wire n16497;
	wire n16498;
	wire n16499;
	wire n16500;
	wire n16501;
	wire n16502;
	wire n16503;
	wire n16504;
	wire n16505;
	wire n16506;
	wire n16507;
	wire n16508;
	wire n16509;
	wire n16510;
	wire n16511;
	wire n16512;
	wire n16513;
	wire n16514;
	wire n16515;
	wire n16516;
	wire n16517;
	wire n16518;
	wire n16519;
	wire n16520;
	wire n16521;
	wire n16522;
	wire n16523;
	wire n16524;
	wire n16525;
	wire n16526;
	wire n16527;
	wire n16528;
	wire n16529;
	wire n16530;
	wire n16531;
	wire n16532;
	wire n16533;
	wire n16534;
	wire n16535;
	wire n16536;
	wire n16537;
	wire n16538;
	wire n16539;
	wire n16540;
	wire n16541;
	wire n16542;
	wire n16543;
	wire n16544;
	wire n16545;
	wire n16546;
	wire n16547;
	wire n16548;
	wire n16549;
	wire n16550;
	wire n16551;
	wire n16552;
	wire n16553;
	wire n16554;
	wire n16555;
	wire n16556;
	wire n16557;
	wire n16558;
	wire n16559;
	wire n16560;
	wire n16561;
	wire n16562;
	wire n16563;
	wire n16564;
	wire n16565;
	wire n16566;
	wire n16567;
	wire n16568;
	wire n16569;
	wire n16570;
	wire n16571;
	wire n16572;
	wire n16573;
	wire n16574;
	wire n16575;
	wire n16576;
	wire n16577;
	wire n16578;
	wire n16579;
	wire n16580;
	wire n16581;
	wire n16582;
	wire n16583;
	wire n16584;
	wire n16585;
	wire n16586;
	wire n16587;
	wire n16588;
	wire n16589;
	wire n16590;
	wire n16591;
	wire n16592;
	wire n16593;
	wire n16594;
	wire n16595;
	wire n16596;
	wire n16597;
	wire n16598;
	wire n16599;
	wire n16600;
	wire n16601;
	wire n16602;
	wire n16603;
	wire n16604;
	wire n16605;
	wire n16606;
	wire n16607;
	wire n16608;
	wire n16609;
	wire n16610;
	wire n16611;
	wire n16612;
	wire n16613;
	wire n16614;
	wire n16615;
	wire n16616;
	wire n16617;
	wire n16618;
	wire n16619;
	wire n16620;
	wire n16621;
	wire n16622;
	wire n16623;
	wire n16624;
	wire n16625;
	wire n16626;
	wire n16627;
	wire n16628;
	wire n16629;
	wire n16630;
	wire n16631;
	wire n16632;
	wire n16633;
	wire n16634;
	wire n16635;
	wire n16636;
	wire n16637;
	wire n16638;
	wire n16639;
	wire n16640;
	wire n16641;
	wire n16642;
	wire n16643;
	wire n16644;
	wire n16645;
	wire n16646;
	wire n16647;
	wire n16648;
	wire n16649;
	wire n16650;
	wire n16651;
	wire n16652;
	wire n16653;
	wire n16654;
	wire n16655;
	wire n16656;
	wire n16657;
	wire n16658;
	wire n16659;
	wire n16660;
	wire n16661;
	wire n16662;
	wire n16663;
	wire n16664;
	wire n16665;
	wire n16666;
	wire n16667;
	wire n16668;
	wire n16669;
	wire n16670;
	wire n16671;
	wire n16672;
	wire n16673;
	wire n16674;
	wire n16675;
	wire n16676;
	wire n16677;
	wire n16678;
	wire n16679;
	wire n16680;
	wire n16681;
	wire n16682;
	wire n16683;
	wire n16684;
	wire n16685;
	wire n16686;
	wire n16687;
	wire n16688;
	wire n16689;
	wire n16690;
	wire n16691;
	wire n16692;
	wire n16693;
	wire n16694;
	wire n16695;
	wire n16696;
	wire n16697;
	wire n16698;
	wire n16699;
	wire n16700;
	wire n16701;
	wire n16702;
	wire n16703;
	wire n16704;
	wire n16705;
	wire n16706;
	wire n16707;
	wire n16708;
	wire n16709;
	wire n16710;
	wire n16711;
	wire n16712;
	wire n16713;
	wire n16714;
	wire n16715;
	wire n16716;
	wire n16717;
	wire n16718;
	wire n16719;
	wire n16720;
	wire n16721;
	wire n16722;
	wire n16723;
	wire n16724;
	wire n16725;
	wire n16726;
	wire n16727;
	wire n16728;
	wire n16729;
	wire n16730;
	wire n16731;
	wire n16732;
	wire n16733;
	wire n16734;
	wire n16735;
	wire n16736;
	wire n16737;
	wire n16738;
	wire n16739;
	wire n16740;
	wire n16741;
	wire n16742;
	wire n16743;
	wire n16744;
	wire n16745;
	wire n16746;
	wire n16747;
	wire n16748;
	wire n16749;
	wire n16750;
	wire n16751;
	wire n16752;
	wire n16753;
	wire n16754;
	wire n16755;
	wire n16756;
	wire n16757;
	wire n16758;
	wire n16759;
	wire n16760;
	wire n16761;
	wire n16762;
	wire n16763;
	wire n16764;
	wire n16765;
	wire n16766;
	wire n16767;
	wire n16768;
	wire n16769;
	wire n16770;
	wire n16771;
	wire n16772;
	wire n16773;
	wire n16774;
	wire n16775;
	wire n16776;
	wire n16777;
	wire n16778;
	wire n16779;
	wire n16780;
	wire n16781;
	wire n16782;
	wire n16783;
	wire n16784;
	wire n16785;
	wire n16786;
	wire n16787;
	wire n16788;
	wire n16789;
	wire n16790;
	wire n16791;
	wire n16792;
	wire n16793;
	wire n16794;
	wire n16795;
	wire n16796;
	wire n16797;
	wire n16798;
	wire n16799;
	wire n16800;
	wire n16801;
	wire n16802;
	wire n16803;
	wire n16804;
	wire n16805;
	wire n16806;
	wire n16807;
	wire n16808;
	wire n16809;
	wire n16810;
	wire n16811;
	wire n16812;
	wire n16813;
	wire n16814;
	wire n16815;
	wire n16816;
	wire n16817;
	wire n16818;
	wire n16819;
	wire n16820;
	wire n16821;
	wire n16822;
	wire n16823;
	wire n16824;
	wire n16825;
	wire n16826;
	wire n16827;
	wire n16828;
	wire n16829;
	wire n16830;
	wire n16831;
	wire n16832;
	wire n16833;
	wire n16834;
	wire n16835;
	wire n16836;
	wire n16837;
	wire n16838;
	wire n16839;
	wire n16840;
	wire n16841;
	wire n16842;
	wire n16843;
	wire n16844;
	wire n16845;
	wire n16846;
	wire n16847;
	wire n16848;
	wire n16849;
	wire n16850;
	wire n16851;
	wire n16852;
	wire n16853;
	wire n16854;
	wire n16855;
	wire n16856;
	wire n16857;
	wire n16858;
	wire n16859;
	wire n16860;
	wire n16861;
	wire n16862;
	wire n16863;
	wire n16864;
	wire n16865;
	wire n16866;
	wire n16867;
	wire n16868;
	wire n16869;
	wire n16871;
	wire n16872;
	wire n16873;
	wire n16874;
	wire n16875;
	wire n16876;
	wire n16877;
	wire n16878;
	wire n16879;
	wire n16880;
	wire n16881;
	wire n16882;
	wire n16885;
	wire n16886;
	wire n16887;
	wire n16888;
	wire n16889;
	wire n16890;
	wire n16891;
	wire n16892;
	wire n16893;
	wire n16894;
	wire n16895;
	wire n16896;
	wire n16898;
	wire n16899;
	wire n16900;
	wire n16901;
	wire n16902;
	wire n16903;
	wire n16904;
	wire n16905;
	wire n16906;
	wire n16907;
	wire n16908;
	wire n16909;
	wire n16910;
	wire n16911;
	wire n16912;
	wire n16913;
	wire n16914;
	wire n16915;
	wire n16916;
	wire n16917;
	wire n16918;
	wire n16919;
	wire n16920;
	wire n16921;
	wire n16922;
	wire n16923;
	wire n16924;
	wire n16925;
	wire n16926;
	wire n16927;
	wire n16928;
	wire n16929;
	wire n16930;
	wire n16931;
	wire n16932;
	wire n16933;
	wire n16934;
	wire n16935;
	wire n16936;
	wire n16937;
	wire n16938;
	wire n16939;
	wire n16940;
	wire n16941;
	wire n16942;
	wire n16943;
	wire n16944;
	wire n16945;
	wire n16946;
	wire n16947;
	wire n16948;
	wire n16949;
	wire n16950;
	wire n16951;
	wire n16952;
	wire n16953;
	wire n16954;
	wire n16955;
	wire n16956;
	wire n16957;
	wire n16958;
	wire n16959;
	wire n16960;
	wire n16961;
	wire n16962;
	wire n16963;
	wire n16964;
	wire n16965;
	wire n16966;
	wire n16967;
	wire n16968;
	wire n16969;
	wire n16970;
	wire n16971;
	wire n16972;
	wire n16973;
	wire n16974;
	wire n16975;
	wire n16976;
	wire n16977;
	wire n16978;
	wire n16979;
	wire n16980;
	wire n16981;
	wire n16982;
	wire n16983;
	wire n16984;
	wire n16985;
	wire n16986;
	wire n16987;
	wire n16988;
	wire n16989;
	wire n16990;
	wire n16991;
	wire n16992;
	wire n16993;
	wire n16994;
	wire n16995;
	wire n16996;
	wire n16997;
	wire n16998;
	wire n16999;
	wire n17000;
	wire n17001;
	wire n17002;
	wire n17003;
	wire n17004;
	wire n17005;
	wire n17006;
	wire n17007;
	wire n17008;
	wire n17009;
	wire n17010;
	wire n17011;
	wire n17012;
	wire n17013;
	wire n17014;
	wire n17015;
	wire n17016;
	wire n17017;
	wire n17018;
	wire n17019;
	wire n17020;
	wire n17021;
	wire n17022;
	wire n17023;
	wire n17024;
	wire n17025;
	wire n17026;
	wire n17027;
	wire n17028;
	wire n17029;
	wire n17030;
	wire n17031;
	wire n17032;
	wire n17033;
	wire n17034;
	wire n17035;
	wire n17036;
	wire n17037;
	wire n17038;
	wire n17039;
	wire n17040;
	wire n17041;
	wire n17042;
	wire n17043;
	wire n17044;
	wire n17045;
	wire n17046;
	wire n17047;
	wire n17048;
	wire n17049;
	wire n17050;
	wire n17051;
	wire n17052;
	wire n17053;
	wire n17054;
	wire n17055;
	wire n17056;
	wire n17057;
	wire n17058;
	wire n17059;
	wire n17060;
	wire n17061;
	wire n17062;
	wire n17063;
	wire n17064;
	wire n17065;
	wire n17066;
	wire n17067;
	wire n17068;
	wire n17069;
	wire n17070;
	wire n17071;
	wire n17072;
	wire n17073;
	wire n17074;
	wire n17075;
	wire n17076;
	wire n17077;
	wire n17078;
	wire n17079;
	wire n17080;
	wire n17081;
	wire n17082;
	wire n17083;
	wire n17084;
	wire n17085;
	wire n17086;
	wire n17087;
	wire n17088;
	wire n17089;
	wire n17090;
	wire n17091;
	wire n17092;
	wire n17093;
	wire n17094;
	wire n17095;
	wire n17096;
	wire n17097;
	wire n17098;
	wire n17099;
	wire n17100;
	wire n17101;
	wire n17102;
	wire n17103;
	wire n17104;
	wire n17105;
	wire n17106;
	wire n17107;
	wire n17108;
	wire n17109;
	wire n17110;
	wire n17111;
	wire n17112;
	wire n17113;
	wire n17114;
	wire n17115;
	wire n17116;
	wire n17117;
	wire n17118;
	wire n17119;
	wire n17120;
	wire n17121;
	wire n17122;
	wire n17123;
	wire n17124;
	wire n17125;
	wire n17126;
	wire n17127;
	wire n17128;
	wire n17129;
	wire n17130;
	wire n17131;
	wire n17132;
	wire n17134;
	wire n17135;
	wire n17136;
	wire n17137;
	wire n17138;
	wire n17139;
	wire n17140;
	wire n17141;
	wire n17142;
	wire n17143;
	wire n17144;
	wire n17145;
	wire n17146;
	wire n17147;
	wire n17148;
	wire n17149;
	wire n17150;
	wire n17151;
	wire n17152;
	wire n17153;
	wire n17154;
	wire n17155;
	wire n17156;
	wire n17157;
	wire n17158;
	wire n17159;
	wire n17160;
	wire n17161;
	wire n17162;
	wire n17163;
	wire n17164;
	wire n17165;
	wire n17166;
	wire n17167;
	wire n17168;
	wire n17169;
	wire n17170;
	wire n17171;
	wire n17172;
	wire n17173;
	wire n17174;
	wire n17175;
	wire n17176;
	wire n17177;
	wire n17178;
	wire n17179;
	wire n17180;
	wire n17181;
	wire n17182;
	wire n17183;
	wire n17184;
	wire n17185;
	wire n17186;
	wire n17187;
	wire n17188;
	wire n17189;
	wire n17190;
	wire n17191;
	wire n17192;
	wire n17193;
	wire n17194;
	wire n17195;
	wire n17196;
	wire n17197;
	wire n17198;
	wire n17199;
	wire n17200;
	wire n17201;
	wire n17202;
	wire n17203;
	wire n17204;
	wire n17205;
	wire n17206;
	wire n17207;
	wire n17208;
	wire n17209;
	wire n17210;
	wire n17211;
	wire n17212;
	wire n17213;
	wire n17214;
	wire n17215;
	wire n17216;
	wire n17217;
	wire n17218;
	wire n17219;
	wire n17220;
	wire n17221;
	wire n17222;
	wire n17223;
	wire n17224;
	wire n17225;
	wire n17226;
	wire n17227;
	wire n17228;
	wire n17229;
	wire n17230;
	wire n17231;
	wire n17232;
	wire n17233;
	wire n17234;
	wire n17235;
	wire n17236;
	wire n17237;
	wire n17238;
	wire n17239;
	wire n17240;
	wire n17241;
	wire n17242;
	wire n17243;
	wire n17244;
	wire n17245;
	wire n17246;
	wire n17247;
	wire n17248;
	wire n17249;
	wire n17250;
	wire n17251;
	wire n17252;
	wire n17253;
	wire n17254;
	wire n17255;
	wire n17256;
	wire n17257;
	wire n17258;
	wire n17259;
	wire n17260;
	wire n17261;
	wire n17262;
	wire n17263;
	wire n17264;
	wire n17265;
	wire n17266;
	wire n17267;
	wire n17268;
	wire n17269;
	wire n17270;
	wire n17271;
	wire n17272;
	wire n17273;
	wire n17274;
	wire n17275;
	wire n17276;
	wire n17277;
	wire n17278;
	wire n17279;
	wire n17280;
	wire n17281;
	wire n17282;
	wire n17283;
	wire n17284;
	wire n17285;
	wire n17286;
	wire n17287;
	wire n17288;
	wire n17289;
	wire n17290;
	wire n17291;
	wire n17292;
	wire n17293;
	wire n17294;
	wire n17295;
	wire n17296;
	wire n17297;
	wire n17298;
	wire n17299;
	wire n17300;
	wire n17301;
	wire n17302;
	wire n17303;
	wire n17304;
	wire n17305;
	wire n17306;
	wire n17307;
	wire n17308;
	wire n17309;
	wire n17310;
	wire n17311;
	wire n17312;
	wire n17313;
	wire n17314;
	wire n17315;
	wire n17316;
	wire n17317;
	wire n17318;
	wire n17319;
	wire n17320;
	wire n17321;
	wire n17322;
	wire n17323;
	wire n17324;
	wire n17325;
	wire n17326;
	wire n17327;
	wire n17328;
	wire n17329;
	wire n17330;
	wire n17331;
	wire n17332;
	wire n17333;
	wire n17334;
	wire n17335;
	wire n17336;
	wire n17337;
	wire n17338;
	wire n17339;
	wire n17340;
	wire n17341;
	wire n17342;
	wire n17343;
	wire n17344;
	wire n17345;
	wire n17346;
	wire n17347;
	wire n17348;
	wire n17349;
	wire n17350;
	wire n17351;
	wire n17352;
	wire n17353;
	wire n17354;
	wire n17355;
	wire n17356;
	wire n17357;
	wire n17358;
	wire n17359;
	wire n17360;
	wire n17361;
	wire n17362;
	wire n17363;
	wire n17364;
	wire n17365;
	wire n17366;
	wire n17367;
	wire n17368;
	wire n17369;
	wire n17370;
	wire n17371;
	wire n17372;
	wire n17373;
	wire n17374;
	wire n17375;
	wire n17376;
	wire n17377;
	wire n17378;
	wire n17379;
	wire n17380;
	wire n17381;
	wire n17382;
	wire n17383;
	wire n17384;
	wire n17385;
	wire n17386;
	wire n17387;
	wire n17388;
	wire n17389;
	wire n17390;
	wire n17391;
	wire n17392;
	wire n17393;
	wire n17394;
	wire n17395;
	wire n17396;
	wire n17397;
	wire n17398;
	wire n17399;
	wire n17400;
	wire n17401;
	wire n17402;
	wire n17403;
	wire n17404;
	wire n17405;
	wire n17406;
	wire n17407;
	wire n17408;
	wire n17409;
	wire n17410;
	wire n17411;
	wire n17412;
	wire n17413;
	wire n17414;
	wire n17415;
	wire n17416;
	wire n17417;
	wire n17418;
	wire n17419;
	wire n17420;
	wire n17421;
	wire n17422;
	wire n17423;
	wire n17424;
	wire n17425;
	wire n17426;
	wire n17427;
	wire n17428;
	wire n17429;
	wire n17430;
	wire n17431;
	wire n17432;
	wire n17433;
	wire n17434;
	wire n17435;
	wire n17436;
	wire n17437;
	wire n17438;
	wire n17439;
	wire n17440;
	wire n17441;
	wire n17442;
	wire n17443;
	wire n17444;
	wire n17445;
	wire n17446;
	wire n17447;
	wire n17448;
	wire n17449;
	wire n17450;
	wire n17451;
	wire n17452;
	wire n17453;
	wire n17454;
	wire n17455;
	wire n17456;
	wire n17457;
	wire n17458;
	wire n17459;
	wire n17460;
	wire n17461;
	wire n17462;
	wire n17463;
	wire n17464;
	wire n17465;
	wire n17466;
	wire n17467;
	wire n17468;
	wire n17469;
	wire n17470;
	wire n17471;
	wire n17472;
	wire n17473;
	wire n17474;
	wire n17475;
	wire n17476;
	wire n17477;
	wire n17478;
	wire n17479;
	wire n17480;
	wire n17481;
	wire n17482;
	wire n17483;
	wire n17484;
	wire n17485;
	wire n17486;
	wire n17487;
	wire n17488;
	wire n17489;
	wire n17490;
	wire n17491;
	wire n17492;
	wire n17493;
	wire n17494;
	wire n17495;
	wire n17496;
	wire n17497;
	wire n17498;
	wire n17499;
	wire n17500;
	wire n17501;
	wire n17502;
	wire n17503;
	wire n17504;
	wire n17505;
	wire n17506;
	wire n17507;
	wire n17508;
	wire n17509;
	wire n17510;
	wire n17511;
	wire n17512;
	wire n17513;
	wire n17514;
	wire n17515;
	wire n17516;
	wire n17517;
	wire n17518;
	wire n17519;
	wire n17520;
	wire n17521;
	wire n17522;
	wire n17523;
	wire n17524;
	wire n17525;
	wire n17526;
	wire n17527;
	wire n17528;
	wire n17529;
	wire n17530;
	wire n17531;
	wire n17532;
	wire n17533;
	wire n17534;
	wire n17535;
	wire n17536;
	wire n17537;
	wire n17538;
	wire n17539;
	wire n17540;
	wire n17541;
	wire n17542;
	wire n17543;
	wire n17544;
	wire n17545;
	wire n17546;
	wire n17547;
	wire n17548;
	wire n17549;
	wire n17550;
	wire n17551;
	wire n17552;
	wire n17553;
	wire n17554;
	wire n17555;
	wire n17556;
	wire n17557;
	wire n17558;
	wire n17559;
	wire n17560;
	wire n17561;
	wire n17562;
	wire n17563;
	wire n17564;
	wire n17565;
	wire n17566;
	wire n17567;
	wire n17568;
	wire n17569;
	wire n17570;
	wire n17571;
	wire n17572;
	wire n17573;
	wire n17574;
	wire n17575;
	wire n17576;
	wire n17577;
	wire n17578;
	wire n17579;
	wire n17580;
	wire n17581;
	wire n17582;
	wire n17583;
	wire n17584;
	wire n17585;
	wire n17586;
	wire n17587;
	wire n17588;
	wire n17589;
	wire n17590;
	wire n17591;
	wire n17592;
	wire n17593;
	wire n17594;
	wire n17595;
	wire n17596;
	wire n17597;
	wire n17598;
	wire n17599;
	wire n17600;
	wire n17601;
	wire n17602;
	wire n17603;
	wire n17604;
	wire n17605;
	wire n17606;
	wire n17607;
	wire n17608;
	wire n17609;
	wire n17610;
	wire n17611;
	wire n17612;
	wire n17613;
	wire n17614;
	wire n17615;
	wire n17616;
	wire n17617;
	wire n17618;
	wire n17619;
	wire n17620;
	wire n17621;
	wire n17622;
	wire n17623;
	wire n17624;
	wire n17625;
	wire n17626;
	wire n17627;
	wire n17628;
	wire n17629;
	wire n17630;
	wire n17631;
	wire n17632;
	wire n17633;
	wire n17634;
	wire n17635;
	wire n17636;
	wire n17637;
	wire n17638;
	wire n17639;
	wire n17640;
	wire n17641;
	wire n17642;
	wire n17643;
	wire n17644;
	wire n17645;
	wire n17646;
	wire n17647;
	wire n17648;
	wire n17649;
	wire n17650;
	wire n17651;
	wire n17652;
	wire n17653;
	wire n17654;
	wire n17655;
	wire n17656;
	wire n17657;
	wire n17658;
	wire n17659;
	wire n17660;
	wire n17661;
	wire n17662;
	wire n17663;
	wire n17664;
	wire n17665;
	wire n17666;
	wire n17667;
	wire n17668;
	wire n17669;
	wire n17670;
	wire n17671;
	wire n17672;
	wire n17673;
	wire n17674;
	wire n17675;
	wire n17676;
	wire n17677;
	wire n17678;
	wire n17679;
	wire n17680;
	wire n17681;
	wire n17682;
	wire n17683;
	wire n17684;
	wire n17685;
	wire n17686;
	wire n17687;
	wire n17688;
	wire n17689;
	wire n17690;
	wire n17691;
	wire n17692;
	wire n17693;
	wire n17694;
	wire n17695;
	wire n17696;
	wire n17697;
	wire n17698;
	wire n17699;
	wire n17700;
	wire n17701;
	wire n17702;
	wire n17703;
	wire n17704;
	wire n17705;
	wire n17706;
	wire n17707;
	wire n17708;
	wire n17709;
	wire n17710;
	wire n17711;
	wire n17712;
	wire n17713;
	wire n17714;
	wire n17715;
	wire n17716;
	wire n17717;
	wire n17718;
	wire n17719;
	wire n17720;
	wire n17721;
	wire n17722;
	wire n17723;
	wire n17724;
	wire n17725;
	wire n17726;
	wire n17727;
	wire n17728;
	wire n17729;
	wire n17730;
	wire n17731;
	wire n17732;
	wire n17733;
	wire n17734;
	wire n17735;
	wire n17736;
	wire n17737;
	wire n17738;
	wire n17739;
	wire n17740;
	wire n17741;
	wire n17742;
	wire n17743;
	wire n17744;
	wire n17745;
	wire n17746;
	wire n17747;
	wire n17748;
	wire n17749;
	wire n17750;
	wire n17751;
	wire n17752;
	wire n17753;
	wire n17754;
	wire n17755;
	wire n17756;
	wire n17757;
	wire n17758;
	wire n17760;
	wire n17761;
	wire n17762;
	wire n17763;
	wire n17764;
	wire n17765;
	wire n17766;
	wire n17767;
	wire n17768;
	wire n17769;
	wire n17770;
	wire n17771;
	wire n17772;
	wire n17773;
	wire n17774;
	wire n17775;
	wire n17776;
	wire n17777;
	wire n17778;
	wire n17779;
	wire n17780;
	wire n17781;
	wire n17782;
	wire n17783;
	wire n17784;
	wire n17785;
	wire n17786;
	wire n17787;
	wire n17788;
	wire n17789;
	wire n17790;
	wire n17791;
	wire n17792;
	wire n17793;
	wire n17794;
	wire n17795;
	wire n17796;
	wire n17797;
	wire n17798;
	wire n17799;
	wire n17800;
	wire n17801;
	wire n17802;
	wire n17803;
	wire n17804;
	wire n17805;
	wire n17806;
	wire n17807;
	wire n17808;
	wire n17809;
	wire n17810;
	wire n17811;
	wire n17812;
	wire n17813;
	wire n17814;
	wire n17815;
	wire n17816;
	wire n17817;
	wire n17818;
	wire n17819;
	wire n17820;
	wire n17821;
	wire n17822;
	wire n17823;
	wire n17824;
	wire n17825;
	wire n17826;
	wire n17827;
	wire n17828;
	wire n17829;
	wire n17830;
	wire n17831;
	wire n17832;
	wire n17833;
	wire n17834;
	wire n17835;
	wire n17836;
	wire n17837;
	wire n17838;
	wire n17839;
	wire n17840;
	wire n17841;
	wire n17842;
	wire n17843;
	wire n17844;
	wire n17845;
	wire n17846;
	wire n17847;
	wire n17848;
	wire n17849;
	wire n17850;
	wire n17851;
	wire n17852;
	wire n17853;
	wire n17854;
	wire n17855;
	wire n17856;
	wire n17857;
	wire n17858;
	wire n17859;
	wire n17860;
	wire n17861;
	wire n17862;
	wire n17863;
	wire n17864;
	wire n17865;
	wire n17866;
	wire n17867;
	wire n17868;
	wire n17869;
	wire n17870;
	wire n17871;
	wire n17872;
	wire n17873;
	wire n17874;
	wire n17875;
	wire n17876;
	wire n17877;
	wire n17878;
	wire n17879;
	wire n17880;
	wire n17881;
	wire n17882;
	wire n17883;
	wire n17884;
	wire n17885;
	wire n17886;
	wire n17887;
	wire n17888;
	wire n17889;
	wire n17890;
	wire n17891;
	wire n17892;
	wire n17893;
	wire n17894;
	wire n17895;
	wire n17896;
	wire n17897;
	wire n17898;
	wire n17899;
	wire n17900;
	wire n17901;
	wire n17902;
	wire n17903;
	wire n17904;
	wire n17905;
	wire n17906;
	wire n17907;
	wire n17908;
	wire n17909;
	wire n17910;
	wire n17911;
	wire n17912;
	wire n17913;
	wire n17914;
	wire n17915;
	wire n17916;
	wire n17917;
	wire n17918;
	wire n17919;
	wire n17920;
	wire n17921;
	wire n17922;
	wire n17923;
	wire n17924;
	wire n17925;
	wire n17926;
	wire n17927;
	wire n17928;
	wire n17929;
	wire n17930;
	wire n17931;
	wire n17932;
	wire n17933;
	wire n17934;
	wire n17935;
	wire n17936;
	wire n17937;
	wire n17938;
	wire n17939;
	wire n17940;
	wire n17941;
	wire n17942;
	wire n17943;
	wire n17944;
	wire n17945;
	wire n17946;
	wire n17947;
	wire n17948;
	wire n17949;
	wire n17950;
	wire n17951;
	wire n17952;
	wire n17953;
	wire n17954;
	wire n17955;
	wire n17956;
	wire n17957;
	wire n17958;
	wire n17959;
	wire n17960;
	wire n17961;
	wire n17962;
	wire n17963;
	wire n17964;
	wire n17965;
	wire n17966;
	wire n17967;
	wire n17968;
	wire n17969;
	wire n17970;
	wire n17971;
	wire n17972;
	wire n17973;
	wire n17974;
	wire n17975;
	wire n17976;
	wire n17977;
	wire n17978;
	wire n17979;
	wire n17980;
	wire n17981;
	wire n17982;
	wire n17983;
	wire n17984;
	wire n17985;
	wire n17986;
	wire n17987;
	wire n17988;
	wire n17989;
	wire n17990;
	wire n17991;
	wire n17992;
	wire n17993;
	wire n17994;
	wire n17995;
	wire n17996;
	wire n17997;
	wire n17998;
	wire n17999;
	wire n18000;
	wire n18001;
	wire n18002;
	wire n18003;
	wire n18004;
	wire n18005;
	wire n18006;
	wire n18007;
	wire n18008;
	wire n18009;
	wire n18010;
	wire n18011;
	wire n18012;
	wire n18013;
	wire n18014;
	wire n18015;
	wire n18016;
	wire n18017;
	wire n18018;
	wire n18019;
	wire n18020;
	wire n18021;
	wire n18022;
	wire n18023;
	wire n18024;
	wire n18025;
	wire n18026;
	wire n18027;
	wire n18028;
	wire n18029;
	wire n18030;
	wire n18031;
	wire n18032;
	wire n18033;
	wire n18034;
	wire n18035;
	wire n18036;
	wire n18037;
	wire n18038;
	wire n18039;
	wire n18040;
	wire n18041;
	wire n18042;
	wire n18043;
	wire n18044;
	wire n18045;
	wire n18046;
	wire n18047;
	wire n18048;
	wire n18049;
	wire n18050;
	wire n18051;
	wire n18052;
	wire n18053;
	wire n18054;
	wire n18055;
	wire n18056;
	wire n18057;
	wire n18058;
	wire n18059;
	wire n18060;
	wire n18061;
	wire n18062;
	wire n18063;
	wire n18064;
	wire n18065;
	wire n18066;
	wire n18067;
	wire n18068;
	wire n18069;
	wire n18070;
	wire n18071;
	wire n18072;
	wire n18073;
	wire n18074;
	wire n18075;
	wire n18076;
	wire n18077;
	wire n18078;
	wire n18079;
	wire n18080;
	wire n18081;
	wire n18082;
	wire n18083;
	wire n18084;
	wire n18085;
	wire n18086;
	wire n18087;
	wire n18088;
	wire n18089;
	wire n18090;
	wire n18091;
	wire n18092;
	wire n18093;
	wire n18094;
	wire n18095;
	wire n18096;
	wire n18097;
	wire n18098;
	wire n18099;
	wire n18100;
	wire n18101;
	wire n18102;
	wire n18103;
	wire n18104;
	wire n18105;
	wire n18106;
	wire n18107;
	wire n18108;
	wire n18109;
	wire n18110;
	wire n18111;
	wire n18112;
	wire n18113;
	wire n18114;
	wire n18115;
	wire n18116;
	wire n18117;
	wire n18118;
	wire n18119;
	wire n18120;
	wire n18121;
	wire n18122;
	wire n18123;
	wire n18124;
	wire n18125;
	wire n18126;
	wire n18127;
	wire n18128;
	wire n18129;
	wire n18130;
	wire n18131;
	wire n18132;
	wire n18133;
	wire n18134;
	wire n18135;
	wire n18136;
	wire n18137;
	wire n18138;
	wire n18139;
	wire n18140;
	wire n18141;
	wire n18142;
	wire n18143;
	wire n18144;
	wire n18145;
	wire n18146;
	wire n18147;
	wire n18148;
	wire n18149;
	wire n18150;
	wire n18151;
	wire n18152;
	wire n18153;
	wire n18154;
	wire n18155;
	wire n18156;
	wire n18157;
	wire n18158;
	wire n18159;
	wire n18160;
	wire n18161;
	wire n18162;
	wire n18163;
	wire n18164;
	wire n18165;
	wire n18166;
	wire n18167;
	wire n18168;
	wire n18169;
	wire n18170;
	wire n18171;
	wire n18172;
	wire n18173;
	wire n18174;
	wire n18175;
	wire n18176;
	wire n18177;
	wire n18178;
	wire n18180;
	wire n18181;
	wire n18182;
	wire n18183;
	wire n18184;
	wire n18185;
	wire n18186;
	wire n18187;
	wire n18188;
	wire n18189;
	wire n18190;
	wire n18191;
	wire n18192;
	wire n18193;
	wire n18194;
	wire n18195;
	wire n18196;
	wire n18197;
	wire n18198;
	wire n18199;
	wire n18200;
	wire n18201;
	wire n18202;
	wire n18203;
	wire n18204;
	wire n18205;
	wire n18206;
	wire n18207;
	wire n18208;
	wire n18209;
	wire n18210;
	wire n18211;
	wire n18212;
	wire n18213;
	wire n18214;
	wire n18215;
	wire n18216;
	wire n18217;
	wire n18218;
	wire n18219;
	wire n18220;
	wire n18221;
	wire n18222;
	wire n18223;
	wire n18224;
	wire n18225;
	wire n18226;
	wire n18227;
	wire n18228;
	wire n18229;
	wire n18230;
	wire n18231;
	wire n18232;
	wire n18233;
	wire n18234;
	wire n18235;
	wire n18236;
	wire n18237;
	wire n18238;
	wire n18239;
	wire n18240;
	wire n18241;
	wire n18242;
	wire n18243;
	wire n18244;
	wire n18245;
	wire n18246;
	wire n18247;
	wire n18248;
	wire n18249;
	wire n18250;
	wire n18251;
	wire n18252;
	wire n18253;
	wire n18254;
	wire n18255;
	wire n18256;
	wire n18257;
	wire n18258;
	wire n18259;
	wire n18260;
	wire n18261;
	wire n18262;
	wire n18263;
	wire n18264;
	wire n18265;
	wire n18266;
	wire n18267;
	wire n18268;
	wire n18269;
	wire n18270;
	wire n18271;
	wire n18272;
	wire n18273;
	wire n18274;
	wire n18275;
	wire n18276;
	wire n18277;
	wire n18278;
	wire n18279;
	wire n18280;
	wire n18281;
	wire n18282;
	wire n18283;
	wire n18284;
	wire n18285;
	wire n18286;
	wire n18287;
	wire n18288;
	wire n18289;
	wire n18290;
	wire n18291;
	wire n18292;
	wire n18293;
	wire n18294;
	wire n18295;
	wire n18296;
	wire n18297;
	wire n18298;
	wire n18299;
	wire n18300;
	wire n18301;
	wire n18302;
	wire n18303;
	wire n18304;
	wire n18305;
	wire n18306;
	wire n18307;
	wire n18308;
	wire n18309;
	wire n18310;
	wire n18311;
	wire n18312;
	wire n18313;
	wire n18314;
	wire n18315;
	wire n18316;
	wire n18317;
	wire n18318;
	wire n18319;
	wire n18320;
	wire n18321;
	wire n18322;
	wire n18323;
	wire n18324;
	wire n18325;
	wire n18326;
	wire n18327;
	wire n18328;
	wire n18329;
	wire n18330;
	wire n18331;
	wire n18332;
	wire n18333;
	wire n18334;
	wire n18335;
	wire n18336;
	wire n18337;
	wire n18338;
	wire n18339;
	wire n18340;
	wire n18341;
	wire n18342;
	wire n18343;
	wire n18344;
	wire n18345;
	wire n18346;
	wire n18347;
	wire n18348;
	wire n18349;
	wire n18350;
	wire n18351;
	wire n18352;
	wire n18353;
	wire n18354;
	wire n18355;
	wire n18356;
	wire n18357;
	wire n18358;
	wire n18359;
	wire n18360;
	wire n18361;
	wire n18362;
	wire n18363;
	wire n18364;
	wire n18365;
	wire n18366;
	wire n18367;
	wire n18368;
	wire n18369;
	wire n18370;
	wire n18371;
	wire n18372;
	wire n18373;
	wire n18374;
	wire n18375;
	wire n18376;
	wire n18377;
	wire n18378;
	wire n18379;
	wire n18380;
	wire n18381;
	wire n18382;
	wire n18383;
	wire n18384;
	wire n18385;
	wire n18386;
	wire n18387;
	wire n18388;
	wire n18389;
	wire n18390;
	wire n18391;
	wire n18392;
	wire n18393;
	wire n18394;
	wire n18395;
	wire n18396;
	wire n18397;
	wire n18398;
	wire n18399;
	wire n18400;
	wire n18401;
	wire n18402;
	wire n18403;
	wire n18404;
	wire n18405;
	wire n18406;
	wire n18407;
	wire n18408;
	wire n18409;
	wire n18410;
	wire n18411;
	wire n18412;
	wire n18413;
	wire n18414;
	wire n18415;
	wire n18416;
	wire n18417;
	wire n18418;
	wire n18419;
	wire n18420;
	wire n18421;
	wire n18422;
	wire n18423;
	wire n18424;
	wire n18425;
	wire n18426;
	wire n18427;
	wire n18428;
	wire n18429;
	wire n18430;
	wire n18431;
	wire n18432;
	wire n18433;
	wire n18434;
	wire n18435;
	wire n18436;
	wire n18437;
	wire n18438;
	wire n18439;
	wire n18440;
	wire n18441;
	wire n18442;
	wire n18443;
	wire n18444;
	wire n18445;
	wire n18446;
	wire n18447;
	wire n18448;
	wire n18449;
	wire n18450;
	wire n18451;
	wire n18452;
	wire n18453;
	wire n18454;
	wire n18455;
	wire n18456;
	wire n18457;
	wire n18458;
	wire n18459;
	wire n18460;
	wire n18461;
	wire n18462;
	wire n18463;
	wire n18464;
	wire n18465;
	wire n18466;
	wire n18467;
	wire n18468;
	wire n18469;
	wire n18470;
	wire n18471;
	wire n18472;
	wire n18473;
	wire n18474;
	wire n18475;
	wire n18476;
	wire n18477;
	wire n18478;
	wire n18479;
	wire n18480;
	wire n18481;
	wire n18482;
	wire n18483;
	wire n18484;
	wire n18485;
	wire n18486;
	wire n18487;
	wire n18488;
	wire n18489;
	wire n18490;
	wire n18491;
	wire n18492;
	wire n18493;
	wire n18494;
	wire n18495;
	wire n18496;
	wire n18497;
	wire n18498;
	wire n18499;
	wire n18500;
	wire n18501;
	wire n18502;
	wire n18503;
	wire n18504;
	wire n18505;
	wire n18506;
	wire n18507;
	wire n18508;
	wire n18509;
	wire n18510;
	wire n18511;
	wire n18512;
	wire n18513;
	wire n18514;
	wire n18515;
	wire n18516;
	wire n18517;
	wire n18518;
	wire n18519;
	wire n18520;
	wire n18521;
	wire n18522;
	wire n18523;
	wire n18524;
	wire n18525;
	wire n18526;
	wire n18527;
	wire n18528;
	wire n18529;
	wire n18530;
	wire n18531;
	wire n18532;
	wire n18533;
	wire n18534;
	wire n18535;
	wire n18536;
	wire n18537;
	wire n18538;
	wire n18539;
	wire n18540;
	wire n18541;
	wire n18542;
	wire n18543;
	wire n18544;
	wire n18545;
	wire n18546;
	wire n18547;
	wire n18548;
	wire n18549;
	wire n18550;
	wire n18551;
	wire n18552;
	wire n18553;
	wire n18554;
	wire n18555;
	wire n18556;
	wire n18557;
	wire n18558;
	wire n18559;
	wire n18560;
	wire n18561;
	wire n18562;
	wire n18563;
	wire n18564;
	wire n18565;
	wire n18566;
	wire n18567;
	wire n18568;
	wire n18569;
	wire n18570;
	wire n18571;
	wire n18572;
	wire n18573;
	wire n18574;
	wire n18575;
	wire n18576;
	wire n18577;
	wire n18578;
	wire n18579;
	wire n18580;
	wire n18581;
	wire n18582;
	wire n18583;
	wire n18584;
	wire n18585;
	wire n18586;
	wire n18587;
	wire n18588;
	wire n18589;
	wire n18590;
	wire n18591;
	wire n18592;
	wire n18593;
	wire n18594;
	wire n18595;
	wire n18596;
	wire n18597;
	wire n18598;
	wire n18599;
	wire n18600;
	wire n18601;
	wire n18602;
	wire n18603;
	wire n18604;
	wire n18605;
	wire n18606;
	wire n18607;
	wire n18608;
	wire n18609;
	wire n18610;
	wire n18611;
	wire n18612;
	wire n18613;
	wire n18614;
	wire n18615;
	wire n18616;
	wire n18617;
	wire n18618;
	wire n18619;
	wire n18620;
	wire n18621;
	wire n18622;
	wire n18623;
	wire n18624;
	wire n18625;
	wire n18626;
	wire n18627;
	wire n18628;
	wire n18629;
	wire n18630;
	wire n18631;
	wire n18632;
	wire n18633;
	wire n18634;
	wire n18635;
	wire n18636;
	wire n18637;
	wire n18638;
	wire n18639;
	wire n18640;
	wire n18641;
	wire n18642;
	wire n18643;
	wire n18644;
	wire n18645;
	wire n18646;
	wire n18647;
	wire n18648;
	wire n18649;
	wire n18650;
	wire n18651;
	wire n18652;
	wire n18653;
	wire n18654;
	wire n18655;
	wire n18656;
	wire n18657;
	wire n18658;
	wire n18659;
	wire n18660;
	wire n18661;
	wire n18662;
	wire n18663;
	wire n18664;
	wire n18665;
	wire n18666;
	wire n18667;
	wire n18668;
	wire n18669;
	wire n18670;
	wire n18671;
	wire n18672;
	wire n18673;
	wire n18674;
	wire n18675;
	wire n18676;
	wire n18677;
	wire n18678;
	wire n18679;
	wire n18680;
	wire n18681;
	wire n18682;
	wire n18683;
	wire n18684;
	wire n18685;
	wire n18686;
	wire n18687;
	wire n18688;
	wire n18689;
	wire n18690;
	wire n18691;
	wire n18692;
	wire n18693;
	wire n18694;
	wire n18695;
	wire n18696;
	wire n18697;
	wire n18698;
	wire n18699;
	wire n18700;
	wire n18701;
	wire n18702;
	wire n18703;
	wire n18704;
	wire n18705;
	wire n18706;
	wire n18707;
	wire n18708;
	wire n18709;
	wire n18710;
	wire n18711;
	wire n18712;
	wire n18713;
	wire n18714;
	wire n18715;
	wire n18716;
	wire n18717;
	wire n18718;
	wire n18719;
	wire n18720;
	wire n18721;
	wire n18722;
	wire n18723;
	wire n18724;
	wire n18725;
	wire n18726;
	wire n18727;
	wire n18728;
	wire n18729;
	wire n18730;
	wire n18731;
	wire n18732;
	wire n18733;
	wire n18734;
	wire n18735;
	wire n18736;
	wire n18737;
	wire n18738;
	wire n18739;
	wire n18740;
	wire n18741;
	wire n18742;
	wire n18743;
	wire n18744;
	wire n18745;
	wire n18746;
	wire n18747;
	wire n18748;
	wire n18749;
	wire n18750;
	wire n18751;
	wire n18752;
	wire n18753;
	wire n18754;
	wire n18755;
	wire n18756;
	wire n18757;
	wire n18758;
	wire n18759;
	wire n18760;
	wire n18761;
	wire n18762;
	wire n18763;
	wire n18764;
	wire n18765;
	wire n18766;
	wire n18767;
	wire n18768;
	wire n18769;
	wire n18770;
	wire n18771;
	wire n18772;
	wire n18773;
	wire n18774;
	wire n18775;
	wire n18776;
	wire n18777;
	wire n18778;
	wire n18779;
	wire n18780;
	wire n18781;
	wire n18782;
	wire n18783;
	wire n18784;
	wire n18785;
	wire n18786;
	wire n18787;
	wire n18788;
	wire n18789;
	wire n18790;
	wire n18791;
	wire n18792;
	wire n18793;
	wire n18794;
	wire n18795;
	wire n18796;
	wire n18797;
	wire n18798;
	wire n18799;
	wire n18800;
	wire n18801;
	wire n18802;
	wire n18803;
	wire n18804;
	wire n18805;
	wire n18806;
	wire n18807;
	wire n18808;
	wire n18809;
	wire n18810;
	wire n18811;
	wire n18812;
	wire n18813;
	wire n18814;
	wire n18815;
	wire n18816;
	wire n18817;
	wire n18818;
	wire n18819;
	wire n18820;
	wire n18821;
	wire n18822;
	wire n18823;
	wire n18824;
	wire n18825;
	wire n18826;
	wire n18827;
	wire n18828;
	wire n18829;
	wire n18830;
	wire n18831;
	wire n18832;
	wire n18833;
	wire n18834;
	wire n18835;
	wire n18836;
	wire n18837;
	wire n18838;
	wire n18839;
	wire n18840;
	wire n18841;
	wire n18842;
	wire n18843;
	wire n18844;
	wire n18845;
	wire n18846;
	wire n18847;
	wire n18848;
	wire n18849;
	wire n18850;
	wire n18851;
	wire n18852;
	wire n18853;
	wire n18854;
	wire n18855;
	wire n18856;
	wire n18857;
	wire n18858;
	wire n18859;
	wire n18860;
	wire n18861;
	wire n18862;
	wire n18863;
	wire n18864;
	wire n18865;
	wire n18866;
	wire n18867;
	wire n18868;
	wire n18869;
	wire n18870;
	wire n18871;
	wire n18872;
	wire n18873;
	wire n18874;
	wire n18875;
	wire n18876;
	wire n18877;
	wire n18878;
	wire n18879;
	wire n18880;
	wire n18881;
	wire n18882;
	wire n18883;
	wire n18884;
	wire n18885;
	wire n18886;
	wire n18887;
	wire n18888;
	wire n18889;
	wire n18890;
	wire n18891;
	wire n18892;
	wire n18893;
	wire n18894;
	wire n18895;
	wire n18896;
	wire n18897;
	wire n18898;
	wire n18899;
	wire n18900;
	wire n18901;
	wire n18902;
	wire n18903;
	wire n18904;
	wire n18905;
	wire n18906;
	wire n18907;
	wire n18908;
	wire n18909;
	wire n18910;
	wire n18911;
	wire n18912;
	wire n18913;
	wire n18914;
	wire n18915;
	wire n18916;
	wire n18917;
	wire n18918;
	wire n18919;
	wire n18920;
	wire n18921;
	wire n18922;
	wire n18923;
	wire n18924;
	wire n18925;
	wire n18926;
	wire n18927;
	wire n18928;
	wire n18929;
	wire n18930;
	wire n18931;
	wire n18932;
	wire n18933;
	wire n18934;
	wire n18935;
	wire n18936;
	wire n18937;
	wire n18938;
	wire n18939;
	wire n18940;
	wire n18941;
	wire n18942;
	wire n18943;
	wire n18944;
	wire n18945;
	wire n18946;
	wire n18947;
	wire n18948;
	wire n18949;
	wire n18950;
	wire n18951;
	wire n18952;
	wire n18953;
	wire n18954;
	wire n18955;
	wire n18956;
	wire n18957;
	wire n18958;
	wire n18959;
	wire n18960;
	wire n18961;
	wire n18962;
	wire n18963;
	wire n18964;
	wire n18965;
	wire n18966;
	wire n18967;
	wire n18968;
	wire n18969;
	wire n18970;
	wire n18971;
	wire n18972;
	wire n18973;
	wire n18974;
	wire n18975;
	wire n18976;
	wire n18977;
	wire n18978;
	wire n18979;
	wire n18980;
	wire n18981;
	wire n18982;
	wire n18983;
	wire n18984;
	wire n18985;
	wire n18986;
	wire n18987;
	wire n18988;
	wire n18989;
	wire n18990;
	wire n18991;
	wire n18992;
	wire n18993;
	wire n18994;
	wire n18995;
	wire n18996;
	wire n18997;
	wire n18998;
	wire n18999;
	wire n19000;
	wire n19001;
	wire n19002;
	wire n19003;
	wire n19004;
	wire n19005;
	wire n19006;
	wire n19007;
	wire n19008;
	wire n19009;
	wire n19010;
	wire n19011;
	wire n19012;
	wire n19013;
	wire n19014;
	wire n19015;
	wire n19016;
	wire n19017;
	wire n19018;
	wire n19019;
	wire n19020;
	wire n19021;
	wire n19022;
	wire n19023;
	wire n19024;
	wire n19025;
	wire n19026;
	wire n19027;
	wire n19028;
	wire n19029;
	wire n19030;
	wire n19031;
	wire n19032;
	wire n19033;
	wire n19034;
	wire n19035;
	wire n19036;
	wire n19037;
	wire n19038;
	wire n19039;
	wire n19040;
	wire n19041;
	wire n19042;
	wire n19043;
	wire n19044;
	wire n19045;
	wire n19046;
	wire n19047;
	wire n19048;
	wire n19049;
	wire n19050;
	wire n19051;
	wire n19052;
	wire n19053;
	wire n19054;
	wire n19055;
	wire n19056;
	wire n19057;
	wire n19058;
	wire n19059;
	wire n19060;
	wire n19061;
	wire n19062;
	wire n19063;
	wire n19064;
	wire n19065;
	wire n19066;
	wire n19067;
	wire n19068;
	wire n19069;
	wire n19070;
	wire n19071;
	wire n19072;
	wire n19073;
	wire n19074;
	wire n19075;
	wire n19076;
	wire n19077;
	wire n19078;
	wire n19079;
	wire n19080;
	wire n19081;
	wire n19083;
	wire n19084;
	wire n19085;
	wire n19086;
	wire n19087;
	wire n19088;
	wire n19089;
	wire n19090;
	wire n19091;
	wire n19092;
	wire n19093;
	wire n19094;
	wire n19095;
	wire n19096;
	wire n19097;
	wire n19098;
	wire n19099;
	wire n19100;
	wire n19101;
	wire n19102;
	wire n19103;
	wire n19104;
	wire n19105;
	wire n19106;
	wire n19107;
	wire n19108;
	wire n19109;
	wire n19110;
	wire n19111;
	wire n19112;
	wire n19113;
	wire n19114;
	wire n19115;
	wire n19116;
	wire n19117;
	wire n19118;
	wire n19119;
	wire n19120;
	wire n19121;
	wire n19122;
	wire n19123;
	wire n19124;
	wire n19125;
	wire n19126;
	wire n19127;
	wire n19128;
	wire n19129;
	wire n19130;
	wire n19131;
	wire n19132;
	wire n19133;
	wire n19134;
	wire n19135;
	wire n19136;
	wire n19137;
	wire n19138;
	wire n19139;
	wire n19140;
	wire n19141;
	wire n19142;
	wire n19143;
	wire n19144;
	wire n19145;
	wire n19146;
	wire n19147;
	wire n19148;
	wire n19149;
	wire n19150;
	wire n19151;
	wire n19152;
	wire n19153;
	wire n19154;
	wire n19155;
	wire n19156;
	wire n19157;
	wire n19158;
	wire n19159;
	wire n19160;
	wire n19161;
	wire n19162;
	wire n19163;
	wire n19164;
	wire n19165;
	wire n19166;
	wire n19167;
	wire n19168;
	wire n19169;
	wire n19170;
	wire n19171;
	wire n19172;
	wire n19173;
	wire n19174;
	wire n19175;
	wire n19176;
	wire n19177;
	wire n19178;
	wire n19179;
	wire n19180;
	wire n19181;
	wire n19182;
	wire n19183;
	wire n19184;
	wire n19185;
	wire n19186;
	wire n19187;
	wire n19188;
	wire n19189;
	wire n19190;
	wire n19191;
	wire n19192;
	wire n19193;
	wire n19194;
	wire n19195;
	wire n19196;
	wire n19197;
	wire n19198;
	wire n19199;
	wire n19200;
	wire n19201;
	wire n19202;
	wire n19203;
	wire n19204;
	wire n19205;
	wire n19206;
	wire n19207;
	wire n19208;
	wire n19209;
	wire n19210;
	wire n19211;
	wire n19212;
	wire n19213;
	wire n19214;
	wire n19215;
	wire n19216;
	wire n19217;
	wire n19218;
	wire n19219;
	wire n19220;
	wire n19221;
	wire n19222;
	wire n19223;
	wire n19224;
	wire n19225;
	wire n19226;
	wire n19227;
	wire n19228;
	wire n19229;
	wire n19230;
	wire n19231;
	wire n19232;
	wire n19233;
	wire n19234;
	wire n19235;
	wire n19236;
	wire n19237;
	wire n19238;
	wire n19239;
	wire n19240;
	wire n19241;
	wire n19242;
	wire n19243;
	wire n19244;
	wire n19245;
	wire n19246;
	wire n19247;
	wire n19248;
	wire n19249;
	wire n19250;
	wire n19251;
	wire n19252;
	wire n19253;
	wire n19254;
	wire n19255;
	wire n19256;
	wire n19257;
	wire n19258;
	wire n19259;
	wire n19260;
	wire n19261;
	wire n19262;
	wire n19263;
	wire n19264;
	wire n19265;
	wire n19266;
	wire n19267;
	wire n19268;
	wire n19269;
	wire n19270;
	wire n19271;
	wire n19272;
	wire n19273;
	wire n19274;
	wire n19275;
	wire n19276;
	wire n19277;
	wire n19278;
	wire n19279;
	wire n19280;
	wire n19281;
	wire n19282;
	wire n19283;
	wire n19284;
	wire n19285;
	wire n19286;
	wire n19287;
	wire n19288;
	wire n19289;
	wire n19290;
	wire n19291;
	wire n19292;
	wire n19293;
	wire n19294;
	wire n19295;
	wire n19296;
	wire n19297;
	wire n19298;
	wire n19299;
	wire n19300;
	wire n19301;
	wire n19302;
	wire n19303;
	wire n19304;
	wire n19305;
	wire n19306;
	wire n19307;
	wire n19308;
	wire n19309;
	wire n19310;
	wire n19311;
	wire n19312;
	wire n19313;
	wire n19314;
	wire n19315;
	wire n19316;
	wire n19317;
	wire n19318;
	wire n19319;
	wire n19320;
	wire n19321;
	wire n19322;
	wire n19323;
	wire n19324;
	wire n19325;
	wire n19326;
	wire n19327;
	wire n19328;
	wire n19329;
	wire n19330;
	wire n19331;
	wire n19332;
	wire n19333;
	wire n19334;
	wire n19335;
	wire n19336;
	wire n19337;
	wire n19338;
	wire n19339;
	wire n19340;
	wire n19341;
	wire n19342;
	wire n19343;
	wire n19344;
	wire n19345;
	wire n19346;
	wire n19347;
	wire n19348;
	wire n19349;
	wire n19350;
	wire n19351;
	wire n19352;
	wire n19353;
	wire n19354;
	wire n19355;
	wire n19356;
	wire n19357;
	wire n19358;
	wire n19359;
	wire n19360;
	wire n19361;
	wire n19362;
	wire n19363;
	wire n19364;
	wire n19365;
	wire n19366;
	wire n19367;
	wire n19368;
	wire n19369;
	wire n19370;
	wire n19371;
	wire n19372;
	wire n19373;
	wire n19374;
	wire n19375;
	wire n19376;
	wire n19377;
	wire n19378;
	wire n19379;
	wire n19380;
	wire n19381;
	wire n19382;
	wire n19383;
	wire n19384;
	wire n19385;
	wire n19386;
	wire n19387;
	wire n19388;
	wire n19389;
	wire n19390;
	wire n19391;
	wire n19392;
	wire n19393;
	wire n19394;
	wire n19395;
	wire n19396;
	wire n19397;
	wire n19398;
	wire n19399;
	wire n19400;
	wire n19401;
	wire n19402;
	wire n19403;
	wire n19404;
	wire n19405;
	wire n19406;
	wire n19407;
	wire n19408;
	wire n19409;
	wire n19410;
	wire n19411;
	wire n19412;
	wire n19413;
	wire n19414;
	wire n19415;
	wire n19416;
	wire n19417;
	wire n19418;
	wire n19419;
	wire n19420;
	wire n19421;
	wire n19422;
	wire n19423;
	wire n19424;
	wire n19425;
	wire n19426;
	wire n19427;
	wire n19428;
	wire n19429;
	wire n19430;
	wire n19431;
	wire n19432;
	wire n19433;
	wire n19434;
	wire n19435;
	wire n19436;
	wire n19437;
	wire n19438;
	wire n19439;
	wire n19440;
	wire n19441;
	wire n19442;
	wire n19443;
	wire n19444;
	wire n19445;
	wire n19446;
	wire n19447;
	wire n19448;
	wire n19449;
	wire n19450;
	wire n19451;
	wire n19452;
	wire n19453;
	wire n19454;
	wire n19455;
	wire n19456;
	wire n19457;
	wire n19458;
	wire n19459;
	wire n19460;
	wire n19461;
	wire n19462;
	wire n19463;
	wire n19464;
	wire n19465;
	wire n19466;
	wire n19467;
	wire n19468;
	wire n19469;
	wire n19470;
	wire n19471;
	wire n19472;
	wire n19473;
	wire n19474;
	wire n19475;
	wire n19476;
	wire n19477;
	wire n19478;
	wire n19479;
	wire n19480;
	wire n19481;
	wire n19482;
	wire n19483;
	wire n19484;
	wire n19485;
	wire n19486;
	wire n19487;
	wire n19488;
	wire n19489;
	wire n19490;
	wire n19491;
	wire n19492;
	wire n19493;
	wire n19494;
	wire n19495;
	wire n19496;
	wire n19497;
	wire n19498;
	wire n19499;
	wire n19500;
	wire n19501;
	wire n19502;
	wire n19503;
	wire n19504;
	wire n19505;
	wire n19506;
	wire n19507;
	wire n19508;
	wire n19509;
	wire n19510;
	wire n19511;
	wire n19512;
	wire n19513;
	wire n19514;
	wire n19515;
	wire n19516;
	wire n19520;
	wire n19521;
	wire n19522;
	wire n19523;
	wire n19524;
	wire n19525;
	wire n19526;
	wire n19527;
	wire n19528;
	wire n19529;
	wire n19530;
	wire n19531;
	wire n19532;
	wire n19533;
	wire n19534;
	wire n19535;
	wire n19536;
	wire n19537;
	wire n19538;
	wire n19539;
	wire n19540;
	wire n19541;
	wire n19542;
	wire n19543;
	wire n19544;
	wire n19545;
	wire n19546;
	wire n19547;
	wire n19548;
	wire n19549;
	wire n19550;
	wire n19551;
	wire n19552;
	wire n19553;
	wire n19554;
	wire n19555;
	wire n19556;
	wire n19557;
	wire n19558;
	wire n19559;
	wire n19560;
	wire n19561;
	wire n19562;
	wire n19563;
	wire n19564;
	wire n19565;
	wire n19566;
	wire n19567;
	wire n19568;
	wire n19569;
	wire n19570;
	wire n19571;
	wire n19572;
	wire n19573;
	wire n19574;
	wire n19575;
	wire n19576;
	wire n19577;
	wire n19578;
	wire n19579;
	wire n19580;
	wire n19581;
	wire n19582;
	wire n19583;
	wire n19584;
	wire n19585;
	wire n19586;
	wire n19587;
	wire n19588;
	wire n19589;
	wire n19590;
	wire n19591;
	wire n19592;
	wire n19593;
	wire n19594;
	wire n19595;
	wire n19596;
	wire n19597;
	wire n19598;
	wire n19599;
	wire n19600;
	wire n19601;
	wire n19602;
	wire n19603;
	wire n19604;
	wire n19605;
	wire n19606;
	wire n19607;
	wire n19608;
	wire n19609;
	wire n19610;
	wire n19611;
	wire n19612;
	wire n19613;
	wire n19614;
	wire n19615;
	wire n19616;
	wire n19617;
	wire n19618;
	wire n19619;
	wire n19620;
	wire n19621;
	wire n19622;
	wire n19623;
	wire n19624;
	wire n19625;
	wire n19626;
	wire n19627;
	wire n19628;
	wire n19629;
	wire n19630;
	wire n19631;
	wire n19632;
	wire n19633;
	wire n19634;
	wire n19635;
	wire n19636;
	wire n19637;
	wire n19638;
	wire n19639;
	wire n19640;
	wire n19641;
	wire n19642;
	wire n19643;
	wire n19644;
	wire n19645;
	wire n19646;
	wire n19647;
	wire n19648;
	wire n19649;
	wire n19650;
	wire n19651;
	wire n19652;
	wire n19653;
	wire n19654;
	wire n19655;
	wire n19656;
	wire n19657;
	wire n19658;
	wire n19659;
	wire n19660;
	wire n19661;
	wire n19662;
	wire n19663;
	wire n19664;
	wire n19665;
	wire n19666;
	wire n19667;
	wire n19668;
	wire n19669;
	wire n19670;
	wire n19671;
	wire n19672;
	wire n19673;
	wire n19674;
	wire n19675;
	wire n19676;
	wire n19677;
	wire n19678;
	wire n19679;
	wire n19680;
	wire n19681;
	wire n19682;
	wire n19683;
	wire n19684;
	wire n19685;
	wire n19686;
	wire n19687;
	wire n19688;
	wire n19689;
	wire n19690;
	wire n19691;
	wire n19692;
	wire n19693;
	wire n19694;
	wire n19695;
	wire n19696;
	wire n19697;
	wire n19698;
	wire n19699;
	wire n19700;
	wire n19701;
	wire n19702;
	wire n19703;
	wire n19704;
	wire n19705;
	wire n19706;
	wire n19707;
	wire n19708;
	wire n19709;
	wire n19710;
	wire n19711;
	wire n19712;
	wire n19713;
	wire n19714;
	wire n19715;
	wire n19716;
	wire n19717;
	wire n19718;
	wire n19719;
	wire n19720;
	wire n19721;
	wire n19722;
	wire n19723;
	wire n19724;
	wire n19725;
	wire n19726;
	wire n19727;
	wire n19728;
	wire n19729;
	wire n19730;
	wire n19731;
	wire n19732;
	wire n19733;
	wire n19734;
	wire n19735;
	wire n19736;
	wire n19737;
	wire n19738;
	wire n19739;
	wire n19740;
	wire n19741;
	wire n19742;
	wire n19743;
	wire n19744;
	wire n19745;
	wire n19746;
	wire n19747;
	wire n19748;
	wire n19749;
	wire n19750;
	wire n19751;
	wire n19752;
	wire n19753;
	wire n19754;
	wire n19755;
	wire n19756;
	wire n19757;
	wire n19758;
	wire n19759;
	wire n19760;
	wire n19761;
	wire n19762;
	wire n19763;
	wire n19764;
	wire n19765;
	wire n19766;
	wire n19767;
	wire n19768;
	wire n19769;
	wire n19770;
	wire n19771;
	wire n19772;
	wire n19773;
	wire n19774;
	wire n19775;
	wire n19776;
	wire n19777;
	wire n19778;
	wire n19779;
	wire n19780;
	wire n19781;
	wire n19782;
	wire n19783;
	wire n19784;
	wire n19785;
	wire n19786;
	wire n19787;
	wire n19788;
	wire n19791;
	wire n19792;
	wire n19793;
	wire n19794;
	wire n19795;
	wire n19796;
	wire n19797;
	wire n19798;
	wire n19799;
	wire n19800;
	wire n19801;
	wire n19802;
	wire n19803;
	wire n19804;
	wire n19805;
	wire n19806;
	wire n19807;
	wire n19808;
	wire n19809;
	wire n19810;
	wire n19811;
	wire n19812;
	wire n19813;
	wire n19814;
	wire n19815;
	wire n19816;
	wire n19817;
	wire n19818;
	wire n19819;
	wire n19820;
	wire n19821;
	wire n19822;
	wire n19823;
	wire n19824;
	wire n19825;
	wire n19826;
	wire n19827;
	wire n19828;
	wire n19829;
	wire n19830;
	wire n19831;
	wire n19832;
	wire n19833;
	wire n19834;
	wire n19835;
	wire n19836;
	wire n19837;
	wire n19838;
	wire n19839;
	wire n19840;
	wire n19841;
	wire n19842;
	wire n19843;
	wire n19844;
	wire n19845;
	wire n19846;
	wire n19847;
	wire n19848;
	wire n19849;
	wire n19850;
	wire n19851;
	wire n19852;
	wire n19853;
	wire n19854;
	wire n19855;
	wire n19856;
	wire n19857;
	wire n19858;
	wire n19859;
	wire n19860;
	wire n19861;
	wire n19862;
	wire n19863;
	wire n19864;
	wire n19865;
	wire n19866;
	wire n19867;
	wire n19868;
	wire n19869;
	wire n19870;
	wire n19871;
	wire n19872;
	wire n19873;
	wire n19874;
	wire n19875;
	wire n19876;
	wire n19877;
	wire n19878;
	wire n19879;
	wire n19880;
	wire n19881;
	wire n19882;
	wire n19883;
	wire n19884;
	wire n19885;
	wire n19886;
	wire n19887;
	wire n19888;
	wire n19889;
	wire n19890;
	wire n19891;
	wire n19892;
	wire n19893;
	wire n19894;
	wire n19895;
	wire n19896;
	wire n19897;
	wire n19898;
	wire n19899;
	wire n19900;
	wire n19901;
	wire n19902;
	wire n19903;
	wire n19904;
	wire n19905;
	wire n19906;
	wire n19907;
	wire n19908;
	wire n19909;
	wire n19910;
	wire n19911;
	wire n19912;
	wire n19913;
	wire n19914;
	wire n19915;
	wire n19916;
	wire n19917;
	wire n19918;
	wire n19919;
	wire n19920;
	wire n19921;
	wire n19922;
	wire n19923;
	wire n19924;
	wire n19925;
	wire n19926;
	wire n19927;
	wire n19928;
	wire n19929;
	wire n19930;
	wire n19931;
	wire n19932;
	wire n19933;
	wire n19934;
	wire n19935;
	wire n19936;
	wire n19937;
	wire n19938;
	wire n19939;
	wire n19940;
	wire n19941;
	wire n19942;
	wire n19943;
	wire n19944;
	wire n19945;
	wire n19946;
	wire n19947;
	wire n19948;
	wire n19949;
	wire n19950;
	wire n19951;
	wire n19952;
	wire n19953;
	wire n19954;
	wire n19955;
	wire n19956;
	wire n19957;
	wire n19958;
	wire n19959;
	wire n19960;
	wire n19961;
	wire n19962;
	wire n19963;
	wire n19964;
	wire n19965;
	wire n19966;
	wire n19967;
	wire n19968;
	wire n19969;
	wire n19970;
	wire n19971;
	wire n19972;
	wire n19973;
	wire n19974;
	wire n19975;
	wire n19976;
	wire n19977;
	wire n19978;
	wire n19979;
	wire n19980;
	wire n19981;
	wire n19982;
	wire n19983;
	wire n19984;
	wire n19985;
	wire n19986;
	wire n19987;
	wire n19988;
	wire n19989;
	wire n19990;
	wire n19991;
	wire n19992;
	wire n19993;
	wire n19994;
	wire n19995;
	wire n19996;
	wire n19997;
	wire n19998;
	wire n19999;
	wire n20000;
	wire n20001;
	wire n20002;
	wire n20003;
	wire n20004;
	wire n20005;
	wire n20006;
	wire n20007;
	wire n20008;
	wire n20009;
	wire n20010;
	wire n20011;
	wire n20012;
	wire n20013;
	wire n20014;
	wire n20015;
	wire n20016;
	wire n20017;
	wire n20018;
	wire n20019;
	wire n20020;
	wire n20021;
	wire n20022;
	wire n20023;
	wire n20024;
	wire n20025;
	wire n20026;
	wire n20027;
	wire n20028;
	wire n20029;
	wire n20030;
	wire n20031;
	wire n20032;
	wire n20033;
	wire n20034;
	wire n20035;
	wire n20036;
	wire n20037;
	wire n20038;
	wire n20039;
	wire n20040;
	wire n20041;
	wire n20042;
	wire n20043;
	wire n20044;
	wire n20045;
	wire n20046;
	wire n20047;
	wire n20048;
	wire n20049;
	wire n20050;
	wire n20051;
	wire n20052;
	wire n20053;
	wire n20054;
	wire n20055;
	wire n20056;
	wire n20057;
	wire n20058;
	wire n20059;
	wire n20060;
	wire n20061;
	wire n20062;
	wire n20063;
	wire n20064;
	wire n20065;
	wire n20066;
	wire n20067;
	wire n20068;
	wire n20069;
	wire n20070;
	wire n20071;
	wire n20072;
	wire n20073;
	wire n20074;
	wire n20075;
	wire n20076;
	wire n20077;
	wire n20078;
	wire n20079;
	wire n20080;
	wire n20081;
	wire n20082;
	wire n20083;
	wire n20084;
	wire n20085;
	wire n20086;
	wire n20087;
	wire n20088;
	wire n20089;
	wire n20090;
	wire n20091;
	wire n20092;
	wire n20093;
	wire n20094;
	wire n20095;
	wire n20096;
	wire n20097;
	wire n20098;
	wire n20099;
	wire n20100;
	wire n20101;
	wire n20102;
	wire n20103;
	wire n20104;
	wire n20105;
	wire n20106;
	wire n20107;
	wire n20108;
	wire n20109;
	wire n20110;
	wire n20111;
	wire n20112;
	wire n20113;
	wire n20114;
	wire n20115;
	wire n20116;
	wire n20117;
	wire n20118;
	wire n20119;
	wire n20120;
	wire n20121;
	wire n20122;
	wire n20123;
	wire n20124;
	wire n20125;
	wire n20126;
	wire n20127;
	wire n20128;
	wire n20129;
	wire n20130;
	wire n20131;
	wire n20132;
	wire n20133;
	wire n20134;
	wire n20135;
	wire n20136;
	wire n20137;
	wire n20138;
	wire n20139;
	wire n20140;
	wire n20141;
	wire n20142;
	wire n20143;
	wire n20144;
	wire n20145;
	wire n20146;
	wire n20147;
	wire n20148;
	wire n20149;
	wire n20150;
	wire n20151;
	wire n20152;
	wire n20153;
	wire n20154;
	wire n20155;
	wire n20156;
	wire n20157;
	wire n20158;
	wire n20159;
	wire n20160;
	wire n20161;
	wire n20162;
	wire n20163;
	wire n20164;
	wire n20165;
	wire n20166;
	wire n20167;
	wire n20168;
	wire n20169;
	wire n20170;
	wire n20171;
	wire n20172;
	wire n20173;
	wire n20174;
	wire n20175;
	wire n20176;
	wire n20177;
	wire n20178;
	wire n20179;
	wire n20180;
	wire n20181;
	wire n20182;
	wire n20183;
	wire n20184;
	wire n20185;
	wire n20186;
	wire n20187;
	wire n20188;
	wire n20189;
	wire n20190;
	wire n20191;
	wire n20192;
	wire n20193;
	wire n20194;
	wire n20195;
	wire n20196;
	wire n20197;
	wire n20198;
	wire n20199;
	wire n20200;
	wire n20201;
	wire n20202;
	wire n20203;
	wire n20204;
	wire n20205;
	wire n20206;
	wire n20207;
	wire n20208;
	wire n20209;
	wire n20210;
	wire n20211;
	wire n20212;
	wire n20213;
	wire n20214;
	wire n20215;
	wire n20216;
	wire n20217;
	wire n20218;
	wire n20219;
	wire n20220;
	wire n20221;
	wire n20222;
	wire n20223;
	wire n20224;
	wire n20225;
	wire n20226;
	wire n20227;
	wire n20228;
	wire n20229;
	wire n20230;
	wire n20231;
	wire n20232;
	wire n20233;
	wire n20234;
	wire n20235;
	wire n20236;
	wire n20237;
	wire n20238;
	wire n20239;
	wire n20240;
	wire n20241;
	wire n20242;
	wire n20243;
	wire n20244;
	wire n20245;
	wire n20246;
	wire n20247;
	wire n20248;
	wire n20249;
	wire n20250;
	wire n20251;
	wire n20252;
	wire n20253;
	wire n20254;
	wire n20255;
	wire n20256;
	wire n20257;
	wire n20258;
	wire n20259;
	wire n20260;
	wire n20261;
	wire n20262;
	wire n20263;
	wire n20264;
	wire n20265;
	wire n20266;
	wire n20267;
	wire n20268;
	wire n20269;
	wire n20270;
	wire n20271;
	wire n20272;
	wire n20273;
	wire n20274;
	wire n20275;
	wire n20276;
	wire n20277;
	wire n20278;
	wire n20279;
	wire n20280;
	wire n20281;
	wire n20282;
	wire n20283;
	wire n20284;
	wire n20285;
	wire n20286;
	wire n20287;
	wire n20288;
	wire n20289;
	wire n20290;
	wire n20291;
	wire n20292;
	wire n20293;
	wire n20294;
	wire n20295;
	wire n20296;
	wire n20297;
	wire n20298;
	wire n20299;
	wire n20300;
	wire n20301;
	wire n20302;
	wire n20303;
	wire n20304;
	wire n20305;
	wire n20306;
	wire n20307;
	wire n20308;
	wire n20309;
	wire n20310;
	wire n20311;
	wire n20312;
	wire n20313;
	wire n20314;
	wire n20315;
	wire n20316;
	wire n20317;
	wire n20318;
	wire n20319;
	wire n20320;
	wire n20321;
	wire n20322;
	wire n20323;
	wire n20324;
	wire n20325;
	wire n20326;
	wire n20327;
	wire n20328;
	wire n20329;
	wire n20330;
	wire n20331;
	wire n20332;
	wire n20333;
	wire n20334;
	wire n20335;
	wire n20336;
	wire n20337;
	wire n20338;
	wire n20339;
	wire n20340;
	wire n20341;
	wire n20342;
	wire n20343;
	wire n20344;
	wire n20345;
	wire n20346;
	wire n20347;
	wire n20348;
	wire n20349;
	wire n20350;
	wire n20351;
	wire n20352;
	wire n20353;
	wire n20354;
	wire n20355;
	wire n20356;
	wire n20357;
	wire n20358;
	wire n20359;
	wire n20360;
	wire n20361;
	wire n20362;
	wire n20363;
	wire n20364;
	wire n20365;
	wire n20366;
	wire n20367;
	wire n20368;
	wire n20369;
	wire n20370;
	wire n20371;
	wire n20372;
	wire n20373;
	wire n20374;
	wire n20375;
	wire n20376;
	wire n20377;
	wire n20378;
	wire n20379;
	wire n20380;
	wire n20381;
	wire n20382;
	wire n20383;
	wire n20384;
	wire n20385;
	wire n20386;
	wire n20387;
	wire n20388;
	wire n20389;
	wire n20390;
	wire n20391;
	wire n20392;
	wire n20393;
	wire n20394;
	wire n20395;
	wire n20396;
	wire n20397;
	wire n20398;
	wire n20399;
	wire n20400;
	wire n20401;
	wire n20402;
	wire n20403;
	wire n20404;
	wire n20405;
	wire n20406;
	wire n20407;
	wire n20408;
	wire n20409;
	wire n20410;
	wire n20411;
	wire n20412;
	wire n20413;
	wire n20414;
	wire n20415;
	wire n20416;
	wire n20417;
	wire n20418;
	wire n20419;
	wire n20420;
	wire n20421;
	wire n20422;
	wire n20423;
	wire n20424;
	wire n20425;
	wire n20426;
	wire n20427;
	wire n20428;
	wire n20429;
	wire n20430;
	wire n20431;
	wire n20432;
	wire n20433;
	wire n20434;
	wire n20435;
	wire n20436;
	wire n20437;
	wire n20438;
	wire n20439;
	wire n20440;
	wire n20441;
	wire n20442;
	wire n20443;
	wire n20444;
	wire n20445;
	wire n20446;
	wire n20447;
	wire n20448;
	wire n20449;
	wire n20450;
	wire n20451;
	wire n20452;
	wire n20453;
	wire n20455;
	wire n20456;
	wire n20457;
	wire n20458;
	wire n20459;
	wire n20460;
	wire n20461;
	wire n20462;
	wire n20463;
	wire n20464;
	wire n20465;
	wire n20466;
	wire n20467;
	wire n20468;
	wire n20469;
	wire n20470;
	wire n20471;
	wire n20472;
	wire n20473;
	wire n20474;
	wire n20475;
	wire n20476;
	wire n20477;
	wire n20478;
	wire n20479;
	wire n20480;
	wire n20481;
	wire n20482;
	wire n20483;
	wire n20484;
	wire n20485;
	wire n20486;
	wire n20487;
	wire n20488;
	wire n20489;
	wire n20490;
	wire n20491;
	wire n20492;
	wire n20493;
	wire n20494;
	wire n20495;
	wire n20496;
	wire n20497;
	wire n20498;
	wire n20499;
	wire n20500;
	wire n20501;
	wire n20502;
	wire n20503;
	wire n20504;
	wire n20505;
	wire n20506;
	wire n20507;
	wire n20508;
	wire n20509;
	wire n20510;
	wire n20511;
	wire n20512;
	wire n20513;
	wire n20514;
	wire n20515;
	wire n20516;
	wire n20517;
	wire n20518;
	wire n20519;
	wire n20520;
	wire n20521;
	wire n20522;
	wire n20523;
	wire n20524;
	wire n20525;
	wire n20526;
	wire n20527;
	wire n20528;
	wire n20529;
	wire n20530;
	wire n20531;
	wire n20532;
	wire n20533;
	wire n20534;
	wire n20535;
	wire n20536;
	wire n20537;
	wire n20538;
	wire n20539;
	wire n20540;
	wire n20541;
	wire n20542;
	wire n20543;
	wire n20544;
	wire n20545;
	wire n20546;
	wire n20547;
	wire n20548;
	wire n20549;
	wire n20550;
	wire n20551;
	wire n20552;
	wire n20553;
	wire n20554;
	wire n20555;
	wire n20556;
	wire n20557;
	wire n20558;
	wire n20559;
	wire n20560;
	wire n20561;
	wire n20562;
	wire n20563;
	wire n20564;
	wire n20565;
	wire n20566;
	wire n20567;
	wire n20568;
	wire n20569;
	wire n20570;
	wire n20571;
	wire n20572;
	wire n20573;
	wire n20574;
	wire n20575;
	wire n20576;
	wire n20577;
	wire n20578;
	wire n20579;
	wire n20580;
	wire n20581;
	wire n20582;
	wire n20583;
	wire n20584;
	wire n20585;
	wire n20586;
	wire n20587;
	wire n20588;
	wire n20589;
	wire n20590;
	wire n20591;
	wire n20592;
	wire n20593;
	wire n20594;
	wire n20595;
	wire n20596;
	wire n20597;
	wire n20598;
	wire n20599;
	wire n20600;
	wire n20601;
	wire n20602;
	wire n20603;
	wire n20604;
	wire n20605;
	wire n20606;
	wire n20607;
	wire n20608;
	wire n20609;
	wire n20610;
	wire n20611;
	wire n20612;
	wire n20613;
	wire n20614;
	wire n20615;
	wire n20616;
	wire n20617;
	wire n20618;
	wire n20619;
	wire n20620;
	wire n20621;
	wire n20622;
	wire n20623;
	wire n20624;
	wire n20625;
	wire n20626;
	wire n20627;
	wire n20628;
	wire n20629;
	wire n20630;
	wire n20631;
	wire n20632;
	wire n20633;
	wire n20634;
	wire n20635;
	wire n20636;
	wire n20637;
	wire n20638;
	wire n20639;
	wire n20640;
	wire n20641;
	wire n20642;
	wire n20643;
	wire n20644;
	wire n20645;
	wire n20646;
	wire n20647;
	wire n20648;
	wire n20649;
	wire n20650;
	wire n20651;
	wire n20652;
	wire n20653;
	wire n20654;
	wire n20655;
	wire n20656;
	wire n20657;
	wire n20658;
	wire n20659;
	wire n20660;
	wire n20661;
	wire n20662;
	wire n20663;
	wire n20664;
	wire n20665;
	wire n20666;
	wire n20667;
	wire n20668;
	wire n20669;
	wire n20670;
	wire n20671;
	wire n20672;
	wire n20673;
	wire n20674;
	wire n20675;
	wire n20676;
	wire n20677;
	wire n20678;
	wire n20679;
	wire n20680;
	wire n20681;
	wire n20682;
	wire n20683;
	wire n20684;
	wire n20685;
	wire n20686;
	wire n20687;
	wire n20688;
	wire n20689;
	wire n20690;
	wire n20691;
	wire n20692;
	wire n20693;
	wire n20694;
	wire n20695;
	wire n20696;
	wire n20697;
	wire n20698;
	wire n20699;
	wire n20700;
	wire n20701;
	wire n20702;
	wire n20703;
	wire n20704;
	wire n20705;
	wire n20706;
	wire n20707;
	wire n20708;
	wire n20709;
	wire n20710;
	wire n20711;
	wire n20712;
	wire n20713;
	wire n20714;
	wire n20715;
	wire n20716;
	wire n20717;
	wire n20718;
	wire n20719;
	wire n20720;
	wire n20721;
	wire n20722;
	wire n20723;
	wire n20724;
	wire n20725;
	wire n20726;
	wire n20727;
	wire n20728;
	wire n20729;
	wire n20730;
	wire n20731;
	wire n20732;
	wire n20733;
	wire n20734;
	wire n20735;
	wire n20736;
	wire n20737;
	wire n20738;
	wire n20739;
	wire n20740;
	wire n20741;
	wire n20742;
	wire n20743;
	wire n20744;
	wire n20745;
	wire n20746;
	wire n20747;
	wire n20748;
	wire n20749;
	wire n20750;
	wire n20751;
	wire n20752;
	wire n20753;
	wire n20754;
	wire n20755;
	wire n20756;
	wire n20757;
	wire n20758;
	wire n20759;
	wire n20760;
	wire n20761;
	wire n20762;
	wire n20763;
	wire n20764;
	wire n20765;
	wire n20766;
	wire n20767;
	wire n20768;
	wire n20769;
	wire n20770;
	wire n20771;
	wire n20772;
	wire n20773;
	wire n20774;
	wire n20775;
	wire n20776;
	wire n20777;
	wire n20778;
	wire n20779;
	wire n20780;
	wire n20781;
	wire n20782;
	wire n20783;
	wire n20784;
	wire n20785;
	wire n20786;
	wire n20787;
	wire n20788;
	wire n20789;
	wire n20790;
	wire n20791;
	wire n20792;
	wire n20793;
	wire n20794;
	wire n20795;
	wire n20796;
	wire n20797;
	wire n20798;
	wire n20799;
	wire n20800;
	wire n20801;
	wire n20802;
	wire n20803;
	wire n20804;
	wire n20805;
	wire n20806;
	wire n20807;
	wire n20808;
	wire n20809;
	wire n20810;
	wire n20811;
	wire n20812;
	wire n20813;
	wire n20814;
	wire n20815;
	wire n20816;
	wire n20817;
	wire n20818;
	wire n20819;
	wire n20820;
	wire n20821;
	wire n20822;
	wire n20823;
	wire n20824;
	wire n20825;
	wire n20826;
	wire n20827;
	wire n20828;
	wire n20829;
	wire n20830;
	wire n20831;
	wire n20832;
	wire n20833;
	wire n20834;
	wire n20835;
	wire n20836;
	wire n20837;
	wire n20838;
	wire n20839;
	wire n20840;
	wire n20841;
	wire n20842;
	wire n20843;
	wire n20844;
	wire n20845;
	wire n20846;
	wire n20847;
	wire n20848;
	wire n20849;
	wire n20850;
	wire n20851;
	wire n20852;
	wire n20853;
	wire n20854;
	wire n20855;
	wire n20856;
	wire n20857;
	wire n20858;
	wire n20859;
	wire n20860;
	wire n20861;
	wire n20862;
	wire n20863;
	wire n20864;
	wire n20865;
	wire n20866;
	wire n20867;
	wire n20868;
	wire n20869;
	wire n20870;
	wire n20871;
	wire n20872;
	wire n20873;
	wire n20874;
	wire n20875;
	wire n20876;
	wire n20877;
	wire n20878;
	wire n20879;
	wire n20880;
	wire n20881;
	wire n20882;
	wire n20883;
	wire n20884;
	wire n20885;
	wire n20886;
	wire n20887;
	wire n20888;
	wire n20889;
	wire n20890;
	wire n20891;
	wire n20892;
	wire n20893;
	wire n20894;
	wire n20895;
	wire n20896;
	wire n20897;
	wire n20898;
	wire n20899;
	wire n20900;
	wire n20901;
	wire n20902;
	wire n20903;
	wire n20904;
	wire n20905;
	wire n20907;
	wire n20908;
	wire n20909;
	wire n20910;
	wire n20911;
	wire n20912;
	wire n20913;
	wire n20914;
	wire n20915;
	wire n20916;
	wire n20917;
	wire n20918;
	wire n20919;
	wire n20920;
	wire n20921;
	wire n20922;
	wire n20923;
	wire n20924;
	wire n20925;
	wire n20926;
	wire n20927;
	wire n20928;
	wire n20929;
	wire n20930;
	wire n20931;
	wire n20932;
	wire n20933;
	wire n20934;
	wire n20935;
	wire n20936;
	wire n20937;
	wire n20938;
	wire n20939;
	wire n20940;
	wire n20941;
	wire n20942;
	wire n20943;
	wire n20944;
	wire n20945;
	wire n20946;
	wire n20947;
	wire n20948;
	wire n20949;
	wire n20950;
	wire n20951;
	wire n20952;
	wire n20953;
	wire n20954;
	wire n20955;
	wire n20956;
	wire n20957;
	wire n20958;
	wire n20959;
	wire n20960;
	wire n20961;
	wire n20962;
	wire n20963;
	wire n20964;
	wire n20965;
	wire n20966;
	wire n20967;
	wire n20968;
	wire n20969;
	wire n20970;
	wire n20971;
	wire n20972;
	wire n20973;
	wire n20974;
	wire n20975;
	wire n20976;
	wire n20977;
	wire n20978;
	wire n20979;
	wire n20980;
	wire n20981;
	wire n20982;
	wire n20983;
	wire n20984;
	wire n20985;
	wire n20986;
	wire n20987;
	wire n20988;
	wire n20989;
	wire n20990;
	wire n20991;
	wire n20992;
	wire n20993;
	wire n20994;
	wire n20995;
	wire n20996;
	wire n20997;
	wire n20998;
	wire n20999;
	wire n21000;
	wire n21001;
	wire n21002;
	wire n21003;
	wire n21004;
	wire n21005;
	wire n21006;
	wire n21007;
	wire n21008;
	wire n21009;
	wire n21010;
	wire n21011;
	wire n21012;
	wire n21013;
	wire n21014;
	wire n21015;
	wire n21016;
	wire n21017;
	wire n21018;
	wire n21019;
	wire n21020;
	wire n21021;
	wire n21022;
	wire n21023;
	wire n21024;
	wire n21025;
	wire n21026;
	wire n21027;
	wire n21028;
	wire n21029;
	wire n21030;
	wire n21031;
	wire n21032;
	wire n21033;
	wire n21034;
	wire n21035;
	wire n21036;
	wire n21037;
	wire n21038;
	wire n21039;
	wire n21040;
	wire n21041;
	wire n21042;
	wire n21043;
	wire n21044;
	wire n21045;
	wire n21046;
	wire n21047;
	wire n21048;
	wire n21049;
	wire n21050;
	wire n21051;
	wire n21052;
	wire n21053;
	wire n21054;
	wire n21055;
	wire n21056;
	wire n21057;
	wire n21058;
	wire n21059;
	wire n21060;
	wire n21061;
	wire n21062;
	wire n21063;
	wire n21064;
	wire n21065;
	wire n21066;
	wire n21067;
	wire n21068;
	wire n21069;
	wire n21070;
	wire n21071;
	wire n21072;
	wire n21073;
	wire n21074;
	wire n21075;
	wire n21076;
	wire n21077;
	wire n21078;
	wire n21079;
	wire n21080;
	wire n21081;
	wire n21082;
	wire n21083;
	wire n21084;
	wire n21085;
	wire n21086;
	wire n21087;
	wire n21088;
	wire n21089;
	wire n21090;
	wire n21091;
	wire n21092;
	wire n21093;
	wire n21094;
	wire n21095;
	wire n21096;
	wire n21097;
	wire n21098;
	wire n21099;
	wire n21100;
	wire n21101;
	wire n21102;
	wire n21103;
	wire n21104;
	wire n21105;
	wire n21106;
	wire n21107;
	wire n21108;
	wire n21109;
	wire n21110;
	wire n21111;
	wire n21112;
	wire n21113;
	wire n21114;
	wire n21115;
	wire n21116;
	wire n21117;
	wire n21118;
	wire n21119;
	wire n21120;
	wire n21121;
	wire n21122;
	wire n21123;
	wire n21124;
	wire n21125;
	wire n21126;
	wire n21127;
	wire n21128;
	wire n21129;
	wire n21130;
	wire n21131;
	wire n21132;
	wire n21133;
	wire n21134;
	wire n21135;
	wire n21136;
	wire n21137;
	wire n21138;
	wire n21139;
	wire n21140;
	wire n21141;
	wire n21142;
	wire n21143;
	wire n21144;
	wire n21145;
	wire n21146;
	wire n21147;
	wire n21148;
	wire n21149;
	wire n21150;
	wire n21151;
	wire n21152;
	wire n21153;
	wire n21154;
	wire n21155;
	wire n21156;
	wire n21157;
	wire n21158;
	wire n21159;
	wire n21160;
	wire n21161;
	wire n21162;
	wire n21163;
	wire n21164;
	wire n21165;
	wire n21166;
	wire n21167;
	wire n21168;
	wire n21169;
	wire n21170;
	wire n21171;
	wire n21172;
	wire n21173;
	wire n21174;
	wire n21175;
	wire n21176;
	wire n21177;
	wire n21178;
	wire n21179;
	wire n21180;
	wire n21181;
	wire n21182;
	wire n21183;
	wire n21184;
	wire n21185;
	wire n21186;
	wire n21187;
	wire n21188;
	wire n21189;
	wire n21190;
	wire n21191;
	wire n21192;
	wire n21193;
	wire n21194;
	wire n21195;
	wire n21196;
	wire n21197;
	wire n21198;
	wire n21199;
	wire n21200;
	wire n21201;
	wire n21202;
	wire n21203;
	wire n21204;
	wire n21205;
	wire n21206;
	wire n21207;
	wire n21208;
	wire n21209;
	wire n21210;
	wire n21211;
	wire n21212;
	wire n21213;
	wire n21214;
	wire n21215;
	wire n21216;
	wire n21217;
	wire n21218;
	wire n21219;
	wire n21220;
	wire n21221;
	wire n21222;
	wire n21223;
	wire n21224;
	wire n21225;
	wire n21226;
	wire n21227;
	wire n21228;
	wire n21229;
	wire n21230;
	wire n21231;
	wire n21232;
	wire n21233;
	wire n21234;
	wire n21235;
	wire n21236;
	wire n21237;
	wire n21238;
	wire n21239;
	wire n21240;
	wire n21241;
	wire n21242;
	wire n21243;
	wire n21244;
	wire n21245;
	wire n21246;
	wire n21247;
	wire n21248;
	wire n21249;
	wire n21250;
	wire n21251;
	wire n21252;
	wire n21253;
	wire n21254;
	wire n21255;
	wire n21256;
	wire n21257;
	wire n21258;
	wire n21259;
	wire n21260;
	wire n21261;
	wire n21262;
	wire n21263;
	wire n21264;
	wire n21265;
	wire n21266;
	wire n21267;
	wire n21268;
	wire n21269;
	wire n21270;
	wire n21271;
	wire n21272;
	wire n21273;
	wire n21274;
	wire n21275;
	wire n21276;
	wire n21277;
	wire n21278;
	wire n21279;
	wire n21280;
	wire n21281;
	wire n21282;
	wire n21283;
	wire n21284;
	wire n21285;
	wire n21286;
	wire n21287;
	wire n21288;
	wire n21289;
	wire n21290;
	wire n21291;
	wire n21292;
	wire n21293;
	wire n21294;
	wire n21295;
	wire n21296;
	wire n21297;
	wire n21298;
	wire n21299;
	wire n21300;
	wire n21301;
	wire n21302;
	wire n21303;
	wire n21304;
	wire n21305;
	wire n21306;
	wire n21307;
	wire n21308;
	wire n21309;
	wire n21310;
	wire n21311;
	wire n21312;
	wire n21313;
	wire n21314;
	wire n21315;
	wire n21316;
	wire n21317;
	wire n21318;
	wire n21319;
	wire n21320;
	wire n21321;
	wire n21322;
	wire n21323;
	wire n21324;
	wire n21325;
	wire n21326;
	wire n21327;
	wire n21328;
	wire n21329;
	wire n21330;
	wire n21331;
	wire n21332;
	wire n21333;
	wire n21334;
	wire n21335;
	wire n21336;
	wire n21337;
	wire n21338;
	wire n21339;
	wire n21340;
	wire n21341;
	wire n21342;
	wire n21343;
	wire n21344;
	wire n21345;
	wire n21346;
	wire n21347;
	wire n21348;
	wire n21349;
	wire n21350;
	wire n21351;
	wire n21352;
	wire n21353;
	wire n21354;
	wire n21355;
	wire n21356;
	wire n21357;
	wire n21358;
	wire n21359;
	wire n21360;
	wire n21361;
	wire n21362;
	wire n21363;
	wire n21364;
	wire n21365;
	wire n21366;
	wire n21367;
	wire n21368;
	wire n21369;
	wire n21370;
	wire n21371;
	wire n21372;
	wire n21373;
	wire n21374;
	wire n21375;
	wire n21376;
	wire n21377;
	wire n21378;
	wire n21379;
	wire n21380;
	wire n21381;
	wire n21382;
	wire n21383;
	wire n21384;
	wire n21385;
	wire n21386;
	wire n21387;
	wire n21388;
	wire n21389;
	wire n21390;
	wire n21391;
	wire n21392;
	wire n21393;
	wire n21394;
	wire n21395;
	wire n21396;
	wire n21397;
	wire n21398;
	wire n21399;
	wire n21400;
	wire n21401;
	wire n21402;
	wire n21403;
	wire n21404;
	wire n21405;
	wire n21406;
	wire n21407;
	wire n21408;
	wire n21409;
	wire n21410;
	wire n21411;
	wire n21412;
	wire n21413;
	wire n21414;
	wire n21415;
	wire n21416;
	wire n21417;
	wire n21418;
	wire n21419;
	wire n21420;
	wire n21421;
	wire n21422;
	wire n21423;
	wire n21424;
	wire n21425;
	wire n21426;
	wire n21427;
	wire n21428;
	wire n21429;
	wire n21430;
	wire n21431;
	wire n21432;
	wire n21433;
	wire n21434;
	wire n21435;
	wire n21436;
	wire n21437;
	wire n21438;
	wire n21439;
	wire n21440;
	wire n21441;
	wire n21442;
	wire n21443;
	wire n21444;
	wire n21445;
	wire n21446;
	wire n21447;
	wire n21448;
	wire n21449;
	wire n21450;
	wire n21451;
	wire n21452;
	wire n21453;
	wire n21454;
	wire n21455;
	wire n21456;
	wire n21457;
	wire n21458;
	wire n21459;
	wire n21460;
	wire n21461;
	wire n21462;
	wire n21463;
	wire n21464;
	wire n21465;
	wire n21466;
	wire n21467;
	wire n21468;
	wire n21469;
	wire n21470;
	wire n21471;
	wire n21472;
	wire n21473;
	wire n21474;
	wire n21475;
	wire n21476;
	wire n21477;
	wire n21478;
	wire n21479;
	wire n21480;
	wire n21481;
	wire n21482;
	wire n21483;
	wire n21484;
	wire n21485;
	wire n21486;
	wire n21487;
	wire n21488;
	wire n21489;
	wire n21490;
	wire n21491;
	wire n21492;
	wire n21493;
	wire n21494;
	wire n21495;
	wire n21496;
	wire n21497;
	wire n21498;
	wire n21499;
	wire n21500;
	wire n21501;
	wire n21502;
	wire n21503;
	wire n21504;
	wire n21505;
	wire n21506;
	wire n21507;
	wire n21508;
	wire n21509;
	wire n21510;
	wire n21511;
	wire n21512;
	wire n21513;
	wire n21514;
	wire n21515;
	wire n21516;
	wire n21517;
	wire n21518;
	wire n21519;
	wire n21520;
	wire n21521;
	wire n21522;
	wire n21523;
	wire n21524;
	wire n21525;
	wire n21526;
	wire n21527;
	wire n21528;
	wire n21529;
	wire n21530;
	wire n21531;
	wire n21532;
	wire n21533;
	wire n21534;
	wire n21535;
	wire n21536;
	wire n21537;
	wire n21538;
	wire n21539;
	wire n21540;
	wire n21541;
	wire n21542;
	wire n21543;
	wire n21544;
	wire n21545;
	wire n21546;
	wire n21547;
	wire n21548;
	wire n21549;
	wire n21550;
	wire n21551;
	wire n21552;
	wire n21553;
	wire n21554;
	wire n21555;
	wire n21556;
	wire n21557;
	wire n21558;
	wire n21559;
	wire n21560;
	wire n21561;
	wire n21562;
	wire n21563;
	wire n21564;
	wire n21565;
	wire n21566;
	wire n21567;
	wire n21568;
	wire n21569;
	wire n21570;
	wire n21571;
	wire n21572;
	wire n21573;
	wire n21574;
	wire n21575;
	wire n21576;
	wire n21577;
	wire n21578;
	wire n21579;
	wire n21580;
	wire n21581;
	wire n21582;
	wire n21583;
	wire n21584;
	wire n21585;
	wire n21586;
	wire n21587;
	wire n21588;
	wire n21589;
	wire n21590;
	wire n21591;
	wire n21592;
	wire n21593;
	wire n21594;
	wire n21595;
	wire n21596;
	wire n21597;
	wire n21598;
	wire n21599;
	wire n21600;
	wire n21601;
	wire n21602;
	wire n21603;
	wire n21604;
	wire n21605;
	wire n21606;
	wire n21607;
	wire n21608;
	wire n21609;
	wire n21610;
	wire n21611;
	wire n21612;
	wire n21613;
	wire n21614;
	wire n21615;
	wire n21616;
	wire n21617;
	wire n21618;
	wire n21619;
	wire n21620;
	wire n21621;
	wire n21622;
	wire n21623;
	wire n21624;
	wire n21625;
	wire n21626;
	wire n21627;
	wire n21628;
	wire n21629;
	wire n21630;
	wire n21631;
	wire n21632;
	wire n21633;
	wire n21634;
	wire n21635;
	wire n21636;
	wire n21637;
	wire n21638;
	wire n21639;
	wire n21640;
	wire n21641;
	wire n21642;
	wire n21643;
	wire n21644;
	wire n21645;
	wire n21646;
	wire n21647;
	wire n21648;
	wire n21649;
	wire n21650;
	wire n21651;
	wire n21652;
	wire n21653;
	wire n21654;
	wire n21655;
	wire n21656;
	wire n21657;
	wire n21658;
	wire n21659;
	wire n21660;
	wire n21661;
	wire n21662;
	wire n21663;
	wire n21664;
	wire n21665;
	wire n21666;
	wire n21667;
	wire n21668;
	wire n21669;
	wire n21670;
	wire n21671;
	wire n21672;
	wire n21673;
	wire n21674;
	wire n21675;
	wire n21676;
	wire n21677;
	wire n21678;
	wire n21679;
	wire n21680;
	wire n21681;
	wire n21682;
	wire n21683;
	wire n21684;
	wire n21685;
	wire n21686;
	wire n21687;
	wire n21688;
	wire n21689;
	wire n21690;
	wire n21691;
	wire n21692;
	wire n21693;
	wire n21694;
	wire n21695;
	wire n21696;
	wire n21697;
	wire n21698;
	wire n21699;
	wire n21700;
	wire n21701;
	wire n21702;
	wire n21703;
	wire n21704;
	wire n21705;
	wire n21706;
	wire n21707;
	wire n21708;
	wire n21709;
	wire n21710;
	wire n21711;
	wire n21712;
	wire n21713;
	wire n21714;
	wire n21715;
	wire n21716;
	wire n21717;
	wire n21718;
	wire n21719;
	wire n21720;
	wire n21721;
	wire n21722;
	wire n21723;
	wire n21724;
	wire n21725;
	wire n21726;
	wire n21727;
	wire n21728;
	wire n21729;
	wire n21730;
	wire n21731;
	wire n21732;
	wire n21733;
	wire n21734;
	wire n21735;
	wire n21736;
	wire n21737;
	wire n21738;
	wire n21739;
	wire n21740;
	wire n21741;
	wire n21742;
	wire n21743;
	wire n21744;
	wire n21745;
	wire n21746;
	wire n21747;
	wire n21748;
	wire n21749;
	wire n21750;
	wire n21751;
	wire n21752;
	wire n21753;
	wire n21754;
	wire n21755;
	wire n21756;
	wire n21757;
	wire n21758;
	wire n21759;
	wire n21760;
	wire n21761;
	wire n21762;
	wire n21763;
	wire n21764;
	wire n21765;
	wire n21766;
	wire n21767;
	wire n21768;
	wire n21769;
	wire n21770;
	wire n21771;
	wire n21772;
	wire n21773;
	wire n21774;
	wire n21775;
	wire n21776;
	wire n21777;
	wire n21778;
	wire n21779;
	wire n21780;
	wire n21781;
	wire n21782;
	wire n21783;
	wire n21784;
	wire n21785;
	wire n21786;
	wire n21787;
	wire n21788;
	wire n21789;
	wire n21790;
	wire n21791;
	wire n21792;
	wire n21793;
	wire n21794;
	wire n21795;
	wire n21796;
	wire n21797;
	wire n21798;
	wire n21799;
	wire n21800;
	wire n21801;
	wire n21802;
	wire n21803;
	wire n21804;
	wire n21805;
	wire n21806;
	wire n21807;
	wire n21808;
	wire n21809;
	wire n21810;
	wire n21811;
	wire n21812;
	wire n21813;
	wire n21814;
	wire n21815;
	wire n21816;
	wire n21817;
	wire n21818;
	wire n21819;
	wire n21820;
	wire n21821;
	wire n21822;
	wire n21823;
	wire n21824;
	wire n21825;
	wire n21826;
	wire n21827;
	wire n21828;
	wire n21829;
	wire n21830;
	wire n21831;
	wire n21832;
	wire n21833;
	wire n21834;
	wire n21835;
	wire n21836;
	wire n21837;
	wire n21838;
	wire n21839;
	wire n21840;
	wire n21841;
	wire n21842;
	wire n21843;
	wire n21844;
	wire n21845;
	wire n21846;
	wire n21847;
	wire n21848;
	wire n21849;
	wire n21850;
	wire n21851;
	wire n21852;
	wire n21853;
	wire n21854;
	wire n21855;
	wire n21856;
	wire n21857;
	wire n21858;
	wire n21859;
	wire n21860;
	wire n21861;
	wire n21862;
	wire n21863;
	wire n21864;
	wire n21865;
	wire n21866;
	wire n21867;
	wire n21868;
	wire n21869;
	wire n21870;
	wire n21871;
	wire n21872;
	wire n21873;
	wire n21874;
	wire n21875;
	wire n21876;
	wire n21877;
	wire n21878;
	wire n21880;
	wire n21881;
	wire n21882;
	wire n21883;
	wire n21884;
	wire n21885;
	wire n21886;
	wire n21887;
	wire n21888;
	wire n21889;
	wire n21890;
	wire n21891;
	wire n21892;
	wire n21893;
	wire n21894;
	wire n21895;
	wire n21896;
	wire n21897;
	wire n21898;
	wire n21899;
	wire n21900;
	wire n21901;
	wire n21902;
	wire n21903;
	wire n21904;
	wire n21905;
	wire n21906;
	wire n21907;
	wire n21908;
	wire n21909;
	wire n21910;
	wire n21911;
	wire n21912;
	wire n21913;
	wire n21914;
	wire n21915;
	wire n21916;
	wire n21917;
	wire n21918;
	wire n21919;
	wire n21920;
	wire n21921;
	wire n21922;
	wire n21923;
	wire n21924;
	wire n21925;
	wire n21926;
	wire n21927;
	wire n21928;
	wire n21929;
	wire n21930;
	wire n21931;
	wire n21932;
	wire n21933;
	wire n21934;
	wire n21935;
	wire n21936;
	wire n21937;
	wire n21938;
	wire n21939;
	wire n21940;
	wire n21941;
	wire n21942;
	wire n21943;
	wire n21944;
	wire n21945;
	wire n21946;
	wire n21947;
	wire n21948;
	wire n21949;
	wire n21950;
	wire n21951;
	wire n21952;
	wire n21953;
	wire n21954;
	wire n21955;
	wire n21956;
	wire n21957;
	wire n21958;
	wire n21959;
	wire n21960;
	wire n21961;
	wire n21962;
	wire n21963;
	wire n21964;
	wire n21965;
	wire n21966;
	wire n21967;
	wire n21968;
	wire n21969;
	wire n21970;
	wire n21971;
	wire n21972;
	wire n21973;
	wire n21974;
	wire n21975;
	wire n21976;
	wire n21977;
	wire n21978;
	wire n21979;
	wire n21980;
	wire n21981;
	wire n21982;
	wire n21983;
	wire n21984;
	wire n21985;
	wire n21986;
	wire n21987;
	wire n21988;
	wire n21989;
	wire n21990;
	wire n21991;
	wire n21992;
	wire n21993;
	wire n21994;
	wire n21995;
	wire n21996;
	wire n21997;
	wire n21998;
	wire n21999;
	wire n22000;
	wire n22001;
	wire n22002;
	wire n22003;
	wire n22004;
	wire n22005;
	wire n22006;
	wire n22007;
	wire n22008;
	wire n22009;
	wire n22010;
	wire n22011;
	wire n22012;
	wire n22013;
	wire n22014;
	wire n22015;
	wire n22016;
	wire n22017;
	wire n22018;
	wire n22019;
	wire n22020;
	wire n22021;
	wire n22022;
	wire n22023;
	wire n22024;
	wire n22025;
	wire n22026;
	wire n22027;
	wire n22028;
	wire n22029;
	wire n22030;
	wire n22031;
	wire n22032;
	wire n22033;
	wire n22034;
	wire n22035;
	wire n22036;
	wire n22037;
	wire n22038;
	wire n22039;
	wire n22040;
	wire n22041;
	wire n22042;
	wire n22043;
	wire n22044;
	wire n22045;
	wire n22046;
	wire n22047;
	wire n22048;
	wire n22049;
	wire n22050;
	wire n22051;
	wire n22052;
	wire n22053;
	wire n22054;
	wire n22055;
	wire n22056;
	wire n22057;
	wire n22058;
	wire n22059;
	wire n22060;
	wire n22061;
	wire n22062;
	wire n22063;
	wire n22064;
	wire n22065;
	wire n22066;
	wire n22067;
	wire n22068;
	wire n22069;
	wire n22070;
	wire n22071;
	wire n22072;
	wire n22073;
	wire n22074;
	wire n22075;
	wire n22076;
	wire n22077;
	wire n22078;
	wire n22079;
	wire n22080;
	wire n22081;
	wire n22082;
	wire n22083;
	wire n22084;
	wire n22085;
	wire n22086;
	wire n22087;
	wire n22088;
	wire n22089;
	wire n22090;
	wire n22091;
	wire n22092;
	wire n22093;
	wire n22094;
	wire n22095;
	wire n22096;
	wire n22097;
	wire n22098;
	wire n22099;
	wire n22100;
	wire n22101;
	wire n22102;
	wire n22103;
	wire n22104;
	wire n22105;
	wire n22106;
	wire n22107;
	wire n22108;
	wire n22109;
	wire n22110;
	wire n22111;
	wire n22112;
	wire n22113;
	wire n22114;
	wire n22115;
	wire n22116;
	wire n22117;
	wire n22118;
	wire n22119;
	wire n22120;
	wire n22121;
	wire n22122;
	wire n22123;
	wire n22124;
	wire n22125;
	wire n22126;
	wire n22127;
	wire n22128;
	wire n22129;
	wire n22130;
	wire n22131;
	wire n22132;
	wire n22133;
	wire n22134;
	wire n22135;
	wire n22136;
	wire n22137;
	wire n22138;
	wire n22139;
	wire n22140;
	wire n22141;
	wire n22142;
	wire n22143;
	wire n22144;
	wire n22145;
	wire n22146;
	wire n22147;
	wire n22148;
	wire n22149;
	wire n22150;
	wire n22151;
	wire n22152;
	wire n22153;
	wire n22154;
	wire n22155;
	wire n22156;
	wire n22157;
	wire n22158;
	wire n22159;
	wire n22160;
	wire n22161;
	wire n22162;
	wire n22163;
	wire n22164;
	wire n22165;
	wire n22166;
	wire n22167;
	wire n22168;
	wire n22169;
	wire n22170;
	wire n22171;
	wire n22172;
	wire n22173;
	wire n22174;
	wire n22175;
	wire n22176;
	wire n22177;
	wire n22178;
	wire n22179;
	wire n22180;
	wire n22181;
	wire n22182;
	wire n22183;
	wire n22184;
	wire n22185;
	wire n22186;
	wire n22187;
	wire n22188;
	wire n22189;
	wire n22190;
	wire n22191;
	wire n22192;
	wire n22193;
	wire n22194;
	wire n22195;
	wire n22196;
	wire n22197;
	wire n22198;
	wire n22199;
	wire n22200;
	wire n22201;
	wire n22202;
	wire n22203;
	wire n22204;
	wire n22205;
	wire n22206;
	wire n22207;
	wire n22208;
	wire n22209;
	wire n22210;
	wire n22211;
	wire n22212;
	wire n22213;
	wire n22214;
	wire n22215;
	wire n22216;
	wire n22217;
	wire n22218;
	wire n22219;
	wire n22220;
	wire n22221;
	wire n22222;
	wire n22223;
	wire n22224;
	wire n22225;
	wire n22226;
	wire n22227;
	wire n22228;
	wire n22229;
	wire n22230;
	wire n22231;
	wire n22232;
	wire n22233;
	wire n22234;
	wire n22235;
	wire n22236;
	wire n22237;
	wire n22238;
	wire n22239;
	wire n22240;
	wire n22241;
	wire n22242;
	wire n22243;
	wire n22244;
	wire n22245;
	wire n22246;
	wire n22247;
	wire n22248;
	wire n22249;
	wire n22250;
	wire n22251;
	wire n22252;
	wire n22253;
	wire n22254;
	wire n22255;
	wire n22256;
	wire n22257;
	wire n22258;
	wire n22259;
	wire n22260;
	wire n22261;
	wire n22262;
	wire n22263;
	wire n22264;
	wire n22265;
	wire n22266;
	wire n22267;
	wire n22268;
	wire n22269;
	wire n22270;
	wire n22271;
	wire n22272;
	wire n22273;
	wire n22274;
	wire n22275;
	wire n22276;
	wire n22277;
	wire n22278;
	wire n22279;
	wire n22280;
	wire n22281;
	wire n22282;
	wire n22283;
	wire n22284;
	wire n22285;
	wire n22286;
	wire n22287;
	wire n22288;
	wire n22289;
	wire n22290;
	wire n22291;
	wire n22292;
	wire n22293;
	wire n22294;
	wire n22295;
	wire n22296;
	wire n22297;
	wire n22298;
	wire n22299;
	wire n22300;
	wire n22301;
	wire n22302;
	wire n22303;
	wire n22304;
	wire n22305;
	wire n22306;
	wire n22307;
	wire n22308;
	wire n22309;
	wire n22310;
	wire n22311;
	wire n22312;
	wire n22313;
	wire n22314;
	wire n22315;
	wire n22316;
	wire n22317;
	wire n22318;
	wire n22319;
	wire n22320;
	wire n22321;
	wire n22322;
	wire n22323;
	wire n22324;
	wire n22325;
	wire n22326;
	wire n22327;
	wire n22328;
	wire n22329;
	wire n22330;
	wire n22331;
	wire n22332;
	wire n22334;
	wire n22335;
	wire n22336;
	wire n22337;
	wire n22338;
	wire n22339;
	wire n22340;
	wire n22341;
	wire n22342;
	wire n22343;
	wire n22344;
	wire n22345;
	wire n22346;
	wire n22347;
	wire n22348;
	wire n22349;
	wire n22350;
	wire n22351;
	wire n22352;
	wire n22353;
	wire n22354;
	wire n22355;
	wire n22356;
	wire n22357;
	wire n22358;
	wire n22359;
	wire n22360;
	wire n22361;
	wire n22362;
	wire n22363;
	wire n22364;
	wire n22365;
	wire n22366;
	wire n22367;
	wire n22368;
	wire n22369;
	wire n22370;
	wire n22371;
	wire n22372;
	wire n22373;
	wire n22374;
	wire n22375;
	wire n22376;
	wire n22377;
	wire n22378;
	wire n22379;
	wire n22380;
	wire n22381;
	wire n22382;
	wire n22383;
	wire n22384;
	wire n22385;
	wire n22386;
	wire n22387;
	wire n22388;
	wire n22389;
	wire n22390;
	wire n22391;
	wire n22392;
	wire n22393;
	wire n22394;
	wire n22395;
	wire n22396;
	wire n22397;
	wire n22398;
	wire n22399;
	wire n22400;
	wire n22401;
	wire n22402;
	wire n22403;
	wire n22404;
	wire n22405;
	wire n22406;
	wire n22407;
	wire n22408;
	wire n22409;
	wire n22410;
	wire n22411;
	wire n22412;
	wire n22413;
	wire n22414;
	wire n22415;
	wire n22416;
	wire n22417;
	wire n22418;
	wire n22419;
	wire n22420;
	wire n22421;
	wire n22422;
	wire n22423;
	wire n22424;
	wire n22425;
	wire n22426;
	wire n22427;
	wire n22428;
	wire n22429;
	wire n22430;
	wire n22431;
	wire n22432;
	wire n22433;
	wire n22434;
	wire n22435;
	wire n22436;
	wire n22437;
	wire n22438;
	wire n22439;
	wire n22440;
	wire n22441;
	wire n22442;
	wire n22443;
	wire n22444;
	wire n22445;
	wire n22446;
	wire n22447;
	wire n22448;
	wire n22449;
	wire n22450;
	wire n22451;
	wire n22452;
	wire n22453;
	wire n22454;
	wire n22455;
	wire n22456;
	wire n22457;
	wire n22458;
	wire n22459;
	wire n22460;
	wire n22461;
	wire n22462;
	wire n22463;
	wire n22464;
	wire n22465;
	wire n22466;
	wire n22467;
	wire n22468;
	wire n22469;
	wire n22470;
	wire n22471;
	wire n22472;
	wire n22473;
	wire n22474;
	wire n22475;
	wire n22476;
	wire n22477;
	wire n22478;
	wire n22479;
	wire n22480;
	wire n22481;
	wire n22482;
	wire n22483;
	wire n22484;
	wire n22485;
	wire n22486;
	wire n22487;
	wire n22488;
	wire n22489;
	wire n22490;
	wire n22491;
	wire n22492;
	wire n22493;
	wire n22494;
	wire n22495;
	wire n22496;
	wire n22497;
	wire n22498;
	wire n22499;
	wire n22500;
	wire n22501;
	wire n22502;
	wire n22503;
	wire n22504;
	wire n22505;
	wire n22506;
	wire n22507;
	wire n22508;
	wire n22509;
	wire n22510;
	wire n22511;
	wire n22512;
	wire n22513;
	wire n22514;
	wire n22515;
	wire n22516;
	wire n22517;
	wire n22518;
	wire n22519;
	wire n22520;
	wire n22521;
	wire n22522;
	wire n22523;
	wire n22524;
	wire n22525;
	wire n22526;
	wire n22527;
	wire n22528;
	wire n22529;
	wire n22530;
	wire n22531;
	wire n22532;
	wire n22533;
	wire n22534;
	wire n22535;
	wire n22536;
	wire n22537;
	wire n22538;
	wire n22539;
	wire n22540;
	wire n22541;
	wire n22542;
	wire n22543;
	wire n22544;
	wire n22545;
	wire n22546;
	wire n22547;
	wire n22548;
	wire n22549;
	wire n22550;
	wire n22551;
	wire n22552;
	wire n22553;
	wire n22554;
	wire n22555;
	wire n22556;
	wire n22557;
	wire n22558;
	wire n22559;
	wire n22560;
	wire n22561;
	wire n22562;
	wire n22563;
	wire n22564;
	wire n22565;
	wire n22566;
	wire n22567;
	wire n22568;
	wire n22569;
	wire n22570;
	wire n22571;
	wire n22572;
	wire n22573;
	wire n22574;
	wire n22575;
	wire n22576;
	wire n22577;
	wire n22578;
	wire n22579;
	wire n22580;
	wire n22581;
	wire n22582;
	wire n22583;
	wire n22584;
	wire n22585;
	wire n22586;
	wire n22587;
	wire n22588;
	wire n22589;
	wire n22590;
	wire n22591;
	wire n22592;
	wire n22593;
	wire n22594;
	wire n22595;
	wire n22596;
	wire n22597;
	wire n22598;
	wire n22599;
	wire n22600;
	wire n22601;
	wire n22602;
	wire n22603;
	wire n22604;
	wire n22605;
	wire n22606;
	wire n22607;
	wire n22608;
	wire n22609;
	wire n22610;
	wire n22611;
	wire n22612;
	wire n22613;
	wire n22614;
	wire n22615;
	wire n22616;
	wire n22617;
	wire n22618;
	wire n22619;
	wire n22620;
	wire n22621;
	wire n22622;
	wire n22623;
	wire n22624;
	wire n22625;
	wire n22626;
	wire n22627;
	wire n22628;
	wire n22629;
	wire n22630;
	wire n22631;
	wire n22632;
	wire n22633;
	wire n22634;
	wire n22635;
	wire n22636;
	wire n22637;
	wire n22638;
	wire n22639;
	wire n22640;
	wire n22641;
	wire n22642;
	wire n22643;
	wire n22644;
	wire n22645;
	wire n22646;
	wire n22647;
	wire n22648;
	wire n22649;
	wire n22650;
	wire n22651;
	wire n22652;
	wire n22653;
	wire n22654;
	wire n22655;
	wire n22656;
	wire n22657;
	wire n22658;
	wire n22659;
	wire n22660;
	wire n22661;
	wire n22662;
	wire n22663;
	wire n22664;
	wire n22665;
	wire n22666;
	wire n22667;
	wire n22668;
	wire n22669;
	wire n22670;
	wire n22671;
	wire n22672;
	wire n22673;
	wire n22674;
	wire n22675;
	wire n22676;
	wire n22677;
	wire n22678;
	wire n22679;
	wire n22680;
	wire n22681;
	wire n22682;
	wire n22683;
	wire n22684;
	wire n22685;
	wire n22686;
	wire n22687;
	wire n22688;
	wire n22689;
	wire n22690;
	wire n22691;
	wire n22692;
	wire n22693;
	wire n22694;
	wire n22695;
	wire n22696;
	wire n22697;
	wire n22698;
	wire n22699;
	wire n22700;
	wire n22701;
	wire n22702;
	wire n22703;
	wire n22704;
	wire n22705;
	wire n22706;
	wire n22707;
	wire n22708;
	wire n22709;
	wire n22710;
	wire n22711;
	wire n22712;
	wire n22713;
	wire n22714;
	wire n22715;
	wire n22716;
	wire n22717;
	wire n22718;
	wire n22719;
	wire n22720;
	wire n22721;
	wire n22722;
	wire n22723;
	wire n22724;
	wire n22725;
	wire n22726;
	wire n22727;
	wire n22728;
	wire n22729;
	wire n22730;
	wire n22731;
	wire n22732;
	wire n22733;
	wire n22734;
	wire n22735;
	wire n22736;
	wire n22737;
	wire n22738;
	wire n22739;
	wire n22740;
	wire n22741;
	wire n22742;
	wire n22743;
	wire n22744;
	wire n22745;
	wire n22746;
	wire n22747;
	wire n22748;
	wire n22749;
	wire n22750;
	wire n22751;
	wire n22752;
	wire n22753;
	wire n22754;
	wire n22755;
	wire n22756;
	wire n22757;
	wire n22758;
	wire n22759;
	wire n22760;
	wire n22761;
	wire n22762;
	wire n22763;
	wire n22764;
	wire n22765;
	wire n22766;
	wire n22767;
	wire n22768;
	wire n22769;
	wire n22770;
	wire n22771;
	wire n22772;
	wire n22773;
	wire n22774;
	wire n22775;
	wire n22776;
	wire n22777;
	wire n22778;
	wire n22779;
	wire n22780;
	wire n22781;
	wire n22782;
	wire n22783;
	wire n22784;
	wire n22785;
	wire n22786;
	wire n22787;
	wire n22788;
	wire n22789;
	wire n22790;
	wire n22791;
	wire n22792;
	wire n22793;
	wire n22794;
	wire n22795;
	wire n22796;
	wire n22797;
	wire n22798;
	wire n22799;
	wire n22800;
	wire n22801;
	wire n22802;
	wire n22803;
	wire n22804;
	wire n22805;
	wire n22806;
	wire n22807;
	wire n22808;
	wire n22809;
	wire n22810;
	wire n22811;
	wire n22812;
	wire n22813;
	wire n22814;
	wire n22815;
	wire n22816;
	wire n22817;
	wire n22818;
	wire n22819;
	wire n22820;
	wire n22821;
	wire n22822;
	wire n22823;
	wire n22824;
	wire n22825;
	wire n22826;
	wire n22827;
	wire n22828;
	wire n22829;
	wire n22830;
	wire n22831;
	wire n22832;
	wire n22833;
	wire n22834;
	wire n22835;
	wire n22836;
	wire n22837;
	wire n22838;
	wire n22839;
	wire n22840;
	wire n22841;
	wire n22842;
	wire n22843;
	wire n22844;
	wire n22845;
	wire n22846;
	wire n22847;
	wire n22848;
	wire n22849;
	wire n22850;
	wire n22851;
	wire n22852;
	wire n22853;
	wire n22854;
	wire n22855;
	wire n22856;
	wire n22857;
	wire n22858;
	wire n22859;
	wire n22860;
	wire n22861;
	wire n22862;
	wire n22863;
	wire n22864;
	wire n22865;
	wire n22866;
	wire n22867;
	wire n22868;
	wire n22869;
	wire n22870;
	wire n22871;
	wire n22872;
	wire n22873;
	wire n22874;
	wire n22875;
	wire n22876;
	wire n22877;
	wire n22878;
	wire n22879;
	wire n22880;
	wire n22881;
	wire n22882;
	wire n22883;
	wire n22884;
	wire n22885;
	wire n22886;
	wire n22887;
	wire n22888;
	wire n22889;
	wire n22890;
	wire n22891;
	wire n22892;
	wire n22893;
	wire n22894;
	wire n22895;
	wire n22896;
	wire n22897;
	wire n22898;
	wire n22899;
	wire n22900;
	wire n22901;
	wire n22902;
	wire n22903;
	wire n22904;
	wire n22905;
	wire n22906;
	wire n22907;
	wire n22908;
	wire n22909;
	wire n22910;
	wire n22911;
	wire n22912;
	wire n22913;
	wire n22914;
	wire n22915;
	wire n22916;
	wire n22917;
	wire n22918;
	wire n22919;
	wire n22920;
	wire n22921;
	wire n22922;
	wire n22923;
	wire n22924;
	wire n22925;
	wire n22926;
	wire n22927;
	wire n22928;
	wire n22929;
	wire n22930;
	wire n22931;
	wire n22932;
	wire n22933;
	wire n22934;
	wire n22935;
	wire n22936;
	wire n22937;
	wire n22938;
	wire n22939;
	wire n22940;
	wire n22941;
	wire n22942;
	wire n22943;
	wire n22944;
	wire n22945;
	wire n22946;
	wire n22947;
	wire n22948;
	wire n22949;
	wire n22950;
	wire n22951;
	wire n22952;
	wire n22953;
	wire n22954;
	wire n22955;
	wire n22956;
	wire n22957;
	wire n22958;
	wire n22959;
	wire n22960;
	wire n22961;
	wire n22962;
	wire n22963;
	wire n22964;
	wire n22965;
	wire n22966;
	wire n22967;
	wire n22968;
	wire n22969;
	wire n22970;
	wire n22971;
	wire n22972;
	wire n22973;
	wire n22974;
	wire n22975;
	wire n22976;
	wire n22977;
	wire n22978;
	wire n22979;
	wire n22980;
	wire n22981;
	wire n22982;
	wire n22983;
	wire n22984;
	wire n22985;
	wire n22986;
	wire n22987;
	wire n22988;
	wire n22989;
	wire n22990;
	wire n22991;
	wire n22992;
	wire n22993;
	wire n22994;
	wire n22995;
	wire n22996;
	wire n22997;
	wire n22998;
	wire n22999;
	wire n23000;
	wire n23001;
	wire n23002;
	wire n23003;
	wire n23004;
	wire n23005;
	wire n23006;
	wire n23007;
	wire n23008;
	wire n23009;
	wire n23010;
	wire n23011;
	wire n23012;
	wire n23013;
	wire n23014;
	wire n23015;
	wire n23016;
	wire n23017;
	wire n23018;
	wire n23019;
	wire n23020;
	wire n23021;
	wire n23022;
	wire n23023;
	wire n23024;
	wire n23025;
	wire n23026;
	wire n23027;
	wire n23028;
	wire n23029;
	wire n23030;
	wire n23031;
	wire n23032;
	wire n23033;
	wire n23034;
	wire n23035;
	wire n23036;
	wire n23037;
	wire n23038;
	wire n23039;
	wire n23040;
	wire n23041;
	wire n23042;
	wire n23043;
	wire n23044;
	wire n23045;
	wire n23046;
	wire n23047;
	wire n23048;
	wire n23049;
	wire n23050;
	wire n23051;
	wire n23052;
	wire n23053;
	wire n23054;
	wire n23055;
	wire n23056;
	wire n23057;
	wire n23058;
	wire n23059;
	wire n23060;
	wire n23061;
	wire n23062;
	wire n23063;
	wire n23064;
	wire n23065;
	wire n23066;
	wire n23067;
	wire n23068;
	wire n23069;
	wire n23070;
	wire n23071;
	wire n23072;
	wire n23073;
	wire n23074;
	wire n23075;
	wire n23076;
	wire n23077;
	wire n23078;
	wire n23079;
	wire n23080;
	wire n23081;
	wire n23082;
	wire n23083;
	wire n23084;
	wire n23085;
	wire n23086;
	wire n23087;
	wire n23088;
	wire n23089;
	wire n23090;
	wire n23091;
	wire n23092;
	wire n23093;
	wire n23094;
	wire n23095;
	wire n23096;
	wire n23097;
	wire n23098;
	wire n23099;
	wire n23100;
	wire n23101;
	wire n23102;
	wire n23103;
	wire n23104;
	wire n23105;
	wire n23106;
	wire n23107;
	wire n23108;
	wire n23109;
	wire n23110;
	wire n23111;
	wire n23112;
	wire n23113;
	wire n23114;
	wire n23115;
	wire n23116;
	wire n23117;
	wire n23118;
	wire n23119;
	wire n23120;
	wire n23121;
	wire n23122;
	wire n23123;
	wire n23124;
	wire n23125;
	wire n23126;
	wire n23127;
	wire n23128;
	wire n23129;
	wire n23130;
	wire n23131;
	wire n23132;
	wire n23133;
	wire n23134;
	wire n23135;
	wire n23136;
	wire n23137;
	wire n23138;
	wire n23139;
	wire n23140;
	wire n23141;
	wire n23142;
	wire n23143;
	wire n23144;
	wire n23145;
	wire n23146;
	wire n23147;
	wire n23148;
	wire n23149;
	wire n23150;
	wire n23151;
	wire n23152;
	wire n23153;
	wire n23154;
	wire n23155;
	wire n23156;
	wire n23157;
	wire n23158;
	wire n23159;
	wire n23160;
	wire n23161;
	wire n23162;
	wire n23163;
	wire n23164;
	wire n23165;
	wire n23166;
	wire n23167;
	wire n23168;
	wire n23169;
	wire n23170;
	wire n23171;
	wire n23172;
	wire n23173;
	wire n23174;
	wire n23175;
	wire n23176;
	wire n23177;
	wire n23178;
	wire n23179;
	wire n23180;
	wire n23181;
	wire n23182;
	wire n23183;
	wire n23184;
	wire n23185;
	wire n23186;
	wire n23187;
	wire n23188;
	wire n23189;
	wire n23190;
	wire n23191;
	wire n23192;
	wire n23193;
	wire n23194;
	wire n23195;
	wire n23196;
	wire n23197;
	wire n23198;
	wire n23199;
	wire n23200;
	wire n23201;
	wire n23202;
	wire n23203;
	wire n23204;
	wire n23205;
	wire n23206;
	wire n23207;
	wire n23208;
	wire n23209;
	wire n23210;
	wire n23211;
	wire n23212;
	wire n23213;
	wire n23214;
	wire n23215;
	wire n23216;
	wire n23217;
	wire n23218;
	wire n23219;
	wire n23220;
	wire n23221;
	wire n23222;
	wire n23223;
	wire n23224;
	wire n23225;
	wire n23226;
	wire n23227;
	wire n23228;
	wire n23229;
	wire n23230;
	wire n23231;
	wire n23232;
	wire n23233;
	wire n23234;
	wire n23235;
	wire n23236;
	wire n23237;
	wire n23238;
	wire n23239;
	wire n23240;
	wire n23241;
	wire n23242;
	wire n23243;
	wire n23244;
	wire n23245;
	wire n23246;
	wire n23247;
	wire n23248;
	wire n23249;
	wire n23250;
	wire n23251;
	wire n23252;
	wire n23253;
	wire n23254;
	wire n23255;
	wire n23256;
	wire n23257;
	wire n23258;
	wire n23259;
	wire n23260;
	wire n23261;
	wire n23262;
	wire n23263;
	wire n23264;
	wire n23265;
	wire n23266;
	wire n23267;
	wire n23268;
	wire n23269;
	wire n23270;
	wire n23271;
	wire n23272;
	wire n23273;
	wire n23274;
	wire n23275;
	wire n23276;
	wire n23277;
	wire n23278;
	wire n23279;
	wire n23280;
	wire n23281;
	wire n23282;
	wire n23283;
	wire n23284;
	wire n23285;
	wire n23286;
	wire n23287;
	wire n23288;
	wire n23289;
	wire n23290;
	wire n23291;
	wire n23292;
	wire n23293;
	wire n23294;
	wire n23295;
	wire n23296;
	wire n23297;
	wire n23298;
	wire n23299;
	wire n23300;
	wire n23301;
	wire n23302;
	wire n23303;
	wire n23304;
	wire n23305;
	wire n23306;
	wire n23307;
	wire n23308;
	wire n23309;
	wire n23310;
	wire n23311;
	wire n23312;
	wire n23313;
	wire n23314;
	wire n23315;
	wire n23316;
	wire n23317;
	wire n23318;
	wire n23319;
	wire n23320;
	wire n23321;
	wire n23322;
	wire n23323;
	wire n23324;
	wire n23325;
	wire n23326;
	wire n23327;
	wire n23328;
	wire n23329;
	wire n23330;
	wire n23331;
	wire n23332;
	wire n23333;
	wire n23334;
	wire n23335;
	wire n23336;
	wire n23338;
	wire n23339;
	wire n23340;
	wire n23341;
	wire n23342;
	wire n23343;
	wire n23344;
	wire n23345;
	wire n23346;
	wire n23347;
	wire n23348;
	wire n23349;
	wire n23350;
	wire n23351;
	wire n23352;
	wire n23353;
	wire n23354;
	wire n23355;
	wire n23356;
	wire n23357;
	wire n23358;
	wire n23359;
	wire n23360;
	wire n23361;
	wire n23362;
	wire n23363;
	wire n23364;
	wire n23365;
	wire n23366;
	wire n23367;
	wire n23368;
	wire n23369;
	wire n23370;
	wire n23371;
	wire n23372;
	wire n23373;
	wire n23374;
	wire n23375;
	wire n23376;
	wire n23377;
	wire n23378;
	wire n23379;
	wire n23380;
	wire n23381;
	wire n23382;
	wire n23383;
	wire n23384;
	wire n23385;
	wire n23386;
	wire n23387;
	wire n23388;
	wire n23389;
	wire n23390;
	wire n23391;
	wire n23392;
	wire n23393;
	wire n23394;
	wire n23395;
	wire n23396;
	wire n23397;
	wire n23398;
	wire n23399;
	wire n23400;
	wire n23401;
	wire n23402;
	wire n23403;
	wire n23404;
	wire n23405;
	wire n23406;
	wire n23407;
	wire n23408;
	wire n23409;
	wire n23410;
	wire n23411;
	wire n23412;
	wire n23413;
	wire n23414;
	wire n23415;
	wire n23416;
	wire n23417;
	wire n23418;
	wire n23419;
	wire n23420;
	wire n23421;
	wire n23422;
	wire n23423;
	wire n23424;
	wire n23425;
	wire n23426;
	wire n23427;
	wire n23428;
	wire n23429;
	wire n23430;
	wire n23431;
	wire n23432;
	wire n23433;
	wire n23434;
	wire n23435;
	wire n23436;
	wire n23437;
	wire n23438;
	wire n23439;
	wire n23440;
	wire n23441;
	wire n23442;
	wire n23443;
	wire n23444;
	wire n23445;
	wire n23446;
	wire n23447;
	wire n23448;
	wire n23449;
	wire n23450;
	wire n23451;
	wire n23452;
	wire n23453;
	wire n23454;
	wire n23455;
	wire n23456;
	wire n23457;
	wire n23458;
	wire n23459;
	wire n23460;
	wire n23461;
	wire n23462;
	wire n23463;
	wire n23464;
	wire n23465;
	wire n23466;
	wire n23467;
	wire n23468;
	wire n23469;
	wire n23470;
	wire n23471;
	wire n23472;
	wire n23473;
	wire n23474;
	wire n23475;
	wire n23476;
	wire n23477;
	wire n23478;
	wire n23479;
	wire n23480;
	wire n23481;
	wire n23482;
	wire n23483;
	wire n23484;
	wire n23485;
	wire n23486;
	wire n23487;
	wire n23488;
	wire n23489;
	wire n23490;
	wire n23491;
	wire n23492;
	wire n23493;
	wire n23494;
	wire n23495;
	wire n23496;
	wire n23497;
	wire n23498;
	wire n23499;
	wire n23500;
	wire n23501;
	wire n23502;
	wire n23503;
	wire n23504;
	wire n23505;
	wire n23506;
	wire n23507;
	wire n23508;
	wire n23509;
	wire n23510;
	wire n23511;
	wire n23512;
	wire n23513;
	wire n23514;
	wire n23515;
	wire n23516;
	wire n23517;
	wire n23518;
	wire n23519;
	wire n23520;
	wire n23521;
	wire n23522;
	wire n23523;
	wire n23524;
	wire n23525;
	wire n23526;
	wire n23527;
	wire n23528;
	wire n23529;
	wire n23530;
	wire n23531;
	wire n23532;
	wire n23533;
	wire n23534;
	wire n23535;
	wire n23536;
	wire n23537;
	wire n23538;
	wire n23539;
	wire n23540;
	wire n23541;
	wire n23542;
	wire n23543;
	wire n23544;
	wire n23545;
	wire n23546;
	wire n23547;
	wire n23548;
	wire n23549;
	wire n23550;
	wire n23551;
	wire n23552;
	wire n23553;
	wire n23554;
	wire n23555;
	wire n23556;
	wire n23557;
	wire n23558;
	wire n23559;
	wire n23560;
	wire n23561;
	wire n23562;
	wire n23563;
	wire n23564;
	wire n23565;
	wire n23566;
	wire n23567;
	wire n23568;
	wire n23569;
	wire n23570;
	wire n23571;
	wire n23572;
	wire n23573;
	wire n23574;
	wire n23575;
	wire n23576;
	wire n23577;
	wire n23578;
	wire n23579;
	wire n23580;
	wire n23581;
	wire n23582;
	wire n23583;
	wire n23584;
	wire n23585;
	wire n23586;
	wire n23587;
	wire n23588;
	wire n23589;
	wire n23590;
	wire n23591;
	wire n23592;
	wire n23593;
	wire n23594;
	wire n23595;
	wire n23596;
	wire n23597;
	wire n23598;
	wire n23599;
	wire n23600;
	wire n23601;
	wire n23602;
	wire n23603;
	wire n23604;
	wire n23605;
	wire n23606;
	wire n23607;
	wire n23608;
	wire n23609;
	wire n23610;
	wire n23611;
	wire n23612;
	wire n23613;
	wire n23614;
	wire n23615;
	wire n23616;
	wire n23617;
	wire n23618;
	wire n23619;
	wire n23620;
	wire n23621;
	wire n23622;
	wire n23623;
	wire n23624;
	wire n23625;
	wire n23626;
	wire n23627;
	wire n23628;
	wire n23629;
	wire n23630;
	wire n23631;
	wire n23632;
	wire n23633;
	wire n23634;
	wire n23635;
	wire n23636;
	wire n23637;
	wire n23638;
	wire n23639;
	wire n23640;
	wire n23641;
	wire n23642;
	wire n23643;
	wire n23644;
	wire n23645;
	wire n23646;
	wire n23647;
	wire n23648;
	wire n23649;
	wire n23650;
	wire n23651;
	wire n23652;
	wire n23653;
	wire n23654;
	wire n23655;
	wire n23656;
	wire n23657;
	wire n23658;
	wire n23659;
	wire n23660;
	wire n23661;
	wire n23662;
	wire n23663;
	wire n23664;
	wire n23665;
	wire n23666;
	wire n23667;
	wire n23668;
	wire n23669;
	wire n23670;
	wire n23671;
	wire n23672;
	wire n23673;
	wire n23674;
	wire n23675;
	wire n23676;
	wire n23677;
	wire n23678;
	wire n23679;
	wire n23680;
	wire n23681;
	wire n23682;
	wire n23683;
	wire n23684;
	wire n23685;
	wire n23686;
	wire n23687;
	wire n23688;
	wire n23689;
	wire n23690;
	wire n23691;
	wire n23692;
	wire n23693;
	wire n23694;
	wire n23695;
	wire n23696;
	wire n23697;
	wire n23698;
	wire n23699;
	wire n23700;
	wire n23701;
	wire n23702;
	wire n23703;
	wire n23704;
	wire n23705;
	wire n23706;
	wire n23707;
	wire n23708;
	wire n23709;
	wire n23710;
	wire n23711;
	wire n23712;
	wire n23713;
	wire n23714;
	wire n23715;
	wire n23716;
	wire n23717;
	wire n23718;
	wire n23719;
	wire n23720;
	wire n23721;
	wire n23722;
	wire n23723;
	wire n23724;
	wire n23725;
	wire n23726;
	wire n23727;
	wire n23728;
	wire n23729;
	wire n23730;
	wire n23731;
	wire n23732;
	wire n23733;
	wire n23734;
	wire n23735;
	wire n23736;
	wire n23737;
	wire n23738;
	wire n23739;
	wire n23740;
	wire n23741;
	wire n23742;
	wire n23743;
	wire n23744;
	wire n23745;
	wire n23746;
	wire n23747;
	wire n23748;
	wire n23749;
	wire n23750;
	wire n23751;
	wire n23752;
	wire n23753;
	wire n23754;
	wire n23755;
	wire n23756;
	wire n23757;
	wire n23758;
	wire n23759;
	wire n23760;
	wire n23761;
	wire n23762;
	wire n23763;
	wire n23764;
	wire n23765;
	wire n23766;
	wire n23767;
	wire n23768;
	wire n23769;
	wire n23770;
	wire n23771;
	wire n23772;
	wire n23773;
	wire n23774;
	wire n23775;
	wire n23776;
	wire n23777;
	wire n23778;
	wire n23779;
	wire n23780;
	wire n23781;
	wire n23782;
	wire n23783;
	wire n23784;
	wire n23785;
	wire n23786;
	wire n23787;
	wire n23788;
	wire n23789;
	wire n23790;
	wire n23791;
	wire n23792;
	wire n23793;
	wire n23794;
	wire n23795;
	wire n23796;
	wire n23797;
	wire n23798;
	wire n23799;
	wire n23800;
	wire n23801;
	wire n23802;
	wire n23803;
	wire n23804;
	wire n23805;
	wire n23806;
	wire n23808;
	wire n23809;
	wire n23810;
	wire n23811;
	wire n23812;
	wire n23813;
	wire n23814;
	wire n23815;
	wire n23816;
	wire n23817;
	wire n23818;
	wire n23819;
	wire n23820;
	wire n23821;
	wire n23822;
	wire n23823;
	wire n23824;
	wire n23825;
	wire n23826;
	wire n23827;
	wire n23828;
	wire n23829;
	wire n23830;
	wire n23831;
	wire n23832;
	wire n23833;
	wire n23834;
	wire n23835;
	wire n23836;
	wire n23837;
	wire n23838;
	wire n23839;
	wire n23840;
	wire n23841;
	wire n23842;
	wire n23843;
	wire n23844;
	wire n23845;
	wire n23846;
	wire n23847;
	wire n23848;
	wire n23849;
	wire n23850;
	wire n23851;
	wire n23852;
	wire n23853;
	wire n23854;
	wire n23855;
	wire n23856;
	wire n23857;
	wire n23858;
	wire n23859;
	wire n23860;
	wire n23861;
	wire n23862;
	wire n23863;
	wire n23864;
	wire n23865;
	wire n23866;
	wire n23867;
	wire n23868;
	wire n23869;
	wire n23870;
	wire n23871;
	wire n23872;
	wire n23873;
	wire n23874;
	wire n23875;
	wire n23876;
	wire n23877;
	wire n23878;
	wire n23879;
	wire n23880;
	wire n23881;
	wire n23882;
	wire n23883;
	wire n23884;
	wire n23885;
	wire n23886;
	wire n23887;
	wire n23888;
	wire n23889;
	wire n23890;
	wire n23891;
	wire n23892;
	wire n23893;
	wire n23894;
	wire n23895;
	wire n23896;
	wire n23897;
	wire n23898;
	wire n23899;
	wire n23900;
	wire n23901;
	wire n23902;
	wire n23903;
	wire n23904;
	wire n23905;
	wire n23906;
	wire n23907;
	wire n23908;
	wire n23909;
	wire n23910;
	wire n23911;
	wire n23912;
	wire n23913;
	wire n23914;
	wire n23915;
	wire n23916;
	wire n23917;
	wire n23918;
	wire n23919;
	wire n23920;
	wire n23921;
	wire n23922;
	wire n23923;
	wire n23924;
	wire n23925;
	wire n23926;
	wire n23927;
	wire n23928;
	wire n23929;
	wire n23930;
	wire n23931;
	wire n23932;
	wire n23933;
	wire n23934;
	wire n23935;
	wire n23936;
	wire n23937;
	wire n23938;
	wire n23939;
	wire n23940;
	wire n23941;
	wire n23942;
	wire n23943;
	wire n23944;
	wire n23945;
	wire n23946;
	wire n23947;
	wire n23948;
	wire n23949;
	wire n23950;
	wire n23951;
	wire n23952;
	wire n23953;
	wire n23954;
	wire n23955;
	wire n23956;
	wire n23957;
	wire n23958;
	wire n23959;
	wire n23960;
	wire n23961;
	wire n23962;
	wire n23963;
	wire n23964;
	wire n23965;
	wire n23966;
	wire n23967;
	wire n23968;
	wire n23969;
	wire n23970;
	wire n23971;
	wire n23972;
	wire n23973;
	wire n23974;
	wire n23975;
	wire n23976;
	wire n23977;
	wire n23978;
	wire n23979;
	wire n23980;
	wire n23981;
	wire n23982;
	wire n23983;
	wire n23984;
	wire n23985;
	wire n23986;
	wire n23987;
	wire n23988;
	wire n23989;
	wire n23990;
	wire n23991;
	wire n23992;
	wire n23993;
	wire n23994;
	wire n23995;
	wire n23996;
	wire n23997;
	wire n23998;
	wire n23999;
	wire n24000;
	wire n24001;
	wire n24002;
	wire n24003;
	wire n24004;
	wire n24005;
	wire n24006;
	wire n24007;
	wire n24008;
	wire n24009;
	wire n24010;
	wire n24011;
	wire n24012;
	wire n24013;
	wire n24014;
	wire n24015;
	wire n24016;
	wire n24017;
	wire n24018;
	wire n24019;
	wire n24020;
	wire n24021;
	wire n24022;
	wire n24023;
	wire n24024;
	wire n24025;
	wire n24026;
	wire n24027;
	wire n24028;
	wire n24029;
	wire n24030;
	wire n24031;
	wire n24032;
	wire n24033;
	wire n24034;
	wire n24035;
	wire n24036;
	wire n24037;
	wire n24038;
	wire n24039;
	wire n24040;
	wire n24041;
	wire n24042;
	wire n24043;
	wire n24044;
	wire n24045;
	wire n24046;
	wire n24047;
	wire n24048;
	wire n24049;
	wire n24050;
	wire n24051;
	wire n24052;
	wire n24053;
	wire n24054;
	wire n24055;
	wire n24056;
	wire n24057;
	wire n24058;
	wire n24059;
	wire n24060;
	wire n24061;
	wire n24062;
	wire n24063;
	wire n24064;
	wire n24065;
	wire n24066;
	wire n24067;
	wire n24068;
	wire n24069;
	wire n24070;
	wire n24071;
	wire n24072;
	wire n24073;
	wire n24074;
	wire n24075;
	wire n24076;
	wire n24077;
	wire n24078;
	wire n24079;
	wire n24080;
	wire n24081;
	wire n24082;
	wire n24083;
	wire n24084;
	wire n24085;
	wire n24086;
	wire n24087;
	wire n24088;
	wire n24089;
	wire n24090;
	wire n24091;
	wire n24092;
	wire n24093;
	wire n24094;
	wire n24095;
	wire n24096;
	wire n24097;
	wire n24098;
	wire n24099;
	wire n24100;
	wire n24101;
	wire n24102;
	wire n24103;
	wire n24104;
	wire n24105;
	wire n24106;
	wire n24107;
	wire n24108;
	wire n24109;
	wire n24110;
	wire n24111;
	wire n24112;
	wire n24113;
	wire n24114;
	wire n24115;
	wire n24116;
	wire n24117;
	wire n24118;
	wire n24119;
	wire n24120;
	wire n24121;
	wire n24122;
	wire n24123;
	wire n24124;
	wire n24125;
	wire n24126;
	wire n24127;
	wire n24128;
	wire n24129;
	wire n24130;
	wire n24131;
	wire n24132;
	wire n24133;
	wire n24134;
	wire n24135;
	wire n24136;
	wire n24137;
	wire n24138;
	wire n24139;
	wire n24140;
	wire n24141;
	wire n24142;
	wire n24143;
	wire n24144;
	wire n24145;
	wire n24146;
	wire n24147;
	wire n24148;
	wire n24149;
	wire n24150;
	wire n24151;
	wire n24152;
	wire n24153;
	wire n24154;
	wire n24155;
	wire n24156;
	wire n24157;
	wire n24158;
	wire n24159;
	wire n24160;
	wire n24161;
	wire n24162;
	wire n24163;
	wire n24164;
	wire n24165;
	wire n24166;
	wire n24167;
	wire n24168;
	wire n24169;
	wire n24170;
	wire n24171;
	wire n24172;
	wire n24173;
	wire n24174;
	wire n24175;
	wire n24176;
	wire n24177;
	wire n24178;
	wire n24179;
	wire n24180;
	wire n24181;
	wire n24182;
	wire n24183;
	wire n24184;
	wire n24185;
	wire n24186;
	wire n24187;
	wire n24188;
	wire n24189;
	wire n24190;
	wire n24191;
	wire n24192;
	wire n24193;
	wire n24194;
	wire n24195;
	wire n24196;
	wire n24197;
	wire n24198;
	wire n24199;
	wire n24200;
	wire n24201;
	wire n24202;
	wire n24203;
	wire n24204;
	wire n24205;
	wire n24206;
	wire n24207;
	wire n24208;
	wire n24209;
	wire n24210;
	wire n24211;
	wire n24212;
	wire n24213;
	wire n24214;
	wire n24215;
	wire n24216;
	wire n24217;
	wire n24218;
	wire n24219;
	wire n24220;
	wire n24221;
	wire n24222;
	wire n24223;
	wire n24224;
	wire n24225;
	wire n24226;
	wire n24227;
	wire n24228;
	wire n24229;
	wire n24230;
	wire n24231;
	wire n24232;
	wire n24233;
	wire n24234;
	wire n24235;
	wire n24236;
	wire n24237;
	wire n24238;
	wire n24239;
	wire n24240;
	wire n24241;
	wire n24242;
	wire n24243;
	wire n24244;
	wire n24245;
	wire n24246;
	wire n24247;
	wire n24248;
	wire n24249;
	wire n24250;
	wire n24251;
	wire n24252;
	wire n24253;
	wire n24254;
	wire n24255;
	wire n24256;
	wire n24257;
	wire n24258;
	wire n24259;
	wire n24260;
	wire n24261;
	wire n24262;
	wire n24263;
	wire n24264;
	wire n24265;
	wire n24266;
	wire n24267;
	wire n24268;
	wire n24269;
	wire n24270;
	wire n24271;
	wire n24272;
	wire n24273;
	wire n24274;
	wire n24275;
	wire n24276;
	wire n24277;
	wire n24278;
	wire n24279;
	wire n24280;
	wire n24281;
	wire n24282;
	wire n24283;
	wire n24284;
	wire n24285;
	wire n24286;
	wire n24287;
	wire n24288;
	wire n24289;
	wire n24290;
	wire n24291;
	wire n24292;
	wire n24293;
	wire n24294;
	wire n24295;
	wire n24296;
	wire n24297;
	wire n24298;
	wire n24299;
	wire n24300;
	wire n24301;
	wire n24302;
	wire n24303;
	wire n24304;
	wire n24305;
	wire n24306;
	wire n24307;
	wire n24308;
	wire n24309;
	wire n24310;
	wire n24311;
	wire n24312;
	wire n24313;
	wire n24314;
	wire n24315;
	wire n24316;
	wire n24317;
	wire n24318;
	wire n24319;
	wire n24320;
	wire n24321;
	wire n24322;
	wire n24323;
	wire n24324;
	wire n24325;
	wire n24326;
	wire n24327;
	wire n24328;
	wire n24329;
	wire n24330;
	wire n24331;
	wire n24332;
	wire n24333;
	wire n24334;
	wire n24335;
	wire n24336;
	wire n24337;
	wire n24338;
	wire n24339;
	wire n24340;
	wire n24341;
	wire n24342;
	wire n24343;
	wire n24344;
	wire n24345;
	wire n24346;
	wire n24347;
	wire n24348;
	wire n24349;
	wire n24350;
	wire n24351;
	wire n24352;
	wire n24353;
	wire n24354;
	wire n24355;
	wire n24356;
	wire n24357;
	wire n24358;
	wire n24359;
	wire n24360;
	wire n24361;
	wire n24362;
	wire n24363;
	wire n24364;
	wire n24365;
	wire n24366;
	wire n24367;
	wire n24368;
	wire n24369;
	wire n24370;
	wire n24371;
	wire n24372;
	wire n24373;
	wire n24374;
	wire n24375;
	wire n24376;
	wire n24377;
	wire n24378;
	wire n24379;
	wire n24380;
	wire n24381;
	wire n24382;
	wire n24383;
	wire n24384;
	wire n24385;
	wire n24386;
	wire n24387;
	wire n24388;
	wire n24389;
	wire n24390;
	wire n24391;
	wire n24392;
	wire n24393;
	wire n24394;
	wire n24395;
	wire n24396;
	wire n24397;
	wire n24398;
	wire n24399;
	wire n24400;
	wire n24401;
	wire n24402;
	wire n24403;
	wire n24404;
	wire n24405;
	wire n24406;
	wire n24407;
	wire n24408;
	wire n24409;
	wire n24410;
	wire n24411;
	wire n24412;
	wire n24413;
	wire n24414;
	wire n24415;
	wire n24416;
	wire n24417;
	wire n24418;
	wire n24419;
	wire n24420;
	wire n24421;
	wire n24422;
	wire n24423;
	wire n24424;
	wire n24425;
	wire n24426;
	wire n24427;
	wire n24428;
	wire n24429;
	wire n24430;
	wire n24431;
	wire n24432;
	wire n24433;
	wire n24434;
	wire n24435;
	wire n24436;
	wire n24437;
	wire n24438;
	wire n24439;
	wire n24440;
	wire n24441;
	wire n24442;
	wire n24443;
	wire n24444;
	wire n24445;
	wire n24446;
	wire n24447;
	wire n24448;
	wire n24449;
	wire n24450;
	wire n24451;
	wire n24452;
	wire n24453;
	wire n24454;
	wire n24455;
	wire n24456;
	wire n24457;
	wire n24458;
	wire n24459;
	wire n24460;
	wire n24461;
	wire n24462;
	wire n24463;
	wire n24464;
	wire n24465;
	wire n24466;
	wire n24467;
	wire n24468;
	wire n24469;
	wire n24470;
	wire n24471;
	wire n24472;
	wire n24473;
	wire n24474;
	wire n24475;
	wire n24476;
	wire n24477;
	wire n24478;
	wire n24479;
	wire n24480;
	wire n24481;
	wire n24482;
	wire n24483;
	wire n24484;
	wire n24485;
	wire n24486;
	wire n24487;
	wire n24488;
	wire n24489;
	wire n24490;
	wire n24491;
	wire n24492;
	wire n24493;
	wire n24494;
	wire n24495;
	wire n24496;
	wire n24497;
	wire n24498;
	wire n24499;
	wire n24500;
	wire n24501;
	wire n24502;
	wire n24503;
	wire n24504;
	wire n24505;
	wire n24506;
	wire n24507;
	wire n24508;
	wire n24509;
	wire n24510;
	wire n24511;
	wire n24512;
	wire n24513;
	wire n24514;
	wire n24515;
	wire n24516;
	wire n24517;
	wire n24518;
	wire n24519;
	wire n24520;
	wire n24521;
	wire n24522;
	wire n24523;
	wire n24524;
	wire n24525;
	wire n24526;
	wire n24527;
	wire n24528;
	wire n24529;
	wire n24530;
	wire n24531;
	wire n24532;
	wire n24533;
	wire n24534;
	wire n24535;
	wire n24536;
	wire n24537;
	wire n24538;
	wire n24539;
	wire n24540;
	wire n24541;
	wire n24542;
	wire n24543;
	wire n24544;
	wire n24545;
	wire n24546;
	wire n24547;
	wire n24548;
	wire n24549;
	wire n24550;
	wire n24551;
	wire n24552;
	wire n24553;
	wire n24554;
	wire n24555;
	wire n24556;
	wire n24557;
	wire n24558;
	wire n24559;
	wire n24560;
	wire n24561;
	wire n24562;
	wire n24563;
	wire n24564;
	wire n24565;
	wire n24566;
	wire n24567;
	wire n24568;
	wire n24569;
	wire n24570;
	wire n24571;
	wire n24572;
	wire n24573;
	wire n24574;
	wire n24575;
	wire n24576;
	wire n24577;
	wire n24578;
	wire n24579;
	wire n24580;
	wire n24581;
	wire n24582;
	wire n24583;
	wire n24584;
	wire n24585;
	wire n24586;
	wire n24587;
	wire n24588;
	wire n24589;
	wire n24590;
	wire n24591;
	wire n24592;
	wire n24593;
	wire n24594;
	wire n24595;
	wire n24596;
	wire n24597;
	wire n24598;
	wire n24599;
	wire n24600;
	wire n24601;
	wire n24602;
	wire n24603;
	wire n24604;
	wire n24605;
	wire n24606;
	wire n24607;
	wire n24608;
	wire n24609;
	wire n24610;
	wire n24611;
	wire n24612;
	wire n24613;
	wire n24614;
	wire n24615;
	wire n24616;
	wire n24617;
	wire n24618;
	wire n24619;
	wire n24620;
	wire n24621;
	wire n24622;
	wire n24623;
	wire n24624;
	wire n24625;
	wire n24626;
	wire n24627;
	wire n24628;
	wire n24629;
	wire n24630;
	wire n24631;
	wire n24632;
	wire n24633;
	wire n24634;
	wire n24635;
	wire n24636;
	wire n24637;
	wire n24638;
	wire n24639;
	wire n24640;
	wire n24641;
	wire n24642;
	wire n24643;
	wire n24644;
	wire n24645;
	wire n24646;
	wire n24647;
	wire n24648;
	wire n24649;
	wire n24650;
	wire n24651;
	wire n24652;
	wire n24653;
	wire n24654;
	wire n24655;
	wire n24656;
	wire n24657;
	wire n24658;
	wire n24659;
	wire n24660;
	wire n24661;
	wire n24662;
	wire n24663;
	wire n24664;
	wire n24665;
	wire n24666;
	wire n24667;
	wire n24668;
	wire n24669;
	wire n24670;
	wire n24671;
	wire n24672;
	wire n24673;
	wire n24674;
	wire n24675;
	wire n24676;
	wire n24677;
	wire n24678;
	wire n24679;
	wire n24680;
	wire n24681;
	wire n24682;
	wire n24683;
	wire n24684;
	wire n24685;
	wire n24686;
	wire n24687;
	wire n24688;
	wire n24689;
	wire n24690;
	wire n24691;
	wire n24692;
	wire n24693;
	wire n24694;
	wire n24695;
	wire n24696;
	wire n24697;
	wire n24698;
	wire n24699;
	wire n24700;
	wire n24701;
	wire n24702;
	wire n24703;
	wire n24704;
	wire n24705;
	wire n24706;
	wire n24707;
	wire n24708;
	wire n24709;
	wire n24710;
	wire n24711;
	wire n24712;
	wire n24713;
	wire n24714;
	wire n24715;
	wire n24716;
	wire n24717;
	wire n24718;
	wire n24719;
	wire n24720;
	wire n24721;
	wire n24722;
	wire n24723;
	wire n24724;
	wire n24725;
	wire n24726;
	wire n24727;
	wire n24728;
	wire n24729;
	wire n24730;
	wire n24731;
	wire n24732;
	wire n24733;
	wire n24734;
	wire n24735;
	wire n24736;
	wire n24737;
	wire n24738;
	wire n24739;
	wire n24740;
	wire n24741;
	wire n24742;
	wire n24743;
	wire n24744;
	wire n24745;
	wire n24746;
	wire n24747;
	wire n24748;
	wire n24749;
	wire n24750;
	wire n24751;
	wire n24752;
	wire n24753;
	wire n24754;
	wire n24755;
	wire n24756;
	wire n24757;
	wire n24758;
	wire n24759;
	wire n24760;
	wire n24761;
	wire n24762;
	wire n24763;
	wire n24764;
	wire n24765;
	wire n24766;
	wire n24767;
	wire n24768;
	wire n24769;
	wire n24770;
	wire n24771;
	wire n24772;
	wire n24773;
	wire n24774;
	wire n24775;
	wire n24776;
	wire n24777;
	wire n24778;
	wire n24779;
	wire n24780;
	wire n24781;
	wire n24782;
	wire n24783;
	wire n24784;
	wire n24785;
	wire n24786;
	wire n24787;
	wire n24788;
	wire n24789;
	wire n24790;
	wire n24791;
	wire n24792;
	wire n24793;
	wire n24794;
	wire n24795;
	wire n24796;
	wire n24797;
	wire n24798;
	wire n24799;
	wire n24800;
	wire n24801;
	wire n24802;
	wire n24803;
	wire n24804;
	wire n24805;
	wire n24806;
	wire n24807;
	wire n24808;
	wire n24809;
	wire n24810;
	wire n24811;
	wire n24812;
	wire n24813;
	wire n24814;
	wire n24815;
	wire n24816;
	wire n24817;
	wire n24818;
	wire n24819;
	wire n24820;
	wire n24821;
	wire n24822;
	wire n24823;
	wire n24824;
	wire n24825;
	wire n24826;
	wire n24827;
	wire n24828;
	wire n24829;
	wire n24830;
	wire n24831;
	wire n24832;
	wire n24833;
	wire n24834;
	wire n24835;
	wire n24836;
	wire n24837;
	wire n24838;
	wire n24839;
	wire n24840;
	wire n24841;
	wire n24842;
	wire n24843;
	wire n24844;
	wire n24845;
	wire n24846;
	wire n24848;
	wire n24849;
	wire n24850;
	wire n24851;
	wire n24852;
	wire n24853;
	wire n24854;
	wire n24855;
	wire n24856;
	wire n24857;
	wire n24858;
	wire n24859;
	wire n24860;
	wire n24861;
	wire n24862;
	wire n24863;
	wire n24864;
	wire n24865;
	wire n24866;
	wire n24867;
	wire n24868;
	wire n24869;
	wire n24870;
	wire n24871;
	wire n24872;
	wire n24873;
	wire n24874;
	wire n24875;
	wire n24876;
	wire n24877;
	wire n24878;
	wire n24879;
	wire n24880;
	wire n24881;
	wire n24882;
	wire n24883;
	wire n24884;
	wire n24885;
	wire n24886;
	wire n24887;
	wire n24888;
	wire n24889;
	wire n24890;
	wire n24891;
	wire n24892;
	wire n24893;
	wire n24894;
	wire n24895;
	wire n24896;
	wire n24897;
	wire n24898;
	wire n24899;
	wire n24900;
	wire n24901;
	wire n24902;
	wire n24903;
	wire n24904;
	wire n24905;
	wire n24906;
	wire n24907;
	wire n24908;
	wire n24909;
	wire n24910;
	wire n24911;
	wire n24912;
	wire n24913;
	wire n24914;
	wire n24915;
	wire n24916;
	wire n24917;
	wire n24918;
	wire n24919;
	wire n24920;
	wire n24921;
	wire n24922;
	wire n24923;
	wire n24924;
	wire n24925;
	wire n24926;
	wire n24927;
	wire n24928;
	wire n24929;
	wire n24930;
	wire n24931;
	wire n24932;
	wire n24933;
	wire n24934;
	wire n24935;
	wire n24936;
	wire n24937;
	wire n24938;
	wire n24939;
	wire n24940;
	wire n24941;
	wire n24942;
	wire n24943;
	wire n24944;
	wire n24945;
	wire n24946;
	wire n24947;
	wire n24948;
	wire n24949;
	wire n24950;
	wire n24951;
	wire n24952;
	wire n24953;
	wire n24954;
	wire n24955;
	wire n24956;
	wire n24957;
	wire n24958;
	wire n24959;
	wire n24960;
	wire n24961;
	wire n24962;
	wire n24963;
	wire n24964;
	wire n24965;
	wire n24966;
	wire n24967;
	wire n24968;
	wire n24969;
	wire n24970;
	wire n24971;
	wire n24972;
	wire n24973;
	wire n24974;
	wire n24975;
	wire n24976;
	wire n24977;
	wire n24978;
	wire n24979;
	wire n24980;
	wire n24981;
	wire n24982;
	wire n24983;
	wire n24984;
	wire n24985;
	wire n24986;
	wire n24987;
	wire n24988;
	wire n24989;
	wire n24990;
	wire n24991;
	wire n24992;
	wire n24993;
	wire n24994;
	wire n24995;
	wire n24996;
	wire n24997;
	wire n24998;
	wire n24999;
	wire n25000;
	wire n25001;
	wire n25002;
	wire n25003;
	wire n25004;
	wire n25005;
	wire n25006;
	wire n25007;
	wire n25008;
	wire n25009;
	wire n25010;
	wire n25011;
	wire n25012;
	wire n25013;
	wire n25014;
	wire n25015;
	wire n25016;
	wire n25017;
	wire n25018;
	wire n25019;
	wire n25020;
	wire n25021;
	wire n25022;
	wire n25023;
	wire n25024;
	wire n25025;
	wire n25026;
	wire n25027;
	wire n25028;
	wire n25029;
	wire n25030;
	wire n25031;
	wire n25032;
	wire n25033;
	wire n25034;
	wire n25035;
	wire n25036;
	wire n25037;
	wire n25038;
	wire n25039;
	wire n25040;
	wire n25041;
	wire n25042;
	wire n25043;
	wire n25044;
	wire n25045;
	wire n25046;
	wire n25047;
	wire n25048;
	wire n25049;
	wire n25050;
	wire n25051;
	wire n25052;
	wire n25053;
	wire n25054;
	wire n25055;
	wire n25056;
	wire n25057;
	wire n25058;
	wire n25059;
	wire n25060;
	wire n25061;
	wire n25062;
	wire n25063;
	wire n25064;
	wire n25065;
	wire n25066;
	wire n25067;
	wire n25068;
	wire n25069;
	wire n25070;
	wire n25071;
	wire n25072;
	wire n25073;
	wire n25074;
	wire n25075;
	wire n25076;
	wire n25077;
	wire n25078;
	wire n25079;
	wire n25080;
	wire n25081;
	wire n25082;
	wire n25083;
	wire n25084;
	wire n25085;
	wire n25086;
	wire n25087;
	wire n25088;
	wire n25089;
	wire n25090;
	wire n25091;
	wire n25092;
	wire n25093;
	wire n25094;
	wire n25095;
	wire n25096;
	wire n25097;
	wire n25098;
	wire n25099;
	wire n25100;
	wire n25101;
	wire n25102;
	wire n25103;
	wire n25104;
	wire n25105;
	wire n25106;
	wire n25107;
	wire n25108;
	wire n25109;
	wire n25110;
	wire n25111;
	wire n25112;
	wire n25113;
	wire n25114;
	wire n25115;
	wire n25116;
	wire n25117;
	wire n25118;
	wire n25119;
	wire n25120;
	wire n25121;
	wire n25122;
	wire n25123;
	wire n25124;
	wire n25125;
	wire n25126;
	wire n25127;
	wire n25128;
	wire n25129;
	wire n25130;
	wire n25131;
	wire n25132;
	wire n25133;
	wire n25134;
	wire n25135;
	wire n25136;
	wire n25137;
	wire n25138;
	wire n25139;
	wire n25140;
	wire n25141;
	wire n25142;
	wire n25143;
	wire n25144;
	wire n25145;
	wire n25146;
	wire n25147;
	wire n25148;
	wire n25149;
	wire n25150;
	wire n25151;
	wire n25152;
	wire n25153;
	wire n25154;
	wire n25155;
	wire n25156;
	wire n25157;
	wire n25158;
	wire n25159;
	wire n25160;
	wire n25161;
	wire n25162;
	wire n25163;
	wire n25164;
	wire n25165;
	wire n25166;
	wire n25167;
	wire n25168;
	wire n25169;
	wire n25170;
	wire n25171;
	wire n25172;
	wire n25173;
	wire n25174;
	wire n25175;
	wire n25176;
	wire n25177;
	wire n25178;
	wire n25179;
	wire n25180;
	wire n25181;
	wire n25182;
	wire n25183;
	wire n25184;
	wire n25185;
	wire n25186;
	wire n25187;
	wire n25188;
	wire n25189;
	wire n25190;
	wire n25191;
	wire n25192;
	wire n25193;
	wire n25194;
	wire n25195;
	wire n25196;
	wire n25197;
	wire n25198;
	wire n25199;
	wire n25200;
	wire n25201;
	wire n25202;
	wire n25203;
	wire n25204;
	wire n25205;
	wire n25206;
	wire n25207;
	wire n25208;
	wire n25209;
	wire n25210;
	wire n25211;
	wire n25212;
	wire n25213;
	wire n25214;
	wire n25215;
	wire n25216;
	wire n25217;
	wire n25218;
	wire n25219;
	wire n25220;
	wire n25221;
	wire n25222;
	wire n25223;
	wire n25224;
	wire n25225;
	wire n25226;
	wire n25227;
	wire n25228;
	wire n25229;
	wire n25230;
	wire n25231;
	wire n25232;
	wire n25233;
	wire n25234;
	wire n25235;
	wire n25236;
	wire n25237;
	wire n25238;
	wire n25239;
	wire n25240;
	wire n25241;
	wire n25242;
	wire n25243;
	wire n25244;
	wire n25245;
	wire n25246;
	wire n25247;
	wire n25248;
	wire n25249;
	wire n25250;
	wire n25251;
	wire n25252;
	wire n25253;
	wire n25254;
	wire n25255;
	wire n25256;
	wire n25257;
	wire n25258;
	wire n25259;
	wire n25260;
	wire n25261;
	wire n25262;
	wire n25263;
	wire n25264;
	wire n25265;
	wire n25266;
	wire n25267;
	wire n25268;
	wire n25269;
	wire n25270;
	wire n25271;
	wire n25272;
	wire n25273;
	wire n25274;
	wire n25275;
	wire n25276;
	wire n25277;
	wire n25278;
	wire n25279;
	wire n25280;
	wire n25281;
	wire n25282;
	wire n25283;
	wire n25284;
	wire n25285;
	wire n25286;
	wire n25287;
	wire n25288;
	wire n25289;
	wire n25290;
	wire n25291;
	wire n25292;
	wire n25293;
	wire n25294;
	wire n25295;
	wire n25296;
	wire n25297;
	wire n25298;
	wire n25299;
	wire n25300;
	wire [2:0] w_a2_0;
	wire [1:0] w_a2_1;
	wire [1:0] w_a3_0;
	wire [2:0] w_a4_0;
	wire [1:0] w_a4_1;
	wire [1:0] w_a5_0;
	wire [2:0] w_a6_0;
	wire [1:0] w_a7_0;
	wire [2:0] w_a8_0;
	wire [1:0] w_a9_0;
	wire [2:0] w_a10_0;
	wire [1:0] w_a11_0;
	wire [2:0] w_a12_0;
	wire [1:0] w_a13_0;
	wire [2:0] w_a14_0;
	wire [1:0] w_a14_1;
	wire [1:0] w_a15_0;
	wire [2:0] w_a16_0;
	wire [1:0] w_a17_0;
	wire [2:0] w_a18_0;
	wire [1:0] w_a18_1;
	wire [1:0] w_a19_0;
	wire [2:0] w_a20_0;
	wire [1:0] w_a21_0;
	wire [2:0] w_a22_0;
	wire [1:0] w_a22_1;
	wire [1:0] w_a23_0;
	wire [2:0] w_a24_0;
	wire [1:0] w_a25_0;
	wire [2:0] w_a26_0;
	wire [1:0] w_a26_1;
	wire [1:0] w_a27_0;
	wire [2:0] w_a28_0;
	wire [1:0] w_a29_0;
	wire [2:0] w_a30_0;
	wire [1:0] w_a30_1;
	wire [1:0] w_a31_0;
	wire [2:0] w_a32_0;
	wire [1:0] w_a33_0;
	wire [2:0] w_a34_0;
	wire [1:0] w_a34_1;
	wire [1:0] w_a35_0;
	wire [2:0] w_a36_0;
	wire [1:0] w_a37_0;
	wire [2:0] w_a38_0;
	wire [1:0] w_a39_0;
	wire [2:0] w_a40_0;
	wire [1:0] w_a41_0;
	wire [2:0] w_a42_0;
	wire [1:0] w_a42_1;
	wire [1:0] w_a43_0;
	wire [2:0] w_a44_0;
	wire [1:0] w_a45_0;
	wire [2:0] w_a46_0;
	wire [1:0] w_a46_1;
	wire [1:0] w_a47_0;
	wire [2:0] w_a48_0;
	wire [1:0] w_a49_0;
	wire [2:0] w_a50_0;
	wire [1:0] w_a51_0;
	wire [2:0] w_a52_0;
	wire [1:0] w_a53_0;
	wire [2:0] w_a54_0;
	wire [1:0] w_a54_1;
	wire [1:0] w_a55_0;
	wire [2:0] w_a56_0;
	wire [1:0] w_a57_0;
	wire [2:0] w_a58_0;
	wire [1:0] w_a59_0;
	wire [2:0] w_a60_0;
	wire [1:0] w_a61_0;
	wire [2:0] w_a62_0;
	wire [1:0] w_a63_0;
	wire [2:0] w_a64_0;
	wire [1:0] w_a65_0;
	wire [2:0] w_a66_0;
	wire [1:0] w_a66_1;
	wire [1:0] w_a67_0;
	wire [2:0] w_a68_0;
	wire [1:0] w_a69_0;
	wire [2:0] w_a70_0;
	wire [1:0] w_a70_1;
	wire [1:0] w_a71_0;
	wire [2:0] w_a72_0;
	wire [1:0] w_a73_0;
	wire [2:0] w_a74_0;
	wire [1:0] w_a74_1;
	wire [1:0] w_a75_0;
	wire [2:0] w_a76_0;
	wire [1:0] w_a77_0;
	wire [2:0] w_a78_0;
	wire [1:0] w_a78_1;
	wire [1:0] w_a79_0;
	wire [2:0] w_a80_0;
	wire [1:0] w_a81_0;
	wire [2:0] w_a82_0;
	wire [1:0] w_a82_1;
	wire [1:0] w_a83_0;
	wire [2:0] w_a84_0;
	wire [1:0] w_a85_0;
	wire [2:0] w_a86_0;
	wire [1:0] w_a86_1;
	wire [1:0] w_a87_0;
	wire [2:0] w_a88_0;
	wire [1:0] w_a89_0;
	wire [2:0] w_a90_0;
	wire [1:0] w_a90_1;
	wire [1:0] w_a91_0;
	wire [2:0] w_a92_0;
	wire [1:0] w_a93_0;
	wire [2:0] w_a94_0;
	wire [1:0] w_a94_1;
	wire [1:0] w_a95_0;
	wire [2:0] w_a96_0;
	wire [1:0] w_a97_0;
	wire [2:0] w_a98_0;
	wire [1:0] w_a98_1;
	wire [1:0] w_a99_0;
	wire [2:0] w_a100_0;
	wire [1:0] w_a101_0;
	wire [2:0] w_a102_0;
	wire [1:0] w_a102_1;
	wire [1:0] w_a103_0;
	wire [2:0] w_a104_0;
	wire [1:0] w_a105_0;
	wire [2:0] w_a106_0;
	wire [1:0] w_a106_1;
	wire [1:0] w_a107_0;
	wire [2:0] w_a108_0;
	wire [1:0] w_a109_0;
	wire [2:0] w_a110_0;
	wire [1:0] w_a110_1;
	wire [1:0] w_a111_0;
	wire [2:0] w_a112_0;
	wire [1:0] w_a113_0;
	wire [2:0] w_a114_0;
	wire [1:0] w_a114_1;
	wire [1:0] w_a115_0;
	wire [2:0] w_a116_0;
	wire [1:0] w_a117_0;
	wire [2:0] w_a118_0;
	wire [1:0] w_a118_1;
	wire [1:0] w_a119_0;
	wire [2:0] w_a120_0;
	wire [1:0] w_a121_0;
	wire [2:0] w_a122_0;
	wire [1:0] w_a123_0;
	wire [2:0] w_a124_0;
	wire [1:0] w_a124_1;
	wire [2:0] w_a125_0;
	wire [2:0] w_a126_0;
	wire [1:0] w_a126_1;
	wire [1:0] w_a127_0;
	wire [2:0] w_asqrt1_0;
	wire w_asqrt1_1;
	wire asqrt_fa_1;
	wire [2:0] w_asqrt2_0;
	wire [2:0] w_asqrt2_1;
	wire [2:0] w_asqrt2_2;
	wire [2:0] w_asqrt2_3;
	wire [2:0] w_asqrt2_4;
	wire [2:0] w_asqrt2_5;
	wire [2:0] w_asqrt2_6;
	wire [2:0] w_asqrt2_7;
	wire [2:0] w_asqrt2_8;
	wire [2:0] w_asqrt2_9;
	wire [2:0] w_asqrt2_10;
	wire [2:0] w_asqrt2_11;
	wire [2:0] w_asqrt2_12;
	wire [2:0] w_asqrt2_13;
	wire [2:0] w_asqrt2_14;
	wire [2:0] w_asqrt2_15;
	wire [2:0] w_asqrt2_16;
	wire [2:0] w_asqrt2_17;
	wire [2:0] w_asqrt2_18;
	wire [2:0] w_asqrt2_19;
	wire [2:0] w_asqrt2_20;
	wire [2:0] w_asqrt2_21;
	wire [2:0] w_asqrt2_22;
	wire [2:0] w_asqrt2_23;
	wire [2:0] w_asqrt2_24;
	wire [2:0] w_asqrt2_25;
	wire [2:0] w_asqrt2_26;
	wire [2:0] w_asqrt2_27;
	wire [2:0] w_asqrt2_28;
	wire [2:0] w_asqrt2_29;
	wire [2:0] w_asqrt2_30;
	wire [1:0] w_asqrt2_31;
	wire asqrt_fa_2;
	wire [2:0] w_asqrt3_0;
	wire [2:0] w_asqrt3_1;
	wire [1:0] w_asqrt3_2;
	wire asqrt_fa_3;
	wire [2:0] w_asqrt4_0;
	wire [2:0] w_asqrt4_1;
	wire [2:0] w_asqrt4_2;
	wire [2:0] w_asqrt4_3;
	wire [2:0] w_asqrt4_4;
	wire [2:0] w_asqrt4_5;
	wire [2:0] w_asqrt4_6;
	wire [2:0] w_asqrt4_7;
	wire [2:0] w_asqrt4_8;
	wire [2:0] w_asqrt4_9;
	wire [2:0] w_asqrt4_10;
	wire [2:0] w_asqrt4_11;
	wire [2:0] w_asqrt4_12;
	wire [2:0] w_asqrt4_13;
	wire [2:0] w_asqrt4_14;
	wire [2:0] w_asqrt4_15;
	wire [2:0] w_asqrt4_16;
	wire [2:0] w_asqrt4_17;
	wire [2:0] w_asqrt4_18;
	wire [2:0] w_asqrt4_19;
	wire [2:0] w_asqrt4_20;
	wire [2:0] w_asqrt4_21;
	wire [2:0] w_asqrt4_22;
	wire [2:0] w_asqrt4_23;
	wire [2:0] w_asqrt4_24;
	wire [2:0] w_asqrt4_25;
	wire [2:0] w_asqrt4_26;
	wire [2:0] w_asqrt4_27;
	wire [2:0] w_asqrt4_28;
	wire [2:0] w_asqrt4_29;
	wire [2:0] w_asqrt4_30;
	wire [1:0] w_asqrt4_31;
	wire asqrt_fa_4;
	wire [2:0] w_asqrt5_0;
	wire [2:0] w_asqrt5_1;
	wire [2:0] w_asqrt5_2;
	wire [2:0] w_asqrt5_3;
	wire [1:0] w_asqrt5_4;
	wire asqrt_fa_5;
	wire [2:0] w_asqrt6_0;
	wire [2:0] w_asqrt6_1;
	wire [2:0] w_asqrt6_2;
	wire [2:0] w_asqrt6_3;
	wire [2:0] w_asqrt6_4;
	wire [2:0] w_asqrt6_5;
	wire [2:0] w_asqrt6_6;
	wire [2:0] w_asqrt6_7;
	wire [2:0] w_asqrt6_8;
	wire [2:0] w_asqrt6_9;
	wire [2:0] w_asqrt6_10;
	wire [2:0] w_asqrt6_11;
	wire [2:0] w_asqrt6_12;
	wire [2:0] w_asqrt6_13;
	wire [2:0] w_asqrt6_14;
	wire [2:0] w_asqrt6_15;
	wire [2:0] w_asqrt6_16;
	wire [2:0] w_asqrt6_17;
	wire [2:0] w_asqrt6_18;
	wire [2:0] w_asqrt6_19;
	wire [2:0] w_asqrt6_20;
	wire [2:0] w_asqrt6_21;
	wire [2:0] w_asqrt6_22;
	wire [2:0] w_asqrt6_23;
	wire [2:0] w_asqrt6_24;
	wire [2:0] w_asqrt6_25;
	wire [2:0] w_asqrt6_26;
	wire [2:0] w_asqrt6_27;
	wire [2:0] w_asqrt6_28;
	wire [2:0] w_asqrt6_29;
	wire [2:0] w_asqrt6_30;
	wire [2:0] w_asqrt6_31;
	wire w_asqrt6_32;
	wire asqrt_fa_6;
	wire [2:0] w_asqrt7_0;
	wire [2:0] w_asqrt7_1;
	wire [2:0] w_asqrt7_2;
	wire [2:0] w_asqrt7_3;
	wire [2:0] w_asqrt7_4;
	wire [2:0] w_asqrt7_5;
	wire w_asqrt7_6;
	wire asqrt_fa_7;
	wire [2:0] w_asqrt8_0;
	wire [2:0] w_asqrt8_1;
	wire [2:0] w_asqrt8_2;
	wire [2:0] w_asqrt8_3;
	wire [2:0] w_asqrt8_4;
	wire [2:0] w_asqrt8_5;
	wire [2:0] w_asqrt8_6;
	wire [2:0] w_asqrt8_7;
	wire [2:0] w_asqrt8_8;
	wire [2:0] w_asqrt8_9;
	wire [2:0] w_asqrt8_10;
	wire [2:0] w_asqrt8_11;
	wire [2:0] w_asqrt8_12;
	wire [2:0] w_asqrt8_13;
	wire [2:0] w_asqrt8_14;
	wire [2:0] w_asqrt8_15;
	wire [2:0] w_asqrt8_16;
	wire [2:0] w_asqrt8_17;
	wire [2:0] w_asqrt8_18;
	wire [2:0] w_asqrt8_19;
	wire [2:0] w_asqrt8_20;
	wire [2:0] w_asqrt8_21;
	wire [2:0] w_asqrt8_22;
	wire [2:0] w_asqrt8_23;
	wire [2:0] w_asqrt8_24;
	wire [2:0] w_asqrt8_25;
	wire [2:0] w_asqrt8_26;
	wire [2:0] w_asqrt8_27;
	wire [2:0] w_asqrt8_28;
	wire [2:0] w_asqrt8_29;
	wire [2:0] w_asqrt8_30;
	wire [2:0] w_asqrt8_31;
	wire [1:0] w_asqrt8_32;
	wire asqrt_fa_8;
	wire [2:0] w_asqrt9_0;
	wire [2:0] w_asqrt9_1;
	wire [2:0] w_asqrt9_2;
	wire [2:0] w_asqrt9_3;
	wire [2:0] w_asqrt9_4;
	wire [2:0] w_asqrt9_5;
	wire [2:0] w_asqrt9_6;
	wire [2:0] w_asqrt9_7;
	wire w_asqrt9_8;
	wire asqrt_fa_9;
	wire [2:0] w_asqrt10_0;
	wire [2:0] w_asqrt10_1;
	wire [2:0] w_asqrt10_2;
	wire [2:0] w_asqrt10_3;
	wire [2:0] w_asqrt10_4;
	wire [2:0] w_asqrt10_5;
	wire [2:0] w_asqrt10_6;
	wire [2:0] w_asqrt10_7;
	wire [2:0] w_asqrt10_8;
	wire [2:0] w_asqrt10_9;
	wire [2:0] w_asqrt10_10;
	wire [2:0] w_asqrt10_11;
	wire [2:0] w_asqrt10_12;
	wire [2:0] w_asqrt10_13;
	wire [2:0] w_asqrt10_14;
	wire [2:0] w_asqrt10_15;
	wire [2:0] w_asqrt10_16;
	wire [2:0] w_asqrt10_17;
	wire [2:0] w_asqrt10_18;
	wire [2:0] w_asqrt10_19;
	wire [2:0] w_asqrt10_20;
	wire [2:0] w_asqrt10_21;
	wire [2:0] w_asqrt10_22;
	wire [2:0] w_asqrt10_23;
	wire [2:0] w_asqrt10_24;
	wire [2:0] w_asqrt10_25;
	wire [2:0] w_asqrt10_26;
	wire [2:0] w_asqrt10_27;
	wire [2:0] w_asqrt10_28;
	wire [2:0] w_asqrt10_29;
	wire [2:0] w_asqrt10_30;
	wire [2:0] w_asqrt10_31;
	wire [1:0] w_asqrt10_32;
	wire asqrt_fa_10;
	wire [2:0] w_asqrt11_0;
	wire [2:0] w_asqrt11_1;
	wire [2:0] w_asqrt11_2;
	wire [2:0] w_asqrt11_3;
	wire [2:0] w_asqrt11_4;
	wire [2:0] w_asqrt11_5;
	wire [2:0] w_asqrt11_6;
	wire [2:0] w_asqrt11_7;
	wire [1:0] w_asqrt11_8;
	wire asqrt_fa_11;
	wire [2:0] w_asqrt12_0;
	wire [2:0] w_asqrt12_1;
	wire [2:0] w_asqrt12_2;
	wire [2:0] w_asqrt12_3;
	wire [2:0] w_asqrt12_4;
	wire [2:0] w_asqrt12_5;
	wire [2:0] w_asqrt12_6;
	wire [2:0] w_asqrt12_7;
	wire [2:0] w_asqrt12_8;
	wire [2:0] w_asqrt12_9;
	wire [2:0] w_asqrt12_10;
	wire [2:0] w_asqrt12_11;
	wire [2:0] w_asqrt12_12;
	wire [2:0] w_asqrt12_13;
	wire [2:0] w_asqrt12_14;
	wire [2:0] w_asqrt12_15;
	wire [2:0] w_asqrt12_16;
	wire [2:0] w_asqrt12_17;
	wire [2:0] w_asqrt12_18;
	wire [2:0] w_asqrt12_19;
	wire [2:0] w_asqrt12_20;
	wire [2:0] w_asqrt12_21;
	wire [2:0] w_asqrt12_22;
	wire [2:0] w_asqrt12_23;
	wire [2:0] w_asqrt12_24;
	wire [2:0] w_asqrt12_25;
	wire [2:0] w_asqrt12_26;
	wire [2:0] w_asqrt12_27;
	wire [2:0] w_asqrt12_28;
	wire [2:0] w_asqrt12_29;
	wire [2:0] w_asqrt12_30;
	wire [2:0] w_asqrt12_31;
	wire [2:0] w_asqrt12_32;
	wire w_asqrt12_33;
	wire asqrt_fa_12;
	wire [2:0] w_asqrt13_0;
	wire [2:0] w_asqrt13_1;
	wire [2:0] w_asqrt13_2;
	wire [2:0] w_asqrt13_3;
	wire [2:0] w_asqrt13_4;
	wire [2:0] w_asqrt13_5;
	wire [2:0] w_asqrt13_6;
	wire [2:0] w_asqrt13_7;
	wire [2:0] w_asqrt13_8;
	wire [2:0] w_asqrt13_9;
	wire [1:0] w_asqrt13_10;
	wire asqrt_fa_13;
	wire [2:0] w_asqrt14_0;
	wire [2:0] w_asqrt14_1;
	wire [2:0] w_asqrt14_2;
	wire [2:0] w_asqrt14_3;
	wire [2:0] w_asqrt14_4;
	wire [2:0] w_asqrt14_5;
	wire [2:0] w_asqrt14_6;
	wire [2:0] w_asqrt14_7;
	wire [2:0] w_asqrt14_8;
	wire [2:0] w_asqrt14_9;
	wire [2:0] w_asqrt14_10;
	wire [2:0] w_asqrt14_11;
	wire [2:0] w_asqrt14_12;
	wire [2:0] w_asqrt14_13;
	wire [2:0] w_asqrt14_14;
	wire [2:0] w_asqrt14_15;
	wire [2:0] w_asqrt14_16;
	wire [2:0] w_asqrt14_17;
	wire [2:0] w_asqrt14_18;
	wire [2:0] w_asqrt14_19;
	wire [2:0] w_asqrt14_20;
	wire [2:0] w_asqrt14_21;
	wire [2:0] w_asqrt14_22;
	wire [2:0] w_asqrt14_23;
	wire [2:0] w_asqrt14_24;
	wire [2:0] w_asqrt14_25;
	wire [2:0] w_asqrt14_26;
	wire [2:0] w_asqrt14_27;
	wire [2:0] w_asqrt14_28;
	wire [2:0] w_asqrt14_29;
	wire [2:0] w_asqrt14_30;
	wire [2:0] w_asqrt14_31;
	wire [2:0] w_asqrt14_32;
	wire [2:0] w_asqrt14_33;
	wire w_asqrt14_34;
	wire asqrt_fa_14;
	wire [2:0] w_asqrt15_0;
	wire [2:0] w_asqrt15_1;
	wire [2:0] w_asqrt15_2;
	wire [2:0] w_asqrt15_3;
	wire [2:0] w_asqrt15_4;
	wire [2:0] w_asqrt15_5;
	wire [2:0] w_asqrt15_6;
	wire [2:0] w_asqrt15_7;
	wire [2:0] w_asqrt15_8;
	wire [2:0] w_asqrt15_9;
	wire [2:0] w_asqrt15_10;
	wire [2:0] w_asqrt15_11;
	wire w_asqrt15_12;
	wire asqrt_fa_15;
	wire [2:0] w_asqrt16_0;
	wire [2:0] w_asqrt16_1;
	wire [2:0] w_asqrt16_2;
	wire [2:0] w_asqrt16_3;
	wire [2:0] w_asqrt16_4;
	wire [2:0] w_asqrt16_5;
	wire [2:0] w_asqrt16_6;
	wire [2:0] w_asqrt16_7;
	wire [2:0] w_asqrt16_8;
	wire [2:0] w_asqrt16_9;
	wire [2:0] w_asqrt16_10;
	wire [2:0] w_asqrt16_11;
	wire [2:0] w_asqrt16_12;
	wire [2:0] w_asqrt16_13;
	wire [2:0] w_asqrt16_14;
	wire [2:0] w_asqrt16_15;
	wire [2:0] w_asqrt16_16;
	wire [2:0] w_asqrt16_17;
	wire [2:0] w_asqrt16_18;
	wire [2:0] w_asqrt16_19;
	wire [2:0] w_asqrt16_20;
	wire [2:0] w_asqrt16_21;
	wire [2:0] w_asqrt16_22;
	wire [2:0] w_asqrt16_23;
	wire [2:0] w_asqrt16_24;
	wire [2:0] w_asqrt16_25;
	wire [2:0] w_asqrt16_26;
	wire [2:0] w_asqrt16_27;
	wire [2:0] w_asqrt16_28;
	wire [2:0] w_asqrt16_29;
	wire [2:0] w_asqrt16_30;
	wire [2:0] w_asqrt16_31;
	wire [2:0] w_asqrt16_32;
	wire [2:0] w_asqrt16_33;
	wire [1:0] w_asqrt16_34;
	wire asqrt_fa_16;
	wire [2:0] w_asqrt17_0;
	wire [2:0] w_asqrt17_1;
	wire [2:0] w_asqrt17_2;
	wire [2:0] w_asqrt17_3;
	wire [2:0] w_asqrt17_4;
	wire [2:0] w_asqrt17_5;
	wire [2:0] w_asqrt17_6;
	wire [2:0] w_asqrt17_7;
	wire [2:0] w_asqrt17_8;
	wire [2:0] w_asqrt17_9;
	wire [2:0] w_asqrt17_10;
	wire [2:0] w_asqrt17_11;
	wire [2:0] w_asqrt17_12;
	wire [1:0] w_asqrt17_13;
	wire asqrt_fa_17;
	wire [2:0] w_asqrt18_0;
	wire [2:0] w_asqrt18_1;
	wire [2:0] w_asqrt18_2;
	wire [2:0] w_asqrt18_3;
	wire [2:0] w_asqrt18_4;
	wire [2:0] w_asqrt18_5;
	wire [2:0] w_asqrt18_6;
	wire [2:0] w_asqrt18_7;
	wire [2:0] w_asqrt18_8;
	wire [2:0] w_asqrt18_9;
	wire [2:0] w_asqrt18_10;
	wire [2:0] w_asqrt18_11;
	wire [2:0] w_asqrt18_12;
	wire [2:0] w_asqrt18_13;
	wire [2:0] w_asqrt18_14;
	wire [2:0] w_asqrt18_15;
	wire [2:0] w_asqrt18_16;
	wire [2:0] w_asqrt18_17;
	wire [2:0] w_asqrt18_18;
	wire [2:0] w_asqrt18_19;
	wire [2:0] w_asqrt18_20;
	wire [2:0] w_asqrt18_21;
	wire [2:0] w_asqrt18_22;
	wire [2:0] w_asqrt18_23;
	wire [2:0] w_asqrt18_24;
	wire [2:0] w_asqrt18_25;
	wire [2:0] w_asqrt18_26;
	wire [2:0] w_asqrt18_27;
	wire [2:0] w_asqrt18_28;
	wire [2:0] w_asqrt18_29;
	wire [2:0] w_asqrt18_30;
	wire [2:0] w_asqrt18_31;
	wire [2:0] w_asqrt18_32;
	wire [2:0] w_asqrt18_33;
	wire [2:0] w_asqrt18_34;
	wire w_asqrt18_35;
	wire asqrt_fa_18;
	wire [2:0] w_asqrt19_0;
	wire [2:0] w_asqrt19_1;
	wire [2:0] w_asqrt19_2;
	wire [2:0] w_asqrt19_3;
	wire [2:0] w_asqrt19_4;
	wire [2:0] w_asqrt19_5;
	wire [2:0] w_asqrt19_6;
	wire [2:0] w_asqrt19_7;
	wire [2:0] w_asqrt19_8;
	wire [2:0] w_asqrt19_9;
	wire [2:0] w_asqrt19_10;
	wire [2:0] w_asqrt19_11;
	wire [2:0] w_asqrt19_12;
	wire [2:0] w_asqrt19_13;
	wire w_asqrt19_14;
	wire asqrt_fa_19;
	wire [2:0] w_asqrt20_0;
	wire [2:0] w_asqrt20_1;
	wire [2:0] w_asqrt20_2;
	wire [2:0] w_asqrt20_3;
	wire [2:0] w_asqrt20_4;
	wire [2:0] w_asqrt20_5;
	wire [2:0] w_asqrt20_6;
	wire [2:0] w_asqrt20_7;
	wire [2:0] w_asqrt20_8;
	wire [2:0] w_asqrt20_9;
	wire [2:0] w_asqrt20_10;
	wire [2:0] w_asqrt20_11;
	wire [2:0] w_asqrt20_12;
	wire [2:0] w_asqrt20_13;
	wire [2:0] w_asqrt20_14;
	wire [2:0] w_asqrt20_15;
	wire [2:0] w_asqrt20_16;
	wire [2:0] w_asqrt20_17;
	wire [2:0] w_asqrt20_18;
	wire [2:0] w_asqrt20_19;
	wire [2:0] w_asqrt20_20;
	wire [2:0] w_asqrt20_21;
	wire [2:0] w_asqrt20_22;
	wire [2:0] w_asqrt20_23;
	wire [2:0] w_asqrt20_24;
	wire [2:0] w_asqrt20_25;
	wire [2:0] w_asqrt20_26;
	wire [2:0] w_asqrt20_27;
	wire [2:0] w_asqrt20_28;
	wire [2:0] w_asqrt20_29;
	wire [2:0] w_asqrt20_30;
	wire [2:0] w_asqrt20_31;
	wire [2:0] w_asqrt20_32;
	wire [2:0] w_asqrt20_33;
	wire [2:0] w_asqrt20_34;
	wire w_asqrt20_35;
	wire asqrt_fa_20;
	wire [2:0] w_asqrt21_0;
	wire [2:0] w_asqrt21_1;
	wire [2:0] w_asqrt21_2;
	wire [2:0] w_asqrt21_3;
	wire [2:0] w_asqrt21_4;
	wire [2:0] w_asqrt21_5;
	wire [2:0] w_asqrt21_6;
	wire [2:0] w_asqrt21_7;
	wire [2:0] w_asqrt21_8;
	wire [2:0] w_asqrt21_9;
	wire [2:0] w_asqrt21_10;
	wire [2:0] w_asqrt21_11;
	wire [2:0] w_asqrt21_12;
	wire [2:0] w_asqrt21_13;
	wire [2:0] w_asqrt21_14;
	wire [2:0] w_asqrt21_15;
	wire w_asqrt21_16;
	wire asqrt_fa_21;
	wire [2:0] w_asqrt22_0;
	wire [2:0] w_asqrt22_1;
	wire [2:0] w_asqrt22_2;
	wire [2:0] w_asqrt22_3;
	wire [2:0] w_asqrt22_4;
	wire [2:0] w_asqrt22_5;
	wire [2:0] w_asqrt22_6;
	wire [2:0] w_asqrt22_7;
	wire [2:0] w_asqrt22_8;
	wire [2:0] w_asqrt22_9;
	wire [2:0] w_asqrt22_10;
	wire [2:0] w_asqrt22_11;
	wire [2:0] w_asqrt22_12;
	wire [2:0] w_asqrt22_13;
	wire [2:0] w_asqrt22_14;
	wire [2:0] w_asqrt22_15;
	wire [2:0] w_asqrt22_16;
	wire [2:0] w_asqrt22_17;
	wire [2:0] w_asqrt22_18;
	wire [2:0] w_asqrt22_19;
	wire [2:0] w_asqrt22_20;
	wire [2:0] w_asqrt22_21;
	wire [2:0] w_asqrt22_22;
	wire [2:0] w_asqrt22_23;
	wire [2:0] w_asqrt22_24;
	wire [2:0] w_asqrt22_25;
	wire [2:0] w_asqrt22_26;
	wire [2:0] w_asqrt22_27;
	wire [2:0] w_asqrt22_28;
	wire [2:0] w_asqrt22_29;
	wire [2:0] w_asqrt22_30;
	wire [2:0] w_asqrt22_31;
	wire [2:0] w_asqrt22_32;
	wire [2:0] w_asqrt22_33;
	wire [2:0] w_asqrt22_34;
	wire [2:0] w_asqrt22_35;
	wire w_asqrt22_36;
	wire asqrt_fa_22;
	wire [2:0] w_asqrt23_0;
	wire [2:0] w_asqrt23_1;
	wire [2:0] w_asqrt23_2;
	wire [2:0] w_asqrt23_3;
	wire [2:0] w_asqrt23_4;
	wire [2:0] w_asqrt23_5;
	wire [2:0] w_asqrt23_6;
	wire [2:0] w_asqrt23_7;
	wire [2:0] w_asqrt23_8;
	wire [2:0] w_asqrt23_9;
	wire [2:0] w_asqrt23_10;
	wire [2:0] w_asqrt23_11;
	wire [2:0] w_asqrt23_12;
	wire [2:0] w_asqrt23_13;
	wire [2:0] w_asqrt23_14;
	wire [2:0] w_asqrt23_15;
	wire [2:0] w_asqrt23_16;
	wire [2:0] w_asqrt23_17;
	wire w_asqrt23_18;
	wire asqrt_fa_23;
	wire [2:0] w_asqrt24_0;
	wire [2:0] w_asqrt24_1;
	wire [2:0] w_asqrt24_2;
	wire [2:0] w_asqrt24_3;
	wire [2:0] w_asqrt24_4;
	wire [2:0] w_asqrt24_5;
	wire [2:0] w_asqrt24_6;
	wire [2:0] w_asqrt24_7;
	wire [2:0] w_asqrt24_8;
	wire [2:0] w_asqrt24_9;
	wire [2:0] w_asqrt24_10;
	wire [2:0] w_asqrt24_11;
	wire [2:0] w_asqrt24_12;
	wire [2:0] w_asqrt24_13;
	wire [2:0] w_asqrt24_14;
	wire [2:0] w_asqrt24_15;
	wire [2:0] w_asqrt24_16;
	wire [2:0] w_asqrt24_17;
	wire [2:0] w_asqrt24_18;
	wire [2:0] w_asqrt24_19;
	wire [2:0] w_asqrt24_20;
	wire [2:0] w_asqrt24_21;
	wire [2:0] w_asqrt24_22;
	wire [2:0] w_asqrt24_23;
	wire [2:0] w_asqrt24_24;
	wire [2:0] w_asqrt24_25;
	wire [2:0] w_asqrt24_26;
	wire [2:0] w_asqrt24_27;
	wire [2:0] w_asqrt24_28;
	wire [2:0] w_asqrt24_29;
	wire [2:0] w_asqrt24_30;
	wire [2:0] w_asqrt24_31;
	wire [2:0] w_asqrt24_32;
	wire [2:0] w_asqrt24_33;
	wire [2:0] w_asqrt24_34;
	wire [2:0] w_asqrt24_35;
	wire [1:0] w_asqrt24_36;
	wire asqrt_fa_24;
	wire [2:0] w_asqrt25_0;
	wire [2:0] w_asqrt25_1;
	wire [2:0] w_asqrt25_2;
	wire [2:0] w_asqrt25_3;
	wire [2:0] w_asqrt25_4;
	wire [2:0] w_asqrt25_5;
	wire [2:0] w_asqrt25_6;
	wire [2:0] w_asqrt25_7;
	wire [2:0] w_asqrt25_8;
	wire [2:0] w_asqrt25_9;
	wire [2:0] w_asqrt25_10;
	wire [2:0] w_asqrt25_11;
	wire [2:0] w_asqrt25_12;
	wire [2:0] w_asqrt25_13;
	wire [2:0] w_asqrt25_14;
	wire [2:0] w_asqrt25_15;
	wire [2:0] w_asqrt25_16;
	wire [2:0] w_asqrt25_17;
	wire [1:0] w_asqrt25_18;
	wire asqrt_fa_25;
	wire [2:0] w_asqrt26_0;
	wire [2:0] w_asqrt26_1;
	wire [2:0] w_asqrt26_2;
	wire [2:0] w_asqrt26_3;
	wire [2:0] w_asqrt26_4;
	wire [2:0] w_asqrt26_5;
	wire [2:0] w_asqrt26_6;
	wire [2:0] w_asqrt26_7;
	wire [2:0] w_asqrt26_8;
	wire [2:0] w_asqrt26_9;
	wire [2:0] w_asqrt26_10;
	wire [2:0] w_asqrt26_11;
	wire [2:0] w_asqrt26_12;
	wire [2:0] w_asqrt26_13;
	wire [2:0] w_asqrt26_14;
	wire [2:0] w_asqrt26_15;
	wire [2:0] w_asqrt26_16;
	wire [2:0] w_asqrt26_17;
	wire [2:0] w_asqrt26_18;
	wire [2:0] w_asqrt26_19;
	wire [2:0] w_asqrt26_20;
	wire [2:0] w_asqrt26_21;
	wire [2:0] w_asqrt26_22;
	wire [2:0] w_asqrt26_23;
	wire [2:0] w_asqrt26_24;
	wire [2:0] w_asqrt26_25;
	wire [2:0] w_asqrt26_26;
	wire [2:0] w_asqrt26_27;
	wire [2:0] w_asqrt26_28;
	wire [2:0] w_asqrt26_29;
	wire [2:0] w_asqrt26_30;
	wire [2:0] w_asqrt26_31;
	wire [2:0] w_asqrt26_32;
	wire [2:0] w_asqrt26_33;
	wire [2:0] w_asqrt26_34;
	wire [2:0] w_asqrt26_35;
	wire [1:0] w_asqrt26_36;
	wire asqrt_fa_26;
	wire [2:0] w_asqrt27_0;
	wire [2:0] w_asqrt27_1;
	wire [2:0] w_asqrt27_2;
	wire [2:0] w_asqrt27_3;
	wire [2:0] w_asqrt27_4;
	wire [2:0] w_asqrt27_5;
	wire [2:0] w_asqrt27_6;
	wire [2:0] w_asqrt27_7;
	wire [2:0] w_asqrt27_8;
	wire [2:0] w_asqrt27_9;
	wire [2:0] w_asqrt27_10;
	wire [2:0] w_asqrt27_11;
	wire [2:0] w_asqrt27_12;
	wire [2:0] w_asqrt27_13;
	wire [2:0] w_asqrt27_14;
	wire [2:0] w_asqrt27_15;
	wire [2:0] w_asqrt27_16;
	wire [2:0] w_asqrt27_17;
	wire [2:0] w_asqrt27_18;
	wire [2:0] w_asqrt27_19;
	wire [1:0] w_asqrt27_20;
	wire asqrt_fa_27;
	wire [2:0] w_asqrt28_0;
	wire [2:0] w_asqrt28_1;
	wire [2:0] w_asqrt28_2;
	wire [2:0] w_asqrt28_3;
	wire [2:0] w_asqrt28_4;
	wire [2:0] w_asqrt28_5;
	wire [2:0] w_asqrt28_6;
	wire [2:0] w_asqrt28_7;
	wire [2:0] w_asqrt28_8;
	wire [2:0] w_asqrt28_9;
	wire [2:0] w_asqrt28_10;
	wire [2:0] w_asqrt28_11;
	wire [2:0] w_asqrt28_12;
	wire [2:0] w_asqrt28_13;
	wire [2:0] w_asqrt28_14;
	wire [2:0] w_asqrt28_15;
	wire [2:0] w_asqrt28_16;
	wire [2:0] w_asqrt28_17;
	wire [2:0] w_asqrt28_18;
	wire [2:0] w_asqrt28_19;
	wire [2:0] w_asqrt28_20;
	wire [2:0] w_asqrt28_21;
	wire [2:0] w_asqrt28_22;
	wire [2:0] w_asqrt28_23;
	wire [2:0] w_asqrt28_24;
	wire [2:0] w_asqrt28_25;
	wire [2:0] w_asqrt28_26;
	wire [2:0] w_asqrt28_27;
	wire [2:0] w_asqrt28_28;
	wire [2:0] w_asqrt28_29;
	wire [2:0] w_asqrt28_30;
	wire [2:0] w_asqrt28_31;
	wire [2:0] w_asqrt28_32;
	wire [2:0] w_asqrt28_33;
	wire [2:0] w_asqrt28_34;
	wire [2:0] w_asqrt28_35;
	wire [2:0] w_asqrt28_36;
	wire [1:0] w_asqrt28_37;
	wire asqrt_fa_28;
	wire [2:0] w_asqrt29_0;
	wire [2:0] w_asqrt29_1;
	wire [2:0] w_asqrt29_2;
	wire [2:0] w_asqrt29_3;
	wire [2:0] w_asqrt29_4;
	wire [2:0] w_asqrt29_5;
	wire [2:0] w_asqrt29_6;
	wire [2:0] w_asqrt29_7;
	wire [2:0] w_asqrt29_8;
	wire [2:0] w_asqrt29_9;
	wire [2:0] w_asqrt29_10;
	wire [2:0] w_asqrt29_11;
	wire [2:0] w_asqrt29_12;
	wire [2:0] w_asqrt29_13;
	wire [2:0] w_asqrt29_14;
	wire [2:0] w_asqrt29_15;
	wire [2:0] w_asqrt29_16;
	wire [2:0] w_asqrt29_17;
	wire [2:0] w_asqrt29_18;
	wire [2:0] w_asqrt29_19;
	wire [2:0] w_asqrt29_20;
	wire [1:0] w_asqrt29_21;
	wire asqrt_fa_29;
	wire [2:0] w_asqrt30_0;
	wire [2:0] w_asqrt30_1;
	wire [2:0] w_asqrt30_2;
	wire [2:0] w_asqrt30_3;
	wire [2:0] w_asqrt30_4;
	wire [2:0] w_asqrt30_5;
	wire [2:0] w_asqrt30_6;
	wire [2:0] w_asqrt30_7;
	wire [2:0] w_asqrt30_8;
	wire [2:0] w_asqrt30_9;
	wire [2:0] w_asqrt30_10;
	wire [2:0] w_asqrt30_11;
	wire [2:0] w_asqrt30_12;
	wire [2:0] w_asqrt30_13;
	wire [2:0] w_asqrt30_14;
	wire [2:0] w_asqrt30_15;
	wire [2:0] w_asqrt30_16;
	wire [2:0] w_asqrt30_17;
	wire [2:0] w_asqrt30_18;
	wire [2:0] w_asqrt30_19;
	wire [2:0] w_asqrt30_20;
	wire [2:0] w_asqrt30_21;
	wire [2:0] w_asqrt30_22;
	wire [2:0] w_asqrt30_23;
	wire [2:0] w_asqrt30_24;
	wire [2:0] w_asqrt30_25;
	wire [2:0] w_asqrt30_26;
	wire [2:0] w_asqrt30_27;
	wire [2:0] w_asqrt30_28;
	wire [2:0] w_asqrt30_29;
	wire [2:0] w_asqrt30_30;
	wire [2:0] w_asqrt30_31;
	wire [2:0] w_asqrt30_32;
	wire [2:0] w_asqrt30_33;
	wire [2:0] w_asqrt30_34;
	wire [2:0] w_asqrt30_35;
	wire [2:0] w_asqrt30_36;
	wire [2:0] w_asqrt30_37;
	wire w_asqrt30_38;
	wire asqrt_fa_30;
	wire [2:0] w_asqrt31_0;
	wire [2:0] w_asqrt31_1;
	wire [2:0] w_asqrt31_2;
	wire [2:0] w_asqrt31_3;
	wire [2:0] w_asqrt31_4;
	wire [2:0] w_asqrt31_5;
	wire [2:0] w_asqrt31_6;
	wire [2:0] w_asqrt31_7;
	wire [2:0] w_asqrt31_8;
	wire [2:0] w_asqrt31_9;
	wire [2:0] w_asqrt31_10;
	wire [2:0] w_asqrt31_11;
	wire [2:0] w_asqrt31_12;
	wire [2:0] w_asqrt31_13;
	wire [2:0] w_asqrt31_14;
	wire [2:0] w_asqrt31_15;
	wire [2:0] w_asqrt31_16;
	wire [2:0] w_asqrt31_17;
	wire [2:0] w_asqrt31_18;
	wire [2:0] w_asqrt31_19;
	wire [2:0] w_asqrt31_20;
	wire [2:0] w_asqrt31_21;
	wire [2:0] w_asqrt31_22;
	wire w_asqrt31_23;
	wire asqrt_fa_31;
	wire [2:0] w_asqrt32_0;
	wire [2:0] w_asqrt32_1;
	wire [2:0] w_asqrt32_2;
	wire [2:0] w_asqrt32_3;
	wire [2:0] w_asqrt32_4;
	wire [2:0] w_asqrt32_5;
	wire [2:0] w_asqrt32_6;
	wire [2:0] w_asqrt32_7;
	wire [2:0] w_asqrt32_8;
	wire [2:0] w_asqrt32_9;
	wire [2:0] w_asqrt32_10;
	wire [2:0] w_asqrt32_11;
	wire [2:0] w_asqrt32_12;
	wire [2:0] w_asqrt32_13;
	wire [2:0] w_asqrt32_14;
	wire [2:0] w_asqrt32_15;
	wire [2:0] w_asqrt32_16;
	wire [2:0] w_asqrt32_17;
	wire [2:0] w_asqrt32_18;
	wire [2:0] w_asqrt32_19;
	wire [2:0] w_asqrt32_20;
	wire [2:0] w_asqrt32_21;
	wire [2:0] w_asqrt32_22;
	wire [2:0] w_asqrt32_23;
	wire [2:0] w_asqrt32_24;
	wire [2:0] w_asqrt32_25;
	wire [2:0] w_asqrt32_26;
	wire [2:0] w_asqrt32_27;
	wire [2:0] w_asqrt32_28;
	wire [2:0] w_asqrt32_29;
	wire [2:0] w_asqrt32_30;
	wire [2:0] w_asqrt32_31;
	wire [2:0] w_asqrt32_32;
	wire [2:0] w_asqrt32_33;
	wire [2:0] w_asqrt32_34;
	wire [2:0] w_asqrt32_35;
	wire [2:0] w_asqrt32_36;
	wire [2:0] w_asqrt32_37;
	wire [1:0] w_asqrt32_38;
	wire asqrt_fa_32;
	wire [2:0] w_asqrt33_0;
	wire [2:0] w_asqrt33_1;
	wire [2:0] w_asqrt33_2;
	wire [2:0] w_asqrt33_3;
	wire [2:0] w_asqrt33_4;
	wire [2:0] w_asqrt33_5;
	wire [2:0] w_asqrt33_6;
	wire [2:0] w_asqrt33_7;
	wire [2:0] w_asqrt33_8;
	wire [2:0] w_asqrt33_9;
	wire [2:0] w_asqrt33_10;
	wire [2:0] w_asqrt33_11;
	wire [2:0] w_asqrt33_12;
	wire [2:0] w_asqrt33_13;
	wire [2:0] w_asqrt33_14;
	wire [2:0] w_asqrt33_15;
	wire [2:0] w_asqrt33_16;
	wire [2:0] w_asqrt33_17;
	wire [2:0] w_asqrt33_18;
	wire [2:0] w_asqrt33_19;
	wire [2:0] w_asqrt33_20;
	wire [2:0] w_asqrt33_21;
	wire [2:0] w_asqrt33_22;
	wire [2:0] w_asqrt33_23;
	wire [2:0] w_asqrt33_24;
	wire w_asqrt33_25;
	wire asqrt_fa_33;
	wire [2:0] w_asqrt34_0;
	wire [2:0] w_asqrt34_1;
	wire [2:0] w_asqrt34_2;
	wire [2:0] w_asqrt34_3;
	wire [2:0] w_asqrt34_4;
	wire [2:0] w_asqrt34_5;
	wire [2:0] w_asqrt34_6;
	wire [2:0] w_asqrt34_7;
	wire [2:0] w_asqrt34_8;
	wire [2:0] w_asqrt34_9;
	wire [2:0] w_asqrt34_10;
	wire [2:0] w_asqrt34_11;
	wire [2:0] w_asqrt34_12;
	wire [2:0] w_asqrt34_13;
	wire [2:0] w_asqrt34_14;
	wire [2:0] w_asqrt34_15;
	wire [2:0] w_asqrt34_16;
	wire [2:0] w_asqrt34_17;
	wire [2:0] w_asqrt34_18;
	wire [2:0] w_asqrt34_19;
	wire [2:0] w_asqrt34_20;
	wire [2:0] w_asqrt34_21;
	wire [2:0] w_asqrt34_22;
	wire [2:0] w_asqrt34_23;
	wire [2:0] w_asqrt34_24;
	wire [2:0] w_asqrt34_25;
	wire [2:0] w_asqrt34_26;
	wire [2:0] w_asqrt34_27;
	wire [2:0] w_asqrt34_28;
	wire [2:0] w_asqrt34_29;
	wire [2:0] w_asqrt34_30;
	wire [2:0] w_asqrt34_31;
	wire [2:0] w_asqrt34_32;
	wire [2:0] w_asqrt34_33;
	wire [2:0] w_asqrt34_34;
	wire [2:0] w_asqrt34_35;
	wire [2:0] w_asqrt34_36;
	wire [2:0] w_asqrt34_37;
	wire [2:0] w_asqrt34_38;
	wire w_asqrt34_39;
	wire asqrt_fa_34;
	wire [2:0] w_asqrt35_0;
	wire [2:0] w_asqrt35_1;
	wire [2:0] w_asqrt35_2;
	wire [2:0] w_asqrt35_3;
	wire [2:0] w_asqrt35_4;
	wire [2:0] w_asqrt35_5;
	wire [2:0] w_asqrt35_6;
	wire [2:0] w_asqrt35_7;
	wire [2:0] w_asqrt35_8;
	wire [2:0] w_asqrt35_9;
	wire [2:0] w_asqrt35_10;
	wire [2:0] w_asqrt35_11;
	wire [2:0] w_asqrt35_12;
	wire [2:0] w_asqrt35_13;
	wire [2:0] w_asqrt35_14;
	wire [2:0] w_asqrt35_15;
	wire [2:0] w_asqrt35_16;
	wire [2:0] w_asqrt35_17;
	wire [2:0] w_asqrt35_18;
	wire [2:0] w_asqrt35_19;
	wire [2:0] w_asqrt35_20;
	wire [2:0] w_asqrt35_21;
	wire [2:0] w_asqrt35_22;
	wire [2:0] w_asqrt35_23;
	wire [2:0] w_asqrt35_24;
	wire [2:0] w_asqrt35_25;
	wire [2:0] w_asqrt35_26;
	wire w_asqrt35_27;
	wire asqrt_fa_35;
	wire [2:0] w_asqrt36_0;
	wire [2:0] w_asqrt36_1;
	wire [2:0] w_asqrt36_2;
	wire [2:0] w_asqrt36_3;
	wire [2:0] w_asqrt36_4;
	wire [2:0] w_asqrt36_5;
	wire [2:0] w_asqrt36_6;
	wire [2:0] w_asqrt36_7;
	wire [2:0] w_asqrt36_8;
	wire [2:0] w_asqrt36_9;
	wire [2:0] w_asqrt36_10;
	wire [2:0] w_asqrt36_11;
	wire [2:0] w_asqrt36_12;
	wire [2:0] w_asqrt36_13;
	wire [2:0] w_asqrt36_14;
	wire [2:0] w_asqrt36_15;
	wire [2:0] w_asqrt36_16;
	wire [2:0] w_asqrt36_17;
	wire [2:0] w_asqrt36_18;
	wire [2:0] w_asqrt36_19;
	wire [2:0] w_asqrt36_20;
	wire [2:0] w_asqrt36_21;
	wire [2:0] w_asqrt36_22;
	wire [2:0] w_asqrt36_23;
	wire [2:0] w_asqrt36_24;
	wire [2:0] w_asqrt36_25;
	wire [2:0] w_asqrt36_26;
	wire [2:0] w_asqrt36_27;
	wire [2:0] w_asqrt36_28;
	wire [2:0] w_asqrt36_29;
	wire [2:0] w_asqrt36_30;
	wire [2:0] w_asqrt36_31;
	wire [2:0] w_asqrt36_32;
	wire [2:0] w_asqrt36_33;
	wire [2:0] w_asqrt36_34;
	wire [2:0] w_asqrt36_35;
	wire [2:0] w_asqrt36_36;
	wire [2:0] w_asqrt36_37;
	wire [2:0] w_asqrt36_38;
	wire w_asqrt36_39;
	wire asqrt_fa_36;
	wire [2:0] w_asqrt37_0;
	wire [2:0] w_asqrt37_1;
	wire [2:0] w_asqrt37_2;
	wire [2:0] w_asqrt37_3;
	wire [2:0] w_asqrt37_4;
	wire [2:0] w_asqrt37_5;
	wire [2:0] w_asqrt37_6;
	wire [2:0] w_asqrt37_7;
	wire [2:0] w_asqrt37_8;
	wire [2:0] w_asqrt37_9;
	wire [2:0] w_asqrt37_10;
	wire [2:0] w_asqrt37_11;
	wire [2:0] w_asqrt37_12;
	wire [2:0] w_asqrt37_13;
	wire [2:0] w_asqrt37_14;
	wire [2:0] w_asqrt37_15;
	wire [2:0] w_asqrt37_16;
	wire [2:0] w_asqrt37_17;
	wire [2:0] w_asqrt37_18;
	wire [2:0] w_asqrt37_19;
	wire [2:0] w_asqrt37_20;
	wire [2:0] w_asqrt37_21;
	wire [2:0] w_asqrt37_22;
	wire [2:0] w_asqrt37_23;
	wire [2:0] w_asqrt37_24;
	wire [2:0] w_asqrt37_25;
	wire [2:0] w_asqrt37_26;
	wire [2:0] w_asqrt37_27;
	wire w_asqrt37_28;
	wire asqrt_fa_37;
	wire [2:0] w_asqrt38_0;
	wire [2:0] w_asqrt38_1;
	wire [2:0] w_asqrt38_2;
	wire [2:0] w_asqrt38_3;
	wire [2:0] w_asqrt38_4;
	wire [2:0] w_asqrt38_5;
	wire [2:0] w_asqrt38_6;
	wire [2:0] w_asqrt38_7;
	wire [2:0] w_asqrt38_8;
	wire [2:0] w_asqrt38_9;
	wire [2:0] w_asqrt38_10;
	wire [2:0] w_asqrt38_11;
	wire [2:0] w_asqrt38_12;
	wire [2:0] w_asqrt38_13;
	wire [2:0] w_asqrt38_14;
	wire [2:0] w_asqrt38_15;
	wire [2:0] w_asqrt38_16;
	wire [2:0] w_asqrt38_17;
	wire [2:0] w_asqrt38_18;
	wire [2:0] w_asqrt38_19;
	wire [2:0] w_asqrt38_20;
	wire [2:0] w_asqrt38_21;
	wire [2:0] w_asqrt38_22;
	wire [2:0] w_asqrt38_23;
	wire [2:0] w_asqrt38_24;
	wire [2:0] w_asqrt38_25;
	wire [2:0] w_asqrt38_26;
	wire [2:0] w_asqrt38_27;
	wire [2:0] w_asqrt38_28;
	wire [2:0] w_asqrt38_29;
	wire [2:0] w_asqrt38_30;
	wire [2:0] w_asqrt38_31;
	wire [2:0] w_asqrt38_32;
	wire [2:0] w_asqrt38_33;
	wire [2:0] w_asqrt38_34;
	wire [2:0] w_asqrt38_35;
	wire [2:0] w_asqrt38_36;
	wire [2:0] w_asqrt38_37;
	wire [2:0] w_asqrt38_38;
	wire [2:0] w_asqrt38_39;
	wire w_asqrt38_40;
	wire asqrt_fa_38;
	wire [2:0] w_asqrt39_0;
	wire [2:0] w_asqrt39_1;
	wire [2:0] w_asqrt39_2;
	wire [2:0] w_asqrt39_3;
	wire [2:0] w_asqrt39_4;
	wire [2:0] w_asqrt39_5;
	wire [2:0] w_asqrt39_6;
	wire [2:0] w_asqrt39_7;
	wire [2:0] w_asqrt39_8;
	wire [2:0] w_asqrt39_9;
	wire [2:0] w_asqrt39_10;
	wire [2:0] w_asqrt39_11;
	wire [2:0] w_asqrt39_12;
	wire [2:0] w_asqrt39_13;
	wire [2:0] w_asqrt39_14;
	wire [2:0] w_asqrt39_15;
	wire [2:0] w_asqrt39_16;
	wire [2:0] w_asqrt39_17;
	wire [2:0] w_asqrt39_18;
	wire [2:0] w_asqrt39_19;
	wire [2:0] w_asqrt39_20;
	wire [2:0] w_asqrt39_21;
	wire [2:0] w_asqrt39_22;
	wire [2:0] w_asqrt39_23;
	wire [2:0] w_asqrt39_24;
	wire [2:0] w_asqrt39_25;
	wire [2:0] w_asqrt39_26;
	wire [2:0] w_asqrt39_27;
	wire [2:0] w_asqrt39_28;
	wire [2:0] w_asqrt39_29;
	wire w_asqrt39_30;
	wire asqrt_fa_39;
	wire [2:0] w_asqrt40_0;
	wire [2:0] w_asqrt40_1;
	wire [2:0] w_asqrt40_2;
	wire [2:0] w_asqrt40_3;
	wire [2:0] w_asqrt40_4;
	wire [2:0] w_asqrt40_5;
	wire [2:0] w_asqrt40_6;
	wire [2:0] w_asqrt40_7;
	wire [2:0] w_asqrt40_8;
	wire [2:0] w_asqrt40_9;
	wire [2:0] w_asqrt40_10;
	wire [2:0] w_asqrt40_11;
	wire [2:0] w_asqrt40_12;
	wire [2:0] w_asqrt40_13;
	wire [2:0] w_asqrt40_14;
	wire [2:0] w_asqrt40_15;
	wire [2:0] w_asqrt40_16;
	wire [2:0] w_asqrt40_17;
	wire [2:0] w_asqrt40_18;
	wire [2:0] w_asqrt40_19;
	wire [2:0] w_asqrt40_20;
	wire [2:0] w_asqrt40_21;
	wire [2:0] w_asqrt40_22;
	wire [2:0] w_asqrt40_23;
	wire [2:0] w_asqrt40_24;
	wire [2:0] w_asqrt40_25;
	wire [2:0] w_asqrt40_26;
	wire [2:0] w_asqrt40_27;
	wire [2:0] w_asqrt40_28;
	wire [2:0] w_asqrt40_29;
	wire [2:0] w_asqrt40_30;
	wire [2:0] w_asqrt40_31;
	wire [2:0] w_asqrt40_32;
	wire [2:0] w_asqrt40_33;
	wire [2:0] w_asqrt40_34;
	wire [2:0] w_asqrt40_35;
	wire [2:0] w_asqrt40_36;
	wire [2:0] w_asqrt40_37;
	wire [2:0] w_asqrt40_38;
	wire [2:0] w_asqrt40_39;
	wire [1:0] w_asqrt40_40;
	wire asqrt_fa_40;
	wire [2:0] w_asqrt41_0;
	wire [2:0] w_asqrt41_1;
	wire [2:0] w_asqrt41_2;
	wire [2:0] w_asqrt41_3;
	wire [2:0] w_asqrt41_4;
	wire [2:0] w_asqrt41_5;
	wire [2:0] w_asqrt41_6;
	wire [2:0] w_asqrt41_7;
	wire [2:0] w_asqrt41_8;
	wire [2:0] w_asqrt41_9;
	wire [2:0] w_asqrt41_10;
	wire [2:0] w_asqrt41_11;
	wire [2:0] w_asqrt41_12;
	wire [2:0] w_asqrt41_13;
	wire [2:0] w_asqrt41_14;
	wire [2:0] w_asqrt41_15;
	wire [2:0] w_asqrt41_16;
	wire [2:0] w_asqrt41_17;
	wire [2:0] w_asqrt41_18;
	wire [2:0] w_asqrt41_19;
	wire [2:0] w_asqrt41_20;
	wire [2:0] w_asqrt41_21;
	wire [2:0] w_asqrt41_22;
	wire [2:0] w_asqrt41_23;
	wire [2:0] w_asqrt41_24;
	wire [2:0] w_asqrt41_25;
	wire [2:0] w_asqrt41_26;
	wire [2:0] w_asqrt41_27;
	wire [2:0] w_asqrt41_28;
	wire [2:0] w_asqrt41_29;
	wire [2:0] w_asqrt41_30;
	wire w_asqrt41_31;
	wire asqrt_fa_41;
	wire [2:0] w_asqrt42_0;
	wire [2:0] w_asqrt42_1;
	wire [2:0] w_asqrt42_2;
	wire [2:0] w_asqrt42_3;
	wire [2:0] w_asqrt42_4;
	wire [2:0] w_asqrt42_5;
	wire [2:0] w_asqrt42_6;
	wire [2:0] w_asqrt42_7;
	wire [2:0] w_asqrt42_8;
	wire [2:0] w_asqrt42_9;
	wire [2:0] w_asqrt42_10;
	wire [2:0] w_asqrt42_11;
	wire [2:0] w_asqrt42_12;
	wire [2:0] w_asqrt42_13;
	wire [2:0] w_asqrt42_14;
	wire [2:0] w_asqrt42_15;
	wire [2:0] w_asqrt42_16;
	wire [2:0] w_asqrt42_17;
	wire [2:0] w_asqrt42_18;
	wire [2:0] w_asqrt42_19;
	wire [2:0] w_asqrt42_20;
	wire [2:0] w_asqrt42_21;
	wire [2:0] w_asqrt42_22;
	wire [2:0] w_asqrt42_23;
	wire [2:0] w_asqrt42_24;
	wire [2:0] w_asqrt42_25;
	wire [2:0] w_asqrt42_26;
	wire [2:0] w_asqrt42_27;
	wire [2:0] w_asqrt42_28;
	wire [2:0] w_asqrt42_29;
	wire [2:0] w_asqrt42_30;
	wire [2:0] w_asqrt42_31;
	wire [2:0] w_asqrt42_32;
	wire [2:0] w_asqrt42_33;
	wire [2:0] w_asqrt42_34;
	wire [2:0] w_asqrt42_35;
	wire [2:0] w_asqrt42_36;
	wire [2:0] w_asqrt42_37;
	wire [2:0] w_asqrt42_38;
	wire [2:0] w_asqrt42_39;
	wire [2:0] w_asqrt42_40;
	wire w_asqrt42_41;
	wire asqrt_fa_42;
	wire [2:0] w_asqrt43_0;
	wire [2:0] w_asqrt43_1;
	wire [2:0] w_asqrt43_2;
	wire [2:0] w_asqrt43_3;
	wire [2:0] w_asqrt43_4;
	wire [2:0] w_asqrt43_5;
	wire [2:0] w_asqrt43_6;
	wire [2:0] w_asqrt43_7;
	wire [2:0] w_asqrt43_8;
	wire [2:0] w_asqrt43_9;
	wire [2:0] w_asqrt43_10;
	wire [2:0] w_asqrt43_11;
	wire [2:0] w_asqrt43_12;
	wire [2:0] w_asqrt43_13;
	wire [2:0] w_asqrt43_14;
	wire [2:0] w_asqrt43_15;
	wire [2:0] w_asqrt43_16;
	wire [2:0] w_asqrt43_17;
	wire [2:0] w_asqrt43_18;
	wire [2:0] w_asqrt43_19;
	wire [2:0] w_asqrt43_20;
	wire [2:0] w_asqrt43_21;
	wire [2:0] w_asqrt43_22;
	wire [2:0] w_asqrt43_23;
	wire [2:0] w_asqrt43_24;
	wire [2:0] w_asqrt43_25;
	wire [2:0] w_asqrt43_26;
	wire [2:0] w_asqrt43_27;
	wire [2:0] w_asqrt43_28;
	wire [2:0] w_asqrt43_29;
	wire [2:0] w_asqrt43_30;
	wire [2:0] w_asqrt43_31;
	wire [1:0] w_asqrt43_32;
	wire asqrt_fa_43;
	wire [2:0] w_asqrt44_0;
	wire [2:0] w_asqrt44_1;
	wire [2:0] w_asqrt44_2;
	wire [2:0] w_asqrt44_3;
	wire [2:0] w_asqrt44_4;
	wire [2:0] w_asqrt44_5;
	wire [2:0] w_asqrt44_6;
	wire [2:0] w_asqrt44_7;
	wire [2:0] w_asqrt44_8;
	wire [2:0] w_asqrt44_9;
	wire [2:0] w_asqrt44_10;
	wire [2:0] w_asqrt44_11;
	wire [2:0] w_asqrt44_12;
	wire [2:0] w_asqrt44_13;
	wire [2:0] w_asqrt44_14;
	wire [2:0] w_asqrt44_15;
	wire [2:0] w_asqrt44_16;
	wire [2:0] w_asqrt44_17;
	wire [2:0] w_asqrt44_18;
	wire [2:0] w_asqrt44_19;
	wire [2:0] w_asqrt44_20;
	wire [2:0] w_asqrt44_21;
	wire [2:0] w_asqrt44_22;
	wire [2:0] w_asqrt44_23;
	wire [2:0] w_asqrt44_24;
	wire [2:0] w_asqrt44_25;
	wire [2:0] w_asqrt44_26;
	wire [2:0] w_asqrt44_27;
	wire [2:0] w_asqrt44_28;
	wire [2:0] w_asqrt44_29;
	wire [2:0] w_asqrt44_30;
	wire [2:0] w_asqrt44_31;
	wire [2:0] w_asqrt44_32;
	wire [2:0] w_asqrt44_33;
	wire [2:0] w_asqrt44_34;
	wire [2:0] w_asqrt44_35;
	wire [2:0] w_asqrt44_36;
	wire [2:0] w_asqrt44_37;
	wire [2:0] w_asqrt44_38;
	wire [2:0] w_asqrt44_39;
	wire [2:0] w_asqrt44_40;
	wire w_asqrt44_41;
	wire asqrt_fa_44;
	wire [2:0] w_asqrt45_0;
	wire [2:0] w_asqrt45_1;
	wire [2:0] w_asqrt45_2;
	wire [2:0] w_asqrt45_3;
	wire [2:0] w_asqrt45_4;
	wire [2:0] w_asqrt45_5;
	wire [2:0] w_asqrt45_6;
	wire [2:0] w_asqrt45_7;
	wire [2:0] w_asqrt45_8;
	wire [2:0] w_asqrt45_9;
	wire [2:0] w_asqrt45_10;
	wire [2:0] w_asqrt45_11;
	wire [2:0] w_asqrt45_12;
	wire [2:0] w_asqrt45_13;
	wire [2:0] w_asqrt45_14;
	wire [2:0] w_asqrt45_15;
	wire [2:0] w_asqrt45_16;
	wire [2:0] w_asqrt45_17;
	wire [2:0] w_asqrt45_18;
	wire [2:0] w_asqrt45_19;
	wire [2:0] w_asqrt45_20;
	wire [2:0] w_asqrt45_21;
	wire [2:0] w_asqrt45_22;
	wire [2:0] w_asqrt45_23;
	wire [2:0] w_asqrt45_24;
	wire [2:0] w_asqrt45_25;
	wire [2:0] w_asqrt45_26;
	wire [2:0] w_asqrt45_27;
	wire [2:0] w_asqrt45_28;
	wire [2:0] w_asqrt45_29;
	wire [2:0] w_asqrt45_30;
	wire [2:0] w_asqrt45_31;
	wire [2:0] w_asqrt45_32;
	wire [2:0] w_asqrt45_33;
	wire w_asqrt45_34;
	wire asqrt_fa_45;
	wire [2:0] w_asqrt46_0;
	wire [2:0] w_asqrt46_1;
	wire [2:0] w_asqrt46_2;
	wire [2:0] w_asqrt46_3;
	wire [2:0] w_asqrt46_4;
	wire [2:0] w_asqrt46_5;
	wire [2:0] w_asqrt46_6;
	wire [2:0] w_asqrt46_7;
	wire [2:0] w_asqrt46_8;
	wire [2:0] w_asqrt46_9;
	wire [2:0] w_asqrt46_10;
	wire [2:0] w_asqrt46_11;
	wire [2:0] w_asqrt46_12;
	wire [2:0] w_asqrt46_13;
	wire [2:0] w_asqrt46_14;
	wire [2:0] w_asqrt46_15;
	wire [2:0] w_asqrt46_16;
	wire [2:0] w_asqrt46_17;
	wire [2:0] w_asqrt46_18;
	wire [2:0] w_asqrt46_19;
	wire [2:0] w_asqrt46_20;
	wire [2:0] w_asqrt46_21;
	wire [2:0] w_asqrt46_22;
	wire [2:0] w_asqrt46_23;
	wire [2:0] w_asqrt46_24;
	wire [2:0] w_asqrt46_25;
	wire [2:0] w_asqrt46_26;
	wire [2:0] w_asqrt46_27;
	wire [2:0] w_asqrt46_28;
	wire [2:0] w_asqrt46_29;
	wire [2:0] w_asqrt46_30;
	wire [2:0] w_asqrt46_31;
	wire [2:0] w_asqrt46_32;
	wire [2:0] w_asqrt46_33;
	wire [2:0] w_asqrt46_34;
	wire [2:0] w_asqrt46_35;
	wire [2:0] w_asqrt46_36;
	wire [2:0] w_asqrt46_37;
	wire [2:0] w_asqrt46_38;
	wire [2:0] w_asqrt46_39;
	wire [2:0] w_asqrt46_40;
	wire [1:0] w_asqrt46_41;
	wire asqrt_fa_46;
	wire [2:0] w_asqrt47_0;
	wire [2:0] w_asqrt47_1;
	wire [2:0] w_asqrt47_2;
	wire [2:0] w_asqrt47_3;
	wire [2:0] w_asqrt47_4;
	wire [2:0] w_asqrt47_5;
	wire [2:0] w_asqrt47_6;
	wire [2:0] w_asqrt47_7;
	wire [2:0] w_asqrt47_8;
	wire [2:0] w_asqrt47_9;
	wire [2:0] w_asqrt47_10;
	wire [2:0] w_asqrt47_11;
	wire [2:0] w_asqrt47_12;
	wire [2:0] w_asqrt47_13;
	wire [2:0] w_asqrt47_14;
	wire [2:0] w_asqrt47_15;
	wire [2:0] w_asqrt47_16;
	wire [2:0] w_asqrt47_17;
	wire [2:0] w_asqrt47_18;
	wire [2:0] w_asqrt47_19;
	wire [2:0] w_asqrt47_20;
	wire [2:0] w_asqrt47_21;
	wire [2:0] w_asqrt47_22;
	wire [2:0] w_asqrt47_23;
	wire [2:0] w_asqrt47_24;
	wire [2:0] w_asqrt47_25;
	wire [2:0] w_asqrt47_26;
	wire [2:0] w_asqrt47_27;
	wire [2:0] w_asqrt47_28;
	wire [2:0] w_asqrt47_29;
	wire [2:0] w_asqrt47_30;
	wire [2:0] w_asqrt47_31;
	wire [2:0] w_asqrt47_32;
	wire [2:0] w_asqrt47_33;
	wire [2:0] w_asqrt47_34;
	wire [2:0] w_asqrt47_35;
	wire w_asqrt47_36;
	wire asqrt_fa_47;
	wire [2:0] w_asqrt48_0;
	wire [2:0] w_asqrt48_1;
	wire [2:0] w_asqrt48_2;
	wire [2:0] w_asqrt48_3;
	wire [2:0] w_asqrt48_4;
	wire [2:0] w_asqrt48_5;
	wire [2:0] w_asqrt48_6;
	wire [2:0] w_asqrt48_7;
	wire [2:0] w_asqrt48_8;
	wire [2:0] w_asqrt48_9;
	wire [2:0] w_asqrt48_10;
	wire [2:0] w_asqrt48_11;
	wire [2:0] w_asqrt48_12;
	wire [2:0] w_asqrt48_13;
	wire [2:0] w_asqrt48_14;
	wire [2:0] w_asqrt48_15;
	wire [2:0] w_asqrt48_16;
	wire [2:0] w_asqrt48_17;
	wire [2:0] w_asqrt48_18;
	wire [2:0] w_asqrt48_19;
	wire [2:0] w_asqrt48_20;
	wire [2:0] w_asqrt48_21;
	wire [2:0] w_asqrt48_22;
	wire [2:0] w_asqrt48_23;
	wire [2:0] w_asqrt48_24;
	wire [2:0] w_asqrt48_25;
	wire [2:0] w_asqrt48_26;
	wire [2:0] w_asqrt48_27;
	wire [2:0] w_asqrt48_28;
	wire [2:0] w_asqrt48_29;
	wire [2:0] w_asqrt48_30;
	wire [2:0] w_asqrt48_31;
	wire [2:0] w_asqrt48_32;
	wire [2:0] w_asqrt48_33;
	wire [2:0] w_asqrt48_34;
	wire [2:0] w_asqrt48_35;
	wire [2:0] w_asqrt48_36;
	wire [2:0] w_asqrt48_37;
	wire [2:0] w_asqrt48_38;
	wire [2:0] w_asqrt48_39;
	wire [2:0] w_asqrt48_40;
	wire [2:0] w_asqrt48_41;
	wire w_asqrt48_42;
	wire asqrt_fa_48;
	wire [2:0] w_asqrt49_0;
	wire [2:0] w_asqrt49_1;
	wire [2:0] w_asqrt49_2;
	wire [2:0] w_asqrt49_3;
	wire [2:0] w_asqrt49_4;
	wire [2:0] w_asqrt49_5;
	wire [2:0] w_asqrt49_6;
	wire [2:0] w_asqrt49_7;
	wire [2:0] w_asqrt49_8;
	wire [2:0] w_asqrt49_9;
	wire [2:0] w_asqrt49_10;
	wire [2:0] w_asqrt49_11;
	wire [2:0] w_asqrt49_12;
	wire [2:0] w_asqrt49_13;
	wire [2:0] w_asqrt49_14;
	wire [2:0] w_asqrt49_15;
	wire [2:0] w_asqrt49_16;
	wire [2:0] w_asqrt49_17;
	wire [2:0] w_asqrt49_18;
	wire [2:0] w_asqrt49_19;
	wire [2:0] w_asqrt49_20;
	wire [2:0] w_asqrt49_21;
	wire [2:0] w_asqrt49_22;
	wire [2:0] w_asqrt49_23;
	wire [2:0] w_asqrt49_24;
	wire [2:0] w_asqrt49_25;
	wire [2:0] w_asqrt49_26;
	wire [2:0] w_asqrt49_27;
	wire [2:0] w_asqrt49_28;
	wire [2:0] w_asqrt49_29;
	wire [2:0] w_asqrt49_30;
	wire [2:0] w_asqrt49_31;
	wire [2:0] w_asqrt49_32;
	wire [2:0] w_asqrt49_33;
	wire [2:0] w_asqrt49_34;
	wire [2:0] w_asqrt49_35;
	wire [2:0] w_asqrt49_36;
	wire [1:0] w_asqrt49_37;
	wire asqrt_fa_49;
	wire [2:0] w_asqrt50_0;
	wire [2:0] w_asqrt50_1;
	wire [2:0] w_asqrt50_2;
	wire [2:0] w_asqrt50_3;
	wire [2:0] w_asqrt50_4;
	wire [2:0] w_asqrt50_5;
	wire [2:0] w_asqrt50_6;
	wire [2:0] w_asqrt50_7;
	wire [2:0] w_asqrt50_8;
	wire [2:0] w_asqrt50_9;
	wire [2:0] w_asqrt50_10;
	wire [2:0] w_asqrt50_11;
	wire [2:0] w_asqrt50_12;
	wire [2:0] w_asqrt50_13;
	wire [2:0] w_asqrt50_14;
	wire [2:0] w_asqrt50_15;
	wire [2:0] w_asqrt50_16;
	wire [2:0] w_asqrt50_17;
	wire [2:0] w_asqrt50_18;
	wire [2:0] w_asqrt50_19;
	wire [2:0] w_asqrt50_20;
	wire [2:0] w_asqrt50_21;
	wire [2:0] w_asqrt50_22;
	wire [2:0] w_asqrt50_23;
	wire [2:0] w_asqrt50_24;
	wire [2:0] w_asqrt50_25;
	wire [2:0] w_asqrt50_26;
	wire [2:0] w_asqrt50_27;
	wire [2:0] w_asqrt50_28;
	wire [2:0] w_asqrt50_29;
	wire [2:0] w_asqrt50_30;
	wire [2:0] w_asqrt50_31;
	wire [2:0] w_asqrt50_32;
	wire [2:0] w_asqrt50_33;
	wire [2:0] w_asqrt50_34;
	wire [2:0] w_asqrt50_35;
	wire [2:0] w_asqrt50_36;
	wire [2:0] w_asqrt50_37;
	wire [2:0] w_asqrt50_38;
	wire [2:0] w_asqrt50_39;
	wire [2:0] w_asqrt50_40;
	wire [2:0] w_asqrt50_41;
	wire [2:0] w_asqrt50_42;
	wire w_asqrt50_43;
	wire asqrt_fa_50;
	wire [2:0] w_asqrt51_0;
	wire [2:0] w_asqrt51_1;
	wire [2:0] w_asqrt51_2;
	wire [2:0] w_asqrt51_3;
	wire [2:0] w_asqrt51_4;
	wire [2:0] w_asqrt51_5;
	wire [2:0] w_asqrt51_6;
	wire [2:0] w_asqrt51_7;
	wire [2:0] w_asqrt51_8;
	wire [2:0] w_asqrt51_9;
	wire [2:0] w_asqrt51_10;
	wire [2:0] w_asqrt51_11;
	wire [2:0] w_asqrt51_12;
	wire [2:0] w_asqrt51_13;
	wire [2:0] w_asqrt51_14;
	wire [2:0] w_asqrt51_15;
	wire [2:0] w_asqrt51_16;
	wire [2:0] w_asqrt51_17;
	wire [2:0] w_asqrt51_18;
	wire [2:0] w_asqrt51_19;
	wire [2:0] w_asqrt51_20;
	wire [2:0] w_asqrt51_21;
	wire [2:0] w_asqrt51_22;
	wire [2:0] w_asqrt51_23;
	wire [2:0] w_asqrt51_24;
	wire [2:0] w_asqrt51_25;
	wire [2:0] w_asqrt51_26;
	wire [2:0] w_asqrt51_27;
	wire [2:0] w_asqrt51_28;
	wire [2:0] w_asqrt51_29;
	wire [2:0] w_asqrt51_30;
	wire [2:0] w_asqrt51_31;
	wire [2:0] w_asqrt51_32;
	wire [2:0] w_asqrt51_33;
	wire [2:0] w_asqrt51_34;
	wire [2:0] w_asqrt51_35;
	wire [2:0] w_asqrt51_36;
	wire [2:0] w_asqrt51_37;
	wire [1:0] w_asqrt51_38;
	wire asqrt_fa_51;
	wire [2:0] w_asqrt52_0;
	wire [2:0] w_asqrt52_1;
	wire [2:0] w_asqrt52_2;
	wire [2:0] w_asqrt52_3;
	wire [2:0] w_asqrt52_4;
	wire [2:0] w_asqrt52_5;
	wire [2:0] w_asqrt52_6;
	wire [2:0] w_asqrt52_7;
	wire [2:0] w_asqrt52_8;
	wire [2:0] w_asqrt52_9;
	wire [2:0] w_asqrt52_10;
	wire [2:0] w_asqrt52_11;
	wire [2:0] w_asqrt52_12;
	wire [2:0] w_asqrt52_13;
	wire [2:0] w_asqrt52_14;
	wire [2:0] w_asqrt52_15;
	wire [2:0] w_asqrt52_16;
	wire [2:0] w_asqrt52_17;
	wire [2:0] w_asqrt52_18;
	wire [2:0] w_asqrt52_19;
	wire [2:0] w_asqrt52_20;
	wire [2:0] w_asqrt52_21;
	wire [2:0] w_asqrt52_22;
	wire [2:0] w_asqrt52_23;
	wire [2:0] w_asqrt52_24;
	wire [2:0] w_asqrt52_25;
	wire [2:0] w_asqrt52_26;
	wire [2:0] w_asqrt52_27;
	wire [2:0] w_asqrt52_28;
	wire [2:0] w_asqrt52_29;
	wire [2:0] w_asqrt52_30;
	wire [2:0] w_asqrt52_31;
	wire [2:0] w_asqrt52_32;
	wire [2:0] w_asqrt52_33;
	wire [2:0] w_asqrt52_34;
	wire [2:0] w_asqrt52_35;
	wire [2:0] w_asqrt52_36;
	wire [2:0] w_asqrt52_37;
	wire [2:0] w_asqrt52_38;
	wire [2:0] w_asqrt52_39;
	wire [2:0] w_asqrt52_40;
	wire [2:0] w_asqrt52_41;
	wire [2:0] w_asqrt52_42;
	wire [1:0] w_asqrt52_43;
	wire asqrt_fa_52;
	wire [2:0] w_asqrt53_0;
	wire [2:0] w_asqrt53_1;
	wire [2:0] w_asqrt53_2;
	wire [2:0] w_asqrt53_3;
	wire [2:0] w_asqrt53_4;
	wire [2:0] w_asqrt53_5;
	wire [2:0] w_asqrt53_6;
	wire [2:0] w_asqrt53_7;
	wire [2:0] w_asqrt53_8;
	wire [2:0] w_asqrt53_9;
	wire [2:0] w_asqrt53_10;
	wire [2:0] w_asqrt53_11;
	wire [2:0] w_asqrt53_12;
	wire [2:0] w_asqrt53_13;
	wire [2:0] w_asqrt53_14;
	wire [2:0] w_asqrt53_15;
	wire [2:0] w_asqrt53_16;
	wire [2:0] w_asqrt53_17;
	wire [2:0] w_asqrt53_18;
	wire [2:0] w_asqrt53_19;
	wire [2:0] w_asqrt53_20;
	wire [2:0] w_asqrt53_21;
	wire [2:0] w_asqrt53_22;
	wire [2:0] w_asqrt53_23;
	wire [2:0] w_asqrt53_24;
	wire [2:0] w_asqrt53_25;
	wire [2:0] w_asqrt53_26;
	wire [2:0] w_asqrt53_27;
	wire [2:0] w_asqrt53_28;
	wire [2:0] w_asqrt53_29;
	wire [2:0] w_asqrt53_30;
	wire [2:0] w_asqrt53_31;
	wire [2:0] w_asqrt53_32;
	wire [2:0] w_asqrt53_33;
	wire [2:0] w_asqrt53_34;
	wire [2:0] w_asqrt53_35;
	wire [2:0] w_asqrt53_36;
	wire [2:0] w_asqrt53_37;
	wire [2:0] w_asqrt53_38;
	wire [2:0] w_asqrt53_39;
	wire [1:0] w_asqrt53_40;
	wire asqrt_fa_53;
	wire [2:0] w_asqrt54_0;
	wire [2:0] w_asqrt54_1;
	wire [2:0] w_asqrt54_2;
	wire [2:0] w_asqrt54_3;
	wire [2:0] w_asqrt54_4;
	wire [2:0] w_asqrt54_5;
	wire [2:0] w_asqrt54_6;
	wire [2:0] w_asqrt54_7;
	wire [2:0] w_asqrt54_8;
	wire [2:0] w_asqrt54_9;
	wire [2:0] w_asqrt54_10;
	wire [2:0] w_asqrt54_11;
	wire [2:0] w_asqrt54_12;
	wire [2:0] w_asqrt54_13;
	wire [2:0] w_asqrt54_14;
	wire [2:0] w_asqrt54_15;
	wire [2:0] w_asqrt54_16;
	wire [2:0] w_asqrt54_17;
	wire [2:0] w_asqrt54_18;
	wire [2:0] w_asqrt54_19;
	wire [2:0] w_asqrt54_20;
	wire [2:0] w_asqrt54_21;
	wire [2:0] w_asqrt54_22;
	wire [2:0] w_asqrt54_23;
	wire [2:0] w_asqrt54_24;
	wire [2:0] w_asqrt54_25;
	wire [2:0] w_asqrt54_26;
	wire [2:0] w_asqrt54_27;
	wire [2:0] w_asqrt54_28;
	wire [2:0] w_asqrt54_29;
	wire [2:0] w_asqrt54_30;
	wire [2:0] w_asqrt54_31;
	wire [2:0] w_asqrt54_32;
	wire [2:0] w_asqrt54_33;
	wire [2:0] w_asqrt54_34;
	wire [2:0] w_asqrt54_35;
	wire [2:0] w_asqrt54_36;
	wire [2:0] w_asqrt54_37;
	wire [2:0] w_asqrt54_38;
	wire [2:0] w_asqrt54_39;
	wire [2:0] w_asqrt54_40;
	wire [2:0] w_asqrt54_41;
	wire [2:0] w_asqrt54_42;
	wire [1:0] w_asqrt54_43;
	wire asqrt_fa_54;
	wire [2:0] w_asqrt55_0;
	wire [2:0] w_asqrt55_1;
	wire [2:0] w_asqrt55_2;
	wire [2:0] w_asqrt55_3;
	wire [2:0] w_asqrt55_4;
	wire [2:0] w_asqrt55_5;
	wire [2:0] w_asqrt55_6;
	wire [2:0] w_asqrt55_7;
	wire [2:0] w_asqrt55_8;
	wire [2:0] w_asqrt55_9;
	wire [2:0] w_asqrt55_10;
	wire [2:0] w_asqrt55_11;
	wire [2:0] w_asqrt55_12;
	wire [2:0] w_asqrt55_13;
	wire [2:0] w_asqrt55_14;
	wire [2:0] w_asqrt55_15;
	wire [2:0] w_asqrt55_16;
	wire [2:0] w_asqrt55_17;
	wire [2:0] w_asqrt55_18;
	wire [2:0] w_asqrt55_19;
	wire [2:0] w_asqrt55_20;
	wire [2:0] w_asqrt55_21;
	wire [2:0] w_asqrt55_22;
	wire [2:0] w_asqrt55_23;
	wire [2:0] w_asqrt55_24;
	wire [2:0] w_asqrt55_25;
	wire [2:0] w_asqrt55_26;
	wire [2:0] w_asqrt55_27;
	wire [2:0] w_asqrt55_28;
	wire [2:0] w_asqrt55_29;
	wire [2:0] w_asqrt55_30;
	wire [2:0] w_asqrt55_31;
	wire [2:0] w_asqrt55_32;
	wire [2:0] w_asqrt55_33;
	wire [2:0] w_asqrt55_34;
	wire [2:0] w_asqrt55_35;
	wire [2:0] w_asqrt55_36;
	wire [2:0] w_asqrt55_37;
	wire [2:0] w_asqrt55_38;
	wire [2:0] w_asqrt55_39;
	wire [2:0] w_asqrt55_40;
	wire [1:0] w_asqrt55_41;
	wire asqrt_fa_55;
	wire [2:0] w_asqrt56_0;
	wire [2:0] w_asqrt56_1;
	wire [2:0] w_asqrt56_2;
	wire [2:0] w_asqrt56_3;
	wire [2:0] w_asqrt56_4;
	wire [2:0] w_asqrt56_5;
	wire [2:0] w_asqrt56_6;
	wire [2:0] w_asqrt56_7;
	wire [2:0] w_asqrt56_8;
	wire [2:0] w_asqrt56_9;
	wire [2:0] w_asqrt56_10;
	wire [2:0] w_asqrt56_11;
	wire [2:0] w_asqrt56_12;
	wire [2:0] w_asqrt56_13;
	wire [2:0] w_asqrt56_14;
	wire [2:0] w_asqrt56_15;
	wire [2:0] w_asqrt56_16;
	wire [2:0] w_asqrt56_17;
	wire [2:0] w_asqrt56_18;
	wire [2:0] w_asqrt56_19;
	wire [2:0] w_asqrt56_20;
	wire [2:0] w_asqrt56_21;
	wire [2:0] w_asqrt56_22;
	wire [2:0] w_asqrt56_23;
	wire [2:0] w_asqrt56_24;
	wire [2:0] w_asqrt56_25;
	wire [2:0] w_asqrt56_26;
	wire [2:0] w_asqrt56_27;
	wire [2:0] w_asqrt56_28;
	wire [2:0] w_asqrt56_29;
	wire [2:0] w_asqrt56_30;
	wire [2:0] w_asqrt56_31;
	wire [2:0] w_asqrt56_32;
	wire [2:0] w_asqrt56_33;
	wire [2:0] w_asqrt56_34;
	wire [2:0] w_asqrt56_35;
	wire [2:0] w_asqrt56_36;
	wire [2:0] w_asqrt56_37;
	wire [2:0] w_asqrt56_38;
	wire [2:0] w_asqrt56_39;
	wire [2:0] w_asqrt56_40;
	wire [2:0] w_asqrt56_41;
	wire [2:0] w_asqrt56_42;
	wire [2:0] w_asqrt56_43;
	wire [1:0] w_asqrt56_44;
	wire asqrt_fa_56;
	wire [2:0] w_asqrt57_0;
	wire [2:0] w_asqrt57_1;
	wire [2:0] w_asqrt57_2;
	wire [2:0] w_asqrt57_3;
	wire [2:0] w_asqrt57_4;
	wire [2:0] w_asqrt57_5;
	wire [2:0] w_asqrt57_6;
	wire [2:0] w_asqrt57_7;
	wire [2:0] w_asqrt57_8;
	wire [2:0] w_asqrt57_9;
	wire [2:0] w_asqrt57_10;
	wire [2:0] w_asqrt57_11;
	wire [2:0] w_asqrt57_12;
	wire [2:0] w_asqrt57_13;
	wire [2:0] w_asqrt57_14;
	wire [2:0] w_asqrt57_15;
	wire [2:0] w_asqrt57_16;
	wire [2:0] w_asqrt57_17;
	wire [2:0] w_asqrt57_18;
	wire [2:0] w_asqrt57_19;
	wire [2:0] w_asqrt57_20;
	wire [2:0] w_asqrt57_21;
	wire [2:0] w_asqrt57_22;
	wire [2:0] w_asqrt57_23;
	wire [2:0] w_asqrt57_24;
	wire [2:0] w_asqrt57_25;
	wire [2:0] w_asqrt57_26;
	wire [2:0] w_asqrt57_27;
	wire [2:0] w_asqrt57_28;
	wire [2:0] w_asqrt57_29;
	wire [2:0] w_asqrt57_30;
	wire [2:0] w_asqrt57_31;
	wire [2:0] w_asqrt57_32;
	wire [2:0] w_asqrt57_33;
	wire [2:0] w_asqrt57_34;
	wire [2:0] w_asqrt57_35;
	wire [2:0] w_asqrt57_36;
	wire [2:0] w_asqrt57_37;
	wire [2:0] w_asqrt57_38;
	wire [2:0] w_asqrt57_39;
	wire [2:0] w_asqrt57_40;
	wire [2:0] w_asqrt57_41;
	wire [2:0] w_asqrt57_42;
	wire [1:0] w_asqrt57_43;
	wire asqrt_fa_57;
	wire [2:0] w_asqrt58_0;
	wire [2:0] w_asqrt58_1;
	wire [2:0] w_asqrt58_2;
	wire [2:0] w_asqrt58_3;
	wire [2:0] w_asqrt58_4;
	wire [2:0] w_asqrt58_5;
	wire [2:0] w_asqrt58_6;
	wire [2:0] w_asqrt58_7;
	wire [2:0] w_asqrt58_8;
	wire [2:0] w_asqrt58_9;
	wire [2:0] w_asqrt58_10;
	wire [2:0] w_asqrt58_11;
	wire [2:0] w_asqrt58_12;
	wire [2:0] w_asqrt58_13;
	wire [2:0] w_asqrt58_14;
	wire [2:0] w_asqrt58_15;
	wire [2:0] w_asqrt58_16;
	wire [2:0] w_asqrt58_17;
	wire [2:0] w_asqrt58_18;
	wire [2:0] w_asqrt58_19;
	wire [2:0] w_asqrt58_20;
	wire [2:0] w_asqrt58_21;
	wire [2:0] w_asqrt58_22;
	wire [2:0] w_asqrt58_23;
	wire [2:0] w_asqrt58_24;
	wire [2:0] w_asqrt58_25;
	wire [2:0] w_asqrt58_26;
	wire [2:0] w_asqrt58_27;
	wire [2:0] w_asqrt58_28;
	wire [2:0] w_asqrt58_29;
	wire [2:0] w_asqrt58_30;
	wire [2:0] w_asqrt58_31;
	wire [2:0] w_asqrt58_32;
	wire [2:0] w_asqrt58_33;
	wire [2:0] w_asqrt58_34;
	wire [2:0] w_asqrt58_35;
	wire [2:0] w_asqrt58_36;
	wire [2:0] w_asqrt58_37;
	wire [2:0] w_asqrt58_38;
	wire [2:0] w_asqrt58_39;
	wire [2:0] w_asqrt58_40;
	wire [2:0] w_asqrt58_41;
	wire [2:0] w_asqrt58_42;
	wire [2:0] w_asqrt58_43;
	wire [2:0] w_asqrt58_44;
	wire w_asqrt58_45;
	wire asqrt_fa_58;
	wire [2:0] w_asqrt59_0;
	wire [2:0] w_asqrt59_1;
	wire [2:0] w_asqrt59_2;
	wire [2:0] w_asqrt59_3;
	wire [2:0] w_asqrt59_4;
	wire [2:0] w_asqrt59_5;
	wire [2:0] w_asqrt59_6;
	wire [2:0] w_asqrt59_7;
	wire [2:0] w_asqrt59_8;
	wire [2:0] w_asqrt59_9;
	wire [2:0] w_asqrt59_10;
	wire [2:0] w_asqrt59_11;
	wire [2:0] w_asqrt59_12;
	wire [2:0] w_asqrt59_13;
	wire [2:0] w_asqrt59_14;
	wire [2:0] w_asqrt59_15;
	wire [2:0] w_asqrt59_16;
	wire [2:0] w_asqrt59_17;
	wire [2:0] w_asqrt59_18;
	wire [2:0] w_asqrt59_19;
	wire [2:0] w_asqrt59_20;
	wire [2:0] w_asqrt59_21;
	wire [2:0] w_asqrt59_22;
	wire [2:0] w_asqrt59_23;
	wire [2:0] w_asqrt59_24;
	wire [2:0] w_asqrt59_25;
	wire [2:0] w_asqrt59_26;
	wire [2:0] w_asqrt59_27;
	wire [2:0] w_asqrt59_28;
	wire [2:0] w_asqrt59_29;
	wire [2:0] w_asqrt59_30;
	wire [2:0] w_asqrt59_31;
	wire [2:0] w_asqrt59_32;
	wire [2:0] w_asqrt59_33;
	wire [2:0] w_asqrt59_34;
	wire [2:0] w_asqrt59_35;
	wire [2:0] w_asqrt59_36;
	wire [2:0] w_asqrt59_37;
	wire [2:0] w_asqrt59_38;
	wire [2:0] w_asqrt59_39;
	wire [2:0] w_asqrt59_40;
	wire [2:0] w_asqrt59_41;
	wire [2:0] w_asqrt59_42;
	wire [2:0] w_asqrt59_43;
	wire [1:0] w_asqrt59_44;
	wire asqrt_fa_59;
	wire [2:0] w_asqrt60_0;
	wire [2:0] w_asqrt60_1;
	wire [2:0] w_asqrt60_2;
	wire [2:0] w_asqrt60_3;
	wire [2:0] w_asqrt60_4;
	wire [2:0] w_asqrt60_5;
	wire [2:0] w_asqrt60_6;
	wire [2:0] w_asqrt60_7;
	wire [2:0] w_asqrt60_8;
	wire [2:0] w_asqrt60_9;
	wire [2:0] w_asqrt60_10;
	wire [2:0] w_asqrt60_11;
	wire [2:0] w_asqrt60_12;
	wire [2:0] w_asqrt60_13;
	wire [2:0] w_asqrt60_14;
	wire [2:0] w_asqrt60_15;
	wire [2:0] w_asqrt60_16;
	wire [2:0] w_asqrt60_17;
	wire [2:0] w_asqrt60_18;
	wire [2:0] w_asqrt60_19;
	wire [2:0] w_asqrt60_20;
	wire [2:0] w_asqrt60_21;
	wire [2:0] w_asqrt60_22;
	wire [2:0] w_asqrt60_23;
	wire [2:0] w_asqrt60_24;
	wire [2:0] w_asqrt60_25;
	wire [2:0] w_asqrt60_26;
	wire [2:0] w_asqrt60_27;
	wire [2:0] w_asqrt60_28;
	wire [2:0] w_asqrt60_29;
	wire [2:0] w_asqrt60_30;
	wire [2:0] w_asqrt60_31;
	wire [2:0] w_asqrt60_32;
	wire [2:0] w_asqrt60_33;
	wire [2:0] w_asqrt60_34;
	wire [2:0] w_asqrt60_35;
	wire [2:0] w_asqrt60_36;
	wire [2:0] w_asqrt60_37;
	wire [2:0] w_asqrt60_38;
	wire [2:0] w_asqrt60_39;
	wire [2:0] w_asqrt60_40;
	wire [2:0] w_asqrt60_41;
	wire [2:0] w_asqrt60_42;
	wire [2:0] w_asqrt60_43;
	wire [2:0] w_asqrt60_44;
	wire [1:0] w_asqrt60_45;
	wire asqrt_fa_60;
	wire [2:0] w_asqrt61_0;
	wire [2:0] w_asqrt61_1;
	wire [2:0] w_asqrt61_2;
	wire [2:0] w_asqrt61_3;
	wire [2:0] w_asqrt61_4;
	wire [2:0] w_asqrt61_5;
	wire [2:0] w_asqrt61_6;
	wire [2:0] w_asqrt61_7;
	wire [2:0] w_asqrt61_8;
	wire [2:0] w_asqrt61_9;
	wire [2:0] w_asqrt61_10;
	wire [2:0] w_asqrt61_11;
	wire [2:0] w_asqrt61_12;
	wire [2:0] w_asqrt61_13;
	wire [2:0] w_asqrt61_14;
	wire [2:0] w_asqrt61_15;
	wire [2:0] w_asqrt61_16;
	wire [2:0] w_asqrt61_17;
	wire [2:0] w_asqrt61_18;
	wire [2:0] w_asqrt61_19;
	wire [2:0] w_asqrt61_20;
	wire [2:0] w_asqrt61_21;
	wire [2:0] w_asqrt61_22;
	wire [2:0] w_asqrt61_23;
	wire [2:0] w_asqrt61_24;
	wire [2:0] w_asqrt61_25;
	wire [2:0] w_asqrt61_26;
	wire [2:0] w_asqrt61_27;
	wire [2:0] w_asqrt61_28;
	wire [2:0] w_asqrt61_29;
	wire [2:0] w_asqrt61_30;
	wire [2:0] w_asqrt61_31;
	wire [2:0] w_asqrt61_32;
	wire [2:0] w_asqrt61_33;
	wire [2:0] w_asqrt61_34;
	wire [2:0] w_asqrt61_35;
	wire [2:0] w_asqrt61_36;
	wire [2:0] w_asqrt61_37;
	wire [2:0] w_asqrt61_38;
	wire [2:0] w_asqrt61_39;
	wire [2:0] w_asqrt61_40;
	wire [2:0] w_asqrt61_41;
	wire [2:0] w_asqrt61_42;
	wire [2:0] w_asqrt61_43;
	wire [2:0] w_asqrt61_44;
	wire w_asqrt61_45;
	wire asqrt_fa_61;
	wire [2:0] w_asqrt62_0;
	wire [2:0] w_asqrt62_1;
	wire [2:0] w_asqrt62_2;
	wire [2:0] w_asqrt62_3;
	wire [2:0] w_asqrt62_4;
	wire [2:0] w_asqrt62_5;
	wire [2:0] w_asqrt62_6;
	wire [2:0] w_asqrt62_7;
	wire [2:0] w_asqrt62_8;
	wire [2:0] w_asqrt62_9;
	wire [2:0] w_asqrt62_10;
	wire [2:0] w_asqrt62_11;
	wire [2:0] w_asqrt62_12;
	wire [2:0] w_asqrt62_13;
	wire [2:0] w_asqrt62_14;
	wire [2:0] w_asqrt62_15;
	wire [2:0] w_asqrt62_16;
	wire [2:0] w_asqrt62_17;
	wire [2:0] w_asqrt62_18;
	wire [2:0] w_asqrt62_19;
	wire [2:0] w_asqrt62_20;
	wire [2:0] w_asqrt62_21;
	wire [2:0] w_asqrt62_22;
	wire [2:0] w_asqrt62_23;
	wire [2:0] w_asqrt62_24;
	wire [2:0] w_asqrt62_25;
	wire [2:0] w_asqrt62_26;
	wire [2:0] w_asqrt62_27;
	wire [2:0] w_asqrt62_28;
	wire [2:0] w_asqrt62_29;
	wire [2:0] w_asqrt62_30;
	wire [2:0] w_asqrt62_31;
	wire [2:0] w_asqrt62_32;
	wire [2:0] w_asqrt62_33;
	wire [2:0] w_asqrt62_34;
	wire [2:0] w_asqrt62_35;
	wire [2:0] w_asqrt62_36;
	wire [2:0] w_asqrt62_37;
	wire [2:0] w_asqrt62_38;
	wire [2:0] w_asqrt62_39;
	wire [2:0] w_asqrt62_40;
	wire [2:0] w_asqrt62_41;
	wire [2:0] w_asqrt62_42;
	wire [2:0] w_asqrt62_43;
	wire [2:0] w_asqrt62_44;
	wire [1:0] w_asqrt62_45;
	wire asqrt_fa_62;
	wire [2:0] w_asqrt63_0;
	wire [2:0] w_asqrt63_1;
	wire [2:0] w_asqrt63_2;
	wire [2:0] w_asqrt63_3;
	wire [2:0] w_asqrt63_4;
	wire [2:0] w_asqrt63_5;
	wire [2:0] w_asqrt63_6;
	wire [2:0] w_asqrt63_7;
	wire [2:0] w_asqrt63_8;
	wire [2:0] w_asqrt63_9;
	wire [2:0] w_asqrt63_10;
	wire [2:0] w_asqrt63_11;
	wire [2:0] w_asqrt63_12;
	wire [2:0] w_asqrt63_13;
	wire [2:0] w_asqrt63_14;
	wire [2:0] w_asqrt63_15;
	wire [2:0] w_asqrt63_16;
	wire [2:0] w_asqrt63_17;
	wire [2:0] w_asqrt63_18;
	wire [2:0] w_asqrt63_19;
	wire [2:0] w_asqrt63_20;
	wire [2:0] w_asqrt63_21;
	wire [2:0] w_asqrt63_22;
	wire [2:0] w_asqrt63_23;
	wire [2:0] w_asqrt63_24;
	wire [2:0] w_asqrt63_25;
	wire [2:0] w_asqrt63_26;
	wire [2:0] w_asqrt63_27;
	wire [2:0] w_asqrt63_28;
	wire [2:0] w_asqrt63_29;
	wire [2:0] w_asqrt63_30;
	wire [2:0] w_asqrt63_31;
	wire [2:0] w_asqrt63_32;
	wire [2:0] w_asqrt63_33;
	wire [2:0] w_asqrt63_34;
	wire [2:0] w_asqrt63_35;
	wire [2:0] w_asqrt63_36;
	wire [2:0] w_asqrt63_37;
	wire [2:0] w_asqrt63_38;
	wire [2:0] w_asqrt63_39;
	wire [2:0] w_asqrt63_40;
	wire [2:0] w_asqrt63_41;
	wire [2:0] w_asqrt63_42;
	wire [2:0] w_asqrt63_43;
	wire [2:0] w_asqrt63_44;
	wire [2:0] w_asqrt63_45;
	wire [2:0] w_asqrt63_46;
	wire [2:0] w_asqrt63_47;
	wire [2:0] w_asqrt63_48;
	wire [2:0] w_asqrt63_49;
	wire [2:0] w_asqrt63_50;
	wire [2:0] w_asqrt63_51;
	wire [2:0] w_asqrt63_52;
	wire [2:0] w_asqrt63_53;
	wire [2:0] w_asqrt63_54;
	wire [2:0] w_asqrt63_55;
	wire [2:0] w_asqrt63_56;
	wire w_asqrt63_57;
	wire asqrt_fa_63;
	wire [2:0] w_n192_0;
	wire [1:0] w_n193_0;
	wire [1:0] w_n195_0;
	wire [1:0] w_n197_0;
	wire [2:0] w_n198_0;
	wire [1:0] w_n198_1;
	wire [1:0] w_n199_0;
	wire [2:0] w_n200_0;
	wire [1:0] w_n203_0;
	wire [2:0] w_n204_0;
	wire [1:0] w_n207_0;
	wire [1:0] w_n209_0;
	wire [2:0] w_n211_0;
	wire [1:0] w_n211_1;
	wire [1:0] w_n212_0;
	wire [2:0] w_n215_0;
	wire [2:0] w_n216_0;
	wire [1:0] w_n216_1;
	wire [1:0] w_n217_0;
	wire [2:0] w_n218_0;
	wire [2:0] w_n218_1;
	wire [2:0] w_n218_2;
	wire [2:0] w_n218_3;
	wire [2:0] w_n218_4;
	wire [2:0] w_n218_5;
	wire [2:0] w_n218_6;
	wire [2:0] w_n218_7;
	wire [2:0] w_n218_8;
	wire [2:0] w_n218_9;
	wire [2:0] w_n218_10;
	wire [2:0] w_n218_11;
	wire [2:0] w_n218_12;
	wire [2:0] w_n218_13;
	wire [2:0] w_n218_14;
	wire [2:0] w_n218_15;
	wire [2:0] w_n218_16;
	wire [2:0] w_n218_17;
	wire [2:0] w_n218_18;
	wire [2:0] w_n218_19;
	wire [2:0] w_n218_20;
	wire [2:0] w_n218_21;
	wire [2:0] w_n218_22;
	wire [2:0] w_n218_23;
	wire [2:0] w_n218_24;
	wire [2:0] w_n218_25;
	wire [2:0] w_n218_26;
	wire [2:0] w_n218_27;
	wire [2:0] w_n218_28;
	wire [2:0] w_n218_29;
	wire [2:0] w_n218_30;
	wire [1:0] w_n218_31;
	wire [2:0] w_n221_0;
	wire [2:0] w_n221_1;
	wire [2:0] w_n221_2;
	wire [2:0] w_n221_3;
	wire [2:0] w_n221_4;
	wire [2:0] w_n221_5;
	wire [2:0] w_n221_6;
	wire [2:0] w_n221_7;
	wire [2:0] w_n221_8;
	wire [2:0] w_n221_9;
	wire [2:0] w_n221_10;
	wire [2:0] w_n221_11;
	wire [2:0] w_n221_12;
	wire [2:0] w_n221_13;
	wire [2:0] w_n221_14;
	wire [2:0] w_n221_15;
	wire [2:0] w_n221_16;
	wire [2:0] w_n221_17;
	wire [2:0] w_n221_18;
	wire [2:0] w_n221_19;
	wire [2:0] w_n221_20;
	wire [2:0] w_n221_21;
	wire [2:0] w_n221_22;
	wire [2:0] w_n221_23;
	wire [2:0] w_n221_24;
	wire [2:0] w_n221_25;
	wire [2:0] w_n221_26;
	wire [2:0] w_n221_27;
	wire [2:0] w_n221_28;
	wire [2:0] w_n221_29;
	wire [2:0] w_n221_30;
	wire [2:0] w_n221_31;
	wire [2:0] w_n221_32;
	wire [2:0] w_n221_33;
	wire [2:0] w_n221_34;
	wire [2:0] w_n221_35;
	wire [2:0] w_n221_36;
	wire [2:0] w_n221_37;
	wire [2:0] w_n221_38;
	wire [2:0] w_n221_39;
	wire [2:0] w_n221_40;
	wire [2:0] w_n221_41;
	wire [2:0] w_n221_42;
	wire [2:0] w_n221_43;
	wire [2:0] w_n221_44;
	wire [2:0] w_n221_45;
	wire [2:0] w_n221_46;
	wire [2:0] w_n221_47;
	wire [2:0] w_n221_48;
	wire [2:0] w_n221_49;
	wire [2:0] w_n221_50;
	wire [2:0] w_n221_51;
	wire [2:0] w_n221_52;
	wire [2:0] w_n221_53;
	wire [2:0] w_n221_54;
	wire [2:0] w_n221_55;
	wire [2:0] w_n221_56;
	wire [2:0] w_n221_57;
	wire [2:0] w_n221_58;
	wire [2:0] w_n221_59;
	wire [2:0] w_n221_60;
	wire [2:0] w_n221_61;
	wire [2:0] w_n221_62;
	wire [2:0] w_n221_63;
	wire [2:0] w_n221_64;
	wire [2:0] w_n221_65;
	wire [2:0] w_n221_66;
	wire [2:0] w_n221_67;
	wire [2:0] w_n221_68;
	wire [2:0] w_n221_69;
	wire [2:0] w_n221_70;
	wire [2:0] w_n221_71;
	wire [2:0] w_n221_72;
	wire [2:0] w_n221_73;
	wire [2:0] w_n221_74;
	wire [2:0] w_n221_75;
	wire [1:0] w_n221_76;
	wire [1:0] w_n224_0;
	wire [1:0] w_n225_0;
	wire [1:0] w_n234_0;
	wire [1:0] w_n235_0;
	wire [1:0] w_n236_0;
	wire [2:0] w_n239_0;
	wire [2:0] w_n239_1;
	wire [2:0] w_n239_2;
	wire [2:0] w_n239_3;
	wire [2:0] w_n239_4;
	wire [2:0] w_n239_5;
	wire [2:0] w_n239_6;
	wire [2:0] w_n239_7;
	wire [2:0] w_n239_8;
	wire [2:0] w_n239_9;
	wire [2:0] w_n239_10;
	wire [2:0] w_n239_11;
	wire [2:0] w_n239_12;
	wire [2:0] w_n239_13;
	wire [2:0] w_n239_14;
	wire [2:0] w_n239_15;
	wire [2:0] w_n239_16;
	wire [2:0] w_n239_17;
	wire [2:0] w_n239_18;
	wire [2:0] w_n239_19;
	wire [2:0] w_n239_20;
	wire [2:0] w_n239_21;
	wire [2:0] w_n239_22;
	wire [2:0] w_n239_23;
	wire [2:0] w_n239_24;
	wire [2:0] w_n239_25;
	wire [2:0] w_n239_26;
	wire [2:0] w_n239_27;
	wire [2:0] w_n239_28;
	wire [2:0] w_n239_29;
	wire [2:0] w_n239_30;
	wire [2:0] w_n239_31;
	wire [2:0] w_n239_32;
	wire [2:0] w_n239_33;
	wire [2:0] w_n239_34;
	wire [2:0] w_n239_35;
	wire [2:0] w_n239_36;
	wire [2:0] w_n239_37;
	wire [2:0] w_n239_38;
	wire [2:0] w_n239_39;
	wire [2:0] w_n239_40;
	wire [2:0] w_n239_41;
	wire [2:0] w_n239_42;
	wire [2:0] w_n239_43;
	wire [2:0] w_n239_44;
	wire [2:0] w_n239_45;
	wire [2:0] w_n239_46;
	wire [2:0] w_n239_47;
	wire [2:0] w_n239_48;
	wire [2:0] w_n239_49;
	wire [2:0] w_n239_50;
	wire [2:0] w_n239_51;
	wire [2:0] w_n239_52;
	wire [2:0] w_n239_53;
	wire [2:0] w_n239_54;
	wire [2:0] w_n239_55;
	wire [2:0] w_n239_56;
	wire [2:0] w_n239_57;
	wire [2:0] w_n239_58;
	wire [2:0] w_n239_59;
	wire [2:0] w_n239_60;
	wire [2:0] w_n239_61;
	wire [2:0] w_n239_62;
	wire [2:0] w_n239_63;
	wire [2:0] w_n239_64;
	wire [2:0] w_n239_65;
	wire [2:0] w_n239_66;
	wire [2:0] w_n239_67;
	wire [2:0] w_n239_68;
	wire [2:0] w_n239_69;
	wire [2:0] w_n239_70;
	wire [2:0] w_n239_71;
	wire [2:0] w_n239_72;
	wire [2:0] w_n239_73;
	wire [2:0] w_n239_74;
	wire [1:0] w_n239_75;
	wire [2:0] w_n241_0;
	wire [2:0] w_n241_1;
	wire [1:0] w_n242_0;
	wire [2:0] w_n243_0;
	wire [1:0] w_n244_0;
	wire [2:0] w_n246_0;
	wire [1:0] w_n247_0;
	wire [1:0] w_n249_0;
	wire [1:0] w_n250_0;
	wire [2:0] w_n252_0;
	wire [2:0] w_n256_0;
	wire [1:0] w_n256_1;
	wire [1:0] w_n260_0;
	wire [1:0] w_n261_0;
	wire [1:0] w_n264_0;
	wire [2:0] w_n267_0;
	wire [1:0] w_n267_1;
	wire [2:0] w_n268_0;
	wire [1:0] w_n268_1;
	wire [1:0] w_n269_0;
	wire [2:0] w_n270_0;
	wire [1:0] w_n271_0;
	wire [2:0] w_n273_0;
	wire [1:0] w_n274_0;
	wire [1:0] w_n287_0;
	wire [2:0] w_n294_0;
	wire [2:0] w_n294_1;
	wire [2:0] w_n294_2;
	wire [2:0] w_n294_3;
	wire [2:0] w_n294_4;
	wire [2:0] w_n294_5;
	wire [2:0] w_n294_6;
	wire [2:0] w_n294_7;
	wire [2:0] w_n294_8;
	wire [2:0] w_n294_9;
	wire [2:0] w_n294_10;
	wire [2:0] w_n294_11;
	wire [2:0] w_n294_12;
	wire [2:0] w_n294_13;
	wire [2:0] w_n294_14;
	wire [2:0] w_n294_15;
	wire [2:0] w_n294_16;
	wire [2:0] w_n294_17;
	wire [2:0] w_n294_18;
	wire [2:0] w_n294_19;
	wire [2:0] w_n294_20;
	wire [2:0] w_n294_21;
	wire [2:0] w_n294_22;
	wire [2:0] w_n294_23;
	wire [2:0] w_n294_24;
	wire [2:0] w_n294_25;
	wire [2:0] w_n294_26;
	wire [2:0] w_n294_27;
	wire [2:0] w_n294_28;
	wire [2:0] w_n294_29;
	wire [2:0] w_n294_30;
	wire [2:0] w_n294_31;
	wire [2:0] w_n294_32;
	wire [2:0] w_n294_33;
	wire [2:0] w_n294_34;
	wire [2:0] w_n294_35;
	wire [2:0] w_n294_36;
	wire [2:0] w_n294_37;
	wire [2:0] w_n294_38;
	wire [2:0] w_n294_39;
	wire [2:0] w_n294_40;
	wire [2:0] w_n294_41;
	wire [2:0] w_n294_42;
	wire [2:0] w_n294_43;
	wire [2:0] w_n294_44;
	wire [2:0] w_n294_45;
	wire [2:0] w_n294_46;
	wire [2:0] w_n294_47;
	wire [2:0] w_n294_48;
	wire [2:0] w_n294_49;
	wire [2:0] w_n294_50;
	wire [2:0] w_n294_51;
	wire [2:0] w_n294_52;
	wire [2:0] w_n294_53;
	wire [2:0] w_n294_54;
	wire [2:0] w_n294_55;
	wire [2:0] w_n294_56;
	wire [2:0] w_n294_57;
	wire [2:0] w_n294_58;
	wire [2:0] w_n294_59;
	wire [2:0] w_n294_60;
	wire [2:0] w_n294_61;
	wire [2:0] w_n294_62;
	wire [2:0] w_n294_63;
	wire [2:0] w_n294_64;
	wire [2:0] w_n294_65;
	wire [2:0] w_n294_66;
	wire [2:0] w_n294_67;
	wire [2:0] w_n294_68;
	wire [2:0] w_n294_69;
	wire [2:0] w_n294_70;
	wire [2:0] w_n294_71;
	wire [2:0] w_n294_72;
	wire [2:0] w_n294_73;
	wire [2:0] w_n294_74;
	wire [1:0] w_n294_75;
	wire [1:0] w_n295_0;
	wire [2:0] w_n298_0;
	wire [1:0] w_n299_0;
	wire [1:0] w_n303_0;
	wire [1:0] w_n304_0;
	wire [1:0] w_n306_0;
	wire [1:0] w_n307_0;
	wire [1:0] w_n308_0;
	wire [1:0] w_n321_0;
	wire [1:0] w_n329_0;
	wire [1:0] w_n330_0;
	wire [2:0] w_n333_0;
	wire [1:0] w_n335_0;
	wire [1:0] w_n337_0;
	wire [1:0] w_n338_0;
	wire [1:0] w_n342_0;
	wire [1:0] w_n343_0;
	wire [1:0] w_n345_0;
	wire [1:0] w_n349_0;
	wire [2:0] w_n352_0;
	wire [2:0] w_n352_1;
	wire [2:0] w_n352_2;
	wire [2:0] w_n352_3;
	wire [2:0] w_n352_4;
	wire [2:0] w_n352_5;
	wire [2:0] w_n352_6;
	wire [2:0] w_n352_7;
	wire [2:0] w_n352_8;
	wire [2:0] w_n352_9;
	wire [2:0] w_n352_10;
	wire [2:0] w_n352_11;
	wire [2:0] w_n352_12;
	wire [2:0] w_n352_13;
	wire [2:0] w_n352_14;
	wire [2:0] w_n352_15;
	wire [2:0] w_n352_16;
	wire [2:0] w_n352_17;
	wire [2:0] w_n352_18;
	wire [2:0] w_n352_19;
	wire [2:0] w_n352_20;
	wire [2:0] w_n352_21;
	wire [2:0] w_n352_22;
	wire [2:0] w_n352_23;
	wire [2:0] w_n352_24;
	wire [2:0] w_n352_25;
	wire [2:0] w_n352_26;
	wire [2:0] w_n352_27;
	wire [2:0] w_n352_28;
	wire [2:0] w_n352_29;
	wire [2:0] w_n352_30;
	wire [2:0] w_n352_31;
	wire [2:0] w_n352_32;
	wire [2:0] w_n352_33;
	wire [2:0] w_n352_34;
	wire [2:0] w_n352_35;
	wire [2:0] w_n352_36;
	wire [2:0] w_n352_37;
	wire [2:0] w_n352_38;
	wire [2:0] w_n352_39;
	wire [2:0] w_n352_40;
	wire [2:0] w_n352_41;
	wire [2:0] w_n352_42;
	wire [2:0] w_n352_43;
	wire [2:0] w_n352_44;
	wire [2:0] w_n352_45;
	wire [2:0] w_n352_46;
	wire [2:0] w_n352_47;
	wire [2:0] w_n352_48;
	wire [2:0] w_n352_49;
	wire [2:0] w_n352_50;
	wire [2:0] w_n352_51;
	wire [2:0] w_n352_52;
	wire [2:0] w_n352_53;
	wire [2:0] w_n352_54;
	wire [2:0] w_n352_55;
	wire [2:0] w_n352_56;
	wire [2:0] w_n352_57;
	wire [2:0] w_n352_58;
	wire [2:0] w_n352_59;
	wire [2:0] w_n352_60;
	wire [2:0] w_n352_61;
	wire [2:0] w_n352_62;
	wire [2:0] w_n352_63;
	wire [2:0] w_n352_64;
	wire [2:0] w_n352_65;
	wire [2:0] w_n352_66;
	wire [2:0] w_n352_67;
	wire [2:0] w_n352_68;
	wire [2:0] w_n352_69;
	wire [2:0] w_n352_70;
	wire [2:0] w_n352_71;
	wire [2:0] w_n352_72;
	wire [2:0] w_n352_73;
	wire [1:0] w_n352_74;
	wire [2:0] w_n354_0;
	wire [2:0] w_n354_1;
	wire [1:0] w_n355_0;
	wire [2:0] w_n356_0;
	wire [1:0] w_n357_0;
	wire [2:0] w_n359_0;
	wire [1:0] w_n360_0;
	wire [2:0] w_n367_0;
	wire [1:0] w_n368_0;
	wire [1:0] w_n371_0;
	wire [2:0] w_n373_0;
	wire [2:0] w_n375_0;
	wire [1:0] w_n376_0;
	wire [2:0] w_n380_0;
	wire [2:0] w_n383_0;
	wire [2:0] w_n386_0;
	wire [1:0] w_n386_1;
	wire [2:0] w_n387_0;
	wire [1:0] w_n388_0;
	wire [1:0] w_n389_0;
	wire [1:0] w_n390_0;
	wire [1:0] w_n393_0;
	wire [1:0] w_n395_0;
	wire [1:0] w_n407_0;
	wire [1:0] w_n418_0;
	wire [1:0] w_n419_0;
	wire [2:0] w_n422_0;
	wire [1:0] w_n423_0;
	wire [2:0] w_n425_0;
	wire [1:0] w_n425_1;
	wire [1:0] w_n426_0;
	wire [2:0] w_n427_0;
	wire [1:0] w_n428_0;
	wire [2:0] w_n429_0;
	wire [1:0] w_n430_0;
	wire [1:0] w_n435_0;
	wire [1:0] w_n440_0;
	wire [1:0] w_n441_0;
	wire [2:0] w_n443_0;
	wire [2:0] w_n443_1;
	wire [2:0] w_n443_2;
	wire [2:0] w_n443_3;
	wire [2:0] w_n443_4;
	wire [2:0] w_n443_5;
	wire [2:0] w_n443_6;
	wire [2:0] w_n443_7;
	wire [2:0] w_n443_8;
	wire [2:0] w_n443_9;
	wire [2:0] w_n443_10;
	wire [2:0] w_n443_11;
	wire [2:0] w_n443_12;
	wire [2:0] w_n443_13;
	wire [2:0] w_n443_14;
	wire [2:0] w_n443_15;
	wire [2:0] w_n443_16;
	wire [2:0] w_n443_17;
	wire [2:0] w_n443_18;
	wire [2:0] w_n443_19;
	wire [2:0] w_n443_20;
	wire [2:0] w_n443_21;
	wire [2:0] w_n443_22;
	wire [2:0] w_n443_23;
	wire [2:0] w_n443_24;
	wire [2:0] w_n443_25;
	wire [2:0] w_n443_26;
	wire [2:0] w_n443_27;
	wire [2:0] w_n443_28;
	wire [2:0] w_n443_29;
	wire [2:0] w_n443_30;
	wire [2:0] w_n443_31;
	wire [2:0] w_n443_32;
	wire [2:0] w_n443_33;
	wire [2:0] w_n443_34;
	wire [2:0] w_n443_35;
	wire [2:0] w_n443_36;
	wire [2:0] w_n443_37;
	wire [2:0] w_n443_38;
	wire [2:0] w_n443_39;
	wire [2:0] w_n443_40;
	wire [2:0] w_n443_41;
	wire [2:0] w_n443_42;
	wire [2:0] w_n443_43;
	wire [2:0] w_n443_44;
	wire [2:0] w_n443_45;
	wire [2:0] w_n443_46;
	wire [2:0] w_n443_47;
	wire [2:0] w_n443_48;
	wire [2:0] w_n443_49;
	wire [2:0] w_n443_50;
	wire [2:0] w_n443_51;
	wire [2:0] w_n443_52;
	wire [2:0] w_n443_53;
	wire [2:0] w_n443_54;
	wire [2:0] w_n443_55;
	wire [2:0] w_n443_56;
	wire [2:0] w_n443_57;
	wire [2:0] w_n443_58;
	wire [2:0] w_n443_59;
	wire [2:0] w_n443_60;
	wire [2:0] w_n443_61;
	wire [2:0] w_n443_62;
	wire [2:0] w_n443_63;
	wire [2:0] w_n443_64;
	wire [2:0] w_n443_65;
	wire [2:0] w_n443_66;
	wire [2:0] w_n443_67;
	wire [2:0] w_n443_68;
	wire [2:0] w_n443_69;
	wire [2:0] w_n443_70;
	wire [2:0] w_n443_71;
	wire [2:0] w_n443_72;
	wire [1:0] w_n443_73;
	wire [2:0] w_n447_0;
	wire [1:0] w_n448_0;
	wire [1:0] w_n450_0;
	wire [1:0] w_n452_0;
	wire [1:0] w_n453_0;
	wire [2:0] w_n455_0;
	wire [1:0] w_n456_0;
	wire [1:0] w_n460_0;
	wire [2:0] w_n462_0;
	wire [1:0] w_n463_0;
	wire [1:0] w_n474_0;
	wire [1:0] w_n481_0;
	wire [2:0] w_n487_0;
	wire [1:0] w_n489_0;
	wire [1:0] w_n490_0;
	wire [1:0] w_n493_0;
	wire [1:0] w_n499_0;
	wire [2:0] w_n500_0;
	wire [1:0] w_n504_0;
	wire [1:0] w_n507_0;
	wire [1:0] w_n511_0;
	wire [2:0] w_n515_0;
	wire [2:0] w_n515_1;
	wire [2:0] w_n515_2;
	wire [2:0] w_n515_3;
	wire [2:0] w_n515_4;
	wire [2:0] w_n515_5;
	wire [2:0] w_n515_6;
	wire [2:0] w_n515_7;
	wire [2:0] w_n515_8;
	wire [2:0] w_n515_9;
	wire [2:0] w_n515_10;
	wire [2:0] w_n515_11;
	wire [2:0] w_n515_12;
	wire [2:0] w_n515_13;
	wire [2:0] w_n515_14;
	wire [2:0] w_n515_15;
	wire [2:0] w_n515_16;
	wire [2:0] w_n515_17;
	wire [2:0] w_n515_18;
	wire [2:0] w_n515_19;
	wire [2:0] w_n515_20;
	wire [2:0] w_n515_21;
	wire [2:0] w_n515_22;
	wire [2:0] w_n515_23;
	wire [2:0] w_n515_24;
	wire [2:0] w_n515_25;
	wire [2:0] w_n515_26;
	wire [2:0] w_n515_27;
	wire [2:0] w_n515_28;
	wire [2:0] w_n515_29;
	wire [2:0] w_n515_30;
	wire [2:0] w_n515_31;
	wire [2:0] w_n515_32;
	wire [2:0] w_n515_33;
	wire [2:0] w_n515_34;
	wire [2:0] w_n515_35;
	wire [2:0] w_n515_36;
	wire [2:0] w_n515_37;
	wire [2:0] w_n515_38;
	wire [2:0] w_n515_39;
	wire [2:0] w_n515_40;
	wire [2:0] w_n515_41;
	wire [2:0] w_n515_42;
	wire [2:0] w_n515_43;
	wire [2:0] w_n515_44;
	wire [2:0] w_n515_45;
	wire [2:0] w_n515_46;
	wire [2:0] w_n515_47;
	wire [2:0] w_n515_48;
	wire [2:0] w_n515_49;
	wire [2:0] w_n515_50;
	wire [2:0] w_n515_51;
	wire [2:0] w_n515_52;
	wire [2:0] w_n515_53;
	wire [2:0] w_n515_54;
	wire [2:0] w_n515_55;
	wire [2:0] w_n515_56;
	wire [2:0] w_n515_57;
	wire [2:0] w_n515_58;
	wire [2:0] w_n515_59;
	wire [2:0] w_n515_60;
	wire [2:0] w_n515_61;
	wire [2:0] w_n515_62;
	wire [2:0] w_n515_63;
	wire [2:0] w_n515_64;
	wire [2:0] w_n515_65;
	wire [2:0] w_n515_66;
	wire [2:0] w_n515_67;
	wire [2:0] w_n515_68;
	wire [2:0] w_n515_69;
	wire [2:0] w_n515_70;
	wire [2:0] w_n515_71;
	wire [2:0] w_n515_72;
	wire [1:0] w_n515_73;
	wire [2:0] w_n518_0;
	wire [2:0] w_n519_0;
	wire [2:0] w_n521_0;
	wire [2:0] w_n521_1;
	wire [1:0] w_n522_0;
	wire [2:0] w_n523_0;
	wire [1:0] w_n524_0;
	wire [2:0] w_n526_0;
	wire [1:0] w_n527_0;
	wire [2:0] w_n534_0;
	wire [1:0] w_n535_0;
	wire [1:0] w_n538_0;
	wire [1:0] w_n539_0;
	wire [2:0] w_n544_0;
	wire [2:0] w_n546_0;
	wire [1:0] w_n547_0;
	wire [2:0] w_n551_0;
	wire [2:0] w_n554_0;
	wire [1:0] w_n555_0;
	wire [2:0] w_n559_0;
	wire [2:0] w_n561_0;
	wire [1:0] w_n562_0;
	wire [2:0] w_n566_0;
	wire [2:0] w_n569_0;
	wire [1:0] w_n570_0;
	wire [1:0] w_n572_0;
	wire [1:0] w_n575_0;
	wire [1:0] w_n576_0;
	wire [1:0] w_n581_0;
	wire [1:0] w_n582_0;
	wire [2:0] w_n588_0;
	wire [2:0] w_n589_0;
	wire [1:0] w_n589_1;
	wire [1:0] w_n590_0;
	wire [2:0] w_n591_0;
	wire [1:0] w_n592_0;
	wire [2:0] w_n594_0;
	wire [1:0] w_n595_0;
	wire [1:0] w_n610_0;
	wire [1:0] w_n626_0;
	wire [1:0] w_n627_0;
	wire [1:0] w_n630_0;
	wire [2:0] w_n632_0;
	wire [2:0] w_n635_0;
	wire [2:0] w_n635_1;
	wire [2:0] w_n635_2;
	wire [2:0] w_n635_3;
	wire [2:0] w_n635_4;
	wire [2:0] w_n635_5;
	wire [2:0] w_n635_6;
	wire [2:0] w_n635_7;
	wire [2:0] w_n635_8;
	wire [2:0] w_n635_9;
	wire [2:0] w_n635_10;
	wire [2:0] w_n635_11;
	wire [2:0] w_n635_12;
	wire [2:0] w_n635_13;
	wire [2:0] w_n635_14;
	wire [2:0] w_n635_15;
	wire [2:0] w_n635_16;
	wire [2:0] w_n635_17;
	wire [2:0] w_n635_18;
	wire [2:0] w_n635_19;
	wire [2:0] w_n635_20;
	wire [2:0] w_n635_21;
	wire [2:0] w_n635_22;
	wire [2:0] w_n635_23;
	wire [2:0] w_n635_24;
	wire [2:0] w_n635_25;
	wire [2:0] w_n635_26;
	wire [2:0] w_n635_27;
	wire [2:0] w_n635_28;
	wire [2:0] w_n635_29;
	wire [2:0] w_n635_30;
	wire [2:0] w_n635_31;
	wire [2:0] w_n635_32;
	wire [2:0] w_n635_33;
	wire [2:0] w_n635_34;
	wire [2:0] w_n635_35;
	wire [2:0] w_n635_36;
	wire [2:0] w_n635_37;
	wire [2:0] w_n635_38;
	wire [2:0] w_n635_39;
	wire [2:0] w_n635_40;
	wire [2:0] w_n635_41;
	wire [2:0] w_n635_42;
	wire [2:0] w_n635_43;
	wire [2:0] w_n635_44;
	wire [2:0] w_n635_45;
	wire [2:0] w_n635_46;
	wire [2:0] w_n635_47;
	wire [2:0] w_n635_48;
	wire [2:0] w_n635_49;
	wire [2:0] w_n635_50;
	wire [2:0] w_n635_51;
	wire [2:0] w_n635_52;
	wire [2:0] w_n635_53;
	wire [2:0] w_n635_54;
	wire [2:0] w_n635_55;
	wire [2:0] w_n635_56;
	wire [2:0] w_n635_57;
	wire [2:0] w_n635_58;
	wire [2:0] w_n635_59;
	wire [2:0] w_n635_60;
	wire [2:0] w_n635_61;
	wire [2:0] w_n635_62;
	wire [2:0] w_n635_63;
	wire [2:0] w_n635_64;
	wire [2:0] w_n635_65;
	wire [2:0] w_n635_66;
	wire [2:0] w_n635_67;
	wire [2:0] w_n635_68;
	wire [2:0] w_n635_69;
	wire [2:0] w_n635_70;
	wire [2:0] w_n639_0;
	wire [1:0] w_n640_0;
	wire [1:0] w_n642_0;
	wire [1:0] w_n647_0;
	wire [1:0] w_n648_0;
	wire [2:0] w_n650_0;
	wire [1:0] w_n651_0;
	wire [1:0] w_n655_0;
	wire [2:0] w_n657_0;
	wire [1:0] w_n658_0;
	wire [1:0] w_n662_0;
	wire [1:0] w_n663_0;
	wire [2:0] w_n665_0;
	wire [1:0] w_n666_0;
	wire [1:0] w_n670_0;
	wire [2:0] w_n672_0;
	wire [1:0] w_n673_0;
	wire [1:0] w_n677_0;
	wire [1:0] w_n678_0;
	wire [1:0] w_n680_0;
	wire [2:0] w_n681_0;
	wire [1:0] w_n681_1;
	wire [2:0] w_n682_0;
	wire [1:0] w_n686_0;
	wire [1:0] w_n687_0;
	wire [1:0] w_n701_0;
	wire [1:0] w_n708_0;
	wire [1:0] w_n715_0;
	wire [1:0] w_n720_0;
	wire [1:0] w_n721_0;
	wire [1:0] w_n723_0;
	wire [1:0] w_n725_0;
	wire [1:0] w_n726_0;
	wire [1:0] w_n728_0;
	wire [2:0] w_n730_0;
	wire [2:0] w_n730_1;
	wire [1:0] w_n731_0;
	wire [2:0] w_n732_0;
	wire [1:0] w_n733_0;
	wire [1:0] w_n736_0;
	wire [1:0] w_n742_0;
	wire [2:0] w_n743_0;
	wire [2:0] w_n743_1;
	wire [2:0] w_n743_2;
	wire [2:0] w_n743_3;
	wire [2:0] w_n743_4;
	wire [2:0] w_n743_5;
	wire [2:0] w_n743_6;
	wire [2:0] w_n743_7;
	wire [2:0] w_n743_8;
	wire [2:0] w_n743_9;
	wire [2:0] w_n743_10;
	wire [2:0] w_n743_11;
	wire [2:0] w_n743_12;
	wire [2:0] w_n743_13;
	wire [2:0] w_n743_14;
	wire [2:0] w_n743_15;
	wire [2:0] w_n743_16;
	wire [2:0] w_n743_17;
	wire [2:0] w_n743_18;
	wire [2:0] w_n743_19;
	wire [2:0] w_n743_20;
	wire [2:0] w_n743_21;
	wire [2:0] w_n743_22;
	wire [2:0] w_n743_23;
	wire [2:0] w_n743_24;
	wire [2:0] w_n743_25;
	wire [2:0] w_n743_26;
	wire [2:0] w_n743_27;
	wire [2:0] w_n743_28;
	wire [2:0] w_n743_29;
	wire [2:0] w_n743_30;
	wire [2:0] w_n743_31;
	wire [2:0] w_n743_32;
	wire [2:0] w_n743_33;
	wire [2:0] w_n743_34;
	wire [2:0] w_n743_35;
	wire [2:0] w_n743_36;
	wire [2:0] w_n743_37;
	wire [2:0] w_n743_38;
	wire [2:0] w_n743_39;
	wire [2:0] w_n743_40;
	wire [2:0] w_n743_41;
	wire [2:0] w_n743_42;
	wire [2:0] w_n743_43;
	wire [2:0] w_n743_44;
	wire [2:0] w_n743_45;
	wire [2:0] w_n743_46;
	wire [2:0] w_n743_47;
	wire [2:0] w_n743_48;
	wire [2:0] w_n743_49;
	wire [2:0] w_n743_50;
	wire [2:0] w_n743_51;
	wire [2:0] w_n743_52;
	wire [2:0] w_n743_53;
	wire [2:0] w_n743_54;
	wire [2:0] w_n743_55;
	wire [2:0] w_n743_56;
	wire [2:0] w_n743_57;
	wire [2:0] w_n743_58;
	wire [2:0] w_n743_59;
	wire [2:0] w_n743_60;
	wire [2:0] w_n743_61;
	wire [2:0] w_n743_62;
	wire [2:0] w_n743_63;
	wire [2:0] w_n743_64;
	wire [2:0] w_n743_65;
	wire [2:0] w_n743_66;
	wire [2:0] w_n743_67;
	wire [2:0] w_n743_68;
	wire [2:0] w_n743_69;
	wire [2:0] w_n743_70;
	wire [2:0] w_n745_0;
	wire [1:0] w_n746_0;
	wire [2:0] w_n753_0;
	wire [1:0] w_n754_0;
	wire [1:0] w_n757_0;
	wire [1:0] w_n762_0;
	wire [2:0] w_n764_0;
	wire [1:0] w_n765_0;
	wire [2:0] w_n769_0;
	wire [2:0] w_n772_0;
	wire [1:0] w_n773_0;
	wire [2:0] w_n777_0;
	wire [2:0] w_n779_0;
	wire [1:0] w_n780_0;
	wire [2:0] w_n784_0;
	wire [2:0] w_n787_0;
	wire [1:0] w_n788_0;
	wire [2:0] w_n792_0;
	wire [2:0] w_n794_0;
	wire [1:0] w_n795_0;
	wire [2:0] w_n799_0;
	wire [2:0] w_n802_0;
	wire [2:0] w_n805_0;
	wire [1:0] w_n805_1;
	wire [2:0] w_n806_0;
	wire [1:0] w_n808_0;
	wire [1:0] w_n809_0;
	wire [1:0] w_n816_0;
	wire [1:0] w_n817_0;
	wire [1:0] w_n819_0;
	wire [1:0] w_n834_0;
	wire [1:0] w_n838_0;
	wire [1:0] w_n859_0;
	wire [1:0] w_n860_0;
	wire [2:0] w_n863_0;
	wire [1:0] w_n864_0;
	wire [2:0] w_n865_0;
	wire [1:0] w_n865_1;
	wire [1:0] w_n866_0;
	wire [2:0] w_n867_0;
	wire [1:0] w_n868_0;
	wire [2:0] w_n870_0;
	wire [1:0] w_n871_0;
	wire [2:0] w_n876_0;
	wire [1:0] w_n876_1;
	wire [1:0] w_n881_0;
	wire [1:0] w_n882_0;
	wire [2:0] w_n884_0;
	wire [2:0] w_n884_1;
	wire [2:0] w_n884_2;
	wire [2:0] w_n884_3;
	wire [2:0] w_n884_4;
	wire [2:0] w_n884_5;
	wire [2:0] w_n884_6;
	wire [2:0] w_n884_7;
	wire [2:0] w_n884_8;
	wire [2:0] w_n884_9;
	wire [2:0] w_n884_10;
	wire [2:0] w_n884_11;
	wire [2:0] w_n884_12;
	wire [2:0] w_n884_13;
	wire [2:0] w_n884_14;
	wire [2:0] w_n884_15;
	wire [2:0] w_n884_16;
	wire [2:0] w_n884_17;
	wire [2:0] w_n884_18;
	wire [2:0] w_n884_19;
	wire [2:0] w_n884_20;
	wire [2:0] w_n884_21;
	wire [2:0] w_n884_22;
	wire [2:0] w_n884_23;
	wire [2:0] w_n884_24;
	wire [2:0] w_n884_25;
	wire [2:0] w_n884_26;
	wire [2:0] w_n884_27;
	wire [2:0] w_n884_28;
	wire [2:0] w_n884_29;
	wire [2:0] w_n884_30;
	wire [2:0] w_n884_31;
	wire [2:0] w_n884_32;
	wire [2:0] w_n884_33;
	wire [2:0] w_n884_34;
	wire [2:0] w_n884_35;
	wire [2:0] w_n884_36;
	wire [2:0] w_n884_37;
	wire [2:0] w_n884_38;
	wire [2:0] w_n884_39;
	wire [2:0] w_n884_40;
	wire [2:0] w_n884_41;
	wire [2:0] w_n884_42;
	wire [2:0] w_n884_43;
	wire [2:0] w_n884_44;
	wire [2:0] w_n884_45;
	wire [2:0] w_n884_46;
	wire [2:0] w_n884_47;
	wire [2:0] w_n884_48;
	wire [2:0] w_n884_49;
	wire [2:0] w_n884_50;
	wire [2:0] w_n884_51;
	wire [2:0] w_n884_52;
	wire [2:0] w_n884_53;
	wire [2:0] w_n884_54;
	wire [2:0] w_n884_55;
	wire [2:0] w_n884_56;
	wire [2:0] w_n884_57;
	wire [2:0] w_n884_58;
	wire [2:0] w_n884_59;
	wire [2:0] w_n884_60;
	wire [2:0] w_n884_61;
	wire [2:0] w_n884_62;
	wire [2:0] w_n884_63;
	wire [2:0] w_n884_64;
	wire [2:0] w_n884_65;
	wire [2:0] w_n884_66;
	wire [2:0] w_n884_67;
	wire [1:0] w_n886_0;
	wire [2:0] w_n888_0;
	wire [1:0] w_n889_0;
	wire [1:0] w_n891_0;
	wire [1:0] w_n896_0;
	wire [1:0] w_n897_0;
	wire [2:0] w_n899_0;
	wire [1:0] w_n900_0;
	wire [1:0] w_n904_0;
	wire [2:0] w_n906_0;
	wire [1:0] w_n907_0;
	wire [1:0] w_n911_0;
	wire [2:0] w_n913_0;
	wire [1:0] w_n914_0;
	wire [1:0] w_n918_0;
	wire [2:0] w_n920_0;
	wire [1:0] w_n921_0;
	wire [1:0] w_n925_0;
	wire [1:0] w_n926_0;
	wire [2:0] w_n928_0;
	wire [1:0] w_n929_0;
	wire [1:0] w_n933_0;
	wire [2:0] w_n935_0;
	wire [1:0] w_n936_0;
	wire [1:0] w_n958_0;
	wire [1:0] w_n962_0;
	wire [1:0] w_n966_0;
	wire [1:0] w_n973_0;
	wire [1:0] w_n979_0;
	wire [1:0] w_n981_0;
	wire [1:0] w_n982_0;
	wire [1:0] w_n985_0;
	wire [1:0] w_n989_0;
	wire [1:0] w_n991_0;
	wire [2:0] w_n992_0;
	wire [1:0] w_n997_0;
	wire [1:0] w_n1000_0;
	wire [1:0] w_n1004_0;
	wire [2:0] w_n1008_0;
	wire [2:0] w_n1008_1;
	wire [2:0] w_n1008_2;
	wire [2:0] w_n1008_3;
	wire [2:0] w_n1008_4;
	wire [2:0] w_n1008_5;
	wire [2:0] w_n1008_6;
	wire [2:0] w_n1008_7;
	wire [2:0] w_n1008_8;
	wire [2:0] w_n1008_9;
	wire [2:0] w_n1008_10;
	wire [2:0] w_n1008_11;
	wire [2:0] w_n1008_12;
	wire [2:0] w_n1008_13;
	wire [2:0] w_n1008_14;
	wire [2:0] w_n1008_15;
	wire [2:0] w_n1008_16;
	wire [2:0] w_n1008_17;
	wire [2:0] w_n1008_18;
	wire [2:0] w_n1008_19;
	wire [2:0] w_n1008_20;
	wire [2:0] w_n1008_21;
	wire [2:0] w_n1008_22;
	wire [2:0] w_n1008_23;
	wire [2:0] w_n1008_24;
	wire [2:0] w_n1008_25;
	wire [2:0] w_n1008_26;
	wire [2:0] w_n1008_27;
	wire [2:0] w_n1008_28;
	wire [2:0] w_n1008_29;
	wire [2:0] w_n1008_30;
	wire [2:0] w_n1008_31;
	wire [2:0] w_n1008_32;
	wire [2:0] w_n1008_33;
	wire [2:0] w_n1008_34;
	wire [2:0] w_n1008_35;
	wire [2:0] w_n1008_36;
	wire [2:0] w_n1008_37;
	wire [2:0] w_n1008_38;
	wire [2:0] w_n1008_39;
	wire [2:0] w_n1008_40;
	wire [2:0] w_n1008_41;
	wire [2:0] w_n1008_42;
	wire [2:0] w_n1008_43;
	wire [2:0] w_n1008_44;
	wire [2:0] w_n1008_45;
	wire [2:0] w_n1008_46;
	wire [2:0] w_n1008_47;
	wire [2:0] w_n1008_48;
	wire [2:0] w_n1008_49;
	wire [2:0] w_n1008_50;
	wire [2:0] w_n1008_51;
	wire [2:0] w_n1008_52;
	wire [2:0] w_n1008_53;
	wire [2:0] w_n1008_54;
	wire [2:0] w_n1008_55;
	wire [2:0] w_n1008_56;
	wire [2:0] w_n1008_57;
	wire [2:0] w_n1008_58;
	wire [2:0] w_n1008_59;
	wire [2:0] w_n1008_60;
	wire [2:0] w_n1008_61;
	wire [2:0] w_n1008_62;
	wire [2:0] w_n1008_63;
	wire [2:0] w_n1008_64;
	wire [2:0] w_n1008_65;
	wire [2:0] w_n1008_66;
	wire [2:0] w_n1008_67;
	wire [2:0] w_n1008_68;
	wire [2:0] w_n1008_69;
	wire [1:0] w_n1008_70;
	wire [2:0] w_n1010_0;
	wire [2:0] w_n1010_1;
	wire [1:0] w_n1011_0;
	wire [2:0] w_n1012_0;
	wire [1:0] w_n1013_0;
	wire [2:0] w_n1015_0;
	wire [1:0] w_n1016_0;
	wire [2:0] w_n1023_0;
	wire [1:0] w_n1024_0;
	wire [1:0] w_n1027_0;
	wire [1:0] w_n1028_0;
	wire [2:0] w_n1033_0;
	wire [2:0] w_n1035_0;
	wire [1:0] w_n1036_0;
	wire [2:0] w_n1040_0;
	wire [2:0] w_n1042_0;
	wire [1:0] w_n1043_0;
	wire [2:0] w_n1047_0;
	wire [2:0] w_n1049_0;
	wire [1:0] w_n1050_0;
	wire [2:0] w_n1054_0;
	wire [2:0] w_n1057_0;
	wire [1:0] w_n1058_0;
	wire [2:0] w_n1062_0;
	wire [2:0] w_n1065_0;
	wire [1:0] w_n1066_0;
	wire [2:0] w_n1070_0;
	wire [2:0] w_n1073_0;
	wire [1:0] w_n1074_0;
	wire [2:0] w_n1078_0;
	wire [2:0] w_n1080_0;
	wire [1:0] w_n1081_0;
	wire [1:0] w_n1085_0;
	wire [1:0] w_n1086_0;
	wire [2:0] w_n1088_0;
	wire [1:0] w_n1088_1;
	wire [2:0] w_n1091_0;
	wire [1:0] w_n1091_1;
	wire [1:0] w_n1092_0;
	wire [1:0] w_n1096_0;
	wire [1:0] w_n1097_0;
	wire [1:0] w_n1101_0;
	wire [1:0] w_n1104_0;
	wire [2:0] w_n1108_0;
	wire [1:0] w_n1108_1;
	wire [1:0] w_n1109_0;
	wire [2:0] w_n1110_0;
	wire [1:0] w_n1111_0;
	wire [2:0] w_n1113_0;
	wire [1:0] w_n1114_0;
	wire [1:0] w_n1119_0;
	wire [1:0] w_n1134_0;
	wire [1:0] w_n1169_0;
	wire [1:0] w_n1172_0;
	wire [2:0] w_n1173_0;
	wire [2:0] w_n1173_1;
	wire [2:0] w_n1173_2;
	wire [2:0] w_n1173_3;
	wire [2:0] w_n1173_4;
	wire [2:0] w_n1173_5;
	wire [2:0] w_n1173_6;
	wire [2:0] w_n1173_7;
	wire [2:0] w_n1173_8;
	wire [2:0] w_n1173_9;
	wire [2:0] w_n1173_10;
	wire [2:0] w_n1173_11;
	wire [2:0] w_n1173_12;
	wire [2:0] w_n1173_13;
	wire [2:0] w_n1173_14;
	wire [2:0] w_n1173_15;
	wire [2:0] w_n1173_16;
	wire [2:0] w_n1173_17;
	wire [2:0] w_n1173_18;
	wire [2:0] w_n1173_19;
	wire [2:0] w_n1173_20;
	wire [2:0] w_n1173_21;
	wire [2:0] w_n1173_22;
	wire [2:0] w_n1173_23;
	wire [2:0] w_n1173_24;
	wire [2:0] w_n1173_25;
	wire [2:0] w_n1173_26;
	wire [2:0] w_n1173_27;
	wire [2:0] w_n1173_28;
	wire [2:0] w_n1173_29;
	wire [2:0] w_n1173_30;
	wire [2:0] w_n1173_31;
	wire [2:0] w_n1173_32;
	wire [2:0] w_n1173_33;
	wire [2:0] w_n1173_34;
	wire [2:0] w_n1173_35;
	wire [2:0] w_n1173_36;
	wire [2:0] w_n1173_37;
	wire [2:0] w_n1173_38;
	wire [2:0] w_n1173_39;
	wire [2:0] w_n1173_40;
	wire [2:0] w_n1173_41;
	wire [2:0] w_n1173_42;
	wire [2:0] w_n1173_43;
	wire [2:0] w_n1173_44;
	wire [2:0] w_n1173_45;
	wire [2:0] w_n1173_46;
	wire [2:0] w_n1173_47;
	wire [2:0] w_n1173_48;
	wire [2:0] w_n1173_49;
	wire [2:0] w_n1173_50;
	wire [2:0] w_n1173_51;
	wire [2:0] w_n1173_52;
	wire [2:0] w_n1173_53;
	wire [2:0] w_n1173_54;
	wire [2:0] w_n1173_55;
	wire [2:0] w_n1173_56;
	wire [2:0] w_n1173_57;
	wire [2:0] w_n1173_58;
	wire [2:0] w_n1173_59;
	wire [2:0] w_n1173_60;
	wire [2:0] w_n1173_61;
	wire [2:0] w_n1173_62;
	wire [2:0] w_n1173_63;
	wire [2:0] w_n1173_64;
	wire [1:0] w_n1175_0;
	wire [2:0] w_n1177_0;
	wire [1:0] w_n1178_0;
	wire [1:0] w_n1180_0;
	wire [1:0] w_n1185_0;
	wire [1:0] w_n1186_0;
	wire [2:0] w_n1188_0;
	wire [1:0] w_n1189_0;
	wire [1:0] w_n1193_0;
	wire [2:0] w_n1195_0;
	wire [1:0] w_n1196_0;
	wire [1:0] w_n1200_0;
	wire [1:0] w_n1201_0;
	wire [2:0] w_n1203_0;
	wire [1:0] w_n1204_0;
	wire [1:0] w_n1208_0;
	wire [1:0] w_n1209_0;
	wire [2:0] w_n1211_0;
	wire [1:0] w_n1212_0;
	wire [1:0] w_n1216_0;
	wire [1:0] w_n1217_0;
	wire [2:0] w_n1219_0;
	wire [1:0] w_n1220_0;
	wire [1:0] w_n1224_0;
	wire [2:0] w_n1226_0;
	wire [1:0] w_n1227_0;
	wire [1:0] w_n1231_0;
	wire [2:0] w_n1233_0;
	wire [1:0] w_n1234_0;
	wire [1:0] w_n1238_0;
	wire [2:0] w_n1240_0;
	wire [1:0] w_n1241_0;
	wire [1:0] w_n1245_0;
	wire [1:0] w_n1246_0;
	wire [1:0] w_n1248_0;
	wire [1:0] w_n1251_0;
	wire [1:0] w_n1252_0;
	wire [2:0] w_n1253_0;
	wire [1:0] w_n1253_1;
	wire [2:0] w_n1254_0;
	wire [1:0] w_n1279_0;
	wire [1:0] w_n1292_0;
	wire [1:0] w_n1296_0;
	wire [1:0] w_n1300_0;
	wire [1:0] w_n1305_0;
	wire [1:0] w_n1306_0;
	wire [1:0] w_n1307_0;
	wire [1:0] w_n1309_0;
	wire [1:0] w_n1311_0;
	wire [1:0] w_n1314_0;
	wire [1:0] w_n1315_0;
	wire [1:0] w_n1316_0;
	wire [2:0] w_n1319_0;
	wire [2:0] w_n1319_1;
	wire [1:0] w_n1320_0;
	wire [2:0] w_n1321_0;
	wire [1:0] w_n1322_0;
	wire [1:0] w_n1325_0;
	wire [1:0] w_n1330_0;
	wire [2:0] w_n1332_0;
	wire [2:0] w_n1332_1;
	wire [2:0] w_n1332_2;
	wire [2:0] w_n1332_3;
	wire [2:0] w_n1332_4;
	wire [2:0] w_n1332_5;
	wire [2:0] w_n1332_6;
	wire [2:0] w_n1332_7;
	wire [2:0] w_n1332_8;
	wire [2:0] w_n1332_9;
	wire [2:0] w_n1332_10;
	wire [2:0] w_n1332_11;
	wire [2:0] w_n1332_12;
	wire [2:0] w_n1332_13;
	wire [2:0] w_n1332_14;
	wire [2:0] w_n1332_15;
	wire [2:0] w_n1332_16;
	wire [2:0] w_n1332_17;
	wire [2:0] w_n1332_18;
	wire [2:0] w_n1332_19;
	wire [2:0] w_n1332_20;
	wire [2:0] w_n1332_21;
	wire [2:0] w_n1332_22;
	wire [2:0] w_n1332_23;
	wire [2:0] w_n1332_24;
	wire [2:0] w_n1332_25;
	wire [2:0] w_n1332_26;
	wire [2:0] w_n1332_27;
	wire [2:0] w_n1332_28;
	wire [2:0] w_n1332_29;
	wire [2:0] w_n1332_30;
	wire [2:0] w_n1332_31;
	wire [2:0] w_n1332_32;
	wire [2:0] w_n1332_33;
	wire [2:0] w_n1332_34;
	wire [2:0] w_n1332_35;
	wire [2:0] w_n1332_36;
	wire [2:0] w_n1332_37;
	wire [2:0] w_n1332_38;
	wire [2:0] w_n1332_39;
	wire [2:0] w_n1332_40;
	wire [2:0] w_n1332_41;
	wire [2:0] w_n1332_42;
	wire [2:0] w_n1332_43;
	wire [2:0] w_n1332_44;
	wire [2:0] w_n1332_45;
	wire [2:0] w_n1332_46;
	wire [2:0] w_n1332_47;
	wire [2:0] w_n1332_48;
	wire [2:0] w_n1332_49;
	wire [2:0] w_n1332_50;
	wire [2:0] w_n1332_51;
	wire [2:0] w_n1332_52;
	wire [2:0] w_n1332_53;
	wire [2:0] w_n1332_54;
	wire [2:0] w_n1332_55;
	wire [2:0] w_n1332_56;
	wire [2:0] w_n1332_57;
	wire [2:0] w_n1332_58;
	wire [2:0] w_n1332_59;
	wire [2:0] w_n1332_60;
	wire [2:0] w_n1332_61;
	wire [2:0] w_n1332_62;
	wire [2:0] w_n1332_63;
	wire [2:0] w_n1332_64;
	wire [2:0] w_n1332_65;
	wire [2:0] w_n1332_66;
	wire [2:0] w_n1332_67;
	wire [2:0] w_n1334_0;
	wire [1:0] w_n1335_0;
	wire [2:0] w_n1342_0;
	wire [1:0] w_n1343_0;
	wire [1:0] w_n1346_0;
	wire [2:0] w_n1351_0;
	wire [2:0] w_n1353_0;
	wire [1:0] w_n1354_0;
	wire [2:0] w_n1358_0;
	wire [2:0] w_n1360_0;
	wire [1:0] w_n1361_0;
	wire [2:0] w_n1365_0;
	wire [2:0] w_n1367_0;
	wire [1:0] w_n1368_0;
	wire [2:0] w_n1372_0;
	wire [2:0] w_n1375_0;
	wire [1:0] w_n1376_0;
	wire [2:0] w_n1380_0;
	wire [2:0] w_n1382_0;
	wire [1:0] w_n1383_0;
	wire [2:0] w_n1387_0;
	wire [2:0] w_n1389_0;
	wire [1:0] w_n1390_0;
	wire [2:0] w_n1394_0;
	wire [2:0] w_n1396_0;
	wire [1:0] w_n1397_0;
	wire [2:0] w_n1401_0;
	wire [2:0] w_n1404_0;
	wire [1:0] w_n1405_0;
	wire [2:0] w_n1409_0;
	wire [2:0] w_n1412_0;
	wire [1:0] w_n1413_0;
	wire [1:0] w_n1417_0;
	wire [1:0] w_n1418_0;
	wire [2:0] w_n1420_0;
	wire [1:0] w_n1420_1;
	wire [2:0] w_n1423_0;
	wire [2:0] w_n1423_1;
	wire [1:0] w_n1424_0;
	wire [1:0] w_n1426_0;
	wire [1:0] w_n1434_0;
	wire [1:0] w_n1435_0;
	wire [2:0] w_n1440_0;
	wire [1:0] w_n1440_1;
	wire [1:0] w_n1441_0;
	wire [2:0] w_n1442_0;
	wire [1:0] w_n1443_0;
	wire [2:0] w_n1445_0;
	wire [1:0] w_n1446_0;
	wire [1:0] w_n1451_0;
	wire [1:0] w_n1470_0;
	wire [1:0] w_n1513_0;
	wire [1:0] w_n1514_0;
	wire [2:0] w_n1516_0;
	wire [2:0] w_n1516_1;
	wire [2:0] w_n1516_2;
	wire [2:0] w_n1516_3;
	wire [2:0] w_n1516_4;
	wire [2:0] w_n1516_5;
	wire [2:0] w_n1516_6;
	wire [2:0] w_n1516_7;
	wire [2:0] w_n1516_8;
	wire [2:0] w_n1516_9;
	wire [2:0] w_n1516_10;
	wire [2:0] w_n1516_11;
	wire [2:0] w_n1516_12;
	wire [2:0] w_n1516_13;
	wire [2:0] w_n1516_14;
	wire [2:0] w_n1516_15;
	wire [2:0] w_n1516_16;
	wire [2:0] w_n1516_17;
	wire [2:0] w_n1516_18;
	wire [2:0] w_n1516_19;
	wire [2:0] w_n1516_20;
	wire [2:0] w_n1516_21;
	wire [2:0] w_n1516_22;
	wire [2:0] w_n1516_23;
	wire [2:0] w_n1516_24;
	wire [2:0] w_n1516_25;
	wire [2:0] w_n1516_26;
	wire [2:0] w_n1516_27;
	wire [2:0] w_n1516_28;
	wire [2:0] w_n1516_29;
	wire [2:0] w_n1516_30;
	wire [2:0] w_n1516_31;
	wire [2:0] w_n1516_32;
	wire [2:0] w_n1516_33;
	wire [2:0] w_n1516_34;
	wire [2:0] w_n1516_35;
	wire [2:0] w_n1516_36;
	wire [2:0] w_n1516_37;
	wire [2:0] w_n1516_38;
	wire [2:0] w_n1516_39;
	wire [2:0] w_n1516_40;
	wire [2:0] w_n1516_41;
	wire [2:0] w_n1516_42;
	wire [2:0] w_n1516_43;
	wire [2:0] w_n1516_44;
	wire [2:0] w_n1516_45;
	wire [2:0] w_n1516_46;
	wire [2:0] w_n1516_47;
	wire [2:0] w_n1516_48;
	wire [2:0] w_n1516_49;
	wire [2:0] w_n1516_50;
	wire [2:0] w_n1516_51;
	wire [2:0] w_n1516_52;
	wire [2:0] w_n1516_53;
	wire [2:0] w_n1516_54;
	wire [2:0] w_n1516_55;
	wire [2:0] w_n1516_56;
	wire [2:0] w_n1516_57;
	wire [2:0] w_n1516_58;
	wire [2:0] w_n1516_59;
	wire [2:0] w_n1516_60;
	wire [2:0] w_n1516_61;
	wire [2:0] w_n1516_62;
	wire [1:0] w_n1518_0;
	wire [2:0] w_n1520_0;
	wire [1:0] w_n1521_0;
	wire [1:0] w_n1523_0;
	wire [2:0] w_n1528_0;
	wire [2:0] w_n1531_0;
	wire [1:0] w_n1532_0;
	wire [1:0] w_n1536_0;
	wire [2:0] w_n1538_0;
	wire [1:0] w_n1539_0;
	wire [1:0] w_n1543_0;
	wire [1:0] w_n1544_0;
	wire [2:0] w_n1546_0;
	wire [1:0] w_n1547_0;
	wire [1:0] w_n1551_0;
	wire [1:0] w_n1552_0;
	wire [2:0] w_n1554_0;
	wire [1:0] w_n1555_0;
	wire [1:0] w_n1559_0;
	wire [1:0] w_n1560_0;
	wire [2:0] w_n1562_0;
	wire [1:0] w_n1563_0;
	wire [1:0] w_n1567_0;
	wire [2:0] w_n1569_0;
	wire [1:0] w_n1570_0;
	wire [1:0] w_n1574_0;
	wire [1:0] w_n1575_0;
	wire [2:0] w_n1577_0;
	wire [1:0] w_n1578_0;
	wire [1:0] w_n1582_0;
	wire [1:0] w_n1583_0;
	wire [2:0] w_n1585_0;
	wire [1:0] w_n1586_0;
	wire [1:0] w_n1590_0;
	wire [1:0] w_n1591_0;
	wire [2:0] w_n1593_0;
	wire [1:0] w_n1594_0;
	wire [1:0] w_n1598_0;
	wire [2:0] w_n1600_0;
	wire [1:0] w_n1601_0;
	wire [1:0] w_n1627_0;
	wire [1:0] w_n1640_0;
	wire [1:0] w_n1653_0;
	wire [2:0] w_n1659_0;
	wire [2:0] w_n1662_0;
	wire [2:0] w_n1665_0;
	wire [1:0] w_n1665_1;
	wire [1:0] w_n1666_0;
	wire [1:0] w_n1667_0;
	wire [1:0] w_n1669_0;
	wire [1:0] w_n1671_0;
	wire [1:0] w_n1672_0;
	wire [2:0] w_n1673_0;
	wire [1:0] w_n1677_0;
	wire [1:0] w_n1678_0;
	wire [2:0] w_n1681_0;
	wire [2:0] w_n1681_1;
	wire [1:0] w_n1682_0;
	wire [2:0] w_n1683_0;
	wire [1:0] w_n1684_0;
	wire [1:0] w_n1688_0;
	wire [1:0] w_n1689_0;
	wire [1:0] w_n1690_0;
	wire [2:0] w_n1695_0;
	wire [2:0] w_n1699_0;
	wire [2:0] w_n1699_1;
	wire [2:0] w_n1699_2;
	wire [2:0] w_n1699_3;
	wire [2:0] w_n1699_4;
	wire [2:0] w_n1699_5;
	wire [2:0] w_n1699_6;
	wire [2:0] w_n1699_7;
	wire [2:0] w_n1699_8;
	wire [2:0] w_n1699_9;
	wire [2:0] w_n1699_10;
	wire [2:0] w_n1699_11;
	wire [2:0] w_n1699_12;
	wire [2:0] w_n1699_13;
	wire [2:0] w_n1699_14;
	wire [2:0] w_n1699_15;
	wire [2:0] w_n1699_16;
	wire [2:0] w_n1699_17;
	wire [2:0] w_n1699_18;
	wire [2:0] w_n1699_19;
	wire [2:0] w_n1699_20;
	wire [2:0] w_n1699_21;
	wire [2:0] w_n1699_22;
	wire [2:0] w_n1699_23;
	wire [2:0] w_n1699_24;
	wire [2:0] w_n1699_25;
	wire [2:0] w_n1699_26;
	wire [2:0] w_n1699_27;
	wire [2:0] w_n1699_28;
	wire [2:0] w_n1699_29;
	wire [2:0] w_n1699_30;
	wire [2:0] w_n1699_31;
	wire [2:0] w_n1699_32;
	wire [2:0] w_n1699_33;
	wire [2:0] w_n1699_34;
	wire [2:0] w_n1699_35;
	wire [2:0] w_n1699_36;
	wire [2:0] w_n1699_37;
	wire [2:0] w_n1699_38;
	wire [2:0] w_n1699_39;
	wire [2:0] w_n1699_40;
	wire [2:0] w_n1699_41;
	wire [2:0] w_n1699_42;
	wire [2:0] w_n1699_43;
	wire [2:0] w_n1699_44;
	wire [2:0] w_n1699_45;
	wire [2:0] w_n1699_46;
	wire [2:0] w_n1699_47;
	wire [2:0] w_n1699_48;
	wire [2:0] w_n1699_49;
	wire [2:0] w_n1699_50;
	wire [2:0] w_n1699_51;
	wire [2:0] w_n1699_52;
	wire [2:0] w_n1699_53;
	wire [2:0] w_n1699_54;
	wire [2:0] w_n1699_55;
	wire [2:0] w_n1699_56;
	wire [2:0] w_n1699_57;
	wire [2:0] w_n1699_58;
	wire [2:0] w_n1699_59;
	wire [2:0] w_n1699_60;
	wire [2:0] w_n1699_61;
	wire [2:0] w_n1699_62;
	wire [2:0] w_n1699_63;
	wire [2:0] w_n1699_64;
	wire [2:0] w_n1699_65;
	wire [2:0] w_n1699_66;
	wire [1:0] w_n1699_67;
	wire [2:0] w_n1701_0;
	wire [1:0] w_n1702_0;
	wire [2:0] w_n1709_0;
	wire [1:0] w_n1710_0;
	wire [1:0] w_n1713_0;
	wire [2:0] w_n1718_0;
	wire [2:0] w_n1720_0;
	wire [1:0] w_n1721_0;
	wire [2:0] w_n1725_0;
	wire [2:0] w_n1727_0;
	wire [1:0] w_n1728_0;
	wire [2:0] w_n1732_0;
	wire [2:0] w_n1735_0;
	wire [1:0] w_n1736_0;
	wire [2:0] w_n1740_0;
	wire [2:0] w_n1743_0;
	wire [1:0] w_n1744_0;
	wire [2:0] w_n1748_0;
	wire [2:0] w_n1750_0;
	wire [1:0] w_n1751_0;
	wire [2:0] w_n1755_0;
	wire [2:0] w_n1757_0;
	wire [1:0] w_n1758_0;
	wire [2:0] w_n1762_0;
	wire [2:0] w_n1764_0;
	wire [1:0] w_n1765_0;
	wire [2:0] w_n1769_0;
	wire [2:0] w_n1772_0;
	wire [1:0] w_n1773_0;
	wire [2:0] w_n1777_0;
	wire [2:0] w_n1779_0;
	wire [1:0] w_n1780_0;
	wire [2:0] w_n1784_0;
	wire [2:0] w_n1786_0;
	wire [1:0] w_n1787_0;
	wire [2:0] w_n1791_0;
	wire [2:0] w_n1793_0;
	wire [1:0] w_n1794_0;
	wire [2:0] w_n1798_0;
	wire [2:0] w_n1801_0;
	wire [2:0] w_n1804_0;
	wire [1:0] w_n1804_1;
	wire [2:0] w_n1805_0;
	wire [1:0] w_n1809_0;
	wire [1:0] w_n1810_0;
	wire [1:0] w_n1812_0;
	wire [1:0] w_n1813_0;
	wire [1:0] w_n1817_0;
	wire [1:0] w_n1819_0;
	wire [1:0] w_n1839_0;
	wire [1:0] w_n1887_0;
	wire [1:0] w_n1888_0;
	wire [2:0] w_n1891_0;
	wire [2:0] w_n1894_0;
	wire [1:0] w_n1894_1;
	wire [1:0] w_n1895_0;
	wire [2:0] w_n1896_0;
	wire [1:0] w_n1897_0;
	wire [2:0] w_n1898_0;
	wire [1:0] w_n1899_0;
	wire [2:0] w_n1904_0;
	wire [1:0] w_n1904_1;
	wire [1:0] w_n1908_0;
	wire [1:0] w_n1911_0;
	wire [2:0] w_n1912_0;
	wire [2:0] w_n1912_1;
	wire [2:0] w_n1912_2;
	wire [2:0] w_n1912_3;
	wire [2:0] w_n1912_4;
	wire [2:0] w_n1912_5;
	wire [2:0] w_n1912_6;
	wire [2:0] w_n1912_7;
	wire [2:0] w_n1912_8;
	wire [2:0] w_n1912_9;
	wire [2:0] w_n1912_10;
	wire [2:0] w_n1912_11;
	wire [2:0] w_n1912_12;
	wire [2:0] w_n1912_13;
	wire [2:0] w_n1912_14;
	wire [2:0] w_n1912_15;
	wire [2:0] w_n1912_16;
	wire [2:0] w_n1912_17;
	wire [2:0] w_n1912_18;
	wire [2:0] w_n1912_19;
	wire [2:0] w_n1912_20;
	wire [2:0] w_n1912_21;
	wire [2:0] w_n1912_22;
	wire [2:0] w_n1912_23;
	wire [2:0] w_n1912_24;
	wire [2:0] w_n1912_25;
	wire [2:0] w_n1912_26;
	wire [2:0] w_n1912_27;
	wire [2:0] w_n1912_28;
	wire [2:0] w_n1912_29;
	wire [2:0] w_n1912_30;
	wire [2:0] w_n1912_31;
	wire [2:0] w_n1912_32;
	wire [2:0] w_n1912_33;
	wire [2:0] w_n1912_34;
	wire [2:0] w_n1912_35;
	wire [2:0] w_n1912_36;
	wire [2:0] w_n1912_37;
	wire [2:0] w_n1912_38;
	wire [2:0] w_n1912_39;
	wire [2:0] w_n1912_40;
	wire [2:0] w_n1912_41;
	wire [2:0] w_n1912_42;
	wire [2:0] w_n1912_43;
	wire [2:0] w_n1912_44;
	wire [2:0] w_n1912_45;
	wire [2:0] w_n1912_46;
	wire [2:0] w_n1912_47;
	wire [2:0] w_n1912_48;
	wire [2:0] w_n1912_49;
	wire [2:0] w_n1912_50;
	wire [2:0] w_n1912_51;
	wire [2:0] w_n1912_52;
	wire [2:0] w_n1912_53;
	wire [2:0] w_n1912_54;
	wire [2:0] w_n1912_55;
	wire [2:0] w_n1912_56;
	wire [2:0] w_n1912_57;
	wire [2:0] w_n1912_58;
	wire [2:0] w_n1912_59;
	wire [1:0] w_n1912_60;
	wire [2:0] w_n1916_0;
	wire [1:0] w_n1917_0;
	wire [1:0] w_n1919_0;
	wire [1:0] w_n1924_0;
	wire [1:0] w_n1925_0;
	wire [2:0] w_n1927_0;
	wire [1:0] w_n1928_0;
	wire [1:0] w_n1932_0;
	wire [2:0] w_n1934_0;
	wire [1:0] w_n1935_0;
	wire [1:0] w_n1939_0;
	wire [1:0] w_n1940_0;
	wire [2:0] w_n1942_0;
	wire [1:0] w_n1943_0;
	wire [1:0] w_n1947_0;
	wire [1:0] w_n1948_0;
	wire [2:0] w_n1950_0;
	wire [1:0] w_n1951_0;
	wire [1:0] w_n1955_0;
	wire [2:0] w_n1957_0;
	wire [1:0] w_n1958_0;
	wire [1:0] w_n1962_0;
	wire [2:0] w_n1964_0;
	wire [1:0] w_n1965_0;
	wire [1:0] w_n1969_0;
	wire [1:0] w_n1970_0;
	wire [2:0] w_n1972_0;
	wire [1:0] w_n1973_0;
	wire [1:0] w_n1977_0;
	wire [1:0] w_n1978_0;
	wire [2:0] w_n1980_0;
	wire [1:0] w_n1981_0;
	wire [2:0] w_n1985_0;
	wire [2:0] w_n1988_0;
	wire [1:0] w_n1989_0;
	wire [1:0] w_n1993_0;
	wire [2:0] w_n1995_0;
	wire [1:0] w_n1996_0;
	wire [1:0] w_n2000_0;
	wire [1:0] w_n2001_0;
	wire [2:0] w_n2003_0;
	wire [1:0] w_n2004_0;
	wire [1:0] w_n2008_0;
	wire [1:0] w_n2009_0;
	wire [2:0] w_n2011_0;
	wire [1:0] w_n2012_0;
	wire [1:0] w_n2033_0;
	wire [1:0] w_n2040_0;
	wire [1:0] w_n2050_0;
	wire [1:0] w_n2054_0;
	wire [1:0] w_n2067_0;
	wire [1:0] w_n2079_0;
	wire [1:0] w_n2081_0;
	wire [1:0] w_n2082_0;
	wire [1:0] w_n2085_0;
	wire [1:0] w_n2089_0;
	wire [1:0] w_n2091_0;
	wire [2:0] w_n2092_0;
	wire [1:0] w_n2097_0;
	wire [1:0] w_n2100_0;
	wire [1:0] w_n2104_0;
	wire [2:0] w_n2108_0;
	wire [2:0] w_n2108_1;
	wire [2:0] w_n2108_2;
	wire [2:0] w_n2108_3;
	wire [2:0] w_n2108_4;
	wire [2:0] w_n2108_5;
	wire [2:0] w_n2108_6;
	wire [2:0] w_n2108_7;
	wire [2:0] w_n2108_8;
	wire [2:0] w_n2108_9;
	wire [2:0] w_n2108_10;
	wire [2:0] w_n2108_11;
	wire [2:0] w_n2108_12;
	wire [2:0] w_n2108_13;
	wire [2:0] w_n2108_14;
	wire [2:0] w_n2108_15;
	wire [2:0] w_n2108_16;
	wire [2:0] w_n2108_17;
	wire [2:0] w_n2108_18;
	wire [2:0] w_n2108_19;
	wire [2:0] w_n2108_20;
	wire [2:0] w_n2108_21;
	wire [2:0] w_n2108_22;
	wire [2:0] w_n2108_23;
	wire [2:0] w_n2108_24;
	wire [2:0] w_n2108_25;
	wire [2:0] w_n2108_26;
	wire [2:0] w_n2108_27;
	wire [2:0] w_n2108_28;
	wire [2:0] w_n2108_29;
	wire [2:0] w_n2108_30;
	wire [2:0] w_n2108_31;
	wire [2:0] w_n2108_32;
	wire [2:0] w_n2108_33;
	wire [2:0] w_n2108_34;
	wire [2:0] w_n2108_35;
	wire [2:0] w_n2108_36;
	wire [2:0] w_n2108_37;
	wire [2:0] w_n2108_38;
	wire [2:0] w_n2108_39;
	wire [2:0] w_n2108_40;
	wire [2:0] w_n2108_41;
	wire [2:0] w_n2108_42;
	wire [2:0] w_n2108_43;
	wire [2:0] w_n2108_44;
	wire [2:0] w_n2108_45;
	wire [2:0] w_n2108_46;
	wire [2:0] w_n2108_47;
	wire [2:0] w_n2108_48;
	wire [2:0] w_n2108_49;
	wire [2:0] w_n2108_50;
	wire [2:0] w_n2108_51;
	wire [2:0] w_n2108_52;
	wire [2:0] w_n2108_53;
	wire [2:0] w_n2108_54;
	wire [2:0] w_n2108_55;
	wire [2:0] w_n2108_56;
	wire [2:0] w_n2108_57;
	wire [2:0] w_n2108_58;
	wire [2:0] w_n2108_59;
	wire [2:0] w_n2108_60;
	wire [2:0] w_n2108_61;
	wire [2:0] w_n2108_62;
	wire [2:0] w_n2108_63;
	wire [2:0] w_n2108_64;
	wire [1:0] w_n2108_65;
	wire [2:0] w_n2110_0;
	wire [2:0] w_n2110_1;
	wire [1:0] w_n2111_0;
	wire [2:0] w_n2112_0;
	wire [1:0] w_n2113_0;
	wire [2:0] w_n2115_0;
	wire [1:0] w_n2116_0;
	wire [2:0] w_n2123_0;
	wire [1:0] w_n2124_0;
	wire [1:0] w_n2127_0;
	wire [1:0] w_n2128_0;
	wire [2:0] w_n2133_0;
	wire [2:0] w_n2135_0;
	wire [1:0] w_n2136_0;
	wire [2:0] w_n2140_0;
	wire [2:0] w_n2143_0;
	wire [1:0] w_n2144_0;
	wire [2:0] w_n2148_0;
	wire [2:0] w_n2150_0;
	wire [1:0] w_n2151_0;
	wire [2:0] w_n2155_0;
	wire [2:0] w_n2158_0;
	wire [1:0] w_n2159_0;
	wire [2:0] w_n2163_0;
	wire [2:0] w_n2165_0;
	wire [1:0] w_n2166_0;
	wire [2:0] w_n2170_0;
	wire [2:0] w_n2172_0;
	wire [1:0] w_n2173_0;
	wire [2:0] w_n2177_0;
	wire [2:0] w_n2180_0;
	wire [1:0] w_n2181_0;
	wire [2:0] w_n2185_0;
	wire [2:0] w_n2188_0;
	wire [1:0] w_n2189_0;
	wire [2:0] w_n2193_0;
	wire [2:0] w_n2195_0;
	wire [1:0] w_n2196_0;
	wire [1:0] w_n2200_0;
	wire [2:0] w_n2202_0;
	wire [1:0] w_n2203_0;
	wire [2:0] w_n2207_0;
	wire [2:0] w_n2210_0;
	wire [1:0] w_n2211_0;
	wire [2:0] w_n2215_0;
	wire [2:0] w_n2218_0;
	wire [1:0] w_n2219_0;
	wire [2:0] w_n2223_0;
	wire [2:0] w_n2225_0;
	wire [1:0] w_n2226_0;
	wire [2:0] w_n2230_0;
	wire [2:0] w_n2232_0;
	wire [2:0] w_n2235_0;
	wire [1:0] w_n2235_1;
	wire [2:0] w_n2236_0;
	wire [1:0] w_n2238_0;
	wire [1:0] w_n2240_0;
	wire [1:0] w_n2246_0;
	wire [1:0] w_n2247_0;
	wire [1:0] w_n2249_0;
	wire [2:0] w_n2252_0;
	wire [1:0] w_n2252_1;
	wire [1:0] w_n2253_0;
	wire [2:0] w_n2254_0;
	wire [1:0] w_n2255_0;
	wire [2:0] w_n2257_0;
	wire [1:0] w_n2258_0;
	wire [2:0] w_n2263_0;
	wire [1:0] w_n2263_1;
	wire [1:0] w_n2285_0;
	wire [1:0] w_n2321_0;
	wire [1:0] w_n2339_0;
	wire [1:0] w_n2342_0;
	wire [1:0] w_n2343_0;
	wire [2:0] w_n2345_0;
	wire [2:0] w_n2345_1;
	wire [2:0] w_n2345_2;
	wire [2:0] w_n2345_3;
	wire [2:0] w_n2345_4;
	wire [2:0] w_n2345_5;
	wire [2:0] w_n2345_6;
	wire [2:0] w_n2345_7;
	wire [2:0] w_n2345_8;
	wire [2:0] w_n2345_9;
	wire [2:0] w_n2345_10;
	wire [2:0] w_n2345_11;
	wire [2:0] w_n2345_12;
	wire [2:0] w_n2345_13;
	wire [2:0] w_n2345_14;
	wire [2:0] w_n2345_15;
	wire [2:0] w_n2345_16;
	wire [2:0] w_n2345_17;
	wire [2:0] w_n2345_18;
	wire [2:0] w_n2345_19;
	wire [2:0] w_n2345_20;
	wire [2:0] w_n2345_21;
	wire [2:0] w_n2345_22;
	wire [2:0] w_n2345_23;
	wire [2:0] w_n2345_24;
	wire [2:0] w_n2345_25;
	wire [2:0] w_n2345_26;
	wire [2:0] w_n2345_27;
	wire [2:0] w_n2345_28;
	wire [2:0] w_n2345_29;
	wire [2:0] w_n2345_30;
	wire [2:0] w_n2345_31;
	wire [2:0] w_n2345_32;
	wire [2:0] w_n2345_33;
	wire [2:0] w_n2345_34;
	wire [2:0] w_n2345_35;
	wire [2:0] w_n2345_36;
	wire [2:0] w_n2345_37;
	wire [2:0] w_n2345_38;
	wire [2:0] w_n2345_39;
	wire [2:0] w_n2345_40;
	wire [2:0] w_n2345_41;
	wire [2:0] w_n2345_42;
	wire [2:0] w_n2345_43;
	wire [2:0] w_n2345_44;
	wire [2:0] w_n2345_45;
	wire [2:0] w_n2345_46;
	wire [2:0] w_n2345_47;
	wire [2:0] w_n2345_48;
	wire [2:0] w_n2345_49;
	wire [2:0] w_n2345_50;
	wire [2:0] w_n2345_51;
	wire [2:0] w_n2345_52;
	wire [2:0] w_n2345_53;
	wire [2:0] w_n2345_54;
	wire [2:0] w_n2345_55;
	wire [2:0] w_n2345_56;
	wire [2:0] w_n2345_57;
	wire [2:0] w_n2349_0;
	wire [1:0] w_n2350_0;
	wire [1:0] w_n2352_0;
	wire [1:0] w_n2357_0;
	wire [1:0] w_n2358_0;
	wire [2:0] w_n2360_0;
	wire [1:0] w_n2361_0;
	wire [1:0] w_n2365_0;
	wire [2:0] w_n2367_0;
	wire [1:0] w_n2368_0;
	wire [1:0] w_n2372_0;
	wire [1:0] w_n2373_0;
	wire [2:0] w_n2375_0;
	wire [1:0] w_n2376_0;
	wire [1:0] w_n2380_0;
	wire [2:0] w_n2382_0;
	wire [1:0] w_n2383_0;
	wire [1:0] w_n2387_0;
	wire [1:0] w_n2388_0;
	wire [2:0] w_n2390_0;
	wire [1:0] w_n2391_0;
	wire [1:0] w_n2395_0;
	wire [2:0] w_n2397_0;
	wire [1:0] w_n2398_0;
	wire [1:0] w_n2402_0;
	wire [1:0] w_n2403_0;
	wire [2:0] w_n2405_0;
	wire [1:0] w_n2406_0;
	wire [1:0] w_n2410_0;
	wire [1:0] w_n2411_0;
	wire [2:0] w_n2413_0;
	wire [1:0] w_n2414_0;
	wire [1:0] w_n2418_0;
	wire [2:0] w_n2420_0;
	wire [1:0] w_n2421_0;
	wire [1:0] w_n2425_0;
	wire [2:0] w_n2427_0;
	wire [1:0] w_n2428_0;
	wire [1:0] w_n2432_0;
	wire [1:0] w_n2433_0;
	wire [2:0] w_n2435_0;
	wire [1:0] w_n2436_0;
	wire [1:0] w_n2440_0;
	wire [2:0] w_n2442_0;
	wire [1:0] w_n2443_0;
	wire [1:0] w_n2447_0;
	wire [2:0] w_n2449_0;
	wire [1:0] w_n2450_0;
	wire [1:0] w_n2454_0;
	wire [2:0] w_n2456_0;
	wire [1:0] w_n2457_0;
	wire [2:0] w_n2461_0;
	wire [1:0] w_n2464_0;
	wire [1:0] w_n2467_0;
	wire [1:0] w_n2468_0;
	wire [2:0] w_n2469_0;
	wire [1:0] w_n2469_1;
	wire [2:0] w_n2470_0;
	wire [1:0] w_n2474_0;
	wire [1:0] w_n2475_0;
	wire [1:0] w_n2476_0;
	wire [1:0] w_n2499_0;
	wire [1:0] w_n2506_0;
	wire [1:0] w_n2513_0;
	wire [1:0] w_n2520_0;
	wire [1:0] w_n2530_0;
	wire [1:0] w_n2534_0;
	wire [1:0] w_n2541_0;
	wire [1:0] w_n2545_0;
	wire [1:0] w_n2549_0;
	wire [1:0] w_n2554_0;
	wire [1:0] w_n2555_0;
	wire [1:0] w_n2558_0;
	wire [1:0] w_n2559_0;
	wire [1:0] w_n2561_0;
	wire [1:0] w_n2565_0;
	wire [1:0] w_n2571_0;
	wire [2:0] w_n2572_0;
	wire [2:0] w_n2572_1;
	wire [2:0] w_n2572_2;
	wire [2:0] w_n2572_3;
	wire [2:0] w_n2572_4;
	wire [2:0] w_n2572_5;
	wire [2:0] w_n2572_6;
	wire [2:0] w_n2572_7;
	wire [2:0] w_n2572_8;
	wire [2:0] w_n2572_9;
	wire [2:0] w_n2572_10;
	wire [2:0] w_n2572_11;
	wire [2:0] w_n2572_12;
	wire [2:0] w_n2572_13;
	wire [2:0] w_n2572_14;
	wire [2:0] w_n2572_15;
	wire [2:0] w_n2572_16;
	wire [2:0] w_n2572_17;
	wire [2:0] w_n2572_18;
	wire [2:0] w_n2572_19;
	wire [2:0] w_n2572_20;
	wire [2:0] w_n2572_21;
	wire [2:0] w_n2572_22;
	wire [2:0] w_n2572_23;
	wire [2:0] w_n2572_24;
	wire [2:0] w_n2572_25;
	wire [2:0] w_n2572_26;
	wire [2:0] w_n2572_27;
	wire [2:0] w_n2572_28;
	wire [2:0] w_n2572_29;
	wire [2:0] w_n2572_30;
	wire [2:0] w_n2572_31;
	wire [2:0] w_n2572_32;
	wire [2:0] w_n2572_33;
	wire [2:0] w_n2572_34;
	wire [2:0] w_n2572_35;
	wire [2:0] w_n2572_36;
	wire [2:0] w_n2572_37;
	wire [2:0] w_n2572_38;
	wire [2:0] w_n2572_39;
	wire [2:0] w_n2572_40;
	wire [2:0] w_n2572_41;
	wire [2:0] w_n2572_42;
	wire [2:0] w_n2572_43;
	wire [2:0] w_n2572_44;
	wire [2:0] w_n2572_45;
	wire [2:0] w_n2572_46;
	wire [2:0] w_n2572_47;
	wire [2:0] w_n2572_48;
	wire [2:0] w_n2572_49;
	wire [2:0] w_n2572_50;
	wire [2:0] w_n2572_51;
	wire [2:0] w_n2572_52;
	wire [2:0] w_n2572_53;
	wire [2:0] w_n2572_54;
	wire [2:0] w_n2572_55;
	wire [2:0] w_n2572_56;
	wire [2:0] w_n2572_57;
	wire [2:0] w_n2572_58;
	wire [2:0] w_n2572_59;
	wire [2:0] w_n2572_60;
	wire [2:0] w_n2572_61;
	wire [2:0] w_n2572_62;
	wire [1:0] w_n2572_63;
	wire [1:0] w_n2575_0;
	wire [2:0] w_n2576_0;
	wire [2:0] w_n2578_0;
	wire [2:0] w_n2578_1;
	wire [1:0] w_n2579_0;
	wire [2:0] w_n2580_0;
	wire [1:0] w_n2581_0;
	wire [2:0] w_n2583_0;
	wire [1:0] w_n2584_0;
	wire [2:0] w_n2591_0;
	wire [1:0] w_n2592_0;
	wire [1:0] w_n2595_0;
	wire [2:0] w_n2600_0;
	wire [2:0] w_n2602_0;
	wire [1:0] w_n2603_0;
	wire [2:0] w_n2607_0;
	wire [2:0] w_n2610_0;
	wire [1:0] w_n2611_0;
	wire [2:0] w_n2615_0;
	wire [2:0] w_n2617_0;
	wire [1:0] w_n2618_0;
	wire [2:0] w_n2622_0;
	wire [2:0] w_n2625_0;
	wire [1:0] w_n2626_0;
	wire [2:0] w_n2630_0;
	wire [2:0] w_n2632_0;
	wire [1:0] w_n2633_0;
	wire [2:0] w_n2637_0;
	wire [2:0] w_n2640_0;
	wire [1:0] w_n2641_0;
	wire [2:0] w_n2645_0;
	wire [2:0] w_n2647_0;
	wire [1:0] w_n2648_0;
	wire [2:0] w_n2652_0;
	wire [2:0] w_n2655_0;
	wire [1:0] w_n2656_0;
	wire [2:0] w_n2660_0;
	wire [2:0] w_n2662_0;
	wire [1:0] w_n2663_0;
	wire [2:0] w_n2667_0;
	wire [2:0] w_n2669_0;
	wire [1:0] w_n2670_0;
	wire [2:0] w_n2674_0;
	wire [2:0] w_n2677_0;
	wire [1:0] w_n2678_0;
	wire [2:0] w_n2682_0;
	wire [2:0] w_n2685_0;
	wire [1:0] w_n2686_0;
	wire [2:0] w_n2690_0;
	wire [2:0] w_n2692_0;
	wire [1:0] w_n2693_0;
	wire [2:0] w_n2697_0;
	wire [2:0] w_n2700_0;
	wire [1:0] w_n2701_0;
	wire [2:0] w_n2705_0;
	wire [2:0] w_n2708_0;
	wire [1:0] w_n2709_0;
	wire [1:0] w_n2713_0;
	wire [1:0] w_n2714_0;
	wire [2:0] w_n2716_0;
	wire [2:0] w_n2717_0;
	wire [1:0] w_n2719_0;
	wire [1:0] w_n2720_0;
	wire [1:0] w_n2727_0;
	wire [1:0] w_n2728_0;
	wire [1:0] w_n2730_0;
	wire [2:0] w_n2734_0;
	wire [1:0] w_n2734_1;
	wire [1:0] w_n2735_0;
	wire [2:0] w_n2736_0;
	wire [1:0] w_n2737_0;
	wire [2:0] w_n2738_0;
	wire [1:0] w_n2739_0;
	wire [2:0] w_n2744_0;
	wire [1:0] w_n2744_1;
	wire [1:0] w_n2769_0;
	wire [1:0] w_n2827_0;
	wire [1:0] w_n2830_0;
	wire [1:0] w_n2831_0;
	wire [2:0] w_n2833_0;
	wire [2:0] w_n2833_1;
	wire [2:0] w_n2833_2;
	wire [2:0] w_n2833_3;
	wire [2:0] w_n2833_4;
	wire [2:0] w_n2833_5;
	wire [2:0] w_n2833_6;
	wire [2:0] w_n2833_7;
	wire [2:0] w_n2833_8;
	wire [2:0] w_n2833_9;
	wire [2:0] w_n2833_10;
	wire [2:0] w_n2833_11;
	wire [2:0] w_n2833_12;
	wire [2:0] w_n2833_13;
	wire [2:0] w_n2833_14;
	wire [2:0] w_n2833_15;
	wire [2:0] w_n2833_16;
	wire [2:0] w_n2833_17;
	wire [2:0] w_n2833_18;
	wire [2:0] w_n2833_19;
	wire [2:0] w_n2833_20;
	wire [2:0] w_n2833_21;
	wire [2:0] w_n2833_22;
	wire [2:0] w_n2833_23;
	wire [2:0] w_n2833_24;
	wire [2:0] w_n2833_25;
	wire [2:0] w_n2833_26;
	wire [2:0] w_n2833_27;
	wire [2:0] w_n2833_28;
	wire [2:0] w_n2833_29;
	wire [2:0] w_n2833_30;
	wire [2:0] w_n2833_31;
	wire [2:0] w_n2833_32;
	wire [2:0] w_n2833_33;
	wire [2:0] w_n2833_34;
	wire [2:0] w_n2833_35;
	wire [2:0] w_n2833_36;
	wire [2:0] w_n2833_37;
	wire [2:0] w_n2833_38;
	wire [2:0] w_n2833_39;
	wire [2:0] w_n2833_40;
	wire [2:0] w_n2833_41;
	wire [2:0] w_n2833_42;
	wire [2:0] w_n2833_43;
	wire [2:0] w_n2833_44;
	wire [2:0] w_n2833_45;
	wire [2:0] w_n2833_46;
	wire [2:0] w_n2833_47;
	wire [2:0] w_n2833_48;
	wire [2:0] w_n2833_49;
	wire [2:0] w_n2833_50;
	wire [2:0] w_n2833_51;
	wire [2:0] w_n2833_52;
	wire [2:0] w_n2833_53;
	wire [2:0] w_n2833_54;
	wire [1:0] w_n2833_55;
	wire [1:0] w_n2835_0;
	wire [2:0] w_n2837_0;
	wire [1:0] w_n2838_0;
	wire [1:0] w_n2840_0;
	wire [1:0] w_n2845_0;
	wire [1:0] w_n2846_0;
	wire [2:0] w_n2848_0;
	wire [1:0] w_n2849_0;
	wire [1:0] w_n2853_0;
	wire [2:0] w_n2855_0;
	wire [1:0] w_n2856_0;
	wire [1:0] w_n2860_0;
	wire [1:0] w_n2861_0;
	wire [2:0] w_n2863_0;
	wire [1:0] w_n2864_0;
	wire [1:0] w_n2868_0;
	wire [2:0] w_n2870_0;
	wire [1:0] w_n2871_0;
	wire [1:0] w_n2875_0;
	wire [1:0] w_n2876_0;
	wire [2:0] w_n2878_0;
	wire [1:0] w_n2879_0;
	wire [1:0] w_n2883_0;
	wire [2:0] w_n2885_0;
	wire [1:0] w_n2886_0;
	wire [1:0] w_n2890_0;
	wire [1:0] w_n2891_0;
	wire [2:0] w_n2893_0;
	wire [1:0] w_n2894_0;
	wire [1:0] w_n2898_0;
	wire [2:0] w_n2900_0;
	wire [1:0] w_n2901_0;
	wire [1:0] w_n2905_0;
	wire [1:0] w_n2906_0;
	wire [2:0] w_n2908_0;
	wire [1:0] w_n2909_0;
	wire [1:0] w_n2913_0;
	wire [2:0] w_n2915_0;
	wire [1:0] w_n2916_0;
	wire [1:0] w_n2920_0;
	wire [1:0] w_n2921_0;
	wire [2:0] w_n2923_0;
	wire [1:0] w_n2924_0;
	wire [1:0] w_n2928_0;
	wire [1:0] w_n2929_0;
	wire [2:0] w_n2931_0;
	wire [1:0] w_n2932_0;
	wire [1:0] w_n2936_0;
	wire [2:0] w_n2938_0;
	wire [1:0] w_n2939_0;
	wire [1:0] w_n2943_0;
	wire [2:0] w_n2945_0;
	wire [1:0] w_n2946_0;
	wire [1:0] w_n2950_0;
	wire [1:0] w_n2951_0;
	wire [2:0] w_n2953_0;
	wire [1:0] w_n2954_0;
	wire [1:0] w_n2958_0;
	wire [2:0] w_n2960_0;
	wire [1:0] w_n2961_0;
	wire [2:0] w_n2965_0;
	wire [1:0] w_n2967_0;
	wire [2:0] w_n2970_0;
	wire [1:0] w_n2971_0;
	wire [2:0] w_n2972_0;
	wire [2:0] w_n2973_0;
	wire [1:0] w_n2977_0;
	wire [1:0] w_n2978_0;
	wire [1:0] w_n2979_0;
	wire [1:0] w_n3011_0;
	wire [1:0] w_n3018_0;
	wire [1:0] w_n3025_0;
	wire [1:0] w_n3032_0;
	wire [1:0] w_n3039_0;
	wire [1:0] w_n3049_0;
	wire [1:0] w_n3053_0;
	wire [1:0] w_n3060_0;
	wire [1:0] w_n3066_0;
	wire [1:0] w_n3067_0;
	wire [1:0] w_n3070_0;
	wire [1:0] w_n3071_0;
	wire [1:0] w_n3073_0;
	wire [2:0] w_n3075_0;
	wire [2:0] w_n3075_1;
	wire [1:0] w_n3076_0;
	wire [2:0] w_n3077_0;
	wire [1:0] w_n3078_0;
	wire [1:0] w_n3082_0;
	wire [1:0] w_n3088_0;
	wire [2:0] w_n3089_0;
	wire [2:0] w_n3089_1;
	wire [2:0] w_n3089_2;
	wire [2:0] w_n3089_3;
	wire [2:0] w_n3089_4;
	wire [2:0] w_n3089_5;
	wire [2:0] w_n3089_6;
	wire [2:0] w_n3089_7;
	wire [2:0] w_n3089_8;
	wire [2:0] w_n3089_9;
	wire [2:0] w_n3089_10;
	wire [2:0] w_n3089_11;
	wire [2:0] w_n3089_12;
	wire [2:0] w_n3089_13;
	wire [2:0] w_n3089_14;
	wire [2:0] w_n3089_15;
	wire [2:0] w_n3089_16;
	wire [2:0] w_n3089_17;
	wire [2:0] w_n3089_18;
	wire [2:0] w_n3089_19;
	wire [2:0] w_n3089_20;
	wire [2:0] w_n3089_21;
	wire [2:0] w_n3089_22;
	wire [2:0] w_n3089_23;
	wire [2:0] w_n3089_24;
	wire [2:0] w_n3089_25;
	wire [2:0] w_n3089_26;
	wire [2:0] w_n3089_27;
	wire [2:0] w_n3089_28;
	wire [2:0] w_n3089_29;
	wire [2:0] w_n3089_30;
	wire [2:0] w_n3089_31;
	wire [2:0] w_n3089_32;
	wire [2:0] w_n3089_33;
	wire [2:0] w_n3089_34;
	wire [2:0] w_n3089_35;
	wire [2:0] w_n3089_36;
	wire [2:0] w_n3089_37;
	wire [2:0] w_n3089_38;
	wire [2:0] w_n3089_39;
	wire [2:0] w_n3089_40;
	wire [2:0] w_n3089_41;
	wire [2:0] w_n3089_42;
	wire [2:0] w_n3089_43;
	wire [2:0] w_n3089_44;
	wire [2:0] w_n3089_45;
	wire [2:0] w_n3089_46;
	wire [2:0] w_n3089_47;
	wire [2:0] w_n3089_48;
	wire [2:0] w_n3089_49;
	wire [2:0] w_n3089_50;
	wire [2:0] w_n3089_51;
	wire [2:0] w_n3089_52;
	wire [2:0] w_n3089_53;
	wire [2:0] w_n3089_54;
	wire [2:0] w_n3089_55;
	wire [2:0] w_n3089_56;
	wire [2:0] w_n3089_57;
	wire [2:0] w_n3089_58;
	wire [2:0] w_n3089_59;
	wire [2:0] w_n3089_60;
	wire [2:0] w_n3089_61;
	wire [1:0] w_n3089_62;
	wire [2:0] w_n3091_0;
	wire [1:0] w_n3092_0;
	wire [2:0] w_n3099_0;
	wire [1:0] w_n3100_0;
	wire [1:0] w_n3103_0;
	wire [1:0] w_n3108_0;
	wire [2:0] w_n3110_0;
	wire [1:0] w_n3111_0;
	wire [2:0] w_n3115_0;
	wire [2:0] w_n3117_0;
	wire [1:0] w_n3118_0;
	wire [2:0] w_n3122_0;
	wire [2:0] w_n3124_0;
	wire [1:0] w_n3125_0;
	wire [2:0] w_n3129_0;
	wire [2:0] w_n3132_0;
	wire [1:0] w_n3133_0;
	wire [2:0] w_n3137_0;
	wire [2:0] w_n3139_0;
	wire [1:0] w_n3140_0;
	wire [2:0] w_n3144_0;
	wire [2:0] w_n3147_0;
	wire [1:0] w_n3148_0;
	wire [2:0] w_n3152_0;
	wire [2:0] w_n3154_0;
	wire [1:0] w_n3155_0;
	wire [2:0] w_n3159_0;
	wire [2:0] w_n3162_0;
	wire [1:0] w_n3163_0;
	wire [2:0] w_n3167_0;
	wire [2:0] w_n3169_0;
	wire [1:0] w_n3170_0;
	wire [2:0] w_n3174_0;
	wire [2:0] w_n3177_0;
	wire [1:0] w_n3178_0;
	wire [2:0] w_n3182_0;
	wire [2:0] w_n3184_0;
	wire [1:0] w_n3185_0;
	wire [2:0] w_n3189_0;
	wire [2:0] w_n3192_0;
	wire [1:0] w_n3193_0;
	wire [2:0] w_n3197_0;
	wire [2:0] w_n3199_0;
	wire [1:0] w_n3200_0;
	wire [2:0] w_n3204_0;
	wire [2:0] w_n3206_0;
	wire [1:0] w_n3207_0;
	wire [2:0] w_n3211_0;
	wire [2:0] w_n3214_0;
	wire [1:0] w_n3215_0;
	wire [2:0] w_n3219_0;
	wire [2:0] w_n3222_0;
	wire [1:0] w_n3223_0;
	wire [2:0] w_n3227_0;
	wire [2:0] w_n3229_0;
	wire [1:0] w_n3230_0;
	wire [1:0] w_n3234_0;
	wire [1:0] w_n3235_0;
	wire [2:0] w_n3237_0;
	wire [1:0] w_n3237_1;
	wire [2:0] w_n3240_0;
	wire [1:0] w_n3240_1;
	wire [1:0] w_n3241_0;
	wire [1:0] w_n3245_0;
	wire [1:0] w_n3246_0;
	wire [1:0] w_n3250_0;
	wire [1:0] w_n3253_0;
	wire [2:0] w_n3258_0;
	wire [1:0] w_n3258_1;
	wire [1:0] w_n3259_0;
	wire [2:0] w_n3260_0;
	wire [1:0] w_n3261_0;
	wire [2:0] w_n3262_0;
	wire [1:0] w_n3263_0;
	wire [1:0] w_n3268_0;
	wire [1:0] w_n3293_0;
	wire [1:0] w_n3297_0;
	wire [1:0] w_n3364_0;
	wire [1:0] w_n3367_0;
	wire [2:0] w_n3368_0;
	wire [2:0] w_n3368_1;
	wire [2:0] w_n3368_2;
	wire [2:0] w_n3368_3;
	wire [2:0] w_n3368_4;
	wire [2:0] w_n3368_5;
	wire [2:0] w_n3368_6;
	wire [2:0] w_n3368_7;
	wire [2:0] w_n3368_8;
	wire [2:0] w_n3368_9;
	wire [2:0] w_n3368_10;
	wire [2:0] w_n3368_11;
	wire [2:0] w_n3368_12;
	wire [2:0] w_n3368_13;
	wire [2:0] w_n3368_14;
	wire [2:0] w_n3368_15;
	wire [2:0] w_n3368_16;
	wire [2:0] w_n3368_17;
	wire [2:0] w_n3368_18;
	wire [2:0] w_n3368_19;
	wire [2:0] w_n3368_20;
	wire [2:0] w_n3368_21;
	wire [2:0] w_n3368_22;
	wire [2:0] w_n3368_23;
	wire [2:0] w_n3368_24;
	wire [2:0] w_n3368_25;
	wire [2:0] w_n3368_26;
	wire [2:0] w_n3368_27;
	wire [2:0] w_n3368_28;
	wire [2:0] w_n3368_29;
	wire [2:0] w_n3368_30;
	wire [2:0] w_n3368_31;
	wire [2:0] w_n3368_32;
	wire [2:0] w_n3368_33;
	wire [2:0] w_n3368_34;
	wire [2:0] w_n3368_35;
	wire [2:0] w_n3368_36;
	wire [2:0] w_n3368_37;
	wire [2:0] w_n3368_38;
	wire [2:0] w_n3368_39;
	wire [2:0] w_n3368_40;
	wire [2:0] w_n3368_41;
	wire [2:0] w_n3368_42;
	wire [2:0] w_n3368_43;
	wire [2:0] w_n3368_44;
	wire [2:0] w_n3368_45;
	wire [2:0] w_n3368_46;
	wire [2:0] w_n3368_47;
	wire [2:0] w_n3368_48;
	wire [2:0] w_n3368_49;
	wire [2:0] w_n3368_50;
	wire [2:0] w_n3368_51;
	wire [1:0] w_n3368_52;
	wire [2:0] w_n3372_0;
	wire [1:0] w_n3373_0;
	wire [1:0] w_n3375_0;
	wire [1:0] w_n3380_0;
	wire [1:0] w_n3381_0;
	wire [2:0] w_n3383_0;
	wire [1:0] w_n3384_0;
	wire [1:0] w_n3388_0;
	wire [2:0] w_n3390_0;
	wire [1:0] w_n3391_0;
	wire [1:0] w_n3395_0;
	wire [2:0] w_n3397_0;
	wire [1:0] w_n3398_0;
	wire [1:0] w_n3402_0;
	wire [1:0] w_n3403_0;
	wire [2:0] w_n3405_0;
	wire [1:0] w_n3406_0;
	wire [1:0] w_n3410_0;
	wire [1:0] w_n3411_0;
	wire [2:0] w_n3413_0;
	wire [1:0] w_n3414_0;
	wire [1:0] w_n3418_0;
	wire [2:0] w_n3420_0;
	wire [1:0] w_n3421_0;
	wire [1:0] w_n3425_0;
	wire [1:0] w_n3426_0;
	wire [2:0] w_n3428_0;
	wire [1:0] w_n3429_0;
	wire [1:0] w_n3433_0;
	wire [2:0] w_n3435_0;
	wire [1:0] w_n3436_0;
	wire [1:0] w_n3440_0;
	wire [1:0] w_n3441_0;
	wire [2:0] w_n3443_0;
	wire [1:0] w_n3444_0;
	wire [1:0] w_n3448_0;
	wire [2:0] w_n3450_0;
	wire [1:0] w_n3451_0;
	wire [1:0] w_n3455_0;
	wire [1:0] w_n3456_0;
	wire [2:0] w_n3458_0;
	wire [1:0] w_n3459_0;
	wire [1:0] w_n3463_0;
	wire [2:0] w_n3465_0;
	wire [1:0] w_n3466_0;
	wire [1:0] w_n3470_0;
	wire [1:0] w_n3471_0;
	wire [2:0] w_n3473_0;
	wire [1:0] w_n3474_0;
	wire [1:0] w_n3478_0;
	wire [2:0] w_n3480_0;
	wire [1:0] w_n3481_0;
	wire [1:0] w_n3485_0;
	wire [1:0] w_n3486_0;
	wire [2:0] w_n3488_0;
	wire [1:0] w_n3489_0;
	wire [1:0] w_n3493_0;
	wire [1:0] w_n3494_0;
	wire [2:0] w_n3496_0;
	wire [1:0] w_n3497_0;
	wire [1:0] w_n3501_0;
	wire [2:0] w_n3503_0;
	wire [1:0] w_n3504_0;
	wire [1:0] w_n3508_0;
	wire [2:0] w_n3510_0;
	wire [1:0] w_n3511_0;
	wire [2:0] w_n3515_0;
	wire [1:0] w_n3518_0;
	wire [2:0] w_n3521_0;
	wire [1:0] w_n3522_0;
	wire [2:0] w_n3523_0;
	wire [1:0] w_n3523_1;
	wire [2:0] w_n3524_0;
	wire [1:0] w_n3552_0;
	wire [1:0] w_n3559_0;
	wire [1:0] w_n3563_0;
	wire [1:0] w_n3573_0;
	wire [1:0] w_n3580_0;
	wire [1:0] w_n3587_0;
	wire [1:0] w_n3594_0;
	wire [1:0] w_n3601_0;
	wire [1:0] w_n3611_0;
	wire [1:0] w_n3615_0;
	wire [1:0] w_n3620_0;
	wire [1:0] w_n3621_0;
	wire [1:0] w_n3622_0;
	wire [1:0] w_n3624_0;
	wire [1:0] w_n3626_0;
	wire [1:0] w_n3629_0;
	wire [1:0] w_n3630_0;
	wire [1:0] w_n3631_0;
	wire [1:0] w_n3635_0;
	wire [1:0] w_n3640_0;
	wire [2:0] w_n3642_0;
	wire [2:0] w_n3642_1;
	wire [2:0] w_n3642_2;
	wire [2:0] w_n3642_3;
	wire [2:0] w_n3642_4;
	wire [2:0] w_n3642_5;
	wire [2:0] w_n3642_6;
	wire [2:0] w_n3642_7;
	wire [2:0] w_n3642_8;
	wire [2:0] w_n3642_9;
	wire [2:0] w_n3642_10;
	wire [2:0] w_n3642_11;
	wire [2:0] w_n3642_12;
	wire [2:0] w_n3642_13;
	wire [2:0] w_n3642_14;
	wire [2:0] w_n3642_15;
	wire [2:0] w_n3642_16;
	wire [2:0] w_n3642_17;
	wire [2:0] w_n3642_18;
	wire [2:0] w_n3642_19;
	wire [2:0] w_n3642_20;
	wire [2:0] w_n3642_21;
	wire [2:0] w_n3642_22;
	wire [2:0] w_n3642_23;
	wire [2:0] w_n3642_24;
	wire [2:0] w_n3642_25;
	wire [2:0] w_n3642_26;
	wire [2:0] w_n3642_27;
	wire [2:0] w_n3642_28;
	wire [2:0] w_n3642_29;
	wire [2:0] w_n3642_30;
	wire [2:0] w_n3642_31;
	wire [2:0] w_n3642_32;
	wire [2:0] w_n3642_33;
	wire [2:0] w_n3642_34;
	wire [2:0] w_n3642_35;
	wire [2:0] w_n3642_36;
	wire [2:0] w_n3642_37;
	wire [2:0] w_n3642_38;
	wire [2:0] w_n3642_39;
	wire [2:0] w_n3642_40;
	wire [2:0] w_n3642_41;
	wire [2:0] w_n3642_42;
	wire [2:0] w_n3642_43;
	wire [2:0] w_n3642_44;
	wire [2:0] w_n3642_45;
	wire [2:0] w_n3642_46;
	wire [2:0] w_n3642_47;
	wire [2:0] w_n3642_48;
	wire [2:0] w_n3642_49;
	wire [2:0] w_n3642_50;
	wire [2:0] w_n3642_51;
	wire [2:0] w_n3642_52;
	wire [2:0] w_n3642_53;
	wire [2:0] w_n3642_54;
	wire [2:0] w_n3642_55;
	wire [2:0] w_n3642_56;
	wire [2:0] w_n3642_57;
	wire [2:0] w_n3642_58;
	wire [2:0] w_n3642_59;
	wire [2:0] w_n3642_60;
	wire [1:0] w_n3645_0;
	wire [2:0] w_n3646_0;
	wire [1:0] w_n3646_1;
	wire [2:0] w_n3648_0;
	wire [2:0] w_n3648_1;
	wire [1:0] w_n3649_0;
	wire [2:0] w_n3650_0;
	wire [1:0] w_n3651_0;
	wire [2:0] w_n3653_0;
	wire [1:0] w_n3654_0;
	wire [2:0] w_n3661_0;
	wire [1:0] w_n3662_0;
	wire [1:0] w_n3665_0;
	wire [2:0] w_n3670_0;
	wire [2:0] w_n3672_0;
	wire [1:0] w_n3673_0;
	wire [2:0] w_n3677_0;
	wire [2:0] w_n3680_0;
	wire [1:0] w_n3681_0;
	wire [2:0] w_n3685_0;
	wire [2:0] w_n3687_0;
	wire [1:0] w_n3688_0;
	wire [2:0] w_n3692_0;
	wire [2:0] w_n3695_0;
	wire [1:0] w_n3696_0;
	wire [2:0] w_n3700_0;
	wire [2:0] w_n3703_0;
	wire [1:0] w_n3704_0;
	wire [2:0] w_n3708_0;
	wire [2:0] w_n3710_0;
	wire [1:0] w_n3711_0;
	wire [2:0] w_n3715_0;
	wire [2:0] w_n3717_0;
	wire [1:0] w_n3718_0;
	wire [2:0] w_n3722_0;
	wire [2:0] w_n3725_0;
	wire [1:0] w_n3726_0;
	wire [2:0] w_n3730_0;
	wire [2:0] w_n3732_0;
	wire [1:0] w_n3733_0;
	wire [2:0] w_n3737_0;
	wire [2:0] w_n3740_0;
	wire [1:0] w_n3741_0;
	wire [2:0] w_n3745_0;
	wire [2:0] w_n3747_0;
	wire [1:0] w_n3748_0;
	wire [2:0] w_n3752_0;
	wire [2:0] w_n3755_0;
	wire [1:0] w_n3756_0;
	wire [2:0] w_n3760_0;
	wire [2:0] w_n3762_0;
	wire [1:0] w_n3763_0;
	wire [2:0] w_n3767_0;
	wire [2:0] w_n3770_0;
	wire [1:0] w_n3771_0;
	wire [2:0] w_n3775_0;
	wire [2:0] w_n3777_0;
	wire [1:0] w_n3778_0;
	wire [2:0] w_n3782_0;
	wire [2:0] w_n3785_0;
	wire [1:0] w_n3786_0;
	wire [2:0] w_n3790_0;
	wire [2:0] w_n3792_0;
	wire [1:0] w_n3793_0;
	wire [2:0] w_n3797_0;
	wire [2:0] w_n3799_0;
	wire [1:0] w_n3800_0;
	wire [2:0] w_n3804_0;
	wire [2:0] w_n3807_0;
	wire [1:0] w_n3808_0;
	wire [2:0] w_n3812_0;
	wire [2:0] w_n3815_0;
	wire [1:0] w_n3815_1;
	wire [1:0] w_n3816_0;
	wire [1:0] w_n3820_0;
	wire [1:0] w_n3821_0;
	wire [1:0] w_n3823_0;
	wire [1:0] w_n3828_0;
	wire [2:0] w_n3834_0;
	wire [2:0] w_n3835_0;
	wire [2:0] w_n3837_0;
	wire [1:0] w_n3837_1;
	wire [1:0] w_n3838_0;
	wire [2:0] w_n3839_0;
	wire [1:0] w_n3840_0;
	wire [2:0] w_n3841_0;
	wire [1:0] w_n3842_0;
	wire [1:0] w_n3847_0;
	wire [1:0] w_n3875_0;
	wire [1:0] w_n3951_0;
	wire [1:0] w_n3954_0;
	wire [2:0] w_n3955_0;
	wire [2:0] w_n3955_1;
	wire [2:0] w_n3955_2;
	wire [2:0] w_n3955_3;
	wire [2:0] w_n3955_4;
	wire [2:0] w_n3955_5;
	wire [2:0] w_n3955_6;
	wire [2:0] w_n3955_7;
	wire [2:0] w_n3955_8;
	wire [2:0] w_n3955_9;
	wire [2:0] w_n3955_10;
	wire [2:0] w_n3955_11;
	wire [2:0] w_n3955_12;
	wire [2:0] w_n3955_13;
	wire [2:0] w_n3955_14;
	wire [2:0] w_n3955_15;
	wire [2:0] w_n3955_16;
	wire [2:0] w_n3955_17;
	wire [2:0] w_n3955_18;
	wire [2:0] w_n3955_19;
	wire [2:0] w_n3955_20;
	wire [2:0] w_n3955_21;
	wire [2:0] w_n3955_22;
	wire [2:0] w_n3955_23;
	wire [2:0] w_n3955_24;
	wire [2:0] w_n3955_25;
	wire [2:0] w_n3955_26;
	wire [2:0] w_n3955_27;
	wire [2:0] w_n3955_28;
	wire [2:0] w_n3955_29;
	wire [2:0] w_n3955_30;
	wire [2:0] w_n3955_31;
	wire [2:0] w_n3955_32;
	wire [2:0] w_n3955_33;
	wire [2:0] w_n3955_34;
	wire [2:0] w_n3955_35;
	wire [2:0] w_n3955_36;
	wire [2:0] w_n3955_37;
	wire [2:0] w_n3955_38;
	wire [2:0] w_n3955_39;
	wire [2:0] w_n3955_40;
	wire [2:0] w_n3955_41;
	wire [2:0] w_n3955_42;
	wire [2:0] w_n3955_43;
	wire [2:0] w_n3955_44;
	wire [2:0] w_n3955_45;
	wire [2:0] w_n3955_46;
	wire [2:0] w_n3955_47;
	wire [2:0] w_n3955_48;
	wire [2:0] w_n3955_49;
	wire [1:0] w_n3955_50;
	wire [1:0] w_n3957_0;
	wire [2:0] w_n3959_0;
	wire [1:0] w_n3960_0;
	wire [1:0] w_n3962_0;
	wire [1:0] w_n3967_0;
	wire [1:0] w_n3968_0;
	wire [2:0] w_n3970_0;
	wire [1:0] w_n3971_0;
	wire [1:0] w_n3975_0;
	wire [2:0] w_n3977_0;
	wire [1:0] w_n3978_0;
	wire [1:0] w_n3982_0;
	wire [1:0] w_n3983_0;
	wire [2:0] w_n3985_0;
	wire [1:0] w_n3986_0;
	wire [1:0] w_n3990_0;
	wire [2:0] w_n3992_0;
	wire [1:0] w_n3993_0;
	wire [1:0] w_n3997_0;
	wire [1:0] w_n3998_0;
	wire [2:0] w_n4000_0;
	wire [1:0] w_n4001_0;
	wire [1:0] w_n4005_0;
	wire [2:0] w_n4007_0;
	wire [1:0] w_n4008_0;
	wire [1:0] w_n4012_0;
	wire [2:0] w_n4014_0;
	wire [1:0] w_n4015_0;
	wire [1:0] w_n4019_0;
	wire [1:0] w_n4020_0;
	wire [2:0] w_n4022_0;
	wire [1:0] w_n4023_0;
	wire [1:0] w_n4027_0;
	wire [1:0] w_n4028_0;
	wire [2:0] w_n4030_0;
	wire [1:0] w_n4031_0;
	wire [1:0] w_n4035_0;
	wire [2:0] w_n4037_0;
	wire [1:0] w_n4038_0;
	wire [1:0] w_n4042_0;
	wire [1:0] w_n4043_0;
	wire [2:0] w_n4045_0;
	wire [1:0] w_n4046_0;
	wire [1:0] w_n4050_0;
	wire [2:0] w_n4052_0;
	wire [1:0] w_n4053_0;
	wire [1:0] w_n4057_0;
	wire [1:0] w_n4058_0;
	wire [2:0] w_n4060_0;
	wire [1:0] w_n4061_0;
	wire [1:0] w_n4065_0;
	wire [2:0] w_n4067_0;
	wire [1:0] w_n4068_0;
	wire [1:0] w_n4072_0;
	wire [1:0] w_n4073_0;
	wire [2:0] w_n4075_0;
	wire [1:0] w_n4076_0;
	wire [1:0] w_n4080_0;
	wire [2:0] w_n4082_0;
	wire [1:0] w_n4083_0;
	wire [1:0] w_n4087_0;
	wire [1:0] w_n4088_0;
	wire [2:0] w_n4090_0;
	wire [1:0] w_n4091_0;
	wire [1:0] w_n4095_0;
	wire [2:0] w_n4097_0;
	wire [1:0] w_n4098_0;
	wire [1:0] w_n4102_0;
	wire [1:0] w_n4103_0;
	wire [2:0] w_n4105_0;
	wire [1:0] w_n4106_0;
	wire [1:0] w_n4110_0;
	wire [1:0] w_n4111_0;
	wire [2:0] w_n4113_0;
	wire [1:0] w_n4114_0;
	wire [1:0] w_n4150_0;
	wire [1:0] w_n4157_0;
	wire [1:0] w_n4164_0;
	wire [1:0] w_n4168_0;
	wire [1:0] w_n4178_0;
	wire [1:0] w_n4185_0;
	wire [1:0] w_n4192_0;
	wire [1:0] w_n4199_0;
	wire [1:0] w_n4206_0;
	wire [1:0] w_n4218_0;
	wire [1:0] w_n4219_0;
	wire [2:0] w_n4221_0;
	wire [1:0] w_n4222_0;
	wire [1:0] w_n4223_0;
	wire [1:0] w_n4225_0;
	wire [1:0] w_n4227_0;
	wire [1:0] w_n4228_0;
	wire [2:0] w_n4229_0;
	wire [1:0] w_n4233_0;
	wire [1:0] w_n4234_0;
	wire [1:0] w_n4239_0;
	wire [1:0] w_n4240_0;
	wire [2:0] w_n4245_0;
	wire [2:0] w_n4249_0;
	wire [2:0] w_n4249_1;
	wire [2:0] w_n4249_2;
	wire [2:0] w_n4249_3;
	wire [2:0] w_n4249_4;
	wire [2:0] w_n4249_5;
	wire [2:0] w_n4249_6;
	wire [2:0] w_n4249_7;
	wire [2:0] w_n4249_8;
	wire [2:0] w_n4249_9;
	wire [2:0] w_n4249_10;
	wire [2:0] w_n4249_11;
	wire [2:0] w_n4249_12;
	wire [2:0] w_n4249_13;
	wire [2:0] w_n4249_14;
	wire [2:0] w_n4249_15;
	wire [2:0] w_n4249_16;
	wire [2:0] w_n4249_17;
	wire [2:0] w_n4249_18;
	wire [2:0] w_n4249_19;
	wire [2:0] w_n4249_20;
	wire [2:0] w_n4249_21;
	wire [2:0] w_n4249_22;
	wire [2:0] w_n4249_23;
	wire [2:0] w_n4249_24;
	wire [2:0] w_n4249_25;
	wire [2:0] w_n4249_26;
	wire [2:0] w_n4249_27;
	wire [2:0] w_n4249_28;
	wire [2:0] w_n4249_29;
	wire [2:0] w_n4249_30;
	wire [2:0] w_n4249_31;
	wire [2:0] w_n4249_32;
	wire [2:0] w_n4249_33;
	wire [2:0] w_n4249_34;
	wire [2:0] w_n4249_35;
	wire [2:0] w_n4249_36;
	wire [2:0] w_n4249_37;
	wire [2:0] w_n4249_38;
	wire [2:0] w_n4249_39;
	wire [2:0] w_n4249_40;
	wire [2:0] w_n4249_41;
	wire [2:0] w_n4249_42;
	wire [2:0] w_n4249_43;
	wire [2:0] w_n4249_44;
	wire [2:0] w_n4249_45;
	wire [2:0] w_n4249_46;
	wire [2:0] w_n4249_47;
	wire [2:0] w_n4249_48;
	wire [2:0] w_n4249_49;
	wire [2:0] w_n4249_50;
	wire [2:0] w_n4249_51;
	wire [2:0] w_n4249_52;
	wire [2:0] w_n4249_53;
	wire [2:0] w_n4249_54;
	wire [2:0] w_n4249_55;
	wire [2:0] w_n4249_56;
	wire [2:0] w_n4249_57;
	wire [2:0] w_n4249_58;
	wire [2:0] w_n4249_59;
	wire [1:0] w_n4252_0;
	wire [2:0] w_n4253_0;
	wire [2:0] w_n4255_0;
	wire [2:0] w_n4255_1;
	wire [1:0] w_n4256_0;
	wire [2:0] w_n4257_0;
	wire [1:0] w_n4258_0;
	wire [2:0] w_n4260_0;
	wire [1:0] w_n4261_0;
	wire [1:0] w_n4266_0;
	wire [2:0] w_n4268_0;
	wire [1:0] w_n4269_0;
	wire [1:0] w_n4272_0;
	wire [2:0] w_n4277_0;
	wire [2:0] w_n4279_0;
	wire [1:0] w_n4280_0;
	wire [2:0] w_n4284_0;
	wire [2:0] w_n4286_0;
	wire [1:0] w_n4287_0;
	wire [2:0] w_n4291_0;
	wire [2:0] w_n4293_0;
	wire [1:0] w_n4294_0;
	wire [2:0] w_n4298_0;
	wire [2:0] w_n4301_0;
	wire [1:0] w_n4302_0;
	wire [2:0] w_n4306_0;
	wire [2:0] w_n4308_0;
	wire [1:0] w_n4309_0;
	wire [2:0] w_n4313_0;
	wire [2:0] w_n4316_0;
	wire [1:0] w_n4317_0;
	wire [2:0] w_n4321_0;
	wire [2:0] w_n4323_0;
	wire [1:0] w_n4324_0;
	wire [2:0] w_n4328_0;
	wire [2:0] w_n4331_0;
	wire [1:0] w_n4332_0;
	wire [2:0] w_n4336_0;
	wire [2:0] w_n4339_0;
	wire [1:0] w_n4340_0;
	wire [2:0] w_n4344_0;
	wire [2:0] w_n4346_0;
	wire [1:0] w_n4347_0;
	wire [2:0] w_n4351_0;
	wire [2:0] w_n4353_0;
	wire [1:0] w_n4354_0;
	wire [2:0] w_n4358_0;
	wire [2:0] w_n4361_0;
	wire [1:0] w_n4362_0;
	wire [2:0] w_n4366_0;
	wire [2:0] w_n4368_0;
	wire [1:0] w_n4369_0;
	wire [2:0] w_n4373_0;
	wire [2:0] w_n4376_0;
	wire [1:0] w_n4377_0;
	wire [2:0] w_n4381_0;
	wire [2:0] w_n4383_0;
	wire [1:0] w_n4384_0;
	wire [2:0] w_n4388_0;
	wire [2:0] w_n4391_0;
	wire [1:0] w_n4392_0;
	wire [2:0] w_n4396_0;
	wire [2:0] w_n4398_0;
	wire [1:0] w_n4399_0;
	wire [2:0] w_n4403_0;
	wire [2:0] w_n4406_0;
	wire [1:0] w_n4407_0;
	wire [2:0] w_n4411_0;
	wire [2:0] w_n4413_0;
	wire [1:0] w_n4414_0;
	wire [2:0] w_n4418_0;
	wire [2:0] w_n4421_0;
	wire [1:0] w_n4422_0;
	wire [2:0] w_n4426_0;
	wire [2:0] w_n4428_0;
	wire [1:0] w_n4429_0;
	wire [1:0] w_n4433_0;
	wire [2:0] w_n4435_0;
	wire [1:0] w_n4436_0;
	wire [1:0] w_n4437_0;
	wire [2:0] w_n4442_0;
	wire [1:0] w_n4447_0;
	wire [1:0] w_n4450_0;
	wire [1:0] w_n4452_0;
	wire [2:0] w_n4455_0;
	wire [2:0] w_n4457_0;
	wire [1:0] w_n4457_1;
	wire [1:0] w_n4458_0;
	wire [2:0] w_n4459_0;
	wire [1:0] w_n4460_0;
	wire [2:0] w_n4461_0;
	wire [1:0] w_n4462_0;
	wire [1:0] w_n4576_0;
	wire [1:0] w_n4580_0;
	wire [2:0] w_n4582_0;
	wire [2:0] w_n4582_1;
	wire [2:0] w_n4582_2;
	wire [2:0] w_n4582_3;
	wire [2:0] w_n4582_4;
	wire [2:0] w_n4582_5;
	wire [2:0] w_n4582_6;
	wire [2:0] w_n4582_7;
	wire [2:0] w_n4582_8;
	wire [2:0] w_n4582_9;
	wire [2:0] w_n4582_10;
	wire [2:0] w_n4582_11;
	wire [2:0] w_n4582_12;
	wire [2:0] w_n4582_13;
	wire [2:0] w_n4582_14;
	wire [2:0] w_n4582_15;
	wire [2:0] w_n4582_16;
	wire [2:0] w_n4582_17;
	wire [2:0] w_n4582_18;
	wire [2:0] w_n4582_19;
	wire [2:0] w_n4582_20;
	wire [2:0] w_n4582_21;
	wire [2:0] w_n4582_22;
	wire [2:0] w_n4582_23;
	wire [2:0] w_n4582_24;
	wire [2:0] w_n4582_25;
	wire [2:0] w_n4582_26;
	wire [2:0] w_n4582_27;
	wire [2:0] w_n4582_28;
	wire [2:0] w_n4582_29;
	wire [2:0] w_n4582_30;
	wire [2:0] w_n4582_31;
	wire [2:0] w_n4582_32;
	wire [2:0] w_n4582_33;
	wire [2:0] w_n4582_34;
	wire [2:0] w_n4582_35;
	wire [2:0] w_n4582_36;
	wire [2:0] w_n4582_37;
	wire [2:0] w_n4582_38;
	wire [2:0] w_n4582_39;
	wire [2:0] w_n4582_40;
	wire [2:0] w_n4582_41;
	wire [2:0] w_n4582_42;
	wire [2:0] w_n4582_43;
	wire [2:0] w_n4582_44;
	wire [2:0] w_n4582_45;
	wire [2:0] w_n4582_46;
	wire [2:0] w_n4582_47;
	wire [1:0] w_n4582_48;
	wire [2:0] w_n4586_0;
	wire [1:0] w_n4587_0;
	wire [1:0] w_n4589_0;
	wire [1:0] w_n4590_0;
	wire [2:0] w_n4595_0;
	wire [2:0] w_n4598_0;
	wire [1:0] w_n4599_0;
	wire [1:0] w_n4603_0;
	wire [1:0] w_n4604_0;
	wire [2:0] w_n4606_0;
	wire [1:0] w_n4607_0;
	wire [1:0] w_n4611_0;
	wire [1:0] w_n4612_0;
	wire [2:0] w_n4614_0;
	wire [1:0] w_n4615_0;
	wire [1:0] w_n4619_0;
	wire [1:0] w_n4620_0;
	wire [2:0] w_n4622_0;
	wire [1:0] w_n4623_0;
	wire [1:0] w_n4627_0;
	wire [1:0] w_n4628_0;
	wire [2:0] w_n4630_0;
	wire [1:0] w_n4631_0;
	wire [1:0] w_n4635_0;
	wire [2:0] w_n4637_0;
	wire [1:0] w_n4638_0;
	wire [1:0] w_n4642_0;
	wire [1:0] w_n4643_0;
	wire [2:0] w_n4645_0;
	wire [1:0] w_n4646_0;
	wire [1:0] w_n4650_0;
	wire [2:0] w_n4652_0;
	wire [1:0] w_n4653_0;
	wire [1:0] w_n4657_0;
	wire [1:0] w_n4658_0;
	wire [2:0] w_n4660_0;
	wire [1:0] w_n4661_0;
	wire [1:0] w_n4665_0;
	wire [2:0] w_n4667_0;
	wire [1:0] w_n4668_0;
	wire [1:0] w_n4672_0;
	wire [2:0] w_n4674_0;
	wire [1:0] w_n4675_0;
	wire [1:0] w_n4679_0;
	wire [1:0] w_n4680_0;
	wire [2:0] w_n4682_0;
	wire [1:0] w_n4683_0;
	wire [1:0] w_n4687_0;
	wire [1:0] w_n4688_0;
	wire [2:0] w_n4690_0;
	wire [1:0] w_n4691_0;
	wire [1:0] w_n4695_0;
	wire [2:0] w_n4697_0;
	wire [1:0] w_n4698_0;
	wire [1:0] w_n4702_0;
	wire [1:0] w_n4703_0;
	wire [2:0] w_n4705_0;
	wire [1:0] w_n4706_0;
	wire [1:0] w_n4710_0;
	wire [2:0] w_n4712_0;
	wire [1:0] w_n4713_0;
	wire [1:0] w_n4717_0;
	wire [1:0] w_n4718_0;
	wire [2:0] w_n4720_0;
	wire [1:0] w_n4721_0;
	wire [1:0] w_n4725_0;
	wire [2:0] w_n4727_0;
	wire [1:0] w_n4728_0;
	wire [1:0] w_n4732_0;
	wire [1:0] w_n4733_0;
	wire [2:0] w_n4735_0;
	wire [1:0] w_n4736_0;
	wire [1:0] w_n4740_0;
	wire [2:0] w_n4742_0;
	wire [1:0] w_n4743_0;
	wire [1:0] w_n4747_0;
	wire [1:0] w_n4748_0;
	wire [2:0] w_n4750_0;
	wire [1:0] w_n4751_0;
	wire [1:0] w_n4755_0;
	wire [2:0] w_n4757_0;
	wire [1:0] w_n4758_0;
	wire [2:0] w_n4762_0;
	wire [1:0] w_n4765_0;
	wire [2:0] w_n4766_0;
	wire [1:0] w_n4766_1;
	wire [2:0] w_n4767_0;
	wire [1:0] w_n4771_0;
	wire [1:0] w_n4772_0;
	wire [1:0] w_n4804_0;
	wire [1:0] w_n4823_0;
	wire [1:0] w_n4830_0;
	wire [1:0] w_n4837_0;
	wire [1:0] w_n4841_0;
	wire [1:0] w_n4851_0;
	wire [1:0] w_n4858_0;
	wire [1:0] w_n4865_0;
	wire [1:0] w_n4872_0;
	wire [1:0] w_n4879_0;
	wire [1:0] w_n4884_0;
	wire [1:0] w_n4885_0;
	wire [1:0] w_n4887_0;
	wire [1:0] w_n4889_0;
	wire [1:0] w_n4890_0;
	wire [1:0] w_n4892_0;
	wire [1:0] w_n4895_0;
	wire [1:0] w_n4901_0;
	wire [2:0] w_n4902_0;
	wire [2:0] w_n4902_1;
	wire [2:0] w_n4902_2;
	wire [2:0] w_n4902_3;
	wire [2:0] w_n4902_4;
	wire [2:0] w_n4902_5;
	wire [2:0] w_n4902_6;
	wire [2:0] w_n4902_7;
	wire [2:0] w_n4902_8;
	wire [2:0] w_n4902_9;
	wire [2:0] w_n4902_10;
	wire [2:0] w_n4902_11;
	wire [2:0] w_n4902_12;
	wire [2:0] w_n4902_13;
	wire [2:0] w_n4902_14;
	wire [2:0] w_n4902_15;
	wire [2:0] w_n4902_16;
	wire [2:0] w_n4902_17;
	wire [2:0] w_n4902_18;
	wire [2:0] w_n4902_19;
	wire [2:0] w_n4902_20;
	wire [2:0] w_n4902_21;
	wire [2:0] w_n4902_22;
	wire [2:0] w_n4902_23;
	wire [2:0] w_n4902_24;
	wire [2:0] w_n4902_25;
	wire [2:0] w_n4902_26;
	wire [2:0] w_n4902_27;
	wire [2:0] w_n4902_28;
	wire [2:0] w_n4902_29;
	wire [2:0] w_n4902_30;
	wire [2:0] w_n4902_31;
	wire [2:0] w_n4902_32;
	wire [2:0] w_n4902_33;
	wire [2:0] w_n4902_34;
	wire [2:0] w_n4902_35;
	wire [2:0] w_n4902_36;
	wire [2:0] w_n4902_37;
	wire [2:0] w_n4902_38;
	wire [2:0] w_n4902_39;
	wire [2:0] w_n4902_40;
	wire [2:0] w_n4902_41;
	wire [2:0] w_n4902_42;
	wire [2:0] w_n4902_43;
	wire [2:0] w_n4902_44;
	wire [2:0] w_n4902_45;
	wire [2:0] w_n4902_46;
	wire [2:0] w_n4902_47;
	wire [2:0] w_n4902_48;
	wire [2:0] w_n4902_49;
	wire [2:0] w_n4902_50;
	wire [2:0] w_n4902_51;
	wire [2:0] w_n4902_52;
	wire [2:0] w_n4902_53;
	wire [2:0] w_n4902_54;
	wire [2:0] w_n4902_55;
	wire [2:0] w_n4902_56;
	wire [1:0] w_n4902_57;
	wire [1:0] w_n4905_0;
	wire [2:0] w_n4906_0;
	wire [2:0] w_n4908_0;
	wire [2:0] w_n4908_1;
	wire [1:0] w_n4909_0;
	wire [2:0] w_n4910_0;
	wire [1:0] w_n4911_0;
	wire [2:0] w_n4913_0;
	wire [1:0] w_n4914_0;
	wire [2:0] w_n4921_0;
	wire [1:0] w_n4922_0;
	wire [1:0] w_n4925_0;
	wire [2:0] w_n4930_0;
	wire [2:0] w_n4932_0;
	wire [1:0] w_n4933_0;
	wire [2:0] w_n4937_0;
	wire [2:0] w_n4940_0;
	wire [1:0] w_n4941_0;
	wire [2:0] w_n4945_0;
	wire [2:0] w_n4948_0;
	wire [1:0] w_n4949_0;
	wire [1:0] w_n4953_0;
	wire [2:0] w_n4955_0;
	wire [1:0] w_n4956_0;
	wire [2:0] w_n4960_0;
	wire [2:0] w_n4962_0;
	wire [1:0] w_n4963_0;
	wire [2:0] w_n4967_0;
	wire [2:0] w_n4969_0;
	wire [1:0] w_n4970_0;
	wire [2:0] w_n4974_0;
	wire [2:0] w_n4976_0;
	wire [1:0] w_n4977_0;
	wire [2:0] w_n4981_0;
	wire [2:0] w_n4984_0;
	wire [1:0] w_n4985_0;
	wire [2:0] w_n4989_0;
	wire [2:0] w_n4991_0;
	wire [1:0] w_n4992_0;
	wire [2:0] w_n4996_0;
	wire [2:0] w_n4999_0;
	wire [1:0] w_n5000_0;
	wire [2:0] w_n5004_0;
	wire [2:0] w_n5006_0;
	wire [1:0] w_n5007_0;
	wire [2:0] w_n5011_0;
	wire [2:0] w_n5014_0;
	wire [1:0] w_n5015_0;
	wire [2:0] w_n5019_0;
	wire [2:0] w_n5022_0;
	wire [1:0] w_n5023_0;
	wire [2:0] w_n5027_0;
	wire [2:0] w_n5029_0;
	wire [1:0] w_n5030_0;
	wire [2:0] w_n5034_0;
	wire [2:0] w_n5036_0;
	wire [1:0] w_n5037_0;
	wire [2:0] w_n5041_0;
	wire [2:0] w_n5044_0;
	wire [1:0] w_n5045_0;
	wire [2:0] w_n5049_0;
	wire [2:0] w_n5051_0;
	wire [1:0] w_n5052_0;
	wire [2:0] w_n5056_0;
	wire [2:0] w_n5059_0;
	wire [1:0] w_n5060_0;
	wire [2:0] w_n5064_0;
	wire [2:0] w_n5066_0;
	wire [1:0] w_n5067_0;
	wire [1:0] w_n5071_0;
	wire [1:0] w_n5072_0;
	wire [2:0] w_n5074_0;
	wire [1:0] w_n5075_0;
	wire [2:0] w_n5079_0;
	wire [2:0] w_n5081_0;
	wire [1:0] w_n5082_0;
	wire [2:0] w_n5086_0;
	wire [2:0] w_n5089_0;
	wire [1:0] w_n5090_0;
	wire [2:0] w_n5094_0;
	wire [2:0] w_n5096_0;
	wire [1:0] w_n5097_0;
	wire [1:0] w_n5101_0;
	wire [1:0] w_n5102_0;
	wire [2:0] w_n5104_0;
	wire [2:0] w_n5105_0;
	wire [1:0] w_n5107_0;
	wire [1:0] w_n5108_0;
	wire [1:0] w_n5115_0;
	wire [1:0] w_n5116_0;
	wire [1:0] w_n5118_0;
	wire [2:0] w_n5121_0;
	wire [1:0] w_n5121_1;
	wire [1:0] w_n5122_0;
	wire [2:0] w_n5123_0;
	wire [1:0] w_n5124_0;
	wire [2:0] w_n5126_0;
	wire [1:0] w_n5127_0;
	wire [2:0] w_n5132_0;
	wire [1:0] w_n5132_1;
	wire [1:0] w_n5165_0;
	wire [1:0] w_n5179_0;
	wire [1:0] w_n5253_0;
	wire [1:0] w_n5256_0;
	wire [1:0] w_n5257_0;
	wire [2:0] w_n5259_0;
	wire [2:0] w_n5259_1;
	wire [2:0] w_n5259_2;
	wire [2:0] w_n5259_3;
	wire [2:0] w_n5259_4;
	wire [2:0] w_n5259_5;
	wire [2:0] w_n5259_6;
	wire [2:0] w_n5259_7;
	wire [2:0] w_n5259_8;
	wire [2:0] w_n5259_9;
	wire [2:0] w_n5259_10;
	wire [2:0] w_n5259_11;
	wire [2:0] w_n5259_12;
	wire [2:0] w_n5259_13;
	wire [2:0] w_n5259_14;
	wire [2:0] w_n5259_15;
	wire [2:0] w_n5259_16;
	wire [2:0] w_n5259_17;
	wire [2:0] w_n5259_18;
	wire [2:0] w_n5259_19;
	wire [2:0] w_n5259_20;
	wire [2:0] w_n5259_21;
	wire [2:0] w_n5259_22;
	wire [2:0] w_n5259_23;
	wire [2:0] w_n5259_24;
	wire [2:0] w_n5259_25;
	wire [2:0] w_n5259_26;
	wire [2:0] w_n5259_27;
	wire [2:0] w_n5259_28;
	wire [2:0] w_n5259_29;
	wire [2:0] w_n5259_30;
	wire [2:0] w_n5259_31;
	wire [2:0] w_n5259_32;
	wire [2:0] w_n5259_33;
	wire [2:0] w_n5259_34;
	wire [2:0] w_n5259_35;
	wire [2:0] w_n5259_36;
	wire [2:0] w_n5259_37;
	wire [2:0] w_n5259_38;
	wire [2:0] w_n5259_39;
	wire [2:0] w_n5259_40;
	wire [2:0] w_n5259_41;
	wire [2:0] w_n5259_42;
	wire [2:0] w_n5259_43;
	wire [2:0] w_n5259_44;
	wire [1:0] w_n5259_45;
	wire [2:0] w_n5263_0;
	wire [1:0] w_n5264_0;
	wire [1:0] w_n5266_0;
	wire [1:0] w_n5271_0;
	wire [1:0] w_n5272_0;
	wire [2:0] w_n5274_0;
	wire [1:0] w_n5275_0;
	wire [1:0] w_n5279_0;
	wire [2:0] w_n5281_0;
	wire [1:0] w_n5282_0;
	wire [1:0] w_n5286_0;
	wire [1:0] w_n5287_0;
	wire [2:0] w_n5289_0;
	wire [1:0] w_n5290_0;
	wire [1:0] w_n5294_0;
	wire [2:0] w_n5296_0;
	wire [1:0] w_n5297_0;
	wire [1:0] w_n5301_0;
	wire [2:0] w_n5303_0;
	wire [1:0] w_n5304_0;
	wire [1:0] w_n5308_0;
	wire [2:0] w_n5310_0;
	wire [1:0] w_n5311_0;
	wire [1:0] w_n5315_0;
	wire [1:0] w_n5316_0;
	wire [2:0] w_n5318_0;
	wire [1:0] w_n5319_0;
	wire [1:0] w_n5323_0;
	wire [1:0] w_n5324_0;
	wire [2:0] w_n5326_0;
	wire [1:0] w_n5327_0;
	wire [1:0] w_n5331_0;
	wire [1:0] w_n5332_0;
	wire [2:0] w_n5334_0;
	wire [1:0] w_n5335_0;
	wire [1:0] w_n5339_0;
	wire [2:0] w_n5341_0;
	wire [1:0] w_n5342_0;
	wire [1:0] w_n5346_0;
	wire [1:0] w_n5347_0;
	wire [2:0] w_n5349_0;
	wire [1:0] w_n5350_0;
	wire [1:0] w_n5354_0;
	wire [2:0] w_n5356_0;
	wire [1:0] w_n5357_0;
	wire [1:0] w_n5361_0;
	wire [1:0] w_n5362_0;
	wire [2:0] w_n5364_0;
	wire [1:0] w_n5365_0;
	wire [1:0] w_n5369_0;
	wire [2:0] w_n5371_0;
	wire [1:0] w_n5372_0;
	wire [1:0] w_n5376_0;
	wire [2:0] w_n5378_0;
	wire [1:0] w_n5379_0;
	wire [1:0] w_n5383_0;
	wire [1:0] w_n5384_0;
	wire [2:0] w_n5386_0;
	wire [1:0] w_n5387_0;
	wire [1:0] w_n5391_0;
	wire [1:0] w_n5392_0;
	wire [2:0] w_n5394_0;
	wire [1:0] w_n5395_0;
	wire [1:0] w_n5399_0;
	wire [2:0] w_n5401_0;
	wire [1:0] w_n5402_0;
	wire [1:0] w_n5406_0;
	wire [1:0] w_n5407_0;
	wire [2:0] w_n5409_0;
	wire [1:0] w_n5410_0;
	wire [1:0] w_n5414_0;
	wire [2:0] w_n5416_0;
	wire [1:0] w_n5417_0;
	wire [1:0] w_n5421_0;
	wire [1:0] w_n5422_0;
	wire [2:0] w_n5424_0;
	wire [1:0] w_n5425_0;
	wire [1:0] w_n5429_0;
	wire [1:0] w_n5430_0;
	wire [2:0] w_n5432_0;
	wire [1:0] w_n5433_0;
	wire [1:0] w_n5437_0;
	wire [1:0] w_n5438_0;
	wire [2:0] w_n5440_0;
	wire [1:0] w_n5441_0;
	wire [1:0] w_n5445_0;
	wire [2:0] w_n5447_0;
	wire [1:0] w_n5448_0;
	wire [2:0] w_n5452_0;
	wire [2:0] w_n5455_0;
	wire [1:0] w_n5458_0;
	wire [2:0] w_n5459_0;
	wire [1:0] w_n5460_0;
	wire [1:0] w_n5461_0;
	wire [1:0] w_n5465_0;
	wire [1:0] w_n5466_0;
	wire [1:0] w_n5467_0;
	wire [1:0] w_n5500_0;
	wire [1:0] w_n5507_0;
	wire [1:0] w_n5514_0;
	wire [1:0] w_n5518_0;
	wire [1:0] w_n5522_0;
	wire [1:0] w_n5535_0;
	wire [1:0] w_n5542_0;
	wire [1:0] w_n5549_0;
	wire [1:0] w_n5553_0;
	wire [1:0] w_n5563_0;
	wire [1:0] w_n5570_0;
	wire [1:0] w_n5583_0;
	wire [1:0] w_n5588_0;
	wire [1:0] w_n5592_0;
	wire [1:0] w_n5593_0;
	wire [1:0] w_n5605_0;
	wire [2:0] w_n5606_0;
	wire [2:0] w_n5606_1;
	wire [2:0] w_n5606_2;
	wire [2:0] w_n5606_3;
	wire [2:0] w_n5606_4;
	wire [2:0] w_n5606_5;
	wire [2:0] w_n5606_6;
	wire [2:0] w_n5606_7;
	wire [2:0] w_n5606_8;
	wire [2:0] w_n5606_9;
	wire [2:0] w_n5606_10;
	wire [2:0] w_n5606_11;
	wire [2:0] w_n5606_12;
	wire [2:0] w_n5606_13;
	wire [2:0] w_n5606_14;
	wire [2:0] w_n5606_15;
	wire [2:0] w_n5606_16;
	wire [2:0] w_n5606_17;
	wire [2:0] w_n5606_18;
	wire [2:0] w_n5606_19;
	wire [2:0] w_n5606_20;
	wire [2:0] w_n5606_21;
	wire [2:0] w_n5606_22;
	wire [2:0] w_n5606_23;
	wire [2:0] w_n5606_24;
	wire [2:0] w_n5606_25;
	wire [2:0] w_n5606_26;
	wire [2:0] w_n5606_27;
	wire [2:0] w_n5606_28;
	wire [2:0] w_n5606_29;
	wire [2:0] w_n5606_30;
	wire [2:0] w_n5606_31;
	wire [2:0] w_n5606_32;
	wire [2:0] w_n5606_33;
	wire [2:0] w_n5606_34;
	wire [2:0] w_n5606_35;
	wire [2:0] w_n5606_36;
	wire [2:0] w_n5606_37;
	wire [2:0] w_n5606_38;
	wire [2:0] w_n5606_39;
	wire [2:0] w_n5606_40;
	wire [2:0] w_n5606_41;
	wire [2:0] w_n5606_42;
	wire [2:0] w_n5606_43;
	wire [2:0] w_n5606_44;
	wire [2:0] w_n5606_45;
	wire [2:0] w_n5606_46;
	wire [2:0] w_n5606_47;
	wire [2:0] w_n5606_48;
	wire [2:0] w_n5606_49;
	wire [2:0] w_n5606_50;
	wire [2:0] w_n5606_51;
	wire [2:0] w_n5606_52;
	wire [2:0] w_n5606_53;
	wire [2:0] w_n5606_54;
	wire [2:0] w_n5606_55;
	wire [1:0] w_n5609_0;
	wire [2:0] w_n5610_0;
	wire [2:0] w_n5612_0;
	wire [2:0] w_n5612_1;
	wire [1:0] w_n5613_0;
	wire [2:0] w_n5614_0;
	wire [1:0] w_n5615_0;
	wire [2:0] w_n5617_0;
	wire [1:0] w_n5618_0;
	wire [2:0] w_n5625_0;
	wire [1:0] w_n5626_0;
	wire [1:0] w_n5629_0;
	wire [2:0] w_n5634_0;
	wire [2:0] w_n5636_0;
	wire [1:0] w_n5637_0;
	wire [2:0] w_n5641_0;
	wire [2:0] w_n5644_0;
	wire [1:0] w_n5645_0;
	wire [2:0] w_n5649_0;
	wire [2:0] w_n5651_0;
	wire [1:0] w_n5652_0;
	wire [2:0] w_n5656_0;
	wire [2:0] w_n5659_0;
	wire [1:0] w_n5660_0;
	wire [2:0] w_n5664_0;
	wire [2:0] w_n5666_0;
	wire [1:0] w_n5667_0;
	wire [2:0] w_n5671_0;
	wire [2:0] w_n5674_0;
	wire [1:0] w_n5675_0;
	wire [2:0] w_n5679_0;
	wire [2:0] w_n5682_0;
	wire [1:0] w_n5683_0;
	wire [2:0] w_n5687_0;
	wire [2:0] w_n5690_0;
	wire [1:0] w_n5691_0;
	wire [2:0] w_n5695_0;
	wire [2:0] w_n5697_0;
	wire [1:0] w_n5698_0;
	wire [2:0] w_n5702_0;
	wire [2:0] w_n5704_0;
	wire [1:0] w_n5705_0;
	wire [2:0] w_n5709_0;
	wire [2:0] w_n5711_0;
	wire [1:0] w_n5712_0;
	wire [2:0] w_n5716_0;
	wire [2:0] w_n5719_0;
	wire [1:0] w_n5720_0;
	wire [2:0] w_n5724_0;
	wire [2:0] w_n5726_0;
	wire [1:0] w_n5727_0;
	wire [2:0] w_n5731_0;
	wire [2:0] w_n5734_0;
	wire [1:0] w_n5735_0;
	wire [2:0] w_n5739_0;
	wire [2:0] w_n5741_0;
	wire [1:0] w_n5742_0;
	wire [2:0] w_n5746_0;
	wire [2:0] w_n5749_0;
	wire [1:0] w_n5750_0;
	wire [2:0] w_n5754_0;
	wire [2:0] w_n5757_0;
	wire [1:0] w_n5758_0;
	wire [2:0] w_n5762_0;
	wire [2:0] w_n5764_0;
	wire [1:0] w_n5765_0;
	wire [2:0] w_n5769_0;
	wire [2:0] w_n5771_0;
	wire [1:0] w_n5772_0;
	wire [2:0] w_n5776_0;
	wire [2:0] w_n5779_0;
	wire [1:0] w_n5780_0;
	wire [2:0] w_n5784_0;
	wire [2:0] w_n5786_0;
	wire [1:0] w_n5787_0;
	wire [2:0] w_n5791_0;
	wire [2:0] w_n5794_0;
	wire [1:0] w_n5795_0;
	wire [2:0] w_n5799_0;
	wire [2:0] w_n5801_0;
	wire [1:0] w_n5802_0;
	wire [2:0] w_n5806_0;
	wire [2:0] w_n5808_0;
	wire [1:0] w_n5809_0;
	wire [2:0] w_n5813_0;
	wire [2:0] w_n5815_0;
	wire [1:0] w_n5816_0;
	wire [2:0] w_n5820_0;
	wire [2:0] w_n5823_0;
	wire [1:0] w_n5823_1;
	wire [1:0] w_n5824_0;
	wire [1:0] w_n5827_0;
	wire [1:0] w_n5829_0;
	wire [1:0] w_n5834_0;
	wire [1:0] w_n5835_0;
	wire [2:0] w_n5842_0;
	wire [2:0] w_n5843_0;
	wire [1:0] w_n5843_1;
	wire [1:0] w_n5844_0;
	wire [2:0] w_n5845_0;
	wire [1:0] w_n5846_0;
	wire [2:0] w_n5848_0;
	wire [1:0] w_n5849_0;
	wire [1:0] w_n5854_0;
	wire [1:0] w_n5888_0;
	wire [1:0] w_n5986_0;
	wire [1:0] w_n5987_0;
	wire [2:0] w_n5989_0;
	wire [2:0] w_n5989_1;
	wire [2:0] w_n5989_2;
	wire [2:0] w_n5989_3;
	wire [2:0] w_n5989_4;
	wire [2:0] w_n5989_5;
	wire [2:0] w_n5989_6;
	wire [2:0] w_n5989_7;
	wire [2:0] w_n5989_8;
	wire [2:0] w_n5989_9;
	wire [2:0] w_n5989_10;
	wire [2:0] w_n5989_11;
	wire [2:0] w_n5989_12;
	wire [2:0] w_n5989_13;
	wire [2:0] w_n5989_14;
	wire [2:0] w_n5989_15;
	wire [2:0] w_n5989_16;
	wire [2:0] w_n5989_17;
	wire [2:0] w_n5989_18;
	wire [2:0] w_n5989_19;
	wire [2:0] w_n5989_20;
	wire [2:0] w_n5989_21;
	wire [2:0] w_n5989_22;
	wire [2:0] w_n5989_23;
	wire [2:0] w_n5989_24;
	wire [2:0] w_n5989_25;
	wire [2:0] w_n5989_26;
	wire [2:0] w_n5989_27;
	wire [2:0] w_n5989_28;
	wire [2:0] w_n5989_29;
	wire [2:0] w_n5989_30;
	wire [2:0] w_n5989_31;
	wire [2:0] w_n5989_32;
	wire [2:0] w_n5989_33;
	wire [2:0] w_n5989_34;
	wire [2:0] w_n5989_35;
	wire [2:0] w_n5989_36;
	wire [2:0] w_n5989_37;
	wire [2:0] w_n5989_38;
	wire [2:0] w_n5989_39;
	wire [2:0] w_n5989_40;
	wire [2:0] w_n5989_41;
	wire [1:0] w_n5989_42;
	wire [2:0] w_n5993_0;
	wire [1:0] w_n5994_0;
	wire [1:0] w_n5996_0;
	wire [1:0] w_n6001_0;
	wire [1:0] w_n6002_0;
	wire [2:0] w_n6004_0;
	wire [1:0] w_n6005_0;
	wire [1:0] w_n6009_0;
	wire [2:0] w_n6011_0;
	wire [1:0] w_n6012_0;
	wire [1:0] w_n6016_0;
	wire [1:0] w_n6017_0;
	wire [2:0] w_n6019_0;
	wire [1:0] w_n6020_0;
	wire [1:0] w_n6024_0;
	wire [2:0] w_n6026_0;
	wire [1:0] w_n6027_0;
	wire [1:0] w_n6031_0;
	wire [1:0] w_n6032_0;
	wire [2:0] w_n6034_0;
	wire [1:0] w_n6035_0;
	wire [1:0] w_n6039_0;
	wire [2:0] w_n6041_0;
	wire [1:0] w_n6042_0;
	wire [1:0] w_n6046_0;
	wire [1:0] w_n6047_0;
	wire [2:0] w_n6049_0;
	wire [1:0] w_n6050_0;
	wire [1:0] w_n6054_0;
	wire [2:0] w_n6056_0;
	wire [1:0] w_n6057_0;
	wire [1:0] w_n6061_0;
	wire [2:0] w_n6063_0;
	wire [1:0] w_n6064_0;
	wire [1:0] w_n6068_0;
	wire [2:0] w_n6070_0;
	wire [1:0] w_n6071_0;
	wire [1:0] w_n6075_0;
	wire [1:0] w_n6076_0;
	wire [2:0] w_n6078_0;
	wire [1:0] w_n6079_0;
	wire [1:0] w_n6083_0;
	wire [1:0] w_n6084_0;
	wire [2:0] w_n6086_0;
	wire [1:0] w_n6087_0;
	wire [1:0] w_n6091_0;
	wire [1:0] w_n6092_0;
	wire [2:0] w_n6094_0;
	wire [1:0] w_n6095_0;
	wire [1:0] w_n6099_0;
	wire [2:0] w_n6101_0;
	wire [1:0] w_n6102_0;
	wire [1:0] w_n6106_0;
	wire [1:0] w_n6107_0;
	wire [2:0] w_n6109_0;
	wire [1:0] w_n6110_0;
	wire [1:0] w_n6114_0;
	wire [2:0] w_n6116_0;
	wire [1:0] w_n6117_0;
	wire [1:0] w_n6121_0;
	wire [1:0] w_n6122_0;
	wire [2:0] w_n6124_0;
	wire [1:0] w_n6125_0;
	wire [1:0] w_n6129_0;
	wire [2:0] w_n6131_0;
	wire [1:0] w_n6132_0;
	wire [1:0] w_n6136_0;
	wire [2:0] w_n6138_0;
	wire [1:0] w_n6139_0;
	wire [1:0] w_n6143_0;
	wire [1:0] w_n6144_0;
	wire [2:0] w_n6146_0;
	wire [1:0] w_n6147_0;
	wire [1:0] w_n6151_0;
	wire [1:0] w_n6152_0;
	wire [2:0] w_n6154_0;
	wire [1:0] w_n6155_0;
	wire [1:0] w_n6159_0;
	wire [2:0] w_n6161_0;
	wire [1:0] w_n6162_0;
	wire [2:0] w_n6166_0;
	wire [2:0] w_n6169_0;
	wire [1:0] w_n6170_0;
	wire [1:0] w_n6174_0;
	wire [2:0] w_n6176_0;
	wire [1:0] w_n6177_0;
	wire [1:0] w_n6181_0;
	wire [1:0] w_n6182_0;
	wire [2:0] w_n6184_0;
	wire [1:0] w_n6185_0;
	wire [1:0] w_n6189_0;
	wire [1:0] w_n6190_0;
	wire [2:0] w_n6192_0;
	wire [1:0] w_n6193_0;
	wire [2:0] w_n6197_0;
	wire [1:0] w_n6200_0;
	wire [2:0] w_n6201_0;
	wire [1:0] w_n6201_1;
	wire [2:0] w_n6202_0;
	wire [1:0] w_n6204_0;
	wire [1:0] w_n6239_0;
	wire [1:0] w_n6246_0;
	wire [1:0] w_n6253_0;
	wire [1:0] w_n6260_0;
	wire [1:0] w_n6267_0;
	wire [1:0] w_n6271_0;
	wire [1:0] w_n6275_0;
	wire [1:0] w_n6288_0;
	wire [1:0] w_n6295_0;
	wire [1:0] w_n6302_0;
	wire [1:0] w_n6306_0;
	wire [1:0] w_n6316_0;
	wire [1:0] w_n6323_0;
	wire [1:0] w_n6334_0;
	wire [1:0] w_n6335_0;
	wire [1:0] w_n6336_0;
	wire [1:0] w_n6338_0;
	wire [1:0] w_n6340_0;
	wire [1:0] w_n6343_0;
	wire [1:0] w_n6344_0;
	wire [1:0] w_n6345_0;
	wire [1:0] w_n6348_0;
	wire [1:0] w_n6349_0;
	wire [1:0] w_n6355_0;
	wire [2:0] w_n6357_0;
	wire [2:0] w_n6357_1;
	wire [2:0] w_n6357_2;
	wire [2:0] w_n6357_3;
	wire [2:0] w_n6357_4;
	wire [2:0] w_n6357_5;
	wire [2:0] w_n6357_6;
	wire [2:0] w_n6357_7;
	wire [2:0] w_n6357_8;
	wire [2:0] w_n6357_9;
	wire [2:0] w_n6357_10;
	wire [2:0] w_n6357_11;
	wire [2:0] w_n6357_12;
	wire [2:0] w_n6357_13;
	wire [2:0] w_n6357_14;
	wire [2:0] w_n6357_15;
	wire [2:0] w_n6357_16;
	wire [2:0] w_n6357_17;
	wire [2:0] w_n6357_18;
	wire [2:0] w_n6357_19;
	wire [2:0] w_n6357_20;
	wire [2:0] w_n6357_21;
	wire [2:0] w_n6357_22;
	wire [2:0] w_n6357_23;
	wire [2:0] w_n6357_24;
	wire [2:0] w_n6357_25;
	wire [2:0] w_n6357_26;
	wire [2:0] w_n6357_27;
	wire [2:0] w_n6357_28;
	wire [2:0] w_n6357_29;
	wire [2:0] w_n6357_30;
	wire [2:0] w_n6357_31;
	wire [2:0] w_n6357_32;
	wire [2:0] w_n6357_33;
	wire [2:0] w_n6357_34;
	wire [2:0] w_n6357_35;
	wire [2:0] w_n6357_36;
	wire [2:0] w_n6357_37;
	wire [2:0] w_n6357_38;
	wire [2:0] w_n6357_39;
	wire [2:0] w_n6357_40;
	wire [2:0] w_n6357_41;
	wire [2:0] w_n6357_42;
	wire [2:0] w_n6357_43;
	wire [2:0] w_n6357_44;
	wire [2:0] w_n6357_45;
	wire [2:0] w_n6357_46;
	wire [2:0] w_n6357_47;
	wire [2:0] w_n6357_48;
	wire [2:0] w_n6357_49;
	wire [2:0] w_n6357_50;
	wire [2:0] w_n6357_51;
	wire [2:0] w_n6357_52;
	wire [2:0] w_n6357_53;
	wire [2:0] w_n6357_54;
	wire [1:0] w_n6360_0;
	wire [2:0] w_n6361_0;
	wire [2:0] w_n6362_0;
	wire [2:0] w_n6362_1;
	wire [1:0] w_n6363_0;
	wire [2:0] w_n6364_0;
	wire [1:0] w_n6365_0;
	wire [2:0] w_n6368_0;
	wire [1:0] w_n6369_0;
	wire [2:0] w_n6376_0;
	wire [1:0] w_n6377_0;
	wire [1:0] w_n6380_0;
	wire [1:0] w_n6385_0;
	wire [2:0] w_n6387_0;
	wire [1:0] w_n6388_0;
	wire [2:0] w_n6392_0;
	wire [2:0] w_n6395_0;
	wire [1:0] w_n6396_0;
	wire [2:0] w_n6400_0;
	wire [2:0] w_n6402_0;
	wire [1:0] w_n6403_0;
	wire [2:0] w_n6407_0;
	wire [2:0] w_n6410_0;
	wire [1:0] w_n6411_0;
	wire [2:0] w_n6415_0;
	wire [2:0] w_n6417_0;
	wire [1:0] w_n6418_0;
	wire [2:0] w_n6422_0;
	wire [2:0] w_n6425_0;
	wire [1:0] w_n6426_0;
	wire [2:0] w_n6430_0;
	wire [2:0] w_n6432_0;
	wire [1:0] w_n6433_0;
	wire [2:0] w_n6437_0;
	wire [2:0] w_n6440_0;
	wire [1:0] w_n6441_0;
	wire [2:0] w_n6445_0;
	wire [2:0] w_n6447_0;
	wire [1:0] w_n6448_0;
	wire [2:0] w_n6452_0;
	wire [2:0] w_n6455_0;
	wire [1:0] w_n6456_0;
	wire [2:0] w_n6460_0;
	wire [2:0] w_n6463_0;
	wire [1:0] w_n6464_0;
	wire [2:0] w_n6468_0;
	wire [2:0] w_n6471_0;
	wire [1:0] w_n6472_0;
	wire [2:0] w_n6476_0;
	wire [2:0] w_n6478_0;
	wire [1:0] w_n6479_0;
	wire [2:0] w_n6483_0;
	wire [2:0] w_n6485_0;
	wire [1:0] w_n6486_0;
	wire [2:0] w_n6490_0;
	wire [2:0] w_n6492_0;
	wire [1:0] w_n6493_0;
	wire [2:0] w_n6497_0;
	wire [2:0] w_n6500_0;
	wire [1:0] w_n6501_0;
	wire [2:0] w_n6505_0;
	wire [2:0] w_n6507_0;
	wire [1:0] w_n6508_0;
	wire [2:0] w_n6512_0;
	wire [2:0] w_n6515_0;
	wire [1:0] w_n6516_0;
	wire [2:0] w_n6520_0;
	wire [2:0] w_n6522_0;
	wire [1:0] w_n6523_0;
	wire [2:0] w_n6527_0;
	wire [2:0] w_n6530_0;
	wire [1:0] w_n6531_0;
	wire [2:0] w_n6535_0;
	wire [2:0] w_n6538_0;
	wire [1:0] w_n6539_0;
	wire [2:0] w_n6543_0;
	wire [2:0] w_n6545_0;
	wire [1:0] w_n6546_0;
	wire [2:0] w_n6550_0;
	wire [2:0] w_n6552_0;
	wire [1:0] w_n6553_0;
	wire [1:0] w_n6557_0;
	wire [1:0] w_n6558_0;
	wire [2:0] w_n6560_0;
	wire [1:0] w_n6561_0;
	wire [2:0] w_n6565_0;
	wire [2:0] w_n6568_0;
	wire [1:0] w_n6569_0;
	wire [2:0] w_n6573_0;
	wire [2:0] w_n6576_0;
	wire [1:0] w_n6577_0;
	wire [2:0] w_n6581_0;
	wire [2:0] w_n6583_0;
	wire [1:0] w_n6584_0;
	wire [2:0] w_n6588_0;
	wire [2:0] w_n6590_0;
	wire [1:0] w_n6591_0;
	wire [2:0] w_n6596_0;
	wire [1:0] w_n6601_0;
	wire [1:0] w_n6604_0;
	wire [2:0] w_n6606_0;
	wire [2:0] w_n6606_1;
	wire [1:0] w_n6607_0;
	wire [2:0] w_n6608_0;
	wire [1:0] w_n6609_0;
	wire [2:0] w_n6611_0;
	wire [1:0] w_n6612_0;
	wire [1:0] w_n6652_0;
	wire [1:0] w_n6656_0;
	wire [1:0] w_n6753_0;
	wire [1:0] w_n6756_0;
	wire [2:0] w_n6758_0;
	wire [2:0] w_n6758_1;
	wire [2:0] w_n6758_2;
	wire [2:0] w_n6758_3;
	wire [2:0] w_n6758_4;
	wire [2:0] w_n6758_5;
	wire [2:0] w_n6758_6;
	wire [2:0] w_n6758_7;
	wire [2:0] w_n6758_8;
	wire [2:0] w_n6758_9;
	wire [2:0] w_n6758_10;
	wire [2:0] w_n6758_11;
	wire [2:0] w_n6758_12;
	wire [2:0] w_n6758_13;
	wire [2:0] w_n6758_14;
	wire [2:0] w_n6758_15;
	wire [2:0] w_n6758_16;
	wire [2:0] w_n6758_17;
	wire [2:0] w_n6758_18;
	wire [2:0] w_n6758_19;
	wire [2:0] w_n6758_20;
	wire [2:0] w_n6758_21;
	wire [2:0] w_n6758_22;
	wire [2:0] w_n6758_23;
	wire [2:0] w_n6758_24;
	wire [2:0] w_n6758_25;
	wire [2:0] w_n6758_26;
	wire [2:0] w_n6758_27;
	wire [2:0] w_n6758_28;
	wire [2:0] w_n6758_29;
	wire [2:0] w_n6758_30;
	wire [2:0] w_n6758_31;
	wire [2:0] w_n6758_32;
	wire [2:0] w_n6758_33;
	wire [2:0] w_n6758_34;
	wire [2:0] w_n6758_35;
	wire [2:0] w_n6758_36;
	wire [2:0] w_n6758_37;
	wire [2:0] w_n6758_38;
	wire [2:0] w_n6758_39;
	wire [2:0] w_n6758_40;
	wire [2:0] w_n6762_0;
	wire [1:0] w_n6763_0;
	wire [1:0] w_n6765_0;
	wire [1:0] w_n6766_0;
	wire [1:0] w_n6771_0;
	wire [1:0] w_n6772_0;
	wire [2:0] w_n6774_0;
	wire [1:0] w_n6775_0;
	wire [1:0] w_n6779_0;
	wire [2:0] w_n6781_0;
	wire [1:0] w_n6782_0;
	wire [1:0] w_n6786_0;
	wire [2:0] w_n6788_0;
	wire [1:0] w_n6789_0;
	wire [1:0] w_n6793_0;
	wire [2:0] w_n6795_0;
	wire [1:0] w_n6796_0;
	wire [1:0] w_n6800_0;
	wire [1:0] w_n6801_0;
	wire [2:0] w_n6803_0;
	wire [1:0] w_n6804_0;
	wire [1:0] w_n6808_0;
	wire [2:0] w_n6810_0;
	wire [1:0] w_n6811_0;
	wire [1:0] w_n6815_0;
	wire [1:0] w_n6816_0;
	wire [2:0] w_n6818_0;
	wire [1:0] w_n6819_0;
	wire [1:0] w_n6823_0;
	wire [2:0] w_n6825_0;
	wire [1:0] w_n6826_0;
	wire [1:0] w_n6830_0;
	wire [1:0] w_n6831_0;
	wire [2:0] w_n6833_0;
	wire [1:0] w_n6834_0;
	wire [1:0] w_n6838_0;
	wire [2:0] w_n6840_0;
	wire [1:0] w_n6841_0;
	wire [1:0] w_n6845_0;
	wire [1:0] w_n6846_0;
	wire [2:0] w_n6848_0;
	wire [1:0] w_n6849_0;
	wire [1:0] w_n6853_0;
	wire [2:0] w_n6855_0;
	wire [1:0] w_n6856_0;
	wire [1:0] w_n6860_0;
	wire [2:0] w_n6862_0;
	wire [1:0] w_n6863_0;
	wire [1:0] w_n6867_0;
	wire [2:0] w_n6869_0;
	wire [1:0] w_n6870_0;
	wire [1:0] w_n6874_0;
	wire [1:0] w_n6875_0;
	wire [2:0] w_n6877_0;
	wire [1:0] w_n6878_0;
	wire [1:0] w_n6882_0;
	wire [1:0] w_n6883_0;
	wire [2:0] w_n6885_0;
	wire [1:0] w_n6886_0;
	wire [1:0] w_n6890_0;
	wire [1:0] w_n6891_0;
	wire [2:0] w_n6893_0;
	wire [1:0] w_n6894_0;
	wire [1:0] w_n6898_0;
	wire [2:0] w_n6900_0;
	wire [1:0] w_n6901_0;
	wire [1:0] w_n6905_0;
	wire [1:0] w_n6906_0;
	wire [2:0] w_n6908_0;
	wire [1:0] w_n6909_0;
	wire [1:0] w_n6913_0;
	wire [2:0] w_n6915_0;
	wire [1:0] w_n6916_0;
	wire [1:0] w_n6920_0;
	wire [1:0] w_n6921_0;
	wire [2:0] w_n6923_0;
	wire [1:0] w_n6924_0;
	wire [1:0] w_n6928_0;
	wire [2:0] w_n6930_0;
	wire [1:0] w_n6931_0;
	wire [1:0] w_n6935_0;
	wire [2:0] w_n6937_0;
	wire [1:0] w_n6938_0;
	wire [1:0] w_n6942_0;
	wire [1:0] w_n6943_0;
	wire [2:0] w_n6945_0;
	wire [1:0] w_n6946_0;
	wire [1:0] w_n6950_0;
	wire [1:0] w_n6951_0;
	wire [2:0] w_n6953_0;
	wire [1:0] w_n6954_0;
	wire [1:0] w_n6958_0;
	wire [1:0] w_n6959_0;
	wire [2:0] w_n6961_0;
	wire [1:0] w_n6962_0;
	wire [1:0] w_n6966_0;
	wire [2:0] w_n6968_0;
	wire [1:0] w_n6969_0;
	wire [1:0] w_n6973_0;
	wire [2:0] w_n6975_0;
	wire [1:0] w_n6976_0;
	wire [1:0] w_n6980_0;
	wire [1:0] w_n6981_0;
	wire [1:0] w_n6983_0;
	wire [2:0] w_n6986_0;
	wire [1:0] w_n6987_0;
	wire [2:0] w_n6988_0;
	wire [1:0] w_n6988_1;
	wire [2:0] w_n6989_0;
	wire [1:0] w_n6993_0;
	wire [1:0] w_n6994_0;
	wire [1:0] w_n7031_0;
	wire [1:0] w_n7038_0;
	wire [1:0] w_n7042_0;
	wire [1:0] w_n7046_0;
	wire [1:0] w_n7053_0;
	wire [1:0] w_n7060_0;
	wire [1:0] w_n7067_0;
	wire [1:0] w_n7074_0;
	wire [1:0] w_n7078_0;
	wire [1:0] w_n7082_0;
	wire [1:0] w_n7095_0;
	wire [1:0] w_n7102_0;
	wire [1:0] w_n7109_0;
	wire [1:0] w_n7113_0;
	wire [1:0] w_n7126_0;
	wire [1:0] w_n7130_0;
	wire [1:0] w_n7135_0;
	wire [1:0] w_n7136_0;
	wire [1:0] w_n7138_0;
	wire [1:0] w_n7140_0;
	wire [1:0] w_n7141_0;
	wire [1:0] w_n7143_0;
	wire [1:0] w_n7145_0;
	wire [1:0] w_n7146_0;
	wire [1:0] w_n7153_0;
	wire [2:0] w_n7154_0;
	wire [2:0] w_n7154_1;
	wire [2:0] w_n7154_2;
	wire [2:0] w_n7154_3;
	wire [2:0] w_n7154_4;
	wire [2:0] w_n7154_5;
	wire [2:0] w_n7154_6;
	wire [2:0] w_n7154_7;
	wire [2:0] w_n7154_8;
	wire [2:0] w_n7154_9;
	wire [2:0] w_n7154_10;
	wire [2:0] w_n7154_11;
	wire [2:0] w_n7154_12;
	wire [2:0] w_n7154_13;
	wire [2:0] w_n7154_14;
	wire [2:0] w_n7154_15;
	wire [2:0] w_n7154_16;
	wire [2:0] w_n7154_17;
	wire [2:0] w_n7154_18;
	wire [2:0] w_n7154_19;
	wire [2:0] w_n7154_20;
	wire [2:0] w_n7154_21;
	wire [2:0] w_n7154_22;
	wire [2:0] w_n7154_23;
	wire [2:0] w_n7154_24;
	wire [2:0] w_n7154_25;
	wire [2:0] w_n7154_26;
	wire [2:0] w_n7154_27;
	wire [2:0] w_n7154_28;
	wire [2:0] w_n7154_29;
	wire [2:0] w_n7154_30;
	wire [2:0] w_n7154_31;
	wire [2:0] w_n7154_32;
	wire [2:0] w_n7154_33;
	wire [2:0] w_n7154_34;
	wire [2:0] w_n7154_35;
	wire [2:0] w_n7154_36;
	wire [2:0] w_n7154_37;
	wire [2:0] w_n7154_38;
	wire [2:0] w_n7154_39;
	wire [2:0] w_n7154_40;
	wire [2:0] w_n7154_41;
	wire [2:0] w_n7154_42;
	wire [2:0] w_n7154_43;
	wire [2:0] w_n7154_44;
	wire [2:0] w_n7154_45;
	wire [2:0] w_n7154_46;
	wire [2:0] w_n7154_47;
	wire [2:0] w_n7154_48;
	wire [2:0] w_n7154_49;
	wire [2:0] w_n7154_50;
	wire [2:0] w_n7154_51;
	wire [2:0] w_n7154_52;
	wire [2:0] w_n7154_53;
	wire [2:0] w_n7156_0;
	wire [2:0] w_n7156_1;
	wire [1:0] w_n7157_0;
	wire [2:0] w_n7158_0;
	wire [1:0] w_n7159_0;
	wire [2:0] w_n7161_0;
	wire [1:0] w_n7162_0;
	wire [2:0] w_n7169_0;
	wire [1:0] w_n7170_0;
	wire [1:0] w_n7173_0;
	wire [2:0] w_n7178_0;
	wire [2:0] w_n7180_0;
	wire [1:0] w_n7181_0;
	wire [2:0] w_n7185_0;
	wire [2:0] w_n7188_0;
	wire [1:0] w_n7189_0;
	wire [2:0] w_n7193_0;
	wire [2:0] w_n7195_0;
	wire [1:0] w_n7196_0;
	wire [2:0] w_n7200_0;
	wire [2:0] w_n7203_0;
	wire [1:0] w_n7204_0;
	wire [2:0] w_n7208_0;
	wire [2:0] w_n7211_0;
	wire [1:0] w_n7212_0;
	wire [2:0] w_n7216_0;
	wire [2:0] w_n7219_0;
	wire [1:0] w_n7220_0;
	wire [2:0] w_n7224_0;
	wire [2:0] w_n7226_0;
	wire [1:0] w_n7227_0;
	wire [2:0] w_n7231_0;
	wire [2:0] w_n7234_0;
	wire [1:0] w_n7235_0;
	wire [2:0] w_n7239_0;
	wire [2:0] w_n7241_0;
	wire [1:0] w_n7242_0;
	wire [2:0] w_n7246_0;
	wire [2:0] w_n7249_0;
	wire [1:0] w_n7250_0;
	wire [2:0] w_n7254_0;
	wire [2:0] w_n7256_0;
	wire [1:0] w_n7257_0;
	wire [2:0] w_n7261_0;
	wire [2:0] w_n7264_0;
	wire [1:0] w_n7265_0;
	wire [2:0] w_n7269_0;
	wire [2:0] w_n7271_0;
	wire [1:0] w_n7272_0;
	wire [2:0] w_n7276_0;
	wire [2:0] w_n7279_0;
	wire [1:0] w_n7280_0;
	wire [2:0] w_n7284_0;
	wire [2:0] w_n7287_0;
	wire [1:0] w_n7288_0;
	wire [2:0] w_n7292_0;
	wire [2:0] w_n7295_0;
	wire [1:0] w_n7296_0;
	wire [2:0] w_n7300_0;
	wire [2:0] w_n7302_0;
	wire [1:0] w_n7303_0;
	wire [2:0] w_n7307_0;
	wire [2:0] w_n7309_0;
	wire [1:0] w_n7310_0;
	wire [2:0] w_n7314_0;
	wire [2:0] w_n7316_0;
	wire [1:0] w_n7317_0;
	wire [2:0] w_n7321_0;
	wire [2:0] w_n7324_0;
	wire [1:0] w_n7325_0;
	wire [2:0] w_n7329_0;
	wire [2:0] w_n7331_0;
	wire [1:0] w_n7332_0;
	wire [2:0] w_n7336_0;
	wire [2:0] w_n7339_0;
	wire [1:0] w_n7340_0;
	wire [2:0] w_n7344_0;
	wire [2:0] w_n7346_0;
	wire [1:0] w_n7347_0;
	wire [2:0] w_n7351_0;
	wire [2:0] w_n7354_0;
	wire [1:0] w_n7355_0;
	wire [2:0] w_n7359_0;
	wire [2:0] w_n7362_0;
	wire [1:0] w_n7363_0;
	wire [2:0] w_n7367_0;
	wire [2:0] w_n7369_0;
	wire [1:0] w_n7370_0;
	wire [2:0] w_n7374_0;
	wire [2:0] w_n7376_0;
	wire [1:0] w_n7377_0;
	wire [2:0] w_n7381_0;
	wire [2:0] w_n7383_0;
	wire [1:0] w_n7384_0;
	wire [2:0] w_n7388_0;
	wire [2:0] w_n7391_0;
	wire [1:0] w_n7392_0;
	wire [2:0] w_n7396_0;
	wire [2:0] w_n7399_0;
	wire [2:0] w_n7402_0;
	wire [1:0] w_n7402_1;
	wire [1:0] w_n7403_0;
	wire [1:0] w_n7406_0;
	wire [2:0] w_n7408_0;
	wire [1:0] w_n7408_1;
	wire [1:0] w_n7413_0;
	wire [1:0] w_n7415_0;
	wire [2:0] w_n7419_0;
	wire [2:0] w_n7421_0;
	wire [2:0] w_n7421_1;
	wire [1:0] w_n7422_0;
	wire [2:0] w_n7423_0;
	wire [1:0] w_n7424_0;
	wire [2:0] w_n7425_0;
	wire [1:0] w_n7426_0;
	wire [1:0] w_n7465_0;
	wire [1:0] w_n7576_0;
	wire [2:0] w_n7581_0;
	wire [2:0] w_n7581_1;
	wire [2:0] w_n7581_2;
	wire [2:0] w_n7581_3;
	wire [2:0] w_n7581_4;
	wire [2:0] w_n7581_5;
	wire [2:0] w_n7581_6;
	wire [2:0] w_n7581_7;
	wire [2:0] w_n7581_8;
	wire [2:0] w_n7581_9;
	wire [2:0] w_n7581_10;
	wire [2:0] w_n7581_11;
	wire [2:0] w_n7581_12;
	wire [2:0] w_n7581_13;
	wire [2:0] w_n7581_14;
	wire [2:0] w_n7581_15;
	wire [2:0] w_n7581_16;
	wire [2:0] w_n7581_17;
	wire [2:0] w_n7581_18;
	wire [2:0] w_n7581_19;
	wire [2:0] w_n7581_20;
	wire [2:0] w_n7581_21;
	wire [2:0] w_n7581_22;
	wire [2:0] w_n7581_23;
	wire [2:0] w_n7581_24;
	wire [2:0] w_n7581_25;
	wire [2:0] w_n7581_26;
	wire [2:0] w_n7581_27;
	wire [2:0] w_n7581_28;
	wire [2:0] w_n7581_29;
	wire [2:0] w_n7581_30;
	wire [2:0] w_n7581_31;
	wire [2:0] w_n7581_32;
	wire [2:0] w_n7581_33;
	wire [2:0] w_n7581_34;
	wire [2:0] w_n7581_35;
	wire [2:0] w_n7581_36;
	wire [2:0] w_n7581_37;
	wire [1:0] w_n7581_38;
	wire [1:0] w_n7582_0;
	wire [1:0] w_n7583_0;
	wire [2:0] w_n7585_0;
	wire [1:0] w_n7586_0;
	wire [1:0] w_n7592_0;
	wire [1:0] w_n7593_0;
	wire [2:0] w_n7595_0;
	wire [1:0] w_n7596_0;
	wire [1:0] w_n7599_0;
	wire [2:0] w_n7602_0;
	wire [1:0] w_n7603_0;
	wire [1:0] w_n7607_0;
	wire [1:0] w_n7608_0;
	wire [2:0] w_n7610_0;
	wire [1:0] w_n7611_0;
	wire [1:0] w_n7615_0;
	wire [2:0] w_n7617_0;
	wire [1:0] w_n7618_0;
	wire [1:0] w_n7622_0;
	wire [1:0] w_n7623_0;
	wire [2:0] w_n7625_0;
	wire [1:0] w_n7626_0;
	wire [1:0] w_n7630_0;
	wire [2:0] w_n7632_0;
	wire [1:0] w_n7633_0;
	wire [1:0] w_n7637_0;
	wire [2:0] w_n7639_0;
	wire [1:0] w_n7640_0;
	wire [1:0] w_n7644_0;
	wire [2:0] w_n7646_0;
	wire [1:0] w_n7647_0;
	wire [1:0] w_n7651_0;
	wire [1:0] w_n7652_0;
	wire [2:0] w_n7654_0;
	wire [1:0] w_n7655_0;
	wire [1:0] w_n7659_0;
	wire [2:0] w_n7661_0;
	wire [1:0] w_n7662_0;
	wire [1:0] w_n7666_0;
	wire [1:0] w_n7667_0;
	wire [2:0] w_n7669_0;
	wire [1:0] w_n7670_0;
	wire [1:0] w_n7674_0;
	wire [2:0] w_n7676_0;
	wire [1:0] w_n7677_0;
	wire [1:0] w_n7681_0;
	wire [1:0] w_n7682_0;
	wire [2:0] w_n7684_0;
	wire [1:0] w_n7685_0;
	wire [1:0] w_n7689_0;
	wire [2:0] w_n7691_0;
	wire [1:0] w_n7692_0;
	wire [1:0] w_n7696_0;
	wire [1:0] w_n7697_0;
	wire [2:0] w_n7699_0;
	wire [1:0] w_n7700_0;
	wire [1:0] w_n7704_0;
	wire [2:0] w_n7706_0;
	wire [1:0] w_n7707_0;
	wire [1:0] w_n7711_0;
	wire [2:0] w_n7713_0;
	wire [1:0] w_n7714_0;
	wire [1:0] w_n7718_0;
	wire [2:0] w_n7720_0;
	wire [1:0] w_n7721_0;
	wire [1:0] w_n7725_0;
	wire [1:0] w_n7726_0;
	wire [2:0] w_n7728_0;
	wire [1:0] w_n7729_0;
	wire [1:0] w_n7733_0;
	wire [1:0] w_n7734_0;
	wire [2:0] w_n7736_0;
	wire [1:0] w_n7737_0;
	wire [1:0] w_n7741_0;
	wire [1:0] w_n7742_0;
	wire [2:0] w_n7744_0;
	wire [1:0] w_n7745_0;
	wire [1:0] w_n7749_0;
	wire [2:0] w_n7751_0;
	wire [1:0] w_n7752_0;
	wire [1:0] w_n7756_0;
	wire [1:0] w_n7757_0;
	wire [2:0] w_n7759_0;
	wire [1:0] w_n7760_0;
	wire [1:0] w_n7764_0;
	wire [2:0] w_n7766_0;
	wire [1:0] w_n7767_0;
	wire [1:0] w_n7771_0;
	wire [1:0] w_n7772_0;
	wire [2:0] w_n7774_0;
	wire [1:0] w_n7775_0;
	wire [1:0] w_n7779_0;
	wire [2:0] w_n7781_0;
	wire [1:0] w_n7782_0;
	wire [1:0] w_n7786_0;
	wire [2:0] w_n7788_0;
	wire [1:0] w_n7789_0;
	wire [1:0] w_n7793_0;
	wire [1:0] w_n7794_0;
	wire [2:0] w_n7796_0;
	wire [1:0] w_n7797_0;
	wire [1:0] w_n7801_0;
	wire [1:0] w_n7802_0;
	wire [2:0] w_n7804_0;
	wire [1:0] w_n7805_0;
	wire [1:0] w_n7809_0;
	wire [1:0] w_n7810_0;
	wire [2:0] w_n7812_0;
	wire [1:0] w_n7813_0;
	wire [2:0] w_n7817_0;
	wire [1:0] w_n7819_0;
	wire [2:0] w_n7820_0;
	wire [1:0] w_n7820_1;
	wire [2:0] w_n7821_0;
	wire [1:0] w_n7826_0;
	wire [1:0] w_n7827_0;
	wire [1:0] w_n7828_0;
	wire [1:0] w_n7859_0;
	wire [1:0] w_n7882_0;
	wire [1:0] w_n7889_0;
	wire [1:0] w_n7893_0;
	wire [1:0] w_n7897_0;
	wire [1:0] w_n7904_0;
	wire [1:0] w_n7911_0;
	wire [1:0] w_n7918_0;
	wire [1:0] w_n7925_0;
	wire [1:0] w_n7929_0;
	wire [1:0] w_n7933_0;
	wire [1:0] w_n7946_0;
	wire [1:0] w_n7953_0;
	wire [1:0] w_n7960_0;
	wire [1:0] w_n7964_0;
	wire [1:0] w_n7979_0;
	wire [1:0] w_n7980_0;
	wire [1:0] w_n7982_0;
	wire [1:0] w_n7984_0;
	wire [1:0] w_n7985_0;
	wire [1:0] w_n7987_0;
	wire [1:0] w_n7989_0;
	wire [1:0] w_n7990_0;
	wire [2:0] w_n7991_0;
	wire [2:0] w_n7991_1;
	wire [1:0] w_n7992_0;
	wire [2:0] w_n7993_0;
	wire [1:0] w_n7994_0;
	wire [1:0] w_n8002_0;
	wire [2:0] w_n8003_0;
	wire [2:0] w_n8003_1;
	wire [2:0] w_n8003_2;
	wire [2:0] w_n8003_3;
	wire [2:0] w_n8003_4;
	wire [2:0] w_n8003_5;
	wire [2:0] w_n8003_6;
	wire [2:0] w_n8003_7;
	wire [2:0] w_n8003_8;
	wire [2:0] w_n8003_9;
	wire [2:0] w_n8003_10;
	wire [2:0] w_n8003_11;
	wire [2:0] w_n8003_12;
	wire [2:0] w_n8003_13;
	wire [2:0] w_n8003_14;
	wire [2:0] w_n8003_15;
	wire [2:0] w_n8003_16;
	wire [2:0] w_n8003_17;
	wire [2:0] w_n8003_18;
	wire [2:0] w_n8003_19;
	wire [2:0] w_n8003_20;
	wire [2:0] w_n8003_21;
	wire [2:0] w_n8003_22;
	wire [2:0] w_n8003_23;
	wire [2:0] w_n8003_24;
	wire [2:0] w_n8003_25;
	wire [2:0] w_n8003_26;
	wire [2:0] w_n8003_27;
	wire [2:0] w_n8003_28;
	wire [2:0] w_n8003_29;
	wire [2:0] w_n8003_30;
	wire [2:0] w_n8003_31;
	wire [2:0] w_n8003_32;
	wire [2:0] w_n8003_33;
	wire [2:0] w_n8003_34;
	wire [2:0] w_n8003_35;
	wire [2:0] w_n8003_36;
	wire [2:0] w_n8003_37;
	wire [2:0] w_n8003_38;
	wire [2:0] w_n8003_39;
	wire [2:0] w_n8003_40;
	wire [2:0] w_n8003_41;
	wire [2:0] w_n8003_42;
	wire [2:0] w_n8003_43;
	wire [2:0] w_n8003_44;
	wire [2:0] w_n8003_45;
	wire [2:0] w_n8003_46;
	wire [2:0] w_n8003_47;
	wire [2:0] w_n8003_48;
	wire [2:0] w_n8003_49;
	wire [2:0] w_n8003_50;
	wire [2:0] w_n8003_51;
	wire [1:0] w_n8003_52;
	wire [2:0] w_n8005_0;
	wire [1:0] w_n8006_0;
	wire [2:0] w_n8013_0;
	wire [1:0] w_n8014_0;
	wire [1:0] w_n8017_0;
	wire [2:0] w_n8022_0;
	wire [2:0] w_n8024_0;
	wire [1:0] w_n8025_0;
	wire [2:0] w_n8029_0;
	wire [2:0] w_n8031_0;
	wire [1:0] w_n8032_0;
	wire [2:0] w_n8036_0;
	wire [2:0] w_n8038_0;
	wire [1:0] w_n8039_0;
	wire [2:0] w_n8042_0;
	wire [2:0] w_n8046_0;
	wire [1:0] w_n8047_0;
	wire [2:0] w_n8051_0;
	wire [2:0] w_n8053_0;
	wire [1:0] w_n8054_0;
	wire [2:0] w_n8058_0;
	wire [2:0] w_n8061_0;
	wire [1:0] w_n8062_0;
	wire [2:0] w_n8066_0;
	wire [2:0] w_n8068_0;
	wire [1:0] w_n8069_0;
	wire [2:0] w_n8073_0;
	wire [2:0] w_n8076_0;
	wire [1:0] w_n8077_0;
	wire [2:0] w_n8081_0;
	wire [2:0] w_n8084_0;
	wire [1:0] w_n8085_0;
	wire [2:0] w_n8089_0;
	wire [2:0] w_n8092_0;
	wire [1:0] w_n8093_0;
	wire [2:0] w_n8097_0;
	wire [2:0] w_n8099_0;
	wire [1:0] w_n8100_0;
	wire [2:0] w_n8104_0;
	wire [2:0] w_n8107_0;
	wire [1:0] w_n8108_0;
	wire [2:0] w_n8112_0;
	wire [2:0] w_n8114_0;
	wire [1:0] w_n8115_0;
	wire [2:0] w_n8119_0;
	wire [2:0] w_n8122_0;
	wire [1:0] w_n8123_0;
	wire [2:0] w_n8127_0;
	wire [2:0] w_n8129_0;
	wire [1:0] w_n8130_0;
	wire [2:0] w_n8134_0;
	wire [2:0] w_n8137_0;
	wire [1:0] w_n8138_0;
	wire [2:0] w_n8142_0;
	wire [2:0] w_n8144_0;
	wire [1:0] w_n8145_0;
	wire [2:0] w_n8149_0;
	wire [2:0] w_n8152_0;
	wire [1:0] w_n8153_0;
	wire [2:0] w_n8157_0;
	wire [2:0] w_n8160_0;
	wire [1:0] w_n8161_0;
	wire [2:0] w_n8165_0;
	wire [2:0] w_n8168_0;
	wire [1:0] w_n8169_0;
	wire [2:0] w_n8173_0;
	wire [2:0] w_n8175_0;
	wire [1:0] w_n8176_0;
	wire [2:0] w_n8180_0;
	wire [2:0] w_n8182_0;
	wire [1:0] w_n8183_0;
	wire [2:0] w_n8187_0;
	wire [2:0] w_n8189_0;
	wire [1:0] w_n8190_0;
	wire [2:0] w_n8194_0;
	wire [2:0] w_n8197_0;
	wire [1:0] w_n8198_0;
	wire [2:0] w_n8202_0;
	wire [2:0] w_n8204_0;
	wire [1:0] w_n8205_0;
	wire [2:0] w_n8209_0;
	wire [2:0] w_n8212_0;
	wire [1:0] w_n8213_0;
	wire [2:0] w_n8217_0;
	wire [2:0] w_n8219_0;
	wire [1:0] w_n8220_0;
	wire [2:0] w_n8224_0;
	wire [2:0] w_n8227_0;
	wire [1:0] w_n8228_0;
	wire [2:0] w_n8232_0;
	wire [2:0] w_n8235_0;
	wire [1:0] w_n8236_0;
	wire [2:0] w_n8240_0;
	wire [2:0] w_n8242_0;
	wire [1:0] w_n8243_0;
	wire [2:0] w_n8247_0;
	wire [2:0] w_n8249_0;
	wire [1:0] w_n8250_0;
	wire [1:0] w_n8254_0;
	wire [2:0] w_n8256_0;
	wire [2:0] w_n8259_0;
	wire [1:0] w_n8260_0;
	wire [1:0] w_n8263_0;
	wire [2:0] w_n8265_0;
	wire [1:0] w_n8265_1;
	wire [1:0] w_n8270_0;
	wire [1:0] w_n8272_0;
	wire [1:0] w_n8274_0;
	wire [2:0] w_n8277_0;
	wire [2:0] w_n8279_0;
	wire [1:0] w_n8279_1;
	wire [1:0] w_n8280_0;
	wire [2:0] w_n8281_0;
	wire [1:0] w_n8282_0;
	wire [2:0] w_n8283_0;
	wire [1:0] w_n8284_0;
	wire [1:0] w_n8328_0;
	wire [1:0] w_n8444_0;
	wire [2:0] w_n8449_0;
	wire [2:0] w_n8449_1;
	wire [2:0] w_n8449_2;
	wire [2:0] w_n8449_3;
	wire [2:0] w_n8449_4;
	wire [2:0] w_n8449_5;
	wire [2:0] w_n8449_6;
	wire [2:0] w_n8449_7;
	wire [2:0] w_n8449_8;
	wire [2:0] w_n8449_9;
	wire [2:0] w_n8449_10;
	wire [2:0] w_n8449_11;
	wire [2:0] w_n8449_12;
	wire [2:0] w_n8449_13;
	wire [2:0] w_n8449_14;
	wire [2:0] w_n8449_15;
	wire [2:0] w_n8449_16;
	wire [2:0] w_n8449_17;
	wire [2:0] w_n8449_18;
	wire [2:0] w_n8449_19;
	wire [2:0] w_n8449_20;
	wire [2:0] w_n8449_21;
	wire [2:0] w_n8449_22;
	wire [2:0] w_n8449_23;
	wire [2:0] w_n8449_24;
	wire [2:0] w_n8449_25;
	wire [2:0] w_n8449_26;
	wire [2:0] w_n8449_27;
	wire [2:0] w_n8449_28;
	wire [2:0] w_n8449_29;
	wire [2:0] w_n8449_30;
	wire [2:0] w_n8449_31;
	wire [2:0] w_n8449_32;
	wire [2:0] w_n8449_33;
	wire [2:0] w_n8449_34;
	wire [1:0] w_n8449_35;
	wire [1:0] w_n8450_0;
	wire [2:0] w_n8453_0;
	wire [1:0] w_n8454_0;
	wire [1:0] w_n8460_0;
	wire [1:0] w_n8461_0;
	wire [2:0] w_n8463_0;
	wire [1:0] w_n8464_0;
	wire [2:0] w_n8468_0;
	wire [2:0] w_n8470_0;
	wire [1:0] w_n8471_0;
	wire [1:0] w_n8475_0;
	wire [1:0] w_n8476_0;
	wire [2:0] w_n8478_0;
	wire [1:0] w_n8479_0;
	wire [1:0] w_n8483_0;
	wire [1:0] w_n8484_0;
	wire [2:0] w_n8486_0;
	wire [1:0] w_n8487_0;
	wire [1:0] w_n8491_0;
	wire [1:0] w_n8492_0;
	wire [2:0] w_n8494_0;
	wire [1:0] w_n8495_0;
	wire [1:0] w_n8498_0;
	wire [2:0] w_n8501_0;
	wire [1:0] w_n8502_0;
	wire [1:0] w_n8506_0;
	wire [1:0] w_n8507_0;
	wire [2:0] w_n8509_0;
	wire [1:0] w_n8510_0;
	wire [1:0] w_n8514_0;
	wire [2:0] w_n8516_0;
	wire [1:0] w_n8517_0;
	wire [1:0] w_n8521_0;
	wire [1:0] w_n8522_0;
	wire [2:0] w_n8524_0;
	wire [1:0] w_n8525_0;
	wire [1:0] w_n8529_0;
	wire [2:0] w_n8531_0;
	wire [1:0] w_n8532_0;
	wire [1:0] w_n8536_0;
	wire [2:0] w_n8538_0;
	wire [1:0] w_n8539_0;
	wire [1:0] w_n8543_0;
	wire [2:0] w_n8545_0;
	wire [1:0] w_n8546_0;
	wire [1:0] w_n8550_0;
	wire [1:0] w_n8551_0;
	wire [2:0] w_n8553_0;
	wire [1:0] w_n8554_0;
	wire [1:0] w_n8558_0;
	wire [2:0] w_n8560_0;
	wire [1:0] w_n8561_0;
	wire [1:0] w_n8565_0;
	wire [1:0] w_n8566_0;
	wire [2:0] w_n8568_0;
	wire [1:0] w_n8569_0;
	wire [1:0] w_n8573_0;
	wire [2:0] w_n8575_0;
	wire [1:0] w_n8576_0;
	wire [1:0] w_n8580_0;
	wire [1:0] w_n8581_0;
	wire [2:0] w_n8583_0;
	wire [1:0] w_n8584_0;
	wire [1:0] w_n8588_0;
	wire [2:0] w_n8590_0;
	wire [1:0] w_n8591_0;
	wire [1:0] w_n8595_0;
	wire [1:0] w_n8596_0;
	wire [2:0] w_n8598_0;
	wire [1:0] w_n8599_0;
	wire [1:0] w_n8603_0;
	wire [2:0] w_n8605_0;
	wire [1:0] w_n8606_0;
	wire [1:0] w_n8610_0;
	wire [2:0] w_n8612_0;
	wire [1:0] w_n8613_0;
	wire [1:0] w_n8617_0;
	wire [2:0] w_n8619_0;
	wire [1:0] w_n8620_0;
	wire [1:0] w_n8624_0;
	wire [1:0] w_n8625_0;
	wire [2:0] w_n8627_0;
	wire [1:0] w_n8628_0;
	wire [1:0] w_n8632_0;
	wire [1:0] w_n8633_0;
	wire [2:0] w_n8635_0;
	wire [1:0] w_n8636_0;
	wire [1:0] w_n8640_0;
	wire [1:0] w_n8641_0;
	wire [2:0] w_n8643_0;
	wire [1:0] w_n8644_0;
	wire [1:0] w_n8648_0;
	wire [2:0] w_n8650_0;
	wire [1:0] w_n8651_0;
	wire [1:0] w_n8655_0;
	wire [1:0] w_n8656_0;
	wire [2:0] w_n8658_0;
	wire [1:0] w_n8659_0;
	wire [1:0] w_n8663_0;
	wire [2:0] w_n8665_0;
	wire [1:0] w_n8666_0;
	wire [1:0] w_n8670_0;
	wire [1:0] w_n8671_0;
	wire [2:0] w_n8673_0;
	wire [1:0] w_n8674_0;
	wire [1:0] w_n8678_0;
	wire [2:0] w_n8680_0;
	wire [1:0] w_n8681_0;
	wire [1:0] w_n8685_0;
	wire [2:0] w_n8687_0;
	wire [1:0] w_n8688_0;
	wire [1:0] w_n8692_0;
	wire [1:0] w_n8693_0;
	wire [2:0] w_n8695_0;
	wire [1:0] w_n8696_0;
	wire [2:0] w_n8700_0;
	wire [1:0] w_n8703_0;
	wire [2:0] w_n8704_0;
	wire [2:0] w_n8705_0;
	wire [1:0] w_n8707_0;
	wire [1:0] w_n8736_0;
	wire [1:0] w_n8750_0;
	wire [1:0] w_n8776_0;
	wire [1:0] w_n8783_0;
	wire [1:0] w_n8787_0;
	wire [1:0] w_n8791_0;
	wire [1:0] w_n8798_0;
	wire [1:0] w_n8805_0;
	wire [1:0] w_n8812_0;
	wire [1:0] w_n8819_0;
	wire [1:0] w_n8823_0;
	wire [1:0] w_n8827_0;
	wire [1:0] w_n8840_0;
	wire [1:0] w_n8847_0;
	wire [1:0] w_n8854_0;
	wire [1:0] w_n8858_0;
	wire [1:0] w_n8866_0;
	wire [1:0] w_n8867_0;
	wire [1:0] w_n8868_0;
	wire [1:0] w_n8871_0;
	wire [1:0] w_n8874_0;
	wire [1:0] w_n8876_0;
	wire [1:0] w_n8877_0;
	wire [1:0] w_n8878_0;
	wire [1:0] w_n8882_0;
	wire [1:0] w_n8888_0;
	wire [2:0] w_n8890_0;
	wire [2:0] w_n8890_1;
	wire [2:0] w_n8890_2;
	wire [2:0] w_n8890_3;
	wire [2:0] w_n8890_4;
	wire [2:0] w_n8890_5;
	wire [2:0] w_n8890_6;
	wire [2:0] w_n8890_7;
	wire [2:0] w_n8890_8;
	wire [2:0] w_n8890_9;
	wire [2:0] w_n8890_10;
	wire [2:0] w_n8890_11;
	wire [2:0] w_n8890_12;
	wire [2:0] w_n8890_13;
	wire [2:0] w_n8890_14;
	wire [2:0] w_n8890_15;
	wire [2:0] w_n8890_16;
	wire [2:0] w_n8890_17;
	wire [2:0] w_n8890_18;
	wire [2:0] w_n8890_19;
	wire [2:0] w_n8890_20;
	wire [2:0] w_n8890_21;
	wire [2:0] w_n8890_22;
	wire [2:0] w_n8890_23;
	wire [2:0] w_n8890_24;
	wire [2:0] w_n8890_25;
	wire [2:0] w_n8890_26;
	wire [2:0] w_n8890_27;
	wire [2:0] w_n8890_28;
	wire [2:0] w_n8890_29;
	wire [2:0] w_n8890_30;
	wire [2:0] w_n8890_31;
	wire [2:0] w_n8890_32;
	wire [2:0] w_n8890_33;
	wire [2:0] w_n8890_34;
	wire [2:0] w_n8890_35;
	wire [2:0] w_n8890_36;
	wire [2:0] w_n8890_37;
	wire [2:0] w_n8890_38;
	wire [2:0] w_n8890_39;
	wire [2:0] w_n8890_40;
	wire [2:0] w_n8890_41;
	wire [2:0] w_n8890_42;
	wire [2:0] w_n8890_43;
	wire [2:0] w_n8890_44;
	wire [2:0] w_n8890_45;
	wire [2:0] w_n8890_46;
	wire [2:0] w_n8890_47;
	wire [2:0] w_n8890_48;
	wire [2:0] w_n8890_49;
	wire [1:0] w_n8890_50;
	wire [1:0] w_n8893_0;
	wire [2:0] w_n8894_0;
	wire [1:0] w_n8894_1;
	wire [2:0] w_n8895_0;
	wire [2:0] w_n8895_1;
	wire [1:0] w_n8896_0;
	wire [2:0] w_n8897_0;
	wire [1:0] w_n8898_0;
	wire [2:0] w_n8901_0;
	wire [1:0] w_n8902_0;
	wire [2:0] w_n8909_0;
	wire [1:0] w_n8910_0;
	wire [1:0] w_n8913_0;
	wire [2:0] w_n8918_0;
	wire [2:0] w_n8920_0;
	wire [1:0] w_n8921_0;
	wire [2:0] w_n8925_0;
	wire [2:0] w_n8928_0;
	wire [1:0] w_n8929_0;
	wire [2:0] w_n8933_0;
	wire [2:0] w_n8935_0;
	wire [1:0] w_n8936_0;
	wire [2:0] w_n8940_0;
	wire [2:0] w_n8942_0;
	wire [1:0] w_n8943_0;
	wire [2:0] w_n8947_0;
	wire [2:0] w_n8949_0;
	wire [1:0] w_n8950_0;
	wire [2:0] w_n8954_0;
	wire [2:0] w_n8956_0;
	wire [1:0] w_n8957_0;
	wire [2:0] w_n8961_0;
	wire [2:0] w_n8963_0;
	wire [1:0] w_n8964_0;
	wire [2:0] w_n8967_0;
	wire [2:0] w_n8971_0;
	wire [1:0] w_n8972_0;
	wire [2:0] w_n8976_0;
	wire [2:0] w_n8978_0;
	wire [1:0] w_n8979_0;
	wire [2:0] w_n8983_0;
	wire [2:0] w_n8986_0;
	wire [1:0] w_n8987_0;
	wire [2:0] w_n8991_0;
	wire [2:0] w_n8993_0;
	wire [1:0] w_n8994_0;
	wire [2:0] w_n8998_0;
	wire [2:0] w_n9001_0;
	wire [1:0] w_n9002_0;
	wire [2:0] w_n9006_0;
	wire [2:0] w_n9009_0;
	wire [1:0] w_n9010_0;
	wire [1:0] w_n9014_0;
	wire [1:0] w_n9015_0;
	wire [2:0] w_n9017_0;
	wire [1:0] w_n9018_0;
	wire [2:0] w_n9022_0;
	wire [2:0] w_n9024_0;
	wire [1:0] w_n9025_0;
	wire [2:0] w_n9029_0;
	wire [2:0] w_n9032_0;
	wire [1:0] w_n9033_0;
	wire [2:0] w_n9037_0;
	wire [2:0] w_n9039_0;
	wire [1:0] w_n9040_0;
	wire [2:0] w_n9044_0;
	wire [2:0] w_n9047_0;
	wire [1:0] w_n9048_0;
	wire [2:0] w_n9052_0;
	wire [2:0] w_n9054_0;
	wire [1:0] w_n9055_0;
	wire [2:0] w_n9059_0;
	wire [2:0] w_n9062_0;
	wire [1:0] w_n9063_0;
	wire [2:0] w_n9067_0;
	wire [2:0] w_n9069_0;
	wire [1:0] w_n9070_0;
	wire [2:0] w_n9074_0;
	wire [2:0] w_n9077_0;
	wire [1:0] w_n9078_0;
	wire [2:0] w_n9082_0;
	wire [2:0] w_n9085_0;
	wire [1:0] w_n9086_0;
	wire [2:0] w_n9090_0;
	wire [2:0] w_n9093_0;
	wire [1:0] w_n9094_0;
	wire [2:0] w_n9098_0;
	wire [2:0] w_n9100_0;
	wire [1:0] w_n9101_0;
	wire [2:0] w_n9105_0;
	wire [2:0] w_n9107_0;
	wire [1:0] w_n9108_0;
	wire [2:0] w_n9112_0;
	wire [2:0] w_n9114_0;
	wire [1:0] w_n9115_0;
	wire [2:0] w_n9119_0;
	wire [2:0] w_n9122_0;
	wire [1:0] w_n9123_0;
	wire [2:0] w_n9127_0;
	wire [2:0] w_n9129_0;
	wire [1:0] w_n9130_0;
	wire [1:0] w_n9134_0;
	wire [1:0] w_n9135_0;
	wire [2:0] w_n9137_0;
	wire [1:0] w_n9138_0;
	wire [2:0] w_n9142_0;
	wire [2:0] w_n9144_0;
	wire [1:0] w_n9145_0;
	wire [2:0] w_n9149_0;
	wire [2:0] w_n9152_0;
	wire [1:0] w_n9153_0;
	wire [2:0] w_n9157_0;
	wire [2:0] w_n9160_0;
	wire [1:0] w_n9161_0;
	wire [1:0] w_n9165_0;
	wire [2:0] w_n9167_0;
	wire [1:0] w_n9167_1;
	wire [1:0] w_n9168_0;
	wire [1:0] w_n9172_0;
	wire [1:0] w_n9173_0;
	wire [1:0] w_n9177_0;
	wire [1:0] w_n9180_0;
	wire [1:0] w_n9184_0;
	wire [2:0] w_n9187_0;
	wire [2:0] w_n9188_0;
	wire [2:0] w_n9188_1;
	wire [1:0] w_n9189_0;
	wire [2:0] w_n9190_0;
	wire [1:0] w_n9191_0;
	wire [2:0] w_n9193_0;
	wire [1:0] w_n9194_0;
	wire [1:0] w_n9199_0;
	wire [1:0] w_n9240_0;
	wire [1:0] w_n9365_0;
	wire [1:0] w_n9368_0;
	wire [2:0] w_n9369_0;
	wire [2:0] w_n9369_1;
	wire [2:0] w_n9369_2;
	wire [2:0] w_n9369_3;
	wire [2:0] w_n9369_4;
	wire [2:0] w_n9369_5;
	wire [2:0] w_n9369_6;
	wire [2:0] w_n9369_7;
	wire [2:0] w_n9369_8;
	wire [2:0] w_n9369_9;
	wire [2:0] w_n9369_10;
	wire [2:0] w_n9369_11;
	wire [2:0] w_n9369_12;
	wire [2:0] w_n9369_13;
	wire [2:0] w_n9369_14;
	wire [2:0] w_n9369_15;
	wire [2:0] w_n9369_16;
	wire [2:0] w_n9369_17;
	wire [2:0] w_n9369_18;
	wire [2:0] w_n9369_19;
	wire [2:0] w_n9369_20;
	wire [2:0] w_n9369_21;
	wire [2:0] w_n9369_22;
	wire [2:0] w_n9369_23;
	wire [2:0] w_n9369_24;
	wire [2:0] w_n9369_25;
	wire [2:0] w_n9369_26;
	wire [2:0] w_n9369_27;
	wire [2:0] w_n9369_28;
	wire [2:0] w_n9369_29;
	wire [2:0] w_n9369_30;
	wire [2:0] w_n9369_31;
	wire [2:0] w_n9369_32;
	wire [1:0] w_n9369_33;
	wire [2:0] w_n9373_0;
	wire [1:0] w_n9374_0;
	wire [1:0] w_n9376_0;
	wire [1:0] w_n9381_0;
	wire [1:0] w_n9382_0;
	wire [2:0] w_n9384_0;
	wire [1:0] w_n9385_0;
	wire [2:0] w_n9389_0;
	wire [2:0] w_n9391_0;
	wire [1:0] w_n9392_0;
	wire [1:0] w_n9396_0;
	wire [1:0] w_n9397_0;
	wire [2:0] w_n9399_0;
	wire [1:0] w_n9400_0;
	wire [1:0] w_n9404_0;
	wire [2:0] w_n9406_0;
	wire [1:0] w_n9407_0;
	wire [1:0] w_n9411_0;
	wire [1:0] w_n9412_0;
	wire [2:0] w_n9414_0;
	wire [1:0] w_n9415_0;
	wire [1:0] w_n9419_0;
	wire [1:0] w_n9420_0;
	wire [2:0] w_n9422_0;
	wire [1:0] w_n9423_0;
	wire [1:0] w_n9427_0;
	wire [1:0] w_n9428_0;
	wire [2:0] w_n9430_0;
	wire [1:0] w_n9431_0;
	wire [1:0] w_n9435_0;
	wire [1:0] w_n9436_0;
	wire [2:0] w_n9438_0;
	wire [1:0] w_n9439_0;
	wire [1:0] w_n9443_0;
	wire [1:0] w_n9444_0;
	wire [2:0] w_n9446_0;
	wire [1:0] w_n9447_0;
	wire [1:0] w_n9450_0;
	wire [2:0] w_n9453_0;
	wire [1:0] w_n9454_0;
	wire [1:0] w_n9458_0;
	wire [1:0] w_n9459_0;
	wire [2:0] w_n9461_0;
	wire [1:0] w_n9462_0;
	wire [1:0] w_n9466_0;
	wire [2:0] w_n9468_0;
	wire [1:0] w_n9469_0;
	wire [1:0] w_n9473_0;
	wire [1:0] w_n9474_0;
	wire [2:0] w_n9476_0;
	wire [1:0] w_n9477_0;
	wire [1:0] w_n9481_0;
	wire [2:0] w_n9483_0;
	wire [1:0] w_n9484_0;
	wire [2:0] w_n9488_0;
	wire [2:0] w_n9490_0;
	wire [1:0] w_n9491_0;
	wire [1:0] w_n9495_0;
	wire [1:0] w_n9496_0;
	wire [2:0] w_n9498_0;
	wire [1:0] w_n9499_0;
	wire [1:0] w_n9503_0;
	wire [1:0] w_n9504_0;
	wire [2:0] w_n9506_0;
	wire [1:0] w_n9507_0;
	wire [1:0] w_n9511_0;
	wire [2:0] w_n9513_0;
	wire [1:0] w_n9514_0;
	wire [1:0] w_n9518_0;
	wire [1:0] w_n9519_0;
	wire [2:0] w_n9521_0;
	wire [1:0] w_n9522_0;
	wire [1:0] w_n9526_0;
	wire [2:0] w_n9528_0;
	wire [1:0] w_n9529_0;
	wire [1:0] w_n9533_0;
	wire [1:0] w_n9534_0;
	wire [2:0] w_n9536_0;
	wire [1:0] w_n9537_0;
	wire [1:0] w_n9541_0;
	wire [2:0] w_n9543_0;
	wire [1:0] w_n9544_0;
	wire [1:0] w_n9548_0;
	wire [1:0] w_n9549_0;
	wire [2:0] w_n9551_0;
	wire [1:0] w_n9552_0;
	wire [1:0] w_n9556_0;
	wire [2:0] w_n9558_0;
	wire [1:0] w_n9559_0;
	wire [1:0] w_n9563_0;
	wire [2:0] w_n9565_0;
	wire [1:0] w_n9566_0;
	wire [1:0] w_n9570_0;
	wire [2:0] w_n9572_0;
	wire [1:0] w_n9573_0;
	wire [1:0] w_n9577_0;
	wire [1:0] w_n9578_0;
	wire [2:0] w_n9580_0;
	wire [1:0] w_n9581_0;
	wire [1:0] w_n9585_0;
	wire [1:0] w_n9586_0;
	wire [2:0] w_n9588_0;
	wire [1:0] w_n9589_0;
	wire [1:0] w_n9593_0;
	wire [1:0] w_n9594_0;
	wire [2:0] w_n9596_0;
	wire [1:0] w_n9597_0;
	wire [1:0] w_n9601_0;
	wire [2:0] w_n9603_0;
	wire [1:0] w_n9604_0;
	wire [1:0] w_n9608_0;
	wire [1:0] w_n9609_0;
	wire [2:0] w_n9611_0;
	wire [1:0] w_n9612_0;
	wire [1:0] w_n9616_0;
	wire [1:0] w_n9617_0;
	wire [2:0] w_n9619_0;
	wire [1:0] w_n9620_0;
	wire [1:0] w_n9624_0;
	wire [1:0] w_n9625_0;
	wire [2:0] w_n9627_0;
	wire [1:0] w_n9628_0;
	wire [1:0] w_n9632_0;
	wire [2:0] w_n9634_0;
	wire [1:0] w_n9635_0;
	wire [2:0] w_n9639_0;
	wire [1:0] w_n9641_0;
	wire [2:0] w_n9642_0;
	wire [1:0] w_n9642_1;
	wire [2:0] w_n9643_0;
	wire [1:0] w_n9646_0;
	wire [1:0] w_n9647_0;
	wire [1:0] w_n9648_0;
	wire [1:0] w_n9649_0;
	wire [1:0] w_n9676_0;
	wire [1:0] w_n9693_0;
	wire [1:0] w_n9707_0;
	wire [1:0] w_n9732_0;
	wire [1:0] w_n9739_0;
	wire [1:0] w_n9753_0;
	wire [1:0] w_n9760_0;
	wire [1:0] w_n9767_0;
	wire [1:0] w_n9774_0;
	wire [1:0] w_n9778_0;
	wire [1:0] w_n9782_0;
	wire [1:0] w_n9795_0;
	wire [1:0] w_n9808_0;
	wire [1:0] w_n9814_0;
	wire [1:0] w_n9815_0;
	wire [1:0] w_n9816_0;
	wire [1:0] w_n9819_0;
	wire [1:0] w_n9820_0;
	wire [1:0] w_n9822_0;
	wire [1:0] w_n9824_0;
	wire [1:0] w_n9825_0;
	wire [1:0] w_n9831_0;
	wire [2:0] w_n9832_0;
	wire [2:0] w_n9832_1;
	wire [2:0] w_n9832_2;
	wire [2:0] w_n9832_3;
	wire [2:0] w_n9832_4;
	wire [2:0] w_n9832_5;
	wire [2:0] w_n9832_6;
	wire [2:0] w_n9832_7;
	wire [2:0] w_n9832_8;
	wire [2:0] w_n9832_9;
	wire [2:0] w_n9832_10;
	wire [2:0] w_n9832_11;
	wire [2:0] w_n9832_12;
	wire [2:0] w_n9832_13;
	wire [2:0] w_n9832_14;
	wire [2:0] w_n9832_15;
	wire [2:0] w_n9832_16;
	wire [2:0] w_n9832_17;
	wire [2:0] w_n9832_18;
	wire [2:0] w_n9832_19;
	wire [2:0] w_n9832_20;
	wire [2:0] w_n9832_21;
	wire [2:0] w_n9832_22;
	wire [2:0] w_n9832_23;
	wire [2:0] w_n9832_24;
	wire [2:0] w_n9832_25;
	wire [2:0] w_n9832_26;
	wire [2:0] w_n9832_27;
	wire [2:0] w_n9832_28;
	wire [2:0] w_n9832_29;
	wire [2:0] w_n9832_30;
	wire [2:0] w_n9832_31;
	wire [2:0] w_n9832_32;
	wire [2:0] w_n9832_33;
	wire [2:0] w_n9832_34;
	wire [2:0] w_n9832_35;
	wire [2:0] w_n9832_36;
	wire [2:0] w_n9832_37;
	wire [2:0] w_n9832_38;
	wire [2:0] w_n9832_39;
	wire [2:0] w_n9832_40;
	wire [2:0] w_n9832_41;
	wire [2:0] w_n9832_42;
	wire [2:0] w_n9832_43;
	wire [2:0] w_n9832_44;
	wire [2:0] w_n9832_45;
	wire [2:0] w_n9832_46;
	wire [2:0] w_n9832_47;
	wire [2:0] w_n9832_48;
	wire [1:0] w_n9832_49;
	wire [2:0] w_n9834_0;
	wire [2:0] w_n9834_1;
	wire [1:0] w_n9835_0;
	wire [2:0] w_n9836_0;
	wire [1:0] w_n9837_0;
	wire [2:0] w_n9839_0;
	wire [1:0] w_n9840_0;
	wire [2:0] w_n9847_0;
	wire [1:0] w_n9848_0;
	wire [1:0] w_n9851_0;
	wire [2:0] w_n9856_0;
	wire [2:0] w_n9858_0;
	wire [1:0] w_n9859_0;
	wire [2:0] w_n9863_0;
	wire [2:0] w_n9866_0;
	wire [1:0] w_n9867_0;
	wire [2:0] w_n9871_0;
	wire [2:0] w_n9873_0;
	wire [1:0] w_n9874_0;
	wire [2:0] w_n9878_0;
	wire [2:0] w_n9880_0;
	wire [1:0] w_n9881_0;
	wire [2:0] w_n9885_0;
	wire [2:0] w_n9887_0;
	wire [1:0] w_n9888_0;
	wire [2:0] w_n9892_0;
	wire [2:0] w_n9895_0;
	wire [1:0] w_n9896_0;
	wire [2:0] w_n9900_0;
	wire [2:0] w_n9902_0;
	wire [1:0] w_n9903_0;
	wire [2:0] w_n9907_0;
	wire [2:0] w_n9909_0;
	wire [1:0] w_n9910_0;
	wire [2:0] w_n9914_0;
	wire [2:0] w_n9916_0;
	wire [1:0] w_n9917_0;
	wire [2:0] w_n9921_0;
	wire [2:0] w_n9923_0;
	wire [1:0] w_n9924_0;
	wire [2:0] w_n9928_0;
	wire [2:0] w_n9930_0;
	wire [1:0] w_n9931_0;
	wire [2:0] w_n9934_0;
	wire [2:0] w_n9938_0;
	wire [1:0] w_n9939_0;
	wire [2:0] w_n9943_0;
	wire [2:0] w_n9945_0;
	wire [1:0] w_n9946_0;
	wire [2:0] w_n9950_0;
	wire [2:0] w_n9953_0;
	wire [1:0] w_n9954_0;
	wire [2:0] w_n9958_0;
	wire [2:0] w_n9960_0;
	wire [1:0] w_n9961_0;
	wire [2:0] w_n9965_0;
	wire [2:0] w_n9968_0;
	wire [1:0] w_n9969_0;
	wire [2:0] w_n9973_0;
	wire [2:0] w_n9975_0;
	wire [1:0] w_n9976_0;
	wire [2:0] w_n9980_0;
	wire [2:0] w_n9982_0;
	wire [1:0] w_n9983_0;
	wire [2:0] w_n9987_0;
	wire [2:0] w_n9989_0;
	wire [1:0] w_n9990_0;
	wire [2:0] w_n9994_0;
	wire [2:0] w_n9997_0;
	wire [1:0] w_n9998_0;
	wire [2:0] w_n10002_0;
	wire [2:0] w_n10004_0;
	wire [1:0] w_n10005_0;
	wire [2:0] w_n10009_0;
	wire [2:0] w_n10012_0;
	wire [1:0] w_n10013_0;
	wire [2:0] w_n10017_0;
	wire [2:0] w_n10019_0;
	wire [1:0] w_n10020_0;
	wire [2:0] w_n10024_0;
	wire [2:0] w_n10027_0;
	wire [1:0] w_n10028_0;
	wire [2:0] w_n10032_0;
	wire [2:0] w_n10034_0;
	wire [1:0] w_n10035_0;
	wire [2:0] w_n10039_0;
	wire [2:0] w_n10042_0;
	wire [1:0] w_n10043_0;
	wire [2:0] w_n10047_0;
	wire [2:0] w_n10050_0;
	wire [1:0] w_n10051_0;
	wire [2:0] w_n10055_0;
	wire [2:0] w_n10058_0;
	wire [1:0] w_n10059_0;
	wire [2:0] w_n10063_0;
	wire [2:0] w_n10065_0;
	wire [1:0] w_n10066_0;
	wire [2:0] w_n10070_0;
	wire [2:0] w_n10072_0;
	wire [1:0] w_n10073_0;
	wire [2:0] w_n10077_0;
	wire [2:0] w_n10079_0;
	wire [1:0] w_n10080_0;
	wire [2:0] w_n10084_0;
	wire [2:0] w_n10087_0;
	wire [1:0] w_n10088_0;
	wire [2:0] w_n10092_0;
	wire [2:0] w_n10094_0;
	wire [1:0] w_n10095_0;
	wire [2:0] w_n10099_0;
	wire [2:0] w_n10101_0;
	wire [1:0] w_n10102_0;
	wire [2:0] w_n10106_0;
	wire [2:0] w_n10108_0;
	wire [1:0] w_n10109_0;
	wire [1:0] w_n10113_0;
	wire [1:0] w_n10114_0;
	wire [2:0] w_n10116_0;
	wire [2:0] w_n10119_0;
	wire [1:0] w_n10119_1;
	wire [1:0] w_n10120_0;
	wire [1:0] w_n10123_0;
	wire [2:0] w_n10125_0;
	wire [1:0] w_n10125_1;
	wire [1:0] w_n10130_0;
	wire [1:0] w_n10132_0;
	wire [2:0] w_n10134_0;
	wire [1:0] w_n10134_1;
	wire [1:0] w_n10135_0;
	wire [2:0] w_n10136_0;
	wire [1:0] w_n10137_0;
	wire [2:0] w_n10139_0;
	wire [1:0] w_n10140_0;
	wire [1:0] w_n10188_0;
	wire [1:0] w_n10323_0;
	wire [2:0] w_n10328_0;
	wire [2:0] w_n10328_1;
	wire [2:0] w_n10328_2;
	wire [2:0] w_n10328_3;
	wire [2:0] w_n10328_4;
	wire [2:0] w_n10328_5;
	wire [2:0] w_n10328_6;
	wire [2:0] w_n10328_7;
	wire [2:0] w_n10328_8;
	wire [2:0] w_n10328_9;
	wire [2:0] w_n10328_10;
	wire [2:0] w_n10328_11;
	wire [2:0] w_n10328_12;
	wire [2:0] w_n10328_13;
	wire [2:0] w_n10328_14;
	wire [2:0] w_n10328_15;
	wire [2:0] w_n10328_16;
	wire [2:0] w_n10328_17;
	wire [2:0] w_n10328_18;
	wire [2:0] w_n10328_19;
	wire [2:0] w_n10328_20;
	wire [2:0] w_n10328_21;
	wire [2:0] w_n10328_22;
	wire [2:0] w_n10328_23;
	wire [2:0] w_n10328_24;
	wire [2:0] w_n10328_25;
	wire [2:0] w_n10328_26;
	wire [2:0] w_n10328_27;
	wire [2:0] w_n10328_28;
	wire [2:0] w_n10328_29;
	wire [2:0] w_n10328_30;
	wire [1:0] w_n10329_0;
	wire [1:0] w_n10330_0;
	wire [2:0] w_n10332_0;
	wire [1:0] w_n10333_0;
	wire [1:0] w_n10339_0;
	wire [1:0] w_n10340_0;
	wire [2:0] w_n10342_0;
	wire [1:0] w_n10343_0;
	wire [1:0] w_n10347_0;
	wire [2:0] w_n10349_0;
	wire [1:0] w_n10350_0;
	wire [1:0] w_n10354_0;
	wire [1:0] w_n10355_0;
	wire [2:0] w_n10357_0;
	wire [1:0] w_n10358_0;
	wire [1:0] w_n10362_0;
	wire [2:0] w_n10364_0;
	wire [1:0] w_n10365_0;
	wire [1:0] w_n10369_0;
	wire [1:0] w_n10370_0;
	wire [2:0] w_n10372_0;
	wire [1:0] w_n10373_0;
	wire [1:0] w_n10377_0;
	wire [1:0] w_n10378_0;
	wire [2:0] w_n10380_0;
	wire [1:0] w_n10381_0;
	wire [1:0] w_n10385_0;
	wire [1:0] w_n10386_0;
	wire [2:0] w_n10388_0;
	wire [1:0] w_n10389_0;
	wire [1:0] w_n10393_0;
	wire [2:0] w_n10395_0;
	wire [1:0] w_n10396_0;
	wire [1:0] w_n10400_0;
	wire [1:0] w_n10401_0;
	wire [2:0] w_n10403_0;
	wire [1:0] w_n10404_0;
	wire [1:0] w_n10408_0;
	wire [1:0] w_n10409_0;
	wire [2:0] w_n10411_0;
	wire [1:0] w_n10412_0;
	wire [1:0] w_n10416_0;
	wire [1:0] w_n10417_0;
	wire [2:0] w_n10419_0;
	wire [1:0] w_n10420_0;
	wire [1:0] w_n10424_0;
	wire [1:0] w_n10425_0;
	wire [2:0] w_n10427_0;
	wire [1:0] w_n10428_0;
	wire [1:0] w_n10432_0;
	wire [1:0] w_n10433_0;
	wire [2:0] w_n10435_0;
	wire [1:0] w_n10436_0;
	wire [1:0] w_n10439_0;
	wire [2:0] w_n10442_0;
	wire [1:0] w_n10443_0;
	wire [1:0] w_n10447_0;
	wire [1:0] w_n10448_0;
	wire [2:0] w_n10450_0;
	wire [1:0] w_n10451_0;
	wire [1:0] w_n10455_0;
	wire [2:0] w_n10457_0;
	wire [1:0] w_n10458_0;
	wire [1:0] w_n10462_0;
	wire [1:0] w_n10463_0;
	wire [2:0] w_n10465_0;
	wire [1:0] w_n10466_0;
	wire [1:0] w_n10470_0;
	wire [2:0] w_n10472_0;
	wire [1:0] w_n10473_0;
	wire [1:0] w_n10477_0;
	wire [1:0] w_n10478_0;
	wire [2:0] w_n10480_0;
	wire [1:0] w_n10481_0;
	wire [1:0] w_n10485_0;
	wire [1:0] w_n10486_0;
	wire [2:0] w_n10488_0;
	wire [1:0] w_n10489_0;
	wire [1:0] w_n10493_0;
	wire [1:0] w_n10494_0;
	wire [2:0] w_n10496_0;
	wire [1:0] w_n10497_0;
	wire [1:0] w_n10501_0;
	wire [2:0] w_n10503_0;
	wire [1:0] w_n10504_0;
	wire [1:0] w_n10508_0;
	wire [1:0] w_n10509_0;
	wire [2:0] w_n10511_0;
	wire [1:0] w_n10512_0;
	wire [1:0] w_n10516_0;
	wire [2:0] w_n10518_0;
	wire [1:0] w_n10519_0;
	wire [1:0] w_n10523_0;
	wire [1:0] w_n10524_0;
	wire [2:0] w_n10526_0;
	wire [1:0] w_n10527_0;
	wire [1:0] w_n10531_0;
	wire [2:0] w_n10533_0;
	wire [1:0] w_n10534_0;
	wire [1:0] w_n10538_0;
	wire [1:0] w_n10539_0;
	wire [2:0] w_n10541_0;
	wire [1:0] w_n10542_0;
	wire [1:0] w_n10546_0;
	wire [2:0] w_n10548_0;
	wire [1:0] w_n10549_0;
	wire [1:0] w_n10553_0;
	wire [2:0] w_n10555_0;
	wire [1:0] w_n10556_0;
	wire [1:0] w_n10560_0;
	wire [2:0] w_n10562_0;
	wire [1:0] w_n10563_0;
	wire [1:0] w_n10567_0;
	wire [1:0] w_n10568_0;
	wire [2:0] w_n10570_0;
	wire [1:0] w_n10571_0;
	wire [1:0] w_n10575_0;
	wire [1:0] w_n10576_0;
	wire [2:0] w_n10578_0;
	wire [1:0] w_n10579_0;
	wire [1:0] w_n10583_0;
	wire [1:0] w_n10584_0;
	wire [2:0] w_n10586_0;
	wire [1:0] w_n10587_0;
	wire [1:0] w_n10591_0;
	wire [2:0] w_n10593_0;
	wire [1:0] w_n10594_0;
	wire [1:0] w_n10598_0;
	wire [1:0] w_n10599_0;
	wire [2:0] w_n10601_0;
	wire [1:0] w_n10602_0;
	wire [1:0] w_n10606_0;
	wire [1:0] w_n10607_0;
	wire [2:0] w_n10609_0;
	wire [1:0] w_n10610_0;
	wire [1:0] w_n10635_0;
	wire [1:0] w_n10664_0;
	wire [1:0] w_n10671_0;
	wire [1:0] w_n10684_0;
	wire [1:0] w_n10709_0;
	wire [1:0] w_n10716_0;
	wire [1:0] w_n10729_0;
	wire [1:0] w_n10736_0;
	wire [1:0] w_n10743_0;
	wire [1:0] w_n10750_0;
	wire [1:0] w_n10754_0;
	wire [1:0] w_n10758_0;
	wire [1:0] w_n10771_0;
	wire [1:0] w_n10783_0;
	wire [2:0] w_n10785_0;
	wire [2:0] w_n10788_0;
	wire [1:0] w_n10788_1;
	wire [1:0] w_n10789_0;
	wire [1:0] w_n10791_0;
	wire [1:0] w_n10793_0;
	wire [1:0] w_n10794_0;
	wire [2:0] w_n10795_0;
	wire [1:0] w_n10801_0;
	wire [1:0] w_n10802_0;
	wire [2:0] w_n10805_0;
	wire [2:0] w_n10805_1;
	wire [1:0] w_n10806_0;
	wire [2:0] w_n10807_0;
	wire [1:0] w_n10808_0;
	wire [1:0] w_n10811_0;
	wire [1:0] w_n10813_0;
	wire [1:0] w_n10814_0;
	wire [1:0] w_n10815_0;
	wire [2:0] w_n10820_0;
	wire [2:0] w_n10824_0;
	wire [2:0] w_n10824_1;
	wire [2:0] w_n10824_2;
	wire [2:0] w_n10824_3;
	wire [2:0] w_n10824_4;
	wire [2:0] w_n10824_5;
	wire [2:0] w_n10824_6;
	wire [2:0] w_n10824_7;
	wire [2:0] w_n10824_8;
	wire [2:0] w_n10824_9;
	wire [2:0] w_n10824_10;
	wire [2:0] w_n10824_11;
	wire [2:0] w_n10824_12;
	wire [2:0] w_n10824_13;
	wire [2:0] w_n10824_14;
	wire [2:0] w_n10824_15;
	wire [2:0] w_n10824_16;
	wire [2:0] w_n10824_17;
	wire [2:0] w_n10824_18;
	wire [2:0] w_n10824_19;
	wire [2:0] w_n10824_20;
	wire [2:0] w_n10824_21;
	wire [2:0] w_n10824_22;
	wire [2:0] w_n10824_23;
	wire [2:0] w_n10824_24;
	wire [2:0] w_n10824_25;
	wire [2:0] w_n10824_26;
	wire [2:0] w_n10824_27;
	wire [2:0] w_n10824_28;
	wire [2:0] w_n10824_29;
	wire [2:0] w_n10824_30;
	wire [2:0] w_n10824_31;
	wire [2:0] w_n10824_32;
	wire [2:0] w_n10824_33;
	wire [2:0] w_n10824_34;
	wire [2:0] w_n10824_35;
	wire [2:0] w_n10824_36;
	wire [2:0] w_n10824_37;
	wire [2:0] w_n10824_38;
	wire [2:0] w_n10824_39;
	wire [2:0] w_n10824_40;
	wire [2:0] w_n10824_41;
	wire [2:0] w_n10824_42;
	wire [2:0] w_n10824_43;
	wire [2:0] w_n10824_44;
	wire [2:0] w_n10824_45;
	wire [2:0] w_n10824_46;
	wire [2:0] w_n10824_47;
	wire [2:0] w_n10826_0;
	wire [1:0] w_n10827_0;
	wire [2:0] w_n10834_0;
	wire [1:0] w_n10835_0;
	wire [1:0] w_n10838_0;
	wire [2:0] w_n10843_0;
	wire [2:0] w_n10845_0;
	wire [1:0] w_n10846_0;
	wire [2:0] w_n10850_0;
	wire [2:0] w_n10852_0;
	wire [1:0] w_n10853_0;
	wire [2:0] w_n10857_0;
	wire [2:0] w_n10859_0;
	wire [1:0] w_n10860_0;
	wire [2:0] w_n10864_0;
	wire [2:0] w_n10867_0;
	wire [1:0] w_n10868_0;
	wire [2:0] w_n10872_0;
	wire [2:0] w_n10874_0;
	wire [1:0] w_n10875_0;
	wire [2:0] w_n10879_0;
	wire [2:0] w_n10882_0;
	wire [1:0] w_n10883_0;
	wire [2:0] w_n10887_0;
	wire [2:0] w_n10889_0;
	wire [1:0] w_n10890_0;
	wire [2:0] w_n10894_0;
	wire [2:0] w_n10896_0;
	wire [1:0] w_n10897_0;
	wire [2:0] w_n10901_0;
	wire [2:0] w_n10903_0;
	wire [1:0] w_n10904_0;
	wire [2:0] w_n10908_0;
	wire [2:0] w_n10911_0;
	wire [1:0] w_n10912_0;
	wire [2:0] w_n10916_0;
	wire [2:0] w_n10918_0;
	wire [1:0] w_n10919_0;
	wire [2:0] w_n10923_0;
	wire [2:0] w_n10925_0;
	wire [1:0] w_n10926_0;
	wire [2:0] w_n10930_0;
	wire [2:0] w_n10932_0;
	wire [1:0] w_n10933_0;
	wire [2:0] w_n10937_0;
	wire [2:0] w_n10939_0;
	wire [1:0] w_n10940_0;
	wire [2:0] w_n10944_0;
	wire [2:0] w_n10946_0;
	wire [1:0] w_n10947_0;
	wire [2:0] w_n10950_0;
	wire [2:0] w_n10954_0;
	wire [1:0] w_n10955_0;
	wire [2:0] w_n10959_0;
	wire [2:0] w_n10961_0;
	wire [1:0] w_n10962_0;
	wire [2:0] w_n10966_0;
	wire [2:0] w_n10969_0;
	wire [1:0] w_n10970_0;
	wire [2:0] w_n10974_0;
	wire [2:0] w_n10976_0;
	wire [1:0] w_n10977_0;
	wire [2:0] w_n10981_0;
	wire [2:0] w_n10984_0;
	wire [1:0] w_n10985_0;
	wire [2:0] w_n10989_0;
	wire [2:0] w_n10991_0;
	wire [1:0] w_n10992_0;
	wire [2:0] w_n10996_0;
	wire [2:0] w_n10998_0;
	wire [1:0] w_n10999_0;
	wire [2:0] w_n11003_0;
	wire [2:0] w_n11005_0;
	wire [1:0] w_n11006_0;
	wire [2:0] w_n11010_0;
	wire [2:0] w_n11013_0;
	wire [1:0] w_n11014_0;
	wire [2:0] w_n11018_0;
	wire [2:0] w_n11020_0;
	wire [1:0] w_n11021_0;
	wire [2:0] w_n11025_0;
	wire [2:0] w_n11028_0;
	wire [1:0] w_n11029_0;
	wire [2:0] w_n11033_0;
	wire [2:0] w_n11035_0;
	wire [1:0] w_n11036_0;
	wire [2:0] w_n11040_0;
	wire [2:0] w_n11043_0;
	wire [1:0] w_n11044_0;
	wire [2:0] w_n11048_0;
	wire [2:0] w_n11050_0;
	wire [1:0] w_n11051_0;
	wire [2:0] w_n11055_0;
	wire [2:0] w_n11058_0;
	wire [1:0] w_n11059_0;
	wire [2:0] w_n11063_0;
	wire [2:0] w_n11066_0;
	wire [1:0] w_n11067_0;
	wire [2:0] w_n11071_0;
	wire [2:0] w_n11074_0;
	wire [1:0] w_n11075_0;
	wire [2:0] w_n11079_0;
	wire [2:0] w_n11081_0;
	wire [1:0] w_n11082_0;
	wire [2:0] w_n11086_0;
	wire [2:0] w_n11088_0;
	wire [1:0] w_n11089_0;
	wire [2:0] w_n11093_0;
	wire [2:0] w_n11095_0;
	wire [1:0] w_n11096_0;
	wire [2:0] w_n11100_0;
	wire [2:0] w_n11103_0;
	wire [1:0] w_n11104_0;
	wire [2:0] w_n11108_0;
	wire [2:0] w_n11110_0;
	wire [1:0] w_n11111_0;
	wire [1:0] w_n11115_0;
	wire [2:0] w_n11117_0;
	wire [1:0] w_n11117_1;
	wire [2:0] w_n11120_0;
	wire [1:0] w_n11120_1;
	wire [1:0] w_n11121_0;
	wire [1:0] w_n11125_0;
	wire [1:0] w_n11126_0;
	wire [1:0] w_n11128_0;
	wire [1:0] w_n11133_0;
	wire [1:0] w_n11137_0;
	wire [2:0] w_n11140_0;
	wire [2:0] w_n11142_0;
	wire [1:0] w_n11142_1;
	wire [1:0] w_n11143_0;
	wire [2:0] w_n11144_0;
	wire [1:0] w_n11145_0;
	wire [2:0] w_n11146_0;
	wire [1:0] w_n11147_0;
	wire [1:0] w_n11152_0;
	wire [1:0] w_n11198_0;
	wire [1:0] w_n11343_0;
	wire [1:0] w_n11346_0;
	wire [2:0] w_n11347_0;
	wire [2:0] w_n11347_1;
	wire [2:0] w_n11347_2;
	wire [2:0] w_n11347_3;
	wire [2:0] w_n11347_4;
	wire [2:0] w_n11347_5;
	wire [2:0] w_n11347_6;
	wire [2:0] w_n11347_7;
	wire [2:0] w_n11347_8;
	wire [2:0] w_n11347_9;
	wire [2:0] w_n11347_10;
	wire [2:0] w_n11347_11;
	wire [2:0] w_n11347_12;
	wire [2:0] w_n11347_13;
	wire [2:0] w_n11347_14;
	wire [2:0] w_n11347_15;
	wire [2:0] w_n11347_16;
	wire [2:0] w_n11347_17;
	wire [2:0] w_n11347_18;
	wire [2:0] w_n11347_19;
	wire [2:0] w_n11347_20;
	wire [2:0] w_n11347_21;
	wire [2:0] w_n11347_22;
	wire [2:0] w_n11347_23;
	wire [2:0] w_n11347_24;
	wire [2:0] w_n11347_25;
	wire [2:0] w_n11347_26;
	wire [1:0] w_n11347_27;
	wire [2:0] w_n11351_0;
	wire [1:0] w_n11352_0;
	wire [1:0] w_n11354_0;
	wire [1:0] w_n11359_0;
	wire [1:0] w_n11360_0;
	wire [2:0] w_n11362_0;
	wire [1:0] w_n11363_0;
	wire [1:0] w_n11367_0;
	wire [2:0] w_n11369_0;
	wire [1:0] w_n11370_0;
	wire [1:0] w_n11374_0;
	wire [1:0] w_n11375_0;
	wire [2:0] w_n11377_0;
	wire [1:0] w_n11378_0;
	wire [1:0] w_n11382_0;
	wire [1:0] w_n11383_0;
	wire [2:0] w_n11385_0;
	wire [1:0] w_n11386_0;
	wire [1:0] w_n11390_0;
	wire [1:0] w_n11391_0;
	wire [2:0] w_n11393_0;
	wire [1:0] w_n11394_0;
	wire [1:0] w_n11398_0;
	wire [2:0] w_n11400_0;
	wire [1:0] w_n11401_0;
	wire [1:0] w_n11405_0;
	wire [1:0] w_n11406_0;
	wire [2:0] w_n11408_0;
	wire [1:0] w_n11409_0;
	wire [1:0] w_n11413_0;
	wire [2:0] w_n11415_0;
	wire [1:0] w_n11416_0;
	wire [1:0] w_n11420_0;
	wire [1:0] w_n11421_0;
	wire [2:0] w_n11423_0;
	wire [1:0] w_n11424_0;
	wire [1:0] w_n11428_0;
	wire [1:0] w_n11429_0;
	wire [2:0] w_n11431_0;
	wire [1:0] w_n11432_0;
	wire [1:0] w_n11436_0;
	wire [1:0] w_n11437_0;
	wire [2:0] w_n11439_0;
	wire [1:0] w_n11440_0;
	wire [1:0] w_n11444_0;
	wire [2:0] w_n11446_0;
	wire [1:0] w_n11447_0;
	wire [1:0] w_n11451_0;
	wire [1:0] w_n11452_0;
	wire [2:0] w_n11454_0;
	wire [1:0] w_n11455_0;
	wire [1:0] w_n11459_0;
	wire [1:0] w_n11460_0;
	wire [2:0] w_n11462_0;
	wire [1:0] w_n11463_0;
	wire [1:0] w_n11467_0;
	wire [1:0] w_n11468_0;
	wire [2:0] w_n11470_0;
	wire [1:0] w_n11471_0;
	wire [1:0] w_n11475_0;
	wire [1:0] w_n11476_0;
	wire [2:0] w_n11478_0;
	wire [1:0] w_n11479_0;
	wire [1:0] w_n11483_0;
	wire [1:0] w_n11484_0;
	wire [2:0] w_n11486_0;
	wire [1:0] w_n11487_0;
	wire [1:0] w_n11490_0;
	wire [2:0] w_n11493_0;
	wire [1:0] w_n11494_0;
	wire [1:0] w_n11498_0;
	wire [1:0] w_n11499_0;
	wire [2:0] w_n11501_0;
	wire [1:0] w_n11502_0;
	wire [1:0] w_n11506_0;
	wire [2:0] w_n11508_0;
	wire [1:0] w_n11509_0;
	wire [1:0] w_n11513_0;
	wire [1:0] w_n11514_0;
	wire [2:0] w_n11516_0;
	wire [1:0] w_n11517_0;
	wire [1:0] w_n11521_0;
	wire [2:0] w_n11523_0;
	wire [1:0] w_n11524_0;
	wire [1:0] w_n11528_0;
	wire [1:0] w_n11529_0;
	wire [2:0] w_n11531_0;
	wire [1:0] w_n11532_0;
	wire [1:0] w_n11536_0;
	wire [1:0] w_n11537_0;
	wire [2:0] w_n11539_0;
	wire [1:0] w_n11540_0;
	wire [1:0] w_n11544_0;
	wire [1:0] w_n11545_0;
	wire [2:0] w_n11547_0;
	wire [1:0] w_n11548_0;
	wire [1:0] w_n11552_0;
	wire [2:0] w_n11554_0;
	wire [1:0] w_n11555_0;
	wire [1:0] w_n11559_0;
	wire [1:0] w_n11560_0;
	wire [2:0] w_n11562_0;
	wire [1:0] w_n11563_0;
	wire [1:0] w_n11567_0;
	wire [2:0] w_n11569_0;
	wire [1:0] w_n11570_0;
	wire [1:0] w_n11574_0;
	wire [1:0] w_n11575_0;
	wire [2:0] w_n11577_0;
	wire [1:0] w_n11578_0;
	wire [1:0] w_n11582_0;
	wire [2:0] w_n11584_0;
	wire [1:0] w_n11585_0;
	wire [1:0] w_n11589_0;
	wire [1:0] w_n11590_0;
	wire [2:0] w_n11592_0;
	wire [1:0] w_n11593_0;
	wire [1:0] w_n11597_0;
	wire [2:0] w_n11599_0;
	wire [1:0] w_n11600_0;
	wire [1:0] w_n11604_0;
	wire [2:0] w_n11606_0;
	wire [1:0] w_n11607_0;
	wire [1:0] w_n11611_0;
	wire [2:0] w_n11613_0;
	wire [1:0] w_n11614_0;
	wire [1:0] w_n11618_0;
	wire [1:0] w_n11619_0;
	wire [2:0] w_n11621_0;
	wire [1:0] w_n11622_0;
	wire [1:0] w_n11626_0;
	wire [1:0] w_n11627_0;
	wire [2:0] w_n11629_0;
	wire [1:0] w_n11630_0;
	wire [1:0] w_n11634_0;
	wire [1:0] w_n11635_0;
	wire [2:0] w_n11637_0;
	wire [1:0] w_n11638_0;
	wire [1:0] w_n11642_0;
	wire [2:0] w_n11644_0;
	wire [1:0] w_n11645_0;
	wire [2:0] w_n11649_0;
	wire [1:0] w_n11652_0;
	wire [2:0] w_n11653_0;
	wire [1:0] w_n11653_1;
	wire [2:0] w_n11654_0;
	wire [1:0] w_n11679_0;
	wire [1:0] w_n11704_0;
	wire [1:0] w_n11711_0;
	wire [1:0] w_n11724_0;
	wire [1:0] w_n11731_0;
	wire [1:0] w_n11744_0;
	wire [1:0] w_n11769_0;
	wire [1:0] w_n11776_0;
	wire [1:0] w_n11789_0;
	wire [1:0] w_n11796_0;
	wire [1:0] w_n11803_0;
	wire [1:0] w_n11810_0;
	wire [1:0] w_n11814_0;
	wire [1:0] w_n11818_0;
	wire [1:0] w_n11831_0;
	wire [1:0] w_n11836_0;
	wire [1:0] w_n11837_0;
	wire [1:0] w_n11838_0;
	wire [1:0] w_n11840_0;
	wire [1:0] w_n11842_0;
	wire [1:0] w_n11845_0;
	wire [1:0] w_n11846_0;
	wire [1:0] w_n11847_0;
	wire [1:0] w_n11851_0;
	wire [1:0] w_n11856_0;
	wire [2:0] w_n11858_0;
	wire [2:0] w_n11858_1;
	wire [2:0] w_n11858_2;
	wire [2:0] w_n11858_3;
	wire [2:0] w_n11858_4;
	wire [2:0] w_n11858_5;
	wire [2:0] w_n11858_6;
	wire [2:0] w_n11858_7;
	wire [2:0] w_n11858_8;
	wire [2:0] w_n11858_9;
	wire [2:0] w_n11858_10;
	wire [2:0] w_n11858_11;
	wire [2:0] w_n11858_12;
	wire [2:0] w_n11858_13;
	wire [2:0] w_n11858_14;
	wire [2:0] w_n11858_15;
	wire [2:0] w_n11858_16;
	wire [2:0] w_n11858_17;
	wire [2:0] w_n11858_18;
	wire [2:0] w_n11858_19;
	wire [2:0] w_n11858_20;
	wire [2:0] w_n11858_21;
	wire [2:0] w_n11858_22;
	wire [2:0] w_n11858_23;
	wire [2:0] w_n11858_24;
	wire [2:0] w_n11858_25;
	wire [2:0] w_n11858_26;
	wire [2:0] w_n11858_27;
	wire [2:0] w_n11858_28;
	wire [2:0] w_n11858_29;
	wire [2:0] w_n11858_30;
	wire [2:0] w_n11858_31;
	wire [2:0] w_n11858_32;
	wire [2:0] w_n11858_33;
	wire [2:0] w_n11858_34;
	wire [2:0] w_n11858_35;
	wire [2:0] w_n11858_36;
	wire [2:0] w_n11858_37;
	wire [2:0] w_n11858_38;
	wire [2:0] w_n11858_39;
	wire [2:0] w_n11858_40;
	wire [2:0] w_n11858_41;
	wire [2:0] w_n11858_42;
	wire [2:0] w_n11858_43;
	wire [2:0] w_n11858_44;
	wire [1:0] w_n11858_45;
	wire [1:0] w_n11861_0;
	wire [2:0] w_n11862_0;
	wire [2:0] w_n11864_0;
	wire [2:0] w_n11864_1;
	wire [1:0] w_n11865_0;
	wire [2:0] w_n11866_0;
	wire [1:0] w_n11867_0;
	wire [2:0] w_n11869_0;
	wire [1:0] w_n11870_0;
	wire [2:0] w_n11877_0;
	wire [1:0] w_n11878_0;
	wire [1:0] w_n11881_0;
	wire [2:0] w_n11886_0;
	wire [2:0] w_n11888_0;
	wire [1:0] w_n11889_0;
	wire [2:0] w_n11893_0;
	wire [2:0] w_n11896_0;
	wire [1:0] w_n11897_0;
	wire [2:0] w_n11901_0;
	wire [2:0] w_n11903_0;
	wire [1:0] w_n11904_0;
	wire [2:0] w_n11908_0;
	wire [2:0] w_n11911_0;
	wire [1:0] w_n11912_0;
	wire [2:0] w_n11916_0;
	wire [2:0] w_n11918_0;
	wire [1:0] w_n11919_0;
	wire [2:0] w_n11923_0;
	wire [2:0] w_n11925_0;
	wire [1:0] w_n11926_0;
	wire [2:0] w_n11930_0;
	wire [2:0] w_n11932_0;
	wire [1:0] w_n11933_0;
	wire [2:0] w_n11937_0;
	wire [2:0] w_n11940_0;
	wire [1:0] w_n11941_0;
	wire [2:0] w_n11945_0;
	wire [2:0] w_n11947_0;
	wire [1:0] w_n11948_0;
	wire [2:0] w_n11952_0;
	wire [2:0] w_n11955_0;
	wire [1:0] w_n11956_0;
	wire [2:0] w_n11960_0;
	wire [2:0] w_n11962_0;
	wire [1:0] w_n11963_0;
	wire [2:0] w_n11967_0;
	wire [2:0] w_n11969_0;
	wire [1:0] w_n11970_0;
	wire [2:0] w_n11974_0;
	wire [2:0] w_n11976_0;
	wire [1:0] w_n11977_0;
	wire [2:0] w_n11981_0;
	wire [2:0] w_n11984_0;
	wire [1:0] w_n11985_0;
	wire [2:0] w_n11989_0;
	wire [2:0] w_n11991_0;
	wire [1:0] w_n11992_0;
	wire [2:0] w_n11996_0;
	wire [2:0] w_n11998_0;
	wire [1:0] w_n11999_0;
	wire [2:0] w_n12003_0;
	wire [2:0] w_n12005_0;
	wire [1:0] w_n12006_0;
	wire [2:0] w_n12010_0;
	wire [2:0] w_n12012_0;
	wire [1:0] w_n12013_0;
	wire [2:0] w_n12017_0;
	wire [2:0] w_n12019_0;
	wire [1:0] w_n12020_0;
	wire [2:0] w_n12023_0;
	wire [2:0] w_n12027_0;
	wire [1:0] w_n12028_0;
	wire [2:0] w_n12032_0;
	wire [2:0] w_n12034_0;
	wire [1:0] w_n12035_0;
	wire [2:0] w_n12039_0;
	wire [2:0] w_n12042_0;
	wire [1:0] w_n12043_0;
	wire [2:0] w_n12047_0;
	wire [2:0] w_n12049_0;
	wire [1:0] w_n12050_0;
	wire [2:0] w_n12054_0;
	wire [2:0] w_n12057_0;
	wire [1:0] w_n12058_0;
	wire [2:0] w_n12062_0;
	wire [2:0] w_n12064_0;
	wire [1:0] w_n12065_0;
	wire [2:0] w_n12069_0;
	wire [2:0] w_n12071_0;
	wire [1:0] w_n12072_0;
	wire [2:0] w_n12076_0;
	wire [2:0] w_n12078_0;
	wire [1:0] w_n12079_0;
	wire [2:0] w_n12083_0;
	wire [2:0] w_n12086_0;
	wire [1:0] w_n12087_0;
	wire [2:0] w_n12091_0;
	wire [2:0] w_n12093_0;
	wire [1:0] w_n12094_0;
	wire [2:0] w_n12098_0;
	wire [2:0] w_n12101_0;
	wire [1:0] w_n12102_0;
	wire [2:0] w_n12106_0;
	wire [2:0] w_n12108_0;
	wire [1:0] w_n12109_0;
	wire [2:0] w_n12113_0;
	wire [2:0] w_n12116_0;
	wire [1:0] w_n12117_0;
	wire [2:0] w_n12121_0;
	wire [2:0] w_n12123_0;
	wire [1:0] w_n12124_0;
	wire [2:0] w_n12128_0;
	wire [2:0] w_n12131_0;
	wire [1:0] w_n12132_0;
	wire [2:0] w_n12136_0;
	wire [2:0] w_n12139_0;
	wire [1:0] w_n12140_0;
	wire [2:0] w_n12144_0;
	wire [2:0] w_n12147_0;
	wire [1:0] w_n12148_0;
	wire [2:0] w_n12152_0;
	wire [2:0] w_n12154_0;
	wire [1:0] w_n12155_0;
	wire [2:0] w_n12159_0;
	wire [2:0] w_n12161_0;
	wire [1:0] w_n12162_0;
	wire [2:0] w_n12166_0;
	wire [2:0] w_n12168_0;
	wire [1:0] w_n12169_0;
	wire [2:0] w_n12173_0;
	wire [2:0] w_n12176_0;
	wire [2:0] w_n12177_0;
	wire [1:0] w_n12179_0;
	wire [1:0] w_n12180_0;
	wire [1:0] w_n12187_0;
	wire [1:0] w_n12188_0;
	wire [1:0] w_n12190_0;
	wire [2:0] w_n12195_0;
	wire [2:0] w_n12196_0;
	wire [2:0] w_n12196_1;
	wire [1:0] w_n12197_0;
	wire [2:0] w_n12198_0;
	wire [1:0] w_n12199_0;
	wire [2:0] w_n12201_0;
	wire [1:0] w_n12202_0;
	wire [2:0] w_n12207_0;
	wire [1:0] w_n12207_1;
	wire [1:0] w_n12256_0;
	wire [1:0] w_n12404_0;
	wire [1:0] w_n12407_0;
	wire [1:0] w_n12408_0;
	wire [2:0] w_n12410_0;
	wire [2:0] w_n12410_1;
	wire [2:0] w_n12410_2;
	wire [2:0] w_n12410_3;
	wire [2:0] w_n12410_4;
	wire [2:0] w_n12410_5;
	wire [2:0] w_n12410_6;
	wire [2:0] w_n12410_7;
	wire [2:0] w_n12410_8;
	wire [2:0] w_n12410_9;
	wire [2:0] w_n12410_10;
	wire [2:0] w_n12410_11;
	wire [2:0] w_n12410_12;
	wire [2:0] w_n12410_13;
	wire [2:0] w_n12410_14;
	wire [2:0] w_n12410_15;
	wire [2:0] w_n12410_16;
	wire [2:0] w_n12410_17;
	wire [2:0] w_n12410_18;
	wire [2:0] w_n12410_19;
	wire [2:0] w_n12410_20;
	wire [2:0] w_n12410_21;
	wire [2:0] w_n12410_22;
	wire [2:0] w_n12410_23;
	wire [2:0] w_n12410_24;
	wire [1:0] w_n12410_25;
	wire [2:0] w_n12414_0;
	wire [1:0] w_n12415_0;
	wire [1:0] w_n12417_0;
	wire [1:0] w_n12422_0;
	wire [1:0] w_n12423_0;
	wire [2:0] w_n12425_0;
	wire [1:0] w_n12426_0;
	wire [1:0] w_n12430_0;
	wire [2:0] w_n12432_0;
	wire [1:0] w_n12433_0;
	wire [1:0] w_n12437_0;
	wire [1:0] w_n12438_0;
	wire [2:0] w_n12440_0;
	wire [1:0] w_n12441_0;
	wire [1:0] w_n12445_0;
	wire [2:0] w_n12447_0;
	wire [1:0] w_n12448_0;
	wire [1:0] w_n12452_0;
	wire [1:0] w_n12453_0;
	wire [2:0] w_n12455_0;
	wire [1:0] w_n12456_0;
	wire [1:0] w_n12460_0;
	wire [2:0] w_n12462_0;
	wire [1:0] w_n12463_0;
	wire [1:0] w_n12467_0;
	wire [1:0] w_n12468_0;
	wire [2:0] w_n12470_0;
	wire [1:0] w_n12471_0;
	wire [1:0] w_n12475_0;
	wire [1:0] w_n12476_0;
	wire [2:0] w_n12478_0;
	wire [1:0] w_n12479_0;
	wire [1:0] w_n12483_0;
	wire [1:0] w_n12484_0;
	wire [2:0] w_n12486_0;
	wire [1:0] w_n12487_0;
	wire [1:0] w_n12491_0;
	wire [2:0] w_n12493_0;
	wire [1:0] w_n12494_0;
	wire [1:0] w_n12498_0;
	wire [1:0] w_n12499_0;
	wire [2:0] w_n12501_0;
	wire [1:0] w_n12502_0;
	wire [1:0] w_n12506_0;
	wire [2:0] w_n12508_0;
	wire [1:0] w_n12509_0;
	wire [1:0] w_n12513_0;
	wire [1:0] w_n12514_0;
	wire [2:0] w_n12516_0;
	wire [1:0] w_n12517_0;
	wire [1:0] w_n12521_0;
	wire [1:0] w_n12522_0;
	wire [2:0] w_n12524_0;
	wire [1:0] w_n12525_0;
	wire [1:0] w_n12529_0;
	wire [1:0] w_n12530_0;
	wire [2:0] w_n12532_0;
	wire [1:0] w_n12533_0;
	wire [1:0] w_n12537_0;
	wire [2:0] w_n12539_0;
	wire [1:0] w_n12540_0;
	wire [1:0] w_n12544_0;
	wire [1:0] w_n12545_0;
	wire [2:0] w_n12547_0;
	wire [1:0] w_n12548_0;
	wire [1:0] w_n12552_0;
	wire [1:0] w_n12553_0;
	wire [2:0] w_n12555_0;
	wire [1:0] w_n12556_0;
	wire [1:0] w_n12560_0;
	wire [1:0] w_n12561_0;
	wire [2:0] w_n12563_0;
	wire [1:0] w_n12564_0;
	wire [1:0] w_n12568_0;
	wire [1:0] w_n12569_0;
	wire [2:0] w_n12571_0;
	wire [1:0] w_n12572_0;
	wire [2:0] w_n12576_0;
	wire [2:0] w_n12579_0;
	wire [1:0] w_n12580_0;
	wire [1:0] w_n12583_0;
	wire [2:0] w_n12586_0;
	wire [1:0] w_n12587_0;
	wire [1:0] w_n12591_0;
	wire [1:0] w_n12592_0;
	wire [2:0] w_n12594_0;
	wire [1:0] w_n12595_0;
	wire [1:0] w_n12599_0;
	wire [2:0] w_n12601_0;
	wire [1:0] w_n12602_0;
	wire [1:0] w_n12606_0;
	wire [1:0] w_n12607_0;
	wire [2:0] w_n12609_0;
	wire [1:0] w_n12610_0;
	wire [1:0] w_n12614_0;
	wire [2:0] w_n12616_0;
	wire [1:0] w_n12617_0;
	wire [1:0] w_n12621_0;
	wire [1:0] w_n12622_0;
	wire [2:0] w_n12624_0;
	wire [1:0] w_n12625_0;
	wire [1:0] w_n12629_0;
	wire [1:0] w_n12630_0;
	wire [2:0] w_n12632_0;
	wire [1:0] w_n12633_0;
	wire [1:0] w_n12637_0;
	wire [1:0] w_n12638_0;
	wire [2:0] w_n12640_0;
	wire [1:0] w_n12641_0;
	wire [1:0] w_n12645_0;
	wire [2:0] w_n12647_0;
	wire [1:0] w_n12648_0;
	wire [1:0] w_n12652_0;
	wire [1:0] w_n12653_0;
	wire [2:0] w_n12655_0;
	wire [1:0] w_n12656_0;
	wire [1:0] w_n12660_0;
	wire [2:0] w_n12662_0;
	wire [1:0] w_n12663_0;
	wire [1:0] w_n12667_0;
	wire [1:0] w_n12668_0;
	wire [2:0] w_n12670_0;
	wire [1:0] w_n12671_0;
	wire [1:0] w_n12675_0;
	wire [2:0] w_n12677_0;
	wire [1:0] w_n12678_0;
	wire [1:0] w_n12682_0;
	wire [1:0] w_n12683_0;
	wire [2:0] w_n12685_0;
	wire [1:0] w_n12686_0;
	wire [1:0] w_n12690_0;
	wire [2:0] w_n12692_0;
	wire [1:0] w_n12693_0;
	wire [1:0] w_n12697_0;
	wire [2:0] w_n12699_0;
	wire [1:0] w_n12700_0;
	wire [1:0] w_n12704_0;
	wire [2:0] w_n12706_0;
	wire [1:0] w_n12707_0;
	wire [1:0] w_n12711_0;
	wire [1:0] w_n12712_0;
	wire [2:0] w_n12714_0;
	wire [1:0] w_n12715_0;
	wire [1:0] w_n12719_0;
	wire [1:0] w_n12720_0;
	wire [2:0] w_n12722_0;
	wire [1:0] w_n12723_0;
	wire [2:0] w_n12727_0;
	wire [1:0] w_n12730_0;
	wire [2:0] w_n12731_0;
	wire [1:0] w_n12731_1;
	wire [2:0] w_n12732_0;
	wire [1:0] w_n12736_0;
	wire [1:0] w_n12737_0;
	wire [1:0] w_n12738_0;
	wire [1:0] w_n12739_0;
	wire [1:0] w_n12760_0;
	wire [1:0] w_n12789_0;
	wire [1:0] w_n12796_0;
	wire [1:0] w_n12803_0;
	wire [1:0] w_n12810_0;
	wire [1:0] w_n12823_0;
	wire [1:0] w_n12830_0;
	wire [1:0] w_n12843_0;
	wire [1:0] w_n12868_0;
	wire [1:0] w_n12875_0;
	wire [1:0] w_n12888_0;
	wire [1:0] w_n12895_0;
	wire [1:0] w_n12902_0;
	wire [1:0] w_n12909_0;
	wire [1:0] w_n12913_0;
	wire [1:0] w_n12917_0;
	wire [1:0] w_n12928_0;
	wire [1:0] w_n12929_0;
	wire [1:0] w_n12932_0;
	wire [1:0] w_n12933_0;
	wire [1:0] w_n12935_0;
	wire [1:0] w_n12937_0;
	wire [1:0] w_n12938_0;
	wire [1:0] w_n12946_0;
	wire [2:0] w_n12947_0;
	wire [2:0] w_n12947_1;
	wire [2:0] w_n12947_2;
	wire [2:0] w_n12947_3;
	wire [2:0] w_n12947_4;
	wire [2:0] w_n12947_5;
	wire [2:0] w_n12947_6;
	wire [2:0] w_n12947_7;
	wire [2:0] w_n12947_8;
	wire [2:0] w_n12947_9;
	wire [2:0] w_n12947_10;
	wire [2:0] w_n12947_11;
	wire [2:0] w_n12947_12;
	wire [2:0] w_n12947_13;
	wire [2:0] w_n12947_14;
	wire [2:0] w_n12947_15;
	wire [2:0] w_n12947_16;
	wire [2:0] w_n12947_17;
	wire [2:0] w_n12947_18;
	wire [2:0] w_n12947_19;
	wire [2:0] w_n12947_20;
	wire [2:0] w_n12947_21;
	wire [2:0] w_n12947_22;
	wire [2:0] w_n12947_23;
	wire [2:0] w_n12947_24;
	wire [2:0] w_n12947_25;
	wire [2:0] w_n12947_26;
	wire [2:0] w_n12947_27;
	wire [2:0] w_n12947_28;
	wire [2:0] w_n12947_29;
	wire [2:0] w_n12947_30;
	wire [2:0] w_n12947_31;
	wire [2:0] w_n12947_32;
	wire [2:0] w_n12947_33;
	wire [2:0] w_n12947_34;
	wire [2:0] w_n12947_35;
	wire [2:0] w_n12947_36;
	wire [2:0] w_n12947_37;
	wire [2:0] w_n12947_38;
	wire [2:0] w_n12947_39;
	wire [2:0] w_n12947_40;
	wire [2:0] w_n12947_41;
	wire [2:0] w_n12947_42;
	wire [2:0] w_n12947_43;
	wire [2:0] w_n12947_44;
	wire [1:0] w_n12950_0;
	wire [2:0] w_n12951_0;
	wire [2:0] w_n12953_0;
	wire [2:0] w_n12953_1;
	wire [1:0] w_n12954_0;
	wire [2:0] w_n12955_0;
	wire [1:0] w_n12956_0;
	wire [2:0] w_n12958_0;
	wire [1:0] w_n12959_0;
	wire [1:0] w_n12964_0;
	wire [2:0] w_n12966_0;
	wire [1:0] w_n12967_0;
	wire [1:0] w_n12970_0;
	wire [2:0] w_n12975_0;
	wire [2:0] w_n12977_0;
	wire [1:0] w_n12978_0;
	wire [2:0] w_n12982_0;
	wire [2:0] w_n12985_0;
	wire [1:0] w_n12986_0;
	wire [2:0] w_n12990_0;
	wire [2:0] w_n12992_0;
	wire [1:0] w_n12993_0;
	wire [2:0] w_n12997_0;
	wire [2:0] w_n13000_0;
	wire [1:0] w_n13001_0;
	wire [2:0] w_n13005_0;
	wire [2:0] w_n13007_0;
	wire [1:0] w_n13008_0;
	wire [2:0] w_n13012_0;
	wire [2:0] w_n13015_0;
	wire [1:0] w_n13016_0;
	wire [2:0] w_n13020_0;
	wire [2:0] w_n13022_0;
	wire [1:0] w_n13023_0;
	wire [2:0] w_n13027_0;
	wire [2:0] w_n13030_0;
	wire [1:0] w_n13031_0;
	wire [2:0] w_n13035_0;
	wire [2:0] w_n13037_0;
	wire [1:0] w_n13038_0;
	wire [2:0] w_n13042_0;
	wire [2:0] w_n13044_0;
	wire [1:0] w_n13045_0;
	wire [2:0] w_n13049_0;
	wire [2:0] w_n13051_0;
	wire [1:0] w_n13052_0;
	wire [2:0] w_n13056_0;
	wire [2:0] w_n13059_0;
	wire [1:0] w_n13060_0;
	wire [2:0] w_n13064_0;
	wire [2:0] w_n13066_0;
	wire [1:0] w_n13067_0;
	wire [2:0] w_n13071_0;
	wire [2:0] w_n13074_0;
	wire [1:0] w_n13075_0;
	wire [2:0] w_n13079_0;
	wire [2:0] w_n13081_0;
	wire [1:0] w_n13082_0;
	wire [2:0] w_n13086_0;
	wire [2:0] w_n13088_0;
	wire [1:0] w_n13089_0;
	wire [2:0] w_n13093_0;
	wire [2:0] w_n13095_0;
	wire [1:0] w_n13096_0;
	wire [2:0] w_n13100_0;
	wire [2:0] w_n13103_0;
	wire [1:0] w_n13104_0;
	wire [2:0] w_n13108_0;
	wire [2:0] w_n13110_0;
	wire [1:0] w_n13111_0;
	wire [2:0] w_n13115_0;
	wire [2:0] w_n13117_0;
	wire [1:0] w_n13118_0;
	wire [2:0] w_n13122_0;
	wire [2:0] w_n13124_0;
	wire [1:0] w_n13125_0;
	wire [2:0] w_n13129_0;
	wire [2:0] w_n13131_0;
	wire [1:0] w_n13132_0;
	wire [2:0] w_n13136_0;
	wire [2:0] w_n13139_0;
	wire [1:0] w_n13140_0;
	wire [2:0] w_n13143_0;
	wire [2:0] w_n13147_0;
	wire [1:0] w_n13148_0;
	wire [2:0] w_n13152_0;
	wire [2:0] w_n13154_0;
	wire [1:0] w_n13155_0;
	wire [2:0] w_n13159_0;
	wire [2:0] w_n13162_0;
	wire [1:0] w_n13163_0;
	wire [2:0] w_n13167_0;
	wire [2:0] w_n13169_0;
	wire [1:0] w_n13170_0;
	wire [2:0] w_n13174_0;
	wire [2:0] w_n13177_0;
	wire [1:0] w_n13178_0;
	wire [2:0] w_n13182_0;
	wire [2:0] w_n13184_0;
	wire [1:0] w_n13185_0;
	wire [2:0] w_n13189_0;
	wire [2:0] w_n13191_0;
	wire [1:0] w_n13192_0;
	wire [2:0] w_n13196_0;
	wire [2:0] w_n13198_0;
	wire [1:0] w_n13199_0;
	wire [2:0] w_n13203_0;
	wire [2:0] w_n13206_0;
	wire [1:0] w_n13207_0;
	wire [2:0] w_n13211_0;
	wire [2:0] w_n13213_0;
	wire [1:0] w_n13214_0;
	wire [2:0] w_n13218_0;
	wire [2:0] w_n13221_0;
	wire [1:0] w_n13222_0;
	wire [2:0] w_n13226_0;
	wire [2:0] w_n13228_0;
	wire [1:0] w_n13229_0;
	wire [2:0] w_n13233_0;
	wire [2:0] w_n13236_0;
	wire [1:0] w_n13237_0;
	wire [2:0] w_n13241_0;
	wire [2:0] w_n13243_0;
	wire [1:0] w_n13244_0;
	wire [2:0] w_n13248_0;
	wire [2:0] w_n13251_0;
	wire [1:0] w_n13252_0;
	wire [2:0] w_n13256_0;
	wire [2:0] w_n13259_0;
	wire [1:0] w_n13260_0;
	wire [2:0] w_n13264_0;
	wire [2:0] w_n13267_0;
	wire [1:0] w_n13268_0;
	wire [2:0] w_n13272_0;
	wire [2:0] w_n13274_0;
	wire [1:0] w_n13275_0;
	wire [2:0] w_n13279_0;
	wire [2:0] w_n13281_0;
	wire [1:0] w_n13282_0;
	wire [1:0] w_n13285_0;
	wire [2:0] w_n13287_0;
	wire [1:0] w_n13287_1;
	wire [1:0] w_n13292_0;
	wire [1:0] w_n13294_0;
	wire [2:0] w_n13296_0;
	wire [1:0] w_n13296_1;
	wire [1:0] w_n13297_0;
	wire [2:0] w_n13298_0;
	wire [1:0] w_n13299_0;
	wire [2:0] w_n13301_0;
	wire [1:0] w_n13302_0;
	wire [1:0] w_n13510_0;
	wire [2:0] w_n13515_0;
	wire [2:0] w_n13515_1;
	wire [2:0] w_n13515_2;
	wire [2:0] w_n13515_3;
	wire [2:0] w_n13515_4;
	wire [2:0] w_n13515_5;
	wire [2:0] w_n13515_6;
	wire [2:0] w_n13515_7;
	wire [2:0] w_n13515_8;
	wire [2:0] w_n13515_9;
	wire [2:0] w_n13515_10;
	wire [2:0] w_n13515_11;
	wire [2:0] w_n13515_12;
	wire [2:0] w_n13515_13;
	wire [2:0] w_n13515_14;
	wire [2:0] w_n13515_15;
	wire [2:0] w_n13515_16;
	wire [2:0] w_n13515_17;
	wire [2:0] w_n13515_18;
	wire [2:0] w_n13515_19;
	wire [2:0] w_n13515_20;
	wire [2:0] w_n13515_21;
	wire [2:0] w_n13515_22;
	wire [1:0] w_n13515_23;
	wire [1:0] w_n13516_0;
	wire [2:0] w_n13519_0;
	wire [1:0] w_n13520_0;
	wire [1:0] w_n13526_0;
	wire [1:0] w_n13527_0;
	wire [2:0] w_n13529_0;
	wire [1:0] w_n13530_0;
	wire [1:0] w_n13534_0;
	wire [1:0] w_n13535_0;
	wire [2:0] w_n13537_0;
	wire [1:0] w_n13538_0;
	wire [1:0] w_n13542_0;
	wire [1:0] w_n13543_0;
	wire [2:0] w_n13545_0;
	wire [1:0] w_n13546_0;
	wire [1:0] w_n13550_0;
	wire [2:0] w_n13552_0;
	wire [1:0] w_n13553_0;
	wire [1:0] w_n13557_0;
	wire [1:0] w_n13558_0;
	wire [2:0] w_n13560_0;
	wire [1:0] w_n13561_0;
	wire [1:0] w_n13565_0;
	wire [2:0] w_n13567_0;
	wire [1:0] w_n13568_0;
	wire [1:0] w_n13572_0;
	wire [1:0] w_n13573_0;
	wire [2:0] w_n13575_0;
	wire [1:0] w_n13576_0;
	wire [1:0] w_n13580_0;
	wire [2:0] w_n13582_0;
	wire [1:0] w_n13583_0;
	wire [1:0] w_n13587_0;
	wire [1:0] w_n13588_0;
	wire [2:0] w_n13590_0;
	wire [1:0] w_n13591_0;
	wire [1:0] w_n13595_0;
	wire [2:0] w_n13597_0;
	wire [1:0] w_n13598_0;
	wire [1:0] w_n13602_0;
	wire [1:0] w_n13603_0;
	wire [2:0] w_n13605_0;
	wire [1:0] w_n13606_0;
	wire [1:0] w_n13610_0;
	wire [1:0] w_n13611_0;
	wire [2:0] w_n13613_0;
	wire [1:0] w_n13614_0;
	wire [1:0] w_n13618_0;
	wire [1:0] w_n13619_0;
	wire [2:0] w_n13621_0;
	wire [1:0] w_n13622_0;
	wire [1:0] w_n13626_0;
	wire [2:0] w_n13628_0;
	wire [1:0] w_n13629_0;
	wire [1:0] w_n13633_0;
	wire [1:0] w_n13634_0;
	wire [2:0] w_n13636_0;
	wire [1:0] w_n13637_0;
	wire [1:0] w_n13641_0;
	wire [2:0] w_n13643_0;
	wire [1:0] w_n13644_0;
	wire [1:0] w_n13648_0;
	wire [1:0] w_n13649_0;
	wire [2:0] w_n13651_0;
	wire [1:0] w_n13652_0;
	wire [1:0] w_n13656_0;
	wire [1:0] w_n13657_0;
	wire [2:0] w_n13659_0;
	wire [1:0] w_n13660_0;
	wire [1:0] w_n13664_0;
	wire [1:0] w_n13665_0;
	wire [2:0] w_n13667_0;
	wire [1:0] w_n13668_0;
	wire [1:0] w_n13672_0;
	wire [2:0] w_n13674_0;
	wire [1:0] w_n13675_0;
	wire [1:0] w_n13679_0;
	wire [1:0] w_n13680_0;
	wire [2:0] w_n13682_0;
	wire [1:0] w_n13683_0;
	wire [1:0] w_n13687_0;
	wire [1:0] w_n13688_0;
	wire [2:0] w_n13690_0;
	wire [1:0] w_n13691_0;
	wire [1:0] w_n13695_0;
	wire [1:0] w_n13696_0;
	wire [2:0] w_n13698_0;
	wire [1:0] w_n13699_0;
	wire [1:0] w_n13703_0;
	wire [1:0] w_n13704_0;
	wire [2:0] w_n13706_0;
	wire [1:0] w_n13707_0;
	wire [1:0] w_n13711_0;
	wire [2:0] w_n13713_0;
	wire [1:0] w_n13714_0;
	wire [1:0] w_n13717_0;
	wire [2:0] w_n13720_0;
	wire [1:0] w_n13721_0;
	wire [1:0] w_n13725_0;
	wire [1:0] w_n13726_0;
	wire [2:0] w_n13728_0;
	wire [1:0] w_n13729_0;
	wire [1:0] w_n13733_0;
	wire [2:0] w_n13735_0;
	wire [1:0] w_n13736_0;
	wire [1:0] w_n13740_0;
	wire [1:0] w_n13741_0;
	wire [2:0] w_n13743_0;
	wire [1:0] w_n13744_0;
	wire [1:0] w_n13748_0;
	wire [2:0] w_n13750_0;
	wire [1:0] w_n13751_0;
	wire [1:0] w_n13755_0;
	wire [1:0] w_n13756_0;
	wire [2:0] w_n13758_0;
	wire [1:0] w_n13759_0;
	wire [1:0] w_n13763_0;
	wire [1:0] w_n13764_0;
	wire [2:0] w_n13766_0;
	wire [1:0] w_n13767_0;
	wire [1:0] w_n13771_0;
	wire [1:0] w_n13772_0;
	wire [2:0] w_n13774_0;
	wire [1:0] w_n13775_0;
	wire [1:0] w_n13779_0;
	wire [2:0] w_n13781_0;
	wire [1:0] w_n13782_0;
	wire [1:0] w_n13786_0;
	wire [1:0] w_n13787_0;
	wire [2:0] w_n13789_0;
	wire [1:0] w_n13790_0;
	wire [1:0] w_n13794_0;
	wire [2:0] w_n13796_0;
	wire [1:0] w_n13797_0;
	wire [1:0] w_n13801_0;
	wire [1:0] w_n13802_0;
	wire [2:0] w_n13804_0;
	wire [1:0] w_n13805_0;
	wire [1:0] w_n13809_0;
	wire [2:0] w_n13811_0;
	wire [1:0] w_n13812_0;
	wire [1:0] w_n13816_0;
	wire [1:0] w_n13817_0;
	wire [2:0] w_n13819_0;
	wire [1:0] w_n13820_0;
	wire [1:0] w_n13824_0;
	wire [2:0] w_n13826_0;
	wire [1:0] w_n13827_0;
	wire [1:0] w_n13831_0;
	wire [2:0] w_n13833_0;
	wire [1:0] w_n13834_0;
	wire [1:0] w_n13838_0;
	wire [2:0] w_n13840_0;
	wire [1:0] w_n13841_0;
	wire [1:0] w_n13845_0;
	wire [1:0] w_n13846_0;
	wire [2:0] w_n13848_0;
	wire [1:0] w_n13851_0;
	wire [2:0] w_n13852_0;
	wire [1:0] w_n13853_0;
	wire [1:0] w_n13854_0;
	wire [1:0] w_n13859_0;
	wire [1:0] w_n13860_0;
	wire [1:0] w_n13879_0;
	wire [1:0] w_n13913_0;
	wire [1:0] w_n13926_0;
	wire [1:0] w_n13933_0;
	wire [1:0] w_n13940_0;
	wire [1:0] w_n13947_0;
	wire [1:0] w_n13960_0;
	wire [1:0] w_n13967_0;
	wire [1:0] w_n13980_0;
	wire [1:0] w_n13996_0;
	wire [1:0] w_n14006_0;
	wire [1:0] w_n14013_0;
	wire [1:0] w_n14026_0;
	wire [1:0] w_n14033_0;
	wire [1:0] w_n14040_0;
	wire [1:0] w_n14047_0;
	wire [1:0] w_n14051_0;
	wire [1:0] w_n14055_0;
	wire [1:0] w_n14060_0;
	wire [1:0] w_n14063_0;
	wire [1:0] w_n14065_0;
	wire [1:0] w_n14066_0;
	wire [1:0] w_n14077_0;
	wire [2:0] w_n14078_0;
	wire [2:0] w_n14078_1;
	wire [2:0] w_n14078_2;
	wire [2:0] w_n14078_3;
	wire [2:0] w_n14078_4;
	wire [2:0] w_n14078_5;
	wire [2:0] w_n14078_6;
	wire [2:0] w_n14078_7;
	wire [2:0] w_n14078_8;
	wire [2:0] w_n14078_9;
	wire [2:0] w_n14078_10;
	wire [2:0] w_n14078_11;
	wire [2:0] w_n14078_12;
	wire [2:0] w_n14078_13;
	wire [2:0] w_n14078_14;
	wire [2:0] w_n14078_15;
	wire [2:0] w_n14078_16;
	wire [2:0] w_n14078_17;
	wire [2:0] w_n14078_18;
	wire [2:0] w_n14078_19;
	wire [2:0] w_n14078_20;
	wire [2:0] w_n14078_21;
	wire [2:0] w_n14078_22;
	wire [2:0] w_n14078_23;
	wire [2:0] w_n14078_24;
	wire [2:0] w_n14078_25;
	wire [2:0] w_n14078_26;
	wire [2:0] w_n14078_27;
	wire [2:0] w_n14078_28;
	wire [2:0] w_n14078_29;
	wire [2:0] w_n14078_30;
	wire [2:0] w_n14078_31;
	wire [2:0] w_n14078_32;
	wire [2:0] w_n14078_33;
	wire [2:0] w_n14078_34;
	wire [2:0] w_n14078_35;
	wire [2:0] w_n14078_36;
	wire [2:0] w_n14078_37;
	wire [2:0] w_n14078_38;
	wire [2:0] w_n14078_39;
	wire [2:0] w_n14078_40;
	wire [2:0] w_n14078_41;
	wire [1:0] w_n14078_42;
	wire [2:0] w_n14080_0;
	wire [2:0] w_n14080_1;
	wire [1:0] w_n14081_0;
	wire [2:0] w_n14082_0;
	wire [1:0] w_n14083_0;
	wire [2:0] w_n14085_0;
	wire [1:0] w_n14086_0;
	wire [2:0] w_n14093_0;
	wire [1:0] w_n14094_0;
	wire [1:0] w_n14097_0;
	wire [2:0] w_n14102_0;
	wire [2:0] w_n14104_0;
	wire [1:0] w_n14105_0;
	wire [2:0] w_n14109_0;
	wire [2:0] w_n14112_0;
	wire [1:0] w_n14113_0;
	wire [2:0] w_n14117_0;
	wire [2:0] w_n14119_0;
	wire [1:0] w_n14120_0;
	wire [2:0] w_n14124_0;
	wire [2:0] w_n14126_0;
	wire [1:0] w_n14127_0;
	wire [2:0] w_n14131_0;
	wire [2:0] w_n14133_0;
	wire [1:0] w_n14134_0;
	wire [2:0] w_n14138_0;
	wire [2:0] w_n14141_0;
	wire [1:0] w_n14142_0;
	wire [2:0] w_n14146_0;
	wire [2:0] w_n14148_0;
	wire [1:0] w_n14149_0;
	wire [2:0] w_n14153_0;
	wire [2:0] w_n14156_0;
	wire [1:0] w_n14157_0;
	wire [2:0] w_n14161_0;
	wire [2:0] w_n14163_0;
	wire [1:0] w_n14164_0;
	wire [2:0] w_n14168_0;
	wire [2:0] w_n14171_0;
	wire [1:0] w_n14172_0;
	wire [2:0] w_n14176_0;
	wire [2:0] w_n14178_0;
	wire [1:0] w_n14179_0;
	wire [2:0] w_n14183_0;
	wire [2:0] w_n14186_0;
	wire [1:0] w_n14187_0;
	wire [2:0] w_n14191_0;
	wire [2:0] w_n14193_0;
	wire [1:0] w_n14194_0;
	wire [2:0] w_n14198_0;
	wire [2:0] w_n14200_0;
	wire [1:0] w_n14201_0;
	wire [2:0] w_n14205_0;
	wire [2:0] w_n14207_0;
	wire [1:0] w_n14208_0;
	wire [2:0] w_n14212_0;
	wire [2:0] w_n14215_0;
	wire [1:0] w_n14216_0;
	wire [2:0] w_n14220_0;
	wire [2:0] w_n14222_0;
	wire [1:0] w_n14223_0;
	wire [2:0] w_n14227_0;
	wire [2:0] w_n14230_0;
	wire [1:0] w_n14231_0;
	wire [2:0] w_n14235_0;
	wire [2:0] w_n14237_0;
	wire [1:0] w_n14238_0;
	wire [2:0] w_n14242_0;
	wire [2:0] w_n14244_0;
	wire [1:0] w_n14245_0;
	wire [2:0] w_n14249_0;
	wire [2:0] w_n14251_0;
	wire [1:0] w_n14252_0;
	wire [2:0] w_n14256_0;
	wire [2:0] w_n14259_0;
	wire [1:0] w_n14260_0;
	wire [2:0] w_n14264_0;
	wire [2:0] w_n14266_0;
	wire [1:0] w_n14267_0;
	wire [1:0] w_n14271_0;
	wire [2:0] w_n14273_0;
	wire [1:0] w_n14274_0;
	wire [2:0] w_n14278_0;
	wire [2:0] w_n14280_0;
	wire [1:0] w_n14281_0;
	wire [2:0] w_n14285_0;
	wire [2:0] w_n14287_0;
	wire [1:0] w_n14288_0;
	wire [2:0] w_n14292_0;
	wire [2:0] w_n14295_0;
	wire [1:0] w_n14296_0;
	wire [2:0] w_n14299_0;
	wire [2:0] w_n14303_0;
	wire [1:0] w_n14304_0;
	wire [2:0] w_n14308_0;
	wire [2:0] w_n14310_0;
	wire [1:0] w_n14311_0;
	wire [2:0] w_n14315_0;
	wire [2:0] w_n14318_0;
	wire [1:0] w_n14319_0;
	wire [2:0] w_n14323_0;
	wire [2:0] w_n14325_0;
	wire [1:0] w_n14326_0;
	wire [2:0] w_n14330_0;
	wire [2:0] w_n14333_0;
	wire [1:0] w_n14334_0;
	wire [2:0] w_n14338_0;
	wire [2:0] w_n14340_0;
	wire [1:0] w_n14341_0;
	wire [2:0] w_n14345_0;
	wire [2:0] w_n14347_0;
	wire [1:0] w_n14348_0;
	wire [2:0] w_n14352_0;
	wire [2:0] w_n14354_0;
	wire [1:0] w_n14355_0;
	wire [2:0] w_n14359_0;
	wire [2:0] w_n14362_0;
	wire [1:0] w_n14363_0;
	wire [2:0] w_n14367_0;
	wire [2:0] w_n14369_0;
	wire [1:0] w_n14370_0;
	wire [2:0] w_n14374_0;
	wire [2:0] w_n14377_0;
	wire [1:0] w_n14378_0;
	wire [2:0] w_n14382_0;
	wire [2:0] w_n14384_0;
	wire [1:0] w_n14385_0;
	wire [2:0] w_n14389_0;
	wire [2:0] w_n14392_0;
	wire [1:0] w_n14393_0;
	wire [2:0] w_n14397_0;
	wire [2:0] w_n14399_0;
	wire [1:0] w_n14400_0;
	wire [2:0] w_n14404_0;
	wire [2:0] w_n14407_0;
	wire [1:0] w_n14408_0;
	wire [2:0] w_n14412_0;
	wire [2:0] w_n14415_0;
	wire [1:0] w_n14416_0;
	wire [1:0] w_n14420_0;
	wire [1:0] w_n14421_0;
	wire [2:0] w_n14423_0;
	wire [1:0] w_n14423_1;
	wire [2:0] w_n14426_0;
	wire [2:0] w_n14426_1;
	wire [1:0] w_n14427_0;
	wire [1:0] w_n14430_0;
	wire [1:0] w_n14432_0;
	wire [1:0] w_n14437_0;
	wire [1:0] w_n14438_0;
	wire [2:0] w_n14443_0;
	wire [1:0] w_n14443_1;
	wire [1:0] w_n14444_0;
	wire [2:0] w_n14445_0;
	wire [1:0] w_n14446_0;
	wire [2:0] w_n14448_0;
	wire [1:0] w_n14449_0;
	wire [1:0] w_n14454_0;
	wire [1:0] w_n14506_0;
	wire [1:0] w_n14594_0;
	wire [1:0] w_n14671_0;
	wire [1:0] w_n14672_0;
	wire [2:0] w_n14674_0;
	wire [2:0] w_n14674_1;
	wire [2:0] w_n14674_2;
	wire [2:0] w_n14674_3;
	wire [2:0] w_n14674_4;
	wire [2:0] w_n14674_5;
	wire [2:0] w_n14674_6;
	wire [2:0] w_n14674_7;
	wire [2:0] w_n14674_8;
	wire [2:0] w_n14674_9;
	wire [2:0] w_n14674_10;
	wire [2:0] w_n14674_11;
	wire [2:0] w_n14674_12;
	wire [2:0] w_n14674_13;
	wire [2:0] w_n14674_14;
	wire [2:0] w_n14674_15;
	wire [2:0] w_n14674_16;
	wire [2:0] w_n14674_17;
	wire [2:0] w_n14674_18;
	wire [2:0] w_n14674_19;
	wire [1:0] w_n14674_20;
	wire [2:0] w_n14678_0;
	wire [1:0] w_n14679_0;
	wire [1:0] w_n14681_0;
	wire [1:0] w_n14686_0;
	wire [1:0] w_n14687_0;
	wire [2:0] w_n14689_0;
	wire [1:0] w_n14690_0;
	wire [1:0] w_n14694_0;
	wire [2:0] w_n14696_0;
	wire [1:0] w_n14697_0;
	wire [1:0] w_n14701_0;
	wire [1:0] w_n14702_0;
	wire [2:0] w_n14704_0;
	wire [1:0] w_n14705_0;
	wire [1:0] w_n14709_0;
	wire [2:0] w_n14711_0;
	wire [1:0] w_n14712_0;
	wire [1:0] w_n14716_0;
	wire [1:0] w_n14717_0;
	wire [2:0] w_n14719_0;
	wire [1:0] w_n14720_0;
	wire [1:0] w_n14724_0;
	wire [1:0] w_n14725_0;
	wire [2:0] w_n14727_0;
	wire [1:0] w_n14728_0;
	wire [1:0] w_n14732_0;
	wire [1:0] w_n14733_0;
	wire [2:0] w_n14735_0;
	wire [1:0] w_n14736_0;
	wire [1:0] w_n14740_0;
	wire [2:0] w_n14742_0;
	wire [1:0] w_n14743_0;
	wire [1:0] w_n14747_0;
	wire [1:0] w_n14748_0;
	wire [2:0] w_n14750_0;
	wire [1:0] w_n14751_0;
	wire [1:0] w_n14755_0;
	wire [2:0] w_n14757_0;
	wire [1:0] w_n14758_0;
	wire [1:0] w_n14762_0;
	wire [1:0] w_n14763_0;
	wire [2:0] w_n14765_0;
	wire [1:0] w_n14766_0;
	wire [1:0] w_n14770_0;
	wire [2:0] w_n14772_0;
	wire [1:0] w_n14773_0;
	wire [1:0] w_n14777_0;
	wire [1:0] w_n14778_0;
	wire [2:0] w_n14780_0;
	wire [1:0] w_n14781_0;
	wire [1:0] w_n14785_0;
	wire [2:0] w_n14787_0;
	wire [1:0] w_n14788_0;
	wire [1:0] w_n14792_0;
	wire [1:0] w_n14793_0;
	wire [2:0] w_n14795_0;
	wire [1:0] w_n14796_0;
	wire [1:0] w_n14800_0;
	wire [1:0] w_n14801_0;
	wire [2:0] w_n14803_0;
	wire [1:0] w_n14804_0;
	wire [1:0] w_n14808_0;
	wire [1:0] w_n14809_0;
	wire [2:0] w_n14811_0;
	wire [1:0] w_n14812_0;
	wire [1:0] w_n14816_0;
	wire [2:0] w_n14818_0;
	wire [1:0] w_n14819_0;
	wire [1:0] w_n14823_0;
	wire [1:0] w_n14824_0;
	wire [2:0] w_n14826_0;
	wire [1:0] w_n14827_0;
	wire [1:0] w_n14831_0;
	wire [2:0] w_n14833_0;
	wire [1:0] w_n14834_0;
	wire [1:0] w_n14838_0;
	wire [1:0] w_n14839_0;
	wire [2:0] w_n14841_0;
	wire [1:0] w_n14842_0;
	wire [1:0] w_n14846_0;
	wire [1:0] w_n14847_0;
	wire [2:0] w_n14849_0;
	wire [1:0] w_n14850_0;
	wire [1:0] w_n14854_0;
	wire [1:0] w_n14855_0;
	wire [2:0] w_n14857_0;
	wire [1:0] w_n14858_0;
	wire [1:0] w_n14862_0;
	wire [2:0] w_n14864_0;
	wire [1:0] w_n14865_0;
	wire [1:0] w_n14869_0;
	wire [1:0] w_n14870_0;
	wire [2:0] w_n14872_0;
	wire [1:0] w_n14873_0;
	wire [1:0] w_n14877_0;
	wire [2:0] w_n14879_0;
	wire [1:0] w_n14880_0;
	wire [1:0] w_n14884_0;
	wire [1:0] w_n14885_0;
	wire [2:0] w_n14887_0;
	wire [1:0] w_n14888_0;
	wire [1:0] w_n14892_0;
	wire [1:0] w_n14893_0;
	wire [2:0] w_n14895_0;
	wire [1:0] w_n14896_0;
	wire [1:0] w_n14900_0;
	wire [2:0] w_n14902_0;
	wire [1:0] w_n14903_0;
	wire [1:0] w_n14906_0;
	wire [2:0] w_n14909_0;
	wire [1:0] w_n14910_0;
	wire [1:0] w_n14914_0;
	wire [1:0] w_n14915_0;
	wire [2:0] w_n14917_0;
	wire [1:0] w_n14918_0;
	wire [1:0] w_n14922_0;
	wire [2:0] w_n14924_0;
	wire [1:0] w_n14925_0;
	wire [1:0] w_n14929_0;
	wire [1:0] w_n14930_0;
	wire [2:0] w_n14932_0;
	wire [1:0] w_n14933_0;
	wire [1:0] w_n14937_0;
	wire [2:0] w_n14939_0;
	wire [1:0] w_n14940_0;
	wire [1:0] w_n14944_0;
	wire [1:0] w_n14945_0;
	wire [2:0] w_n14947_0;
	wire [1:0] w_n14948_0;
	wire [1:0] w_n14952_0;
	wire [1:0] w_n14953_0;
	wire [2:0] w_n14955_0;
	wire [1:0] w_n14956_0;
	wire [1:0] w_n14960_0;
	wire [1:0] w_n14961_0;
	wire [2:0] w_n14963_0;
	wire [1:0] w_n14964_0;
	wire [1:0] w_n14968_0;
	wire [2:0] w_n14970_0;
	wire [1:0] w_n14971_0;
	wire [1:0] w_n14975_0;
	wire [1:0] w_n14976_0;
	wire [2:0] w_n14978_0;
	wire [1:0] w_n14979_0;
	wire [1:0] w_n14983_0;
	wire [2:0] w_n14985_0;
	wire [1:0] w_n14986_0;
	wire [1:0] w_n14990_0;
	wire [1:0] w_n14991_0;
	wire [2:0] w_n14993_0;
	wire [1:0] w_n14994_0;
	wire [1:0] w_n14998_0;
	wire [2:0] w_n15000_0;
	wire [1:0] w_n15001_0;
	wire [1:0] w_n15005_0;
	wire [1:0] w_n15006_0;
	wire [2:0] w_n15008_0;
	wire [1:0] w_n15009_0;
	wire [1:0] w_n15013_0;
	wire [2:0] w_n15015_0;
	wire [1:0] w_n15016_0;
	wire [1:0] w_n15033_0;
	wire [1:0] w_n15070_0;
	wire [1:0] w_n15077_0;
	wire [1:0] w_n15084_0;
	wire [1:0] w_n15097_0;
	wire [1:0] w_n15104_0;
	wire [1:0] w_n15111_0;
	wire [1:0] w_n15118_0;
	wire [1:0] w_n15131_0;
	wire [1:0] w_n15138_0;
	wire [1:0] w_n15151_0;
	wire [1:0] w_n15158_0;
	wire [1:0] w_n15168_0;
	wire [1:0] w_n15178_0;
	wire [1:0] w_n15185_0;
	wire [1:0] w_n15198_0;
	wire [1:0] w_n15205_0;
	wire [1:0] w_n15212_0;
	wire [1:0] w_n15219_0;
	wire [1:0] w_n15225_0;
	wire [1:0] w_n15226_0;
	wire [2:0] w_n15228_0;
	wire [2:0] w_n15231_0;
	wire [1:0] w_n15231_1;
	wire [1:0] w_n15232_0;
	wire [1:0] w_n15233_0;
	wire [1:0] w_n15235_0;
	wire [1:0] w_n15237_0;
	wire [1:0] w_n15238_0;
	wire [2:0] w_n15239_0;
	wire [1:0] w_n15243_0;
	wire [1:0] w_n15244_0;
	wire [1:0] w_n15249_0;
	wire [1:0] w_n15250_0;
	wire [1:0] w_n15251_0;
	wire [2:0] w_n15256_0;
	wire [2:0] w_n15260_0;
	wire [2:0] w_n15260_1;
	wire [2:0] w_n15260_2;
	wire [2:0] w_n15260_3;
	wire [2:0] w_n15260_4;
	wire [2:0] w_n15260_5;
	wire [2:0] w_n15260_6;
	wire [2:0] w_n15260_7;
	wire [2:0] w_n15260_8;
	wire [2:0] w_n15260_9;
	wire [2:0] w_n15260_10;
	wire [2:0] w_n15260_11;
	wire [2:0] w_n15260_12;
	wire [2:0] w_n15260_13;
	wire [2:0] w_n15260_14;
	wire [2:0] w_n15260_15;
	wire [2:0] w_n15260_16;
	wire [2:0] w_n15260_17;
	wire [2:0] w_n15260_18;
	wire [2:0] w_n15260_19;
	wire [2:0] w_n15260_20;
	wire [2:0] w_n15260_21;
	wire [2:0] w_n15260_22;
	wire [2:0] w_n15260_23;
	wire [2:0] w_n15260_24;
	wire [2:0] w_n15260_25;
	wire [2:0] w_n15260_26;
	wire [2:0] w_n15260_27;
	wire [2:0] w_n15260_28;
	wire [2:0] w_n15260_29;
	wire [2:0] w_n15260_30;
	wire [2:0] w_n15260_31;
	wire [2:0] w_n15260_32;
	wire [2:0] w_n15260_33;
	wire [2:0] w_n15260_34;
	wire [2:0] w_n15260_35;
	wire [2:0] w_n15260_36;
	wire [2:0] w_n15260_37;
	wire [2:0] w_n15260_38;
	wire [2:0] w_n15260_39;
	wire [2:0] w_n15260_40;
	wire [2:0] w_n15260_41;
	wire [1:0] w_n15263_0;
	wire [2:0] w_n15264_0;
	wire [2:0] w_n15265_0;
	wire [2:0] w_n15265_1;
	wire [1:0] w_n15266_0;
	wire [2:0] w_n15267_0;
	wire [1:0] w_n15268_0;
	wire [2:0] w_n15271_0;
	wire [1:0] w_n15272_0;
	wire [2:0] w_n15279_0;
	wire [1:0] w_n15280_0;
	wire [1:0] w_n15283_0;
	wire [1:0] w_n15288_0;
	wire [2:0] w_n15290_0;
	wire [1:0] w_n15291_0;
	wire [2:0] w_n15295_0;
	wire [2:0] w_n15298_0;
	wire [1:0] w_n15299_0;
	wire [2:0] w_n15303_0;
	wire [2:0] w_n15305_0;
	wire [1:0] w_n15306_0;
	wire [2:0] w_n15310_0;
	wire [2:0] w_n15313_0;
	wire [1:0] w_n15314_0;
	wire [2:0] w_n15318_0;
	wire [2:0] w_n15320_0;
	wire [1:0] w_n15321_0;
	wire [2:0] w_n15325_0;
	wire [2:0] w_n15328_0;
	wire [1:0] w_n15329_0;
	wire [2:0] w_n15333_0;
	wire [2:0] w_n15335_0;
	wire [1:0] w_n15336_0;
	wire [2:0] w_n15340_0;
	wire [2:0] w_n15342_0;
	wire [1:0] w_n15343_0;
	wire [2:0] w_n15347_0;
	wire [2:0] w_n15349_0;
	wire [1:0] w_n15350_0;
	wire [2:0] w_n15354_0;
	wire [2:0] w_n15357_0;
	wire [1:0] w_n15358_0;
	wire [2:0] w_n15362_0;
	wire [2:0] w_n15364_0;
	wire [1:0] w_n15365_0;
	wire [2:0] w_n15369_0;
	wire [2:0] w_n15372_0;
	wire [1:0] w_n15373_0;
	wire [2:0] w_n15377_0;
	wire [2:0] w_n15379_0;
	wire [1:0] w_n15380_0;
	wire [2:0] w_n15384_0;
	wire [2:0] w_n15387_0;
	wire [1:0] w_n15388_0;
	wire [2:0] w_n15392_0;
	wire [2:0] w_n15394_0;
	wire [1:0] w_n15395_0;
	wire [2:0] w_n15399_0;
	wire [2:0] w_n15402_0;
	wire [1:0] w_n15403_0;
	wire [2:0] w_n15407_0;
	wire [2:0] w_n15409_0;
	wire [1:0] w_n15410_0;
	wire [2:0] w_n15414_0;
	wire [2:0] w_n15416_0;
	wire [1:0] w_n15417_0;
	wire [2:0] w_n15421_0;
	wire [2:0] w_n15423_0;
	wire [1:0] w_n15424_0;
	wire [2:0] w_n15428_0;
	wire [2:0] w_n15431_0;
	wire [1:0] w_n15432_0;
	wire [2:0] w_n15436_0;
	wire [2:0] w_n15438_0;
	wire [1:0] w_n15439_0;
	wire [2:0] w_n15443_0;
	wire [2:0] w_n15446_0;
	wire [1:0] w_n15447_0;
	wire [2:0] w_n15451_0;
	wire [2:0] w_n15453_0;
	wire [1:0] w_n15454_0;
	wire [2:0] w_n15458_0;
	wire [2:0] w_n15460_0;
	wire [1:0] w_n15461_0;
	wire [2:0] w_n15465_0;
	wire [2:0] w_n15467_0;
	wire [1:0] w_n15468_0;
	wire [2:0] w_n15472_0;
	wire [2:0] w_n15475_0;
	wire [1:0] w_n15476_0;
	wire [2:0] w_n15480_0;
	wire [2:0] w_n15482_0;
	wire [1:0] w_n15483_0;
	wire [2:0] w_n15487_0;
	wire [2:0] w_n15490_0;
	wire [1:0] w_n15491_0;
	wire [2:0] w_n15495_0;
	wire [2:0] w_n15497_0;
	wire [1:0] w_n15498_0;
	wire [2:0] w_n15502_0;
	wire [2:0] w_n15504_0;
	wire [1:0] w_n15505_0;
	wire [2:0] w_n15509_0;
	wire [2:0] w_n15512_0;
	wire [1:0] w_n15513_0;
	wire [2:0] w_n15516_0;
	wire [2:0] w_n15520_0;
	wire [1:0] w_n15521_0;
	wire [2:0] w_n15525_0;
	wire [2:0] w_n15527_0;
	wire [1:0] w_n15528_0;
	wire [2:0] w_n15532_0;
	wire [2:0] w_n15535_0;
	wire [1:0] w_n15536_0;
	wire [2:0] w_n15540_0;
	wire [2:0] w_n15542_0;
	wire [1:0] w_n15543_0;
	wire [2:0] w_n15547_0;
	wire [2:0] w_n15550_0;
	wire [1:0] w_n15551_0;
	wire [2:0] w_n15555_0;
	wire [2:0] w_n15557_0;
	wire [1:0] w_n15558_0;
	wire [2:0] w_n15562_0;
	wire [2:0] w_n15564_0;
	wire [1:0] w_n15565_0;
	wire [2:0] w_n15569_0;
	wire [2:0] w_n15571_0;
	wire [1:0] w_n15572_0;
	wire [2:0] w_n15576_0;
	wire [2:0] w_n15579_0;
	wire [1:0] w_n15580_0;
	wire [2:0] w_n15584_0;
	wire [2:0] w_n15586_0;
	wire [1:0] w_n15587_0;
	wire [2:0] w_n15591_0;
	wire [2:0] w_n15594_0;
	wire [1:0] w_n15595_0;
	wire [2:0] w_n15599_0;
	wire [2:0] w_n15601_0;
	wire [1:0] w_n15602_0;
	wire [2:0] w_n15606_0;
	wire [2:0] w_n15609_0;
	wire [1:0] w_n15610_0;
	wire [2:0] w_n15614_0;
	wire [2:0] w_n15616_0;
	wire [1:0] w_n15617_0;
	wire [1:0] w_n15621_0;
	wire [1:0] w_n15622_0;
	wire [2:0] w_n15624_0;
	wire [1:0] w_n15625_0;
	wire [1:0] w_n15626_0;
	wire [2:0] w_n15631_0;
	wire [1:0] w_n15636_0;
	wire [1:0] w_n15639_0;
	wire [2:0] w_n15642_0;
	wire [1:0] w_n15642_1;
	wire [1:0] w_n15643_0;
	wire [2:0] w_n15644_0;
	wire [1:0] w_n15645_0;
	wire [2:0] w_n15646_0;
	wire [1:0] w_n15647_0;
	wire [1:0] w_n15704_0;
	wire [1:0] w_n15708_0;
	wire [1:0] w_n15872_0;
	wire [1:0] w_n15876_0;
	wire [2:0] w_n15878_0;
	wire [2:0] w_n15878_1;
	wire [2:0] w_n15878_2;
	wire [2:0] w_n15878_3;
	wire [2:0] w_n15878_4;
	wire [2:0] w_n15878_5;
	wire [2:0] w_n15878_6;
	wire [2:0] w_n15878_7;
	wire [2:0] w_n15878_8;
	wire [2:0] w_n15878_9;
	wire [2:0] w_n15878_10;
	wire [2:0] w_n15878_11;
	wire [2:0] w_n15878_12;
	wire [2:0] w_n15878_13;
	wire [2:0] w_n15878_14;
	wire [2:0] w_n15878_15;
	wire [2:0] w_n15878_16;
	wire [2:0] w_n15878_17;
	wire [1:0] w_n15878_18;
	wire [2:0] w_n15882_0;
	wire [1:0] w_n15883_0;
	wire [1:0] w_n15885_0;
	wire [1:0] w_n15886_0;
	wire [1:0] w_n15891_0;
	wire [1:0] w_n15892_0;
	wire [2:0] w_n15894_0;
	wire [1:0] w_n15895_0;
	wire [2:0] w_n15899_0;
	wire [2:0] w_n15901_0;
	wire [1:0] w_n15902_0;
	wire [1:0] w_n15906_0;
	wire [2:0] w_n15908_0;
	wire [1:0] w_n15909_0;
	wire [1:0] w_n15913_0;
	wire [2:0] w_n15915_0;
	wire [1:0] w_n15916_0;
	wire [1:0] w_n15920_0;
	wire [1:0] w_n15921_0;
	wire [2:0] w_n15923_0;
	wire [1:0] w_n15924_0;
	wire [1:0] w_n15928_0;
	wire [2:0] w_n15930_0;
	wire [1:0] w_n15931_0;
	wire [1:0] w_n15935_0;
	wire [1:0] w_n15936_0;
	wire [2:0] w_n15938_0;
	wire [1:0] w_n15939_0;
	wire [1:0] w_n15943_0;
	wire [2:0] w_n15945_0;
	wire [1:0] w_n15946_0;
	wire [1:0] w_n15950_0;
	wire [1:0] w_n15951_0;
	wire [2:0] w_n15953_0;
	wire [1:0] w_n15954_0;
	wire [1:0] w_n15958_0;
	wire [1:0] w_n15959_0;
	wire [2:0] w_n15961_0;
	wire [1:0] w_n15962_0;
	wire [1:0] w_n15966_0;
	wire [1:0] w_n15967_0;
	wire [2:0] w_n15969_0;
	wire [1:0] w_n15970_0;
	wire [1:0] w_n15974_0;
	wire [2:0] w_n15976_0;
	wire [1:0] w_n15977_0;
	wire [1:0] w_n15981_0;
	wire [1:0] w_n15982_0;
	wire [2:0] w_n15984_0;
	wire [1:0] w_n15985_0;
	wire [1:0] w_n15989_0;
	wire [2:0] w_n15991_0;
	wire [1:0] w_n15992_0;
	wire [1:0] w_n15996_0;
	wire [1:0] w_n15997_0;
	wire [2:0] w_n15999_0;
	wire [1:0] w_n16000_0;
	wire [1:0] w_n16004_0;
	wire [2:0] w_n16006_0;
	wire [1:0] w_n16007_0;
	wire [1:0] w_n16011_0;
	wire [1:0] w_n16012_0;
	wire [2:0] w_n16014_0;
	wire [1:0] w_n16015_0;
	wire [1:0] w_n16019_0;
	wire [2:0] w_n16021_0;
	wire [1:0] w_n16022_0;
	wire [1:0] w_n16026_0;
	wire [1:0] w_n16027_0;
	wire [2:0] w_n16029_0;
	wire [1:0] w_n16030_0;
	wire [1:0] w_n16034_0;
	wire [1:0] w_n16035_0;
	wire [2:0] w_n16037_0;
	wire [1:0] w_n16038_0;
	wire [1:0] w_n16042_0;
	wire [1:0] w_n16043_0;
	wire [2:0] w_n16045_0;
	wire [1:0] w_n16046_0;
	wire [1:0] w_n16050_0;
	wire [2:0] w_n16052_0;
	wire [1:0] w_n16053_0;
	wire [1:0] w_n16057_0;
	wire [1:0] w_n16058_0;
	wire [2:0] w_n16060_0;
	wire [1:0] w_n16061_0;
	wire [1:0] w_n16065_0;
	wire [2:0] w_n16067_0;
	wire [1:0] w_n16068_0;
	wire [1:0] w_n16072_0;
	wire [1:0] w_n16073_0;
	wire [2:0] w_n16075_0;
	wire [1:0] w_n16076_0;
	wire [1:0] w_n16080_0;
	wire [1:0] w_n16081_0;
	wire [2:0] w_n16083_0;
	wire [1:0] w_n16084_0;
	wire [1:0] w_n16088_0;
	wire [1:0] w_n16089_0;
	wire [2:0] w_n16091_0;
	wire [1:0] w_n16092_0;
	wire [1:0] w_n16096_0;
	wire [2:0] w_n16098_0;
	wire [1:0] w_n16099_0;
	wire [1:0] w_n16103_0;
	wire [1:0] w_n16104_0;
	wire [2:0] w_n16106_0;
	wire [1:0] w_n16107_0;
	wire [1:0] w_n16111_0;
	wire [2:0] w_n16113_0;
	wire [1:0] w_n16114_0;
	wire [1:0] w_n16118_0;
	wire [1:0] w_n16119_0;
	wire [2:0] w_n16121_0;
	wire [1:0] w_n16122_0;
	wire [1:0] w_n16126_0;
	wire [1:0] w_n16127_0;
	wire [2:0] w_n16129_0;
	wire [1:0] w_n16130_0;
	wire [1:0] w_n16134_0;
	wire [2:0] w_n16136_0;
	wire [1:0] w_n16137_0;
	wire [1:0] w_n16140_0;
	wire [2:0] w_n16143_0;
	wire [1:0] w_n16144_0;
	wire [1:0] w_n16148_0;
	wire [1:0] w_n16149_0;
	wire [2:0] w_n16151_0;
	wire [1:0] w_n16152_0;
	wire [1:0] w_n16156_0;
	wire [2:0] w_n16158_0;
	wire [1:0] w_n16159_0;
	wire [1:0] w_n16163_0;
	wire [1:0] w_n16164_0;
	wire [2:0] w_n16166_0;
	wire [1:0] w_n16167_0;
	wire [1:0] w_n16171_0;
	wire [2:0] w_n16173_0;
	wire [1:0] w_n16174_0;
	wire [1:0] w_n16178_0;
	wire [1:0] w_n16179_0;
	wire [2:0] w_n16181_0;
	wire [1:0] w_n16182_0;
	wire [1:0] w_n16186_0;
	wire [1:0] w_n16187_0;
	wire [2:0] w_n16189_0;
	wire [1:0] w_n16190_0;
	wire [1:0] w_n16194_0;
	wire [1:0] w_n16195_0;
	wire [2:0] w_n16197_0;
	wire [1:0] w_n16198_0;
	wire [1:0] w_n16202_0;
	wire [2:0] w_n16204_0;
	wire [1:0] w_n16205_0;
	wire [1:0] w_n16209_0;
	wire [1:0] w_n16210_0;
	wire [2:0] w_n16212_0;
	wire [1:0] w_n16213_0;
	wire [1:0] w_n16217_0;
	wire [2:0] w_n16219_0;
	wire [1:0] w_n16220_0;
	wire [1:0] w_n16224_0;
	wire [1:0] w_n16225_0;
	wire [2:0] w_n16227_0;
	wire [1:0] w_n16228_0;
	wire [1:0] w_n16232_0;
	wire [2:0] w_n16234_0;
	wire [1:0] w_n16235_0;
	wire [1:0] w_n16250_0;
	wire [1:0] w_n16291_0;
	wire [1:0] w_n16302_0;
	wire [1:0] w_n16306_0;
	wire [1:0] w_n16313_0;
	wire [1:0] w_n16320_0;
	wire [1:0] w_n16333_0;
	wire [1:0] w_n16340_0;
	wire [1:0] w_n16347_0;
	wire [1:0] w_n16354_0;
	wire [1:0] w_n16367_0;
	wire [1:0] w_n16374_0;
	wire [1:0] w_n16387_0;
	wire [1:0] w_n16394_0;
	wire [1:0] w_n16404_0;
	wire [1:0] w_n16414_0;
	wire [1:0] w_n16421_0;
	wire [1:0] w_n16434_0;
	wire [1:0] w_n16441_0;
	wire [1:0] w_n16448_0;
	wire [2:0] w_n16454_0;
	wire [2:0] w_n16456_0;
	wire [2:0] w_n16459_0;
	wire [1:0] w_n16460_0;
	wire [1:0] w_n16462_0;
	wire [1:0] w_n16464_0;
	wire [1:0] w_n16465_0;
	wire [2:0] w_n16466_0;
	wire [1:0] w_n16471_0;
	wire [1:0] w_n16472_0;
	wire [1:0] w_n16478_0;
	wire [1:0] w_n16479_0;
	wire [1:0] w_n16480_0;
	wire [2:0] w_n16485_0;
	wire [2:0] w_n16489_0;
	wire [2:0] w_n16489_1;
	wire [2:0] w_n16489_2;
	wire [2:0] w_n16489_3;
	wire [2:0] w_n16489_4;
	wire [2:0] w_n16489_5;
	wire [2:0] w_n16489_6;
	wire [2:0] w_n16489_7;
	wire [2:0] w_n16489_8;
	wire [2:0] w_n16489_9;
	wire [2:0] w_n16489_10;
	wire [2:0] w_n16489_11;
	wire [2:0] w_n16489_12;
	wire [2:0] w_n16489_13;
	wire [2:0] w_n16489_14;
	wire [2:0] w_n16489_15;
	wire [2:0] w_n16489_16;
	wire [2:0] w_n16489_17;
	wire [2:0] w_n16489_18;
	wire [2:0] w_n16489_19;
	wire [2:0] w_n16489_20;
	wire [2:0] w_n16489_21;
	wire [2:0] w_n16489_22;
	wire [2:0] w_n16489_23;
	wire [2:0] w_n16489_24;
	wire [2:0] w_n16489_25;
	wire [2:0] w_n16489_26;
	wire [2:0] w_n16489_27;
	wire [2:0] w_n16489_28;
	wire [2:0] w_n16489_29;
	wire [2:0] w_n16489_30;
	wire [2:0] w_n16489_31;
	wire [2:0] w_n16489_32;
	wire [2:0] w_n16489_33;
	wire [2:0] w_n16489_34;
	wire [2:0] w_n16489_35;
	wire [2:0] w_n16489_36;
	wire [2:0] w_n16489_37;
	wire [2:0] w_n16489_38;
	wire [2:0] w_n16489_39;
	wire [1:0] w_n16492_0;
	wire [2:0] w_n16493_0;
	wire [2:0] w_n16494_0;
	wire [2:0] w_n16494_1;
	wire [1:0] w_n16495_0;
	wire [2:0] w_n16496_0;
	wire [1:0] w_n16497_0;
	wire [2:0] w_n16500_0;
	wire [1:0] w_n16501_0;
	wire [2:0] w_n16508_0;
	wire [1:0] w_n16509_0;
	wire [1:0] w_n16512_0;
	wire [2:0] w_n16517_0;
	wire [2:0] w_n16519_0;
	wire [1:0] w_n16520_0;
	wire [2:0] w_n16524_0;
	wire [2:0] w_n16527_0;
	wire [1:0] w_n16528_0;
	wire [2:0] w_n16532_0;
	wire [2:0] w_n16534_0;
	wire [1:0] w_n16535_0;
	wire [2:0] w_n16539_0;
	wire [2:0] w_n16541_0;
	wire [1:0] w_n16542_0;
	wire [2:0] w_n16546_0;
	wire [2:0] w_n16549_0;
	wire [1:0] w_n16550_0;
	wire [2:0] w_n16554_0;
	wire [2:0] w_n16557_0;
	wire [1:0] w_n16558_0;
	wire [2:0] w_n16562_0;
	wire [2:0] w_n16564_0;
	wire [1:0] w_n16565_0;
	wire [2:0] w_n16569_0;
	wire [2:0] w_n16572_0;
	wire [1:0] w_n16573_0;
	wire [2:0] w_n16577_0;
	wire [2:0] w_n16579_0;
	wire [1:0] w_n16580_0;
	wire [2:0] w_n16584_0;
	wire [2:0] w_n16587_0;
	wire [1:0] w_n16588_0;
	wire [2:0] w_n16592_0;
	wire [2:0] w_n16594_0;
	wire [1:0] w_n16595_0;
	wire [2:0] w_n16599_0;
	wire [2:0] w_n16601_0;
	wire [1:0] w_n16602_0;
	wire [2:0] w_n16606_0;
	wire [2:0] w_n16608_0;
	wire [1:0] w_n16609_0;
	wire [2:0] w_n16613_0;
	wire [2:0] w_n16616_0;
	wire [1:0] w_n16617_0;
	wire [2:0] w_n16621_0;
	wire [2:0] w_n16623_0;
	wire [1:0] w_n16624_0;
	wire [2:0] w_n16628_0;
	wire [2:0] w_n16631_0;
	wire [1:0] w_n16632_0;
	wire [2:0] w_n16636_0;
	wire [2:0] w_n16638_0;
	wire [1:0] w_n16639_0;
	wire [2:0] w_n16643_0;
	wire [2:0] w_n16646_0;
	wire [1:0] w_n16647_0;
	wire [2:0] w_n16651_0;
	wire [2:0] w_n16653_0;
	wire [1:0] w_n16654_0;
	wire [2:0] w_n16658_0;
	wire [2:0] w_n16661_0;
	wire [1:0] w_n16662_0;
	wire [2:0] w_n16666_0;
	wire [2:0] w_n16668_0;
	wire [1:0] w_n16669_0;
	wire [2:0] w_n16673_0;
	wire [2:0] w_n16675_0;
	wire [1:0] w_n16676_0;
	wire [2:0] w_n16680_0;
	wire [2:0] w_n16682_0;
	wire [1:0] w_n16683_0;
	wire [2:0] w_n16687_0;
	wire [2:0] w_n16690_0;
	wire [1:0] w_n16691_0;
	wire [2:0] w_n16695_0;
	wire [2:0] w_n16697_0;
	wire [1:0] w_n16698_0;
	wire [2:0] w_n16702_0;
	wire [2:0] w_n16705_0;
	wire [1:0] w_n16706_0;
	wire [2:0] w_n16710_0;
	wire [2:0] w_n16712_0;
	wire [1:0] w_n16713_0;
	wire [2:0] w_n16717_0;
	wire [2:0] w_n16719_0;
	wire [1:0] w_n16720_0;
	wire [2:0] w_n16724_0;
	wire [2:0] w_n16726_0;
	wire [1:0] w_n16727_0;
	wire [2:0] w_n16731_0;
	wire [2:0] w_n16734_0;
	wire [1:0] w_n16735_0;
	wire [2:0] w_n16739_0;
	wire [2:0] w_n16741_0;
	wire [1:0] w_n16742_0;
	wire [2:0] w_n16746_0;
	wire [2:0] w_n16749_0;
	wire [1:0] w_n16750_0;
	wire [2:0] w_n16754_0;
	wire [2:0] w_n16756_0;
	wire [1:0] w_n16757_0;
	wire [2:0] w_n16761_0;
	wire [2:0] w_n16763_0;
	wire [1:0] w_n16764_0;
	wire [2:0] w_n16768_0;
	wire [2:0] w_n16771_0;
	wire [1:0] w_n16772_0;
	wire [2:0] w_n16775_0;
	wire [2:0] w_n16779_0;
	wire [1:0] w_n16780_0;
	wire [2:0] w_n16784_0;
	wire [2:0] w_n16786_0;
	wire [1:0] w_n16787_0;
	wire [2:0] w_n16791_0;
	wire [2:0] w_n16794_0;
	wire [1:0] w_n16795_0;
	wire [2:0] w_n16799_0;
	wire [2:0] w_n16801_0;
	wire [1:0] w_n16802_0;
	wire [2:0] w_n16806_0;
	wire [2:0] w_n16809_0;
	wire [1:0] w_n16810_0;
	wire [2:0] w_n16814_0;
	wire [2:0] w_n16816_0;
	wire [1:0] w_n16817_0;
	wire [2:0] w_n16821_0;
	wire [2:0] w_n16823_0;
	wire [1:0] w_n16824_0;
	wire [2:0] w_n16828_0;
	wire [2:0] w_n16830_0;
	wire [1:0] w_n16831_0;
	wire [2:0] w_n16835_0;
	wire [2:0] w_n16838_0;
	wire [1:0] w_n16839_0;
	wire [2:0] w_n16843_0;
	wire [2:0] w_n16845_0;
	wire [1:0] w_n16846_0;
	wire [2:0] w_n16850_0;
	wire [2:0] w_n16853_0;
	wire [1:0] w_n16854_0;
	wire [2:0] w_n16858_0;
	wire [2:0] w_n16860_0;
	wire [1:0] w_n16861_0;
	wire [1:0] w_n16865_0;
	wire [1:0] w_n16866_0;
	wire [2:0] w_n16868_0;
	wire [2:0] w_n16869_0;
	wire [1:0] w_n16871_0;
	wire [1:0] w_n16872_0;
	wire [1:0] w_n16879_0;
	wire [1:0] w_n16880_0;
	wire [1:0] w_n16882_0;
	wire [2:0] w_n16885_0;
	wire [1:0] w_n16885_1;
	wire [1:0] w_n16886_0;
	wire [2:0] w_n16887_0;
	wire [1:0] w_n16888_0;
	wire [2:0] w_n16890_0;
	wire [1:0] w_n16891_0;
	wire [2:0] w_n16896_0;
	wire [1:0] w_n16896_1;
	wire [1:0] w_n16952_0;
	wire [1:0] w_n17127_0;
	wire [1:0] w_n17131_0;
	wire [1:0] w_n17132_0;
	wire [2:0] w_n17134_0;
	wire [2:0] w_n17134_1;
	wire [2:0] w_n17134_2;
	wire [2:0] w_n17134_3;
	wire [2:0] w_n17134_4;
	wire [2:0] w_n17134_5;
	wire [2:0] w_n17134_6;
	wire [2:0] w_n17134_7;
	wire [2:0] w_n17134_8;
	wire [2:0] w_n17134_9;
	wire [2:0] w_n17134_10;
	wire [2:0] w_n17134_11;
	wire [2:0] w_n17134_12;
	wire [2:0] w_n17134_13;
	wire [2:0] w_n17134_14;
	wire [1:0] w_n17134_15;
	wire [2:0] w_n17138_0;
	wire [1:0] w_n17139_0;
	wire [1:0] w_n17141_0;
	wire [1:0] w_n17146_0;
	wire [1:0] w_n17147_0;
	wire [2:0] w_n17149_0;
	wire [1:0] w_n17150_0;
	wire [1:0] w_n17154_0;
	wire [2:0] w_n17156_0;
	wire [1:0] w_n17157_0;
	wire [1:0] w_n17161_0;
	wire [1:0] w_n17162_0;
	wire [2:0] w_n17164_0;
	wire [1:0] w_n17165_0;
	wire [1:0] w_n17169_0;
	wire [2:0] w_n17171_0;
	wire [1:0] w_n17172_0;
	wire [1:0] w_n17176_0;
	wire [1:0] w_n17177_0;
	wire [2:0] w_n17179_0;
	wire [1:0] w_n17180_0;
	wire [1:0] w_n17184_0;
	wire [1:0] w_n17185_0;
	wire [2:0] w_n17187_0;
	wire [1:0] w_n17188_0;
	wire [1:0] w_n17192_0;
	wire [2:0] w_n17194_0;
	wire [1:0] w_n17195_0;
	wire [1:0] w_n17199_0;
	wire [2:0] w_n17201_0;
	wire [1:0] w_n17202_0;
	wire [1:0] w_n17206_0;
	wire [1:0] w_n17207_0;
	wire [2:0] w_n17209_0;
	wire [1:0] w_n17210_0;
	wire [1:0] w_n17214_0;
	wire [2:0] w_n17216_0;
	wire [1:0] w_n17217_0;
	wire [1:0] w_n17221_0;
	wire [1:0] w_n17222_0;
	wire [2:0] w_n17224_0;
	wire [1:0] w_n17225_0;
	wire [1:0] w_n17229_0;
	wire [2:0] w_n17231_0;
	wire [1:0] w_n17232_0;
	wire [1:0] w_n17236_0;
	wire [1:0] w_n17237_0;
	wire [2:0] w_n17239_0;
	wire [1:0] w_n17240_0;
	wire [1:0] w_n17244_0;
	wire [1:0] w_n17245_0;
	wire [2:0] w_n17247_0;
	wire [1:0] w_n17248_0;
	wire [1:0] w_n17252_0;
	wire [1:0] w_n17253_0;
	wire [2:0] w_n17255_0;
	wire [1:0] w_n17256_0;
	wire [1:0] w_n17260_0;
	wire [2:0] w_n17262_0;
	wire [1:0] w_n17263_0;
	wire [1:0] w_n17267_0;
	wire [1:0] w_n17268_0;
	wire [2:0] w_n17270_0;
	wire [1:0] w_n17271_0;
	wire [1:0] w_n17275_0;
	wire [2:0] w_n17277_0;
	wire [1:0] w_n17278_0;
	wire [1:0] w_n17282_0;
	wire [1:0] w_n17283_0;
	wire [2:0] w_n17285_0;
	wire [1:0] w_n17286_0;
	wire [1:0] w_n17290_0;
	wire [2:0] w_n17292_0;
	wire [1:0] w_n17293_0;
	wire [1:0] w_n17297_0;
	wire [1:0] w_n17298_0;
	wire [2:0] w_n17300_0;
	wire [1:0] w_n17301_0;
	wire [1:0] w_n17305_0;
	wire [2:0] w_n17307_0;
	wire [1:0] w_n17308_0;
	wire [1:0] w_n17312_0;
	wire [1:0] w_n17313_0;
	wire [2:0] w_n17315_0;
	wire [1:0] w_n17316_0;
	wire [1:0] w_n17320_0;
	wire [1:0] w_n17321_0;
	wire [2:0] w_n17323_0;
	wire [1:0] w_n17324_0;
	wire [1:0] w_n17328_0;
	wire [1:0] w_n17329_0;
	wire [2:0] w_n17331_0;
	wire [1:0] w_n17332_0;
	wire [1:0] w_n17336_0;
	wire [2:0] w_n17338_0;
	wire [1:0] w_n17339_0;
	wire [1:0] w_n17343_0;
	wire [1:0] w_n17344_0;
	wire [2:0] w_n17346_0;
	wire [1:0] w_n17347_0;
	wire [1:0] w_n17351_0;
	wire [2:0] w_n17353_0;
	wire [1:0] w_n17354_0;
	wire [1:0] w_n17358_0;
	wire [1:0] w_n17359_0;
	wire [2:0] w_n17361_0;
	wire [1:0] w_n17362_0;
	wire [1:0] w_n17366_0;
	wire [1:0] w_n17367_0;
	wire [2:0] w_n17369_0;
	wire [1:0] w_n17370_0;
	wire [1:0] w_n17374_0;
	wire [1:0] w_n17375_0;
	wire [2:0] w_n17377_0;
	wire [1:0] w_n17378_0;
	wire [1:0] w_n17382_0;
	wire [2:0] w_n17384_0;
	wire [1:0] w_n17385_0;
	wire [1:0] w_n17389_0;
	wire [1:0] w_n17390_0;
	wire [2:0] w_n17392_0;
	wire [1:0] w_n17393_0;
	wire [1:0] w_n17397_0;
	wire [2:0] w_n17399_0;
	wire [1:0] w_n17400_0;
	wire [1:0] w_n17404_0;
	wire [1:0] w_n17405_0;
	wire [2:0] w_n17407_0;
	wire [1:0] w_n17408_0;
	wire [1:0] w_n17412_0;
	wire [1:0] w_n17413_0;
	wire [2:0] w_n17415_0;
	wire [1:0] w_n17416_0;
	wire [1:0] w_n17420_0;
	wire [2:0] w_n17422_0;
	wire [1:0] w_n17423_0;
	wire [1:0] w_n17426_0;
	wire [2:0] w_n17429_0;
	wire [1:0] w_n17430_0;
	wire [1:0] w_n17434_0;
	wire [1:0] w_n17435_0;
	wire [2:0] w_n17437_0;
	wire [1:0] w_n17438_0;
	wire [1:0] w_n17442_0;
	wire [2:0] w_n17444_0;
	wire [1:0] w_n17445_0;
	wire [1:0] w_n17449_0;
	wire [1:0] w_n17450_0;
	wire [2:0] w_n17452_0;
	wire [1:0] w_n17453_0;
	wire [1:0] w_n17457_0;
	wire [2:0] w_n17459_0;
	wire [1:0] w_n17460_0;
	wire [1:0] w_n17464_0;
	wire [1:0] w_n17465_0;
	wire [2:0] w_n17467_0;
	wire [1:0] w_n17468_0;
	wire [1:0] w_n17472_0;
	wire [1:0] w_n17473_0;
	wire [2:0] w_n17475_0;
	wire [1:0] w_n17476_0;
	wire [1:0] w_n17480_0;
	wire [1:0] w_n17481_0;
	wire [2:0] w_n17483_0;
	wire [1:0] w_n17484_0;
	wire [1:0] w_n17488_0;
	wire [2:0] w_n17490_0;
	wire [1:0] w_n17491_0;
	wire [1:0] w_n17495_0;
	wire [1:0] w_n17496_0;
	wire [2:0] w_n17498_0;
	wire [1:0] w_n17499_0;
	wire [1:0] w_n17503_0;
	wire [2:0] w_n17505_0;
	wire [1:0] w_n17506_0;
	wire [2:0] w_n17510_0;
	wire [1:0] w_n17513_0;
	wire [2:0] w_n17516_0;
	wire [1:0] w_n17517_0;
	wire [2:0] w_n17518_0;
	wire [1:0] w_n17518_1;
	wire [2:0] w_n17519_0;
	wire [1:0] w_n17523_0;
	wire [1:0] w_n17524_0;
	wire [1:0] w_n17525_0;
	wire [1:0] w_n17538_0;
	wire [1:0] w_n17583_0;
	wire [1:0] w_n17590_0;
	wire [1:0] w_n17597_0;
	wire [1:0] w_n17607_0;
	wire [1:0] w_n17611_0;
	wire [1:0] w_n17618_0;
	wire [1:0] w_n17625_0;
	wire [1:0] w_n17638_0;
	wire [1:0] w_n17645_0;
	wire [1:0] w_n17652_0;
	wire [1:0] w_n17659_0;
	wire [1:0] w_n17672_0;
	wire [1:0] w_n17679_0;
	wire [1:0] w_n17692_0;
	wire [1:0] w_n17699_0;
	wire [1:0] w_n17709_0;
	wire [1:0] w_n17719_0;
	wire [1:0] w_n17726_0;
	wire [1:0] w_n17739_0;
	wire [1:0] w_n17746_0;
	wire [1:0] w_n17751_0;
	wire [1:0] w_n17752_0;
	wire [1:0] w_n17755_0;
	wire [1:0] w_n17756_0;
	wire [1:0] w_n17758_0;
	wire [1:0] w_n17762_0;
	wire [1:0] w_n17768_0;
	wire [2:0] w_n17769_0;
	wire [2:0] w_n17769_1;
	wire [2:0] w_n17769_2;
	wire [2:0] w_n17769_3;
	wire [2:0] w_n17769_4;
	wire [2:0] w_n17769_5;
	wire [2:0] w_n17769_6;
	wire [2:0] w_n17769_7;
	wire [2:0] w_n17769_8;
	wire [2:0] w_n17769_9;
	wire [2:0] w_n17769_10;
	wire [2:0] w_n17769_11;
	wire [2:0] w_n17769_12;
	wire [2:0] w_n17769_13;
	wire [2:0] w_n17769_14;
	wire [2:0] w_n17769_15;
	wire [2:0] w_n17769_16;
	wire [2:0] w_n17769_17;
	wire [2:0] w_n17769_18;
	wire [2:0] w_n17769_19;
	wire [2:0] w_n17769_20;
	wire [2:0] w_n17769_21;
	wire [2:0] w_n17769_22;
	wire [2:0] w_n17769_23;
	wire [2:0] w_n17769_24;
	wire [2:0] w_n17769_25;
	wire [2:0] w_n17769_26;
	wire [2:0] w_n17769_27;
	wire [2:0] w_n17769_28;
	wire [2:0] w_n17769_29;
	wire [2:0] w_n17769_30;
	wire [2:0] w_n17769_31;
	wire [2:0] w_n17769_32;
	wire [2:0] w_n17769_33;
	wire [2:0] w_n17769_34;
	wire [2:0] w_n17769_35;
	wire [2:0] w_n17769_36;
	wire [2:0] w_n17769_37;
	wire [1:0] w_n17769_38;
	wire [1:0] w_n17772_0;
	wire [2:0] w_n17773_0;
	wire [2:0] w_n17774_0;
	wire [2:0] w_n17774_1;
	wire [1:0] w_n17775_0;
	wire [2:0] w_n17776_0;
	wire [1:0] w_n17777_0;
	wire [2:0] w_n17780_0;
	wire [1:0] w_n17781_0;
	wire [2:0] w_n17788_0;
	wire [1:0] w_n17789_0;
	wire [1:0] w_n17792_0;
	wire [2:0] w_n17797_0;
	wire [2:0] w_n17799_0;
	wire [1:0] w_n17800_0;
	wire [2:0] w_n17804_0;
	wire [2:0] w_n17807_0;
	wire [1:0] w_n17808_0;
	wire [2:0] w_n17812_0;
	wire [2:0] w_n17814_0;
	wire [1:0] w_n17815_0;
	wire [2:0] w_n17819_0;
	wire [2:0] w_n17822_0;
	wire [1:0] w_n17823_0;
	wire [2:0] w_n17827_0;
	wire [2:0] w_n17829_0;
	wire [1:0] w_n17830_0;
	wire [2:0] w_n17834_0;
	wire [2:0] w_n17837_0;
	wire [1:0] w_n17838_0;
	wire [2:0] w_n17842_0;
	wire [2:0] w_n17844_0;
	wire [1:0] w_n17845_0;
	wire [2:0] w_n17849_0;
	wire [2:0] w_n17851_0;
	wire [1:0] w_n17852_0;
	wire [2:0] w_n17856_0;
	wire [2:0] w_n17859_0;
	wire [1:0] w_n17860_0;
	wire [2:0] w_n17864_0;
	wire [2:0] w_n17867_0;
	wire [1:0] w_n17868_0;
	wire [2:0] w_n17872_0;
	wire [2:0] w_n17874_0;
	wire [1:0] w_n17875_0;
	wire [2:0] w_n17879_0;
	wire [2:0] w_n17882_0;
	wire [1:0] w_n17883_0;
	wire [2:0] w_n17887_0;
	wire [2:0] w_n17889_0;
	wire [1:0] w_n17890_0;
	wire [2:0] w_n17894_0;
	wire [2:0] w_n17897_0;
	wire [1:0] w_n17898_0;
	wire [2:0] w_n17902_0;
	wire [2:0] w_n17904_0;
	wire [1:0] w_n17905_0;
	wire [2:0] w_n17909_0;
	wire [2:0] w_n17911_0;
	wire [1:0] w_n17912_0;
	wire [2:0] w_n17916_0;
	wire [2:0] w_n17918_0;
	wire [1:0] w_n17919_0;
	wire [2:0] w_n17923_0;
	wire [2:0] w_n17926_0;
	wire [1:0] w_n17927_0;
	wire [2:0] w_n17931_0;
	wire [2:0] w_n17933_0;
	wire [1:0] w_n17934_0;
	wire [2:0] w_n17938_0;
	wire [2:0] w_n17941_0;
	wire [1:0] w_n17942_0;
	wire [2:0] w_n17946_0;
	wire [2:0] w_n17948_0;
	wire [1:0] w_n17949_0;
	wire [2:0] w_n17953_0;
	wire [2:0] w_n17956_0;
	wire [1:0] w_n17957_0;
	wire [2:0] w_n17961_0;
	wire [2:0] w_n17963_0;
	wire [1:0] w_n17964_0;
	wire [2:0] w_n17968_0;
	wire [2:0] w_n17971_0;
	wire [1:0] w_n17972_0;
	wire [2:0] w_n17976_0;
	wire [2:0] w_n17978_0;
	wire [1:0] w_n17979_0;
	wire [2:0] w_n17983_0;
	wire [2:0] w_n17985_0;
	wire [1:0] w_n17986_0;
	wire [2:0] w_n17990_0;
	wire [2:0] w_n17992_0;
	wire [1:0] w_n17993_0;
	wire [2:0] w_n17997_0;
	wire [2:0] w_n18000_0;
	wire [1:0] w_n18001_0;
	wire [2:0] w_n18005_0;
	wire [2:0] w_n18007_0;
	wire [1:0] w_n18008_0;
	wire [1:0] w_n18012_0;
	wire [1:0] w_n18013_0;
	wire [2:0] w_n18015_0;
	wire [1:0] w_n18016_0;
	wire [2:0] w_n18020_0;
	wire [2:0] w_n18022_0;
	wire [1:0] w_n18023_0;
	wire [2:0] w_n18027_0;
	wire [2:0] w_n18029_0;
	wire [1:0] w_n18030_0;
	wire [2:0] w_n18034_0;
	wire [2:0] w_n18036_0;
	wire [1:0] w_n18037_0;
	wire [2:0] w_n18041_0;
	wire [2:0] w_n18044_0;
	wire [1:0] w_n18045_0;
	wire [2:0] w_n18049_0;
	wire [2:0] w_n18051_0;
	wire [1:0] w_n18052_0;
	wire [2:0] w_n18056_0;
	wire [2:0] w_n18059_0;
	wire [1:0] w_n18060_0;
	wire [2:0] w_n18064_0;
	wire [2:0] w_n18066_0;
	wire [1:0] w_n18067_0;
	wire [2:0] w_n18071_0;
	wire [2:0] w_n18073_0;
	wire [1:0] w_n18074_0;
	wire [2:0] w_n18078_0;
	wire [2:0] w_n18081_0;
	wire [1:0] w_n18082_0;
	wire [2:0] w_n18085_0;
	wire [2:0] w_n18089_0;
	wire [1:0] w_n18090_0;
	wire [2:0] w_n18094_0;
	wire [2:0] w_n18096_0;
	wire [1:0] w_n18097_0;
	wire [2:0] w_n18101_0;
	wire [2:0] w_n18104_0;
	wire [1:0] w_n18105_0;
	wire [2:0] w_n18109_0;
	wire [2:0] w_n18111_0;
	wire [1:0] w_n18112_0;
	wire [2:0] w_n18116_0;
	wire [2:0] w_n18119_0;
	wire [1:0] w_n18120_0;
	wire [2:0] w_n18124_0;
	wire [2:0] w_n18126_0;
	wire [1:0] w_n18127_0;
	wire [2:0] w_n18131_0;
	wire [2:0] w_n18133_0;
	wire [1:0] w_n18134_0;
	wire [2:0] w_n18138_0;
	wire [2:0] w_n18140_0;
	wire [1:0] w_n18141_0;
	wire [2:0] w_n18145_0;
	wire [2:0] w_n18148_0;
	wire [1:0] w_n18149_0;
	wire [2:0] w_n18153_0;
	wire [2:0] w_n18155_0;
	wire [1:0] w_n18156_0;
	wire [2:0] w_n18160_0;
	wire [2:0] w_n18163_0;
	wire [2:0] w_n18164_0;
	wire [1:0] w_n18168_0;
	wire [1:0] w_n18169_0;
	wire [1:0] w_n18171_0;
	wire [1:0] w_n18172_0;
	wire [1:0] w_n18176_0;
	wire [1:0] w_n18178_0;
	wire [2:0] w_n18182_0;
	wire [1:0] w_n18182_1;
	wire [1:0] w_n18183_0;
	wire [2:0] w_n18185_0;
	wire [1:0] w_n18185_1;
	wire [1:0] w_n18186_0;
	wire [2:0] w_n18187_0;
	wire [1:0] w_n18188_0;
	wire [2:0] w_n18189_0;
	wire [1:0] w_n18190_0;
	wire [2:0] w_n18195_0;
	wire [1:0] w_n18253_0;
	wire [1:0] w_n18435_0;
	wire [1:0] w_n18438_0;
	wire [1:0] w_n18441_0;
	wire [2:0] w_n18442_0;
	wire [2:0] w_n18442_1;
	wire [2:0] w_n18442_2;
	wire [2:0] w_n18442_3;
	wire [2:0] w_n18442_4;
	wire [2:0] w_n18442_5;
	wire [2:0] w_n18442_6;
	wire [2:0] w_n18442_7;
	wire [2:0] w_n18442_8;
	wire [2:0] w_n18442_9;
	wire [2:0] w_n18442_10;
	wire [2:0] w_n18442_11;
	wire [2:0] w_n18442_12;
	wire [2:0] w_n18446_0;
	wire [1:0] w_n18447_0;
	wire [1:0] w_n18449_0;
	wire [1:0] w_n18454_0;
	wire [1:0] w_n18455_0;
	wire [2:0] w_n18457_0;
	wire [1:0] w_n18458_0;
	wire [1:0] w_n18462_0;
	wire [2:0] w_n18464_0;
	wire [1:0] w_n18465_0;
	wire [1:0] w_n18469_0;
	wire [1:0] w_n18470_0;
	wire [2:0] w_n18472_0;
	wire [1:0] w_n18473_0;
	wire [1:0] w_n18477_0;
	wire [2:0] w_n18479_0;
	wire [1:0] w_n18480_0;
	wire [1:0] w_n18484_0;
	wire [1:0] w_n18485_0;
	wire [2:0] w_n18487_0;
	wire [1:0] w_n18488_0;
	wire [1:0] w_n18492_0;
	wire [2:0] w_n18494_0;
	wire [1:0] w_n18495_0;
	wire [1:0] w_n18499_0;
	wire [1:0] w_n18500_0;
	wire [2:0] w_n18502_0;
	wire [1:0] w_n18503_0;
	wire [1:0] w_n18507_0;
	wire [2:0] w_n18509_0;
	wire [1:0] w_n18510_0;
	wire [1:0] w_n18514_0;
	wire [1:0] w_n18515_0;
	wire [2:0] w_n18517_0;
	wire [1:0] w_n18518_0;
	wire [1:0] w_n18522_0;
	wire [1:0] w_n18523_0;
	wire [2:0] w_n18525_0;
	wire [1:0] w_n18526_0;
	wire [1:0] w_n18530_0;
	wire [2:0] w_n18532_0;
	wire [1:0] w_n18533_0;
	wire [1:0] w_n18537_0;
	wire [2:0] w_n18539_0;
	wire [1:0] w_n18540_0;
	wire [1:0] w_n18544_0;
	wire [1:0] w_n18545_0;
	wire [2:0] w_n18547_0;
	wire [1:0] w_n18548_0;
	wire [1:0] w_n18552_0;
	wire [2:0] w_n18554_0;
	wire [1:0] w_n18555_0;
	wire [1:0] w_n18559_0;
	wire [1:0] w_n18560_0;
	wire [2:0] w_n18562_0;
	wire [1:0] w_n18563_0;
	wire [1:0] w_n18567_0;
	wire [2:0] w_n18569_0;
	wire [1:0] w_n18570_0;
	wire [1:0] w_n18574_0;
	wire [1:0] w_n18575_0;
	wire [2:0] w_n18577_0;
	wire [1:0] w_n18578_0;
	wire [1:0] w_n18582_0;
	wire [1:0] w_n18583_0;
	wire [2:0] w_n18585_0;
	wire [1:0] w_n18586_0;
	wire [1:0] w_n18590_0;
	wire [1:0] w_n18591_0;
	wire [2:0] w_n18593_0;
	wire [1:0] w_n18594_0;
	wire [1:0] w_n18598_0;
	wire [2:0] w_n18600_0;
	wire [1:0] w_n18601_0;
	wire [1:0] w_n18605_0;
	wire [1:0] w_n18606_0;
	wire [2:0] w_n18608_0;
	wire [1:0] w_n18609_0;
	wire [1:0] w_n18613_0;
	wire [2:0] w_n18615_0;
	wire [1:0] w_n18616_0;
	wire [1:0] w_n18620_0;
	wire [1:0] w_n18621_0;
	wire [2:0] w_n18623_0;
	wire [1:0] w_n18624_0;
	wire [1:0] w_n18628_0;
	wire [2:0] w_n18630_0;
	wire [1:0] w_n18631_0;
	wire [1:0] w_n18635_0;
	wire [1:0] w_n18636_0;
	wire [2:0] w_n18638_0;
	wire [1:0] w_n18639_0;
	wire [1:0] w_n18643_0;
	wire [2:0] w_n18645_0;
	wire [1:0] w_n18646_0;
	wire [1:0] w_n18650_0;
	wire [1:0] w_n18651_0;
	wire [2:0] w_n18653_0;
	wire [1:0] w_n18654_0;
	wire [1:0] w_n18658_0;
	wire [1:0] w_n18659_0;
	wire [2:0] w_n18661_0;
	wire [1:0] w_n18662_0;
	wire [1:0] w_n18666_0;
	wire [1:0] w_n18667_0;
	wire [2:0] w_n18669_0;
	wire [1:0] w_n18670_0;
	wire [1:0] w_n18674_0;
	wire [2:0] w_n18676_0;
	wire [1:0] w_n18677_0;
	wire [1:0] w_n18681_0;
	wire [1:0] w_n18682_0;
	wire [2:0] w_n18684_0;
	wire [1:0] w_n18685_0;
	wire [1:0] w_n18689_0;
	wire [1:0] w_n18690_0;
	wire [2:0] w_n18692_0;
	wire [1:0] w_n18693_0;
	wire [1:0] w_n18697_0;
	wire [1:0] w_n18698_0;
	wire [2:0] w_n18700_0;
	wire [1:0] w_n18701_0;
	wire [1:0] w_n18705_0;
	wire [1:0] w_n18706_0;
	wire [2:0] w_n18708_0;
	wire [1:0] w_n18709_0;
	wire [1:0] w_n18713_0;
	wire [1:0] w_n18714_0;
	wire [2:0] w_n18716_0;
	wire [1:0] w_n18717_0;
	wire [1:0] w_n18721_0;
	wire [2:0] w_n18723_0;
	wire [1:0] w_n18724_0;
	wire [1:0] w_n18728_0;
	wire [1:0] w_n18729_0;
	wire [2:0] w_n18731_0;
	wire [1:0] w_n18732_0;
	wire [1:0] w_n18736_0;
	wire [2:0] w_n18738_0;
	wire [1:0] w_n18739_0;
	wire [1:0] w_n18743_0;
	wire [1:0] w_n18744_0;
	wire [2:0] w_n18746_0;
	wire [1:0] w_n18747_0;
	wire [1:0] w_n18751_0;
	wire [1:0] w_n18752_0;
	wire [2:0] w_n18754_0;
	wire [1:0] w_n18755_0;
	wire [1:0] w_n18759_0;
	wire [2:0] w_n18761_0;
	wire [1:0] w_n18762_0;
	wire [1:0] w_n18765_0;
	wire [2:0] w_n18768_0;
	wire [1:0] w_n18769_0;
	wire [1:0] w_n18773_0;
	wire [1:0] w_n18774_0;
	wire [2:0] w_n18776_0;
	wire [1:0] w_n18777_0;
	wire [1:0] w_n18781_0;
	wire [2:0] w_n18783_0;
	wire [1:0] w_n18784_0;
	wire [1:0] w_n18788_0;
	wire [1:0] w_n18789_0;
	wire [2:0] w_n18791_0;
	wire [1:0] w_n18792_0;
	wire [1:0] w_n18796_0;
	wire [2:0] w_n18798_0;
	wire [1:0] w_n18799_0;
	wire [2:0] w_n18803_0;
	wire [2:0] w_n18806_0;
	wire [1:0] w_n18807_0;
	wire [1:0] w_n18811_0;
	wire [1:0] w_n18812_0;
	wire [2:0] w_n18814_0;
	wire [1:0] w_n18815_0;
	wire [1:0] w_n18819_0;
	wire [1:0] w_n18820_0;
	wire [2:0] w_n18822_0;
	wire [1:0] w_n18823_0;
	wire [1:0] w_n18827_0;
	wire [2:0] w_n18829_0;
	wire [1:0] w_n18830_0;
	wire [1:0] w_n18841_0;
	wire [1:0] w_n18890_0;
	wire [1:0] w_n18897_0;
	wire [1:0] w_n18904_0;
	wire [1:0] w_n18911_0;
	wire [1:0] w_n18918_0;
	wire [1:0] w_n18928_0;
	wire [1:0] w_n18932_0;
	wire [1:0] w_n18939_0;
	wire [1:0] w_n18946_0;
	wire [1:0] w_n18959_0;
	wire [1:0] w_n18966_0;
	wire [1:0] w_n18973_0;
	wire [1:0] w_n18980_0;
	wire [1:0] w_n18993_0;
	wire [1:0] w_n19012_0;
	wire [1:0] w_n19019_0;
	wire [1:0] w_n19029_0;
	wire [1:0] w_n19039_0;
	wire [1:0] w_n19046_0;
	wire [1:0] w_n19059_0;
	wire [2:0] w_n19065_0;
	wire [1:0] w_n19067_0;
	wire [1:0] w_n19068_0;
	wire [1:0] w_n19070_0;
	wire [1:0] w_n19072_0;
	wire [1:0] w_n19073_0;
	wire [2:0] w_n19074_0;
	wire [1:0] w_n19079_0;
	wire [1:0] w_n19080_0;
	wire [2:0] w_n19086_0;
	wire [1:0] w_n19087_0;
	wire [2:0] w_n19096_0;
	wire [2:0] w_n19096_1;
	wire [2:0] w_n19096_2;
	wire [2:0] w_n19096_3;
	wire [2:0] w_n19096_4;
	wire [2:0] w_n19096_5;
	wire [2:0] w_n19096_6;
	wire [2:0] w_n19096_7;
	wire [2:0] w_n19096_8;
	wire [2:0] w_n19096_9;
	wire [2:0] w_n19096_10;
	wire [2:0] w_n19096_11;
	wire [2:0] w_n19096_12;
	wire [2:0] w_n19096_13;
	wire [2:0] w_n19096_14;
	wire [2:0] w_n19096_15;
	wire [2:0] w_n19096_16;
	wire [2:0] w_n19096_17;
	wire [2:0] w_n19096_18;
	wire [2:0] w_n19096_19;
	wire [2:0] w_n19096_20;
	wire [2:0] w_n19096_21;
	wire [2:0] w_n19096_22;
	wire [2:0] w_n19096_23;
	wire [2:0] w_n19096_24;
	wire [2:0] w_n19096_25;
	wire [2:0] w_n19096_26;
	wire [2:0] w_n19096_27;
	wire [2:0] w_n19096_28;
	wire [2:0] w_n19096_29;
	wire [2:0] w_n19096_30;
	wire [2:0] w_n19096_31;
	wire [2:0] w_n19096_32;
	wire [2:0] w_n19096_33;
	wire [2:0] w_n19096_34;
	wire [2:0] w_n19096_35;
	wire [1:0] w_n19096_36;
	wire [2:0] w_n19099_0;
	wire [2:0] w_n19100_0;
	wire [2:0] w_n19101_0;
	wire [2:0] w_n19101_1;
	wire [1:0] w_n19102_0;
	wire [2:0] w_n19103_0;
	wire [1:0] w_n19104_0;
	wire [2:0] w_n19107_0;
	wire [1:0] w_n19108_0;
	wire [1:0] w_n19113_0;
	wire [2:0] w_n19115_0;
	wire [1:0] w_n19116_0;
	wire [1:0] w_n19119_0;
	wire [2:0] w_n19124_0;
	wire [2:0] w_n19126_0;
	wire [1:0] w_n19127_0;
	wire [2:0] w_n19131_0;
	wire [2:0] w_n19134_0;
	wire [1:0] w_n19135_0;
	wire [2:0] w_n19139_0;
	wire [2:0] w_n19141_0;
	wire [1:0] w_n19142_0;
	wire [2:0] w_n19146_0;
	wire [2:0] w_n19149_0;
	wire [1:0] w_n19150_0;
	wire [2:0] w_n19154_0;
	wire [2:0] w_n19156_0;
	wire [1:0] w_n19157_0;
	wire [2:0] w_n19161_0;
	wire [2:0] w_n19164_0;
	wire [1:0] w_n19165_0;
	wire [2:0] w_n19169_0;
	wire [2:0] w_n19171_0;
	wire [1:0] w_n19172_0;
	wire [2:0] w_n19176_0;
	wire [2:0] w_n19179_0;
	wire [1:0] w_n19180_0;
	wire [2:0] w_n19184_0;
	wire [2:0] w_n19186_0;
	wire [1:0] w_n19187_0;
	wire [2:0] w_n19191_0;
	wire [2:0] w_n19194_0;
	wire [1:0] w_n19195_0;
	wire [2:0] w_n19199_0;
	wire [2:0] w_n19201_0;
	wire [1:0] w_n19202_0;
	wire [2:0] w_n19206_0;
	wire [2:0] w_n19208_0;
	wire [1:0] w_n19209_0;
	wire [2:0] w_n19213_0;
	wire [2:0] w_n19216_0;
	wire [1:0] w_n19217_0;
	wire [2:0] w_n19221_0;
	wire [2:0] w_n19224_0;
	wire [1:0] w_n19225_0;
	wire [2:0] w_n19229_0;
	wire [2:0] w_n19231_0;
	wire [1:0] w_n19232_0;
	wire [2:0] w_n19236_0;
	wire [2:0] w_n19239_0;
	wire [1:0] w_n19240_0;
	wire [2:0] w_n19244_0;
	wire [2:0] w_n19246_0;
	wire [1:0] w_n19247_0;
	wire [2:0] w_n19251_0;
	wire [2:0] w_n19254_0;
	wire [1:0] w_n19255_0;
	wire [2:0] w_n19259_0;
	wire [2:0] w_n19261_0;
	wire [1:0] w_n19262_0;
	wire [2:0] w_n19266_0;
	wire [2:0] w_n19268_0;
	wire [1:0] w_n19269_0;
	wire [2:0] w_n19273_0;
	wire [2:0] w_n19275_0;
	wire [1:0] w_n19276_0;
	wire [2:0] w_n19280_0;
	wire [2:0] w_n19283_0;
	wire [1:0] w_n19284_0;
	wire [2:0] w_n19288_0;
	wire [2:0] w_n19290_0;
	wire [1:0] w_n19291_0;
	wire [2:0] w_n19295_0;
	wire [2:0] w_n19298_0;
	wire [1:0] w_n19299_0;
	wire [2:0] w_n19303_0;
	wire [2:0] w_n19305_0;
	wire [1:0] w_n19306_0;
	wire [2:0] w_n19310_0;
	wire [2:0] w_n19313_0;
	wire [1:0] w_n19314_0;
	wire [2:0] w_n19318_0;
	wire [2:0] w_n19320_0;
	wire [1:0] w_n19321_0;
	wire [2:0] w_n19325_0;
	wire [2:0] w_n19328_0;
	wire [1:0] w_n19329_0;
	wire [2:0] w_n19333_0;
	wire [2:0] w_n19335_0;
	wire [1:0] w_n19336_0;
	wire [2:0] w_n19340_0;
	wire [2:0] w_n19342_0;
	wire [1:0] w_n19343_0;
	wire [2:0] w_n19347_0;
	wire [2:0] w_n19349_0;
	wire [1:0] w_n19350_0;
	wire [2:0] w_n19354_0;
	wire [2:0] w_n19357_0;
	wire [1:0] w_n19358_0;
	wire [2:0] w_n19362_0;
	wire [2:0] w_n19364_0;
	wire [1:0] w_n19365_0;
	wire [2:0] w_n19369_0;
	wire [2:0] w_n19371_0;
	wire [1:0] w_n19372_0;
	wire [2:0] w_n19376_0;
	wire [2:0] w_n19378_0;
	wire [1:0] w_n19379_0;
	wire [2:0] w_n19383_0;
	wire [2:0] w_n19385_0;
	wire [1:0] w_n19386_0;
	wire [2:0] w_n19390_0;
	wire [2:0] w_n19392_0;
	wire [1:0] w_n19393_0;
	wire [2:0] w_n19397_0;
	wire [2:0] w_n19400_0;
	wire [1:0] w_n19401_0;
	wire [2:0] w_n19405_0;
	wire [2:0] w_n19407_0;
	wire [1:0] w_n19408_0;
	wire [2:0] w_n19412_0;
	wire [2:0] w_n19415_0;
	wire [1:0] w_n19416_0;
	wire [2:0] w_n19420_0;
	wire [2:0] w_n19422_0;
	wire [1:0] w_n19423_0;
	wire [2:0] w_n19427_0;
	wire [2:0] w_n19429_0;
	wire [1:0] w_n19430_0;
	wire [2:0] w_n19434_0;
	wire [2:0] w_n19437_0;
	wire [1:0] w_n19438_0;
	wire [2:0] w_n19441_0;
	wire [2:0] w_n19445_0;
	wire [1:0] w_n19446_0;
	wire [2:0] w_n19450_0;
	wire [2:0] w_n19452_0;
	wire [1:0] w_n19453_0;
	wire [2:0] w_n19457_0;
	wire [2:0] w_n19460_0;
	wire [1:0] w_n19461_0;
	wire [2:0] w_n19465_0;
	wire [2:0] w_n19467_0;
	wire [1:0] w_n19468_0;
	wire [1:0] w_n19472_0;
	wire [1:0] w_n19473_0;
	wire [2:0] w_n19475_0;
	wire [1:0] w_n19476_0;
	wire [2:0] w_n19480_0;
	wire [2:0] w_n19483_0;
	wire [1:0] w_n19484_0;
	wire [2:0] w_n19488_0;
	wire [2:0] w_n19490_0;
	wire [1:0] w_n19491_0;
	wire [2:0] w_n19495_0;
	wire [2:0] w_n19497_0;
	wire [1:0] w_n19498_0;
	wire [2:0] w_n19502_0;
	wire [2:0] w_n19505_0;
	wire [1:0] w_n19506_0;
	wire [1:0] w_n19508_0;
	wire [1:0] w_n19511_0;
	wire [1:0] w_n19515_0;
	wire [2:0] w_n19522_0;
	wire [2:0] w_n19523_0;
	wire [2:0] w_n19524_0;
	wire [1:0] w_n19524_1;
	wire [1:0] w_n19525_0;
	wire [2:0] w_n19526_0;
	wire [1:0] w_n19527_0;
	wire [2:0] w_n19529_0;
	wire [1:0] w_n19530_0;
	wire [1:0] w_n19781_0;
	wire [1:0] w_n19782_0;
	wire [1:0] w_n19785_0;
	wire [1:0] w_n19786_0;
	wire [1:0] w_n19788_0;
	wire [2:0] w_n19791_0;
	wire [2:0] w_n19791_1;
	wire [2:0] w_n19791_2;
	wire [2:0] w_n19791_3;
	wire [2:0] w_n19791_4;
	wire [2:0] w_n19791_5;
	wire [2:0] w_n19791_6;
	wire [2:0] w_n19791_7;
	wire [2:0] w_n19791_8;
	wire [2:0] w_n19791_9;
	wire [2:0] w_n19791_10;
	wire [2:0] w_n19795_0;
	wire [1:0] w_n19796_0;
	wire [1:0] w_n19798_0;
	wire [1:0] w_n19802_0;
	wire [1:0] w_n19803_0;
	wire [2:0] w_n19805_0;
	wire [1:0] w_n19806_0;
	wire [1:0] w_n19810_0;
	wire [1:0] w_n19811_0;
	wire [2:0] w_n19813_0;
	wire [1:0] w_n19814_0;
	wire [1:0] w_n19818_0;
	wire [1:0] w_n19819_0;
	wire [2:0] w_n19821_0;
	wire [1:0] w_n19822_0;
	wire [1:0] w_n19826_0;
	wire [2:0] w_n19828_0;
	wire [1:0] w_n19829_0;
	wire [1:0] w_n19833_0;
	wire [1:0] w_n19834_0;
	wire [2:0] w_n19836_0;
	wire [1:0] w_n19837_0;
	wire [1:0] w_n19841_0;
	wire [2:0] w_n19843_0;
	wire [1:0] w_n19844_0;
	wire [1:0] w_n19848_0;
	wire [1:0] w_n19849_0;
	wire [2:0] w_n19851_0;
	wire [1:0] w_n19852_0;
	wire [1:0] w_n19856_0;
	wire [2:0] w_n19858_0;
	wire [1:0] w_n19859_0;
	wire [1:0] w_n19863_0;
	wire [1:0] w_n19864_0;
	wire [2:0] w_n19866_0;
	wire [1:0] w_n19867_0;
	wire [1:0] w_n19871_0;
	wire [2:0] w_n19873_0;
	wire [1:0] w_n19874_0;
	wire [1:0] w_n19878_0;
	wire [1:0] w_n19879_0;
	wire [2:0] w_n19881_0;
	wire [1:0] w_n19882_0;
	wire [1:0] w_n19886_0;
	wire [2:0] w_n19888_0;
	wire [1:0] w_n19889_0;
	wire [1:0] w_n19893_0;
	wire [1:0] w_n19894_0;
	wire [2:0] w_n19896_0;
	wire [1:0] w_n19897_0;
	wire [1:0] w_n19901_0;
	wire [1:0] w_n19902_0;
	wire [2:0] w_n19904_0;
	wire [1:0] w_n19905_0;
	wire [1:0] w_n19909_0;
	wire [2:0] w_n19911_0;
	wire [1:0] w_n19912_0;
	wire [1:0] w_n19916_0;
	wire [2:0] w_n19918_0;
	wire [1:0] w_n19919_0;
	wire [1:0] w_n19923_0;
	wire [1:0] w_n19924_0;
	wire [2:0] w_n19926_0;
	wire [1:0] w_n19927_0;
	wire [1:0] w_n19931_0;
	wire [2:0] w_n19933_0;
	wire [1:0] w_n19934_0;
	wire [1:0] w_n19938_0;
	wire [1:0] w_n19939_0;
	wire [2:0] w_n19941_0;
	wire [1:0] w_n19942_0;
	wire [1:0] w_n19946_0;
	wire [2:0] w_n19948_0;
	wire [1:0] w_n19949_0;
	wire [1:0] w_n19953_0;
	wire [1:0] w_n19954_0;
	wire [2:0] w_n19956_0;
	wire [1:0] w_n19957_0;
	wire [1:0] w_n19961_0;
	wire [1:0] w_n19962_0;
	wire [2:0] w_n19964_0;
	wire [1:0] w_n19965_0;
	wire [1:0] w_n19969_0;
	wire [1:0] w_n19970_0;
	wire [2:0] w_n19972_0;
	wire [1:0] w_n19973_0;
	wire [1:0] w_n19977_0;
	wire [2:0] w_n19979_0;
	wire [1:0] w_n19980_0;
	wire [1:0] w_n19984_0;
	wire [1:0] w_n19985_0;
	wire [2:0] w_n19987_0;
	wire [1:0] w_n19988_0;
	wire [1:0] w_n19992_0;
	wire [2:0] w_n19994_0;
	wire [1:0] w_n19995_0;
	wire [1:0] w_n19999_0;
	wire [1:0] w_n20000_0;
	wire [2:0] w_n20002_0;
	wire [1:0] w_n20003_0;
	wire [1:0] w_n20007_0;
	wire [2:0] w_n20009_0;
	wire [1:0] w_n20010_0;
	wire [1:0] w_n20014_0;
	wire [1:0] w_n20015_0;
	wire [2:0] w_n20017_0;
	wire [1:0] w_n20018_0;
	wire [1:0] w_n20022_0;
	wire [2:0] w_n20024_0;
	wire [1:0] w_n20025_0;
	wire [1:0] w_n20029_0;
	wire [1:0] w_n20030_0;
	wire [2:0] w_n20032_0;
	wire [1:0] w_n20033_0;
	wire [1:0] w_n20037_0;
	wire [1:0] w_n20038_0;
	wire [2:0] w_n20040_0;
	wire [1:0] w_n20041_0;
	wire [1:0] w_n20045_0;
	wire [1:0] w_n20046_0;
	wire [2:0] w_n20048_0;
	wire [1:0] w_n20049_0;
	wire [1:0] w_n20053_0;
	wire [2:0] w_n20055_0;
	wire [1:0] w_n20056_0;
	wire [1:0] w_n20060_0;
	wire [1:0] w_n20061_0;
	wire [2:0] w_n20063_0;
	wire [1:0] w_n20064_0;
	wire [1:0] w_n20068_0;
	wire [1:0] w_n20069_0;
	wire [2:0] w_n20071_0;
	wire [1:0] w_n20072_0;
	wire [1:0] w_n20076_0;
	wire [1:0] w_n20077_0;
	wire [2:0] w_n20079_0;
	wire [1:0] w_n20080_0;
	wire [1:0] w_n20084_0;
	wire [1:0] w_n20085_0;
	wire [2:0] w_n20087_0;
	wire [1:0] w_n20088_0;
	wire [1:0] w_n20092_0;
	wire [1:0] w_n20093_0;
	wire [2:0] w_n20095_0;
	wire [1:0] w_n20096_0;
	wire [1:0] w_n20100_0;
	wire [2:0] w_n20102_0;
	wire [1:0] w_n20103_0;
	wire [1:0] w_n20107_0;
	wire [1:0] w_n20108_0;
	wire [2:0] w_n20110_0;
	wire [1:0] w_n20111_0;
	wire [1:0] w_n20115_0;
	wire [2:0] w_n20117_0;
	wire [1:0] w_n20118_0;
	wire [1:0] w_n20122_0;
	wire [1:0] w_n20123_0;
	wire [2:0] w_n20125_0;
	wire [1:0] w_n20126_0;
	wire [1:0] w_n20130_0;
	wire [1:0] w_n20131_0;
	wire [2:0] w_n20133_0;
	wire [1:0] w_n20134_0;
	wire [1:0] w_n20138_0;
	wire [2:0] w_n20140_0;
	wire [1:0] w_n20141_0;
	wire [1:0] w_n20144_0;
	wire [2:0] w_n20147_0;
	wire [1:0] w_n20148_0;
	wire [1:0] w_n20152_0;
	wire [1:0] w_n20153_0;
	wire [2:0] w_n20155_0;
	wire [1:0] w_n20156_0;
	wire [1:0] w_n20160_0;
	wire [2:0] w_n20162_0;
	wire [1:0] w_n20163_0;
	wire [1:0] w_n20167_0;
	wire [1:0] w_n20168_0;
	wire [2:0] w_n20170_0;
	wire [1:0] w_n20171_0;
	wire [1:0] w_n20175_0;
	wire [1:0] w_n20176_0;
	wire [2:0] w_n20178_0;
	wire [1:0] w_n20179_0;
	wire [1:0] w_n20183_0;
	wire [2:0] w_n20185_0;
	wire [1:0] w_n20186_0;
	wire [1:0] w_n20190_0;
	wire [1:0] w_n20191_0;
	wire [2:0] w_n20193_0;
	wire [1:0] w_n20194_0;
	wire [1:0] w_n20203_0;
	wire [1:0] w_n20256_0;
	wire [1:0] w_n20269_0;
	wire [1:0] w_n20276_0;
	wire [1:0] w_n20283_0;
	wire [1:0] w_n20290_0;
	wire [1:0] w_n20297_0;
	wire [1:0] w_n20307_0;
	wire [1:0] w_n20311_0;
	wire [1:0] w_n20318_0;
	wire [1:0] w_n20325_0;
	wire [1:0] w_n20338_0;
	wire [1:0] w_n20345_0;
	wire [1:0] w_n20352_0;
	wire [1:0] w_n20359_0;
	wire [1:0] w_n20372_0;
	wire [1:0] w_n20391_0;
	wire [1:0] w_n20398_0;
	wire [1:0] w_n20408_0;
	wire [1:0] w_n20418_0;
	wire [1:0] w_n20428_0;
	wire [2:0] w_n20437_0;
	wire [2:0] w_n20439_0;
	wire [1:0] w_n20440_0;
	wire [1:0] w_n20442_0;
	wire [1:0] w_n20444_0;
	wire [1:0] w_n20445_0;
	wire [2:0] w_n20446_0;
	wire [1:0] w_n20451_0;
	wire [1:0] w_n20452_0;
	wire [1:0] w_n20458_0;
	wire [1:0] w_n20459_0;
	wire [1:0] w_n20464_0;
	wire [2:0] w_n20468_0;
	wire [2:0] w_n20468_1;
	wire [2:0] w_n20468_2;
	wire [2:0] w_n20468_3;
	wire [2:0] w_n20468_4;
	wire [2:0] w_n20468_5;
	wire [2:0] w_n20468_6;
	wire [2:0] w_n20468_7;
	wire [2:0] w_n20468_8;
	wire [2:0] w_n20468_9;
	wire [2:0] w_n20468_10;
	wire [2:0] w_n20468_11;
	wire [2:0] w_n20468_12;
	wire [2:0] w_n20468_13;
	wire [2:0] w_n20468_14;
	wire [2:0] w_n20468_15;
	wire [2:0] w_n20468_16;
	wire [2:0] w_n20468_17;
	wire [2:0] w_n20468_18;
	wire [2:0] w_n20468_19;
	wire [2:0] w_n20468_20;
	wire [2:0] w_n20468_21;
	wire [2:0] w_n20468_22;
	wire [2:0] w_n20468_23;
	wire [2:0] w_n20468_24;
	wire [2:0] w_n20468_25;
	wire [2:0] w_n20468_26;
	wire [2:0] w_n20468_27;
	wire [2:0] w_n20468_28;
	wire [2:0] w_n20468_29;
	wire [2:0] w_n20468_30;
	wire [2:0] w_n20468_31;
	wire [2:0] w_n20468_32;
	wire [2:0] w_n20468_33;
	wire [2:0] w_n20468_34;
	wire [2:0] w_n20468_35;
	wire [2:0] w_n20471_0;
	wire [1:0] w_n20472_0;
	wire [2:0] w_n20473_0;
	wire [2:0] w_n20473_1;
	wire [1:0] w_n20474_0;
	wire [2:0] w_n20475_0;
	wire [1:0] w_n20476_0;
	wire [2:0] w_n20479_0;
	wire [1:0] w_n20480_0;
	wire [2:0] w_n20487_0;
	wire [1:0] w_n20488_0;
	wire [1:0] w_n20491_0;
	wire [2:0] w_n20496_0;
	wire [2:0] w_n20498_0;
	wire [1:0] w_n20499_0;
	wire [2:0] w_n20503_0;
	wire [2:0] w_n20506_0;
	wire [1:0] w_n20507_0;
	wire [2:0] w_n20511_0;
	wire [2:0] w_n20513_0;
	wire [1:0] w_n20514_0;
	wire [2:0] w_n20518_0;
	wire [2:0] w_n20520_0;
	wire [1:0] w_n20521_0;
	wire [2:0] w_n20525_0;
	wire [2:0] w_n20527_0;
	wire [1:0] w_n20528_0;
	wire [2:0] w_n20532_0;
	wire [2:0] w_n20535_0;
	wire [1:0] w_n20536_0;
	wire [2:0] w_n20540_0;
	wire [2:0] w_n20542_0;
	wire [1:0] w_n20543_0;
	wire [1:0] w_n20547_0;
	wire [1:0] w_n20548_0;
	wire [2:0] w_n20550_0;
	wire [1:0] w_n20551_0;
	wire [2:0] w_n20555_0;
	wire [2:0] w_n20557_0;
	wire [1:0] w_n20558_0;
	wire [2:0] w_n20562_0;
	wire [2:0] w_n20565_0;
	wire [1:0] w_n20566_0;
	wire [2:0] w_n20570_0;
	wire [2:0] w_n20572_0;
	wire [1:0] w_n20573_0;
	wire [2:0] w_n20577_0;
	wire [2:0] w_n20580_0;
	wire [1:0] w_n20581_0;
	wire [2:0] w_n20585_0;
	wire [2:0] w_n20587_0;
	wire [1:0] w_n20588_0;
	wire [2:0] w_n20592_0;
	wire [2:0] w_n20595_0;
	wire [1:0] w_n20596_0;
	wire [2:0] w_n20600_0;
	wire [2:0] w_n20602_0;
	wire [1:0] w_n20603_0;
	wire [2:0] w_n20607_0;
	wire [2:0] w_n20609_0;
	wire [1:0] w_n20610_0;
	wire [2:0] w_n20614_0;
	wire [2:0] w_n20617_0;
	wire [1:0] w_n20618_0;
	wire [2:0] w_n20622_0;
	wire [2:0] w_n20625_0;
	wire [1:0] w_n20626_0;
	wire [2:0] w_n20630_0;
	wire [2:0] w_n20632_0;
	wire [1:0] w_n20633_0;
	wire [2:0] w_n20637_0;
	wire [2:0] w_n20640_0;
	wire [1:0] w_n20641_0;
	wire [2:0] w_n20645_0;
	wire [2:0] w_n20647_0;
	wire [1:0] w_n20648_0;
	wire [2:0] w_n20652_0;
	wire [2:0] w_n20655_0;
	wire [1:0] w_n20656_0;
	wire [2:0] w_n20660_0;
	wire [2:0] w_n20662_0;
	wire [1:0] w_n20663_0;
	wire [2:0] w_n20667_0;
	wire [2:0] w_n20669_0;
	wire [1:0] w_n20670_0;
	wire [2:0] w_n20674_0;
	wire [2:0] w_n20676_0;
	wire [1:0] w_n20677_0;
	wire [2:0] w_n20681_0;
	wire [2:0] w_n20684_0;
	wire [1:0] w_n20685_0;
	wire [2:0] w_n20689_0;
	wire [2:0] w_n20691_0;
	wire [1:0] w_n20692_0;
	wire [2:0] w_n20696_0;
	wire [2:0] w_n20699_0;
	wire [1:0] w_n20700_0;
	wire [2:0] w_n20704_0;
	wire [2:0] w_n20706_0;
	wire [1:0] w_n20707_0;
	wire [2:0] w_n20711_0;
	wire [2:0] w_n20714_0;
	wire [1:0] w_n20715_0;
	wire [2:0] w_n20719_0;
	wire [2:0] w_n20721_0;
	wire [1:0] w_n20722_0;
	wire [2:0] w_n20726_0;
	wire [2:0] w_n20729_0;
	wire [1:0] w_n20730_0;
	wire [2:0] w_n20734_0;
	wire [2:0] w_n20736_0;
	wire [1:0] w_n20737_0;
	wire [2:0] w_n20741_0;
	wire [2:0] w_n20743_0;
	wire [1:0] w_n20744_0;
	wire [2:0] w_n20748_0;
	wire [2:0] w_n20750_0;
	wire [1:0] w_n20751_0;
	wire [2:0] w_n20755_0;
	wire [2:0] w_n20758_0;
	wire [1:0] w_n20759_0;
	wire [2:0] w_n20763_0;
	wire [2:0] w_n20765_0;
	wire [1:0] w_n20766_0;
	wire [2:0] w_n20770_0;
	wire [2:0] w_n20772_0;
	wire [1:0] w_n20773_0;
	wire [2:0] w_n20777_0;
	wire [2:0] w_n20779_0;
	wire [1:0] w_n20780_0;
	wire [2:0] w_n20784_0;
	wire [2:0] w_n20786_0;
	wire [1:0] w_n20787_0;
	wire [2:0] w_n20791_0;
	wire [2:0] w_n20793_0;
	wire [1:0] w_n20794_0;
	wire [2:0] w_n20798_0;
	wire [2:0] w_n20801_0;
	wire [1:0] w_n20802_0;
	wire [2:0] w_n20806_0;
	wire [2:0] w_n20808_0;
	wire [1:0] w_n20809_0;
	wire [2:0] w_n20813_0;
	wire [2:0] w_n20816_0;
	wire [1:0] w_n20817_0;
	wire [2:0] w_n20821_0;
	wire [2:0] w_n20823_0;
	wire [1:0] w_n20824_0;
	wire [2:0] w_n20828_0;
	wire [2:0] w_n20830_0;
	wire [1:0] w_n20831_0;
	wire [2:0] w_n20835_0;
	wire [2:0] w_n20838_0;
	wire [1:0] w_n20839_0;
	wire [2:0] w_n20842_0;
	wire [2:0] w_n20846_0;
	wire [1:0] w_n20847_0;
	wire [2:0] w_n20851_0;
	wire [2:0] w_n20853_0;
	wire [1:0] w_n20854_0;
	wire [1:0] w_n20858_0;
	wire [1:0] w_n20859_0;
	wire [2:0] w_n20861_0;
	wire [1:0] w_n20862_0;
	wire [2:0] w_n20866_0;
	wire [2:0] w_n20868_0;
	wire [1:0] w_n20869_0;
	wire [2:0] w_n20873_0;
	wire [2:0] w_n20875_0;
	wire [1:0] w_n20876_0;
	wire [2:0] w_n20880_0;
	wire [2:0] w_n20883_0;
	wire [1:0] w_n20884_0;
	wire [2:0] w_n20888_0;
	wire [2:0] w_n20890_0;
	wire [1:0] w_n20891_0;
	wire [1:0] w_n20893_0;
	wire [1:0] w_n20896_0;
	wire [1:0] w_n20897_0;
	wire [1:0] w_n20902_0;
	wire [1:0] w_n20903_0;
	wire [2:0] w_n20907_0;
	wire [2:0] w_n20907_1;
	wire [1:0] w_n20908_0;
	wire [2:0] w_n20909_0;
	wire [1:0] w_n20910_0;
	wire [2:0] w_n20912_0;
	wire [1:0] w_n20913_0;
	wire [1:0] w_n20978_0;
	wire [1:0] w_n21175_0;
	wire [1:0] w_n21176_0;
	wire [1:0] w_n21179_0;
	wire [2:0] w_n21181_0;
	wire [1:0] w_n21181_1;
	wire [2:0] w_n21184_0;
	wire [2:0] w_n21184_1;
	wire [2:0] w_n21184_2;
	wire [2:0] w_n21184_3;
	wire [2:0] w_n21184_4;
	wire [2:0] w_n21184_5;
	wire [2:0] w_n21184_6;
	wire [2:0] w_n21184_7;
	wire [2:0] w_n21188_0;
	wire [1:0] w_n21189_0;
	wire [1:0] w_n21191_0;
	wire [1:0] w_n21196_0;
	wire [1:0] w_n21197_0;
	wire [2:0] w_n21199_0;
	wire [1:0] w_n21200_0;
	wire [1:0] w_n21204_0;
	wire [2:0] w_n21206_0;
	wire [1:0] w_n21207_0;
	wire [1:0] w_n21211_0;
	wire [1:0] w_n21212_0;
	wire [2:0] w_n21214_0;
	wire [1:0] w_n21215_0;
	wire [1:0] w_n21219_0;
	wire [2:0] w_n21221_0;
	wire [1:0] w_n21222_0;
	wire [1:0] w_n21226_0;
	wire [1:0] w_n21227_0;
	wire [2:0] w_n21229_0;
	wire [1:0] w_n21230_0;
	wire [1:0] w_n21234_0;
	wire [1:0] w_n21235_0;
	wire [2:0] w_n21237_0;
	wire [1:0] w_n21238_0;
	wire [1:0] w_n21242_0;
	wire [1:0] w_n21243_0;
	wire [2:0] w_n21245_0;
	wire [1:0] w_n21246_0;
	wire [1:0] w_n21250_0;
	wire [2:0] w_n21252_0;
	wire [1:0] w_n21253_0;
	wire [1:0] w_n21257_0;
	wire [1:0] w_n21258_0;
	wire [2:0] w_n21260_0;
	wire [1:0] w_n21261_0;
	wire [1:0] w_n21265_0;
	wire [1:0] w_n21266_0;
	wire [2:0] w_n21268_0;
	wire [1:0] w_n21269_0;
	wire [1:0] w_n21273_0;
	wire [1:0] w_n21274_0;
	wire [2:0] w_n21276_0;
	wire [1:0] w_n21277_0;
	wire [1:0] w_n21281_0;
	wire [2:0] w_n21283_0;
	wire [1:0] w_n21284_0;
	wire [1:0] w_n21288_0;
	wire [1:0] w_n21289_0;
	wire [2:0] w_n21291_0;
	wire [1:0] w_n21292_0;
	wire [1:0] w_n21296_0;
	wire [2:0] w_n21298_0;
	wire [1:0] w_n21299_0;
	wire [1:0] w_n21303_0;
	wire [1:0] w_n21304_0;
	wire [2:0] w_n21306_0;
	wire [1:0] w_n21307_0;
	wire [1:0] w_n21311_0;
	wire [2:0] w_n21313_0;
	wire [1:0] w_n21314_0;
	wire [1:0] w_n21318_0;
	wire [1:0] w_n21319_0;
	wire [2:0] w_n21321_0;
	wire [1:0] w_n21322_0;
	wire [1:0] w_n21326_0;
	wire [1:0] w_n21327_0;
	wire [2:0] w_n21329_0;
	wire [1:0] w_n21330_0;
	wire [1:0] w_n21334_0;
	wire [2:0] w_n21336_0;
	wire [1:0] w_n21337_0;
	wire [1:0] w_n21341_0;
	wire [2:0] w_n21343_0;
	wire [1:0] w_n21344_0;
	wire [1:0] w_n21348_0;
	wire [1:0] w_n21349_0;
	wire [2:0] w_n21351_0;
	wire [1:0] w_n21352_0;
	wire [1:0] w_n21356_0;
	wire [2:0] w_n21358_0;
	wire [1:0] w_n21359_0;
	wire [1:0] w_n21363_0;
	wire [1:0] w_n21364_0;
	wire [2:0] w_n21366_0;
	wire [1:0] w_n21367_0;
	wire [1:0] w_n21371_0;
	wire [2:0] w_n21373_0;
	wire [1:0] w_n21374_0;
	wire [1:0] w_n21378_0;
	wire [1:0] w_n21379_0;
	wire [2:0] w_n21381_0;
	wire [1:0] w_n21382_0;
	wire [1:0] w_n21386_0;
	wire [1:0] w_n21387_0;
	wire [2:0] w_n21389_0;
	wire [1:0] w_n21390_0;
	wire [1:0] w_n21394_0;
	wire [1:0] w_n21395_0;
	wire [2:0] w_n21397_0;
	wire [1:0] w_n21398_0;
	wire [1:0] w_n21402_0;
	wire [2:0] w_n21404_0;
	wire [1:0] w_n21405_0;
	wire [1:0] w_n21409_0;
	wire [1:0] w_n21410_0;
	wire [2:0] w_n21412_0;
	wire [1:0] w_n21413_0;
	wire [1:0] w_n21417_0;
	wire [2:0] w_n21419_0;
	wire [1:0] w_n21420_0;
	wire [1:0] w_n21424_0;
	wire [1:0] w_n21425_0;
	wire [2:0] w_n21427_0;
	wire [1:0] w_n21428_0;
	wire [1:0] w_n21432_0;
	wire [2:0] w_n21434_0;
	wire [1:0] w_n21435_0;
	wire [1:0] w_n21439_0;
	wire [1:0] w_n21440_0;
	wire [2:0] w_n21442_0;
	wire [1:0] w_n21443_0;
	wire [1:0] w_n21447_0;
	wire [2:0] w_n21449_0;
	wire [1:0] w_n21450_0;
	wire [1:0] w_n21454_0;
	wire [1:0] w_n21455_0;
	wire [2:0] w_n21457_0;
	wire [1:0] w_n21458_0;
	wire [1:0] w_n21462_0;
	wire [1:0] w_n21463_0;
	wire [2:0] w_n21465_0;
	wire [1:0] w_n21466_0;
	wire [1:0] w_n21470_0;
	wire [1:0] w_n21471_0;
	wire [2:0] w_n21473_0;
	wire [1:0] w_n21474_0;
	wire [1:0] w_n21478_0;
	wire [2:0] w_n21480_0;
	wire [1:0] w_n21481_0;
	wire [1:0] w_n21485_0;
	wire [1:0] w_n21486_0;
	wire [2:0] w_n21488_0;
	wire [1:0] w_n21489_0;
	wire [1:0] w_n21493_0;
	wire [1:0] w_n21494_0;
	wire [2:0] w_n21496_0;
	wire [1:0] w_n21497_0;
	wire [1:0] w_n21501_0;
	wire [1:0] w_n21502_0;
	wire [2:0] w_n21504_0;
	wire [1:0] w_n21505_0;
	wire [1:0] w_n21509_0;
	wire [1:0] w_n21510_0;
	wire [2:0] w_n21512_0;
	wire [1:0] w_n21513_0;
	wire [1:0] w_n21517_0;
	wire [1:0] w_n21518_0;
	wire [2:0] w_n21520_0;
	wire [1:0] w_n21521_0;
	wire [1:0] w_n21525_0;
	wire [2:0] w_n21527_0;
	wire [1:0] w_n21528_0;
	wire [1:0] w_n21532_0;
	wire [1:0] w_n21533_0;
	wire [2:0] w_n21535_0;
	wire [1:0] w_n21536_0;
	wire [1:0] w_n21540_0;
	wire [2:0] w_n21542_0;
	wire [1:0] w_n21543_0;
	wire [1:0] w_n21547_0;
	wire [1:0] w_n21548_0;
	wire [2:0] w_n21550_0;
	wire [1:0] w_n21551_0;
	wire [1:0] w_n21555_0;
	wire [1:0] w_n21556_0;
	wire [2:0] w_n21558_0;
	wire [1:0] w_n21559_0;
	wire [1:0] w_n21563_0;
	wire [2:0] w_n21565_0;
	wire [1:0] w_n21566_0;
	wire [1:0] w_n21570_0;
	wire [2:0] w_n21572_0;
	wire [1:0] w_n21573_0;
	wire [1:0] w_n21577_0;
	wire [1:0] w_n21578_0;
	wire [2:0] w_n21580_0;
	wire [1:0] w_n21581_0;
	wire [1:0] w_n21585_0;
	wire [1:0] w_n21586_0;
	wire [2:0] w_n21588_0;
	wire [1:0] w_n21589_0;
	wire [1:0] w_n21593_0;
	wire [1:0] w_n21594_0;
	wire [2:0] w_n21596_0;
	wire [1:0] w_n21597_0;
	wire [2:0] w_n21601_0;
	wire [2:0] w_n21604_0;
	wire [1:0] w_n21605_0;
	wire [2:0] w_n21609_0;
	wire [2:0] w_n21611_0;
	wire [1:0] w_n21614_0;
	wire [2:0] w_n21615_0;
	wire [1:0] w_n21616_0;
	wire [1:0] w_n21618_0;
	wire [1:0] w_n21681_0;
	wire [1:0] w_n21688_0;
	wire [1:0] w_n21695_0;
	wire [1:0] w_n21708_0;
	wire [1:0] w_n21721_0;
	wire [1:0] w_n21728_0;
	wire [1:0] w_n21735_0;
	wire [1:0] w_n21745_0;
	wire [1:0] w_n21749_0;
	wire [1:0] w_n21756_0;
	wire [1:0] w_n21763_0;
	wire [1:0] w_n21776_0;
	wire [1:0] w_n21783_0;
	wire [1:0] w_n21790_0;
	wire [1:0] w_n21797_0;
	wire [1:0] w_n21810_0;
	wire [1:0] w_n21829_0;
	wire [1:0] w_n21836_0;
	wire [1:0] w_n21846_0;
	wire [1:0] w_n21850_0;
	wire [1:0] w_n21868_0;
	wire [1:0] w_n21877_0;
	wire [2:0] w_n21887_0;
	wire [2:0] w_n21887_1;
	wire [2:0] w_n21887_2;
	wire [2:0] w_n21887_3;
	wire [2:0] w_n21887_4;
	wire [2:0] w_n21887_5;
	wire [2:0] w_n21887_6;
	wire [2:0] w_n21887_7;
	wire [2:0] w_n21887_8;
	wire [2:0] w_n21887_9;
	wire [2:0] w_n21887_10;
	wire [2:0] w_n21887_11;
	wire [2:0] w_n21887_12;
	wire [2:0] w_n21887_13;
	wire [2:0] w_n21887_14;
	wire [2:0] w_n21887_15;
	wire [2:0] w_n21887_16;
	wire [2:0] w_n21887_17;
	wire [2:0] w_n21887_18;
	wire [2:0] w_n21887_19;
	wire [2:0] w_n21887_20;
	wire [2:0] w_n21887_21;
	wire [2:0] w_n21887_22;
	wire [2:0] w_n21887_23;
	wire [2:0] w_n21887_24;
	wire [2:0] w_n21887_25;
	wire [2:0] w_n21887_26;
	wire [2:0] w_n21887_27;
	wire [2:0] w_n21887_28;
	wire [2:0] w_n21887_29;
	wire [2:0] w_n21887_30;
	wire [2:0] w_n21887_31;
	wire [2:0] w_n21887_32;
	wire [2:0] w_n21887_33;
	wire [1:0] w_n21887_34;
	wire [2:0] w_n21889_0;
	wire [2:0] w_n21889_1;
	wire [1:0] w_n21890_0;
	wire [2:0] w_n21891_0;
	wire [1:0] w_n21892_0;
	wire [2:0] w_n21894_0;
	wire [1:0] w_n21895_0;
	wire [2:0] w_n21902_0;
	wire [1:0] w_n21903_0;
	wire [1:0] w_n21906_0;
	wire [1:0] w_n21909_0;
	wire [2:0] w_n21911_0;
	wire [1:0] w_n21912_0;
	wire [2:0] w_n21916_0;
	wire [2:0] w_n21919_0;
	wire [1:0] w_n21920_0;
	wire [2:0] w_n21924_0;
	wire [2:0] w_n21926_0;
	wire [1:0] w_n21927_0;
	wire [2:0] w_n21931_0;
	wire [2:0] w_n21934_0;
	wire [1:0] w_n21935_0;
	wire [2:0] w_n21939_0;
	wire [2:0] w_n21941_0;
	wire [1:0] w_n21942_0;
	wire [2:0] w_n21946_0;
	wire [2:0] w_n21949_0;
	wire [1:0] w_n21950_0;
	wire [2:0] w_n21954_0;
	wire [2:0] w_n21956_0;
	wire [1:0] w_n21957_0;
	wire [2:0] w_n21961_0;
	wire [2:0] w_n21963_0;
	wire [1:0] w_n21964_0;
	wire [2:0] w_n21968_0;
	wire [2:0] w_n21970_0;
	wire [1:0] w_n21971_0;
	wire [2:0] w_n21975_0;
	wire [2:0] w_n21978_0;
	wire [1:0] w_n21979_0;
	wire [2:0] w_n21983_0;
	wire [2:0] w_n21985_0;
	wire [1:0] w_n21986_0;
	wire [2:0] w_n21990_0;
	wire [2:0] w_n21992_0;
	wire [1:0] w_n21993_0;
	wire [2:0] w_n21997_0;
	wire [2:0] w_n21999_0;
	wire [1:0] w_n22000_0;
	wire [2:0] w_n22004_0;
	wire [2:0] w_n22007_0;
	wire [1:0] w_n22008_0;
	wire [2:0] w_n22012_0;
	wire [2:0] w_n22014_0;
	wire [1:0] w_n22015_0;
	wire [2:0] w_n22019_0;
	wire [2:0] w_n22022_0;
	wire [1:0] w_n22023_0;
	wire [2:0] w_n22027_0;
	wire [2:0] w_n22029_0;
	wire [1:0] w_n22030_0;
	wire [2:0] w_n22034_0;
	wire [2:0] w_n22037_0;
	wire [1:0] w_n22038_0;
	wire [2:0] w_n22042_0;
	wire [2:0] w_n22044_0;
	wire [1:0] w_n22045_0;
	wire [2:0] w_n22049_0;
	wire [2:0] w_n22051_0;
	wire [1:0] w_n22052_0;
	wire [2:0] w_n22056_0;
	wire [2:0] w_n22059_0;
	wire [1:0] w_n22060_0;
	wire [2:0] w_n22064_0;
	wire [2:0] w_n22067_0;
	wire [1:0] w_n22068_0;
	wire [2:0] w_n22072_0;
	wire [2:0] w_n22074_0;
	wire [1:0] w_n22075_0;
	wire [2:0] w_n22079_0;
	wire [2:0] w_n22082_0;
	wire [1:0] w_n22083_0;
	wire [2:0] w_n22087_0;
	wire [2:0] w_n22089_0;
	wire [1:0] w_n22090_0;
	wire [2:0] w_n22094_0;
	wire [2:0] w_n22097_0;
	wire [1:0] w_n22098_0;
	wire [2:0] w_n22102_0;
	wire [2:0] w_n22104_0;
	wire [1:0] w_n22105_0;
	wire [2:0] w_n22109_0;
	wire [2:0] w_n22111_0;
	wire [1:0] w_n22112_0;
	wire [2:0] w_n22116_0;
	wire [2:0] w_n22118_0;
	wire [1:0] w_n22119_0;
	wire [2:0] w_n22123_0;
	wire [2:0] w_n22126_0;
	wire [1:0] w_n22127_0;
	wire [2:0] w_n22131_0;
	wire [2:0] w_n22133_0;
	wire [1:0] w_n22134_0;
	wire [2:0] w_n22138_0;
	wire [2:0] w_n22141_0;
	wire [1:0] w_n22142_0;
	wire [2:0] w_n22146_0;
	wire [2:0] w_n22148_0;
	wire [1:0] w_n22149_0;
	wire [2:0] w_n22153_0;
	wire [2:0] w_n22156_0;
	wire [1:0] w_n22157_0;
	wire [2:0] w_n22161_0;
	wire [2:0] w_n22163_0;
	wire [1:0] w_n22164_0;
	wire [2:0] w_n22168_0;
	wire [2:0] w_n22171_0;
	wire [1:0] w_n22172_0;
	wire [2:0] w_n22176_0;
	wire [2:0] w_n22178_0;
	wire [1:0] w_n22179_0;
	wire [2:0] w_n22183_0;
	wire [2:0] w_n22185_0;
	wire [1:0] w_n22186_0;
	wire [2:0] w_n22190_0;
	wire [2:0] w_n22192_0;
	wire [1:0] w_n22193_0;
	wire [2:0] w_n22197_0;
	wire [2:0] w_n22200_0;
	wire [1:0] w_n22201_0;
	wire [2:0] w_n22205_0;
	wire [2:0] w_n22207_0;
	wire [1:0] w_n22208_0;
	wire [2:0] w_n22212_0;
	wire [2:0] w_n22214_0;
	wire [1:0] w_n22215_0;
	wire [2:0] w_n22219_0;
	wire [2:0] w_n22221_0;
	wire [1:0] w_n22222_0;
	wire [2:0] w_n22226_0;
	wire [2:0] w_n22228_0;
	wire [1:0] w_n22229_0;
	wire [2:0] w_n22233_0;
	wire [2:0] w_n22235_0;
	wire [1:0] w_n22236_0;
	wire [2:0] w_n22240_0;
	wire [2:0] w_n22243_0;
	wire [1:0] w_n22244_0;
	wire [2:0] w_n22248_0;
	wire [2:0] w_n22250_0;
	wire [1:0] w_n22251_0;
	wire [2:0] w_n22255_0;
	wire [2:0] w_n22258_0;
	wire [1:0] w_n22259_0;
	wire [2:0] w_n22263_0;
	wire [2:0] w_n22265_0;
	wire [1:0] w_n22266_0;
	wire [2:0] w_n22270_0;
	wire [2:0] w_n22272_0;
	wire [1:0] w_n22273_0;
	wire [2:0] w_n22277_0;
	wire [2:0] w_n22280_0;
	wire [1:0] w_n22281_0;
	wire [2:0] w_n22285_0;
	wire [2:0] w_n22288_0;
	wire [1:0] w_n22289_0;
	wire [2:0] w_n22293_0;
	wire [2:0] w_n22295_0;
	wire [1:0] w_n22296_0;
	wire [2:0] w_n22300_0;
	wire [2:0] w_n22302_0;
	wire [1:0] w_n22303_0;
	wire [2:0] w_n22307_0;
	wire [2:0] w_n22309_0;
	wire [1:0] w_n22310_0;
	wire [1:0] w_n22314_0;
	wire [1:0] w_n22315_0;
	wire [2:0] w_n22317_0;
	wire [1:0] w_n22317_1;
	wire [2:0] w_n22320_0;
	wire [1:0] w_n22320_1;
	wire [2:0] w_n22321_0;
	wire [1:0] w_n22324_0;
	wire [1:0] w_n22325_0;
	wire [1:0] w_n22330_0;
	wire [1:0] w_n22332_0;
	wire [2:0] w_n22334_0;
	wire [2:0] w_n22334_1;
	wire [1:0] w_n22335_0;
	wire [2:0] w_n22336_0;
	wire [1:0] w_n22337_0;
	wire [2:0] w_n22339_0;
	wire [1:0] w_n22340_0;
	wire [1:0] w_n22345_0;
	wire [1:0] w_n22408_0;
	wire [1:0] w_n22412_0;
	wire [1:0] w_n22615_0;
	wire [1:0] w_n22619_0;
	wire [2:0] w_n22620_0;
	wire [2:0] w_n22620_1;
	wire [2:0] w_n22620_2;
	wire [2:0] w_n22620_3;
	wire [2:0] w_n22620_4;
	wire [1:0] w_n22621_0;
	wire [1:0] w_n22622_0;
	wire [2:0] w_n22624_0;
	wire [1:0] w_n22625_0;
	wire [1:0] w_n22629_0;
	wire [1:0] w_n22630_0;
	wire [2:0] w_n22632_0;
	wire [1:0] w_n22633_0;
	wire [1:0] w_n22637_0;
	wire [2:0] w_n22639_0;
	wire [1:0] w_n22640_0;
	wire [1:0] w_n22644_0;
	wire [2:0] w_n22646_0;
	wire [1:0] w_n22647_0;
	wire [1:0] w_n22651_0;
	wire [2:0] w_n22653_0;
	wire [1:0] w_n22654_0;
	wire [1:0] w_n22658_0;
	wire [1:0] w_n22659_0;
	wire [2:0] w_n22661_0;
	wire [1:0] w_n22662_0;
	wire [1:0] w_n22666_0;
	wire [2:0] w_n22668_0;
	wire [1:0] w_n22669_0;
	wire [1:0] w_n22673_0;
	wire [1:0] w_n22674_0;
	wire [2:0] w_n22676_0;
	wire [1:0] w_n22677_0;
	wire [1:0] w_n22681_0;
	wire [2:0] w_n22683_0;
	wire [1:0] w_n22684_0;
	wire [1:0] w_n22688_0;
	wire [1:0] w_n22689_0;
	wire [2:0] w_n22691_0;
	wire [1:0] w_n22692_0;
	wire [1:0] w_n22696_0;
	wire [1:0] w_n22697_0;
	wire [2:0] w_n22699_0;
	wire [1:0] w_n22700_0;
	wire [1:0] w_n22704_0;
	wire [1:0] w_n22705_0;
	wire [2:0] w_n22707_0;
	wire [1:0] w_n22708_0;
	wire [1:0] w_n22712_0;
	wire [2:0] w_n22714_0;
	wire [1:0] w_n22715_0;
	wire [1:0] w_n22719_0;
	wire [1:0] w_n22720_0;
	wire [2:0] w_n22722_0;
	wire [1:0] w_n22723_0;
	wire [1:0] w_n22727_0;
	wire [1:0] w_n22728_0;
	wire [2:0] w_n22730_0;
	wire [1:0] w_n22731_0;
	wire [1:0] w_n22735_0;
	wire [1:0] w_n22736_0;
	wire [2:0] w_n22738_0;
	wire [1:0] w_n22739_0;
	wire [1:0] w_n22743_0;
	wire [2:0] w_n22745_0;
	wire [1:0] w_n22746_0;
	wire [1:0] w_n22750_0;
	wire [1:0] w_n22751_0;
	wire [2:0] w_n22753_0;
	wire [1:0] w_n22754_0;
	wire [1:0] w_n22758_0;
	wire [2:0] w_n22760_0;
	wire [1:0] w_n22761_0;
	wire [1:0] w_n22765_0;
	wire [1:0] w_n22766_0;
	wire [2:0] w_n22768_0;
	wire [1:0] w_n22769_0;
	wire [1:0] w_n22773_0;
	wire [2:0] w_n22775_0;
	wire [1:0] w_n22776_0;
	wire [1:0] w_n22780_0;
	wire [1:0] w_n22781_0;
	wire [2:0] w_n22783_0;
	wire [1:0] w_n22784_0;
	wire [1:0] w_n22788_0;
	wire [1:0] w_n22789_0;
	wire [2:0] w_n22791_0;
	wire [1:0] w_n22792_0;
	wire [1:0] w_n22796_0;
	wire [2:0] w_n22798_0;
	wire [1:0] w_n22799_0;
	wire [1:0] w_n22803_0;
	wire [2:0] w_n22805_0;
	wire [1:0] w_n22806_0;
	wire [1:0] w_n22810_0;
	wire [1:0] w_n22811_0;
	wire [2:0] w_n22813_0;
	wire [1:0] w_n22814_0;
	wire [1:0] w_n22818_0;
	wire [2:0] w_n22820_0;
	wire [1:0] w_n22821_0;
	wire [1:0] w_n22825_0;
	wire [1:0] w_n22826_0;
	wire [2:0] w_n22828_0;
	wire [1:0] w_n22829_0;
	wire [1:0] w_n22833_0;
	wire [2:0] w_n22835_0;
	wire [1:0] w_n22836_0;
	wire [1:0] w_n22840_0;
	wire [1:0] w_n22841_0;
	wire [2:0] w_n22843_0;
	wire [1:0] w_n22844_0;
	wire [1:0] w_n22848_0;
	wire [1:0] w_n22849_0;
	wire [2:0] w_n22851_0;
	wire [1:0] w_n22852_0;
	wire [1:0] w_n22856_0;
	wire [1:0] w_n22857_0;
	wire [2:0] w_n22859_0;
	wire [1:0] w_n22860_0;
	wire [1:0] w_n22864_0;
	wire [2:0] w_n22866_0;
	wire [1:0] w_n22867_0;
	wire [1:0] w_n22871_0;
	wire [1:0] w_n22872_0;
	wire [2:0] w_n22874_0;
	wire [1:0] w_n22875_0;
	wire [1:0] w_n22879_0;
	wire [2:0] w_n22881_0;
	wire [1:0] w_n22882_0;
	wire [1:0] w_n22886_0;
	wire [1:0] w_n22887_0;
	wire [2:0] w_n22889_0;
	wire [1:0] w_n22890_0;
	wire [1:0] w_n22894_0;
	wire [2:0] w_n22896_0;
	wire [1:0] w_n22897_0;
	wire [1:0] w_n22901_0;
	wire [1:0] w_n22902_0;
	wire [2:0] w_n22904_0;
	wire [1:0] w_n22905_0;
	wire [1:0] w_n22909_0;
	wire [2:0] w_n22911_0;
	wire [1:0] w_n22912_0;
	wire [1:0] w_n22916_0;
	wire [1:0] w_n22917_0;
	wire [2:0] w_n22919_0;
	wire [1:0] w_n22920_0;
	wire [1:0] w_n22924_0;
	wire [1:0] w_n22925_0;
	wire [2:0] w_n22927_0;
	wire [1:0] w_n22928_0;
	wire [1:0] w_n22932_0;
	wire [1:0] w_n22933_0;
	wire [2:0] w_n22935_0;
	wire [1:0] w_n22936_0;
	wire [1:0] w_n22940_0;
	wire [2:0] w_n22942_0;
	wire [1:0] w_n22943_0;
	wire [1:0] w_n22947_0;
	wire [1:0] w_n22948_0;
	wire [2:0] w_n22950_0;
	wire [1:0] w_n22951_0;
	wire [1:0] w_n22955_0;
	wire [1:0] w_n22956_0;
	wire [2:0] w_n22958_0;
	wire [1:0] w_n22959_0;
	wire [1:0] w_n22963_0;
	wire [1:0] w_n22964_0;
	wire [2:0] w_n22966_0;
	wire [1:0] w_n22967_0;
	wire [1:0] w_n22971_0;
	wire [1:0] w_n22972_0;
	wire [2:0] w_n22974_0;
	wire [1:0] w_n22975_0;
	wire [1:0] w_n22979_0;
	wire [1:0] w_n22980_0;
	wire [2:0] w_n22982_0;
	wire [1:0] w_n22983_0;
	wire [1:0] w_n22987_0;
	wire [2:0] w_n22989_0;
	wire [1:0] w_n22990_0;
	wire [1:0] w_n22994_0;
	wire [1:0] w_n22995_0;
	wire [2:0] w_n22997_0;
	wire [1:0] w_n22998_0;
	wire [1:0] w_n23002_0;
	wire [2:0] w_n23004_0;
	wire [1:0] w_n23005_0;
	wire [1:0] w_n23009_0;
	wire [1:0] w_n23010_0;
	wire [2:0] w_n23012_0;
	wire [1:0] w_n23013_0;
	wire [1:0] w_n23017_0;
	wire [1:0] w_n23018_0;
	wire [2:0] w_n23020_0;
	wire [1:0] w_n23021_0;
	wire [1:0] w_n23025_0;
	wire [2:0] w_n23027_0;
	wire [1:0] w_n23028_0;
	wire [1:0] w_n23032_0;
	wire [2:0] w_n23034_0;
	wire [1:0] w_n23035_0;
	wire [1:0] w_n23039_0;
	wire [1:0] w_n23040_0;
	wire [2:0] w_n23042_0;
	wire [1:0] w_n23043_0;
	wire [1:0] w_n23047_0;
	wire [1:0] w_n23048_0;
	wire [2:0] w_n23050_0;
	wire [1:0] w_n23051_0;
	wire [2:0] w_n23055_0;
	wire [1:0] w_n23058_0;
	wire [1:0] w_n23061_0;
	wire [1:0] w_n23062_0;
	wire [2:0] w_n23063_0;
	wire [1:0] w_n23063_1;
	wire [1:0] w_n23064_0;
	wire [1:0] w_n23065_0;
	wire [1:0] w_n23138_0;
	wire [1:0] w_n23142_0;
	wire [1:0] w_n23146_0;
	wire [1:0] w_n23153_0;
	wire [1:0] w_n23160_0;
	wire [1:0] w_n23173_0;
	wire [1:0] w_n23186_0;
	wire [1:0] w_n23193_0;
	wire [1:0] w_n23200_0;
	wire [1:0] w_n23210_0;
	wire [1:0] w_n23214_0;
	wire [1:0] w_n23221_0;
	wire [1:0] w_n23228_0;
	wire [1:0] w_n23241_0;
	wire [1:0] w_n23248_0;
	wire [1:0] w_n23255_0;
	wire [1:0] w_n23262_0;
	wire [1:0] w_n23275_0;
	wire [1:0] w_n23294_0;
	wire [1:0] w_n23301_0;
	wire [1:0] w_n23311_0;
	wire [1:0] w_n23315_0;
	wire [1:0] w_n23326_0;
	wire [1:0] w_n23327_0;
	wire [1:0] w_n23335_0;
	wire [1:0] w_n23336_0;
	wire [1:0] w_n23339_0;
	wire [1:0] w_n23344_0;
	wire [2:0] w_n23345_0;
	wire [2:0] w_n23345_1;
	wire [2:0] w_n23345_2;
	wire [2:0] w_n23345_3;
	wire [2:0] w_n23345_4;
	wire [2:0] w_n23345_5;
	wire [2:0] w_n23345_6;
	wire [2:0] w_n23345_7;
	wire [2:0] w_n23345_8;
	wire [2:0] w_n23345_9;
	wire [2:0] w_n23345_10;
	wire [2:0] w_n23345_11;
	wire [2:0] w_n23345_12;
	wire [2:0] w_n23345_13;
	wire [2:0] w_n23345_14;
	wire [2:0] w_n23345_15;
	wire [2:0] w_n23345_16;
	wire [2:0] w_n23345_17;
	wire [2:0] w_n23345_18;
	wire [2:0] w_n23345_19;
	wire [2:0] w_n23345_20;
	wire [2:0] w_n23345_21;
	wire [2:0] w_n23345_22;
	wire [2:0] w_n23345_23;
	wire [2:0] w_n23345_24;
	wire [2:0] w_n23345_25;
	wire [2:0] w_n23345_26;
	wire [2:0] w_n23345_27;
	wire [2:0] w_n23345_28;
	wire [2:0] w_n23345_29;
	wire [2:0] w_n23345_30;
	wire [2:0] w_n23345_31;
	wire [1:0] w_n23345_32;
	wire [1:0] w_n23348_0;
	wire [2:0] w_n23349_0;
	wire [2:0] w_n23351_0;
	wire [1:0] w_n23351_1;
	wire [1:0] w_n23352_0;
	wire [2:0] w_n23353_0;
	wire [1:0] w_n23354_0;
	wire [2:0] w_n23356_0;
	wire [1:0] w_n23357_0;
	wire [2:0] w_n23364_0;
	wire [1:0] w_n23365_0;
	wire [1:0] w_n23368_0;
	wire [1:0] w_n23371_0;
	wire [2:0] w_n23373_0;
	wire [1:0] w_n23374_0;
	wire [2:0] w_n23378_0;
	wire [2:0] w_n23380_0;
	wire [1:0] w_n23381_0;
	wire [2:0] w_n23385_0;
	wire [2:0] w_n23387_0;
	wire [1:0] w_n23388_0;
	wire [2:0] w_n23392_0;
	wire [2:0] w_n23395_0;
	wire [1:0] w_n23396_0;
	wire [2:0] w_n23400_0;
	wire [2:0] w_n23403_0;
	wire [1:0] w_n23404_0;
	wire [2:0] w_n23408_0;
	wire [2:0] w_n23411_0;
	wire [1:0] w_n23412_0;
	wire [2:0] w_n23416_0;
	wire [2:0] w_n23418_0;
	wire [1:0] w_n23419_0;
	wire [2:0] w_n23423_0;
	wire [2:0] w_n23426_0;
	wire [1:0] w_n23427_0;
	wire [2:0] w_n23431_0;
	wire [2:0] w_n23433_0;
	wire [1:0] w_n23434_0;
	wire [2:0] w_n23438_0;
	wire [2:0] w_n23441_0;
	wire [1:0] w_n23442_0;
	wire [2:0] w_n23446_0;
	wire [2:0] w_n23448_0;
	wire [1:0] w_n23449_0;
	wire [2:0] w_n23453_0;
	wire [2:0] w_n23455_0;
	wire [1:0] w_n23456_0;
	wire [2:0] w_n23460_0;
	wire [2:0] w_n23462_0;
	wire [1:0] w_n23463_0;
	wire [2:0] w_n23467_0;
	wire [2:0] w_n23470_0;
	wire [1:0] w_n23471_0;
	wire [2:0] w_n23475_0;
	wire [2:0] w_n23477_0;
	wire [1:0] w_n23478_0;
	wire [2:0] w_n23482_0;
	wire [2:0] w_n23484_0;
	wire [1:0] w_n23485_0;
	wire [2:0] w_n23489_0;
	wire [2:0] w_n23491_0;
	wire [1:0] w_n23492_0;
	wire [2:0] w_n23496_0;
	wire [2:0] w_n23499_0;
	wire [1:0] w_n23500_0;
	wire [2:0] w_n23504_0;
	wire [2:0] w_n23506_0;
	wire [1:0] w_n23507_0;
	wire [2:0] w_n23511_0;
	wire [2:0] w_n23514_0;
	wire [1:0] w_n23515_0;
	wire [2:0] w_n23519_0;
	wire [2:0] w_n23521_0;
	wire [1:0] w_n23522_0;
	wire [2:0] w_n23526_0;
	wire [2:0] w_n23529_0;
	wire [1:0] w_n23530_0;
	wire [2:0] w_n23534_0;
	wire [2:0] w_n23536_0;
	wire [1:0] w_n23537_0;
	wire [2:0] w_n23541_0;
	wire [2:0] w_n23543_0;
	wire [1:0] w_n23544_0;
	wire [2:0] w_n23548_0;
	wire [2:0] w_n23551_0;
	wire [1:0] w_n23552_0;
	wire [2:0] w_n23556_0;
	wire [2:0] w_n23559_0;
	wire [1:0] w_n23560_0;
	wire [2:0] w_n23564_0;
	wire [2:0] w_n23566_0;
	wire [1:0] w_n23567_0;
	wire [2:0] w_n23571_0;
	wire [2:0] w_n23574_0;
	wire [1:0] w_n23575_0;
	wire [2:0] w_n23579_0;
	wire [2:0] w_n23581_0;
	wire [1:0] w_n23582_0;
	wire [2:0] w_n23586_0;
	wire [2:0] w_n23589_0;
	wire [1:0] w_n23590_0;
	wire [2:0] w_n23594_0;
	wire [2:0] w_n23596_0;
	wire [1:0] w_n23597_0;
	wire [2:0] w_n23601_0;
	wire [2:0] w_n23603_0;
	wire [1:0] w_n23604_0;
	wire [2:0] w_n23608_0;
	wire [2:0] w_n23610_0;
	wire [1:0] w_n23611_0;
	wire [2:0] w_n23615_0;
	wire [2:0] w_n23618_0;
	wire [1:0] w_n23619_0;
	wire [2:0] w_n23623_0;
	wire [2:0] w_n23625_0;
	wire [1:0] w_n23626_0;
	wire [2:0] w_n23630_0;
	wire [2:0] w_n23633_0;
	wire [1:0] w_n23634_0;
	wire [2:0] w_n23638_0;
	wire [2:0] w_n23640_0;
	wire [1:0] w_n23641_0;
	wire [2:0] w_n23645_0;
	wire [2:0] w_n23648_0;
	wire [1:0] w_n23649_0;
	wire [2:0] w_n23653_0;
	wire [2:0] w_n23655_0;
	wire [1:0] w_n23656_0;
	wire [2:0] w_n23660_0;
	wire [2:0] w_n23663_0;
	wire [1:0] w_n23664_0;
	wire [2:0] w_n23668_0;
	wire [2:0] w_n23670_0;
	wire [1:0] w_n23671_0;
	wire [2:0] w_n23675_0;
	wire [2:0] w_n23677_0;
	wire [1:0] w_n23678_0;
	wire [2:0] w_n23682_0;
	wire [2:0] w_n23684_0;
	wire [1:0] w_n23685_0;
	wire [2:0] w_n23689_0;
	wire [2:0] w_n23692_0;
	wire [1:0] w_n23693_0;
	wire [2:0] w_n23697_0;
	wire [2:0] w_n23699_0;
	wire [1:0] w_n23700_0;
	wire [2:0] w_n23704_0;
	wire [2:0] w_n23706_0;
	wire [1:0] w_n23707_0;
	wire [2:0] w_n23711_0;
	wire [2:0] w_n23713_0;
	wire [1:0] w_n23714_0;
	wire [2:0] w_n23718_0;
	wire [2:0] w_n23720_0;
	wire [1:0] w_n23721_0;
	wire [2:0] w_n23725_0;
	wire [2:0] w_n23727_0;
	wire [1:0] w_n23728_0;
	wire [2:0] w_n23732_0;
	wire [2:0] w_n23735_0;
	wire [1:0] w_n23736_0;
	wire [2:0] w_n23740_0;
	wire [2:0] w_n23742_0;
	wire [1:0] w_n23743_0;
	wire [2:0] w_n23747_0;
	wire [2:0] w_n23750_0;
	wire [1:0] w_n23751_0;
	wire [2:0] w_n23755_0;
	wire [2:0] w_n23757_0;
	wire [1:0] w_n23758_0;
	wire [1:0] w_n23762_0;
	wire [2:0] w_n23764_0;
	wire [1:0] w_n23765_0;
	wire [2:0] w_n23769_0;
	wire [2:0] w_n23772_0;
	wire [1:0] w_n23773_0;
	wire [2:0] w_n23777_0;
	wire [2:0] w_n23780_0;
	wire [1:0] w_n23781_0;
	wire [2:0] w_n23785_0;
	wire [2:0] w_n23787_0;
	wire [1:0] w_n23788_0;
	wire [2:0] w_n23792_0;
	wire [2:0] w_n23794_0;
	wire [1:0] w_n23794_1;
	wire [2:0] w_n23795_0;
	wire [1:0] w_n23796_0;
	wire [1:0] w_n23805_0;
	wire [1:0] w_n23806_0;
	wire [1:0] w_n23810_0;
	wire [1:0] w_n23811_0;
	wire [2:0] w_n23812_0;
	wire [1:0] w_n23813_0;
	wire [1:0] w_n23818_0;
	wire [1:0] w_n23884_0;
	wire [1:0] w_n23888_0;
	wire [1:0] w_n24080_0;
	wire [1:0] w_n24097_0;
	wire [1:0] w_n24102_0;
	wire [2:0] w_n24103_0;
	wire [2:0] w_n24103_1;
	wire [1:0] w_n24104_0;
	wire [1:0] w_n24105_0;
	wire [2:0] w_n24107_0;
	wire [1:0] w_n24108_0;
	wire [1:0] w_n24112_0;
	wire [1:0] w_n24113_0;
	wire [2:0] w_n24115_0;
	wire [1:0] w_n24116_0;
	wire [2:0] w_n24120_0;
	wire [2:0] w_n24122_0;
	wire [1:0] w_n24123_0;
	wire [2:0] w_n24127_0;
	wire [2:0] w_n24129_0;
	wire [1:0] w_n24130_0;
	wire [1:0] w_n24134_0;
	wire [1:0] w_n24135_0;
	wire [2:0] w_n24137_0;
	wire [1:0] w_n24138_0;
	wire [1:0] w_n24142_0;
	wire [1:0] w_n24143_0;
	wire [2:0] w_n24145_0;
	wire [1:0] w_n24146_0;
	wire [2:0] w_n24150_0;
	wire [2:0] w_n24152_0;
	wire [1:0] w_n24153_0;
	wire [2:0] w_n24157_0;
	wire [2:0] w_n24159_0;
	wire [1:0] w_n24160_0;
	wire [2:0] w_n24164_0;
	wire [2:0] w_n24166_0;
	wire [1:0] w_n24167_0;
	wire [1:0] w_n24171_0;
	wire [1:0] w_n24172_0;
	wire [2:0] w_n24174_0;
	wire [1:0] w_n24175_0;
	wire [2:0] w_n24179_0;
	wire [2:0] w_n24181_0;
	wire [1:0] w_n24182_0;
	wire [1:0] w_n24186_0;
	wire [1:0] w_n24187_0;
	wire [2:0] w_n24189_0;
	wire [1:0] w_n24190_0;
	wire [2:0] w_n24194_0;
	wire [2:0] w_n24196_0;
	wire [1:0] w_n24197_0;
	wire [1:0] w_n24201_0;
	wire [1:0] w_n24202_0;
	wire [2:0] w_n24204_0;
	wire [1:0] w_n24205_0;
	wire [1:0] w_n24209_0;
	wire [1:0] w_n24210_0;
	wire [2:0] w_n24212_0;
	wire [1:0] w_n24213_0;
	wire [1:0] w_n24217_0;
	wire [1:0] w_n24218_0;
	wire [2:0] w_n24220_0;
	wire [1:0] w_n24221_0;
	wire [2:0] w_n24225_0;
	wire [2:0] w_n24227_0;
	wire [1:0] w_n24228_0;
	wire [1:0] w_n24232_0;
	wire [1:0] w_n24233_0;
	wire [2:0] w_n24235_0;
	wire [1:0] w_n24236_0;
	wire [1:0] w_n24240_0;
	wire [1:0] w_n24241_0;
	wire [2:0] w_n24243_0;
	wire [1:0] w_n24244_0;
	wire [1:0] w_n24248_0;
	wire [1:0] w_n24249_0;
	wire [2:0] w_n24251_0;
	wire [1:0] w_n24252_0;
	wire [2:0] w_n24256_0;
	wire [2:0] w_n24258_0;
	wire [1:0] w_n24259_0;
	wire [1:0] w_n24263_0;
	wire [1:0] w_n24264_0;
	wire [2:0] w_n24266_0;
	wire [1:0] w_n24267_0;
	wire [2:0] w_n24271_0;
	wire [2:0] w_n24273_0;
	wire [1:0] w_n24274_0;
	wire [1:0] w_n24278_0;
	wire [1:0] w_n24279_0;
	wire [2:0] w_n24281_0;
	wire [1:0] w_n24282_0;
	wire [2:0] w_n24286_0;
	wire [2:0] w_n24288_0;
	wire [1:0] w_n24289_0;
	wire [1:0] w_n24293_0;
	wire [1:0] w_n24294_0;
	wire [2:0] w_n24296_0;
	wire [1:0] w_n24297_0;
	wire [1:0] w_n24301_0;
	wire [1:0] w_n24302_0;
	wire [2:0] w_n24304_0;
	wire [1:0] w_n24305_0;
	wire [2:0] w_n24309_0;
	wire [2:0] w_n24311_0;
	wire [1:0] w_n24312_0;
	wire [2:0] w_n24316_0;
	wire [2:0] w_n24318_0;
	wire [1:0] w_n24319_0;
	wire [1:0] w_n24323_0;
	wire [1:0] w_n24324_0;
	wire [2:0] w_n24326_0;
	wire [1:0] w_n24327_0;
	wire [2:0] w_n24331_0;
	wire [2:0] w_n24333_0;
	wire [1:0] w_n24334_0;
	wire [1:0] w_n24338_0;
	wire [1:0] w_n24339_0;
	wire [2:0] w_n24341_0;
	wire [1:0] w_n24342_0;
	wire [2:0] w_n24346_0;
	wire [2:0] w_n24348_0;
	wire [1:0] w_n24349_0;
	wire [1:0] w_n24353_0;
	wire [1:0] w_n24354_0;
	wire [2:0] w_n24356_0;
	wire [1:0] w_n24357_0;
	wire [1:0] w_n24361_0;
	wire [1:0] w_n24362_0;
	wire [2:0] w_n24364_0;
	wire [1:0] w_n24365_0;
	wire [1:0] w_n24369_0;
	wire [1:0] w_n24370_0;
	wire [2:0] w_n24372_0;
	wire [1:0] w_n24373_0;
	wire [2:0] w_n24377_0;
	wire [2:0] w_n24379_0;
	wire [1:0] w_n24380_0;
	wire [1:0] w_n24384_0;
	wire [1:0] w_n24385_0;
	wire [2:0] w_n24387_0;
	wire [1:0] w_n24388_0;
	wire [2:0] w_n24392_0;
	wire [2:0] w_n24394_0;
	wire [1:0] w_n24395_0;
	wire [1:0] w_n24399_0;
	wire [1:0] w_n24400_0;
	wire [2:0] w_n24402_0;
	wire [1:0] w_n24403_0;
	wire [2:0] w_n24407_0;
	wire [2:0] w_n24409_0;
	wire [1:0] w_n24410_0;
	wire [1:0] w_n24414_0;
	wire [1:0] w_n24415_0;
	wire [2:0] w_n24417_0;
	wire [1:0] w_n24418_0;
	wire [2:0] w_n24422_0;
	wire [2:0] w_n24424_0;
	wire [1:0] w_n24425_0;
	wire [1:0] w_n24429_0;
	wire [1:0] w_n24430_0;
	wire [2:0] w_n24432_0;
	wire [1:0] w_n24433_0;
	wire [1:0] w_n24437_0;
	wire [1:0] w_n24438_0;
	wire [2:0] w_n24440_0;
	wire [1:0] w_n24441_0;
	wire [1:0] w_n24445_0;
	wire [1:0] w_n24446_0;
	wire [2:0] w_n24448_0;
	wire [1:0] w_n24449_0;
	wire [2:0] w_n24453_0;
	wire [2:0] w_n24455_0;
	wire [1:0] w_n24456_0;
	wire [1:0] w_n24460_0;
	wire [1:0] w_n24461_0;
	wire [2:0] w_n24463_0;
	wire [1:0] w_n24464_0;
	wire [1:0] w_n24468_0;
	wire [1:0] w_n24469_0;
	wire [2:0] w_n24471_0;
	wire [1:0] w_n24472_0;
	wire [1:0] w_n24476_0;
	wire [1:0] w_n24477_0;
	wire [2:0] w_n24479_0;
	wire [1:0] w_n24480_0;
	wire [1:0] w_n24484_0;
	wire [1:0] w_n24485_0;
	wire [2:0] w_n24487_0;
	wire [1:0] w_n24488_0;
	wire [1:0] w_n24492_0;
	wire [1:0] w_n24493_0;
	wire [2:0] w_n24495_0;
	wire [1:0] w_n24496_0;
	wire [2:0] w_n24500_0;
	wire [2:0] w_n24502_0;
	wire [1:0] w_n24503_0;
	wire [1:0] w_n24507_0;
	wire [1:0] w_n24508_0;
	wire [2:0] w_n24510_0;
	wire [1:0] w_n24511_0;
	wire [2:0] w_n24515_0;
	wire [2:0] w_n24517_0;
	wire [1:0] w_n24518_0;
	wire [1:0] w_n24522_0;
	wire [1:0] w_n24523_0;
	wire [2:0] w_n24525_0;
	wire [1:0] w_n24526_0;
	wire [2:0] w_n24530_0;
	wire [2:0] w_n24532_0;
	wire [1:0] w_n24533_0;
	wire [2:0] w_n24537_0;
	wire [2:0] w_n24539_0;
	wire [1:0] w_n24540_0;
	wire [2:0] w_n24544_0;
	wire [2:0] w_n24546_0;
	wire [1:0] w_n24547_0;
	wire [1:0] w_n24551_0;
	wire [1:0] w_n24552_0;
	wire [2:0] w_n24554_0;
	wire [1:0] w_n24555_0;
	wire [1:0] w_n24830_0;
	wire [1:0] w_n24831_0;
	wire [1:0] w_n24834_0;
	wire [2:0] w_n24835_0;
	wire [1:0] w_n24836_0;
	wire [1:0] w_n24839_0;
	wire [1:0] w_n24845_0;
	wire [1:0] w_n24852_0;
	wire [2:0] w_n24856_0;
	wire [2:0] w_n24856_1;
	wire [2:0] w_n24856_2;
	wire [2:0] w_n24856_3;
	wire [2:0] w_n24856_4;
	wire [2:0] w_n24856_5;
	wire [2:0] w_n24856_6;
	wire [2:0] w_n24856_7;
	wire [2:0] w_n24856_8;
	wire [2:0] w_n24856_9;
	wire [2:0] w_n24856_10;
	wire [2:0] w_n24856_11;
	wire [2:0] w_n24856_12;
	wire [2:0] w_n24856_13;
	wire [2:0] w_n24856_14;
	wire [2:0] w_n24856_15;
	wire [2:0] w_n24856_16;
	wire [2:0] w_n24856_17;
	wire [2:0] w_n24856_18;
	wire [2:0] w_n24856_19;
	wire [2:0] w_n24856_20;
	wire [2:0] w_n24856_21;
	wire [2:0] w_n24856_22;
	wire [2:0] w_n24856_23;
	wire [2:0] w_n24856_24;
	wire [2:0] w_n24856_25;
	wire [2:0] w_n24856_26;
	wire [2:0] w_n24856_27;
	wire [2:0] w_n24856_28;
	wire [2:0] w_n24856_29;
	wire [2:0] w_n24856_30;
	wire [1:0] w_n24859_0;
	wire [1:0] w_n24863_0;
	wire [1:0] w_n24867_0;
	wire [1:0] w_n24873_0;
	wire [1:0] w_n24877_0;
	wire [1:0] w_n24881_0;
	wire [1:0] w_n24885_0;
	wire [1:0] w_n24889_0;
	wire [1:0] w_n24893_0;
	wire [1:0] w_n24897_0;
	wire [1:0] w_n24901_0;
	wire [1:0] w_n24905_0;
	wire [1:0] w_n24909_0;
	wire [1:0] w_n24913_0;
	wire [1:0] w_n24917_0;
	wire [1:0] w_n24921_0;
	wire [1:0] w_n24925_0;
	wire [1:0] w_n24929_0;
	wire [1:0] w_n24933_0;
	wire [1:0] w_n24937_0;
	wire [1:0] w_n24941_0;
	wire [1:0] w_n24945_0;
	wire [1:0] w_n24949_0;
	wire [1:0] w_n24953_0;
	wire [1:0] w_n24958_0;
	wire [1:0] w_n24962_0;
	wire [1:0] w_n24966_0;
	wire [1:0] w_n24968_0;
	wire [1:0] w_n24971_0;
	wire [1:0] w_n24977_0;
	wire [1:0] w_n24988_0;
	wire [1:0] w_n24995_0;
	wire [1:0] w_n25014_0;
	wire [1:0] w_n25021_0;
	wire [1:0] w_n25037_0;
	wire [1:0] w_n25050_0;
	wire [1:0] w_n25057_0;
	wire [1:0] w_n25070_0;
	wire [1:0] w_n25083_0;
	wire [1:0] w_n25090_0;
	wire [1:0] w_n25097_0;
	wire [1:0] w_n25113_0;
	wire [1:0] w_n25119_0;
	wire [1:0] w_n25130_0;
	wire [1:0] w_n25137_0;
	wire [1:0] w_n25143_0;
	wire [1:0] w_n25151_0;
	wire [1:0] w_n25164_0;
	wire [1:0] w_n25171_0;
	wire [1:0] w_n25178_0;
	wire [1:0] w_n25189_0;
	wire [1:0] w_n25195_0;
	wire [1:0] w_n25208_0;
	wire [1:0] w_n25215_0;
	wire [1:0] w_n25222_0;
	wire [1:0] w_n25235_0;
	wire [1:0] w_n25246_0;
	wire [1:0] w_n25253_0;
	wire [1:0] w_n25260_0;
	wire [1:0] w_n25267_0;
	wire [1:0] w_n25273_0;
	wire [1:0] w_n25281_0;
	wire [1:0] w_n25292_0;
	jand g00000(.dina(w_a127_0[1]),.dinb(w_a126_1[1]),.dout(n192),.clk(gclk));
	jnot g00001(.din(w_a126_1[0]),.dout(n193),.clk(gclk));
	jor g00002(.dina(w_a125_0[2]),.dinb(w_a124_1[1]),.dout(n194),.clk(gclk));
	jand g00003(.dina(n194),.dinb(w_n193_0[1]),.dout(n195),.clk(gclk));
	jor g00004(.dina(w_n195_0[1]),.dinb(w_n192_0[2]),.dout(asqrt_fa_63),.clk(gclk));
	jnot g00005(.din(w_a127_0[0]),.dout(n197),.clk(gclk));
	jnot g00006(.din(w_a124_1[0]),.dout(n198),.clk(gclk));
	jnot g00007(.din(w_a125_0[1]),.dout(n199),.clk(gclk));
	jand g00008(.dina(w_n199_0[1]),.dinb(w_n198_1[1]),.dout(n200),.clk(gclk));
	jand g00009(.dina(w_n200_0[2]),.dinb(w_a126_0[2]),.dout(n201),.clk(gclk));
	jor g00010(.dina(n201),.dinb(w_n197_0[1]),.dout(n202),.clk(gclk));
	jor g00011(.dina(n202),.dinb(w_n195_0[0]),.dout(n203),.clk(gclk));
	jnot g00012(.din(w_n203_0[1]),.dout(n204),.clk(gclk));
	jand g00013(.dina(w_asqrt62_45[1]),.dinb(w_n198_1[0]),.dout(n205),.clk(gclk));
	jor g00014(.dina(n205),.dinb(w_n199_0[0]),.dout(n206),.clk(gclk));
	jand g00015(.dina(w_n200_0[1]),.dinb(w_n192_0[1]),.dout(n207),.clk(gclk));
	jnot g00016(.din(w_n207_0[1]),.dout(n208),.clk(gclk));
	jand g00017(.dina(n208),.dinb(n206),.dout(n209),.clk(gclk));
	jand g00018(.dina(w_asqrt62_45[0]),.dinb(w_a124_0[2]),.dout(n210),.clk(gclk));
	jnot g00019(.din(w_a122_0[2]),.dout(n211),.clk(gclk));
	jnot g00020(.din(w_a123_0[1]),.dout(n212),.clk(gclk));
	jand g00021(.dina(w_n198_0[2]),.dinb(w_n212_0[1]),.dout(n213),.clk(gclk));
	jand g00022(.dina(n213),.dinb(w_n211_1[1]),.dout(n214),.clk(gclk));
	jor g00023(.dina(n214),.dinb(n210),.dout(n215),.clk(gclk));
	jor g00024(.dina(w_n215_0[2]),.dinb(w_n209_0[1]),.dout(n216),.clk(gclk));
	jnot g00025(.din(w_n216_1[1]),.dout(n217),.clk(gclk));
	jand g00026(.dina(w_n197_0[0]),.dinb(w_n193_0[0]),.dout(n218),.clk(gclk));
	jnot g00027(.din(w_n192_0[0]),.dout(n219),.clk(gclk));
	jor g00028(.dina(w_n200_0[0]),.dinb(w_a126_0[1]),.dout(n220),.clk(gclk));
	jand g00029(.dina(n220),.dinb(n219),.dout(n221),.clk(gclk));
	jor g00030(.dina(w_n221_76[1]),.dinb(w_a124_0[1]),.dout(n222),.clk(gclk));
	jand g00031(.dina(n222),.dinb(w_a125_0[0]),.dout(n223),.clk(gclk));
	jor g00032(.dina(w_n207_0[0]),.dinb(n223),.dout(n224),.clk(gclk));
	jnot g00033(.din(w_n215_0[1]),.dout(n225),.clk(gclk));
	jor g00034(.dina(w_n225_0[1]),.dinb(w_n224_0[1]),.dout(n226),.clk(gclk));
	jand g00035(.dina(n226),.dinb(w_n218_31[1]),.dout(n227),.clk(gclk));
	jor g00036(.dina(n227),.dinb(w_n217_0[1]),.dout(n228),.clk(gclk));
	jor g00037(.dina(n228),.dinb(w_n204_0[2]),.dout(asqrt_fa_62),.clk(gclk));
	jnot g00038(.din(w_n218_31[0]),.dout(asqrt[63]),.clk(gclk));
	jand g00039(.dina(w_n225_0[0]),.dinb(w_n204_0[1]),.dout(n231),.clk(gclk));
	jor g00040(.dina(n231),.dinb(w_n224_0[0]),.dout(n232),.clk(gclk));
	jand g00041(.dina(n232),.dinb(w_asqrt63_57),.dout(n233),.clk(gclk));
	jand g00042(.dina(n233),.dinb(w_n216_1[0]),.dout(n234),.clk(gclk));
	jand g00043(.dina(w_n215_0[0]),.dinb(w_n209_0[0]),.dout(n235),.clk(gclk));
	jand g00044(.dina(w_n235_0[1]),.dinb(w_n204_0[0]),.dout(n236),.clk(gclk));
	jor g00045(.dina(w_n235_0[0]),.dinb(w_asqrt63_56[2]),.dout(n237),.clk(gclk));
	jand g00046(.dina(n237),.dinb(w_n216_0[2]),.dout(n238),.clk(gclk));
	jand g00047(.dina(n238),.dinb(w_n203_0[0]),.dout(n239),.clk(gclk));
	jor g00048(.dina(w_n239_75[1]),.dinb(w_n211_1[0]),.dout(n240),.clk(gclk));
	jnot g00049(.din(w_a120_0[2]),.dout(n241),.clk(gclk));
	jnot g00050(.din(w_a121_0[1]),.dout(n242),.clk(gclk));
	jand g00051(.dina(w_n242_0[1]),.dinb(w_n241_1[2]),.dout(n243),.clk(gclk));
	jand g00052(.dina(w_n243_0[2]),.dinb(w_n211_0[2]),.dout(n244),.clk(gclk));
	jnot g00053(.din(w_n244_0[1]),.dout(n245),.clk(gclk));
	jand g00054(.dina(n245),.dinb(n240),.dout(n246),.clk(gclk));
	jor g00055(.dina(w_n246_0[2]),.dinb(w_n221_76[0]),.dout(n247),.clk(gclk));
	jand g00056(.dina(w_n246_0[1]),.dinb(w_n221_75[2]),.dout(n248),.clk(gclk));
	jor g00057(.dina(w_n239_75[0]),.dinb(w_a122_0[1]),.dout(n249),.clk(gclk));
	jxor g00058(.dina(w_n249_0[1]),.dinb(w_n212_0[0]),.dout(n250),.clk(gclk));
	jor g00059(.dina(w_n250_0[1]),.dinb(n248),.dout(n251),.clk(gclk));
	jand g00060(.dina(n251),.dinb(w_n247_0[1]),.dout(n252),.clk(gclk));
	jor g00061(.dina(w_n249_0[0]),.dinb(w_a123_0[0]),.dout(n253),.clk(gclk));
	jor g00062(.dina(w_asqrt61_45),.dinb(w_n221_75[1]),.dout(n254),.clk(gclk));
	jand g00063(.dina(n254),.dinb(n253),.dout(n255),.clk(gclk));
	jxor g00064(.dina(n255),.dinb(w_n198_0[1]),.dout(n256),.clk(gclk));
	jor g00065(.dina(w_n256_1[1]),.dinb(w_n252_0[2]),.dout(n257),.clk(gclk));
	jor g00066(.dina(n257),.dinb(w_n217_0[0]),.dout(n258),.clk(gclk));
	jor g00067(.dina(n258),.dinb(w_n236_0[1]),.dout(n259),.clk(gclk));
	jand g00068(.dina(n259),.dinb(w_n218_30[2]),.dout(n260),.clk(gclk));
	jand g00069(.dina(w_n256_1[0]),.dinb(w_n252_0[1]),.dout(n261),.clk(gclk));
	jor g00070(.dina(w_n261_0[1]),.dinb(w_n260_0[1]),.dout(n262),.clk(gclk));
	jor g00071(.dina(n262),.dinb(w_n234_0[1]),.dout(asqrt_fa_61),.clk(gclk));
	jnot g00072(.din(w_n250_0[0]),.dout(n264),.clk(gclk));
	jxor g00073(.dina(w_n246_0[0]),.dinb(w_n221_75[0]),.dout(n265),.clk(gclk));
	jand g00074(.dina(n265),.dinb(w_asqrt60_45[1]),.dout(n266),.clk(gclk));
	jxor g00075(.dina(n266),.dinb(w_n264_0[1]),.dout(n267),.clk(gclk));
	jnot g00076(.din(w_a118_1[1]),.dout(n268),.clk(gclk));
	jnot g00077(.din(w_a119_0[1]),.dout(n269),.clk(gclk));
	jand g00078(.dina(w_n269_0[1]),.dinb(w_n268_1[1]),.dout(n270),.clk(gclk));
	jand g00079(.dina(w_n270_0[2]),.dinb(w_n241_1[1]),.dout(n271),.clk(gclk));
	jand g00080(.dina(w_asqrt60_45[0]),.dinb(w_a120_0[1]),.dout(n272),.clk(gclk));
	jor g00081(.dina(n272),.dinb(w_n271_0[1]),.dout(n273),.clk(gclk));
	jand g00082(.dina(w_n273_0[2]),.dinb(w_asqrt61_44[2]),.dout(n274),.clk(gclk));
	jor g00083(.dina(w_n273_0[1]),.dinb(w_asqrt61_44[1]),.dout(n275),.clk(gclk));
	jand g00084(.dina(w_asqrt60_44[2]),.dinb(w_n241_1[0]),.dout(n276),.clk(gclk));
	jor g00085(.dina(n276),.dinb(w_n242_0[0]),.dout(n277),.clk(gclk));
	jnot g00086(.din(w_n243_0[1]),.dout(n278),.clk(gclk));
	jnot g00087(.din(w_n234_0[0]),.dout(n279),.clk(gclk));
	jnot g00088(.din(w_n236_0[0]),.dout(n280),.clk(gclk));
	jnot g00089(.din(w_n247_0[0]),.dout(n281),.clk(gclk));
	jand g00090(.dina(w_asqrt61_44[0]),.dinb(w_a122_0[0]),.dout(n282),.clk(gclk));
	jor g00091(.dina(w_n244_0[0]),.dinb(n282),.dout(n283),.clk(gclk));
	jor g00092(.dina(n283),.dinb(w_asqrt62_44[2]),.dout(n284),.clk(gclk));
	jand g00093(.dina(w_n264_0[0]),.dinb(n284),.dout(n285),.clk(gclk));
	jor g00094(.dina(n285),.dinb(n281),.dout(n286),.clk(gclk));
	jnot g00095(.din(w_n256_0[2]),.dout(n287),.clk(gclk));
	jand g00096(.dina(w_n287_0[1]),.dinb(n286),.dout(n288),.clk(gclk));
	jand g00097(.dina(n288),.dinb(w_n216_0[1]),.dout(n289),.clk(gclk));
	jand g00098(.dina(n289),.dinb(n280),.dout(n290),.clk(gclk));
	jor g00099(.dina(n290),.dinb(w_asqrt63_56[1]),.dout(n291),.clk(gclk));
	jnot g00100(.din(w_n261_0[0]),.dout(n292),.clk(gclk));
	jand g00101(.dina(n292),.dinb(n291),.dout(n293),.clk(gclk));
	jand g00102(.dina(n293),.dinb(n279),.dout(n294),.clk(gclk));
	jor g00103(.dina(w_n294_75[1]),.dinb(n278),.dout(n295),.clk(gclk));
	jand g00104(.dina(w_n295_0[1]),.dinb(n277),.dout(n296),.clk(gclk));
	jand g00105(.dina(n296),.dinb(n275),.dout(n297),.clk(gclk));
	jor g00106(.dina(n297),.dinb(w_n274_0[1]),.dout(n298),.clk(gclk));
	jand g00107(.dina(w_n298_0[2]),.dinb(w_asqrt62_44[1]),.dout(n299),.clk(gclk));
	jor g00108(.dina(w_n298_0[1]),.dinb(w_asqrt62_44[0]),.dout(n300),.clk(gclk));
	jor g00109(.dina(w_asqrt60_44[1]),.dinb(w_n239_74[2]),.dout(n301),.clk(gclk));
	jand g00110(.dina(n301),.dinb(w_n295_0[0]),.dout(n302),.clk(gclk));
	jxor g00111(.dina(n302),.dinb(w_n211_0[1]),.dout(n303),.clk(gclk));
	jnot g00112(.din(w_n303_0[1]),.dout(n304),.clk(gclk));
	jand g00113(.dina(w_n304_0[1]),.dinb(n300),.dout(n305),.clk(gclk));
	jor g00114(.dina(n305),.dinb(w_n299_0[1]),.dout(n306),.clk(gclk));
	jor g00115(.dina(w_n306_0[1]),.dinb(w_n267_1[1]),.dout(n307),.clk(gclk));
	jand g00116(.dina(w_n307_0[1]),.dinb(w_asqrt63_56[0]),.dout(n308),.clk(gclk));
	jnot g00117(.din(w_n308_0[1]),.dout(n309),.clk(gclk));
	jnot g00118(.din(w_n307_0[0]),.dout(n310),.clk(gclk));
	jnot g00119(.din(w_n267_1[0]),.dout(n311),.clk(gclk));
	jnot g00120(.din(w_n299_0[0]),.dout(n312),.clk(gclk));
	jnot g00121(.din(w_n274_0[0]),.dout(n313),.clk(gclk));
	jnot g00122(.din(w_n271_0[0]),.dout(n314),.clk(gclk));
	jor g00123(.dina(w_n294_75[0]),.dinb(w_n241_0[2]),.dout(n315),.clk(gclk));
	jand g00124(.dina(n315),.dinb(n314),.dout(n316),.clk(gclk));
	jand g00125(.dina(n316),.dinb(w_n239_74[1]),.dout(n317),.clk(gclk));
	jor g00126(.dina(w_n294_74[2]),.dinb(w_a120_0[0]),.dout(n318),.clk(gclk));
	jand g00127(.dina(n318),.dinb(w_a121_0[0]),.dout(n319),.clk(gclk));
	jand g00128(.dina(w_asqrt60_44[0]),.dinb(w_n243_0[0]),.dout(n320),.clk(gclk));
	jor g00129(.dina(n320),.dinb(n319),.dout(n321),.clk(gclk));
	jor g00130(.dina(w_n321_0[1]),.dinb(n317),.dout(n322),.clk(gclk));
	jand g00131(.dina(n322),.dinb(n313),.dout(n323),.clk(gclk));
	jand g00132(.dina(n323),.dinb(w_n221_74[2]),.dout(n324),.clk(gclk));
	jor g00133(.dina(w_n303_0[0]),.dinb(n324),.dout(n325),.clk(gclk));
	jand g00134(.dina(n325),.dinb(n312),.dout(n326),.clk(gclk));
	jor g00135(.dina(n326),.dinb(n311),.dout(n327),.clk(gclk));
	jxor g00136(.dina(w_n256_0[1]),.dinb(w_n252_0[0]),.dout(n328),.clk(gclk));
	jor g00137(.dina(n328),.dinb(w_n294_74[1]),.dout(n329),.clk(gclk));
	jnot g00138(.din(w_n329_0[1]),.dout(n330),.clk(gclk));
	jor g00139(.dina(w_n330_0[1]),.dinb(n327),.dout(n331),.clk(gclk));
	jand g00140(.dina(n331),.dinb(n309),.dout(n333),.clk(gclk));
	jor g00141(.dina(w_n260_0[0]),.dinb(w_n330_0[0]),.dout(n335),.clk(gclk));
	jnot g00142(.din(w_n335_0[1]),.dout(n336),.clk(gclk));
	jor g00143(.dina(n336),.dinb(w_n333_0[2]),.dout(n337),.clk(gclk));
	jand g00144(.dina(w_n294_74[0]),.dinb(w_n287_0[0]),.dout(n338),.clk(gclk));
	jnot g00145(.din(w_n338_0[1]),.dout(n339),.clk(gclk));
	jor g00146(.dina(n339),.dinb(w_n333_0[1]),.dout(n340),.clk(gclk));
	jand g00147(.dina(n340),.dinb(w_n337_0[1]),.dout(asqrt_fa_60),.clk(gclk));
	jand g00148(.dina(w_n306_0[0]),.dinb(w_n267_0[2]),.dout(n342),.clk(gclk));
	jand g00149(.dina(w_asqrt59_44[1]),.dinb(w_n342_0[1]),.dout(n343),.clk(gclk));
	jor g00150(.dina(w_n333_0[0]),.dinb(w_n343_0[1]),.dout(n345),.clk(gclk));
	jnot g00151(.din(w_n345_0[1]),.dout(n346),.clk(gclk));
	jand g00152(.dina(w_n329_0[0]),.dinb(w_n342_0[0]),.dout(n347),.clk(gclk));
	jor g00153(.dina(n347),.dinb(w_n308_0[0]),.dout(n349),.clk(gclk));
	jand g00154(.dina(w_n335_0[0]),.dinb(w_n349_0[1]),.dout(n350),.clk(gclk));
	jand g00155(.dina(w_n338_0[0]),.dinb(w_n349_0[0]),.dout(n351),.clk(gclk));
	jor g00156(.dina(n351),.dinb(n350),.dout(n352),.clk(gclk));
	jor g00157(.dina(w_n352_74[1]),.dinb(w_n268_1[0]),.dout(n353),.clk(gclk));
	jnot g00158(.din(w_a116_0[2]),.dout(n354),.clk(gclk));
	jnot g00159(.din(w_a117_0[1]),.dout(n355),.clk(gclk));
	jand g00160(.dina(w_n355_0[1]),.dinb(w_n354_1[2]),.dout(n356),.clk(gclk));
	jand g00161(.dina(w_n356_0[2]),.dinb(w_n268_0[2]),.dout(n357),.clk(gclk));
	jnot g00162(.din(w_n357_0[1]),.dout(n358),.clk(gclk));
	jand g00163(.dina(n358),.dinb(n353),.dout(n359),.clk(gclk));
	jor g00164(.dina(w_n359_0[2]),.dinb(w_n294_73[2]),.dout(n360),.clk(gclk));
	jand g00165(.dina(w_n359_0[1]),.dinb(w_n294_73[1]),.dout(n361),.clk(gclk));
	jor g00166(.dina(w_n352_74[0]),.dinb(w_a118_1[0]),.dout(n362),.clk(gclk));
	jand g00167(.dina(n362),.dinb(w_a119_0[0]),.dout(n363),.clk(gclk));
	jand g00168(.dina(w_asqrt59_44[0]),.dinb(w_n270_0[1]),.dout(n364),.clk(gclk));
	jor g00169(.dina(n364),.dinb(n363),.dout(n365),.clk(gclk));
	jor g00170(.dina(n365),.dinb(n361),.dout(n366),.clk(gclk));
	jand g00171(.dina(n366),.dinb(w_n360_0[1]),.dout(n367),.clk(gclk));
	jor g00172(.dina(w_n367_0[2]),.dinb(w_n239_74[0]),.dout(n368),.clk(gclk));
	jand g00173(.dina(w_n367_0[1]),.dinb(w_n239_73[2]),.dout(n369),.clk(gclk));
	jnot g00174(.din(w_n270_0[0]),.dout(n370),.clk(gclk));
	jor g00175(.dina(w_n352_73[2]),.dinb(n370),.dout(n371),.clk(gclk));
	jand g00176(.dina(w_n371_0[1]),.dinb(w_n337_0[0]),.dout(n372),.clk(gclk));
	jxor g00177(.dina(n372),.dinb(w_n241_0[1]),.dout(n373),.clk(gclk));
	jor g00178(.dina(w_n373_0[2]),.dinb(n369),.dout(n374),.clk(gclk));
	jand g00179(.dina(n374),.dinb(w_n368_0[1]),.dout(n375),.clk(gclk));
	jor g00180(.dina(w_n375_0[2]),.dinb(w_n221_74[1]),.dout(n376),.clk(gclk));
	jand g00181(.dina(w_n375_0[1]),.dinb(w_n221_74[0]),.dout(n377),.clk(gclk));
	jxor g00182(.dina(w_n273_0[0]),.dinb(w_n239_73[1]),.dout(n378),.clk(gclk));
	jor g00183(.dina(n378),.dinb(w_n352_73[1]),.dout(n379),.clk(gclk));
	jxor g00184(.dina(n379),.dinb(w_n321_0[0]),.dout(n380),.clk(gclk));
	jnot g00185(.din(w_n380_0[2]),.dout(n381),.clk(gclk));
	jor g00186(.dina(n381),.dinb(n377),.dout(n382),.clk(gclk));
	jand g00187(.dina(n382),.dinb(w_n376_0[1]),.dout(n383),.clk(gclk));
	jxor g00188(.dina(w_n298_0[0]),.dinb(w_n221_73[2]),.dout(n384),.clk(gclk));
	jor g00189(.dina(n384),.dinb(w_n352_73[0]),.dout(n385),.clk(gclk));
	jxor g00190(.dina(n385),.dinb(w_n304_0[0]),.dout(n386),.clk(gclk));
	jand g00191(.dina(w_n386_1[1]),.dinb(w_n383_0[2]),.dout(n387),.clk(gclk));
	jor g00192(.dina(w_n387_0[2]),.dinb(w_n218_30[1]),.dout(n388),.clk(gclk));
	jor g00193(.dina(w_n386_1[0]),.dinb(w_n383_0[1]),.dout(n389),.clk(gclk));
	jor g00194(.dina(w_n343_0[0]),.dinb(n310),.dout(n390),.clk(gclk));
	jor g00195(.dina(w_n390_0[1]),.dinb(w_n389_0[1]),.dout(n391),.clk(gclk));
	jand g00196(.dina(n391),.dinb(w_n388_0[1]),.dout(n393),.clk(gclk));
	jor g00197(.dina(w_n393_0[1]),.dinb(n346),.dout(n394),.clk(gclk));
	jand g00198(.dina(w_n352_72[2]),.dinb(w_n267_0[1]),.dout(n395),.clk(gclk));
	jnot g00199(.din(w_n395_0[1]),.dout(n396),.clk(gclk));
	jor g00200(.dina(n396),.dinb(w_n393_0[0]),.dout(n397),.clk(gclk));
	jand g00201(.dina(n397),.dinb(n394),.dout(asqrt_fa_59),.clk(gclk));
	jnot g00202(.din(w_n376_0[0]),.dout(n399),.clk(gclk));
	jnot g00203(.din(w_n368_0[0]),.dout(n400),.clk(gclk));
	jnot g00204(.din(w_n360_0[0]),.dout(n401),.clk(gclk));
	jand g00205(.dina(w_asqrt59_43[2]),.dinb(w_a118_0[2]),.dout(n402),.clk(gclk));
	jor g00206(.dina(w_n357_0[0]),.dinb(n402),.dout(n403),.clk(gclk));
	jor g00207(.dina(n403),.dinb(w_asqrt60_43[2]),.dout(n404),.clk(gclk));
	jand g00208(.dina(w_asqrt59_43[1]),.dinb(w_n268_0[1]),.dout(n405),.clk(gclk));
	jor g00209(.dina(n405),.dinb(w_n269_0[0]),.dout(n406),.clk(gclk));
	jand g00210(.dina(w_n371_0[0]),.dinb(n406),.dout(n407),.clk(gclk));
	jand g00211(.dina(w_n407_0[1]),.dinb(n404),.dout(n408),.clk(gclk));
	jor g00212(.dina(n408),.dinb(n401),.dout(n409),.clk(gclk));
	jor g00213(.dina(n409),.dinb(w_asqrt61_43[2]),.dout(n410),.clk(gclk));
	jnot g00214(.din(w_n373_0[1]),.dout(n411),.clk(gclk));
	jand g00215(.dina(n411),.dinb(n410),.dout(n412),.clk(gclk));
	jor g00216(.dina(n412),.dinb(n400),.dout(n413),.clk(gclk));
	jor g00217(.dina(n413),.dinb(w_asqrt62_43[2]),.dout(n414),.clk(gclk));
	jand g00218(.dina(w_n380_0[1]),.dinb(n414),.dout(n415),.clk(gclk));
	jor g00219(.dina(n415),.dinb(n399),.dout(n416),.clk(gclk));
	jnot g00220(.din(w_n386_0[2]),.dout(n417),.clk(gclk));
	jand g00221(.dina(n417),.dinb(n416),.dout(n418),.clk(gclk));
	jand g00222(.dina(w_asqrt58_45),.dinb(w_n418_0[1]),.dout(n419),.clk(gclk));
	jxor g00223(.dina(w_n375_0[0]),.dinb(w_n221_73[1]),.dout(n420),.clk(gclk));
	jand g00224(.dina(n420),.dinb(w_asqrt58_44[2]),.dout(n421),.clk(gclk));
	jxor g00225(.dina(n421),.dinb(w_n380_0[0]),.dout(n422),.clk(gclk));
	jnot g00226(.din(w_n422_0[2]),.dout(n423),.clk(gclk));
	jand g00227(.dina(w_asqrt58_44[1]),.dinb(w_a116_0[1]),.dout(n424),.clk(gclk));
	jnot g00228(.din(w_a114_1[1]),.dout(n425),.clk(gclk));
	jnot g00229(.din(w_a115_0[1]),.dout(n426),.clk(gclk));
	jand g00230(.dina(w_n426_0[1]),.dinb(w_n425_1[1]),.dout(n427),.clk(gclk));
	jand g00231(.dina(w_n427_0[2]),.dinb(w_n354_1[1]),.dout(n428),.clk(gclk));
	jor g00232(.dina(w_n428_0[1]),.dinb(n424),.dout(n429),.clk(gclk));
	jand g00233(.dina(w_n429_0[2]),.dinb(w_asqrt59_43[0]),.dout(n430),.clk(gclk));
	jor g00234(.dina(w_n429_0[1]),.dinb(w_asqrt59_42[2]),.dout(n431),.clk(gclk));
	jand g00235(.dina(w_asqrt58_44[0]),.dinb(w_n354_1[0]),.dout(n432),.clk(gclk));
	jor g00236(.dina(n432),.dinb(w_n355_0[0]),.dout(n433),.clk(gclk));
	jnot g00237(.din(w_n356_0[1]),.dout(n434),.clk(gclk));
	jnot g00238(.din(w_n388_0[0]),.dout(n435),.clk(gclk));
	jnot g00239(.din(w_n387_0[1]),.dout(n436),.clk(gclk));
	jnot g00240(.din(w_n390_0[0]),.dout(n437),.clk(gclk));
	jand g00241(.dina(n437),.dinb(w_n418_0[0]),.dout(n438),.clk(gclk));
	jor g00242(.dina(n438),.dinb(w_n435_0[1]),.dout(n440),.clk(gclk));
	jand g00243(.dina(w_n440_0[1]),.dinb(w_n345_0[0]),.dout(n441),.clk(gclk));
	jand g00244(.dina(w_n395_0[0]),.dinb(w_n440_0[0]),.dout(n442),.clk(gclk));
	jor g00245(.dina(n442),.dinb(w_n441_0[1]),.dout(n443),.clk(gclk));
	jor g00246(.dina(w_n443_73[1]),.dinb(n434),.dout(n444),.clk(gclk));
	jand g00247(.dina(n444),.dinb(n433),.dout(n445),.clk(gclk));
	jand g00248(.dina(n445),.dinb(n431),.dout(n446),.clk(gclk));
	jor g00249(.dina(n446),.dinb(w_n430_0[1]),.dout(n447),.clk(gclk));
	jand g00250(.dina(w_n447_0[2]),.dinb(w_asqrt60_43[1]),.dout(n448),.clk(gclk));
	jor g00251(.dina(w_n447_0[1]),.dinb(w_asqrt60_43[0]),.dout(n449),.clk(gclk));
	jand g00252(.dina(w_asqrt58_43[2]),.dinb(w_n356_0[0]),.dout(n450),.clk(gclk));
	jor g00253(.dina(w_n450_0[1]),.dinb(w_n441_0[0]),.dout(n451),.clk(gclk));
	jxor g00254(.dina(n451),.dinb(w_a118_0[1]),.dout(n452),.clk(gclk));
	jnot g00255(.din(w_n452_0[1]),.dout(n453),.clk(gclk));
	jand g00256(.dina(w_n453_0[1]),.dinb(n449),.dout(n454),.clk(gclk));
	jor g00257(.dina(n454),.dinb(w_n448_0[1]),.dout(n455),.clk(gclk));
	jand g00258(.dina(w_n455_0[2]),.dinb(w_asqrt61_43[1]),.dout(n456),.clk(gclk));
	jor g00259(.dina(w_n455_0[1]),.dinb(w_asqrt61_43[0]),.dout(n457),.clk(gclk));
	jxor g00260(.dina(w_n359_0[0]),.dinb(w_n294_73[0]),.dout(n458),.clk(gclk));
	jand g00261(.dina(n458),.dinb(w_asqrt58_43[1]),.dout(n459),.clk(gclk));
	jxor g00262(.dina(n459),.dinb(w_n407_0[0]),.dout(n460),.clk(gclk));
	jand g00263(.dina(w_n460_0[1]),.dinb(n457),.dout(n461),.clk(gclk));
	jor g00264(.dina(n461),.dinb(w_n456_0[1]),.dout(n462),.clk(gclk));
	jand g00265(.dina(w_n462_0[2]),.dinb(w_asqrt62_43[1]),.dout(n463),.clk(gclk));
	jnot g00266(.din(w_n463_0[1]),.dout(n464),.clk(gclk));
	jnot g00267(.din(w_n456_0[0]),.dout(n465),.clk(gclk));
	jnot g00268(.din(w_n448_0[0]),.dout(n466),.clk(gclk));
	jnot g00269(.din(w_n430_0[0]),.dout(n467),.clk(gclk));
	jor g00270(.dina(w_n443_73[0]),.dinb(w_n354_0[2]),.dout(n468),.clk(gclk));
	jnot g00271(.din(w_n428_0[0]),.dout(n469),.clk(gclk));
	jand g00272(.dina(n469),.dinb(n468),.dout(n470),.clk(gclk));
	jand g00273(.dina(n470),.dinb(w_n352_72[1]),.dout(n471),.clk(gclk));
	jor g00274(.dina(w_n443_72[2]),.dinb(w_a116_0[0]),.dout(n472),.clk(gclk));
	jand g00275(.dina(n472),.dinb(w_a117_0[0]),.dout(n473),.clk(gclk));
	jor g00276(.dina(w_n450_0[0]),.dinb(n473),.dout(n474),.clk(gclk));
	jor g00277(.dina(w_n474_0[1]),.dinb(n471),.dout(n475),.clk(gclk));
	jand g00278(.dina(n475),.dinb(n467),.dout(n476),.clk(gclk));
	jand g00279(.dina(n476),.dinb(w_n294_72[2]),.dout(n477),.clk(gclk));
	jor g00280(.dina(w_n452_0[0]),.dinb(n477),.dout(n478),.clk(gclk));
	jand g00281(.dina(n478),.dinb(n466),.dout(n479),.clk(gclk));
	jand g00282(.dina(n479),.dinb(w_n239_73[0]),.dout(n480),.clk(gclk));
	jnot g00283(.din(w_n460_0[0]),.dout(n481),.clk(gclk));
	jor g00284(.dina(w_n481_0[1]),.dinb(n480),.dout(n482),.clk(gclk));
	jand g00285(.dina(n482),.dinb(n465),.dout(n483),.clk(gclk));
	jand g00286(.dina(n483),.dinb(w_n221_73[0]),.dout(n484),.clk(gclk));
	jxor g00287(.dina(w_n367_0[0]),.dinb(w_n239_72[2]),.dout(n485),.clk(gclk));
	jand g00288(.dina(n485),.dinb(w_asqrt58_43[0]),.dout(n486),.clk(gclk));
	jxor g00289(.dina(n486),.dinb(w_n373_0[0]),.dout(n487),.clk(gclk));
	jor g00290(.dina(w_n487_0[2]),.dinb(n484),.dout(n488),.clk(gclk));
	jand g00291(.dina(n488),.dinb(n464),.dout(n489),.clk(gclk));
	jor g00292(.dina(w_n489_0[1]),.dinb(w_n423_0[1]),.dout(n490),.clk(gclk));
	jor g00293(.dina(w_n490_0[1]),.dinb(w_n387_0[0]),.dout(n491),.clk(gclk));
	jor g00294(.dina(n491),.dinb(w_n419_0[1]),.dout(n492),.clk(gclk));
	jand g00295(.dina(n492),.dinb(w_n218_30[0]),.dout(n493),.clk(gclk));
	jand g00296(.dina(w_n443_72[1]),.dinb(w_n386_0[1]),.dout(n494),.clk(gclk));
	jnot g00297(.din(n494),.dout(n495),.clk(gclk));
	jor g00298(.dina(w_n462_0[1]),.dinb(w_asqrt62_43[0]),.dout(n496),.clk(gclk));
	jnot g00299(.din(w_n487_0[1]),.dout(n497),.clk(gclk));
	jand g00300(.dina(n497),.dinb(n496),.dout(n498),.clk(gclk));
	jor g00301(.dina(n498),.dinb(w_n463_0[0]),.dout(n499),.clk(gclk));
	jor g00302(.dina(w_n499_0[1]),.dinb(w_n422_0[1]),.dout(n500),.clk(gclk));
	jand g00303(.dina(w_n500_0[2]),.dinb(n495),.dout(n501),.clk(gclk));
	jand g00304(.dina(w_n443_72[0]),.dinb(w_n383_0[0]),.dout(n502),.clk(gclk));
	jnot g00305(.din(n502),.dout(n503),.clk(gclk));
	jand g00306(.dina(w_n389_0[0]),.dinb(w_n435_0[0]),.dout(n504),.clk(gclk));
	jand g00307(.dina(w_n504_0[1]),.dinb(n503),.dout(n505),.clk(gclk));
	jnot g00308(.din(n505),.dout(n506),.clk(gclk));
	jand g00309(.dina(n506),.dinb(n501),.dout(n507),.clk(gclk));
	jnot g00310(.din(w_n507_0[1]),.dout(n508),.clk(gclk));
	jor g00311(.dina(n508),.dinb(w_n493_0[1]),.dout(asqrt_fa_58),.clk(gclk));
	jnot g00312(.din(w_n419_0[0]),.dout(n510),.clk(gclk));
	jand g00313(.dina(w_n499_0[0]),.dinb(w_n422_0[0]),.dout(n511),.clk(gclk));
	jand g00314(.dina(w_n511_0[1]),.dinb(n436),.dout(n512),.clk(gclk));
	jand g00315(.dina(n512),.dinb(n510),.dout(n513),.clk(gclk));
	jor g00316(.dina(n513),.dinb(w_asqrt63_55[2]),.dout(n514),.clk(gclk));
	jand g00317(.dina(w_n507_0[0]),.dinb(n514),.dout(n515),.clk(gclk));
	jxor g00318(.dina(w_n462_0[0]),.dinb(w_n221_72[2]),.dout(n516),.clk(gclk));
	jor g00319(.dina(n516),.dinb(w_n515_73[1]),.dout(n517),.clk(gclk));
	jxor g00320(.dina(n517),.dinb(w_n487_0[0]),.dout(n518),.clk(gclk));
	jnot g00321(.din(w_n518_0[2]),.dout(n519),.clk(gclk));
	jor g00322(.dina(w_n515_73[0]),.dinb(w_n425_1[0]),.dout(n520),.clk(gclk));
	jnot g00323(.din(w_a112_0[2]),.dout(n521),.clk(gclk));
	jnot g00324(.din(w_a113_0[1]),.dout(n522),.clk(gclk));
	jand g00325(.dina(w_n522_0[1]),.dinb(w_n521_1[2]),.dout(n523),.clk(gclk));
	jand g00326(.dina(w_n523_0[2]),.dinb(w_n425_0[2]),.dout(n524),.clk(gclk));
	jnot g00327(.din(w_n524_0[1]),.dout(n525),.clk(gclk));
	jand g00328(.dina(n525),.dinb(n520),.dout(n526),.clk(gclk));
	jor g00329(.dina(w_n526_0[2]),.dinb(w_n443_71[2]),.dout(n527),.clk(gclk));
	jand g00330(.dina(w_n526_0[1]),.dinb(w_n443_71[1]),.dout(n528),.clk(gclk));
	jor g00331(.dina(w_n515_72[2]),.dinb(w_a114_1[0]),.dout(n529),.clk(gclk));
	jand g00332(.dina(n529),.dinb(w_a115_0[0]),.dout(n530),.clk(gclk));
	jand g00333(.dina(w_asqrt57_43[1]),.dinb(w_n427_0[1]),.dout(n531),.clk(gclk));
	jor g00334(.dina(n531),.dinb(n530),.dout(n532),.clk(gclk));
	jor g00335(.dina(n532),.dinb(n528),.dout(n533),.clk(gclk));
	jand g00336(.dina(n533),.dinb(w_n527_0[1]),.dout(n534),.clk(gclk));
	jor g00337(.dina(w_n534_0[2]),.dinb(w_n352_72[0]),.dout(n535),.clk(gclk));
	jand g00338(.dina(w_n534_0[1]),.dinb(w_n352_71[2]),.dout(n536),.clk(gclk));
	jnot g00339(.din(w_n427_0[0]),.dout(n537),.clk(gclk));
	jor g00340(.dina(w_n515_72[1]),.dinb(n537),.dout(n538),.clk(gclk));
	jnot g00341(.din(w_n500_0[1]),.dout(n539),.clk(gclk));
	jor g00342(.dina(w_n504_0[0]),.dinb(w_n443_71[0]),.dout(n540),.clk(gclk));
	jor g00343(.dina(n540),.dinb(w_n539_0[1]),.dout(n541),.clk(gclk));
	jor g00344(.dina(n541),.dinb(w_n493_0[0]),.dout(n542),.clk(gclk));
	jand g00345(.dina(n542),.dinb(w_n538_0[1]),.dout(n543),.clk(gclk));
	jxor g00346(.dina(n543),.dinb(w_n354_0[1]),.dout(n544),.clk(gclk));
	jor g00347(.dina(w_n544_0[2]),.dinb(n536),.dout(n545),.clk(gclk));
	jand g00348(.dina(n545),.dinb(w_n535_0[1]),.dout(n546),.clk(gclk));
	jor g00349(.dina(w_n546_0[2]),.dinb(w_n294_72[1]),.dout(n547),.clk(gclk));
	jand g00350(.dina(w_n546_0[1]),.dinb(w_n294_72[0]),.dout(n548),.clk(gclk));
	jxor g00351(.dina(w_n429_0[0]),.dinb(w_n352_71[1]),.dout(n549),.clk(gclk));
	jor g00352(.dina(n549),.dinb(w_n515_72[0]),.dout(n550),.clk(gclk));
	jxor g00353(.dina(n550),.dinb(w_n474_0[0]),.dout(n551),.clk(gclk));
	jnot g00354(.din(w_n551_0[2]),.dout(n552),.clk(gclk));
	jor g00355(.dina(n552),.dinb(n548),.dout(n553),.clk(gclk));
	jand g00356(.dina(n553),.dinb(w_n547_0[1]),.dout(n554),.clk(gclk));
	jor g00357(.dina(w_n554_0[2]),.dinb(w_n239_72[1]),.dout(n555),.clk(gclk));
	jand g00358(.dina(w_n554_0[1]),.dinb(w_n239_72[0]),.dout(n556),.clk(gclk));
	jxor g00359(.dina(w_n447_0[0]),.dinb(w_n294_71[2]),.dout(n557),.clk(gclk));
	jor g00360(.dina(n557),.dinb(w_n515_71[2]),.dout(n558),.clk(gclk));
	jxor g00361(.dina(n558),.dinb(w_n453_0[0]),.dout(n559),.clk(gclk));
	jor g00362(.dina(w_n559_0[2]),.dinb(n556),.dout(n560),.clk(gclk));
	jand g00363(.dina(n560),.dinb(w_n555_0[1]),.dout(n561),.clk(gclk));
	jor g00364(.dina(w_n561_0[2]),.dinb(w_n221_72[1]),.dout(n562),.clk(gclk));
	jand g00365(.dina(w_n561_0[1]),.dinb(w_n221_72[0]),.dout(n563),.clk(gclk));
	jxor g00366(.dina(w_n455_0[0]),.dinb(w_n239_71[2]),.dout(n564),.clk(gclk));
	jor g00367(.dina(n564),.dinb(w_n515_71[1]),.dout(n565),.clk(gclk));
	jxor g00368(.dina(n565),.dinb(w_n481_0[0]),.dout(n566),.clk(gclk));
	jnot g00369(.din(w_n566_0[2]),.dout(n567),.clk(gclk));
	jor g00370(.dina(n567),.dinb(n563),.dout(n568),.clk(gclk));
	jand g00371(.dina(n568),.dinb(w_n562_0[1]),.dout(n569),.clk(gclk));
	jor g00372(.dina(w_n569_0[2]),.dinb(w_n519_0[2]),.dout(n570),.clk(gclk));
	jand g00373(.dina(w_asqrt57_43[0]),.dinb(w_n511_0[0]),.dout(n571),.clk(gclk));
	jor g00374(.dina(n571),.dinb(w_n539_0[0]),.dout(n572),.clk(gclk));
	jor g00375(.dina(w_n572_0[1]),.dinb(w_n570_0[1]),.dout(n573),.clk(gclk));
	jand g00376(.dina(n573),.dinb(w_n218_29[2]),.dout(n574),.clk(gclk));
	jand g00377(.dina(w_n515_71[0]),.dinb(w_n423_0[0]),.dout(n575),.clk(gclk));
	jand g00378(.dina(w_n569_0[1]),.dinb(w_n519_0[1]),.dout(n576),.clk(gclk));
	jor g00379(.dina(w_n576_0[1]),.dinb(w_n575_0[1]),.dout(n577),.clk(gclk));
	jand g00380(.dina(w_n515_70[2]),.dinb(w_n489_0[0]),.dout(n578),.clk(gclk));
	jand g00381(.dina(w_n490_0[0]),.dinb(w_asqrt63_55[1]),.dout(n579),.clk(gclk));
	jand g00382(.dina(n579),.dinb(w_n500_0[0]),.dout(n580),.clk(gclk));
	jnot g00383(.din(n580),.dout(n581),.clk(gclk));
	jor g00384(.dina(w_n581_0[1]),.dinb(n578),.dout(n582),.clk(gclk));
	jnot g00385(.din(w_n582_0[1]),.dout(n583),.clk(gclk));
	jor g00386(.dina(n583),.dinb(n577),.dout(n584),.clk(gclk));
	jor g00387(.dina(n584),.dinb(n574),.dout(asqrt_fa_57),.clk(gclk));
	jxor g00388(.dina(w_n561_0[0]),.dinb(w_n221_71[2]),.dout(n586),.clk(gclk));
	jand g00389(.dina(n586),.dinb(w_asqrt56_44[1]),.dout(n587),.clk(gclk));
	jxor g00390(.dina(n587),.dinb(w_n566_0[1]),.dout(n588),.clk(gclk));
	jnot g00391(.din(w_a110_1[1]),.dout(n589),.clk(gclk));
	jnot g00392(.din(w_a111_0[1]),.dout(n590),.clk(gclk));
	jand g00393(.dina(w_n590_0[1]),.dinb(w_n589_1[1]),.dout(n591),.clk(gclk));
	jand g00394(.dina(w_n591_0[2]),.dinb(w_n521_1[1]),.dout(n592),.clk(gclk));
	jand g00395(.dina(w_asqrt56_44[0]),.dinb(w_a112_0[1]),.dout(n593),.clk(gclk));
	jor g00396(.dina(n593),.dinb(w_n592_0[1]),.dout(n594),.clk(gclk));
	jand g00397(.dina(w_n594_0[2]),.dinb(w_asqrt57_42[2]),.dout(n595),.clk(gclk));
	jor g00398(.dina(w_n594_0[1]),.dinb(w_asqrt57_42[1]),.dout(n596),.clk(gclk));
	jand g00399(.dina(w_asqrt56_43[2]),.dinb(w_n521_1[0]),.dout(n597),.clk(gclk));
	jor g00400(.dina(n597),.dinb(w_n522_0[0]),.dout(n598),.clk(gclk));
	jnot g00401(.din(w_n523_0[1]),.dout(n599),.clk(gclk));
	jnot g00402(.din(w_n562_0[0]),.dout(n600),.clk(gclk));
	jnot g00403(.din(w_n555_0[0]),.dout(n601),.clk(gclk));
	jnot g00404(.din(w_n547_0[0]),.dout(n602),.clk(gclk));
	jnot g00405(.din(w_n535_0[0]),.dout(n603),.clk(gclk));
	jnot g00406(.din(w_n527_0[0]),.dout(n604),.clk(gclk));
	jand g00407(.dina(w_asqrt57_42[0]),.dinb(w_a114_0[2]),.dout(n605),.clk(gclk));
	jor g00408(.dina(w_n524_0[0]),.dinb(n605),.dout(n606),.clk(gclk));
	jor g00409(.dina(n606),.dinb(w_asqrt58_42[2]),.dout(n607),.clk(gclk));
	jand g00410(.dina(w_asqrt57_41[2]),.dinb(w_n425_0[1]),.dout(n608),.clk(gclk));
	jor g00411(.dina(n608),.dinb(w_n426_0[0]),.dout(n609),.clk(gclk));
	jand g00412(.dina(w_n538_0[0]),.dinb(n609),.dout(n610),.clk(gclk));
	jand g00413(.dina(w_n610_0[1]),.dinb(n607),.dout(n611),.clk(gclk));
	jor g00414(.dina(n611),.dinb(n604),.dout(n612),.clk(gclk));
	jor g00415(.dina(n612),.dinb(w_asqrt59_42[1]),.dout(n613),.clk(gclk));
	jnot g00416(.din(w_n544_0[1]),.dout(n614),.clk(gclk));
	jand g00417(.dina(n614),.dinb(n613),.dout(n615),.clk(gclk));
	jor g00418(.dina(n615),.dinb(n603),.dout(n616),.clk(gclk));
	jor g00419(.dina(n616),.dinb(w_asqrt60_42[2]),.dout(n617),.clk(gclk));
	jand g00420(.dina(w_n551_0[1]),.dinb(n617),.dout(n618),.clk(gclk));
	jor g00421(.dina(n618),.dinb(n602),.dout(n619),.clk(gclk));
	jor g00422(.dina(n619),.dinb(w_asqrt61_42[2]),.dout(n620),.clk(gclk));
	jnot g00423(.din(w_n559_0[1]),.dout(n621),.clk(gclk));
	jand g00424(.dina(n621),.dinb(n620),.dout(n622),.clk(gclk));
	jor g00425(.dina(n622),.dinb(n601),.dout(n623),.clk(gclk));
	jor g00426(.dina(n623),.dinb(w_asqrt62_42[2]),.dout(n624),.clk(gclk));
	jand g00427(.dina(w_n566_0[0]),.dinb(n624),.dout(n625),.clk(gclk));
	jor g00428(.dina(n625),.dinb(n600),.dout(n626),.clk(gclk));
	jand g00429(.dina(w_n626_0[1]),.dinb(w_n518_0[1]),.dout(n627),.clk(gclk));
	jnot g00430(.din(w_n572_0[0]),.dout(n628),.clk(gclk));
	jand g00431(.dina(n628),.dinb(w_n627_0[1]),.dout(n629),.clk(gclk));
	jor g00432(.dina(n629),.dinb(w_asqrt63_55[0]),.dout(n630),.clk(gclk));
	jnot g00433(.din(w_n575_0[0]),.dout(n631),.clk(gclk));
	jor g00434(.dina(w_n626_0[0]),.dinb(w_n518_0[0]),.dout(n632),.clk(gclk));
	jand g00435(.dina(w_n632_0[2]),.dinb(n631),.dout(n633),.clk(gclk));
	jand g00436(.dina(w_n582_0[0]),.dinb(n633),.dout(n634),.clk(gclk));
	jand g00437(.dina(n634),.dinb(w_n630_0[1]),.dout(n635),.clk(gclk));
	jor g00438(.dina(w_n635_70[2]),.dinb(n599),.dout(n636),.clk(gclk));
	jand g00439(.dina(n636),.dinb(n598),.dout(n637),.clk(gclk));
	jand g00440(.dina(n637),.dinb(n596),.dout(n638),.clk(gclk));
	jor g00441(.dina(n638),.dinb(w_n595_0[1]),.dout(n639),.clk(gclk));
	jand g00442(.dina(w_n639_0[2]),.dinb(w_asqrt58_42[1]),.dout(n640),.clk(gclk));
	jor g00443(.dina(w_n639_0[1]),.dinb(w_asqrt58_42[0]),.dout(n641),.clk(gclk));
	jand g00444(.dina(w_asqrt56_43[1]),.dinb(w_n523_0[0]),.dout(n642),.clk(gclk));
	jand g00445(.dina(w_n581_0[0]),.dinb(w_asqrt57_41[1]),.dout(n643),.clk(gclk));
	jand g00446(.dina(n643),.dinb(w_n632_0[1]),.dout(n644),.clk(gclk));
	jand g00447(.dina(n644),.dinb(w_n630_0[0]),.dout(n645),.clk(gclk));
	jor g00448(.dina(n645),.dinb(w_n642_0[1]),.dout(n646),.clk(gclk));
	jxor g00449(.dina(n646),.dinb(w_a114_0[1]),.dout(n647),.clk(gclk));
	jnot g00450(.din(w_n647_0[1]),.dout(n648),.clk(gclk));
	jand g00451(.dina(w_n648_0[1]),.dinb(n641),.dout(n649),.clk(gclk));
	jor g00452(.dina(n649),.dinb(w_n640_0[1]),.dout(n650),.clk(gclk));
	jand g00453(.dina(w_n650_0[2]),.dinb(w_asqrt59_42[0]),.dout(n651),.clk(gclk));
	jor g00454(.dina(w_n650_0[1]),.dinb(w_asqrt59_41[2]),.dout(n652),.clk(gclk));
	jxor g00455(.dina(w_n526_0[0]),.dinb(w_n443_70[2]),.dout(n653),.clk(gclk));
	jand g00456(.dina(n653),.dinb(w_asqrt56_43[0]),.dout(n654),.clk(gclk));
	jxor g00457(.dina(n654),.dinb(w_n610_0[0]),.dout(n655),.clk(gclk));
	jand g00458(.dina(w_n655_0[1]),.dinb(n652),.dout(n656),.clk(gclk));
	jor g00459(.dina(n656),.dinb(w_n651_0[1]),.dout(n657),.clk(gclk));
	jand g00460(.dina(w_n657_0[2]),.dinb(w_asqrt60_42[1]),.dout(n658),.clk(gclk));
	jor g00461(.dina(w_n657_0[1]),.dinb(w_asqrt60_42[0]),.dout(n659),.clk(gclk));
	jxor g00462(.dina(w_n534_0[0]),.dinb(w_n352_71[0]),.dout(n660),.clk(gclk));
	jand g00463(.dina(n660),.dinb(w_asqrt56_42[2]),.dout(n661),.clk(gclk));
	jxor g00464(.dina(n661),.dinb(w_n544_0[0]),.dout(n662),.clk(gclk));
	jnot g00465(.din(w_n662_0[1]),.dout(n663),.clk(gclk));
	jand g00466(.dina(w_n663_0[1]),.dinb(n659),.dout(n664),.clk(gclk));
	jor g00467(.dina(n664),.dinb(w_n658_0[1]),.dout(n665),.clk(gclk));
	jand g00468(.dina(w_n665_0[2]),.dinb(w_asqrt61_42[1]),.dout(n666),.clk(gclk));
	jor g00469(.dina(w_n665_0[1]),.dinb(w_asqrt61_42[0]),.dout(n667),.clk(gclk));
	jxor g00470(.dina(w_n546_0[0]),.dinb(w_n294_71[1]),.dout(n668),.clk(gclk));
	jand g00471(.dina(n668),.dinb(w_asqrt56_42[1]),.dout(n669),.clk(gclk));
	jxor g00472(.dina(n669),.dinb(w_n551_0[0]),.dout(n670),.clk(gclk));
	jand g00473(.dina(w_n670_0[1]),.dinb(n667),.dout(n671),.clk(gclk));
	jor g00474(.dina(n671),.dinb(w_n666_0[1]),.dout(n672),.clk(gclk));
	jand g00475(.dina(w_n672_0[2]),.dinb(w_asqrt62_42[1]),.dout(n673),.clk(gclk));
	jor g00476(.dina(w_n672_0[1]),.dinb(w_asqrt62_42[0]),.dout(n674),.clk(gclk));
	jxor g00477(.dina(w_n554_0[0]),.dinb(w_n239_71[1]),.dout(n675),.clk(gclk));
	jand g00478(.dina(n675),.dinb(w_asqrt56_42[0]),.dout(n676),.clk(gclk));
	jxor g00479(.dina(n676),.dinb(w_n559_0[0]),.dout(n677),.clk(gclk));
	jnot g00480(.din(w_n677_0[1]),.dout(n678),.clk(gclk));
	jand g00481(.dina(w_n678_0[1]),.dinb(n674),.dout(n679),.clk(gclk));
	jor g00482(.dina(n679),.dinb(w_n673_0[1]),.dout(n680),.clk(gclk));
	jor g00483(.dina(w_n680_0[1]),.dinb(w_n588_0[2]),.dout(n681),.clk(gclk));
	jnot g00484(.din(w_n681_1[1]),.dout(n682),.clk(gclk));
	jand g00485(.dina(w_n635_70[1]),.dinb(w_n569_0[0]),.dout(n683),.clk(gclk));
	jnot g00486(.din(n683),.dout(n684),.clk(gclk));
	jand g00487(.dina(w_n570_0[0]),.dinb(w_asqrt63_54[2]),.dout(n685),.clk(gclk));
	jand g00488(.dina(n685),.dinb(w_n632_0[0]),.dout(n686),.clk(gclk));
	jand g00489(.dina(w_n686_0[1]),.dinb(n684),.dout(n687),.clk(gclk));
	jnot g00490(.din(w_n588_0[1]),.dout(n688),.clk(gclk));
	jnot g00491(.din(w_n673_0[0]),.dout(n689),.clk(gclk));
	jnot g00492(.din(w_n666_0[0]),.dout(n690),.clk(gclk));
	jnot g00493(.din(w_n658_0[0]),.dout(n691),.clk(gclk));
	jnot g00494(.din(w_n651_0[0]),.dout(n692),.clk(gclk));
	jnot g00495(.din(w_n640_0[0]),.dout(n693),.clk(gclk));
	jnot g00496(.din(w_n595_0[0]),.dout(n694),.clk(gclk));
	jnot g00497(.din(w_n592_0[0]),.dout(n695),.clk(gclk));
	jor g00498(.dina(w_n635_70[0]),.dinb(w_n521_0[2]),.dout(n696),.clk(gclk));
	jand g00499(.dina(n696),.dinb(n695),.dout(n697),.clk(gclk));
	jand g00500(.dina(n697),.dinb(w_n515_70[1]),.dout(n698),.clk(gclk));
	jor g00501(.dina(w_n635_69[2]),.dinb(w_a112_0[0]),.dout(n699),.clk(gclk));
	jand g00502(.dina(n699),.dinb(w_a113_0[0]),.dout(n700),.clk(gclk));
	jor g00503(.dina(w_n642_0[0]),.dinb(n700),.dout(n701),.clk(gclk));
	jor g00504(.dina(w_n701_0[1]),.dinb(n698),.dout(n702),.clk(gclk));
	jand g00505(.dina(n702),.dinb(n694),.dout(n703),.clk(gclk));
	jand g00506(.dina(n703),.dinb(w_n443_70[1]),.dout(n704),.clk(gclk));
	jor g00507(.dina(w_n647_0[0]),.dinb(n704),.dout(n705),.clk(gclk));
	jand g00508(.dina(n705),.dinb(n693),.dout(n706),.clk(gclk));
	jand g00509(.dina(n706),.dinb(w_n352_70[2]),.dout(n707),.clk(gclk));
	jnot g00510(.din(w_n655_0[0]),.dout(n708),.clk(gclk));
	jor g00511(.dina(w_n708_0[1]),.dinb(n707),.dout(n709),.clk(gclk));
	jand g00512(.dina(n709),.dinb(n692),.dout(n710),.clk(gclk));
	jand g00513(.dina(n710),.dinb(w_n294_71[0]),.dout(n711),.clk(gclk));
	jor g00514(.dina(w_n662_0[0]),.dinb(n711),.dout(n712),.clk(gclk));
	jand g00515(.dina(n712),.dinb(n691),.dout(n713),.clk(gclk));
	jand g00516(.dina(n713),.dinb(w_n239_71[0]),.dout(n714),.clk(gclk));
	jnot g00517(.din(w_n670_0[0]),.dout(n715),.clk(gclk));
	jor g00518(.dina(w_n715_0[1]),.dinb(n714),.dout(n716),.clk(gclk));
	jand g00519(.dina(n716),.dinb(n690),.dout(n717),.clk(gclk));
	jand g00520(.dina(n717),.dinb(w_n221_71[1]),.dout(n718),.clk(gclk));
	jor g00521(.dina(w_n677_0[0]),.dinb(n718),.dout(n719),.clk(gclk));
	jand g00522(.dina(n719),.dinb(n689),.dout(n720),.clk(gclk));
	jor g00523(.dina(w_n720_0[1]),.dinb(n688),.dout(n721),.clk(gclk));
	jand g00524(.dina(w_asqrt56_41[2]),.dinb(w_n627_0[0]),.dout(n722),.clk(gclk));
	jor g00525(.dina(n722),.dinb(w_n576_0[0]),.dout(n723),.clk(gclk));
	jor g00526(.dina(w_n723_0[1]),.dinb(w_n721_0[1]),.dout(n724),.clk(gclk));
	jand g00527(.dina(n724),.dinb(w_n218_29[1]),.dout(n725),.clk(gclk));
	jand g00528(.dina(w_n635_69[1]),.dinb(w_n519_0[0]),.dout(n726),.clk(gclk));
	jor g00529(.dina(w_n726_0[1]),.dinb(w_n725_0[1]),.dout(n727),.clk(gclk));
	jor g00530(.dina(n727),.dinb(w_n687_0[1]),.dout(n728),.clk(gclk));
	jor g00531(.dina(w_n728_0[1]),.dinb(w_n682_0[2]),.dout(asqrt_fa_56),.clk(gclk));
	jnot g00532(.din(w_a108_0[2]),.dout(n730),.clk(gclk));
	jnot g00533(.din(w_a109_0[1]),.dout(n731),.clk(gclk));
	jand g00534(.dina(w_n731_0[1]),.dinb(w_n730_1[2]),.dout(n732),.clk(gclk));
	jand g00535(.dina(w_n732_0[2]),.dinb(w_n589_1[0]),.dout(n733),.clk(gclk));
	jnot g00536(.din(w_n733_0[1]),.dout(n734),.clk(gclk));
	jnot g00537(.din(w_n687_0[0]),.dout(n735),.clk(gclk));
	jand g00538(.dina(w_n680_0[0]),.dinb(w_n588_0[0]),.dout(n736),.clk(gclk));
	jnot g00539(.din(w_n723_0[0]),.dout(n737),.clk(gclk));
	jand g00540(.dina(n737),.dinb(w_n736_0[1]),.dout(n738),.clk(gclk));
	jor g00541(.dina(n738),.dinb(w_asqrt63_54[1]),.dout(n739),.clk(gclk));
	jnot g00542(.din(w_n726_0[0]),.dout(n740),.clk(gclk));
	jand g00543(.dina(n740),.dinb(n739),.dout(n741),.clk(gclk));
	jand g00544(.dina(n741),.dinb(n735),.dout(n742),.clk(gclk));
	jand g00545(.dina(w_n742_0[1]),.dinb(w_n681_1[0]),.dout(n743),.clk(gclk));
	jor g00546(.dina(w_n743_70[2]),.dinb(w_n589_0[2]),.dout(n744),.clk(gclk));
	jand g00547(.dina(n744),.dinb(n734),.dout(n745),.clk(gclk));
	jor g00548(.dina(w_n745_0[2]),.dinb(w_n635_69[0]),.dout(n746),.clk(gclk));
	jand g00549(.dina(w_n745_0[1]),.dinb(w_n635_68[2]),.dout(n747),.clk(gclk));
	jor g00550(.dina(w_n743_70[1]),.dinb(w_a110_1[0]),.dout(n748),.clk(gclk));
	jand g00551(.dina(n748),.dinb(w_a111_0[0]),.dout(n749),.clk(gclk));
	jand g00552(.dina(w_asqrt55_41[1]),.dinb(w_n591_0[1]),.dout(n750),.clk(gclk));
	jor g00553(.dina(n750),.dinb(n749),.dout(n751),.clk(gclk));
	jor g00554(.dina(n751),.dinb(n747),.dout(n752),.clk(gclk));
	jand g00555(.dina(n752),.dinb(w_n746_0[1]),.dout(n753),.clk(gclk));
	jor g00556(.dina(w_n753_0[2]),.dinb(w_n515_70[0]),.dout(n754),.clk(gclk));
	jand g00557(.dina(w_n753_0[1]),.dinb(w_n515_69[2]),.dout(n755),.clk(gclk));
	jnot g00558(.din(w_n591_0[0]),.dout(n756),.clk(gclk));
	jor g00559(.dina(w_n743_70[0]),.dinb(n756),.dout(n757),.clk(gclk));
	jor g00560(.dina(w_n682_0[1]),.dinb(w_n635_68[1]),.dout(n758),.clk(gclk));
	jor g00561(.dina(n758),.dinb(w_n686_0[0]),.dout(n759),.clk(gclk));
	jor g00562(.dina(n759),.dinb(w_n725_0[0]),.dout(n760),.clk(gclk));
	jand g00563(.dina(n760),.dinb(w_n757_0[1]),.dout(n761),.clk(gclk));
	jxor g00564(.dina(n761),.dinb(w_n521_0[1]),.dout(n762),.clk(gclk));
	jor g00565(.dina(w_n762_0[1]),.dinb(n755),.dout(n763),.clk(gclk));
	jand g00566(.dina(n763),.dinb(w_n754_0[1]),.dout(n764),.clk(gclk));
	jor g00567(.dina(w_n764_0[2]),.dinb(w_n443_70[0]),.dout(n765),.clk(gclk));
	jand g00568(.dina(w_n764_0[1]),.dinb(w_n443_69[2]),.dout(n766),.clk(gclk));
	jxor g00569(.dina(w_n594_0[0]),.dinb(w_n515_69[1]),.dout(n767),.clk(gclk));
	jor g00570(.dina(n767),.dinb(w_n743_69[2]),.dout(n768),.clk(gclk));
	jxor g00571(.dina(n768),.dinb(w_n701_0[0]),.dout(n769),.clk(gclk));
	jnot g00572(.din(w_n769_0[2]),.dout(n770),.clk(gclk));
	jor g00573(.dina(n770),.dinb(n766),.dout(n771),.clk(gclk));
	jand g00574(.dina(n771),.dinb(w_n765_0[1]),.dout(n772),.clk(gclk));
	jor g00575(.dina(w_n772_0[2]),.dinb(w_n352_70[1]),.dout(n773),.clk(gclk));
	jand g00576(.dina(w_n772_0[1]),.dinb(w_n352_70[0]),.dout(n774),.clk(gclk));
	jxor g00577(.dina(w_n639_0[0]),.dinb(w_n443_69[1]),.dout(n775),.clk(gclk));
	jor g00578(.dina(n775),.dinb(w_n743_69[1]),.dout(n776),.clk(gclk));
	jxor g00579(.dina(n776),.dinb(w_n648_0[0]),.dout(n777),.clk(gclk));
	jor g00580(.dina(w_n777_0[2]),.dinb(n774),.dout(n778),.clk(gclk));
	jand g00581(.dina(n778),.dinb(w_n773_0[1]),.dout(n779),.clk(gclk));
	jor g00582(.dina(w_n779_0[2]),.dinb(w_n294_70[2]),.dout(n780),.clk(gclk));
	jand g00583(.dina(w_n779_0[1]),.dinb(w_n294_70[1]),.dout(n781),.clk(gclk));
	jxor g00584(.dina(w_n650_0[0]),.dinb(w_n352_69[2]),.dout(n782),.clk(gclk));
	jor g00585(.dina(n782),.dinb(w_n743_69[0]),.dout(n783),.clk(gclk));
	jxor g00586(.dina(n783),.dinb(w_n708_0[0]),.dout(n784),.clk(gclk));
	jnot g00587(.din(w_n784_0[2]),.dout(n785),.clk(gclk));
	jor g00588(.dina(n785),.dinb(n781),.dout(n786),.clk(gclk));
	jand g00589(.dina(n786),.dinb(w_n780_0[1]),.dout(n787),.clk(gclk));
	jor g00590(.dina(w_n787_0[2]),.dinb(w_n239_70[2]),.dout(n788),.clk(gclk));
	jand g00591(.dina(w_n787_0[1]),.dinb(w_n239_70[1]),.dout(n789),.clk(gclk));
	jxor g00592(.dina(w_n657_0[0]),.dinb(w_n294_70[0]),.dout(n790),.clk(gclk));
	jor g00593(.dina(n790),.dinb(w_n743_68[2]),.dout(n791),.clk(gclk));
	jxor g00594(.dina(n791),.dinb(w_n663_0[0]),.dout(n792),.clk(gclk));
	jor g00595(.dina(w_n792_0[2]),.dinb(n789),.dout(n793),.clk(gclk));
	jand g00596(.dina(n793),.dinb(w_n788_0[1]),.dout(n794),.clk(gclk));
	jor g00597(.dina(w_n794_0[2]),.dinb(w_n221_71[0]),.dout(n795),.clk(gclk));
	jand g00598(.dina(w_n794_0[1]),.dinb(w_n221_70[2]),.dout(n796),.clk(gclk));
	jxor g00599(.dina(w_n665_0[0]),.dinb(w_n239_70[0]),.dout(n797),.clk(gclk));
	jor g00600(.dina(n797),.dinb(w_n743_68[1]),.dout(n798),.clk(gclk));
	jxor g00601(.dina(n798),.dinb(w_n715_0[0]),.dout(n799),.clk(gclk));
	jnot g00602(.din(w_n799_0[2]),.dout(n800),.clk(gclk));
	jor g00603(.dina(n800),.dinb(n796),.dout(n801),.clk(gclk));
	jand g00604(.dina(n801),.dinb(w_n795_0[1]),.dout(n802),.clk(gclk));
	jxor g00605(.dina(w_n672_0[0]),.dinb(w_n221_70[1]),.dout(n803),.clk(gclk));
	jor g00606(.dina(n803),.dinb(w_n743_68[0]),.dout(n804),.clk(gclk));
	jxor g00607(.dina(n804),.dinb(w_n678_0[0]),.dout(n805),.clk(gclk));
	jand g00608(.dina(w_n805_1[1]),.dinb(w_n802_0[2]),.dout(n806),.clk(gclk));
	jand g00609(.dina(w_n728_0[0]),.dinb(w_n736_0[0]),.dout(n808),.clk(gclk));
	jor g00610(.dina(w_n805_1[0]),.dinb(w_n802_0[1]),.dout(n809),.clk(gclk));
	jor g00611(.dina(w_n809_0[1]),.dinb(w_n682_0[0]),.dout(n810),.clk(gclk));
	jor g00612(.dina(n810),.dinb(w_n808_0[1]),.dout(n811),.clk(gclk));
	jand g00613(.dina(n811),.dinb(w_n218_29[0]),.dout(n812),.clk(gclk));
	jand g00614(.dina(w_n742_0[0]),.dinb(w_n720_0[0]),.dout(n813),.clk(gclk));
	jand g00615(.dina(w_n721_0[0]),.dinb(w_asqrt63_54[0]),.dout(n814),.clk(gclk));
	jand g00616(.dina(n814),.dinb(w_n681_0[2]),.dout(n815),.clk(gclk));
	jnot g00617(.din(n815),.dout(n816),.clk(gclk));
	jor g00618(.dina(w_n816_0[1]),.dinb(n813),.dout(n817),.clk(gclk));
	jnot g00619(.din(w_n817_0[1]),.dout(n818),.clk(gclk));
	jor g00620(.dina(n818),.dinb(n812),.dout(n819),.clk(gclk));
	jor g00621(.dina(w_n819_0[1]),.dinb(w_n806_0[2]),.dout(asqrt_fa_55),.clk(gclk));
	jnot g00622(.din(w_n795_0[0]),.dout(n822),.clk(gclk));
	jnot g00623(.din(w_n788_0[0]),.dout(n823),.clk(gclk));
	jnot g00624(.din(w_n780_0[0]),.dout(n824),.clk(gclk));
	jnot g00625(.din(w_n773_0[0]),.dout(n825),.clk(gclk));
	jnot g00626(.din(w_n765_0[0]),.dout(n826),.clk(gclk));
	jnot g00627(.din(w_n754_0[0]),.dout(n827),.clk(gclk));
	jnot g00628(.din(w_n746_0[0]),.dout(n828),.clk(gclk));
	jand g00629(.dina(w_asqrt55_41[0]),.dinb(w_a110_0[2]),.dout(n829),.clk(gclk));
	jor g00630(.dina(n829),.dinb(w_n733_0[0]),.dout(n830),.clk(gclk));
	jor g00631(.dina(n830),.dinb(w_asqrt56_41[1]),.dout(n831),.clk(gclk));
	jand g00632(.dina(w_asqrt55_40[2]),.dinb(w_n589_0[1]),.dout(n832),.clk(gclk));
	jor g00633(.dina(n832),.dinb(w_n590_0[0]),.dout(n833),.clk(gclk));
	jand g00634(.dina(w_n757_0[0]),.dinb(n833),.dout(n834),.clk(gclk));
	jand g00635(.dina(w_n834_0[1]),.dinb(n831),.dout(n835),.clk(gclk));
	jor g00636(.dina(n835),.dinb(n828),.dout(n836),.clk(gclk));
	jor g00637(.dina(n836),.dinb(w_asqrt57_41[0]),.dout(n837),.clk(gclk));
	jnot g00638(.din(w_n762_0[0]),.dout(n838),.clk(gclk));
	jand g00639(.dina(w_n838_0[1]),.dinb(n837),.dout(n839),.clk(gclk));
	jor g00640(.dina(n839),.dinb(n827),.dout(n840),.clk(gclk));
	jor g00641(.dina(n840),.dinb(w_asqrt58_41[2]),.dout(n841),.clk(gclk));
	jand g00642(.dina(w_n769_0[1]),.dinb(n841),.dout(n842),.clk(gclk));
	jor g00643(.dina(n842),.dinb(n826),.dout(n843),.clk(gclk));
	jor g00644(.dina(n843),.dinb(w_asqrt59_41[1]),.dout(n844),.clk(gclk));
	jnot g00645(.din(w_n777_0[1]),.dout(n845),.clk(gclk));
	jand g00646(.dina(n845),.dinb(n844),.dout(n846),.clk(gclk));
	jor g00647(.dina(n846),.dinb(n825),.dout(n847),.clk(gclk));
	jor g00648(.dina(n847),.dinb(w_asqrt60_41[2]),.dout(n848),.clk(gclk));
	jand g00649(.dina(w_n784_0[1]),.dinb(n848),.dout(n849),.clk(gclk));
	jor g00650(.dina(n849),.dinb(n824),.dout(n850),.clk(gclk));
	jor g00651(.dina(n850),.dinb(w_asqrt61_41[2]),.dout(n851),.clk(gclk));
	jnot g00652(.din(w_n792_0[1]),.dout(n852),.clk(gclk));
	jand g00653(.dina(n852),.dinb(n851),.dout(n853),.clk(gclk));
	jor g00654(.dina(n853),.dinb(n823),.dout(n854),.clk(gclk));
	jor g00655(.dina(n854),.dinb(w_asqrt62_41[2]),.dout(n855),.clk(gclk));
	jand g00656(.dina(w_n799_0[1]),.dinb(n855),.dout(n856),.clk(gclk));
	jor g00657(.dina(n856),.dinb(n822),.dout(n857),.clk(gclk));
	jnot g00658(.din(w_n805_0[2]),.dout(n858),.clk(gclk));
	jand g00659(.dina(n858),.dinb(n857),.dout(n859),.clk(gclk));
	jand g00660(.dina(w_n819_0[0]),.dinb(w_n859_0[1]),.dout(n860),.clk(gclk));
	jxor g00661(.dina(w_n794_0[0]),.dinb(w_n221_70[0]),.dout(n861),.clk(gclk));
	jand g00662(.dina(n861),.dinb(w_asqrt54_43[1]),.dout(n862),.clk(gclk));
	jxor g00663(.dina(n862),.dinb(w_n799_0[0]),.dout(n863),.clk(gclk));
	jnot g00664(.din(w_n863_0[2]),.dout(n864),.clk(gclk));
	jnot g00665(.din(w_a106_1[1]),.dout(n865),.clk(gclk));
	jnot g00666(.din(w_a107_0[1]),.dout(n866),.clk(gclk));
	jand g00667(.dina(w_n866_0[1]),.dinb(w_n865_1[1]),.dout(n867),.clk(gclk));
	jand g00668(.dina(w_n867_0[2]),.dinb(w_n730_1[1]),.dout(n868),.clk(gclk));
	jand g00669(.dina(w_asqrt54_43[0]),.dinb(w_a108_0[1]),.dout(n869),.clk(gclk));
	jor g00670(.dina(n869),.dinb(w_n868_0[1]),.dout(n870),.clk(gclk));
	jand g00671(.dina(w_n870_0[2]),.dinb(w_asqrt55_40[1]),.dout(n871),.clk(gclk));
	jor g00672(.dina(w_n870_0[1]),.dinb(w_asqrt55_40[0]),.dout(n872),.clk(gclk));
	jand g00673(.dina(w_asqrt54_42[2]),.dinb(w_n730_1[0]),.dout(n873),.clk(gclk));
	jor g00674(.dina(n873),.dinb(w_n731_0[0]),.dout(n874),.clk(gclk));
	jnot g00675(.din(w_n732_0[1]),.dout(n875),.clk(gclk));
	jnot g00676(.din(w_n806_0[1]),.dout(n876),.clk(gclk));
	jnot g00677(.din(w_n808_0[0]),.dout(n878),.clk(gclk));
	jand g00678(.dina(w_n859_0[0]),.dinb(w_n681_0[1]),.dout(n879),.clk(gclk));
	jand g00679(.dina(n879),.dinb(n878),.dout(n880),.clk(gclk));
	jor g00680(.dina(n880),.dinb(w_asqrt63_53[2]),.dout(n881),.clk(gclk));
	jand g00681(.dina(w_n817_0[0]),.dinb(w_n881_0[1]),.dout(n882),.clk(gclk));
	jand g00682(.dina(w_n882_0[1]),.dinb(w_n876_1[1]),.dout(n884),.clk(gclk));
	jor g00683(.dina(w_n884_67[2]),.dinb(n875),.dout(n885),.clk(gclk));
	jand g00684(.dina(n885),.dinb(n874),.dout(n886),.clk(gclk));
	jand g00685(.dina(w_n886_0[1]),.dinb(n872),.dout(n887),.clk(gclk));
	jor g00686(.dina(n887),.dinb(w_n871_0[1]),.dout(n888),.clk(gclk));
	jand g00687(.dina(w_n888_0[2]),.dinb(w_asqrt56_41[0]),.dout(n889),.clk(gclk));
	jor g00688(.dina(w_n888_0[1]),.dinb(w_asqrt56_40[2]),.dout(n890),.clk(gclk));
	jand g00689(.dina(w_asqrt54_42[1]),.dinb(w_n732_0[0]),.dout(n891),.clk(gclk));
	jand g00690(.dina(w_n816_0[0]),.dinb(w_n876_1[0]),.dout(n892),.clk(gclk));
	jand g00691(.dina(n892),.dinb(w_n881_0[0]),.dout(n893),.clk(gclk));
	jand g00692(.dina(n893),.dinb(w_asqrt55_39[2]),.dout(n894),.clk(gclk));
	jor g00693(.dina(n894),.dinb(w_n891_0[1]),.dout(n895),.clk(gclk));
	jxor g00694(.dina(n895),.dinb(w_a110_0[1]),.dout(n896),.clk(gclk));
	jnot g00695(.din(w_n896_0[1]),.dout(n897),.clk(gclk));
	jand g00696(.dina(w_n897_0[1]),.dinb(n890),.dout(n898),.clk(gclk));
	jor g00697(.dina(n898),.dinb(w_n889_0[1]),.dout(n899),.clk(gclk));
	jand g00698(.dina(w_n899_0[2]),.dinb(w_asqrt57_40[2]),.dout(n900),.clk(gclk));
	jor g00699(.dina(w_n899_0[1]),.dinb(w_asqrt57_40[1]),.dout(n901),.clk(gclk));
	jxor g00700(.dina(w_n745_0[0]),.dinb(w_n635_68[0]),.dout(n902),.clk(gclk));
	jand g00701(.dina(n902),.dinb(w_asqrt54_42[0]),.dout(n903),.clk(gclk));
	jxor g00702(.dina(n903),.dinb(w_n834_0[0]),.dout(n904),.clk(gclk));
	jand g00703(.dina(w_n904_0[1]),.dinb(n901),.dout(n905),.clk(gclk));
	jor g00704(.dina(n905),.dinb(w_n900_0[1]),.dout(n906),.clk(gclk));
	jand g00705(.dina(w_n906_0[2]),.dinb(w_asqrt58_41[1]),.dout(n907),.clk(gclk));
	jor g00706(.dina(w_n906_0[1]),.dinb(w_asqrt58_41[0]),.dout(n908),.clk(gclk));
	jxor g00707(.dina(w_n753_0[0]),.dinb(w_n515_69[0]),.dout(n909),.clk(gclk));
	jand g00708(.dina(n909),.dinb(w_asqrt54_41[2]),.dout(n910),.clk(gclk));
	jxor g00709(.dina(n910),.dinb(w_n838_0[0]),.dout(n911),.clk(gclk));
	jand g00710(.dina(w_n911_0[1]),.dinb(n908),.dout(n912),.clk(gclk));
	jor g00711(.dina(n912),.dinb(w_n907_0[1]),.dout(n913),.clk(gclk));
	jand g00712(.dina(w_n913_0[2]),.dinb(w_asqrt59_41[0]),.dout(n914),.clk(gclk));
	jor g00713(.dina(w_n913_0[1]),.dinb(w_asqrt59_40[2]),.dout(n915),.clk(gclk));
	jxor g00714(.dina(w_n764_0[0]),.dinb(w_n443_69[0]),.dout(n916),.clk(gclk));
	jand g00715(.dina(n916),.dinb(w_asqrt54_41[1]),.dout(n917),.clk(gclk));
	jxor g00716(.dina(n917),.dinb(w_n769_0[0]),.dout(n918),.clk(gclk));
	jand g00717(.dina(w_n918_0[1]),.dinb(n915),.dout(n919),.clk(gclk));
	jor g00718(.dina(n919),.dinb(w_n914_0[1]),.dout(n920),.clk(gclk));
	jand g00719(.dina(w_n920_0[2]),.dinb(w_asqrt60_41[1]),.dout(n921),.clk(gclk));
	jor g00720(.dina(w_n920_0[1]),.dinb(w_asqrt60_41[0]),.dout(n922),.clk(gclk));
	jxor g00721(.dina(w_n772_0[0]),.dinb(w_n352_69[1]),.dout(n923),.clk(gclk));
	jand g00722(.dina(n923),.dinb(w_asqrt54_41[0]),.dout(n924),.clk(gclk));
	jxor g00723(.dina(n924),.dinb(w_n777_0[0]),.dout(n925),.clk(gclk));
	jnot g00724(.din(w_n925_0[1]),.dout(n926),.clk(gclk));
	jand g00725(.dina(w_n926_0[1]),.dinb(n922),.dout(n927),.clk(gclk));
	jor g00726(.dina(n927),.dinb(w_n921_0[1]),.dout(n928),.clk(gclk));
	jand g00727(.dina(w_n928_0[2]),.dinb(w_asqrt61_41[1]),.dout(n929),.clk(gclk));
	jor g00728(.dina(w_n928_0[1]),.dinb(w_asqrt61_41[0]),.dout(n930),.clk(gclk));
	jxor g00729(.dina(w_n779_0[0]),.dinb(w_n294_69[2]),.dout(n931),.clk(gclk));
	jand g00730(.dina(n931),.dinb(w_asqrt54_40[2]),.dout(n932),.clk(gclk));
	jxor g00731(.dina(n932),.dinb(w_n784_0[0]),.dout(n933),.clk(gclk));
	jand g00732(.dina(w_n933_0[1]),.dinb(n930),.dout(n934),.clk(gclk));
	jor g00733(.dina(n934),.dinb(w_n929_0[1]),.dout(n935),.clk(gclk));
	jand g00734(.dina(w_n935_0[2]),.dinb(w_asqrt62_41[1]),.dout(n936),.clk(gclk));
	jnot g00735(.din(w_n936_0[1]),.dout(n937),.clk(gclk));
	jnot g00736(.din(w_n929_0[0]),.dout(n938),.clk(gclk));
	jnot g00737(.din(w_n921_0[0]),.dout(n939),.clk(gclk));
	jnot g00738(.din(w_n914_0[0]),.dout(n940),.clk(gclk));
	jnot g00739(.din(w_n907_0[0]),.dout(n941),.clk(gclk));
	jnot g00740(.din(w_n900_0[0]),.dout(n942),.clk(gclk));
	jnot g00741(.din(w_n889_0[0]),.dout(n943),.clk(gclk));
	jnot g00742(.din(w_n871_0[0]),.dout(n944),.clk(gclk));
	jnot g00743(.din(w_n868_0[0]),.dout(n945),.clk(gclk));
	jor g00744(.dina(w_n884_67[1]),.dinb(w_n730_0[2]),.dout(n946),.clk(gclk));
	jand g00745(.dina(n946),.dinb(n945),.dout(n947),.clk(gclk));
	jand g00746(.dina(n947),.dinb(w_n743_67[2]),.dout(n948),.clk(gclk));
	jor g00747(.dina(w_n884_67[0]),.dinb(w_a108_0[0]),.dout(n949),.clk(gclk));
	jand g00748(.dina(n949),.dinb(w_a109_0[0]),.dout(n950),.clk(gclk));
	jor g00749(.dina(w_n891_0[0]),.dinb(n950),.dout(n951),.clk(gclk));
	jor g00750(.dina(n951),.dinb(n948),.dout(n952),.clk(gclk));
	jand g00751(.dina(n952),.dinb(n944),.dout(n953),.clk(gclk));
	jand g00752(.dina(n953),.dinb(w_n635_67[2]),.dout(n954),.clk(gclk));
	jor g00753(.dina(w_n896_0[0]),.dinb(n954),.dout(n955),.clk(gclk));
	jand g00754(.dina(n955),.dinb(n943),.dout(n956),.clk(gclk));
	jand g00755(.dina(n956),.dinb(w_n515_68[2]),.dout(n957),.clk(gclk));
	jnot g00756(.din(w_n904_0[0]),.dout(n958),.clk(gclk));
	jor g00757(.dina(w_n958_0[1]),.dinb(n957),.dout(n959),.clk(gclk));
	jand g00758(.dina(n959),.dinb(n942),.dout(n960),.clk(gclk));
	jand g00759(.dina(n960),.dinb(w_n443_68[2]),.dout(n961),.clk(gclk));
	jnot g00760(.din(w_n911_0[0]),.dout(n962),.clk(gclk));
	jor g00761(.dina(w_n962_0[1]),.dinb(n961),.dout(n963),.clk(gclk));
	jand g00762(.dina(n963),.dinb(n941),.dout(n964),.clk(gclk));
	jand g00763(.dina(n964),.dinb(w_n352_69[0]),.dout(n965),.clk(gclk));
	jnot g00764(.din(w_n918_0[0]),.dout(n966),.clk(gclk));
	jor g00765(.dina(w_n966_0[1]),.dinb(n965),.dout(n967),.clk(gclk));
	jand g00766(.dina(n967),.dinb(n940),.dout(n968),.clk(gclk));
	jand g00767(.dina(n968),.dinb(w_n294_69[1]),.dout(n969),.clk(gclk));
	jor g00768(.dina(w_n925_0[0]),.dinb(n969),.dout(n970),.clk(gclk));
	jand g00769(.dina(n970),.dinb(n939),.dout(n971),.clk(gclk));
	jand g00770(.dina(n971),.dinb(w_n239_69[2]),.dout(n972),.clk(gclk));
	jnot g00771(.din(w_n933_0[0]),.dout(n973),.clk(gclk));
	jor g00772(.dina(w_n973_0[1]),.dinb(n972),.dout(n974),.clk(gclk));
	jand g00773(.dina(n974),.dinb(n938),.dout(n975),.clk(gclk));
	jand g00774(.dina(n975),.dinb(w_n221_69[2]),.dout(n976),.clk(gclk));
	jxor g00775(.dina(w_n787_0[0]),.dinb(w_n239_69[1]),.dout(n977),.clk(gclk));
	jand g00776(.dina(n977),.dinb(w_asqrt54_40[1]),.dout(n978),.clk(gclk));
	jxor g00777(.dina(n978),.dinb(w_n792_0[0]),.dout(n979),.clk(gclk));
	jor g00778(.dina(w_n979_0[1]),.dinb(n976),.dout(n980),.clk(gclk));
	jand g00779(.dina(n980),.dinb(n937),.dout(n981),.clk(gclk));
	jor g00780(.dina(w_n981_0[1]),.dinb(w_n864_0[1]),.dout(n982),.clk(gclk));
	jor g00781(.dina(w_n982_0[1]),.dinb(w_n806_0[0]),.dout(n983),.clk(gclk));
	jor g00782(.dina(n983),.dinb(w_n860_0[1]),.dout(n984),.clk(gclk));
	jand g00783(.dina(n984),.dinb(w_n218_28[2]),.dout(n985),.clk(gclk));
	jand g00784(.dina(w_n884_66[2]),.dinb(w_n805_0[1]),.dout(n986),.clk(gclk));
	jnot g00785(.din(n986),.dout(n987),.clk(gclk));
	jor g00786(.dina(w_n935_0[1]),.dinb(w_asqrt62_41[0]),.dout(n988),.clk(gclk));
	jnot g00787(.din(w_n979_0[0]),.dout(n989),.clk(gclk));
	jand g00788(.dina(w_n989_0[1]),.dinb(n988),.dout(n990),.clk(gclk));
	jor g00789(.dina(n990),.dinb(w_n936_0[0]),.dout(n991),.clk(gclk));
	jor g00790(.dina(w_n991_0[1]),.dinb(w_n863_0[1]),.dout(n992),.clk(gclk));
	jand g00791(.dina(w_n992_0[2]),.dinb(n987),.dout(n993),.clk(gclk));
	jand g00792(.dina(w_n882_0[0]),.dinb(w_n802_0[0]),.dout(n994),.clk(gclk));
	jnot g00793(.din(n994),.dout(n995),.clk(gclk));
	jand g00794(.dina(w_n809_0[0]),.dinb(w_asqrt63_53[1]),.dout(n996),.clk(gclk));
	jand g00795(.dina(n996),.dinb(w_n876_0[2]),.dout(n997),.clk(gclk));
	jand g00796(.dina(w_n997_0[1]),.dinb(n995),.dout(n998),.clk(gclk));
	jnot g00797(.din(n998),.dout(n999),.clk(gclk));
	jand g00798(.dina(n999),.dinb(n993),.dout(n1000),.clk(gclk));
	jnot g00799(.din(w_n1000_0[1]),.dout(n1001),.clk(gclk));
	jor g00800(.dina(n1001),.dinb(w_n985_0[1]),.dout(asqrt_fa_54),.clk(gclk));
	jnot g00801(.din(w_n860_0[0]),.dout(n1003),.clk(gclk));
	jand g00802(.dina(w_n991_0[0]),.dinb(w_n863_0[0]),.dout(n1004),.clk(gclk));
	jand g00803(.dina(w_n1004_0[1]),.dinb(w_n876_0[1]),.dout(n1005),.clk(gclk));
	jand g00804(.dina(n1005),.dinb(n1003),.dout(n1006),.clk(gclk));
	jor g00805(.dina(n1006),.dinb(w_asqrt63_53[0]),.dout(n1007),.clk(gclk));
	jand g00806(.dina(w_n1000_0[0]),.dinb(n1007),.dout(n1008),.clk(gclk));
	jor g00807(.dina(w_n1008_70[1]),.dinb(w_n865_1[0]),.dout(n1009),.clk(gclk));
	jnot g00808(.din(w_a104_0[2]),.dout(n1010),.clk(gclk));
	jnot g00809(.din(w_a105_0[1]),.dout(n1011),.clk(gclk));
	jand g00810(.dina(w_n1011_0[1]),.dinb(w_n1010_1[2]),.dout(n1012),.clk(gclk));
	jand g00811(.dina(w_n1012_0[2]),.dinb(w_n865_0[2]),.dout(n1013),.clk(gclk));
	jnot g00812(.din(w_n1013_0[1]),.dout(n1014),.clk(gclk));
	jand g00813(.dina(n1014),.dinb(n1009),.dout(n1015),.clk(gclk));
	jor g00814(.dina(w_n1015_0[2]),.dinb(w_n884_66[1]),.dout(n1016),.clk(gclk));
	jand g00815(.dina(w_n1015_0[1]),.dinb(w_n884_66[0]),.dout(n1017),.clk(gclk));
	jor g00816(.dina(w_n1008_70[0]),.dinb(w_a106_1[0]),.dout(n1018),.clk(gclk));
	jand g00817(.dina(n1018),.dinb(w_a107_0[0]),.dout(n1019),.clk(gclk));
	jand g00818(.dina(w_asqrt53_40[1]),.dinb(w_n867_0[1]),.dout(n1020),.clk(gclk));
	jor g00819(.dina(n1020),.dinb(n1019),.dout(n1021),.clk(gclk));
	jor g00820(.dina(n1021),.dinb(n1017),.dout(n1022),.clk(gclk));
	jand g00821(.dina(n1022),.dinb(w_n1016_0[1]),.dout(n1023),.clk(gclk));
	jor g00822(.dina(w_n1023_0[2]),.dinb(w_n743_67[1]),.dout(n1024),.clk(gclk));
	jand g00823(.dina(w_n1023_0[1]),.dinb(w_n743_67[0]),.dout(n1025),.clk(gclk));
	jnot g00824(.din(w_n867_0[0]),.dout(n1026),.clk(gclk));
	jor g00825(.dina(w_n1008_69[2]),.dinb(n1026),.dout(n1027),.clk(gclk));
	jnot g00826(.din(w_n992_0[1]),.dout(n1028),.clk(gclk));
	jor g00827(.dina(w_n997_0[0]),.dinb(w_n884_65[2]),.dout(n1029),.clk(gclk));
	jor g00828(.dina(n1029),.dinb(w_n985_0[0]),.dout(n1030),.clk(gclk));
	jor g00829(.dina(n1030),.dinb(w_n1028_0[1]),.dout(n1031),.clk(gclk));
	jand g00830(.dina(n1031),.dinb(w_n1027_0[1]),.dout(n1032),.clk(gclk));
	jxor g00831(.dina(n1032),.dinb(w_n730_0[1]),.dout(n1033),.clk(gclk));
	jor g00832(.dina(w_n1033_0[2]),.dinb(n1025),.dout(n1034),.clk(gclk));
	jand g00833(.dina(n1034),.dinb(w_n1024_0[1]),.dout(n1035),.clk(gclk));
	jor g00834(.dina(w_n1035_0[2]),.dinb(w_n635_67[1]),.dout(n1036),.clk(gclk));
	jand g00835(.dina(w_n1035_0[1]),.dinb(w_n635_67[0]),.dout(n1037),.clk(gclk));
	jxor g00836(.dina(w_n870_0[0]),.dinb(w_n743_66[2]),.dout(n1038),.clk(gclk));
	jor g00837(.dina(n1038),.dinb(w_n1008_69[1]),.dout(n1039),.clk(gclk));
	jxor g00838(.dina(n1039),.dinb(w_n886_0[0]),.dout(n1040),.clk(gclk));
	jor g00839(.dina(w_n1040_0[2]),.dinb(n1037),.dout(n1041),.clk(gclk));
	jand g00840(.dina(n1041),.dinb(w_n1036_0[1]),.dout(n1042),.clk(gclk));
	jor g00841(.dina(w_n1042_0[2]),.dinb(w_n515_68[1]),.dout(n1043),.clk(gclk));
	jand g00842(.dina(w_n1042_0[1]),.dinb(w_n515_68[0]),.dout(n1044),.clk(gclk));
	jxor g00843(.dina(w_n888_0[0]),.dinb(w_n635_66[2]),.dout(n1045),.clk(gclk));
	jor g00844(.dina(n1045),.dinb(w_n1008_69[0]),.dout(n1046),.clk(gclk));
	jxor g00845(.dina(n1046),.dinb(w_n897_0[0]),.dout(n1047),.clk(gclk));
	jor g00846(.dina(w_n1047_0[2]),.dinb(n1044),.dout(n1048),.clk(gclk));
	jand g00847(.dina(n1048),.dinb(w_n1043_0[1]),.dout(n1049),.clk(gclk));
	jor g00848(.dina(w_n1049_0[2]),.dinb(w_n443_68[1]),.dout(n1050),.clk(gclk));
	jand g00849(.dina(w_n1049_0[1]),.dinb(w_n443_68[0]),.dout(n1051),.clk(gclk));
	jxor g00850(.dina(w_n899_0[0]),.dinb(w_n515_67[2]),.dout(n1052),.clk(gclk));
	jor g00851(.dina(n1052),.dinb(w_n1008_68[2]),.dout(n1053),.clk(gclk));
	jxor g00852(.dina(n1053),.dinb(w_n958_0[0]),.dout(n1054),.clk(gclk));
	jnot g00853(.din(w_n1054_0[2]),.dout(n1055),.clk(gclk));
	jor g00854(.dina(n1055),.dinb(n1051),.dout(n1056),.clk(gclk));
	jand g00855(.dina(n1056),.dinb(w_n1050_0[1]),.dout(n1057),.clk(gclk));
	jor g00856(.dina(w_n1057_0[2]),.dinb(w_n352_68[2]),.dout(n1058),.clk(gclk));
	jand g00857(.dina(w_n1057_0[1]),.dinb(w_n352_68[1]),.dout(n1059),.clk(gclk));
	jxor g00858(.dina(w_n906_0[0]),.dinb(w_n443_67[2]),.dout(n1060),.clk(gclk));
	jor g00859(.dina(n1060),.dinb(w_n1008_68[1]),.dout(n1061),.clk(gclk));
	jxor g00860(.dina(n1061),.dinb(w_n962_0[0]),.dout(n1062),.clk(gclk));
	jnot g00861(.din(w_n1062_0[2]),.dout(n1063),.clk(gclk));
	jor g00862(.dina(n1063),.dinb(n1059),.dout(n1064),.clk(gclk));
	jand g00863(.dina(n1064),.dinb(w_n1058_0[1]),.dout(n1065),.clk(gclk));
	jor g00864(.dina(w_n1065_0[2]),.dinb(w_n294_69[0]),.dout(n1066),.clk(gclk));
	jand g00865(.dina(w_n1065_0[1]),.dinb(w_n294_68[2]),.dout(n1067),.clk(gclk));
	jxor g00866(.dina(w_n913_0[0]),.dinb(w_n352_68[0]),.dout(n1068),.clk(gclk));
	jor g00867(.dina(n1068),.dinb(w_n1008_68[0]),.dout(n1069),.clk(gclk));
	jxor g00868(.dina(n1069),.dinb(w_n966_0[0]),.dout(n1070),.clk(gclk));
	jnot g00869(.din(w_n1070_0[2]),.dout(n1071),.clk(gclk));
	jor g00870(.dina(n1071),.dinb(n1067),.dout(n1072),.clk(gclk));
	jand g00871(.dina(n1072),.dinb(w_n1066_0[1]),.dout(n1073),.clk(gclk));
	jor g00872(.dina(w_n1073_0[2]),.dinb(w_n239_69[0]),.dout(n1074),.clk(gclk));
	jand g00873(.dina(w_n1073_0[1]),.dinb(w_n239_68[2]),.dout(n1075),.clk(gclk));
	jxor g00874(.dina(w_n920_0[0]),.dinb(w_n294_68[1]),.dout(n1076),.clk(gclk));
	jor g00875(.dina(n1076),.dinb(w_n1008_67[2]),.dout(n1077),.clk(gclk));
	jxor g00876(.dina(n1077),.dinb(w_n926_0[0]),.dout(n1078),.clk(gclk));
	jor g00877(.dina(w_n1078_0[2]),.dinb(n1075),.dout(n1079),.clk(gclk));
	jand g00878(.dina(n1079),.dinb(w_n1074_0[1]),.dout(n1080),.clk(gclk));
	jor g00879(.dina(w_n1080_0[2]),.dinb(w_n221_69[1]),.dout(n1081),.clk(gclk));
	jand g00880(.dina(w_n1080_0[1]),.dinb(w_n221_69[0]),.dout(n1082),.clk(gclk));
	jxor g00881(.dina(w_n928_0[0]),.dinb(w_n239_68[1]),.dout(n1083),.clk(gclk));
	jor g00882(.dina(n1083),.dinb(w_n1008_67[1]),.dout(n1084),.clk(gclk));
	jxor g00883(.dina(n1084),.dinb(w_n973_0[0]),.dout(n1085),.clk(gclk));
	jnot g00884(.din(w_n1085_0[1]),.dout(n1086),.clk(gclk));
	jor g00885(.dina(w_n1086_0[1]),.dinb(n1082),.dout(n1087),.clk(gclk));
	jand g00886(.dina(n1087),.dinb(w_n1081_0[1]),.dout(n1088),.clk(gclk));
	jxor g00887(.dina(w_n935_0[0]),.dinb(w_n221_68[2]),.dout(n1089),.clk(gclk));
	jor g00888(.dina(n1089),.dinb(w_n1008_67[0]),.dout(n1090),.clk(gclk));
	jxor g00889(.dina(n1090),.dinb(w_n989_0[0]),.dout(n1091),.clk(gclk));
	jand g00890(.dina(w_n1091_1[1]),.dinb(w_n1088_1[1]),.dout(n1092),.clk(gclk));
	jand g00891(.dina(w_n1008_66[2]),.dinb(w_n981_0[0]),.dout(n1093),.clk(gclk));
	jand g00892(.dina(w_n982_0[0]),.dinb(w_asqrt63_52[2]),.dout(n1094),.clk(gclk));
	jand g00893(.dina(n1094),.dinb(w_n992_0[0]),.dout(n1095),.clk(gclk));
	jnot g00894(.din(n1095),.dout(n1096),.clk(gclk));
	jor g00895(.dina(w_n1096_0[1]),.dinb(n1093),.dout(n1097),.clk(gclk));
	jnot g00896(.din(w_n1097_0[1]),.dout(n1098),.clk(gclk));
	jor g00897(.dina(w_n1091_1[0]),.dinb(w_n1088_1[0]),.dout(n1099),.clk(gclk));
	jand g00898(.dina(w_asqrt53_40[0]),.dinb(w_n1004_0[0]),.dout(n1100),.clk(gclk));
	jor g00899(.dina(n1100),.dinb(w_n1028_0[0]),.dout(n1101),.clk(gclk));
	jor g00900(.dina(w_n1101_0[1]),.dinb(n1099),.dout(n1102),.clk(gclk));
	jand g00901(.dina(n1102),.dinb(w_n218_28[1]),.dout(n1103),.clk(gclk));
	jand g00902(.dina(w_n1008_66[1]),.dinb(w_n864_0[0]),.dout(n1104),.clk(gclk));
	jor g00903(.dina(w_n1104_0[1]),.dinb(n1103),.dout(n1105),.clk(gclk));
	jor g00904(.dina(n1105),.dinb(n1098),.dout(n1106),.clk(gclk));
	jor g00905(.dina(n1106),.dinb(w_n1092_0[1]),.dout(asqrt_fa_53),.clk(gclk));
	jnot g00906(.din(w_a102_1[1]),.dout(n1108),.clk(gclk));
	jnot g00907(.din(w_a103_0[1]),.dout(n1109),.clk(gclk));
	jand g00908(.dina(w_n1109_0[1]),.dinb(w_n1108_1[1]),.dout(n1110),.clk(gclk));
	jand g00909(.dina(w_n1110_0[2]),.dinb(w_n1010_1[1]),.dout(n1111),.clk(gclk));
	jand g00910(.dina(w_asqrt52_43[1]),.dinb(w_a104_0[1]),.dout(n1112),.clk(gclk));
	jor g00911(.dina(n1112),.dinb(w_n1111_0[1]),.dout(n1113),.clk(gclk));
	jand g00912(.dina(w_n1113_0[2]),.dinb(w_asqrt53_39[2]),.dout(n1114),.clk(gclk));
	jor g00913(.dina(w_n1113_0[1]),.dinb(w_asqrt53_39[1]),.dout(n1115),.clk(gclk));
	jand g00914(.dina(w_asqrt52_43[0]),.dinb(w_n1010_1[0]),.dout(n1116),.clk(gclk));
	jor g00915(.dina(n1116),.dinb(w_n1011_0[0]),.dout(n1117),.clk(gclk));
	jnot g00916(.din(w_n1012_0[1]),.dout(n1118),.clk(gclk));
	jnot g00917(.din(w_n1092_0[0]),.dout(n1119),.clk(gclk));
	jnot g00918(.din(w_n1081_0[0]),.dout(n1120),.clk(gclk));
	jnot g00919(.din(w_n1074_0[0]),.dout(n1121),.clk(gclk));
	jnot g00920(.din(w_n1066_0[0]),.dout(n1122),.clk(gclk));
	jnot g00921(.din(w_n1058_0[0]),.dout(n1123),.clk(gclk));
	jnot g00922(.din(w_n1050_0[0]),.dout(n1124),.clk(gclk));
	jnot g00923(.din(w_n1043_0[0]),.dout(n1125),.clk(gclk));
	jnot g00924(.din(w_n1036_0[0]),.dout(n1126),.clk(gclk));
	jnot g00925(.din(w_n1024_0[0]),.dout(n1127),.clk(gclk));
	jnot g00926(.din(w_n1016_0[0]),.dout(n1128),.clk(gclk));
	jand g00927(.dina(w_asqrt53_39[0]),.dinb(w_a106_0[2]),.dout(n1129),.clk(gclk));
	jor g00928(.dina(w_n1013_0[0]),.dinb(n1129),.dout(n1130),.clk(gclk));
	jor g00929(.dina(n1130),.dinb(w_asqrt54_40[0]),.dout(n1131),.clk(gclk));
	jand g00930(.dina(w_asqrt53_38[2]),.dinb(w_n865_0[1]),.dout(n1132),.clk(gclk));
	jor g00931(.dina(n1132),.dinb(w_n866_0[0]),.dout(n1133),.clk(gclk));
	jand g00932(.dina(w_n1027_0[0]),.dinb(n1133),.dout(n1134),.clk(gclk));
	jand g00933(.dina(w_n1134_0[1]),.dinb(n1131),.dout(n1135),.clk(gclk));
	jor g00934(.dina(n1135),.dinb(n1128),.dout(n1136),.clk(gclk));
	jor g00935(.dina(n1136),.dinb(w_asqrt55_39[1]),.dout(n1137),.clk(gclk));
	jnot g00936(.din(w_n1033_0[1]),.dout(n1138),.clk(gclk));
	jand g00937(.dina(n1138),.dinb(n1137),.dout(n1139),.clk(gclk));
	jor g00938(.dina(n1139),.dinb(n1127),.dout(n1140),.clk(gclk));
	jor g00939(.dina(n1140),.dinb(w_asqrt56_40[1]),.dout(n1141),.clk(gclk));
	jnot g00940(.din(w_n1040_0[1]),.dout(n1142),.clk(gclk));
	jand g00941(.dina(n1142),.dinb(n1141),.dout(n1143),.clk(gclk));
	jor g00942(.dina(n1143),.dinb(n1126),.dout(n1144),.clk(gclk));
	jor g00943(.dina(n1144),.dinb(w_asqrt57_40[0]),.dout(n1145),.clk(gclk));
	jnot g00944(.din(w_n1047_0[1]),.dout(n1146),.clk(gclk));
	jand g00945(.dina(n1146),.dinb(n1145),.dout(n1147),.clk(gclk));
	jor g00946(.dina(n1147),.dinb(n1125),.dout(n1148),.clk(gclk));
	jor g00947(.dina(n1148),.dinb(w_asqrt58_40[2]),.dout(n1149),.clk(gclk));
	jand g00948(.dina(w_n1054_0[1]),.dinb(n1149),.dout(n1150),.clk(gclk));
	jor g00949(.dina(n1150),.dinb(n1124),.dout(n1151),.clk(gclk));
	jor g00950(.dina(n1151),.dinb(w_asqrt59_40[1]),.dout(n1152),.clk(gclk));
	jand g00951(.dina(w_n1062_0[1]),.dinb(n1152),.dout(n1153),.clk(gclk));
	jor g00952(.dina(n1153),.dinb(n1123),.dout(n1154),.clk(gclk));
	jor g00953(.dina(n1154),.dinb(w_asqrt60_40[2]),.dout(n1155),.clk(gclk));
	jand g00954(.dina(w_n1070_0[1]),.dinb(n1155),.dout(n1156),.clk(gclk));
	jor g00955(.dina(n1156),.dinb(n1122),.dout(n1157),.clk(gclk));
	jor g00956(.dina(n1157),.dinb(w_asqrt61_40[2]),.dout(n1158),.clk(gclk));
	jnot g00957(.din(w_n1078_0[1]),.dout(n1159),.clk(gclk));
	jand g00958(.dina(n1159),.dinb(n1158),.dout(n1160),.clk(gclk));
	jor g00959(.dina(n1160),.dinb(n1121),.dout(n1161),.clk(gclk));
	jor g00960(.dina(n1161),.dinb(w_asqrt62_40[2]),.dout(n1162),.clk(gclk));
	jand g00961(.dina(w_n1085_0[0]),.dinb(n1162),.dout(n1163),.clk(gclk));
	jor g00962(.dina(n1163),.dinb(n1120),.dout(n1164),.clk(gclk));
	jnot g00963(.din(w_n1091_0[2]),.dout(n1165),.clk(gclk));
	jand g00964(.dina(n1165),.dinb(n1164),.dout(n1166),.clk(gclk));
	jnot g00965(.din(w_n1101_0[0]),.dout(n1167),.clk(gclk));
	jand g00966(.dina(n1167),.dinb(n1166),.dout(n1168),.clk(gclk));
	jor g00967(.dina(n1168),.dinb(w_asqrt63_52[1]),.dout(n1169),.clk(gclk));
	jnot g00968(.din(w_n1104_0[0]),.dout(n1170),.clk(gclk));
	jand g00969(.dina(n1170),.dinb(w_n1169_0[1]),.dout(n1171),.clk(gclk));
	jand g00970(.dina(n1171),.dinb(w_n1097_0[0]),.dout(n1172),.clk(gclk));
	jand g00971(.dina(w_n1172_0[1]),.dinb(w_n1119_0[1]),.dout(n1173),.clk(gclk));
	jor g00972(.dina(w_n1173_64[2]),.dinb(n1118),.dout(n1174),.clk(gclk));
	jand g00973(.dina(n1174),.dinb(n1117),.dout(n1175),.clk(gclk));
	jand g00974(.dina(w_n1175_0[1]),.dinb(n1115),.dout(n1176),.clk(gclk));
	jor g00975(.dina(n1176),.dinb(w_n1114_0[1]),.dout(n1177),.clk(gclk));
	jand g00976(.dina(w_n1177_0[2]),.dinb(w_asqrt54_39[2]),.dout(n1178),.clk(gclk));
	jor g00977(.dina(w_n1177_0[1]),.dinb(w_asqrt54_39[1]),.dout(n1179),.clk(gclk));
	jand g00978(.dina(w_asqrt52_42[2]),.dinb(w_n1012_0[0]),.dout(n1180),.clk(gclk));
	jand g00979(.dina(w_n1119_0[0]),.dinb(w_asqrt53_38[1]),.dout(n1181),.clk(gclk));
	jand g00980(.dina(n1181),.dinb(w_n1096_0[0]),.dout(n1182),.clk(gclk));
	jand g00981(.dina(n1182),.dinb(w_n1169_0[0]),.dout(n1183),.clk(gclk));
	jor g00982(.dina(n1183),.dinb(w_n1180_0[1]),.dout(n1184),.clk(gclk));
	jxor g00983(.dina(n1184),.dinb(w_a106_0[1]),.dout(n1185),.clk(gclk));
	jnot g00984(.din(w_n1185_0[1]),.dout(n1186),.clk(gclk));
	jand g00985(.dina(w_n1186_0[1]),.dinb(n1179),.dout(n1187),.clk(gclk));
	jor g00986(.dina(n1187),.dinb(w_n1178_0[1]),.dout(n1188),.clk(gclk));
	jand g00987(.dina(w_n1188_0[2]),.dinb(w_asqrt55_39[0]),.dout(n1189),.clk(gclk));
	jor g00988(.dina(w_n1188_0[1]),.dinb(w_asqrt55_38[2]),.dout(n1190),.clk(gclk));
	jxor g00989(.dina(w_n1015_0[0]),.dinb(w_n884_65[1]),.dout(n1191),.clk(gclk));
	jand g00990(.dina(n1191),.dinb(w_asqrt52_42[1]),.dout(n1192),.clk(gclk));
	jxor g00991(.dina(n1192),.dinb(w_n1134_0[0]),.dout(n1193),.clk(gclk));
	jand g00992(.dina(w_n1193_0[1]),.dinb(n1190),.dout(n1194),.clk(gclk));
	jor g00993(.dina(n1194),.dinb(w_n1189_0[1]),.dout(n1195),.clk(gclk));
	jand g00994(.dina(w_n1195_0[2]),.dinb(w_asqrt56_40[0]),.dout(n1196),.clk(gclk));
	jor g00995(.dina(w_n1195_0[1]),.dinb(w_asqrt56_39[2]),.dout(n1197),.clk(gclk));
	jxor g00996(.dina(w_n1023_0[0]),.dinb(w_n743_66[1]),.dout(n1198),.clk(gclk));
	jand g00997(.dina(n1198),.dinb(w_asqrt52_42[0]),.dout(n1199),.clk(gclk));
	jxor g00998(.dina(n1199),.dinb(w_n1033_0[0]),.dout(n1200),.clk(gclk));
	jnot g00999(.din(w_n1200_0[1]),.dout(n1201),.clk(gclk));
	jand g01000(.dina(w_n1201_0[1]),.dinb(n1197),.dout(n1202),.clk(gclk));
	jor g01001(.dina(n1202),.dinb(w_n1196_0[1]),.dout(n1203),.clk(gclk));
	jand g01002(.dina(w_n1203_0[2]),.dinb(w_asqrt57_39[2]),.dout(n1204),.clk(gclk));
	jor g01003(.dina(w_n1203_0[1]),.dinb(w_asqrt57_39[1]),.dout(n1205),.clk(gclk));
	jxor g01004(.dina(w_n1035_0[0]),.dinb(w_n635_66[1]),.dout(n1206),.clk(gclk));
	jand g01005(.dina(n1206),.dinb(w_asqrt52_41[2]),.dout(n1207),.clk(gclk));
	jxor g01006(.dina(n1207),.dinb(w_n1040_0[0]),.dout(n1208),.clk(gclk));
	jnot g01007(.din(w_n1208_0[1]),.dout(n1209),.clk(gclk));
	jand g01008(.dina(w_n1209_0[1]),.dinb(n1205),.dout(n1210),.clk(gclk));
	jor g01009(.dina(n1210),.dinb(w_n1204_0[1]),.dout(n1211),.clk(gclk));
	jand g01010(.dina(w_n1211_0[2]),.dinb(w_asqrt58_40[1]),.dout(n1212),.clk(gclk));
	jor g01011(.dina(w_n1211_0[1]),.dinb(w_asqrt58_40[0]),.dout(n1213),.clk(gclk));
	jxor g01012(.dina(w_n1042_0[0]),.dinb(w_n515_67[1]),.dout(n1214),.clk(gclk));
	jand g01013(.dina(n1214),.dinb(w_asqrt52_41[1]),.dout(n1215),.clk(gclk));
	jxor g01014(.dina(n1215),.dinb(w_n1047_0[0]),.dout(n1216),.clk(gclk));
	jnot g01015(.din(w_n1216_0[1]),.dout(n1217),.clk(gclk));
	jand g01016(.dina(w_n1217_0[1]),.dinb(n1213),.dout(n1218),.clk(gclk));
	jor g01017(.dina(n1218),.dinb(w_n1212_0[1]),.dout(n1219),.clk(gclk));
	jand g01018(.dina(w_n1219_0[2]),.dinb(w_asqrt59_40[0]),.dout(n1220),.clk(gclk));
	jor g01019(.dina(w_n1219_0[1]),.dinb(w_asqrt59_39[2]),.dout(n1221),.clk(gclk));
	jxor g01020(.dina(w_n1049_0[0]),.dinb(w_n443_67[1]),.dout(n1222),.clk(gclk));
	jand g01021(.dina(n1222),.dinb(w_asqrt52_41[0]),.dout(n1223),.clk(gclk));
	jxor g01022(.dina(n1223),.dinb(w_n1054_0[0]),.dout(n1224),.clk(gclk));
	jand g01023(.dina(w_n1224_0[1]),.dinb(n1221),.dout(n1225),.clk(gclk));
	jor g01024(.dina(n1225),.dinb(w_n1220_0[1]),.dout(n1226),.clk(gclk));
	jand g01025(.dina(w_n1226_0[2]),.dinb(w_asqrt60_40[1]),.dout(n1227),.clk(gclk));
	jor g01026(.dina(w_n1226_0[1]),.dinb(w_asqrt60_40[0]),.dout(n1228),.clk(gclk));
	jxor g01027(.dina(w_n1057_0[0]),.dinb(w_n352_67[2]),.dout(n1229),.clk(gclk));
	jand g01028(.dina(n1229),.dinb(w_asqrt52_40[2]),.dout(n1230),.clk(gclk));
	jxor g01029(.dina(n1230),.dinb(w_n1062_0[0]),.dout(n1231),.clk(gclk));
	jand g01030(.dina(w_n1231_0[1]),.dinb(n1228),.dout(n1232),.clk(gclk));
	jor g01031(.dina(n1232),.dinb(w_n1227_0[1]),.dout(n1233),.clk(gclk));
	jand g01032(.dina(w_n1233_0[2]),.dinb(w_asqrt61_40[1]),.dout(n1234),.clk(gclk));
	jor g01033(.dina(w_n1233_0[1]),.dinb(w_asqrt61_40[0]),.dout(n1235),.clk(gclk));
	jxor g01034(.dina(w_n1065_0[0]),.dinb(w_n294_68[0]),.dout(n1236),.clk(gclk));
	jand g01035(.dina(n1236),.dinb(w_asqrt52_40[1]),.dout(n1237),.clk(gclk));
	jxor g01036(.dina(n1237),.dinb(w_n1070_0[0]),.dout(n1238),.clk(gclk));
	jand g01037(.dina(w_n1238_0[1]),.dinb(n1235),.dout(n1239),.clk(gclk));
	jor g01038(.dina(n1239),.dinb(w_n1234_0[1]),.dout(n1240),.clk(gclk));
	jand g01039(.dina(w_n1240_0[2]),.dinb(w_asqrt62_40[1]),.dout(n1241),.clk(gclk));
	jor g01040(.dina(w_n1240_0[1]),.dinb(w_asqrt62_40[0]),.dout(n1242),.clk(gclk));
	jxor g01041(.dina(w_n1073_0[0]),.dinb(w_n239_68[0]),.dout(n1243),.clk(gclk));
	jand g01042(.dina(n1243),.dinb(w_asqrt52_40[0]),.dout(n1244),.clk(gclk));
	jxor g01043(.dina(n1244),.dinb(w_n1078_0[0]),.dout(n1245),.clk(gclk));
	jnot g01044(.din(w_n1245_0[1]),.dout(n1246),.clk(gclk));
	jand g01045(.dina(w_n1246_0[1]),.dinb(n1242),.dout(n1247),.clk(gclk));
	jor g01046(.dina(n1247),.dinb(w_n1241_0[1]),.dout(n1248),.clk(gclk));
	jxor g01047(.dina(w_n1080_0[0]),.dinb(w_n221_68[1]),.dout(n1249),.clk(gclk));
	jand g01048(.dina(n1249),.dinb(w_asqrt52_39[2]),.dout(n1250),.clk(gclk));
	jxor g01049(.dina(n1250),.dinb(w_n1086_0[0]),.dout(n1251),.clk(gclk));
	jnot g01050(.din(w_n1251_0[1]),.dout(n1252),.clk(gclk));
	jor g01051(.dina(w_n1252_0[1]),.dinb(w_n1248_0[1]),.dout(n1253),.clk(gclk));
	jnot g01052(.din(w_n1253_1[1]),.dout(n1254),.clk(gclk));
	jnot g01053(.din(w_n1241_0[0]),.dout(n1256),.clk(gclk));
	jnot g01054(.din(w_n1234_0[0]),.dout(n1257),.clk(gclk));
	jnot g01055(.din(w_n1227_0[0]),.dout(n1258),.clk(gclk));
	jnot g01056(.din(w_n1220_0[0]),.dout(n1259),.clk(gclk));
	jnot g01057(.din(w_n1212_0[0]),.dout(n1260),.clk(gclk));
	jnot g01058(.din(w_n1204_0[0]),.dout(n1261),.clk(gclk));
	jnot g01059(.din(w_n1196_0[0]),.dout(n1262),.clk(gclk));
	jnot g01060(.din(w_n1189_0[0]),.dout(n1263),.clk(gclk));
	jnot g01061(.din(w_n1178_0[0]),.dout(n1264),.clk(gclk));
	jnot g01062(.din(w_n1114_0[0]),.dout(n1265),.clk(gclk));
	jnot g01063(.din(w_n1111_0[0]),.dout(n1266),.clk(gclk));
	jor g01064(.dina(w_n1173_64[1]),.dinb(w_n1010_0[2]),.dout(n1267),.clk(gclk));
	jand g01065(.dina(n1267),.dinb(n1266),.dout(n1268),.clk(gclk));
	jand g01066(.dina(n1268),.dinb(w_n1008_66[0]),.dout(n1269),.clk(gclk));
	jor g01067(.dina(w_n1173_64[0]),.dinb(w_a104_0[0]),.dout(n1270),.clk(gclk));
	jand g01068(.dina(n1270),.dinb(w_a105_0[0]),.dout(n1271),.clk(gclk));
	jor g01069(.dina(w_n1180_0[0]),.dinb(n1271),.dout(n1272),.clk(gclk));
	jor g01070(.dina(n1272),.dinb(n1269),.dout(n1273),.clk(gclk));
	jand g01071(.dina(n1273),.dinb(n1265),.dout(n1274),.clk(gclk));
	jand g01072(.dina(n1274),.dinb(w_n884_65[0]),.dout(n1275),.clk(gclk));
	jor g01073(.dina(w_n1185_0[0]),.dinb(n1275),.dout(n1276),.clk(gclk));
	jand g01074(.dina(n1276),.dinb(n1264),.dout(n1277),.clk(gclk));
	jand g01075(.dina(n1277),.dinb(w_n743_66[0]),.dout(n1278),.clk(gclk));
	jnot g01076(.din(w_n1193_0[0]),.dout(n1279),.clk(gclk));
	jor g01077(.dina(w_n1279_0[1]),.dinb(n1278),.dout(n1280),.clk(gclk));
	jand g01078(.dina(n1280),.dinb(n1263),.dout(n1281),.clk(gclk));
	jand g01079(.dina(n1281),.dinb(w_n635_66[0]),.dout(n1282),.clk(gclk));
	jor g01080(.dina(w_n1200_0[0]),.dinb(n1282),.dout(n1283),.clk(gclk));
	jand g01081(.dina(n1283),.dinb(n1262),.dout(n1284),.clk(gclk));
	jand g01082(.dina(n1284),.dinb(w_n515_67[0]),.dout(n1285),.clk(gclk));
	jor g01083(.dina(w_n1208_0[0]),.dinb(n1285),.dout(n1286),.clk(gclk));
	jand g01084(.dina(n1286),.dinb(n1261),.dout(n1287),.clk(gclk));
	jand g01085(.dina(n1287),.dinb(w_n443_67[0]),.dout(n1288),.clk(gclk));
	jor g01086(.dina(w_n1216_0[0]),.dinb(n1288),.dout(n1289),.clk(gclk));
	jand g01087(.dina(n1289),.dinb(n1260),.dout(n1290),.clk(gclk));
	jand g01088(.dina(n1290),.dinb(w_n352_67[1]),.dout(n1291),.clk(gclk));
	jnot g01089(.din(w_n1224_0[0]),.dout(n1292),.clk(gclk));
	jor g01090(.dina(w_n1292_0[1]),.dinb(n1291),.dout(n1293),.clk(gclk));
	jand g01091(.dina(n1293),.dinb(n1259),.dout(n1294),.clk(gclk));
	jand g01092(.dina(n1294),.dinb(w_n294_67[2]),.dout(n1295),.clk(gclk));
	jnot g01093(.din(w_n1231_0[0]),.dout(n1296),.clk(gclk));
	jor g01094(.dina(w_n1296_0[1]),.dinb(n1295),.dout(n1297),.clk(gclk));
	jand g01095(.dina(n1297),.dinb(n1258),.dout(n1298),.clk(gclk));
	jand g01096(.dina(n1298),.dinb(w_n239_67[2]),.dout(n1299),.clk(gclk));
	jnot g01097(.din(w_n1238_0[0]),.dout(n1300),.clk(gclk));
	jor g01098(.dina(w_n1300_0[1]),.dinb(n1299),.dout(n1301),.clk(gclk));
	jand g01099(.dina(n1301),.dinb(n1257),.dout(n1302),.clk(gclk));
	jand g01100(.dina(n1302),.dinb(w_n221_68[0]),.dout(n1303),.clk(gclk));
	jor g01101(.dina(w_n1245_0[0]),.dinb(n1303),.dout(n1304),.clk(gclk));
	jand g01102(.dina(n1304),.dinb(n1256),.dout(n1305),.clk(gclk));
	jor g01103(.dina(w_n1251_0[0]),.dinb(w_n1305_0[1]),.dout(n1306),.clk(gclk));
	jxor g01104(.dina(w_n1091_0[1]),.dinb(w_n1088_0[2]),.dout(n1307),.clk(gclk));
	jnot g01105(.din(w_n1307_0[1]),.dout(n1308),.clk(gclk));
	jand g01106(.dina(n1308),.dinb(w_asqrt52_39[1]),.dout(n1309),.clk(gclk));
	jor g01107(.dina(w_n1309_0[1]),.dinb(w_n1306_0[1]),.dout(n1310),.clk(gclk));
	jand g01108(.dina(n1310),.dinb(w_n218_28[0]),.dout(n1311),.clk(gclk));
	jand g01109(.dina(w_n1172_0[0]),.dinb(w_n1088_0[1]),.dout(n1312),.clk(gclk));
	jnot g01110(.din(n1312),.dout(n1313),.clk(gclk));
	jand g01111(.dina(w_n1307_0[0]),.dinb(w_asqrt63_52[0]),.dout(n1314),.clk(gclk));
	jand g01112(.dina(w_n1314_0[1]),.dinb(n1313),.dout(n1315),.clk(gclk));
	jor g01113(.dina(w_n1315_0[1]),.dinb(w_n1311_0[1]),.dout(n1316),.clk(gclk));
	jor g01114(.dina(w_n1316_0[1]),.dinb(w_n1254_0[2]),.dout(asqrt_fa_52),.clk(gclk));
	jnot g01115(.din(w_a100_0[2]),.dout(n1319),.clk(gclk));
	jnot g01116(.din(w_a101_0[1]),.dout(n1320),.clk(gclk));
	jand g01117(.dina(w_n1320_0[1]),.dinb(w_n1319_1[2]),.dout(n1321),.clk(gclk));
	jand g01118(.dina(w_n1321_0[2]),.dinb(w_n1108_1[0]),.dout(n1322),.clk(gclk));
	jnot g01119(.din(w_n1322_0[1]),.dout(n1323),.clk(gclk));
	jand g01120(.dina(w_n1252_0[0]),.dinb(w_n1248_0[0]),.dout(n1325),.clk(gclk));
	jnot g01121(.din(w_n1309_0[0]),.dout(n1326),.clk(gclk));
	jand g01122(.dina(n1326),.dinb(w_n1325_0[1]),.dout(n1327),.clk(gclk));
	jor g01123(.dina(n1327),.dinb(w_asqrt63_51[2]),.dout(n1328),.clk(gclk));
	jnot g01124(.din(w_n1315_0[0]),.dout(n1329),.clk(gclk));
	jand g01125(.dina(n1329),.dinb(n1328),.dout(n1330),.clk(gclk));
	jand g01126(.dina(w_n1330_0[1]),.dinb(w_n1253_1[0]),.dout(n1332),.clk(gclk));
	jor g01127(.dina(w_n1332_67[2]),.dinb(w_n1108_0[2]),.dout(n1333),.clk(gclk));
	jand g01128(.dina(n1333),.dinb(n1323),.dout(n1334),.clk(gclk));
	jor g01129(.dina(w_n1334_0[2]),.dinb(w_n1173_63[2]),.dout(n1335),.clk(gclk));
	jand g01130(.dina(w_n1334_0[1]),.dinb(w_n1173_63[1]),.dout(n1336),.clk(gclk));
	jor g01131(.dina(w_n1332_67[1]),.dinb(w_a102_1[0]),.dout(n1337),.clk(gclk));
	jand g01132(.dina(n1337),.dinb(w_a103_0[0]),.dout(n1338),.clk(gclk));
	jand g01133(.dina(w_asqrt51_38[1]),.dinb(w_n1110_0[1]),.dout(n1339),.clk(gclk));
	jor g01134(.dina(n1339),.dinb(n1338),.dout(n1340),.clk(gclk));
	jor g01135(.dina(n1340),.dinb(n1336),.dout(n1341),.clk(gclk));
	jand g01136(.dina(n1341),.dinb(w_n1335_0[1]),.dout(n1342),.clk(gclk));
	jor g01137(.dina(w_n1342_0[2]),.dinb(w_n1008_65[2]),.dout(n1343),.clk(gclk));
	jand g01138(.dina(w_n1342_0[1]),.dinb(w_n1008_65[1]),.dout(n1344),.clk(gclk));
	jnot g01139(.din(w_n1110_0[0]),.dout(n1345),.clk(gclk));
	jor g01140(.dina(w_n1332_67[0]),.dinb(n1345),.dout(n1346),.clk(gclk));
	jor g01141(.dina(w_n1314_0[0]),.dinb(w_n1254_0[1]),.dout(n1347),.clk(gclk));
	jor g01142(.dina(n1347),.dinb(w_n1311_0[0]),.dout(n1348),.clk(gclk));
	jor g01143(.dina(n1348),.dinb(w_n1173_63[0]),.dout(n1349),.clk(gclk));
	jand g01144(.dina(n1349),.dinb(w_n1346_0[1]),.dout(n1350),.clk(gclk));
	jxor g01145(.dina(n1350),.dinb(w_n1010_0[1]),.dout(n1351),.clk(gclk));
	jor g01146(.dina(w_n1351_0[2]),.dinb(n1344),.dout(n1352),.clk(gclk));
	jand g01147(.dina(n1352),.dinb(w_n1343_0[1]),.dout(n1353),.clk(gclk));
	jor g01148(.dina(w_n1353_0[2]),.dinb(w_n884_64[2]),.dout(n1354),.clk(gclk));
	jand g01149(.dina(w_n1353_0[1]),.dinb(w_n884_64[1]),.dout(n1355),.clk(gclk));
	jxor g01150(.dina(w_n1113_0[0]),.dinb(w_n1008_65[0]),.dout(n1356),.clk(gclk));
	jor g01151(.dina(n1356),.dinb(w_n1332_66[2]),.dout(n1357),.clk(gclk));
	jxor g01152(.dina(n1357),.dinb(w_n1175_0[0]),.dout(n1358),.clk(gclk));
	jor g01153(.dina(w_n1358_0[2]),.dinb(n1355),.dout(n1359),.clk(gclk));
	jand g01154(.dina(n1359),.dinb(w_n1354_0[1]),.dout(n1360),.clk(gclk));
	jor g01155(.dina(w_n1360_0[2]),.dinb(w_n743_65[2]),.dout(n1361),.clk(gclk));
	jand g01156(.dina(w_n1360_0[1]),.dinb(w_n743_65[1]),.dout(n1362),.clk(gclk));
	jxor g01157(.dina(w_n1177_0[0]),.dinb(w_n884_64[0]),.dout(n1363),.clk(gclk));
	jor g01158(.dina(n1363),.dinb(w_n1332_66[1]),.dout(n1364),.clk(gclk));
	jxor g01159(.dina(n1364),.dinb(w_n1186_0[0]),.dout(n1365),.clk(gclk));
	jor g01160(.dina(w_n1365_0[2]),.dinb(n1362),.dout(n1366),.clk(gclk));
	jand g01161(.dina(n1366),.dinb(w_n1361_0[1]),.dout(n1367),.clk(gclk));
	jor g01162(.dina(w_n1367_0[2]),.dinb(w_n635_65[2]),.dout(n1368),.clk(gclk));
	jand g01163(.dina(w_n1367_0[1]),.dinb(w_n635_65[1]),.dout(n1369),.clk(gclk));
	jxor g01164(.dina(w_n1188_0[0]),.dinb(w_n743_65[0]),.dout(n1370),.clk(gclk));
	jor g01165(.dina(n1370),.dinb(w_n1332_66[0]),.dout(n1371),.clk(gclk));
	jxor g01166(.dina(n1371),.dinb(w_n1279_0[0]),.dout(n1372),.clk(gclk));
	jnot g01167(.din(w_n1372_0[2]),.dout(n1373),.clk(gclk));
	jor g01168(.dina(n1373),.dinb(n1369),.dout(n1374),.clk(gclk));
	jand g01169(.dina(n1374),.dinb(w_n1368_0[1]),.dout(n1375),.clk(gclk));
	jor g01170(.dina(w_n1375_0[2]),.dinb(w_n515_66[2]),.dout(n1376),.clk(gclk));
	jand g01171(.dina(w_n1375_0[1]),.dinb(w_n515_66[1]),.dout(n1377),.clk(gclk));
	jxor g01172(.dina(w_n1195_0[0]),.dinb(w_n635_65[0]),.dout(n1378),.clk(gclk));
	jor g01173(.dina(n1378),.dinb(w_n1332_65[2]),.dout(n1379),.clk(gclk));
	jxor g01174(.dina(n1379),.dinb(w_n1201_0[0]),.dout(n1380),.clk(gclk));
	jor g01175(.dina(w_n1380_0[2]),.dinb(n1377),.dout(n1381),.clk(gclk));
	jand g01176(.dina(n1381),.dinb(w_n1376_0[1]),.dout(n1382),.clk(gclk));
	jor g01177(.dina(w_n1382_0[2]),.dinb(w_n443_66[2]),.dout(n1383),.clk(gclk));
	jand g01178(.dina(w_n1382_0[1]),.dinb(w_n443_66[1]),.dout(n1384),.clk(gclk));
	jxor g01179(.dina(w_n1203_0[0]),.dinb(w_n515_66[0]),.dout(n1385),.clk(gclk));
	jor g01180(.dina(n1385),.dinb(w_n1332_65[1]),.dout(n1386),.clk(gclk));
	jxor g01181(.dina(n1386),.dinb(w_n1209_0[0]),.dout(n1387),.clk(gclk));
	jor g01182(.dina(w_n1387_0[2]),.dinb(n1384),.dout(n1388),.clk(gclk));
	jand g01183(.dina(n1388),.dinb(w_n1383_0[1]),.dout(n1389),.clk(gclk));
	jor g01184(.dina(w_n1389_0[2]),.dinb(w_n352_67[0]),.dout(n1390),.clk(gclk));
	jand g01185(.dina(w_n1389_0[1]),.dinb(w_n352_66[2]),.dout(n1391),.clk(gclk));
	jxor g01186(.dina(w_n1211_0[0]),.dinb(w_n443_66[0]),.dout(n1392),.clk(gclk));
	jor g01187(.dina(n1392),.dinb(w_n1332_65[0]),.dout(n1393),.clk(gclk));
	jxor g01188(.dina(n1393),.dinb(w_n1217_0[0]),.dout(n1394),.clk(gclk));
	jor g01189(.dina(w_n1394_0[2]),.dinb(n1391),.dout(n1395),.clk(gclk));
	jand g01190(.dina(n1395),.dinb(w_n1390_0[1]),.dout(n1396),.clk(gclk));
	jor g01191(.dina(w_n1396_0[2]),.dinb(w_n294_67[1]),.dout(n1397),.clk(gclk));
	jand g01192(.dina(w_n1396_0[1]),.dinb(w_n294_67[0]),.dout(n1398),.clk(gclk));
	jxor g01193(.dina(w_n1219_0[0]),.dinb(w_n352_66[1]),.dout(n1399),.clk(gclk));
	jor g01194(.dina(n1399),.dinb(w_n1332_64[2]),.dout(n1400),.clk(gclk));
	jxor g01195(.dina(n1400),.dinb(w_n1292_0[0]),.dout(n1401),.clk(gclk));
	jnot g01196(.din(w_n1401_0[2]),.dout(n1402),.clk(gclk));
	jor g01197(.dina(n1402),.dinb(n1398),.dout(n1403),.clk(gclk));
	jand g01198(.dina(n1403),.dinb(w_n1397_0[1]),.dout(n1404),.clk(gclk));
	jor g01199(.dina(w_n1404_0[2]),.dinb(w_n239_67[1]),.dout(n1405),.clk(gclk));
	jand g01200(.dina(w_n1404_0[1]),.dinb(w_n239_67[0]),.dout(n1406),.clk(gclk));
	jxor g01201(.dina(w_n1226_0[0]),.dinb(w_n294_66[2]),.dout(n1407),.clk(gclk));
	jor g01202(.dina(n1407),.dinb(w_n1332_64[1]),.dout(n1408),.clk(gclk));
	jxor g01203(.dina(n1408),.dinb(w_n1296_0[0]),.dout(n1409),.clk(gclk));
	jnot g01204(.din(w_n1409_0[2]),.dout(n1410),.clk(gclk));
	jor g01205(.dina(n1410),.dinb(n1406),.dout(n1411),.clk(gclk));
	jand g01206(.dina(n1411),.dinb(w_n1405_0[1]),.dout(n1412),.clk(gclk));
	jor g01207(.dina(w_n1412_0[2]),.dinb(w_n221_67[2]),.dout(n1413),.clk(gclk));
	jand g01208(.dina(w_n1412_0[1]),.dinb(w_n221_67[1]),.dout(n1414),.clk(gclk));
	jxor g01209(.dina(w_n1233_0[0]),.dinb(w_n239_66[2]),.dout(n1415),.clk(gclk));
	jor g01210(.dina(n1415),.dinb(w_n1332_64[0]),.dout(n1416),.clk(gclk));
	jxor g01211(.dina(n1416),.dinb(w_n1300_0[0]),.dout(n1417),.clk(gclk));
	jnot g01212(.din(w_n1417_0[1]),.dout(n1418),.clk(gclk));
	jor g01213(.dina(w_n1418_0[1]),.dinb(n1414),.dout(n1419),.clk(gclk));
	jand g01214(.dina(n1419),.dinb(w_n1413_0[1]),.dout(n1420),.clk(gclk));
	jxor g01215(.dina(w_n1240_0[0]),.dinb(w_n221_67[0]),.dout(n1421),.clk(gclk));
	jor g01216(.dina(n1421),.dinb(w_n1332_63[2]),.dout(n1422),.clk(gclk));
	jxor g01217(.dina(n1422),.dinb(w_n1246_0[0]),.dout(n1423),.clk(gclk));
	jand g01218(.dina(w_n1423_1[2]),.dinb(w_n1420_1[1]),.dout(n1424),.clk(gclk));
	jand g01219(.dina(w_n1316_0[0]),.dinb(w_n1325_0[0]),.dout(n1426),.clk(gclk));
	jor g01220(.dina(w_n1423_1[1]),.dinb(w_n1420_1[0]),.dout(n1427),.clk(gclk));
	jor g01221(.dina(n1427),.dinb(w_n1254_0[0]),.dout(n1428),.clk(gclk));
	jor g01222(.dina(n1428),.dinb(w_n1426_0[1]),.dout(n1429),.clk(gclk));
	jand g01223(.dina(n1429),.dinb(w_n218_27[2]),.dout(n1430),.clk(gclk));
	jand g01224(.dina(w_n1330_0[0]),.dinb(w_n1305_0[0]),.dout(n1431),.clk(gclk));
	jand g01225(.dina(w_n1306_0[0]),.dinb(w_asqrt63_51[1]),.dout(n1432),.clk(gclk));
	jand g01226(.dina(n1432),.dinb(w_n1253_0[2]),.dout(n1433),.clk(gclk));
	jnot g01227(.din(n1433),.dout(n1434),.clk(gclk));
	jor g01228(.dina(w_n1434_0[1]),.dinb(n1431),.dout(n1435),.clk(gclk));
	jnot g01229(.din(w_n1435_0[1]),.dout(n1436),.clk(gclk));
	jor g01230(.dina(n1436),.dinb(n1430),.dout(n1437),.clk(gclk));
	jor g01231(.dina(n1437),.dinb(w_n1424_0[1]),.dout(asqrt_fa_51),.clk(gclk));
	jnot g01232(.din(w_a98_1[1]),.dout(n1440),.clk(gclk));
	jnot g01233(.din(w_a99_0[1]),.dout(n1441),.clk(gclk));
	jand g01234(.dina(w_n1441_0[1]),.dinb(w_n1440_1[1]),.dout(n1442),.clk(gclk));
	jand g01235(.dina(w_n1442_0[2]),.dinb(w_n1319_1[1]),.dout(n1443),.clk(gclk));
	jand g01236(.dina(w_asqrt50_43),.dinb(w_a100_0[1]),.dout(n1444),.clk(gclk));
	jor g01237(.dina(n1444),.dinb(w_n1443_0[1]),.dout(n1445),.clk(gclk));
	jand g01238(.dina(w_n1445_0[2]),.dinb(w_asqrt51_38[0]),.dout(n1446),.clk(gclk));
	jor g01239(.dina(w_n1445_0[1]),.dinb(w_asqrt51_37[2]),.dout(n1447),.clk(gclk));
	jand g01240(.dina(w_asqrt50_42[2]),.dinb(w_n1319_1[0]),.dout(n1448),.clk(gclk));
	jor g01241(.dina(n1448),.dinb(w_n1320_0[0]),.dout(n1449),.clk(gclk));
	jnot g01242(.din(w_n1321_0[1]),.dout(n1450),.clk(gclk));
	jnot g01243(.din(w_n1424_0[0]),.dout(n1451),.clk(gclk));
	jnot g01244(.din(w_n1426_0[0]),.dout(n1453),.clk(gclk));
	jnot g01245(.din(w_n1413_0[0]),.dout(n1454),.clk(gclk));
	jnot g01246(.din(w_n1405_0[0]),.dout(n1455),.clk(gclk));
	jnot g01247(.din(w_n1397_0[0]),.dout(n1456),.clk(gclk));
	jnot g01248(.din(w_n1390_0[0]),.dout(n1457),.clk(gclk));
	jnot g01249(.din(w_n1383_0[0]),.dout(n1458),.clk(gclk));
	jnot g01250(.din(w_n1376_0[0]),.dout(n1459),.clk(gclk));
	jnot g01251(.din(w_n1368_0[0]),.dout(n1460),.clk(gclk));
	jnot g01252(.din(w_n1361_0[0]),.dout(n1461),.clk(gclk));
	jnot g01253(.din(w_n1354_0[0]),.dout(n1462),.clk(gclk));
	jnot g01254(.din(w_n1343_0[0]),.dout(n1463),.clk(gclk));
	jnot g01255(.din(w_n1335_0[0]),.dout(n1464),.clk(gclk));
	jand g01256(.dina(w_asqrt51_37[1]),.dinb(w_a102_0[2]),.dout(n1465),.clk(gclk));
	jor g01257(.dina(n1465),.dinb(w_n1322_0[0]),.dout(n1466),.clk(gclk));
	jor g01258(.dina(n1466),.dinb(w_asqrt52_39[0]),.dout(n1467),.clk(gclk));
	jand g01259(.dina(w_asqrt51_37[0]),.dinb(w_n1108_0[1]),.dout(n1468),.clk(gclk));
	jor g01260(.dina(n1468),.dinb(w_n1109_0[0]),.dout(n1469),.clk(gclk));
	jand g01261(.dina(w_n1346_0[0]),.dinb(n1469),.dout(n1470),.clk(gclk));
	jand g01262(.dina(w_n1470_0[1]),.dinb(n1467),.dout(n1471),.clk(gclk));
	jor g01263(.dina(n1471),.dinb(n1464),.dout(n1472),.clk(gclk));
	jor g01264(.dina(n1472),.dinb(w_asqrt53_38[0]),.dout(n1473),.clk(gclk));
	jnot g01265(.din(w_n1351_0[1]),.dout(n1474),.clk(gclk));
	jand g01266(.dina(n1474),.dinb(n1473),.dout(n1475),.clk(gclk));
	jor g01267(.dina(n1475),.dinb(n1463),.dout(n1476),.clk(gclk));
	jor g01268(.dina(n1476),.dinb(w_asqrt54_39[0]),.dout(n1477),.clk(gclk));
	jnot g01269(.din(w_n1358_0[1]),.dout(n1478),.clk(gclk));
	jand g01270(.dina(n1478),.dinb(n1477),.dout(n1479),.clk(gclk));
	jor g01271(.dina(n1479),.dinb(n1462),.dout(n1480),.clk(gclk));
	jor g01272(.dina(n1480),.dinb(w_asqrt55_38[1]),.dout(n1481),.clk(gclk));
	jnot g01273(.din(w_n1365_0[1]),.dout(n1482),.clk(gclk));
	jand g01274(.dina(n1482),.dinb(n1481),.dout(n1483),.clk(gclk));
	jor g01275(.dina(n1483),.dinb(n1461),.dout(n1484),.clk(gclk));
	jor g01276(.dina(n1484),.dinb(w_asqrt56_39[1]),.dout(n1485),.clk(gclk));
	jand g01277(.dina(w_n1372_0[1]),.dinb(n1485),.dout(n1486),.clk(gclk));
	jor g01278(.dina(n1486),.dinb(n1460),.dout(n1487),.clk(gclk));
	jor g01279(.dina(n1487),.dinb(w_asqrt57_39[0]),.dout(n1488),.clk(gclk));
	jnot g01280(.din(w_n1380_0[1]),.dout(n1489),.clk(gclk));
	jand g01281(.dina(n1489),.dinb(n1488),.dout(n1490),.clk(gclk));
	jor g01282(.dina(n1490),.dinb(n1459),.dout(n1491),.clk(gclk));
	jor g01283(.dina(n1491),.dinb(w_asqrt58_39[2]),.dout(n1492),.clk(gclk));
	jnot g01284(.din(w_n1387_0[1]),.dout(n1493),.clk(gclk));
	jand g01285(.dina(n1493),.dinb(n1492),.dout(n1494),.clk(gclk));
	jor g01286(.dina(n1494),.dinb(n1458),.dout(n1495),.clk(gclk));
	jor g01287(.dina(n1495),.dinb(w_asqrt59_39[1]),.dout(n1496),.clk(gclk));
	jnot g01288(.din(w_n1394_0[1]),.dout(n1497),.clk(gclk));
	jand g01289(.dina(n1497),.dinb(n1496),.dout(n1498),.clk(gclk));
	jor g01290(.dina(n1498),.dinb(n1457),.dout(n1499),.clk(gclk));
	jor g01291(.dina(n1499),.dinb(w_asqrt60_39[2]),.dout(n1500),.clk(gclk));
	jand g01292(.dina(w_n1401_0[1]),.dinb(n1500),.dout(n1501),.clk(gclk));
	jor g01293(.dina(n1501),.dinb(n1456),.dout(n1502),.clk(gclk));
	jor g01294(.dina(n1502),.dinb(w_asqrt61_39[2]),.dout(n1503),.clk(gclk));
	jand g01295(.dina(w_n1409_0[1]),.dinb(n1503),.dout(n1504),.clk(gclk));
	jor g01296(.dina(n1504),.dinb(n1455),.dout(n1505),.clk(gclk));
	jor g01297(.dina(n1505),.dinb(w_asqrt62_39[2]),.dout(n1506),.clk(gclk));
	jand g01298(.dina(w_n1417_0[0]),.dinb(n1506),.dout(n1507),.clk(gclk));
	jor g01299(.dina(n1507),.dinb(n1454),.dout(n1508),.clk(gclk));
	jnot g01300(.din(w_n1423_1[0]),.dout(n1509),.clk(gclk));
	jand g01301(.dina(n1509),.dinb(n1508),.dout(n1510),.clk(gclk));
	jand g01302(.dina(n1510),.dinb(w_n1253_0[1]),.dout(n1511),.clk(gclk));
	jand g01303(.dina(n1511),.dinb(n1453),.dout(n1512),.clk(gclk));
	jor g01304(.dina(n1512),.dinb(w_asqrt63_51[0]),.dout(n1513),.clk(gclk));
	jand g01305(.dina(w_n1435_0[0]),.dinb(w_n1513_0[1]),.dout(n1514),.clk(gclk));
	jand g01306(.dina(w_n1514_0[1]),.dinb(w_n1451_0[1]),.dout(n1516),.clk(gclk));
	jor g01307(.dina(w_n1516_62[2]),.dinb(n1450),.dout(n1517),.clk(gclk));
	jand g01308(.dina(n1517),.dinb(n1449),.dout(n1518),.clk(gclk));
	jand g01309(.dina(w_n1518_0[1]),.dinb(n1447),.dout(n1519),.clk(gclk));
	jor g01310(.dina(n1519),.dinb(w_n1446_0[1]),.dout(n1520),.clk(gclk));
	jand g01311(.dina(w_n1520_0[2]),.dinb(w_asqrt52_38[2]),.dout(n1521),.clk(gclk));
	jor g01312(.dina(w_n1520_0[1]),.dinb(w_asqrt52_38[1]),.dout(n1522),.clk(gclk));
	jand g01313(.dina(w_asqrt50_42[1]),.dinb(w_n1321_0[0]),.dout(n1523),.clk(gclk));
	jand g01314(.dina(w_n1451_0[0]),.dinb(w_asqrt51_36[2]),.dout(n1524),.clk(gclk));
	jand g01315(.dina(n1524),.dinb(w_n1434_0[0]),.dout(n1525),.clk(gclk));
	jand g01316(.dina(n1525),.dinb(w_n1513_0[0]),.dout(n1526),.clk(gclk));
	jor g01317(.dina(n1526),.dinb(w_n1523_0[1]),.dout(n1527),.clk(gclk));
	jxor g01318(.dina(n1527),.dinb(w_a102_0[1]),.dout(n1528),.clk(gclk));
	jnot g01319(.din(w_n1528_0[2]),.dout(n1529),.clk(gclk));
	jand g01320(.dina(n1529),.dinb(n1522),.dout(n1530),.clk(gclk));
	jor g01321(.dina(n1530),.dinb(w_n1521_0[1]),.dout(n1531),.clk(gclk));
	jand g01322(.dina(w_n1531_0[2]),.dinb(w_asqrt53_37[2]),.dout(n1532),.clk(gclk));
	jor g01323(.dina(w_n1531_0[1]),.dinb(w_asqrt53_37[1]),.dout(n1533),.clk(gclk));
	jxor g01324(.dina(w_n1334_0[0]),.dinb(w_n1173_62[2]),.dout(n1534),.clk(gclk));
	jand g01325(.dina(n1534),.dinb(w_asqrt50_42[0]),.dout(n1535),.clk(gclk));
	jxor g01326(.dina(n1535),.dinb(w_n1470_0[0]),.dout(n1536),.clk(gclk));
	jand g01327(.dina(w_n1536_0[1]),.dinb(n1533),.dout(n1537),.clk(gclk));
	jor g01328(.dina(n1537),.dinb(w_n1532_0[1]),.dout(n1538),.clk(gclk));
	jand g01329(.dina(w_n1538_0[2]),.dinb(w_asqrt54_38[2]),.dout(n1539),.clk(gclk));
	jor g01330(.dina(w_n1538_0[1]),.dinb(w_asqrt54_38[1]),.dout(n1540),.clk(gclk));
	jxor g01331(.dina(w_n1342_0[0]),.dinb(w_n1008_64[2]),.dout(n1541),.clk(gclk));
	jand g01332(.dina(n1541),.dinb(w_asqrt50_41[2]),.dout(n1542),.clk(gclk));
	jxor g01333(.dina(n1542),.dinb(w_n1351_0[0]),.dout(n1543),.clk(gclk));
	jnot g01334(.din(w_n1543_0[1]),.dout(n1544),.clk(gclk));
	jand g01335(.dina(w_n1544_0[1]),.dinb(n1540),.dout(n1545),.clk(gclk));
	jor g01336(.dina(n1545),.dinb(w_n1539_0[1]),.dout(n1546),.clk(gclk));
	jand g01337(.dina(w_n1546_0[2]),.dinb(w_asqrt55_38[0]),.dout(n1547),.clk(gclk));
	jor g01338(.dina(w_n1546_0[1]),.dinb(w_asqrt55_37[2]),.dout(n1548),.clk(gclk));
	jxor g01339(.dina(w_n1353_0[0]),.dinb(w_n884_63[2]),.dout(n1549),.clk(gclk));
	jand g01340(.dina(n1549),.dinb(w_asqrt50_41[1]),.dout(n1550),.clk(gclk));
	jxor g01341(.dina(n1550),.dinb(w_n1358_0[0]),.dout(n1551),.clk(gclk));
	jnot g01342(.din(w_n1551_0[1]),.dout(n1552),.clk(gclk));
	jand g01343(.dina(w_n1552_0[1]),.dinb(n1548),.dout(n1553),.clk(gclk));
	jor g01344(.dina(n1553),.dinb(w_n1547_0[1]),.dout(n1554),.clk(gclk));
	jand g01345(.dina(w_n1554_0[2]),.dinb(w_asqrt56_39[0]),.dout(n1555),.clk(gclk));
	jor g01346(.dina(w_n1554_0[1]),.dinb(w_asqrt56_38[2]),.dout(n1556),.clk(gclk));
	jxor g01347(.dina(w_n1360_0[0]),.dinb(w_n743_64[2]),.dout(n1557),.clk(gclk));
	jand g01348(.dina(n1557),.dinb(w_asqrt50_41[0]),.dout(n1558),.clk(gclk));
	jxor g01349(.dina(n1558),.dinb(w_n1365_0[0]),.dout(n1559),.clk(gclk));
	jnot g01350(.din(w_n1559_0[1]),.dout(n1560),.clk(gclk));
	jand g01351(.dina(w_n1560_0[1]),.dinb(n1556),.dout(n1561),.clk(gclk));
	jor g01352(.dina(n1561),.dinb(w_n1555_0[1]),.dout(n1562),.clk(gclk));
	jand g01353(.dina(w_n1562_0[2]),.dinb(w_asqrt57_38[2]),.dout(n1563),.clk(gclk));
	jor g01354(.dina(w_n1562_0[1]),.dinb(w_asqrt57_38[1]),.dout(n1564),.clk(gclk));
	jxor g01355(.dina(w_n1367_0[0]),.dinb(w_n635_64[2]),.dout(n1565),.clk(gclk));
	jand g01356(.dina(n1565),.dinb(w_asqrt50_40[2]),.dout(n1566),.clk(gclk));
	jxor g01357(.dina(n1566),.dinb(w_n1372_0[0]),.dout(n1567),.clk(gclk));
	jand g01358(.dina(w_n1567_0[1]),.dinb(n1564),.dout(n1568),.clk(gclk));
	jor g01359(.dina(n1568),.dinb(w_n1563_0[1]),.dout(n1569),.clk(gclk));
	jand g01360(.dina(w_n1569_0[2]),.dinb(w_asqrt58_39[1]),.dout(n1570),.clk(gclk));
	jor g01361(.dina(w_n1569_0[1]),.dinb(w_asqrt58_39[0]),.dout(n1571),.clk(gclk));
	jxor g01362(.dina(w_n1375_0[0]),.dinb(w_n515_65[2]),.dout(n1572),.clk(gclk));
	jand g01363(.dina(n1572),.dinb(w_asqrt50_40[1]),.dout(n1573),.clk(gclk));
	jxor g01364(.dina(n1573),.dinb(w_n1380_0[0]),.dout(n1574),.clk(gclk));
	jnot g01365(.din(w_n1574_0[1]),.dout(n1575),.clk(gclk));
	jand g01366(.dina(w_n1575_0[1]),.dinb(n1571),.dout(n1576),.clk(gclk));
	jor g01367(.dina(n1576),.dinb(w_n1570_0[1]),.dout(n1577),.clk(gclk));
	jand g01368(.dina(w_n1577_0[2]),.dinb(w_asqrt59_39[0]),.dout(n1578),.clk(gclk));
	jor g01369(.dina(w_n1577_0[1]),.dinb(w_asqrt59_38[2]),.dout(n1579),.clk(gclk));
	jxor g01370(.dina(w_n1382_0[0]),.dinb(w_n443_65[2]),.dout(n1580),.clk(gclk));
	jand g01371(.dina(n1580),.dinb(w_asqrt50_40[0]),.dout(n1581),.clk(gclk));
	jxor g01372(.dina(n1581),.dinb(w_n1387_0[0]),.dout(n1582),.clk(gclk));
	jnot g01373(.din(w_n1582_0[1]),.dout(n1583),.clk(gclk));
	jand g01374(.dina(w_n1583_0[1]),.dinb(n1579),.dout(n1584),.clk(gclk));
	jor g01375(.dina(n1584),.dinb(w_n1578_0[1]),.dout(n1585),.clk(gclk));
	jand g01376(.dina(w_n1585_0[2]),.dinb(w_asqrt60_39[1]),.dout(n1586),.clk(gclk));
	jor g01377(.dina(w_n1585_0[1]),.dinb(w_asqrt60_39[0]),.dout(n1587),.clk(gclk));
	jxor g01378(.dina(w_n1389_0[0]),.dinb(w_n352_66[0]),.dout(n1588),.clk(gclk));
	jand g01379(.dina(n1588),.dinb(w_asqrt50_39[2]),.dout(n1589),.clk(gclk));
	jxor g01380(.dina(n1589),.dinb(w_n1394_0[0]),.dout(n1590),.clk(gclk));
	jnot g01381(.din(w_n1590_0[1]),.dout(n1591),.clk(gclk));
	jand g01382(.dina(w_n1591_0[1]),.dinb(n1587),.dout(n1592),.clk(gclk));
	jor g01383(.dina(n1592),.dinb(w_n1586_0[1]),.dout(n1593),.clk(gclk));
	jand g01384(.dina(w_n1593_0[2]),.dinb(w_asqrt61_39[1]),.dout(n1594),.clk(gclk));
	jor g01385(.dina(w_n1593_0[1]),.dinb(w_asqrt61_39[0]),.dout(n1595),.clk(gclk));
	jxor g01386(.dina(w_n1396_0[0]),.dinb(w_n294_66[1]),.dout(n1596),.clk(gclk));
	jand g01387(.dina(n1596),.dinb(w_asqrt50_39[1]),.dout(n1597),.clk(gclk));
	jxor g01388(.dina(n1597),.dinb(w_n1401_0[0]),.dout(n1598),.clk(gclk));
	jand g01389(.dina(w_n1598_0[1]),.dinb(n1595),.dout(n1599),.clk(gclk));
	jor g01390(.dina(n1599),.dinb(w_n1594_0[1]),.dout(n1600),.clk(gclk));
	jand g01391(.dina(w_n1600_0[2]),.dinb(w_asqrt62_39[1]),.dout(n1601),.clk(gclk));
	jnot g01392(.din(w_n1601_0[1]),.dout(n1602),.clk(gclk));
	jnot g01393(.din(w_n1594_0[0]),.dout(n1603),.clk(gclk));
	jnot g01394(.din(w_n1586_0[0]),.dout(n1604),.clk(gclk));
	jnot g01395(.din(w_n1578_0[0]),.dout(n1605),.clk(gclk));
	jnot g01396(.din(w_n1570_0[0]),.dout(n1606),.clk(gclk));
	jnot g01397(.din(w_n1563_0[0]),.dout(n1607),.clk(gclk));
	jnot g01398(.din(w_n1555_0[0]),.dout(n1608),.clk(gclk));
	jnot g01399(.din(w_n1547_0[0]),.dout(n1609),.clk(gclk));
	jnot g01400(.din(w_n1539_0[0]),.dout(n1610),.clk(gclk));
	jnot g01401(.din(w_n1532_0[0]),.dout(n1611),.clk(gclk));
	jnot g01402(.din(w_n1521_0[0]),.dout(n1612),.clk(gclk));
	jnot g01403(.din(w_n1446_0[0]),.dout(n1613),.clk(gclk));
	jnot g01404(.din(w_n1443_0[0]),.dout(n1614),.clk(gclk));
	jor g01405(.dina(w_n1516_62[1]),.dinb(w_n1319_0[2]),.dout(n1615),.clk(gclk));
	jand g01406(.dina(n1615),.dinb(n1614),.dout(n1616),.clk(gclk));
	jand g01407(.dina(n1616),.dinb(w_n1332_63[1]),.dout(n1617),.clk(gclk));
	jor g01408(.dina(w_n1516_62[0]),.dinb(w_a100_0[0]),.dout(n1618),.clk(gclk));
	jand g01409(.dina(n1618),.dinb(w_a101_0[0]),.dout(n1619),.clk(gclk));
	jor g01410(.dina(w_n1523_0[0]),.dinb(n1619),.dout(n1620),.clk(gclk));
	jor g01411(.dina(n1620),.dinb(n1617),.dout(n1621),.clk(gclk));
	jand g01412(.dina(n1621),.dinb(n1613),.dout(n1622),.clk(gclk));
	jand g01413(.dina(n1622),.dinb(w_n1173_62[1]),.dout(n1623),.clk(gclk));
	jor g01414(.dina(w_n1528_0[1]),.dinb(n1623),.dout(n1624),.clk(gclk));
	jand g01415(.dina(n1624),.dinb(n1612),.dout(n1625),.clk(gclk));
	jand g01416(.dina(n1625),.dinb(w_n1008_64[1]),.dout(n1626),.clk(gclk));
	jnot g01417(.din(w_n1536_0[0]),.dout(n1627),.clk(gclk));
	jor g01418(.dina(w_n1627_0[1]),.dinb(n1626),.dout(n1628),.clk(gclk));
	jand g01419(.dina(n1628),.dinb(n1611),.dout(n1629),.clk(gclk));
	jand g01420(.dina(n1629),.dinb(w_n884_63[1]),.dout(n1630),.clk(gclk));
	jor g01421(.dina(w_n1543_0[0]),.dinb(n1630),.dout(n1631),.clk(gclk));
	jand g01422(.dina(n1631),.dinb(n1610),.dout(n1632),.clk(gclk));
	jand g01423(.dina(n1632),.dinb(w_n743_64[1]),.dout(n1633),.clk(gclk));
	jor g01424(.dina(w_n1551_0[0]),.dinb(n1633),.dout(n1634),.clk(gclk));
	jand g01425(.dina(n1634),.dinb(n1609),.dout(n1635),.clk(gclk));
	jand g01426(.dina(n1635),.dinb(w_n635_64[1]),.dout(n1636),.clk(gclk));
	jor g01427(.dina(w_n1559_0[0]),.dinb(n1636),.dout(n1637),.clk(gclk));
	jand g01428(.dina(n1637),.dinb(n1608),.dout(n1638),.clk(gclk));
	jand g01429(.dina(n1638),.dinb(w_n515_65[1]),.dout(n1639),.clk(gclk));
	jnot g01430(.din(w_n1567_0[0]),.dout(n1640),.clk(gclk));
	jor g01431(.dina(w_n1640_0[1]),.dinb(n1639),.dout(n1641),.clk(gclk));
	jand g01432(.dina(n1641),.dinb(n1607),.dout(n1642),.clk(gclk));
	jand g01433(.dina(n1642),.dinb(w_n443_65[1]),.dout(n1643),.clk(gclk));
	jor g01434(.dina(w_n1574_0[0]),.dinb(n1643),.dout(n1644),.clk(gclk));
	jand g01435(.dina(n1644),.dinb(n1606),.dout(n1645),.clk(gclk));
	jand g01436(.dina(n1645),.dinb(w_n352_65[2]),.dout(n1646),.clk(gclk));
	jor g01437(.dina(w_n1582_0[0]),.dinb(n1646),.dout(n1647),.clk(gclk));
	jand g01438(.dina(n1647),.dinb(n1605),.dout(n1648),.clk(gclk));
	jand g01439(.dina(n1648),.dinb(w_n294_66[0]),.dout(n1649),.clk(gclk));
	jor g01440(.dina(w_n1590_0[0]),.dinb(n1649),.dout(n1650),.clk(gclk));
	jand g01441(.dina(n1650),.dinb(n1604),.dout(n1651),.clk(gclk));
	jand g01442(.dina(n1651),.dinb(w_n239_66[1]),.dout(n1652),.clk(gclk));
	jnot g01443(.din(w_n1598_0[0]),.dout(n1653),.clk(gclk));
	jor g01444(.dina(w_n1653_0[1]),.dinb(n1652),.dout(n1654),.clk(gclk));
	jand g01445(.dina(n1654),.dinb(n1603),.dout(n1655),.clk(gclk));
	jand g01446(.dina(n1655),.dinb(w_n221_66[2]),.dout(n1656),.clk(gclk));
	jxor g01447(.dina(w_n1404_0[0]),.dinb(w_n239_66[0]),.dout(n1657),.clk(gclk));
	jand g01448(.dina(n1657),.dinb(w_asqrt50_39[0]),.dout(n1658),.clk(gclk));
	jxor g01449(.dina(n1658),.dinb(w_n1409_0[0]),.dout(n1659),.clk(gclk));
	jnot g01450(.din(w_n1659_0[2]),.dout(n1660),.clk(gclk));
	jor g01451(.dina(n1660),.dinb(n1656),.dout(n1661),.clk(gclk));
	jand g01452(.dina(n1661),.dinb(n1602),.dout(n1662),.clk(gclk));
	jxor g01453(.dina(w_n1412_0[0]),.dinb(w_n221_66[1]),.dout(n1663),.clk(gclk));
	jand g01454(.dina(n1663),.dinb(w_asqrt50_38[2]),.dout(n1664),.clk(gclk));
	jxor g01455(.dina(n1664),.dinb(w_n1418_0[0]),.dout(n1665),.clk(gclk));
	jor g01456(.dina(w_n1665_1[1]),.dinb(w_n1662_0[2]),.dout(n1666),.clk(gclk));
	jxor g01457(.dina(w_n1423_0[2]),.dinb(w_n1420_0[2]),.dout(n1667),.clk(gclk));
	jnot g01458(.din(w_n1667_0[1]),.dout(n1668),.clk(gclk));
	jand g01459(.dina(n1668),.dinb(w_asqrt50_38[1]),.dout(n1669),.clk(gclk));
	jor g01460(.dina(w_n1669_0[1]),.dinb(w_n1666_0[1]),.dout(n1670),.clk(gclk));
	jand g01461(.dina(n1670),.dinb(w_n218_27[1]),.dout(n1671),.clk(gclk));
	jand g01462(.dina(w_n1516_61[2]),.dinb(w_n1423_0[1]),.dout(n1672),.clk(gclk));
	jand g01463(.dina(w_n1665_1[0]),.dinb(w_n1662_0[1]),.dout(n1673),.clk(gclk));
	jor g01464(.dina(w_n1673_0[2]),.dinb(w_n1672_0[1]),.dout(n1674),.clk(gclk));
	jand g01465(.dina(w_n1514_0[0]),.dinb(w_n1420_0[1]),.dout(n1675),.clk(gclk));
	jnot g01466(.din(n1675),.dout(n1676),.clk(gclk));
	jand g01467(.dina(w_n1667_0[0]),.dinb(w_asqrt63_50[2]),.dout(n1677),.clk(gclk));
	jand g01468(.dina(w_n1677_0[1]),.dinb(n1676),.dout(n1678),.clk(gclk));
	jor g01469(.dina(w_n1678_0[1]),.dinb(n1674),.dout(n1679),.clk(gclk));
	jor g01470(.dina(n1679),.dinb(w_n1671_0[1]),.dout(asqrt_fa_50),.clk(gclk));
	jnot g01471(.din(w_a96_0[2]),.dout(n1681),.clk(gclk));
	jnot g01472(.din(w_a97_0[1]),.dout(n1682),.clk(gclk));
	jand g01473(.dina(w_n1682_0[1]),.dinb(w_n1681_1[2]),.dout(n1683),.clk(gclk));
	jand g01474(.dina(w_n1683_0[2]),.dinb(w_n1440_1[0]),.dout(n1684),.clk(gclk));
	jnot g01475(.din(w_n1684_0[1]),.dout(n1685),.clk(gclk));
	jor g01476(.dina(w_n1600_0[1]),.dinb(w_asqrt62_39[0]),.dout(n1686),.clk(gclk));
	jand g01477(.dina(w_n1659_0[1]),.dinb(n1686),.dout(n1687),.clk(gclk));
	jor g01478(.dina(n1687),.dinb(w_n1601_0[0]),.dout(n1688),.clk(gclk));
	jnot g01479(.din(w_n1665_0[2]),.dout(n1689),.clk(gclk));
	jand g01480(.dina(w_n1689_0[1]),.dinb(w_n1688_0[1]),.dout(n1690),.clk(gclk));
	jnot g01481(.din(w_n1669_0[0]),.dout(n1691),.clk(gclk));
	jand g01482(.dina(n1691),.dinb(w_n1690_0[1]),.dout(n1692),.clk(gclk));
	jor g01483(.dina(n1692),.dinb(w_asqrt63_50[1]),.dout(n1693),.clk(gclk));
	jnot g01484(.din(w_n1672_0[0]),.dout(n1694),.clk(gclk));
	jor g01485(.dina(w_n1689_0[0]),.dinb(w_n1688_0[0]),.dout(n1695),.clk(gclk));
	jand g01486(.dina(w_n1695_0[2]),.dinb(n1694),.dout(n1696),.clk(gclk));
	jnot g01487(.din(w_n1678_0[0]),.dout(n1697),.clk(gclk));
	jand g01488(.dina(n1697),.dinb(n1696),.dout(n1698),.clk(gclk));
	jand g01489(.dina(n1698),.dinb(n1693),.dout(n1699),.clk(gclk));
	jor g01490(.dina(w_n1699_67[1]),.dinb(w_n1440_0[2]),.dout(n1700),.clk(gclk));
	jand g01491(.dina(n1700),.dinb(n1685),.dout(n1701),.clk(gclk));
	jor g01492(.dina(w_n1701_0[2]),.dinb(w_n1516_61[1]),.dout(n1702),.clk(gclk));
	jand g01493(.dina(w_n1701_0[1]),.dinb(w_n1516_61[0]),.dout(n1703),.clk(gclk));
	jor g01494(.dina(w_n1699_67[0]),.dinb(w_a98_1[0]),.dout(n1704),.clk(gclk));
	jand g01495(.dina(n1704),.dinb(w_a99_0[0]),.dout(n1705),.clk(gclk));
	jand g01496(.dina(w_asqrt49_37[1]),.dinb(w_n1442_0[1]),.dout(n1706),.clk(gclk));
	jor g01497(.dina(n1706),.dinb(n1705),.dout(n1707),.clk(gclk));
	jor g01498(.dina(n1707),.dinb(n1703),.dout(n1708),.clk(gclk));
	jand g01499(.dina(n1708),.dinb(w_n1702_0[1]),.dout(n1709),.clk(gclk));
	jor g01500(.dina(w_n1709_0[2]),.dinb(w_n1332_63[0]),.dout(n1710),.clk(gclk));
	jand g01501(.dina(w_n1709_0[1]),.dinb(w_n1332_62[2]),.dout(n1711),.clk(gclk));
	jnot g01502(.din(w_n1442_0[0]),.dout(n1712),.clk(gclk));
	jor g01503(.dina(w_n1699_66[2]),.dinb(n1712),.dout(n1713),.clk(gclk));
	jor g01504(.dina(w_n1673_0[1]),.dinb(w_n1516_60[2]),.dout(n1714),.clk(gclk));
	jor g01505(.dina(n1714),.dinb(w_n1671_0[0]),.dout(n1715),.clk(gclk));
	jor g01506(.dina(n1715),.dinb(w_n1677_0[0]),.dout(n1716),.clk(gclk));
	jand g01507(.dina(n1716),.dinb(w_n1713_0[1]),.dout(n1717),.clk(gclk));
	jxor g01508(.dina(n1717),.dinb(w_n1319_0[1]),.dout(n1718),.clk(gclk));
	jor g01509(.dina(w_n1718_0[2]),.dinb(n1711),.dout(n1719),.clk(gclk));
	jand g01510(.dina(n1719),.dinb(w_n1710_0[1]),.dout(n1720),.clk(gclk));
	jor g01511(.dina(w_n1720_0[2]),.dinb(w_n1173_62[0]),.dout(n1721),.clk(gclk));
	jand g01512(.dina(w_n1720_0[1]),.dinb(w_n1173_61[2]),.dout(n1722),.clk(gclk));
	jxor g01513(.dina(w_n1445_0[0]),.dinb(w_n1332_62[1]),.dout(n1723),.clk(gclk));
	jor g01514(.dina(n1723),.dinb(w_n1699_66[1]),.dout(n1724),.clk(gclk));
	jxor g01515(.dina(n1724),.dinb(w_n1518_0[0]),.dout(n1725),.clk(gclk));
	jor g01516(.dina(w_n1725_0[2]),.dinb(n1722),.dout(n1726),.clk(gclk));
	jand g01517(.dina(n1726),.dinb(w_n1721_0[1]),.dout(n1727),.clk(gclk));
	jor g01518(.dina(w_n1727_0[2]),.dinb(w_n1008_64[0]),.dout(n1728),.clk(gclk));
	jand g01519(.dina(w_n1727_0[1]),.dinb(w_n1008_63[2]),.dout(n1729),.clk(gclk));
	jxor g01520(.dina(w_n1520_0[0]),.dinb(w_n1173_61[1]),.dout(n1730),.clk(gclk));
	jor g01521(.dina(n1730),.dinb(w_n1699_66[0]),.dout(n1731),.clk(gclk));
	jxor g01522(.dina(n1731),.dinb(w_n1528_0[0]),.dout(n1732),.clk(gclk));
	jnot g01523(.din(w_n1732_0[2]),.dout(n1733),.clk(gclk));
	jor g01524(.dina(n1733),.dinb(n1729),.dout(n1734),.clk(gclk));
	jand g01525(.dina(n1734),.dinb(w_n1728_0[1]),.dout(n1735),.clk(gclk));
	jor g01526(.dina(w_n1735_0[2]),.dinb(w_n884_63[0]),.dout(n1736),.clk(gclk));
	jand g01527(.dina(w_n1735_0[1]),.dinb(w_n884_62[2]),.dout(n1737),.clk(gclk));
	jxor g01528(.dina(w_n1531_0[0]),.dinb(w_n1008_63[1]),.dout(n1738),.clk(gclk));
	jor g01529(.dina(n1738),.dinb(w_n1699_65[2]),.dout(n1739),.clk(gclk));
	jxor g01530(.dina(n1739),.dinb(w_n1627_0[0]),.dout(n1740),.clk(gclk));
	jnot g01531(.din(w_n1740_0[2]),.dout(n1741),.clk(gclk));
	jor g01532(.dina(n1741),.dinb(n1737),.dout(n1742),.clk(gclk));
	jand g01533(.dina(n1742),.dinb(w_n1736_0[1]),.dout(n1743),.clk(gclk));
	jor g01534(.dina(w_n1743_0[2]),.dinb(w_n743_64[0]),.dout(n1744),.clk(gclk));
	jand g01535(.dina(w_n1743_0[1]),.dinb(w_n743_63[2]),.dout(n1745),.clk(gclk));
	jxor g01536(.dina(w_n1538_0[0]),.dinb(w_n884_62[1]),.dout(n1746),.clk(gclk));
	jor g01537(.dina(n1746),.dinb(w_n1699_65[1]),.dout(n1747),.clk(gclk));
	jxor g01538(.dina(n1747),.dinb(w_n1544_0[0]),.dout(n1748),.clk(gclk));
	jor g01539(.dina(w_n1748_0[2]),.dinb(n1745),.dout(n1749),.clk(gclk));
	jand g01540(.dina(n1749),.dinb(w_n1744_0[1]),.dout(n1750),.clk(gclk));
	jor g01541(.dina(w_n1750_0[2]),.dinb(w_n635_64[0]),.dout(n1751),.clk(gclk));
	jand g01542(.dina(w_n1750_0[1]),.dinb(w_n635_63[2]),.dout(n1752),.clk(gclk));
	jxor g01543(.dina(w_n1546_0[0]),.dinb(w_n743_63[1]),.dout(n1753),.clk(gclk));
	jor g01544(.dina(n1753),.dinb(w_n1699_65[0]),.dout(n1754),.clk(gclk));
	jxor g01545(.dina(n1754),.dinb(w_n1552_0[0]),.dout(n1755),.clk(gclk));
	jor g01546(.dina(w_n1755_0[2]),.dinb(n1752),.dout(n1756),.clk(gclk));
	jand g01547(.dina(n1756),.dinb(w_n1751_0[1]),.dout(n1757),.clk(gclk));
	jor g01548(.dina(w_n1757_0[2]),.dinb(w_n515_65[0]),.dout(n1758),.clk(gclk));
	jand g01549(.dina(w_n1757_0[1]),.dinb(w_n515_64[2]),.dout(n1759),.clk(gclk));
	jxor g01550(.dina(w_n1554_0[0]),.dinb(w_n635_63[1]),.dout(n1760),.clk(gclk));
	jor g01551(.dina(n1760),.dinb(w_n1699_64[2]),.dout(n1761),.clk(gclk));
	jxor g01552(.dina(n1761),.dinb(w_n1560_0[0]),.dout(n1762),.clk(gclk));
	jor g01553(.dina(w_n1762_0[2]),.dinb(n1759),.dout(n1763),.clk(gclk));
	jand g01554(.dina(n1763),.dinb(w_n1758_0[1]),.dout(n1764),.clk(gclk));
	jor g01555(.dina(w_n1764_0[2]),.dinb(w_n443_65[0]),.dout(n1765),.clk(gclk));
	jand g01556(.dina(w_n1764_0[1]),.dinb(w_n443_64[2]),.dout(n1766),.clk(gclk));
	jxor g01557(.dina(w_n1562_0[0]),.dinb(w_n515_64[1]),.dout(n1767),.clk(gclk));
	jor g01558(.dina(n1767),.dinb(w_n1699_64[1]),.dout(n1768),.clk(gclk));
	jxor g01559(.dina(n1768),.dinb(w_n1640_0[0]),.dout(n1769),.clk(gclk));
	jnot g01560(.din(w_n1769_0[2]),.dout(n1770),.clk(gclk));
	jor g01561(.dina(n1770),.dinb(n1766),.dout(n1771),.clk(gclk));
	jand g01562(.dina(n1771),.dinb(w_n1765_0[1]),.dout(n1772),.clk(gclk));
	jor g01563(.dina(w_n1772_0[2]),.dinb(w_n352_65[1]),.dout(n1773),.clk(gclk));
	jand g01564(.dina(w_n1772_0[1]),.dinb(w_n352_65[0]),.dout(n1774),.clk(gclk));
	jxor g01565(.dina(w_n1569_0[0]),.dinb(w_n443_64[1]),.dout(n1775),.clk(gclk));
	jor g01566(.dina(n1775),.dinb(w_n1699_64[0]),.dout(n1776),.clk(gclk));
	jxor g01567(.dina(n1776),.dinb(w_n1575_0[0]),.dout(n1777),.clk(gclk));
	jor g01568(.dina(w_n1777_0[2]),.dinb(n1774),.dout(n1778),.clk(gclk));
	jand g01569(.dina(n1778),.dinb(w_n1773_0[1]),.dout(n1779),.clk(gclk));
	jor g01570(.dina(w_n1779_0[2]),.dinb(w_n294_65[2]),.dout(n1780),.clk(gclk));
	jand g01571(.dina(w_n1779_0[1]),.dinb(w_n294_65[1]),.dout(n1781),.clk(gclk));
	jxor g01572(.dina(w_n1577_0[0]),.dinb(w_n352_64[2]),.dout(n1782),.clk(gclk));
	jor g01573(.dina(n1782),.dinb(w_n1699_63[2]),.dout(n1783),.clk(gclk));
	jxor g01574(.dina(n1783),.dinb(w_n1583_0[0]),.dout(n1784),.clk(gclk));
	jor g01575(.dina(w_n1784_0[2]),.dinb(n1781),.dout(n1785),.clk(gclk));
	jand g01576(.dina(n1785),.dinb(w_n1780_0[1]),.dout(n1786),.clk(gclk));
	jor g01577(.dina(w_n1786_0[2]),.dinb(w_n239_65[2]),.dout(n1787),.clk(gclk));
	jand g01578(.dina(w_n1786_0[1]),.dinb(w_n239_65[1]),.dout(n1788),.clk(gclk));
	jxor g01579(.dina(w_n1585_0[0]),.dinb(w_n294_65[0]),.dout(n1789),.clk(gclk));
	jor g01580(.dina(n1789),.dinb(w_n1699_63[1]),.dout(n1790),.clk(gclk));
	jxor g01581(.dina(n1790),.dinb(w_n1591_0[0]),.dout(n1791),.clk(gclk));
	jor g01582(.dina(w_n1791_0[2]),.dinb(n1788),.dout(n1792),.clk(gclk));
	jand g01583(.dina(n1792),.dinb(w_n1787_0[1]),.dout(n1793),.clk(gclk));
	jor g01584(.dina(w_n1793_0[2]),.dinb(w_n221_66[0]),.dout(n1794),.clk(gclk));
	jand g01585(.dina(w_n1793_0[1]),.dinb(w_n221_65[2]),.dout(n1795),.clk(gclk));
	jxor g01586(.dina(w_n1593_0[0]),.dinb(w_n239_65[0]),.dout(n1796),.clk(gclk));
	jor g01587(.dina(n1796),.dinb(w_n1699_63[0]),.dout(n1797),.clk(gclk));
	jxor g01588(.dina(n1797),.dinb(w_n1653_0[0]),.dout(n1798),.clk(gclk));
	jnot g01589(.din(w_n1798_0[2]),.dout(n1799),.clk(gclk));
	jor g01590(.dina(n1799),.dinb(n1795),.dout(n1800),.clk(gclk));
	jand g01591(.dina(n1800),.dinb(w_n1794_0[1]),.dout(n1801),.clk(gclk));
	jxor g01592(.dina(w_n1600_0[0]),.dinb(w_n221_65[1]),.dout(n1802),.clk(gclk));
	jor g01593(.dina(n1802),.dinb(w_n1699_62[2]),.dout(n1803),.clk(gclk));
	jxor g01594(.dina(n1803),.dinb(w_n1659_0[0]),.dout(n1804),.clk(gclk));
	jand g01595(.dina(w_n1804_1[1]),.dinb(w_n1801_0[2]),.dout(n1805),.clk(gclk));
	jand g01596(.dina(w_n1699_62[1]),.dinb(w_n1662_0[0]),.dout(n1806),.clk(gclk));
	jand g01597(.dina(w_n1666_0[0]),.dinb(w_asqrt63_50[0]),.dout(n1807),.clk(gclk));
	jand g01598(.dina(n1807),.dinb(w_n1695_0[1]),.dout(n1808),.clk(gclk));
	jnot g01599(.din(n1808),.dout(n1809),.clk(gclk));
	jor g01600(.dina(w_n1809_0[1]),.dinb(n1806),.dout(n1810),.clk(gclk));
	jnot g01601(.din(w_n1810_0[1]),.dout(n1811),.clk(gclk));
	jor g01602(.dina(w_n1804_1[0]),.dinb(w_n1801_0[1]),.dout(n1812),.clk(gclk));
	jand g01603(.dina(w_asqrt49_37[0]),.dinb(w_n1690_0[0]),.dout(n1813),.clk(gclk));
	jor g01604(.dina(w_n1813_0[1]),.dinb(w_n1812_0[1]),.dout(n1814),.clk(gclk));
	jor g01605(.dina(n1814),.dinb(w_n1673_0[0]),.dout(n1815),.clk(gclk));
	jand g01606(.dina(n1815),.dinb(w_n218_27[0]),.dout(n1816),.clk(gclk));
	jand g01607(.dina(w_n1699_62[0]),.dinb(w_n1665_0[1]),.dout(n1817),.clk(gclk));
	jor g01608(.dina(w_n1817_0[1]),.dinb(n1816),.dout(n1818),.clk(gclk));
	jor g01609(.dina(n1818),.dinb(n1811),.dout(n1819),.clk(gclk));
	jor g01610(.dina(w_n1819_0[1]),.dinb(w_n1805_0[2]),.dout(asqrt_fa_49),.clk(gclk));
	jnot g01611(.din(w_n1794_0[0]),.dout(n1821),.clk(gclk));
	jnot g01612(.din(w_n1787_0[0]),.dout(n1822),.clk(gclk));
	jnot g01613(.din(w_n1780_0[0]),.dout(n1823),.clk(gclk));
	jnot g01614(.din(w_n1773_0[0]),.dout(n1824),.clk(gclk));
	jnot g01615(.din(w_n1765_0[0]),.dout(n1825),.clk(gclk));
	jnot g01616(.din(w_n1758_0[0]),.dout(n1826),.clk(gclk));
	jnot g01617(.din(w_n1751_0[0]),.dout(n1827),.clk(gclk));
	jnot g01618(.din(w_n1744_0[0]),.dout(n1828),.clk(gclk));
	jnot g01619(.din(w_n1736_0[0]),.dout(n1829),.clk(gclk));
	jnot g01620(.din(w_n1728_0[0]),.dout(n1830),.clk(gclk));
	jnot g01621(.din(w_n1721_0[0]),.dout(n1831),.clk(gclk));
	jnot g01622(.din(w_n1710_0[0]),.dout(n1832),.clk(gclk));
	jnot g01623(.din(w_n1702_0[0]),.dout(n1833),.clk(gclk));
	jand g01624(.dina(w_asqrt49_36[2]),.dinb(w_a98_0[2]),.dout(n1834),.clk(gclk));
	jor g01625(.dina(n1834),.dinb(w_n1684_0[0]),.dout(n1835),.clk(gclk));
	jor g01626(.dina(n1835),.dinb(w_asqrt50_38[0]),.dout(n1836),.clk(gclk));
	jand g01627(.dina(w_asqrt49_36[1]),.dinb(w_n1440_0[1]),.dout(n1837),.clk(gclk));
	jor g01628(.dina(n1837),.dinb(w_n1441_0[0]),.dout(n1838),.clk(gclk));
	jand g01629(.dina(w_n1713_0[0]),.dinb(n1838),.dout(n1839),.clk(gclk));
	jand g01630(.dina(w_n1839_0[1]),.dinb(n1836),.dout(n1840),.clk(gclk));
	jor g01631(.dina(n1840),.dinb(n1833),.dout(n1841),.clk(gclk));
	jor g01632(.dina(n1841),.dinb(w_asqrt51_36[1]),.dout(n1842),.clk(gclk));
	jnot g01633(.din(w_n1718_0[1]),.dout(n1843),.clk(gclk));
	jand g01634(.dina(n1843),.dinb(n1842),.dout(n1844),.clk(gclk));
	jor g01635(.dina(n1844),.dinb(n1832),.dout(n1845),.clk(gclk));
	jor g01636(.dina(n1845),.dinb(w_asqrt52_38[0]),.dout(n1846),.clk(gclk));
	jnot g01637(.din(w_n1725_0[1]),.dout(n1847),.clk(gclk));
	jand g01638(.dina(n1847),.dinb(n1846),.dout(n1848),.clk(gclk));
	jor g01639(.dina(n1848),.dinb(n1831),.dout(n1849),.clk(gclk));
	jor g01640(.dina(n1849),.dinb(w_asqrt53_37[0]),.dout(n1850),.clk(gclk));
	jand g01641(.dina(w_n1732_0[1]),.dinb(n1850),.dout(n1851),.clk(gclk));
	jor g01642(.dina(n1851),.dinb(n1830),.dout(n1852),.clk(gclk));
	jor g01643(.dina(n1852),.dinb(w_asqrt54_38[0]),.dout(n1853),.clk(gclk));
	jand g01644(.dina(w_n1740_0[1]),.dinb(n1853),.dout(n1854),.clk(gclk));
	jor g01645(.dina(n1854),.dinb(n1829),.dout(n1855),.clk(gclk));
	jor g01646(.dina(n1855),.dinb(w_asqrt55_37[1]),.dout(n1856),.clk(gclk));
	jnot g01647(.din(w_n1748_0[1]),.dout(n1857),.clk(gclk));
	jand g01648(.dina(n1857),.dinb(n1856),.dout(n1858),.clk(gclk));
	jor g01649(.dina(n1858),.dinb(n1828),.dout(n1859),.clk(gclk));
	jor g01650(.dina(n1859),.dinb(w_asqrt56_38[1]),.dout(n1860),.clk(gclk));
	jnot g01651(.din(w_n1755_0[1]),.dout(n1861),.clk(gclk));
	jand g01652(.dina(n1861),.dinb(n1860),.dout(n1862),.clk(gclk));
	jor g01653(.dina(n1862),.dinb(n1827),.dout(n1863),.clk(gclk));
	jor g01654(.dina(n1863),.dinb(w_asqrt57_38[0]),.dout(n1864),.clk(gclk));
	jnot g01655(.din(w_n1762_0[1]),.dout(n1865),.clk(gclk));
	jand g01656(.dina(n1865),.dinb(n1864),.dout(n1866),.clk(gclk));
	jor g01657(.dina(n1866),.dinb(n1826),.dout(n1867),.clk(gclk));
	jor g01658(.dina(n1867),.dinb(w_asqrt58_38[2]),.dout(n1868),.clk(gclk));
	jand g01659(.dina(w_n1769_0[1]),.dinb(n1868),.dout(n1869),.clk(gclk));
	jor g01660(.dina(n1869),.dinb(n1825),.dout(n1870),.clk(gclk));
	jor g01661(.dina(n1870),.dinb(w_asqrt59_38[1]),.dout(n1871),.clk(gclk));
	jnot g01662(.din(w_n1777_0[1]),.dout(n1872),.clk(gclk));
	jand g01663(.dina(n1872),.dinb(n1871),.dout(n1873),.clk(gclk));
	jor g01664(.dina(n1873),.dinb(n1824),.dout(n1874),.clk(gclk));
	jor g01665(.dina(n1874),.dinb(w_asqrt60_38[2]),.dout(n1875),.clk(gclk));
	jnot g01666(.din(w_n1784_0[1]),.dout(n1876),.clk(gclk));
	jand g01667(.dina(n1876),.dinb(n1875),.dout(n1877),.clk(gclk));
	jor g01668(.dina(n1877),.dinb(n1823),.dout(n1878),.clk(gclk));
	jor g01669(.dina(n1878),.dinb(w_asqrt61_38[2]),.dout(n1879),.clk(gclk));
	jnot g01670(.din(w_n1791_0[1]),.dout(n1880),.clk(gclk));
	jand g01671(.dina(n1880),.dinb(n1879),.dout(n1881),.clk(gclk));
	jor g01672(.dina(n1881),.dinb(n1822),.dout(n1882),.clk(gclk));
	jor g01673(.dina(n1882),.dinb(w_asqrt62_38[2]),.dout(n1883),.clk(gclk));
	jand g01674(.dina(w_n1798_0[1]),.dinb(n1883),.dout(n1884),.clk(gclk));
	jor g01675(.dina(n1884),.dinb(n1821),.dout(n1885),.clk(gclk));
	jnot g01676(.din(w_n1804_0[2]),.dout(n1886),.clk(gclk));
	jand g01677(.dina(n1886),.dinb(n1885),.dout(n1887),.clk(gclk));
	jand g01678(.dina(w_n1819_0[0]),.dinb(w_n1887_0[1]),.dout(n1888),.clk(gclk));
	jxor g01679(.dina(w_n1793_0[0]),.dinb(w_n221_65[0]),.dout(n1889),.clk(gclk));
	jand g01680(.dina(n1889),.dinb(w_asqrt48_42),.dout(n1890),.clk(gclk));
	jxor g01681(.dina(n1890),.dinb(w_n1798_0[0]),.dout(n1891),.clk(gclk));
	jnot g01682(.din(w_n1891_0[2]),.dout(n1892),.clk(gclk));
	jand g01683(.dina(w_asqrt48_41[2]),.dinb(w_a96_0[1]),.dout(n1893),.clk(gclk));
	jnot g01684(.din(w_a94_1[1]),.dout(n1894),.clk(gclk));
	jnot g01685(.din(w_a95_0[1]),.dout(n1895),.clk(gclk));
	jand g01686(.dina(w_n1895_0[1]),.dinb(w_n1894_1[1]),.dout(n1896),.clk(gclk));
	jand g01687(.dina(w_n1896_0[2]),.dinb(w_n1681_1[1]),.dout(n1897),.clk(gclk));
	jor g01688(.dina(w_n1897_0[1]),.dinb(n1893),.dout(n1898),.clk(gclk));
	jand g01689(.dina(w_n1898_0[2]),.dinb(w_asqrt49_36[0]),.dout(n1899),.clk(gclk));
	jor g01690(.dina(w_n1898_0[1]),.dinb(w_asqrt49_35[2]),.dout(n1900),.clk(gclk));
	jand g01691(.dina(w_asqrt48_41[1]),.dinb(w_n1681_1[0]),.dout(n1901),.clk(gclk));
	jor g01692(.dina(n1901),.dinb(w_n1682_0[0]),.dout(n1902),.clk(gclk));
	jnot g01693(.din(w_n1683_0[1]),.dout(n1903),.clk(gclk));
	jnot g01694(.din(w_n1805_0[1]),.dout(n1904),.clk(gclk));
	jnot g01695(.din(w_n1813_0[0]),.dout(n1905),.clk(gclk));
	jand g01696(.dina(n1905),.dinb(w_n1887_0[0]),.dout(n1906),.clk(gclk));
	jand g01697(.dina(n1906),.dinb(w_n1695_0[0]),.dout(n1907),.clk(gclk));
	jor g01698(.dina(n1907),.dinb(w_asqrt63_49[2]),.dout(n1908),.clk(gclk));
	jnot g01699(.din(w_n1817_0[0]),.dout(n1909),.clk(gclk));
	jand g01700(.dina(n1909),.dinb(w_n1908_0[1]),.dout(n1910),.clk(gclk));
	jand g01701(.dina(n1910),.dinb(w_n1810_0[0]),.dout(n1911),.clk(gclk));
	jand g01702(.dina(w_n1911_0[1]),.dinb(w_n1904_1[1]),.dout(n1912),.clk(gclk));
	jor g01703(.dina(w_n1912_60[1]),.dinb(n1903),.dout(n1913),.clk(gclk));
	jand g01704(.dina(n1913),.dinb(n1902),.dout(n1914),.clk(gclk));
	jand g01705(.dina(n1914),.dinb(n1900),.dout(n1915),.clk(gclk));
	jor g01706(.dina(n1915),.dinb(w_n1899_0[1]),.dout(n1916),.clk(gclk));
	jand g01707(.dina(w_n1916_0[2]),.dinb(w_asqrt50_37[2]),.dout(n1917),.clk(gclk));
	jor g01708(.dina(w_n1916_0[1]),.dinb(w_asqrt50_37[1]),.dout(n1918),.clk(gclk));
	jand g01709(.dina(w_asqrt48_41[0]),.dinb(w_n1683_0[0]),.dout(n1919),.clk(gclk));
	jand g01710(.dina(w_n1904_1[0]),.dinb(w_asqrt49_35[1]),.dout(n1920),.clk(gclk));
	jand g01711(.dina(n1920),.dinb(w_n1809_0[0]),.dout(n1921),.clk(gclk));
	jand g01712(.dina(n1921),.dinb(w_n1908_0[0]),.dout(n1922),.clk(gclk));
	jor g01713(.dina(n1922),.dinb(w_n1919_0[1]),.dout(n1923),.clk(gclk));
	jxor g01714(.dina(n1923),.dinb(w_a98_0[1]),.dout(n1924),.clk(gclk));
	jnot g01715(.din(w_n1924_0[1]),.dout(n1925),.clk(gclk));
	jand g01716(.dina(w_n1925_0[1]),.dinb(n1918),.dout(n1926),.clk(gclk));
	jor g01717(.dina(n1926),.dinb(w_n1917_0[1]),.dout(n1927),.clk(gclk));
	jand g01718(.dina(w_n1927_0[2]),.dinb(w_asqrt51_36[0]),.dout(n1928),.clk(gclk));
	jor g01719(.dina(w_n1927_0[1]),.dinb(w_asqrt51_35[2]),.dout(n1929),.clk(gclk));
	jxor g01720(.dina(w_n1701_0[0]),.dinb(w_n1516_60[1]),.dout(n1930),.clk(gclk));
	jand g01721(.dina(n1930),.dinb(w_asqrt48_40[2]),.dout(n1931),.clk(gclk));
	jxor g01722(.dina(n1931),.dinb(w_n1839_0[0]),.dout(n1932),.clk(gclk));
	jand g01723(.dina(w_n1932_0[1]),.dinb(n1929),.dout(n1933),.clk(gclk));
	jor g01724(.dina(n1933),.dinb(w_n1928_0[1]),.dout(n1934),.clk(gclk));
	jand g01725(.dina(w_n1934_0[2]),.dinb(w_asqrt52_37[2]),.dout(n1935),.clk(gclk));
	jor g01726(.dina(w_n1934_0[1]),.dinb(w_asqrt52_37[1]),.dout(n1936),.clk(gclk));
	jxor g01727(.dina(w_n1709_0[0]),.dinb(w_n1332_62[0]),.dout(n1937),.clk(gclk));
	jand g01728(.dina(n1937),.dinb(w_asqrt48_40[1]),.dout(n1938),.clk(gclk));
	jxor g01729(.dina(n1938),.dinb(w_n1718_0[0]),.dout(n1939),.clk(gclk));
	jnot g01730(.din(w_n1939_0[1]),.dout(n1940),.clk(gclk));
	jand g01731(.dina(w_n1940_0[1]),.dinb(n1936),.dout(n1941),.clk(gclk));
	jor g01732(.dina(n1941),.dinb(w_n1935_0[1]),.dout(n1942),.clk(gclk));
	jand g01733(.dina(w_n1942_0[2]),.dinb(w_asqrt53_36[2]),.dout(n1943),.clk(gclk));
	jor g01734(.dina(w_n1942_0[1]),.dinb(w_asqrt53_36[1]),.dout(n1944),.clk(gclk));
	jxor g01735(.dina(w_n1720_0[0]),.dinb(w_n1173_61[0]),.dout(n1945),.clk(gclk));
	jand g01736(.dina(n1945),.dinb(w_asqrt48_40[0]),.dout(n1946),.clk(gclk));
	jxor g01737(.dina(n1946),.dinb(w_n1725_0[0]),.dout(n1947),.clk(gclk));
	jnot g01738(.din(w_n1947_0[1]),.dout(n1948),.clk(gclk));
	jand g01739(.dina(w_n1948_0[1]),.dinb(n1944),.dout(n1949),.clk(gclk));
	jor g01740(.dina(n1949),.dinb(w_n1943_0[1]),.dout(n1950),.clk(gclk));
	jand g01741(.dina(w_n1950_0[2]),.dinb(w_asqrt54_37[2]),.dout(n1951),.clk(gclk));
	jor g01742(.dina(w_n1950_0[1]),.dinb(w_asqrt54_37[1]),.dout(n1952),.clk(gclk));
	jxor g01743(.dina(w_n1727_0[0]),.dinb(w_n1008_63[0]),.dout(n1953),.clk(gclk));
	jand g01744(.dina(n1953),.dinb(w_asqrt48_39[2]),.dout(n1954),.clk(gclk));
	jxor g01745(.dina(n1954),.dinb(w_n1732_0[0]),.dout(n1955),.clk(gclk));
	jand g01746(.dina(w_n1955_0[1]),.dinb(n1952),.dout(n1956),.clk(gclk));
	jor g01747(.dina(n1956),.dinb(w_n1951_0[1]),.dout(n1957),.clk(gclk));
	jand g01748(.dina(w_n1957_0[2]),.dinb(w_asqrt55_37[0]),.dout(n1958),.clk(gclk));
	jor g01749(.dina(w_n1957_0[1]),.dinb(w_asqrt55_36[2]),.dout(n1959),.clk(gclk));
	jxor g01750(.dina(w_n1735_0[0]),.dinb(w_n884_62[0]),.dout(n1960),.clk(gclk));
	jand g01751(.dina(n1960),.dinb(w_asqrt48_39[1]),.dout(n1961),.clk(gclk));
	jxor g01752(.dina(n1961),.dinb(w_n1740_0[0]),.dout(n1962),.clk(gclk));
	jand g01753(.dina(w_n1962_0[1]),.dinb(n1959),.dout(n1963),.clk(gclk));
	jor g01754(.dina(n1963),.dinb(w_n1958_0[1]),.dout(n1964),.clk(gclk));
	jand g01755(.dina(w_n1964_0[2]),.dinb(w_asqrt56_38[0]),.dout(n1965),.clk(gclk));
	jor g01756(.dina(w_n1964_0[1]),.dinb(w_asqrt56_37[2]),.dout(n1966),.clk(gclk));
	jxor g01757(.dina(w_n1743_0[0]),.dinb(w_n743_63[0]),.dout(n1967),.clk(gclk));
	jand g01758(.dina(n1967),.dinb(w_asqrt48_39[0]),.dout(n1968),.clk(gclk));
	jxor g01759(.dina(n1968),.dinb(w_n1748_0[0]),.dout(n1969),.clk(gclk));
	jnot g01760(.din(w_n1969_0[1]),.dout(n1970),.clk(gclk));
	jand g01761(.dina(w_n1970_0[1]),.dinb(n1966),.dout(n1971),.clk(gclk));
	jor g01762(.dina(n1971),.dinb(w_n1965_0[1]),.dout(n1972),.clk(gclk));
	jand g01763(.dina(w_n1972_0[2]),.dinb(w_asqrt57_37[2]),.dout(n1973),.clk(gclk));
	jor g01764(.dina(w_n1972_0[1]),.dinb(w_asqrt57_37[1]),.dout(n1974),.clk(gclk));
	jxor g01765(.dina(w_n1750_0[0]),.dinb(w_n635_63[0]),.dout(n1975),.clk(gclk));
	jand g01766(.dina(n1975),.dinb(w_asqrt48_38[2]),.dout(n1976),.clk(gclk));
	jxor g01767(.dina(n1976),.dinb(w_n1755_0[0]),.dout(n1977),.clk(gclk));
	jnot g01768(.din(w_n1977_0[1]),.dout(n1978),.clk(gclk));
	jand g01769(.dina(w_n1978_0[1]),.dinb(n1974),.dout(n1979),.clk(gclk));
	jor g01770(.dina(n1979),.dinb(w_n1973_0[1]),.dout(n1980),.clk(gclk));
	jand g01771(.dina(w_n1980_0[2]),.dinb(w_asqrt58_38[1]),.dout(n1981),.clk(gclk));
	jor g01772(.dina(w_n1980_0[1]),.dinb(w_asqrt58_38[0]),.dout(n1982),.clk(gclk));
	jxor g01773(.dina(w_n1757_0[0]),.dinb(w_n515_64[0]),.dout(n1983),.clk(gclk));
	jand g01774(.dina(n1983),.dinb(w_asqrt48_38[1]),.dout(n1984),.clk(gclk));
	jxor g01775(.dina(n1984),.dinb(w_n1762_0[0]),.dout(n1985),.clk(gclk));
	jnot g01776(.din(w_n1985_0[2]),.dout(n1986),.clk(gclk));
	jand g01777(.dina(n1986),.dinb(n1982),.dout(n1987),.clk(gclk));
	jor g01778(.dina(n1987),.dinb(w_n1981_0[1]),.dout(n1988),.clk(gclk));
	jand g01779(.dina(w_n1988_0[2]),.dinb(w_asqrt59_38[0]),.dout(n1989),.clk(gclk));
	jor g01780(.dina(w_n1988_0[1]),.dinb(w_asqrt59_37[2]),.dout(n1990),.clk(gclk));
	jxor g01781(.dina(w_n1764_0[0]),.dinb(w_n443_64[0]),.dout(n1991),.clk(gclk));
	jand g01782(.dina(n1991),.dinb(w_asqrt48_38[0]),.dout(n1992),.clk(gclk));
	jxor g01783(.dina(n1992),.dinb(w_n1769_0[0]),.dout(n1993),.clk(gclk));
	jand g01784(.dina(w_n1993_0[1]),.dinb(n1990),.dout(n1994),.clk(gclk));
	jor g01785(.dina(n1994),.dinb(w_n1989_0[1]),.dout(n1995),.clk(gclk));
	jand g01786(.dina(w_n1995_0[2]),.dinb(w_asqrt60_38[1]),.dout(n1996),.clk(gclk));
	jor g01787(.dina(w_n1995_0[1]),.dinb(w_asqrt60_38[0]),.dout(n1997),.clk(gclk));
	jxor g01788(.dina(w_n1772_0[0]),.dinb(w_n352_64[1]),.dout(n1998),.clk(gclk));
	jand g01789(.dina(n1998),.dinb(w_asqrt48_37[2]),.dout(n1999),.clk(gclk));
	jxor g01790(.dina(n1999),.dinb(w_n1777_0[0]),.dout(n2000),.clk(gclk));
	jnot g01791(.din(w_n2000_0[1]),.dout(n2001),.clk(gclk));
	jand g01792(.dina(w_n2001_0[1]),.dinb(n1997),.dout(n2002),.clk(gclk));
	jor g01793(.dina(n2002),.dinb(w_n1996_0[1]),.dout(n2003),.clk(gclk));
	jand g01794(.dina(w_n2003_0[2]),.dinb(w_asqrt61_38[1]),.dout(n2004),.clk(gclk));
	jor g01795(.dina(w_n2003_0[1]),.dinb(w_asqrt61_38[0]),.dout(n2005),.clk(gclk));
	jxor g01796(.dina(w_n1779_0[0]),.dinb(w_n294_64[2]),.dout(n2006),.clk(gclk));
	jand g01797(.dina(n2006),.dinb(w_asqrt48_37[1]),.dout(n2007),.clk(gclk));
	jxor g01798(.dina(n2007),.dinb(w_n1784_0[0]),.dout(n2008),.clk(gclk));
	jnot g01799(.din(w_n2008_0[1]),.dout(n2009),.clk(gclk));
	jand g01800(.dina(w_n2009_0[1]),.dinb(n2005),.dout(n2010),.clk(gclk));
	jor g01801(.dina(n2010),.dinb(w_n2004_0[1]),.dout(n2011),.clk(gclk));
	jand g01802(.dina(w_n2011_0[2]),.dinb(w_asqrt62_38[1]),.dout(n2012),.clk(gclk));
	jnot g01803(.din(w_n2012_0[1]),.dout(n2013),.clk(gclk));
	jnot g01804(.din(w_n2004_0[0]),.dout(n2014),.clk(gclk));
	jnot g01805(.din(w_n1996_0[0]),.dout(n2015),.clk(gclk));
	jnot g01806(.din(w_n1989_0[0]),.dout(n2016),.clk(gclk));
	jnot g01807(.din(w_n1981_0[0]),.dout(n2017),.clk(gclk));
	jnot g01808(.din(w_n1973_0[0]),.dout(n2018),.clk(gclk));
	jnot g01809(.din(w_n1965_0[0]),.dout(n2019),.clk(gclk));
	jnot g01810(.din(w_n1958_0[0]),.dout(n2020),.clk(gclk));
	jnot g01811(.din(w_n1951_0[0]),.dout(n2021),.clk(gclk));
	jnot g01812(.din(w_n1943_0[0]),.dout(n2022),.clk(gclk));
	jnot g01813(.din(w_n1935_0[0]),.dout(n2023),.clk(gclk));
	jnot g01814(.din(w_n1928_0[0]),.dout(n2024),.clk(gclk));
	jnot g01815(.din(w_n1917_0[0]),.dout(n2025),.clk(gclk));
	jnot g01816(.din(w_n1899_0[0]),.dout(n2026),.clk(gclk));
	jor g01817(.dina(w_n1912_60[0]),.dinb(w_n1681_0[2]),.dout(n2027),.clk(gclk));
	jnot g01818(.din(w_n1897_0[0]),.dout(n2028),.clk(gclk));
	jand g01819(.dina(n2028),.dinb(n2027),.dout(n2029),.clk(gclk));
	jand g01820(.dina(n2029),.dinb(w_n1699_61[2]),.dout(n2030),.clk(gclk));
	jor g01821(.dina(w_n1912_59[2]),.dinb(w_a96_0[0]),.dout(n2031),.clk(gclk));
	jand g01822(.dina(n2031),.dinb(w_a97_0[0]),.dout(n2032),.clk(gclk));
	jor g01823(.dina(w_n1919_0[0]),.dinb(n2032),.dout(n2033),.clk(gclk));
	jor g01824(.dina(w_n2033_0[1]),.dinb(n2030),.dout(n2034),.clk(gclk));
	jand g01825(.dina(n2034),.dinb(n2026),.dout(n2035),.clk(gclk));
	jand g01826(.dina(n2035),.dinb(w_n1516_60[0]),.dout(n2036),.clk(gclk));
	jor g01827(.dina(w_n1924_0[0]),.dinb(n2036),.dout(n2037),.clk(gclk));
	jand g01828(.dina(n2037),.dinb(n2025),.dout(n2038),.clk(gclk));
	jand g01829(.dina(n2038),.dinb(w_n1332_61[2]),.dout(n2039),.clk(gclk));
	jnot g01830(.din(w_n1932_0[0]),.dout(n2040),.clk(gclk));
	jor g01831(.dina(w_n2040_0[1]),.dinb(n2039),.dout(n2041),.clk(gclk));
	jand g01832(.dina(n2041),.dinb(n2024),.dout(n2042),.clk(gclk));
	jand g01833(.dina(n2042),.dinb(w_n1173_60[2]),.dout(n2043),.clk(gclk));
	jor g01834(.dina(w_n1939_0[0]),.dinb(n2043),.dout(n2044),.clk(gclk));
	jand g01835(.dina(n2044),.dinb(n2023),.dout(n2045),.clk(gclk));
	jand g01836(.dina(n2045),.dinb(w_n1008_62[2]),.dout(n2046),.clk(gclk));
	jor g01837(.dina(w_n1947_0[0]),.dinb(n2046),.dout(n2047),.clk(gclk));
	jand g01838(.dina(n2047),.dinb(n2022),.dout(n2048),.clk(gclk));
	jand g01839(.dina(n2048),.dinb(w_n884_61[2]),.dout(n2049),.clk(gclk));
	jnot g01840(.din(w_n1955_0[0]),.dout(n2050),.clk(gclk));
	jor g01841(.dina(w_n2050_0[1]),.dinb(n2049),.dout(n2051),.clk(gclk));
	jand g01842(.dina(n2051),.dinb(n2021),.dout(n2052),.clk(gclk));
	jand g01843(.dina(n2052),.dinb(w_n743_62[2]),.dout(n2053),.clk(gclk));
	jnot g01844(.din(w_n1962_0[0]),.dout(n2054),.clk(gclk));
	jor g01845(.dina(w_n2054_0[1]),.dinb(n2053),.dout(n2055),.clk(gclk));
	jand g01846(.dina(n2055),.dinb(n2020),.dout(n2056),.clk(gclk));
	jand g01847(.dina(n2056),.dinb(w_n635_62[2]),.dout(n2057),.clk(gclk));
	jor g01848(.dina(w_n1969_0[0]),.dinb(n2057),.dout(n2058),.clk(gclk));
	jand g01849(.dina(n2058),.dinb(n2019),.dout(n2059),.clk(gclk));
	jand g01850(.dina(n2059),.dinb(w_n515_63[2]),.dout(n2060),.clk(gclk));
	jor g01851(.dina(w_n1977_0[0]),.dinb(n2060),.dout(n2061),.clk(gclk));
	jand g01852(.dina(n2061),.dinb(n2018),.dout(n2062),.clk(gclk));
	jand g01853(.dina(n2062),.dinb(w_n443_63[2]),.dout(n2063),.clk(gclk));
	jor g01854(.dina(w_n1985_0[1]),.dinb(n2063),.dout(n2064),.clk(gclk));
	jand g01855(.dina(n2064),.dinb(n2017),.dout(n2065),.clk(gclk));
	jand g01856(.dina(n2065),.dinb(w_n352_64[0]),.dout(n2066),.clk(gclk));
	jnot g01857(.din(w_n1993_0[0]),.dout(n2067),.clk(gclk));
	jor g01858(.dina(w_n2067_0[1]),.dinb(n2066),.dout(n2068),.clk(gclk));
	jand g01859(.dina(n2068),.dinb(n2016),.dout(n2069),.clk(gclk));
	jand g01860(.dina(n2069),.dinb(w_n294_64[1]),.dout(n2070),.clk(gclk));
	jor g01861(.dina(w_n2000_0[0]),.dinb(n2070),.dout(n2071),.clk(gclk));
	jand g01862(.dina(n2071),.dinb(n2015),.dout(n2072),.clk(gclk));
	jand g01863(.dina(n2072),.dinb(w_n239_64[2]),.dout(n2073),.clk(gclk));
	jor g01864(.dina(w_n2008_0[0]),.dinb(n2073),.dout(n2074),.clk(gclk));
	jand g01865(.dina(n2074),.dinb(n2014),.dout(n2075),.clk(gclk));
	jand g01866(.dina(n2075),.dinb(w_n221_64[2]),.dout(n2076),.clk(gclk));
	jxor g01867(.dina(w_n1786_0[0]),.dinb(w_n239_64[1]),.dout(n2077),.clk(gclk));
	jand g01868(.dina(n2077),.dinb(w_asqrt48_37[0]),.dout(n2078),.clk(gclk));
	jxor g01869(.dina(n2078),.dinb(w_n1791_0[0]),.dout(n2079),.clk(gclk));
	jor g01870(.dina(w_n2079_0[1]),.dinb(n2076),.dout(n2080),.clk(gclk));
	jand g01871(.dina(n2080),.dinb(n2013),.dout(n2081),.clk(gclk));
	jor g01872(.dina(w_n2081_0[1]),.dinb(n1892),.dout(n2082),.clk(gclk));
	jor g01873(.dina(w_n2082_0[1]),.dinb(w_n1805_0[0]),.dout(n2083),.clk(gclk));
	jor g01874(.dina(n2083),.dinb(w_n1888_0[1]),.dout(n2084),.clk(gclk));
	jand g01875(.dina(n2084),.dinb(w_n218_26[2]),.dout(n2085),.clk(gclk));
	jand g01876(.dina(w_n1912_59[1]),.dinb(w_n1804_0[1]),.dout(n2086),.clk(gclk));
	jnot g01877(.din(n2086),.dout(n2087),.clk(gclk));
	jor g01878(.dina(w_n2011_0[1]),.dinb(w_asqrt62_38[0]),.dout(n2088),.clk(gclk));
	jnot g01879(.din(w_n2079_0[0]),.dout(n2089),.clk(gclk));
	jand g01880(.dina(w_n2089_0[1]),.dinb(n2088),.dout(n2090),.clk(gclk));
	jor g01881(.dina(n2090),.dinb(w_n2012_0[0]),.dout(n2091),.clk(gclk));
	jor g01882(.dina(w_n2091_0[1]),.dinb(w_n1891_0[1]),.dout(n2092),.clk(gclk));
	jand g01883(.dina(w_n2092_0[2]),.dinb(n2087),.dout(n2093),.clk(gclk));
	jand g01884(.dina(w_n1911_0[0]),.dinb(w_n1801_0[0]),.dout(n2094),.clk(gclk));
	jnot g01885(.din(n2094),.dout(n2095),.clk(gclk));
	jand g01886(.dina(w_n1812_0[0]),.dinb(w_asqrt63_49[1]),.dout(n2096),.clk(gclk));
	jand g01887(.dina(n2096),.dinb(w_n1904_0[2]),.dout(n2097),.clk(gclk));
	jand g01888(.dina(w_n2097_0[1]),.dinb(n2095),.dout(n2098),.clk(gclk));
	jnot g01889(.din(n2098),.dout(n2099),.clk(gclk));
	jand g01890(.dina(n2099),.dinb(n2093),.dout(n2100),.clk(gclk));
	jnot g01891(.din(w_n2100_0[1]),.dout(n2101),.clk(gclk));
	jor g01892(.dina(n2101),.dinb(w_n2085_0[1]),.dout(asqrt_fa_48),.clk(gclk));
	jnot g01893(.din(w_n1888_0[0]),.dout(n2103),.clk(gclk));
	jand g01894(.dina(w_n2091_0[0]),.dinb(w_n1891_0[0]),.dout(n2104),.clk(gclk));
	jand g01895(.dina(w_n2104_0[1]),.dinb(w_n1904_0[1]),.dout(n2105),.clk(gclk));
	jand g01896(.dina(n2105),.dinb(n2103),.dout(n2106),.clk(gclk));
	jor g01897(.dina(n2106),.dinb(w_asqrt63_49[0]),.dout(n2107),.clk(gclk));
	jand g01898(.dina(w_n2100_0[0]),.dinb(n2107),.dout(n2108),.clk(gclk));
	jor g01899(.dina(w_n2108_65[1]),.dinb(w_n1894_1[0]),.dout(n2109),.clk(gclk));
	jnot g01900(.din(w_a92_0[2]),.dout(n2110),.clk(gclk));
	jnot g01901(.din(w_a93_0[1]),.dout(n2111),.clk(gclk));
	jand g01902(.dina(w_n2111_0[1]),.dinb(w_n2110_1[2]),.dout(n2112),.clk(gclk));
	jand g01903(.dina(w_n2112_0[2]),.dinb(w_n1894_0[2]),.dout(n2113),.clk(gclk));
	jnot g01904(.din(w_n2113_0[1]),.dout(n2114),.clk(gclk));
	jand g01905(.dina(n2114),.dinb(n2109),.dout(n2115),.clk(gclk));
	jor g01906(.dina(w_n2115_0[2]),.dinb(w_n1912_59[0]),.dout(n2116),.clk(gclk));
	jand g01907(.dina(w_n2115_0[1]),.dinb(w_n1912_58[2]),.dout(n2117),.clk(gclk));
	jor g01908(.dina(w_n2108_65[0]),.dinb(w_a94_1[0]),.dout(n2118),.clk(gclk));
	jand g01909(.dina(n2118),.dinb(w_a95_0[0]),.dout(n2119),.clk(gclk));
	jand g01910(.dina(w_asqrt47_36),.dinb(w_n1896_0[1]),.dout(n2120),.clk(gclk));
	jor g01911(.dina(n2120),.dinb(n2119),.dout(n2121),.clk(gclk));
	jor g01912(.dina(n2121),.dinb(n2117),.dout(n2122),.clk(gclk));
	jand g01913(.dina(n2122),.dinb(w_n2116_0[1]),.dout(n2123),.clk(gclk));
	jor g01914(.dina(w_n2123_0[2]),.dinb(w_n1699_61[1]),.dout(n2124),.clk(gclk));
	jand g01915(.dina(w_n2123_0[1]),.dinb(w_n1699_61[0]),.dout(n2125),.clk(gclk));
	jnot g01916(.din(w_n1896_0[0]),.dout(n2126),.clk(gclk));
	jor g01917(.dina(w_n2108_64[2]),.dinb(n2126),.dout(n2127),.clk(gclk));
	jnot g01918(.din(w_n2092_0[1]),.dout(n2128),.clk(gclk));
	jor g01919(.dina(w_n2097_0[0]),.dinb(w_n2128_0[1]),.dout(n2129),.clk(gclk));
	jor g01920(.dina(n2129),.dinb(w_n2085_0[0]),.dout(n2130),.clk(gclk));
	jor g01921(.dina(n2130),.dinb(w_n1912_58[1]),.dout(n2131),.clk(gclk));
	jand g01922(.dina(n2131),.dinb(w_n2127_0[1]),.dout(n2132),.clk(gclk));
	jxor g01923(.dina(n2132),.dinb(w_n1681_0[1]),.dout(n2133),.clk(gclk));
	jor g01924(.dina(w_n2133_0[2]),.dinb(n2125),.dout(n2134),.clk(gclk));
	jand g01925(.dina(n2134),.dinb(w_n2124_0[1]),.dout(n2135),.clk(gclk));
	jor g01926(.dina(w_n2135_0[2]),.dinb(w_n1516_59[2]),.dout(n2136),.clk(gclk));
	jand g01927(.dina(w_n2135_0[1]),.dinb(w_n1516_59[1]),.dout(n2137),.clk(gclk));
	jxor g01928(.dina(w_n1898_0[0]),.dinb(w_n1699_60[2]),.dout(n2138),.clk(gclk));
	jor g01929(.dina(n2138),.dinb(w_n2108_64[1]),.dout(n2139),.clk(gclk));
	jxor g01930(.dina(n2139),.dinb(w_n2033_0[0]),.dout(n2140),.clk(gclk));
	jnot g01931(.din(w_n2140_0[2]),.dout(n2141),.clk(gclk));
	jor g01932(.dina(n2141),.dinb(n2137),.dout(n2142),.clk(gclk));
	jand g01933(.dina(n2142),.dinb(w_n2136_0[1]),.dout(n2143),.clk(gclk));
	jor g01934(.dina(w_n2143_0[2]),.dinb(w_n1332_61[1]),.dout(n2144),.clk(gclk));
	jand g01935(.dina(w_n2143_0[1]),.dinb(w_n1332_61[0]),.dout(n2145),.clk(gclk));
	jxor g01936(.dina(w_n1916_0[0]),.dinb(w_n1516_59[0]),.dout(n2146),.clk(gclk));
	jor g01937(.dina(n2146),.dinb(w_n2108_64[0]),.dout(n2147),.clk(gclk));
	jxor g01938(.dina(n2147),.dinb(w_n1925_0[0]),.dout(n2148),.clk(gclk));
	jor g01939(.dina(w_n2148_0[2]),.dinb(n2145),.dout(n2149),.clk(gclk));
	jand g01940(.dina(n2149),.dinb(w_n2144_0[1]),.dout(n2150),.clk(gclk));
	jor g01941(.dina(w_n2150_0[2]),.dinb(w_n1173_60[1]),.dout(n2151),.clk(gclk));
	jand g01942(.dina(w_n2150_0[1]),.dinb(w_n1173_60[0]),.dout(n2152),.clk(gclk));
	jxor g01943(.dina(w_n1927_0[0]),.dinb(w_n1332_60[2]),.dout(n2153),.clk(gclk));
	jor g01944(.dina(n2153),.dinb(w_n2108_63[2]),.dout(n2154),.clk(gclk));
	jxor g01945(.dina(n2154),.dinb(w_n2040_0[0]),.dout(n2155),.clk(gclk));
	jnot g01946(.din(w_n2155_0[2]),.dout(n2156),.clk(gclk));
	jor g01947(.dina(n2156),.dinb(n2152),.dout(n2157),.clk(gclk));
	jand g01948(.dina(n2157),.dinb(w_n2151_0[1]),.dout(n2158),.clk(gclk));
	jor g01949(.dina(w_n2158_0[2]),.dinb(w_n1008_62[1]),.dout(n2159),.clk(gclk));
	jand g01950(.dina(w_n2158_0[1]),.dinb(w_n1008_62[0]),.dout(n2160),.clk(gclk));
	jxor g01951(.dina(w_n1934_0[0]),.dinb(w_n1173_59[2]),.dout(n2161),.clk(gclk));
	jor g01952(.dina(n2161),.dinb(w_n2108_63[1]),.dout(n2162),.clk(gclk));
	jxor g01953(.dina(n2162),.dinb(w_n1940_0[0]),.dout(n2163),.clk(gclk));
	jor g01954(.dina(w_n2163_0[2]),.dinb(n2160),.dout(n2164),.clk(gclk));
	jand g01955(.dina(n2164),.dinb(w_n2159_0[1]),.dout(n2165),.clk(gclk));
	jor g01956(.dina(w_n2165_0[2]),.dinb(w_n884_61[1]),.dout(n2166),.clk(gclk));
	jand g01957(.dina(w_n2165_0[1]),.dinb(w_n884_61[0]),.dout(n2167),.clk(gclk));
	jxor g01958(.dina(w_n1942_0[0]),.dinb(w_n1008_61[2]),.dout(n2168),.clk(gclk));
	jor g01959(.dina(n2168),.dinb(w_n2108_63[0]),.dout(n2169),.clk(gclk));
	jxor g01960(.dina(n2169),.dinb(w_n1948_0[0]),.dout(n2170),.clk(gclk));
	jor g01961(.dina(w_n2170_0[2]),.dinb(n2167),.dout(n2171),.clk(gclk));
	jand g01962(.dina(n2171),.dinb(w_n2166_0[1]),.dout(n2172),.clk(gclk));
	jor g01963(.dina(w_n2172_0[2]),.dinb(w_n743_62[1]),.dout(n2173),.clk(gclk));
	jand g01964(.dina(w_n2172_0[1]),.dinb(w_n743_62[0]),.dout(n2174),.clk(gclk));
	jxor g01965(.dina(w_n1950_0[0]),.dinb(w_n884_60[2]),.dout(n2175),.clk(gclk));
	jor g01966(.dina(n2175),.dinb(w_n2108_62[2]),.dout(n2176),.clk(gclk));
	jxor g01967(.dina(n2176),.dinb(w_n2050_0[0]),.dout(n2177),.clk(gclk));
	jnot g01968(.din(w_n2177_0[2]),.dout(n2178),.clk(gclk));
	jor g01969(.dina(n2178),.dinb(n2174),.dout(n2179),.clk(gclk));
	jand g01970(.dina(n2179),.dinb(w_n2173_0[1]),.dout(n2180),.clk(gclk));
	jor g01971(.dina(w_n2180_0[2]),.dinb(w_n635_62[1]),.dout(n2181),.clk(gclk));
	jand g01972(.dina(w_n2180_0[1]),.dinb(w_n635_62[0]),.dout(n2182),.clk(gclk));
	jxor g01973(.dina(w_n1957_0[0]),.dinb(w_n743_61[2]),.dout(n2183),.clk(gclk));
	jor g01974(.dina(n2183),.dinb(w_n2108_62[1]),.dout(n2184),.clk(gclk));
	jxor g01975(.dina(n2184),.dinb(w_n2054_0[0]),.dout(n2185),.clk(gclk));
	jnot g01976(.din(w_n2185_0[2]),.dout(n2186),.clk(gclk));
	jor g01977(.dina(n2186),.dinb(n2182),.dout(n2187),.clk(gclk));
	jand g01978(.dina(n2187),.dinb(w_n2181_0[1]),.dout(n2188),.clk(gclk));
	jor g01979(.dina(w_n2188_0[2]),.dinb(w_n515_63[1]),.dout(n2189),.clk(gclk));
	jand g01980(.dina(w_n2188_0[1]),.dinb(w_n515_63[0]),.dout(n2190),.clk(gclk));
	jxor g01981(.dina(w_n1964_0[0]),.dinb(w_n635_61[2]),.dout(n2191),.clk(gclk));
	jor g01982(.dina(n2191),.dinb(w_n2108_62[0]),.dout(n2192),.clk(gclk));
	jxor g01983(.dina(n2192),.dinb(w_n1970_0[0]),.dout(n2193),.clk(gclk));
	jor g01984(.dina(w_n2193_0[2]),.dinb(n2190),.dout(n2194),.clk(gclk));
	jand g01985(.dina(n2194),.dinb(w_n2189_0[1]),.dout(n2195),.clk(gclk));
	jor g01986(.dina(w_n2195_0[2]),.dinb(w_n443_63[1]),.dout(n2196),.clk(gclk));
	jand g01987(.dina(w_n2195_0[1]),.dinb(w_n443_63[0]),.dout(n2197),.clk(gclk));
	jxor g01988(.dina(w_n1972_0[0]),.dinb(w_n515_62[2]),.dout(n2198),.clk(gclk));
	jor g01989(.dina(n2198),.dinb(w_n2108_61[2]),.dout(n2199),.clk(gclk));
	jxor g01990(.dina(n2199),.dinb(w_n1978_0[0]),.dout(n2200),.clk(gclk));
	jor g01991(.dina(w_n2200_0[1]),.dinb(n2197),.dout(n2201),.clk(gclk));
	jand g01992(.dina(n2201),.dinb(w_n2196_0[1]),.dout(n2202),.clk(gclk));
	jor g01993(.dina(w_n2202_0[2]),.dinb(w_n352_63[2]),.dout(n2203),.clk(gclk));
	jand g01994(.dina(w_n2202_0[1]),.dinb(w_n352_63[1]),.dout(n2204),.clk(gclk));
	jxor g01995(.dina(w_n1980_0[0]),.dinb(w_n443_62[2]),.dout(n2205),.clk(gclk));
	jor g01996(.dina(n2205),.dinb(w_n2108_61[1]),.dout(n2206),.clk(gclk));
	jxor g01997(.dina(n2206),.dinb(w_n1985_0[0]),.dout(n2207),.clk(gclk));
	jnot g01998(.din(w_n2207_0[2]),.dout(n2208),.clk(gclk));
	jor g01999(.dina(n2208),.dinb(n2204),.dout(n2209),.clk(gclk));
	jand g02000(.dina(n2209),.dinb(w_n2203_0[1]),.dout(n2210),.clk(gclk));
	jor g02001(.dina(w_n2210_0[2]),.dinb(w_n294_64[0]),.dout(n2211),.clk(gclk));
	jand g02002(.dina(w_n2210_0[1]),.dinb(w_n294_63[2]),.dout(n2212),.clk(gclk));
	jxor g02003(.dina(w_n1988_0[0]),.dinb(w_n352_63[0]),.dout(n2213),.clk(gclk));
	jor g02004(.dina(n2213),.dinb(w_n2108_61[0]),.dout(n2214),.clk(gclk));
	jxor g02005(.dina(n2214),.dinb(w_n2067_0[0]),.dout(n2215),.clk(gclk));
	jnot g02006(.din(w_n2215_0[2]),.dout(n2216),.clk(gclk));
	jor g02007(.dina(n2216),.dinb(n2212),.dout(n2217),.clk(gclk));
	jand g02008(.dina(n2217),.dinb(w_n2211_0[1]),.dout(n2218),.clk(gclk));
	jor g02009(.dina(w_n2218_0[2]),.dinb(w_n239_64[0]),.dout(n2219),.clk(gclk));
	jand g02010(.dina(w_n2218_0[1]),.dinb(w_n239_63[2]),.dout(n2220),.clk(gclk));
	jxor g02011(.dina(w_n1995_0[0]),.dinb(w_n294_63[1]),.dout(n2221),.clk(gclk));
	jor g02012(.dina(n2221),.dinb(w_n2108_60[2]),.dout(n2222),.clk(gclk));
	jxor g02013(.dina(n2222),.dinb(w_n2001_0[0]),.dout(n2223),.clk(gclk));
	jor g02014(.dina(w_n2223_0[2]),.dinb(n2220),.dout(n2224),.clk(gclk));
	jand g02015(.dina(n2224),.dinb(w_n2219_0[1]),.dout(n2225),.clk(gclk));
	jor g02016(.dina(w_n2225_0[2]),.dinb(w_n221_64[1]),.dout(n2226),.clk(gclk));
	jand g02017(.dina(w_n2225_0[1]),.dinb(w_n221_64[0]),.dout(n2227),.clk(gclk));
	jxor g02018(.dina(w_n2003_0[0]),.dinb(w_n239_63[1]),.dout(n2228),.clk(gclk));
	jor g02019(.dina(n2228),.dinb(w_n2108_60[1]),.dout(n2229),.clk(gclk));
	jxor g02020(.dina(n2229),.dinb(w_n2009_0[0]),.dout(n2230),.clk(gclk));
	jor g02021(.dina(w_n2230_0[2]),.dinb(n2227),.dout(n2231),.clk(gclk));
	jand g02022(.dina(n2231),.dinb(w_n2226_0[1]),.dout(n2232),.clk(gclk));
	jxor g02023(.dina(w_n2011_0[0]),.dinb(w_n221_63[2]),.dout(n2233),.clk(gclk));
	jor g02024(.dina(n2233),.dinb(w_n2108_60[0]),.dout(n2234),.clk(gclk));
	jxor g02025(.dina(n2234),.dinb(w_n2089_0[0]),.dout(n2235),.clk(gclk));
	jand g02026(.dina(w_n2235_1[1]),.dinb(w_n2232_0[2]),.dout(n2236),.clk(gclk));
	jor g02027(.dina(w_n2235_1[0]),.dinb(w_n2232_0[1]),.dout(n2238),.clk(gclk));
	jand g02028(.dina(w_asqrt47_35[2]),.dinb(w_n2104_0[0]),.dout(n2239),.clk(gclk));
	jor g02029(.dina(n2239),.dinb(w_n2128_0[0]),.dout(n2240),.clk(gclk));
	jor g02030(.dina(w_n2240_0[1]),.dinb(w_n2238_0[1]),.dout(n2241),.clk(gclk));
	jand g02031(.dina(n2241),.dinb(w_n218_26[1]),.dout(n2242),.clk(gclk));
	jand g02032(.dina(w_n2108_59[2]),.dinb(w_n2081_0[0]),.dout(n2243),.clk(gclk));
	jand g02033(.dina(w_n2082_0[0]),.dinb(w_asqrt63_48[2]),.dout(n2244),.clk(gclk));
	jand g02034(.dina(n2244),.dinb(w_n2092_0[0]),.dout(n2245),.clk(gclk));
	jnot g02035(.din(n2245),.dout(n2246),.clk(gclk));
	jor g02036(.dina(w_n2246_0[1]),.dinb(n2243),.dout(n2247),.clk(gclk));
	jnot g02037(.din(w_n2247_0[1]),.dout(n2248),.clk(gclk));
	jor g02038(.dina(n2248),.dinb(n2242),.dout(n2249),.clk(gclk));
	jor g02039(.dina(w_n2249_0[1]),.dinb(w_n2236_0[2]),.dout(asqrt_fa_47),.clk(gclk));
	jnot g02040(.din(w_a90_1[1]),.dout(n2252),.clk(gclk));
	jnot g02041(.din(w_a91_0[1]),.dout(n2253),.clk(gclk));
	jand g02042(.dina(w_n2253_0[1]),.dinb(w_n2252_1[1]),.dout(n2254),.clk(gclk));
	jand g02043(.dina(w_n2254_0[2]),.dinb(w_n2110_1[1]),.dout(n2255),.clk(gclk));
	jand g02044(.dina(w_asqrt46_41[1]),.dinb(w_a92_0[1]),.dout(n2256),.clk(gclk));
	jor g02045(.dina(n2256),.dinb(w_n2255_0[1]),.dout(n2257),.clk(gclk));
	jand g02046(.dina(w_n2257_0[2]),.dinb(w_asqrt47_35[1]),.dout(n2258),.clk(gclk));
	jor g02047(.dina(w_n2257_0[1]),.dinb(w_asqrt47_35[0]),.dout(n2259),.clk(gclk));
	jand g02048(.dina(w_asqrt46_41[0]),.dinb(w_n2110_1[0]),.dout(n2260),.clk(gclk));
	jor g02049(.dina(n2260),.dinb(w_n2111_0[0]),.dout(n2261),.clk(gclk));
	jnot g02050(.din(w_n2112_0[1]),.dout(n2262),.clk(gclk));
	jnot g02051(.din(w_n2236_0[1]),.dout(n2263),.clk(gclk));
	jnot g02052(.din(w_n2226_0[0]),.dout(n2265),.clk(gclk));
	jnot g02053(.din(w_n2219_0[0]),.dout(n2266),.clk(gclk));
	jnot g02054(.din(w_n2211_0[0]),.dout(n2267),.clk(gclk));
	jnot g02055(.din(w_n2203_0[0]),.dout(n2268),.clk(gclk));
	jnot g02056(.din(w_n2196_0[0]),.dout(n2269),.clk(gclk));
	jnot g02057(.din(w_n2189_0[0]),.dout(n2270),.clk(gclk));
	jnot g02058(.din(w_n2181_0[0]),.dout(n2271),.clk(gclk));
	jnot g02059(.din(w_n2173_0[0]),.dout(n2272),.clk(gclk));
	jnot g02060(.din(w_n2166_0[0]),.dout(n2273),.clk(gclk));
	jnot g02061(.din(w_n2159_0[0]),.dout(n2274),.clk(gclk));
	jnot g02062(.din(w_n2151_0[0]),.dout(n2275),.clk(gclk));
	jnot g02063(.din(w_n2144_0[0]),.dout(n2276),.clk(gclk));
	jnot g02064(.din(w_n2136_0[0]),.dout(n2277),.clk(gclk));
	jnot g02065(.din(w_n2124_0[0]),.dout(n2278),.clk(gclk));
	jnot g02066(.din(w_n2116_0[0]),.dout(n2279),.clk(gclk));
	jand g02067(.dina(w_asqrt47_34[2]),.dinb(w_a94_0[2]),.dout(n2280),.clk(gclk));
	jor g02068(.dina(w_n2113_0[0]),.dinb(n2280),.dout(n2281),.clk(gclk));
	jor g02069(.dina(n2281),.dinb(w_asqrt48_36[2]),.dout(n2282),.clk(gclk));
	jand g02070(.dina(w_asqrt47_34[1]),.dinb(w_n1894_0[1]),.dout(n2283),.clk(gclk));
	jor g02071(.dina(n2283),.dinb(w_n1895_0[0]),.dout(n2284),.clk(gclk));
	jand g02072(.dina(w_n2127_0[0]),.dinb(n2284),.dout(n2285),.clk(gclk));
	jand g02073(.dina(w_n2285_0[1]),.dinb(n2282),.dout(n2286),.clk(gclk));
	jor g02074(.dina(n2286),.dinb(n2279),.dout(n2287),.clk(gclk));
	jor g02075(.dina(n2287),.dinb(w_asqrt49_35[0]),.dout(n2288),.clk(gclk));
	jnot g02076(.din(w_n2133_0[1]),.dout(n2289),.clk(gclk));
	jand g02077(.dina(n2289),.dinb(n2288),.dout(n2290),.clk(gclk));
	jor g02078(.dina(n2290),.dinb(n2278),.dout(n2291),.clk(gclk));
	jor g02079(.dina(n2291),.dinb(w_asqrt50_37[0]),.dout(n2292),.clk(gclk));
	jand g02080(.dina(w_n2140_0[1]),.dinb(n2292),.dout(n2293),.clk(gclk));
	jor g02081(.dina(n2293),.dinb(n2277),.dout(n2294),.clk(gclk));
	jor g02082(.dina(n2294),.dinb(w_asqrt51_35[1]),.dout(n2295),.clk(gclk));
	jnot g02083(.din(w_n2148_0[1]),.dout(n2296),.clk(gclk));
	jand g02084(.dina(n2296),.dinb(n2295),.dout(n2297),.clk(gclk));
	jor g02085(.dina(n2297),.dinb(n2276),.dout(n2298),.clk(gclk));
	jor g02086(.dina(n2298),.dinb(w_asqrt52_37[0]),.dout(n2299),.clk(gclk));
	jand g02087(.dina(w_n2155_0[1]),.dinb(n2299),.dout(n2300),.clk(gclk));
	jor g02088(.dina(n2300),.dinb(n2275),.dout(n2301),.clk(gclk));
	jor g02089(.dina(n2301),.dinb(w_asqrt53_36[0]),.dout(n2302),.clk(gclk));
	jnot g02090(.din(w_n2163_0[1]),.dout(n2303),.clk(gclk));
	jand g02091(.dina(n2303),.dinb(n2302),.dout(n2304),.clk(gclk));
	jor g02092(.dina(n2304),.dinb(n2274),.dout(n2305),.clk(gclk));
	jor g02093(.dina(n2305),.dinb(w_asqrt54_37[0]),.dout(n2306),.clk(gclk));
	jnot g02094(.din(w_n2170_0[1]),.dout(n2307),.clk(gclk));
	jand g02095(.dina(n2307),.dinb(n2306),.dout(n2308),.clk(gclk));
	jor g02096(.dina(n2308),.dinb(n2273),.dout(n2309),.clk(gclk));
	jor g02097(.dina(n2309),.dinb(w_asqrt55_36[1]),.dout(n2310),.clk(gclk));
	jand g02098(.dina(w_n2177_0[1]),.dinb(n2310),.dout(n2311),.clk(gclk));
	jor g02099(.dina(n2311),.dinb(n2272),.dout(n2312),.clk(gclk));
	jor g02100(.dina(n2312),.dinb(w_asqrt56_37[1]),.dout(n2313),.clk(gclk));
	jand g02101(.dina(w_n2185_0[1]),.dinb(n2313),.dout(n2314),.clk(gclk));
	jor g02102(.dina(n2314),.dinb(n2271),.dout(n2315),.clk(gclk));
	jor g02103(.dina(n2315),.dinb(w_asqrt57_37[0]),.dout(n2316),.clk(gclk));
	jnot g02104(.din(w_n2193_0[1]),.dout(n2317),.clk(gclk));
	jand g02105(.dina(n2317),.dinb(n2316),.dout(n2318),.clk(gclk));
	jor g02106(.dina(n2318),.dinb(n2270),.dout(n2319),.clk(gclk));
	jor g02107(.dina(n2319),.dinb(w_asqrt58_37[2]),.dout(n2320),.clk(gclk));
	jnot g02108(.din(w_n2200_0[0]),.dout(n2321),.clk(gclk));
	jand g02109(.dina(w_n2321_0[1]),.dinb(n2320),.dout(n2322),.clk(gclk));
	jor g02110(.dina(n2322),.dinb(n2269),.dout(n2323),.clk(gclk));
	jor g02111(.dina(n2323),.dinb(w_asqrt59_37[1]),.dout(n2324),.clk(gclk));
	jand g02112(.dina(w_n2207_0[1]),.dinb(n2324),.dout(n2325),.clk(gclk));
	jor g02113(.dina(n2325),.dinb(n2268),.dout(n2326),.clk(gclk));
	jor g02114(.dina(n2326),.dinb(w_asqrt60_37[2]),.dout(n2327),.clk(gclk));
	jand g02115(.dina(w_n2215_0[1]),.dinb(n2327),.dout(n2328),.clk(gclk));
	jor g02116(.dina(n2328),.dinb(n2267),.dout(n2329),.clk(gclk));
	jor g02117(.dina(n2329),.dinb(w_asqrt61_37[2]),.dout(n2330),.clk(gclk));
	jnot g02118(.din(w_n2223_0[1]),.dout(n2331),.clk(gclk));
	jand g02119(.dina(n2331),.dinb(n2330),.dout(n2332),.clk(gclk));
	jor g02120(.dina(n2332),.dinb(n2266),.dout(n2333),.clk(gclk));
	jor g02121(.dina(n2333),.dinb(w_asqrt62_37[2]),.dout(n2334),.clk(gclk));
	jnot g02122(.din(w_n2230_0[1]),.dout(n2335),.clk(gclk));
	jand g02123(.dina(n2335),.dinb(n2334),.dout(n2336),.clk(gclk));
	jor g02124(.dina(n2336),.dinb(n2265),.dout(n2337),.clk(gclk));
	jnot g02125(.din(w_n2235_0[2]),.dout(n2338),.clk(gclk));
	jand g02126(.dina(n2338),.dinb(n2337),.dout(n2339),.clk(gclk));
	jnot g02127(.din(w_n2240_0[0]),.dout(n2340),.clk(gclk));
	jand g02128(.dina(n2340),.dinb(w_n2339_0[1]),.dout(n2341),.clk(gclk));
	jor g02129(.dina(n2341),.dinb(w_asqrt63_48[1]),.dout(n2342),.clk(gclk));
	jand g02130(.dina(w_n2247_0[0]),.dinb(w_n2342_0[1]),.dout(n2343),.clk(gclk));
	jand g02131(.dina(w_n2343_0[1]),.dinb(w_n2263_1[1]),.dout(n2345),.clk(gclk));
	jor g02132(.dina(w_n2345_57[2]),.dinb(n2262),.dout(n2346),.clk(gclk));
	jand g02133(.dina(n2346),.dinb(n2261),.dout(n2347),.clk(gclk));
	jand g02134(.dina(n2347),.dinb(n2259),.dout(n2348),.clk(gclk));
	jor g02135(.dina(n2348),.dinb(w_n2258_0[1]),.dout(n2349),.clk(gclk));
	jand g02136(.dina(w_n2349_0[2]),.dinb(w_asqrt48_36[1]),.dout(n2350),.clk(gclk));
	jor g02137(.dina(w_n2349_0[1]),.dinb(w_asqrt48_36[0]),.dout(n2351),.clk(gclk));
	jand g02138(.dina(w_asqrt46_40[2]),.dinb(w_n2112_0[0]),.dout(n2352),.clk(gclk));
	jand g02139(.dina(w_n2263_1[0]),.dinb(w_asqrt47_34[0]),.dout(n2353),.clk(gclk));
	jand g02140(.dina(n2353),.dinb(w_n2246_0[0]),.dout(n2354),.clk(gclk));
	jand g02141(.dina(n2354),.dinb(w_n2342_0[0]),.dout(n2355),.clk(gclk));
	jor g02142(.dina(n2355),.dinb(w_n2352_0[1]),.dout(n2356),.clk(gclk));
	jxor g02143(.dina(n2356),.dinb(w_a94_0[1]),.dout(n2357),.clk(gclk));
	jnot g02144(.din(w_n2357_0[1]),.dout(n2358),.clk(gclk));
	jand g02145(.dina(w_n2358_0[1]),.dinb(n2351),.dout(n2359),.clk(gclk));
	jor g02146(.dina(n2359),.dinb(w_n2350_0[1]),.dout(n2360),.clk(gclk));
	jand g02147(.dina(w_n2360_0[2]),.dinb(w_asqrt49_34[2]),.dout(n2361),.clk(gclk));
	jor g02148(.dina(w_n2360_0[1]),.dinb(w_asqrt49_34[1]),.dout(n2362),.clk(gclk));
	jxor g02149(.dina(w_n2115_0[0]),.dinb(w_n1912_58[0]),.dout(n2363),.clk(gclk));
	jand g02150(.dina(n2363),.dinb(w_asqrt46_40[1]),.dout(n2364),.clk(gclk));
	jxor g02151(.dina(n2364),.dinb(w_n2285_0[0]),.dout(n2365),.clk(gclk));
	jand g02152(.dina(w_n2365_0[1]),.dinb(n2362),.dout(n2366),.clk(gclk));
	jor g02153(.dina(n2366),.dinb(w_n2361_0[1]),.dout(n2367),.clk(gclk));
	jand g02154(.dina(w_n2367_0[2]),.dinb(w_asqrt50_36[2]),.dout(n2368),.clk(gclk));
	jor g02155(.dina(w_n2367_0[1]),.dinb(w_asqrt50_36[1]),.dout(n2369),.clk(gclk));
	jxor g02156(.dina(w_n2123_0[0]),.dinb(w_n1699_60[1]),.dout(n2370),.clk(gclk));
	jand g02157(.dina(n2370),.dinb(w_asqrt46_40[0]),.dout(n2371),.clk(gclk));
	jxor g02158(.dina(n2371),.dinb(w_n2133_0[0]),.dout(n2372),.clk(gclk));
	jnot g02159(.din(w_n2372_0[1]),.dout(n2373),.clk(gclk));
	jand g02160(.dina(w_n2373_0[1]),.dinb(n2369),.dout(n2374),.clk(gclk));
	jor g02161(.dina(n2374),.dinb(w_n2368_0[1]),.dout(n2375),.clk(gclk));
	jand g02162(.dina(w_n2375_0[2]),.dinb(w_asqrt51_35[0]),.dout(n2376),.clk(gclk));
	jor g02163(.dina(w_n2375_0[1]),.dinb(w_asqrt51_34[2]),.dout(n2377),.clk(gclk));
	jxor g02164(.dina(w_n2135_0[0]),.dinb(w_n1516_58[2]),.dout(n2378),.clk(gclk));
	jand g02165(.dina(n2378),.dinb(w_asqrt46_39[2]),.dout(n2379),.clk(gclk));
	jxor g02166(.dina(n2379),.dinb(w_n2140_0[0]),.dout(n2380),.clk(gclk));
	jand g02167(.dina(w_n2380_0[1]),.dinb(n2377),.dout(n2381),.clk(gclk));
	jor g02168(.dina(n2381),.dinb(w_n2376_0[1]),.dout(n2382),.clk(gclk));
	jand g02169(.dina(w_n2382_0[2]),.dinb(w_asqrt52_36[2]),.dout(n2383),.clk(gclk));
	jor g02170(.dina(w_n2382_0[1]),.dinb(w_asqrt52_36[1]),.dout(n2384),.clk(gclk));
	jxor g02171(.dina(w_n2143_0[0]),.dinb(w_n1332_60[1]),.dout(n2385),.clk(gclk));
	jand g02172(.dina(n2385),.dinb(w_asqrt46_39[1]),.dout(n2386),.clk(gclk));
	jxor g02173(.dina(n2386),.dinb(w_n2148_0[0]),.dout(n2387),.clk(gclk));
	jnot g02174(.din(w_n2387_0[1]),.dout(n2388),.clk(gclk));
	jand g02175(.dina(w_n2388_0[1]),.dinb(n2384),.dout(n2389),.clk(gclk));
	jor g02176(.dina(n2389),.dinb(w_n2383_0[1]),.dout(n2390),.clk(gclk));
	jand g02177(.dina(w_n2390_0[2]),.dinb(w_asqrt53_35[2]),.dout(n2391),.clk(gclk));
	jor g02178(.dina(w_n2390_0[1]),.dinb(w_asqrt53_35[1]),.dout(n2392),.clk(gclk));
	jxor g02179(.dina(w_n2150_0[0]),.dinb(w_n1173_59[1]),.dout(n2393),.clk(gclk));
	jand g02180(.dina(n2393),.dinb(w_asqrt46_39[0]),.dout(n2394),.clk(gclk));
	jxor g02181(.dina(n2394),.dinb(w_n2155_0[0]),.dout(n2395),.clk(gclk));
	jand g02182(.dina(w_n2395_0[1]),.dinb(n2392),.dout(n2396),.clk(gclk));
	jor g02183(.dina(n2396),.dinb(w_n2391_0[1]),.dout(n2397),.clk(gclk));
	jand g02184(.dina(w_n2397_0[2]),.dinb(w_asqrt54_36[2]),.dout(n2398),.clk(gclk));
	jor g02185(.dina(w_n2397_0[1]),.dinb(w_asqrt54_36[1]),.dout(n2399),.clk(gclk));
	jxor g02186(.dina(w_n2158_0[0]),.dinb(w_n1008_61[1]),.dout(n2400),.clk(gclk));
	jand g02187(.dina(n2400),.dinb(w_asqrt46_38[2]),.dout(n2401),.clk(gclk));
	jxor g02188(.dina(n2401),.dinb(w_n2163_0[0]),.dout(n2402),.clk(gclk));
	jnot g02189(.din(w_n2402_0[1]),.dout(n2403),.clk(gclk));
	jand g02190(.dina(w_n2403_0[1]),.dinb(n2399),.dout(n2404),.clk(gclk));
	jor g02191(.dina(n2404),.dinb(w_n2398_0[1]),.dout(n2405),.clk(gclk));
	jand g02192(.dina(w_n2405_0[2]),.dinb(w_asqrt55_36[0]),.dout(n2406),.clk(gclk));
	jor g02193(.dina(w_n2405_0[1]),.dinb(w_asqrt55_35[2]),.dout(n2407),.clk(gclk));
	jxor g02194(.dina(w_n2165_0[0]),.dinb(w_n884_60[1]),.dout(n2408),.clk(gclk));
	jand g02195(.dina(n2408),.dinb(w_asqrt46_38[1]),.dout(n2409),.clk(gclk));
	jxor g02196(.dina(n2409),.dinb(w_n2170_0[0]),.dout(n2410),.clk(gclk));
	jnot g02197(.din(w_n2410_0[1]),.dout(n2411),.clk(gclk));
	jand g02198(.dina(w_n2411_0[1]),.dinb(n2407),.dout(n2412),.clk(gclk));
	jor g02199(.dina(n2412),.dinb(w_n2406_0[1]),.dout(n2413),.clk(gclk));
	jand g02200(.dina(w_n2413_0[2]),.dinb(w_asqrt56_37[0]),.dout(n2414),.clk(gclk));
	jor g02201(.dina(w_n2413_0[1]),.dinb(w_asqrt56_36[2]),.dout(n2415),.clk(gclk));
	jxor g02202(.dina(w_n2172_0[0]),.dinb(w_n743_61[1]),.dout(n2416),.clk(gclk));
	jand g02203(.dina(n2416),.dinb(w_asqrt46_38[0]),.dout(n2417),.clk(gclk));
	jxor g02204(.dina(n2417),.dinb(w_n2177_0[0]),.dout(n2418),.clk(gclk));
	jand g02205(.dina(w_n2418_0[1]),.dinb(n2415),.dout(n2419),.clk(gclk));
	jor g02206(.dina(n2419),.dinb(w_n2414_0[1]),.dout(n2420),.clk(gclk));
	jand g02207(.dina(w_n2420_0[2]),.dinb(w_asqrt57_36[2]),.dout(n2421),.clk(gclk));
	jor g02208(.dina(w_n2420_0[1]),.dinb(w_asqrt57_36[1]),.dout(n2422),.clk(gclk));
	jxor g02209(.dina(w_n2180_0[0]),.dinb(w_n635_61[1]),.dout(n2423),.clk(gclk));
	jand g02210(.dina(n2423),.dinb(w_asqrt46_37[2]),.dout(n2424),.clk(gclk));
	jxor g02211(.dina(n2424),.dinb(w_n2185_0[0]),.dout(n2425),.clk(gclk));
	jand g02212(.dina(w_n2425_0[1]),.dinb(n2422),.dout(n2426),.clk(gclk));
	jor g02213(.dina(n2426),.dinb(w_n2421_0[1]),.dout(n2427),.clk(gclk));
	jand g02214(.dina(w_n2427_0[2]),.dinb(w_asqrt58_37[1]),.dout(n2428),.clk(gclk));
	jor g02215(.dina(w_n2427_0[1]),.dinb(w_asqrt58_37[0]),.dout(n2429),.clk(gclk));
	jxor g02216(.dina(w_n2188_0[0]),.dinb(w_n515_62[1]),.dout(n2430),.clk(gclk));
	jand g02217(.dina(n2430),.dinb(w_asqrt46_37[1]),.dout(n2431),.clk(gclk));
	jxor g02218(.dina(n2431),.dinb(w_n2193_0[0]),.dout(n2432),.clk(gclk));
	jnot g02219(.din(w_n2432_0[1]),.dout(n2433),.clk(gclk));
	jand g02220(.dina(w_n2433_0[1]),.dinb(n2429),.dout(n2434),.clk(gclk));
	jor g02221(.dina(n2434),.dinb(w_n2428_0[1]),.dout(n2435),.clk(gclk));
	jand g02222(.dina(w_n2435_0[2]),.dinb(w_asqrt59_37[0]),.dout(n2436),.clk(gclk));
	jor g02223(.dina(w_n2435_0[1]),.dinb(w_asqrt59_36[2]),.dout(n2437),.clk(gclk));
	jxor g02224(.dina(w_n2195_0[0]),.dinb(w_n443_62[1]),.dout(n2438),.clk(gclk));
	jand g02225(.dina(n2438),.dinb(w_asqrt46_37[0]),.dout(n2439),.clk(gclk));
	jxor g02226(.dina(n2439),.dinb(w_n2321_0[0]),.dout(n2440),.clk(gclk));
	jand g02227(.dina(w_n2440_0[1]),.dinb(n2437),.dout(n2441),.clk(gclk));
	jor g02228(.dina(n2441),.dinb(w_n2436_0[1]),.dout(n2442),.clk(gclk));
	jand g02229(.dina(w_n2442_0[2]),.dinb(w_asqrt60_37[1]),.dout(n2443),.clk(gclk));
	jor g02230(.dina(w_n2442_0[1]),.dinb(w_asqrt60_37[0]),.dout(n2444),.clk(gclk));
	jxor g02231(.dina(w_n2202_0[0]),.dinb(w_n352_62[2]),.dout(n2445),.clk(gclk));
	jand g02232(.dina(n2445),.dinb(w_asqrt46_36[2]),.dout(n2446),.clk(gclk));
	jxor g02233(.dina(n2446),.dinb(w_n2207_0[0]),.dout(n2447),.clk(gclk));
	jand g02234(.dina(w_n2447_0[1]),.dinb(n2444),.dout(n2448),.clk(gclk));
	jor g02235(.dina(n2448),.dinb(w_n2443_0[1]),.dout(n2449),.clk(gclk));
	jand g02236(.dina(w_n2449_0[2]),.dinb(w_asqrt61_37[1]),.dout(n2450),.clk(gclk));
	jor g02237(.dina(w_n2449_0[1]),.dinb(w_asqrt61_37[0]),.dout(n2451),.clk(gclk));
	jxor g02238(.dina(w_n2210_0[0]),.dinb(w_n294_63[0]),.dout(n2452),.clk(gclk));
	jand g02239(.dina(n2452),.dinb(w_asqrt46_36[1]),.dout(n2453),.clk(gclk));
	jxor g02240(.dina(n2453),.dinb(w_n2215_0[0]),.dout(n2454),.clk(gclk));
	jand g02241(.dina(w_n2454_0[1]),.dinb(n2451),.dout(n2455),.clk(gclk));
	jor g02242(.dina(n2455),.dinb(w_n2450_0[1]),.dout(n2456),.clk(gclk));
	jand g02243(.dina(w_n2456_0[2]),.dinb(w_asqrt62_37[1]),.dout(n2457),.clk(gclk));
	jor g02244(.dina(w_n2456_0[1]),.dinb(w_asqrt62_37[0]),.dout(n2458),.clk(gclk));
	jxor g02245(.dina(w_n2218_0[0]),.dinb(w_n239_63[0]),.dout(n2459),.clk(gclk));
	jand g02246(.dina(n2459),.dinb(w_asqrt46_36[0]),.dout(n2460),.clk(gclk));
	jxor g02247(.dina(n2460),.dinb(w_n2223_0[0]),.dout(n2461),.clk(gclk));
	jnot g02248(.din(w_n2461_0[2]),.dout(n2462),.clk(gclk));
	jand g02249(.dina(n2462),.dinb(n2458),.dout(n2463),.clk(gclk));
	jor g02250(.dina(n2463),.dinb(w_n2457_0[1]),.dout(n2464),.clk(gclk));
	jxor g02251(.dina(w_n2225_0[0]),.dinb(w_n221_63[1]),.dout(n2465),.clk(gclk));
	jand g02252(.dina(n2465),.dinb(w_asqrt46_35[2]),.dout(n2466),.clk(gclk));
	jxor g02253(.dina(n2466),.dinb(w_n2230_0[0]),.dout(n2467),.clk(gclk));
	jnot g02254(.din(w_n2467_0[1]),.dout(n2468),.clk(gclk));
	jor g02255(.dina(w_n2468_0[1]),.dinb(w_n2464_0[1]),.dout(n2469),.clk(gclk));
	jnot g02256(.din(w_n2469_1[1]),.dout(n2470),.clk(gclk));
	jand g02257(.dina(w_n2343_0[0]),.dinb(w_n2232_0[0]),.dout(n2471),.clk(gclk));
	jnot g02258(.din(n2471),.dout(n2472),.clk(gclk));
	jand g02259(.dina(w_n2238_0[0]),.dinb(w_asqrt63_48[0]),.dout(n2473),.clk(gclk));
	jand g02260(.dina(n2473),.dinb(w_n2263_0[2]),.dout(n2474),.clk(gclk));
	jand g02261(.dina(w_n2474_0[1]),.dinb(n2472),.dout(n2475),.clk(gclk));
	jand g02262(.dina(w_n2249_0[0]),.dinb(w_n2339_0[0]),.dout(n2476),.clk(gclk));
	jnot g02263(.din(w_n2457_0[0]),.dout(n2477),.clk(gclk));
	jnot g02264(.din(w_n2450_0[0]),.dout(n2478),.clk(gclk));
	jnot g02265(.din(w_n2443_0[0]),.dout(n2479),.clk(gclk));
	jnot g02266(.din(w_n2436_0[0]),.dout(n2480),.clk(gclk));
	jnot g02267(.din(w_n2428_0[0]),.dout(n2481),.clk(gclk));
	jnot g02268(.din(w_n2421_0[0]),.dout(n2482),.clk(gclk));
	jnot g02269(.din(w_n2414_0[0]),.dout(n2483),.clk(gclk));
	jnot g02270(.din(w_n2406_0[0]),.dout(n2484),.clk(gclk));
	jnot g02271(.din(w_n2398_0[0]),.dout(n2485),.clk(gclk));
	jnot g02272(.din(w_n2391_0[0]),.dout(n2486),.clk(gclk));
	jnot g02273(.din(w_n2383_0[0]),.dout(n2487),.clk(gclk));
	jnot g02274(.din(w_n2376_0[0]),.dout(n2488),.clk(gclk));
	jnot g02275(.din(w_n2368_0[0]),.dout(n2489),.clk(gclk));
	jnot g02276(.din(w_n2361_0[0]),.dout(n2490),.clk(gclk));
	jnot g02277(.din(w_n2350_0[0]),.dout(n2491),.clk(gclk));
	jnot g02278(.din(w_n2258_0[0]),.dout(n2492),.clk(gclk));
	jnot g02279(.din(w_n2255_0[0]),.dout(n2493),.clk(gclk));
	jor g02280(.dina(w_n2345_57[1]),.dinb(w_n2110_0[2]),.dout(n2494),.clk(gclk));
	jand g02281(.dina(n2494),.dinb(n2493),.dout(n2495),.clk(gclk));
	jand g02282(.dina(n2495),.dinb(w_n2108_59[1]),.dout(n2496),.clk(gclk));
	jor g02283(.dina(w_n2345_57[0]),.dinb(w_a92_0[0]),.dout(n2497),.clk(gclk));
	jand g02284(.dina(n2497),.dinb(w_a93_0[0]),.dout(n2498),.clk(gclk));
	jor g02285(.dina(w_n2352_0[0]),.dinb(n2498),.dout(n2499),.clk(gclk));
	jor g02286(.dina(w_n2499_0[1]),.dinb(n2496),.dout(n2500),.clk(gclk));
	jand g02287(.dina(n2500),.dinb(n2492),.dout(n2501),.clk(gclk));
	jand g02288(.dina(n2501),.dinb(w_n1912_57[2]),.dout(n2502),.clk(gclk));
	jor g02289(.dina(w_n2357_0[0]),.dinb(n2502),.dout(n2503),.clk(gclk));
	jand g02290(.dina(n2503),.dinb(n2491),.dout(n2504),.clk(gclk));
	jand g02291(.dina(n2504),.dinb(w_n1699_60[0]),.dout(n2505),.clk(gclk));
	jnot g02292(.din(w_n2365_0[0]),.dout(n2506),.clk(gclk));
	jor g02293(.dina(w_n2506_0[1]),.dinb(n2505),.dout(n2507),.clk(gclk));
	jand g02294(.dina(n2507),.dinb(n2490),.dout(n2508),.clk(gclk));
	jand g02295(.dina(n2508),.dinb(w_n1516_58[1]),.dout(n2509),.clk(gclk));
	jor g02296(.dina(w_n2372_0[0]),.dinb(n2509),.dout(n2510),.clk(gclk));
	jand g02297(.dina(n2510),.dinb(n2489),.dout(n2511),.clk(gclk));
	jand g02298(.dina(n2511),.dinb(w_n1332_60[0]),.dout(n2512),.clk(gclk));
	jnot g02299(.din(w_n2380_0[0]),.dout(n2513),.clk(gclk));
	jor g02300(.dina(w_n2513_0[1]),.dinb(n2512),.dout(n2514),.clk(gclk));
	jand g02301(.dina(n2514),.dinb(n2488),.dout(n2515),.clk(gclk));
	jand g02302(.dina(n2515),.dinb(w_n1173_59[0]),.dout(n2516),.clk(gclk));
	jor g02303(.dina(w_n2387_0[0]),.dinb(n2516),.dout(n2517),.clk(gclk));
	jand g02304(.dina(n2517),.dinb(n2487),.dout(n2518),.clk(gclk));
	jand g02305(.dina(n2518),.dinb(w_n1008_61[0]),.dout(n2519),.clk(gclk));
	jnot g02306(.din(w_n2395_0[0]),.dout(n2520),.clk(gclk));
	jor g02307(.dina(w_n2520_0[1]),.dinb(n2519),.dout(n2521),.clk(gclk));
	jand g02308(.dina(n2521),.dinb(n2486),.dout(n2522),.clk(gclk));
	jand g02309(.dina(n2522),.dinb(w_n884_60[0]),.dout(n2523),.clk(gclk));
	jor g02310(.dina(w_n2402_0[0]),.dinb(n2523),.dout(n2524),.clk(gclk));
	jand g02311(.dina(n2524),.dinb(n2485),.dout(n2525),.clk(gclk));
	jand g02312(.dina(n2525),.dinb(w_n743_61[0]),.dout(n2526),.clk(gclk));
	jor g02313(.dina(w_n2410_0[0]),.dinb(n2526),.dout(n2527),.clk(gclk));
	jand g02314(.dina(n2527),.dinb(n2484),.dout(n2528),.clk(gclk));
	jand g02315(.dina(n2528),.dinb(w_n635_61[0]),.dout(n2529),.clk(gclk));
	jnot g02316(.din(w_n2418_0[0]),.dout(n2530),.clk(gclk));
	jor g02317(.dina(w_n2530_0[1]),.dinb(n2529),.dout(n2531),.clk(gclk));
	jand g02318(.dina(n2531),.dinb(n2483),.dout(n2532),.clk(gclk));
	jand g02319(.dina(n2532),.dinb(w_n515_62[0]),.dout(n2533),.clk(gclk));
	jnot g02320(.din(w_n2425_0[0]),.dout(n2534),.clk(gclk));
	jor g02321(.dina(w_n2534_0[1]),.dinb(n2533),.dout(n2535),.clk(gclk));
	jand g02322(.dina(n2535),.dinb(n2482),.dout(n2536),.clk(gclk));
	jand g02323(.dina(n2536),.dinb(w_n443_62[0]),.dout(n2537),.clk(gclk));
	jor g02324(.dina(w_n2432_0[0]),.dinb(n2537),.dout(n2538),.clk(gclk));
	jand g02325(.dina(n2538),.dinb(n2481),.dout(n2539),.clk(gclk));
	jand g02326(.dina(n2539),.dinb(w_n352_62[1]),.dout(n2540),.clk(gclk));
	jnot g02327(.din(w_n2440_0[0]),.dout(n2541),.clk(gclk));
	jor g02328(.dina(w_n2541_0[1]),.dinb(n2540),.dout(n2542),.clk(gclk));
	jand g02329(.dina(n2542),.dinb(n2480),.dout(n2543),.clk(gclk));
	jand g02330(.dina(n2543),.dinb(w_n294_62[2]),.dout(n2544),.clk(gclk));
	jnot g02331(.din(w_n2447_0[0]),.dout(n2545),.clk(gclk));
	jor g02332(.dina(w_n2545_0[1]),.dinb(n2544),.dout(n2546),.clk(gclk));
	jand g02333(.dina(n2546),.dinb(n2479),.dout(n2547),.clk(gclk));
	jand g02334(.dina(n2547),.dinb(w_n239_62[2]),.dout(n2548),.clk(gclk));
	jnot g02335(.din(w_n2454_0[0]),.dout(n2549),.clk(gclk));
	jor g02336(.dina(w_n2549_0[1]),.dinb(n2548),.dout(n2550),.clk(gclk));
	jand g02337(.dina(n2550),.dinb(n2478),.dout(n2551),.clk(gclk));
	jand g02338(.dina(n2551),.dinb(w_n221_63[0]),.dout(n2552),.clk(gclk));
	jor g02339(.dina(w_n2461_0[1]),.dinb(n2552),.dout(n2553),.clk(gclk));
	jand g02340(.dina(n2553),.dinb(n2477),.dout(n2554),.clk(gclk));
	jor g02341(.dina(w_n2467_0[0]),.dinb(w_n2554_0[1]),.dout(n2555),.clk(gclk));
	jor g02342(.dina(w_n2555_0[1]),.dinb(w_n2236_0[0]),.dout(n2556),.clk(gclk));
	jor g02343(.dina(n2556),.dinb(w_n2476_0[1]),.dout(n2557),.clk(gclk));
	jand g02344(.dina(n2557),.dinb(w_n218_26[0]),.dout(n2558),.clk(gclk));
	jand g02345(.dina(w_n2345_56[2]),.dinb(w_n2235_0[1]),.dout(n2559),.clk(gclk));
	jor g02346(.dina(w_n2559_0[1]),.dinb(w_n2558_0[1]),.dout(n2560),.clk(gclk));
	jor g02347(.dina(n2560),.dinb(w_n2475_0[1]),.dout(n2561),.clk(gclk));
	jor g02348(.dina(w_n2561_0[1]),.dinb(w_n2470_0[2]),.dout(asqrt_fa_46),.clk(gclk));
	jnot g02349(.din(w_n2475_0[0]),.dout(n2563),.clk(gclk));
	jnot g02350(.din(w_n2476_0[0]),.dout(n2564),.clk(gclk));
	jand g02351(.dina(w_n2468_0[0]),.dinb(w_n2464_0[0]),.dout(n2565),.clk(gclk));
	jand g02352(.dina(w_n2565_0[1]),.dinb(w_n2263_0[1]),.dout(n2566),.clk(gclk));
	jand g02353(.dina(n2566),.dinb(n2564),.dout(n2567),.clk(gclk));
	jor g02354(.dina(n2567),.dinb(w_asqrt63_47[2]),.dout(n2568),.clk(gclk));
	jnot g02355(.din(w_n2559_0[0]),.dout(n2569),.clk(gclk));
	jand g02356(.dina(n2569),.dinb(n2568),.dout(n2570),.clk(gclk));
	jand g02357(.dina(n2570),.dinb(n2563),.dout(n2571),.clk(gclk));
	jand g02358(.dina(w_n2571_0[1]),.dinb(w_n2469_1[0]),.dout(n2572),.clk(gclk));
	jxor g02359(.dina(w_n2456_0[0]),.dinb(w_n221_62[2]),.dout(n2573),.clk(gclk));
	jor g02360(.dina(n2573),.dinb(w_n2572_63[1]),.dout(n2574),.clk(gclk));
	jxor g02361(.dina(n2574),.dinb(w_n2461_0[0]),.dout(n2575),.clk(gclk));
	jnot g02362(.din(w_n2575_0[1]),.dout(n2576),.clk(gclk));
	jor g02363(.dina(w_n2572_63[0]),.dinb(w_n2252_1[0]),.dout(n2577),.clk(gclk));
	jnot g02364(.din(w_a88_0[2]),.dout(n2578),.clk(gclk));
	jnot g02365(.din(w_a89_0[1]),.dout(n2579),.clk(gclk));
	jand g02366(.dina(w_n2579_0[1]),.dinb(w_n2578_1[2]),.dout(n2580),.clk(gclk));
	jand g02367(.dina(w_n2580_0[2]),.dinb(w_n2252_0[2]),.dout(n2581),.clk(gclk));
	jnot g02368(.din(w_n2581_0[1]),.dout(n2582),.clk(gclk));
	jand g02369(.dina(n2582),.dinb(n2577),.dout(n2583),.clk(gclk));
	jor g02370(.dina(w_n2583_0[2]),.dinb(w_n2345_56[1]),.dout(n2584),.clk(gclk));
	jand g02371(.dina(w_n2583_0[1]),.dinb(w_n2345_56[0]),.dout(n2585),.clk(gclk));
	jor g02372(.dina(w_n2572_62[2]),.dinb(w_a90_1[0]),.dout(n2586),.clk(gclk));
	jand g02373(.dina(n2586),.dinb(w_a91_0[0]),.dout(n2587),.clk(gclk));
	jand g02374(.dina(w_asqrt45_34),.dinb(w_n2254_0[1]),.dout(n2588),.clk(gclk));
	jor g02375(.dina(n2588),.dinb(n2587),.dout(n2589),.clk(gclk));
	jor g02376(.dina(n2589),.dinb(n2585),.dout(n2590),.clk(gclk));
	jand g02377(.dina(n2590),.dinb(w_n2584_0[1]),.dout(n2591),.clk(gclk));
	jor g02378(.dina(w_n2591_0[2]),.dinb(w_n2108_59[0]),.dout(n2592),.clk(gclk));
	jand g02379(.dina(w_n2591_0[1]),.dinb(w_n2108_58[2]),.dout(n2593),.clk(gclk));
	jnot g02380(.din(w_n2254_0[0]),.dout(n2594),.clk(gclk));
	jor g02381(.dina(w_n2572_62[1]),.dinb(n2594),.dout(n2595),.clk(gclk));
	jor g02382(.dina(w_n2470_0[1]),.dinb(w_n2345_55[2]),.dout(n2596),.clk(gclk));
	jor g02383(.dina(n2596),.dinb(w_n2474_0[0]),.dout(n2597),.clk(gclk));
	jor g02384(.dina(n2597),.dinb(w_n2558_0[0]),.dout(n2598),.clk(gclk));
	jand g02385(.dina(n2598),.dinb(w_n2595_0[1]),.dout(n2599),.clk(gclk));
	jxor g02386(.dina(n2599),.dinb(w_n2110_0[1]),.dout(n2600),.clk(gclk));
	jor g02387(.dina(w_n2600_0[2]),.dinb(n2593),.dout(n2601),.clk(gclk));
	jand g02388(.dina(n2601),.dinb(w_n2592_0[1]),.dout(n2602),.clk(gclk));
	jor g02389(.dina(w_n2602_0[2]),.dinb(w_n1912_57[1]),.dout(n2603),.clk(gclk));
	jand g02390(.dina(w_n2602_0[1]),.dinb(w_n1912_57[0]),.dout(n2604),.clk(gclk));
	jxor g02391(.dina(w_n2257_0[0]),.dinb(w_n2108_58[1]),.dout(n2605),.clk(gclk));
	jor g02392(.dina(n2605),.dinb(w_n2572_62[0]),.dout(n2606),.clk(gclk));
	jxor g02393(.dina(n2606),.dinb(w_n2499_0[0]),.dout(n2607),.clk(gclk));
	jnot g02394(.din(w_n2607_0[2]),.dout(n2608),.clk(gclk));
	jor g02395(.dina(n2608),.dinb(n2604),.dout(n2609),.clk(gclk));
	jand g02396(.dina(n2609),.dinb(w_n2603_0[1]),.dout(n2610),.clk(gclk));
	jor g02397(.dina(w_n2610_0[2]),.dinb(w_n1699_59[2]),.dout(n2611),.clk(gclk));
	jand g02398(.dina(w_n2610_0[1]),.dinb(w_n1699_59[1]),.dout(n2612),.clk(gclk));
	jxor g02399(.dina(w_n2349_0[0]),.dinb(w_n1912_56[2]),.dout(n2613),.clk(gclk));
	jor g02400(.dina(n2613),.dinb(w_n2572_61[2]),.dout(n2614),.clk(gclk));
	jxor g02401(.dina(n2614),.dinb(w_n2358_0[0]),.dout(n2615),.clk(gclk));
	jor g02402(.dina(w_n2615_0[2]),.dinb(n2612),.dout(n2616),.clk(gclk));
	jand g02403(.dina(n2616),.dinb(w_n2611_0[1]),.dout(n2617),.clk(gclk));
	jor g02404(.dina(w_n2617_0[2]),.dinb(w_n1516_58[0]),.dout(n2618),.clk(gclk));
	jand g02405(.dina(w_n2617_0[1]),.dinb(w_n1516_57[2]),.dout(n2619),.clk(gclk));
	jxor g02406(.dina(w_n2360_0[0]),.dinb(w_n1699_59[0]),.dout(n2620),.clk(gclk));
	jor g02407(.dina(n2620),.dinb(w_n2572_61[1]),.dout(n2621),.clk(gclk));
	jxor g02408(.dina(n2621),.dinb(w_n2506_0[0]),.dout(n2622),.clk(gclk));
	jnot g02409(.din(w_n2622_0[2]),.dout(n2623),.clk(gclk));
	jor g02410(.dina(n2623),.dinb(n2619),.dout(n2624),.clk(gclk));
	jand g02411(.dina(n2624),.dinb(w_n2618_0[1]),.dout(n2625),.clk(gclk));
	jor g02412(.dina(w_n2625_0[2]),.dinb(w_n1332_59[2]),.dout(n2626),.clk(gclk));
	jand g02413(.dina(w_n2625_0[1]),.dinb(w_n1332_59[1]),.dout(n2627),.clk(gclk));
	jxor g02414(.dina(w_n2367_0[0]),.dinb(w_n1516_57[1]),.dout(n2628),.clk(gclk));
	jor g02415(.dina(n2628),.dinb(w_n2572_61[0]),.dout(n2629),.clk(gclk));
	jxor g02416(.dina(n2629),.dinb(w_n2373_0[0]),.dout(n2630),.clk(gclk));
	jor g02417(.dina(w_n2630_0[2]),.dinb(n2627),.dout(n2631),.clk(gclk));
	jand g02418(.dina(n2631),.dinb(w_n2626_0[1]),.dout(n2632),.clk(gclk));
	jor g02419(.dina(w_n2632_0[2]),.dinb(w_n1173_58[2]),.dout(n2633),.clk(gclk));
	jand g02420(.dina(w_n2632_0[1]),.dinb(w_n1173_58[1]),.dout(n2634),.clk(gclk));
	jxor g02421(.dina(w_n2375_0[0]),.dinb(w_n1332_59[0]),.dout(n2635),.clk(gclk));
	jor g02422(.dina(n2635),.dinb(w_n2572_60[2]),.dout(n2636),.clk(gclk));
	jxor g02423(.dina(n2636),.dinb(w_n2513_0[0]),.dout(n2637),.clk(gclk));
	jnot g02424(.din(w_n2637_0[2]),.dout(n2638),.clk(gclk));
	jor g02425(.dina(n2638),.dinb(n2634),.dout(n2639),.clk(gclk));
	jand g02426(.dina(n2639),.dinb(w_n2633_0[1]),.dout(n2640),.clk(gclk));
	jor g02427(.dina(w_n2640_0[2]),.dinb(w_n1008_60[2]),.dout(n2641),.clk(gclk));
	jand g02428(.dina(w_n2640_0[1]),.dinb(w_n1008_60[1]),.dout(n2642),.clk(gclk));
	jxor g02429(.dina(w_n2382_0[0]),.dinb(w_n1173_58[0]),.dout(n2643),.clk(gclk));
	jor g02430(.dina(n2643),.dinb(w_n2572_60[1]),.dout(n2644),.clk(gclk));
	jxor g02431(.dina(n2644),.dinb(w_n2388_0[0]),.dout(n2645),.clk(gclk));
	jor g02432(.dina(w_n2645_0[2]),.dinb(n2642),.dout(n2646),.clk(gclk));
	jand g02433(.dina(n2646),.dinb(w_n2641_0[1]),.dout(n2647),.clk(gclk));
	jor g02434(.dina(w_n2647_0[2]),.dinb(w_n884_59[2]),.dout(n2648),.clk(gclk));
	jand g02435(.dina(w_n2647_0[1]),.dinb(w_n884_59[1]),.dout(n2649),.clk(gclk));
	jxor g02436(.dina(w_n2390_0[0]),.dinb(w_n1008_60[0]),.dout(n2650),.clk(gclk));
	jor g02437(.dina(n2650),.dinb(w_n2572_60[0]),.dout(n2651),.clk(gclk));
	jxor g02438(.dina(n2651),.dinb(w_n2520_0[0]),.dout(n2652),.clk(gclk));
	jnot g02439(.din(w_n2652_0[2]),.dout(n2653),.clk(gclk));
	jor g02440(.dina(n2653),.dinb(n2649),.dout(n2654),.clk(gclk));
	jand g02441(.dina(n2654),.dinb(w_n2648_0[1]),.dout(n2655),.clk(gclk));
	jor g02442(.dina(w_n2655_0[2]),.dinb(w_n743_60[2]),.dout(n2656),.clk(gclk));
	jand g02443(.dina(w_n2655_0[1]),.dinb(w_n743_60[1]),.dout(n2657),.clk(gclk));
	jxor g02444(.dina(w_n2397_0[0]),.dinb(w_n884_59[0]),.dout(n2658),.clk(gclk));
	jor g02445(.dina(n2658),.dinb(w_n2572_59[2]),.dout(n2659),.clk(gclk));
	jxor g02446(.dina(n2659),.dinb(w_n2403_0[0]),.dout(n2660),.clk(gclk));
	jor g02447(.dina(w_n2660_0[2]),.dinb(n2657),.dout(n2661),.clk(gclk));
	jand g02448(.dina(n2661),.dinb(w_n2656_0[1]),.dout(n2662),.clk(gclk));
	jor g02449(.dina(w_n2662_0[2]),.dinb(w_n635_60[2]),.dout(n2663),.clk(gclk));
	jand g02450(.dina(w_n2662_0[1]),.dinb(w_n635_60[1]),.dout(n2664),.clk(gclk));
	jxor g02451(.dina(w_n2405_0[0]),.dinb(w_n743_60[0]),.dout(n2665),.clk(gclk));
	jor g02452(.dina(n2665),.dinb(w_n2572_59[1]),.dout(n2666),.clk(gclk));
	jxor g02453(.dina(n2666),.dinb(w_n2411_0[0]),.dout(n2667),.clk(gclk));
	jor g02454(.dina(w_n2667_0[2]),.dinb(n2664),.dout(n2668),.clk(gclk));
	jand g02455(.dina(n2668),.dinb(w_n2663_0[1]),.dout(n2669),.clk(gclk));
	jor g02456(.dina(w_n2669_0[2]),.dinb(w_n515_61[2]),.dout(n2670),.clk(gclk));
	jand g02457(.dina(w_n2669_0[1]),.dinb(w_n515_61[1]),.dout(n2671),.clk(gclk));
	jxor g02458(.dina(w_n2413_0[0]),.dinb(w_n635_60[0]),.dout(n2672),.clk(gclk));
	jor g02459(.dina(n2672),.dinb(w_n2572_59[0]),.dout(n2673),.clk(gclk));
	jxor g02460(.dina(n2673),.dinb(w_n2530_0[0]),.dout(n2674),.clk(gclk));
	jnot g02461(.din(w_n2674_0[2]),.dout(n2675),.clk(gclk));
	jor g02462(.dina(n2675),.dinb(n2671),.dout(n2676),.clk(gclk));
	jand g02463(.dina(n2676),.dinb(w_n2670_0[1]),.dout(n2677),.clk(gclk));
	jor g02464(.dina(w_n2677_0[2]),.dinb(w_n443_61[2]),.dout(n2678),.clk(gclk));
	jand g02465(.dina(w_n2677_0[1]),.dinb(w_n443_61[1]),.dout(n2679),.clk(gclk));
	jxor g02466(.dina(w_n2420_0[0]),.dinb(w_n515_61[0]),.dout(n2680),.clk(gclk));
	jor g02467(.dina(n2680),.dinb(w_n2572_58[2]),.dout(n2681),.clk(gclk));
	jxor g02468(.dina(n2681),.dinb(w_n2534_0[0]),.dout(n2682),.clk(gclk));
	jnot g02469(.din(w_n2682_0[2]),.dout(n2683),.clk(gclk));
	jor g02470(.dina(n2683),.dinb(n2679),.dout(n2684),.clk(gclk));
	jand g02471(.dina(n2684),.dinb(w_n2678_0[1]),.dout(n2685),.clk(gclk));
	jor g02472(.dina(w_n2685_0[2]),.dinb(w_n352_62[0]),.dout(n2686),.clk(gclk));
	jand g02473(.dina(w_n2685_0[1]),.dinb(w_n352_61[2]),.dout(n2687),.clk(gclk));
	jxor g02474(.dina(w_n2427_0[0]),.dinb(w_n443_61[0]),.dout(n2688),.clk(gclk));
	jor g02475(.dina(n2688),.dinb(w_n2572_58[1]),.dout(n2689),.clk(gclk));
	jxor g02476(.dina(n2689),.dinb(w_n2433_0[0]),.dout(n2690),.clk(gclk));
	jor g02477(.dina(w_n2690_0[2]),.dinb(n2687),.dout(n2691),.clk(gclk));
	jand g02478(.dina(n2691),.dinb(w_n2686_0[1]),.dout(n2692),.clk(gclk));
	jor g02479(.dina(w_n2692_0[2]),.dinb(w_n294_62[1]),.dout(n2693),.clk(gclk));
	jand g02480(.dina(w_n2692_0[1]),.dinb(w_n294_62[0]),.dout(n2694),.clk(gclk));
	jxor g02481(.dina(w_n2435_0[0]),.dinb(w_n352_61[1]),.dout(n2695),.clk(gclk));
	jor g02482(.dina(n2695),.dinb(w_n2572_58[0]),.dout(n2696),.clk(gclk));
	jxor g02483(.dina(n2696),.dinb(w_n2541_0[0]),.dout(n2697),.clk(gclk));
	jnot g02484(.din(w_n2697_0[2]),.dout(n2698),.clk(gclk));
	jor g02485(.dina(n2698),.dinb(n2694),.dout(n2699),.clk(gclk));
	jand g02486(.dina(n2699),.dinb(w_n2693_0[1]),.dout(n2700),.clk(gclk));
	jor g02487(.dina(w_n2700_0[2]),.dinb(w_n239_62[1]),.dout(n2701),.clk(gclk));
	jand g02488(.dina(w_n2700_0[1]),.dinb(w_n239_62[0]),.dout(n2702),.clk(gclk));
	jxor g02489(.dina(w_n2442_0[0]),.dinb(w_n294_61[2]),.dout(n2703),.clk(gclk));
	jor g02490(.dina(n2703),.dinb(w_n2572_57[2]),.dout(n2704),.clk(gclk));
	jxor g02491(.dina(n2704),.dinb(w_n2545_0[0]),.dout(n2705),.clk(gclk));
	jnot g02492(.din(w_n2705_0[2]),.dout(n2706),.clk(gclk));
	jor g02493(.dina(n2706),.dinb(n2702),.dout(n2707),.clk(gclk));
	jand g02494(.dina(n2707),.dinb(w_n2701_0[1]),.dout(n2708),.clk(gclk));
	jor g02495(.dina(w_n2708_0[2]),.dinb(w_n221_62[1]),.dout(n2709),.clk(gclk));
	jand g02496(.dina(w_n2708_0[1]),.dinb(w_n221_62[0]),.dout(n2710),.clk(gclk));
	jxor g02497(.dina(w_n2449_0[0]),.dinb(w_n239_61[2]),.dout(n2711),.clk(gclk));
	jor g02498(.dina(n2711),.dinb(w_n2572_57[1]),.dout(n2712),.clk(gclk));
	jxor g02499(.dina(n2712),.dinb(w_n2549_0[0]),.dout(n2713),.clk(gclk));
	jnot g02500(.din(w_n2713_0[1]),.dout(n2714),.clk(gclk));
	jor g02501(.dina(w_n2714_0[1]),.dinb(n2710),.dout(n2715),.clk(gclk));
	jand g02502(.dina(n2715),.dinb(w_n2709_0[1]),.dout(n2716),.clk(gclk));
	jand g02503(.dina(w_n2716_0[2]),.dinb(w_n2576_0[2]),.dout(n2717),.clk(gclk));
	jand g02504(.dina(w_n2561_0[0]),.dinb(w_n2565_0[0]),.dout(n2719),.clk(gclk));
	jor g02505(.dina(w_n2716_0[1]),.dinb(w_n2576_0[1]),.dout(n2720),.clk(gclk));
	jor g02506(.dina(w_n2720_0[1]),.dinb(w_n2470_0[0]),.dout(n2721),.clk(gclk));
	jor g02507(.dina(n2721),.dinb(w_n2719_0[1]),.dout(n2722),.clk(gclk));
	jand g02508(.dina(n2722),.dinb(w_n218_25[2]),.dout(n2723),.clk(gclk));
	jand g02509(.dina(w_n2571_0[0]),.dinb(w_n2554_0[0]),.dout(n2724),.clk(gclk));
	jand g02510(.dina(w_n2555_0[0]),.dinb(w_asqrt63_47[1]),.dout(n2725),.clk(gclk));
	jand g02511(.dina(n2725),.dinb(w_n2469_0[2]),.dout(n2726),.clk(gclk));
	jnot g02512(.din(n2726),.dout(n2727),.clk(gclk));
	jor g02513(.dina(w_n2727_0[1]),.dinb(n2724),.dout(n2728),.clk(gclk));
	jnot g02514(.din(w_n2728_0[1]),.dout(n2729),.clk(gclk));
	jor g02515(.dina(n2729),.dinb(n2723),.dout(n2730),.clk(gclk));
	jor g02516(.dina(w_n2730_0[1]),.dinb(w_n2717_0[2]),.dout(asqrt_fa_45),.clk(gclk));
	jand g02517(.dina(w_asqrt44_41),.dinb(w_a88_0[1]),.dout(n2733),.clk(gclk));
	jnot g02518(.din(w_a86_1[1]),.dout(n2734),.clk(gclk));
	jnot g02519(.din(w_a87_0[1]),.dout(n2735),.clk(gclk));
	jand g02520(.dina(w_n2735_0[1]),.dinb(w_n2734_1[1]),.dout(n2736),.clk(gclk));
	jand g02521(.dina(w_n2736_0[2]),.dinb(w_n2578_1[1]),.dout(n2737),.clk(gclk));
	jor g02522(.dina(w_n2737_0[1]),.dinb(n2733),.dout(n2738),.clk(gclk));
	jand g02523(.dina(w_n2738_0[2]),.dinb(w_asqrt45_33[2]),.dout(n2739),.clk(gclk));
	jor g02524(.dina(w_n2738_0[1]),.dinb(w_asqrt45_33[1]),.dout(n2740),.clk(gclk));
	jand g02525(.dina(w_asqrt44_40[2]),.dinb(w_n2578_1[0]),.dout(n2741),.clk(gclk));
	jor g02526(.dina(n2741),.dinb(w_n2579_0[0]),.dout(n2742),.clk(gclk));
	jnot g02527(.din(w_n2580_0[1]),.dout(n2743),.clk(gclk));
	jnot g02528(.din(w_n2717_0[1]),.dout(n2744),.clk(gclk));
	jnot g02529(.din(w_n2719_0[0]),.dout(n2746),.clk(gclk));
	jnot g02530(.din(w_n2709_0[0]),.dout(n2747),.clk(gclk));
	jnot g02531(.din(w_n2701_0[0]),.dout(n2748),.clk(gclk));
	jnot g02532(.din(w_n2693_0[0]),.dout(n2749),.clk(gclk));
	jnot g02533(.din(w_n2686_0[0]),.dout(n2750),.clk(gclk));
	jnot g02534(.din(w_n2678_0[0]),.dout(n2751),.clk(gclk));
	jnot g02535(.din(w_n2670_0[0]),.dout(n2752),.clk(gclk));
	jnot g02536(.din(w_n2663_0[0]),.dout(n2753),.clk(gclk));
	jnot g02537(.din(w_n2656_0[0]),.dout(n2754),.clk(gclk));
	jnot g02538(.din(w_n2648_0[0]),.dout(n2755),.clk(gclk));
	jnot g02539(.din(w_n2641_0[0]),.dout(n2756),.clk(gclk));
	jnot g02540(.din(w_n2633_0[0]),.dout(n2757),.clk(gclk));
	jnot g02541(.din(w_n2626_0[0]),.dout(n2758),.clk(gclk));
	jnot g02542(.din(w_n2618_0[0]),.dout(n2759),.clk(gclk));
	jnot g02543(.din(w_n2611_0[0]),.dout(n2760),.clk(gclk));
	jnot g02544(.din(w_n2603_0[0]),.dout(n2761),.clk(gclk));
	jnot g02545(.din(w_n2592_0[0]),.dout(n2762),.clk(gclk));
	jnot g02546(.din(w_n2584_0[0]),.dout(n2763),.clk(gclk));
	jand g02547(.dina(w_asqrt45_33[0]),.dinb(w_a90_0[2]),.dout(n2764),.clk(gclk));
	jor g02548(.dina(w_n2581_0[0]),.dinb(n2764),.dout(n2765),.clk(gclk));
	jor g02549(.dina(n2765),.dinb(w_asqrt46_35[1]),.dout(n2766),.clk(gclk));
	jand g02550(.dina(w_asqrt45_32[2]),.dinb(w_n2252_0[1]),.dout(n2767),.clk(gclk));
	jor g02551(.dina(n2767),.dinb(w_n2253_0[0]),.dout(n2768),.clk(gclk));
	jand g02552(.dina(w_n2595_0[0]),.dinb(n2768),.dout(n2769),.clk(gclk));
	jand g02553(.dina(w_n2769_0[1]),.dinb(n2766),.dout(n2770),.clk(gclk));
	jor g02554(.dina(n2770),.dinb(n2763),.dout(n2771),.clk(gclk));
	jor g02555(.dina(n2771),.dinb(w_asqrt47_33[2]),.dout(n2772),.clk(gclk));
	jnot g02556(.din(w_n2600_0[1]),.dout(n2773),.clk(gclk));
	jand g02557(.dina(n2773),.dinb(n2772),.dout(n2774),.clk(gclk));
	jor g02558(.dina(n2774),.dinb(n2762),.dout(n2775),.clk(gclk));
	jor g02559(.dina(n2775),.dinb(w_asqrt48_35[2]),.dout(n2776),.clk(gclk));
	jand g02560(.dina(w_n2607_0[1]),.dinb(n2776),.dout(n2777),.clk(gclk));
	jor g02561(.dina(n2777),.dinb(n2761),.dout(n2778),.clk(gclk));
	jor g02562(.dina(n2778),.dinb(w_asqrt49_34[0]),.dout(n2779),.clk(gclk));
	jnot g02563(.din(w_n2615_0[1]),.dout(n2780),.clk(gclk));
	jand g02564(.dina(n2780),.dinb(n2779),.dout(n2781),.clk(gclk));
	jor g02565(.dina(n2781),.dinb(n2760),.dout(n2782),.clk(gclk));
	jor g02566(.dina(n2782),.dinb(w_asqrt50_36[0]),.dout(n2783),.clk(gclk));
	jand g02567(.dina(w_n2622_0[1]),.dinb(n2783),.dout(n2784),.clk(gclk));
	jor g02568(.dina(n2784),.dinb(n2759),.dout(n2785),.clk(gclk));
	jor g02569(.dina(n2785),.dinb(w_asqrt51_34[1]),.dout(n2786),.clk(gclk));
	jnot g02570(.din(w_n2630_0[1]),.dout(n2787),.clk(gclk));
	jand g02571(.dina(n2787),.dinb(n2786),.dout(n2788),.clk(gclk));
	jor g02572(.dina(n2788),.dinb(n2758),.dout(n2789),.clk(gclk));
	jor g02573(.dina(n2789),.dinb(w_asqrt52_36[0]),.dout(n2790),.clk(gclk));
	jand g02574(.dina(w_n2637_0[1]),.dinb(n2790),.dout(n2791),.clk(gclk));
	jor g02575(.dina(n2791),.dinb(n2757),.dout(n2792),.clk(gclk));
	jor g02576(.dina(n2792),.dinb(w_asqrt53_35[0]),.dout(n2793),.clk(gclk));
	jnot g02577(.din(w_n2645_0[1]),.dout(n2794),.clk(gclk));
	jand g02578(.dina(n2794),.dinb(n2793),.dout(n2795),.clk(gclk));
	jor g02579(.dina(n2795),.dinb(n2756),.dout(n2796),.clk(gclk));
	jor g02580(.dina(n2796),.dinb(w_asqrt54_36[0]),.dout(n2797),.clk(gclk));
	jand g02581(.dina(w_n2652_0[1]),.dinb(n2797),.dout(n2798),.clk(gclk));
	jor g02582(.dina(n2798),.dinb(n2755),.dout(n2799),.clk(gclk));
	jor g02583(.dina(n2799),.dinb(w_asqrt55_35[1]),.dout(n2800),.clk(gclk));
	jnot g02584(.din(w_n2660_0[1]),.dout(n2801),.clk(gclk));
	jand g02585(.dina(n2801),.dinb(n2800),.dout(n2802),.clk(gclk));
	jor g02586(.dina(n2802),.dinb(n2754),.dout(n2803),.clk(gclk));
	jor g02587(.dina(n2803),.dinb(w_asqrt56_36[1]),.dout(n2804),.clk(gclk));
	jnot g02588(.din(w_n2667_0[1]),.dout(n2805),.clk(gclk));
	jand g02589(.dina(n2805),.dinb(n2804),.dout(n2806),.clk(gclk));
	jor g02590(.dina(n2806),.dinb(n2753),.dout(n2807),.clk(gclk));
	jor g02591(.dina(n2807),.dinb(w_asqrt57_36[0]),.dout(n2808),.clk(gclk));
	jand g02592(.dina(w_n2674_0[1]),.dinb(n2808),.dout(n2809),.clk(gclk));
	jor g02593(.dina(n2809),.dinb(n2752),.dout(n2810),.clk(gclk));
	jor g02594(.dina(n2810),.dinb(w_asqrt58_36[2]),.dout(n2811),.clk(gclk));
	jand g02595(.dina(w_n2682_0[1]),.dinb(n2811),.dout(n2812),.clk(gclk));
	jor g02596(.dina(n2812),.dinb(n2751),.dout(n2813),.clk(gclk));
	jor g02597(.dina(n2813),.dinb(w_asqrt59_36[1]),.dout(n2814),.clk(gclk));
	jnot g02598(.din(w_n2690_0[1]),.dout(n2815),.clk(gclk));
	jand g02599(.dina(n2815),.dinb(n2814),.dout(n2816),.clk(gclk));
	jor g02600(.dina(n2816),.dinb(n2750),.dout(n2817),.clk(gclk));
	jor g02601(.dina(n2817),.dinb(w_asqrt60_36[2]),.dout(n2818),.clk(gclk));
	jand g02602(.dina(w_n2697_0[1]),.dinb(n2818),.dout(n2819),.clk(gclk));
	jor g02603(.dina(n2819),.dinb(n2749),.dout(n2820),.clk(gclk));
	jor g02604(.dina(n2820),.dinb(w_asqrt61_36[2]),.dout(n2821),.clk(gclk));
	jand g02605(.dina(w_n2705_0[1]),.dinb(n2821),.dout(n2822),.clk(gclk));
	jor g02606(.dina(n2822),.dinb(n2748),.dout(n2823),.clk(gclk));
	jor g02607(.dina(n2823),.dinb(w_asqrt62_36[2]),.dout(n2824),.clk(gclk));
	jand g02608(.dina(w_n2713_0[0]),.dinb(n2824),.dout(n2825),.clk(gclk));
	jor g02609(.dina(n2825),.dinb(n2747),.dout(n2826),.clk(gclk));
	jand g02610(.dina(n2826),.dinb(w_n2575_0[0]),.dout(n2827),.clk(gclk));
	jand g02611(.dina(w_n2827_0[1]),.dinb(w_n2469_0[1]),.dout(n2828),.clk(gclk));
	jand g02612(.dina(n2828),.dinb(n2746),.dout(n2829),.clk(gclk));
	jor g02613(.dina(n2829),.dinb(w_asqrt63_47[0]),.dout(n2830),.clk(gclk));
	jand g02614(.dina(w_n2728_0[0]),.dinb(w_n2830_0[1]),.dout(n2831),.clk(gclk));
	jand g02615(.dina(w_n2831_0[1]),.dinb(w_n2744_1[1]),.dout(n2833),.clk(gclk));
	jor g02616(.dina(w_n2833_55[1]),.dinb(n2743),.dout(n2834),.clk(gclk));
	jand g02617(.dina(n2834),.dinb(n2742),.dout(n2835),.clk(gclk));
	jand g02618(.dina(w_n2835_0[1]),.dinb(n2740),.dout(n2836),.clk(gclk));
	jor g02619(.dina(n2836),.dinb(w_n2739_0[1]),.dout(n2837),.clk(gclk));
	jand g02620(.dina(w_n2837_0[2]),.dinb(w_asqrt46_35[0]),.dout(n2838),.clk(gclk));
	jor g02621(.dina(w_n2837_0[1]),.dinb(w_asqrt46_34[2]),.dout(n2839),.clk(gclk));
	jand g02622(.dina(w_asqrt44_40[1]),.dinb(w_n2580_0[0]),.dout(n2840),.clk(gclk));
	jand g02623(.dina(w_n2744_1[0]),.dinb(w_asqrt45_32[1]),.dout(n2841),.clk(gclk));
	jand g02624(.dina(n2841),.dinb(w_n2727_0[0]),.dout(n2842),.clk(gclk));
	jand g02625(.dina(n2842),.dinb(w_n2830_0[0]),.dout(n2843),.clk(gclk));
	jor g02626(.dina(n2843),.dinb(w_n2840_0[1]),.dout(n2844),.clk(gclk));
	jxor g02627(.dina(n2844),.dinb(w_a90_0[1]),.dout(n2845),.clk(gclk));
	jnot g02628(.din(w_n2845_0[1]),.dout(n2846),.clk(gclk));
	jand g02629(.dina(w_n2846_0[1]),.dinb(n2839),.dout(n2847),.clk(gclk));
	jor g02630(.dina(n2847),.dinb(w_n2838_0[1]),.dout(n2848),.clk(gclk));
	jand g02631(.dina(w_n2848_0[2]),.dinb(w_asqrt47_33[1]),.dout(n2849),.clk(gclk));
	jor g02632(.dina(w_n2848_0[1]),.dinb(w_asqrt47_33[0]),.dout(n2850),.clk(gclk));
	jxor g02633(.dina(w_n2583_0[0]),.dinb(w_n2345_55[1]),.dout(n2851),.clk(gclk));
	jand g02634(.dina(n2851),.dinb(w_asqrt44_40[0]),.dout(n2852),.clk(gclk));
	jxor g02635(.dina(n2852),.dinb(w_n2769_0[0]),.dout(n2853),.clk(gclk));
	jand g02636(.dina(w_n2853_0[1]),.dinb(n2850),.dout(n2854),.clk(gclk));
	jor g02637(.dina(n2854),.dinb(w_n2849_0[1]),.dout(n2855),.clk(gclk));
	jand g02638(.dina(w_n2855_0[2]),.dinb(w_asqrt48_35[1]),.dout(n2856),.clk(gclk));
	jor g02639(.dina(w_n2855_0[1]),.dinb(w_asqrt48_35[0]),.dout(n2857),.clk(gclk));
	jxor g02640(.dina(w_n2591_0[0]),.dinb(w_n2108_58[0]),.dout(n2858),.clk(gclk));
	jand g02641(.dina(n2858),.dinb(w_asqrt44_39[2]),.dout(n2859),.clk(gclk));
	jxor g02642(.dina(n2859),.dinb(w_n2600_0[0]),.dout(n2860),.clk(gclk));
	jnot g02643(.din(w_n2860_0[1]),.dout(n2861),.clk(gclk));
	jand g02644(.dina(w_n2861_0[1]),.dinb(n2857),.dout(n2862),.clk(gclk));
	jor g02645(.dina(n2862),.dinb(w_n2856_0[1]),.dout(n2863),.clk(gclk));
	jand g02646(.dina(w_n2863_0[2]),.dinb(w_asqrt49_33[2]),.dout(n2864),.clk(gclk));
	jor g02647(.dina(w_n2863_0[1]),.dinb(w_asqrt49_33[1]),.dout(n2865),.clk(gclk));
	jxor g02648(.dina(w_n2602_0[0]),.dinb(w_n1912_56[1]),.dout(n2866),.clk(gclk));
	jand g02649(.dina(n2866),.dinb(w_asqrt44_39[1]),.dout(n2867),.clk(gclk));
	jxor g02650(.dina(n2867),.dinb(w_n2607_0[0]),.dout(n2868),.clk(gclk));
	jand g02651(.dina(w_n2868_0[1]),.dinb(n2865),.dout(n2869),.clk(gclk));
	jor g02652(.dina(n2869),.dinb(w_n2864_0[1]),.dout(n2870),.clk(gclk));
	jand g02653(.dina(w_n2870_0[2]),.dinb(w_asqrt50_35[2]),.dout(n2871),.clk(gclk));
	jor g02654(.dina(w_n2870_0[1]),.dinb(w_asqrt50_35[1]),.dout(n2872),.clk(gclk));
	jxor g02655(.dina(w_n2610_0[0]),.dinb(w_n1699_58[2]),.dout(n2873),.clk(gclk));
	jand g02656(.dina(n2873),.dinb(w_asqrt44_39[0]),.dout(n2874),.clk(gclk));
	jxor g02657(.dina(n2874),.dinb(w_n2615_0[0]),.dout(n2875),.clk(gclk));
	jnot g02658(.din(w_n2875_0[1]),.dout(n2876),.clk(gclk));
	jand g02659(.dina(w_n2876_0[1]),.dinb(n2872),.dout(n2877),.clk(gclk));
	jor g02660(.dina(n2877),.dinb(w_n2871_0[1]),.dout(n2878),.clk(gclk));
	jand g02661(.dina(w_n2878_0[2]),.dinb(w_asqrt51_34[0]),.dout(n2879),.clk(gclk));
	jor g02662(.dina(w_n2878_0[1]),.dinb(w_asqrt51_33[2]),.dout(n2880),.clk(gclk));
	jxor g02663(.dina(w_n2617_0[0]),.dinb(w_n1516_57[0]),.dout(n2881),.clk(gclk));
	jand g02664(.dina(n2881),.dinb(w_asqrt44_38[2]),.dout(n2882),.clk(gclk));
	jxor g02665(.dina(n2882),.dinb(w_n2622_0[0]),.dout(n2883),.clk(gclk));
	jand g02666(.dina(w_n2883_0[1]),.dinb(n2880),.dout(n2884),.clk(gclk));
	jor g02667(.dina(n2884),.dinb(w_n2879_0[1]),.dout(n2885),.clk(gclk));
	jand g02668(.dina(w_n2885_0[2]),.dinb(w_asqrt52_35[2]),.dout(n2886),.clk(gclk));
	jor g02669(.dina(w_n2885_0[1]),.dinb(w_asqrt52_35[1]),.dout(n2887),.clk(gclk));
	jxor g02670(.dina(w_n2625_0[0]),.dinb(w_n1332_58[2]),.dout(n2888),.clk(gclk));
	jand g02671(.dina(n2888),.dinb(w_asqrt44_38[1]),.dout(n2889),.clk(gclk));
	jxor g02672(.dina(n2889),.dinb(w_n2630_0[0]),.dout(n2890),.clk(gclk));
	jnot g02673(.din(w_n2890_0[1]),.dout(n2891),.clk(gclk));
	jand g02674(.dina(w_n2891_0[1]),.dinb(n2887),.dout(n2892),.clk(gclk));
	jor g02675(.dina(n2892),.dinb(w_n2886_0[1]),.dout(n2893),.clk(gclk));
	jand g02676(.dina(w_n2893_0[2]),.dinb(w_asqrt53_34[2]),.dout(n2894),.clk(gclk));
	jor g02677(.dina(w_n2893_0[1]),.dinb(w_asqrt53_34[1]),.dout(n2895),.clk(gclk));
	jxor g02678(.dina(w_n2632_0[0]),.dinb(w_n1173_57[2]),.dout(n2896),.clk(gclk));
	jand g02679(.dina(n2896),.dinb(w_asqrt44_38[0]),.dout(n2897),.clk(gclk));
	jxor g02680(.dina(n2897),.dinb(w_n2637_0[0]),.dout(n2898),.clk(gclk));
	jand g02681(.dina(w_n2898_0[1]),.dinb(n2895),.dout(n2899),.clk(gclk));
	jor g02682(.dina(n2899),.dinb(w_n2894_0[1]),.dout(n2900),.clk(gclk));
	jand g02683(.dina(w_n2900_0[2]),.dinb(w_asqrt54_35[2]),.dout(n2901),.clk(gclk));
	jor g02684(.dina(w_n2900_0[1]),.dinb(w_asqrt54_35[1]),.dout(n2902),.clk(gclk));
	jxor g02685(.dina(w_n2640_0[0]),.dinb(w_n1008_59[2]),.dout(n2903),.clk(gclk));
	jand g02686(.dina(n2903),.dinb(w_asqrt44_37[2]),.dout(n2904),.clk(gclk));
	jxor g02687(.dina(n2904),.dinb(w_n2645_0[0]),.dout(n2905),.clk(gclk));
	jnot g02688(.din(w_n2905_0[1]),.dout(n2906),.clk(gclk));
	jand g02689(.dina(w_n2906_0[1]),.dinb(n2902),.dout(n2907),.clk(gclk));
	jor g02690(.dina(n2907),.dinb(w_n2901_0[1]),.dout(n2908),.clk(gclk));
	jand g02691(.dina(w_n2908_0[2]),.dinb(w_asqrt55_35[0]),.dout(n2909),.clk(gclk));
	jor g02692(.dina(w_n2908_0[1]),.dinb(w_asqrt55_34[2]),.dout(n2910),.clk(gclk));
	jxor g02693(.dina(w_n2647_0[0]),.dinb(w_n884_58[2]),.dout(n2911),.clk(gclk));
	jand g02694(.dina(n2911),.dinb(w_asqrt44_37[1]),.dout(n2912),.clk(gclk));
	jxor g02695(.dina(n2912),.dinb(w_n2652_0[0]),.dout(n2913),.clk(gclk));
	jand g02696(.dina(w_n2913_0[1]),.dinb(n2910),.dout(n2914),.clk(gclk));
	jor g02697(.dina(n2914),.dinb(w_n2909_0[1]),.dout(n2915),.clk(gclk));
	jand g02698(.dina(w_n2915_0[2]),.dinb(w_asqrt56_36[0]),.dout(n2916),.clk(gclk));
	jor g02699(.dina(w_n2915_0[1]),.dinb(w_asqrt56_35[2]),.dout(n2917),.clk(gclk));
	jxor g02700(.dina(w_n2655_0[0]),.dinb(w_n743_59[2]),.dout(n2918),.clk(gclk));
	jand g02701(.dina(n2918),.dinb(w_asqrt44_37[0]),.dout(n2919),.clk(gclk));
	jxor g02702(.dina(n2919),.dinb(w_n2660_0[0]),.dout(n2920),.clk(gclk));
	jnot g02703(.din(w_n2920_0[1]),.dout(n2921),.clk(gclk));
	jand g02704(.dina(w_n2921_0[1]),.dinb(n2917),.dout(n2922),.clk(gclk));
	jor g02705(.dina(n2922),.dinb(w_n2916_0[1]),.dout(n2923),.clk(gclk));
	jand g02706(.dina(w_n2923_0[2]),.dinb(w_asqrt57_35[2]),.dout(n2924),.clk(gclk));
	jor g02707(.dina(w_n2923_0[1]),.dinb(w_asqrt57_35[1]),.dout(n2925),.clk(gclk));
	jxor g02708(.dina(w_n2662_0[0]),.dinb(w_n635_59[2]),.dout(n2926),.clk(gclk));
	jand g02709(.dina(n2926),.dinb(w_asqrt44_36[2]),.dout(n2927),.clk(gclk));
	jxor g02710(.dina(n2927),.dinb(w_n2667_0[0]),.dout(n2928),.clk(gclk));
	jnot g02711(.din(w_n2928_0[1]),.dout(n2929),.clk(gclk));
	jand g02712(.dina(w_n2929_0[1]),.dinb(n2925),.dout(n2930),.clk(gclk));
	jor g02713(.dina(n2930),.dinb(w_n2924_0[1]),.dout(n2931),.clk(gclk));
	jand g02714(.dina(w_n2931_0[2]),.dinb(w_asqrt58_36[1]),.dout(n2932),.clk(gclk));
	jor g02715(.dina(w_n2931_0[1]),.dinb(w_asqrt58_36[0]),.dout(n2933),.clk(gclk));
	jxor g02716(.dina(w_n2669_0[0]),.dinb(w_n515_60[2]),.dout(n2934),.clk(gclk));
	jand g02717(.dina(n2934),.dinb(w_asqrt44_36[1]),.dout(n2935),.clk(gclk));
	jxor g02718(.dina(n2935),.dinb(w_n2674_0[0]),.dout(n2936),.clk(gclk));
	jand g02719(.dina(w_n2936_0[1]),.dinb(n2933),.dout(n2937),.clk(gclk));
	jor g02720(.dina(n2937),.dinb(w_n2932_0[1]),.dout(n2938),.clk(gclk));
	jand g02721(.dina(w_n2938_0[2]),.dinb(w_asqrt59_36[0]),.dout(n2939),.clk(gclk));
	jor g02722(.dina(w_n2938_0[1]),.dinb(w_asqrt59_35[2]),.dout(n2940),.clk(gclk));
	jxor g02723(.dina(w_n2677_0[0]),.dinb(w_n443_60[2]),.dout(n2941),.clk(gclk));
	jand g02724(.dina(n2941),.dinb(w_asqrt44_36[0]),.dout(n2942),.clk(gclk));
	jxor g02725(.dina(n2942),.dinb(w_n2682_0[0]),.dout(n2943),.clk(gclk));
	jand g02726(.dina(w_n2943_0[1]),.dinb(n2940),.dout(n2944),.clk(gclk));
	jor g02727(.dina(n2944),.dinb(w_n2939_0[1]),.dout(n2945),.clk(gclk));
	jand g02728(.dina(w_n2945_0[2]),.dinb(w_asqrt60_36[1]),.dout(n2946),.clk(gclk));
	jor g02729(.dina(w_n2945_0[1]),.dinb(w_asqrt60_36[0]),.dout(n2947),.clk(gclk));
	jxor g02730(.dina(w_n2685_0[0]),.dinb(w_n352_61[0]),.dout(n2948),.clk(gclk));
	jand g02731(.dina(n2948),.dinb(w_asqrt44_35[2]),.dout(n2949),.clk(gclk));
	jxor g02732(.dina(n2949),.dinb(w_n2690_0[0]),.dout(n2950),.clk(gclk));
	jnot g02733(.din(w_n2950_0[1]),.dout(n2951),.clk(gclk));
	jand g02734(.dina(w_n2951_0[1]),.dinb(n2947),.dout(n2952),.clk(gclk));
	jor g02735(.dina(n2952),.dinb(w_n2946_0[1]),.dout(n2953),.clk(gclk));
	jand g02736(.dina(w_n2953_0[2]),.dinb(w_asqrt61_36[1]),.dout(n2954),.clk(gclk));
	jor g02737(.dina(w_n2953_0[1]),.dinb(w_asqrt61_36[0]),.dout(n2955),.clk(gclk));
	jxor g02738(.dina(w_n2692_0[0]),.dinb(w_n294_61[1]),.dout(n2956),.clk(gclk));
	jand g02739(.dina(n2956),.dinb(w_asqrt44_35[1]),.dout(n2957),.clk(gclk));
	jxor g02740(.dina(n2957),.dinb(w_n2697_0[0]),.dout(n2958),.clk(gclk));
	jand g02741(.dina(w_n2958_0[1]),.dinb(n2955),.dout(n2959),.clk(gclk));
	jor g02742(.dina(n2959),.dinb(w_n2954_0[1]),.dout(n2960),.clk(gclk));
	jand g02743(.dina(w_n2960_0[2]),.dinb(w_asqrt62_36[1]),.dout(n2961),.clk(gclk));
	jor g02744(.dina(w_n2960_0[1]),.dinb(w_asqrt62_36[0]),.dout(n2962),.clk(gclk));
	jxor g02745(.dina(w_n2700_0[0]),.dinb(w_n239_61[1]),.dout(n2963),.clk(gclk));
	jand g02746(.dina(n2963),.dinb(w_asqrt44_35[0]),.dout(n2964),.clk(gclk));
	jxor g02747(.dina(n2964),.dinb(w_n2705_0[0]),.dout(n2965),.clk(gclk));
	jand g02748(.dina(w_n2965_0[2]),.dinb(n2962),.dout(n2966),.clk(gclk));
	jor g02749(.dina(n2966),.dinb(w_n2961_0[1]),.dout(n2967),.clk(gclk));
	jxor g02750(.dina(w_n2708_0[0]),.dinb(w_n221_61[2]),.dout(n2968),.clk(gclk));
	jand g02751(.dina(n2968),.dinb(w_asqrt44_34[2]),.dout(n2969),.clk(gclk));
	jxor g02752(.dina(n2969),.dinb(w_n2714_0[0]),.dout(n2970),.clk(gclk));
	jnot g02753(.din(w_n2970_0[2]),.dout(n2971),.clk(gclk));
	jor g02754(.dina(w_n2971_0[1]),.dinb(w_n2967_0[1]),.dout(n2972),.clk(gclk));
	jnot g02755(.din(w_n2972_0[2]),.dout(n2973),.clk(gclk));
	jand g02756(.dina(w_n2831_0[0]),.dinb(w_n2716_0[0]),.dout(n2974),.clk(gclk));
	jnot g02757(.din(n2974),.dout(n2975),.clk(gclk));
	jand g02758(.dina(w_n2720_0[0]),.dinb(w_asqrt63_46[2]),.dout(n2976),.clk(gclk));
	jand g02759(.dina(n2976),.dinb(w_n2744_0[2]),.dout(n2977),.clk(gclk));
	jand g02760(.dina(w_n2977_0[1]),.dinb(n2975),.dout(n2978),.clk(gclk));
	jand g02761(.dina(w_n2730_0[0]),.dinb(w_n2827_0[0]),.dout(n2979),.clk(gclk));
	jnot g02762(.din(w_n2961_0[0]),.dout(n2980),.clk(gclk));
	jnot g02763(.din(w_n2954_0[0]),.dout(n2981),.clk(gclk));
	jnot g02764(.din(w_n2946_0[0]),.dout(n2982),.clk(gclk));
	jnot g02765(.din(w_n2939_0[0]),.dout(n2983),.clk(gclk));
	jnot g02766(.din(w_n2932_0[0]),.dout(n2984),.clk(gclk));
	jnot g02767(.din(w_n2924_0[0]),.dout(n2985),.clk(gclk));
	jnot g02768(.din(w_n2916_0[0]),.dout(n2986),.clk(gclk));
	jnot g02769(.din(w_n2909_0[0]),.dout(n2987),.clk(gclk));
	jnot g02770(.din(w_n2901_0[0]),.dout(n2988),.clk(gclk));
	jnot g02771(.din(w_n2894_0[0]),.dout(n2989),.clk(gclk));
	jnot g02772(.din(w_n2886_0[0]),.dout(n2990),.clk(gclk));
	jnot g02773(.din(w_n2879_0[0]),.dout(n2991),.clk(gclk));
	jnot g02774(.din(w_n2871_0[0]),.dout(n2992),.clk(gclk));
	jnot g02775(.din(w_n2864_0[0]),.dout(n2993),.clk(gclk));
	jnot g02776(.din(w_n2856_0[0]),.dout(n2994),.clk(gclk));
	jnot g02777(.din(w_n2849_0[0]),.dout(n2995),.clk(gclk));
	jnot g02778(.din(w_n2838_0[0]),.dout(n2996),.clk(gclk));
	jnot g02779(.din(w_n2739_0[0]),.dout(n2997),.clk(gclk));
	jor g02780(.dina(w_n2833_55[0]),.dinb(w_n2578_0[2]),.dout(n2998),.clk(gclk));
	jnot g02781(.din(w_n2737_0[0]),.dout(n2999),.clk(gclk));
	jand g02782(.dina(n2999),.dinb(n2998),.dout(n3000),.clk(gclk));
	jand g02783(.dina(n3000),.dinb(w_n2572_57[0]),.dout(n3001),.clk(gclk));
	jor g02784(.dina(w_n2833_54[2]),.dinb(w_a88_0[0]),.dout(n3002),.clk(gclk));
	jand g02785(.dina(n3002),.dinb(w_a89_0[0]),.dout(n3003),.clk(gclk));
	jor g02786(.dina(w_n2840_0[0]),.dinb(n3003),.dout(n3004),.clk(gclk));
	jor g02787(.dina(n3004),.dinb(n3001),.dout(n3005),.clk(gclk));
	jand g02788(.dina(n3005),.dinb(n2997),.dout(n3006),.clk(gclk));
	jand g02789(.dina(n3006),.dinb(w_n2345_55[0]),.dout(n3007),.clk(gclk));
	jor g02790(.dina(w_n2845_0[0]),.dinb(n3007),.dout(n3008),.clk(gclk));
	jand g02791(.dina(n3008),.dinb(n2996),.dout(n3009),.clk(gclk));
	jand g02792(.dina(n3009),.dinb(w_n2108_57[2]),.dout(n3010),.clk(gclk));
	jnot g02793(.din(w_n2853_0[0]),.dout(n3011),.clk(gclk));
	jor g02794(.dina(w_n3011_0[1]),.dinb(n3010),.dout(n3012),.clk(gclk));
	jand g02795(.dina(n3012),.dinb(n2995),.dout(n3013),.clk(gclk));
	jand g02796(.dina(n3013),.dinb(w_n1912_56[0]),.dout(n3014),.clk(gclk));
	jor g02797(.dina(w_n2860_0[0]),.dinb(n3014),.dout(n3015),.clk(gclk));
	jand g02798(.dina(n3015),.dinb(n2994),.dout(n3016),.clk(gclk));
	jand g02799(.dina(n3016),.dinb(w_n1699_58[1]),.dout(n3017),.clk(gclk));
	jnot g02800(.din(w_n2868_0[0]),.dout(n3018),.clk(gclk));
	jor g02801(.dina(w_n3018_0[1]),.dinb(n3017),.dout(n3019),.clk(gclk));
	jand g02802(.dina(n3019),.dinb(n2993),.dout(n3020),.clk(gclk));
	jand g02803(.dina(n3020),.dinb(w_n1516_56[2]),.dout(n3021),.clk(gclk));
	jor g02804(.dina(w_n2875_0[0]),.dinb(n3021),.dout(n3022),.clk(gclk));
	jand g02805(.dina(n3022),.dinb(n2992),.dout(n3023),.clk(gclk));
	jand g02806(.dina(n3023),.dinb(w_n1332_58[1]),.dout(n3024),.clk(gclk));
	jnot g02807(.din(w_n2883_0[0]),.dout(n3025),.clk(gclk));
	jor g02808(.dina(w_n3025_0[1]),.dinb(n3024),.dout(n3026),.clk(gclk));
	jand g02809(.dina(n3026),.dinb(n2991),.dout(n3027),.clk(gclk));
	jand g02810(.dina(n3027),.dinb(w_n1173_57[1]),.dout(n3028),.clk(gclk));
	jor g02811(.dina(w_n2890_0[0]),.dinb(n3028),.dout(n3029),.clk(gclk));
	jand g02812(.dina(n3029),.dinb(n2990),.dout(n3030),.clk(gclk));
	jand g02813(.dina(n3030),.dinb(w_n1008_59[1]),.dout(n3031),.clk(gclk));
	jnot g02814(.din(w_n2898_0[0]),.dout(n3032),.clk(gclk));
	jor g02815(.dina(w_n3032_0[1]),.dinb(n3031),.dout(n3033),.clk(gclk));
	jand g02816(.dina(n3033),.dinb(n2989),.dout(n3034),.clk(gclk));
	jand g02817(.dina(n3034),.dinb(w_n884_58[1]),.dout(n3035),.clk(gclk));
	jor g02818(.dina(w_n2905_0[0]),.dinb(n3035),.dout(n3036),.clk(gclk));
	jand g02819(.dina(n3036),.dinb(n2988),.dout(n3037),.clk(gclk));
	jand g02820(.dina(n3037),.dinb(w_n743_59[1]),.dout(n3038),.clk(gclk));
	jnot g02821(.din(w_n2913_0[0]),.dout(n3039),.clk(gclk));
	jor g02822(.dina(w_n3039_0[1]),.dinb(n3038),.dout(n3040),.clk(gclk));
	jand g02823(.dina(n3040),.dinb(n2987),.dout(n3041),.clk(gclk));
	jand g02824(.dina(n3041),.dinb(w_n635_59[1]),.dout(n3042),.clk(gclk));
	jor g02825(.dina(w_n2920_0[0]),.dinb(n3042),.dout(n3043),.clk(gclk));
	jand g02826(.dina(n3043),.dinb(n2986),.dout(n3044),.clk(gclk));
	jand g02827(.dina(n3044),.dinb(w_n515_60[1]),.dout(n3045),.clk(gclk));
	jor g02828(.dina(w_n2928_0[0]),.dinb(n3045),.dout(n3046),.clk(gclk));
	jand g02829(.dina(n3046),.dinb(n2985),.dout(n3047),.clk(gclk));
	jand g02830(.dina(n3047),.dinb(w_n443_60[1]),.dout(n3048),.clk(gclk));
	jnot g02831(.din(w_n2936_0[0]),.dout(n3049),.clk(gclk));
	jor g02832(.dina(w_n3049_0[1]),.dinb(n3048),.dout(n3050),.clk(gclk));
	jand g02833(.dina(n3050),.dinb(n2984),.dout(n3051),.clk(gclk));
	jand g02834(.dina(n3051),.dinb(w_n352_60[2]),.dout(n3052),.clk(gclk));
	jnot g02835(.din(w_n2943_0[0]),.dout(n3053),.clk(gclk));
	jor g02836(.dina(w_n3053_0[1]),.dinb(n3052),.dout(n3054),.clk(gclk));
	jand g02837(.dina(n3054),.dinb(n2983),.dout(n3055),.clk(gclk));
	jand g02838(.dina(n3055),.dinb(w_n294_61[0]),.dout(n3056),.clk(gclk));
	jor g02839(.dina(w_n2950_0[0]),.dinb(n3056),.dout(n3057),.clk(gclk));
	jand g02840(.dina(n3057),.dinb(n2982),.dout(n3058),.clk(gclk));
	jand g02841(.dina(n3058),.dinb(w_n239_61[0]),.dout(n3059),.clk(gclk));
	jnot g02842(.din(w_n2958_0[0]),.dout(n3060),.clk(gclk));
	jor g02843(.dina(w_n3060_0[1]),.dinb(n3059),.dout(n3061),.clk(gclk));
	jand g02844(.dina(n3061),.dinb(n2981),.dout(n3062),.clk(gclk));
	jand g02845(.dina(n3062),.dinb(w_n221_61[1]),.dout(n3063),.clk(gclk));
	jnot g02846(.din(w_n2965_0[1]),.dout(n3064),.clk(gclk));
	jor g02847(.dina(n3064),.dinb(n3063),.dout(n3065),.clk(gclk));
	jand g02848(.dina(n3065),.dinb(n2980),.dout(n3066),.clk(gclk));
	jor g02849(.dina(w_n2970_0[1]),.dinb(w_n3066_0[1]),.dout(n3067),.clk(gclk));
	jor g02850(.dina(w_n3067_0[1]),.dinb(w_n2717_0[0]),.dout(n3068),.clk(gclk));
	jor g02851(.dina(n3068),.dinb(w_n2979_0[1]),.dout(n3069),.clk(gclk));
	jand g02852(.dina(n3069),.dinb(w_n218_25[1]),.dout(n3070),.clk(gclk));
	jand g02853(.dina(w_n2833_54[1]),.dinb(w_n2576_0[0]),.dout(n3071),.clk(gclk));
	jor g02854(.dina(w_n3071_0[1]),.dinb(w_n3070_0[1]),.dout(n3072),.clk(gclk));
	jor g02855(.dina(n3072),.dinb(w_n2978_0[1]),.dout(n3073),.clk(gclk));
	jor g02856(.dina(w_n3073_0[1]),.dinb(w_n2973_0[2]),.dout(asqrt_fa_44),.clk(gclk));
	jnot g02857(.din(w_a84_0[2]),.dout(n3075),.clk(gclk));
	jnot g02858(.din(w_a85_0[1]),.dout(n3076),.clk(gclk));
	jand g02859(.dina(w_n3076_0[1]),.dinb(w_n3075_1[2]),.dout(n3077),.clk(gclk));
	jand g02860(.dina(w_n3077_0[2]),.dinb(w_n2734_1[0]),.dout(n3078),.clk(gclk));
	jnot g02861(.din(w_n3078_0[1]),.dout(n3079),.clk(gclk));
	jnot g02862(.din(w_n2978_0[0]),.dout(n3080),.clk(gclk));
	jnot g02863(.din(w_n2979_0[0]),.dout(n3081),.clk(gclk));
	jand g02864(.dina(w_n2971_0[0]),.dinb(w_n2967_0[0]),.dout(n3082),.clk(gclk));
	jand g02865(.dina(w_n3082_0[1]),.dinb(w_n2744_0[1]),.dout(n3083),.clk(gclk));
	jand g02866(.dina(n3083),.dinb(n3081),.dout(n3084),.clk(gclk));
	jor g02867(.dina(n3084),.dinb(w_asqrt63_46[1]),.dout(n3085),.clk(gclk));
	jnot g02868(.din(w_n3071_0[0]),.dout(n3086),.clk(gclk));
	jand g02869(.dina(n3086),.dinb(n3085),.dout(n3087),.clk(gclk));
	jand g02870(.dina(n3087),.dinb(n3080),.dout(n3088),.clk(gclk));
	jand g02871(.dina(w_n3088_0[1]),.dinb(w_n2972_0[1]),.dout(n3089),.clk(gclk));
	jor g02872(.dina(w_n3089_62[1]),.dinb(w_n2734_0[2]),.dout(n3090),.clk(gclk));
	jand g02873(.dina(n3090),.dinb(n3079),.dout(n3091),.clk(gclk));
	jor g02874(.dina(w_n3091_0[2]),.dinb(w_n2833_54[0]),.dout(n3092),.clk(gclk));
	jand g02875(.dina(w_n3091_0[1]),.dinb(w_n2833_53[2]),.dout(n3093),.clk(gclk));
	jor g02876(.dina(w_n3089_62[0]),.dinb(w_a86_1[0]),.dout(n3094),.clk(gclk));
	jand g02877(.dina(n3094),.dinb(w_a87_0[0]),.dout(n3095),.clk(gclk));
	jand g02878(.dina(w_asqrt43_32[1]),.dinb(w_n2736_0[1]),.dout(n3096),.clk(gclk));
	jor g02879(.dina(n3096),.dinb(n3095),.dout(n3097),.clk(gclk));
	jor g02880(.dina(n3097),.dinb(n3093),.dout(n3098),.clk(gclk));
	jand g02881(.dina(n3098),.dinb(w_n3092_0[1]),.dout(n3099),.clk(gclk));
	jor g02882(.dina(w_n3099_0[2]),.dinb(w_n2572_56[2]),.dout(n3100),.clk(gclk));
	jand g02883(.dina(w_n3099_0[1]),.dinb(w_n2572_56[1]),.dout(n3101),.clk(gclk));
	jnot g02884(.din(w_n2736_0[0]),.dout(n3102),.clk(gclk));
	jor g02885(.dina(w_n3089_61[2]),.dinb(n3102),.dout(n3103),.clk(gclk));
	jor g02886(.dina(w_n2977_0[0]),.dinb(w_n2973_0[1]),.dout(n3104),.clk(gclk));
	jor g02887(.dina(n3104),.dinb(w_n3070_0[0]),.dout(n3105),.clk(gclk));
	jor g02888(.dina(n3105),.dinb(w_n2833_53[1]),.dout(n3106),.clk(gclk));
	jand g02889(.dina(n3106),.dinb(w_n3103_0[1]),.dout(n3107),.clk(gclk));
	jxor g02890(.dina(n3107),.dinb(w_n2578_0[1]),.dout(n3108),.clk(gclk));
	jor g02891(.dina(w_n3108_0[1]),.dinb(n3101),.dout(n3109),.clk(gclk));
	jand g02892(.dina(n3109),.dinb(w_n3100_0[1]),.dout(n3110),.clk(gclk));
	jor g02893(.dina(w_n3110_0[2]),.dinb(w_n2345_54[2]),.dout(n3111),.clk(gclk));
	jand g02894(.dina(w_n3110_0[1]),.dinb(w_n2345_54[1]),.dout(n3112),.clk(gclk));
	jxor g02895(.dina(w_n2738_0[0]),.dinb(w_n2572_56[0]),.dout(n3113),.clk(gclk));
	jor g02896(.dina(n3113),.dinb(w_n3089_61[1]),.dout(n3114),.clk(gclk));
	jxor g02897(.dina(n3114),.dinb(w_n2835_0[0]),.dout(n3115),.clk(gclk));
	jor g02898(.dina(w_n3115_0[2]),.dinb(n3112),.dout(n3116),.clk(gclk));
	jand g02899(.dina(n3116),.dinb(w_n3111_0[1]),.dout(n3117),.clk(gclk));
	jor g02900(.dina(w_n3117_0[2]),.dinb(w_n2108_57[1]),.dout(n3118),.clk(gclk));
	jand g02901(.dina(w_n3117_0[1]),.dinb(w_n2108_57[0]),.dout(n3119),.clk(gclk));
	jxor g02902(.dina(w_n2837_0[0]),.dinb(w_n2345_54[0]),.dout(n3120),.clk(gclk));
	jor g02903(.dina(n3120),.dinb(w_n3089_61[0]),.dout(n3121),.clk(gclk));
	jxor g02904(.dina(n3121),.dinb(w_n2846_0[0]),.dout(n3122),.clk(gclk));
	jor g02905(.dina(w_n3122_0[2]),.dinb(n3119),.dout(n3123),.clk(gclk));
	jand g02906(.dina(n3123),.dinb(w_n3118_0[1]),.dout(n3124),.clk(gclk));
	jor g02907(.dina(w_n3124_0[2]),.dinb(w_n1912_55[2]),.dout(n3125),.clk(gclk));
	jand g02908(.dina(w_n3124_0[1]),.dinb(w_n1912_55[1]),.dout(n3126),.clk(gclk));
	jxor g02909(.dina(w_n2848_0[0]),.dinb(w_n2108_56[2]),.dout(n3127),.clk(gclk));
	jor g02910(.dina(n3127),.dinb(w_n3089_60[2]),.dout(n3128),.clk(gclk));
	jxor g02911(.dina(n3128),.dinb(w_n3011_0[0]),.dout(n3129),.clk(gclk));
	jnot g02912(.din(w_n3129_0[2]),.dout(n3130),.clk(gclk));
	jor g02913(.dina(n3130),.dinb(n3126),.dout(n3131),.clk(gclk));
	jand g02914(.dina(n3131),.dinb(w_n3125_0[1]),.dout(n3132),.clk(gclk));
	jor g02915(.dina(w_n3132_0[2]),.dinb(w_n1699_58[0]),.dout(n3133),.clk(gclk));
	jand g02916(.dina(w_n3132_0[1]),.dinb(w_n1699_57[2]),.dout(n3134),.clk(gclk));
	jxor g02917(.dina(w_n2855_0[0]),.dinb(w_n1912_55[0]),.dout(n3135),.clk(gclk));
	jor g02918(.dina(n3135),.dinb(w_n3089_60[1]),.dout(n3136),.clk(gclk));
	jxor g02919(.dina(n3136),.dinb(w_n2861_0[0]),.dout(n3137),.clk(gclk));
	jor g02920(.dina(w_n3137_0[2]),.dinb(n3134),.dout(n3138),.clk(gclk));
	jand g02921(.dina(n3138),.dinb(w_n3133_0[1]),.dout(n3139),.clk(gclk));
	jor g02922(.dina(w_n3139_0[2]),.dinb(w_n1516_56[1]),.dout(n3140),.clk(gclk));
	jand g02923(.dina(w_n3139_0[1]),.dinb(w_n1516_56[0]),.dout(n3141),.clk(gclk));
	jxor g02924(.dina(w_n2863_0[0]),.dinb(w_n1699_57[1]),.dout(n3142),.clk(gclk));
	jor g02925(.dina(n3142),.dinb(w_n3089_60[0]),.dout(n3143),.clk(gclk));
	jxor g02926(.dina(n3143),.dinb(w_n3018_0[0]),.dout(n3144),.clk(gclk));
	jnot g02927(.din(w_n3144_0[2]),.dout(n3145),.clk(gclk));
	jor g02928(.dina(n3145),.dinb(n3141),.dout(n3146),.clk(gclk));
	jand g02929(.dina(n3146),.dinb(w_n3140_0[1]),.dout(n3147),.clk(gclk));
	jor g02930(.dina(w_n3147_0[2]),.dinb(w_n1332_58[0]),.dout(n3148),.clk(gclk));
	jand g02931(.dina(w_n3147_0[1]),.dinb(w_n1332_57[2]),.dout(n3149),.clk(gclk));
	jxor g02932(.dina(w_n2870_0[0]),.dinb(w_n1516_55[2]),.dout(n3150),.clk(gclk));
	jor g02933(.dina(n3150),.dinb(w_n3089_59[2]),.dout(n3151),.clk(gclk));
	jxor g02934(.dina(n3151),.dinb(w_n2876_0[0]),.dout(n3152),.clk(gclk));
	jor g02935(.dina(w_n3152_0[2]),.dinb(n3149),.dout(n3153),.clk(gclk));
	jand g02936(.dina(n3153),.dinb(w_n3148_0[1]),.dout(n3154),.clk(gclk));
	jor g02937(.dina(w_n3154_0[2]),.dinb(w_n1173_57[0]),.dout(n3155),.clk(gclk));
	jand g02938(.dina(w_n3154_0[1]),.dinb(w_n1173_56[2]),.dout(n3156),.clk(gclk));
	jxor g02939(.dina(w_n2878_0[0]),.dinb(w_n1332_57[1]),.dout(n3157),.clk(gclk));
	jor g02940(.dina(n3157),.dinb(w_n3089_59[1]),.dout(n3158),.clk(gclk));
	jxor g02941(.dina(n3158),.dinb(w_n3025_0[0]),.dout(n3159),.clk(gclk));
	jnot g02942(.din(w_n3159_0[2]),.dout(n3160),.clk(gclk));
	jor g02943(.dina(n3160),.dinb(n3156),.dout(n3161),.clk(gclk));
	jand g02944(.dina(n3161),.dinb(w_n3155_0[1]),.dout(n3162),.clk(gclk));
	jor g02945(.dina(w_n3162_0[2]),.dinb(w_n1008_59[0]),.dout(n3163),.clk(gclk));
	jand g02946(.dina(w_n3162_0[1]),.dinb(w_n1008_58[2]),.dout(n3164),.clk(gclk));
	jxor g02947(.dina(w_n2885_0[0]),.dinb(w_n1173_56[1]),.dout(n3165),.clk(gclk));
	jor g02948(.dina(n3165),.dinb(w_n3089_59[0]),.dout(n3166),.clk(gclk));
	jxor g02949(.dina(n3166),.dinb(w_n2891_0[0]),.dout(n3167),.clk(gclk));
	jor g02950(.dina(w_n3167_0[2]),.dinb(n3164),.dout(n3168),.clk(gclk));
	jand g02951(.dina(n3168),.dinb(w_n3163_0[1]),.dout(n3169),.clk(gclk));
	jor g02952(.dina(w_n3169_0[2]),.dinb(w_n884_58[0]),.dout(n3170),.clk(gclk));
	jand g02953(.dina(w_n3169_0[1]),.dinb(w_n884_57[2]),.dout(n3171),.clk(gclk));
	jxor g02954(.dina(w_n2893_0[0]),.dinb(w_n1008_58[1]),.dout(n3172),.clk(gclk));
	jor g02955(.dina(n3172),.dinb(w_n3089_58[2]),.dout(n3173),.clk(gclk));
	jxor g02956(.dina(n3173),.dinb(w_n3032_0[0]),.dout(n3174),.clk(gclk));
	jnot g02957(.din(w_n3174_0[2]),.dout(n3175),.clk(gclk));
	jor g02958(.dina(n3175),.dinb(n3171),.dout(n3176),.clk(gclk));
	jand g02959(.dina(n3176),.dinb(w_n3170_0[1]),.dout(n3177),.clk(gclk));
	jor g02960(.dina(w_n3177_0[2]),.dinb(w_n743_59[0]),.dout(n3178),.clk(gclk));
	jand g02961(.dina(w_n3177_0[1]),.dinb(w_n743_58[2]),.dout(n3179),.clk(gclk));
	jxor g02962(.dina(w_n2900_0[0]),.dinb(w_n884_57[1]),.dout(n3180),.clk(gclk));
	jor g02963(.dina(n3180),.dinb(w_n3089_58[1]),.dout(n3181),.clk(gclk));
	jxor g02964(.dina(n3181),.dinb(w_n2906_0[0]),.dout(n3182),.clk(gclk));
	jor g02965(.dina(w_n3182_0[2]),.dinb(n3179),.dout(n3183),.clk(gclk));
	jand g02966(.dina(n3183),.dinb(w_n3178_0[1]),.dout(n3184),.clk(gclk));
	jor g02967(.dina(w_n3184_0[2]),.dinb(w_n635_59[0]),.dout(n3185),.clk(gclk));
	jand g02968(.dina(w_n3184_0[1]),.dinb(w_n635_58[2]),.dout(n3186),.clk(gclk));
	jxor g02969(.dina(w_n2908_0[0]),.dinb(w_n743_58[1]),.dout(n3187),.clk(gclk));
	jor g02970(.dina(n3187),.dinb(w_n3089_58[0]),.dout(n3188),.clk(gclk));
	jxor g02971(.dina(n3188),.dinb(w_n3039_0[0]),.dout(n3189),.clk(gclk));
	jnot g02972(.din(w_n3189_0[2]),.dout(n3190),.clk(gclk));
	jor g02973(.dina(n3190),.dinb(n3186),.dout(n3191),.clk(gclk));
	jand g02974(.dina(n3191),.dinb(w_n3185_0[1]),.dout(n3192),.clk(gclk));
	jor g02975(.dina(w_n3192_0[2]),.dinb(w_n515_60[0]),.dout(n3193),.clk(gclk));
	jand g02976(.dina(w_n3192_0[1]),.dinb(w_n515_59[2]),.dout(n3194),.clk(gclk));
	jxor g02977(.dina(w_n2915_0[0]),.dinb(w_n635_58[1]),.dout(n3195),.clk(gclk));
	jor g02978(.dina(n3195),.dinb(w_n3089_57[2]),.dout(n3196),.clk(gclk));
	jxor g02979(.dina(n3196),.dinb(w_n2921_0[0]),.dout(n3197),.clk(gclk));
	jor g02980(.dina(w_n3197_0[2]),.dinb(n3194),.dout(n3198),.clk(gclk));
	jand g02981(.dina(n3198),.dinb(w_n3193_0[1]),.dout(n3199),.clk(gclk));
	jor g02982(.dina(w_n3199_0[2]),.dinb(w_n443_60[0]),.dout(n3200),.clk(gclk));
	jand g02983(.dina(w_n3199_0[1]),.dinb(w_n443_59[2]),.dout(n3201),.clk(gclk));
	jxor g02984(.dina(w_n2923_0[0]),.dinb(w_n515_59[1]),.dout(n3202),.clk(gclk));
	jor g02985(.dina(n3202),.dinb(w_n3089_57[1]),.dout(n3203),.clk(gclk));
	jxor g02986(.dina(n3203),.dinb(w_n2929_0[0]),.dout(n3204),.clk(gclk));
	jor g02987(.dina(w_n3204_0[2]),.dinb(n3201),.dout(n3205),.clk(gclk));
	jand g02988(.dina(n3205),.dinb(w_n3200_0[1]),.dout(n3206),.clk(gclk));
	jor g02989(.dina(w_n3206_0[2]),.dinb(w_n352_60[1]),.dout(n3207),.clk(gclk));
	jand g02990(.dina(w_n3206_0[1]),.dinb(w_n352_60[0]),.dout(n3208),.clk(gclk));
	jxor g02991(.dina(w_n2931_0[0]),.dinb(w_n443_59[1]),.dout(n3209),.clk(gclk));
	jor g02992(.dina(n3209),.dinb(w_n3089_57[0]),.dout(n3210),.clk(gclk));
	jxor g02993(.dina(n3210),.dinb(w_n3049_0[0]),.dout(n3211),.clk(gclk));
	jnot g02994(.din(w_n3211_0[2]),.dout(n3212),.clk(gclk));
	jor g02995(.dina(n3212),.dinb(n3208),.dout(n3213),.clk(gclk));
	jand g02996(.dina(n3213),.dinb(w_n3207_0[1]),.dout(n3214),.clk(gclk));
	jor g02997(.dina(w_n3214_0[2]),.dinb(w_n294_60[2]),.dout(n3215),.clk(gclk));
	jand g02998(.dina(w_n3214_0[1]),.dinb(w_n294_60[1]),.dout(n3216),.clk(gclk));
	jxor g02999(.dina(w_n2938_0[0]),.dinb(w_n352_59[2]),.dout(n3217),.clk(gclk));
	jor g03000(.dina(n3217),.dinb(w_n3089_56[2]),.dout(n3218),.clk(gclk));
	jxor g03001(.dina(n3218),.dinb(w_n3053_0[0]),.dout(n3219),.clk(gclk));
	jnot g03002(.din(w_n3219_0[2]),.dout(n3220),.clk(gclk));
	jor g03003(.dina(n3220),.dinb(n3216),.dout(n3221),.clk(gclk));
	jand g03004(.dina(n3221),.dinb(w_n3215_0[1]),.dout(n3222),.clk(gclk));
	jor g03005(.dina(w_n3222_0[2]),.dinb(w_n239_60[2]),.dout(n3223),.clk(gclk));
	jand g03006(.dina(w_n3222_0[1]),.dinb(w_n239_60[1]),.dout(n3224),.clk(gclk));
	jxor g03007(.dina(w_n2945_0[0]),.dinb(w_n294_60[0]),.dout(n3225),.clk(gclk));
	jor g03008(.dina(n3225),.dinb(w_n3089_56[1]),.dout(n3226),.clk(gclk));
	jxor g03009(.dina(n3226),.dinb(w_n2951_0[0]),.dout(n3227),.clk(gclk));
	jor g03010(.dina(w_n3227_0[2]),.dinb(n3224),.dout(n3228),.clk(gclk));
	jand g03011(.dina(n3228),.dinb(w_n3223_0[1]),.dout(n3229),.clk(gclk));
	jor g03012(.dina(w_n3229_0[2]),.dinb(w_n221_61[0]),.dout(n3230),.clk(gclk));
	jand g03013(.dina(w_n3229_0[1]),.dinb(w_n221_60[2]),.dout(n3231),.clk(gclk));
	jxor g03014(.dina(w_n2953_0[0]),.dinb(w_n239_60[0]),.dout(n3232),.clk(gclk));
	jor g03015(.dina(n3232),.dinb(w_n3089_56[0]),.dout(n3233),.clk(gclk));
	jxor g03016(.dina(n3233),.dinb(w_n3060_0[0]),.dout(n3234),.clk(gclk));
	jnot g03017(.din(w_n3234_0[1]),.dout(n3235),.clk(gclk));
	jor g03018(.dina(w_n3235_0[1]),.dinb(n3231),.dout(n3236),.clk(gclk));
	jand g03019(.dina(n3236),.dinb(w_n3230_0[1]),.dout(n3237),.clk(gclk));
	jxor g03020(.dina(w_n2960_0[0]),.dinb(w_n221_60[1]),.dout(n3238),.clk(gclk));
	jor g03021(.dina(n3238),.dinb(w_n3089_55[2]),.dout(n3239),.clk(gclk));
	jxor g03022(.dina(n3239),.dinb(w_n2965_0[0]),.dout(n3240),.clk(gclk));
	jand g03023(.dina(w_n3240_1[1]),.dinb(w_n3237_1[1]),.dout(n3241),.clk(gclk));
	jand g03024(.dina(w_n3088_0[0]),.dinb(w_n3066_0[0]),.dout(n3242),.clk(gclk));
	jand g03025(.dina(w_n3067_0[0]),.dinb(w_asqrt63_46[0]),.dout(n3243),.clk(gclk));
	jand g03026(.dina(n3243),.dinb(w_n2972_0[0]),.dout(n3244),.clk(gclk));
	jnot g03027(.din(n3244),.dout(n3245),.clk(gclk));
	jor g03028(.dina(w_n3245_0[1]),.dinb(n3242),.dout(n3246),.clk(gclk));
	jnot g03029(.din(w_n3246_0[1]),.dout(n3247),.clk(gclk));
	jor g03030(.dina(w_n3240_1[0]),.dinb(w_n3237_1[0]),.dout(n3248),.clk(gclk));
	jand g03031(.dina(w_n3073_0[0]),.dinb(w_n3082_0[0]),.dout(n3249),.clk(gclk));
	jor g03032(.dina(n3249),.dinb(w_n2973_0[0]),.dout(n3250),.clk(gclk));
	jor g03033(.dina(w_n3250_0[1]),.dinb(n3248),.dout(n3251),.clk(gclk));
	jand g03034(.dina(n3251),.dinb(w_n218_25[0]),.dout(n3252),.clk(gclk));
	jand g03035(.dina(w_n3089_55[1]),.dinb(w_n2970_0[0]),.dout(n3253),.clk(gclk));
	jor g03036(.dina(w_n3253_0[1]),.dinb(n3252),.dout(n3254),.clk(gclk));
	jor g03037(.dina(n3254),.dinb(n3247),.dout(n3255),.clk(gclk));
	jor g03038(.dina(n3255),.dinb(w_n3241_0[1]),.dout(asqrt_fa_43),.clk(gclk));
	jand g03039(.dina(w_asqrt42_41),.dinb(w_a84_0[1]),.dout(n3257),.clk(gclk));
	jnot g03040(.din(w_a82_1[1]),.dout(n3258),.clk(gclk));
	jnot g03041(.din(w_a83_0[1]),.dout(n3259),.clk(gclk));
	jand g03042(.dina(w_n3259_0[1]),.dinb(w_n3258_1[1]),.dout(n3260),.clk(gclk));
	jand g03043(.dina(w_n3260_0[2]),.dinb(w_n3075_1[1]),.dout(n3261),.clk(gclk));
	jor g03044(.dina(w_n3261_0[1]),.dinb(n3257),.dout(n3262),.clk(gclk));
	jand g03045(.dina(w_n3262_0[2]),.dinb(w_asqrt43_32[0]),.dout(n3263),.clk(gclk));
	jor g03046(.dina(w_n3262_0[1]),.dinb(w_asqrt43_31[2]),.dout(n3264),.clk(gclk));
	jand g03047(.dina(w_asqrt42_40[2]),.dinb(w_n3075_1[0]),.dout(n3265),.clk(gclk));
	jor g03048(.dina(n3265),.dinb(w_n3076_0[0]),.dout(n3266),.clk(gclk));
	jnot g03049(.din(w_n3077_0[1]),.dout(n3267),.clk(gclk));
	jnot g03050(.din(w_n3241_0[0]),.dout(n3268),.clk(gclk));
	jnot g03051(.din(w_n3230_0[0]),.dout(n3269),.clk(gclk));
	jnot g03052(.din(w_n3223_0[0]),.dout(n3270),.clk(gclk));
	jnot g03053(.din(w_n3215_0[0]),.dout(n3271),.clk(gclk));
	jnot g03054(.din(w_n3207_0[0]),.dout(n3272),.clk(gclk));
	jnot g03055(.din(w_n3200_0[0]),.dout(n3273),.clk(gclk));
	jnot g03056(.din(w_n3193_0[0]),.dout(n3274),.clk(gclk));
	jnot g03057(.din(w_n3185_0[0]),.dout(n3275),.clk(gclk));
	jnot g03058(.din(w_n3178_0[0]),.dout(n3276),.clk(gclk));
	jnot g03059(.din(w_n3170_0[0]),.dout(n3277),.clk(gclk));
	jnot g03060(.din(w_n3163_0[0]),.dout(n3278),.clk(gclk));
	jnot g03061(.din(w_n3155_0[0]),.dout(n3279),.clk(gclk));
	jnot g03062(.din(w_n3148_0[0]),.dout(n3280),.clk(gclk));
	jnot g03063(.din(w_n3140_0[0]),.dout(n3281),.clk(gclk));
	jnot g03064(.din(w_n3133_0[0]),.dout(n3282),.clk(gclk));
	jnot g03065(.din(w_n3125_0[0]),.dout(n3283),.clk(gclk));
	jnot g03066(.din(w_n3118_0[0]),.dout(n3284),.clk(gclk));
	jnot g03067(.din(w_n3111_0[0]),.dout(n3285),.clk(gclk));
	jnot g03068(.din(w_n3100_0[0]),.dout(n3286),.clk(gclk));
	jnot g03069(.din(w_n3092_0[0]),.dout(n3287),.clk(gclk));
	jand g03070(.dina(w_asqrt43_31[1]),.dinb(w_a86_0[2]),.dout(n3288),.clk(gclk));
	jor g03071(.dina(n3288),.dinb(w_n3078_0[0]),.dout(n3289),.clk(gclk));
	jor g03072(.dina(n3289),.dinb(w_asqrt44_34[1]),.dout(n3290),.clk(gclk));
	jand g03073(.dina(w_asqrt43_31[0]),.dinb(w_n2734_0[1]),.dout(n3291),.clk(gclk));
	jor g03074(.dina(n3291),.dinb(w_n2735_0[0]),.dout(n3292),.clk(gclk));
	jand g03075(.dina(w_n3103_0[0]),.dinb(n3292),.dout(n3293),.clk(gclk));
	jand g03076(.dina(w_n3293_0[1]),.dinb(n3290),.dout(n3294),.clk(gclk));
	jor g03077(.dina(n3294),.dinb(n3287),.dout(n3295),.clk(gclk));
	jor g03078(.dina(n3295),.dinb(w_asqrt45_32[0]),.dout(n3296),.clk(gclk));
	jnot g03079(.din(w_n3108_0[0]),.dout(n3297),.clk(gclk));
	jand g03080(.dina(w_n3297_0[1]),.dinb(n3296),.dout(n3298),.clk(gclk));
	jor g03081(.dina(n3298),.dinb(n3286),.dout(n3299),.clk(gclk));
	jor g03082(.dina(n3299),.dinb(w_asqrt46_34[1]),.dout(n3300),.clk(gclk));
	jnot g03083(.din(w_n3115_0[1]),.dout(n3301),.clk(gclk));
	jand g03084(.dina(n3301),.dinb(n3300),.dout(n3302),.clk(gclk));
	jor g03085(.dina(n3302),.dinb(n3285),.dout(n3303),.clk(gclk));
	jor g03086(.dina(n3303),.dinb(w_asqrt47_32[2]),.dout(n3304),.clk(gclk));
	jnot g03087(.din(w_n3122_0[1]),.dout(n3305),.clk(gclk));
	jand g03088(.dina(n3305),.dinb(n3304),.dout(n3306),.clk(gclk));
	jor g03089(.dina(n3306),.dinb(n3284),.dout(n3307),.clk(gclk));
	jor g03090(.dina(n3307),.dinb(w_asqrt48_34[2]),.dout(n3308),.clk(gclk));
	jand g03091(.dina(w_n3129_0[1]),.dinb(n3308),.dout(n3309),.clk(gclk));
	jor g03092(.dina(n3309),.dinb(n3283),.dout(n3310),.clk(gclk));
	jor g03093(.dina(n3310),.dinb(w_asqrt49_33[0]),.dout(n3311),.clk(gclk));
	jnot g03094(.din(w_n3137_0[1]),.dout(n3312),.clk(gclk));
	jand g03095(.dina(n3312),.dinb(n3311),.dout(n3313),.clk(gclk));
	jor g03096(.dina(n3313),.dinb(n3282),.dout(n3314),.clk(gclk));
	jor g03097(.dina(n3314),.dinb(w_asqrt50_35[0]),.dout(n3315),.clk(gclk));
	jand g03098(.dina(w_n3144_0[1]),.dinb(n3315),.dout(n3316),.clk(gclk));
	jor g03099(.dina(n3316),.dinb(n3281),.dout(n3317),.clk(gclk));
	jor g03100(.dina(n3317),.dinb(w_asqrt51_33[1]),.dout(n3318),.clk(gclk));
	jnot g03101(.din(w_n3152_0[1]),.dout(n3319),.clk(gclk));
	jand g03102(.dina(n3319),.dinb(n3318),.dout(n3320),.clk(gclk));
	jor g03103(.dina(n3320),.dinb(n3280),.dout(n3321),.clk(gclk));
	jor g03104(.dina(n3321),.dinb(w_asqrt52_35[0]),.dout(n3322),.clk(gclk));
	jand g03105(.dina(w_n3159_0[1]),.dinb(n3322),.dout(n3323),.clk(gclk));
	jor g03106(.dina(n3323),.dinb(n3279),.dout(n3324),.clk(gclk));
	jor g03107(.dina(n3324),.dinb(w_asqrt53_34[0]),.dout(n3325),.clk(gclk));
	jnot g03108(.din(w_n3167_0[1]),.dout(n3326),.clk(gclk));
	jand g03109(.dina(n3326),.dinb(n3325),.dout(n3327),.clk(gclk));
	jor g03110(.dina(n3327),.dinb(n3278),.dout(n3328),.clk(gclk));
	jor g03111(.dina(n3328),.dinb(w_asqrt54_35[0]),.dout(n3329),.clk(gclk));
	jand g03112(.dina(w_n3174_0[1]),.dinb(n3329),.dout(n3330),.clk(gclk));
	jor g03113(.dina(n3330),.dinb(n3277),.dout(n3331),.clk(gclk));
	jor g03114(.dina(n3331),.dinb(w_asqrt55_34[1]),.dout(n3332),.clk(gclk));
	jnot g03115(.din(w_n3182_0[1]),.dout(n3333),.clk(gclk));
	jand g03116(.dina(n3333),.dinb(n3332),.dout(n3334),.clk(gclk));
	jor g03117(.dina(n3334),.dinb(n3276),.dout(n3335),.clk(gclk));
	jor g03118(.dina(n3335),.dinb(w_asqrt56_35[1]),.dout(n3336),.clk(gclk));
	jand g03119(.dina(w_n3189_0[1]),.dinb(n3336),.dout(n3337),.clk(gclk));
	jor g03120(.dina(n3337),.dinb(n3275),.dout(n3338),.clk(gclk));
	jor g03121(.dina(n3338),.dinb(w_asqrt57_35[0]),.dout(n3339),.clk(gclk));
	jnot g03122(.din(w_n3197_0[1]),.dout(n3340),.clk(gclk));
	jand g03123(.dina(n3340),.dinb(n3339),.dout(n3341),.clk(gclk));
	jor g03124(.dina(n3341),.dinb(n3274),.dout(n3342),.clk(gclk));
	jor g03125(.dina(n3342),.dinb(w_asqrt58_35[2]),.dout(n3343),.clk(gclk));
	jnot g03126(.din(w_n3204_0[1]),.dout(n3344),.clk(gclk));
	jand g03127(.dina(n3344),.dinb(n3343),.dout(n3345),.clk(gclk));
	jor g03128(.dina(n3345),.dinb(n3273),.dout(n3346),.clk(gclk));
	jor g03129(.dina(n3346),.dinb(w_asqrt59_35[1]),.dout(n3347),.clk(gclk));
	jand g03130(.dina(w_n3211_0[1]),.dinb(n3347),.dout(n3348),.clk(gclk));
	jor g03131(.dina(n3348),.dinb(n3272),.dout(n3349),.clk(gclk));
	jor g03132(.dina(n3349),.dinb(w_asqrt60_35[2]),.dout(n3350),.clk(gclk));
	jand g03133(.dina(w_n3219_0[1]),.dinb(n3350),.dout(n3351),.clk(gclk));
	jor g03134(.dina(n3351),.dinb(n3271),.dout(n3352),.clk(gclk));
	jor g03135(.dina(n3352),.dinb(w_asqrt61_35[2]),.dout(n3353),.clk(gclk));
	jnot g03136(.din(w_n3227_0[1]),.dout(n3354),.clk(gclk));
	jand g03137(.dina(n3354),.dinb(n3353),.dout(n3355),.clk(gclk));
	jor g03138(.dina(n3355),.dinb(n3270),.dout(n3356),.clk(gclk));
	jor g03139(.dina(n3356),.dinb(w_asqrt62_35[2]),.dout(n3357),.clk(gclk));
	jand g03140(.dina(w_n3234_0[0]),.dinb(n3357),.dout(n3358),.clk(gclk));
	jor g03141(.dina(n3358),.dinb(n3269),.dout(n3359),.clk(gclk));
	jnot g03142(.din(w_n3240_0[2]),.dout(n3360),.clk(gclk));
	jand g03143(.dina(n3360),.dinb(n3359),.dout(n3361),.clk(gclk));
	jnot g03144(.din(w_n3250_0[0]),.dout(n3362),.clk(gclk));
	jand g03145(.dina(n3362),.dinb(n3361),.dout(n3363),.clk(gclk));
	jor g03146(.dina(n3363),.dinb(w_asqrt63_45[2]),.dout(n3364),.clk(gclk));
	jnot g03147(.din(w_n3253_0[0]),.dout(n3365),.clk(gclk));
	jand g03148(.dina(n3365),.dinb(w_n3364_0[1]),.dout(n3366),.clk(gclk));
	jand g03149(.dina(n3366),.dinb(w_n3246_0[0]),.dout(n3367),.clk(gclk));
	jand g03150(.dina(w_n3367_0[1]),.dinb(w_n3268_0[1]),.dout(n3368),.clk(gclk));
	jor g03151(.dina(w_n3368_52[1]),.dinb(n3267),.dout(n3369),.clk(gclk));
	jand g03152(.dina(n3369),.dinb(n3266),.dout(n3370),.clk(gclk));
	jand g03153(.dina(n3370),.dinb(n3264),.dout(n3371),.clk(gclk));
	jor g03154(.dina(n3371),.dinb(w_n3263_0[1]),.dout(n3372),.clk(gclk));
	jand g03155(.dina(w_n3372_0[2]),.dinb(w_asqrt44_34[0]),.dout(n3373),.clk(gclk));
	jor g03156(.dina(w_n3372_0[1]),.dinb(w_asqrt44_33[2]),.dout(n3374),.clk(gclk));
	jand g03157(.dina(w_asqrt42_40[1]),.dinb(w_n3077_0[0]),.dout(n3375),.clk(gclk));
	jand g03158(.dina(w_n3268_0[0]),.dinb(w_asqrt43_30[2]),.dout(n3376),.clk(gclk));
	jand g03159(.dina(n3376),.dinb(w_n3245_0[0]),.dout(n3377),.clk(gclk));
	jand g03160(.dina(n3377),.dinb(w_n3364_0[0]),.dout(n3378),.clk(gclk));
	jor g03161(.dina(n3378),.dinb(w_n3375_0[1]),.dout(n3379),.clk(gclk));
	jxor g03162(.dina(n3379),.dinb(w_a86_0[1]),.dout(n3380),.clk(gclk));
	jnot g03163(.din(w_n3380_0[1]),.dout(n3381),.clk(gclk));
	jand g03164(.dina(w_n3381_0[1]),.dinb(n3374),.dout(n3382),.clk(gclk));
	jor g03165(.dina(n3382),.dinb(w_n3373_0[1]),.dout(n3383),.clk(gclk));
	jand g03166(.dina(w_n3383_0[2]),.dinb(w_asqrt45_31[2]),.dout(n3384),.clk(gclk));
	jor g03167(.dina(w_n3383_0[1]),.dinb(w_asqrt45_31[1]),.dout(n3385),.clk(gclk));
	jxor g03168(.dina(w_n3091_0[0]),.dinb(w_n2833_53[0]),.dout(n3386),.clk(gclk));
	jand g03169(.dina(n3386),.dinb(w_asqrt42_40[0]),.dout(n3387),.clk(gclk));
	jxor g03170(.dina(n3387),.dinb(w_n3293_0[0]),.dout(n3388),.clk(gclk));
	jand g03171(.dina(w_n3388_0[1]),.dinb(n3385),.dout(n3389),.clk(gclk));
	jor g03172(.dina(n3389),.dinb(w_n3384_0[1]),.dout(n3390),.clk(gclk));
	jand g03173(.dina(w_n3390_0[2]),.dinb(w_asqrt46_34[0]),.dout(n3391),.clk(gclk));
	jor g03174(.dina(w_n3390_0[1]),.dinb(w_asqrt46_33[2]),.dout(n3392),.clk(gclk));
	jxor g03175(.dina(w_n3099_0[0]),.dinb(w_n2572_55[2]),.dout(n3393),.clk(gclk));
	jand g03176(.dina(n3393),.dinb(w_asqrt42_39[2]),.dout(n3394),.clk(gclk));
	jxor g03177(.dina(n3394),.dinb(w_n3297_0[0]),.dout(n3395),.clk(gclk));
	jand g03178(.dina(w_n3395_0[1]),.dinb(n3392),.dout(n3396),.clk(gclk));
	jor g03179(.dina(n3396),.dinb(w_n3391_0[1]),.dout(n3397),.clk(gclk));
	jand g03180(.dina(w_n3397_0[2]),.dinb(w_asqrt47_32[1]),.dout(n3398),.clk(gclk));
	jor g03181(.dina(w_n3397_0[1]),.dinb(w_asqrt47_32[0]),.dout(n3399),.clk(gclk));
	jxor g03182(.dina(w_n3110_0[0]),.dinb(w_n2345_53[2]),.dout(n3400),.clk(gclk));
	jand g03183(.dina(n3400),.dinb(w_asqrt42_39[1]),.dout(n3401),.clk(gclk));
	jxor g03184(.dina(n3401),.dinb(w_n3115_0[0]),.dout(n3402),.clk(gclk));
	jnot g03185(.din(w_n3402_0[1]),.dout(n3403),.clk(gclk));
	jand g03186(.dina(w_n3403_0[1]),.dinb(n3399),.dout(n3404),.clk(gclk));
	jor g03187(.dina(n3404),.dinb(w_n3398_0[1]),.dout(n3405),.clk(gclk));
	jand g03188(.dina(w_n3405_0[2]),.dinb(w_asqrt48_34[1]),.dout(n3406),.clk(gclk));
	jor g03189(.dina(w_n3405_0[1]),.dinb(w_asqrt48_34[0]),.dout(n3407),.clk(gclk));
	jxor g03190(.dina(w_n3117_0[0]),.dinb(w_n2108_56[1]),.dout(n3408),.clk(gclk));
	jand g03191(.dina(n3408),.dinb(w_asqrt42_39[0]),.dout(n3409),.clk(gclk));
	jxor g03192(.dina(n3409),.dinb(w_n3122_0[0]),.dout(n3410),.clk(gclk));
	jnot g03193(.din(w_n3410_0[1]),.dout(n3411),.clk(gclk));
	jand g03194(.dina(w_n3411_0[1]),.dinb(n3407),.dout(n3412),.clk(gclk));
	jor g03195(.dina(n3412),.dinb(w_n3406_0[1]),.dout(n3413),.clk(gclk));
	jand g03196(.dina(w_n3413_0[2]),.dinb(w_asqrt49_32[2]),.dout(n3414),.clk(gclk));
	jor g03197(.dina(w_n3413_0[1]),.dinb(w_asqrt49_32[1]),.dout(n3415),.clk(gclk));
	jxor g03198(.dina(w_n3124_0[0]),.dinb(w_n1912_54[2]),.dout(n3416),.clk(gclk));
	jand g03199(.dina(n3416),.dinb(w_asqrt42_38[2]),.dout(n3417),.clk(gclk));
	jxor g03200(.dina(n3417),.dinb(w_n3129_0[0]),.dout(n3418),.clk(gclk));
	jand g03201(.dina(w_n3418_0[1]),.dinb(n3415),.dout(n3419),.clk(gclk));
	jor g03202(.dina(n3419),.dinb(w_n3414_0[1]),.dout(n3420),.clk(gclk));
	jand g03203(.dina(w_n3420_0[2]),.dinb(w_asqrt50_34[2]),.dout(n3421),.clk(gclk));
	jor g03204(.dina(w_n3420_0[1]),.dinb(w_asqrt50_34[1]),.dout(n3422),.clk(gclk));
	jxor g03205(.dina(w_n3132_0[0]),.dinb(w_n1699_57[0]),.dout(n3423),.clk(gclk));
	jand g03206(.dina(n3423),.dinb(w_asqrt42_38[1]),.dout(n3424),.clk(gclk));
	jxor g03207(.dina(n3424),.dinb(w_n3137_0[0]),.dout(n3425),.clk(gclk));
	jnot g03208(.din(w_n3425_0[1]),.dout(n3426),.clk(gclk));
	jand g03209(.dina(w_n3426_0[1]),.dinb(n3422),.dout(n3427),.clk(gclk));
	jor g03210(.dina(n3427),.dinb(w_n3421_0[1]),.dout(n3428),.clk(gclk));
	jand g03211(.dina(w_n3428_0[2]),.dinb(w_asqrt51_33[0]),.dout(n3429),.clk(gclk));
	jor g03212(.dina(w_n3428_0[1]),.dinb(w_asqrt51_32[2]),.dout(n3430),.clk(gclk));
	jxor g03213(.dina(w_n3139_0[0]),.dinb(w_n1516_55[1]),.dout(n3431),.clk(gclk));
	jand g03214(.dina(n3431),.dinb(w_asqrt42_38[0]),.dout(n3432),.clk(gclk));
	jxor g03215(.dina(n3432),.dinb(w_n3144_0[0]),.dout(n3433),.clk(gclk));
	jand g03216(.dina(w_n3433_0[1]),.dinb(n3430),.dout(n3434),.clk(gclk));
	jor g03217(.dina(n3434),.dinb(w_n3429_0[1]),.dout(n3435),.clk(gclk));
	jand g03218(.dina(w_n3435_0[2]),.dinb(w_asqrt52_34[2]),.dout(n3436),.clk(gclk));
	jor g03219(.dina(w_n3435_0[1]),.dinb(w_asqrt52_34[1]),.dout(n3437),.clk(gclk));
	jxor g03220(.dina(w_n3147_0[0]),.dinb(w_n1332_57[0]),.dout(n3438),.clk(gclk));
	jand g03221(.dina(n3438),.dinb(w_asqrt42_37[2]),.dout(n3439),.clk(gclk));
	jxor g03222(.dina(n3439),.dinb(w_n3152_0[0]),.dout(n3440),.clk(gclk));
	jnot g03223(.din(w_n3440_0[1]),.dout(n3441),.clk(gclk));
	jand g03224(.dina(w_n3441_0[1]),.dinb(n3437),.dout(n3442),.clk(gclk));
	jor g03225(.dina(n3442),.dinb(w_n3436_0[1]),.dout(n3443),.clk(gclk));
	jand g03226(.dina(w_n3443_0[2]),.dinb(w_asqrt53_33[2]),.dout(n3444),.clk(gclk));
	jor g03227(.dina(w_n3443_0[1]),.dinb(w_asqrt53_33[1]),.dout(n3445),.clk(gclk));
	jxor g03228(.dina(w_n3154_0[0]),.dinb(w_n1173_56[0]),.dout(n3446),.clk(gclk));
	jand g03229(.dina(n3446),.dinb(w_asqrt42_37[1]),.dout(n3447),.clk(gclk));
	jxor g03230(.dina(n3447),.dinb(w_n3159_0[0]),.dout(n3448),.clk(gclk));
	jand g03231(.dina(w_n3448_0[1]),.dinb(n3445),.dout(n3449),.clk(gclk));
	jor g03232(.dina(n3449),.dinb(w_n3444_0[1]),.dout(n3450),.clk(gclk));
	jand g03233(.dina(w_n3450_0[2]),.dinb(w_asqrt54_34[2]),.dout(n3451),.clk(gclk));
	jor g03234(.dina(w_n3450_0[1]),.dinb(w_asqrt54_34[1]),.dout(n3452),.clk(gclk));
	jxor g03235(.dina(w_n3162_0[0]),.dinb(w_n1008_58[0]),.dout(n3453),.clk(gclk));
	jand g03236(.dina(n3453),.dinb(w_asqrt42_37[0]),.dout(n3454),.clk(gclk));
	jxor g03237(.dina(n3454),.dinb(w_n3167_0[0]),.dout(n3455),.clk(gclk));
	jnot g03238(.din(w_n3455_0[1]),.dout(n3456),.clk(gclk));
	jand g03239(.dina(w_n3456_0[1]),.dinb(n3452),.dout(n3457),.clk(gclk));
	jor g03240(.dina(n3457),.dinb(w_n3451_0[1]),.dout(n3458),.clk(gclk));
	jand g03241(.dina(w_n3458_0[2]),.dinb(w_asqrt55_34[0]),.dout(n3459),.clk(gclk));
	jor g03242(.dina(w_n3458_0[1]),.dinb(w_asqrt55_33[2]),.dout(n3460),.clk(gclk));
	jxor g03243(.dina(w_n3169_0[0]),.dinb(w_n884_57[0]),.dout(n3461),.clk(gclk));
	jand g03244(.dina(n3461),.dinb(w_asqrt42_36[2]),.dout(n3462),.clk(gclk));
	jxor g03245(.dina(n3462),.dinb(w_n3174_0[0]),.dout(n3463),.clk(gclk));
	jand g03246(.dina(w_n3463_0[1]),.dinb(n3460),.dout(n3464),.clk(gclk));
	jor g03247(.dina(n3464),.dinb(w_n3459_0[1]),.dout(n3465),.clk(gclk));
	jand g03248(.dina(w_n3465_0[2]),.dinb(w_asqrt56_35[0]),.dout(n3466),.clk(gclk));
	jor g03249(.dina(w_n3465_0[1]),.dinb(w_asqrt56_34[2]),.dout(n3467),.clk(gclk));
	jxor g03250(.dina(w_n3177_0[0]),.dinb(w_n743_58[0]),.dout(n3468),.clk(gclk));
	jand g03251(.dina(n3468),.dinb(w_asqrt42_36[1]),.dout(n3469),.clk(gclk));
	jxor g03252(.dina(n3469),.dinb(w_n3182_0[0]),.dout(n3470),.clk(gclk));
	jnot g03253(.din(w_n3470_0[1]),.dout(n3471),.clk(gclk));
	jand g03254(.dina(w_n3471_0[1]),.dinb(n3467),.dout(n3472),.clk(gclk));
	jor g03255(.dina(n3472),.dinb(w_n3466_0[1]),.dout(n3473),.clk(gclk));
	jand g03256(.dina(w_n3473_0[2]),.dinb(w_asqrt57_34[2]),.dout(n3474),.clk(gclk));
	jor g03257(.dina(w_n3473_0[1]),.dinb(w_asqrt57_34[1]),.dout(n3475),.clk(gclk));
	jxor g03258(.dina(w_n3184_0[0]),.dinb(w_n635_58[0]),.dout(n3476),.clk(gclk));
	jand g03259(.dina(n3476),.dinb(w_asqrt42_36[0]),.dout(n3477),.clk(gclk));
	jxor g03260(.dina(n3477),.dinb(w_n3189_0[0]),.dout(n3478),.clk(gclk));
	jand g03261(.dina(w_n3478_0[1]),.dinb(n3475),.dout(n3479),.clk(gclk));
	jor g03262(.dina(n3479),.dinb(w_n3474_0[1]),.dout(n3480),.clk(gclk));
	jand g03263(.dina(w_n3480_0[2]),.dinb(w_asqrt58_35[1]),.dout(n3481),.clk(gclk));
	jor g03264(.dina(w_n3480_0[1]),.dinb(w_asqrt58_35[0]),.dout(n3482),.clk(gclk));
	jxor g03265(.dina(w_n3192_0[0]),.dinb(w_n515_59[0]),.dout(n3483),.clk(gclk));
	jand g03266(.dina(n3483),.dinb(w_asqrt42_35[2]),.dout(n3484),.clk(gclk));
	jxor g03267(.dina(n3484),.dinb(w_n3197_0[0]),.dout(n3485),.clk(gclk));
	jnot g03268(.din(w_n3485_0[1]),.dout(n3486),.clk(gclk));
	jand g03269(.dina(w_n3486_0[1]),.dinb(n3482),.dout(n3487),.clk(gclk));
	jor g03270(.dina(n3487),.dinb(w_n3481_0[1]),.dout(n3488),.clk(gclk));
	jand g03271(.dina(w_n3488_0[2]),.dinb(w_asqrt59_35[0]),.dout(n3489),.clk(gclk));
	jor g03272(.dina(w_n3488_0[1]),.dinb(w_asqrt59_34[2]),.dout(n3490),.clk(gclk));
	jxor g03273(.dina(w_n3199_0[0]),.dinb(w_n443_59[0]),.dout(n3491),.clk(gclk));
	jand g03274(.dina(n3491),.dinb(w_asqrt42_35[1]),.dout(n3492),.clk(gclk));
	jxor g03275(.dina(n3492),.dinb(w_n3204_0[0]),.dout(n3493),.clk(gclk));
	jnot g03276(.din(w_n3493_0[1]),.dout(n3494),.clk(gclk));
	jand g03277(.dina(w_n3494_0[1]),.dinb(n3490),.dout(n3495),.clk(gclk));
	jor g03278(.dina(n3495),.dinb(w_n3489_0[1]),.dout(n3496),.clk(gclk));
	jand g03279(.dina(w_n3496_0[2]),.dinb(w_asqrt60_35[1]),.dout(n3497),.clk(gclk));
	jor g03280(.dina(w_n3496_0[1]),.dinb(w_asqrt60_35[0]),.dout(n3498),.clk(gclk));
	jxor g03281(.dina(w_n3206_0[0]),.dinb(w_n352_59[1]),.dout(n3499),.clk(gclk));
	jand g03282(.dina(n3499),.dinb(w_asqrt42_35[0]),.dout(n3500),.clk(gclk));
	jxor g03283(.dina(n3500),.dinb(w_n3211_0[0]),.dout(n3501),.clk(gclk));
	jand g03284(.dina(w_n3501_0[1]),.dinb(n3498),.dout(n3502),.clk(gclk));
	jor g03285(.dina(n3502),.dinb(w_n3497_0[1]),.dout(n3503),.clk(gclk));
	jand g03286(.dina(w_n3503_0[2]),.dinb(w_asqrt61_35[1]),.dout(n3504),.clk(gclk));
	jor g03287(.dina(w_n3503_0[1]),.dinb(w_asqrt61_35[0]),.dout(n3505),.clk(gclk));
	jxor g03288(.dina(w_n3214_0[0]),.dinb(w_n294_59[2]),.dout(n3506),.clk(gclk));
	jand g03289(.dina(n3506),.dinb(w_asqrt42_34[2]),.dout(n3507),.clk(gclk));
	jxor g03290(.dina(n3507),.dinb(w_n3219_0[0]),.dout(n3508),.clk(gclk));
	jand g03291(.dina(w_n3508_0[1]),.dinb(n3505),.dout(n3509),.clk(gclk));
	jor g03292(.dina(n3509),.dinb(w_n3504_0[1]),.dout(n3510),.clk(gclk));
	jand g03293(.dina(w_n3510_0[2]),.dinb(w_asqrt62_35[1]),.dout(n3511),.clk(gclk));
	jor g03294(.dina(w_n3510_0[1]),.dinb(w_asqrt62_35[0]),.dout(n3512),.clk(gclk));
	jxor g03295(.dina(w_n3222_0[0]),.dinb(w_n239_59[2]),.dout(n3513),.clk(gclk));
	jand g03296(.dina(n3513),.dinb(w_asqrt42_34[1]),.dout(n3514),.clk(gclk));
	jxor g03297(.dina(n3514),.dinb(w_n3227_0[0]),.dout(n3515),.clk(gclk));
	jnot g03298(.din(w_n3515_0[2]),.dout(n3516),.clk(gclk));
	jand g03299(.dina(n3516),.dinb(n3512),.dout(n3517),.clk(gclk));
	jor g03300(.dina(n3517),.dinb(w_n3511_0[1]),.dout(n3518),.clk(gclk));
	jxor g03301(.dina(w_n3229_0[0]),.dinb(w_n221_60[0]),.dout(n3519),.clk(gclk));
	jand g03302(.dina(n3519),.dinb(w_asqrt42_34[0]),.dout(n3520),.clk(gclk));
	jxor g03303(.dina(n3520),.dinb(w_n3235_0[0]),.dout(n3521),.clk(gclk));
	jnot g03304(.din(w_n3521_0[2]),.dout(n3522),.clk(gclk));
	jor g03305(.dina(w_n3522_0[1]),.dinb(w_n3518_0[1]),.dout(n3523),.clk(gclk));
	jnot g03306(.din(w_n3523_1[1]),.dout(n3524),.clk(gclk));
	jnot g03307(.din(w_n3511_0[0]),.dout(n3526),.clk(gclk));
	jnot g03308(.din(w_n3504_0[0]),.dout(n3527),.clk(gclk));
	jnot g03309(.din(w_n3497_0[0]),.dout(n3528),.clk(gclk));
	jnot g03310(.din(w_n3489_0[0]),.dout(n3529),.clk(gclk));
	jnot g03311(.din(w_n3481_0[0]),.dout(n3530),.clk(gclk));
	jnot g03312(.din(w_n3474_0[0]),.dout(n3531),.clk(gclk));
	jnot g03313(.din(w_n3466_0[0]),.dout(n3532),.clk(gclk));
	jnot g03314(.din(w_n3459_0[0]),.dout(n3533),.clk(gclk));
	jnot g03315(.din(w_n3451_0[0]),.dout(n3534),.clk(gclk));
	jnot g03316(.din(w_n3444_0[0]),.dout(n3535),.clk(gclk));
	jnot g03317(.din(w_n3436_0[0]),.dout(n3536),.clk(gclk));
	jnot g03318(.din(w_n3429_0[0]),.dout(n3537),.clk(gclk));
	jnot g03319(.din(w_n3421_0[0]),.dout(n3538),.clk(gclk));
	jnot g03320(.din(w_n3414_0[0]),.dout(n3539),.clk(gclk));
	jnot g03321(.din(w_n3406_0[0]),.dout(n3540),.clk(gclk));
	jnot g03322(.din(w_n3398_0[0]),.dout(n3541),.clk(gclk));
	jnot g03323(.din(w_n3391_0[0]),.dout(n3542),.clk(gclk));
	jnot g03324(.din(w_n3384_0[0]),.dout(n3543),.clk(gclk));
	jnot g03325(.din(w_n3373_0[0]),.dout(n3544),.clk(gclk));
	jnot g03326(.din(w_n3263_0[0]),.dout(n3545),.clk(gclk));
	jor g03327(.dina(w_n3368_52[0]),.dinb(w_n3075_0[2]),.dout(n3546),.clk(gclk));
	jnot g03328(.din(w_n3261_0[0]),.dout(n3547),.clk(gclk));
	jand g03329(.dina(n3547),.dinb(n3546),.dout(n3548),.clk(gclk));
	jand g03330(.dina(n3548),.dinb(w_n3089_55[0]),.dout(n3549),.clk(gclk));
	jor g03331(.dina(w_n3368_51[2]),.dinb(w_a84_0[0]),.dout(n3550),.clk(gclk));
	jand g03332(.dina(n3550),.dinb(w_a85_0[0]),.dout(n3551),.clk(gclk));
	jor g03333(.dina(w_n3375_0[0]),.dinb(n3551),.dout(n3552),.clk(gclk));
	jor g03334(.dina(w_n3552_0[1]),.dinb(n3549),.dout(n3553),.clk(gclk));
	jand g03335(.dina(n3553),.dinb(n3545),.dout(n3554),.clk(gclk));
	jand g03336(.dina(n3554),.dinb(w_n2833_52[2]),.dout(n3555),.clk(gclk));
	jor g03337(.dina(w_n3380_0[0]),.dinb(n3555),.dout(n3556),.clk(gclk));
	jand g03338(.dina(n3556),.dinb(n3544),.dout(n3557),.clk(gclk));
	jand g03339(.dina(n3557),.dinb(w_n2572_55[1]),.dout(n3558),.clk(gclk));
	jnot g03340(.din(w_n3388_0[0]),.dout(n3559),.clk(gclk));
	jor g03341(.dina(w_n3559_0[1]),.dinb(n3558),.dout(n3560),.clk(gclk));
	jand g03342(.dina(n3560),.dinb(n3543),.dout(n3561),.clk(gclk));
	jand g03343(.dina(n3561),.dinb(w_n2345_53[1]),.dout(n3562),.clk(gclk));
	jnot g03344(.din(w_n3395_0[0]),.dout(n3563),.clk(gclk));
	jor g03345(.dina(w_n3563_0[1]),.dinb(n3562),.dout(n3564),.clk(gclk));
	jand g03346(.dina(n3564),.dinb(n3542),.dout(n3565),.clk(gclk));
	jand g03347(.dina(n3565),.dinb(w_n2108_56[0]),.dout(n3566),.clk(gclk));
	jor g03348(.dina(w_n3402_0[0]),.dinb(n3566),.dout(n3567),.clk(gclk));
	jand g03349(.dina(n3567),.dinb(n3541),.dout(n3568),.clk(gclk));
	jand g03350(.dina(n3568),.dinb(w_n1912_54[1]),.dout(n3569),.clk(gclk));
	jor g03351(.dina(w_n3410_0[0]),.dinb(n3569),.dout(n3570),.clk(gclk));
	jand g03352(.dina(n3570),.dinb(n3540),.dout(n3571),.clk(gclk));
	jand g03353(.dina(n3571),.dinb(w_n1699_56[2]),.dout(n3572),.clk(gclk));
	jnot g03354(.din(w_n3418_0[0]),.dout(n3573),.clk(gclk));
	jor g03355(.dina(w_n3573_0[1]),.dinb(n3572),.dout(n3574),.clk(gclk));
	jand g03356(.dina(n3574),.dinb(n3539),.dout(n3575),.clk(gclk));
	jand g03357(.dina(n3575),.dinb(w_n1516_55[0]),.dout(n3576),.clk(gclk));
	jor g03358(.dina(w_n3425_0[0]),.dinb(n3576),.dout(n3577),.clk(gclk));
	jand g03359(.dina(n3577),.dinb(n3538),.dout(n3578),.clk(gclk));
	jand g03360(.dina(n3578),.dinb(w_n1332_56[2]),.dout(n3579),.clk(gclk));
	jnot g03361(.din(w_n3433_0[0]),.dout(n3580),.clk(gclk));
	jor g03362(.dina(w_n3580_0[1]),.dinb(n3579),.dout(n3581),.clk(gclk));
	jand g03363(.dina(n3581),.dinb(n3537),.dout(n3582),.clk(gclk));
	jand g03364(.dina(n3582),.dinb(w_n1173_55[2]),.dout(n3583),.clk(gclk));
	jor g03365(.dina(w_n3440_0[0]),.dinb(n3583),.dout(n3584),.clk(gclk));
	jand g03366(.dina(n3584),.dinb(n3536),.dout(n3585),.clk(gclk));
	jand g03367(.dina(n3585),.dinb(w_n1008_57[2]),.dout(n3586),.clk(gclk));
	jnot g03368(.din(w_n3448_0[0]),.dout(n3587),.clk(gclk));
	jor g03369(.dina(w_n3587_0[1]),.dinb(n3586),.dout(n3588),.clk(gclk));
	jand g03370(.dina(n3588),.dinb(n3535),.dout(n3589),.clk(gclk));
	jand g03371(.dina(n3589),.dinb(w_n884_56[2]),.dout(n3590),.clk(gclk));
	jor g03372(.dina(w_n3455_0[0]),.dinb(n3590),.dout(n3591),.clk(gclk));
	jand g03373(.dina(n3591),.dinb(n3534),.dout(n3592),.clk(gclk));
	jand g03374(.dina(n3592),.dinb(w_n743_57[2]),.dout(n3593),.clk(gclk));
	jnot g03375(.din(w_n3463_0[0]),.dout(n3594),.clk(gclk));
	jor g03376(.dina(w_n3594_0[1]),.dinb(n3593),.dout(n3595),.clk(gclk));
	jand g03377(.dina(n3595),.dinb(n3533),.dout(n3596),.clk(gclk));
	jand g03378(.dina(n3596),.dinb(w_n635_57[2]),.dout(n3597),.clk(gclk));
	jor g03379(.dina(w_n3470_0[0]),.dinb(n3597),.dout(n3598),.clk(gclk));
	jand g03380(.dina(n3598),.dinb(n3532),.dout(n3599),.clk(gclk));
	jand g03381(.dina(n3599),.dinb(w_n515_58[2]),.dout(n3600),.clk(gclk));
	jnot g03382(.din(w_n3478_0[0]),.dout(n3601),.clk(gclk));
	jor g03383(.dina(w_n3601_0[1]),.dinb(n3600),.dout(n3602),.clk(gclk));
	jand g03384(.dina(n3602),.dinb(n3531),.dout(n3603),.clk(gclk));
	jand g03385(.dina(n3603),.dinb(w_n443_58[2]),.dout(n3604),.clk(gclk));
	jor g03386(.dina(w_n3485_0[0]),.dinb(n3604),.dout(n3605),.clk(gclk));
	jand g03387(.dina(n3605),.dinb(n3530),.dout(n3606),.clk(gclk));
	jand g03388(.dina(n3606),.dinb(w_n352_59[0]),.dout(n3607),.clk(gclk));
	jor g03389(.dina(w_n3493_0[0]),.dinb(n3607),.dout(n3608),.clk(gclk));
	jand g03390(.dina(n3608),.dinb(n3529),.dout(n3609),.clk(gclk));
	jand g03391(.dina(n3609),.dinb(w_n294_59[1]),.dout(n3610),.clk(gclk));
	jnot g03392(.din(w_n3501_0[0]),.dout(n3611),.clk(gclk));
	jor g03393(.dina(w_n3611_0[1]),.dinb(n3610),.dout(n3612),.clk(gclk));
	jand g03394(.dina(n3612),.dinb(n3528),.dout(n3613),.clk(gclk));
	jand g03395(.dina(n3613),.dinb(w_n239_59[1]),.dout(n3614),.clk(gclk));
	jnot g03396(.din(w_n3508_0[0]),.dout(n3615),.clk(gclk));
	jor g03397(.dina(w_n3615_0[1]),.dinb(n3614),.dout(n3616),.clk(gclk));
	jand g03398(.dina(n3616),.dinb(n3527),.dout(n3617),.clk(gclk));
	jand g03399(.dina(n3617),.dinb(w_n221_59[2]),.dout(n3618),.clk(gclk));
	jor g03400(.dina(w_n3515_0[1]),.dinb(n3618),.dout(n3619),.clk(gclk));
	jand g03401(.dina(n3619),.dinb(n3526),.dout(n3620),.clk(gclk));
	jor g03402(.dina(w_n3521_0[1]),.dinb(w_n3620_0[1]),.dout(n3621),.clk(gclk));
	jxor g03403(.dina(w_n3240_0[1]),.dinb(w_n3237_0[2]),.dout(n3622),.clk(gclk));
	jnot g03404(.din(w_n3622_0[1]),.dout(n3623),.clk(gclk));
	jand g03405(.dina(n3623),.dinb(w_asqrt42_33[2]),.dout(n3624),.clk(gclk));
	jor g03406(.dina(w_n3624_0[1]),.dinb(w_n3621_0[1]),.dout(n3625),.clk(gclk));
	jand g03407(.dina(n3625),.dinb(w_n218_24[2]),.dout(n3626),.clk(gclk));
	jand g03408(.dina(w_n3367_0[0]),.dinb(w_n3237_0[1]),.dout(n3627),.clk(gclk));
	jnot g03409(.din(n3627),.dout(n3628),.clk(gclk));
	jand g03410(.dina(w_n3622_0[0]),.dinb(w_asqrt63_45[1]),.dout(n3629),.clk(gclk));
	jand g03411(.dina(w_n3629_0[1]),.dinb(n3628),.dout(n3630),.clk(gclk));
	jor g03412(.dina(w_n3630_0[1]),.dinb(w_n3626_0[1]),.dout(n3631),.clk(gclk));
	jor g03413(.dina(w_n3631_0[1]),.dinb(w_n3524_0[2]),.dout(asqrt_fa_42),.clk(gclk));
	jand g03414(.dina(w_n3522_0[0]),.dinb(w_n3518_0[0]),.dout(n3635),.clk(gclk));
	jnot g03415(.din(w_n3624_0[0]),.dout(n3636),.clk(gclk));
	jand g03416(.dina(n3636),.dinb(w_n3635_0[1]),.dout(n3637),.clk(gclk));
	jor g03417(.dina(n3637),.dinb(w_asqrt63_45[0]),.dout(n3638),.clk(gclk));
	jnot g03418(.din(w_n3630_0[0]),.dout(n3639),.clk(gclk));
	jand g03419(.dina(n3639),.dinb(n3638),.dout(n3640),.clk(gclk));
	jand g03420(.dina(w_n3640_0[1]),.dinb(w_n3523_1[0]),.dout(n3642),.clk(gclk));
	jxor g03421(.dina(w_n3510_0[0]),.dinb(w_n221_59[1]),.dout(n3643),.clk(gclk));
	jor g03422(.dina(n3643),.dinb(w_n3642_60[2]),.dout(n3644),.clk(gclk));
	jxor g03423(.dina(n3644),.dinb(w_n3515_0[0]),.dout(n3645),.clk(gclk));
	jnot g03424(.din(w_n3645_0[1]),.dout(n3646),.clk(gclk));
	jor g03425(.dina(w_n3642_60[1]),.dinb(w_n3258_1[0]),.dout(n3647),.clk(gclk));
	jnot g03426(.din(w_a80_0[2]),.dout(n3648),.clk(gclk));
	jnot g03427(.din(w_a81_0[1]),.dout(n3649),.clk(gclk));
	jand g03428(.dina(w_n3649_0[1]),.dinb(w_n3648_1[2]),.dout(n3650),.clk(gclk));
	jand g03429(.dina(w_n3650_0[2]),.dinb(w_n3258_0[2]),.dout(n3651),.clk(gclk));
	jnot g03430(.din(w_n3651_0[1]),.dout(n3652),.clk(gclk));
	jand g03431(.dina(n3652),.dinb(n3647),.dout(n3653),.clk(gclk));
	jor g03432(.dina(w_n3653_0[2]),.dinb(w_n3368_51[1]),.dout(n3654),.clk(gclk));
	jand g03433(.dina(w_n3653_0[1]),.dinb(w_n3368_51[0]),.dout(n3655),.clk(gclk));
	jor g03434(.dina(w_n3642_60[0]),.dinb(w_a82_1[0]),.dout(n3656),.clk(gclk));
	jand g03435(.dina(n3656),.dinb(w_a83_0[0]),.dout(n3657),.clk(gclk));
	jand g03436(.dina(w_asqrt41_31),.dinb(w_n3260_0[1]),.dout(n3658),.clk(gclk));
	jor g03437(.dina(n3658),.dinb(n3657),.dout(n3659),.clk(gclk));
	jor g03438(.dina(n3659),.dinb(n3655),.dout(n3660),.clk(gclk));
	jand g03439(.dina(n3660),.dinb(w_n3654_0[1]),.dout(n3661),.clk(gclk));
	jor g03440(.dina(w_n3661_0[2]),.dinb(w_n3089_54[2]),.dout(n3662),.clk(gclk));
	jand g03441(.dina(w_n3661_0[1]),.dinb(w_n3089_54[1]),.dout(n3663),.clk(gclk));
	jnot g03442(.din(w_n3260_0[0]),.dout(n3664),.clk(gclk));
	jor g03443(.dina(w_n3642_59[2]),.dinb(n3664),.dout(n3665),.clk(gclk));
	jor g03444(.dina(w_n3629_0[0]),.dinb(w_n3524_0[1]),.dout(n3666),.clk(gclk));
	jor g03445(.dina(n3666),.dinb(w_n3626_0[0]),.dout(n3667),.clk(gclk));
	jor g03446(.dina(n3667),.dinb(w_n3368_50[2]),.dout(n3668),.clk(gclk));
	jand g03447(.dina(n3668),.dinb(w_n3665_0[1]),.dout(n3669),.clk(gclk));
	jxor g03448(.dina(n3669),.dinb(w_n3075_0[1]),.dout(n3670),.clk(gclk));
	jor g03449(.dina(w_n3670_0[2]),.dinb(n3663),.dout(n3671),.clk(gclk));
	jand g03450(.dina(n3671),.dinb(w_n3662_0[1]),.dout(n3672),.clk(gclk));
	jor g03451(.dina(w_n3672_0[2]),.dinb(w_n2833_52[1]),.dout(n3673),.clk(gclk));
	jand g03452(.dina(w_n3672_0[1]),.dinb(w_n2833_52[0]),.dout(n3674),.clk(gclk));
	jxor g03453(.dina(w_n3262_0[0]),.dinb(w_n3089_54[0]),.dout(n3675),.clk(gclk));
	jor g03454(.dina(n3675),.dinb(w_n3642_59[1]),.dout(n3676),.clk(gclk));
	jxor g03455(.dina(n3676),.dinb(w_n3552_0[0]),.dout(n3677),.clk(gclk));
	jnot g03456(.din(w_n3677_0[2]),.dout(n3678),.clk(gclk));
	jor g03457(.dina(n3678),.dinb(n3674),.dout(n3679),.clk(gclk));
	jand g03458(.dina(n3679),.dinb(w_n3673_0[1]),.dout(n3680),.clk(gclk));
	jor g03459(.dina(w_n3680_0[2]),.dinb(w_n2572_55[0]),.dout(n3681),.clk(gclk));
	jand g03460(.dina(w_n3680_0[1]),.dinb(w_n2572_54[2]),.dout(n3682),.clk(gclk));
	jxor g03461(.dina(w_n3372_0[0]),.dinb(w_n2833_51[2]),.dout(n3683),.clk(gclk));
	jor g03462(.dina(n3683),.dinb(w_n3642_59[0]),.dout(n3684),.clk(gclk));
	jxor g03463(.dina(n3684),.dinb(w_n3381_0[0]),.dout(n3685),.clk(gclk));
	jor g03464(.dina(w_n3685_0[2]),.dinb(n3682),.dout(n3686),.clk(gclk));
	jand g03465(.dina(n3686),.dinb(w_n3681_0[1]),.dout(n3687),.clk(gclk));
	jor g03466(.dina(w_n3687_0[2]),.dinb(w_n2345_53[0]),.dout(n3688),.clk(gclk));
	jand g03467(.dina(w_n3687_0[1]),.dinb(w_n2345_52[2]),.dout(n3689),.clk(gclk));
	jxor g03468(.dina(w_n3383_0[0]),.dinb(w_n2572_54[1]),.dout(n3690),.clk(gclk));
	jor g03469(.dina(n3690),.dinb(w_n3642_58[2]),.dout(n3691),.clk(gclk));
	jxor g03470(.dina(n3691),.dinb(w_n3559_0[0]),.dout(n3692),.clk(gclk));
	jnot g03471(.din(w_n3692_0[2]),.dout(n3693),.clk(gclk));
	jor g03472(.dina(n3693),.dinb(n3689),.dout(n3694),.clk(gclk));
	jand g03473(.dina(n3694),.dinb(w_n3688_0[1]),.dout(n3695),.clk(gclk));
	jor g03474(.dina(w_n3695_0[2]),.dinb(w_n2108_55[2]),.dout(n3696),.clk(gclk));
	jand g03475(.dina(w_n3695_0[1]),.dinb(w_n2108_55[1]),.dout(n3697),.clk(gclk));
	jxor g03476(.dina(w_n3390_0[0]),.dinb(w_n2345_52[1]),.dout(n3698),.clk(gclk));
	jor g03477(.dina(n3698),.dinb(w_n3642_58[1]),.dout(n3699),.clk(gclk));
	jxor g03478(.dina(n3699),.dinb(w_n3563_0[0]),.dout(n3700),.clk(gclk));
	jnot g03479(.din(w_n3700_0[2]),.dout(n3701),.clk(gclk));
	jor g03480(.dina(n3701),.dinb(n3697),.dout(n3702),.clk(gclk));
	jand g03481(.dina(n3702),.dinb(w_n3696_0[1]),.dout(n3703),.clk(gclk));
	jor g03482(.dina(w_n3703_0[2]),.dinb(w_n1912_54[0]),.dout(n3704),.clk(gclk));
	jand g03483(.dina(w_n3703_0[1]),.dinb(w_n1912_53[2]),.dout(n3705),.clk(gclk));
	jxor g03484(.dina(w_n3397_0[0]),.dinb(w_n2108_55[0]),.dout(n3706),.clk(gclk));
	jor g03485(.dina(n3706),.dinb(w_n3642_58[0]),.dout(n3707),.clk(gclk));
	jxor g03486(.dina(n3707),.dinb(w_n3403_0[0]),.dout(n3708),.clk(gclk));
	jor g03487(.dina(w_n3708_0[2]),.dinb(n3705),.dout(n3709),.clk(gclk));
	jand g03488(.dina(n3709),.dinb(w_n3704_0[1]),.dout(n3710),.clk(gclk));
	jor g03489(.dina(w_n3710_0[2]),.dinb(w_n1699_56[1]),.dout(n3711),.clk(gclk));
	jand g03490(.dina(w_n3710_0[1]),.dinb(w_n1699_56[0]),.dout(n3712),.clk(gclk));
	jxor g03491(.dina(w_n3405_0[0]),.dinb(w_n1912_53[1]),.dout(n3713),.clk(gclk));
	jor g03492(.dina(n3713),.dinb(w_n3642_57[2]),.dout(n3714),.clk(gclk));
	jxor g03493(.dina(n3714),.dinb(w_n3411_0[0]),.dout(n3715),.clk(gclk));
	jor g03494(.dina(w_n3715_0[2]),.dinb(n3712),.dout(n3716),.clk(gclk));
	jand g03495(.dina(n3716),.dinb(w_n3711_0[1]),.dout(n3717),.clk(gclk));
	jor g03496(.dina(w_n3717_0[2]),.dinb(w_n1516_54[2]),.dout(n3718),.clk(gclk));
	jand g03497(.dina(w_n3717_0[1]),.dinb(w_n1516_54[1]),.dout(n3719),.clk(gclk));
	jxor g03498(.dina(w_n3413_0[0]),.dinb(w_n1699_55[2]),.dout(n3720),.clk(gclk));
	jor g03499(.dina(n3720),.dinb(w_n3642_57[1]),.dout(n3721),.clk(gclk));
	jxor g03500(.dina(n3721),.dinb(w_n3573_0[0]),.dout(n3722),.clk(gclk));
	jnot g03501(.din(w_n3722_0[2]),.dout(n3723),.clk(gclk));
	jor g03502(.dina(n3723),.dinb(n3719),.dout(n3724),.clk(gclk));
	jand g03503(.dina(n3724),.dinb(w_n3718_0[1]),.dout(n3725),.clk(gclk));
	jor g03504(.dina(w_n3725_0[2]),.dinb(w_n1332_56[1]),.dout(n3726),.clk(gclk));
	jand g03505(.dina(w_n3725_0[1]),.dinb(w_n1332_56[0]),.dout(n3727),.clk(gclk));
	jxor g03506(.dina(w_n3420_0[0]),.dinb(w_n1516_54[0]),.dout(n3728),.clk(gclk));
	jor g03507(.dina(n3728),.dinb(w_n3642_57[0]),.dout(n3729),.clk(gclk));
	jxor g03508(.dina(n3729),.dinb(w_n3426_0[0]),.dout(n3730),.clk(gclk));
	jor g03509(.dina(w_n3730_0[2]),.dinb(n3727),.dout(n3731),.clk(gclk));
	jand g03510(.dina(n3731),.dinb(w_n3726_0[1]),.dout(n3732),.clk(gclk));
	jor g03511(.dina(w_n3732_0[2]),.dinb(w_n1173_55[1]),.dout(n3733),.clk(gclk));
	jand g03512(.dina(w_n3732_0[1]),.dinb(w_n1173_55[0]),.dout(n3734),.clk(gclk));
	jxor g03513(.dina(w_n3428_0[0]),.dinb(w_n1332_55[2]),.dout(n3735),.clk(gclk));
	jor g03514(.dina(n3735),.dinb(w_n3642_56[2]),.dout(n3736),.clk(gclk));
	jxor g03515(.dina(n3736),.dinb(w_n3580_0[0]),.dout(n3737),.clk(gclk));
	jnot g03516(.din(w_n3737_0[2]),.dout(n3738),.clk(gclk));
	jor g03517(.dina(n3738),.dinb(n3734),.dout(n3739),.clk(gclk));
	jand g03518(.dina(n3739),.dinb(w_n3733_0[1]),.dout(n3740),.clk(gclk));
	jor g03519(.dina(w_n3740_0[2]),.dinb(w_n1008_57[1]),.dout(n3741),.clk(gclk));
	jand g03520(.dina(w_n3740_0[1]),.dinb(w_n1008_57[0]),.dout(n3742),.clk(gclk));
	jxor g03521(.dina(w_n3435_0[0]),.dinb(w_n1173_54[2]),.dout(n3743),.clk(gclk));
	jor g03522(.dina(n3743),.dinb(w_n3642_56[1]),.dout(n3744),.clk(gclk));
	jxor g03523(.dina(n3744),.dinb(w_n3441_0[0]),.dout(n3745),.clk(gclk));
	jor g03524(.dina(w_n3745_0[2]),.dinb(n3742),.dout(n3746),.clk(gclk));
	jand g03525(.dina(n3746),.dinb(w_n3741_0[1]),.dout(n3747),.clk(gclk));
	jor g03526(.dina(w_n3747_0[2]),.dinb(w_n884_56[1]),.dout(n3748),.clk(gclk));
	jand g03527(.dina(w_n3747_0[1]),.dinb(w_n884_56[0]),.dout(n3749),.clk(gclk));
	jxor g03528(.dina(w_n3443_0[0]),.dinb(w_n1008_56[2]),.dout(n3750),.clk(gclk));
	jor g03529(.dina(n3750),.dinb(w_n3642_56[0]),.dout(n3751),.clk(gclk));
	jxor g03530(.dina(n3751),.dinb(w_n3587_0[0]),.dout(n3752),.clk(gclk));
	jnot g03531(.din(w_n3752_0[2]),.dout(n3753),.clk(gclk));
	jor g03532(.dina(n3753),.dinb(n3749),.dout(n3754),.clk(gclk));
	jand g03533(.dina(n3754),.dinb(w_n3748_0[1]),.dout(n3755),.clk(gclk));
	jor g03534(.dina(w_n3755_0[2]),.dinb(w_n743_57[1]),.dout(n3756),.clk(gclk));
	jand g03535(.dina(w_n3755_0[1]),.dinb(w_n743_57[0]),.dout(n3757),.clk(gclk));
	jxor g03536(.dina(w_n3450_0[0]),.dinb(w_n884_55[2]),.dout(n3758),.clk(gclk));
	jor g03537(.dina(n3758),.dinb(w_n3642_55[2]),.dout(n3759),.clk(gclk));
	jxor g03538(.dina(n3759),.dinb(w_n3456_0[0]),.dout(n3760),.clk(gclk));
	jor g03539(.dina(w_n3760_0[2]),.dinb(n3757),.dout(n3761),.clk(gclk));
	jand g03540(.dina(n3761),.dinb(w_n3756_0[1]),.dout(n3762),.clk(gclk));
	jor g03541(.dina(w_n3762_0[2]),.dinb(w_n635_57[1]),.dout(n3763),.clk(gclk));
	jand g03542(.dina(w_n3762_0[1]),.dinb(w_n635_57[0]),.dout(n3764),.clk(gclk));
	jxor g03543(.dina(w_n3458_0[0]),.dinb(w_n743_56[2]),.dout(n3765),.clk(gclk));
	jor g03544(.dina(n3765),.dinb(w_n3642_55[1]),.dout(n3766),.clk(gclk));
	jxor g03545(.dina(n3766),.dinb(w_n3594_0[0]),.dout(n3767),.clk(gclk));
	jnot g03546(.din(w_n3767_0[2]),.dout(n3768),.clk(gclk));
	jor g03547(.dina(n3768),.dinb(n3764),.dout(n3769),.clk(gclk));
	jand g03548(.dina(n3769),.dinb(w_n3763_0[1]),.dout(n3770),.clk(gclk));
	jor g03549(.dina(w_n3770_0[2]),.dinb(w_n515_58[1]),.dout(n3771),.clk(gclk));
	jand g03550(.dina(w_n3770_0[1]),.dinb(w_n515_58[0]),.dout(n3772),.clk(gclk));
	jxor g03551(.dina(w_n3465_0[0]),.dinb(w_n635_56[2]),.dout(n3773),.clk(gclk));
	jor g03552(.dina(n3773),.dinb(w_n3642_55[0]),.dout(n3774),.clk(gclk));
	jxor g03553(.dina(n3774),.dinb(w_n3471_0[0]),.dout(n3775),.clk(gclk));
	jor g03554(.dina(w_n3775_0[2]),.dinb(n3772),.dout(n3776),.clk(gclk));
	jand g03555(.dina(n3776),.dinb(w_n3771_0[1]),.dout(n3777),.clk(gclk));
	jor g03556(.dina(w_n3777_0[2]),.dinb(w_n443_58[1]),.dout(n3778),.clk(gclk));
	jand g03557(.dina(w_n3777_0[1]),.dinb(w_n443_58[0]),.dout(n3779),.clk(gclk));
	jxor g03558(.dina(w_n3473_0[0]),.dinb(w_n515_57[2]),.dout(n3780),.clk(gclk));
	jor g03559(.dina(n3780),.dinb(w_n3642_54[2]),.dout(n3781),.clk(gclk));
	jxor g03560(.dina(n3781),.dinb(w_n3601_0[0]),.dout(n3782),.clk(gclk));
	jnot g03561(.din(w_n3782_0[2]),.dout(n3783),.clk(gclk));
	jor g03562(.dina(n3783),.dinb(n3779),.dout(n3784),.clk(gclk));
	jand g03563(.dina(n3784),.dinb(w_n3778_0[1]),.dout(n3785),.clk(gclk));
	jor g03564(.dina(w_n3785_0[2]),.dinb(w_n352_58[2]),.dout(n3786),.clk(gclk));
	jand g03565(.dina(w_n3785_0[1]),.dinb(w_n352_58[1]),.dout(n3787),.clk(gclk));
	jxor g03566(.dina(w_n3480_0[0]),.dinb(w_n443_57[2]),.dout(n3788),.clk(gclk));
	jor g03567(.dina(n3788),.dinb(w_n3642_54[1]),.dout(n3789),.clk(gclk));
	jxor g03568(.dina(n3789),.dinb(w_n3486_0[0]),.dout(n3790),.clk(gclk));
	jor g03569(.dina(w_n3790_0[2]),.dinb(n3787),.dout(n3791),.clk(gclk));
	jand g03570(.dina(n3791),.dinb(w_n3786_0[1]),.dout(n3792),.clk(gclk));
	jor g03571(.dina(w_n3792_0[2]),.dinb(w_n294_59[0]),.dout(n3793),.clk(gclk));
	jand g03572(.dina(w_n3792_0[1]),.dinb(w_n294_58[2]),.dout(n3794),.clk(gclk));
	jxor g03573(.dina(w_n3488_0[0]),.dinb(w_n352_58[0]),.dout(n3795),.clk(gclk));
	jor g03574(.dina(n3795),.dinb(w_n3642_54[0]),.dout(n3796),.clk(gclk));
	jxor g03575(.dina(n3796),.dinb(w_n3494_0[0]),.dout(n3797),.clk(gclk));
	jor g03576(.dina(w_n3797_0[2]),.dinb(n3794),.dout(n3798),.clk(gclk));
	jand g03577(.dina(n3798),.dinb(w_n3793_0[1]),.dout(n3799),.clk(gclk));
	jor g03578(.dina(w_n3799_0[2]),.dinb(w_n239_59[0]),.dout(n3800),.clk(gclk));
	jand g03579(.dina(w_n3799_0[1]),.dinb(w_n239_58[2]),.dout(n3801),.clk(gclk));
	jxor g03580(.dina(w_n3496_0[0]),.dinb(w_n294_58[1]),.dout(n3802),.clk(gclk));
	jor g03581(.dina(n3802),.dinb(w_n3642_53[2]),.dout(n3803),.clk(gclk));
	jxor g03582(.dina(n3803),.dinb(w_n3611_0[0]),.dout(n3804),.clk(gclk));
	jnot g03583(.din(w_n3804_0[2]),.dout(n3805),.clk(gclk));
	jor g03584(.dina(n3805),.dinb(n3801),.dout(n3806),.clk(gclk));
	jand g03585(.dina(n3806),.dinb(w_n3800_0[1]),.dout(n3807),.clk(gclk));
	jor g03586(.dina(w_n3807_0[2]),.dinb(w_n221_59[0]),.dout(n3808),.clk(gclk));
	jand g03587(.dina(w_n3807_0[1]),.dinb(w_n221_58[2]),.dout(n3809),.clk(gclk));
	jxor g03588(.dina(w_n3503_0[0]),.dinb(w_n239_58[1]),.dout(n3810),.clk(gclk));
	jor g03589(.dina(n3810),.dinb(w_n3642_53[1]),.dout(n3811),.clk(gclk));
	jxor g03590(.dina(n3811),.dinb(w_n3615_0[0]),.dout(n3812),.clk(gclk));
	jnot g03591(.din(w_n3812_0[2]),.dout(n3813),.clk(gclk));
	jor g03592(.dina(n3813),.dinb(n3809),.dout(n3814),.clk(gclk));
	jand g03593(.dina(n3814),.dinb(w_n3808_0[1]),.dout(n3815),.clk(gclk));
	jand g03594(.dina(w_n3815_1[1]),.dinb(w_n3646_1[1]),.dout(n3816),.clk(gclk));
	jand g03595(.dina(w_n3640_0[0]),.dinb(w_n3620_0[0]),.dout(n3817),.clk(gclk));
	jand g03596(.dina(w_n3621_0[0]),.dinb(w_asqrt63_44[2]),.dout(n3818),.clk(gclk));
	jand g03597(.dina(n3818),.dinb(w_n3523_0[2]),.dout(n3819),.clk(gclk));
	jnot g03598(.din(n3819),.dout(n3820),.clk(gclk));
	jor g03599(.dina(w_n3820_0[1]),.dinb(n3817),.dout(n3821),.clk(gclk));
	jnot g03600(.din(w_n3821_0[1]),.dout(n3822),.clk(gclk));
	jand g03601(.dina(w_n3631_0[0]),.dinb(w_n3635_0[0]),.dout(n3823),.clk(gclk));
	jor g03602(.dina(w_n3815_1[0]),.dinb(w_n3646_1[0]),.dout(n3824),.clk(gclk));
	jor g03603(.dina(n3824),.dinb(w_n3524_0[0]),.dout(n3825),.clk(gclk));
	jor g03604(.dina(n3825),.dinb(w_n3823_0[1]),.dout(n3826),.clk(gclk));
	jand g03605(.dina(n3826),.dinb(w_n218_24[1]),.dout(n3827),.clk(gclk));
	jand g03606(.dina(w_n3642_53[0]),.dinb(w_n3521_0[0]),.dout(n3828),.clk(gclk));
	jor g03607(.dina(w_n3828_0[1]),.dinb(n3827),.dout(n3829),.clk(gclk));
	jor g03608(.dina(n3829),.dinb(n3822),.dout(n3830),.clk(gclk));
	jor g03609(.dina(n3830),.dinb(w_n3816_0[1]),.dout(asqrt_fa_41),.clk(gclk));
	jxor g03610(.dina(w_n3807_0[0]),.dinb(w_n221_58[1]),.dout(n3832),.clk(gclk));
	jand g03611(.dina(n3832),.dinb(w_asqrt40_40[1]),.dout(n3833),.clk(gclk));
	jxor g03612(.dina(n3833),.dinb(w_n3812_0[1]),.dout(n3834),.clk(gclk));
	jnot g03613(.din(w_n3834_0[2]),.dout(n3835),.clk(gclk));
	jand g03614(.dina(w_asqrt40_40[0]),.dinb(w_a80_0[1]),.dout(n3836),.clk(gclk));
	jnot g03615(.din(w_a78_1[1]),.dout(n3837),.clk(gclk));
	jnot g03616(.din(w_a79_0[1]),.dout(n3838),.clk(gclk));
	jand g03617(.dina(w_n3838_0[1]),.dinb(w_n3837_1[1]),.dout(n3839),.clk(gclk));
	jand g03618(.dina(w_n3839_0[2]),.dinb(w_n3648_1[1]),.dout(n3840),.clk(gclk));
	jor g03619(.dina(w_n3840_0[1]),.dinb(n3836),.dout(n3841),.clk(gclk));
	jand g03620(.dina(w_n3841_0[2]),.dinb(w_asqrt41_30[2]),.dout(n3842),.clk(gclk));
	jor g03621(.dina(w_n3841_0[1]),.dinb(w_asqrt41_30[1]),.dout(n3843),.clk(gclk));
	jand g03622(.dina(w_asqrt40_39[2]),.dinb(w_n3648_1[0]),.dout(n3844),.clk(gclk));
	jor g03623(.dina(n3844),.dinb(w_n3649_0[0]),.dout(n3845),.clk(gclk));
	jnot g03624(.din(w_n3650_0[1]),.dout(n3846),.clk(gclk));
	jnot g03625(.din(w_n3816_0[0]),.dout(n3847),.clk(gclk));
	jnot g03626(.din(w_n3823_0[0]),.dout(n3848),.clk(gclk));
	jnot g03627(.din(w_n3808_0[0]),.dout(n3849),.clk(gclk));
	jnot g03628(.din(w_n3800_0[0]),.dout(n3850),.clk(gclk));
	jnot g03629(.din(w_n3793_0[0]),.dout(n3851),.clk(gclk));
	jnot g03630(.din(w_n3786_0[0]),.dout(n3852),.clk(gclk));
	jnot g03631(.din(w_n3778_0[0]),.dout(n3853),.clk(gclk));
	jnot g03632(.din(w_n3771_0[0]),.dout(n3854),.clk(gclk));
	jnot g03633(.din(w_n3763_0[0]),.dout(n3855),.clk(gclk));
	jnot g03634(.din(w_n3756_0[0]),.dout(n3856),.clk(gclk));
	jnot g03635(.din(w_n3748_0[0]),.dout(n3857),.clk(gclk));
	jnot g03636(.din(w_n3741_0[0]),.dout(n3858),.clk(gclk));
	jnot g03637(.din(w_n3733_0[0]),.dout(n3859),.clk(gclk));
	jnot g03638(.din(w_n3726_0[0]),.dout(n3860),.clk(gclk));
	jnot g03639(.din(w_n3718_0[0]),.dout(n3861),.clk(gclk));
	jnot g03640(.din(w_n3711_0[0]),.dout(n3862),.clk(gclk));
	jnot g03641(.din(w_n3704_0[0]),.dout(n3863),.clk(gclk));
	jnot g03642(.din(w_n3696_0[0]),.dout(n3864),.clk(gclk));
	jnot g03643(.din(w_n3688_0[0]),.dout(n3865),.clk(gclk));
	jnot g03644(.din(w_n3681_0[0]),.dout(n3866),.clk(gclk));
	jnot g03645(.din(w_n3673_0[0]),.dout(n3867),.clk(gclk));
	jnot g03646(.din(w_n3662_0[0]),.dout(n3868),.clk(gclk));
	jnot g03647(.din(w_n3654_0[0]),.dout(n3869),.clk(gclk));
	jand g03648(.dina(w_asqrt41_30[0]),.dinb(w_a82_0[2]),.dout(n3870),.clk(gclk));
	jor g03649(.dina(w_n3651_0[0]),.dinb(n3870),.dout(n3871),.clk(gclk));
	jor g03650(.dina(n3871),.dinb(w_asqrt42_33[1]),.dout(n3872),.clk(gclk));
	jand g03651(.dina(w_asqrt41_29[2]),.dinb(w_n3258_0[1]),.dout(n3873),.clk(gclk));
	jor g03652(.dina(n3873),.dinb(w_n3259_0[0]),.dout(n3874),.clk(gclk));
	jand g03653(.dina(w_n3665_0[0]),.dinb(n3874),.dout(n3875),.clk(gclk));
	jand g03654(.dina(w_n3875_0[1]),.dinb(n3872),.dout(n3876),.clk(gclk));
	jor g03655(.dina(n3876),.dinb(n3869),.dout(n3877),.clk(gclk));
	jor g03656(.dina(n3877),.dinb(w_asqrt43_30[1]),.dout(n3878),.clk(gclk));
	jnot g03657(.din(w_n3670_0[1]),.dout(n3879),.clk(gclk));
	jand g03658(.dina(n3879),.dinb(n3878),.dout(n3880),.clk(gclk));
	jor g03659(.dina(n3880),.dinb(n3868),.dout(n3881),.clk(gclk));
	jor g03660(.dina(n3881),.dinb(w_asqrt44_33[1]),.dout(n3882),.clk(gclk));
	jand g03661(.dina(w_n3677_0[1]),.dinb(n3882),.dout(n3883),.clk(gclk));
	jor g03662(.dina(n3883),.dinb(n3867),.dout(n3884),.clk(gclk));
	jor g03663(.dina(n3884),.dinb(w_asqrt45_31[0]),.dout(n3885),.clk(gclk));
	jnot g03664(.din(w_n3685_0[1]),.dout(n3886),.clk(gclk));
	jand g03665(.dina(n3886),.dinb(n3885),.dout(n3887),.clk(gclk));
	jor g03666(.dina(n3887),.dinb(n3866),.dout(n3888),.clk(gclk));
	jor g03667(.dina(n3888),.dinb(w_asqrt46_33[1]),.dout(n3889),.clk(gclk));
	jand g03668(.dina(w_n3692_0[1]),.dinb(n3889),.dout(n3890),.clk(gclk));
	jor g03669(.dina(n3890),.dinb(n3865),.dout(n3891),.clk(gclk));
	jor g03670(.dina(n3891),.dinb(w_asqrt47_31[2]),.dout(n3892),.clk(gclk));
	jand g03671(.dina(w_n3700_0[1]),.dinb(n3892),.dout(n3893),.clk(gclk));
	jor g03672(.dina(n3893),.dinb(n3864),.dout(n3894),.clk(gclk));
	jor g03673(.dina(n3894),.dinb(w_asqrt48_33[2]),.dout(n3895),.clk(gclk));
	jnot g03674(.din(w_n3708_0[1]),.dout(n3896),.clk(gclk));
	jand g03675(.dina(n3896),.dinb(n3895),.dout(n3897),.clk(gclk));
	jor g03676(.dina(n3897),.dinb(n3863),.dout(n3898),.clk(gclk));
	jor g03677(.dina(n3898),.dinb(w_asqrt49_32[0]),.dout(n3899),.clk(gclk));
	jnot g03678(.din(w_n3715_0[1]),.dout(n3900),.clk(gclk));
	jand g03679(.dina(n3900),.dinb(n3899),.dout(n3901),.clk(gclk));
	jor g03680(.dina(n3901),.dinb(n3862),.dout(n3902),.clk(gclk));
	jor g03681(.dina(n3902),.dinb(w_asqrt50_34[0]),.dout(n3903),.clk(gclk));
	jand g03682(.dina(w_n3722_0[1]),.dinb(n3903),.dout(n3904),.clk(gclk));
	jor g03683(.dina(n3904),.dinb(n3861),.dout(n3905),.clk(gclk));
	jor g03684(.dina(n3905),.dinb(w_asqrt51_32[1]),.dout(n3906),.clk(gclk));
	jnot g03685(.din(w_n3730_0[1]),.dout(n3907),.clk(gclk));
	jand g03686(.dina(n3907),.dinb(n3906),.dout(n3908),.clk(gclk));
	jor g03687(.dina(n3908),.dinb(n3860),.dout(n3909),.clk(gclk));
	jor g03688(.dina(n3909),.dinb(w_asqrt52_34[0]),.dout(n3910),.clk(gclk));
	jand g03689(.dina(w_n3737_0[1]),.dinb(n3910),.dout(n3911),.clk(gclk));
	jor g03690(.dina(n3911),.dinb(n3859),.dout(n3912),.clk(gclk));
	jor g03691(.dina(n3912),.dinb(w_asqrt53_33[0]),.dout(n3913),.clk(gclk));
	jnot g03692(.din(w_n3745_0[1]),.dout(n3914),.clk(gclk));
	jand g03693(.dina(n3914),.dinb(n3913),.dout(n3915),.clk(gclk));
	jor g03694(.dina(n3915),.dinb(n3858),.dout(n3916),.clk(gclk));
	jor g03695(.dina(n3916),.dinb(w_asqrt54_34[0]),.dout(n3917),.clk(gclk));
	jand g03696(.dina(w_n3752_0[1]),.dinb(n3917),.dout(n3918),.clk(gclk));
	jor g03697(.dina(n3918),.dinb(n3857),.dout(n3919),.clk(gclk));
	jor g03698(.dina(n3919),.dinb(w_asqrt55_33[1]),.dout(n3920),.clk(gclk));
	jnot g03699(.din(w_n3760_0[1]),.dout(n3921),.clk(gclk));
	jand g03700(.dina(n3921),.dinb(n3920),.dout(n3922),.clk(gclk));
	jor g03701(.dina(n3922),.dinb(n3856),.dout(n3923),.clk(gclk));
	jor g03702(.dina(n3923),.dinb(w_asqrt56_34[1]),.dout(n3924),.clk(gclk));
	jand g03703(.dina(w_n3767_0[1]),.dinb(n3924),.dout(n3925),.clk(gclk));
	jor g03704(.dina(n3925),.dinb(n3855),.dout(n3926),.clk(gclk));
	jor g03705(.dina(n3926),.dinb(w_asqrt57_34[0]),.dout(n3927),.clk(gclk));
	jnot g03706(.din(w_n3775_0[1]),.dout(n3928),.clk(gclk));
	jand g03707(.dina(n3928),.dinb(n3927),.dout(n3929),.clk(gclk));
	jor g03708(.dina(n3929),.dinb(n3854),.dout(n3930),.clk(gclk));
	jor g03709(.dina(n3930),.dinb(w_asqrt58_34[2]),.dout(n3931),.clk(gclk));
	jand g03710(.dina(w_n3782_0[1]),.dinb(n3931),.dout(n3932),.clk(gclk));
	jor g03711(.dina(n3932),.dinb(n3853),.dout(n3933),.clk(gclk));
	jor g03712(.dina(n3933),.dinb(w_asqrt59_34[1]),.dout(n3934),.clk(gclk));
	jnot g03713(.din(w_n3790_0[1]),.dout(n3935),.clk(gclk));
	jand g03714(.dina(n3935),.dinb(n3934),.dout(n3936),.clk(gclk));
	jor g03715(.dina(n3936),.dinb(n3852),.dout(n3937),.clk(gclk));
	jor g03716(.dina(n3937),.dinb(w_asqrt60_34[2]),.dout(n3938),.clk(gclk));
	jnot g03717(.din(w_n3797_0[1]),.dout(n3939),.clk(gclk));
	jand g03718(.dina(n3939),.dinb(n3938),.dout(n3940),.clk(gclk));
	jor g03719(.dina(n3940),.dinb(n3851),.dout(n3941),.clk(gclk));
	jor g03720(.dina(n3941),.dinb(w_asqrt61_34[2]),.dout(n3942),.clk(gclk));
	jand g03721(.dina(w_n3804_0[1]),.dinb(n3942),.dout(n3943),.clk(gclk));
	jor g03722(.dina(n3943),.dinb(n3850),.dout(n3944),.clk(gclk));
	jor g03723(.dina(n3944),.dinb(w_asqrt62_34[2]),.dout(n3945),.clk(gclk));
	jand g03724(.dina(w_n3812_0[0]),.dinb(n3945),.dout(n3946),.clk(gclk));
	jor g03725(.dina(n3946),.dinb(n3849),.dout(n3947),.clk(gclk));
	jand g03726(.dina(n3947),.dinb(w_n3645_0[0]),.dout(n3948),.clk(gclk));
	jand g03727(.dina(n3948),.dinb(w_n3523_0[1]),.dout(n3949),.clk(gclk));
	jand g03728(.dina(n3949),.dinb(n3848),.dout(n3950),.clk(gclk));
	jor g03729(.dina(n3950),.dinb(w_asqrt63_44[1]),.dout(n3951),.clk(gclk));
	jnot g03730(.din(w_n3828_0[0]),.dout(n3952),.clk(gclk));
	jand g03731(.dina(n3952),.dinb(w_n3951_0[1]),.dout(n3953),.clk(gclk));
	jand g03732(.dina(n3953),.dinb(w_n3821_0[0]),.dout(n3954),.clk(gclk));
	jand g03733(.dina(w_n3954_0[1]),.dinb(w_n3847_0[1]),.dout(n3955),.clk(gclk));
	jor g03734(.dina(w_n3955_50[1]),.dinb(n3846),.dout(n3956),.clk(gclk));
	jand g03735(.dina(n3956),.dinb(n3845),.dout(n3957),.clk(gclk));
	jand g03736(.dina(w_n3957_0[1]),.dinb(n3843),.dout(n3958),.clk(gclk));
	jor g03737(.dina(n3958),.dinb(w_n3842_0[1]),.dout(n3959),.clk(gclk));
	jand g03738(.dina(w_n3959_0[2]),.dinb(w_asqrt42_33[0]),.dout(n3960),.clk(gclk));
	jor g03739(.dina(w_n3959_0[1]),.dinb(w_asqrt42_32[2]),.dout(n3961),.clk(gclk));
	jand g03740(.dina(w_asqrt40_39[1]),.dinb(w_n3650_0[0]),.dout(n3962),.clk(gclk));
	jand g03741(.dina(w_n3847_0[0]),.dinb(w_asqrt41_29[1]),.dout(n3963),.clk(gclk));
	jand g03742(.dina(n3963),.dinb(w_n3820_0[0]),.dout(n3964),.clk(gclk));
	jand g03743(.dina(n3964),.dinb(w_n3951_0[0]),.dout(n3965),.clk(gclk));
	jor g03744(.dina(n3965),.dinb(w_n3962_0[1]),.dout(n3966),.clk(gclk));
	jxor g03745(.dina(n3966),.dinb(w_a82_0[1]),.dout(n3967),.clk(gclk));
	jnot g03746(.din(w_n3967_0[1]),.dout(n3968),.clk(gclk));
	jand g03747(.dina(w_n3968_0[1]),.dinb(n3961),.dout(n3969),.clk(gclk));
	jor g03748(.dina(n3969),.dinb(w_n3960_0[1]),.dout(n3970),.clk(gclk));
	jand g03749(.dina(w_n3970_0[2]),.dinb(w_asqrt43_30[0]),.dout(n3971),.clk(gclk));
	jor g03750(.dina(w_n3970_0[1]),.dinb(w_asqrt43_29[2]),.dout(n3972),.clk(gclk));
	jxor g03751(.dina(w_n3653_0[0]),.dinb(w_n3368_50[1]),.dout(n3973),.clk(gclk));
	jand g03752(.dina(n3973),.dinb(w_asqrt40_39[0]),.dout(n3974),.clk(gclk));
	jxor g03753(.dina(n3974),.dinb(w_n3875_0[0]),.dout(n3975),.clk(gclk));
	jand g03754(.dina(w_n3975_0[1]),.dinb(n3972),.dout(n3976),.clk(gclk));
	jor g03755(.dina(n3976),.dinb(w_n3971_0[1]),.dout(n3977),.clk(gclk));
	jand g03756(.dina(w_n3977_0[2]),.dinb(w_asqrt44_33[0]),.dout(n3978),.clk(gclk));
	jor g03757(.dina(w_n3977_0[1]),.dinb(w_asqrt44_32[2]),.dout(n3979),.clk(gclk));
	jxor g03758(.dina(w_n3661_0[0]),.dinb(w_n3089_53[2]),.dout(n3980),.clk(gclk));
	jand g03759(.dina(n3980),.dinb(w_asqrt40_38[2]),.dout(n3981),.clk(gclk));
	jxor g03760(.dina(n3981),.dinb(w_n3670_0[0]),.dout(n3982),.clk(gclk));
	jnot g03761(.din(w_n3982_0[1]),.dout(n3983),.clk(gclk));
	jand g03762(.dina(w_n3983_0[1]),.dinb(n3979),.dout(n3984),.clk(gclk));
	jor g03763(.dina(n3984),.dinb(w_n3978_0[1]),.dout(n3985),.clk(gclk));
	jand g03764(.dina(w_n3985_0[2]),.dinb(w_asqrt45_30[2]),.dout(n3986),.clk(gclk));
	jor g03765(.dina(w_n3985_0[1]),.dinb(w_asqrt45_30[1]),.dout(n3987),.clk(gclk));
	jxor g03766(.dina(w_n3672_0[0]),.dinb(w_n2833_51[1]),.dout(n3988),.clk(gclk));
	jand g03767(.dina(n3988),.dinb(w_asqrt40_38[1]),.dout(n3989),.clk(gclk));
	jxor g03768(.dina(n3989),.dinb(w_n3677_0[0]),.dout(n3990),.clk(gclk));
	jand g03769(.dina(w_n3990_0[1]),.dinb(n3987),.dout(n3991),.clk(gclk));
	jor g03770(.dina(n3991),.dinb(w_n3986_0[1]),.dout(n3992),.clk(gclk));
	jand g03771(.dina(w_n3992_0[2]),.dinb(w_asqrt46_33[0]),.dout(n3993),.clk(gclk));
	jor g03772(.dina(w_n3992_0[1]),.dinb(w_asqrt46_32[2]),.dout(n3994),.clk(gclk));
	jxor g03773(.dina(w_n3680_0[0]),.dinb(w_n2572_54[0]),.dout(n3995),.clk(gclk));
	jand g03774(.dina(n3995),.dinb(w_asqrt40_38[0]),.dout(n3996),.clk(gclk));
	jxor g03775(.dina(n3996),.dinb(w_n3685_0[0]),.dout(n3997),.clk(gclk));
	jnot g03776(.din(w_n3997_0[1]),.dout(n3998),.clk(gclk));
	jand g03777(.dina(w_n3998_0[1]),.dinb(n3994),.dout(n3999),.clk(gclk));
	jor g03778(.dina(n3999),.dinb(w_n3993_0[1]),.dout(n4000),.clk(gclk));
	jand g03779(.dina(w_n4000_0[2]),.dinb(w_asqrt47_31[1]),.dout(n4001),.clk(gclk));
	jor g03780(.dina(w_n4000_0[1]),.dinb(w_asqrt47_31[0]),.dout(n4002),.clk(gclk));
	jxor g03781(.dina(w_n3687_0[0]),.dinb(w_n2345_52[0]),.dout(n4003),.clk(gclk));
	jand g03782(.dina(n4003),.dinb(w_asqrt40_37[2]),.dout(n4004),.clk(gclk));
	jxor g03783(.dina(n4004),.dinb(w_n3692_0[0]),.dout(n4005),.clk(gclk));
	jand g03784(.dina(w_n4005_0[1]),.dinb(n4002),.dout(n4006),.clk(gclk));
	jor g03785(.dina(n4006),.dinb(w_n4001_0[1]),.dout(n4007),.clk(gclk));
	jand g03786(.dina(w_n4007_0[2]),.dinb(w_asqrt48_33[1]),.dout(n4008),.clk(gclk));
	jor g03787(.dina(w_n4007_0[1]),.dinb(w_asqrt48_33[0]),.dout(n4009),.clk(gclk));
	jxor g03788(.dina(w_n3695_0[0]),.dinb(w_n2108_54[2]),.dout(n4010),.clk(gclk));
	jand g03789(.dina(n4010),.dinb(w_asqrt40_37[1]),.dout(n4011),.clk(gclk));
	jxor g03790(.dina(n4011),.dinb(w_n3700_0[0]),.dout(n4012),.clk(gclk));
	jand g03791(.dina(w_n4012_0[1]),.dinb(n4009),.dout(n4013),.clk(gclk));
	jor g03792(.dina(n4013),.dinb(w_n4008_0[1]),.dout(n4014),.clk(gclk));
	jand g03793(.dina(w_n4014_0[2]),.dinb(w_asqrt49_31[2]),.dout(n4015),.clk(gclk));
	jor g03794(.dina(w_n4014_0[1]),.dinb(w_asqrt49_31[1]),.dout(n4016),.clk(gclk));
	jxor g03795(.dina(w_n3703_0[0]),.dinb(w_n1912_53[0]),.dout(n4017),.clk(gclk));
	jand g03796(.dina(n4017),.dinb(w_asqrt40_37[0]),.dout(n4018),.clk(gclk));
	jxor g03797(.dina(n4018),.dinb(w_n3708_0[0]),.dout(n4019),.clk(gclk));
	jnot g03798(.din(w_n4019_0[1]),.dout(n4020),.clk(gclk));
	jand g03799(.dina(w_n4020_0[1]),.dinb(n4016),.dout(n4021),.clk(gclk));
	jor g03800(.dina(n4021),.dinb(w_n4015_0[1]),.dout(n4022),.clk(gclk));
	jand g03801(.dina(w_n4022_0[2]),.dinb(w_asqrt50_33[2]),.dout(n4023),.clk(gclk));
	jor g03802(.dina(w_n4022_0[1]),.dinb(w_asqrt50_33[1]),.dout(n4024),.clk(gclk));
	jxor g03803(.dina(w_n3710_0[0]),.dinb(w_n1699_55[1]),.dout(n4025),.clk(gclk));
	jand g03804(.dina(n4025),.dinb(w_asqrt40_36[2]),.dout(n4026),.clk(gclk));
	jxor g03805(.dina(n4026),.dinb(w_n3715_0[0]),.dout(n4027),.clk(gclk));
	jnot g03806(.din(w_n4027_0[1]),.dout(n4028),.clk(gclk));
	jand g03807(.dina(w_n4028_0[1]),.dinb(n4024),.dout(n4029),.clk(gclk));
	jor g03808(.dina(n4029),.dinb(w_n4023_0[1]),.dout(n4030),.clk(gclk));
	jand g03809(.dina(w_n4030_0[2]),.dinb(w_asqrt51_32[0]),.dout(n4031),.clk(gclk));
	jor g03810(.dina(w_n4030_0[1]),.dinb(w_asqrt51_31[2]),.dout(n4032),.clk(gclk));
	jxor g03811(.dina(w_n3717_0[0]),.dinb(w_n1516_53[2]),.dout(n4033),.clk(gclk));
	jand g03812(.dina(n4033),.dinb(w_asqrt40_36[1]),.dout(n4034),.clk(gclk));
	jxor g03813(.dina(n4034),.dinb(w_n3722_0[0]),.dout(n4035),.clk(gclk));
	jand g03814(.dina(w_n4035_0[1]),.dinb(n4032),.dout(n4036),.clk(gclk));
	jor g03815(.dina(n4036),.dinb(w_n4031_0[1]),.dout(n4037),.clk(gclk));
	jand g03816(.dina(w_n4037_0[2]),.dinb(w_asqrt52_33[2]),.dout(n4038),.clk(gclk));
	jor g03817(.dina(w_n4037_0[1]),.dinb(w_asqrt52_33[1]),.dout(n4039),.clk(gclk));
	jxor g03818(.dina(w_n3725_0[0]),.dinb(w_n1332_55[1]),.dout(n4040),.clk(gclk));
	jand g03819(.dina(n4040),.dinb(w_asqrt40_36[0]),.dout(n4041),.clk(gclk));
	jxor g03820(.dina(n4041),.dinb(w_n3730_0[0]),.dout(n4042),.clk(gclk));
	jnot g03821(.din(w_n4042_0[1]),.dout(n4043),.clk(gclk));
	jand g03822(.dina(w_n4043_0[1]),.dinb(n4039),.dout(n4044),.clk(gclk));
	jor g03823(.dina(n4044),.dinb(w_n4038_0[1]),.dout(n4045),.clk(gclk));
	jand g03824(.dina(w_n4045_0[2]),.dinb(w_asqrt53_32[2]),.dout(n4046),.clk(gclk));
	jor g03825(.dina(w_n4045_0[1]),.dinb(w_asqrt53_32[1]),.dout(n4047),.clk(gclk));
	jxor g03826(.dina(w_n3732_0[0]),.dinb(w_n1173_54[1]),.dout(n4048),.clk(gclk));
	jand g03827(.dina(n4048),.dinb(w_asqrt40_35[2]),.dout(n4049),.clk(gclk));
	jxor g03828(.dina(n4049),.dinb(w_n3737_0[0]),.dout(n4050),.clk(gclk));
	jand g03829(.dina(w_n4050_0[1]),.dinb(n4047),.dout(n4051),.clk(gclk));
	jor g03830(.dina(n4051),.dinb(w_n4046_0[1]),.dout(n4052),.clk(gclk));
	jand g03831(.dina(w_n4052_0[2]),.dinb(w_asqrt54_33[2]),.dout(n4053),.clk(gclk));
	jor g03832(.dina(w_n4052_0[1]),.dinb(w_asqrt54_33[1]),.dout(n4054),.clk(gclk));
	jxor g03833(.dina(w_n3740_0[0]),.dinb(w_n1008_56[1]),.dout(n4055),.clk(gclk));
	jand g03834(.dina(n4055),.dinb(w_asqrt40_35[1]),.dout(n4056),.clk(gclk));
	jxor g03835(.dina(n4056),.dinb(w_n3745_0[0]),.dout(n4057),.clk(gclk));
	jnot g03836(.din(w_n4057_0[1]),.dout(n4058),.clk(gclk));
	jand g03837(.dina(w_n4058_0[1]),.dinb(n4054),.dout(n4059),.clk(gclk));
	jor g03838(.dina(n4059),.dinb(w_n4053_0[1]),.dout(n4060),.clk(gclk));
	jand g03839(.dina(w_n4060_0[2]),.dinb(w_asqrt55_33[0]),.dout(n4061),.clk(gclk));
	jor g03840(.dina(w_n4060_0[1]),.dinb(w_asqrt55_32[2]),.dout(n4062),.clk(gclk));
	jxor g03841(.dina(w_n3747_0[0]),.dinb(w_n884_55[1]),.dout(n4063),.clk(gclk));
	jand g03842(.dina(n4063),.dinb(w_asqrt40_35[0]),.dout(n4064),.clk(gclk));
	jxor g03843(.dina(n4064),.dinb(w_n3752_0[0]),.dout(n4065),.clk(gclk));
	jand g03844(.dina(w_n4065_0[1]),.dinb(n4062),.dout(n4066),.clk(gclk));
	jor g03845(.dina(n4066),.dinb(w_n4061_0[1]),.dout(n4067),.clk(gclk));
	jand g03846(.dina(w_n4067_0[2]),.dinb(w_asqrt56_34[0]),.dout(n4068),.clk(gclk));
	jor g03847(.dina(w_n4067_0[1]),.dinb(w_asqrt56_33[2]),.dout(n4069),.clk(gclk));
	jxor g03848(.dina(w_n3755_0[0]),.dinb(w_n743_56[1]),.dout(n4070),.clk(gclk));
	jand g03849(.dina(n4070),.dinb(w_asqrt40_34[2]),.dout(n4071),.clk(gclk));
	jxor g03850(.dina(n4071),.dinb(w_n3760_0[0]),.dout(n4072),.clk(gclk));
	jnot g03851(.din(w_n4072_0[1]),.dout(n4073),.clk(gclk));
	jand g03852(.dina(w_n4073_0[1]),.dinb(n4069),.dout(n4074),.clk(gclk));
	jor g03853(.dina(n4074),.dinb(w_n4068_0[1]),.dout(n4075),.clk(gclk));
	jand g03854(.dina(w_n4075_0[2]),.dinb(w_asqrt57_33[2]),.dout(n4076),.clk(gclk));
	jor g03855(.dina(w_n4075_0[1]),.dinb(w_asqrt57_33[1]),.dout(n4077),.clk(gclk));
	jxor g03856(.dina(w_n3762_0[0]),.dinb(w_n635_56[1]),.dout(n4078),.clk(gclk));
	jand g03857(.dina(n4078),.dinb(w_asqrt40_34[1]),.dout(n4079),.clk(gclk));
	jxor g03858(.dina(n4079),.dinb(w_n3767_0[0]),.dout(n4080),.clk(gclk));
	jand g03859(.dina(w_n4080_0[1]),.dinb(n4077),.dout(n4081),.clk(gclk));
	jor g03860(.dina(n4081),.dinb(w_n4076_0[1]),.dout(n4082),.clk(gclk));
	jand g03861(.dina(w_n4082_0[2]),.dinb(w_asqrt58_34[1]),.dout(n4083),.clk(gclk));
	jor g03862(.dina(w_n4082_0[1]),.dinb(w_asqrt58_34[0]),.dout(n4084),.clk(gclk));
	jxor g03863(.dina(w_n3770_0[0]),.dinb(w_n515_57[1]),.dout(n4085),.clk(gclk));
	jand g03864(.dina(n4085),.dinb(w_asqrt40_34[0]),.dout(n4086),.clk(gclk));
	jxor g03865(.dina(n4086),.dinb(w_n3775_0[0]),.dout(n4087),.clk(gclk));
	jnot g03866(.din(w_n4087_0[1]),.dout(n4088),.clk(gclk));
	jand g03867(.dina(w_n4088_0[1]),.dinb(n4084),.dout(n4089),.clk(gclk));
	jor g03868(.dina(n4089),.dinb(w_n4083_0[1]),.dout(n4090),.clk(gclk));
	jand g03869(.dina(w_n4090_0[2]),.dinb(w_asqrt59_34[0]),.dout(n4091),.clk(gclk));
	jor g03870(.dina(w_n4090_0[1]),.dinb(w_asqrt59_33[2]),.dout(n4092),.clk(gclk));
	jxor g03871(.dina(w_n3777_0[0]),.dinb(w_n443_57[1]),.dout(n4093),.clk(gclk));
	jand g03872(.dina(n4093),.dinb(w_asqrt40_33[2]),.dout(n4094),.clk(gclk));
	jxor g03873(.dina(n4094),.dinb(w_n3782_0[0]),.dout(n4095),.clk(gclk));
	jand g03874(.dina(w_n4095_0[1]),.dinb(n4092),.dout(n4096),.clk(gclk));
	jor g03875(.dina(n4096),.dinb(w_n4091_0[1]),.dout(n4097),.clk(gclk));
	jand g03876(.dina(w_n4097_0[2]),.dinb(w_asqrt60_34[1]),.dout(n4098),.clk(gclk));
	jor g03877(.dina(w_n4097_0[1]),.dinb(w_asqrt60_34[0]),.dout(n4099),.clk(gclk));
	jxor g03878(.dina(w_n3785_0[0]),.dinb(w_n352_57[2]),.dout(n4100),.clk(gclk));
	jand g03879(.dina(n4100),.dinb(w_asqrt40_33[1]),.dout(n4101),.clk(gclk));
	jxor g03880(.dina(n4101),.dinb(w_n3790_0[0]),.dout(n4102),.clk(gclk));
	jnot g03881(.din(w_n4102_0[1]),.dout(n4103),.clk(gclk));
	jand g03882(.dina(w_n4103_0[1]),.dinb(n4099),.dout(n4104),.clk(gclk));
	jor g03883(.dina(n4104),.dinb(w_n4098_0[1]),.dout(n4105),.clk(gclk));
	jand g03884(.dina(w_n4105_0[2]),.dinb(w_asqrt61_34[1]),.dout(n4106),.clk(gclk));
	jor g03885(.dina(w_n4105_0[1]),.dinb(w_asqrt61_34[0]),.dout(n4107),.clk(gclk));
	jxor g03886(.dina(w_n3792_0[0]),.dinb(w_n294_58[0]),.dout(n4108),.clk(gclk));
	jand g03887(.dina(n4108),.dinb(w_asqrt40_33[0]),.dout(n4109),.clk(gclk));
	jxor g03888(.dina(n4109),.dinb(w_n3797_0[0]),.dout(n4110),.clk(gclk));
	jnot g03889(.din(w_n4110_0[1]),.dout(n4111),.clk(gclk));
	jand g03890(.dina(w_n4111_0[1]),.dinb(n4107),.dout(n4112),.clk(gclk));
	jor g03891(.dina(n4112),.dinb(w_n4106_0[1]),.dout(n4113),.clk(gclk));
	jand g03892(.dina(w_n4113_0[2]),.dinb(w_asqrt62_34[1]),.dout(n4114),.clk(gclk));
	jnot g03893(.din(w_n4114_0[1]),.dout(n4115),.clk(gclk));
	jnot g03894(.din(w_n4106_0[0]),.dout(n4116),.clk(gclk));
	jnot g03895(.din(w_n4098_0[0]),.dout(n4117),.clk(gclk));
	jnot g03896(.din(w_n4091_0[0]),.dout(n4118),.clk(gclk));
	jnot g03897(.din(w_n4083_0[0]),.dout(n4119),.clk(gclk));
	jnot g03898(.din(w_n4076_0[0]),.dout(n4120),.clk(gclk));
	jnot g03899(.din(w_n4068_0[0]),.dout(n4121),.clk(gclk));
	jnot g03900(.din(w_n4061_0[0]),.dout(n4122),.clk(gclk));
	jnot g03901(.din(w_n4053_0[0]),.dout(n4123),.clk(gclk));
	jnot g03902(.din(w_n4046_0[0]),.dout(n4124),.clk(gclk));
	jnot g03903(.din(w_n4038_0[0]),.dout(n4125),.clk(gclk));
	jnot g03904(.din(w_n4031_0[0]),.dout(n4126),.clk(gclk));
	jnot g03905(.din(w_n4023_0[0]),.dout(n4127),.clk(gclk));
	jnot g03906(.din(w_n4015_0[0]),.dout(n4128),.clk(gclk));
	jnot g03907(.din(w_n4008_0[0]),.dout(n4129),.clk(gclk));
	jnot g03908(.din(w_n4001_0[0]),.dout(n4130),.clk(gclk));
	jnot g03909(.din(w_n3993_0[0]),.dout(n4131),.clk(gclk));
	jnot g03910(.din(w_n3986_0[0]),.dout(n4132),.clk(gclk));
	jnot g03911(.din(w_n3978_0[0]),.dout(n4133),.clk(gclk));
	jnot g03912(.din(w_n3971_0[0]),.dout(n4134),.clk(gclk));
	jnot g03913(.din(w_n3960_0[0]),.dout(n4135),.clk(gclk));
	jnot g03914(.din(w_n3842_0[0]),.dout(n4136),.clk(gclk));
	jor g03915(.dina(w_n3955_50[0]),.dinb(w_n3648_0[2]),.dout(n4137),.clk(gclk));
	jnot g03916(.din(w_n3840_0[0]),.dout(n4138),.clk(gclk));
	jand g03917(.dina(n4138),.dinb(n4137),.dout(n4139),.clk(gclk));
	jand g03918(.dina(n4139),.dinb(w_n3642_52[2]),.dout(n4140),.clk(gclk));
	jor g03919(.dina(w_n3955_49[2]),.dinb(w_a80_0[0]),.dout(n4141),.clk(gclk));
	jand g03920(.dina(n4141),.dinb(w_a81_0[0]),.dout(n4142),.clk(gclk));
	jor g03921(.dina(w_n3962_0[0]),.dinb(n4142),.dout(n4143),.clk(gclk));
	jor g03922(.dina(n4143),.dinb(n4140),.dout(n4144),.clk(gclk));
	jand g03923(.dina(n4144),.dinb(n4136),.dout(n4145),.clk(gclk));
	jand g03924(.dina(n4145),.dinb(w_n3368_50[0]),.dout(n4146),.clk(gclk));
	jor g03925(.dina(w_n3967_0[0]),.dinb(n4146),.dout(n4147),.clk(gclk));
	jand g03926(.dina(n4147),.dinb(n4135),.dout(n4148),.clk(gclk));
	jand g03927(.dina(n4148),.dinb(w_n3089_53[1]),.dout(n4149),.clk(gclk));
	jnot g03928(.din(w_n3975_0[0]),.dout(n4150),.clk(gclk));
	jor g03929(.dina(w_n4150_0[1]),.dinb(n4149),.dout(n4151),.clk(gclk));
	jand g03930(.dina(n4151),.dinb(n4134),.dout(n4152),.clk(gclk));
	jand g03931(.dina(n4152),.dinb(w_n2833_51[0]),.dout(n4153),.clk(gclk));
	jor g03932(.dina(w_n3982_0[0]),.dinb(n4153),.dout(n4154),.clk(gclk));
	jand g03933(.dina(n4154),.dinb(n4133),.dout(n4155),.clk(gclk));
	jand g03934(.dina(n4155),.dinb(w_n2572_53[2]),.dout(n4156),.clk(gclk));
	jnot g03935(.din(w_n3990_0[0]),.dout(n4157),.clk(gclk));
	jor g03936(.dina(w_n4157_0[1]),.dinb(n4156),.dout(n4158),.clk(gclk));
	jand g03937(.dina(n4158),.dinb(n4132),.dout(n4159),.clk(gclk));
	jand g03938(.dina(n4159),.dinb(w_n2345_51[2]),.dout(n4160),.clk(gclk));
	jor g03939(.dina(w_n3997_0[0]),.dinb(n4160),.dout(n4161),.clk(gclk));
	jand g03940(.dina(n4161),.dinb(n4131),.dout(n4162),.clk(gclk));
	jand g03941(.dina(n4162),.dinb(w_n2108_54[1]),.dout(n4163),.clk(gclk));
	jnot g03942(.din(w_n4005_0[0]),.dout(n4164),.clk(gclk));
	jor g03943(.dina(w_n4164_0[1]),.dinb(n4163),.dout(n4165),.clk(gclk));
	jand g03944(.dina(n4165),.dinb(n4130),.dout(n4166),.clk(gclk));
	jand g03945(.dina(n4166),.dinb(w_n1912_52[2]),.dout(n4167),.clk(gclk));
	jnot g03946(.din(w_n4012_0[0]),.dout(n4168),.clk(gclk));
	jor g03947(.dina(w_n4168_0[1]),.dinb(n4167),.dout(n4169),.clk(gclk));
	jand g03948(.dina(n4169),.dinb(n4129),.dout(n4170),.clk(gclk));
	jand g03949(.dina(n4170),.dinb(w_n1699_55[0]),.dout(n4171),.clk(gclk));
	jor g03950(.dina(w_n4019_0[0]),.dinb(n4171),.dout(n4172),.clk(gclk));
	jand g03951(.dina(n4172),.dinb(n4128),.dout(n4173),.clk(gclk));
	jand g03952(.dina(n4173),.dinb(w_n1516_53[1]),.dout(n4174),.clk(gclk));
	jor g03953(.dina(w_n4027_0[0]),.dinb(n4174),.dout(n4175),.clk(gclk));
	jand g03954(.dina(n4175),.dinb(n4127),.dout(n4176),.clk(gclk));
	jand g03955(.dina(n4176),.dinb(w_n1332_55[0]),.dout(n4177),.clk(gclk));
	jnot g03956(.din(w_n4035_0[0]),.dout(n4178),.clk(gclk));
	jor g03957(.dina(w_n4178_0[1]),.dinb(n4177),.dout(n4179),.clk(gclk));
	jand g03958(.dina(n4179),.dinb(n4126),.dout(n4180),.clk(gclk));
	jand g03959(.dina(n4180),.dinb(w_n1173_54[0]),.dout(n4181),.clk(gclk));
	jor g03960(.dina(w_n4042_0[0]),.dinb(n4181),.dout(n4182),.clk(gclk));
	jand g03961(.dina(n4182),.dinb(n4125),.dout(n4183),.clk(gclk));
	jand g03962(.dina(n4183),.dinb(w_n1008_56[0]),.dout(n4184),.clk(gclk));
	jnot g03963(.din(w_n4050_0[0]),.dout(n4185),.clk(gclk));
	jor g03964(.dina(w_n4185_0[1]),.dinb(n4184),.dout(n4186),.clk(gclk));
	jand g03965(.dina(n4186),.dinb(n4124),.dout(n4187),.clk(gclk));
	jand g03966(.dina(n4187),.dinb(w_n884_55[0]),.dout(n4188),.clk(gclk));
	jor g03967(.dina(w_n4057_0[0]),.dinb(n4188),.dout(n4189),.clk(gclk));
	jand g03968(.dina(n4189),.dinb(n4123),.dout(n4190),.clk(gclk));
	jand g03969(.dina(n4190),.dinb(w_n743_56[0]),.dout(n4191),.clk(gclk));
	jnot g03970(.din(w_n4065_0[0]),.dout(n4192),.clk(gclk));
	jor g03971(.dina(w_n4192_0[1]),.dinb(n4191),.dout(n4193),.clk(gclk));
	jand g03972(.dina(n4193),.dinb(n4122),.dout(n4194),.clk(gclk));
	jand g03973(.dina(n4194),.dinb(w_n635_56[0]),.dout(n4195),.clk(gclk));
	jor g03974(.dina(w_n4072_0[0]),.dinb(n4195),.dout(n4196),.clk(gclk));
	jand g03975(.dina(n4196),.dinb(n4121),.dout(n4197),.clk(gclk));
	jand g03976(.dina(n4197),.dinb(w_n515_57[0]),.dout(n4198),.clk(gclk));
	jnot g03977(.din(w_n4080_0[0]),.dout(n4199),.clk(gclk));
	jor g03978(.dina(w_n4199_0[1]),.dinb(n4198),.dout(n4200),.clk(gclk));
	jand g03979(.dina(n4200),.dinb(n4120),.dout(n4201),.clk(gclk));
	jand g03980(.dina(n4201),.dinb(w_n443_57[0]),.dout(n4202),.clk(gclk));
	jor g03981(.dina(w_n4087_0[0]),.dinb(n4202),.dout(n4203),.clk(gclk));
	jand g03982(.dina(n4203),.dinb(n4119),.dout(n4204),.clk(gclk));
	jand g03983(.dina(n4204),.dinb(w_n352_57[1]),.dout(n4205),.clk(gclk));
	jnot g03984(.din(w_n4095_0[0]),.dout(n4206),.clk(gclk));
	jor g03985(.dina(w_n4206_0[1]),.dinb(n4205),.dout(n4207),.clk(gclk));
	jand g03986(.dina(n4207),.dinb(n4118),.dout(n4208),.clk(gclk));
	jand g03987(.dina(n4208),.dinb(w_n294_57[2]),.dout(n4209),.clk(gclk));
	jor g03988(.dina(w_n4102_0[0]),.dinb(n4209),.dout(n4210),.clk(gclk));
	jand g03989(.dina(n4210),.dinb(n4117),.dout(n4211),.clk(gclk));
	jand g03990(.dina(n4211),.dinb(w_n239_58[0]),.dout(n4212),.clk(gclk));
	jor g03991(.dina(w_n4110_0[0]),.dinb(n4212),.dout(n4213),.clk(gclk));
	jand g03992(.dina(n4213),.dinb(n4116),.dout(n4214),.clk(gclk));
	jand g03993(.dina(n4214),.dinb(w_n221_58[0]),.dout(n4215),.clk(gclk));
	jxor g03994(.dina(w_n3799_0[0]),.dinb(w_n239_57[2]),.dout(n4216),.clk(gclk));
	jand g03995(.dina(n4216),.dinb(w_asqrt40_32[2]),.dout(n4217),.clk(gclk));
	jxor g03996(.dina(n4217),.dinb(w_n3804_0[0]),.dout(n4218),.clk(gclk));
	jnot g03997(.din(w_n4218_0[1]),.dout(n4219),.clk(gclk));
	jor g03998(.dina(w_n4219_0[1]),.dinb(n4215),.dout(n4220),.clk(gclk));
	jand g03999(.dina(n4220),.dinb(n4115),.dout(n4221),.clk(gclk));
	jor g04000(.dina(w_n4221_0[2]),.dinb(w_n3835_0[2]),.dout(n4222),.clk(gclk));
	jxor g04001(.dina(w_n3815_0[2]),.dinb(w_n3646_0[2]),.dout(n4223),.clk(gclk));
	jnot g04002(.din(w_n4223_0[1]),.dout(n4224),.clk(gclk));
	jand g04003(.dina(n4224),.dinb(w_asqrt40_32[1]),.dout(n4225),.clk(gclk));
	jor g04004(.dina(w_n4225_0[1]),.dinb(w_n4222_0[1]),.dout(n4226),.clk(gclk));
	jand g04005(.dina(n4226),.dinb(w_n218_24[0]),.dout(n4227),.clk(gclk));
	jand g04006(.dina(w_n3955_49[1]),.dinb(w_n3646_0[1]),.dout(n4228),.clk(gclk));
	jand g04007(.dina(w_n4221_0[1]),.dinb(w_n3835_0[1]),.dout(n4229),.clk(gclk));
	jor g04008(.dina(w_n4229_0[2]),.dinb(w_n4228_0[1]),.dout(n4230),.clk(gclk));
	jand g04009(.dina(w_n3954_0[0]),.dinb(w_n3815_0[1]),.dout(n4231),.clk(gclk));
	jnot g04010(.din(n4231),.dout(n4232),.clk(gclk));
	jand g04011(.dina(w_n4223_0[0]),.dinb(w_asqrt63_44[0]),.dout(n4233),.clk(gclk));
	jand g04012(.dina(w_n4233_0[1]),.dinb(n4232),.dout(n4234),.clk(gclk));
	jor g04013(.dina(w_n4234_0[1]),.dinb(n4230),.dout(n4235),.clk(gclk));
	jor g04014(.dina(n4235),.dinb(w_n4227_0[1]),.dout(asqrt_fa_40),.clk(gclk));
	jor g04015(.dina(w_n4113_0[1]),.dinb(w_asqrt62_34[0]),.dout(n4237),.clk(gclk));
	jand g04016(.dina(w_n4218_0[0]),.dinb(n4237),.dout(n4238),.clk(gclk));
	jor g04017(.dina(n4238),.dinb(w_n4114_0[0]),.dout(n4239),.clk(gclk));
	jand g04018(.dina(w_n4239_0[1]),.dinb(w_n3834_0[1]),.dout(n4240),.clk(gclk));
	jnot g04019(.din(w_n4225_0[0]),.dout(n4241),.clk(gclk));
	jand g04020(.dina(n4241),.dinb(w_n4240_0[1]),.dout(n4242),.clk(gclk));
	jor g04021(.dina(n4242),.dinb(w_asqrt63_43[2]),.dout(n4243),.clk(gclk));
	jnot g04022(.din(w_n4228_0[0]),.dout(n4244),.clk(gclk));
	jor g04023(.dina(w_n4239_0[0]),.dinb(w_n3834_0[0]),.dout(n4245),.clk(gclk));
	jand g04024(.dina(w_n4245_0[2]),.dinb(n4244),.dout(n4246),.clk(gclk));
	jnot g04025(.din(w_n4234_0[0]),.dout(n4247),.clk(gclk));
	jand g04026(.dina(n4247),.dinb(n4246),.dout(n4248),.clk(gclk));
	jand g04027(.dina(n4248),.dinb(n4243),.dout(n4249),.clk(gclk));
	jxor g04028(.dina(w_n4113_0[0]),.dinb(w_n221_57[2]),.dout(n4250),.clk(gclk));
	jor g04029(.dina(n4250),.dinb(w_n4249_59[2]),.dout(n4251),.clk(gclk));
	jxor g04030(.dina(n4251),.dinb(w_n4219_0[0]),.dout(n4252),.clk(gclk));
	jnot g04031(.din(w_n4252_0[1]),.dout(n4253),.clk(gclk));
	jor g04032(.dina(w_n4249_59[1]),.dinb(w_n3837_1[0]),.dout(n4254),.clk(gclk));
	jnot g04033(.din(w_a76_0[2]),.dout(n4255),.clk(gclk));
	jnot g04034(.din(w_a77_0[1]),.dout(n4256),.clk(gclk));
	jand g04035(.dina(w_n4256_0[1]),.dinb(w_n4255_1[2]),.dout(n4257),.clk(gclk));
	jand g04036(.dina(w_n4257_0[2]),.dinb(w_n3837_0[2]),.dout(n4258),.clk(gclk));
	jnot g04037(.din(w_n4258_0[1]),.dout(n4259),.clk(gclk));
	jand g04038(.dina(n4259),.dinb(n4254),.dout(n4260),.clk(gclk));
	jor g04039(.dina(w_n4260_0[2]),.dinb(w_n3955_49[0]),.dout(n4261),.clk(gclk));
	jand g04040(.dina(w_n4260_0[1]),.dinb(w_n3955_48[2]),.dout(n4262),.clk(gclk));
	jor g04041(.dina(w_n4249_59[0]),.dinb(w_a78_1[0]),.dout(n4263),.clk(gclk));
	jand g04042(.dina(n4263),.dinb(w_a79_0[0]),.dout(n4264),.clk(gclk));
	jand g04043(.dina(w_asqrt39_30),.dinb(w_n3839_0[1]),.dout(n4265),.clk(gclk));
	jor g04044(.dina(n4265),.dinb(n4264),.dout(n4266),.clk(gclk));
	jor g04045(.dina(w_n4266_0[1]),.dinb(n4262),.dout(n4267),.clk(gclk));
	jand g04046(.dina(n4267),.dinb(w_n4261_0[1]),.dout(n4268),.clk(gclk));
	jor g04047(.dina(w_n4268_0[2]),.dinb(w_n3642_52[1]),.dout(n4269),.clk(gclk));
	jand g04048(.dina(w_n4268_0[1]),.dinb(w_n3642_52[0]),.dout(n4270),.clk(gclk));
	jnot g04049(.din(w_n3839_0[0]),.dout(n4271),.clk(gclk));
	jor g04050(.dina(w_n4249_58[2]),.dinb(n4271),.dout(n4272),.clk(gclk));
	jor g04051(.dina(w_n4229_0[1]),.dinb(w_n3955_48[1]),.dout(n4273),.clk(gclk));
	jor g04052(.dina(n4273),.dinb(w_n4227_0[0]),.dout(n4274),.clk(gclk));
	jor g04053(.dina(n4274),.dinb(w_n4233_0[0]),.dout(n4275),.clk(gclk));
	jand g04054(.dina(n4275),.dinb(w_n4272_0[1]),.dout(n4276),.clk(gclk));
	jxor g04055(.dina(n4276),.dinb(w_n3648_0[1]),.dout(n4277),.clk(gclk));
	jor g04056(.dina(w_n4277_0[2]),.dinb(n4270),.dout(n4278),.clk(gclk));
	jand g04057(.dina(n4278),.dinb(w_n4269_0[1]),.dout(n4279),.clk(gclk));
	jor g04058(.dina(w_n4279_0[2]),.dinb(w_n3368_49[2]),.dout(n4280),.clk(gclk));
	jand g04059(.dina(w_n4279_0[1]),.dinb(w_n3368_49[1]),.dout(n4281),.clk(gclk));
	jxor g04060(.dina(w_n3841_0[0]),.dinb(w_n3642_51[2]),.dout(n4282),.clk(gclk));
	jor g04061(.dina(n4282),.dinb(w_n4249_58[1]),.dout(n4283),.clk(gclk));
	jxor g04062(.dina(n4283),.dinb(w_n3957_0[0]),.dout(n4284),.clk(gclk));
	jor g04063(.dina(w_n4284_0[2]),.dinb(n4281),.dout(n4285),.clk(gclk));
	jand g04064(.dina(n4285),.dinb(w_n4280_0[1]),.dout(n4286),.clk(gclk));
	jor g04065(.dina(w_n4286_0[2]),.dinb(w_n3089_53[0]),.dout(n4287),.clk(gclk));
	jand g04066(.dina(w_n4286_0[1]),.dinb(w_n3089_52[2]),.dout(n4288),.clk(gclk));
	jxor g04067(.dina(w_n3959_0[0]),.dinb(w_n3368_49[0]),.dout(n4289),.clk(gclk));
	jor g04068(.dina(n4289),.dinb(w_n4249_58[0]),.dout(n4290),.clk(gclk));
	jxor g04069(.dina(n4290),.dinb(w_n3968_0[0]),.dout(n4291),.clk(gclk));
	jor g04070(.dina(w_n4291_0[2]),.dinb(n4288),.dout(n4292),.clk(gclk));
	jand g04071(.dina(n4292),.dinb(w_n4287_0[1]),.dout(n4293),.clk(gclk));
	jor g04072(.dina(w_n4293_0[2]),.dinb(w_n2833_50[2]),.dout(n4294),.clk(gclk));
	jand g04073(.dina(w_n4293_0[1]),.dinb(w_n2833_50[1]),.dout(n4295),.clk(gclk));
	jxor g04074(.dina(w_n3970_0[0]),.dinb(w_n3089_52[1]),.dout(n4296),.clk(gclk));
	jor g04075(.dina(n4296),.dinb(w_n4249_57[2]),.dout(n4297),.clk(gclk));
	jxor g04076(.dina(n4297),.dinb(w_n4150_0[0]),.dout(n4298),.clk(gclk));
	jnot g04077(.din(w_n4298_0[2]),.dout(n4299),.clk(gclk));
	jor g04078(.dina(n4299),.dinb(n4295),.dout(n4300),.clk(gclk));
	jand g04079(.dina(n4300),.dinb(w_n4294_0[1]),.dout(n4301),.clk(gclk));
	jor g04080(.dina(w_n4301_0[2]),.dinb(w_n2572_53[1]),.dout(n4302),.clk(gclk));
	jand g04081(.dina(w_n4301_0[1]),.dinb(w_n2572_53[0]),.dout(n4303),.clk(gclk));
	jxor g04082(.dina(w_n3977_0[0]),.dinb(w_n2833_50[0]),.dout(n4304),.clk(gclk));
	jor g04083(.dina(n4304),.dinb(w_n4249_57[1]),.dout(n4305),.clk(gclk));
	jxor g04084(.dina(n4305),.dinb(w_n3983_0[0]),.dout(n4306),.clk(gclk));
	jor g04085(.dina(w_n4306_0[2]),.dinb(n4303),.dout(n4307),.clk(gclk));
	jand g04086(.dina(n4307),.dinb(w_n4302_0[1]),.dout(n4308),.clk(gclk));
	jor g04087(.dina(w_n4308_0[2]),.dinb(w_n2345_51[1]),.dout(n4309),.clk(gclk));
	jand g04088(.dina(w_n4308_0[1]),.dinb(w_n2345_51[0]),.dout(n4310),.clk(gclk));
	jxor g04089(.dina(w_n3985_0[0]),.dinb(w_n2572_52[2]),.dout(n4311),.clk(gclk));
	jor g04090(.dina(n4311),.dinb(w_n4249_57[0]),.dout(n4312),.clk(gclk));
	jxor g04091(.dina(n4312),.dinb(w_n4157_0[0]),.dout(n4313),.clk(gclk));
	jnot g04092(.din(w_n4313_0[2]),.dout(n4314),.clk(gclk));
	jor g04093(.dina(n4314),.dinb(n4310),.dout(n4315),.clk(gclk));
	jand g04094(.dina(n4315),.dinb(w_n4309_0[1]),.dout(n4316),.clk(gclk));
	jor g04095(.dina(w_n4316_0[2]),.dinb(w_n2108_54[0]),.dout(n4317),.clk(gclk));
	jand g04096(.dina(w_n4316_0[1]),.dinb(w_n2108_53[2]),.dout(n4318),.clk(gclk));
	jxor g04097(.dina(w_n3992_0[0]),.dinb(w_n2345_50[2]),.dout(n4319),.clk(gclk));
	jor g04098(.dina(n4319),.dinb(w_n4249_56[2]),.dout(n4320),.clk(gclk));
	jxor g04099(.dina(n4320),.dinb(w_n3998_0[0]),.dout(n4321),.clk(gclk));
	jor g04100(.dina(w_n4321_0[2]),.dinb(n4318),.dout(n4322),.clk(gclk));
	jand g04101(.dina(n4322),.dinb(w_n4317_0[1]),.dout(n4323),.clk(gclk));
	jor g04102(.dina(w_n4323_0[2]),.dinb(w_n1912_52[1]),.dout(n4324),.clk(gclk));
	jand g04103(.dina(w_n4323_0[1]),.dinb(w_n1912_52[0]),.dout(n4325),.clk(gclk));
	jxor g04104(.dina(w_n4000_0[0]),.dinb(w_n2108_53[1]),.dout(n4326),.clk(gclk));
	jor g04105(.dina(n4326),.dinb(w_n4249_56[1]),.dout(n4327),.clk(gclk));
	jxor g04106(.dina(n4327),.dinb(w_n4164_0[0]),.dout(n4328),.clk(gclk));
	jnot g04107(.din(w_n4328_0[2]),.dout(n4329),.clk(gclk));
	jor g04108(.dina(n4329),.dinb(n4325),.dout(n4330),.clk(gclk));
	jand g04109(.dina(n4330),.dinb(w_n4324_0[1]),.dout(n4331),.clk(gclk));
	jor g04110(.dina(w_n4331_0[2]),.dinb(w_n1699_54[2]),.dout(n4332),.clk(gclk));
	jand g04111(.dina(w_n4331_0[1]),.dinb(w_n1699_54[1]),.dout(n4333),.clk(gclk));
	jxor g04112(.dina(w_n4007_0[0]),.dinb(w_n1912_51[2]),.dout(n4334),.clk(gclk));
	jor g04113(.dina(n4334),.dinb(w_n4249_56[0]),.dout(n4335),.clk(gclk));
	jxor g04114(.dina(n4335),.dinb(w_n4168_0[0]),.dout(n4336),.clk(gclk));
	jnot g04115(.din(w_n4336_0[2]),.dout(n4337),.clk(gclk));
	jor g04116(.dina(n4337),.dinb(n4333),.dout(n4338),.clk(gclk));
	jand g04117(.dina(n4338),.dinb(w_n4332_0[1]),.dout(n4339),.clk(gclk));
	jor g04118(.dina(w_n4339_0[2]),.dinb(w_n1516_53[0]),.dout(n4340),.clk(gclk));
	jand g04119(.dina(w_n4339_0[1]),.dinb(w_n1516_52[2]),.dout(n4341),.clk(gclk));
	jxor g04120(.dina(w_n4014_0[0]),.dinb(w_n1699_54[0]),.dout(n4342),.clk(gclk));
	jor g04121(.dina(n4342),.dinb(w_n4249_55[2]),.dout(n4343),.clk(gclk));
	jxor g04122(.dina(n4343),.dinb(w_n4020_0[0]),.dout(n4344),.clk(gclk));
	jor g04123(.dina(w_n4344_0[2]),.dinb(n4341),.dout(n4345),.clk(gclk));
	jand g04124(.dina(n4345),.dinb(w_n4340_0[1]),.dout(n4346),.clk(gclk));
	jor g04125(.dina(w_n4346_0[2]),.dinb(w_n1332_54[2]),.dout(n4347),.clk(gclk));
	jand g04126(.dina(w_n4346_0[1]),.dinb(w_n1332_54[1]),.dout(n4348),.clk(gclk));
	jxor g04127(.dina(w_n4022_0[0]),.dinb(w_n1516_52[1]),.dout(n4349),.clk(gclk));
	jor g04128(.dina(n4349),.dinb(w_n4249_55[1]),.dout(n4350),.clk(gclk));
	jxor g04129(.dina(n4350),.dinb(w_n4028_0[0]),.dout(n4351),.clk(gclk));
	jor g04130(.dina(w_n4351_0[2]),.dinb(n4348),.dout(n4352),.clk(gclk));
	jand g04131(.dina(n4352),.dinb(w_n4347_0[1]),.dout(n4353),.clk(gclk));
	jor g04132(.dina(w_n4353_0[2]),.dinb(w_n1173_53[2]),.dout(n4354),.clk(gclk));
	jand g04133(.dina(w_n4353_0[1]),.dinb(w_n1173_53[1]),.dout(n4355),.clk(gclk));
	jxor g04134(.dina(w_n4030_0[0]),.dinb(w_n1332_54[0]),.dout(n4356),.clk(gclk));
	jor g04135(.dina(n4356),.dinb(w_n4249_55[0]),.dout(n4357),.clk(gclk));
	jxor g04136(.dina(n4357),.dinb(w_n4178_0[0]),.dout(n4358),.clk(gclk));
	jnot g04137(.din(w_n4358_0[2]),.dout(n4359),.clk(gclk));
	jor g04138(.dina(n4359),.dinb(n4355),.dout(n4360),.clk(gclk));
	jand g04139(.dina(n4360),.dinb(w_n4354_0[1]),.dout(n4361),.clk(gclk));
	jor g04140(.dina(w_n4361_0[2]),.dinb(w_n1008_55[2]),.dout(n4362),.clk(gclk));
	jand g04141(.dina(w_n4361_0[1]),.dinb(w_n1008_55[1]),.dout(n4363),.clk(gclk));
	jxor g04142(.dina(w_n4037_0[0]),.dinb(w_n1173_53[0]),.dout(n4364),.clk(gclk));
	jor g04143(.dina(n4364),.dinb(w_n4249_54[2]),.dout(n4365),.clk(gclk));
	jxor g04144(.dina(n4365),.dinb(w_n4043_0[0]),.dout(n4366),.clk(gclk));
	jor g04145(.dina(w_n4366_0[2]),.dinb(n4363),.dout(n4367),.clk(gclk));
	jand g04146(.dina(n4367),.dinb(w_n4362_0[1]),.dout(n4368),.clk(gclk));
	jor g04147(.dina(w_n4368_0[2]),.dinb(w_n884_54[2]),.dout(n4369),.clk(gclk));
	jand g04148(.dina(w_n4368_0[1]),.dinb(w_n884_54[1]),.dout(n4370),.clk(gclk));
	jxor g04149(.dina(w_n4045_0[0]),.dinb(w_n1008_55[0]),.dout(n4371),.clk(gclk));
	jor g04150(.dina(n4371),.dinb(w_n4249_54[1]),.dout(n4372),.clk(gclk));
	jxor g04151(.dina(n4372),.dinb(w_n4185_0[0]),.dout(n4373),.clk(gclk));
	jnot g04152(.din(w_n4373_0[2]),.dout(n4374),.clk(gclk));
	jor g04153(.dina(n4374),.dinb(n4370),.dout(n4375),.clk(gclk));
	jand g04154(.dina(n4375),.dinb(w_n4369_0[1]),.dout(n4376),.clk(gclk));
	jor g04155(.dina(w_n4376_0[2]),.dinb(w_n743_55[2]),.dout(n4377),.clk(gclk));
	jand g04156(.dina(w_n4376_0[1]),.dinb(w_n743_55[1]),.dout(n4378),.clk(gclk));
	jxor g04157(.dina(w_n4052_0[0]),.dinb(w_n884_54[0]),.dout(n4379),.clk(gclk));
	jor g04158(.dina(n4379),.dinb(w_n4249_54[0]),.dout(n4380),.clk(gclk));
	jxor g04159(.dina(n4380),.dinb(w_n4058_0[0]),.dout(n4381),.clk(gclk));
	jor g04160(.dina(w_n4381_0[2]),.dinb(n4378),.dout(n4382),.clk(gclk));
	jand g04161(.dina(n4382),.dinb(w_n4377_0[1]),.dout(n4383),.clk(gclk));
	jor g04162(.dina(w_n4383_0[2]),.dinb(w_n635_55[2]),.dout(n4384),.clk(gclk));
	jand g04163(.dina(w_n4383_0[1]),.dinb(w_n635_55[1]),.dout(n4385),.clk(gclk));
	jxor g04164(.dina(w_n4060_0[0]),.dinb(w_n743_55[0]),.dout(n4386),.clk(gclk));
	jor g04165(.dina(n4386),.dinb(w_n4249_53[2]),.dout(n4387),.clk(gclk));
	jxor g04166(.dina(n4387),.dinb(w_n4192_0[0]),.dout(n4388),.clk(gclk));
	jnot g04167(.din(w_n4388_0[2]),.dout(n4389),.clk(gclk));
	jor g04168(.dina(n4389),.dinb(n4385),.dout(n4390),.clk(gclk));
	jand g04169(.dina(n4390),.dinb(w_n4384_0[1]),.dout(n4391),.clk(gclk));
	jor g04170(.dina(w_n4391_0[2]),.dinb(w_n515_56[2]),.dout(n4392),.clk(gclk));
	jand g04171(.dina(w_n4391_0[1]),.dinb(w_n515_56[1]),.dout(n4393),.clk(gclk));
	jxor g04172(.dina(w_n4067_0[0]),.dinb(w_n635_55[0]),.dout(n4394),.clk(gclk));
	jor g04173(.dina(n4394),.dinb(w_n4249_53[1]),.dout(n4395),.clk(gclk));
	jxor g04174(.dina(n4395),.dinb(w_n4073_0[0]),.dout(n4396),.clk(gclk));
	jor g04175(.dina(w_n4396_0[2]),.dinb(n4393),.dout(n4397),.clk(gclk));
	jand g04176(.dina(n4397),.dinb(w_n4392_0[1]),.dout(n4398),.clk(gclk));
	jor g04177(.dina(w_n4398_0[2]),.dinb(w_n443_56[2]),.dout(n4399),.clk(gclk));
	jand g04178(.dina(w_n4398_0[1]),.dinb(w_n443_56[1]),.dout(n4400),.clk(gclk));
	jxor g04179(.dina(w_n4075_0[0]),.dinb(w_n515_56[0]),.dout(n4401),.clk(gclk));
	jor g04180(.dina(n4401),.dinb(w_n4249_53[0]),.dout(n4402),.clk(gclk));
	jxor g04181(.dina(n4402),.dinb(w_n4199_0[0]),.dout(n4403),.clk(gclk));
	jnot g04182(.din(w_n4403_0[2]),.dout(n4404),.clk(gclk));
	jor g04183(.dina(n4404),.dinb(n4400),.dout(n4405),.clk(gclk));
	jand g04184(.dina(n4405),.dinb(w_n4399_0[1]),.dout(n4406),.clk(gclk));
	jor g04185(.dina(w_n4406_0[2]),.dinb(w_n352_57[0]),.dout(n4407),.clk(gclk));
	jand g04186(.dina(w_n4406_0[1]),.dinb(w_n352_56[2]),.dout(n4408),.clk(gclk));
	jxor g04187(.dina(w_n4082_0[0]),.dinb(w_n443_56[0]),.dout(n4409),.clk(gclk));
	jor g04188(.dina(n4409),.dinb(w_n4249_52[2]),.dout(n4410),.clk(gclk));
	jxor g04189(.dina(n4410),.dinb(w_n4088_0[0]),.dout(n4411),.clk(gclk));
	jor g04190(.dina(w_n4411_0[2]),.dinb(n4408),.dout(n4412),.clk(gclk));
	jand g04191(.dina(n4412),.dinb(w_n4407_0[1]),.dout(n4413),.clk(gclk));
	jor g04192(.dina(w_n4413_0[2]),.dinb(w_n294_57[1]),.dout(n4414),.clk(gclk));
	jand g04193(.dina(w_n4413_0[1]),.dinb(w_n294_57[0]),.dout(n4415),.clk(gclk));
	jxor g04194(.dina(w_n4090_0[0]),.dinb(w_n352_56[1]),.dout(n4416),.clk(gclk));
	jor g04195(.dina(n4416),.dinb(w_n4249_52[1]),.dout(n4417),.clk(gclk));
	jxor g04196(.dina(n4417),.dinb(w_n4206_0[0]),.dout(n4418),.clk(gclk));
	jnot g04197(.din(w_n4418_0[2]),.dout(n4419),.clk(gclk));
	jor g04198(.dina(n4419),.dinb(n4415),.dout(n4420),.clk(gclk));
	jand g04199(.dina(n4420),.dinb(w_n4414_0[1]),.dout(n4421),.clk(gclk));
	jor g04200(.dina(w_n4421_0[2]),.dinb(w_n239_57[1]),.dout(n4422),.clk(gclk));
	jand g04201(.dina(w_n4421_0[1]),.dinb(w_n239_57[0]),.dout(n4423),.clk(gclk));
	jxor g04202(.dina(w_n4097_0[0]),.dinb(w_n294_56[2]),.dout(n4424),.clk(gclk));
	jor g04203(.dina(n4424),.dinb(w_n4249_52[0]),.dout(n4425),.clk(gclk));
	jxor g04204(.dina(n4425),.dinb(w_n4103_0[0]),.dout(n4426),.clk(gclk));
	jor g04205(.dina(w_n4426_0[2]),.dinb(n4423),.dout(n4427),.clk(gclk));
	jand g04206(.dina(n4427),.dinb(w_n4422_0[1]),.dout(n4428),.clk(gclk));
	jor g04207(.dina(w_n4428_0[2]),.dinb(w_n221_57[1]),.dout(n4429),.clk(gclk));
	jand g04208(.dina(w_n4428_0[1]),.dinb(w_n221_57[0]),.dout(n4430),.clk(gclk));
	jxor g04209(.dina(w_n4105_0[0]),.dinb(w_n239_56[2]),.dout(n4431),.clk(gclk));
	jor g04210(.dina(n4431),.dinb(w_n4249_51[2]),.dout(n4432),.clk(gclk));
	jxor g04211(.dina(n4432),.dinb(w_n4111_0[0]),.dout(n4433),.clk(gclk));
	jor g04212(.dina(w_n4433_0[1]),.dinb(n4430),.dout(n4434),.clk(gclk));
	jand g04213(.dina(n4434),.dinb(w_n4429_0[1]),.dout(n4435),.clk(gclk));
	jor g04214(.dina(w_n4435_0[2]),.dinb(w_n4253_0[2]),.dout(n4436),.clk(gclk));
	jand g04215(.dina(w_asqrt39_29[2]),.dinb(w_n4240_0[0]),.dout(n4437),.clk(gclk));
	jor g04216(.dina(w_n4437_0[1]),.dinb(w_n4436_0[1]),.dout(n4438),.clk(gclk));
	jor g04217(.dina(n4438),.dinb(w_n4229_0[0]),.dout(n4439),.clk(gclk));
	jand g04218(.dina(n4439),.dinb(w_n218_23[2]),.dout(n4440),.clk(gclk));
	jand g04219(.dina(w_n4249_51[1]),.dinb(w_n3835_0[0]),.dout(n4441),.clk(gclk));
	jand g04220(.dina(w_n4435_0[1]),.dinb(w_n4253_0[1]),.dout(n4442),.clk(gclk));
	jor g04221(.dina(w_n4442_0[2]),.dinb(n4441),.dout(n4443),.clk(gclk));
	jand g04222(.dina(w_n4249_51[0]),.dinb(w_n4221_0[0]),.dout(n4444),.clk(gclk));
	jand g04223(.dina(w_n4222_0[0]),.dinb(w_asqrt63_43[1]),.dout(n4445),.clk(gclk));
	jand g04224(.dina(n4445),.dinb(w_n4245_0[1]),.dout(n4446),.clk(gclk));
	jnot g04225(.din(n4446),.dout(n4447),.clk(gclk));
	jor g04226(.dina(w_n4447_0[1]),.dinb(n4444),.dout(n4448),.clk(gclk));
	jnot g04227(.din(n4448),.dout(n4449),.clk(gclk));
	jor g04228(.dina(n4449),.dinb(n4443),.dout(n4450),.clk(gclk));
	jor g04229(.dina(w_n4450_0[1]),.dinb(n4440),.dout(asqrt_fa_39),.clk(gclk));
	jnot g04230(.din(w_n4433_0[0]),.dout(n4452),.clk(gclk));
	jxor g04231(.dina(w_n4428_0[0]),.dinb(w_n221_56[2]),.dout(n4453),.clk(gclk));
	jand g04232(.dina(n4453),.dinb(w_asqrt38_40),.dout(n4454),.clk(gclk));
	jxor g04233(.dina(n4454),.dinb(w_n4452_0[1]),.dout(n4455),.clk(gclk));
	jand g04234(.dina(w_asqrt38_39[2]),.dinb(w_a76_0[1]),.dout(n4456),.clk(gclk));
	jnot g04235(.din(w_a74_1[1]),.dout(n4457),.clk(gclk));
	jnot g04236(.din(w_a75_0[1]),.dout(n4458),.clk(gclk));
	jand g04237(.dina(w_n4458_0[1]),.dinb(w_n4457_1[1]),.dout(n4459),.clk(gclk));
	jand g04238(.dina(w_n4459_0[2]),.dinb(w_n4255_1[1]),.dout(n4460),.clk(gclk));
	jor g04239(.dina(w_n4460_0[1]),.dinb(n4456),.dout(n4461),.clk(gclk));
	jand g04240(.dina(w_n4461_0[2]),.dinb(w_asqrt39_29[1]),.dout(n4462),.clk(gclk));
	jor g04241(.dina(w_n4461_0[1]),.dinb(w_asqrt39_29[0]),.dout(n4463),.clk(gclk));
	jand g04242(.dina(w_asqrt38_39[1]),.dinb(w_n4255_1[0]),.dout(n4464),.clk(gclk));
	jor g04243(.dina(n4464),.dinb(w_n4256_0[0]),.dout(n4465),.clk(gclk));
	jnot g04244(.din(w_n4257_0[1]),.dout(n4466),.clk(gclk));
	jnot g04245(.din(w_n4429_0[0]),.dout(n4467),.clk(gclk));
	jnot g04246(.din(w_n4422_0[0]),.dout(n4468),.clk(gclk));
	jnot g04247(.din(w_n4414_0[0]),.dout(n4469),.clk(gclk));
	jnot g04248(.din(w_n4407_0[0]),.dout(n4470),.clk(gclk));
	jnot g04249(.din(w_n4399_0[0]),.dout(n4471),.clk(gclk));
	jnot g04250(.din(w_n4392_0[0]),.dout(n4472),.clk(gclk));
	jnot g04251(.din(w_n4384_0[0]),.dout(n4473),.clk(gclk));
	jnot g04252(.din(w_n4377_0[0]),.dout(n4474),.clk(gclk));
	jnot g04253(.din(w_n4369_0[0]),.dout(n4475),.clk(gclk));
	jnot g04254(.din(w_n4362_0[0]),.dout(n4476),.clk(gclk));
	jnot g04255(.din(w_n4354_0[0]),.dout(n4477),.clk(gclk));
	jnot g04256(.din(w_n4347_0[0]),.dout(n4478),.clk(gclk));
	jnot g04257(.din(w_n4340_0[0]),.dout(n4479),.clk(gclk));
	jnot g04258(.din(w_n4332_0[0]),.dout(n4480),.clk(gclk));
	jnot g04259(.din(w_n4324_0[0]),.dout(n4481),.clk(gclk));
	jnot g04260(.din(w_n4317_0[0]),.dout(n4482),.clk(gclk));
	jnot g04261(.din(w_n4309_0[0]),.dout(n4483),.clk(gclk));
	jnot g04262(.din(w_n4302_0[0]),.dout(n4484),.clk(gclk));
	jnot g04263(.din(w_n4294_0[0]),.dout(n4485),.clk(gclk));
	jnot g04264(.din(w_n4287_0[0]),.dout(n4486),.clk(gclk));
	jnot g04265(.din(w_n4280_0[0]),.dout(n4487),.clk(gclk));
	jnot g04266(.din(w_n4269_0[0]),.dout(n4488),.clk(gclk));
	jnot g04267(.din(w_n4261_0[0]),.dout(n4489),.clk(gclk));
	jand g04268(.dina(w_asqrt39_28[2]),.dinb(w_a78_0[2]),.dout(n4490),.clk(gclk));
	jor g04269(.dina(w_n4258_0[0]),.dinb(n4490),.dout(n4491),.clk(gclk));
	jor g04270(.dina(n4491),.dinb(w_asqrt40_32[0]),.dout(n4492),.clk(gclk));
	jand g04271(.dina(w_asqrt39_28[1]),.dinb(w_n3837_0[1]),.dout(n4493),.clk(gclk));
	jor g04272(.dina(n4493),.dinb(w_n3838_0[0]),.dout(n4494),.clk(gclk));
	jand g04273(.dina(w_n4272_0[0]),.dinb(n4494),.dout(n4495),.clk(gclk));
	jand g04274(.dina(n4495),.dinb(n4492),.dout(n4496),.clk(gclk));
	jor g04275(.dina(n4496),.dinb(n4489),.dout(n4497),.clk(gclk));
	jor g04276(.dina(n4497),.dinb(w_asqrt41_29[0]),.dout(n4498),.clk(gclk));
	jnot g04277(.din(w_n4277_0[1]),.dout(n4499),.clk(gclk));
	jand g04278(.dina(n4499),.dinb(n4498),.dout(n4500),.clk(gclk));
	jor g04279(.dina(n4500),.dinb(n4488),.dout(n4501),.clk(gclk));
	jor g04280(.dina(n4501),.dinb(w_asqrt42_32[1]),.dout(n4502),.clk(gclk));
	jnot g04281(.din(w_n4284_0[1]),.dout(n4503),.clk(gclk));
	jand g04282(.dina(n4503),.dinb(n4502),.dout(n4504),.clk(gclk));
	jor g04283(.dina(n4504),.dinb(n4487),.dout(n4505),.clk(gclk));
	jor g04284(.dina(n4505),.dinb(w_asqrt43_29[1]),.dout(n4506),.clk(gclk));
	jnot g04285(.din(w_n4291_0[1]),.dout(n4507),.clk(gclk));
	jand g04286(.dina(n4507),.dinb(n4506),.dout(n4508),.clk(gclk));
	jor g04287(.dina(n4508),.dinb(n4486),.dout(n4509),.clk(gclk));
	jor g04288(.dina(n4509),.dinb(w_asqrt44_32[1]),.dout(n4510),.clk(gclk));
	jand g04289(.dina(w_n4298_0[1]),.dinb(n4510),.dout(n4511),.clk(gclk));
	jor g04290(.dina(n4511),.dinb(n4485),.dout(n4512),.clk(gclk));
	jor g04291(.dina(n4512),.dinb(w_asqrt45_30[0]),.dout(n4513),.clk(gclk));
	jnot g04292(.din(w_n4306_0[1]),.dout(n4514),.clk(gclk));
	jand g04293(.dina(n4514),.dinb(n4513),.dout(n4515),.clk(gclk));
	jor g04294(.dina(n4515),.dinb(n4484),.dout(n4516),.clk(gclk));
	jor g04295(.dina(n4516),.dinb(w_asqrt46_32[1]),.dout(n4517),.clk(gclk));
	jand g04296(.dina(w_n4313_0[1]),.dinb(n4517),.dout(n4518),.clk(gclk));
	jor g04297(.dina(n4518),.dinb(n4483),.dout(n4519),.clk(gclk));
	jor g04298(.dina(n4519),.dinb(w_asqrt47_30[2]),.dout(n4520),.clk(gclk));
	jnot g04299(.din(w_n4321_0[1]),.dout(n4521),.clk(gclk));
	jand g04300(.dina(n4521),.dinb(n4520),.dout(n4522),.clk(gclk));
	jor g04301(.dina(n4522),.dinb(n4482),.dout(n4523),.clk(gclk));
	jor g04302(.dina(n4523),.dinb(w_asqrt48_32[2]),.dout(n4524),.clk(gclk));
	jand g04303(.dina(w_n4328_0[1]),.dinb(n4524),.dout(n4525),.clk(gclk));
	jor g04304(.dina(n4525),.dinb(n4481),.dout(n4526),.clk(gclk));
	jor g04305(.dina(n4526),.dinb(w_asqrt49_31[0]),.dout(n4527),.clk(gclk));
	jand g04306(.dina(w_n4336_0[1]),.dinb(n4527),.dout(n4528),.clk(gclk));
	jor g04307(.dina(n4528),.dinb(n4480),.dout(n4529),.clk(gclk));
	jor g04308(.dina(n4529),.dinb(w_asqrt50_33[0]),.dout(n4530),.clk(gclk));
	jnot g04309(.din(w_n4344_0[1]),.dout(n4531),.clk(gclk));
	jand g04310(.dina(n4531),.dinb(n4530),.dout(n4532),.clk(gclk));
	jor g04311(.dina(n4532),.dinb(n4479),.dout(n4533),.clk(gclk));
	jor g04312(.dina(n4533),.dinb(w_asqrt51_31[1]),.dout(n4534),.clk(gclk));
	jnot g04313(.din(w_n4351_0[1]),.dout(n4535),.clk(gclk));
	jand g04314(.dina(n4535),.dinb(n4534),.dout(n4536),.clk(gclk));
	jor g04315(.dina(n4536),.dinb(n4478),.dout(n4537),.clk(gclk));
	jor g04316(.dina(n4537),.dinb(w_asqrt52_33[0]),.dout(n4538),.clk(gclk));
	jand g04317(.dina(w_n4358_0[1]),.dinb(n4538),.dout(n4539),.clk(gclk));
	jor g04318(.dina(n4539),.dinb(n4477),.dout(n4540),.clk(gclk));
	jor g04319(.dina(n4540),.dinb(w_asqrt53_32[0]),.dout(n4541),.clk(gclk));
	jnot g04320(.din(w_n4366_0[1]),.dout(n4542),.clk(gclk));
	jand g04321(.dina(n4542),.dinb(n4541),.dout(n4543),.clk(gclk));
	jor g04322(.dina(n4543),.dinb(n4476),.dout(n4544),.clk(gclk));
	jor g04323(.dina(n4544),.dinb(w_asqrt54_33[0]),.dout(n4545),.clk(gclk));
	jand g04324(.dina(w_n4373_0[1]),.dinb(n4545),.dout(n4546),.clk(gclk));
	jor g04325(.dina(n4546),.dinb(n4475),.dout(n4547),.clk(gclk));
	jor g04326(.dina(n4547),.dinb(w_asqrt55_32[1]),.dout(n4548),.clk(gclk));
	jnot g04327(.din(w_n4381_0[1]),.dout(n4549),.clk(gclk));
	jand g04328(.dina(n4549),.dinb(n4548),.dout(n4550),.clk(gclk));
	jor g04329(.dina(n4550),.dinb(n4474),.dout(n4551),.clk(gclk));
	jor g04330(.dina(n4551),.dinb(w_asqrt56_33[1]),.dout(n4552),.clk(gclk));
	jand g04331(.dina(w_n4388_0[1]),.dinb(n4552),.dout(n4553),.clk(gclk));
	jor g04332(.dina(n4553),.dinb(n4473),.dout(n4554),.clk(gclk));
	jor g04333(.dina(n4554),.dinb(w_asqrt57_33[0]),.dout(n4555),.clk(gclk));
	jnot g04334(.din(w_n4396_0[1]),.dout(n4556),.clk(gclk));
	jand g04335(.dina(n4556),.dinb(n4555),.dout(n4557),.clk(gclk));
	jor g04336(.dina(n4557),.dinb(n4472),.dout(n4558),.clk(gclk));
	jor g04337(.dina(n4558),.dinb(w_asqrt58_33[2]),.dout(n4559),.clk(gclk));
	jand g04338(.dina(w_n4403_0[1]),.dinb(n4559),.dout(n4560),.clk(gclk));
	jor g04339(.dina(n4560),.dinb(n4471),.dout(n4561),.clk(gclk));
	jor g04340(.dina(n4561),.dinb(w_asqrt59_33[1]),.dout(n4562),.clk(gclk));
	jnot g04341(.din(w_n4411_0[1]),.dout(n4563),.clk(gclk));
	jand g04342(.dina(n4563),.dinb(n4562),.dout(n4564),.clk(gclk));
	jor g04343(.dina(n4564),.dinb(n4470),.dout(n4565),.clk(gclk));
	jor g04344(.dina(n4565),.dinb(w_asqrt60_33[2]),.dout(n4566),.clk(gclk));
	jand g04345(.dina(w_n4418_0[1]),.dinb(n4566),.dout(n4567),.clk(gclk));
	jor g04346(.dina(n4567),.dinb(n4469),.dout(n4568),.clk(gclk));
	jor g04347(.dina(n4568),.dinb(w_asqrt61_33[2]),.dout(n4569),.clk(gclk));
	jnot g04348(.din(w_n4426_0[1]),.dout(n4570),.clk(gclk));
	jand g04349(.dina(n4570),.dinb(n4569),.dout(n4571),.clk(gclk));
	jor g04350(.dina(n4571),.dinb(n4468),.dout(n4572),.clk(gclk));
	jor g04351(.dina(n4572),.dinb(w_asqrt62_33[2]),.dout(n4573),.clk(gclk));
	jand g04352(.dina(w_n4452_0[0]),.dinb(n4573),.dout(n4574),.clk(gclk));
	jor g04353(.dina(n4574),.dinb(n4467),.dout(n4575),.clk(gclk));
	jand g04354(.dina(n4575),.dinb(w_n4252_0[0]),.dout(n4576),.clk(gclk));
	jnot g04355(.din(w_n4437_0[0]),.dout(n4577),.clk(gclk));
	jand g04356(.dina(n4577),.dinb(w_n4576_0[1]),.dout(n4578),.clk(gclk));
	jand g04357(.dina(n4578),.dinb(w_n4245_0[0]),.dout(n4579),.clk(gclk));
	jor g04358(.dina(n4579),.dinb(w_asqrt63_43[0]),.dout(n4580),.clk(gclk));
	jnot g04359(.din(w_n4450_0[0]),.dout(n4581),.clk(gclk));
	jand g04360(.dina(n4581),.dinb(w_n4580_0[1]),.dout(n4582),.clk(gclk));
	jor g04361(.dina(w_n4582_48[1]),.dinb(n4466),.dout(n4583),.clk(gclk));
	jand g04362(.dina(n4583),.dinb(n4465),.dout(n4584),.clk(gclk));
	jand g04363(.dina(n4584),.dinb(n4463),.dout(n4585),.clk(gclk));
	jor g04364(.dina(n4585),.dinb(w_n4462_0[1]),.dout(n4586),.clk(gclk));
	jand g04365(.dina(w_n4586_0[2]),.dinb(w_asqrt40_31[2]),.dout(n4587),.clk(gclk));
	jor g04366(.dina(w_n4586_0[1]),.dinb(w_asqrt40_31[1]),.dout(n4588),.clk(gclk));
	jand g04367(.dina(w_asqrt38_39[0]),.dinb(w_n4257_0[0]),.dout(n4589),.clk(gclk));
	jnot g04368(.din(w_n4442_0[1]),.dout(n4590),.clk(gclk));
	jand g04369(.dina(w_n4447_0[0]),.dinb(w_asqrt39_28[0]),.dout(n4591),.clk(gclk));
	jand g04370(.dina(n4591),.dinb(w_n4590_0[1]),.dout(n4592),.clk(gclk));
	jand g04371(.dina(n4592),.dinb(w_n4580_0[0]),.dout(n4593),.clk(gclk));
	jor g04372(.dina(n4593),.dinb(w_n4589_0[1]),.dout(n4594),.clk(gclk));
	jxor g04373(.dina(n4594),.dinb(w_a78_0[1]),.dout(n4595),.clk(gclk));
	jnot g04374(.din(w_n4595_0[2]),.dout(n4596),.clk(gclk));
	jand g04375(.dina(n4596),.dinb(n4588),.dout(n4597),.clk(gclk));
	jor g04376(.dina(n4597),.dinb(w_n4587_0[1]),.dout(n4598),.clk(gclk));
	jand g04377(.dina(w_n4598_0[2]),.dinb(w_asqrt41_28[2]),.dout(n4599),.clk(gclk));
	jor g04378(.dina(w_n4598_0[1]),.dinb(w_asqrt41_28[1]),.dout(n4600),.clk(gclk));
	jxor g04379(.dina(w_n4260_0[0]),.dinb(w_n3955_48[0]),.dout(n4601),.clk(gclk));
	jand g04380(.dina(n4601),.dinb(w_asqrt38_38[2]),.dout(n4602),.clk(gclk));
	jxor g04381(.dina(n4602),.dinb(w_n4266_0[0]),.dout(n4603),.clk(gclk));
	jnot g04382(.din(w_n4603_0[1]),.dout(n4604),.clk(gclk));
	jand g04383(.dina(w_n4604_0[1]),.dinb(n4600),.dout(n4605),.clk(gclk));
	jor g04384(.dina(n4605),.dinb(w_n4599_0[1]),.dout(n4606),.clk(gclk));
	jand g04385(.dina(w_n4606_0[2]),.dinb(w_asqrt42_32[0]),.dout(n4607),.clk(gclk));
	jor g04386(.dina(w_n4606_0[1]),.dinb(w_asqrt42_31[2]),.dout(n4608),.clk(gclk));
	jxor g04387(.dina(w_n4268_0[0]),.dinb(w_n3642_51[1]),.dout(n4609),.clk(gclk));
	jand g04388(.dina(n4609),.dinb(w_asqrt38_38[1]),.dout(n4610),.clk(gclk));
	jxor g04389(.dina(n4610),.dinb(w_n4277_0[0]),.dout(n4611),.clk(gclk));
	jnot g04390(.din(w_n4611_0[1]),.dout(n4612),.clk(gclk));
	jand g04391(.dina(w_n4612_0[1]),.dinb(n4608),.dout(n4613),.clk(gclk));
	jor g04392(.dina(n4613),.dinb(w_n4607_0[1]),.dout(n4614),.clk(gclk));
	jand g04393(.dina(w_n4614_0[2]),.dinb(w_asqrt43_29[0]),.dout(n4615),.clk(gclk));
	jor g04394(.dina(w_n4614_0[1]),.dinb(w_asqrt43_28[2]),.dout(n4616),.clk(gclk));
	jxor g04395(.dina(w_n4279_0[0]),.dinb(w_n3368_48[2]),.dout(n4617),.clk(gclk));
	jand g04396(.dina(n4617),.dinb(w_asqrt38_38[0]),.dout(n4618),.clk(gclk));
	jxor g04397(.dina(n4618),.dinb(w_n4284_0[0]),.dout(n4619),.clk(gclk));
	jnot g04398(.din(w_n4619_0[1]),.dout(n4620),.clk(gclk));
	jand g04399(.dina(w_n4620_0[1]),.dinb(n4616),.dout(n4621),.clk(gclk));
	jor g04400(.dina(n4621),.dinb(w_n4615_0[1]),.dout(n4622),.clk(gclk));
	jand g04401(.dina(w_n4622_0[2]),.dinb(w_asqrt44_32[0]),.dout(n4623),.clk(gclk));
	jor g04402(.dina(w_n4622_0[1]),.dinb(w_asqrt44_31[2]),.dout(n4624),.clk(gclk));
	jxor g04403(.dina(w_n4286_0[0]),.dinb(w_n3089_52[0]),.dout(n4625),.clk(gclk));
	jand g04404(.dina(n4625),.dinb(w_asqrt38_37[2]),.dout(n4626),.clk(gclk));
	jxor g04405(.dina(n4626),.dinb(w_n4291_0[0]),.dout(n4627),.clk(gclk));
	jnot g04406(.din(w_n4627_0[1]),.dout(n4628),.clk(gclk));
	jand g04407(.dina(w_n4628_0[1]),.dinb(n4624),.dout(n4629),.clk(gclk));
	jor g04408(.dina(n4629),.dinb(w_n4623_0[1]),.dout(n4630),.clk(gclk));
	jand g04409(.dina(w_n4630_0[2]),.dinb(w_asqrt45_29[2]),.dout(n4631),.clk(gclk));
	jor g04410(.dina(w_n4630_0[1]),.dinb(w_asqrt45_29[1]),.dout(n4632),.clk(gclk));
	jxor g04411(.dina(w_n4293_0[0]),.dinb(w_n2833_49[2]),.dout(n4633),.clk(gclk));
	jand g04412(.dina(n4633),.dinb(w_asqrt38_37[1]),.dout(n4634),.clk(gclk));
	jxor g04413(.dina(n4634),.dinb(w_n4298_0[0]),.dout(n4635),.clk(gclk));
	jand g04414(.dina(w_n4635_0[1]),.dinb(n4632),.dout(n4636),.clk(gclk));
	jor g04415(.dina(n4636),.dinb(w_n4631_0[1]),.dout(n4637),.clk(gclk));
	jand g04416(.dina(w_n4637_0[2]),.dinb(w_asqrt46_32[0]),.dout(n4638),.clk(gclk));
	jor g04417(.dina(w_n4637_0[1]),.dinb(w_asqrt46_31[2]),.dout(n4639),.clk(gclk));
	jxor g04418(.dina(w_n4301_0[0]),.dinb(w_n2572_52[1]),.dout(n4640),.clk(gclk));
	jand g04419(.dina(n4640),.dinb(w_asqrt38_37[0]),.dout(n4641),.clk(gclk));
	jxor g04420(.dina(n4641),.dinb(w_n4306_0[0]),.dout(n4642),.clk(gclk));
	jnot g04421(.din(w_n4642_0[1]),.dout(n4643),.clk(gclk));
	jand g04422(.dina(w_n4643_0[1]),.dinb(n4639),.dout(n4644),.clk(gclk));
	jor g04423(.dina(n4644),.dinb(w_n4638_0[1]),.dout(n4645),.clk(gclk));
	jand g04424(.dina(w_n4645_0[2]),.dinb(w_asqrt47_30[1]),.dout(n4646),.clk(gclk));
	jor g04425(.dina(w_n4645_0[1]),.dinb(w_asqrt47_30[0]),.dout(n4647),.clk(gclk));
	jxor g04426(.dina(w_n4308_0[0]),.dinb(w_n2345_50[1]),.dout(n4648),.clk(gclk));
	jand g04427(.dina(n4648),.dinb(w_asqrt38_36[2]),.dout(n4649),.clk(gclk));
	jxor g04428(.dina(n4649),.dinb(w_n4313_0[0]),.dout(n4650),.clk(gclk));
	jand g04429(.dina(w_n4650_0[1]),.dinb(n4647),.dout(n4651),.clk(gclk));
	jor g04430(.dina(n4651),.dinb(w_n4646_0[1]),.dout(n4652),.clk(gclk));
	jand g04431(.dina(w_n4652_0[2]),.dinb(w_asqrt48_32[1]),.dout(n4653),.clk(gclk));
	jor g04432(.dina(w_n4652_0[1]),.dinb(w_asqrt48_32[0]),.dout(n4654),.clk(gclk));
	jxor g04433(.dina(w_n4316_0[0]),.dinb(w_n2108_53[0]),.dout(n4655),.clk(gclk));
	jand g04434(.dina(n4655),.dinb(w_asqrt38_36[1]),.dout(n4656),.clk(gclk));
	jxor g04435(.dina(n4656),.dinb(w_n4321_0[0]),.dout(n4657),.clk(gclk));
	jnot g04436(.din(w_n4657_0[1]),.dout(n4658),.clk(gclk));
	jand g04437(.dina(w_n4658_0[1]),.dinb(n4654),.dout(n4659),.clk(gclk));
	jor g04438(.dina(n4659),.dinb(w_n4653_0[1]),.dout(n4660),.clk(gclk));
	jand g04439(.dina(w_n4660_0[2]),.dinb(w_asqrt49_30[2]),.dout(n4661),.clk(gclk));
	jor g04440(.dina(w_n4660_0[1]),.dinb(w_asqrt49_30[1]),.dout(n4662),.clk(gclk));
	jxor g04441(.dina(w_n4323_0[0]),.dinb(w_n1912_51[1]),.dout(n4663),.clk(gclk));
	jand g04442(.dina(n4663),.dinb(w_asqrt38_36[0]),.dout(n4664),.clk(gclk));
	jxor g04443(.dina(n4664),.dinb(w_n4328_0[0]),.dout(n4665),.clk(gclk));
	jand g04444(.dina(w_n4665_0[1]),.dinb(n4662),.dout(n4666),.clk(gclk));
	jor g04445(.dina(n4666),.dinb(w_n4661_0[1]),.dout(n4667),.clk(gclk));
	jand g04446(.dina(w_n4667_0[2]),.dinb(w_asqrt50_32[2]),.dout(n4668),.clk(gclk));
	jor g04447(.dina(w_n4667_0[1]),.dinb(w_asqrt50_32[1]),.dout(n4669),.clk(gclk));
	jxor g04448(.dina(w_n4331_0[0]),.dinb(w_n1699_53[2]),.dout(n4670),.clk(gclk));
	jand g04449(.dina(n4670),.dinb(w_asqrt38_35[2]),.dout(n4671),.clk(gclk));
	jxor g04450(.dina(n4671),.dinb(w_n4336_0[0]),.dout(n4672),.clk(gclk));
	jand g04451(.dina(w_n4672_0[1]),.dinb(n4669),.dout(n4673),.clk(gclk));
	jor g04452(.dina(n4673),.dinb(w_n4668_0[1]),.dout(n4674),.clk(gclk));
	jand g04453(.dina(w_n4674_0[2]),.dinb(w_asqrt51_31[0]),.dout(n4675),.clk(gclk));
	jor g04454(.dina(w_n4674_0[1]),.dinb(w_asqrt51_30[2]),.dout(n4676),.clk(gclk));
	jxor g04455(.dina(w_n4339_0[0]),.dinb(w_n1516_52[0]),.dout(n4677),.clk(gclk));
	jand g04456(.dina(n4677),.dinb(w_asqrt38_35[1]),.dout(n4678),.clk(gclk));
	jxor g04457(.dina(n4678),.dinb(w_n4344_0[0]),.dout(n4679),.clk(gclk));
	jnot g04458(.din(w_n4679_0[1]),.dout(n4680),.clk(gclk));
	jand g04459(.dina(w_n4680_0[1]),.dinb(n4676),.dout(n4681),.clk(gclk));
	jor g04460(.dina(n4681),.dinb(w_n4675_0[1]),.dout(n4682),.clk(gclk));
	jand g04461(.dina(w_n4682_0[2]),.dinb(w_asqrt52_32[2]),.dout(n4683),.clk(gclk));
	jor g04462(.dina(w_n4682_0[1]),.dinb(w_asqrt52_32[1]),.dout(n4684),.clk(gclk));
	jxor g04463(.dina(w_n4346_0[0]),.dinb(w_n1332_53[2]),.dout(n4685),.clk(gclk));
	jand g04464(.dina(n4685),.dinb(w_asqrt38_35[0]),.dout(n4686),.clk(gclk));
	jxor g04465(.dina(n4686),.dinb(w_n4351_0[0]),.dout(n4687),.clk(gclk));
	jnot g04466(.din(w_n4687_0[1]),.dout(n4688),.clk(gclk));
	jand g04467(.dina(w_n4688_0[1]),.dinb(n4684),.dout(n4689),.clk(gclk));
	jor g04468(.dina(n4689),.dinb(w_n4683_0[1]),.dout(n4690),.clk(gclk));
	jand g04469(.dina(w_n4690_0[2]),.dinb(w_asqrt53_31[2]),.dout(n4691),.clk(gclk));
	jor g04470(.dina(w_n4690_0[1]),.dinb(w_asqrt53_31[1]),.dout(n4692),.clk(gclk));
	jxor g04471(.dina(w_n4353_0[0]),.dinb(w_n1173_52[2]),.dout(n4693),.clk(gclk));
	jand g04472(.dina(n4693),.dinb(w_asqrt38_34[2]),.dout(n4694),.clk(gclk));
	jxor g04473(.dina(n4694),.dinb(w_n4358_0[0]),.dout(n4695),.clk(gclk));
	jand g04474(.dina(w_n4695_0[1]),.dinb(n4692),.dout(n4696),.clk(gclk));
	jor g04475(.dina(n4696),.dinb(w_n4691_0[1]),.dout(n4697),.clk(gclk));
	jand g04476(.dina(w_n4697_0[2]),.dinb(w_asqrt54_32[2]),.dout(n4698),.clk(gclk));
	jor g04477(.dina(w_n4697_0[1]),.dinb(w_asqrt54_32[1]),.dout(n4699),.clk(gclk));
	jxor g04478(.dina(w_n4361_0[0]),.dinb(w_n1008_54[2]),.dout(n4700),.clk(gclk));
	jand g04479(.dina(n4700),.dinb(w_asqrt38_34[1]),.dout(n4701),.clk(gclk));
	jxor g04480(.dina(n4701),.dinb(w_n4366_0[0]),.dout(n4702),.clk(gclk));
	jnot g04481(.din(w_n4702_0[1]),.dout(n4703),.clk(gclk));
	jand g04482(.dina(w_n4703_0[1]),.dinb(n4699),.dout(n4704),.clk(gclk));
	jor g04483(.dina(n4704),.dinb(w_n4698_0[1]),.dout(n4705),.clk(gclk));
	jand g04484(.dina(w_n4705_0[2]),.dinb(w_asqrt55_32[0]),.dout(n4706),.clk(gclk));
	jor g04485(.dina(w_n4705_0[1]),.dinb(w_asqrt55_31[2]),.dout(n4707),.clk(gclk));
	jxor g04486(.dina(w_n4368_0[0]),.dinb(w_n884_53[2]),.dout(n4708),.clk(gclk));
	jand g04487(.dina(n4708),.dinb(w_asqrt38_34[0]),.dout(n4709),.clk(gclk));
	jxor g04488(.dina(n4709),.dinb(w_n4373_0[0]),.dout(n4710),.clk(gclk));
	jand g04489(.dina(w_n4710_0[1]),.dinb(n4707),.dout(n4711),.clk(gclk));
	jor g04490(.dina(n4711),.dinb(w_n4706_0[1]),.dout(n4712),.clk(gclk));
	jand g04491(.dina(w_n4712_0[2]),.dinb(w_asqrt56_33[0]),.dout(n4713),.clk(gclk));
	jor g04492(.dina(w_n4712_0[1]),.dinb(w_asqrt56_32[2]),.dout(n4714),.clk(gclk));
	jxor g04493(.dina(w_n4376_0[0]),.dinb(w_n743_54[2]),.dout(n4715),.clk(gclk));
	jand g04494(.dina(n4715),.dinb(w_asqrt38_33[2]),.dout(n4716),.clk(gclk));
	jxor g04495(.dina(n4716),.dinb(w_n4381_0[0]),.dout(n4717),.clk(gclk));
	jnot g04496(.din(w_n4717_0[1]),.dout(n4718),.clk(gclk));
	jand g04497(.dina(w_n4718_0[1]),.dinb(n4714),.dout(n4719),.clk(gclk));
	jor g04498(.dina(n4719),.dinb(w_n4713_0[1]),.dout(n4720),.clk(gclk));
	jand g04499(.dina(w_n4720_0[2]),.dinb(w_asqrt57_32[2]),.dout(n4721),.clk(gclk));
	jor g04500(.dina(w_n4720_0[1]),.dinb(w_asqrt57_32[1]),.dout(n4722),.clk(gclk));
	jxor g04501(.dina(w_n4383_0[0]),.dinb(w_n635_54[2]),.dout(n4723),.clk(gclk));
	jand g04502(.dina(n4723),.dinb(w_asqrt38_33[1]),.dout(n4724),.clk(gclk));
	jxor g04503(.dina(n4724),.dinb(w_n4388_0[0]),.dout(n4725),.clk(gclk));
	jand g04504(.dina(w_n4725_0[1]),.dinb(n4722),.dout(n4726),.clk(gclk));
	jor g04505(.dina(n4726),.dinb(w_n4721_0[1]),.dout(n4727),.clk(gclk));
	jand g04506(.dina(w_n4727_0[2]),.dinb(w_asqrt58_33[1]),.dout(n4728),.clk(gclk));
	jor g04507(.dina(w_n4727_0[1]),.dinb(w_asqrt58_33[0]),.dout(n4729),.clk(gclk));
	jxor g04508(.dina(w_n4391_0[0]),.dinb(w_n515_55[2]),.dout(n4730),.clk(gclk));
	jand g04509(.dina(n4730),.dinb(w_asqrt38_33[0]),.dout(n4731),.clk(gclk));
	jxor g04510(.dina(n4731),.dinb(w_n4396_0[0]),.dout(n4732),.clk(gclk));
	jnot g04511(.din(w_n4732_0[1]),.dout(n4733),.clk(gclk));
	jand g04512(.dina(w_n4733_0[1]),.dinb(n4729),.dout(n4734),.clk(gclk));
	jor g04513(.dina(n4734),.dinb(w_n4728_0[1]),.dout(n4735),.clk(gclk));
	jand g04514(.dina(w_n4735_0[2]),.dinb(w_asqrt59_33[0]),.dout(n4736),.clk(gclk));
	jor g04515(.dina(w_n4735_0[1]),.dinb(w_asqrt59_32[2]),.dout(n4737),.clk(gclk));
	jxor g04516(.dina(w_n4398_0[0]),.dinb(w_n443_55[2]),.dout(n4738),.clk(gclk));
	jand g04517(.dina(n4738),.dinb(w_asqrt38_32[2]),.dout(n4739),.clk(gclk));
	jxor g04518(.dina(n4739),.dinb(w_n4403_0[0]),.dout(n4740),.clk(gclk));
	jand g04519(.dina(w_n4740_0[1]),.dinb(n4737),.dout(n4741),.clk(gclk));
	jor g04520(.dina(n4741),.dinb(w_n4736_0[1]),.dout(n4742),.clk(gclk));
	jand g04521(.dina(w_n4742_0[2]),.dinb(w_asqrt60_33[1]),.dout(n4743),.clk(gclk));
	jor g04522(.dina(w_n4742_0[1]),.dinb(w_asqrt60_33[0]),.dout(n4744),.clk(gclk));
	jxor g04523(.dina(w_n4406_0[0]),.dinb(w_n352_56[0]),.dout(n4745),.clk(gclk));
	jand g04524(.dina(n4745),.dinb(w_asqrt38_32[1]),.dout(n4746),.clk(gclk));
	jxor g04525(.dina(n4746),.dinb(w_n4411_0[0]),.dout(n4747),.clk(gclk));
	jnot g04526(.din(w_n4747_0[1]),.dout(n4748),.clk(gclk));
	jand g04527(.dina(w_n4748_0[1]),.dinb(n4744),.dout(n4749),.clk(gclk));
	jor g04528(.dina(n4749),.dinb(w_n4743_0[1]),.dout(n4750),.clk(gclk));
	jand g04529(.dina(w_n4750_0[2]),.dinb(w_asqrt61_33[1]),.dout(n4751),.clk(gclk));
	jor g04530(.dina(w_n4750_0[1]),.dinb(w_asqrt61_33[0]),.dout(n4752),.clk(gclk));
	jxor g04531(.dina(w_n4413_0[0]),.dinb(w_n294_56[1]),.dout(n4753),.clk(gclk));
	jand g04532(.dina(n4753),.dinb(w_asqrt38_32[0]),.dout(n4754),.clk(gclk));
	jxor g04533(.dina(n4754),.dinb(w_n4418_0[0]),.dout(n4755),.clk(gclk));
	jand g04534(.dina(w_n4755_0[1]),.dinb(n4752),.dout(n4756),.clk(gclk));
	jor g04535(.dina(n4756),.dinb(w_n4751_0[1]),.dout(n4757),.clk(gclk));
	jand g04536(.dina(w_n4757_0[2]),.dinb(w_asqrt62_33[1]),.dout(n4758),.clk(gclk));
	jor g04537(.dina(w_n4757_0[1]),.dinb(w_asqrt62_33[0]),.dout(n4759),.clk(gclk));
	jxor g04538(.dina(w_n4421_0[0]),.dinb(w_n239_56[1]),.dout(n4760),.clk(gclk));
	jand g04539(.dina(n4760),.dinb(w_asqrt38_31[2]),.dout(n4761),.clk(gclk));
	jxor g04540(.dina(n4761),.dinb(w_n4426_0[0]),.dout(n4762),.clk(gclk));
	jnot g04541(.din(w_n4762_0[2]),.dout(n4763),.clk(gclk));
	jand g04542(.dina(n4763),.dinb(n4759),.dout(n4764),.clk(gclk));
	jor g04543(.dina(n4764),.dinb(w_n4758_0[1]),.dout(n4765),.clk(gclk));
	jor g04544(.dina(w_n4765_0[1]),.dinb(w_n4455_0[2]),.dout(n4766),.clk(gclk));
	jnot g04545(.din(w_n4766_1[1]),.dout(n4767),.clk(gclk));
	jand g04546(.dina(w_n4582_48[0]),.dinb(w_n4435_0[0]),.dout(n4768),.clk(gclk));
	jnot g04547(.din(n4768),.dout(n4769),.clk(gclk));
	jand g04548(.dina(w_n4436_0[0]),.dinb(w_asqrt63_42[2]),.dout(n4770),.clk(gclk));
	jand g04549(.dina(n4770),.dinb(w_n4590_0[0]),.dout(n4771),.clk(gclk));
	jand g04550(.dina(w_n4771_0[1]),.dinb(n4769),.dout(n4772),.clk(gclk));
	jnot g04551(.din(w_n4455_0[1]),.dout(n4773),.clk(gclk));
	jnot g04552(.din(w_n4758_0[0]),.dout(n4774),.clk(gclk));
	jnot g04553(.din(w_n4751_0[0]),.dout(n4775),.clk(gclk));
	jnot g04554(.din(w_n4743_0[0]),.dout(n4776),.clk(gclk));
	jnot g04555(.din(w_n4736_0[0]),.dout(n4777),.clk(gclk));
	jnot g04556(.din(w_n4728_0[0]),.dout(n4778),.clk(gclk));
	jnot g04557(.din(w_n4721_0[0]),.dout(n4779),.clk(gclk));
	jnot g04558(.din(w_n4713_0[0]),.dout(n4780),.clk(gclk));
	jnot g04559(.din(w_n4706_0[0]),.dout(n4781),.clk(gclk));
	jnot g04560(.din(w_n4698_0[0]),.dout(n4782),.clk(gclk));
	jnot g04561(.din(w_n4691_0[0]),.dout(n4783),.clk(gclk));
	jnot g04562(.din(w_n4683_0[0]),.dout(n4784),.clk(gclk));
	jnot g04563(.din(w_n4675_0[0]),.dout(n4785),.clk(gclk));
	jnot g04564(.din(w_n4668_0[0]),.dout(n4786),.clk(gclk));
	jnot g04565(.din(w_n4661_0[0]),.dout(n4787),.clk(gclk));
	jnot g04566(.din(w_n4653_0[0]),.dout(n4788),.clk(gclk));
	jnot g04567(.din(w_n4646_0[0]),.dout(n4789),.clk(gclk));
	jnot g04568(.din(w_n4638_0[0]),.dout(n4790),.clk(gclk));
	jnot g04569(.din(w_n4631_0[0]),.dout(n4791),.clk(gclk));
	jnot g04570(.din(w_n4623_0[0]),.dout(n4792),.clk(gclk));
	jnot g04571(.din(w_n4615_0[0]),.dout(n4793),.clk(gclk));
	jnot g04572(.din(w_n4607_0[0]),.dout(n4794),.clk(gclk));
	jnot g04573(.din(w_n4599_0[0]),.dout(n4795),.clk(gclk));
	jnot g04574(.din(w_n4587_0[0]),.dout(n4796),.clk(gclk));
	jnot g04575(.din(w_n4462_0[0]),.dout(n4797),.clk(gclk));
	jor g04576(.dina(w_n4582_47[2]),.dinb(w_n4255_0[2]),.dout(n4798),.clk(gclk));
	jnot g04577(.din(w_n4460_0[0]),.dout(n4799),.clk(gclk));
	jand g04578(.dina(n4799),.dinb(n4798),.dout(n4800),.clk(gclk));
	jand g04579(.dina(n4800),.dinb(w_n4249_50[2]),.dout(n4801),.clk(gclk));
	jor g04580(.dina(w_n4582_47[1]),.dinb(w_a76_0[0]),.dout(n4802),.clk(gclk));
	jand g04581(.dina(n4802),.dinb(w_a77_0[0]),.dout(n4803),.clk(gclk));
	jor g04582(.dina(w_n4589_0[0]),.dinb(n4803),.dout(n4804),.clk(gclk));
	jor g04583(.dina(w_n4804_0[1]),.dinb(n4801),.dout(n4805),.clk(gclk));
	jand g04584(.dina(n4805),.dinb(n4797),.dout(n4806),.clk(gclk));
	jand g04585(.dina(n4806),.dinb(w_n3955_47[2]),.dout(n4807),.clk(gclk));
	jor g04586(.dina(w_n4595_0[1]),.dinb(n4807),.dout(n4808),.clk(gclk));
	jand g04587(.dina(n4808),.dinb(n4796),.dout(n4809),.clk(gclk));
	jand g04588(.dina(n4809),.dinb(w_n3642_51[0]),.dout(n4810),.clk(gclk));
	jor g04589(.dina(w_n4603_0[0]),.dinb(n4810),.dout(n4811),.clk(gclk));
	jand g04590(.dina(n4811),.dinb(n4795),.dout(n4812),.clk(gclk));
	jand g04591(.dina(n4812),.dinb(w_n3368_48[1]),.dout(n4813),.clk(gclk));
	jor g04592(.dina(w_n4611_0[0]),.dinb(n4813),.dout(n4814),.clk(gclk));
	jand g04593(.dina(n4814),.dinb(n4794),.dout(n4815),.clk(gclk));
	jand g04594(.dina(n4815),.dinb(w_n3089_51[2]),.dout(n4816),.clk(gclk));
	jor g04595(.dina(w_n4619_0[0]),.dinb(n4816),.dout(n4817),.clk(gclk));
	jand g04596(.dina(n4817),.dinb(n4793),.dout(n4818),.clk(gclk));
	jand g04597(.dina(n4818),.dinb(w_n2833_49[1]),.dout(n4819),.clk(gclk));
	jor g04598(.dina(w_n4627_0[0]),.dinb(n4819),.dout(n4820),.clk(gclk));
	jand g04599(.dina(n4820),.dinb(n4792),.dout(n4821),.clk(gclk));
	jand g04600(.dina(n4821),.dinb(w_n2572_52[0]),.dout(n4822),.clk(gclk));
	jnot g04601(.din(w_n4635_0[0]),.dout(n4823),.clk(gclk));
	jor g04602(.dina(w_n4823_0[1]),.dinb(n4822),.dout(n4824),.clk(gclk));
	jand g04603(.dina(n4824),.dinb(n4791),.dout(n4825),.clk(gclk));
	jand g04604(.dina(n4825),.dinb(w_n2345_50[0]),.dout(n4826),.clk(gclk));
	jor g04605(.dina(w_n4642_0[0]),.dinb(n4826),.dout(n4827),.clk(gclk));
	jand g04606(.dina(n4827),.dinb(n4790),.dout(n4828),.clk(gclk));
	jand g04607(.dina(n4828),.dinb(w_n2108_52[2]),.dout(n4829),.clk(gclk));
	jnot g04608(.din(w_n4650_0[0]),.dout(n4830),.clk(gclk));
	jor g04609(.dina(w_n4830_0[1]),.dinb(n4829),.dout(n4831),.clk(gclk));
	jand g04610(.dina(n4831),.dinb(n4789),.dout(n4832),.clk(gclk));
	jand g04611(.dina(n4832),.dinb(w_n1912_51[0]),.dout(n4833),.clk(gclk));
	jor g04612(.dina(w_n4657_0[0]),.dinb(n4833),.dout(n4834),.clk(gclk));
	jand g04613(.dina(n4834),.dinb(n4788),.dout(n4835),.clk(gclk));
	jand g04614(.dina(n4835),.dinb(w_n1699_53[1]),.dout(n4836),.clk(gclk));
	jnot g04615(.din(w_n4665_0[0]),.dout(n4837),.clk(gclk));
	jor g04616(.dina(w_n4837_0[1]),.dinb(n4836),.dout(n4838),.clk(gclk));
	jand g04617(.dina(n4838),.dinb(n4787),.dout(n4839),.clk(gclk));
	jand g04618(.dina(n4839),.dinb(w_n1516_51[2]),.dout(n4840),.clk(gclk));
	jnot g04619(.din(w_n4672_0[0]),.dout(n4841),.clk(gclk));
	jor g04620(.dina(w_n4841_0[1]),.dinb(n4840),.dout(n4842),.clk(gclk));
	jand g04621(.dina(n4842),.dinb(n4786),.dout(n4843),.clk(gclk));
	jand g04622(.dina(n4843),.dinb(w_n1332_53[1]),.dout(n4844),.clk(gclk));
	jor g04623(.dina(w_n4679_0[0]),.dinb(n4844),.dout(n4845),.clk(gclk));
	jand g04624(.dina(n4845),.dinb(n4785),.dout(n4846),.clk(gclk));
	jand g04625(.dina(n4846),.dinb(w_n1173_52[1]),.dout(n4847),.clk(gclk));
	jor g04626(.dina(w_n4687_0[0]),.dinb(n4847),.dout(n4848),.clk(gclk));
	jand g04627(.dina(n4848),.dinb(n4784),.dout(n4849),.clk(gclk));
	jand g04628(.dina(n4849),.dinb(w_n1008_54[1]),.dout(n4850),.clk(gclk));
	jnot g04629(.din(w_n4695_0[0]),.dout(n4851),.clk(gclk));
	jor g04630(.dina(w_n4851_0[1]),.dinb(n4850),.dout(n4852),.clk(gclk));
	jand g04631(.dina(n4852),.dinb(n4783),.dout(n4853),.clk(gclk));
	jand g04632(.dina(n4853),.dinb(w_n884_53[1]),.dout(n4854),.clk(gclk));
	jor g04633(.dina(w_n4702_0[0]),.dinb(n4854),.dout(n4855),.clk(gclk));
	jand g04634(.dina(n4855),.dinb(n4782),.dout(n4856),.clk(gclk));
	jand g04635(.dina(n4856),.dinb(w_n743_54[1]),.dout(n4857),.clk(gclk));
	jnot g04636(.din(w_n4710_0[0]),.dout(n4858),.clk(gclk));
	jor g04637(.dina(w_n4858_0[1]),.dinb(n4857),.dout(n4859),.clk(gclk));
	jand g04638(.dina(n4859),.dinb(n4781),.dout(n4860),.clk(gclk));
	jand g04639(.dina(n4860),.dinb(w_n635_54[1]),.dout(n4861),.clk(gclk));
	jor g04640(.dina(w_n4717_0[0]),.dinb(n4861),.dout(n4862),.clk(gclk));
	jand g04641(.dina(n4862),.dinb(n4780),.dout(n4863),.clk(gclk));
	jand g04642(.dina(n4863),.dinb(w_n515_55[1]),.dout(n4864),.clk(gclk));
	jnot g04643(.din(w_n4725_0[0]),.dout(n4865),.clk(gclk));
	jor g04644(.dina(w_n4865_0[1]),.dinb(n4864),.dout(n4866),.clk(gclk));
	jand g04645(.dina(n4866),.dinb(n4779),.dout(n4867),.clk(gclk));
	jand g04646(.dina(n4867),.dinb(w_n443_55[1]),.dout(n4868),.clk(gclk));
	jor g04647(.dina(w_n4732_0[0]),.dinb(n4868),.dout(n4869),.clk(gclk));
	jand g04648(.dina(n4869),.dinb(n4778),.dout(n4870),.clk(gclk));
	jand g04649(.dina(n4870),.dinb(w_n352_55[2]),.dout(n4871),.clk(gclk));
	jnot g04650(.din(w_n4740_0[0]),.dout(n4872),.clk(gclk));
	jor g04651(.dina(w_n4872_0[1]),.dinb(n4871),.dout(n4873),.clk(gclk));
	jand g04652(.dina(n4873),.dinb(n4777),.dout(n4874),.clk(gclk));
	jand g04653(.dina(n4874),.dinb(w_n294_56[0]),.dout(n4875),.clk(gclk));
	jor g04654(.dina(w_n4747_0[0]),.dinb(n4875),.dout(n4876),.clk(gclk));
	jand g04655(.dina(n4876),.dinb(n4776),.dout(n4877),.clk(gclk));
	jand g04656(.dina(n4877),.dinb(w_n239_56[0]),.dout(n4878),.clk(gclk));
	jnot g04657(.din(w_n4755_0[0]),.dout(n4879),.clk(gclk));
	jor g04658(.dina(w_n4879_0[1]),.dinb(n4878),.dout(n4880),.clk(gclk));
	jand g04659(.dina(n4880),.dinb(n4775),.dout(n4881),.clk(gclk));
	jand g04660(.dina(n4881),.dinb(w_n221_56[1]),.dout(n4882),.clk(gclk));
	jor g04661(.dina(w_n4762_0[1]),.dinb(n4882),.dout(n4883),.clk(gclk));
	jand g04662(.dina(n4883),.dinb(n4774),.dout(n4884),.clk(gclk));
	jor g04663(.dina(w_n4884_0[1]),.dinb(n4773),.dout(n4885),.clk(gclk));
	jand g04664(.dina(w_asqrt38_31[1]),.dinb(w_n4576_0[0]),.dout(n4886),.clk(gclk));
	jor g04665(.dina(n4886),.dinb(w_n4442_0[0]),.dout(n4887),.clk(gclk));
	jor g04666(.dina(w_n4887_0[1]),.dinb(w_n4885_0[1]),.dout(n4888),.clk(gclk));
	jand g04667(.dina(n4888),.dinb(w_n218_23[1]),.dout(n4889),.clk(gclk));
	jand g04668(.dina(w_n4582_47[0]),.dinb(w_n4253_0[0]),.dout(n4890),.clk(gclk));
	jor g04669(.dina(w_n4890_0[1]),.dinb(w_n4889_0[1]),.dout(n4891),.clk(gclk));
	jor g04670(.dina(n4891),.dinb(w_n4772_0[1]),.dout(n4892),.clk(gclk));
	jor g04671(.dina(w_n4892_0[1]),.dinb(w_n4767_0[2]),.dout(asqrt_fa_38),.clk(gclk));
	jnot g04672(.din(w_n4772_0[0]),.dout(n4894),.clk(gclk));
	jand g04673(.dina(w_n4765_0[0]),.dinb(w_n4455_0[0]),.dout(n4895),.clk(gclk));
	jnot g04674(.din(w_n4887_0[0]),.dout(n4896),.clk(gclk));
	jand g04675(.dina(n4896),.dinb(w_n4895_0[1]),.dout(n4897),.clk(gclk));
	jor g04676(.dina(n4897),.dinb(w_asqrt63_42[1]),.dout(n4898),.clk(gclk));
	jnot g04677(.din(w_n4890_0[0]),.dout(n4899),.clk(gclk));
	jand g04678(.dina(n4899),.dinb(n4898),.dout(n4900),.clk(gclk));
	jand g04679(.dina(n4900),.dinb(n4894),.dout(n4901),.clk(gclk));
	jand g04680(.dina(w_n4901_0[1]),.dinb(w_n4766_1[0]),.dout(n4902),.clk(gclk));
	jxor g04681(.dina(w_n4757_0[0]),.dinb(w_n221_56[0]),.dout(n4903),.clk(gclk));
	jor g04682(.dina(n4903),.dinb(w_n4902_57[1]),.dout(n4904),.clk(gclk));
	jxor g04683(.dina(n4904),.dinb(w_n4762_0[0]),.dout(n4905),.clk(gclk));
	jnot g04684(.din(w_n4905_0[1]),.dout(n4906),.clk(gclk));
	jor g04685(.dina(w_n4902_57[0]),.dinb(w_n4457_1[0]),.dout(n4907),.clk(gclk));
	jnot g04686(.din(w_a72_0[2]),.dout(n4908),.clk(gclk));
	jnot g04687(.din(w_a73_0[1]),.dout(n4909),.clk(gclk));
	jand g04688(.dina(w_n4909_0[1]),.dinb(w_n4908_1[2]),.dout(n4910),.clk(gclk));
	jand g04689(.dina(w_n4910_0[2]),.dinb(w_n4457_0[2]),.dout(n4911),.clk(gclk));
	jnot g04690(.din(w_n4911_0[1]),.dout(n4912),.clk(gclk));
	jand g04691(.dina(n4912),.dinb(n4907),.dout(n4913),.clk(gclk));
	jor g04692(.dina(w_n4913_0[2]),.dinb(w_n4582_46[2]),.dout(n4914),.clk(gclk));
	jand g04693(.dina(w_n4913_0[1]),.dinb(w_n4582_46[1]),.dout(n4915),.clk(gclk));
	jor g04694(.dina(w_n4902_56[2]),.dinb(w_a74_1[0]),.dout(n4916),.clk(gclk));
	jand g04695(.dina(n4916),.dinb(w_a75_0[0]),.dout(n4917),.clk(gclk));
	jand g04696(.dina(w_asqrt37_28),.dinb(w_n4459_0[1]),.dout(n4918),.clk(gclk));
	jor g04697(.dina(n4918),.dinb(n4917),.dout(n4919),.clk(gclk));
	jor g04698(.dina(n4919),.dinb(n4915),.dout(n4920),.clk(gclk));
	jand g04699(.dina(n4920),.dinb(w_n4914_0[1]),.dout(n4921),.clk(gclk));
	jor g04700(.dina(w_n4921_0[2]),.dinb(w_n4249_50[1]),.dout(n4922),.clk(gclk));
	jand g04701(.dina(w_n4921_0[1]),.dinb(w_n4249_50[0]),.dout(n4923),.clk(gclk));
	jnot g04702(.din(w_n4459_0[0]),.dout(n4924),.clk(gclk));
	jor g04703(.dina(w_n4902_56[1]),.dinb(n4924),.dout(n4925),.clk(gclk));
	jor g04704(.dina(w_n4767_0[1]),.dinb(w_n4582_46[0]),.dout(n4926),.clk(gclk));
	jor g04705(.dina(n4926),.dinb(w_n4771_0[0]),.dout(n4927),.clk(gclk));
	jor g04706(.dina(n4927),.dinb(w_n4889_0[0]),.dout(n4928),.clk(gclk));
	jand g04707(.dina(n4928),.dinb(w_n4925_0[1]),.dout(n4929),.clk(gclk));
	jxor g04708(.dina(n4929),.dinb(w_n4255_0[1]),.dout(n4930),.clk(gclk));
	jor g04709(.dina(w_n4930_0[2]),.dinb(n4923),.dout(n4931),.clk(gclk));
	jand g04710(.dina(n4931),.dinb(w_n4922_0[1]),.dout(n4932),.clk(gclk));
	jor g04711(.dina(w_n4932_0[2]),.dinb(w_n3955_47[1]),.dout(n4933),.clk(gclk));
	jand g04712(.dina(w_n4932_0[1]),.dinb(w_n3955_47[0]),.dout(n4934),.clk(gclk));
	jxor g04713(.dina(w_n4461_0[0]),.dinb(w_n4249_49[2]),.dout(n4935),.clk(gclk));
	jor g04714(.dina(n4935),.dinb(w_n4902_56[0]),.dout(n4936),.clk(gclk));
	jxor g04715(.dina(n4936),.dinb(w_n4804_0[0]),.dout(n4937),.clk(gclk));
	jnot g04716(.din(w_n4937_0[2]),.dout(n4938),.clk(gclk));
	jor g04717(.dina(n4938),.dinb(n4934),.dout(n4939),.clk(gclk));
	jand g04718(.dina(n4939),.dinb(w_n4933_0[1]),.dout(n4940),.clk(gclk));
	jor g04719(.dina(w_n4940_0[2]),.dinb(w_n3642_50[2]),.dout(n4941),.clk(gclk));
	jand g04720(.dina(w_n4940_0[1]),.dinb(w_n3642_50[1]),.dout(n4942),.clk(gclk));
	jxor g04721(.dina(w_n4586_0[0]),.dinb(w_n3955_46[2]),.dout(n4943),.clk(gclk));
	jor g04722(.dina(n4943),.dinb(w_n4902_55[2]),.dout(n4944),.clk(gclk));
	jxor g04723(.dina(n4944),.dinb(w_n4595_0[0]),.dout(n4945),.clk(gclk));
	jnot g04724(.din(w_n4945_0[2]),.dout(n4946),.clk(gclk));
	jor g04725(.dina(n4946),.dinb(n4942),.dout(n4947),.clk(gclk));
	jand g04726(.dina(n4947),.dinb(w_n4941_0[1]),.dout(n4948),.clk(gclk));
	jor g04727(.dina(w_n4948_0[2]),.dinb(w_n3368_48[0]),.dout(n4949),.clk(gclk));
	jand g04728(.dina(w_n4948_0[1]),.dinb(w_n3368_47[2]),.dout(n4950),.clk(gclk));
	jxor g04729(.dina(w_n4598_0[0]),.dinb(w_n3642_50[0]),.dout(n4951),.clk(gclk));
	jor g04730(.dina(n4951),.dinb(w_n4902_55[1]),.dout(n4952),.clk(gclk));
	jxor g04731(.dina(n4952),.dinb(w_n4604_0[0]),.dout(n4953),.clk(gclk));
	jor g04732(.dina(w_n4953_0[1]),.dinb(n4950),.dout(n4954),.clk(gclk));
	jand g04733(.dina(n4954),.dinb(w_n4949_0[1]),.dout(n4955),.clk(gclk));
	jor g04734(.dina(w_n4955_0[2]),.dinb(w_n3089_51[1]),.dout(n4956),.clk(gclk));
	jand g04735(.dina(w_n4955_0[1]),.dinb(w_n3089_51[0]),.dout(n4957),.clk(gclk));
	jxor g04736(.dina(w_n4606_0[0]),.dinb(w_n3368_47[1]),.dout(n4958),.clk(gclk));
	jor g04737(.dina(n4958),.dinb(w_n4902_55[0]),.dout(n4959),.clk(gclk));
	jxor g04738(.dina(n4959),.dinb(w_n4612_0[0]),.dout(n4960),.clk(gclk));
	jor g04739(.dina(w_n4960_0[2]),.dinb(n4957),.dout(n4961),.clk(gclk));
	jand g04740(.dina(n4961),.dinb(w_n4956_0[1]),.dout(n4962),.clk(gclk));
	jor g04741(.dina(w_n4962_0[2]),.dinb(w_n2833_49[0]),.dout(n4963),.clk(gclk));
	jand g04742(.dina(w_n4962_0[1]),.dinb(w_n2833_48[2]),.dout(n4964),.clk(gclk));
	jxor g04743(.dina(w_n4614_0[0]),.dinb(w_n3089_50[2]),.dout(n4965),.clk(gclk));
	jor g04744(.dina(n4965),.dinb(w_n4902_54[2]),.dout(n4966),.clk(gclk));
	jxor g04745(.dina(n4966),.dinb(w_n4620_0[0]),.dout(n4967),.clk(gclk));
	jor g04746(.dina(w_n4967_0[2]),.dinb(n4964),.dout(n4968),.clk(gclk));
	jand g04747(.dina(n4968),.dinb(w_n4963_0[1]),.dout(n4969),.clk(gclk));
	jor g04748(.dina(w_n4969_0[2]),.dinb(w_n2572_51[2]),.dout(n4970),.clk(gclk));
	jand g04749(.dina(w_n4969_0[1]),.dinb(w_n2572_51[1]),.dout(n4971),.clk(gclk));
	jxor g04750(.dina(w_n4622_0[0]),.dinb(w_n2833_48[1]),.dout(n4972),.clk(gclk));
	jor g04751(.dina(n4972),.dinb(w_n4902_54[1]),.dout(n4973),.clk(gclk));
	jxor g04752(.dina(n4973),.dinb(w_n4628_0[0]),.dout(n4974),.clk(gclk));
	jor g04753(.dina(w_n4974_0[2]),.dinb(n4971),.dout(n4975),.clk(gclk));
	jand g04754(.dina(n4975),.dinb(w_n4970_0[1]),.dout(n4976),.clk(gclk));
	jor g04755(.dina(w_n4976_0[2]),.dinb(w_n2345_49[2]),.dout(n4977),.clk(gclk));
	jand g04756(.dina(w_n4976_0[1]),.dinb(w_n2345_49[1]),.dout(n4978),.clk(gclk));
	jxor g04757(.dina(w_n4630_0[0]),.dinb(w_n2572_51[0]),.dout(n4979),.clk(gclk));
	jor g04758(.dina(n4979),.dinb(w_n4902_54[0]),.dout(n4980),.clk(gclk));
	jxor g04759(.dina(n4980),.dinb(w_n4823_0[0]),.dout(n4981),.clk(gclk));
	jnot g04760(.din(w_n4981_0[2]),.dout(n4982),.clk(gclk));
	jor g04761(.dina(n4982),.dinb(n4978),.dout(n4983),.clk(gclk));
	jand g04762(.dina(n4983),.dinb(w_n4977_0[1]),.dout(n4984),.clk(gclk));
	jor g04763(.dina(w_n4984_0[2]),.dinb(w_n2108_52[1]),.dout(n4985),.clk(gclk));
	jand g04764(.dina(w_n4984_0[1]),.dinb(w_n2108_52[0]),.dout(n4986),.clk(gclk));
	jxor g04765(.dina(w_n4637_0[0]),.dinb(w_n2345_49[0]),.dout(n4987),.clk(gclk));
	jor g04766(.dina(n4987),.dinb(w_n4902_53[2]),.dout(n4988),.clk(gclk));
	jxor g04767(.dina(n4988),.dinb(w_n4643_0[0]),.dout(n4989),.clk(gclk));
	jor g04768(.dina(w_n4989_0[2]),.dinb(n4986),.dout(n4990),.clk(gclk));
	jand g04769(.dina(n4990),.dinb(w_n4985_0[1]),.dout(n4991),.clk(gclk));
	jor g04770(.dina(w_n4991_0[2]),.dinb(w_n1912_50[2]),.dout(n4992),.clk(gclk));
	jand g04771(.dina(w_n4991_0[1]),.dinb(w_n1912_50[1]),.dout(n4993),.clk(gclk));
	jxor g04772(.dina(w_n4645_0[0]),.dinb(w_n2108_51[2]),.dout(n4994),.clk(gclk));
	jor g04773(.dina(n4994),.dinb(w_n4902_53[1]),.dout(n4995),.clk(gclk));
	jxor g04774(.dina(n4995),.dinb(w_n4830_0[0]),.dout(n4996),.clk(gclk));
	jnot g04775(.din(w_n4996_0[2]),.dout(n4997),.clk(gclk));
	jor g04776(.dina(n4997),.dinb(n4993),.dout(n4998),.clk(gclk));
	jand g04777(.dina(n4998),.dinb(w_n4992_0[1]),.dout(n4999),.clk(gclk));
	jor g04778(.dina(w_n4999_0[2]),.dinb(w_n1699_53[0]),.dout(n5000),.clk(gclk));
	jand g04779(.dina(w_n4999_0[1]),.dinb(w_n1699_52[2]),.dout(n5001),.clk(gclk));
	jxor g04780(.dina(w_n4652_0[0]),.dinb(w_n1912_50[0]),.dout(n5002),.clk(gclk));
	jor g04781(.dina(n5002),.dinb(w_n4902_53[0]),.dout(n5003),.clk(gclk));
	jxor g04782(.dina(n5003),.dinb(w_n4658_0[0]),.dout(n5004),.clk(gclk));
	jor g04783(.dina(w_n5004_0[2]),.dinb(n5001),.dout(n5005),.clk(gclk));
	jand g04784(.dina(n5005),.dinb(w_n5000_0[1]),.dout(n5006),.clk(gclk));
	jor g04785(.dina(w_n5006_0[2]),.dinb(w_n1516_51[1]),.dout(n5007),.clk(gclk));
	jand g04786(.dina(w_n5006_0[1]),.dinb(w_n1516_51[0]),.dout(n5008),.clk(gclk));
	jxor g04787(.dina(w_n4660_0[0]),.dinb(w_n1699_52[1]),.dout(n5009),.clk(gclk));
	jor g04788(.dina(n5009),.dinb(w_n4902_52[2]),.dout(n5010),.clk(gclk));
	jxor g04789(.dina(n5010),.dinb(w_n4837_0[0]),.dout(n5011),.clk(gclk));
	jnot g04790(.din(w_n5011_0[2]),.dout(n5012),.clk(gclk));
	jor g04791(.dina(n5012),.dinb(n5008),.dout(n5013),.clk(gclk));
	jand g04792(.dina(n5013),.dinb(w_n5007_0[1]),.dout(n5014),.clk(gclk));
	jor g04793(.dina(w_n5014_0[2]),.dinb(w_n1332_53[0]),.dout(n5015),.clk(gclk));
	jand g04794(.dina(w_n5014_0[1]),.dinb(w_n1332_52[2]),.dout(n5016),.clk(gclk));
	jxor g04795(.dina(w_n4667_0[0]),.dinb(w_n1516_50[2]),.dout(n5017),.clk(gclk));
	jor g04796(.dina(n5017),.dinb(w_n4902_52[1]),.dout(n5018),.clk(gclk));
	jxor g04797(.dina(n5018),.dinb(w_n4841_0[0]),.dout(n5019),.clk(gclk));
	jnot g04798(.din(w_n5019_0[2]),.dout(n5020),.clk(gclk));
	jor g04799(.dina(n5020),.dinb(n5016),.dout(n5021),.clk(gclk));
	jand g04800(.dina(n5021),.dinb(w_n5015_0[1]),.dout(n5022),.clk(gclk));
	jor g04801(.dina(w_n5022_0[2]),.dinb(w_n1173_52[0]),.dout(n5023),.clk(gclk));
	jand g04802(.dina(w_n5022_0[1]),.dinb(w_n1173_51[2]),.dout(n5024),.clk(gclk));
	jxor g04803(.dina(w_n4674_0[0]),.dinb(w_n1332_52[1]),.dout(n5025),.clk(gclk));
	jor g04804(.dina(n5025),.dinb(w_n4902_52[0]),.dout(n5026),.clk(gclk));
	jxor g04805(.dina(n5026),.dinb(w_n4680_0[0]),.dout(n5027),.clk(gclk));
	jor g04806(.dina(w_n5027_0[2]),.dinb(n5024),.dout(n5028),.clk(gclk));
	jand g04807(.dina(n5028),.dinb(w_n5023_0[1]),.dout(n5029),.clk(gclk));
	jor g04808(.dina(w_n5029_0[2]),.dinb(w_n1008_54[0]),.dout(n5030),.clk(gclk));
	jand g04809(.dina(w_n5029_0[1]),.dinb(w_n1008_53[2]),.dout(n5031),.clk(gclk));
	jxor g04810(.dina(w_n4682_0[0]),.dinb(w_n1173_51[1]),.dout(n5032),.clk(gclk));
	jor g04811(.dina(n5032),.dinb(w_n4902_51[2]),.dout(n5033),.clk(gclk));
	jxor g04812(.dina(n5033),.dinb(w_n4688_0[0]),.dout(n5034),.clk(gclk));
	jor g04813(.dina(w_n5034_0[2]),.dinb(n5031),.dout(n5035),.clk(gclk));
	jand g04814(.dina(n5035),.dinb(w_n5030_0[1]),.dout(n5036),.clk(gclk));
	jor g04815(.dina(w_n5036_0[2]),.dinb(w_n884_53[0]),.dout(n5037),.clk(gclk));
	jand g04816(.dina(w_n5036_0[1]),.dinb(w_n884_52[2]),.dout(n5038),.clk(gclk));
	jxor g04817(.dina(w_n4690_0[0]),.dinb(w_n1008_53[1]),.dout(n5039),.clk(gclk));
	jor g04818(.dina(n5039),.dinb(w_n4902_51[1]),.dout(n5040),.clk(gclk));
	jxor g04819(.dina(n5040),.dinb(w_n4851_0[0]),.dout(n5041),.clk(gclk));
	jnot g04820(.din(w_n5041_0[2]),.dout(n5042),.clk(gclk));
	jor g04821(.dina(n5042),.dinb(n5038),.dout(n5043),.clk(gclk));
	jand g04822(.dina(n5043),.dinb(w_n5037_0[1]),.dout(n5044),.clk(gclk));
	jor g04823(.dina(w_n5044_0[2]),.dinb(w_n743_54[0]),.dout(n5045),.clk(gclk));
	jand g04824(.dina(w_n5044_0[1]),.dinb(w_n743_53[2]),.dout(n5046),.clk(gclk));
	jxor g04825(.dina(w_n4697_0[0]),.dinb(w_n884_52[1]),.dout(n5047),.clk(gclk));
	jor g04826(.dina(n5047),.dinb(w_n4902_51[0]),.dout(n5048),.clk(gclk));
	jxor g04827(.dina(n5048),.dinb(w_n4703_0[0]),.dout(n5049),.clk(gclk));
	jor g04828(.dina(w_n5049_0[2]),.dinb(n5046),.dout(n5050),.clk(gclk));
	jand g04829(.dina(n5050),.dinb(w_n5045_0[1]),.dout(n5051),.clk(gclk));
	jor g04830(.dina(w_n5051_0[2]),.dinb(w_n635_54[0]),.dout(n5052),.clk(gclk));
	jand g04831(.dina(w_n5051_0[1]),.dinb(w_n635_53[2]),.dout(n5053),.clk(gclk));
	jxor g04832(.dina(w_n4705_0[0]),.dinb(w_n743_53[1]),.dout(n5054),.clk(gclk));
	jor g04833(.dina(n5054),.dinb(w_n4902_50[2]),.dout(n5055),.clk(gclk));
	jxor g04834(.dina(n5055),.dinb(w_n4858_0[0]),.dout(n5056),.clk(gclk));
	jnot g04835(.din(w_n5056_0[2]),.dout(n5057),.clk(gclk));
	jor g04836(.dina(n5057),.dinb(n5053),.dout(n5058),.clk(gclk));
	jand g04837(.dina(n5058),.dinb(w_n5052_0[1]),.dout(n5059),.clk(gclk));
	jor g04838(.dina(w_n5059_0[2]),.dinb(w_n515_55[0]),.dout(n5060),.clk(gclk));
	jand g04839(.dina(w_n5059_0[1]),.dinb(w_n515_54[2]),.dout(n5061),.clk(gclk));
	jxor g04840(.dina(w_n4712_0[0]),.dinb(w_n635_53[1]),.dout(n5062),.clk(gclk));
	jor g04841(.dina(n5062),.dinb(w_n4902_50[1]),.dout(n5063),.clk(gclk));
	jxor g04842(.dina(n5063),.dinb(w_n4718_0[0]),.dout(n5064),.clk(gclk));
	jor g04843(.dina(w_n5064_0[2]),.dinb(n5061),.dout(n5065),.clk(gclk));
	jand g04844(.dina(n5065),.dinb(w_n5060_0[1]),.dout(n5066),.clk(gclk));
	jor g04845(.dina(w_n5066_0[2]),.dinb(w_n443_55[0]),.dout(n5067),.clk(gclk));
	jand g04846(.dina(w_n5066_0[1]),.dinb(w_n443_54[2]),.dout(n5068),.clk(gclk));
	jxor g04847(.dina(w_n4720_0[0]),.dinb(w_n515_54[1]),.dout(n5069),.clk(gclk));
	jor g04848(.dina(n5069),.dinb(w_n4902_50[0]),.dout(n5070),.clk(gclk));
	jxor g04849(.dina(n5070),.dinb(w_n4865_0[0]),.dout(n5071),.clk(gclk));
	jnot g04850(.din(w_n5071_0[1]),.dout(n5072),.clk(gclk));
	jor g04851(.dina(w_n5072_0[1]),.dinb(n5068),.dout(n5073),.clk(gclk));
	jand g04852(.dina(n5073),.dinb(w_n5067_0[1]),.dout(n5074),.clk(gclk));
	jor g04853(.dina(w_n5074_0[2]),.dinb(w_n352_55[1]),.dout(n5075),.clk(gclk));
	jand g04854(.dina(w_n5074_0[1]),.dinb(w_n352_55[0]),.dout(n5076),.clk(gclk));
	jxor g04855(.dina(w_n4727_0[0]),.dinb(w_n443_54[1]),.dout(n5077),.clk(gclk));
	jor g04856(.dina(n5077),.dinb(w_n4902_49[2]),.dout(n5078),.clk(gclk));
	jxor g04857(.dina(n5078),.dinb(w_n4733_0[0]),.dout(n5079),.clk(gclk));
	jor g04858(.dina(w_n5079_0[2]),.dinb(n5076),.dout(n5080),.clk(gclk));
	jand g04859(.dina(n5080),.dinb(w_n5075_0[1]),.dout(n5081),.clk(gclk));
	jor g04860(.dina(w_n5081_0[2]),.dinb(w_n294_55[2]),.dout(n5082),.clk(gclk));
	jand g04861(.dina(w_n5081_0[1]),.dinb(w_n294_55[1]),.dout(n5083),.clk(gclk));
	jxor g04862(.dina(w_n4735_0[0]),.dinb(w_n352_54[2]),.dout(n5084),.clk(gclk));
	jor g04863(.dina(n5084),.dinb(w_n4902_49[1]),.dout(n5085),.clk(gclk));
	jxor g04864(.dina(n5085),.dinb(w_n4872_0[0]),.dout(n5086),.clk(gclk));
	jnot g04865(.din(w_n5086_0[2]),.dout(n5087),.clk(gclk));
	jor g04866(.dina(n5087),.dinb(n5083),.dout(n5088),.clk(gclk));
	jand g04867(.dina(n5088),.dinb(w_n5082_0[1]),.dout(n5089),.clk(gclk));
	jor g04868(.dina(w_n5089_0[2]),.dinb(w_n239_55[2]),.dout(n5090),.clk(gclk));
	jand g04869(.dina(w_n5089_0[1]),.dinb(w_n239_55[1]),.dout(n5091),.clk(gclk));
	jxor g04870(.dina(w_n4742_0[0]),.dinb(w_n294_55[0]),.dout(n5092),.clk(gclk));
	jor g04871(.dina(n5092),.dinb(w_n4902_49[0]),.dout(n5093),.clk(gclk));
	jxor g04872(.dina(n5093),.dinb(w_n4748_0[0]),.dout(n5094),.clk(gclk));
	jor g04873(.dina(w_n5094_0[2]),.dinb(n5091),.dout(n5095),.clk(gclk));
	jand g04874(.dina(n5095),.dinb(w_n5090_0[1]),.dout(n5096),.clk(gclk));
	jor g04875(.dina(w_n5096_0[2]),.dinb(w_n221_55[2]),.dout(n5097),.clk(gclk));
	jand g04876(.dina(w_n5096_0[1]),.dinb(w_n221_55[1]),.dout(n5098),.clk(gclk));
	jxor g04877(.dina(w_n4750_0[0]),.dinb(w_n239_55[0]),.dout(n5099),.clk(gclk));
	jor g04878(.dina(n5099),.dinb(w_n4902_48[2]),.dout(n5100),.clk(gclk));
	jxor g04879(.dina(n5100),.dinb(w_n4879_0[0]),.dout(n5101),.clk(gclk));
	jnot g04880(.din(w_n5101_0[1]),.dout(n5102),.clk(gclk));
	jor g04881(.dina(w_n5102_0[1]),.dinb(n5098),.dout(n5103),.clk(gclk));
	jand g04882(.dina(n5103),.dinb(w_n5097_0[1]),.dout(n5104),.clk(gclk));
	jand g04883(.dina(w_n5104_0[2]),.dinb(w_n4906_0[2]),.dout(n5105),.clk(gclk));
	jand g04884(.dina(w_n4892_0[0]),.dinb(w_n4895_0[0]),.dout(n5107),.clk(gclk));
	jor g04885(.dina(w_n5104_0[1]),.dinb(w_n4906_0[1]),.dout(n5108),.clk(gclk));
	jor g04886(.dina(w_n5108_0[1]),.dinb(w_n4767_0[0]),.dout(n5109),.clk(gclk));
	jor g04887(.dina(n5109),.dinb(w_n5107_0[1]),.dout(n5110),.clk(gclk));
	jand g04888(.dina(n5110),.dinb(w_n218_23[0]),.dout(n5111),.clk(gclk));
	jand g04889(.dina(w_n4901_0[0]),.dinb(w_n4884_0[0]),.dout(n5112),.clk(gclk));
	jand g04890(.dina(w_n4885_0[0]),.dinb(w_asqrt63_42[0]),.dout(n5113),.clk(gclk));
	jand g04891(.dina(n5113),.dinb(w_n4766_0[2]),.dout(n5114),.clk(gclk));
	jnot g04892(.din(n5114),.dout(n5115),.clk(gclk));
	jor g04893(.dina(w_n5115_0[1]),.dinb(n5112),.dout(n5116),.clk(gclk));
	jnot g04894(.din(w_n5116_0[1]),.dout(n5117),.clk(gclk));
	jor g04895(.dina(n5117),.dinb(n5111),.dout(n5118),.clk(gclk));
	jor g04896(.dina(w_n5118_0[1]),.dinb(w_n5105_0[2]),.dout(asqrt_fa_37),.clk(gclk));
	jnot g04897(.din(w_a70_1[1]),.dout(n5121),.clk(gclk));
	jnot g04898(.din(w_a71_0[1]),.dout(n5122),.clk(gclk));
	jand g04899(.dina(w_n5122_0[1]),.dinb(w_n5121_1[1]),.dout(n5123),.clk(gclk));
	jand g04900(.dina(w_n5123_0[2]),.dinb(w_n4908_1[1]),.dout(n5124),.clk(gclk));
	jand g04901(.dina(w_asqrt36_39),.dinb(w_a72_0[1]),.dout(n5125),.clk(gclk));
	jor g04902(.dina(n5125),.dinb(w_n5124_0[1]),.dout(n5126),.clk(gclk));
	jand g04903(.dina(w_n5126_0[2]),.dinb(w_asqrt37_27[2]),.dout(n5127),.clk(gclk));
	jor g04904(.dina(w_n5126_0[1]),.dinb(w_asqrt37_27[1]),.dout(n5128),.clk(gclk));
	jand g04905(.dina(w_asqrt36_38[2]),.dinb(w_n4908_1[0]),.dout(n5129),.clk(gclk));
	jor g04906(.dina(n5129),.dinb(w_n4909_0[0]),.dout(n5130),.clk(gclk));
	jnot g04907(.din(w_n4910_0[1]),.dout(n5131),.clk(gclk));
	jnot g04908(.din(w_n5105_0[1]),.dout(n5132),.clk(gclk));
	jnot g04909(.din(w_n5107_0[0]),.dout(n5134),.clk(gclk));
	jnot g04910(.din(w_n5097_0[0]),.dout(n5135),.clk(gclk));
	jnot g04911(.din(w_n5090_0[0]),.dout(n5136),.clk(gclk));
	jnot g04912(.din(w_n5082_0[0]),.dout(n5137),.clk(gclk));
	jnot g04913(.din(w_n5075_0[0]),.dout(n5138),.clk(gclk));
	jnot g04914(.din(w_n5067_0[0]),.dout(n5139),.clk(gclk));
	jnot g04915(.din(w_n5060_0[0]),.dout(n5140),.clk(gclk));
	jnot g04916(.din(w_n5052_0[0]),.dout(n5141),.clk(gclk));
	jnot g04917(.din(w_n5045_0[0]),.dout(n5142),.clk(gclk));
	jnot g04918(.din(w_n5037_0[0]),.dout(n5143),.clk(gclk));
	jnot g04919(.din(w_n5030_0[0]),.dout(n5144),.clk(gclk));
	jnot g04920(.din(w_n5023_0[0]),.dout(n5145),.clk(gclk));
	jnot g04921(.din(w_n5015_0[0]),.dout(n5146),.clk(gclk));
	jnot g04922(.din(w_n5007_0[0]),.dout(n5147),.clk(gclk));
	jnot g04923(.din(w_n5000_0[0]),.dout(n5148),.clk(gclk));
	jnot g04924(.din(w_n4992_0[0]),.dout(n5149),.clk(gclk));
	jnot g04925(.din(w_n4985_0[0]),.dout(n5150),.clk(gclk));
	jnot g04926(.din(w_n4977_0[0]),.dout(n5151),.clk(gclk));
	jnot g04927(.din(w_n4970_0[0]),.dout(n5152),.clk(gclk));
	jnot g04928(.din(w_n4963_0[0]),.dout(n5153),.clk(gclk));
	jnot g04929(.din(w_n4956_0[0]),.dout(n5154),.clk(gclk));
	jnot g04930(.din(w_n4949_0[0]),.dout(n5155),.clk(gclk));
	jnot g04931(.din(w_n4941_0[0]),.dout(n5156),.clk(gclk));
	jnot g04932(.din(w_n4933_0[0]),.dout(n5157),.clk(gclk));
	jnot g04933(.din(w_n4922_0[0]),.dout(n5158),.clk(gclk));
	jnot g04934(.din(w_n4914_0[0]),.dout(n5159),.clk(gclk));
	jand g04935(.dina(w_asqrt37_27[0]),.dinb(w_a74_0[2]),.dout(n5160),.clk(gclk));
	jor g04936(.dina(w_n4911_0[0]),.dinb(n5160),.dout(n5161),.clk(gclk));
	jor g04937(.dina(n5161),.dinb(w_asqrt38_31[0]),.dout(n5162),.clk(gclk));
	jand g04938(.dina(w_asqrt37_26[2]),.dinb(w_n4457_0[1]),.dout(n5163),.clk(gclk));
	jor g04939(.dina(n5163),.dinb(w_n4458_0[0]),.dout(n5164),.clk(gclk));
	jand g04940(.dina(w_n4925_0[0]),.dinb(n5164),.dout(n5165),.clk(gclk));
	jand g04941(.dina(w_n5165_0[1]),.dinb(n5162),.dout(n5166),.clk(gclk));
	jor g04942(.dina(n5166),.dinb(n5159),.dout(n5167),.clk(gclk));
	jor g04943(.dina(n5167),.dinb(w_asqrt39_27[2]),.dout(n5168),.clk(gclk));
	jnot g04944(.din(w_n4930_0[1]),.dout(n5169),.clk(gclk));
	jand g04945(.dina(n5169),.dinb(n5168),.dout(n5170),.clk(gclk));
	jor g04946(.dina(n5170),.dinb(n5158),.dout(n5171),.clk(gclk));
	jor g04947(.dina(n5171),.dinb(w_asqrt40_31[0]),.dout(n5172),.clk(gclk));
	jand g04948(.dina(w_n4937_0[1]),.dinb(n5172),.dout(n5173),.clk(gclk));
	jor g04949(.dina(n5173),.dinb(n5157),.dout(n5174),.clk(gclk));
	jor g04950(.dina(n5174),.dinb(w_asqrt41_28[0]),.dout(n5175),.clk(gclk));
	jand g04951(.dina(w_n4945_0[1]),.dinb(n5175),.dout(n5176),.clk(gclk));
	jor g04952(.dina(n5176),.dinb(n5156),.dout(n5177),.clk(gclk));
	jor g04953(.dina(n5177),.dinb(w_asqrt42_31[1]),.dout(n5178),.clk(gclk));
	jnot g04954(.din(w_n4953_0[0]),.dout(n5179),.clk(gclk));
	jand g04955(.dina(w_n5179_0[1]),.dinb(n5178),.dout(n5180),.clk(gclk));
	jor g04956(.dina(n5180),.dinb(n5155),.dout(n5181),.clk(gclk));
	jor g04957(.dina(n5181),.dinb(w_asqrt43_28[1]),.dout(n5182),.clk(gclk));
	jnot g04958(.din(w_n4960_0[1]),.dout(n5183),.clk(gclk));
	jand g04959(.dina(n5183),.dinb(n5182),.dout(n5184),.clk(gclk));
	jor g04960(.dina(n5184),.dinb(n5154),.dout(n5185),.clk(gclk));
	jor g04961(.dina(n5185),.dinb(w_asqrt44_31[1]),.dout(n5186),.clk(gclk));
	jnot g04962(.din(w_n4967_0[1]),.dout(n5187),.clk(gclk));
	jand g04963(.dina(n5187),.dinb(n5186),.dout(n5188),.clk(gclk));
	jor g04964(.dina(n5188),.dinb(n5153),.dout(n5189),.clk(gclk));
	jor g04965(.dina(n5189),.dinb(w_asqrt45_29[0]),.dout(n5190),.clk(gclk));
	jnot g04966(.din(w_n4974_0[1]),.dout(n5191),.clk(gclk));
	jand g04967(.dina(n5191),.dinb(n5190),.dout(n5192),.clk(gclk));
	jor g04968(.dina(n5192),.dinb(n5152),.dout(n5193),.clk(gclk));
	jor g04969(.dina(n5193),.dinb(w_asqrt46_31[1]),.dout(n5194),.clk(gclk));
	jand g04970(.dina(w_n4981_0[1]),.dinb(n5194),.dout(n5195),.clk(gclk));
	jor g04971(.dina(n5195),.dinb(n5151),.dout(n5196),.clk(gclk));
	jor g04972(.dina(n5196),.dinb(w_asqrt47_29[2]),.dout(n5197),.clk(gclk));
	jnot g04973(.din(w_n4989_0[1]),.dout(n5198),.clk(gclk));
	jand g04974(.dina(n5198),.dinb(n5197),.dout(n5199),.clk(gclk));
	jor g04975(.dina(n5199),.dinb(n5150),.dout(n5200),.clk(gclk));
	jor g04976(.dina(n5200),.dinb(w_asqrt48_31[2]),.dout(n5201),.clk(gclk));
	jand g04977(.dina(w_n4996_0[1]),.dinb(n5201),.dout(n5202),.clk(gclk));
	jor g04978(.dina(n5202),.dinb(n5149),.dout(n5203),.clk(gclk));
	jor g04979(.dina(n5203),.dinb(w_asqrt49_30[0]),.dout(n5204),.clk(gclk));
	jnot g04980(.din(w_n5004_0[1]),.dout(n5205),.clk(gclk));
	jand g04981(.dina(n5205),.dinb(n5204),.dout(n5206),.clk(gclk));
	jor g04982(.dina(n5206),.dinb(n5148),.dout(n5207),.clk(gclk));
	jor g04983(.dina(n5207),.dinb(w_asqrt50_32[0]),.dout(n5208),.clk(gclk));
	jand g04984(.dina(w_n5011_0[1]),.dinb(n5208),.dout(n5209),.clk(gclk));
	jor g04985(.dina(n5209),.dinb(n5147),.dout(n5210),.clk(gclk));
	jor g04986(.dina(n5210),.dinb(w_asqrt51_30[1]),.dout(n5211),.clk(gclk));
	jand g04987(.dina(w_n5019_0[1]),.dinb(n5211),.dout(n5212),.clk(gclk));
	jor g04988(.dina(n5212),.dinb(n5146),.dout(n5213),.clk(gclk));
	jor g04989(.dina(n5213),.dinb(w_asqrt52_32[0]),.dout(n5214),.clk(gclk));
	jnot g04990(.din(w_n5027_0[1]),.dout(n5215),.clk(gclk));
	jand g04991(.dina(n5215),.dinb(n5214),.dout(n5216),.clk(gclk));
	jor g04992(.dina(n5216),.dinb(n5145),.dout(n5217),.clk(gclk));
	jor g04993(.dina(n5217),.dinb(w_asqrt53_31[0]),.dout(n5218),.clk(gclk));
	jnot g04994(.din(w_n5034_0[1]),.dout(n5219),.clk(gclk));
	jand g04995(.dina(n5219),.dinb(n5218),.dout(n5220),.clk(gclk));
	jor g04996(.dina(n5220),.dinb(n5144),.dout(n5221),.clk(gclk));
	jor g04997(.dina(n5221),.dinb(w_asqrt54_32[0]),.dout(n5222),.clk(gclk));
	jand g04998(.dina(w_n5041_0[1]),.dinb(n5222),.dout(n5223),.clk(gclk));
	jor g04999(.dina(n5223),.dinb(n5143),.dout(n5224),.clk(gclk));
	jor g05000(.dina(n5224),.dinb(w_asqrt55_31[1]),.dout(n5225),.clk(gclk));
	jnot g05001(.din(w_n5049_0[1]),.dout(n5226),.clk(gclk));
	jand g05002(.dina(n5226),.dinb(n5225),.dout(n5227),.clk(gclk));
	jor g05003(.dina(n5227),.dinb(n5142),.dout(n5228),.clk(gclk));
	jor g05004(.dina(n5228),.dinb(w_asqrt56_32[1]),.dout(n5229),.clk(gclk));
	jand g05005(.dina(w_n5056_0[1]),.dinb(n5229),.dout(n5230),.clk(gclk));
	jor g05006(.dina(n5230),.dinb(n5141),.dout(n5231),.clk(gclk));
	jor g05007(.dina(n5231),.dinb(w_asqrt57_32[0]),.dout(n5232),.clk(gclk));
	jnot g05008(.din(w_n5064_0[1]),.dout(n5233),.clk(gclk));
	jand g05009(.dina(n5233),.dinb(n5232),.dout(n5234),.clk(gclk));
	jor g05010(.dina(n5234),.dinb(n5140),.dout(n5235),.clk(gclk));
	jor g05011(.dina(n5235),.dinb(w_asqrt58_32[2]),.dout(n5236),.clk(gclk));
	jand g05012(.dina(w_n5071_0[0]),.dinb(n5236),.dout(n5237),.clk(gclk));
	jor g05013(.dina(n5237),.dinb(n5139),.dout(n5238),.clk(gclk));
	jor g05014(.dina(n5238),.dinb(w_asqrt59_32[1]),.dout(n5239),.clk(gclk));
	jnot g05015(.din(w_n5079_0[1]),.dout(n5240),.clk(gclk));
	jand g05016(.dina(n5240),.dinb(n5239),.dout(n5241),.clk(gclk));
	jor g05017(.dina(n5241),.dinb(n5138),.dout(n5242),.clk(gclk));
	jor g05018(.dina(n5242),.dinb(w_asqrt60_32[2]),.dout(n5243),.clk(gclk));
	jand g05019(.dina(w_n5086_0[1]),.dinb(n5243),.dout(n5244),.clk(gclk));
	jor g05020(.dina(n5244),.dinb(n5137),.dout(n5245),.clk(gclk));
	jor g05021(.dina(n5245),.dinb(w_asqrt61_32[2]),.dout(n5246),.clk(gclk));
	jnot g05022(.din(w_n5094_0[1]),.dout(n5247),.clk(gclk));
	jand g05023(.dina(n5247),.dinb(n5246),.dout(n5248),.clk(gclk));
	jor g05024(.dina(n5248),.dinb(n5136),.dout(n5249),.clk(gclk));
	jor g05025(.dina(n5249),.dinb(w_asqrt62_32[2]),.dout(n5250),.clk(gclk));
	jand g05026(.dina(w_n5101_0[0]),.dinb(n5250),.dout(n5251),.clk(gclk));
	jor g05027(.dina(n5251),.dinb(n5135),.dout(n5252),.clk(gclk));
	jand g05028(.dina(n5252),.dinb(w_n4905_0[0]),.dout(n5253),.clk(gclk));
	jand g05029(.dina(w_n5253_0[1]),.dinb(w_n4766_0[1]),.dout(n5254),.clk(gclk));
	jand g05030(.dina(n5254),.dinb(n5134),.dout(n5255),.clk(gclk));
	jor g05031(.dina(n5255),.dinb(w_asqrt63_41[2]),.dout(n5256),.clk(gclk));
	jand g05032(.dina(w_n5116_0[0]),.dinb(w_n5256_0[1]),.dout(n5257),.clk(gclk));
	jand g05033(.dina(w_n5257_0[1]),.dinb(w_n5132_1[1]),.dout(n5259),.clk(gclk));
	jor g05034(.dina(w_n5259_45[1]),.dinb(n5131),.dout(n5260),.clk(gclk));
	jand g05035(.dina(n5260),.dinb(n5130),.dout(n5261),.clk(gclk));
	jand g05036(.dina(n5261),.dinb(n5128),.dout(n5262),.clk(gclk));
	jor g05037(.dina(n5262),.dinb(w_n5127_0[1]),.dout(n5263),.clk(gclk));
	jand g05038(.dina(w_n5263_0[2]),.dinb(w_asqrt38_30[2]),.dout(n5264),.clk(gclk));
	jor g05039(.dina(w_n5263_0[1]),.dinb(w_asqrt38_30[1]),.dout(n5265),.clk(gclk));
	jand g05040(.dina(w_asqrt36_38[1]),.dinb(w_n4910_0[0]),.dout(n5266),.clk(gclk));
	jand g05041(.dina(w_n5115_0[0]),.dinb(w_n5132_1[0]),.dout(n5267),.clk(gclk));
	jand g05042(.dina(n5267),.dinb(w_n5256_0[0]),.dout(n5268),.clk(gclk));
	jand g05043(.dina(n5268),.dinb(w_asqrt37_26[1]),.dout(n5269),.clk(gclk));
	jor g05044(.dina(n5269),.dinb(w_n5266_0[1]),.dout(n5270),.clk(gclk));
	jxor g05045(.dina(n5270),.dinb(w_a74_0[1]),.dout(n5271),.clk(gclk));
	jnot g05046(.din(w_n5271_0[1]),.dout(n5272),.clk(gclk));
	jand g05047(.dina(w_n5272_0[1]),.dinb(n5265),.dout(n5273),.clk(gclk));
	jor g05048(.dina(n5273),.dinb(w_n5264_0[1]),.dout(n5274),.clk(gclk));
	jand g05049(.dina(w_n5274_0[2]),.dinb(w_asqrt39_27[1]),.dout(n5275),.clk(gclk));
	jor g05050(.dina(w_n5274_0[1]),.dinb(w_asqrt39_27[0]),.dout(n5276),.clk(gclk));
	jxor g05051(.dina(w_n4913_0[0]),.dinb(w_n4582_45[2]),.dout(n5277),.clk(gclk));
	jand g05052(.dina(n5277),.dinb(w_asqrt36_38[0]),.dout(n5278),.clk(gclk));
	jxor g05053(.dina(n5278),.dinb(w_n5165_0[0]),.dout(n5279),.clk(gclk));
	jand g05054(.dina(w_n5279_0[1]),.dinb(n5276),.dout(n5280),.clk(gclk));
	jor g05055(.dina(n5280),.dinb(w_n5275_0[1]),.dout(n5281),.clk(gclk));
	jand g05056(.dina(w_n5281_0[2]),.dinb(w_asqrt40_30[2]),.dout(n5282),.clk(gclk));
	jor g05057(.dina(w_n5281_0[1]),.dinb(w_asqrt40_30[1]),.dout(n5283),.clk(gclk));
	jxor g05058(.dina(w_n4921_0[0]),.dinb(w_n4249_49[1]),.dout(n5284),.clk(gclk));
	jand g05059(.dina(n5284),.dinb(w_asqrt36_37[2]),.dout(n5285),.clk(gclk));
	jxor g05060(.dina(n5285),.dinb(w_n4930_0[0]),.dout(n5286),.clk(gclk));
	jnot g05061(.din(w_n5286_0[1]),.dout(n5287),.clk(gclk));
	jand g05062(.dina(w_n5287_0[1]),.dinb(n5283),.dout(n5288),.clk(gclk));
	jor g05063(.dina(n5288),.dinb(w_n5282_0[1]),.dout(n5289),.clk(gclk));
	jand g05064(.dina(w_n5289_0[2]),.dinb(w_asqrt41_27[2]),.dout(n5290),.clk(gclk));
	jor g05065(.dina(w_n5289_0[1]),.dinb(w_asqrt41_27[1]),.dout(n5291),.clk(gclk));
	jxor g05066(.dina(w_n4932_0[0]),.dinb(w_n3955_46[1]),.dout(n5292),.clk(gclk));
	jand g05067(.dina(n5292),.dinb(w_asqrt36_37[1]),.dout(n5293),.clk(gclk));
	jxor g05068(.dina(n5293),.dinb(w_n4937_0[0]),.dout(n5294),.clk(gclk));
	jand g05069(.dina(w_n5294_0[1]),.dinb(n5291),.dout(n5295),.clk(gclk));
	jor g05070(.dina(n5295),.dinb(w_n5290_0[1]),.dout(n5296),.clk(gclk));
	jand g05071(.dina(w_n5296_0[2]),.dinb(w_asqrt42_31[0]),.dout(n5297),.clk(gclk));
	jor g05072(.dina(w_n5296_0[1]),.dinb(w_asqrt42_30[2]),.dout(n5298),.clk(gclk));
	jxor g05073(.dina(w_n4940_0[0]),.dinb(w_n3642_49[2]),.dout(n5299),.clk(gclk));
	jand g05074(.dina(n5299),.dinb(w_asqrt36_37[0]),.dout(n5300),.clk(gclk));
	jxor g05075(.dina(n5300),.dinb(w_n4945_0[0]),.dout(n5301),.clk(gclk));
	jand g05076(.dina(w_n5301_0[1]),.dinb(n5298),.dout(n5302),.clk(gclk));
	jor g05077(.dina(n5302),.dinb(w_n5297_0[1]),.dout(n5303),.clk(gclk));
	jand g05078(.dina(w_n5303_0[2]),.dinb(w_asqrt43_28[0]),.dout(n5304),.clk(gclk));
	jor g05079(.dina(w_n5303_0[1]),.dinb(w_asqrt43_27[2]),.dout(n5305),.clk(gclk));
	jxor g05080(.dina(w_n4948_0[0]),.dinb(w_n3368_47[0]),.dout(n5306),.clk(gclk));
	jand g05081(.dina(n5306),.dinb(w_asqrt36_36[2]),.dout(n5307),.clk(gclk));
	jxor g05082(.dina(n5307),.dinb(w_n5179_0[0]),.dout(n5308),.clk(gclk));
	jand g05083(.dina(w_n5308_0[1]),.dinb(n5305),.dout(n5309),.clk(gclk));
	jor g05084(.dina(n5309),.dinb(w_n5304_0[1]),.dout(n5310),.clk(gclk));
	jand g05085(.dina(w_n5310_0[2]),.dinb(w_asqrt44_31[0]),.dout(n5311),.clk(gclk));
	jor g05086(.dina(w_n5310_0[1]),.dinb(w_asqrt44_30[2]),.dout(n5312),.clk(gclk));
	jxor g05087(.dina(w_n4955_0[0]),.dinb(w_n3089_50[1]),.dout(n5313),.clk(gclk));
	jand g05088(.dina(n5313),.dinb(w_asqrt36_36[1]),.dout(n5314),.clk(gclk));
	jxor g05089(.dina(n5314),.dinb(w_n4960_0[0]),.dout(n5315),.clk(gclk));
	jnot g05090(.din(w_n5315_0[1]),.dout(n5316),.clk(gclk));
	jand g05091(.dina(w_n5316_0[1]),.dinb(n5312),.dout(n5317),.clk(gclk));
	jor g05092(.dina(n5317),.dinb(w_n5311_0[1]),.dout(n5318),.clk(gclk));
	jand g05093(.dina(w_n5318_0[2]),.dinb(w_asqrt45_28[2]),.dout(n5319),.clk(gclk));
	jor g05094(.dina(w_n5318_0[1]),.dinb(w_asqrt45_28[1]),.dout(n5320),.clk(gclk));
	jxor g05095(.dina(w_n4962_0[0]),.dinb(w_n2833_48[0]),.dout(n5321),.clk(gclk));
	jand g05096(.dina(n5321),.dinb(w_asqrt36_36[0]),.dout(n5322),.clk(gclk));
	jxor g05097(.dina(n5322),.dinb(w_n4967_0[0]),.dout(n5323),.clk(gclk));
	jnot g05098(.din(w_n5323_0[1]),.dout(n5324),.clk(gclk));
	jand g05099(.dina(w_n5324_0[1]),.dinb(n5320),.dout(n5325),.clk(gclk));
	jor g05100(.dina(n5325),.dinb(w_n5319_0[1]),.dout(n5326),.clk(gclk));
	jand g05101(.dina(w_n5326_0[2]),.dinb(w_asqrt46_31[0]),.dout(n5327),.clk(gclk));
	jor g05102(.dina(w_n5326_0[1]),.dinb(w_asqrt46_30[2]),.dout(n5328),.clk(gclk));
	jxor g05103(.dina(w_n4969_0[0]),.dinb(w_n2572_50[2]),.dout(n5329),.clk(gclk));
	jand g05104(.dina(n5329),.dinb(w_asqrt36_35[2]),.dout(n5330),.clk(gclk));
	jxor g05105(.dina(n5330),.dinb(w_n4974_0[0]),.dout(n5331),.clk(gclk));
	jnot g05106(.din(w_n5331_0[1]),.dout(n5332),.clk(gclk));
	jand g05107(.dina(w_n5332_0[1]),.dinb(n5328),.dout(n5333),.clk(gclk));
	jor g05108(.dina(n5333),.dinb(w_n5327_0[1]),.dout(n5334),.clk(gclk));
	jand g05109(.dina(w_n5334_0[2]),.dinb(w_asqrt47_29[1]),.dout(n5335),.clk(gclk));
	jor g05110(.dina(w_n5334_0[1]),.dinb(w_asqrt47_29[0]),.dout(n5336),.clk(gclk));
	jxor g05111(.dina(w_n4976_0[0]),.dinb(w_n2345_48[2]),.dout(n5337),.clk(gclk));
	jand g05112(.dina(n5337),.dinb(w_asqrt36_35[1]),.dout(n5338),.clk(gclk));
	jxor g05113(.dina(n5338),.dinb(w_n4981_0[0]),.dout(n5339),.clk(gclk));
	jand g05114(.dina(w_n5339_0[1]),.dinb(n5336),.dout(n5340),.clk(gclk));
	jor g05115(.dina(n5340),.dinb(w_n5335_0[1]),.dout(n5341),.clk(gclk));
	jand g05116(.dina(w_n5341_0[2]),.dinb(w_asqrt48_31[1]),.dout(n5342),.clk(gclk));
	jor g05117(.dina(w_n5341_0[1]),.dinb(w_asqrt48_31[0]),.dout(n5343),.clk(gclk));
	jxor g05118(.dina(w_n4984_0[0]),.dinb(w_n2108_51[1]),.dout(n5344),.clk(gclk));
	jand g05119(.dina(n5344),.dinb(w_asqrt36_35[0]),.dout(n5345),.clk(gclk));
	jxor g05120(.dina(n5345),.dinb(w_n4989_0[0]),.dout(n5346),.clk(gclk));
	jnot g05121(.din(w_n5346_0[1]),.dout(n5347),.clk(gclk));
	jand g05122(.dina(w_n5347_0[1]),.dinb(n5343),.dout(n5348),.clk(gclk));
	jor g05123(.dina(n5348),.dinb(w_n5342_0[1]),.dout(n5349),.clk(gclk));
	jand g05124(.dina(w_n5349_0[2]),.dinb(w_asqrt49_29[2]),.dout(n5350),.clk(gclk));
	jor g05125(.dina(w_n5349_0[1]),.dinb(w_asqrt49_29[1]),.dout(n5351),.clk(gclk));
	jxor g05126(.dina(w_n4991_0[0]),.dinb(w_n1912_49[2]),.dout(n5352),.clk(gclk));
	jand g05127(.dina(n5352),.dinb(w_asqrt36_34[2]),.dout(n5353),.clk(gclk));
	jxor g05128(.dina(n5353),.dinb(w_n4996_0[0]),.dout(n5354),.clk(gclk));
	jand g05129(.dina(w_n5354_0[1]),.dinb(n5351),.dout(n5355),.clk(gclk));
	jor g05130(.dina(n5355),.dinb(w_n5350_0[1]),.dout(n5356),.clk(gclk));
	jand g05131(.dina(w_n5356_0[2]),.dinb(w_asqrt50_31[2]),.dout(n5357),.clk(gclk));
	jor g05132(.dina(w_n5356_0[1]),.dinb(w_asqrt50_31[1]),.dout(n5358),.clk(gclk));
	jxor g05133(.dina(w_n4999_0[0]),.dinb(w_n1699_52[0]),.dout(n5359),.clk(gclk));
	jand g05134(.dina(n5359),.dinb(w_asqrt36_34[1]),.dout(n5360),.clk(gclk));
	jxor g05135(.dina(n5360),.dinb(w_n5004_0[0]),.dout(n5361),.clk(gclk));
	jnot g05136(.din(w_n5361_0[1]),.dout(n5362),.clk(gclk));
	jand g05137(.dina(w_n5362_0[1]),.dinb(n5358),.dout(n5363),.clk(gclk));
	jor g05138(.dina(n5363),.dinb(w_n5357_0[1]),.dout(n5364),.clk(gclk));
	jand g05139(.dina(w_n5364_0[2]),.dinb(w_asqrt51_30[0]),.dout(n5365),.clk(gclk));
	jor g05140(.dina(w_n5364_0[1]),.dinb(w_asqrt51_29[2]),.dout(n5366),.clk(gclk));
	jxor g05141(.dina(w_n5006_0[0]),.dinb(w_n1516_50[1]),.dout(n5367),.clk(gclk));
	jand g05142(.dina(n5367),.dinb(w_asqrt36_34[0]),.dout(n5368),.clk(gclk));
	jxor g05143(.dina(n5368),.dinb(w_n5011_0[0]),.dout(n5369),.clk(gclk));
	jand g05144(.dina(w_n5369_0[1]),.dinb(n5366),.dout(n5370),.clk(gclk));
	jor g05145(.dina(n5370),.dinb(w_n5365_0[1]),.dout(n5371),.clk(gclk));
	jand g05146(.dina(w_n5371_0[2]),.dinb(w_asqrt52_31[2]),.dout(n5372),.clk(gclk));
	jor g05147(.dina(w_n5371_0[1]),.dinb(w_asqrt52_31[1]),.dout(n5373),.clk(gclk));
	jxor g05148(.dina(w_n5014_0[0]),.dinb(w_n1332_52[0]),.dout(n5374),.clk(gclk));
	jand g05149(.dina(n5374),.dinb(w_asqrt36_33[2]),.dout(n5375),.clk(gclk));
	jxor g05150(.dina(n5375),.dinb(w_n5019_0[0]),.dout(n5376),.clk(gclk));
	jand g05151(.dina(w_n5376_0[1]),.dinb(n5373),.dout(n5377),.clk(gclk));
	jor g05152(.dina(n5377),.dinb(w_n5372_0[1]),.dout(n5378),.clk(gclk));
	jand g05153(.dina(w_n5378_0[2]),.dinb(w_asqrt53_30[2]),.dout(n5379),.clk(gclk));
	jor g05154(.dina(w_n5378_0[1]),.dinb(w_asqrt53_30[1]),.dout(n5380),.clk(gclk));
	jxor g05155(.dina(w_n5022_0[0]),.dinb(w_n1173_51[0]),.dout(n5381),.clk(gclk));
	jand g05156(.dina(n5381),.dinb(w_asqrt36_33[1]),.dout(n5382),.clk(gclk));
	jxor g05157(.dina(n5382),.dinb(w_n5027_0[0]),.dout(n5383),.clk(gclk));
	jnot g05158(.din(w_n5383_0[1]),.dout(n5384),.clk(gclk));
	jand g05159(.dina(w_n5384_0[1]),.dinb(n5380),.dout(n5385),.clk(gclk));
	jor g05160(.dina(n5385),.dinb(w_n5379_0[1]),.dout(n5386),.clk(gclk));
	jand g05161(.dina(w_n5386_0[2]),.dinb(w_asqrt54_31[2]),.dout(n5387),.clk(gclk));
	jor g05162(.dina(w_n5386_0[1]),.dinb(w_asqrt54_31[1]),.dout(n5388),.clk(gclk));
	jxor g05163(.dina(w_n5029_0[0]),.dinb(w_n1008_53[0]),.dout(n5389),.clk(gclk));
	jand g05164(.dina(n5389),.dinb(w_asqrt36_33[0]),.dout(n5390),.clk(gclk));
	jxor g05165(.dina(n5390),.dinb(w_n5034_0[0]),.dout(n5391),.clk(gclk));
	jnot g05166(.din(w_n5391_0[1]),.dout(n5392),.clk(gclk));
	jand g05167(.dina(w_n5392_0[1]),.dinb(n5388),.dout(n5393),.clk(gclk));
	jor g05168(.dina(n5393),.dinb(w_n5387_0[1]),.dout(n5394),.clk(gclk));
	jand g05169(.dina(w_n5394_0[2]),.dinb(w_asqrt55_31[0]),.dout(n5395),.clk(gclk));
	jor g05170(.dina(w_n5394_0[1]),.dinb(w_asqrt55_30[2]),.dout(n5396),.clk(gclk));
	jxor g05171(.dina(w_n5036_0[0]),.dinb(w_n884_52[0]),.dout(n5397),.clk(gclk));
	jand g05172(.dina(n5397),.dinb(w_asqrt36_32[2]),.dout(n5398),.clk(gclk));
	jxor g05173(.dina(n5398),.dinb(w_n5041_0[0]),.dout(n5399),.clk(gclk));
	jand g05174(.dina(w_n5399_0[1]),.dinb(n5396),.dout(n5400),.clk(gclk));
	jor g05175(.dina(n5400),.dinb(w_n5395_0[1]),.dout(n5401),.clk(gclk));
	jand g05176(.dina(w_n5401_0[2]),.dinb(w_asqrt56_32[0]),.dout(n5402),.clk(gclk));
	jor g05177(.dina(w_n5401_0[1]),.dinb(w_asqrt56_31[2]),.dout(n5403),.clk(gclk));
	jxor g05178(.dina(w_n5044_0[0]),.dinb(w_n743_53[0]),.dout(n5404),.clk(gclk));
	jand g05179(.dina(n5404),.dinb(w_asqrt36_32[1]),.dout(n5405),.clk(gclk));
	jxor g05180(.dina(n5405),.dinb(w_n5049_0[0]),.dout(n5406),.clk(gclk));
	jnot g05181(.din(w_n5406_0[1]),.dout(n5407),.clk(gclk));
	jand g05182(.dina(w_n5407_0[1]),.dinb(n5403),.dout(n5408),.clk(gclk));
	jor g05183(.dina(n5408),.dinb(w_n5402_0[1]),.dout(n5409),.clk(gclk));
	jand g05184(.dina(w_n5409_0[2]),.dinb(w_asqrt57_31[2]),.dout(n5410),.clk(gclk));
	jor g05185(.dina(w_n5409_0[1]),.dinb(w_asqrt57_31[1]),.dout(n5411),.clk(gclk));
	jxor g05186(.dina(w_n5051_0[0]),.dinb(w_n635_53[0]),.dout(n5412),.clk(gclk));
	jand g05187(.dina(n5412),.dinb(w_asqrt36_32[0]),.dout(n5413),.clk(gclk));
	jxor g05188(.dina(n5413),.dinb(w_n5056_0[0]),.dout(n5414),.clk(gclk));
	jand g05189(.dina(w_n5414_0[1]),.dinb(n5411),.dout(n5415),.clk(gclk));
	jor g05190(.dina(n5415),.dinb(w_n5410_0[1]),.dout(n5416),.clk(gclk));
	jand g05191(.dina(w_n5416_0[2]),.dinb(w_asqrt58_32[1]),.dout(n5417),.clk(gclk));
	jor g05192(.dina(w_n5416_0[1]),.dinb(w_asqrt58_32[0]),.dout(n5418),.clk(gclk));
	jxor g05193(.dina(w_n5059_0[0]),.dinb(w_n515_54[0]),.dout(n5419),.clk(gclk));
	jand g05194(.dina(n5419),.dinb(w_asqrt36_31[2]),.dout(n5420),.clk(gclk));
	jxor g05195(.dina(n5420),.dinb(w_n5064_0[0]),.dout(n5421),.clk(gclk));
	jnot g05196(.din(w_n5421_0[1]),.dout(n5422),.clk(gclk));
	jand g05197(.dina(w_n5422_0[1]),.dinb(n5418),.dout(n5423),.clk(gclk));
	jor g05198(.dina(n5423),.dinb(w_n5417_0[1]),.dout(n5424),.clk(gclk));
	jand g05199(.dina(w_n5424_0[2]),.dinb(w_asqrt59_32[0]),.dout(n5425),.clk(gclk));
	jor g05200(.dina(w_n5424_0[1]),.dinb(w_asqrt59_31[2]),.dout(n5426),.clk(gclk));
	jxor g05201(.dina(w_n5066_0[0]),.dinb(w_n443_54[0]),.dout(n5427),.clk(gclk));
	jand g05202(.dina(n5427),.dinb(w_asqrt36_31[1]),.dout(n5428),.clk(gclk));
	jxor g05203(.dina(n5428),.dinb(w_n5072_0[0]),.dout(n5429),.clk(gclk));
	jnot g05204(.din(w_n5429_0[1]),.dout(n5430),.clk(gclk));
	jand g05205(.dina(w_n5430_0[1]),.dinb(n5426),.dout(n5431),.clk(gclk));
	jor g05206(.dina(n5431),.dinb(w_n5425_0[1]),.dout(n5432),.clk(gclk));
	jand g05207(.dina(w_n5432_0[2]),.dinb(w_asqrt60_32[1]),.dout(n5433),.clk(gclk));
	jor g05208(.dina(w_n5432_0[1]),.dinb(w_asqrt60_32[0]),.dout(n5434),.clk(gclk));
	jxor g05209(.dina(w_n5074_0[0]),.dinb(w_n352_54[1]),.dout(n5435),.clk(gclk));
	jand g05210(.dina(n5435),.dinb(w_asqrt36_31[0]),.dout(n5436),.clk(gclk));
	jxor g05211(.dina(n5436),.dinb(w_n5079_0[0]),.dout(n5437),.clk(gclk));
	jnot g05212(.din(w_n5437_0[1]),.dout(n5438),.clk(gclk));
	jand g05213(.dina(w_n5438_0[1]),.dinb(n5434),.dout(n5439),.clk(gclk));
	jor g05214(.dina(n5439),.dinb(w_n5433_0[1]),.dout(n5440),.clk(gclk));
	jand g05215(.dina(w_n5440_0[2]),.dinb(w_asqrt61_32[1]),.dout(n5441),.clk(gclk));
	jor g05216(.dina(w_n5440_0[1]),.dinb(w_asqrt61_32[0]),.dout(n5442),.clk(gclk));
	jxor g05217(.dina(w_n5081_0[0]),.dinb(w_n294_54[2]),.dout(n5443),.clk(gclk));
	jand g05218(.dina(n5443),.dinb(w_asqrt36_30[2]),.dout(n5444),.clk(gclk));
	jxor g05219(.dina(n5444),.dinb(w_n5086_0[0]),.dout(n5445),.clk(gclk));
	jand g05220(.dina(w_n5445_0[1]),.dinb(n5442),.dout(n5446),.clk(gclk));
	jor g05221(.dina(n5446),.dinb(w_n5441_0[1]),.dout(n5447),.clk(gclk));
	jand g05222(.dina(w_n5447_0[2]),.dinb(w_asqrt62_32[1]),.dout(n5448),.clk(gclk));
	jor g05223(.dina(w_n5447_0[1]),.dinb(w_asqrt62_32[0]),.dout(n5449),.clk(gclk));
	jxor g05224(.dina(w_n5089_0[0]),.dinb(w_n239_54[2]),.dout(n5450),.clk(gclk));
	jand g05225(.dina(n5450),.dinb(w_asqrt36_30[1]),.dout(n5451),.clk(gclk));
	jxor g05226(.dina(n5451),.dinb(w_n5094_0[0]),.dout(n5452),.clk(gclk));
	jnot g05227(.din(w_n5452_0[2]),.dout(n5453),.clk(gclk));
	jand g05228(.dina(n5453),.dinb(n5449),.dout(n5454),.clk(gclk));
	jor g05229(.dina(n5454),.dinb(w_n5448_0[1]),.dout(n5455),.clk(gclk));
	jxor g05230(.dina(w_n5096_0[0]),.dinb(w_n221_55[0]),.dout(n5456),.clk(gclk));
	jand g05231(.dina(n5456),.dinb(w_asqrt36_30[0]),.dout(n5457),.clk(gclk));
	jxor g05232(.dina(n5457),.dinb(w_n5102_0[0]),.dout(n5458),.clk(gclk));
	jnot g05233(.din(w_n5458_0[1]),.dout(n5459),.clk(gclk));
	jor g05234(.dina(w_n5459_0[2]),.dinb(w_n5455_0[2]),.dout(n5460),.clk(gclk));
	jnot g05235(.din(w_n5460_0[1]),.dout(n5461),.clk(gclk));
	jand g05236(.dina(w_n5257_0[0]),.dinb(w_n5104_0[0]),.dout(n5462),.clk(gclk));
	jnot g05237(.din(n5462),.dout(n5463),.clk(gclk));
	jand g05238(.dina(w_n5108_0[0]),.dinb(w_asqrt63_41[1]),.dout(n5464),.clk(gclk));
	jand g05239(.dina(n5464),.dinb(w_n5132_0[2]),.dout(n5465),.clk(gclk));
	jand g05240(.dina(w_n5465_0[1]),.dinb(n5463),.dout(n5466),.clk(gclk));
	jand g05241(.dina(w_n5118_0[0]),.dinb(w_n5253_0[0]),.dout(n5467),.clk(gclk));
	jnot g05242(.din(w_n5448_0[0]),.dout(n5468),.clk(gclk));
	jnot g05243(.din(w_n5441_0[0]),.dout(n5469),.clk(gclk));
	jnot g05244(.din(w_n5433_0[0]),.dout(n5470),.clk(gclk));
	jnot g05245(.din(w_n5425_0[0]),.dout(n5471),.clk(gclk));
	jnot g05246(.din(w_n5417_0[0]),.dout(n5472),.clk(gclk));
	jnot g05247(.din(w_n5410_0[0]),.dout(n5473),.clk(gclk));
	jnot g05248(.din(w_n5402_0[0]),.dout(n5474),.clk(gclk));
	jnot g05249(.din(w_n5395_0[0]),.dout(n5475),.clk(gclk));
	jnot g05250(.din(w_n5387_0[0]),.dout(n5476),.clk(gclk));
	jnot g05251(.din(w_n5379_0[0]),.dout(n5477),.clk(gclk));
	jnot g05252(.din(w_n5372_0[0]),.dout(n5478),.clk(gclk));
	jnot g05253(.din(w_n5365_0[0]),.dout(n5479),.clk(gclk));
	jnot g05254(.din(w_n5357_0[0]),.dout(n5480),.clk(gclk));
	jnot g05255(.din(w_n5350_0[0]),.dout(n5481),.clk(gclk));
	jnot g05256(.din(w_n5342_0[0]),.dout(n5482),.clk(gclk));
	jnot g05257(.din(w_n5335_0[0]),.dout(n5483),.clk(gclk));
	jnot g05258(.din(w_n5327_0[0]),.dout(n5484),.clk(gclk));
	jnot g05259(.din(w_n5319_0[0]),.dout(n5485),.clk(gclk));
	jnot g05260(.din(w_n5311_0[0]),.dout(n5486),.clk(gclk));
	jnot g05261(.din(w_n5304_0[0]),.dout(n5487),.clk(gclk));
	jnot g05262(.din(w_n5297_0[0]),.dout(n5488),.clk(gclk));
	jnot g05263(.din(w_n5290_0[0]),.dout(n5489),.clk(gclk));
	jnot g05264(.din(w_n5282_0[0]),.dout(n5490),.clk(gclk));
	jnot g05265(.din(w_n5275_0[0]),.dout(n5491),.clk(gclk));
	jnot g05266(.din(w_n5264_0[0]),.dout(n5492),.clk(gclk));
	jnot g05267(.din(w_n5127_0[0]),.dout(n5493),.clk(gclk));
	jnot g05268(.din(w_n5124_0[0]),.dout(n5494),.clk(gclk));
	jor g05269(.dina(w_n5259_45[0]),.dinb(w_n4908_0[2]),.dout(n5495),.clk(gclk));
	jand g05270(.dina(n5495),.dinb(n5494),.dout(n5496),.clk(gclk));
	jand g05271(.dina(n5496),.dinb(w_n4902_48[1]),.dout(n5497),.clk(gclk));
	jor g05272(.dina(w_n5259_44[2]),.dinb(w_a72_0[0]),.dout(n5498),.clk(gclk));
	jand g05273(.dina(n5498),.dinb(w_a73_0[0]),.dout(n5499),.clk(gclk));
	jor g05274(.dina(w_n5266_0[0]),.dinb(n5499),.dout(n5500),.clk(gclk));
	jor g05275(.dina(w_n5500_0[1]),.dinb(n5497),.dout(n5501),.clk(gclk));
	jand g05276(.dina(n5501),.dinb(n5493),.dout(n5502),.clk(gclk));
	jand g05277(.dina(n5502),.dinb(w_n4582_45[1]),.dout(n5503),.clk(gclk));
	jor g05278(.dina(w_n5271_0[0]),.dinb(n5503),.dout(n5504),.clk(gclk));
	jand g05279(.dina(n5504),.dinb(n5492),.dout(n5505),.clk(gclk));
	jand g05280(.dina(n5505),.dinb(w_n4249_49[0]),.dout(n5506),.clk(gclk));
	jnot g05281(.din(w_n5279_0[0]),.dout(n5507),.clk(gclk));
	jor g05282(.dina(w_n5507_0[1]),.dinb(n5506),.dout(n5508),.clk(gclk));
	jand g05283(.dina(n5508),.dinb(n5491),.dout(n5509),.clk(gclk));
	jand g05284(.dina(n5509),.dinb(w_n3955_46[0]),.dout(n5510),.clk(gclk));
	jor g05285(.dina(w_n5286_0[0]),.dinb(n5510),.dout(n5511),.clk(gclk));
	jand g05286(.dina(n5511),.dinb(n5490),.dout(n5512),.clk(gclk));
	jand g05287(.dina(n5512),.dinb(w_n3642_49[1]),.dout(n5513),.clk(gclk));
	jnot g05288(.din(w_n5294_0[0]),.dout(n5514),.clk(gclk));
	jor g05289(.dina(w_n5514_0[1]),.dinb(n5513),.dout(n5515),.clk(gclk));
	jand g05290(.dina(n5515),.dinb(n5489),.dout(n5516),.clk(gclk));
	jand g05291(.dina(n5516),.dinb(w_n3368_46[2]),.dout(n5517),.clk(gclk));
	jnot g05292(.din(w_n5301_0[0]),.dout(n5518),.clk(gclk));
	jor g05293(.dina(w_n5518_0[1]),.dinb(n5517),.dout(n5519),.clk(gclk));
	jand g05294(.dina(n5519),.dinb(n5488),.dout(n5520),.clk(gclk));
	jand g05295(.dina(n5520),.dinb(w_n3089_50[0]),.dout(n5521),.clk(gclk));
	jnot g05296(.din(w_n5308_0[0]),.dout(n5522),.clk(gclk));
	jor g05297(.dina(w_n5522_0[1]),.dinb(n5521),.dout(n5523),.clk(gclk));
	jand g05298(.dina(n5523),.dinb(n5487),.dout(n5524),.clk(gclk));
	jand g05299(.dina(n5524),.dinb(w_n2833_47[2]),.dout(n5525),.clk(gclk));
	jor g05300(.dina(w_n5315_0[0]),.dinb(n5525),.dout(n5526),.clk(gclk));
	jand g05301(.dina(n5526),.dinb(n5486),.dout(n5527),.clk(gclk));
	jand g05302(.dina(n5527),.dinb(w_n2572_50[1]),.dout(n5528),.clk(gclk));
	jor g05303(.dina(w_n5323_0[0]),.dinb(n5528),.dout(n5529),.clk(gclk));
	jand g05304(.dina(n5529),.dinb(n5485),.dout(n5530),.clk(gclk));
	jand g05305(.dina(n5530),.dinb(w_n2345_48[1]),.dout(n5531),.clk(gclk));
	jor g05306(.dina(w_n5331_0[0]),.dinb(n5531),.dout(n5532),.clk(gclk));
	jand g05307(.dina(n5532),.dinb(n5484),.dout(n5533),.clk(gclk));
	jand g05308(.dina(n5533),.dinb(w_n2108_51[0]),.dout(n5534),.clk(gclk));
	jnot g05309(.din(w_n5339_0[0]),.dout(n5535),.clk(gclk));
	jor g05310(.dina(w_n5535_0[1]),.dinb(n5534),.dout(n5536),.clk(gclk));
	jand g05311(.dina(n5536),.dinb(n5483),.dout(n5537),.clk(gclk));
	jand g05312(.dina(n5537),.dinb(w_n1912_49[1]),.dout(n5538),.clk(gclk));
	jor g05313(.dina(w_n5346_0[0]),.dinb(n5538),.dout(n5539),.clk(gclk));
	jand g05314(.dina(n5539),.dinb(n5482),.dout(n5540),.clk(gclk));
	jand g05315(.dina(n5540),.dinb(w_n1699_51[2]),.dout(n5541),.clk(gclk));
	jnot g05316(.din(w_n5354_0[0]),.dout(n5542),.clk(gclk));
	jor g05317(.dina(w_n5542_0[1]),.dinb(n5541),.dout(n5543),.clk(gclk));
	jand g05318(.dina(n5543),.dinb(n5481),.dout(n5544),.clk(gclk));
	jand g05319(.dina(n5544),.dinb(w_n1516_50[0]),.dout(n5545),.clk(gclk));
	jor g05320(.dina(w_n5361_0[0]),.dinb(n5545),.dout(n5546),.clk(gclk));
	jand g05321(.dina(n5546),.dinb(n5480),.dout(n5547),.clk(gclk));
	jand g05322(.dina(n5547),.dinb(w_n1332_51[2]),.dout(n5548),.clk(gclk));
	jnot g05323(.din(w_n5369_0[0]),.dout(n5549),.clk(gclk));
	jor g05324(.dina(w_n5549_0[1]),.dinb(n5548),.dout(n5550),.clk(gclk));
	jand g05325(.dina(n5550),.dinb(n5479),.dout(n5551),.clk(gclk));
	jand g05326(.dina(n5551),.dinb(w_n1173_50[2]),.dout(n5552),.clk(gclk));
	jnot g05327(.din(w_n5376_0[0]),.dout(n5553),.clk(gclk));
	jor g05328(.dina(w_n5553_0[1]),.dinb(n5552),.dout(n5554),.clk(gclk));
	jand g05329(.dina(n5554),.dinb(n5478),.dout(n5555),.clk(gclk));
	jand g05330(.dina(n5555),.dinb(w_n1008_52[2]),.dout(n5556),.clk(gclk));
	jor g05331(.dina(w_n5383_0[0]),.dinb(n5556),.dout(n5557),.clk(gclk));
	jand g05332(.dina(n5557),.dinb(n5477),.dout(n5558),.clk(gclk));
	jand g05333(.dina(n5558),.dinb(w_n884_51[2]),.dout(n5559),.clk(gclk));
	jor g05334(.dina(w_n5391_0[0]),.dinb(n5559),.dout(n5560),.clk(gclk));
	jand g05335(.dina(n5560),.dinb(n5476),.dout(n5561),.clk(gclk));
	jand g05336(.dina(n5561),.dinb(w_n743_52[2]),.dout(n5562),.clk(gclk));
	jnot g05337(.din(w_n5399_0[0]),.dout(n5563),.clk(gclk));
	jor g05338(.dina(w_n5563_0[1]),.dinb(n5562),.dout(n5564),.clk(gclk));
	jand g05339(.dina(n5564),.dinb(n5475),.dout(n5565),.clk(gclk));
	jand g05340(.dina(n5565),.dinb(w_n635_52[2]),.dout(n5566),.clk(gclk));
	jor g05341(.dina(w_n5406_0[0]),.dinb(n5566),.dout(n5567),.clk(gclk));
	jand g05342(.dina(n5567),.dinb(n5474),.dout(n5568),.clk(gclk));
	jand g05343(.dina(n5568),.dinb(w_n515_53[2]),.dout(n5569),.clk(gclk));
	jnot g05344(.din(w_n5414_0[0]),.dout(n5570),.clk(gclk));
	jor g05345(.dina(w_n5570_0[1]),.dinb(n5569),.dout(n5571),.clk(gclk));
	jand g05346(.dina(n5571),.dinb(n5473),.dout(n5572),.clk(gclk));
	jand g05347(.dina(n5572),.dinb(w_n443_53[2]),.dout(n5573),.clk(gclk));
	jor g05348(.dina(w_n5421_0[0]),.dinb(n5573),.dout(n5574),.clk(gclk));
	jand g05349(.dina(n5574),.dinb(n5472),.dout(n5575),.clk(gclk));
	jand g05350(.dina(n5575),.dinb(w_n352_54[0]),.dout(n5576),.clk(gclk));
	jor g05351(.dina(w_n5429_0[0]),.dinb(n5576),.dout(n5577),.clk(gclk));
	jand g05352(.dina(n5577),.dinb(n5471),.dout(n5578),.clk(gclk));
	jand g05353(.dina(n5578),.dinb(w_n294_54[1]),.dout(n5579),.clk(gclk));
	jor g05354(.dina(w_n5437_0[0]),.dinb(n5579),.dout(n5580),.clk(gclk));
	jand g05355(.dina(n5580),.dinb(n5470),.dout(n5581),.clk(gclk));
	jand g05356(.dina(n5581),.dinb(w_n239_54[1]),.dout(n5582),.clk(gclk));
	jnot g05357(.din(w_n5445_0[0]),.dout(n5583),.clk(gclk));
	jor g05358(.dina(w_n5583_0[1]),.dinb(n5582),.dout(n5584),.clk(gclk));
	jand g05359(.dina(n5584),.dinb(n5469),.dout(n5585),.clk(gclk));
	jand g05360(.dina(n5585),.dinb(w_n221_54[2]),.dout(n5586),.clk(gclk));
	jor g05361(.dina(w_n5452_0[1]),.dinb(n5586),.dout(n5587),.clk(gclk));
	jand g05362(.dina(n5587),.dinb(n5468),.dout(n5588),.clk(gclk));
	jor g05363(.dina(w_n5458_0[0]),.dinb(w_n5588_0[1]),.dout(n5589),.clk(gclk));
	jor g05364(.dina(n5589),.dinb(w_n5105_0[0]),.dout(n5590),.clk(gclk));
	jor g05365(.dina(n5590),.dinb(w_n5467_0[1]),.dout(n5591),.clk(gclk));
	jand g05366(.dina(n5591),.dinb(w_n218_22[2]),.dout(n5592),.clk(gclk));
	jand g05367(.dina(w_n5259_44[1]),.dinb(w_n4906_0[0]),.dout(n5593),.clk(gclk));
	jor g05368(.dina(w_n5593_0[1]),.dinb(w_n5592_0[1]),.dout(n5594),.clk(gclk));
	jor g05369(.dina(n5594),.dinb(w_n5466_0[1]),.dout(n5595),.clk(gclk));
	jor g05370(.dina(n5595),.dinb(w_n5461_0[1]),.dout(asqrt_fa_36),.clk(gclk));
	jnot g05371(.din(w_n5466_0[0]),.dout(n5597),.clk(gclk));
	jnot g05372(.din(w_n5467_0[0]),.dout(n5598),.clk(gclk));
	jand g05373(.dina(w_n5459_0[1]),.dinb(w_n5455_0[1]),.dout(n5599),.clk(gclk));
	jand g05374(.dina(n5599),.dinb(w_n5132_0[1]),.dout(n5600),.clk(gclk));
	jand g05375(.dina(n5600),.dinb(n5598),.dout(n5601),.clk(gclk));
	jor g05376(.dina(n5601),.dinb(w_asqrt63_41[0]),.dout(n5602),.clk(gclk));
	jnot g05377(.din(w_n5593_0[0]),.dout(n5603),.clk(gclk));
	jand g05378(.dina(n5603),.dinb(n5602),.dout(n5604),.clk(gclk));
	jand g05379(.dina(n5604),.dinb(n5597),.dout(n5605),.clk(gclk));
	jand g05380(.dina(w_n5605_0[1]),.dinb(w_n5460_0[0]),.dout(n5606),.clk(gclk));
	jxor g05381(.dina(w_n5447_0[0]),.dinb(w_n221_54[1]),.dout(n5607),.clk(gclk));
	jor g05382(.dina(n5607),.dinb(w_n5606_55[2]),.dout(n5608),.clk(gclk));
	jxor g05383(.dina(n5608),.dinb(w_n5452_0[0]),.dout(n5609),.clk(gclk));
	jnot g05384(.din(w_n5609_0[1]),.dout(n5610),.clk(gclk));
	jor g05385(.dina(w_n5606_55[1]),.dinb(w_n5121_1[0]),.dout(n5611),.clk(gclk));
	jnot g05386(.din(w_a68_0[2]),.dout(n5612),.clk(gclk));
	jnot g05387(.din(w_a69_0[1]),.dout(n5613),.clk(gclk));
	jand g05388(.dina(w_n5613_0[1]),.dinb(w_n5612_1[2]),.dout(n5614),.clk(gclk));
	jand g05389(.dina(w_n5614_0[2]),.dinb(w_n5121_0[2]),.dout(n5615),.clk(gclk));
	jnot g05390(.din(w_n5615_0[1]),.dout(n5616),.clk(gclk));
	jand g05391(.dina(n5616),.dinb(n5611),.dout(n5617),.clk(gclk));
	jor g05392(.dina(w_n5617_0[2]),.dinb(w_n5259_44[0]),.dout(n5618),.clk(gclk));
	jand g05393(.dina(w_n5617_0[1]),.dinb(w_n5259_43[2]),.dout(n5619),.clk(gclk));
	jor g05394(.dina(w_n5606_55[0]),.dinb(w_a70_1[0]),.dout(n5620),.clk(gclk));
	jand g05395(.dina(n5620),.dinb(w_a71_0[0]),.dout(n5621),.clk(gclk));
	jand g05396(.dina(w_asqrt35_27),.dinb(w_n5123_0[1]),.dout(n5622),.clk(gclk));
	jor g05397(.dina(n5622),.dinb(n5621),.dout(n5623),.clk(gclk));
	jor g05398(.dina(n5623),.dinb(n5619),.dout(n5624),.clk(gclk));
	jand g05399(.dina(n5624),.dinb(w_n5618_0[1]),.dout(n5625),.clk(gclk));
	jor g05400(.dina(w_n5625_0[2]),.dinb(w_n4902_48[0]),.dout(n5626),.clk(gclk));
	jand g05401(.dina(w_n5625_0[1]),.dinb(w_n4902_47[2]),.dout(n5627),.clk(gclk));
	jnot g05402(.din(w_n5123_0[0]),.dout(n5628),.clk(gclk));
	jor g05403(.dina(w_n5606_54[2]),.dinb(n5628),.dout(n5629),.clk(gclk));
	jor g05404(.dina(w_n5461_0[0]),.dinb(w_n5259_43[1]),.dout(n5630),.clk(gclk));
	jor g05405(.dina(n5630),.dinb(w_n5465_0[0]),.dout(n5631),.clk(gclk));
	jor g05406(.dina(n5631),.dinb(w_n5592_0[0]),.dout(n5632),.clk(gclk));
	jand g05407(.dina(n5632),.dinb(w_n5629_0[1]),.dout(n5633),.clk(gclk));
	jxor g05408(.dina(n5633),.dinb(w_n4908_0[1]),.dout(n5634),.clk(gclk));
	jor g05409(.dina(w_n5634_0[2]),.dinb(n5627),.dout(n5635),.clk(gclk));
	jand g05410(.dina(n5635),.dinb(w_n5626_0[1]),.dout(n5636),.clk(gclk));
	jor g05411(.dina(w_n5636_0[2]),.dinb(w_n4582_45[0]),.dout(n5637),.clk(gclk));
	jand g05412(.dina(w_n5636_0[1]),.dinb(w_n4582_44[2]),.dout(n5638),.clk(gclk));
	jxor g05413(.dina(w_n5126_0[0]),.dinb(w_n4902_47[1]),.dout(n5639),.clk(gclk));
	jor g05414(.dina(n5639),.dinb(w_n5606_54[1]),.dout(n5640),.clk(gclk));
	jxor g05415(.dina(n5640),.dinb(w_n5500_0[0]),.dout(n5641),.clk(gclk));
	jnot g05416(.din(w_n5641_0[2]),.dout(n5642),.clk(gclk));
	jor g05417(.dina(n5642),.dinb(n5638),.dout(n5643),.clk(gclk));
	jand g05418(.dina(n5643),.dinb(w_n5637_0[1]),.dout(n5644),.clk(gclk));
	jor g05419(.dina(w_n5644_0[2]),.dinb(w_n4249_48[2]),.dout(n5645),.clk(gclk));
	jand g05420(.dina(w_n5644_0[1]),.dinb(w_n4249_48[1]),.dout(n5646),.clk(gclk));
	jxor g05421(.dina(w_n5263_0[0]),.dinb(w_n4582_44[1]),.dout(n5647),.clk(gclk));
	jor g05422(.dina(n5647),.dinb(w_n5606_54[0]),.dout(n5648),.clk(gclk));
	jxor g05423(.dina(n5648),.dinb(w_n5272_0[0]),.dout(n5649),.clk(gclk));
	jor g05424(.dina(w_n5649_0[2]),.dinb(n5646),.dout(n5650),.clk(gclk));
	jand g05425(.dina(n5650),.dinb(w_n5645_0[1]),.dout(n5651),.clk(gclk));
	jor g05426(.dina(w_n5651_0[2]),.dinb(w_n3955_45[2]),.dout(n5652),.clk(gclk));
	jand g05427(.dina(w_n5651_0[1]),.dinb(w_n3955_45[1]),.dout(n5653),.clk(gclk));
	jxor g05428(.dina(w_n5274_0[0]),.dinb(w_n4249_48[0]),.dout(n5654),.clk(gclk));
	jor g05429(.dina(n5654),.dinb(w_n5606_53[2]),.dout(n5655),.clk(gclk));
	jxor g05430(.dina(n5655),.dinb(w_n5507_0[0]),.dout(n5656),.clk(gclk));
	jnot g05431(.din(w_n5656_0[2]),.dout(n5657),.clk(gclk));
	jor g05432(.dina(n5657),.dinb(n5653),.dout(n5658),.clk(gclk));
	jand g05433(.dina(n5658),.dinb(w_n5652_0[1]),.dout(n5659),.clk(gclk));
	jor g05434(.dina(w_n5659_0[2]),.dinb(w_n3642_49[0]),.dout(n5660),.clk(gclk));
	jand g05435(.dina(w_n5659_0[1]),.dinb(w_n3642_48[2]),.dout(n5661),.clk(gclk));
	jxor g05436(.dina(w_n5281_0[0]),.dinb(w_n3955_45[0]),.dout(n5662),.clk(gclk));
	jor g05437(.dina(n5662),.dinb(w_n5606_53[1]),.dout(n5663),.clk(gclk));
	jxor g05438(.dina(n5663),.dinb(w_n5287_0[0]),.dout(n5664),.clk(gclk));
	jor g05439(.dina(w_n5664_0[2]),.dinb(n5661),.dout(n5665),.clk(gclk));
	jand g05440(.dina(n5665),.dinb(w_n5660_0[1]),.dout(n5666),.clk(gclk));
	jor g05441(.dina(w_n5666_0[2]),.dinb(w_n3368_46[1]),.dout(n5667),.clk(gclk));
	jand g05442(.dina(w_n5666_0[1]),.dinb(w_n3368_46[0]),.dout(n5668),.clk(gclk));
	jxor g05443(.dina(w_n5289_0[0]),.dinb(w_n3642_48[1]),.dout(n5669),.clk(gclk));
	jor g05444(.dina(n5669),.dinb(w_n5606_53[0]),.dout(n5670),.clk(gclk));
	jxor g05445(.dina(n5670),.dinb(w_n5514_0[0]),.dout(n5671),.clk(gclk));
	jnot g05446(.din(w_n5671_0[2]),.dout(n5672),.clk(gclk));
	jor g05447(.dina(n5672),.dinb(n5668),.dout(n5673),.clk(gclk));
	jand g05448(.dina(n5673),.dinb(w_n5667_0[1]),.dout(n5674),.clk(gclk));
	jor g05449(.dina(w_n5674_0[2]),.dinb(w_n3089_49[2]),.dout(n5675),.clk(gclk));
	jand g05450(.dina(w_n5674_0[1]),.dinb(w_n3089_49[1]),.dout(n5676),.clk(gclk));
	jxor g05451(.dina(w_n5296_0[0]),.dinb(w_n3368_45[2]),.dout(n5677),.clk(gclk));
	jor g05452(.dina(n5677),.dinb(w_n5606_52[2]),.dout(n5678),.clk(gclk));
	jxor g05453(.dina(n5678),.dinb(w_n5518_0[0]),.dout(n5679),.clk(gclk));
	jnot g05454(.din(w_n5679_0[2]),.dout(n5680),.clk(gclk));
	jor g05455(.dina(n5680),.dinb(n5676),.dout(n5681),.clk(gclk));
	jand g05456(.dina(n5681),.dinb(w_n5675_0[1]),.dout(n5682),.clk(gclk));
	jor g05457(.dina(w_n5682_0[2]),.dinb(w_n2833_47[1]),.dout(n5683),.clk(gclk));
	jand g05458(.dina(w_n5682_0[1]),.dinb(w_n2833_47[0]),.dout(n5684),.clk(gclk));
	jxor g05459(.dina(w_n5303_0[0]),.dinb(w_n3089_49[0]),.dout(n5685),.clk(gclk));
	jor g05460(.dina(n5685),.dinb(w_n5606_52[1]),.dout(n5686),.clk(gclk));
	jxor g05461(.dina(n5686),.dinb(w_n5522_0[0]),.dout(n5687),.clk(gclk));
	jnot g05462(.din(w_n5687_0[2]),.dout(n5688),.clk(gclk));
	jor g05463(.dina(n5688),.dinb(n5684),.dout(n5689),.clk(gclk));
	jand g05464(.dina(n5689),.dinb(w_n5683_0[1]),.dout(n5690),.clk(gclk));
	jor g05465(.dina(w_n5690_0[2]),.dinb(w_n2572_50[0]),.dout(n5691),.clk(gclk));
	jand g05466(.dina(w_n5690_0[1]),.dinb(w_n2572_49[2]),.dout(n5692),.clk(gclk));
	jxor g05467(.dina(w_n5310_0[0]),.dinb(w_n2833_46[2]),.dout(n5693),.clk(gclk));
	jor g05468(.dina(n5693),.dinb(w_n5606_52[0]),.dout(n5694),.clk(gclk));
	jxor g05469(.dina(n5694),.dinb(w_n5316_0[0]),.dout(n5695),.clk(gclk));
	jor g05470(.dina(w_n5695_0[2]),.dinb(n5692),.dout(n5696),.clk(gclk));
	jand g05471(.dina(n5696),.dinb(w_n5691_0[1]),.dout(n5697),.clk(gclk));
	jor g05472(.dina(w_n5697_0[2]),.dinb(w_n2345_48[0]),.dout(n5698),.clk(gclk));
	jand g05473(.dina(w_n5697_0[1]),.dinb(w_n2345_47[2]),.dout(n5699),.clk(gclk));
	jxor g05474(.dina(w_n5318_0[0]),.dinb(w_n2572_49[1]),.dout(n5700),.clk(gclk));
	jor g05475(.dina(n5700),.dinb(w_n5606_51[2]),.dout(n5701),.clk(gclk));
	jxor g05476(.dina(n5701),.dinb(w_n5324_0[0]),.dout(n5702),.clk(gclk));
	jor g05477(.dina(w_n5702_0[2]),.dinb(n5699),.dout(n5703),.clk(gclk));
	jand g05478(.dina(n5703),.dinb(w_n5698_0[1]),.dout(n5704),.clk(gclk));
	jor g05479(.dina(w_n5704_0[2]),.dinb(w_n2108_50[2]),.dout(n5705),.clk(gclk));
	jand g05480(.dina(w_n5704_0[1]),.dinb(w_n2108_50[1]),.dout(n5706),.clk(gclk));
	jxor g05481(.dina(w_n5326_0[0]),.dinb(w_n2345_47[1]),.dout(n5707),.clk(gclk));
	jor g05482(.dina(n5707),.dinb(w_n5606_51[1]),.dout(n5708),.clk(gclk));
	jxor g05483(.dina(n5708),.dinb(w_n5332_0[0]),.dout(n5709),.clk(gclk));
	jor g05484(.dina(w_n5709_0[2]),.dinb(n5706),.dout(n5710),.clk(gclk));
	jand g05485(.dina(n5710),.dinb(w_n5705_0[1]),.dout(n5711),.clk(gclk));
	jor g05486(.dina(w_n5711_0[2]),.dinb(w_n1912_49[0]),.dout(n5712),.clk(gclk));
	jand g05487(.dina(w_n5711_0[1]),.dinb(w_n1912_48[2]),.dout(n5713),.clk(gclk));
	jxor g05488(.dina(w_n5334_0[0]),.dinb(w_n2108_50[0]),.dout(n5714),.clk(gclk));
	jor g05489(.dina(n5714),.dinb(w_n5606_51[0]),.dout(n5715),.clk(gclk));
	jxor g05490(.dina(n5715),.dinb(w_n5535_0[0]),.dout(n5716),.clk(gclk));
	jnot g05491(.din(w_n5716_0[2]),.dout(n5717),.clk(gclk));
	jor g05492(.dina(n5717),.dinb(n5713),.dout(n5718),.clk(gclk));
	jand g05493(.dina(n5718),.dinb(w_n5712_0[1]),.dout(n5719),.clk(gclk));
	jor g05494(.dina(w_n5719_0[2]),.dinb(w_n1699_51[1]),.dout(n5720),.clk(gclk));
	jand g05495(.dina(w_n5719_0[1]),.dinb(w_n1699_51[0]),.dout(n5721),.clk(gclk));
	jxor g05496(.dina(w_n5341_0[0]),.dinb(w_n1912_48[1]),.dout(n5722),.clk(gclk));
	jor g05497(.dina(n5722),.dinb(w_n5606_50[2]),.dout(n5723),.clk(gclk));
	jxor g05498(.dina(n5723),.dinb(w_n5347_0[0]),.dout(n5724),.clk(gclk));
	jor g05499(.dina(w_n5724_0[2]),.dinb(n5721),.dout(n5725),.clk(gclk));
	jand g05500(.dina(n5725),.dinb(w_n5720_0[1]),.dout(n5726),.clk(gclk));
	jor g05501(.dina(w_n5726_0[2]),.dinb(w_n1516_49[2]),.dout(n5727),.clk(gclk));
	jand g05502(.dina(w_n5726_0[1]),.dinb(w_n1516_49[1]),.dout(n5728),.clk(gclk));
	jxor g05503(.dina(w_n5349_0[0]),.dinb(w_n1699_50[2]),.dout(n5729),.clk(gclk));
	jor g05504(.dina(n5729),.dinb(w_n5606_50[1]),.dout(n5730),.clk(gclk));
	jxor g05505(.dina(n5730),.dinb(w_n5542_0[0]),.dout(n5731),.clk(gclk));
	jnot g05506(.din(w_n5731_0[2]),.dout(n5732),.clk(gclk));
	jor g05507(.dina(n5732),.dinb(n5728),.dout(n5733),.clk(gclk));
	jand g05508(.dina(n5733),.dinb(w_n5727_0[1]),.dout(n5734),.clk(gclk));
	jor g05509(.dina(w_n5734_0[2]),.dinb(w_n1332_51[1]),.dout(n5735),.clk(gclk));
	jand g05510(.dina(w_n5734_0[1]),.dinb(w_n1332_51[0]),.dout(n5736),.clk(gclk));
	jxor g05511(.dina(w_n5356_0[0]),.dinb(w_n1516_49[0]),.dout(n5737),.clk(gclk));
	jor g05512(.dina(n5737),.dinb(w_n5606_50[0]),.dout(n5738),.clk(gclk));
	jxor g05513(.dina(n5738),.dinb(w_n5362_0[0]),.dout(n5739),.clk(gclk));
	jor g05514(.dina(w_n5739_0[2]),.dinb(n5736),.dout(n5740),.clk(gclk));
	jand g05515(.dina(n5740),.dinb(w_n5735_0[1]),.dout(n5741),.clk(gclk));
	jor g05516(.dina(w_n5741_0[2]),.dinb(w_n1173_50[1]),.dout(n5742),.clk(gclk));
	jand g05517(.dina(w_n5741_0[1]),.dinb(w_n1173_50[0]),.dout(n5743),.clk(gclk));
	jxor g05518(.dina(w_n5364_0[0]),.dinb(w_n1332_50[2]),.dout(n5744),.clk(gclk));
	jor g05519(.dina(n5744),.dinb(w_n5606_49[2]),.dout(n5745),.clk(gclk));
	jxor g05520(.dina(n5745),.dinb(w_n5549_0[0]),.dout(n5746),.clk(gclk));
	jnot g05521(.din(w_n5746_0[2]),.dout(n5747),.clk(gclk));
	jor g05522(.dina(n5747),.dinb(n5743),.dout(n5748),.clk(gclk));
	jand g05523(.dina(n5748),.dinb(w_n5742_0[1]),.dout(n5749),.clk(gclk));
	jor g05524(.dina(w_n5749_0[2]),.dinb(w_n1008_52[1]),.dout(n5750),.clk(gclk));
	jand g05525(.dina(w_n5749_0[1]),.dinb(w_n1008_52[0]),.dout(n5751),.clk(gclk));
	jxor g05526(.dina(w_n5371_0[0]),.dinb(w_n1173_49[2]),.dout(n5752),.clk(gclk));
	jor g05527(.dina(n5752),.dinb(w_n5606_49[1]),.dout(n5753),.clk(gclk));
	jxor g05528(.dina(n5753),.dinb(w_n5553_0[0]),.dout(n5754),.clk(gclk));
	jnot g05529(.din(w_n5754_0[2]),.dout(n5755),.clk(gclk));
	jor g05530(.dina(n5755),.dinb(n5751),.dout(n5756),.clk(gclk));
	jand g05531(.dina(n5756),.dinb(w_n5750_0[1]),.dout(n5757),.clk(gclk));
	jor g05532(.dina(w_n5757_0[2]),.dinb(w_n884_51[1]),.dout(n5758),.clk(gclk));
	jand g05533(.dina(w_n5757_0[1]),.dinb(w_n884_51[0]),.dout(n5759),.clk(gclk));
	jxor g05534(.dina(w_n5378_0[0]),.dinb(w_n1008_51[2]),.dout(n5760),.clk(gclk));
	jor g05535(.dina(n5760),.dinb(w_n5606_49[0]),.dout(n5761),.clk(gclk));
	jxor g05536(.dina(n5761),.dinb(w_n5384_0[0]),.dout(n5762),.clk(gclk));
	jor g05537(.dina(w_n5762_0[2]),.dinb(n5759),.dout(n5763),.clk(gclk));
	jand g05538(.dina(n5763),.dinb(w_n5758_0[1]),.dout(n5764),.clk(gclk));
	jor g05539(.dina(w_n5764_0[2]),.dinb(w_n743_52[1]),.dout(n5765),.clk(gclk));
	jand g05540(.dina(w_n5764_0[1]),.dinb(w_n743_52[0]),.dout(n5766),.clk(gclk));
	jxor g05541(.dina(w_n5386_0[0]),.dinb(w_n884_50[2]),.dout(n5767),.clk(gclk));
	jor g05542(.dina(n5767),.dinb(w_n5606_48[2]),.dout(n5768),.clk(gclk));
	jxor g05543(.dina(n5768),.dinb(w_n5392_0[0]),.dout(n5769),.clk(gclk));
	jor g05544(.dina(w_n5769_0[2]),.dinb(n5766),.dout(n5770),.clk(gclk));
	jand g05545(.dina(n5770),.dinb(w_n5765_0[1]),.dout(n5771),.clk(gclk));
	jor g05546(.dina(w_n5771_0[2]),.dinb(w_n635_52[1]),.dout(n5772),.clk(gclk));
	jand g05547(.dina(w_n5771_0[1]),.dinb(w_n635_52[0]),.dout(n5773),.clk(gclk));
	jxor g05548(.dina(w_n5394_0[0]),.dinb(w_n743_51[2]),.dout(n5774),.clk(gclk));
	jor g05549(.dina(n5774),.dinb(w_n5606_48[1]),.dout(n5775),.clk(gclk));
	jxor g05550(.dina(n5775),.dinb(w_n5563_0[0]),.dout(n5776),.clk(gclk));
	jnot g05551(.din(w_n5776_0[2]),.dout(n5777),.clk(gclk));
	jor g05552(.dina(n5777),.dinb(n5773),.dout(n5778),.clk(gclk));
	jand g05553(.dina(n5778),.dinb(w_n5772_0[1]),.dout(n5779),.clk(gclk));
	jor g05554(.dina(w_n5779_0[2]),.dinb(w_n515_53[1]),.dout(n5780),.clk(gclk));
	jand g05555(.dina(w_n5779_0[1]),.dinb(w_n515_53[0]),.dout(n5781),.clk(gclk));
	jxor g05556(.dina(w_n5401_0[0]),.dinb(w_n635_51[2]),.dout(n5782),.clk(gclk));
	jor g05557(.dina(n5782),.dinb(w_n5606_48[0]),.dout(n5783),.clk(gclk));
	jxor g05558(.dina(n5783),.dinb(w_n5407_0[0]),.dout(n5784),.clk(gclk));
	jor g05559(.dina(w_n5784_0[2]),.dinb(n5781),.dout(n5785),.clk(gclk));
	jand g05560(.dina(n5785),.dinb(w_n5780_0[1]),.dout(n5786),.clk(gclk));
	jor g05561(.dina(w_n5786_0[2]),.dinb(w_n443_53[1]),.dout(n5787),.clk(gclk));
	jand g05562(.dina(w_n5786_0[1]),.dinb(w_n443_53[0]),.dout(n5788),.clk(gclk));
	jxor g05563(.dina(w_n5409_0[0]),.dinb(w_n515_52[2]),.dout(n5789),.clk(gclk));
	jor g05564(.dina(n5789),.dinb(w_n5606_47[2]),.dout(n5790),.clk(gclk));
	jxor g05565(.dina(n5790),.dinb(w_n5570_0[0]),.dout(n5791),.clk(gclk));
	jnot g05566(.din(w_n5791_0[2]),.dout(n5792),.clk(gclk));
	jor g05567(.dina(n5792),.dinb(n5788),.dout(n5793),.clk(gclk));
	jand g05568(.dina(n5793),.dinb(w_n5787_0[1]),.dout(n5794),.clk(gclk));
	jor g05569(.dina(w_n5794_0[2]),.dinb(w_n352_53[2]),.dout(n5795),.clk(gclk));
	jand g05570(.dina(w_n5794_0[1]),.dinb(w_n352_53[1]),.dout(n5796),.clk(gclk));
	jxor g05571(.dina(w_n5416_0[0]),.dinb(w_n443_52[2]),.dout(n5797),.clk(gclk));
	jor g05572(.dina(n5797),.dinb(w_n5606_47[1]),.dout(n5798),.clk(gclk));
	jxor g05573(.dina(n5798),.dinb(w_n5422_0[0]),.dout(n5799),.clk(gclk));
	jor g05574(.dina(w_n5799_0[2]),.dinb(n5796),.dout(n5800),.clk(gclk));
	jand g05575(.dina(n5800),.dinb(w_n5795_0[1]),.dout(n5801),.clk(gclk));
	jor g05576(.dina(w_n5801_0[2]),.dinb(w_n294_54[0]),.dout(n5802),.clk(gclk));
	jand g05577(.dina(w_n5801_0[1]),.dinb(w_n294_53[2]),.dout(n5803),.clk(gclk));
	jxor g05578(.dina(w_n5424_0[0]),.dinb(w_n352_53[0]),.dout(n5804),.clk(gclk));
	jor g05579(.dina(n5804),.dinb(w_n5606_47[0]),.dout(n5805),.clk(gclk));
	jxor g05580(.dina(n5805),.dinb(w_n5430_0[0]),.dout(n5806),.clk(gclk));
	jor g05581(.dina(w_n5806_0[2]),.dinb(n5803),.dout(n5807),.clk(gclk));
	jand g05582(.dina(n5807),.dinb(w_n5802_0[1]),.dout(n5808),.clk(gclk));
	jor g05583(.dina(w_n5808_0[2]),.dinb(w_n239_54[0]),.dout(n5809),.clk(gclk));
	jand g05584(.dina(w_n5808_0[1]),.dinb(w_n239_53[2]),.dout(n5810),.clk(gclk));
	jxor g05585(.dina(w_n5432_0[0]),.dinb(w_n294_53[1]),.dout(n5811),.clk(gclk));
	jor g05586(.dina(n5811),.dinb(w_n5606_46[2]),.dout(n5812),.clk(gclk));
	jxor g05587(.dina(n5812),.dinb(w_n5438_0[0]),.dout(n5813),.clk(gclk));
	jor g05588(.dina(w_n5813_0[2]),.dinb(n5810),.dout(n5814),.clk(gclk));
	jand g05589(.dina(n5814),.dinb(w_n5809_0[1]),.dout(n5815),.clk(gclk));
	jor g05590(.dina(w_n5815_0[2]),.dinb(w_n221_54[0]),.dout(n5816),.clk(gclk));
	jand g05591(.dina(w_n5815_0[1]),.dinb(w_n221_53[2]),.dout(n5817),.clk(gclk));
	jxor g05592(.dina(w_n5440_0[0]),.dinb(w_n239_53[1]),.dout(n5818),.clk(gclk));
	jor g05593(.dina(n5818),.dinb(w_n5606_46[1]),.dout(n5819),.clk(gclk));
	jxor g05594(.dina(n5819),.dinb(w_n5583_0[0]),.dout(n5820),.clk(gclk));
	jnot g05595(.din(w_n5820_0[2]),.dout(n5821),.clk(gclk));
	jor g05596(.dina(n5821),.dinb(n5817),.dout(n5822),.clk(gclk));
	jand g05597(.dina(n5822),.dinb(w_n5816_0[1]),.dout(n5823),.clk(gclk));
	jand g05598(.dina(w_n5823_1[1]),.dinb(w_n5610_0[2]),.dout(n5824),.clk(gclk));
	jor g05599(.dina(w_n5823_1[0]),.dinb(w_n5610_0[1]),.dout(n5826),.clk(gclk));
	jxor g05600(.dina(w_n5459_0[0]),.dinb(w_n5455_0[0]),.dout(n5827),.clk(gclk));
	jnot g05601(.din(w_n5827_0[1]),.dout(n5828),.clk(gclk));
	jand g05602(.dina(n5828),.dinb(w_asqrt35_26[2]),.dout(n5829),.clk(gclk));
	jor g05603(.dina(w_n5829_0[1]),.dinb(n5826),.dout(n5830),.clk(gclk));
	jand g05604(.dina(n5830),.dinb(w_n218_22[1]),.dout(n5831),.clk(gclk));
	jand g05605(.dina(w_n5605_0[0]),.dinb(w_n5588_0[0]),.dout(n5832),.clk(gclk));
	jand g05606(.dina(w_n5827_0[0]),.dinb(w_asqrt63_40[2]),.dout(n5833),.clk(gclk));
	jnot g05607(.din(n5833),.dout(n5834),.clk(gclk));
	jor g05608(.dina(w_n5834_0[1]),.dinb(n5832),.dout(n5835),.clk(gclk));
	jnot g05609(.din(w_n5835_0[1]),.dout(n5836),.clk(gclk));
	jor g05610(.dina(n5836),.dinb(n5831),.dout(n5837),.clk(gclk));
	jor g05611(.dina(n5837),.dinb(w_n5824_0[1]),.dout(asqrt_fa_35),.clk(gclk));
	jxor g05612(.dina(w_n5815_0[0]),.dinb(w_n221_53[1]),.dout(n5840),.clk(gclk));
	jand g05613(.dina(n5840),.dinb(w_asqrt34_39),.dout(n5841),.clk(gclk));
	jxor g05614(.dina(n5841),.dinb(w_n5820_0[1]),.dout(n5842),.clk(gclk));
	jnot g05615(.din(w_a66_1[1]),.dout(n5843),.clk(gclk));
	jnot g05616(.din(w_a67_0[1]),.dout(n5844),.clk(gclk));
	jand g05617(.dina(w_n5844_0[1]),.dinb(w_n5843_1[1]),.dout(n5845),.clk(gclk));
	jand g05618(.dina(w_n5845_0[2]),.dinb(w_n5612_1[1]),.dout(n5846),.clk(gclk));
	jand g05619(.dina(w_asqrt34_38[2]),.dinb(w_a68_0[1]),.dout(n5847),.clk(gclk));
	jor g05620(.dina(n5847),.dinb(w_n5846_0[1]),.dout(n5848),.clk(gclk));
	jand g05621(.dina(w_n5848_0[2]),.dinb(w_asqrt35_26[1]),.dout(n5849),.clk(gclk));
	jor g05622(.dina(w_n5848_0[1]),.dinb(w_asqrt35_26[0]),.dout(n5850),.clk(gclk));
	jand g05623(.dina(w_asqrt34_38[1]),.dinb(w_n5612_1[0]),.dout(n5851),.clk(gclk));
	jor g05624(.dina(n5851),.dinb(w_n5613_0[0]),.dout(n5852),.clk(gclk));
	jnot g05625(.din(w_n5614_0[1]),.dout(n5853),.clk(gclk));
	jnot g05626(.din(w_n5824_0[0]),.dout(n5854),.clk(gclk));
	jnot g05627(.din(w_n5816_0[0]),.dout(n5856),.clk(gclk));
	jnot g05628(.din(w_n5809_0[0]),.dout(n5857),.clk(gclk));
	jnot g05629(.din(w_n5802_0[0]),.dout(n5858),.clk(gclk));
	jnot g05630(.din(w_n5795_0[0]),.dout(n5859),.clk(gclk));
	jnot g05631(.din(w_n5787_0[0]),.dout(n5860),.clk(gclk));
	jnot g05632(.din(w_n5780_0[0]),.dout(n5861),.clk(gclk));
	jnot g05633(.din(w_n5772_0[0]),.dout(n5862),.clk(gclk));
	jnot g05634(.din(w_n5765_0[0]),.dout(n5863),.clk(gclk));
	jnot g05635(.din(w_n5758_0[0]),.dout(n5864),.clk(gclk));
	jnot g05636(.din(w_n5750_0[0]),.dout(n5865),.clk(gclk));
	jnot g05637(.din(w_n5742_0[0]),.dout(n5866),.clk(gclk));
	jnot g05638(.din(w_n5735_0[0]),.dout(n5867),.clk(gclk));
	jnot g05639(.din(w_n5727_0[0]),.dout(n5868),.clk(gclk));
	jnot g05640(.din(w_n5720_0[0]),.dout(n5869),.clk(gclk));
	jnot g05641(.din(w_n5712_0[0]),.dout(n5870),.clk(gclk));
	jnot g05642(.din(w_n5705_0[0]),.dout(n5871),.clk(gclk));
	jnot g05643(.din(w_n5698_0[0]),.dout(n5872),.clk(gclk));
	jnot g05644(.din(w_n5691_0[0]),.dout(n5873),.clk(gclk));
	jnot g05645(.din(w_n5683_0[0]),.dout(n5874),.clk(gclk));
	jnot g05646(.din(w_n5675_0[0]),.dout(n5875),.clk(gclk));
	jnot g05647(.din(w_n5667_0[0]),.dout(n5876),.clk(gclk));
	jnot g05648(.din(w_n5660_0[0]),.dout(n5877),.clk(gclk));
	jnot g05649(.din(w_n5652_0[0]),.dout(n5878),.clk(gclk));
	jnot g05650(.din(w_n5645_0[0]),.dout(n5879),.clk(gclk));
	jnot g05651(.din(w_n5637_0[0]),.dout(n5880),.clk(gclk));
	jnot g05652(.din(w_n5626_0[0]),.dout(n5881),.clk(gclk));
	jnot g05653(.din(w_n5618_0[0]),.dout(n5882),.clk(gclk));
	jand g05654(.dina(w_asqrt35_25[2]),.dinb(w_a70_0[2]),.dout(n5883),.clk(gclk));
	jor g05655(.dina(w_n5615_0[0]),.dinb(n5883),.dout(n5884),.clk(gclk));
	jor g05656(.dina(n5884),.dinb(w_asqrt36_29[2]),.dout(n5885),.clk(gclk));
	jand g05657(.dina(w_asqrt35_25[1]),.dinb(w_n5121_0[1]),.dout(n5886),.clk(gclk));
	jor g05658(.dina(n5886),.dinb(w_n5122_0[0]),.dout(n5887),.clk(gclk));
	jand g05659(.dina(w_n5629_0[0]),.dinb(n5887),.dout(n5888),.clk(gclk));
	jand g05660(.dina(w_n5888_0[1]),.dinb(n5885),.dout(n5889),.clk(gclk));
	jor g05661(.dina(n5889),.dinb(n5882),.dout(n5890),.clk(gclk));
	jor g05662(.dina(n5890),.dinb(w_asqrt37_26[0]),.dout(n5891),.clk(gclk));
	jnot g05663(.din(w_n5634_0[1]),.dout(n5892),.clk(gclk));
	jand g05664(.dina(n5892),.dinb(n5891),.dout(n5893),.clk(gclk));
	jor g05665(.dina(n5893),.dinb(n5881),.dout(n5894),.clk(gclk));
	jor g05666(.dina(n5894),.dinb(w_asqrt38_30[0]),.dout(n5895),.clk(gclk));
	jand g05667(.dina(w_n5641_0[1]),.dinb(n5895),.dout(n5896),.clk(gclk));
	jor g05668(.dina(n5896),.dinb(n5880),.dout(n5897),.clk(gclk));
	jor g05669(.dina(n5897),.dinb(w_asqrt39_26[2]),.dout(n5898),.clk(gclk));
	jnot g05670(.din(w_n5649_0[1]),.dout(n5899),.clk(gclk));
	jand g05671(.dina(n5899),.dinb(n5898),.dout(n5900),.clk(gclk));
	jor g05672(.dina(n5900),.dinb(n5879),.dout(n5901),.clk(gclk));
	jor g05673(.dina(n5901),.dinb(w_asqrt40_30[0]),.dout(n5902),.clk(gclk));
	jand g05674(.dina(w_n5656_0[1]),.dinb(n5902),.dout(n5903),.clk(gclk));
	jor g05675(.dina(n5903),.dinb(n5878),.dout(n5904),.clk(gclk));
	jor g05676(.dina(n5904),.dinb(w_asqrt41_27[0]),.dout(n5905),.clk(gclk));
	jnot g05677(.din(w_n5664_0[1]),.dout(n5906),.clk(gclk));
	jand g05678(.dina(n5906),.dinb(n5905),.dout(n5907),.clk(gclk));
	jor g05679(.dina(n5907),.dinb(n5877),.dout(n5908),.clk(gclk));
	jor g05680(.dina(n5908),.dinb(w_asqrt42_30[1]),.dout(n5909),.clk(gclk));
	jand g05681(.dina(w_n5671_0[1]),.dinb(n5909),.dout(n5910),.clk(gclk));
	jor g05682(.dina(n5910),.dinb(n5876),.dout(n5911),.clk(gclk));
	jor g05683(.dina(n5911),.dinb(w_asqrt43_27[1]),.dout(n5912),.clk(gclk));
	jand g05684(.dina(w_n5679_0[1]),.dinb(n5912),.dout(n5913),.clk(gclk));
	jor g05685(.dina(n5913),.dinb(n5875),.dout(n5914),.clk(gclk));
	jor g05686(.dina(n5914),.dinb(w_asqrt44_30[1]),.dout(n5915),.clk(gclk));
	jand g05687(.dina(w_n5687_0[1]),.dinb(n5915),.dout(n5916),.clk(gclk));
	jor g05688(.dina(n5916),.dinb(n5874),.dout(n5917),.clk(gclk));
	jor g05689(.dina(n5917),.dinb(w_asqrt45_28[0]),.dout(n5918),.clk(gclk));
	jnot g05690(.din(w_n5695_0[1]),.dout(n5919),.clk(gclk));
	jand g05691(.dina(n5919),.dinb(n5918),.dout(n5920),.clk(gclk));
	jor g05692(.dina(n5920),.dinb(n5873),.dout(n5921),.clk(gclk));
	jor g05693(.dina(n5921),.dinb(w_asqrt46_30[1]),.dout(n5922),.clk(gclk));
	jnot g05694(.din(w_n5702_0[1]),.dout(n5923),.clk(gclk));
	jand g05695(.dina(n5923),.dinb(n5922),.dout(n5924),.clk(gclk));
	jor g05696(.dina(n5924),.dinb(n5872),.dout(n5925),.clk(gclk));
	jor g05697(.dina(n5925),.dinb(w_asqrt47_28[2]),.dout(n5926),.clk(gclk));
	jnot g05698(.din(w_n5709_0[1]),.dout(n5927),.clk(gclk));
	jand g05699(.dina(n5927),.dinb(n5926),.dout(n5928),.clk(gclk));
	jor g05700(.dina(n5928),.dinb(n5871),.dout(n5929),.clk(gclk));
	jor g05701(.dina(n5929),.dinb(w_asqrt48_30[2]),.dout(n5930),.clk(gclk));
	jand g05702(.dina(w_n5716_0[1]),.dinb(n5930),.dout(n5931),.clk(gclk));
	jor g05703(.dina(n5931),.dinb(n5870),.dout(n5932),.clk(gclk));
	jor g05704(.dina(n5932),.dinb(w_asqrt49_29[0]),.dout(n5933),.clk(gclk));
	jnot g05705(.din(w_n5724_0[1]),.dout(n5934),.clk(gclk));
	jand g05706(.dina(n5934),.dinb(n5933),.dout(n5935),.clk(gclk));
	jor g05707(.dina(n5935),.dinb(n5869),.dout(n5936),.clk(gclk));
	jor g05708(.dina(n5936),.dinb(w_asqrt50_31[0]),.dout(n5937),.clk(gclk));
	jand g05709(.dina(w_n5731_0[1]),.dinb(n5937),.dout(n5938),.clk(gclk));
	jor g05710(.dina(n5938),.dinb(n5868),.dout(n5939),.clk(gclk));
	jor g05711(.dina(n5939),.dinb(w_asqrt51_29[1]),.dout(n5940),.clk(gclk));
	jnot g05712(.din(w_n5739_0[1]),.dout(n5941),.clk(gclk));
	jand g05713(.dina(n5941),.dinb(n5940),.dout(n5942),.clk(gclk));
	jor g05714(.dina(n5942),.dinb(n5867),.dout(n5943),.clk(gclk));
	jor g05715(.dina(n5943),.dinb(w_asqrt52_31[0]),.dout(n5944),.clk(gclk));
	jand g05716(.dina(w_n5746_0[1]),.dinb(n5944),.dout(n5945),.clk(gclk));
	jor g05717(.dina(n5945),.dinb(n5866),.dout(n5946),.clk(gclk));
	jor g05718(.dina(n5946),.dinb(w_asqrt53_30[0]),.dout(n5947),.clk(gclk));
	jand g05719(.dina(w_n5754_0[1]),.dinb(n5947),.dout(n5948),.clk(gclk));
	jor g05720(.dina(n5948),.dinb(n5865),.dout(n5949),.clk(gclk));
	jor g05721(.dina(n5949),.dinb(w_asqrt54_31[0]),.dout(n5950),.clk(gclk));
	jnot g05722(.din(w_n5762_0[1]),.dout(n5951),.clk(gclk));
	jand g05723(.dina(n5951),.dinb(n5950),.dout(n5952),.clk(gclk));
	jor g05724(.dina(n5952),.dinb(n5864),.dout(n5953),.clk(gclk));
	jor g05725(.dina(n5953),.dinb(w_asqrt55_30[1]),.dout(n5954),.clk(gclk));
	jnot g05726(.din(w_n5769_0[1]),.dout(n5955),.clk(gclk));
	jand g05727(.dina(n5955),.dinb(n5954),.dout(n5956),.clk(gclk));
	jor g05728(.dina(n5956),.dinb(n5863),.dout(n5957),.clk(gclk));
	jor g05729(.dina(n5957),.dinb(w_asqrt56_31[1]),.dout(n5958),.clk(gclk));
	jand g05730(.dina(w_n5776_0[1]),.dinb(n5958),.dout(n5959),.clk(gclk));
	jor g05731(.dina(n5959),.dinb(n5862),.dout(n5960),.clk(gclk));
	jor g05732(.dina(n5960),.dinb(w_asqrt57_31[0]),.dout(n5961),.clk(gclk));
	jnot g05733(.din(w_n5784_0[1]),.dout(n5962),.clk(gclk));
	jand g05734(.dina(n5962),.dinb(n5961),.dout(n5963),.clk(gclk));
	jor g05735(.dina(n5963),.dinb(n5861),.dout(n5964),.clk(gclk));
	jor g05736(.dina(n5964),.dinb(w_asqrt58_31[2]),.dout(n5965),.clk(gclk));
	jand g05737(.dina(w_n5791_0[1]),.dinb(n5965),.dout(n5966),.clk(gclk));
	jor g05738(.dina(n5966),.dinb(n5860),.dout(n5967),.clk(gclk));
	jor g05739(.dina(n5967),.dinb(w_asqrt59_31[1]),.dout(n5968),.clk(gclk));
	jnot g05740(.din(w_n5799_0[1]),.dout(n5969),.clk(gclk));
	jand g05741(.dina(n5969),.dinb(n5968),.dout(n5970),.clk(gclk));
	jor g05742(.dina(n5970),.dinb(n5859),.dout(n5971),.clk(gclk));
	jor g05743(.dina(n5971),.dinb(w_asqrt60_31[2]),.dout(n5972),.clk(gclk));
	jnot g05744(.din(w_n5806_0[1]),.dout(n5973),.clk(gclk));
	jand g05745(.dina(n5973),.dinb(n5972),.dout(n5974),.clk(gclk));
	jor g05746(.dina(n5974),.dinb(n5858),.dout(n5975),.clk(gclk));
	jor g05747(.dina(n5975),.dinb(w_asqrt61_31[2]),.dout(n5976),.clk(gclk));
	jnot g05748(.din(w_n5813_0[1]),.dout(n5977),.clk(gclk));
	jand g05749(.dina(n5977),.dinb(n5976),.dout(n5978),.clk(gclk));
	jor g05750(.dina(n5978),.dinb(n5857),.dout(n5979),.clk(gclk));
	jor g05751(.dina(n5979),.dinb(w_asqrt62_31[2]),.dout(n5980),.clk(gclk));
	jand g05752(.dina(w_n5820_0[0]),.dinb(n5980),.dout(n5981),.clk(gclk));
	jor g05753(.dina(n5981),.dinb(n5856),.dout(n5982),.clk(gclk));
	jand g05754(.dina(n5982),.dinb(w_n5609_0[0]),.dout(n5983),.clk(gclk));
	jnot g05755(.din(w_n5829_0[0]),.dout(n5984),.clk(gclk));
	jand g05756(.dina(n5984),.dinb(n5983),.dout(n5985),.clk(gclk));
	jor g05757(.dina(n5985),.dinb(w_asqrt63_40[1]),.dout(n5986),.clk(gclk));
	jand g05758(.dina(w_n5835_0[0]),.dinb(w_n5986_0[1]),.dout(n5987),.clk(gclk));
	jand g05759(.dina(w_n5987_0[1]),.dinb(w_n5854_0[1]),.dout(n5989),.clk(gclk));
	jor g05760(.dina(w_n5989_42[1]),.dinb(n5853),.dout(n5990),.clk(gclk));
	jand g05761(.dina(n5990),.dinb(n5852),.dout(n5991),.clk(gclk));
	jand g05762(.dina(n5991),.dinb(n5850),.dout(n5992),.clk(gclk));
	jor g05763(.dina(n5992),.dinb(w_n5849_0[1]),.dout(n5993),.clk(gclk));
	jand g05764(.dina(w_n5993_0[2]),.dinb(w_asqrt36_29[1]),.dout(n5994),.clk(gclk));
	jor g05765(.dina(w_n5993_0[1]),.dinb(w_asqrt36_29[0]),.dout(n5995),.clk(gclk));
	jand g05766(.dina(w_asqrt34_38[0]),.dinb(w_n5614_0[0]),.dout(n5996),.clk(gclk));
	jand g05767(.dina(w_n5986_0[0]),.dinb(w_asqrt35_25[0]),.dout(n5997),.clk(gclk));
	jand g05768(.dina(n5997),.dinb(w_n5834_0[0]),.dout(n5998),.clk(gclk));
	jand g05769(.dina(n5998),.dinb(w_n5854_0[0]),.dout(n5999),.clk(gclk));
	jor g05770(.dina(n5999),.dinb(w_n5996_0[1]),.dout(n6000),.clk(gclk));
	jxor g05771(.dina(n6000),.dinb(w_a70_0[1]),.dout(n6001),.clk(gclk));
	jnot g05772(.din(w_n6001_0[1]),.dout(n6002),.clk(gclk));
	jand g05773(.dina(w_n6002_0[1]),.dinb(n5995),.dout(n6003),.clk(gclk));
	jor g05774(.dina(n6003),.dinb(w_n5994_0[1]),.dout(n6004),.clk(gclk));
	jand g05775(.dina(w_n6004_0[2]),.dinb(w_asqrt37_25[2]),.dout(n6005),.clk(gclk));
	jor g05776(.dina(w_n6004_0[1]),.dinb(w_asqrt37_25[1]),.dout(n6006),.clk(gclk));
	jxor g05777(.dina(w_n5617_0[0]),.dinb(w_n5259_43[0]),.dout(n6007),.clk(gclk));
	jand g05778(.dina(n6007),.dinb(w_asqrt34_37[2]),.dout(n6008),.clk(gclk));
	jxor g05779(.dina(n6008),.dinb(w_n5888_0[0]),.dout(n6009),.clk(gclk));
	jand g05780(.dina(w_n6009_0[1]),.dinb(n6006),.dout(n6010),.clk(gclk));
	jor g05781(.dina(n6010),.dinb(w_n6005_0[1]),.dout(n6011),.clk(gclk));
	jand g05782(.dina(w_n6011_0[2]),.dinb(w_asqrt38_29[2]),.dout(n6012),.clk(gclk));
	jor g05783(.dina(w_n6011_0[1]),.dinb(w_asqrt38_29[1]),.dout(n6013),.clk(gclk));
	jxor g05784(.dina(w_n5625_0[0]),.dinb(w_n4902_47[0]),.dout(n6014),.clk(gclk));
	jand g05785(.dina(n6014),.dinb(w_asqrt34_37[1]),.dout(n6015),.clk(gclk));
	jxor g05786(.dina(n6015),.dinb(w_n5634_0[0]),.dout(n6016),.clk(gclk));
	jnot g05787(.din(w_n6016_0[1]),.dout(n6017),.clk(gclk));
	jand g05788(.dina(w_n6017_0[1]),.dinb(n6013),.dout(n6018),.clk(gclk));
	jor g05789(.dina(n6018),.dinb(w_n6012_0[1]),.dout(n6019),.clk(gclk));
	jand g05790(.dina(w_n6019_0[2]),.dinb(w_asqrt39_26[1]),.dout(n6020),.clk(gclk));
	jor g05791(.dina(w_n6019_0[1]),.dinb(w_asqrt39_26[0]),.dout(n6021),.clk(gclk));
	jxor g05792(.dina(w_n5636_0[0]),.dinb(w_n4582_44[0]),.dout(n6022),.clk(gclk));
	jand g05793(.dina(n6022),.dinb(w_asqrt34_37[0]),.dout(n6023),.clk(gclk));
	jxor g05794(.dina(n6023),.dinb(w_n5641_0[0]),.dout(n6024),.clk(gclk));
	jand g05795(.dina(w_n6024_0[1]),.dinb(n6021),.dout(n6025),.clk(gclk));
	jor g05796(.dina(n6025),.dinb(w_n6020_0[1]),.dout(n6026),.clk(gclk));
	jand g05797(.dina(w_n6026_0[2]),.dinb(w_asqrt40_29[2]),.dout(n6027),.clk(gclk));
	jor g05798(.dina(w_n6026_0[1]),.dinb(w_asqrt40_29[1]),.dout(n6028),.clk(gclk));
	jxor g05799(.dina(w_n5644_0[0]),.dinb(w_n4249_47[2]),.dout(n6029),.clk(gclk));
	jand g05800(.dina(n6029),.dinb(w_asqrt34_36[2]),.dout(n6030),.clk(gclk));
	jxor g05801(.dina(n6030),.dinb(w_n5649_0[0]),.dout(n6031),.clk(gclk));
	jnot g05802(.din(w_n6031_0[1]),.dout(n6032),.clk(gclk));
	jand g05803(.dina(w_n6032_0[1]),.dinb(n6028),.dout(n6033),.clk(gclk));
	jor g05804(.dina(n6033),.dinb(w_n6027_0[1]),.dout(n6034),.clk(gclk));
	jand g05805(.dina(w_n6034_0[2]),.dinb(w_asqrt41_26[2]),.dout(n6035),.clk(gclk));
	jor g05806(.dina(w_n6034_0[1]),.dinb(w_asqrt41_26[1]),.dout(n6036),.clk(gclk));
	jxor g05807(.dina(w_n5651_0[0]),.dinb(w_n3955_44[2]),.dout(n6037),.clk(gclk));
	jand g05808(.dina(n6037),.dinb(w_asqrt34_36[1]),.dout(n6038),.clk(gclk));
	jxor g05809(.dina(n6038),.dinb(w_n5656_0[0]),.dout(n6039),.clk(gclk));
	jand g05810(.dina(w_n6039_0[1]),.dinb(n6036),.dout(n6040),.clk(gclk));
	jor g05811(.dina(n6040),.dinb(w_n6035_0[1]),.dout(n6041),.clk(gclk));
	jand g05812(.dina(w_n6041_0[2]),.dinb(w_asqrt42_30[0]),.dout(n6042),.clk(gclk));
	jor g05813(.dina(w_n6041_0[1]),.dinb(w_asqrt42_29[2]),.dout(n6043),.clk(gclk));
	jxor g05814(.dina(w_n5659_0[0]),.dinb(w_n3642_48[0]),.dout(n6044),.clk(gclk));
	jand g05815(.dina(n6044),.dinb(w_asqrt34_36[0]),.dout(n6045),.clk(gclk));
	jxor g05816(.dina(n6045),.dinb(w_n5664_0[0]),.dout(n6046),.clk(gclk));
	jnot g05817(.din(w_n6046_0[1]),.dout(n6047),.clk(gclk));
	jand g05818(.dina(w_n6047_0[1]),.dinb(n6043),.dout(n6048),.clk(gclk));
	jor g05819(.dina(n6048),.dinb(w_n6042_0[1]),.dout(n6049),.clk(gclk));
	jand g05820(.dina(w_n6049_0[2]),.dinb(w_asqrt43_27[0]),.dout(n6050),.clk(gclk));
	jor g05821(.dina(w_n6049_0[1]),.dinb(w_asqrt43_26[2]),.dout(n6051),.clk(gclk));
	jxor g05822(.dina(w_n5666_0[0]),.dinb(w_n3368_45[1]),.dout(n6052),.clk(gclk));
	jand g05823(.dina(n6052),.dinb(w_asqrt34_35[2]),.dout(n6053),.clk(gclk));
	jxor g05824(.dina(n6053),.dinb(w_n5671_0[0]),.dout(n6054),.clk(gclk));
	jand g05825(.dina(w_n6054_0[1]),.dinb(n6051),.dout(n6055),.clk(gclk));
	jor g05826(.dina(n6055),.dinb(w_n6050_0[1]),.dout(n6056),.clk(gclk));
	jand g05827(.dina(w_n6056_0[2]),.dinb(w_asqrt44_30[0]),.dout(n6057),.clk(gclk));
	jor g05828(.dina(w_n6056_0[1]),.dinb(w_asqrt44_29[2]),.dout(n6058),.clk(gclk));
	jxor g05829(.dina(w_n5674_0[0]),.dinb(w_n3089_48[2]),.dout(n6059),.clk(gclk));
	jand g05830(.dina(n6059),.dinb(w_asqrt34_35[1]),.dout(n6060),.clk(gclk));
	jxor g05831(.dina(n6060),.dinb(w_n5679_0[0]),.dout(n6061),.clk(gclk));
	jand g05832(.dina(w_n6061_0[1]),.dinb(n6058),.dout(n6062),.clk(gclk));
	jor g05833(.dina(n6062),.dinb(w_n6057_0[1]),.dout(n6063),.clk(gclk));
	jand g05834(.dina(w_n6063_0[2]),.dinb(w_asqrt45_27[2]),.dout(n6064),.clk(gclk));
	jor g05835(.dina(w_n6063_0[1]),.dinb(w_asqrt45_27[1]),.dout(n6065),.clk(gclk));
	jxor g05836(.dina(w_n5682_0[0]),.dinb(w_n2833_46[1]),.dout(n6066),.clk(gclk));
	jand g05837(.dina(n6066),.dinb(w_asqrt34_35[0]),.dout(n6067),.clk(gclk));
	jxor g05838(.dina(n6067),.dinb(w_n5687_0[0]),.dout(n6068),.clk(gclk));
	jand g05839(.dina(w_n6068_0[1]),.dinb(n6065),.dout(n6069),.clk(gclk));
	jor g05840(.dina(n6069),.dinb(w_n6064_0[1]),.dout(n6070),.clk(gclk));
	jand g05841(.dina(w_n6070_0[2]),.dinb(w_asqrt46_30[0]),.dout(n6071),.clk(gclk));
	jor g05842(.dina(w_n6070_0[1]),.dinb(w_asqrt46_29[2]),.dout(n6072),.clk(gclk));
	jxor g05843(.dina(w_n5690_0[0]),.dinb(w_n2572_49[0]),.dout(n6073),.clk(gclk));
	jand g05844(.dina(n6073),.dinb(w_asqrt34_34[2]),.dout(n6074),.clk(gclk));
	jxor g05845(.dina(n6074),.dinb(w_n5695_0[0]),.dout(n6075),.clk(gclk));
	jnot g05846(.din(w_n6075_0[1]),.dout(n6076),.clk(gclk));
	jand g05847(.dina(w_n6076_0[1]),.dinb(n6072),.dout(n6077),.clk(gclk));
	jor g05848(.dina(n6077),.dinb(w_n6071_0[1]),.dout(n6078),.clk(gclk));
	jand g05849(.dina(w_n6078_0[2]),.dinb(w_asqrt47_28[1]),.dout(n6079),.clk(gclk));
	jor g05850(.dina(w_n6078_0[1]),.dinb(w_asqrt47_28[0]),.dout(n6080),.clk(gclk));
	jxor g05851(.dina(w_n5697_0[0]),.dinb(w_n2345_47[0]),.dout(n6081),.clk(gclk));
	jand g05852(.dina(n6081),.dinb(w_asqrt34_34[1]),.dout(n6082),.clk(gclk));
	jxor g05853(.dina(n6082),.dinb(w_n5702_0[0]),.dout(n6083),.clk(gclk));
	jnot g05854(.din(w_n6083_0[1]),.dout(n6084),.clk(gclk));
	jand g05855(.dina(w_n6084_0[1]),.dinb(n6080),.dout(n6085),.clk(gclk));
	jor g05856(.dina(n6085),.dinb(w_n6079_0[1]),.dout(n6086),.clk(gclk));
	jand g05857(.dina(w_n6086_0[2]),.dinb(w_asqrt48_30[1]),.dout(n6087),.clk(gclk));
	jor g05858(.dina(w_n6086_0[1]),.dinb(w_asqrt48_30[0]),.dout(n6088),.clk(gclk));
	jxor g05859(.dina(w_n5704_0[0]),.dinb(w_n2108_49[2]),.dout(n6089),.clk(gclk));
	jand g05860(.dina(n6089),.dinb(w_asqrt34_34[0]),.dout(n6090),.clk(gclk));
	jxor g05861(.dina(n6090),.dinb(w_n5709_0[0]),.dout(n6091),.clk(gclk));
	jnot g05862(.din(w_n6091_0[1]),.dout(n6092),.clk(gclk));
	jand g05863(.dina(w_n6092_0[1]),.dinb(n6088),.dout(n6093),.clk(gclk));
	jor g05864(.dina(n6093),.dinb(w_n6087_0[1]),.dout(n6094),.clk(gclk));
	jand g05865(.dina(w_n6094_0[2]),.dinb(w_asqrt49_28[2]),.dout(n6095),.clk(gclk));
	jor g05866(.dina(w_n6094_0[1]),.dinb(w_asqrt49_28[1]),.dout(n6096),.clk(gclk));
	jxor g05867(.dina(w_n5711_0[0]),.dinb(w_n1912_48[0]),.dout(n6097),.clk(gclk));
	jand g05868(.dina(n6097),.dinb(w_asqrt34_33[2]),.dout(n6098),.clk(gclk));
	jxor g05869(.dina(n6098),.dinb(w_n5716_0[0]),.dout(n6099),.clk(gclk));
	jand g05870(.dina(w_n6099_0[1]),.dinb(n6096),.dout(n6100),.clk(gclk));
	jor g05871(.dina(n6100),.dinb(w_n6095_0[1]),.dout(n6101),.clk(gclk));
	jand g05872(.dina(w_n6101_0[2]),.dinb(w_asqrt50_30[2]),.dout(n6102),.clk(gclk));
	jor g05873(.dina(w_n6101_0[1]),.dinb(w_asqrt50_30[1]),.dout(n6103),.clk(gclk));
	jxor g05874(.dina(w_n5719_0[0]),.dinb(w_n1699_50[1]),.dout(n6104),.clk(gclk));
	jand g05875(.dina(n6104),.dinb(w_asqrt34_33[1]),.dout(n6105),.clk(gclk));
	jxor g05876(.dina(n6105),.dinb(w_n5724_0[0]),.dout(n6106),.clk(gclk));
	jnot g05877(.din(w_n6106_0[1]),.dout(n6107),.clk(gclk));
	jand g05878(.dina(w_n6107_0[1]),.dinb(n6103),.dout(n6108),.clk(gclk));
	jor g05879(.dina(n6108),.dinb(w_n6102_0[1]),.dout(n6109),.clk(gclk));
	jand g05880(.dina(w_n6109_0[2]),.dinb(w_asqrt51_29[0]),.dout(n6110),.clk(gclk));
	jor g05881(.dina(w_n6109_0[1]),.dinb(w_asqrt51_28[2]),.dout(n6111),.clk(gclk));
	jxor g05882(.dina(w_n5726_0[0]),.dinb(w_n1516_48[2]),.dout(n6112),.clk(gclk));
	jand g05883(.dina(n6112),.dinb(w_asqrt34_33[0]),.dout(n6113),.clk(gclk));
	jxor g05884(.dina(n6113),.dinb(w_n5731_0[0]),.dout(n6114),.clk(gclk));
	jand g05885(.dina(w_n6114_0[1]),.dinb(n6111),.dout(n6115),.clk(gclk));
	jor g05886(.dina(n6115),.dinb(w_n6110_0[1]),.dout(n6116),.clk(gclk));
	jand g05887(.dina(w_n6116_0[2]),.dinb(w_asqrt52_30[2]),.dout(n6117),.clk(gclk));
	jor g05888(.dina(w_n6116_0[1]),.dinb(w_asqrt52_30[1]),.dout(n6118),.clk(gclk));
	jxor g05889(.dina(w_n5734_0[0]),.dinb(w_n1332_50[1]),.dout(n6119),.clk(gclk));
	jand g05890(.dina(n6119),.dinb(w_asqrt34_32[2]),.dout(n6120),.clk(gclk));
	jxor g05891(.dina(n6120),.dinb(w_n5739_0[0]),.dout(n6121),.clk(gclk));
	jnot g05892(.din(w_n6121_0[1]),.dout(n6122),.clk(gclk));
	jand g05893(.dina(w_n6122_0[1]),.dinb(n6118),.dout(n6123),.clk(gclk));
	jor g05894(.dina(n6123),.dinb(w_n6117_0[1]),.dout(n6124),.clk(gclk));
	jand g05895(.dina(w_n6124_0[2]),.dinb(w_asqrt53_29[2]),.dout(n6125),.clk(gclk));
	jor g05896(.dina(w_n6124_0[1]),.dinb(w_asqrt53_29[1]),.dout(n6126),.clk(gclk));
	jxor g05897(.dina(w_n5741_0[0]),.dinb(w_n1173_49[1]),.dout(n6127),.clk(gclk));
	jand g05898(.dina(n6127),.dinb(w_asqrt34_32[1]),.dout(n6128),.clk(gclk));
	jxor g05899(.dina(n6128),.dinb(w_n5746_0[0]),.dout(n6129),.clk(gclk));
	jand g05900(.dina(w_n6129_0[1]),.dinb(n6126),.dout(n6130),.clk(gclk));
	jor g05901(.dina(n6130),.dinb(w_n6125_0[1]),.dout(n6131),.clk(gclk));
	jand g05902(.dina(w_n6131_0[2]),.dinb(w_asqrt54_30[2]),.dout(n6132),.clk(gclk));
	jor g05903(.dina(w_n6131_0[1]),.dinb(w_asqrt54_30[1]),.dout(n6133),.clk(gclk));
	jxor g05904(.dina(w_n5749_0[0]),.dinb(w_n1008_51[1]),.dout(n6134),.clk(gclk));
	jand g05905(.dina(n6134),.dinb(w_asqrt34_32[0]),.dout(n6135),.clk(gclk));
	jxor g05906(.dina(n6135),.dinb(w_n5754_0[0]),.dout(n6136),.clk(gclk));
	jand g05907(.dina(w_n6136_0[1]),.dinb(n6133),.dout(n6137),.clk(gclk));
	jor g05908(.dina(n6137),.dinb(w_n6132_0[1]),.dout(n6138),.clk(gclk));
	jand g05909(.dina(w_n6138_0[2]),.dinb(w_asqrt55_30[0]),.dout(n6139),.clk(gclk));
	jor g05910(.dina(w_n6138_0[1]),.dinb(w_asqrt55_29[2]),.dout(n6140),.clk(gclk));
	jxor g05911(.dina(w_n5757_0[0]),.dinb(w_n884_50[1]),.dout(n6141),.clk(gclk));
	jand g05912(.dina(n6141),.dinb(w_asqrt34_31[2]),.dout(n6142),.clk(gclk));
	jxor g05913(.dina(n6142),.dinb(w_n5762_0[0]),.dout(n6143),.clk(gclk));
	jnot g05914(.din(w_n6143_0[1]),.dout(n6144),.clk(gclk));
	jand g05915(.dina(w_n6144_0[1]),.dinb(n6140),.dout(n6145),.clk(gclk));
	jor g05916(.dina(n6145),.dinb(w_n6139_0[1]),.dout(n6146),.clk(gclk));
	jand g05917(.dina(w_n6146_0[2]),.dinb(w_asqrt56_31[0]),.dout(n6147),.clk(gclk));
	jor g05918(.dina(w_n6146_0[1]),.dinb(w_asqrt56_30[2]),.dout(n6148),.clk(gclk));
	jxor g05919(.dina(w_n5764_0[0]),.dinb(w_n743_51[1]),.dout(n6149),.clk(gclk));
	jand g05920(.dina(n6149),.dinb(w_asqrt34_31[1]),.dout(n6150),.clk(gclk));
	jxor g05921(.dina(n6150),.dinb(w_n5769_0[0]),.dout(n6151),.clk(gclk));
	jnot g05922(.din(w_n6151_0[1]),.dout(n6152),.clk(gclk));
	jand g05923(.dina(w_n6152_0[1]),.dinb(n6148),.dout(n6153),.clk(gclk));
	jor g05924(.dina(n6153),.dinb(w_n6147_0[1]),.dout(n6154),.clk(gclk));
	jand g05925(.dina(w_n6154_0[2]),.dinb(w_asqrt57_30[2]),.dout(n6155),.clk(gclk));
	jor g05926(.dina(w_n6154_0[1]),.dinb(w_asqrt57_30[1]),.dout(n6156),.clk(gclk));
	jxor g05927(.dina(w_n5771_0[0]),.dinb(w_n635_51[1]),.dout(n6157),.clk(gclk));
	jand g05928(.dina(n6157),.dinb(w_asqrt34_31[0]),.dout(n6158),.clk(gclk));
	jxor g05929(.dina(n6158),.dinb(w_n5776_0[0]),.dout(n6159),.clk(gclk));
	jand g05930(.dina(w_n6159_0[1]),.dinb(n6156),.dout(n6160),.clk(gclk));
	jor g05931(.dina(n6160),.dinb(w_n6155_0[1]),.dout(n6161),.clk(gclk));
	jand g05932(.dina(w_n6161_0[2]),.dinb(w_asqrt58_31[1]),.dout(n6162),.clk(gclk));
	jor g05933(.dina(w_n6161_0[1]),.dinb(w_asqrt58_31[0]),.dout(n6163),.clk(gclk));
	jxor g05934(.dina(w_n5779_0[0]),.dinb(w_n515_52[1]),.dout(n6164),.clk(gclk));
	jand g05935(.dina(n6164),.dinb(w_asqrt34_30[2]),.dout(n6165),.clk(gclk));
	jxor g05936(.dina(n6165),.dinb(w_n5784_0[0]),.dout(n6166),.clk(gclk));
	jnot g05937(.din(w_n6166_0[2]),.dout(n6167),.clk(gclk));
	jand g05938(.dina(n6167),.dinb(n6163),.dout(n6168),.clk(gclk));
	jor g05939(.dina(n6168),.dinb(w_n6162_0[1]),.dout(n6169),.clk(gclk));
	jand g05940(.dina(w_n6169_0[2]),.dinb(w_asqrt59_31[0]),.dout(n6170),.clk(gclk));
	jor g05941(.dina(w_n6169_0[1]),.dinb(w_asqrt59_30[2]),.dout(n6171),.clk(gclk));
	jxor g05942(.dina(w_n5786_0[0]),.dinb(w_n443_52[1]),.dout(n6172),.clk(gclk));
	jand g05943(.dina(n6172),.dinb(w_asqrt34_30[1]),.dout(n6173),.clk(gclk));
	jxor g05944(.dina(n6173),.dinb(w_n5791_0[0]),.dout(n6174),.clk(gclk));
	jand g05945(.dina(w_n6174_0[1]),.dinb(n6171),.dout(n6175),.clk(gclk));
	jor g05946(.dina(n6175),.dinb(w_n6170_0[1]),.dout(n6176),.clk(gclk));
	jand g05947(.dina(w_n6176_0[2]),.dinb(w_asqrt60_31[1]),.dout(n6177),.clk(gclk));
	jor g05948(.dina(w_n6176_0[1]),.dinb(w_asqrt60_31[0]),.dout(n6178),.clk(gclk));
	jxor g05949(.dina(w_n5794_0[0]),.dinb(w_n352_52[2]),.dout(n6179),.clk(gclk));
	jand g05950(.dina(n6179),.dinb(w_asqrt34_30[0]),.dout(n6180),.clk(gclk));
	jxor g05951(.dina(n6180),.dinb(w_n5799_0[0]),.dout(n6181),.clk(gclk));
	jnot g05952(.din(w_n6181_0[1]),.dout(n6182),.clk(gclk));
	jand g05953(.dina(w_n6182_0[1]),.dinb(n6178),.dout(n6183),.clk(gclk));
	jor g05954(.dina(n6183),.dinb(w_n6177_0[1]),.dout(n6184),.clk(gclk));
	jand g05955(.dina(w_n6184_0[2]),.dinb(w_asqrt61_31[1]),.dout(n6185),.clk(gclk));
	jor g05956(.dina(w_n6184_0[1]),.dinb(w_asqrt61_31[0]),.dout(n6186),.clk(gclk));
	jxor g05957(.dina(w_n5801_0[0]),.dinb(w_n294_53[0]),.dout(n6187),.clk(gclk));
	jand g05958(.dina(n6187),.dinb(w_asqrt34_29[2]),.dout(n6188),.clk(gclk));
	jxor g05959(.dina(n6188),.dinb(w_n5806_0[0]),.dout(n6189),.clk(gclk));
	jnot g05960(.din(w_n6189_0[1]),.dout(n6190),.clk(gclk));
	jand g05961(.dina(w_n6190_0[1]),.dinb(n6186),.dout(n6191),.clk(gclk));
	jor g05962(.dina(n6191),.dinb(w_n6185_0[1]),.dout(n6192),.clk(gclk));
	jand g05963(.dina(w_n6192_0[2]),.dinb(w_asqrt62_31[1]),.dout(n6193),.clk(gclk));
	jor g05964(.dina(w_n6192_0[1]),.dinb(w_asqrt62_31[0]),.dout(n6194),.clk(gclk));
	jxor g05965(.dina(w_n5808_0[0]),.dinb(w_n239_53[0]),.dout(n6195),.clk(gclk));
	jand g05966(.dina(n6195),.dinb(w_asqrt34_29[1]),.dout(n6196),.clk(gclk));
	jxor g05967(.dina(n6196),.dinb(w_n5813_0[0]),.dout(n6197),.clk(gclk));
	jnot g05968(.din(w_n6197_0[2]),.dout(n6198),.clk(gclk));
	jand g05969(.dina(n6198),.dinb(n6194),.dout(n6199),.clk(gclk));
	jor g05970(.dina(n6199),.dinb(w_n6193_0[1]),.dout(n6200),.clk(gclk));
	jor g05971(.dina(w_n6200_0[1]),.dinb(w_n5842_0[2]),.dout(n6201),.clk(gclk));
	jnot g05972(.din(w_n6201_1[1]),.dout(n6202),.clk(gclk));
	jnot g05973(.din(w_n5842_0[1]),.dout(n6204),.clk(gclk));
	jnot g05974(.din(w_n6193_0[0]),.dout(n6205),.clk(gclk));
	jnot g05975(.din(w_n6185_0[0]),.dout(n6206),.clk(gclk));
	jnot g05976(.din(w_n6177_0[0]),.dout(n6207),.clk(gclk));
	jnot g05977(.din(w_n6170_0[0]),.dout(n6208),.clk(gclk));
	jnot g05978(.din(w_n6162_0[0]),.dout(n6209),.clk(gclk));
	jnot g05979(.din(w_n6155_0[0]),.dout(n6210),.clk(gclk));
	jnot g05980(.din(w_n6147_0[0]),.dout(n6211),.clk(gclk));
	jnot g05981(.din(w_n6139_0[0]),.dout(n6212),.clk(gclk));
	jnot g05982(.din(w_n6132_0[0]),.dout(n6213),.clk(gclk));
	jnot g05983(.din(w_n6125_0[0]),.dout(n6214),.clk(gclk));
	jnot g05984(.din(w_n6117_0[0]),.dout(n6215),.clk(gclk));
	jnot g05985(.din(w_n6110_0[0]),.dout(n6216),.clk(gclk));
	jnot g05986(.din(w_n6102_0[0]),.dout(n6217),.clk(gclk));
	jnot g05987(.din(w_n6095_0[0]),.dout(n6218),.clk(gclk));
	jnot g05988(.din(w_n6087_0[0]),.dout(n6219),.clk(gclk));
	jnot g05989(.din(w_n6079_0[0]),.dout(n6220),.clk(gclk));
	jnot g05990(.din(w_n6071_0[0]),.dout(n6221),.clk(gclk));
	jnot g05991(.din(w_n6064_0[0]),.dout(n6222),.clk(gclk));
	jnot g05992(.din(w_n6057_0[0]),.dout(n6223),.clk(gclk));
	jnot g05993(.din(w_n6050_0[0]),.dout(n6224),.clk(gclk));
	jnot g05994(.din(w_n6042_0[0]),.dout(n6225),.clk(gclk));
	jnot g05995(.din(w_n6035_0[0]),.dout(n6226),.clk(gclk));
	jnot g05996(.din(w_n6027_0[0]),.dout(n6227),.clk(gclk));
	jnot g05997(.din(w_n6020_0[0]),.dout(n6228),.clk(gclk));
	jnot g05998(.din(w_n6012_0[0]),.dout(n6229),.clk(gclk));
	jnot g05999(.din(w_n6005_0[0]),.dout(n6230),.clk(gclk));
	jnot g06000(.din(w_n5994_0[0]),.dout(n6231),.clk(gclk));
	jnot g06001(.din(w_n5849_0[0]),.dout(n6232),.clk(gclk));
	jnot g06002(.din(w_n5846_0[0]),.dout(n6233),.clk(gclk));
	jor g06003(.dina(w_n5989_42[0]),.dinb(w_n5612_0[2]),.dout(n6234),.clk(gclk));
	jand g06004(.dina(n6234),.dinb(n6233),.dout(n6235),.clk(gclk));
	jand g06005(.dina(n6235),.dinb(w_n5606_46[0]),.dout(n6236),.clk(gclk));
	jor g06006(.dina(w_n5989_41[2]),.dinb(w_a68_0[0]),.dout(n6237),.clk(gclk));
	jand g06007(.dina(n6237),.dinb(w_a69_0[0]),.dout(n6238),.clk(gclk));
	jor g06008(.dina(w_n5996_0[0]),.dinb(n6238),.dout(n6239),.clk(gclk));
	jor g06009(.dina(w_n6239_0[1]),.dinb(n6236),.dout(n6240),.clk(gclk));
	jand g06010(.dina(n6240),.dinb(n6232),.dout(n6241),.clk(gclk));
	jand g06011(.dina(n6241),.dinb(w_n5259_42[2]),.dout(n6242),.clk(gclk));
	jor g06012(.dina(w_n6001_0[0]),.dinb(n6242),.dout(n6243),.clk(gclk));
	jand g06013(.dina(n6243),.dinb(n6231),.dout(n6244),.clk(gclk));
	jand g06014(.dina(n6244),.dinb(w_n4902_46[2]),.dout(n6245),.clk(gclk));
	jnot g06015(.din(w_n6009_0[0]),.dout(n6246),.clk(gclk));
	jor g06016(.dina(w_n6246_0[1]),.dinb(n6245),.dout(n6247),.clk(gclk));
	jand g06017(.dina(n6247),.dinb(n6230),.dout(n6248),.clk(gclk));
	jand g06018(.dina(n6248),.dinb(w_n4582_43[2]),.dout(n6249),.clk(gclk));
	jor g06019(.dina(w_n6016_0[0]),.dinb(n6249),.dout(n6250),.clk(gclk));
	jand g06020(.dina(n6250),.dinb(n6229),.dout(n6251),.clk(gclk));
	jand g06021(.dina(n6251),.dinb(w_n4249_47[1]),.dout(n6252),.clk(gclk));
	jnot g06022(.din(w_n6024_0[0]),.dout(n6253),.clk(gclk));
	jor g06023(.dina(w_n6253_0[1]),.dinb(n6252),.dout(n6254),.clk(gclk));
	jand g06024(.dina(n6254),.dinb(n6228),.dout(n6255),.clk(gclk));
	jand g06025(.dina(n6255),.dinb(w_n3955_44[1]),.dout(n6256),.clk(gclk));
	jor g06026(.dina(w_n6031_0[0]),.dinb(n6256),.dout(n6257),.clk(gclk));
	jand g06027(.dina(n6257),.dinb(n6227),.dout(n6258),.clk(gclk));
	jand g06028(.dina(n6258),.dinb(w_n3642_47[2]),.dout(n6259),.clk(gclk));
	jnot g06029(.din(w_n6039_0[0]),.dout(n6260),.clk(gclk));
	jor g06030(.dina(w_n6260_0[1]),.dinb(n6259),.dout(n6261),.clk(gclk));
	jand g06031(.dina(n6261),.dinb(n6226),.dout(n6262),.clk(gclk));
	jand g06032(.dina(n6262),.dinb(w_n3368_45[0]),.dout(n6263),.clk(gclk));
	jor g06033(.dina(w_n6046_0[0]),.dinb(n6263),.dout(n6264),.clk(gclk));
	jand g06034(.dina(n6264),.dinb(n6225),.dout(n6265),.clk(gclk));
	jand g06035(.dina(n6265),.dinb(w_n3089_48[1]),.dout(n6266),.clk(gclk));
	jnot g06036(.din(w_n6054_0[0]),.dout(n6267),.clk(gclk));
	jor g06037(.dina(w_n6267_0[1]),.dinb(n6266),.dout(n6268),.clk(gclk));
	jand g06038(.dina(n6268),.dinb(n6224),.dout(n6269),.clk(gclk));
	jand g06039(.dina(n6269),.dinb(w_n2833_46[0]),.dout(n6270),.clk(gclk));
	jnot g06040(.din(w_n6061_0[0]),.dout(n6271),.clk(gclk));
	jor g06041(.dina(w_n6271_0[1]),.dinb(n6270),.dout(n6272),.clk(gclk));
	jand g06042(.dina(n6272),.dinb(n6223),.dout(n6273),.clk(gclk));
	jand g06043(.dina(n6273),.dinb(w_n2572_48[2]),.dout(n6274),.clk(gclk));
	jnot g06044(.din(w_n6068_0[0]),.dout(n6275),.clk(gclk));
	jor g06045(.dina(w_n6275_0[1]),.dinb(n6274),.dout(n6276),.clk(gclk));
	jand g06046(.dina(n6276),.dinb(n6222),.dout(n6277),.clk(gclk));
	jand g06047(.dina(n6277),.dinb(w_n2345_46[2]),.dout(n6278),.clk(gclk));
	jor g06048(.dina(w_n6075_0[0]),.dinb(n6278),.dout(n6279),.clk(gclk));
	jand g06049(.dina(n6279),.dinb(n6221),.dout(n6280),.clk(gclk));
	jand g06050(.dina(n6280),.dinb(w_n2108_49[1]),.dout(n6281),.clk(gclk));
	jor g06051(.dina(w_n6083_0[0]),.dinb(n6281),.dout(n6282),.clk(gclk));
	jand g06052(.dina(n6282),.dinb(n6220),.dout(n6283),.clk(gclk));
	jand g06053(.dina(n6283),.dinb(w_n1912_47[2]),.dout(n6284),.clk(gclk));
	jor g06054(.dina(w_n6091_0[0]),.dinb(n6284),.dout(n6285),.clk(gclk));
	jand g06055(.dina(n6285),.dinb(n6219),.dout(n6286),.clk(gclk));
	jand g06056(.dina(n6286),.dinb(w_n1699_50[0]),.dout(n6287),.clk(gclk));
	jnot g06057(.din(w_n6099_0[0]),.dout(n6288),.clk(gclk));
	jor g06058(.dina(w_n6288_0[1]),.dinb(n6287),.dout(n6289),.clk(gclk));
	jand g06059(.dina(n6289),.dinb(n6218),.dout(n6290),.clk(gclk));
	jand g06060(.dina(n6290),.dinb(w_n1516_48[1]),.dout(n6291),.clk(gclk));
	jor g06061(.dina(w_n6106_0[0]),.dinb(n6291),.dout(n6292),.clk(gclk));
	jand g06062(.dina(n6292),.dinb(n6217),.dout(n6293),.clk(gclk));
	jand g06063(.dina(n6293),.dinb(w_n1332_50[0]),.dout(n6294),.clk(gclk));
	jnot g06064(.din(w_n6114_0[0]),.dout(n6295),.clk(gclk));
	jor g06065(.dina(w_n6295_0[1]),.dinb(n6294),.dout(n6296),.clk(gclk));
	jand g06066(.dina(n6296),.dinb(n6216),.dout(n6297),.clk(gclk));
	jand g06067(.dina(n6297),.dinb(w_n1173_49[0]),.dout(n6298),.clk(gclk));
	jor g06068(.dina(w_n6121_0[0]),.dinb(n6298),.dout(n6299),.clk(gclk));
	jand g06069(.dina(n6299),.dinb(n6215),.dout(n6300),.clk(gclk));
	jand g06070(.dina(n6300),.dinb(w_n1008_51[0]),.dout(n6301),.clk(gclk));
	jnot g06071(.din(w_n6129_0[0]),.dout(n6302),.clk(gclk));
	jor g06072(.dina(w_n6302_0[1]),.dinb(n6301),.dout(n6303),.clk(gclk));
	jand g06073(.dina(n6303),.dinb(n6214),.dout(n6304),.clk(gclk));
	jand g06074(.dina(n6304),.dinb(w_n884_50[0]),.dout(n6305),.clk(gclk));
	jnot g06075(.din(w_n6136_0[0]),.dout(n6306),.clk(gclk));
	jor g06076(.dina(w_n6306_0[1]),.dinb(n6305),.dout(n6307),.clk(gclk));
	jand g06077(.dina(n6307),.dinb(n6213),.dout(n6308),.clk(gclk));
	jand g06078(.dina(n6308),.dinb(w_n743_51[0]),.dout(n6309),.clk(gclk));
	jor g06079(.dina(w_n6143_0[0]),.dinb(n6309),.dout(n6310),.clk(gclk));
	jand g06080(.dina(n6310),.dinb(n6212),.dout(n6311),.clk(gclk));
	jand g06081(.dina(n6311),.dinb(w_n635_51[0]),.dout(n6312),.clk(gclk));
	jor g06082(.dina(w_n6151_0[0]),.dinb(n6312),.dout(n6313),.clk(gclk));
	jand g06083(.dina(n6313),.dinb(n6211),.dout(n6314),.clk(gclk));
	jand g06084(.dina(n6314),.dinb(w_n515_52[0]),.dout(n6315),.clk(gclk));
	jnot g06085(.din(w_n6159_0[0]),.dout(n6316),.clk(gclk));
	jor g06086(.dina(w_n6316_0[1]),.dinb(n6315),.dout(n6317),.clk(gclk));
	jand g06087(.dina(n6317),.dinb(n6210),.dout(n6318),.clk(gclk));
	jand g06088(.dina(n6318),.dinb(w_n443_52[0]),.dout(n6319),.clk(gclk));
	jor g06089(.dina(w_n6166_0[1]),.dinb(n6319),.dout(n6320),.clk(gclk));
	jand g06090(.dina(n6320),.dinb(n6209),.dout(n6321),.clk(gclk));
	jand g06091(.dina(n6321),.dinb(w_n352_52[1]),.dout(n6322),.clk(gclk));
	jnot g06092(.din(w_n6174_0[0]),.dout(n6323),.clk(gclk));
	jor g06093(.dina(w_n6323_0[1]),.dinb(n6322),.dout(n6324),.clk(gclk));
	jand g06094(.dina(n6324),.dinb(n6208),.dout(n6325),.clk(gclk));
	jand g06095(.dina(n6325),.dinb(w_n294_52[2]),.dout(n6326),.clk(gclk));
	jor g06096(.dina(w_n6181_0[0]),.dinb(n6326),.dout(n6327),.clk(gclk));
	jand g06097(.dina(n6327),.dinb(n6207),.dout(n6328),.clk(gclk));
	jand g06098(.dina(n6328),.dinb(w_n239_52[2]),.dout(n6329),.clk(gclk));
	jor g06099(.dina(w_n6189_0[0]),.dinb(n6329),.dout(n6330),.clk(gclk));
	jand g06100(.dina(n6330),.dinb(n6206),.dout(n6331),.clk(gclk));
	jand g06101(.dina(n6331),.dinb(w_n221_53[0]),.dout(n6332),.clk(gclk));
	jor g06102(.dina(w_n6197_0[1]),.dinb(n6332),.dout(n6333),.clk(gclk));
	jand g06103(.dina(n6333),.dinb(n6205),.dout(n6334),.clk(gclk));
	jor g06104(.dina(w_n6334_0[1]),.dinb(w_n6204_0[1]),.dout(n6335),.clk(gclk));
	jxor g06105(.dina(w_n5823_0[2]),.dinb(w_n5610_0[0]),.dout(n6336),.clk(gclk));
	jnot g06106(.din(w_n6336_0[1]),.dout(n6337),.clk(gclk));
	jand g06107(.dina(n6337),.dinb(w_asqrt34_29[0]),.dout(n6338),.clk(gclk));
	jor g06108(.dina(w_n6338_0[1]),.dinb(w_n6335_0[1]),.dout(n6339),.clk(gclk));
	jand g06109(.dina(n6339),.dinb(w_n218_22[0]),.dout(n6340),.clk(gclk));
	jand g06110(.dina(w_n5987_0[0]),.dinb(w_n5823_0[1]),.dout(n6341),.clk(gclk));
	jnot g06111(.din(n6341),.dout(n6342),.clk(gclk));
	jand g06112(.dina(w_n6336_0[0]),.dinb(w_asqrt63_40[0]),.dout(n6343),.clk(gclk));
	jand g06113(.dina(w_n6343_0[1]),.dinb(n6342),.dout(n6344),.clk(gclk));
	jor g06114(.dina(w_n6344_0[1]),.dinb(w_n6340_0[1]),.dout(n6345),.clk(gclk));
	jor g06115(.dina(w_n6345_0[1]),.dinb(w_n6202_0[2]),.dout(asqrt_fa_34),.clk(gclk));
	jand g06116(.dina(w_n6200_0[0]),.dinb(w_n5842_0[0]),.dout(n6348),.clk(gclk));
	jand g06117(.dina(w_n6345_0[0]),.dinb(w_n6348_0[1]),.dout(n6349),.clk(gclk));
	jnot g06118(.din(w_n6338_0[0]),.dout(n6351),.clk(gclk));
	jand g06119(.dina(n6351),.dinb(w_n6348_0[0]),.dout(n6352),.clk(gclk));
	jor g06120(.dina(n6352),.dinb(w_asqrt63_39[2]),.dout(n6353),.clk(gclk));
	jnot g06121(.din(w_n6344_0[0]),.dout(n6354),.clk(gclk));
	jand g06122(.dina(n6354),.dinb(n6353),.dout(n6355),.clk(gclk));
	jand g06123(.dina(w_n6355_0[1]),.dinb(w_n6201_1[0]),.dout(n6357),.clk(gclk));
	jxor g06124(.dina(w_n6192_0[0]),.dinb(w_n221_52[2]),.dout(n6358),.clk(gclk));
	jor g06125(.dina(n6358),.dinb(w_n6357_54[2]),.dout(n6359),.clk(gclk));
	jxor g06126(.dina(n6359),.dinb(w_n6197_0[0]),.dout(n6360),.clk(gclk));
	jnot g06127(.din(w_n6360_0[1]),.dout(n6361),.clk(gclk));
	jnot g06128(.din(w_a64_0[2]),.dout(n6362),.clk(gclk));
	jnot g06129(.din(w_a65_0[1]),.dout(n6363),.clk(gclk));
	jand g06130(.dina(w_n6363_0[1]),.dinb(w_n6362_1[2]),.dout(n6364),.clk(gclk));
	jand g06131(.dina(w_n6364_0[2]),.dinb(w_n5843_1[0]),.dout(n6365),.clk(gclk));
	jnot g06132(.din(w_n6365_0[1]),.dout(n6366),.clk(gclk));
	jor g06133(.dina(w_n6357_54[1]),.dinb(w_n5843_0[2]),.dout(n6367),.clk(gclk));
	jand g06134(.dina(n6367),.dinb(n6366),.dout(n6368),.clk(gclk));
	jor g06135(.dina(w_n6368_0[2]),.dinb(w_n5989_41[1]),.dout(n6369),.clk(gclk));
	jand g06136(.dina(w_n6368_0[1]),.dinb(w_n5989_41[0]),.dout(n6370),.clk(gclk));
	jor g06137(.dina(w_n6357_54[0]),.dinb(w_a66_1[0]),.dout(n6371),.clk(gclk));
	jand g06138(.dina(n6371),.dinb(w_a67_0[0]),.dout(n6372),.clk(gclk));
	jand g06139(.dina(w_asqrt33_25),.dinb(w_n5845_0[1]),.dout(n6373),.clk(gclk));
	jor g06140(.dina(n6373),.dinb(n6372),.dout(n6374),.clk(gclk));
	jor g06141(.dina(n6374),.dinb(n6370),.dout(n6375),.clk(gclk));
	jand g06142(.dina(n6375),.dinb(w_n6369_0[1]),.dout(n6376),.clk(gclk));
	jor g06143(.dina(w_n6376_0[2]),.dinb(w_n5606_45[2]),.dout(n6377),.clk(gclk));
	jand g06144(.dina(w_n6376_0[1]),.dinb(w_n5606_45[1]),.dout(n6378),.clk(gclk));
	jnot g06145(.din(w_n5845_0[0]),.dout(n6379),.clk(gclk));
	jor g06146(.dina(w_n6357_53[2]),.dinb(n6379),.dout(n6380),.clk(gclk));
	jor g06147(.dina(w_n6343_0[0]),.dinb(w_n6202_0[1]),.dout(n6381),.clk(gclk));
	jor g06148(.dina(n6381),.dinb(w_n6340_0[0]),.dout(n6382),.clk(gclk));
	jor g06149(.dina(n6382),.dinb(w_n5989_40[2]),.dout(n6383),.clk(gclk));
	jand g06150(.dina(n6383),.dinb(w_n6380_0[1]),.dout(n6384),.clk(gclk));
	jxor g06151(.dina(n6384),.dinb(w_n5612_0[1]),.dout(n6385),.clk(gclk));
	jor g06152(.dina(w_n6385_0[1]),.dinb(n6378),.dout(n6386),.clk(gclk));
	jand g06153(.dina(n6386),.dinb(w_n6377_0[1]),.dout(n6387),.clk(gclk));
	jor g06154(.dina(w_n6387_0[2]),.dinb(w_n5259_42[1]),.dout(n6388),.clk(gclk));
	jand g06155(.dina(w_n6387_0[1]),.dinb(w_n5259_42[0]),.dout(n6389),.clk(gclk));
	jxor g06156(.dina(w_n5848_0[0]),.dinb(w_n5606_45[0]),.dout(n6390),.clk(gclk));
	jor g06157(.dina(n6390),.dinb(w_n6357_53[1]),.dout(n6391),.clk(gclk));
	jxor g06158(.dina(n6391),.dinb(w_n6239_0[0]),.dout(n6392),.clk(gclk));
	jnot g06159(.din(w_n6392_0[2]),.dout(n6393),.clk(gclk));
	jor g06160(.dina(n6393),.dinb(n6389),.dout(n6394),.clk(gclk));
	jand g06161(.dina(n6394),.dinb(w_n6388_0[1]),.dout(n6395),.clk(gclk));
	jor g06162(.dina(w_n6395_0[2]),.dinb(w_n4902_46[1]),.dout(n6396),.clk(gclk));
	jand g06163(.dina(w_n6395_0[1]),.dinb(w_n4902_46[0]),.dout(n6397),.clk(gclk));
	jxor g06164(.dina(w_n5993_0[0]),.dinb(w_n5259_41[2]),.dout(n6398),.clk(gclk));
	jor g06165(.dina(n6398),.dinb(w_n6357_53[0]),.dout(n6399),.clk(gclk));
	jxor g06166(.dina(n6399),.dinb(w_n6002_0[0]),.dout(n6400),.clk(gclk));
	jor g06167(.dina(w_n6400_0[2]),.dinb(n6397),.dout(n6401),.clk(gclk));
	jand g06168(.dina(n6401),.dinb(w_n6396_0[1]),.dout(n6402),.clk(gclk));
	jor g06169(.dina(w_n6402_0[2]),.dinb(w_n4582_43[1]),.dout(n6403),.clk(gclk));
	jand g06170(.dina(w_n6402_0[1]),.dinb(w_n4582_43[0]),.dout(n6404),.clk(gclk));
	jxor g06171(.dina(w_n6004_0[0]),.dinb(w_n4902_45[2]),.dout(n6405),.clk(gclk));
	jor g06172(.dina(n6405),.dinb(w_n6357_52[2]),.dout(n6406),.clk(gclk));
	jxor g06173(.dina(n6406),.dinb(w_n6246_0[0]),.dout(n6407),.clk(gclk));
	jnot g06174(.din(w_n6407_0[2]),.dout(n6408),.clk(gclk));
	jor g06175(.dina(n6408),.dinb(n6404),.dout(n6409),.clk(gclk));
	jand g06176(.dina(n6409),.dinb(w_n6403_0[1]),.dout(n6410),.clk(gclk));
	jor g06177(.dina(w_n6410_0[2]),.dinb(w_n4249_47[0]),.dout(n6411),.clk(gclk));
	jand g06178(.dina(w_n6410_0[1]),.dinb(w_n4249_46[2]),.dout(n6412),.clk(gclk));
	jxor g06179(.dina(w_n6011_0[0]),.dinb(w_n4582_42[2]),.dout(n6413),.clk(gclk));
	jor g06180(.dina(n6413),.dinb(w_n6357_52[1]),.dout(n6414),.clk(gclk));
	jxor g06181(.dina(n6414),.dinb(w_n6017_0[0]),.dout(n6415),.clk(gclk));
	jor g06182(.dina(w_n6415_0[2]),.dinb(n6412),.dout(n6416),.clk(gclk));
	jand g06183(.dina(n6416),.dinb(w_n6411_0[1]),.dout(n6417),.clk(gclk));
	jor g06184(.dina(w_n6417_0[2]),.dinb(w_n3955_44[0]),.dout(n6418),.clk(gclk));
	jand g06185(.dina(w_n6417_0[1]),.dinb(w_n3955_43[2]),.dout(n6419),.clk(gclk));
	jxor g06186(.dina(w_n6019_0[0]),.dinb(w_n4249_46[1]),.dout(n6420),.clk(gclk));
	jor g06187(.dina(n6420),.dinb(w_n6357_52[0]),.dout(n6421),.clk(gclk));
	jxor g06188(.dina(n6421),.dinb(w_n6253_0[0]),.dout(n6422),.clk(gclk));
	jnot g06189(.din(w_n6422_0[2]),.dout(n6423),.clk(gclk));
	jor g06190(.dina(n6423),.dinb(n6419),.dout(n6424),.clk(gclk));
	jand g06191(.dina(n6424),.dinb(w_n6418_0[1]),.dout(n6425),.clk(gclk));
	jor g06192(.dina(w_n6425_0[2]),.dinb(w_n3642_47[1]),.dout(n6426),.clk(gclk));
	jand g06193(.dina(w_n6425_0[1]),.dinb(w_n3642_47[0]),.dout(n6427),.clk(gclk));
	jxor g06194(.dina(w_n6026_0[0]),.dinb(w_n3955_43[1]),.dout(n6428),.clk(gclk));
	jor g06195(.dina(n6428),.dinb(w_n6357_51[2]),.dout(n6429),.clk(gclk));
	jxor g06196(.dina(n6429),.dinb(w_n6032_0[0]),.dout(n6430),.clk(gclk));
	jor g06197(.dina(w_n6430_0[2]),.dinb(n6427),.dout(n6431),.clk(gclk));
	jand g06198(.dina(n6431),.dinb(w_n6426_0[1]),.dout(n6432),.clk(gclk));
	jor g06199(.dina(w_n6432_0[2]),.dinb(w_n3368_44[2]),.dout(n6433),.clk(gclk));
	jand g06200(.dina(w_n6432_0[1]),.dinb(w_n3368_44[1]),.dout(n6434),.clk(gclk));
	jxor g06201(.dina(w_n6034_0[0]),.dinb(w_n3642_46[2]),.dout(n6435),.clk(gclk));
	jor g06202(.dina(n6435),.dinb(w_n6357_51[1]),.dout(n6436),.clk(gclk));
	jxor g06203(.dina(n6436),.dinb(w_n6260_0[0]),.dout(n6437),.clk(gclk));
	jnot g06204(.din(w_n6437_0[2]),.dout(n6438),.clk(gclk));
	jor g06205(.dina(n6438),.dinb(n6434),.dout(n6439),.clk(gclk));
	jand g06206(.dina(n6439),.dinb(w_n6433_0[1]),.dout(n6440),.clk(gclk));
	jor g06207(.dina(w_n6440_0[2]),.dinb(w_n3089_48[0]),.dout(n6441),.clk(gclk));
	jand g06208(.dina(w_n6440_0[1]),.dinb(w_n3089_47[2]),.dout(n6442),.clk(gclk));
	jxor g06209(.dina(w_n6041_0[0]),.dinb(w_n3368_44[0]),.dout(n6443),.clk(gclk));
	jor g06210(.dina(n6443),.dinb(w_n6357_51[0]),.dout(n6444),.clk(gclk));
	jxor g06211(.dina(n6444),.dinb(w_n6047_0[0]),.dout(n6445),.clk(gclk));
	jor g06212(.dina(w_n6445_0[2]),.dinb(n6442),.dout(n6446),.clk(gclk));
	jand g06213(.dina(n6446),.dinb(w_n6441_0[1]),.dout(n6447),.clk(gclk));
	jor g06214(.dina(w_n6447_0[2]),.dinb(w_n2833_45[2]),.dout(n6448),.clk(gclk));
	jand g06215(.dina(w_n6447_0[1]),.dinb(w_n2833_45[1]),.dout(n6449),.clk(gclk));
	jxor g06216(.dina(w_n6049_0[0]),.dinb(w_n3089_47[1]),.dout(n6450),.clk(gclk));
	jor g06217(.dina(n6450),.dinb(w_n6357_50[2]),.dout(n6451),.clk(gclk));
	jxor g06218(.dina(n6451),.dinb(w_n6267_0[0]),.dout(n6452),.clk(gclk));
	jnot g06219(.din(w_n6452_0[2]),.dout(n6453),.clk(gclk));
	jor g06220(.dina(n6453),.dinb(n6449),.dout(n6454),.clk(gclk));
	jand g06221(.dina(n6454),.dinb(w_n6448_0[1]),.dout(n6455),.clk(gclk));
	jor g06222(.dina(w_n6455_0[2]),.dinb(w_n2572_48[1]),.dout(n6456),.clk(gclk));
	jand g06223(.dina(w_n6455_0[1]),.dinb(w_n2572_48[0]),.dout(n6457),.clk(gclk));
	jxor g06224(.dina(w_n6056_0[0]),.dinb(w_n2833_45[0]),.dout(n6458),.clk(gclk));
	jor g06225(.dina(n6458),.dinb(w_n6357_50[1]),.dout(n6459),.clk(gclk));
	jxor g06226(.dina(n6459),.dinb(w_n6271_0[0]),.dout(n6460),.clk(gclk));
	jnot g06227(.din(w_n6460_0[2]),.dout(n6461),.clk(gclk));
	jor g06228(.dina(n6461),.dinb(n6457),.dout(n6462),.clk(gclk));
	jand g06229(.dina(n6462),.dinb(w_n6456_0[1]),.dout(n6463),.clk(gclk));
	jor g06230(.dina(w_n6463_0[2]),.dinb(w_n2345_46[1]),.dout(n6464),.clk(gclk));
	jand g06231(.dina(w_n6463_0[1]),.dinb(w_n2345_46[0]),.dout(n6465),.clk(gclk));
	jxor g06232(.dina(w_n6063_0[0]),.dinb(w_n2572_47[2]),.dout(n6466),.clk(gclk));
	jor g06233(.dina(n6466),.dinb(w_n6357_50[0]),.dout(n6467),.clk(gclk));
	jxor g06234(.dina(n6467),.dinb(w_n6275_0[0]),.dout(n6468),.clk(gclk));
	jnot g06235(.din(w_n6468_0[2]),.dout(n6469),.clk(gclk));
	jor g06236(.dina(n6469),.dinb(n6465),.dout(n6470),.clk(gclk));
	jand g06237(.dina(n6470),.dinb(w_n6464_0[1]),.dout(n6471),.clk(gclk));
	jor g06238(.dina(w_n6471_0[2]),.dinb(w_n2108_49[0]),.dout(n6472),.clk(gclk));
	jand g06239(.dina(w_n6471_0[1]),.dinb(w_n2108_48[2]),.dout(n6473),.clk(gclk));
	jxor g06240(.dina(w_n6070_0[0]),.dinb(w_n2345_45[2]),.dout(n6474),.clk(gclk));
	jor g06241(.dina(n6474),.dinb(w_n6357_49[2]),.dout(n6475),.clk(gclk));
	jxor g06242(.dina(n6475),.dinb(w_n6076_0[0]),.dout(n6476),.clk(gclk));
	jor g06243(.dina(w_n6476_0[2]),.dinb(n6473),.dout(n6477),.clk(gclk));
	jand g06244(.dina(n6477),.dinb(w_n6472_0[1]),.dout(n6478),.clk(gclk));
	jor g06245(.dina(w_n6478_0[2]),.dinb(w_n1912_47[1]),.dout(n6479),.clk(gclk));
	jand g06246(.dina(w_n6478_0[1]),.dinb(w_n1912_47[0]),.dout(n6480),.clk(gclk));
	jxor g06247(.dina(w_n6078_0[0]),.dinb(w_n2108_48[1]),.dout(n6481),.clk(gclk));
	jor g06248(.dina(n6481),.dinb(w_n6357_49[1]),.dout(n6482),.clk(gclk));
	jxor g06249(.dina(n6482),.dinb(w_n6084_0[0]),.dout(n6483),.clk(gclk));
	jor g06250(.dina(w_n6483_0[2]),.dinb(n6480),.dout(n6484),.clk(gclk));
	jand g06251(.dina(n6484),.dinb(w_n6479_0[1]),.dout(n6485),.clk(gclk));
	jor g06252(.dina(w_n6485_0[2]),.dinb(w_n1699_49[2]),.dout(n6486),.clk(gclk));
	jand g06253(.dina(w_n6485_0[1]),.dinb(w_n1699_49[1]),.dout(n6487),.clk(gclk));
	jxor g06254(.dina(w_n6086_0[0]),.dinb(w_n1912_46[2]),.dout(n6488),.clk(gclk));
	jor g06255(.dina(n6488),.dinb(w_n6357_49[0]),.dout(n6489),.clk(gclk));
	jxor g06256(.dina(n6489),.dinb(w_n6092_0[0]),.dout(n6490),.clk(gclk));
	jor g06257(.dina(w_n6490_0[2]),.dinb(n6487),.dout(n6491),.clk(gclk));
	jand g06258(.dina(n6491),.dinb(w_n6486_0[1]),.dout(n6492),.clk(gclk));
	jor g06259(.dina(w_n6492_0[2]),.dinb(w_n1516_48[0]),.dout(n6493),.clk(gclk));
	jand g06260(.dina(w_n6492_0[1]),.dinb(w_n1516_47[2]),.dout(n6494),.clk(gclk));
	jxor g06261(.dina(w_n6094_0[0]),.dinb(w_n1699_49[0]),.dout(n6495),.clk(gclk));
	jor g06262(.dina(n6495),.dinb(w_n6357_48[2]),.dout(n6496),.clk(gclk));
	jxor g06263(.dina(n6496),.dinb(w_n6288_0[0]),.dout(n6497),.clk(gclk));
	jnot g06264(.din(w_n6497_0[2]),.dout(n6498),.clk(gclk));
	jor g06265(.dina(n6498),.dinb(n6494),.dout(n6499),.clk(gclk));
	jand g06266(.dina(n6499),.dinb(w_n6493_0[1]),.dout(n6500),.clk(gclk));
	jor g06267(.dina(w_n6500_0[2]),.dinb(w_n1332_49[2]),.dout(n6501),.clk(gclk));
	jand g06268(.dina(w_n6500_0[1]),.dinb(w_n1332_49[1]),.dout(n6502),.clk(gclk));
	jxor g06269(.dina(w_n6101_0[0]),.dinb(w_n1516_47[1]),.dout(n6503),.clk(gclk));
	jor g06270(.dina(n6503),.dinb(w_n6357_48[1]),.dout(n6504),.clk(gclk));
	jxor g06271(.dina(n6504),.dinb(w_n6107_0[0]),.dout(n6505),.clk(gclk));
	jor g06272(.dina(w_n6505_0[2]),.dinb(n6502),.dout(n6506),.clk(gclk));
	jand g06273(.dina(n6506),.dinb(w_n6501_0[1]),.dout(n6507),.clk(gclk));
	jor g06274(.dina(w_n6507_0[2]),.dinb(w_n1173_48[2]),.dout(n6508),.clk(gclk));
	jand g06275(.dina(w_n6507_0[1]),.dinb(w_n1173_48[1]),.dout(n6509),.clk(gclk));
	jxor g06276(.dina(w_n6109_0[0]),.dinb(w_n1332_49[0]),.dout(n6510),.clk(gclk));
	jor g06277(.dina(n6510),.dinb(w_n6357_48[0]),.dout(n6511),.clk(gclk));
	jxor g06278(.dina(n6511),.dinb(w_n6295_0[0]),.dout(n6512),.clk(gclk));
	jnot g06279(.din(w_n6512_0[2]),.dout(n6513),.clk(gclk));
	jor g06280(.dina(n6513),.dinb(n6509),.dout(n6514),.clk(gclk));
	jand g06281(.dina(n6514),.dinb(w_n6508_0[1]),.dout(n6515),.clk(gclk));
	jor g06282(.dina(w_n6515_0[2]),.dinb(w_n1008_50[2]),.dout(n6516),.clk(gclk));
	jand g06283(.dina(w_n6515_0[1]),.dinb(w_n1008_50[1]),.dout(n6517),.clk(gclk));
	jxor g06284(.dina(w_n6116_0[0]),.dinb(w_n1173_48[0]),.dout(n6518),.clk(gclk));
	jor g06285(.dina(n6518),.dinb(w_n6357_47[2]),.dout(n6519),.clk(gclk));
	jxor g06286(.dina(n6519),.dinb(w_n6122_0[0]),.dout(n6520),.clk(gclk));
	jor g06287(.dina(w_n6520_0[2]),.dinb(n6517),.dout(n6521),.clk(gclk));
	jand g06288(.dina(n6521),.dinb(w_n6516_0[1]),.dout(n6522),.clk(gclk));
	jor g06289(.dina(w_n6522_0[2]),.dinb(w_n884_49[2]),.dout(n6523),.clk(gclk));
	jand g06290(.dina(w_n6522_0[1]),.dinb(w_n884_49[1]),.dout(n6524),.clk(gclk));
	jxor g06291(.dina(w_n6124_0[0]),.dinb(w_n1008_50[0]),.dout(n6525),.clk(gclk));
	jor g06292(.dina(n6525),.dinb(w_n6357_47[1]),.dout(n6526),.clk(gclk));
	jxor g06293(.dina(n6526),.dinb(w_n6302_0[0]),.dout(n6527),.clk(gclk));
	jnot g06294(.din(w_n6527_0[2]),.dout(n6528),.clk(gclk));
	jor g06295(.dina(n6528),.dinb(n6524),.dout(n6529),.clk(gclk));
	jand g06296(.dina(n6529),.dinb(w_n6523_0[1]),.dout(n6530),.clk(gclk));
	jor g06297(.dina(w_n6530_0[2]),.dinb(w_n743_50[2]),.dout(n6531),.clk(gclk));
	jand g06298(.dina(w_n6530_0[1]),.dinb(w_n743_50[1]),.dout(n6532),.clk(gclk));
	jxor g06299(.dina(w_n6131_0[0]),.dinb(w_n884_49[0]),.dout(n6533),.clk(gclk));
	jor g06300(.dina(n6533),.dinb(w_n6357_47[0]),.dout(n6534),.clk(gclk));
	jxor g06301(.dina(n6534),.dinb(w_n6306_0[0]),.dout(n6535),.clk(gclk));
	jnot g06302(.din(w_n6535_0[2]),.dout(n6536),.clk(gclk));
	jor g06303(.dina(n6536),.dinb(n6532),.dout(n6537),.clk(gclk));
	jand g06304(.dina(n6537),.dinb(w_n6531_0[1]),.dout(n6538),.clk(gclk));
	jor g06305(.dina(w_n6538_0[2]),.dinb(w_n635_50[2]),.dout(n6539),.clk(gclk));
	jand g06306(.dina(w_n6538_0[1]),.dinb(w_n635_50[1]),.dout(n6540),.clk(gclk));
	jxor g06307(.dina(w_n6138_0[0]),.dinb(w_n743_50[0]),.dout(n6541),.clk(gclk));
	jor g06308(.dina(n6541),.dinb(w_n6357_46[2]),.dout(n6542),.clk(gclk));
	jxor g06309(.dina(n6542),.dinb(w_n6144_0[0]),.dout(n6543),.clk(gclk));
	jor g06310(.dina(w_n6543_0[2]),.dinb(n6540),.dout(n6544),.clk(gclk));
	jand g06311(.dina(n6544),.dinb(w_n6539_0[1]),.dout(n6545),.clk(gclk));
	jor g06312(.dina(w_n6545_0[2]),.dinb(w_n515_51[2]),.dout(n6546),.clk(gclk));
	jand g06313(.dina(w_n6545_0[1]),.dinb(w_n515_51[1]),.dout(n6547),.clk(gclk));
	jxor g06314(.dina(w_n6146_0[0]),.dinb(w_n635_50[0]),.dout(n6548),.clk(gclk));
	jor g06315(.dina(n6548),.dinb(w_n6357_46[1]),.dout(n6549),.clk(gclk));
	jxor g06316(.dina(n6549),.dinb(w_n6152_0[0]),.dout(n6550),.clk(gclk));
	jor g06317(.dina(w_n6550_0[2]),.dinb(n6547),.dout(n6551),.clk(gclk));
	jand g06318(.dina(n6551),.dinb(w_n6546_0[1]),.dout(n6552),.clk(gclk));
	jor g06319(.dina(w_n6552_0[2]),.dinb(w_n443_51[2]),.dout(n6553),.clk(gclk));
	jand g06320(.dina(w_n6552_0[1]),.dinb(w_n443_51[1]),.dout(n6554),.clk(gclk));
	jxor g06321(.dina(w_n6154_0[0]),.dinb(w_n515_51[0]),.dout(n6555),.clk(gclk));
	jor g06322(.dina(n6555),.dinb(w_n6357_46[0]),.dout(n6556),.clk(gclk));
	jxor g06323(.dina(n6556),.dinb(w_n6316_0[0]),.dout(n6557),.clk(gclk));
	jnot g06324(.din(w_n6557_0[1]),.dout(n6558),.clk(gclk));
	jor g06325(.dina(w_n6558_0[1]),.dinb(n6554),.dout(n6559),.clk(gclk));
	jand g06326(.dina(n6559),.dinb(w_n6553_0[1]),.dout(n6560),.clk(gclk));
	jor g06327(.dina(w_n6560_0[2]),.dinb(w_n352_52[0]),.dout(n6561),.clk(gclk));
	jand g06328(.dina(w_n6560_0[1]),.dinb(w_n352_51[2]),.dout(n6562),.clk(gclk));
	jxor g06329(.dina(w_n6161_0[0]),.dinb(w_n443_51[0]),.dout(n6563),.clk(gclk));
	jor g06330(.dina(n6563),.dinb(w_n6357_45[2]),.dout(n6564),.clk(gclk));
	jxor g06331(.dina(n6564),.dinb(w_n6166_0[0]),.dout(n6565),.clk(gclk));
	jnot g06332(.din(w_n6565_0[2]),.dout(n6566),.clk(gclk));
	jor g06333(.dina(n6566),.dinb(n6562),.dout(n6567),.clk(gclk));
	jand g06334(.dina(n6567),.dinb(w_n6561_0[1]),.dout(n6568),.clk(gclk));
	jor g06335(.dina(w_n6568_0[2]),.dinb(w_n294_52[1]),.dout(n6569),.clk(gclk));
	jand g06336(.dina(w_n6568_0[1]),.dinb(w_n294_52[0]),.dout(n6570),.clk(gclk));
	jxor g06337(.dina(w_n6169_0[0]),.dinb(w_n352_51[1]),.dout(n6571),.clk(gclk));
	jor g06338(.dina(n6571),.dinb(w_n6357_45[1]),.dout(n6572),.clk(gclk));
	jxor g06339(.dina(n6572),.dinb(w_n6323_0[0]),.dout(n6573),.clk(gclk));
	jnot g06340(.din(w_n6573_0[2]),.dout(n6574),.clk(gclk));
	jor g06341(.dina(n6574),.dinb(n6570),.dout(n6575),.clk(gclk));
	jand g06342(.dina(n6575),.dinb(w_n6569_0[1]),.dout(n6576),.clk(gclk));
	jor g06343(.dina(w_n6576_0[2]),.dinb(w_n239_52[1]),.dout(n6577),.clk(gclk));
	jand g06344(.dina(w_n6576_0[1]),.dinb(w_n239_52[0]),.dout(n6578),.clk(gclk));
	jxor g06345(.dina(w_n6176_0[0]),.dinb(w_n294_51[2]),.dout(n6579),.clk(gclk));
	jor g06346(.dina(n6579),.dinb(w_n6357_45[0]),.dout(n6580),.clk(gclk));
	jxor g06347(.dina(n6580),.dinb(w_n6182_0[0]),.dout(n6581),.clk(gclk));
	jor g06348(.dina(w_n6581_0[2]),.dinb(n6578),.dout(n6582),.clk(gclk));
	jand g06349(.dina(n6582),.dinb(w_n6577_0[1]),.dout(n6583),.clk(gclk));
	jor g06350(.dina(w_n6583_0[2]),.dinb(w_n221_52[1]),.dout(n6584),.clk(gclk));
	jand g06351(.dina(w_n6583_0[1]),.dinb(w_n221_52[0]),.dout(n6585),.clk(gclk));
	jxor g06352(.dina(w_n6184_0[0]),.dinb(w_n239_51[2]),.dout(n6586),.clk(gclk));
	jor g06353(.dina(n6586),.dinb(w_n6357_44[2]),.dout(n6587),.clk(gclk));
	jxor g06354(.dina(n6587),.dinb(w_n6190_0[0]),.dout(n6588),.clk(gclk));
	jor g06355(.dina(w_n6588_0[2]),.dinb(n6585),.dout(n6589),.clk(gclk));
	jand g06356(.dina(n6589),.dinb(w_n6584_0[1]),.dout(n6590),.clk(gclk));
	jor g06357(.dina(w_n6590_0[2]),.dinb(w_n6361_0[2]),.dout(n6591),.clk(gclk));
	jor g06358(.dina(w_n6591_0[1]),.dinb(w_n6202_0[0]),.dout(n6592),.clk(gclk));
	jor g06359(.dina(n6592),.dinb(w_n6349_0[1]),.dout(n6593),.clk(gclk));
	jand g06360(.dina(n6593),.dinb(w_n218_21[2]),.dout(n6594),.clk(gclk));
	jand g06361(.dina(w_n6357_44[1]),.dinb(w_n6204_0[0]),.dout(n6595),.clk(gclk));
	jand g06362(.dina(w_n6590_0[1]),.dinb(w_n6361_0[1]),.dout(n6596),.clk(gclk));
	jor g06363(.dina(w_n6596_0[2]),.dinb(n6595),.dout(n6597),.clk(gclk));
	jand g06364(.dina(w_n6355_0[0]),.dinb(w_n6334_0[0]),.dout(n6598),.clk(gclk));
	jand g06365(.dina(w_n6335_0[0]),.dinb(w_asqrt63_39[1]),.dout(n6599),.clk(gclk));
	jand g06366(.dina(n6599),.dinb(w_n6201_0[2]),.dout(n6600),.clk(gclk));
	jnot g06367(.din(n6600),.dout(n6601),.clk(gclk));
	jor g06368(.dina(w_n6601_0[1]),.dinb(n6598),.dout(n6602),.clk(gclk));
	jnot g06369(.din(n6602),.dout(n6603),.clk(gclk));
	jor g06370(.dina(n6603),.dinb(n6597),.dout(n6604),.clk(gclk));
	jor g06371(.dina(w_n6604_0[1]),.dinb(n6594),.dout(asqrt_fa_33),.clk(gclk));
	jnot g06372(.din(w_a62_0[2]),.dout(n6606),.clk(gclk));
	jnot g06373(.din(w_a63_0[1]),.dout(n6607),.clk(gclk));
	jand g06374(.dina(w_n6607_0[1]),.dinb(w_n6606_1[2]),.dout(n6608),.clk(gclk));
	jand g06375(.dina(w_n6608_0[2]),.dinb(w_n6362_1[1]),.dout(n6609),.clk(gclk));
	jand g06376(.dina(w_asqrt32_38[1]),.dinb(w_a64_0[1]),.dout(n6610),.clk(gclk));
	jor g06377(.dina(n6610),.dinb(w_n6609_0[1]),.dout(n6611),.clk(gclk));
	jand g06378(.dina(w_n6611_0[2]),.dinb(w_asqrt33_24[2]),.dout(n6612),.clk(gclk));
	jor g06379(.dina(w_n6611_0[1]),.dinb(w_asqrt33_24[1]),.dout(n6613),.clk(gclk));
	jand g06380(.dina(w_asqrt32_38[0]),.dinb(w_n6362_1[0]),.dout(n6614),.clk(gclk));
	jor g06381(.dina(n6614),.dinb(w_n6363_0[0]),.dout(n6615),.clk(gclk));
	jnot g06382(.din(w_n6364_0[1]),.dout(n6616),.clk(gclk));
	jnot g06383(.din(w_n6349_0[0]),.dout(n6617),.clk(gclk));
	jnot g06384(.din(w_n6584_0[0]),.dout(n6618),.clk(gclk));
	jnot g06385(.din(w_n6577_0[0]),.dout(n6619),.clk(gclk));
	jnot g06386(.din(w_n6569_0[0]),.dout(n6620),.clk(gclk));
	jnot g06387(.din(w_n6561_0[0]),.dout(n6621),.clk(gclk));
	jnot g06388(.din(w_n6553_0[0]),.dout(n6622),.clk(gclk));
	jnot g06389(.din(w_n6546_0[0]),.dout(n6623),.clk(gclk));
	jnot g06390(.din(w_n6539_0[0]),.dout(n6624),.clk(gclk));
	jnot g06391(.din(w_n6531_0[0]),.dout(n6625),.clk(gclk));
	jnot g06392(.din(w_n6523_0[0]),.dout(n6626),.clk(gclk));
	jnot g06393(.din(w_n6516_0[0]),.dout(n6627),.clk(gclk));
	jnot g06394(.din(w_n6508_0[0]),.dout(n6628),.clk(gclk));
	jnot g06395(.din(w_n6501_0[0]),.dout(n6629),.clk(gclk));
	jnot g06396(.din(w_n6493_0[0]),.dout(n6630),.clk(gclk));
	jnot g06397(.din(w_n6486_0[0]),.dout(n6631),.clk(gclk));
	jnot g06398(.din(w_n6479_0[0]),.dout(n6632),.clk(gclk));
	jnot g06399(.din(w_n6472_0[0]),.dout(n6633),.clk(gclk));
	jnot g06400(.din(w_n6464_0[0]),.dout(n6634),.clk(gclk));
	jnot g06401(.din(w_n6456_0[0]),.dout(n6635),.clk(gclk));
	jnot g06402(.din(w_n6448_0[0]),.dout(n6636),.clk(gclk));
	jnot g06403(.din(w_n6441_0[0]),.dout(n6637),.clk(gclk));
	jnot g06404(.din(w_n6433_0[0]),.dout(n6638),.clk(gclk));
	jnot g06405(.din(w_n6426_0[0]),.dout(n6639),.clk(gclk));
	jnot g06406(.din(w_n6418_0[0]),.dout(n6640),.clk(gclk));
	jnot g06407(.din(w_n6411_0[0]),.dout(n6641),.clk(gclk));
	jnot g06408(.din(w_n6403_0[0]),.dout(n6642),.clk(gclk));
	jnot g06409(.din(w_n6396_0[0]),.dout(n6643),.clk(gclk));
	jnot g06410(.din(w_n6388_0[0]),.dout(n6644),.clk(gclk));
	jnot g06411(.din(w_n6377_0[0]),.dout(n6645),.clk(gclk));
	jnot g06412(.din(w_n6369_0[0]),.dout(n6646),.clk(gclk));
	jand g06413(.dina(w_asqrt33_24[0]),.dinb(w_a66_0[2]),.dout(n6647),.clk(gclk));
	jor g06414(.dina(n6647),.dinb(w_n6365_0[0]),.dout(n6648),.clk(gclk));
	jor g06415(.dina(n6648),.dinb(w_asqrt34_28[2]),.dout(n6649),.clk(gclk));
	jand g06416(.dina(w_asqrt33_23[2]),.dinb(w_n5843_0[1]),.dout(n6650),.clk(gclk));
	jor g06417(.dina(n6650),.dinb(w_n5844_0[0]),.dout(n6651),.clk(gclk));
	jand g06418(.dina(w_n6380_0[0]),.dinb(n6651),.dout(n6652),.clk(gclk));
	jand g06419(.dina(w_n6652_0[1]),.dinb(n6649),.dout(n6653),.clk(gclk));
	jor g06420(.dina(n6653),.dinb(n6646),.dout(n6654),.clk(gclk));
	jor g06421(.dina(n6654),.dinb(w_asqrt35_24[2]),.dout(n6655),.clk(gclk));
	jnot g06422(.din(w_n6385_0[0]),.dout(n6656),.clk(gclk));
	jand g06423(.dina(w_n6656_0[1]),.dinb(n6655),.dout(n6657),.clk(gclk));
	jor g06424(.dina(n6657),.dinb(n6645),.dout(n6658),.clk(gclk));
	jor g06425(.dina(n6658),.dinb(w_asqrt36_28[2]),.dout(n6659),.clk(gclk));
	jand g06426(.dina(w_n6392_0[1]),.dinb(n6659),.dout(n6660),.clk(gclk));
	jor g06427(.dina(n6660),.dinb(n6644),.dout(n6661),.clk(gclk));
	jor g06428(.dina(n6661),.dinb(w_asqrt37_25[0]),.dout(n6662),.clk(gclk));
	jnot g06429(.din(w_n6400_0[1]),.dout(n6663),.clk(gclk));
	jand g06430(.dina(n6663),.dinb(n6662),.dout(n6664),.clk(gclk));
	jor g06431(.dina(n6664),.dinb(n6643),.dout(n6665),.clk(gclk));
	jor g06432(.dina(n6665),.dinb(w_asqrt38_29[0]),.dout(n6666),.clk(gclk));
	jand g06433(.dina(w_n6407_0[1]),.dinb(n6666),.dout(n6667),.clk(gclk));
	jor g06434(.dina(n6667),.dinb(n6642),.dout(n6668),.clk(gclk));
	jor g06435(.dina(n6668),.dinb(w_asqrt39_25[2]),.dout(n6669),.clk(gclk));
	jnot g06436(.din(w_n6415_0[1]),.dout(n6670),.clk(gclk));
	jand g06437(.dina(n6670),.dinb(n6669),.dout(n6671),.clk(gclk));
	jor g06438(.dina(n6671),.dinb(n6641),.dout(n6672),.clk(gclk));
	jor g06439(.dina(n6672),.dinb(w_asqrt40_29[0]),.dout(n6673),.clk(gclk));
	jand g06440(.dina(w_n6422_0[1]),.dinb(n6673),.dout(n6674),.clk(gclk));
	jor g06441(.dina(n6674),.dinb(n6640),.dout(n6675),.clk(gclk));
	jor g06442(.dina(n6675),.dinb(w_asqrt41_26[0]),.dout(n6676),.clk(gclk));
	jnot g06443(.din(w_n6430_0[1]),.dout(n6677),.clk(gclk));
	jand g06444(.dina(n6677),.dinb(n6676),.dout(n6678),.clk(gclk));
	jor g06445(.dina(n6678),.dinb(n6639),.dout(n6679),.clk(gclk));
	jor g06446(.dina(n6679),.dinb(w_asqrt42_29[1]),.dout(n6680),.clk(gclk));
	jand g06447(.dina(w_n6437_0[1]),.dinb(n6680),.dout(n6681),.clk(gclk));
	jor g06448(.dina(n6681),.dinb(n6638),.dout(n6682),.clk(gclk));
	jor g06449(.dina(n6682),.dinb(w_asqrt43_26[1]),.dout(n6683),.clk(gclk));
	jnot g06450(.din(w_n6445_0[1]),.dout(n6684),.clk(gclk));
	jand g06451(.dina(n6684),.dinb(n6683),.dout(n6685),.clk(gclk));
	jor g06452(.dina(n6685),.dinb(n6637),.dout(n6686),.clk(gclk));
	jor g06453(.dina(n6686),.dinb(w_asqrt44_29[1]),.dout(n6687),.clk(gclk));
	jand g06454(.dina(w_n6452_0[1]),.dinb(n6687),.dout(n6688),.clk(gclk));
	jor g06455(.dina(n6688),.dinb(n6636),.dout(n6689),.clk(gclk));
	jor g06456(.dina(n6689),.dinb(w_asqrt45_27[0]),.dout(n6690),.clk(gclk));
	jand g06457(.dina(w_n6460_0[1]),.dinb(n6690),.dout(n6691),.clk(gclk));
	jor g06458(.dina(n6691),.dinb(n6635),.dout(n6692),.clk(gclk));
	jor g06459(.dina(n6692),.dinb(w_asqrt46_29[1]),.dout(n6693),.clk(gclk));
	jand g06460(.dina(w_n6468_0[1]),.dinb(n6693),.dout(n6694),.clk(gclk));
	jor g06461(.dina(n6694),.dinb(n6634),.dout(n6695),.clk(gclk));
	jor g06462(.dina(n6695),.dinb(w_asqrt47_27[2]),.dout(n6696),.clk(gclk));
	jnot g06463(.din(w_n6476_0[1]),.dout(n6697),.clk(gclk));
	jand g06464(.dina(n6697),.dinb(n6696),.dout(n6698),.clk(gclk));
	jor g06465(.dina(n6698),.dinb(n6633),.dout(n6699),.clk(gclk));
	jor g06466(.dina(n6699),.dinb(w_asqrt48_29[2]),.dout(n6700),.clk(gclk));
	jnot g06467(.din(w_n6483_0[1]),.dout(n6701),.clk(gclk));
	jand g06468(.dina(n6701),.dinb(n6700),.dout(n6702),.clk(gclk));
	jor g06469(.dina(n6702),.dinb(n6632),.dout(n6703),.clk(gclk));
	jor g06470(.dina(n6703),.dinb(w_asqrt49_28[0]),.dout(n6704),.clk(gclk));
	jnot g06471(.din(w_n6490_0[1]),.dout(n6705),.clk(gclk));
	jand g06472(.dina(n6705),.dinb(n6704),.dout(n6706),.clk(gclk));
	jor g06473(.dina(n6706),.dinb(n6631),.dout(n6707),.clk(gclk));
	jor g06474(.dina(n6707),.dinb(w_asqrt50_30[0]),.dout(n6708),.clk(gclk));
	jand g06475(.dina(w_n6497_0[1]),.dinb(n6708),.dout(n6709),.clk(gclk));
	jor g06476(.dina(n6709),.dinb(n6630),.dout(n6710),.clk(gclk));
	jor g06477(.dina(n6710),.dinb(w_asqrt51_28[1]),.dout(n6711),.clk(gclk));
	jnot g06478(.din(w_n6505_0[1]),.dout(n6712),.clk(gclk));
	jand g06479(.dina(n6712),.dinb(n6711),.dout(n6713),.clk(gclk));
	jor g06480(.dina(n6713),.dinb(n6629),.dout(n6714),.clk(gclk));
	jor g06481(.dina(n6714),.dinb(w_asqrt52_30[0]),.dout(n6715),.clk(gclk));
	jand g06482(.dina(w_n6512_0[1]),.dinb(n6715),.dout(n6716),.clk(gclk));
	jor g06483(.dina(n6716),.dinb(n6628),.dout(n6717),.clk(gclk));
	jor g06484(.dina(n6717),.dinb(w_asqrt53_29[0]),.dout(n6718),.clk(gclk));
	jnot g06485(.din(w_n6520_0[1]),.dout(n6719),.clk(gclk));
	jand g06486(.dina(n6719),.dinb(n6718),.dout(n6720),.clk(gclk));
	jor g06487(.dina(n6720),.dinb(n6627),.dout(n6721),.clk(gclk));
	jor g06488(.dina(n6721),.dinb(w_asqrt54_30[0]),.dout(n6722),.clk(gclk));
	jand g06489(.dina(w_n6527_0[1]),.dinb(n6722),.dout(n6723),.clk(gclk));
	jor g06490(.dina(n6723),.dinb(n6626),.dout(n6724),.clk(gclk));
	jor g06491(.dina(n6724),.dinb(w_asqrt55_29[1]),.dout(n6725),.clk(gclk));
	jand g06492(.dina(w_n6535_0[1]),.dinb(n6725),.dout(n6726),.clk(gclk));
	jor g06493(.dina(n6726),.dinb(n6625),.dout(n6727),.clk(gclk));
	jor g06494(.dina(n6727),.dinb(w_asqrt56_30[1]),.dout(n6728),.clk(gclk));
	jnot g06495(.din(w_n6543_0[1]),.dout(n6729),.clk(gclk));
	jand g06496(.dina(n6729),.dinb(n6728),.dout(n6730),.clk(gclk));
	jor g06497(.dina(n6730),.dinb(n6624),.dout(n6731),.clk(gclk));
	jor g06498(.dina(n6731),.dinb(w_asqrt57_30[0]),.dout(n6732),.clk(gclk));
	jnot g06499(.din(w_n6550_0[1]),.dout(n6733),.clk(gclk));
	jand g06500(.dina(n6733),.dinb(n6732),.dout(n6734),.clk(gclk));
	jor g06501(.dina(n6734),.dinb(n6623),.dout(n6735),.clk(gclk));
	jor g06502(.dina(n6735),.dinb(w_asqrt58_30[2]),.dout(n6736),.clk(gclk));
	jand g06503(.dina(w_n6557_0[0]),.dinb(n6736),.dout(n6737),.clk(gclk));
	jor g06504(.dina(n6737),.dinb(n6622),.dout(n6738),.clk(gclk));
	jor g06505(.dina(n6738),.dinb(w_asqrt59_30[1]),.dout(n6739),.clk(gclk));
	jand g06506(.dina(w_n6565_0[1]),.dinb(n6739),.dout(n6740),.clk(gclk));
	jor g06507(.dina(n6740),.dinb(n6621),.dout(n6741),.clk(gclk));
	jor g06508(.dina(n6741),.dinb(w_asqrt60_30[2]),.dout(n6742),.clk(gclk));
	jand g06509(.dina(w_n6573_0[1]),.dinb(n6742),.dout(n6743),.clk(gclk));
	jor g06510(.dina(n6743),.dinb(n6620),.dout(n6744),.clk(gclk));
	jor g06511(.dina(n6744),.dinb(w_asqrt61_30[2]),.dout(n6745),.clk(gclk));
	jnot g06512(.din(w_n6581_0[1]),.dout(n6746),.clk(gclk));
	jand g06513(.dina(n6746),.dinb(n6745),.dout(n6747),.clk(gclk));
	jor g06514(.dina(n6747),.dinb(n6619),.dout(n6748),.clk(gclk));
	jor g06515(.dina(n6748),.dinb(w_asqrt62_30[2]),.dout(n6749),.clk(gclk));
	jnot g06516(.din(w_n6588_0[1]),.dout(n6750),.clk(gclk));
	jand g06517(.dina(n6750),.dinb(n6749),.dout(n6751),.clk(gclk));
	jor g06518(.dina(n6751),.dinb(n6618),.dout(n6752),.clk(gclk));
	jand g06519(.dina(n6752),.dinb(w_n6360_0[0]),.dout(n6753),.clk(gclk));
	jand g06520(.dina(w_n6753_0[1]),.dinb(w_n6201_0[1]),.dout(n6754),.clk(gclk));
	jand g06521(.dina(n6754),.dinb(n6617),.dout(n6755),.clk(gclk));
	jor g06522(.dina(n6755),.dinb(w_asqrt63_39[0]),.dout(n6756),.clk(gclk));
	jnot g06523(.din(w_n6604_0[0]),.dout(n6757),.clk(gclk));
	jand g06524(.dina(n6757),.dinb(w_n6756_0[1]),.dout(n6758),.clk(gclk));
	jor g06525(.dina(w_n6758_40[2]),.dinb(n6616),.dout(n6759),.clk(gclk));
	jand g06526(.dina(n6759),.dinb(n6615),.dout(n6760),.clk(gclk));
	jand g06527(.dina(n6760),.dinb(n6613),.dout(n6761),.clk(gclk));
	jor g06528(.dina(n6761),.dinb(w_n6612_0[1]),.dout(n6762),.clk(gclk));
	jand g06529(.dina(w_n6762_0[2]),.dinb(w_asqrt34_28[1]),.dout(n6763),.clk(gclk));
	jor g06530(.dina(w_n6762_0[1]),.dinb(w_asqrt34_28[0]),.dout(n6764),.clk(gclk));
	jand g06531(.dina(w_asqrt32_37[2]),.dinb(w_n6364_0[0]),.dout(n6765),.clk(gclk));
	jnot g06532(.din(w_n6596_0[1]),.dout(n6766),.clk(gclk));
	jand g06533(.dina(w_n6601_0[0]),.dinb(w_asqrt33_23[1]),.dout(n6767),.clk(gclk));
	jand g06534(.dina(n6767),.dinb(w_n6766_0[1]),.dout(n6768),.clk(gclk));
	jand g06535(.dina(n6768),.dinb(w_n6756_0[0]),.dout(n6769),.clk(gclk));
	jor g06536(.dina(n6769),.dinb(w_n6765_0[1]),.dout(n6770),.clk(gclk));
	jxor g06537(.dina(n6770),.dinb(w_a66_0[1]),.dout(n6771),.clk(gclk));
	jnot g06538(.din(w_n6771_0[1]),.dout(n6772),.clk(gclk));
	jand g06539(.dina(w_n6772_0[1]),.dinb(n6764),.dout(n6773),.clk(gclk));
	jor g06540(.dina(n6773),.dinb(w_n6763_0[1]),.dout(n6774),.clk(gclk));
	jand g06541(.dina(w_n6774_0[2]),.dinb(w_asqrt35_24[1]),.dout(n6775),.clk(gclk));
	jor g06542(.dina(w_n6774_0[1]),.dinb(w_asqrt35_24[0]),.dout(n6776),.clk(gclk));
	jxor g06543(.dina(w_n6368_0[0]),.dinb(w_n5989_40[1]),.dout(n6777),.clk(gclk));
	jand g06544(.dina(n6777),.dinb(w_asqrt32_37[1]),.dout(n6778),.clk(gclk));
	jxor g06545(.dina(n6778),.dinb(w_n6652_0[0]),.dout(n6779),.clk(gclk));
	jand g06546(.dina(w_n6779_0[1]),.dinb(n6776),.dout(n6780),.clk(gclk));
	jor g06547(.dina(n6780),.dinb(w_n6775_0[1]),.dout(n6781),.clk(gclk));
	jand g06548(.dina(w_n6781_0[2]),.dinb(w_asqrt36_28[1]),.dout(n6782),.clk(gclk));
	jor g06549(.dina(w_n6781_0[1]),.dinb(w_asqrt36_28[0]),.dout(n6783),.clk(gclk));
	jxor g06550(.dina(w_n6376_0[0]),.dinb(w_n5606_44[2]),.dout(n6784),.clk(gclk));
	jand g06551(.dina(n6784),.dinb(w_asqrt32_37[0]),.dout(n6785),.clk(gclk));
	jxor g06552(.dina(n6785),.dinb(w_n6656_0[0]),.dout(n6786),.clk(gclk));
	jand g06553(.dina(w_n6786_0[1]),.dinb(n6783),.dout(n6787),.clk(gclk));
	jor g06554(.dina(n6787),.dinb(w_n6782_0[1]),.dout(n6788),.clk(gclk));
	jand g06555(.dina(w_n6788_0[2]),.dinb(w_asqrt37_24[2]),.dout(n6789),.clk(gclk));
	jor g06556(.dina(w_n6788_0[1]),.dinb(w_asqrt37_24[1]),.dout(n6790),.clk(gclk));
	jxor g06557(.dina(w_n6387_0[0]),.dinb(w_n5259_41[1]),.dout(n6791),.clk(gclk));
	jand g06558(.dina(n6791),.dinb(w_asqrt32_36[2]),.dout(n6792),.clk(gclk));
	jxor g06559(.dina(n6792),.dinb(w_n6392_0[0]),.dout(n6793),.clk(gclk));
	jand g06560(.dina(w_n6793_0[1]),.dinb(n6790),.dout(n6794),.clk(gclk));
	jor g06561(.dina(n6794),.dinb(w_n6789_0[1]),.dout(n6795),.clk(gclk));
	jand g06562(.dina(w_n6795_0[2]),.dinb(w_asqrt38_28[2]),.dout(n6796),.clk(gclk));
	jor g06563(.dina(w_n6795_0[1]),.dinb(w_asqrt38_28[1]),.dout(n6797),.clk(gclk));
	jxor g06564(.dina(w_n6395_0[0]),.dinb(w_n4902_45[1]),.dout(n6798),.clk(gclk));
	jand g06565(.dina(n6798),.dinb(w_asqrt32_36[1]),.dout(n6799),.clk(gclk));
	jxor g06566(.dina(n6799),.dinb(w_n6400_0[0]),.dout(n6800),.clk(gclk));
	jnot g06567(.din(w_n6800_0[1]),.dout(n6801),.clk(gclk));
	jand g06568(.dina(w_n6801_0[1]),.dinb(n6797),.dout(n6802),.clk(gclk));
	jor g06569(.dina(n6802),.dinb(w_n6796_0[1]),.dout(n6803),.clk(gclk));
	jand g06570(.dina(w_n6803_0[2]),.dinb(w_asqrt39_25[1]),.dout(n6804),.clk(gclk));
	jor g06571(.dina(w_n6803_0[1]),.dinb(w_asqrt39_25[0]),.dout(n6805),.clk(gclk));
	jxor g06572(.dina(w_n6402_0[0]),.dinb(w_n4582_42[1]),.dout(n6806),.clk(gclk));
	jand g06573(.dina(n6806),.dinb(w_asqrt32_36[0]),.dout(n6807),.clk(gclk));
	jxor g06574(.dina(n6807),.dinb(w_n6407_0[0]),.dout(n6808),.clk(gclk));
	jand g06575(.dina(w_n6808_0[1]),.dinb(n6805),.dout(n6809),.clk(gclk));
	jor g06576(.dina(n6809),.dinb(w_n6804_0[1]),.dout(n6810),.clk(gclk));
	jand g06577(.dina(w_n6810_0[2]),.dinb(w_asqrt40_28[2]),.dout(n6811),.clk(gclk));
	jor g06578(.dina(w_n6810_0[1]),.dinb(w_asqrt40_28[1]),.dout(n6812),.clk(gclk));
	jxor g06579(.dina(w_n6410_0[0]),.dinb(w_n4249_46[0]),.dout(n6813),.clk(gclk));
	jand g06580(.dina(n6813),.dinb(w_asqrt32_35[2]),.dout(n6814),.clk(gclk));
	jxor g06581(.dina(n6814),.dinb(w_n6415_0[0]),.dout(n6815),.clk(gclk));
	jnot g06582(.din(w_n6815_0[1]),.dout(n6816),.clk(gclk));
	jand g06583(.dina(w_n6816_0[1]),.dinb(n6812),.dout(n6817),.clk(gclk));
	jor g06584(.dina(n6817),.dinb(w_n6811_0[1]),.dout(n6818),.clk(gclk));
	jand g06585(.dina(w_n6818_0[2]),.dinb(w_asqrt41_25[2]),.dout(n6819),.clk(gclk));
	jor g06586(.dina(w_n6818_0[1]),.dinb(w_asqrt41_25[1]),.dout(n6820),.clk(gclk));
	jxor g06587(.dina(w_n6417_0[0]),.dinb(w_n3955_43[0]),.dout(n6821),.clk(gclk));
	jand g06588(.dina(n6821),.dinb(w_asqrt32_35[1]),.dout(n6822),.clk(gclk));
	jxor g06589(.dina(n6822),.dinb(w_n6422_0[0]),.dout(n6823),.clk(gclk));
	jand g06590(.dina(w_n6823_0[1]),.dinb(n6820),.dout(n6824),.clk(gclk));
	jor g06591(.dina(n6824),.dinb(w_n6819_0[1]),.dout(n6825),.clk(gclk));
	jand g06592(.dina(w_n6825_0[2]),.dinb(w_asqrt42_29[0]),.dout(n6826),.clk(gclk));
	jor g06593(.dina(w_n6825_0[1]),.dinb(w_asqrt42_28[2]),.dout(n6827),.clk(gclk));
	jxor g06594(.dina(w_n6425_0[0]),.dinb(w_n3642_46[1]),.dout(n6828),.clk(gclk));
	jand g06595(.dina(n6828),.dinb(w_asqrt32_35[0]),.dout(n6829),.clk(gclk));
	jxor g06596(.dina(n6829),.dinb(w_n6430_0[0]),.dout(n6830),.clk(gclk));
	jnot g06597(.din(w_n6830_0[1]),.dout(n6831),.clk(gclk));
	jand g06598(.dina(w_n6831_0[1]),.dinb(n6827),.dout(n6832),.clk(gclk));
	jor g06599(.dina(n6832),.dinb(w_n6826_0[1]),.dout(n6833),.clk(gclk));
	jand g06600(.dina(w_n6833_0[2]),.dinb(w_asqrt43_26[0]),.dout(n6834),.clk(gclk));
	jor g06601(.dina(w_n6833_0[1]),.dinb(w_asqrt43_25[2]),.dout(n6835),.clk(gclk));
	jxor g06602(.dina(w_n6432_0[0]),.dinb(w_n3368_43[2]),.dout(n6836),.clk(gclk));
	jand g06603(.dina(n6836),.dinb(w_asqrt32_34[2]),.dout(n6837),.clk(gclk));
	jxor g06604(.dina(n6837),.dinb(w_n6437_0[0]),.dout(n6838),.clk(gclk));
	jand g06605(.dina(w_n6838_0[1]),.dinb(n6835),.dout(n6839),.clk(gclk));
	jor g06606(.dina(n6839),.dinb(w_n6834_0[1]),.dout(n6840),.clk(gclk));
	jand g06607(.dina(w_n6840_0[2]),.dinb(w_asqrt44_29[0]),.dout(n6841),.clk(gclk));
	jor g06608(.dina(w_n6840_0[1]),.dinb(w_asqrt44_28[2]),.dout(n6842),.clk(gclk));
	jxor g06609(.dina(w_n6440_0[0]),.dinb(w_n3089_47[0]),.dout(n6843),.clk(gclk));
	jand g06610(.dina(n6843),.dinb(w_asqrt32_34[1]),.dout(n6844),.clk(gclk));
	jxor g06611(.dina(n6844),.dinb(w_n6445_0[0]),.dout(n6845),.clk(gclk));
	jnot g06612(.din(w_n6845_0[1]),.dout(n6846),.clk(gclk));
	jand g06613(.dina(w_n6846_0[1]),.dinb(n6842),.dout(n6847),.clk(gclk));
	jor g06614(.dina(n6847),.dinb(w_n6841_0[1]),.dout(n6848),.clk(gclk));
	jand g06615(.dina(w_n6848_0[2]),.dinb(w_asqrt45_26[2]),.dout(n6849),.clk(gclk));
	jor g06616(.dina(w_n6848_0[1]),.dinb(w_asqrt45_26[1]),.dout(n6850),.clk(gclk));
	jxor g06617(.dina(w_n6447_0[0]),.dinb(w_n2833_44[2]),.dout(n6851),.clk(gclk));
	jand g06618(.dina(n6851),.dinb(w_asqrt32_34[0]),.dout(n6852),.clk(gclk));
	jxor g06619(.dina(n6852),.dinb(w_n6452_0[0]),.dout(n6853),.clk(gclk));
	jand g06620(.dina(w_n6853_0[1]),.dinb(n6850),.dout(n6854),.clk(gclk));
	jor g06621(.dina(n6854),.dinb(w_n6849_0[1]),.dout(n6855),.clk(gclk));
	jand g06622(.dina(w_n6855_0[2]),.dinb(w_asqrt46_29[0]),.dout(n6856),.clk(gclk));
	jor g06623(.dina(w_n6855_0[1]),.dinb(w_asqrt46_28[2]),.dout(n6857),.clk(gclk));
	jxor g06624(.dina(w_n6455_0[0]),.dinb(w_n2572_47[1]),.dout(n6858),.clk(gclk));
	jand g06625(.dina(n6858),.dinb(w_asqrt32_33[2]),.dout(n6859),.clk(gclk));
	jxor g06626(.dina(n6859),.dinb(w_n6460_0[0]),.dout(n6860),.clk(gclk));
	jand g06627(.dina(w_n6860_0[1]),.dinb(n6857),.dout(n6861),.clk(gclk));
	jor g06628(.dina(n6861),.dinb(w_n6856_0[1]),.dout(n6862),.clk(gclk));
	jand g06629(.dina(w_n6862_0[2]),.dinb(w_asqrt47_27[1]),.dout(n6863),.clk(gclk));
	jor g06630(.dina(w_n6862_0[1]),.dinb(w_asqrt47_27[0]),.dout(n6864),.clk(gclk));
	jxor g06631(.dina(w_n6463_0[0]),.dinb(w_n2345_45[1]),.dout(n6865),.clk(gclk));
	jand g06632(.dina(n6865),.dinb(w_asqrt32_33[1]),.dout(n6866),.clk(gclk));
	jxor g06633(.dina(n6866),.dinb(w_n6468_0[0]),.dout(n6867),.clk(gclk));
	jand g06634(.dina(w_n6867_0[1]),.dinb(n6864),.dout(n6868),.clk(gclk));
	jor g06635(.dina(n6868),.dinb(w_n6863_0[1]),.dout(n6869),.clk(gclk));
	jand g06636(.dina(w_n6869_0[2]),.dinb(w_asqrt48_29[1]),.dout(n6870),.clk(gclk));
	jor g06637(.dina(w_n6869_0[1]),.dinb(w_asqrt48_29[0]),.dout(n6871),.clk(gclk));
	jxor g06638(.dina(w_n6471_0[0]),.dinb(w_n2108_48[0]),.dout(n6872),.clk(gclk));
	jand g06639(.dina(n6872),.dinb(w_asqrt32_33[0]),.dout(n6873),.clk(gclk));
	jxor g06640(.dina(n6873),.dinb(w_n6476_0[0]),.dout(n6874),.clk(gclk));
	jnot g06641(.din(w_n6874_0[1]),.dout(n6875),.clk(gclk));
	jand g06642(.dina(w_n6875_0[1]),.dinb(n6871),.dout(n6876),.clk(gclk));
	jor g06643(.dina(n6876),.dinb(w_n6870_0[1]),.dout(n6877),.clk(gclk));
	jand g06644(.dina(w_n6877_0[2]),.dinb(w_asqrt49_27[2]),.dout(n6878),.clk(gclk));
	jor g06645(.dina(w_n6877_0[1]),.dinb(w_asqrt49_27[1]),.dout(n6879),.clk(gclk));
	jxor g06646(.dina(w_n6478_0[0]),.dinb(w_n1912_46[1]),.dout(n6880),.clk(gclk));
	jand g06647(.dina(n6880),.dinb(w_asqrt32_32[2]),.dout(n6881),.clk(gclk));
	jxor g06648(.dina(n6881),.dinb(w_n6483_0[0]),.dout(n6882),.clk(gclk));
	jnot g06649(.din(w_n6882_0[1]),.dout(n6883),.clk(gclk));
	jand g06650(.dina(w_n6883_0[1]),.dinb(n6879),.dout(n6884),.clk(gclk));
	jor g06651(.dina(n6884),.dinb(w_n6878_0[1]),.dout(n6885),.clk(gclk));
	jand g06652(.dina(w_n6885_0[2]),.dinb(w_asqrt50_29[2]),.dout(n6886),.clk(gclk));
	jor g06653(.dina(w_n6885_0[1]),.dinb(w_asqrt50_29[1]),.dout(n6887),.clk(gclk));
	jxor g06654(.dina(w_n6485_0[0]),.dinb(w_n1699_48[2]),.dout(n6888),.clk(gclk));
	jand g06655(.dina(n6888),.dinb(w_asqrt32_32[1]),.dout(n6889),.clk(gclk));
	jxor g06656(.dina(n6889),.dinb(w_n6490_0[0]),.dout(n6890),.clk(gclk));
	jnot g06657(.din(w_n6890_0[1]),.dout(n6891),.clk(gclk));
	jand g06658(.dina(w_n6891_0[1]),.dinb(n6887),.dout(n6892),.clk(gclk));
	jor g06659(.dina(n6892),.dinb(w_n6886_0[1]),.dout(n6893),.clk(gclk));
	jand g06660(.dina(w_n6893_0[2]),.dinb(w_asqrt51_28[0]),.dout(n6894),.clk(gclk));
	jor g06661(.dina(w_n6893_0[1]),.dinb(w_asqrt51_27[2]),.dout(n6895),.clk(gclk));
	jxor g06662(.dina(w_n6492_0[0]),.dinb(w_n1516_47[0]),.dout(n6896),.clk(gclk));
	jand g06663(.dina(n6896),.dinb(w_asqrt32_32[0]),.dout(n6897),.clk(gclk));
	jxor g06664(.dina(n6897),.dinb(w_n6497_0[0]),.dout(n6898),.clk(gclk));
	jand g06665(.dina(w_n6898_0[1]),.dinb(n6895),.dout(n6899),.clk(gclk));
	jor g06666(.dina(n6899),.dinb(w_n6894_0[1]),.dout(n6900),.clk(gclk));
	jand g06667(.dina(w_n6900_0[2]),.dinb(w_asqrt52_29[2]),.dout(n6901),.clk(gclk));
	jor g06668(.dina(w_n6900_0[1]),.dinb(w_asqrt52_29[1]),.dout(n6902),.clk(gclk));
	jxor g06669(.dina(w_n6500_0[0]),.dinb(w_n1332_48[2]),.dout(n6903),.clk(gclk));
	jand g06670(.dina(n6903),.dinb(w_asqrt32_31[2]),.dout(n6904),.clk(gclk));
	jxor g06671(.dina(n6904),.dinb(w_n6505_0[0]),.dout(n6905),.clk(gclk));
	jnot g06672(.din(w_n6905_0[1]),.dout(n6906),.clk(gclk));
	jand g06673(.dina(w_n6906_0[1]),.dinb(n6902),.dout(n6907),.clk(gclk));
	jor g06674(.dina(n6907),.dinb(w_n6901_0[1]),.dout(n6908),.clk(gclk));
	jand g06675(.dina(w_n6908_0[2]),.dinb(w_asqrt53_28[2]),.dout(n6909),.clk(gclk));
	jor g06676(.dina(w_n6908_0[1]),.dinb(w_asqrt53_28[1]),.dout(n6910),.clk(gclk));
	jxor g06677(.dina(w_n6507_0[0]),.dinb(w_n1173_47[2]),.dout(n6911),.clk(gclk));
	jand g06678(.dina(n6911),.dinb(w_asqrt32_31[1]),.dout(n6912),.clk(gclk));
	jxor g06679(.dina(n6912),.dinb(w_n6512_0[0]),.dout(n6913),.clk(gclk));
	jand g06680(.dina(w_n6913_0[1]),.dinb(n6910),.dout(n6914),.clk(gclk));
	jor g06681(.dina(n6914),.dinb(w_n6909_0[1]),.dout(n6915),.clk(gclk));
	jand g06682(.dina(w_n6915_0[2]),.dinb(w_asqrt54_29[2]),.dout(n6916),.clk(gclk));
	jor g06683(.dina(w_n6915_0[1]),.dinb(w_asqrt54_29[1]),.dout(n6917),.clk(gclk));
	jxor g06684(.dina(w_n6515_0[0]),.dinb(w_n1008_49[2]),.dout(n6918),.clk(gclk));
	jand g06685(.dina(n6918),.dinb(w_asqrt32_31[0]),.dout(n6919),.clk(gclk));
	jxor g06686(.dina(n6919),.dinb(w_n6520_0[0]),.dout(n6920),.clk(gclk));
	jnot g06687(.din(w_n6920_0[1]),.dout(n6921),.clk(gclk));
	jand g06688(.dina(w_n6921_0[1]),.dinb(n6917),.dout(n6922),.clk(gclk));
	jor g06689(.dina(n6922),.dinb(w_n6916_0[1]),.dout(n6923),.clk(gclk));
	jand g06690(.dina(w_n6923_0[2]),.dinb(w_asqrt55_29[0]),.dout(n6924),.clk(gclk));
	jor g06691(.dina(w_n6923_0[1]),.dinb(w_asqrt55_28[2]),.dout(n6925),.clk(gclk));
	jxor g06692(.dina(w_n6522_0[0]),.dinb(w_n884_48[2]),.dout(n6926),.clk(gclk));
	jand g06693(.dina(n6926),.dinb(w_asqrt32_30[2]),.dout(n6927),.clk(gclk));
	jxor g06694(.dina(n6927),.dinb(w_n6527_0[0]),.dout(n6928),.clk(gclk));
	jand g06695(.dina(w_n6928_0[1]),.dinb(n6925),.dout(n6929),.clk(gclk));
	jor g06696(.dina(n6929),.dinb(w_n6924_0[1]),.dout(n6930),.clk(gclk));
	jand g06697(.dina(w_n6930_0[2]),.dinb(w_asqrt56_30[0]),.dout(n6931),.clk(gclk));
	jor g06698(.dina(w_n6930_0[1]),.dinb(w_asqrt56_29[2]),.dout(n6932),.clk(gclk));
	jxor g06699(.dina(w_n6530_0[0]),.dinb(w_n743_49[2]),.dout(n6933),.clk(gclk));
	jand g06700(.dina(n6933),.dinb(w_asqrt32_30[1]),.dout(n6934),.clk(gclk));
	jxor g06701(.dina(n6934),.dinb(w_n6535_0[0]),.dout(n6935),.clk(gclk));
	jand g06702(.dina(w_n6935_0[1]),.dinb(n6932),.dout(n6936),.clk(gclk));
	jor g06703(.dina(n6936),.dinb(w_n6931_0[1]),.dout(n6937),.clk(gclk));
	jand g06704(.dina(w_n6937_0[2]),.dinb(w_asqrt57_29[2]),.dout(n6938),.clk(gclk));
	jor g06705(.dina(w_n6937_0[1]),.dinb(w_asqrt57_29[1]),.dout(n6939),.clk(gclk));
	jxor g06706(.dina(w_n6538_0[0]),.dinb(w_n635_49[2]),.dout(n6940),.clk(gclk));
	jand g06707(.dina(n6940),.dinb(w_asqrt32_30[0]),.dout(n6941),.clk(gclk));
	jxor g06708(.dina(n6941),.dinb(w_n6543_0[0]),.dout(n6942),.clk(gclk));
	jnot g06709(.din(w_n6942_0[1]),.dout(n6943),.clk(gclk));
	jand g06710(.dina(w_n6943_0[1]),.dinb(n6939),.dout(n6944),.clk(gclk));
	jor g06711(.dina(n6944),.dinb(w_n6938_0[1]),.dout(n6945),.clk(gclk));
	jand g06712(.dina(w_n6945_0[2]),.dinb(w_asqrt58_30[1]),.dout(n6946),.clk(gclk));
	jor g06713(.dina(w_n6945_0[1]),.dinb(w_asqrt58_30[0]),.dout(n6947),.clk(gclk));
	jxor g06714(.dina(w_n6545_0[0]),.dinb(w_n515_50[2]),.dout(n6948),.clk(gclk));
	jand g06715(.dina(n6948),.dinb(w_asqrt32_29[2]),.dout(n6949),.clk(gclk));
	jxor g06716(.dina(n6949),.dinb(w_n6550_0[0]),.dout(n6950),.clk(gclk));
	jnot g06717(.din(w_n6950_0[1]),.dout(n6951),.clk(gclk));
	jand g06718(.dina(w_n6951_0[1]),.dinb(n6947),.dout(n6952),.clk(gclk));
	jor g06719(.dina(n6952),.dinb(w_n6946_0[1]),.dout(n6953),.clk(gclk));
	jand g06720(.dina(w_n6953_0[2]),.dinb(w_asqrt59_30[0]),.dout(n6954),.clk(gclk));
	jor g06721(.dina(w_n6953_0[1]),.dinb(w_asqrt59_29[2]),.dout(n6955),.clk(gclk));
	jxor g06722(.dina(w_n6552_0[0]),.dinb(w_n443_50[2]),.dout(n6956),.clk(gclk));
	jand g06723(.dina(n6956),.dinb(w_asqrt32_29[1]),.dout(n6957),.clk(gclk));
	jxor g06724(.dina(n6957),.dinb(w_n6558_0[0]),.dout(n6958),.clk(gclk));
	jnot g06725(.din(w_n6958_0[1]),.dout(n6959),.clk(gclk));
	jand g06726(.dina(w_n6959_0[1]),.dinb(n6955),.dout(n6960),.clk(gclk));
	jor g06727(.dina(n6960),.dinb(w_n6954_0[1]),.dout(n6961),.clk(gclk));
	jand g06728(.dina(w_n6961_0[2]),.dinb(w_asqrt60_30[1]),.dout(n6962),.clk(gclk));
	jor g06729(.dina(w_n6961_0[1]),.dinb(w_asqrt60_30[0]),.dout(n6963),.clk(gclk));
	jxor g06730(.dina(w_n6560_0[0]),.dinb(w_n352_51[0]),.dout(n6964),.clk(gclk));
	jand g06731(.dina(n6964),.dinb(w_asqrt32_29[0]),.dout(n6965),.clk(gclk));
	jxor g06732(.dina(n6965),.dinb(w_n6565_0[0]),.dout(n6966),.clk(gclk));
	jand g06733(.dina(w_n6966_0[1]),.dinb(n6963),.dout(n6967),.clk(gclk));
	jor g06734(.dina(n6967),.dinb(w_n6962_0[1]),.dout(n6968),.clk(gclk));
	jand g06735(.dina(w_n6968_0[2]),.dinb(w_asqrt61_30[1]),.dout(n6969),.clk(gclk));
	jor g06736(.dina(w_n6968_0[1]),.dinb(w_asqrt61_30[0]),.dout(n6970),.clk(gclk));
	jxor g06737(.dina(w_n6568_0[0]),.dinb(w_n294_51[1]),.dout(n6971),.clk(gclk));
	jand g06738(.dina(n6971),.dinb(w_asqrt32_28[2]),.dout(n6972),.clk(gclk));
	jxor g06739(.dina(n6972),.dinb(w_n6573_0[0]),.dout(n6973),.clk(gclk));
	jand g06740(.dina(w_n6973_0[1]),.dinb(n6970),.dout(n6974),.clk(gclk));
	jor g06741(.dina(n6974),.dinb(w_n6969_0[1]),.dout(n6975),.clk(gclk));
	jand g06742(.dina(w_n6975_0[2]),.dinb(w_asqrt62_30[1]),.dout(n6976),.clk(gclk));
	jor g06743(.dina(w_n6975_0[1]),.dinb(w_asqrt62_30[0]),.dout(n6977),.clk(gclk));
	jxor g06744(.dina(w_n6576_0[0]),.dinb(w_n239_51[1]),.dout(n6978),.clk(gclk));
	jand g06745(.dina(n6978),.dinb(w_asqrt32_28[1]),.dout(n6979),.clk(gclk));
	jxor g06746(.dina(n6979),.dinb(w_n6581_0[0]),.dout(n6980),.clk(gclk));
	jnot g06747(.din(w_n6980_0[1]),.dout(n6981),.clk(gclk));
	jand g06748(.dina(w_n6981_0[1]),.dinb(n6977),.dout(n6982),.clk(gclk));
	jor g06749(.dina(n6982),.dinb(w_n6976_0[1]),.dout(n6983),.clk(gclk));
	jxor g06750(.dina(w_n6583_0[0]),.dinb(w_n221_51[2]),.dout(n6984),.clk(gclk));
	jand g06751(.dina(n6984),.dinb(w_asqrt32_28[0]),.dout(n6985),.clk(gclk));
	jxor g06752(.dina(n6985),.dinb(w_n6588_0[0]),.dout(n6986),.clk(gclk));
	jnot g06753(.din(w_n6986_0[2]),.dout(n6987),.clk(gclk));
	jor g06754(.dina(w_n6987_0[1]),.dinb(w_n6983_0[1]),.dout(n6988),.clk(gclk));
	jnot g06755(.din(w_n6988_1[1]),.dout(n6989),.clk(gclk));
	jand g06756(.dina(w_n6758_40[1]),.dinb(w_n6590_0[0]),.dout(n6990),.clk(gclk));
	jnot g06757(.din(n6990),.dout(n6991),.clk(gclk));
	jand g06758(.dina(w_n6591_0[0]),.dinb(w_asqrt63_38[2]),.dout(n6992),.clk(gclk));
	jand g06759(.dina(n6992),.dinb(w_n6766_0[0]),.dout(n6993),.clk(gclk));
	jand g06760(.dina(w_n6993_0[1]),.dinb(n6991),.dout(n6994),.clk(gclk));
	jnot g06761(.din(w_n6976_0[0]),.dout(n6995),.clk(gclk));
	jnot g06762(.din(w_n6969_0[0]),.dout(n6996),.clk(gclk));
	jnot g06763(.din(w_n6962_0[0]),.dout(n6997),.clk(gclk));
	jnot g06764(.din(w_n6954_0[0]),.dout(n6998),.clk(gclk));
	jnot g06765(.din(w_n6946_0[0]),.dout(n6999),.clk(gclk));
	jnot g06766(.din(w_n6938_0[0]),.dout(n7000),.clk(gclk));
	jnot g06767(.din(w_n6931_0[0]),.dout(n7001),.clk(gclk));
	jnot g06768(.din(w_n6924_0[0]),.dout(n7002),.clk(gclk));
	jnot g06769(.din(w_n6916_0[0]),.dout(n7003),.clk(gclk));
	jnot g06770(.din(w_n6909_0[0]),.dout(n7004),.clk(gclk));
	jnot g06771(.din(w_n6901_0[0]),.dout(n7005),.clk(gclk));
	jnot g06772(.din(w_n6894_0[0]),.dout(n7006),.clk(gclk));
	jnot g06773(.din(w_n6886_0[0]),.dout(n7007),.clk(gclk));
	jnot g06774(.din(w_n6878_0[0]),.dout(n7008),.clk(gclk));
	jnot g06775(.din(w_n6870_0[0]),.dout(n7009),.clk(gclk));
	jnot g06776(.din(w_n6863_0[0]),.dout(n7010),.clk(gclk));
	jnot g06777(.din(w_n6856_0[0]),.dout(n7011),.clk(gclk));
	jnot g06778(.din(w_n6849_0[0]),.dout(n7012),.clk(gclk));
	jnot g06779(.din(w_n6841_0[0]),.dout(n7013),.clk(gclk));
	jnot g06780(.din(w_n6834_0[0]),.dout(n7014),.clk(gclk));
	jnot g06781(.din(w_n6826_0[0]),.dout(n7015),.clk(gclk));
	jnot g06782(.din(w_n6819_0[0]),.dout(n7016),.clk(gclk));
	jnot g06783(.din(w_n6811_0[0]),.dout(n7017),.clk(gclk));
	jnot g06784(.din(w_n6804_0[0]),.dout(n7018),.clk(gclk));
	jnot g06785(.din(w_n6796_0[0]),.dout(n7019),.clk(gclk));
	jnot g06786(.din(w_n6789_0[0]),.dout(n7020),.clk(gclk));
	jnot g06787(.din(w_n6782_0[0]),.dout(n7021),.clk(gclk));
	jnot g06788(.din(w_n6775_0[0]),.dout(n7022),.clk(gclk));
	jnot g06789(.din(w_n6763_0[0]),.dout(n7023),.clk(gclk));
	jnot g06790(.din(w_n6612_0[0]),.dout(n7024),.clk(gclk));
	jnot g06791(.din(w_n6609_0[0]),.dout(n7025),.clk(gclk));
	jor g06792(.dina(w_n6758_40[0]),.dinb(w_n6362_0[2]),.dout(n7026),.clk(gclk));
	jand g06793(.dina(n7026),.dinb(n7025),.dout(n7027),.clk(gclk));
	jand g06794(.dina(n7027),.dinb(w_n6357_44[0]),.dout(n7028),.clk(gclk));
	jor g06795(.dina(w_n6758_39[2]),.dinb(w_a64_0[0]),.dout(n7029),.clk(gclk));
	jand g06796(.dina(n7029),.dinb(w_a65_0[0]),.dout(n7030),.clk(gclk));
	jor g06797(.dina(w_n6765_0[0]),.dinb(n7030),.dout(n7031),.clk(gclk));
	jor g06798(.dina(w_n7031_0[1]),.dinb(n7028),.dout(n7032),.clk(gclk));
	jand g06799(.dina(n7032),.dinb(n7024),.dout(n7033),.clk(gclk));
	jand g06800(.dina(n7033),.dinb(w_n5989_40[0]),.dout(n7034),.clk(gclk));
	jor g06801(.dina(w_n6771_0[0]),.dinb(n7034),.dout(n7035),.clk(gclk));
	jand g06802(.dina(n7035),.dinb(n7023),.dout(n7036),.clk(gclk));
	jand g06803(.dina(n7036),.dinb(w_n5606_44[1]),.dout(n7037),.clk(gclk));
	jnot g06804(.din(w_n6779_0[0]),.dout(n7038),.clk(gclk));
	jor g06805(.dina(w_n7038_0[1]),.dinb(n7037),.dout(n7039),.clk(gclk));
	jand g06806(.dina(n7039),.dinb(n7022),.dout(n7040),.clk(gclk));
	jand g06807(.dina(n7040),.dinb(w_n5259_41[0]),.dout(n7041),.clk(gclk));
	jnot g06808(.din(w_n6786_0[0]),.dout(n7042),.clk(gclk));
	jor g06809(.dina(w_n7042_0[1]),.dinb(n7041),.dout(n7043),.clk(gclk));
	jand g06810(.dina(n7043),.dinb(n7021),.dout(n7044),.clk(gclk));
	jand g06811(.dina(n7044),.dinb(w_n4902_45[0]),.dout(n7045),.clk(gclk));
	jnot g06812(.din(w_n6793_0[0]),.dout(n7046),.clk(gclk));
	jor g06813(.dina(w_n7046_0[1]),.dinb(n7045),.dout(n7047),.clk(gclk));
	jand g06814(.dina(n7047),.dinb(n7020),.dout(n7048),.clk(gclk));
	jand g06815(.dina(n7048),.dinb(w_n4582_42[0]),.dout(n7049),.clk(gclk));
	jor g06816(.dina(w_n6800_0[0]),.dinb(n7049),.dout(n7050),.clk(gclk));
	jand g06817(.dina(n7050),.dinb(n7019),.dout(n7051),.clk(gclk));
	jand g06818(.dina(n7051),.dinb(w_n4249_45[2]),.dout(n7052),.clk(gclk));
	jnot g06819(.din(w_n6808_0[0]),.dout(n7053),.clk(gclk));
	jor g06820(.dina(w_n7053_0[1]),.dinb(n7052),.dout(n7054),.clk(gclk));
	jand g06821(.dina(n7054),.dinb(n7018),.dout(n7055),.clk(gclk));
	jand g06822(.dina(n7055),.dinb(w_n3955_42[2]),.dout(n7056),.clk(gclk));
	jor g06823(.dina(w_n6815_0[0]),.dinb(n7056),.dout(n7057),.clk(gclk));
	jand g06824(.dina(n7057),.dinb(n7017),.dout(n7058),.clk(gclk));
	jand g06825(.dina(n7058),.dinb(w_n3642_46[0]),.dout(n7059),.clk(gclk));
	jnot g06826(.din(w_n6823_0[0]),.dout(n7060),.clk(gclk));
	jor g06827(.dina(w_n7060_0[1]),.dinb(n7059),.dout(n7061),.clk(gclk));
	jand g06828(.dina(n7061),.dinb(n7016),.dout(n7062),.clk(gclk));
	jand g06829(.dina(n7062),.dinb(w_n3368_43[1]),.dout(n7063),.clk(gclk));
	jor g06830(.dina(w_n6830_0[0]),.dinb(n7063),.dout(n7064),.clk(gclk));
	jand g06831(.dina(n7064),.dinb(n7015),.dout(n7065),.clk(gclk));
	jand g06832(.dina(n7065),.dinb(w_n3089_46[2]),.dout(n7066),.clk(gclk));
	jnot g06833(.din(w_n6838_0[0]),.dout(n7067),.clk(gclk));
	jor g06834(.dina(w_n7067_0[1]),.dinb(n7066),.dout(n7068),.clk(gclk));
	jand g06835(.dina(n7068),.dinb(n7014),.dout(n7069),.clk(gclk));
	jand g06836(.dina(n7069),.dinb(w_n2833_44[1]),.dout(n7070),.clk(gclk));
	jor g06837(.dina(w_n6845_0[0]),.dinb(n7070),.dout(n7071),.clk(gclk));
	jand g06838(.dina(n7071),.dinb(n7013),.dout(n7072),.clk(gclk));
	jand g06839(.dina(n7072),.dinb(w_n2572_47[0]),.dout(n7073),.clk(gclk));
	jnot g06840(.din(w_n6853_0[0]),.dout(n7074),.clk(gclk));
	jor g06841(.dina(w_n7074_0[1]),.dinb(n7073),.dout(n7075),.clk(gclk));
	jand g06842(.dina(n7075),.dinb(n7012),.dout(n7076),.clk(gclk));
	jand g06843(.dina(n7076),.dinb(w_n2345_45[0]),.dout(n7077),.clk(gclk));
	jnot g06844(.din(w_n6860_0[0]),.dout(n7078),.clk(gclk));
	jor g06845(.dina(w_n7078_0[1]),.dinb(n7077),.dout(n7079),.clk(gclk));
	jand g06846(.dina(n7079),.dinb(n7011),.dout(n7080),.clk(gclk));
	jand g06847(.dina(n7080),.dinb(w_n2108_47[2]),.dout(n7081),.clk(gclk));
	jnot g06848(.din(w_n6867_0[0]),.dout(n7082),.clk(gclk));
	jor g06849(.dina(w_n7082_0[1]),.dinb(n7081),.dout(n7083),.clk(gclk));
	jand g06850(.dina(n7083),.dinb(n7010),.dout(n7084),.clk(gclk));
	jand g06851(.dina(n7084),.dinb(w_n1912_46[0]),.dout(n7085),.clk(gclk));
	jor g06852(.dina(w_n6874_0[0]),.dinb(n7085),.dout(n7086),.clk(gclk));
	jand g06853(.dina(n7086),.dinb(n7009),.dout(n7087),.clk(gclk));
	jand g06854(.dina(n7087),.dinb(w_n1699_48[1]),.dout(n7088),.clk(gclk));
	jor g06855(.dina(w_n6882_0[0]),.dinb(n7088),.dout(n7089),.clk(gclk));
	jand g06856(.dina(n7089),.dinb(n7008),.dout(n7090),.clk(gclk));
	jand g06857(.dina(n7090),.dinb(w_n1516_46[2]),.dout(n7091),.clk(gclk));
	jor g06858(.dina(w_n6890_0[0]),.dinb(n7091),.dout(n7092),.clk(gclk));
	jand g06859(.dina(n7092),.dinb(n7007),.dout(n7093),.clk(gclk));
	jand g06860(.dina(n7093),.dinb(w_n1332_48[1]),.dout(n7094),.clk(gclk));
	jnot g06861(.din(w_n6898_0[0]),.dout(n7095),.clk(gclk));
	jor g06862(.dina(w_n7095_0[1]),.dinb(n7094),.dout(n7096),.clk(gclk));
	jand g06863(.dina(n7096),.dinb(n7006),.dout(n7097),.clk(gclk));
	jand g06864(.dina(n7097),.dinb(w_n1173_47[1]),.dout(n7098),.clk(gclk));
	jor g06865(.dina(w_n6905_0[0]),.dinb(n7098),.dout(n7099),.clk(gclk));
	jand g06866(.dina(n7099),.dinb(n7005),.dout(n7100),.clk(gclk));
	jand g06867(.dina(n7100),.dinb(w_n1008_49[1]),.dout(n7101),.clk(gclk));
	jnot g06868(.din(w_n6913_0[0]),.dout(n7102),.clk(gclk));
	jor g06869(.dina(w_n7102_0[1]),.dinb(n7101),.dout(n7103),.clk(gclk));
	jand g06870(.dina(n7103),.dinb(n7004),.dout(n7104),.clk(gclk));
	jand g06871(.dina(n7104),.dinb(w_n884_48[1]),.dout(n7105),.clk(gclk));
	jor g06872(.dina(w_n6920_0[0]),.dinb(n7105),.dout(n7106),.clk(gclk));
	jand g06873(.dina(n7106),.dinb(n7003),.dout(n7107),.clk(gclk));
	jand g06874(.dina(n7107),.dinb(w_n743_49[1]),.dout(n7108),.clk(gclk));
	jnot g06875(.din(w_n6928_0[0]),.dout(n7109),.clk(gclk));
	jor g06876(.dina(w_n7109_0[1]),.dinb(n7108),.dout(n7110),.clk(gclk));
	jand g06877(.dina(n7110),.dinb(n7002),.dout(n7111),.clk(gclk));
	jand g06878(.dina(n7111),.dinb(w_n635_49[1]),.dout(n7112),.clk(gclk));
	jnot g06879(.din(w_n6935_0[0]),.dout(n7113),.clk(gclk));
	jor g06880(.dina(w_n7113_0[1]),.dinb(n7112),.dout(n7114),.clk(gclk));
	jand g06881(.dina(n7114),.dinb(n7001),.dout(n7115),.clk(gclk));
	jand g06882(.dina(n7115),.dinb(w_n515_50[1]),.dout(n7116),.clk(gclk));
	jor g06883(.dina(w_n6942_0[0]),.dinb(n7116),.dout(n7117),.clk(gclk));
	jand g06884(.dina(n7117),.dinb(n7000),.dout(n7118),.clk(gclk));
	jand g06885(.dina(n7118),.dinb(w_n443_50[1]),.dout(n7119),.clk(gclk));
	jor g06886(.dina(w_n6950_0[0]),.dinb(n7119),.dout(n7120),.clk(gclk));
	jand g06887(.dina(n7120),.dinb(n6999),.dout(n7121),.clk(gclk));
	jand g06888(.dina(n7121),.dinb(w_n352_50[2]),.dout(n7122),.clk(gclk));
	jor g06889(.dina(w_n6958_0[0]),.dinb(n7122),.dout(n7123),.clk(gclk));
	jand g06890(.dina(n7123),.dinb(n6998),.dout(n7124),.clk(gclk));
	jand g06891(.dina(n7124),.dinb(w_n294_51[0]),.dout(n7125),.clk(gclk));
	jnot g06892(.din(w_n6966_0[0]),.dout(n7126),.clk(gclk));
	jor g06893(.dina(w_n7126_0[1]),.dinb(n7125),.dout(n7127),.clk(gclk));
	jand g06894(.dina(n7127),.dinb(n6997),.dout(n7128),.clk(gclk));
	jand g06895(.dina(n7128),.dinb(w_n239_51[0]),.dout(n7129),.clk(gclk));
	jnot g06896(.din(w_n6973_0[0]),.dout(n7130),.clk(gclk));
	jor g06897(.dina(w_n7130_0[1]),.dinb(n7129),.dout(n7131),.clk(gclk));
	jand g06898(.dina(n7131),.dinb(n6996),.dout(n7132),.clk(gclk));
	jand g06899(.dina(n7132),.dinb(w_n221_51[1]),.dout(n7133),.clk(gclk));
	jor g06900(.dina(w_n6980_0[0]),.dinb(n7133),.dout(n7134),.clk(gclk));
	jand g06901(.dina(n7134),.dinb(n6995),.dout(n7135),.clk(gclk));
	jor g06902(.dina(w_n6986_0[1]),.dinb(w_n7135_0[1]),.dout(n7136),.clk(gclk));
	jand g06903(.dina(w_asqrt32_27[2]),.dinb(w_n6753_0[0]),.dout(n7137),.clk(gclk));
	jor g06904(.dina(n7137),.dinb(w_n6596_0[0]),.dout(n7138),.clk(gclk));
	jor g06905(.dina(w_n7138_0[1]),.dinb(w_n7136_0[1]),.dout(n7139),.clk(gclk));
	jand g06906(.dina(n7139),.dinb(w_n218_21[1]),.dout(n7140),.clk(gclk));
	jand g06907(.dina(w_n6758_39[1]),.dinb(w_n6361_0[0]),.dout(n7141),.clk(gclk));
	jor g06908(.dina(w_n7141_0[1]),.dinb(w_n7140_0[1]),.dout(n7142),.clk(gclk));
	jor g06909(.dina(n7142),.dinb(w_n6994_0[1]),.dout(n7143),.clk(gclk));
	jor g06910(.dina(w_n7143_0[1]),.dinb(w_n6989_0[2]),.dout(asqrt_fa_32),.clk(gclk));
	jand g06911(.dina(w_n6987_0[0]),.dinb(w_n6983_0[0]),.dout(n7145),.clk(gclk));
	jand g06912(.dina(w_n7143_0[0]),.dinb(w_n7145_0[1]),.dout(n7146),.clk(gclk));
	jnot g06913(.din(w_n6994_0[0]),.dout(n7147),.clk(gclk));
	jnot g06914(.din(w_n7138_0[0]),.dout(n7148),.clk(gclk));
	jand g06915(.dina(n7148),.dinb(w_n7145_0[0]),.dout(n7149),.clk(gclk));
	jor g06916(.dina(n7149),.dinb(w_asqrt63_38[1]),.dout(n7150),.clk(gclk));
	jnot g06917(.din(w_n7141_0[0]),.dout(n7151),.clk(gclk));
	jand g06918(.dina(n7151),.dinb(n7150),.dout(n7152),.clk(gclk));
	jand g06919(.dina(n7152),.dinb(n7147),.dout(n7153),.clk(gclk));
	jand g06920(.dina(w_n7153_0[1]),.dinb(w_n6988_1[0]),.dout(n7154),.clk(gclk));
	jor g06921(.dina(w_n7154_53[2]),.dinb(w_n6606_1[1]),.dout(n7155),.clk(gclk));
	jnot g06922(.din(w_a60_0[2]),.dout(n7156),.clk(gclk));
	jnot g06923(.din(w_a61_0[1]),.dout(n7157),.clk(gclk));
	jand g06924(.dina(w_n7157_0[1]),.dinb(w_n7156_1[2]),.dout(n7158),.clk(gclk));
	jand g06925(.dina(w_n7158_0[2]),.dinb(w_n6606_1[0]),.dout(n7159),.clk(gclk));
	jnot g06926(.din(w_n7159_0[1]),.dout(n7160),.clk(gclk));
	jand g06927(.dina(n7160),.dinb(n7155),.dout(n7161),.clk(gclk));
	jor g06928(.dina(w_n7161_0[2]),.dinb(w_n6758_39[0]),.dout(n7162),.clk(gclk));
	jand g06929(.dina(w_asqrt31_23),.dinb(w_n6608_0[1]),.dout(n7163),.clk(gclk));
	jor g06930(.dina(w_n7154_53[1]),.dinb(w_a62_0[1]),.dout(n7164),.clk(gclk));
	jand g06931(.dina(n7164),.dinb(w_a63_0[0]),.dout(n7165),.clk(gclk));
	jor g06932(.dina(n7165),.dinb(n7163),.dout(n7166),.clk(gclk));
	jand g06933(.dina(w_n7161_0[1]),.dinb(w_n6758_38[2]),.dout(n7167),.clk(gclk));
	jor g06934(.dina(n7167),.dinb(n7166),.dout(n7168),.clk(gclk));
	jand g06935(.dina(n7168),.dinb(w_n7162_0[1]),.dout(n7169),.clk(gclk));
	jor g06936(.dina(w_n7169_0[2]),.dinb(w_n6357_43[2]),.dout(n7170),.clk(gclk));
	jand g06937(.dina(w_n7169_0[1]),.dinb(w_n6357_43[1]),.dout(n7171),.clk(gclk));
	jnot g06938(.din(w_n6608_0[0]),.dout(n7172),.clk(gclk));
	jor g06939(.dina(w_n7154_53[0]),.dinb(n7172),.dout(n7173),.clk(gclk));
	jor g06940(.dina(w_n6989_0[1]),.dinb(w_n6758_38[1]),.dout(n7174),.clk(gclk));
	jor g06941(.dina(n7174),.dinb(w_n6993_0[0]),.dout(n7175),.clk(gclk));
	jor g06942(.dina(n7175),.dinb(w_n7140_0[0]),.dout(n7176),.clk(gclk));
	jand g06943(.dina(n7176),.dinb(w_n7173_0[1]),.dout(n7177),.clk(gclk));
	jxor g06944(.dina(n7177),.dinb(w_n6362_0[1]),.dout(n7178),.clk(gclk));
	jor g06945(.dina(w_n7178_0[2]),.dinb(n7171),.dout(n7179),.clk(gclk));
	jand g06946(.dina(n7179),.dinb(w_n7170_0[1]),.dout(n7180),.clk(gclk));
	jor g06947(.dina(w_n7180_0[2]),.dinb(w_n5989_39[2]),.dout(n7181),.clk(gclk));
	jand g06948(.dina(w_n7180_0[1]),.dinb(w_n5989_39[1]),.dout(n7182),.clk(gclk));
	jxor g06949(.dina(w_n6611_0[0]),.dinb(w_n6357_43[0]),.dout(n7183),.clk(gclk));
	jor g06950(.dina(n7183),.dinb(w_n7154_52[2]),.dout(n7184),.clk(gclk));
	jxor g06951(.dina(n7184),.dinb(w_n7031_0[0]),.dout(n7185),.clk(gclk));
	jnot g06952(.din(w_n7185_0[2]),.dout(n7186),.clk(gclk));
	jor g06953(.dina(n7186),.dinb(n7182),.dout(n7187),.clk(gclk));
	jand g06954(.dina(n7187),.dinb(w_n7181_0[1]),.dout(n7188),.clk(gclk));
	jor g06955(.dina(w_n7188_0[2]),.dinb(w_n5606_44[0]),.dout(n7189),.clk(gclk));
	jand g06956(.dina(w_n7188_0[1]),.dinb(w_n5606_43[2]),.dout(n7190),.clk(gclk));
	jxor g06957(.dina(w_n6762_0[0]),.dinb(w_n5989_39[0]),.dout(n7191),.clk(gclk));
	jor g06958(.dina(n7191),.dinb(w_n7154_52[1]),.dout(n7192),.clk(gclk));
	jxor g06959(.dina(n7192),.dinb(w_n6772_0[0]),.dout(n7193),.clk(gclk));
	jor g06960(.dina(w_n7193_0[2]),.dinb(n7190),.dout(n7194),.clk(gclk));
	jand g06961(.dina(n7194),.dinb(w_n7189_0[1]),.dout(n7195),.clk(gclk));
	jor g06962(.dina(w_n7195_0[2]),.dinb(w_n5259_40[2]),.dout(n7196),.clk(gclk));
	jand g06963(.dina(w_n7195_0[1]),.dinb(w_n5259_40[1]),.dout(n7197),.clk(gclk));
	jxor g06964(.dina(w_n6774_0[0]),.dinb(w_n5606_43[1]),.dout(n7198),.clk(gclk));
	jor g06965(.dina(n7198),.dinb(w_n7154_52[0]),.dout(n7199),.clk(gclk));
	jxor g06966(.dina(n7199),.dinb(w_n7038_0[0]),.dout(n7200),.clk(gclk));
	jnot g06967(.din(w_n7200_0[2]),.dout(n7201),.clk(gclk));
	jor g06968(.dina(n7201),.dinb(n7197),.dout(n7202),.clk(gclk));
	jand g06969(.dina(n7202),.dinb(w_n7196_0[1]),.dout(n7203),.clk(gclk));
	jor g06970(.dina(w_n7203_0[2]),.dinb(w_n4902_44[2]),.dout(n7204),.clk(gclk));
	jand g06971(.dina(w_n7203_0[1]),.dinb(w_n4902_44[1]),.dout(n7205),.clk(gclk));
	jxor g06972(.dina(w_n6781_0[0]),.dinb(w_n5259_40[0]),.dout(n7206),.clk(gclk));
	jor g06973(.dina(n7206),.dinb(w_n7154_51[2]),.dout(n7207),.clk(gclk));
	jxor g06974(.dina(n7207),.dinb(w_n7042_0[0]),.dout(n7208),.clk(gclk));
	jnot g06975(.din(w_n7208_0[2]),.dout(n7209),.clk(gclk));
	jor g06976(.dina(n7209),.dinb(n7205),.dout(n7210),.clk(gclk));
	jand g06977(.dina(n7210),.dinb(w_n7204_0[1]),.dout(n7211),.clk(gclk));
	jor g06978(.dina(w_n7211_0[2]),.dinb(w_n4582_41[2]),.dout(n7212),.clk(gclk));
	jand g06979(.dina(w_n7211_0[1]),.dinb(w_n4582_41[1]),.dout(n7213),.clk(gclk));
	jxor g06980(.dina(w_n6788_0[0]),.dinb(w_n4902_44[0]),.dout(n7214),.clk(gclk));
	jor g06981(.dina(n7214),.dinb(w_n7154_51[1]),.dout(n7215),.clk(gclk));
	jxor g06982(.dina(n7215),.dinb(w_n7046_0[0]),.dout(n7216),.clk(gclk));
	jnot g06983(.din(w_n7216_0[2]),.dout(n7217),.clk(gclk));
	jor g06984(.dina(n7217),.dinb(n7213),.dout(n7218),.clk(gclk));
	jand g06985(.dina(n7218),.dinb(w_n7212_0[1]),.dout(n7219),.clk(gclk));
	jor g06986(.dina(w_n7219_0[2]),.dinb(w_n4249_45[1]),.dout(n7220),.clk(gclk));
	jand g06987(.dina(w_n7219_0[1]),.dinb(w_n4249_45[0]),.dout(n7221),.clk(gclk));
	jxor g06988(.dina(w_n6795_0[0]),.dinb(w_n4582_41[0]),.dout(n7222),.clk(gclk));
	jor g06989(.dina(n7222),.dinb(w_n7154_51[0]),.dout(n7223),.clk(gclk));
	jxor g06990(.dina(n7223),.dinb(w_n6801_0[0]),.dout(n7224),.clk(gclk));
	jor g06991(.dina(w_n7224_0[2]),.dinb(n7221),.dout(n7225),.clk(gclk));
	jand g06992(.dina(n7225),.dinb(w_n7220_0[1]),.dout(n7226),.clk(gclk));
	jor g06993(.dina(w_n7226_0[2]),.dinb(w_n3955_42[1]),.dout(n7227),.clk(gclk));
	jand g06994(.dina(w_n7226_0[1]),.dinb(w_n3955_42[0]),.dout(n7228),.clk(gclk));
	jxor g06995(.dina(w_n6803_0[0]),.dinb(w_n4249_44[2]),.dout(n7229),.clk(gclk));
	jor g06996(.dina(n7229),.dinb(w_n7154_50[2]),.dout(n7230),.clk(gclk));
	jxor g06997(.dina(n7230),.dinb(w_n7053_0[0]),.dout(n7231),.clk(gclk));
	jnot g06998(.din(w_n7231_0[2]),.dout(n7232),.clk(gclk));
	jor g06999(.dina(n7232),.dinb(n7228),.dout(n7233),.clk(gclk));
	jand g07000(.dina(n7233),.dinb(w_n7227_0[1]),.dout(n7234),.clk(gclk));
	jor g07001(.dina(w_n7234_0[2]),.dinb(w_n3642_45[2]),.dout(n7235),.clk(gclk));
	jand g07002(.dina(w_n7234_0[1]),.dinb(w_n3642_45[1]),.dout(n7236),.clk(gclk));
	jxor g07003(.dina(w_n6810_0[0]),.dinb(w_n3955_41[2]),.dout(n7237),.clk(gclk));
	jor g07004(.dina(n7237),.dinb(w_n7154_50[1]),.dout(n7238),.clk(gclk));
	jxor g07005(.dina(n7238),.dinb(w_n6816_0[0]),.dout(n7239),.clk(gclk));
	jor g07006(.dina(w_n7239_0[2]),.dinb(n7236),.dout(n7240),.clk(gclk));
	jand g07007(.dina(n7240),.dinb(w_n7235_0[1]),.dout(n7241),.clk(gclk));
	jor g07008(.dina(w_n7241_0[2]),.dinb(w_n3368_43[0]),.dout(n7242),.clk(gclk));
	jand g07009(.dina(w_n7241_0[1]),.dinb(w_n3368_42[2]),.dout(n7243),.clk(gclk));
	jxor g07010(.dina(w_n6818_0[0]),.dinb(w_n3642_45[0]),.dout(n7244),.clk(gclk));
	jor g07011(.dina(n7244),.dinb(w_n7154_50[0]),.dout(n7245),.clk(gclk));
	jxor g07012(.dina(n7245),.dinb(w_n7060_0[0]),.dout(n7246),.clk(gclk));
	jnot g07013(.din(w_n7246_0[2]),.dout(n7247),.clk(gclk));
	jor g07014(.dina(n7247),.dinb(n7243),.dout(n7248),.clk(gclk));
	jand g07015(.dina(n7248),.dinb(w_n7242_0[1]),.dout(n7249),.clk(gclk));
	jor g07016(.dina(w_n7249_0[2]),.dinb(w_n3089_46[1]),.dout(n7250),.clk(gclk));
	jand g07017(.dina(w_n7249_0[1]),.dinb(w_n3089_46[0]),.dout(n7251),.clk(gclk));
	jxor g07018(.dina(w_n6825_0[0]),.dinb(w_n3368_42[1]),.dout(n7252),.clk(gclk));
	jor g07019(.dina(n7252),.dinb(w_n7154_49[2]),.dout(n7253),.clk(gclk));
	jxor g07020(.dina(n7253),.dinb(w_n6831_0[0]),.dout(n7254),.clk(gclk));
	jor g07021(.dina(w_n7254_0[2]),.dinb(n7251),.dout(n7255),.clk(gclk));
	jand g07022(.dina(n7255),.dinb(w_n7250_0[1]),.dout(n7256),.clk(gclk));
	jor g07023(.dina(w_n7256_0[2]),.dinb(w_n2833_44[0]),.dout(n7257),.clk(gclk));
	jand g07024(.dina(w_n7256_0[1]),.dinb(w_n2833_43[2]),.dout(n7258),.clk(gclk));
	jxor g07025(.dina(w_n6833_0[0]),.dinb(w_n3089_45[2]),.dout(n7259),.clk(gclk));
	jor g07026(.dina(n7259),.dinb(w_n7154_49[1]),.dout(n7260),.clk(gclk));
	jxor g07027(.dina(n7260),.dinb(w_n7067_0[0]),.dout(n7261),.clk(gclk));
	jnot g07028(.din(w_n7261_0[2]),.dout(n7262),.clk(gclk));
	jor g07029(.dina(n7262),.dinb(n7258),.dout(n7263),.clk(gclk));
	jand g07030(.dina(n7263),.dinb(w_n7257_0[1]),.dout(n7264),.clk(gclk));
	jor g07031(.dina(w_n7264_0[2]),.dinb(w_n2572_46[2]),.dout(n7265),.clk(gclk));
	jand g07032(.dina(w_n7264_0[1]),.dinb(w_n2572_46[1]),.dout(n7266),.clk(gclk));
	jxor g07033(.dina(w_n6840_0[0]),.dinb(w_n2833_43[1]),.dout(n7267),.clk(gclk));
	jor g07034(.dina(n7267),.dinb(w_n7154_49[0]),.dout(n7268),.clk(gclk));
	jxor g07035(.dina(n7268),.dinb(w_n6846_0[0]),.dout(n7269),.clk(gclk));
	jor g07036(.dina(w_n7269_0[2]),.dinb(n7266),.dout(n7270),.clk(gclk));
	jand g07037(.dina(n7270),.dinb(w_n7265_0[1]),.dout(n7271),.clk(gclk));
	jor g07038(.dina(w_n7271_0[2]),.dinb(w_n2345_44[2]),.dout(n7272),.clk(gclk));
	jand g07039(.dina(w_n7271_0[1]),.dinb(w_n2345_44[1]),.dout(n7273),.clk(gclk));
	jxor g07040(.dina(w_n6848_0[0]),.dinb(w_n2572_46[0]),.dout(n7274),.clk(gclk));
	jor g07041(.dina(n7274),.dinb(w_n7154_48[2]),.dout(n7275),.clk(gclk));
	jxor g07042(.dina(n7275),.dinb(w_n7074_0[0]),.dout(n7276),.clk(gclk));
	jnot g07043(.din(w_n7276_0[2]),.dout(n7277),.clk(gclk));
	jor g07044(.dina(n7277),.dinb(n7273),.dout(n7278),.clk(gclk));
	jand g07045(.dina(n7278),.dinb(w_n7272_0[1]),.dout(n7279),.clk(gclk));
	jor g07046(.dina(w_n7279_0[2]),.dinb(w_n2108_47[1]),.dout(n7280),.clk(gclk));
	jand g07047(.dina(w_n7279_0[1]),.dinb(w_n2108_47[0]),.dout(n7281),.clk(gclk));
	jxor g07048(.dina(w_n6855_0[0]),.dinb(w_n2345_44[0]),.dout(n7282),.clk(gclk));
	jor g07049(.dina(n7282),.dinb(w_n7154_48[1]),.dout(n7283),.clk(gclk));
	jxor g07050(.dina(n7283),.dinb(w_n7078_0[0]),.dout(n7284),.clk(gclk));
	jnot g07051(.din(w_n7284_0[2]),.dout(n7285),.clk(gclk));
	jor g07052(.dina(n7285),.dinb(n7281),.dout(n7286),.clk(gclk));
	jand g07053(.dina(n7286),.dinb(w_n7280_0[1]),.dout(n7287),.clk(gclk));
	jor g07054(.dina(w_n7287_0[2]),.dinb(w_n1912_45[2]),.dout(n7288),.clk(gclk));
	jand g07055(.dina(w_n7287_0[1]),.dinb(w_n1912_45[1]),.dout(n7289),.clk(gclk));
	jxor g07056(.dina(w_n6862_0[0]),.dinb(w_n2108_46[2]),.dout(n7290),.clk(gclk));
	jor g07057(.dina(n7290),.dinb(w_n7154_48[0]),.dout(n7291),.clk(gclk));
	jxor g07058(.dina(n7291),.dinb(w_n7082_0[0]),.dout(n7292),.clk(gclk));
	jnot g07059(.din(w_n7292_0[2]),.dout(n7293),.clk(gclk));
	jor g07060(.dina(n7293),.dinb(n7289),.dout(n7294),.clk(gclk));
	jand g07061(.dina(n7294),.dinb(w_n7288_0[1]),.dout(n7295),.clk(gclk));
	jor g07062(.dina(w_n7295_0[2]),.dinb(w_n1699_48[0]),.dout(n7296),.clk(gclk));
	jand g07063(.dina(w_n7295_0[1]),.dinb(w_n1699_47[2]),.dout(n7297),.clk(gclk));
	jxor g07064(.dina(w_n6869_0[0]),.dinb(w_n1912_45[0]),.dout(n7298),.clk(gclk));
	jor g07065(.dina(n7298),.dinb(w_n7154_47[2]),.dout(n7299),.clk(gclk));
	jxor g07066(.dina(n7299),.dinb(w_n6875_0[0]),.dout(n7300),.clk(gclk));
	jor g07067(.dina(w_n7300_0[2]),.dinb(n7297),.dout(n7301),.clk(gclk));
	jand g07068(.dina(n7301),.dinb(w_n7296_0[1]),.dout(n7302),.clk(gclk));
	jor g07069(.dina(w_n7302_0[2]),.dinb(w_n1516_46[1]),.dout(n7303),.clk(gclk));
	jand g07070(.dina(w_n7302_0[1]),.dinb(w_n1516_46[0]),.dout(n7304),.clk(gclk));
	jxor g07071(.dina(w_n6877_0[0]),.dinb(w_n1699_47[1]),.dout(n7305),.clk(gclk));
	jor g07072(.dina(n7305),.dinb(w_n7154_47[1]),.dout(n7306),.clk(gclk));
	jxor g07073(.dina(n7306),.dinb(w_n6883_0[0]),.dout(n7307),.clk(gclk));
	jor g07074(.dina(w_n7307_0[2]),.dinb(n7304),.dout(n7308),.clk(gclk));
	jand g07075(.dina(n7308),.dinb(w_n7303_0[1]),.dout(n7309),.clk(gclk));
	jor g07076(.dina(w_n7309_0[2]),.dinb(w_n1332_48[0]),.dout(n7310),.clk(gclk));
	jand g07077(.dina(w_n7309_0[1]),.dinb(w_n1332_47[2]),.dout(n7311),.clk(gclk));
	jxor g07078(.dina(w_n6885_0[0]),.dinb(w_n1516_45[2]),.dout(n7312),.clk(gclk));
	jor g07079(.dina(n7312),.dinb(w_n7154_47[0]),.dout(n7313),.clk(gclk));
	jxor g07080(.dina(n7313),.dinb(w_n6891_0[0]),.dout(n7314),.clk(gclk));
	jor g07081(.dina(w_n7314_0[2]),.dinb(n7311),.dout(n7315),.clk(gclk));
	jand g07082(.dina(n7315),.dinb(w_n7310_0[1]),.dout(n7316),.clk(gclk));
	jor g07083(.dina(w_n7316_0[2]),.dinb(w_n1173_47[0]),.dout(n7317),.clk(gclk));
	jand g07084(.dina(w_n7316_0[1]),.dinb(w_n1173_46[2]),.dout(n7318),.clk(gclk));
	jxor g07085(.dina(w_n6893_0[0]),.dinb(w_n1332_47[1]),.dout(n7319),.clk(gclk));
	jor g07086(.dina(n7319),.dinb(w_n7154_46[2]),.dout(n7320),.clk(gclk));
	jxor g07087(.dina(n7320),.dinb(w_n7095_0[0]),.dout(n7321),.clk(gclk));
	jnot g07088(.din(w_n7321_0[2]),.dout(n7322),.clk(gclk));
	jor g07089(.dina(n7322),.dinb(n7318),.dout(n7323),.clk(gclk));
	jand g07090(.dina(n7323),.dinb(w_n7317_0[1]),.dout(n7324),.clk(gclk));
	jor g07091(.dina(w_n7324_0[2]),.dinb(w_n1008_49[0]),.dout(n7325),.clk(gclk));
	jand g07092(.dina(w_n7324_0[1]),.dinb(w_n1008_48[2]),.dout(n7326),.clk(gclk));
	jxor g07093(.dina(w_n6900_0[0]),.dinb(w_n1173_46[1]),.dout(n7327),.clk(gclk));
	jor g07094(.dina(n7327),.dinb(w_n7154_46[1]),.dout(n7328),.clk(gclk));
	jxor g07095(.dina(n7328),.dinb(w_n6906_0[0]),.dout(n7329),.clk(gclk));
	jor g07096(.dina(w_n7329_0[2]),.dinb(n7326),.dout(n7330),.clk(gclk));
	jand g07097(.dina(n7330),.dinb(w_n7325_0[1]),.dout(n7331),.clk(gclk));
	jor g07098(.dina(w_n7331_0[2]),.dinb(w_n884_48[0]),.dout(n7332),.clk(gclk));
	jand g07099(.dina(w_n7331_0[1]),.dinb(w_n884_47[2]),.dout(n7333),.clk(gclk));
	jxor g07100(.dina(w_n6908_0[0]),.dinb(w_n1008_48[1]),.dout(n7334),.clk(gclk));
	jor g07101(.dina(n7334),.dinb(w_n7154_46[0]),.dout(n7335),.clk(gclk));
	jxor g07102(.dina(n7335),.dinb(w_n7102_0[0]),.dout(n7336),.clk(gclk));
	jnot g07103(.din(w_n7336_0[2]),.dout(n7337),.clk(gclk));
	jor g07104(.dina(n7337),.dinb(n7333),.dout(n7338),.clk(gclk));
	jand g07105(.dina(n7338),.dinb(w_n7332_0[1]),.dout(n7339),.clk(gclk));
	jor g07106(.dina(w_n7339_0[2]),.dinb(w_n743_49[0]),.dout(n7340),.clk(gclk));
	jand g07107(.dina(w_n7339_0[1]),.dinb(w_n743_48[2]),.dout(n7341),.clk(gclk));
	jxor g07108(.dina(w_n6915_0[0]),.dinb(w_n884_47[1]),.dout(n7342),.clk(gclk));
	jor g07109(.dina(n7342),.dinb(w_n7154_45[2]),.dout(n7343),.clk(gclk));
	jxor g07110(.dina(n7343),.dinb(w_n6921_0[0]),.dout(n7344),.clk(gclk));
	jor g07111(.dina(w_n7344_0[2]),.dinb(n7341),.dout(n7345),.clk(gclk));
	jand g07112(.dina(n7345),.dinb(w_n7340_0[1]),.dout(n7346),.clk(gclk));
	jor g07113(.dina(w_n7346_0[2]),.dinb(w_n635_49[0]),.dout(n7347),.clk(gclk));
	jand g07114(.dina(w_n7346_0[1]),.dinb(w_n635_48[2]),.dout(n7348),.clk(gclk));
	jxor g07115(.dina(w_n6923_0[0]),.dinb(w_n743_48[1]),.dout(n7349),.clk(gclk));
	jor g07116(.dina(n7349),.dinb(w_n7154_45[1]),.dout(n7350),.clk(gclk));
	jxor g07117(.dina(n7350),.dinb(w_n7109_0[0]),.dout(n7351),.clk(gclk));
	jnot g07118(.din(w_n7351_0[2]),.dout(n7352),.clk(gclk));
	jor g07119(.dina(n7352),.dinb(n7348),.dout(n7353),.clk(gclk));
	jand g07120(.dina(n7353),.dinb(w_n7347_0[1]),.dout(n7354),.clk(gclk));
	jor g07121(.dina(w_n7354_0[2]),.dinb(w_n515_50[0]),.dout(n7355),.clk(gclk));
	jand g07122(.dina(w_n7354_0[1]),.dinb(w_n515_49[2]),.dout(n7356),.clk(gclk));
	jxor g07123(.dina(w_n6930_0[0]),.dinb(w_n635_48[1]),.dout(n7357),.clk(gclk));
	jor g07124(.dina(n7357),.dinb(w_n7154_45[0]),.dout(n7358),.clk(gclk));
	jxor g07125(.dina(n7358),.dinb(w_n7113_0[0]),.dout(n7359),.clk(gclk));
	jnot g07126(.din(w_n7359_0[2]),.dout(n7360),.clk(gclk));
	jor g07127(.dina(n7360),.dinb(n7356),.dout(n7361),.clk(gclk));
	jand g07128(.dina(n7361),.dinb(w_n7355_0[1]),.dout(n7362),.clk(gclk));
	jor g07129(.dina(w_n7362_0[2]),.dinb(w_n443_50[0]),.dout(n7363),.clk(gclk));
	jand g07130(.dina(w_n7362_0[1]),.dinb(w_n443_49[2]),.dout(n7364),.clk(gclk));
	jxor g07131(.dina(w_n6937_0[0]),.dinb(w_n515_49[1]),.dout(n7365),.clk(gclk));
	jor g07132(.dina(n7365),.dinb(w_n7154_44[2]),.dout(n7366),.clk(gclk));
	jxor g07133(.dina(n7366),.dinb(w_n6943_0[0]),.dout(n7367),.clk(gclk));
	jor g07134(.dina(w_n7367_0[2]),.dinb(n7364),.dout(n7368),.clk(gclk));
	jand g07135(.dina(n7368),.dinb(w_n7363_0[1]),.dout(n7369),.clk(gclk));
	jor g07136(.dina(w_n7369_0[2]),.dinb(w_n352_50[1]),.dout(n7370),.clk(gclk));
	jand g07137(.dina(w_n7369_0[1]),.dinb(w_n352_50[0]),.dout(n7371),.clk(gclk));
	jxor g07138(.dina(w_n6945_0[0]),.dinb(w_n443_49[1]),.dout(n7372),.clk(gclk));
	jor g07139(.dina(n7372),.dinb(w_n7154_44[1]),.dout(n7373),.clk(gclk));
	jxor g07140(.dina(n7373),.dinb(w_n6951_0[0]),.dout(n7374),.clk(gclk));
	jor g07141(.dina(w_n7374_0[2]),.dinb(n7371),.dout(n7375),.clk(gclk));
	jand g07142(.dina(n7375),.dinb(w_n7370_0[1]),.dout(n7376),.clk(gclk));
	jor g07143(.dina(w_n7376_0[2]),.dinb(w_n294_50[2]),.dout(n7377),.clk(gclk));
	jand g07144(.dina(w_n7376_0[1]),.dinb(w_n294_50[1]),.dout(n7378),.clk(gclk));
	jxor g07145(.dina(w_n6953_0[0]),.dinb(w_n352_49[2]),.dout(n7379),.clk(gclk));
	jor g07146(.dina(n7379),.dinb(w_n7154_44[0]),.dout(n7380),.clk(gclk));
	jxor g07147(.dina(n7380),.dinb(w_n6959_0[0]),.dout(n7381),.clk(gclk));
	jor g07148(.dina(w_n7381_0[2]),.dinb(n7378),.dout(n7382),.clk(gclk));
	jand g07149(.dina(n7382),.dinb(w_n7377_0[1]),.dout(n7383),.clk(gclk));
	jor g07150(.dina(w_n7383_0[2]),.dinb(w_n239_50[2]),.dout(n7384),.clk(gclk));
	jand g07151(.dina(w_n7383_0[1]),.dinb(w_n239_50[1]),.dout(n7385),.clk(gclk));
	jxor g07152(.dina(w_n6961_0[0]),.dinb(w_n294_50[0]),.dout(n7386),.clk(gclk));
	jor g07153(.dina(n7386),.dinb(w_n7154_43[2]),.dout(n7387),.clk(gclk));
	jxor g07154(.dina(n7387),.dinb(w_n7126_0[0]),.dout(n7388),.clk(gclk));
	jnot g07155(.din(w_n7388_0[2]),.dout(n7389),.clk(gclk));
	jor g07156(.dina(n7389),.dinb(n7385),.dout(n7390),.clk(gclk));
	jand g07157(.dina(n7390),.dinb(w_n7384_0[1]),.dout(n7391),.clk(gclk));
	jor g07158(.dina(w_n7391_0[2]),.dinb(w_n221_51[0]),.dout(n7392),.clk(gclk));
	jand g07159(.dina(w_n7391_0[1]),.dinb(w_n221_50[2]),.dout(n7393),.clk(gclk));
	jxor g07160(.dina(w_n6968_0[0]),.dinb(w_n239_50[0]),.dout(n7394),.clk(gclk));
	jor g07161(.dina(n7394),.dinb(w_n7154_43[1]),.dout(n7395),.clk(gclk));
	jxor g07162(.dina(n7395),.dinb(w_n7130_0[0]),.dout(n7396),.clk(gclk));
	jnot g07163(.din(w_n7396_0[2]),.dout(n7397),.clk(gclk));
	jor g07164(.dina(n7397),.dinb(n7393),.dout(n7398),.clk(gclk));
	jand g07165(.dina(n7398),.dinb(w_n7392_0[1]),.dout(n7399),.clk(gclk));
	jxor g07166(.dina(w_n6975_0[0]),.dinb(w_n221_50[1]),.dout(n7400),.clk(gclk));
	jor g07167(.dina(n7400),.dinb(w_n7154_43[0]),.dout(n7401),.clk(gclk));
	jxor g07168(.dina(n7401),.dinb(w_n6981_0[0]),.dout(n7402),.clk(gclk));
	jor g07169(.dina(w_n7402_1[1]),.dinb(w_n7399_0[2]),.dout(n7403),.clk(gclk));
	jor g07170(.dina(w_n7403_0[1]),.dinb(w_n6989_0[0]),.dout(n7404),.clk(gclk));
	jor g07171(.dina(n7404),.dinb(w_n7146_0[1]),.dout(n7405),.clk(gclk));
	jand g07172(.dina(n7405),.dinb(w_n218_21[0]),.dout(n7406),.clk(gclk));
	jand g07173(.dina(w_n7154_42[2]),.dinb(w_n6986_0[0]),.dout(n7407),.clk(gclk));
	jand g07174(.dina(w_n7402_1[0]),.dinb(w_n7399_0[1]),.dout(n7408),.clk(gclk));
	jor g07175(.dina(w_n7408_1[1]),.dinb(n7407),.dout(n7409),.clk(gclk));
	jand g07176(.dina(w_n7153_0[0]),.dinb(w_n7135_0[0]),.dout(n7410),.clk(gclk));
	jnot g07177(.din(n7410),.dout(n7411),.clk(gclk));
	jand g07178(.dina(w_n7136_0[0]),.dinb(w_asqrt63_38[0]),.dout(n7412),.clk(gclk));
	jand g07179(.dina(n7412),.dinb(w_n6988_0[2]),.dout(n7413),.clk(gclk));
	jand g07180(.dina(w_n7413_0[1]),.dinb(n7411),.dout(n7414),.clk(gclk));
	jor g07181(.dina(n7414),.dinb(n7409),.dout(n7415),.clk(gclk));
	jor g07182(.dina(w_n7415_0[1]),.dinb(w_n7406_0[1]),.dout(asqrt_fa_31),.clk(gclk));
	jxor g07183(.dina(w_n7391_0[0]),.dinb(w_n221_50[0]),.dout(n7417),.clk(gclk));
	jand g07184(.dina(n7417),.dinb(w_asqrt30_38),.dout(n7418),.clk(gclk));
	jxor g07185(.dina(n7418),.dinb(w_n7396_0[1]),.dout(n7419),.clk(gclk));
	jand g07186(.dina(w_asqrt30_37[2]),.dinb(w_a60_0[1]),.dout(n7420),.clk(gclk));
	jnot g07187(.din(w_a58_0[2]),.dout(n7421),.clk(gclk));
	jnot g07188(.din(w_a59_0[1]),.dout(n7422),.clk(gclk));
	jand g07189(.dina(w_n7422_0[1]),.dinb(w_n7421_1[2]),.dout(n7423),.clk(gclk));
	jand g07190(.dina(w_n7423_0[2]),.dinb(w_n7156_1[1]),.dout(n7424),.clk(gclk));
	jor g07191(.dina(w_n7424_0[1]),.dinb(n7420),.dout(n7425),.clk(gclk));
	jand g07192(.dina(w_n7425_0[2]),.dinb(w_asqrt31_22[2]),.dout(n7426),.clk(gclk));
	jor g07193(.dina(w_n7425_0[1]),.dinb(w_asqrt31_22[1]),.dout(n7427),.clk(gclk));
	jand g07194(.dina(w_asqrt30_37[1]),.dinb(w_n7156_1[0]),.dout(n7428),.clk(gclk));
	jor g07195(.dina(n7428),.dinb(w_n7157_0[0]),.dout(n7429),.clk(gclk));
	jnot g07196(.din(w_n7158_0[1]),.dout(n7430),.clk(gclk));
	jnot g07197(.din(w_n7146_0[0]),.dout(n7431),.clk(gclk));
	jnot g07198(.din(w_n7392_0[0]),.dout(n7432),.clk(gclk));
	jnot g07199(.din(w_n7384_0[0]),.dout(n7433),.clk(gclk));
	jnot g07200(.din(w_n7377_0[0]),.dout(n7434),.clk(gclk));
	jnot g07201(.din(w_n7370_0[0]),.dout(n7435),.clk(gclk));
	jnot g07202(.din(w_n7363_0[0]),.dout(n7436),.clk(gclk));
	jnot g07203(.din(w_n7355_0[0]),.dout(n7437),.clk(gclk));
	jnot g07204(.din(w_n7347_0[0]),.dout(n7438),.clk(gclk));
	jnot g07205(.din(w_n7340_0[0]),.dout(n7439),.clk(gclk));
	jnot g07206(.din(w_n7332_0[0]),.dout(n7440),.clk(gclk));
	jnot g07207(.din(w_n7325_0[0]),.dout(n7441),.clk(gclk));
	jnot g07208(.din(w_n7317_0[0]),.dout(n7442),.clk(gclk));
	jnot g07209(.din(w_n7310_0[0]),.dout(n7443),.clk(gclk));
	jnot g07210(.din(w_n7303_0[0]),.dout(n7444),.clk(gclk));
	jnot g07211(.din(w_n7296_0[0]),.dout(n7445),.clk(gclk));
	jnot g07212(.din(w_n7288_0[0]),.dout(n7446),.clk(gclk));
	jnot g07213(.din(w_n7280_0[0]),.dout(n7447),.clk(gclk));
	jnot g07214(.din(w_n7272_0[0]),.dout(n7448),.clk(gclk));
	jnot g07215(.din(w_n7265_0[0]),.dout(n7449),.clk(gclk));
	jnot g07216(.din(w_n7257_0[0]),.dout(n7450),.clk(gclk));
	jnot g07217(.din(w_n7250_0[0]),.dout(n7451),.clk(gclk));
	jnot g07218(.din(w_n7242_0[0]),.dout(n7452),.clk(gclk));
	jnot g07219(.din(w_n7235_0[0]),.dout(n7453),.clk(gclk));
	jnot g07220(.din(w_n7227_0[0]),.dout(n7454),.clk(gclk));
	jnot g07221(.din(w_n7220_0[0]),.dout(n7455),.clk(gclk));
	jnot g07222(.din(w_n7212_0[0]),.dout(n7456),.clk(gclk));
	jnot g07223(.din(w_n7204_0[0]),.dout(n7457),.clk(gclk));
	jnot g07224(.din(w_n7196_0[0]),.dout(n7458),.clk(gclk));
	jnot g07225(.din(w_n7189_0[0]),.dout(n7459),.clk(gclk));
	jnot g07226(.din(w_n7181_0[0]),.dout(n7460),.clk(gclk));
	jnot g07227(.din(w_n7170_0[0]),.dout(n7461),.clk(gclk));
	jnot g07228(.din(w_n7162_0[0]),.dout(n7462),.clk(gclk));
	jand g07229(.dina(w_asqrt31_22[0]),.dinb(w_n6606_0[2]),.dout(n7463),.clk(gclk));
	jor g07230(.dina(n7463),.dinb(w_n6607_0[0]),.dout(n7464),.clk(gclk));
	jand g07231(.dina(n7464),.dinb(w_n7173_0[0]),.dout(n7465),.clk(gclk));
	jand g07232(.dina(w_asqrt31_21[2]),.dinb(w_a62_0[0]),.dout(n7466),.clk(gclk));
	jor g07233(.dina(w_n7159_0[0]),.dinb(n7466),.dout(n7467),.clk(gclk));
	jor g07234(.dina(n7467),.dinb(w_asqrt32_27[1]),.dout(n7468),.clk(gclk));
	jand g07235(.dina(n7468),.dinb(w_n7465_0[1]),.dout(n7469),.clk(gclk));
	jor g07236(.dina(n7469),.dinb(n7462),.dout(n7470),.clk(gclk));
	jor g07237(.dina(n7470),.dinb(w_asqrt33_23[0]),.dout(n7471),.clk(gclk));
	jnot g07238(.din(w_n7178_0[1]),.dout(n7472),.clk(gclk));
	jand g07239(.dina(n7472),.dinb(n7471),.dout(n7473),.clk(gclk));
	jor g07240(.dina(n7473),.dinb(n7461),.dout(n7474),.clk(gclk));
	jor g07241(.dina(n7474),.dinb(w_asqrt34_27[2]),.dout(n7475),.clk(gclk));
	jand g07242(.dina(w_n7185_0[1]),.dinb(n7475),.dout(n7476),.clk(gclk));
	jor g07243(.dina(n7476),.dinb(n7460),.dout(n7477),.clk(gclk));
	jor g07244(.dina(n7477),.dinb(w_asqrt35_23[2]),.dout(n7478),.clk(gclk));
	jnot g07245(.din(w_n7193_0[1]),.dout(n7479),.clk(gclk));
	jand g07246(.dina(n7479),.dinb(n7478),.dout(n7480),.clk(gclk));
	jor g07247(.dina(n7480),.dinb(n7459),.dout(n7481),.clk(gclk));
	jor g07248(.dina(n7481),.dinb(w_asqrt36_27[2]),.dout(n7482),.clk(gclk));
	jand g07249(.dina(w_n7200_0[1]),.dinb(n7482),.dout(n7483),.clk(gclk));
	jor g07250(.dina(n7483),.dinb(n7458),.dout(n7484),.clk(gclk));
	jor g07251(.dina(n7484),.dinb(w_asqrt37_24[0]),.dout(n7485),.clk(gclk));
	jand g07252(.dina(w_n7208_0[1]),.dinb(n7485),.dout(n7486),.clk(gclk));
	jor g07253(.dina(n7486),.dinb(n7457),.dout(n7487),.clk(gclk));
	jor g07254(.dina(n7487),.dinb(w_asqrt38_28[0]),.dout(n7488),.clk(gclk));
	jand g07255(.dina(w_n7216_0[1]),.dinb(n7488),.dout(n7489),.clk(gclk));
	jor g07256(.dina(n7489),.dinb(n7456),.dout(n7490),.clk(gclk));
	jor g07257(.dina(n7490),.dinb(w_asqrt39_24[2]),.dout(n7491),.clk(gclk));
	jnot g07258(.din(w_n7224_0[1]),.dout(n7492),.clk(gclk));
	jand g07259(.dina(n7492),.dinb(n7491),.dout(n7493),.clk(gclk));
	jor g07260(.dina(n7493),.dinb(n7455),.dout(n7494),.clk(gclk));
	jor g07261(.dina(n7494),.dinb(w_asqrt40_28[0]),.dout(n7495),.clk(gclk));
	jand g07262(.dina(w_n7231_0[1]),.dinb(n7495),.dout(n7496),.clk(gclk));
	jor g07263(.dina(n7496),.dinb(n7454),.dout(n7497),.clk(gclk));
	jor g07264(.dina(n7497),.dinb(w_asqrt41_25[0]),.dout(n7498),.clk(gclk));
	jnot g07265(.din(w_n7239_0[1]),.dout(n7499),.clk(gclk));
	jand g07266(.dina(n7499),.dinb(n7498),.dout(n7500),.clk(gclk));
	jor g07267(.dina(n7500),.dinb(n7453),.dout(n7501),.clk(gclk));
	jor g07268(.dina(n7501),.dinb(w_asqrt42_28[1]),.dout(n7502),.clk(gclk));
	jand g07269(.dina(w_n7246_0[1]),.dinb(n7502),.dout(n7503),.clk(gclk));
	jor g07270(.dina(n7503),.dinb(n7452),.dout(n7504),.clk(gclk));
	jor g07271(.dina(n7504),.dinb(w_asqrt43_25[1]),.dout(n7505),.clk(gclk));
	jnot g07272(.din(w_n7254_0[1]),.dout(n7506),.clk(gclk));
	jand g07273(.dina(n7506),.dinb(n7505),.dout(n7507),.clk(gclk));
	jor g07274(.dina(n7507),.dinb(n7451),.dout(n7508),.clk(gclk));
	jor g07275(.dina(n7508),.dinb(w_asqrt44_28[1]),.dout(n7509),.clk(gclk));
	jand g07276(.dina(w_n7261_0[1]),.dinb(n7509),.dout(n7510),.clk(gclk));
	jor g07277(.dina(n7510),.dinb(n7450),.dout(n7511),.clk(gclk));
	jor g07278(.dina(n7511),.dinb(w_asqrt45_26[0]),.dout(n7512),.clk(gclk));
	jnot g07279(.din(w_n7269_0[1]),.dout(n7513),.clk(gclk));
	jand g07280(.dina(n7513),.dinb(n7512),.dout(n7514),.clk(gclk));
	jor g07281(.dina(n7514),.dinb(n7449),.dout(n7515),.clk(gclk));
	jor g07282(.dina(n7515),.dinb(w_asqrt46_28[1]),.dout(n7516),.clk(gclk));
	jand g07283(.dina(w_n7276_0[1]),.dinb(n7516),.dout(n7517),.clk(gclk));
	jor g07284(.dina(n7517),.dinb(n7448),.dout(n7518),.clk(gclk));
	jor g07285(.dina(n7518),.dinb(w_asqrt47_26[2]),.dout(n7519),.clk(gclk));
	jand g07286(.dina(w_n7284_0[1]),.dinb(n7519),.dout(n7520),.clk(gclk));
	jor g07287(.dina(n7520),.dinb(n7447),.dout(n7521),.clk(gclk));
	jor g07288(.dina(n7521),.dinb(w_asqrt48_28[2]),.dout(n7522),.clk(gclk));
	jand g07289(.dina(w_n7292_0[1]),.dinb(n7522),.dout(n7523),.clk(gclk));
	jor g07290(.dina(n7523),.dinb(n7446),.dout(n7524),.clk(gclk));
	jor g07291(.dina(n7524),.dinb(w_asqrt49_27[0]),.dout(n7525),.clk(gclk));
	jnot g07292(.din(w_n7300_0[1]),.dout(n7526),.clk(gclk));
	jand g07293(.dina(n7526),.dinb(n7525),.dout(n7527),.clk(gclk));
	jor g07294(.dina(n7527),.dinb(n7445),.dout(n7528),.clk(gclk));
	jor g07295(.dina(n7528),.dinb(w_asqrt50_29[0]),.dout(n7529),.clk(gclk));
	jnot g07296(.din(w_n7307_0[1]),.dout(n7530),.clk(gclk));
	jand g07297(.dina(n7530),.dinb(n7529),.dout(n7531),.clk(gclk));
	jor g07298(.dina(n7531),.dinb(n7444),.dout(n7532),.clk(gclk));
	jor g07299(.dina(n7532),.dinb(w_asqrt51_27[1]),.dout(n7533),.clk(gclk));
	jnot g07300(.din(w_n7314_0[1]),.dout(n7534),.clk(gclk));
	jand g07301(.dina(n7534),.dinb(n7533),.dout(n7535),.clk(gclk));
	jor g07302(.dina(n7535),.dinb(n7443),.dout(n7536),.clk(gclk));
	jor g07303(.dina(n7536),.dinb(w_asqrt52_29[0]),.dout(n7537),.clk(gclk));
	jand g07304(.dina(w_n7321_0[1]),.dinb(n7537),.dout(n7538),.clk(gclk));
	jor g07305(.dina(n7538),.dinb(n7442),.dout(n7539),.clk(gclk));
	jor g07306(.dina(n7539),.dinb(w_asqrt53_28[0]),.dout(n7540),.clk(gclk));
	jnot g07307(.din(w_n7329_0[1]),.dout(n7541),.clk(gclk));
	jand g07308(.dina(n7541),.dinb(n7540),.dout(n7542),.clk(gclk));
	jor g07309(.dina(n7542),.dinb(n7441),.dout(n7543),.clk(gclk));
	jor g07310(.dina(n7543),.dinb(w_asqrt54_29[0]),.dout(n7544),.clk(gclk));
	jand g07311(.dina(w_n7336_0[1]),.dinb(n7544),.dout(n7545),.clk(gclk));
	jor g07312(.dina(n7545),.dinb(n7440),.dout(n7546),.clk(gclk));
	jor g07313(.dina(n7546),.dinb(w_asqrt55_28[1]),.dout(n7547),.clk(gclk));
	jnot g07314(.din(w_n7344_0[1]),.dout(n7548),.clk(gclk));
	jand g07315(.dina(n7548),.dinb(n7547),.dout(n7549),.clk(gclk));
	jor g07316(.dina(n7549),.dinb(n7439),.dout(n7550),.clk(gclk));
	jor g07317(.dina(n7550),.dinb(w_asqrt56_29[1]),.dout(n7551),.clk(gclk));
	jand g07318(.dina(w_n7351_0[1]),.dinb(n7551),.dout(n7552),.clk(gclk));
	jor g07319(.dina(n7552),.dinb(n7438),.dout(n7553),.clk(gclk));
	jor g07320(.dina(n7553),.dinb(w_asqrt57_29[0]),.dout(n7554),.clk(gclk));
	jand g07321(.dina(w_n7359_0[1]),.dinb(n7554),.dout(n7555),.clk(gclk));
	jor g07322(.dina(n7555),.dinb(n7437),.dout(n7556),.clk(gclk));
	jor g07323(.dina(n7556),.dinb(w_asqrt58_29[2]),.dout(n7557),.clk(gclk));
	jnot g07324(.din(w_n7367_0[1]),.dout(n7558),.clk(gclk));
	jand g07325(.dina(n7558),.dinb(n7557),.dout(n7559),.clk(gclk));
	jor g07326(.dina(n7559),.dinb(n7436),.dout(n7560),.clk(gclk));
	jor g07327(.dina(n7560),.dinb(w_asqrt59_29[1]),.dout(n7561),.clk(gclk));
	jnot g07328(.din(w_n7374_0[1]),.dout(n7562),.clk(gclk));
	jand g07329(.dina(n7562),.dinb(n7561),.dout(n7563),.clk(gclk));
	jor g07330(.dina(n7563),.dinb(n7435),.dout(n7564),.clk(gclk));
	jor g07331(.dina(n7564),.dinb(w_asqrt60_29[2]),.dout(n7565),.clk(gclk));
	jnot g07332(.din(w_n7381_0[1]),.dout(n7566),.clk(gclk));
	jand g07333(.dina(n7566),.dinb(n7565),.dout(n7567),.clk(gclk));
	jor g07334(.dina(n7567),.dinb(n7434),.dout(n7568),.clk(gclk));
	jor g07335(.dina(n7568),.dinb(w_asqrt61_29[2]),.dout(n7569),.clk(gclk));
	jand g07336(.dina(w_n7388_0[1]),.dinb(n7569),.dout(n7570),.clk(gclk));
	jor g07337(.dina(n7570),.dinb(n7433),.dout(n7571),.clk(gclk));
	jor g07338(.dina(n7571),.dinb(w_asqrt62_29[2]),.dout(n7572),.clk(gclk));
	jand g07339(.dina(w_n7396_0[0]),.dinb(n7572),.dout(n7573),.clk(gclk));
	jor g07340(.dina(n7573),.dinb(n7432),.dout(n7574),.clk(gclk));
	jnot g07341(.din(w_n7402_0[2]),.dout(n7575),.clk(gclk));
	jand g07342(.dina(n7575),.dinb(n7574),.dout(n7576),.clk(gclk));
	jand g07343(.dina(w_n7576_0[1]),.dinb(w_n6988_0[1]),.dout(n7577),.clk(gclk));
	jand g07344(.dina(n7577),.dinb(n7431),.dout(n7578),.clk(gclk));
	jor g07345(.dina(n7578),.dinb(w_asqrt63_37[2]),.dout(n7579),.clk(gclk));
	jnot g07346(.din(w_n7415_0[0]),.dout(n7580),.clk(gclk));
	jand g07347(.dina(n7580),.dinb(n7579),.dout(n7581),.clk(gclk));
	jor g07348(.dina(w_n7581_38[1]),.dinb(n7430),.dout(n7582),.clk(gclk));
	jand g07349(.dina(w_n7582_0[1]),.dinb(n7429),.dout(n7583),.clk(gclk));
	jand g07350(.dina(w_n7583_0[1]),.dinb(n7427),.dout(n7584),.clk(gclk));
	jor g07351(.dina(n7584),.dinb(w_n7426_0[1]),.dout(n7585),.clk(gclk));
	jand g07352(.dina(w_n7585_0[2]),.dinb(w_asqrt32_27[0]),.dout(n7586),.clk(gclk));
	jor g07353(.dina(w_n7585_0[1]),.dinb(w_asqrt32_26[2]),.dout(n7587),.clk(gclk));
	jor g07354(.dina(w_n7413_0[0]),.dinb(w_n7408_1[0]),.dout(n7588),.clk(gclk));
	jor g07355(.dina(n7588),.dinb(w_n7406_0[0]),.dout(n7589),.clk(gclk));
	jor g07356(.dina(n7589),.dinb(w_n7154_42[1]),.dout(n7590),.clk(gclk));
	jand g07357(.dina(n7590),.dinb(w_n7582_0[0]),.dout(n7591),.clk(gclk));
	jxor g07358(.dina(n7591),.dinb(w_n6606_0[1]),.dout(n7592),.clk(gclk));
	jnot g07359(.din(w_n7592_0[1]),.dout(n7593),.clk(gclk));
	jand g07360(.dina(w_n7593_0[1]),.dinb(n7587),.dout(n7594),.clk(gclk));
	jor g07361(.dina(n7594),.dinb(w_n7586_0[1]),.dout(n7595),.clk(gclk));
	jand g07362(.dina(w_n7595_0[2]),.dinb(w_asqrt33_22[2]),.dout(n7596),.clk(gclk));
	jxor g07363(.dina(w_n7161_0[0]),.dinb(w_n6758_38[0]),.dout(n7597),.clk(gclk));
	jand g07364(.dina(n7597),.dinb(w_asqrt30_37[0]),.dout(n7598),.clk(gclk));
	jxor g07365(.dina(n7598),.dinb(w_n7465_0[0]),.dout(n7599),.clk(gclk));
	jor g07366(.dina(w_n7595_0[1]),.dinb(w_asqrt33_22[1]),.dout(n7600),.clk(gclk));
	jand g07367(.dina(n7600),.dinb(w_n7599_0[1]),.dout(n7601),.clk(gclk));
	jor g07368(.dina(n7601),.dinb(w_n7596_0[1]),.dout(n7602),.clk(gclk));
	jand g07369(.dina(w_n7602_0[2]),.dinb(w_asqrt34_27[1]),.dout(n7603),.clk(gclk));
	jor g07370(.dina(w_n7602_0[1]),.dinb(w_asqrt34_27[0]),.dout(n7604),.clk(gclk));
	jxor g07371(.dina(w_n7169_0[0]),.dinb(w_n6357_42[2]),.dout(n7605),.clk(gclk));
	jand g07372(.dina(n7605),.dinb(w_asqrt30_36[2]),.dout(n7606),.clk(gclk));
	jxor g07373(.dina(n7606),.dinb(w_n7178_0[0]),.dout(n7607),.clk(gclk));
	jnot g07374(.din(w_n7607_0[1]),.dout(n7608),.clk(gclk));
	jand g07375(.dina(w_n7608_0[1]),.dinb(n7604),.dout(n7609),.clk(gclk));
	jor g07376(.dina(n7609),.dinb(w_n7603_0[1]),.dout(n7610),.clk(gclk));
	jand g07377(.dina(w_n7610_0[2]),.dinb(w_asqrt35_23[1]),.dout(n7611),.clk(gclk));
	jor g07378(.dina(w_n7610_0[1]),.dinb(w_asqrt35_23[0]),.dout(n7612),.clk(gclk));
	jxor g07379(.dina(w_n7180_0[0]),.dinb(w_n5989_38[2]),.dout(n7613),.clk(gclk));
	jand g07380(.dina(n7613),.dinb(w_asqrt30_36[1]),.dout(n7614),.clk(gclk));
	jxor g07381(.dina(n7614),.dinb(w_n7185_0[0]),.dout(n7615),.clk(gclk));
	jand g07382(.dina(w_n7615_0[1]),.dinb(n7612),.dout(n7616),.clk(gclk));
	jor g07383(.dina(n7616),.dinb(w_n7611_0[1]),.dout(n7617),.clk(gclk));
	jand g07384(.dina(w_n7617_0[2]),.dinb(w_asqrt36_27[1]),.dout(n7618),.clk(gclk));
	jor g07385(.dina(w_n7617_0[1]),.dinb(w_asqrt36_27[0]),.dout(n7619),.clk(gclk));
	jxor g07386(.dina(w_n7188_0[0]),.dinb(w_n5606_43[0]),.dout(n7620),.clk(gclk));
	jand g07387(.dina(n7620),.dinb(w_asqrt30_36[0]),.dout(n7621),.clk(gclk));
	jxor g07388(.dina(n7621),.dinb(w_n7193_0[0]),.dout(n7622),.clk(gclk));
	jnot g07389(.din(w_n7622_0[1]),.dout(n7623),.clk(gclk));
	jand g07390(.dina(w_n7623_0[1]),.dinb(n7619),.dout(n7624),.clk(gclk));
	jor g07391(.dina(n7624),.dinb(w_n7618_0[1]),.dout(n7625),.clk(gclk));
	jand g07392(.dina(w_n7625_0[2]),.dinb(w_asqrt37_23[2]),.dout(n7626),.clk(gclk));
	jor g07393(.dina(w_n7625_0[1]),.dinb(w_asqrt37_23[1]),.dout(n7627),.clk(gclk));
	jxor g07394(.dina(w_n7195_0[0]),.dinb(w_n5259_39[2]),.dout(n7628),.clk(gclk));
	jand g07395(.dina(n7628),.dinb(w_asqrt30_35[2]),.dout(n7629),.clk(gclk));
	jxor g07396(.dina(n7629),.dinb(w_n7200_0[0]),.dout(n7630),.clk(gclk));
	jand g07397(.dina(w_n7630_0[1]),.dinb(n7627),.dout(n7631),.clk(gclk));
	jor g07398(.dina(n7631),.dinb(w_n7626_0[1]),.dout(n7632),.clk(gclk));
	jand g07399(.dina(w_n7632_0[2]),.dinb(w_asqrt38_27[2]),.dout(n7633),.clk(gclk));
	jor g07400(.dina(w_n7632_0[1]),.dinb(w_asqrt38_27[1]),.dout(n7634),.clk(gclk));
	jxor g07401(.dina(w_n7203_0[0]),.dinb(w_n4902_43[2]),.dout(n7635),.clk(gclk));
	jand g07402(.dina(n7635),.dinb(w_asqrt30_35[1]),.dout(n7636),.clk(gclk));
	jxor g07403(.dina(n7636),.dinb(w_n7208_0[0]),.dout(n7637),.clk(gclk));
	jand g07404(.dina(w_n7637_0[1]),.dinb(n7634),.dout(n7638),.clk(gclk));
	jor g07405(.dina(n7638),.dinb(w_n7633_0[1]),.dout(n7639),.clk(gclk));
	jand g07406(.dina(w_n7639_0[2]),.dinb(w_asqrt39_24[1]),.dout(n7640),.clk(gclk));
	jor g07407(.dina(w_n7639_0[1]),.dinb(w_asqrt39_24[0]),.dout(n7641),.clk(gclk));
	jxor g07408(.dina(w_n7211_0[0]),.dinb(w_n4582_40[2]),.dout(n7642),.clk(gclk));
	jand g07409(.dina(n7642),.dinb(w_asqrt30_35[0]),.dout(n7643),.clk(gclk));
	jxor g07410(.dina(n7643),.dinb(w_n7216_0[0]),.dout(n7644),.clk(gclk));
	jand g07411(.dina(w_n7644_0[1]),.dinb(n7641),.dout(n7645),.clk(gclk));
	jor g07412(.dina(n7645),.dinb(w_n7640_0[1]),.dout(n7646),.clk(gclk));
	jand g07413(.dina(w_n7646_0[2]),.dinb(w_asqrt40_27[2]),.dout(n7647),.clk(gclk));
	jor g07414(.dina(w_n7646_0[1]),.dinb(w_asqrt40_27[1]),.dout(n7648),.clk(gclk));
	jxor g07415(.dina(w_n7219_0[0]),.dinb(w_n4249_44[1]),.dout(n7649),.clk(gclk));
	jand g07416(.dina(n7649),.dinb(w_asqrt30_34[2]),.dout(n7650),.clk(gclk));
	jxor g07417(.dina(n7650),.dinb(w_n7224_0[0]),.dout(n7651),.clk(gclk));
	jnot g07418(.din(w_n7651_0[1]),.dout(n7652),.clk(gclk));
	jand g07419(.dina(w_n7652_0[1]),.dinb(n7648),.dout(n7653),.clk(gclk));
	jor g07420(.dina(n7653),.dinb(w_n7647_0[1]),.dout(n7654),.clk(gclk));
	jand g07421(.dina(w_n7654_0[2]),.dinb(w_asqrt41_24[2]),.dout(n7655),.clk(gclk));
	jor g07422(.dina(w_n7654_0[1]),.dinb(w_asqrt41_24[1]),.dout(n7656),.clk(gclk));
	jxor g07423(.dina(w_n7226_0[0]),.dinb(w_n3955_41[1]),.dout(n7657),.clk(gclk));
	jand g07424(.dina(n7657),.dinb(w_asqrt30_34[1]),.dout(n7658),.clk(gclk));
	jxor g07425(.dina(n7658),.dinb(w_n7231_0[0]),.dout(n7659),.clk(gclk));
	jand g07426(.dina(w_n7659_0[1]),.dinb(n7656),.dout(n7660),.clk(gclk));
	jor g07427(.dina(n7660),.dinb(w_n7655_0[1]),.dout(n7661),.clk(gclk));
	jand g07428(.dina(w_n7661_0[2]),.dinb(w_asqrt42_28[0]),.dout(n7662),.clk(gclk));
	jor g07429(.dina(w_n7661_0[1]),.dinb(w_asqrt42_27[2]),.dout(n7663),.clk(gclk));
	jxor g07430(.dina(w_n7234_0[0]),.dinb(w_n3642_44[2]),.dout(n7664),.clk(gclk));
	jand g07431(.dina(n7664),.dinb(w_asqrt30_34[0]),.dout(n7665),.clk(gclk));
	jxor g07432(.dina(n7665),.dinb(w_n7239_0[0]),.dout(n7666),.clk(gclk));
	jnot g07433(.din(w_n7666_0[1]),.dout(n7667),.clk(gclk));
	jand g07434(.dina(w_n7667_0[1]),.dinb(n7663),.dout(n7668),.clk(gclk));
	jor g07435(.dina(n7668),.dinb(w_n7662_0[1]),.dout(n7669),.clk(gclk));
	jand g07436(.dina(w_n7669_0[2]),.dinb(w_asqrt43_25[0]),.dout(n7670),.clk(gclk));
	jor g07437(.dina(w_n7669_0[1]),.dinb(w_asqrt43_24[2]),.dout(n7671),.clk(gclk));
	jxor g07438(.dina(w_n7241_0[0]),.dinb(w_n3368_42[0]),.dout(n7672),.clk(gclk));
	jand g07439(.dina(n7672),.dinb(w_asqrt30_33[2]),.dout(n7673),.clk(gclk));
	jxor g07440(.dina(n7673),.dinb(w_n7246_0[0]),.dout(n7674),.clk(gclk));
	jand g07441(.dina(w_n7674_0[1]),.dinb(n7671),.dout(n7675),.clk(gclk));
	jor g07442(.dina(n7675),.dinb(w_n7670_0[1]),.dout(n7676),.clk(gclk));
	jand g07443(.dina(w_n7676_0[2]),.dinb(w_asqrt44_28[0]),.dout(n7677),.clk(gclk));
	jor g07444(.dina(w_n7676_0[1]),.dinb(w_asqrt44_27[2]),.dout(n7678),.clk(gclk));
	jxor g07445(.dina(w_n7249_0[0]),.dinb(w_n3089_45[1]),.dout(n7679),.clk(gclk));
	jand g07446(.dina(n7679),.dinb(w_asqrt30_33[1]),.dout(n7680),.clk(gclk));
	jxor g07447(.dina(n7680),.dinb(w_n7254_0[0]),.dout(n7681),.clk(gclk));
	jnot g07448(.din(w_n7681_0[1]),.dout(n7682),.clk(gclk));
	jand g07449(.dina(w_n7682_0[1]),.dinb(n7678),.dout(n7683),.clk(gclk));
	jor g07450(.dina(n7683),.dinb(w_n7677_0[1]),.dout(n7684),.clk(gclk));
	jand g07451(.dina(w_n7684_0[2]),.dinb(w_asqrt45_25[2]),.dout(n7685),.clk(gclk));
	jor g07452(.dina(w_n7684_0[1]),.dinb(w_asqrt45_25[1]),.dout(n7686),.clk(gclk));
	jxor g07453(.dina(w_n7256_0[0]),.dinb(w_n2833_43[0]),.dout(n7687),.clk(gclk));
	jand g07454(.dina(n7687),.dinb(w_asqrt30_33[0]),.dout(n7688),.clk(gclk));
	jxor g07455(.dina(n7688),.dinb(w_n7261_0[0]),.dout(n7689),.clk(gclk));
	jand g07456(.dina(w_n7689_0[1]),.dinb(n7686),.dout(n7690),.clk(gclk));
	jor g07457(.dina(n7690),.dinb(w_n7685_0[1]),.dout(n7691),.clk(gclk));
	jand g07458(.dina(w_n7691_0[2]),.dinb(w_asqrt46_28[0]),.dout(n7692),.clk(gclk));
	jor g07459(.dina(w_n7691_0[1]),.dinb(w_asqrt46_27[2]),.dout(n7693),.clk(gclk));
	jxor g07460(.dina(w_n7264_0[0]),.dinb(w_n2572_45[2]),.dout(n7694),.clk(gclk));
	jand g07461(.dina(n7694),.dinb(w_asqrt30_32[2]),.dout(n7695),.clk(gclk));
	jxor g07462(.dina(n7695),.dinb(w_n7269_0[0]),.dout(n7696),.clk(gclk));
	jnot g07463(.din(w_n7696_0[1]),.dout(n7697),.clk(gclk));
	jand g07464(.dina(w_n7697_0[1]),.dinb(n7693),.dout(n7698),.clk(gclk));
	jor g07465(.dina(n7698),.dinb(w_n7692_0[1]),.dout(n7699),.clk(gclk));
	jand g07466(.dina(w_n7699_0[2]),.dinb(w_asqrt47_26[1]),.dout(n7700),.clk(gclk));
	jor g07467(.dina(w_n7699_0[1]),.dinb(w_asqrt47_26[0]),.dout(n7701),.clk(gclk));
	jxor g07468(.dina(w_n7271_0[0]),.dinb(w_n2345_43[2]),.dout(n7702),.clk(gclk));
	jand g07469(.dina(n7702),.dinb(w_asqrt30_32[1]),.dout(n7703),.clk(gclk));
	jxor g07470(.dina(n7703),.dinb(w_n7276_0[0]),.dout(n7704),.clk(gclk));
	jand g07471(.dina(w_n7704_0[1]),.dinb(n7701),.dout(n7705),.clk(gclk));
	jor g07472(.dina(n7705),.dinb(w_n7700_0[1]),.dout(n7706),.clk(gclk));
	jand g07473(.dina(w_n7706_0[2]),.dinb(w_asqrt48_28[1]),.dout(n7707),.clk(gclk));
	jor g07474(.dina(w_n7706_0[1]),.dinb(w_asqrt48_28[0]),.dout(n7708),.clk(gclk));
	jxor g07475(.dina(w_n7279_0[0]),.dinb(w_n2108_46[1]),.dout(n7709),.clk(gclk));
	jand g07476(.dina(n7709),.dinb(w_asqrt30_32[0]),.dout(n7710),.clk(gclk));
	jxor g07477(.dina(n7710),.dinb(w_n7284_0[0]),.dout(n7711),.clk(gclk));
	jand g07478(.dina(w_n7711_0[1]),.dinb(n7708),.dout(n7712),.clk(gclk));
	jor g07479(.dina(n7712),.dinb(w_n7707_0[1]),.dout(n7713),.clk(gclk));
	jand g07480(.dina(w_n7713_0[2]),.dinb(w_asqrt49_26[2]),.dout(n7714),.clk(gclk));
	jor g07481(.dina(w_n7713_0[1]),.dinb(w_asqrt49_26[1]),.dout(n7715),.clk(gclk));
	jxor g07482(.dina(w_n7287_0[0]),.dinb(w_n1912_44[2]),.dout(n7716),.clk(gclk));
	jand g07483(.dina(n7716),.dinb(w_asqrt30_31[2]),.dout(n7717),.clk(gclk));
	jxor g07484(.dina(n7717),.dinb(w_n7292_0[0]),.dout(n7718),.clk(gclk));
	jand g07485(.dina(w_n7718_0[1]),.dinb(n7715),.dout(n7719),.clk(gclk));
	jor g07486(.dina(n7719),.dinb(w_n7714_0[1]),.dout(n7720),.clk(gclk));
	jand g07487(.dina(w_n7720_0[2]),.dinb(w_asqrt50_28[2]),.dout(n7721),.clk(gclk));
	jor g07488(.dina(w_n7720_0[1]),.dinb(w_asqrt50_28[1]),.dout(n7722),.clk(gclk));
	jxor g07489(.dina(w_n7295_0[0]),.dinb(w_n1699_47[0]),.dout(n7723),.clk(gclk));
	jand g07490(.dina(n7723),.dinb(w_asqrt30_31[1]),.dout(n7724),.clk(gclk));
	jxor g07491(.dina(n7724),.dinb(w_n7300_0[0]),.dout(n7725),.clk(gclk));
	jnot g07492(.din(w_n7725_0[1]),.dout(n7726),.clk(gclk));
	jand g07493(.dina(w_n7726_0[1]),.dinb(n7722),.dout(n7727),.clk(gclk));
	jor g07494(.dina(n7727),.dinb(w_n7721_0[1]),.dout(n7728),.clk(gclk));
	jand g07495(.dina(w_n7728_0[2]),.dinb(w_asqrt51_27[0]),.dout(n7729),.clk(gclk));
	jor g07496(.dina(w_n7728_0[1]),.dinb(w_asqrt51_26[2]),.dout(n7730),.clk(gclk));
	jxor g07497(.dina(w_n7302_0[0]),.dinb(w_n1516_45[1]),.dout(n7731),.clk(gclk));
	jand g07498(.dina(n7731),.dinb(w_asqrt30_31[0]),.dout(n7732),.clk(gclk));
	jxor g07499(.dina(n7732),.dinb(w_n7307_0[0]),.dout(n7733),.clk(gclk));
	jnot g07500(.din(w_n7733_0[1]),.dout(n7734),.clk(gclk));
	jand g07501(.dina(w_n7734_0[1]),.dinb(n7730),.dout(n7735),.clk(gclk));
	jor g07502(.dina(n7735),.dinb(w_n7729_0[1]),.dout(n7736),.clk(gclk));
	jand g07503(.dina(w_n7736_0[2]),.dinb(w_asqrt52_28[2]),.dout(n7737),.clk(gclk));
	jor g07504(.dina(w_n7736_0[1]),.dinb(w_asqrt52_28[1]),.dout(n7738),.clk(gclk));
	jxor g07505(.dina(w_n7309_0[0]),.dinb(w_n1332_47[0]),.dout(n7739),.clk(gclk));
	jand g07506(.dina(n7739),.dinb(w_asqrt30_30[2]),.dout(n7740),.clk(gclk));
	jxor g07507(.dina(n7740),.dinb(w_n7314_0[0]),.dout(n7741),.clk(gclk));
	jnot g07508(.din(w_n7741_0[1]),.dout(n7742),.clk(gclk));
	jand g07509(.dina(w_n7742_0[1]),.dinb(n7738),.dout(n7743),.clk(gclk));
	jor g07510(.dina(n7743),.dinb(w_n7737_0[1]),.dout(n7744),.clk(gclk));
	jand g07511(.dina(w_n7744_0[2]),.dinb(w_asqrt53_27[2]),.dout(n7745),.clk(gclk));
	jor g07512(.dina(w_n7744_0[1]),.dinb(w_asqrt53_27[1]),.dout(n7746),.clk(gclk));
	jxor g07513(.dina(w_n7316_0[0]),.dinb(w_n1173_46[0]),.dout(n7747),.clk(gclk));
	jand g07514(.dina(n7747),.dinb(w_asqrt30_30[1]),.dout(n7748),.clk(gclk));
	jxor g07515(.dina(n7748),.dinb(w_n7321_0[0]),.dout(n7749),.clk(gclk));
	jand g07516(.dina(w_n7749_0[1]),.dinb(n7746),.dout(n7750),.clk(gclk));
	jor g07517(.dina(n7750),.dinb(w_n7745_0[1]),.dout(n7751),.clk(gclk));
	jand g07518(.dina(w_n7751_0[2]),.dinb(w_asqrt54_28[2]),.dout(n7752),.clk(gclk));
	jor g07519(.dina(w_n7751_0[1]),.dinb(w_asqrt54_28[1]),.dout(n7753),.clk(gclk));
	jxor g07520(.dina(w_n7324_0[0]),.dinb(w_n1008_48[0]),.dout(n7754),.clk(gclk));
	jand g07521(.dina(n7754),.dinb(w_asqrt30_30[0]),.dout(n7755),.clk(gclk));
	jxor g07522(.dina(n7755),.dinb(w_n7329_0[0]),.dout(n7756),.clk(gclk));
	jnot g07523(.din(w_n7756_0[1]),.dout(n7757),.clk(gclk));
	jand g07524(.dina(w_n7757_0[1]),.dinb(n7753),.dout(n7758),.clk(gclk));
	jor g07525(.dina(n7758),.dinb(w_n7752_0[1]),.dout(n7759),.clk(gclk));
	jand g07526(.dina(w_n7759_0[2]),.dinb(w_asqrt55_28[0]),.dout(n7760),.clk(gclk));
	jor g07527(.dina(w_n7759_0[1]),.dinb(w_asqrt55_27[2]),.dout(n7761),.clk(gclk));
	jxor g07528(.dina(w_n7331_0[0]),.dinb(w_n884_47[0]),.dout(n7762),.clk(gclk));
	jand g07529(.dina(n7762),.dinb(w_asqrt30_29[2]),.dout(n7763),.clk(gclk));
	jxor g07530(.dina(n7763),.dinb(w_n7336_0[0]),.dout(n7764),.clk(gclk));
	jand g07531(.dina(w_n7764_0[1]),.dinb(n7761),.dout(n7765),.clk(gclk));
	jor g07532(.dina(n7765),.dinb(w_n7760_0[1]),.dout(n7766),.clk(gclk));
	jand g07533(.dina(w_n7766_0[2]),.dinb(w_asqrt56_29[0]),.dout(n7767),.clk(gclk));
	jor g07534(.dina(w_n7766_0[1]),.dinb(w_asqrt56_28[2]),.dout(n7768),.clk(gclk));
	jxor g07535(.dina(w_n7339_0[0]),.dinb(w_n743_48[0]),.dout(n7769),.clk(gclk));
	jand g07536(.dina(n7769),.dinb(w_asqrt30_29[1]),.dout(n7770),.clk(gclk));
	jxor g07537(.dina(n7770),.dinb(w_n7344_0[0]),.dout(n7771),.clk(gclk));
	jnot g07538(.din(w_n7771_0[1]),.dout(n7772),.clk(gclk));
	jand g07539(.dina(w_n7772_0[1]),.dinb(n7768),.dout(n7773),.clk(gclk));
	jor g07540(.dina(n7773),.dinb(w_n7767_0[1]),.dout(n7774),.clk(gclk));
	jand g07541(.dina(w_n7774_0[2]),.dinb(w_asqrt57_28[2]),.dout(n7775),.clk(gclk));
	jor g07542(.dina(w_n7774_0[1]),.dinb(w_asqrt57_28[1]),.dout(n7776),.clk(gclk));
	jxor g07543(.dina(w_n7346_0[0]),.dinb(w_n635_48[0]),.dout(n7777),.clk(gclk));
	jand g07544(.dina(n7777),.dinb(w_asqrt30_29[0]),.dout(n7778),.clk(gclk));
	jxor g07545(.dina(n7778),.dinb(w_n7351_0[0]),.dout(n7779),.clk(gclk));
	jand g07546(.dina(w_n7779_0[1]),.dinb(n7776),.dout(n7780),.clk(gclk));
	jor g07547(.dina(n7780),.dinb(w_n7775_0[1]),.dout(n7781),.clk(gclk));
	jand g07548(.dina(w_n7781_0[2]),.dinb(w_asqrt58_29[1]),.dout(n7782),.clk(gclk));
	jor g07549(.dina(w_n7781_0[1]),.dinb(w_asqrt58_29[0]),.dout(n7783),.clk(gclk));
	jxor g07550(.dina(w_n7354_0[0]),.dinb(w_n515_49[0]),.dout(n7784),.clk(gclk));
	jand g07551(.dina(n7784),.dinb(w_asqrt30_28[2]),.dout(n7785),.clk(gclk));
	jxor g07552(.dina(n7785),.dinb(w_n7359_0[0]),.dout(n7786),.clk(gclk));
	jand g07553(.dina(w_n7786_0[1]),.dinb(n7783),.dout(n7787),.clk(gclk));
	jor g07554(.dina(n7787),.dinb(w_n7782_0[1]),.dout(n7788),.clk(gclk));
	jand g07555(.dina(w_n7788_0[2]),.dinb(w_asqrt59_29[0]),.dout(n7789),.clk(gclk));
	jor g07556(.dina(w_n7788_0[1]),.dinb(w_asqrt59_28[2]),.dout(n7790),.clk(gclk));
	jxor g07557(.dina(w_n7362_0[0]),.dinb(w_n443_49[0]),.dout(n7791),.clk(gclk));
	jand g07558(.dina(n7791),.dinb(w_asqrt30_28[1]),.dout(n7792),.clk(gclk));
	jxor g07559(.dina(n7792),.dinb(w_n7367_0[0]),.dout(n7793),.clk(gclk));
	jnot g07560(.din(w_n7793_0[1]),.dout(n7794),.clk(gclk));
	jand g07561(.dina(w_n7794_0[1]),.dinb(n7790),.dout(n7795),.clk(gclk));
	jor g07562(.dina(n7795),.dinb(w_n7789_0[1]),.dout(n7796),.clk(gclk));
	jand g07563(.dina(w_n7796_0[2]),.dinb(w_asqrt60_29[1]),.dout(n7797),.clk(gclk));
	jor g07564(.dina(w_n7796_0[1]),.dinb(w_asqrt60_29[0]),.dout(n7798),.clk(gclk));
	jxor g07565(.dina(w_n7369_0[0]),.dinb(w_n352_49[1]),.dout(n7799),.clk(gclk));
	jand g07566(.dina(n7799),.dinb(w_asqrt30_28[0]),.dout(n7800),.clk(gclk));
	jxor g07567(.dina(n7800),.dinb(w_n7374_0[0]),.dout(n7801),.clk(gclk));
	jnot g07568(.din(w_n7801_0[1]),.dout(n7802),.clk(gclk));
	jand g07569(.dina(w_n7802_0[1]),.dinb(n7798),.dout(n7803),.clk(gclk));
	jor g07570(.dina(n7803),.dinb(w_n7797_0[1]),.dout(n7804),.clk(gclk));
	jand g07571(.dina(w_n7804_0[2]),.dinb(w_asqrt61_29[1]),.dout(n7805),.clk(gclk));
	jor g07572(.dina(w_n7804_0[1]),.dinb(w_asqrt61_29[0]),.dout(n7806),.clk(gclk));
	jxor g07573(.dina(w_n7376_0[0]),.dinb(w_n294_49[2]),.dout(n7807),.clk(gclk));
	jand g07574(.dina(n7807),.dinb(w_asqrt30_27[2]),.dout(n7808),.clk(gclk));
	jxor g07575(.dina(n7808),.dinb(w_n7381_0[0]),.dout(n7809),.clk(gclk));
	jnot g07576(.din(w_n7809_0[1]),.dout(n7810),.clk(gclk));
	jand g07577(.dina(w_n7810_0[1]),.dinb(n7806),.dout(n7811),.clk(gclk));
	jor g07578(.dina(n7811),.dinb(w_n7805_0[1]),.dout(n7812),.clk(gclk));
	jand g07579(.dina(w_n7812_0[2]),.dinb(w_asqrt62_29[1]),.dout(n7813),.clk(gclk));
	jor g07580(.dina(w_n7812_0[1]),.dinb(w_asqrt62_29[0]),.dout(n7814),.clk(gclk));
	jxor g07581(.dina(w_n7383_0[0]),.dinb(w_n239_49[2]),.dout(n7815),.clk(gclk));
	jand g07582(.dina(n7815),.dinb(w_asqrt30_27[1]),.dout(n7816),.clk(gclk));
	jxor g07583(.dina(n7816),.dinb(w_n7388_0[0]),.dout(n7817),.clk(gclk));
	jand g07584(.dina(w_n7817_0[2]),.dinb(n7814),.dout(n7818),.clk(gclk));
	jor g07585(.dina(n7818),.dinb(w_n7813_0[1]),.dout(n7819),.clk(gclk));
	jor g07586(.dina(w_n7819_0[1]),.dinb(w_n7419_0[2]),.dout(n7820),.clk(gclk));
	jnot g07587(.din(w_n7820_1[1]),.dout(n7821),.clk(gclk));
	jand g07588(.dina(w_n7581_38[0]),.dinb(w_n7399_0[0]),.dout(n7822),.clk(gclk));
	jnot g07589(.din(n7822),.dout(n7823),.clk(gclk));
	jnot g07590(.din(w_n7408_0[2]),.dout(n7824),.clk(gclk));
	jand g07591(.dina(w_n7403_0[0]),.dinb(w_asqrt63_37[1]),.dout(n7825),.clk(gclk));
	jand g07592(.dina(n7825),.dinb(n7824),.dout(n7826),.clk(gclk));
	jand g07593(.dina(w_n7826_0[1]),.dinb(n7823),.dout(n7827),.clk(gclk));
	jnot g07594(.din(w_n7419_0[1]),.dout(n7828),.clk(gclk));
	jnot g07595(.din(w_n7813_0[0]),.dout(n7829),.clk(gclk));
	jnot g07596(.din(w_n7805_0[0]),.dout(n7830),.clk(gclk));
	jnot g07597(.din(w_n7797_0[0]),.dout(n7831),.clk(gclk));
	jnot g07598(.din(w_n7789_0[0]),.dout(n7832),.clk(gclk));
	jnot g07599(.din(w_n7782_0[0]),.dout(n7833),.clk(gclk));
	jnot g07600(.din(w_n7775_0[0]),.dout(n7834),.clk(gclk));
	jnot g07601(.din(w_n7767_0[0]),.dout(n7835),.clk(gclk));
	jnot g07602(.din(w_n7760_0[0]),.dout(n7836),.clk(gclk));
	jnot g07603(.din(w_n7752_0[0]),.dout(n7837),.clk(gclk));
	jnot g07604(.din(w_n7745_0[0]),.dout(n7838),.clk(gclk));
	jnot g07605(.din(w_n7737_0[0]),.dout(n7839),.clk(gclk));
	jnot g07606(.din(w_n7729_0[0]),.dout(n7840),.clk(gclk));
	jnot g07607(.din(w_n7721_0[0]),.dout(n7841),.clk(gclk));
	jnot g07608(.din(w_n7714_0[0]),.dout(n7842),.clk(gclk));
	jnot g07609(.din(w_n7707_0[0]),.dout(n7843),.clk(gclk));
	jnot g07610(.din(w_n7700_0[0]),.dout(n7844),.clk(gclk));
	jnot g07611(.din(w_n7692_0[0]),.dout(n7845),.clk(gclk));
	jnot g07612(.din(w_n7685_0[0]),.dout(n7846),.clk(gclk));
	jnot g07613(.din(w_n7677_0[0]),.dout(n7847),.clk(gclk));
	jnot g07614(.din(w_n7670_0[0]),.dout(n7848),.clk(gclk));
	jnot g07615(.din(w_n7662_0[0]),.dout(n7849),.clk(gclk));
	jnot g07616(.din(w_n7655_0[0]),.dout(n7850),.clk(gclk));
	jnot g07617(.din(w_n7647_0[0]),.dout(n7851),.clk(gclk));
	jnot g07618(.din(w_n7640_0[0]),.dout(n7852),.clk(gclk));
	jnot g07619(.din(w_n7633_0[0]),.dout(n7853),.clk(gclk));
	jnot g07620(.din(w_n7626_0[0]),.dout(n7854),.clk(gclk));
	jnot g07621(.din(w_n7618_0[0]),.dout(n7855),.clk(gclk));
	jnot g07622(.din(w_n7611_0[0]),.dout(n7856),.clk(gclk));
	jnot g07623(.din(w_n7603_0[0]),.dout(n7857),.clk(gclk));
	jnot g07624(.din(w_n7596_0[0]),.dout(n7858),.clk(gclk));
	jnot g07625(.din(w_n7599_0[0]),.dout(n7859),.clk(gclk));
	jnot g07626(.din(w_n7586_0[0]),.dout(n7860),.clk(gclk));
	jnot g07627(.din(w_n7426_0[0]),.dout(n7861),.clk(gclk));
	jor g07628(.dina(w_n7581_37[2]),.dinb(w_n7156_0[2]),.dout(n7862),.clk(gclk));
	jnot g07629(.din(w_n7424_0[0]),.dout(n7863),.clk(gclk));
	jand g07630(.dina(n7863),.dinb(n7862),.dout(n7864),.clk(gclk));
	jand g07631(.dina(n7864),.dinb(w_n7154_42[0]),.dout(n7865),.clk(gclk));
	jor g07632(.dina(w_n7581_37[1]),.dinb(w_a60_0[0]),.dout(n7866),.clk(gclk));
	jand g07633(.dina(n7866),.dinb(w_a61_0[0]),.dout(n7867),.clk(gclk));
	jand g07634(.dina(w_asqrt30_27[0]),.dinb(w_n7158_0[0]),.dout(n7868),.clk(gclk));
	jor g07635(.dina(n7868),.dinb(n7867),.dout(n7869),.clk(gclk));
	jor g07636(.dina(n7869),.dinb(n7865),.dout(n7870),.clk(gclk));
	jand g07637(.dina(n7870),.dinb(n7861),.dout(n7871),.clk(gclk));
	jand g07638(.dina(n7871),.dinb(w_n6758_37[2]),.dout(n7872),.clk(gclk));
	jor g07639(.dina(w_n7592_0[0]),.dinb(n7872),.dout(n7873),.clk(gclk));
	jand g07640(.dina(n7873),.dinb(n7860),.dout(n7874),.clk(gclk));
	jand g07641(.dina(n7874),.dinb(w_n6357_42[1]),.dout(n7875),.clk(gclk));
	jor g07642(.dina(n7875),.dinb(w_n7859_0[1]),.dout(n7876),.clk(gclk));
	jand g07643(.dina(n7876),.dinb(n7858),.dout(n7877),.clk(gclk));
	jand g07644(.dina(n7877),.dinb(w_n5989_38[1]),.dout(n7878),.clk(gclk));
	jor g07645(.dina(w_n7607_0[0]),.dinb(n7878),.dout(n7879),.clk(gclk));
	jand g07646(.dina(n7879),.dinb(n7857),.dout(n7880),.clk(gclk));
	jand g07647(.dina(n7880),.dinb(w_n5606_42[2]),.dout(n7881),.clk(gclk));
	jnot g07648(.din(w_n7615_0[0]),.dout(n7882),.clk(gclk));
	jor g07649(.dina(w_n7882_0[1]),.dinb(n7881),.dout(n7883),.clk(gclk));
	jand g07650(.dina(n7883),.dinb(n7856),.dout(n7884),.clk(gclk));
	jand g07651(.dina(n7884),.dinb(w_n5259_39[1]),.dout(n7885),.clk(gclk));
	jor g07652(.dina(w_n7622_0[0]),.dinb(n7885),.dout(n7886),.clk(gclk));
	jand g07653(.dina(n7886),.dinb(n7855),.dout(n7887),.clk(gclk));
	jand g07654(.dina(n7887),.dinb(w_n4902_43[1]),.dout(n7888),.clk(gclk));
	jnot g07655(.din(w_n7630_0[0]),.dout(n7889),.clk(gclk));
	jor g07656(.dina(w_n7889_0[1]),.dinb(n7888),.dout(n7890),.clk(gclk));
	jand g07657(.dina(n7890),.dinb(n7854),.dout(n7891),.clk(gclk));
	jand g07658(.dina(n7891),.dinb(w_n4582_40[1]),.dout(n7892),.clk(gclk));
	jnot g07659(.din(w_n7637_0[0]),.dout(n7893),.clk(gclk));
	jor g07660(.dina(w_n7893_0[1]),.dinb(n7892),.dout(n7894),.clk(gclk));
	jand g07661(.dina(n7894),.dinb(n7853),.dout(n7895),.clk(gclk));
	jand g07662(.dina(n7895),.dinb(w_n4249_44[0]),.dout(n7896),.clk(gclk));
	jnot g07663(.din(w_n7644_0[0]),.dout(n7897),.clk(gclk));
	jor g07664(.dina(w_n7897_0[1]),.dinb(n7896),.dout(n7898),.clk(gclk));
	jand g07665(.dina(n7898),.dinb(n7852),.dout(n7899),.clk(gclk));
	jand g07666(.dina(n7899),.dinb(w_n3955_41[0]),.dout(n7900),.clk(gclk));
	jor g07667(.dina(w_n7651_0[0]),.dinb(n7900),.dout(n7901),.clk(gclk));
	jand g07668(.dina(n7901),.dinb(n7851),.dout(n7902),.clk(gclk));
	jand g07669(.dina(n7902),.dinb(w_n3642_44[1]),.dout(n7903),.clk(gclk));
	jnot g07670(.din(w_n7659_0[0]),.dout(n7904),.clk(gclk));
	jor g07671(.dina(w_n7904_0[1]),.dinb(n7903),.dout(n7905),.clk(gclk));
	jand g07672(.dina(n7905),.dinb(n7850),.dout(n7906),.clk(gclk));
	jand g07673(.dina(n7906),.dinb(w_n3368_41[2]),.dout(n7907),.clk(gclk));
	jor g07674(.dina(w_n7666_0[0]),.dinb(n7907),.dout(n7908),.clk(gclk));
	jand g07675(.dina(n7908),.dinb(n7849),.dout(n7909),.clk(gclk));
	jand g07676(.dina(n7909),.dinb(w_n3089_45[0]),.dout(n7910),.clk(gclk));
	jnot g07677(.din(w_n7674_0[0]),.dout(n7911),.clk(gclk));
	jor g07678(.dina(w_n7911_0[1]),.dinb(n7910),.dout(n7912),.clk(gclk));
	jand g07679(.dina(n7912),.dinb(n7848),.dout(n7913),.clk(gclk));
	jand g07680(.dina(n7913),.dinb(w_n2833_42[2]),.dout(n7914),.clk(gclk));
	jor g07681(.dina(w_n7681_0[0]),.dinb(n7914),.dout(n7915),.clk(gclk));
	jand g07682(.dina(n7915),.dinb(n7847),.dout(n7916),.clk(gclk));
	jand g07683(.dina(n7916),.dinb(w_n2572_45[1]),.dout(n7917),.clk(gclk));
	jnot g07684(.din(w_n7689_0[0]),.dout(n7918),.clk(gclk));
	jor g07685(.dina(w_n7918_0[1]),.dinb(n7917),.dout(n7919),.clk(gclk));
	jand g07686(.dina(n7919),.dinb(n7846),.dout(n7920),.clk(gclk));
	jand g07687(.dina(n7920),.dinb(w_n2345_43[1]),.dout(n7921),.clk(gclk));
	jor g07688(.dina(w_n7696_0[0]),.dinb(n7921),.dout(n7922),.clk(gclk));
	jand g07689(.dina(n7922),.dinb(n7845),.dout(n7923),.clk(gclk));
	jand g07690(.dina(n7923),.dinb(w_n2108_46[0]),.dout(n7924),.clk(gclk));
	jnot g07691(.din(w_n7704_0[0]),.dout(n7925),.clk(gclk));
	jor g07692(.dina(w_n7925_0[1]),.dinb(n7924),.dout(n7926),.clk(gclk));
	jand g07693(.dina(n7926),.dinb(n7844),.dout(n7927),.clk(gclk));
	jand g07694(.dina(n7927),.dinb(w_n1912_44[1]),.dout(n7928),.clk(gclk));
	jnot g07695(.din(w_n7711_0[0]),.dout(n7929),.clk(gclk));
	jor g07696(.dina(w_n7929_0[1]),.dinb(n7928),.dout(n7930),.clk(gclk));
	jand g07697(.dina(n7930),.dinb(n7843),.dout(n7931),.clk(gclk));
	jand g07698(.dina(n7931),.dinb(w_n1699_46[2]),.dout(n7932),.clk(gclk));
	jnot g07699(.din(w_n7718_0[0]),.dout(n7933),.clk(gclk));
	jor g07700(.dina(w_n7933_0[1]),.dinb(n7932),.dout(n7934),.clk(gclk));
	jand g07701(.dina(n7934),.dinb(n7842),.dout(n7935),.clk(gclk));
	jand g07702(.dina(n7935),.dinb(w_n1516_45[0]),.dout(n7936),.clk(gclk));
	jor g07703(.dina(w_n7725_0[0]),.dinb(n7936),.dout(n7937),.clk(gclk));
	jand g07704(.dina(n7937),.dinb(n7841),.dout(n7938),.clk(gclk));
	jand g07705(.dina(n7938),.dinb(w_n1332_46[2]),.dout(n7939),.clk(gclk));
	jor g07706(.dina(w_n7733_0[0]),.dinb(n7939),.dout(n7940),.clk(gclk));
	jand g07707(.dina(n7940),.dinb(n7840),.dout(n7941),.clk(gclk));
	jand g07708(.dina(n7941),.dinb(w_n1173_45[2]),.dout(n7942),.clk(gclk));
	jor g07709(.dina(w_n7741_0[0]),.dinb(n7942),.dout(n7943),.clk(gclk));
	jand g07710(.dina(n7943),.dinb(n7839),.dout(n7944),.clk(gclk));
	jand g07711(.dina(n7944),.dinb(w_n1008_47[2]),.dout(n7945),.clk(gclk));
	jnot g07712(.din(w_n7749_0[0]),.dout(n7946),.clk(gclk));
	jor g07713(.dina(w_n7946_0[1]),.dinb(n7945),.dout(n7947),.clk(gclk));
	jand g07714(.dina(n7947),.dinb(n7838),.dout(n7948),.clk(gclk));
	jand g07715(.dina(n7948),.dinb(w_n884_46[2]),.dout(n7949),.clk(gclk));
	jor g07716(.dina(w_n7756_0[0]),.dinb(n7949),.dout(n7950),.clk(gclk));
	jand g07717(.dina(n7950),.dinb(n7837),.dout(n7951),.clk(gclk));
	jand g07718(.dina(n7951),.dinb(w_n743_47[2]),.dout(n7952),.clk(gclk));
	jnot g07719(.din(w_n7764_0[0]),.dout(n7953),.clk(gclk));
	jor g07720(.dina(w_n7953_0[1]),.dinb(n7952),.dout(n7954),.clk(gclk));
	jand g07721(.dina(n7954),.dinb(n7836),.dout(n7955),.clk(gclk));
	jand g07722(.dina(n7955),.dinb(w_n635_47[2]),.dout(n7956),.clk(gclk));
	jor g07723(.dina(w_n7771_0[0]),.dinb(n7956),.dout(n7957),.clk(gclk));
	jand g07724(.dina(n7957),.dinb(n7835),.dout(n7958),.clk(gclk));
	jand g07725(.dina(n7958),.dinb(w_n515_48[2]),.dout(n7959),.clk(gclk));
	jnot g07726(.din(w_n7779_0[0]),.dout(n7960),.clk(gclk));
	jor g07727(.dina(w_n7960_0[1]),.dinb(n7959),.dout(n7961),.clk(gclk));
	jand g07728(.dina(n7961),.dinb(n7834),.dout(n7962),.clk(gclk));
	jand g07729(.dina(n7962),.dinb(w_n443_48[2]),.dout(n7963),.clk(gclk));
	jnot g07730(.din(w_n7786_0[0]),.dout(n7964),.clk(gclk));
	jor g07731(.dina(w_n7964_0[1]),.dinb(n7963),.dout(n7965),.clk(gclk));
	jand g07732(.dina(n7965),.dinb(n7833),.dout(n7966),.clk(gclk));
	jand g07733(.dina(n7966),.dinb(w_n352_49[0]),.dout(n7967),.clk(gclk));
	jor g07734(.dina(w_n7793_0[0]),.dinb(n7967),.dout(n7968),.clk(gclk));
	jand g07735(.dina(n7968),.dinb(n7832),.dout(n7969),.clk(gclk));
	jand g07736(.dina(n7969),.dinb(w_n294_49[1]),.dout(n7970),.clk(gclk));
	jor g07737(.dina(w_n7801_0[0]),.dinb(n7970),.dout(n7971),.clk(gclk));
	jand g07738(.dina(n7971),.dinb(n7831),.dout(n7972),.clk(gclk));
	jand g07739(.dina(n7972),.dinb(w_n239_49[1]),.dout(n7973),.clk(gclk));
	jor g07740(.dina(w_n7809_0[0]),.dinb(n7973),.dout(n7974),.clk(gclk));
	jand g07741(.dina(n7974),.dinb(n7830),.dout(n7975),.clk(gclk));
	jand g07742(.dina(n7975),.dinb(w_n221_49[2]),.dout(n7976),.clk(gclk));
	jnot g07743(.din(w_n7817_0[1]),.dout(n7977),.clk(gclk));
	jor g07744(.dina(n7977),.dinb(n7976),.dout(n7978),.clk(gclk));
	jand g07745(.dina(n7978),.dinb(n7829),.dout(n7979),.clk(gclk));
	jor g07746(.dina(w_n7979_0[1]),.dinb(w_n7828_0[1]),.dout(n7980),.clk(gclk));
	jand g07747(.dina(w_asqrt30_26[2]),.dinb(w_n7576_0[0]),.dout(n7981),.clk(gclk));
	jor g07748(.dina(n7981),.dinb(w_n7408_0[1]),.dout(n7982),.clk(gclk));
	jor g07749(.dina(w_n7982_0[1]),.dinb(w_n7980_0[1]),.dout(n7983),.clk(gclk));
	jand g07750(.dina(n7983),.dinb(w_n218_20[2]),.dout(n7984),.clk(gclk));
	jand g07751(.dina(w_n7581_37[0]),.dinb(w_n7402_0[1]),.dout(n7985),.clk(gclk));
	jor g07752(.dina(w_n7985_0[1]),.dinb(w_n7984_0[1]),.dout(n7986),.clk(gclk));
	jor g07753(.dina(n7986),.dinb(w_n7827_0[1]),.dout(n7987),.clk(gclk));
	jor g07754(.dina(w_n7987_0[1]),.dinb(w_n7821_0[2]),.dout(asqrt_fa_30),.clk(gclk));
	jand g07755(.dina(w_n7819_0[0]),.dinb(w_n7419_0[0]),.dout(n7989),.clk(gclk));
	jand g07756(.dina(w_n7987_0[0]),.dinb(w_n7989_0[1]),.dout(n7990),.clk(gclk));
	jnot g07757(.din(w_a56_0[2]),.dout(n7991),.clk(gclk));
	jnot g07758(.din(w_a57_0[1]),.dout(n7992),.clk(gclk));
	jand g07759(.dina(w_n7992_0[1]),.dinb(w_n7991_1[2]),.dout(n7993),.clk(gclk));
	jand g07760(.dina(w_n7993_0[2]),.dinb(w_n7421_1[1]),.dout(n7994),.clk(gclk));
	jnot g07761(.din(w_n7994_0[1]),.dout(n7995),.clk(gclk));
	jnot g07762(.din(w_n7827_0[0]),.dout(n7996),.clk(gclk));
	jnot g07763(.din(w_n7982_0[0]),.dout(n7997),.clk(gclk));
	jand g07764(.dina(n7997),.dinb(w_n7989_0[0]),.dout(n7998),.clk(gclk));
	jor g07765(.dina(n7998),.dinb(w_asqrt63_37[0]),.dout(n7999),.clk(gclk));
	jnot g07766(.din(w_n7985_0[0]),.dout(n8000),.clk(gclk));
	jand g07767(.dina(n8000),.dinb(n7999),.dout(n8001),.clk(gclk));
	jand g07768(.dina(n8001),.dinb(n7996),.dout(n8002),.clk(gclk));
	jand g07769(.dina(w_n8002_0[1]),.dinb(w_n7820_1[0]),.dout(n8003),.clk(gclk));
	jor g07770(.dina(w_n8003_52[1]),.dinb(w_n7421_1[0]),.dout(n8004),.clk(gclk));
	jand g07771(.dina(n8004),.dinb(n7995),.dout(n8005),.clk(gclk));
	jor g07772(.dina(w_n8005_0[2]),.dinb(w_n7581_36[2]),.dout(n8006),.clk(gclk));
	jand g07773(.dina(w_n8005_0[1]),.dinb(w_n7581_36[1]),.dout(n8007),.clk(gclk));
	jor g07774(.dina(w_n8003_52[0]),.dinb(w_a58_0[1]),.dout(n8008),.clk(gclk));
	jand g07775(.dina(n8008),.dinb(w_a59_0[0]),.dout(n8009),.clk(gclk));
	jand g07776(.dina(w_asqrt29_21[1]),.dinb(w_n7423_0[1]),.dout(n8010),.clk(gclk));
	jor g07777(.dina(n8010),.dinb(n8009),.dout(n8011),.clk(gclk));
	jor g07778(.dina(n8011),.dinb(n8007),.dout(n8012),.clk(gclk));
	jand g07779(.dina(n8012),.dinb(w_n8006_0[1]),.dout(n8013),.clk(gclk));
	jor g07780(.dina(w_n8013_0[2]),.dinb(w_n7154_41[2]),.dout(n8014),.clk(gclk));
	jand g07781(.dina(w_n8013_0[1]),.dinb(w_n7154_41[1]),.dout(n8015),.clk(gclk));
	jnot g07782(.din(w_n7423_0[0]),.dout(n8016),.clk(gclk));
	jor g07783(.dina(w_n8003_51[2]),.dinb(n8016),.dout(n8017),.clk(gclk));
	jor g07784(.dina(w_n7821_0[1]),.dinb(w_n7581_36[0]),.dout(n8018),.clk(gclk));
	jor g07785(.dina(n8018),.dinb(w_n7826_0[0]),.dout(n8019),.clk(gclk));
	jor g07786(.dina(n8019),.dinb(w_n7984_0[0]),.dout(n8020),.clk(gclk));
	jand g07787(.dina(n8020),.dinb(w_n8017_0[1]),.dout(n8021),.clk(gclk));
	jxor g07788(.dina(n8021),.dinb(w_n7156_0[1]),.dout(n8022),.clk(gclk));
	jor g07789(.dina(w_n8022_0[2]),.dinb(n8015),.dout(n8023),.clk(gclk));
	jand g07790(.dina(n8023),.dinb(w_n8014_0[1]),.dout(n8024),.clk(gclk));
	jor g07791(.dina(w_n8024_0[2]),.dinb(w_n6758_37[1]),.dout(n8025),.clk(gclk));
	jand g07792(.dina(w_n8024_0[1]),.dinb(w_n6758_37[0]),.dout(n8026),.clk(gclk));
	jxor g07793(.dina(w_n7425_0[0]),.dinb(w_n7154_41[0]),.dout(n8027),.clk(gclk));
	jor g07794(.dina(n8027),.dinb(w_n8003_51[1]),.dout(n8028),.clk(gclk));
	jxor g07795(.dina(n8028),.dinb(w_n7583_0[0]),.dout(n8029),.clk(gclk));
	jor g07796(.dina(w_n8029_0[2]),.dinb(n8026),.dout(n8030),.clk(gclk));
	jand g07797(.dina(n8030),.dinb(w_n8025_0[1]),.dout(n8031),.clk(gclk));
	jor g07798(.dina(w_n8031_0[2]),.dinb(w_n6357_42[0]),.dout(n8032),.clk(gclk));
	jand g07799(.dina(w_n8031_0[1]),.dinb(w_n6357_41[2]),.dout(n8033),.clk(gclk));
	jxor g07800(.dina(w_n7585_0[0]),.dinb(w_n6758_36[2]),.dout(n8034),.clk(gclk));
	jor g07801(.dina(n8034),.dinb(w_n8003_51[0]),.dout(n8035),.clk(gclk));
	jxor g07802(.dina(n8035),.dinb(w_n7593_0[0]),.dout(n8036),.clk(gclk));
	jor g07803(.dina(w_n8036_0[2]),.dinb(n8033),.dout(n8037),.clk(gclk));
	jand g07804(.dina(n8037),.dinb(w_n8032_0[1]),.dout(n8038),.clk(gclk));
	jor g07805(.dina(w_n8038_0[2]),.dinb(w_n5989_38[0]),.dout(n8039),.clk(gclk));
	jxor g07806(.dina(w_n7595_0[0]),.dinb(w_n6357_41[1]),.dout(n8040),.clk(gclk));
	jor g07807(.dina(n8040),.dinb(w_n8003_50[2]),.dout(n8041),.clk(gclk));
	jxor g07808(.dina(n8041),.dinb(w_n7859_0[0]),.dout(n8042),.clk(gclk));
	jnot g07809(.din(w_n8042_0[2]),.dout(n8043),.clk(gclk));
	jand g07810(.dina(w_n8038_0[1]),.dinb(w_n5989_37[2]),.dout(n8044),.clk(gclk));
	jor g07811(.dina(n8044),.dinb(n8043),.dout(n8045),.clk(gclk));
	jand g07812(.dina(n8045),.dinb(w_n8039_0[1]),.dout(n8046),.clk(gclk));
	jor g07813(.dina(w_n8046_0[2]),.dinb(w_n5606_42[1]),.dout(n8047),.clk(gclk));
	jand g07814(.dina(w_n8046_0[1]),.dinb(w_n5606_42[0]),.dout(n8048),.clk(gclk));
	jxor g07815(.dina(w_n7602_0[0]),.dinb(w_n5989_37[1]),.dout(n8049),.clk(gclk));
	jor g07816(.dina(n8049),.dinb(w_n8003_50[1]),.dout(n8050),.clk(gclk));
	jxor g07817(.dina(n8050),.dinb(w_n7608_0[0]),.dout(n8051),.clk(gclk));
	jor g07818(.dina(w_n8051_0[2]),.dinb(n8048),.dout(n8052),.clk(gclk));
	jand g07819(.dina(n8052),.dinb(w_n8047_0[1]),.dout(n8053),.clk(gclk));
	jor g07820(.dina(w_n8053_0[2]),.dinb(w_n5259_39[0]),.dout(n8054),.clk(gclk));
	jand g07821(.dina(w_n8053_0[1]),.dinb(w_n5259_38[2]),.dout(n8055),.clk(gclk));
	jxor g07822(.dina(w_n7610_0[0]),.dinb(w_n5606_41[2]),.dout(n8056),.clk(gclk));
	jor g07823(.dina(n8056),.dinb(w_n8003_50[0]),.dout(n8057),.clk(gclk));
	jxor g07824(.dina(n8057),.dinb(w_n7882_0[0]),.dout(n8058),.clk(gclk));
	jnot g07825(.din(w_n8058_0[2]),.dout(n8059),.clk(gclk));
	jor g07826(.dina(n8059),.dinb(n8055),.dout(n8060),.clk(gclk));
	jand g07827(.dina(n8060),.dinb(w_n8054_0[1]),.dout(n8061),.clk(gclk));
	jor g07828(.dina(w_n8061_0[2]),.dinb(w_n4902_43[0]),.dout(n8062),.clk(gclk));
	jand g07829(.dina(w_n8061_0[1]),.dinb(w_n4902_42[2]),.dout(n8063),.clk(gclk));
	jxor g07830(.dina(w_n7617_0[0]),.dinb(w_n5259_38[1]),.dout(n8064),.clk(gclk));
	jor g07831(.dina(n8064),.dinb(w_n8003_49[2]),.dout(n8065),.clk(gclk));
	jxor g07832(.dina(n8065),.dinb(w_n7623_0[0]),.dout(n8066),.clk(gclk));
	jor g07833(.dina(w_n8066_0[2]),.dinb(n8063),.dout(n8067),.clk(gclk));
	jand g07834(.dina(n8067),.dinb(w_n8062_0[1]),.dout(n8068),.clk(gclk));
	jor g07835(.dina(w_n8068_0[2]),.dinb(w_n4582_40[0]),.dout(n8069),.clk(gclk));
	jand g07836(.dina(w_n8068_0[1]),.dinb(w_n4582_39[2]),.dout(n8070),.clk(gclk));
	jxor g07837(.dina(w_n7625_0[0]),.dinb(w_n4902_42[1]),.dout(n8071),.clk(gclk));
	jor g07838(.dina(n8071),.dinb(w_n8003_49[1]),.dout(n8072),.clk(gclk));
	jxor g07839(.dina(n8072),.dinb(w_n7889_0[0]),.dout(n8073),.clk(gclk));
	jnot g07840(.din(w_n8073_0[2]),.dout(n8074),.clk(gclk));
	jor g07841(.dina(n8074),.dinb(n8070),.dout(n8075),.clk(gclk));
	jand g07842(.dina(n8075),.dinb(w_n8069_0[1]),.dout(n8076),.clk(gclk));
	jor g07843(.dina(w_n8076_0[2]),.dinb(w_n4249_43[2]),.dout(n8077),.clk(gclk));
	jand g07844(.dina(w_n8076_0[1]),.dinb(w_n4249_43[1]),.dout(n8078),.clk(gclk));
	jxor g07845(.dina(w_n7632_0[0]),.dinb(w_n4582_39[1]),.dout(n8079),.clk(gclk));
	jor g07846(.dina(n8079),.dinb(w_n8003_49[0]),.dout(n8080),.clk(gclk));
	jxor g07847(.dina(n8080),.dinb(w_n7893_0[0]),.dout(n8081),.clk(gclk));
	jnot g07848(.din(w_n8081_0[2]),.dout(n8082),.clk(gclk));
	jor g07849(.dina(n8082),.dinb(n8078),.dout(n8083),.clk(gclk));
	jand g07850(.dina(n8083),.dinb(w_n8077_0[1]),.dout(n8084),.clk(gclk));
	jor g07851(.dina(w_n8084_0[2]),.dinb(w_n3955_40[2]),.dout(n8085),.clk(gclk));
	jand g07852(.dina(w_n8084_0[1]),.dinb(w_n3955_40[1]),.dout(n8086),.clk(gclk));
	jxor g07853(.dina(w_n7639_0[0]),.dinb(w_n4249_43[0]),.dout(n8087),.clk(gclk));
	jor g07854(.dina(n8087),.dinb(w_n8003_48[2]),.dout(n8088),.clk(gclk));
	jxor g07855(.dina(n8088),.dinb(w_n7897_0[0]),.dout(n8089),.clk(gclk));
	jnot g07856(.din(w_n8089_0[2]),.dout(n8090),.clk(gclk));
	jor g07857(.dina(n8090),.dinb(n8086),.dout(n8091),.clk(gclk));
	jand g07858(.dina(n8091),.dinb(w_n8085_0[1]),.dout(n8092),.clk(gclk));
	jor g07859(.dina(w_n8092_0[2]),.dinb(w_n3642_44[0]),.dout(n8093),.clk(gclk));
	jand g07860(.dina(w_n8092_0[1]),.dinb(w_n3642_43[2]),.dout(n8094),.clk(gclk));
	jxor g07861(.dina(w_n7646_0[0]),.dinb(w_n3955_40[0]),.dout(n8095),.clk(gclk));
	jor g07862(.dina(n8095),.dinb(w_n8003_48[1]),.dout(n8096),.clk(gclk));
	jxor g07863(.dina(n8096),.dinb(w_n7652_0[0]),.dout(n8097),.clk(gclk));
	jor g07864(.dina(w_n8097_0[2]),.dinb(n8094),.dout(n8098),.clk(gclk));
	jand g07865(.dina(n8098),.dinb(w_n8093_0[1]),.dout(n8099),.clk(gclk));
	jor g07866(.dina(w_n8099_0[2]),.dinb(w_n3368_41[1]),.dout(n8100),.clk(gclk));
	jand g07867(.dina(w_n8099_0[1]),.dinb(w_n3368_41[0]),.dout(n8101),.clk(gclk));
	jxor g07868(.dina(w_n7654_0[0]),.dinb(w_n3642_43[1]),.dout(n8102),.clk(gclk));
	jor g07869(.dina(n8102),.dinb(w_n8003_48[0]),.dout(n8103),.clk(gclk));
	jxor g07870(.dina(n8103),.dinb(w_n7904_0[0]),.dout(n8104),.clk(gclk));
	jnot g07871(.din(w_n8104_0[2]),.dout(n8105),.clk(gclk));
	jor g07872(.dina(n8105),.dinb(n8101),.dout(n8106),.clk(gclk));
	jand g07873(.dina(n8106),.dinb(w_n8100_0[1]),.dout(n8107),.clk(gclk));
	jor g07874(.dina(w_n8107_0[2]),.dinb(w_n3089_44[2]),.dout(n8108),.clk(gclk));
	jand g07875(.dina(w_n8107_0[1]),.dinb(w_n3089_44[1]),.dout(n8109),.clk(gclk));
	jxor g07876(.dina(w_n7661_0[0]),.dinb(w_n3368_40[2]),.dout(n8110),.clk(gclk));
	jor g07877(.dina(n8110),.dinb(w_n8003_47[2]),.dout(n8111),.clk(gclk));
	jxor g07878(.dina(n8111),.dinb(w_n7667_0[0]),.dout(n8112),.clk(gclk));
	jor g07879(.dina(w_n8112_0[2]),.dinb(n8109),.dout(n8113),.clk(gclk));
	jand g07880(.dina(n8113),.dinb(w_n8108_0[1]),.dout(n8114),.clk(gclk));
	jor g07881(.dina(w_n8114_0[2]),.dinb(w_n2833_42[1]),.dout(n8115),.clk(gclk));
	jand g07882(.dina(w_n8114_0[1]),.dinb(w_n2833_42[0]),.dout(n8116),.clk(gclk));
	jxor g07883(.dina(w_n7669_0[0]),.dinb(w_n3089_44[0]),.dout(n8117),.clk(gclk));
	jor g07884(.dina(n8117),.dinb(w_n8003_47[1]),.dout(n8118),.clk(gclk));
	jxor g07885(.dina(n8118),.dinb(w_n7911_0[0]),.dout(n8119),.clk(gclk));
	jnot g07886(.din(w_n8119_0[2]),.dout(n8120),.clk(gclk));
	jor g07887(.dina(n8120),.dinb(n8116),.dout(n8121),.clk(gclk));
	jand g07888(.dina(n8121),.dinb(w_n8115_0[1]),.dout(n8122),.clk(gclk));
	jor g07889(.dina(w_n8122_0[2]),.dinb(w_n2572_45[0]),.dout(n8123),.clk(gclk));
	jand g07890(.dina(w_n8122_0[1]),.dinb(w_n2572_44[2]),.dout(n8124),.clk(gclk));
	jxor g07891(.dina(w_n7676_0[0]),.dinb(w_n2833_41[2]),.dout(n8125),.clk(gclk));
	jor g07892(.dina(n8125),.dinb(w_n8003_47[0]),.dout(n8126),.clk(gclk));
	jxor g07893(.dina(n8126),.dinb(w_n7682_0[0]),.dout(n8127),.clk(gclk));
	jor g07894(.dina(w_n8127_0[2]),.dinb(n8124),.dout(n8128),.clk(gclk));
	jand g07895(.dina(n8128),.dinb(w_n8123_0[1]),.dout(n8129),.clk(gclk));
	jor g07896(.dina(w_n8129_0[2]),.dinb(w_n2345_43[0]),.dout(n8130),.clk(gclk));
	jand g07897(.dina(w_n8129_0[1]),.dinb(w_n2345_42[2]),.dout(n8131),.clk(gclk));
	jxor g07898(.dina(w_n7684_0[0]),.dinb(w_n2572_44[1]),.dout(n8132),.clk(gclk));
	jor g07899(.dina(n8132),.dinb(w_n8003_46[2]),.dout(n8133),.clk(gclk));
	jxor g07900(.dina(n8133),.dinb(w_n7918_0[0]),.dout(n8134),.clk(gclk));
	jnot g07901(.din(w_n8134_0[2]),.dout(n8135),.clk(gclk));
	jor g07902(.dina(n8135),.dinb(n8131),.dout(n8136),.clk(gclk));
	jand g07903(.dina(n8136),.dinb(w_n8130_0[1]),.dout(n8137),.clk(gclk));
	jor g07904(.dina(w_n8137_0[2]),.dinb(w_n2108_45[2]),.dout(n8138),.clk(gclk));
	jand g07905(.dina(w_n8137_0[1]),.dinb(w_n2108_45[1]),.dout(n8139),.clk(gclk));
	jxor g07906(.dina(w_n7691_0[0]),.dinb(w_n2345_42[1]),.dout(n8140),.clk(gclk));
	jor g07907(.dina(n8140),.dinb(w_n8003_46[1]),.dout(n8141),.clk(gclk));
	jxor g07908(.dina(n8141),.dinb(w_n7697_0[0]),.dout(n8142),.clk(gclk));
	jor g07909(.dina(w_n8142_0[2]),.dinb(n8139),.dout(n8143),.clk(gclk));
	jand g07910(.dina(n8143),.dinb(w_n8138_0[1]),.dout(n8144),.clk(gclk));
	jor g07911(.dina(w_n8144_0[2]),.dinb(w_n1912_44[0]),.dout(n8145),.clk(gclk));
	jand g07912(.dina(w_n8144_0[1]),.dinb(w_n1912_43[2]),.dout(n8146),.clk(gclk));
	jxor g07913(.dina(w_n7699_0[0]),.dinb(w_n2108_45[0]),.dout(n8147),.clk(gclk));
	jor g07914(.dina(n8147),.dinb(w_n8003_46[0]),.dout(n8148),.clk(gclk));
	jxor g07915(.dina(n8148),.dinb(w_n7925_0[0]),.dout(n8149),.clk(gclk));
	jnot g07916(.din(w_n8149_0[2]),.dout(n8150),.clk(gclk));
	jor g07917(.dina(n8150),.dinb(n8146),.dout(n8151),.clk(gclk));
	jand g07918(.dina(n8151),.dinb(w_n8145_0[1]),.dout(n8152),.clk(gclk));
	jor g07919(.dina(w_n8152_0[2]),.dinb(w_n1699_46[1]),.dout(n8153),.clk(gclk));
	jand g07920(.dina(w_n8152_0[1]),.dinb(w_n1699_46[0]),.dout(n8154),.clk(gclk));
	jxor g07921(.dina(w_n7706_0[0]),.dinb(w_n1912_43[1]),.dout(n8155),.clk(gclk));
	jor g07922(.dina(n8155),.dinb(w_n8003_45[2]),.dout(n8156),.clk(gclk));
	jxor g07923(.dina(n8156),.dinb(w_n7929_0[0]),.dout(n8157),.clk(gclk));
	jnot g07924(.din(w_n8157_0[2]),.dout(n8158),.clk(gclk));
	jor g07925(.dina(n8158),.dinb(n8154),.dout(n8159),.clk(gclk));
	jand g07926(.dina(n8159),.dinb(w_n8153_0[1]),.dout(n8160),.clk(gclk));
	jor g07927(.dina(w_n8160_0[2]),.dinb(w_n1516_44[2]),.dout(n8161),.clk(gclk));
	jand g07928(.dina(w_n8160_0[1]),.dinb(w_n1516_44[1]),.dout(n8162),.clk(gclk));
	jxor g07929(.dina(w_n7713_0[0]),.dinb(w_n1699_45[2]),.dout(n8163),.clk(gclk));
	jor g07930(.dina(n8163),.dinb(w_n8003_45[1]),.dout(n8164),.clk(gclk));
	jxor g07931(.dina(n8164),.dinb(w_n7933_0[0]),.dout(n8165),.clk(gclk));
	jnot g07932(.din(w_n8165_0[2]),.dout(n8166),.clk(gclk));
	jor g07933(.dina(n8166),.dinb(n8162),.dout(n8167),.clk(gclk));
	jand g07934(.dina(n8167),.dinb(w_n8161_0[1]),.dout(n8168),.clk(gclk));
	jor g07935(.dina(w_n8168_0[2]),.dinb(w_n1332_46[1]),.dout(n8169),.clk(gclk));
	jand g07936(.dina(w_n8168_0[1]),.dinb(w_n1332_46[0]),.dout(n8170),.clk(gclk));
	jxor g07937(.dina(w_n7720_0[0]),.dinb(w_n1516_44[0]),.dout(n8171),.clk(gclk));
	jor g07938(.dina(n8171),.dinb(w_n8003_45[0]),.dout(n8172),.clk(gclk));
	jxor g07939(.dina(n8172),.dinb(w_n7726_0[0]),.dout(n8173),.clk(gclk));
	jor g07940(.dina(w_n8173_0[2]),.dinb(n8170),.dout(n8174),.clk(gclk));
	jand g07941(.dina(n8174),.dinb(w_n8169_0[1]),.dout(n8175),.clk(gclk));
	jor g07942(.dina(w_n8175_0[2]),.dinb(w_n1173_45[1]),.dout(n8176),.clk(gclk));
	jand g07943(.dina(w_n8175_0[1]),.dinb(w_n1173_45[0]),.dout(n8177),.clk(gclk));
	jxor g07944(.dina(w_n7728_0[0]),.dinb(w_n1332_45[2]),.dout(n8178),.clk(gclk));
	jor g07945(.dina(n8178),.dinb(w_n8003_44[2]),.dout(n8179),.clk(gclk));
	jxor g07946(.dina(n8179),.dinb(w_n7734_0[0]),.dout(n8180),.clk(gclk));
	jor g07947(.dina(w_n8180_0[2]),.dinb(n8177),.dout(n8181),.clk(gclk));
	jand g07948(.dina(n8181),.dinb(w_n8176_0[1]),.dout(n8182),.clk(gclk));
	jor g07949(.dina(w_n8182_0[2]),.dinb(w_n1008_47[1]),.dout(n8183),.clk(gclk));
	jand g07950(.dina(w_n8182_0[1]),.dinb(w_n1008_47[0]),.dout(n8184),.clk(gclk));
	jxor g07951(.dina(w_n7736_0[0]),.dinb(w_n1173_44[2]),.dout(n8185),.clk(gclk));
	jor g07952(.dina(n8185),.dinb(w_n8003_44[1]),.dout(n8186),.clk(gclk));
	jxor g07953(.dina(n8186),.dinb(w_n7742_0[0]),.dout(n8187),.clk(gclk));
	jor g07954(.dina(w_n8187_0[2]),.dinb(n8184),.dout(n8188),.clk(gclk));
	jand g07955(.dina(n8188),.dinb(w_n8183_0[1]),.dout(n8189),.clk(gclk));
	jor g07956(.dina(w_n8189_0[2]),.dinb(w_n884_46[1]),.dout(n8190),.clk(gclk));
	jand g07957(.dina(w_n8189_0[1]),.dinb(w_n884_46[0]),.dout(n8191),.clk(gclk));
	jxor g07958(.dina(w_n7744_0[0]),.dinb(w_n1008_46[2]),.dout(n8192),.clk(gclk));
	jor g07959(.dina(n8192),.dinb(w_n8003_44[0]),.dout(n8193),.clk(gclk));
	jxor g07960(.dina(n8193),.dinb(w_n7946_0[0]),.dout(n8194),.clk(gclk));
	jnot g07961(.din(w_n8194_0[2]),.dout(n8195),.clk(gclk));
	jor g07962(.dina(n8195),.dinb(n8191),.dout(n8196),.clk(gclk));
	jand g07963(.dina(n8196),.dinb(w_n8190_0[1]),.dout(n8197),.clk(gclk));
	jor g07964(.dina(w_n8197_0[2]),.dinb(w_n743_47[1]),.dout(n8198),.clk(gclk));
	jand g07965(.dina(w_n8197_0[1]),.dinb(w_n743_47[0]),.dout(n8199),.clk(gclk));
	jxor g07966(.dina(w_n7751_0[0]),.dinb(w_n884_45[2]),.dout(n8200),.clk(gclk));
	jor g07967(.dina(n8200),.dinb(w_n8003_43[2]),.dout(n8201),.clk(gclk));
	jxor g07968(.dina(n8201),.dinb(w_n7757_0[0]),.dout(n8202),.clk(gclk));
	jor g07969(.dina(w_n8202_0[2]),.dinb(n8199),.dout(n8203),.clk(gclk));
	jand g07970(.dina(n8203),.dinb(w_n8198_0[1]),.dout(n8204),.clk(gclk));
	jor g07971(.dina(w_n8204_0[2]),.dinb(w_n635_47[1]),.dout(n8205),.clk(gclk));
	jand g07972(.dina(w_n8204_0[1]),.dinb(w_n635_47[0]),.dout(n8206),.clk(gclk));
	jxor g07973(.dina(w_n7759_0[0]),.dinb(w_n743_46[2]),.dout(n8207),.clk(gclk));
	jor g07974(.dina(n8207),.dinb(w_n8003_43[1]),.dout(n8208),.clk(gclk));
	jxor g07975(.dina(n8208),.dinb(w_n7953_0[0]),.dout(n8209),.clk(gclk));
	jnot g07976(.din(w_n8209_0[2]),.dout(n8210),.clk(gclk));
	jor g07977(.dina(n8210),.dinb(n8206),.dout(n8211),.clk(gclk));
	jand g07978(.dina(n8211),.dinb(w_n8205_0[1]),.dout(n8212),.clk(gclk));
	jor g07979(.dina(w_n8212_0[2]),.dinb(w_n515_48[1]),.dout(n8213),.clk(gclk));
	jand g07980(.dina(w_n8212_0[1]),.dinb(w_n515_48[0]),.dout(n8214),.clk(gclk));
	jxor g07981(.dina(w_n7766_0[0]),.dinb(w_n635_46[2]),.dout(n8215),.clk(gclk));
	jor g07982(.dina(n8215),.dinb(w_n8003_43[0]),.dout(n8216),.clk(gclk));
	jxor g07983(.dina(n8216),.dinb(w_n7772_0[0]),.dout(n8217),.clk(gclk));
	jor g07984(.dina(w_n8217_0[2]),.dinb(n8214),.dout(n8218),.clk(gclk));
	jand g07985(.dina(n8218),.dinb(w_n8213_0[1]),.dout(n8219),.clk(gclk));
	jor g07986(.dina(w_n8219_0[2]),.dinb(w_n443_48[1]),.dout(n8220),.clk(gclk));
	jand g07987(.dina(w_n8219_0[1]),.dinb(w_n443_48[0]),.dout(n8221),.clk(gclk));
	jxor g07988(.dina(w_n7774_0[0]),.dinb(w_n515_47[2]),.dout(n8222),.clk(gclk));
	jor g07989(.dina(n8222),.dinb(w_n8003_42[2]),.dout(n8223),.clk(gclk));
	jxor g07990(.dina(n8223),.dinb(w_n7960_0[0]),.dout(n8224),.clk(gclk));
	jnot g07991(.din(w_n8224_0[2]),.dout(n8225),.clk(gclk));
	jor g07992(.dina(n8225),.dinb(n8221),.dout(n8226),.clk(gclk));
	jand g07993(.dina(n8226),.dinb(w_n8220_0[1]),.dout(n8227),.clk(gclk));
	jor g07994(.dina(w_n8227_0[2]),.dinb(w_n352_48[2]),.dout(n8228),.clk(gclk));
	jand g07995(.dina(w_n8227_0[1]),.dinb(w_n352_48[1]),.dout(n8229),.clk(gclk));
	jxor g07996(.dina(w_n7781_0[0]),.dinb(w_n443_47[2]),.dout(n8230),.clk(gclk));
	jor g07997(.dina(n8230),.dinb(w_n8003_42[1]),.dout(n8231),.clk(gclk));
	jxor g07998(.dina(n8231),.dinb(w_n7964_0[0]),.dout(n8232),.clk(gclk));
	jnot g07999(.din(w_n8232_0[2]),.dout(n8233),.clk(gclk));
	jor g08000(.dina(n8233),.dinb(n8229),.dout(n8234),.clk(gclk));
	jand g08001(.dina(n8234),.dinb(w_n8228_0[1]),.dout(n8235),.clk(gclk));
	jor g08002(.dina(w_n8235_0[2]),.dinb(w_n294_49[0]),.dout(n8236),.clk(gclk));
	jand g08003(.dina(w_n8235_0[1]),.dinb(w_n294_48[2]),.dout(n8237),.clk(gclk));
	jxor g08004(.dina(w_n7788_0[0]),.dinb(w_n352_48[0]),.dout(n8238),.clk(gclk));
	jor g08005(.dina(n8238),.dinb(w_n8003_42[0]),.dout(n8239),.clk(gclk));
	jxor g08006(.dina(n8239),.dinb(w_n7794_0[0]),.dout(n8240),.clk(gclk));
	jor g08007(.dina(w_n8240_0[2]),.dinb(n8237),.dout(n8241),.clk(gclk));
	jand g08008(.dina(n8241),.dinb(w_n8236_0[1]),.dout(n8242),.clk(gclk));
	jor g08009(.dina(w_n8242_0[2]),.dinb(w_n239_49[0]),.dout(n8243),.clk(gclk));
	jand g08010(.dina(w_n8242_0[1]),.dinb(w_n239_48[2]),.dout(n8244),.clk(gclk));
	jxor g08011(.dina(w_n7796_0[0]),.dinb(w_n294_48[1]),.dout(n8245),.clk(gclk));
	jor g08012(.dina(n8245),.dinb(w_n8003_41[2]),.dout(n8246),.clk(gclk));
	jxor g08013(.dina(n8246),.dinb(w_n7802_0[0]),.dout(n8247),.clk(gclk));
	jor g08014(.dina(w_n8247_0[2]),.dinb(n8244),.dout(n8248),.clk(gclk));
	jand g08015(.dina(n8248),.dinb(w_n8243_0[1]),.dout(n8249),.clk(gclk));
	jor g08016(.dina(w_n8249_0[2]),.dinb(w_n221_49[1]),.dout(n8250),.clk(gclk));
	jand g08017(.dina(w_n8249_0[1]),.dinb(w_n221_49[0]),.dout(n8251),.clk(gclk));
	jxor g08018(.dina(w_n7804_0[0]),.dinb(w_n239_48[1]),.dout(n8252),.clk(gclk));
	jor g08019(.dina(n8252),.dinb(w_n8003_41[1]),.dout(n8253),.clk(gclk));
	jxor g08020(.dina(n8253),.dinb(w_n7810_0[0]),.dout(n8254),.clk(gclk));
	jor g08021(.dina(w_n8254_0[1]),.dinb(n8251),.dout(n8255),.clk(gclk));
	jand g08022(.dina(n8255),.dinb(w_n8250_0[1]),.dout(n8256),.clk(gclk));
	jxor g08023(.dina(w_n7812_0[0]),.dinb(w_n221_48[2]),.dout(n8257),.clk(gclk));
	jor g08024(.dina(n8257),.dinb(w_n8003_41[0]),.dout(n8258),.clk(gclk));
	jxor g08025(.dina(n8258),.dinb(w_n7817_0[0]),.dout(n8259),.clk(gclk));
	jor g08026(.dina(w_n8259_0[2]),.dinb(w_n8256_0[2]),.dout(n8260),.clk(gclk));
	jor g08027(.dina(w_n8260_0[1]),.dinb(w_n7821_0[0]),.dout(n8261),.clk(gclk));
	jor g08028(.dina(n8261),.dinb(w_n7990_0[1]),.dout(n8262),.clk(gclk));
	jand g08029(.dina(n8262),.dinb(w_n218_20[1]),.dout(n8263),.clk(gclk));
	jand g08030(.dina(w_n8003_40[2]),.dinb(w_n7828_0[0]),.dout(n8264),.clk(gclk));
	jand g08031(.dina(w_n8259_0[1]),.dinb(w_n8256_0[1]),.dout(n8265),.clk(gclk));
	jor g08032(.dina(w_n8265_1[1]),.dinb(n8264),.dout(n8266),.clk(gclk));
	jand g08033(.dina(w_n8002_0[0]),.dinb(w_n7979_0[0]),.dout(n8267),.clk(gclk));
	jnot g08034(.din(n8267),.dout(n8268),.clk(gclk));
	jand g08035(.dina(w_n7980_0[0]),.dinb(w_asqrt63_36[2]),.dout(n8269),.clk(gclk));
	jand g08036(.dina(n8269),.dinb(w_n7820_0[2]),.dout(n8270),.clk(gclk));
	jand g08037(.dina(w_n8270_0[1]),.dinb(n8268),.dout(n8271),.clk(gclk));
	jor g08038(.dina(n8271),.dinb(n8266),.dout(n8272),.clk(gclk));
	jor g08039(.dina(w_n8272_0[1]),.dinb(w_n8263_0[1]),.dout(asqrt_fa_29),.clk(gclk));
	jnot g08040(.din(w_n8254_0[0]),.dout(n8274),.clk(gclk));
	jxor g08041(.dina(w_n8249_0[0]),.dinb(w_n221_48[1]),.dout(n8275),.clk(gclk));
	jand g08042(.dina(n8275),.dinb(w_asqrt28_37[1]),.dout(n8276),.clk(gclk));
	jxor g08043(.dina(n8276),.dinb(w_n8274_0[1]),.dout(n8277),.clk(gclk));
	jand g08044(.dina(w_asqrt28_37[0]),.dinb(w_a56_0[1]),.dout(n8278),.clk(gclk));
	jnot g08045(.din(w_a54_1[1]),.dout(n8279),.clk(gclk));
	jnot g08046(.din(w_a55_0[1]),.dout(n8280),.clk(gclk));
	jand g08047(.dina(w_n8280_0[1]),.dinb(w_n8279_1[1]),.dout(n8281),.clk(gclk));
	jand g08048(.dina(w_n8281_0[2]),.dinb(w_n7991_1[1]),.dout(n8282),.clk(gclk));
	jor g08049(.dina(w_n8282_0[1]),.dinb(n8278),.dout(n8283),.clk(gclk));
	jand g08050(.dina(w_n8283_0[2]),.dinb(w_asqrt29_21[0]),.dout(n8284),.clk(gclk));
	jor g08051(.dina(w_n8283_0[1]),.dinb(w_asqrt29_20[2]),.dout(n8285),.clk(gclk));
	jand g08052(.dina(w_asqrt28_36[2]),.dinb(w_n7991_1[0]),.dout(n8286),.clk(gclk));
	jor g08053(.dina(n8286),.dinb(w_n7992_0[0]),.dout(n8287),.clk(gclk));
	jnot g08054(.din(w_n7993_0[1]),.dout(n8288),.clk(gclk));
	jnot g08055(.din(w_n7990_0[0]),.dout(n8289),.clk(gclk));
	jnot g08056(.din(w_n8250_0[0]),.dout(n8290),.clk(gclk));
	jnot g08057(.din(w_n8243_0[0]),.dout(n8291),.clk(gclk));
	jnot g08058(.din(w_n8236_0[0]),.dout(n8292),.clk(gclk));
	jnot g08059(.din(w_n8228_0[0]),.dout(n8293),.clk(gclk));
	jnot g08060(.din(w_n8220_0[0]),.dout(n8294),.clk(gclk));
	jnot g08061(.din(w_n8213_0[0]),.dout(n8295),.clk(gclk));
	jnot g08062(.din(w_n8205_0[0]),.dout(n8296),.clk(gclk));
	jnot g08063(.din(w_n8198_0[0]),.dout(n8297),.clk(gclk));
	jnot g08064(.din(w_n8190_0[0]),.dout(n8298),.clk(gclk));
	jnot g08065(.din(w_n8183_0[0]),.dout(n8299),.clk(gclk));
	jnot g08066(.din(w_n8176_0[0]),.dout(n8300),.clk(gclk));
	jnot g08067(.din(w_n8169_0[0]),.dout(n8301),.clk(gclk));
	jnot g08068(.din(w_n8161_0[0]),.dout(n8302),.clk(gclk));
	jnot g08069(.din(w_n8153_0[0]),.dout(n8303),.clk(gclk));
	jnot g08070(.din(w_n8145_0[0]),.dout(n8304),.clk(gclk));
	jnot g08071(.din(w_n8138_0[0]),.dout(n8305),.clk(gclk));
	jnot g08072(.din(w_n8130_0[0]),.dout(n8306),.clk(gclk));
	jnot g08073(.din(w_n8123_0[0]),.dout(n8307),.clk(gclk));
	jnot g08074(.din(w_n8115_0[0]),.dout(n8308),.clk(gclk));
	jnot g08075(.din(w_n8108_0[0]),.dout(n8309),.clk(gclk));
	jnot g08076(.din(w_n8100_0[0]),.dout(n8310),.clk(gclk));
	jnot g08077(.din(w_n8093_0[0]),.dout(n8311),.clk(gclk));
	jnot g08078(.din(w_n8085_0[0]),.dout(n8312),.clk(gclk));
	jnot g08079(.din(w_n8077_0[0]),.dout(n8313),.clk(gclk));
	jnot g08080(.din(w_n8069_0[0]),.dout(n8314),.clk(gclk));
	jnot g08081(.din(w_n8062_0[0]),.dout(n8315),.clk(gclk));
	jnot g08082(.din(w_n8054_0[0]),.dout(n8316),.clk(gclk));
	jnot g08083(.din(w_n8047_0[0]),.dout(n8317),.clk(gclk));
	jnot g08084(.din(w_n8039_0[0]),.dout(n8318),.clk(gclk));
	jnot g08085(.din(w_n8032_0[0]),.dout(n8319),.clk(gclk));
	jnot g08086(.din(w_n8025_0[0]),.dout(n8320),.clk(gclk));
	jnot g08087(.din(w_n8014_0[0]),.dout(n8321),.clk(gclk));
	jnot g08088(.din(w_n8006_0[0]),.dout(n8322),.clk(gclk));
	jand g08089(.dina(w_asqrt29_20[1]),.dinb(w_a58_0[0]),.dout(n8323),.clk(gclk));
	jor g08090(.dina(n8323),.dinb(w_n7994_0[0]),.dout(n8324),.clk(gclk));
	jor g08091(.dina(n8324),.dinb(w_asqrt30_26[1]),.dout(n8325),.clk(gclk));
	jand g08092(.dina(w_asqrt29_20[0]),.dinb(w_n7421_0[2]),.dout(n8326),.clk(gclk));
	jor g08093(.dina(n8326),.dinb(w_n7422_0[0]),.dout(n8327),.clk(gclk));
	jand g08094(.dina(w_n8017_0[0]),.dinb(n8327),.dout(n8328),.clk(gclk));
	jand g08095(.dina(w_n8328_0[1]),.dinb(n8325),.dout(n8329),.clk(gclk));
	jor g08096(.dina(n8329),.dinb(n8322),.dout(n8330),.clk(gclk));
	jor g08097(.dina(n8330),.dinb(w_asqrt31_21[1]),.dout(n8331),.clk(gclk));
	jnot g08098(.din(w_n8022_0[1]),.dout(n8332),.clk(gclk));
	jand g08099(.dina(n8332),.dinb(n8331),.dout(n8333),.clk(gclk));
	jor g08100(.dina(n8333),.dinb(n8321),.dout(n8334),.clk(gclk));
	jor g08101(.dina(n8334),.dinb(w_asqrt32_26[1]),.dout(n8335),.clk(gclk));
	jnot g08102(.din(w_n8029_0[1]),.dout(n8336),.clk(gclk));
	jand g08103(.dina(n8336),.dinb(n8335),.dout(n8337),.clk(gclk));
	jor g08104(.dina(n8337),.dinb(n8320),.dout(n8338),.clk(gclk));
	jor g08105(.dina(n8338),.dinb(w_asqrt33_22[0]),.dout(n8339),.clk(gclk));
	jnot g08106(.din(w_n8036_0[1]),.dout(n8340),.clk(gclk));
	jand g08107(.dina(n8340),.dinb(n8339),.dout(n8341),.clk(gclk));
	jor g08108(.dina(n8341),.dinb(n8319),.dout(n8342),.clk(gclk));
	jor g08109(.dina(n8342),.dinb(w_asqrt34_26[2]),.dout(n8343),.clk(gclk));
	jand g08110(.dina(n8343),.dinb(w_n8042_0[1]),.dout(n8344),.clk(gclk));
	jor g08111(.dina(n8344),.dinb(n8318),.dout(n8345),.clk(gclk));
	jor g08112(.dina(n8345),.dinb(w_asqrt35_22[2]),.dout(n8346),.clk(gclk));
	jnot g08113(.din(w_n8051_0[1]),.dout(n8347),.clk(gclk));
	jand g08114(.dina(n8347),.dinb(n8346),.dout(n8348),.clk(gclk));
	jor g08115(.dina(n8348),.dinb(n8317),.dout(n8349),.clk(gclk));
	jor g08116(.dina(n8349),.dinb(w_asqrt36_26[2]),.dout(n8350),.clk(gclk));
	jand g08117(.dina(w_n8058_0[1]),.dinb(n8350),.dout(n8351),.clk(gclk));
	jor g08118(.dina(n8351),.dinb(n8316),.dout(n8352),.clk(gclk));
	jor g08119(.dina(n8352),.dinb(w_asqrt37_23[0]),.dout(n8353),.clk(gclk));
	jnot g08120(.din(w_n8066_0[1]),.dout(n8354),.clk(gclk));
	jand g08121(.dina(n8354),.dinb(n8353),.dout(n8355),.clk(gclk));
	jor g08122(.dina(n8355),.dinb(n8315),.dout(n8356),.clk(gclk));
	jor g08123(.dina(n8356),.dinb(w_asqrt38_27[0]),.dout(n8357),.clk(gclk));
	jand g08124(.dina(w_n8073_0[1]),.dinb(n8357),.dout(n8358),.clk(gclk));
	jor g08125(.dina(n8358),.dinb(n8314),.dout(n8359),.clk(gclk));
	jor g08126(.dina(n8359),.dinb(w_asqrt39_23[2]),.dout(n8360),.clk(gclk));
	jand g08127(.dina(w_n8081_0[1]),.dinb(n8360),.dout(n8361),.clk(gclk));
	jor g08128(.dina(n8361),.dinb(n8313),.dout(n8362),.clk(gclk));
	jor g08129(.dina(n8362),.dinb(w_asqrt40_27[0]),.dout(n8363),.clk(gclk));
	jand g08130(.dina(w_n8089_0[1]),.dinb(n8363),.dout(n8364),.clk(gclk));
	jor g08131(.dina(n8364),.dinb(n8312),.dout(n8365),.clk(gclk));
	jor g08132(.dina(n8365),.dinb(w_asqrt41_24[0]),.dout(n8366),.clk(gclk));
	jnot g08133(.din(w_n8097_0[1]),.dout(n8367),.clk(gclk));
	jand g08134(.dina(n8367),.dinb(n8366),.dout(n8368),.clk(gclk));
	jor g08135(.dina(n8368),.dinb(n8311),.dout(n8369),.clk(gclk));
	jor g08136(.dina(n8369),.dinb(w_asqrt42_27[1]),.dout(n8370),.clk(gclk));
	jand g08137(.dina(w_n8104_0[1]),.dinb(n8370),.dout(n8371),.clk(gclk));
	jor g08138(.dina(n8371),.dinb(n8310),.dout(n8372),.clk(gclk));
	jor g08139(.dina(n8372),.dinb(w_asqrt43_24[1]),.dout(n8373),.clk(gclk));
	jnot g08140(.din(w_n8112_0[1]),.dout(n8374),.clk(gclk));
	jand g08141(.dina(n8374),.dinb(n8373),.dout(n8375),.clk(gclk));
	jor g08142(.dina(n8375),.dinb(n8309),.dout(n8376),.clk(gclk));
	jor g08143(.dina(n8376),.dinb(w_asqrt44_27[1]),.dout(n8377),.clk(gclk));
	jand g08144(.dina(w_n8119_0[1]),.dinb(n8377),.dout(n8378),.clk(gclk));
	jor g08145(.dina(n8378),.dinb(n8308),.dout(n8379),.clk(gclk));
	jor g08146(.dina(n8379),.dinb(w_asqrt45_25[0]),.dout(n8380),.clk(gclk));
	jnot g08147(.din(w_n8127_0[1]),.dout(n8381),.clk(gclk));
	jand g08148(.dina(n8381),.dinb(n8380),.dout(n8382),.clk(gclk));
	jor g08149(.dina(n8382),.dinb(n8307),.dout(n8383),.clk(gclk));
	jor g08150(.dina(n8383),.dinb(w_asqrt46_27[1]),.dout(n8384),.clk(gclk));
	jand g08151(.dina(w_n8134_0[1]),.dinb(n8384),.dout(n8385),.clk(gclk));
	jor g08152(.dina(n8385),.dinb(n8306),.dout(n8386),.clk(gclk));
	jor g08153(.dina(n8386),.dinb(w_asqrt47_25[2]),.dout(n8387),.clk(gclk));
	jnot g08154(.din(w_n8142_0[1]),.dout(n8388),.clk(gclk));
	jand g08155(.dina(n8388),.dinb(n8387),.dout(n8389),.clk(gclk));
	jor g08156(.dina(n8389),.dinb(n8305),.dout(n8390),.clk(gclk));
	jor g08157(.dina(n8390),.dinb(w_asqrt48_27[2]),.dout(n8391),.clk(gclk));
	jand g08158(.dina(w_n8149_0[1]),.dinb(n8391),.dout(n8392),.clk(gclk));
	jor g08159(.dina(n8392),.dinb(n8304),.dout(n8393),.clk(gclk));
	jor g08160(.dina(n8393),.dinb(w_asqrt49_26[0]),.dout(n8394),.clk(gclk));
	jand g08161(.dina(w_n8157_0[1]),.dinb(n8394),.dout(n8395),.clk(gclk));
	jor g08162(.dina(n8395),.dinb(n8303),.dout(n8396),.clk(gclk));
	jor g08163(.dina(n8396),.dinb(w_asqrt50_28[0]),.dout(n8397),.clk(gclk));
	jand g08164(.dina(w_n8165_0[1]),.dinb(n8397),.dout(n8398),.clk(gclk));
	jor g08165(.dina(n8398),.dinb(n8302),.dout(n8399),.clk(gclk));
	jor g08166(.dina(n8399),.dinb(w_asqrt51_26[1]),.dout(n8400),.clk(gclk));
	jnot g08167(.din(w_n8173_0[1]),.dout(n8401),.clk(gclk));
	jand g08168(.dina(n8401),.dinb(n8400),.dout(n8402),.clk(gclk));
	jor g08169(.dina(n8402),.dinb(n8301),.dout(n8403),.clk(gclk));
	jor g08170(.dina(n8403),.dinb(w_asqrt52_28[0]),.dout(n8404),.clk(gclk));
	jnot g08171(.din(w_n8180_0[1]),.dout(n8405),.clk(gclk));
	jand g08172(.dina(n8405),.dinb(n8404),.dout(n8406),.clk(gclk));
	jor g08173(.dina(n8406),.dinb(n8300),.dout(n8407),.clk(gclk));
	jor g08174(.dina(n8407),.dinb(w_asqrt53_27[0]),.dout(n8408),.clk(gclk));
	jnot g08175(.din(w_n8187_0[1]),.dout(n8409),.clk(gclk));
	jand g08176(.dina(n8409),.dinb(n8408),.dout(n8410),.clk(gclk));
	jor g08177(.dina(n8410),.dinb(n8299),.dout(n8411),.clk(gclk));
	jor g08178(.dina(n8411),.dinb(w_asqrt54_28[0]),.dout(n8412),.clk(gclk));
	jand g08179(.dina(w_n8194_0[1]),.dinb(n8412),.dout(n8413),.clk(gclk));
	jor g08180(.dina(n8413),.dinb(n8298),.dout(n8414),.clk(gclk));
	jor g08181(.dina(n8414),.dinb(w_asqrt55_27[1]),.dout(n8415),.clk(gclk));
	jnot g08182(.din(w_n8202_0[1]),.dout(n8416),.clk(gclk));
	jand g08183(.dina(n8416),.dinb(n8415),.dout(n8417),.clk(gclk));
	jor g08184(.dina(n8417),.dinb(n8297),.dout(n8418),.clk(gclk));
	jor g08185(.dina(n8418),.dinb(w_asqrt56_28[1]),.dout(n8419),.clk(gclk));
	jand g08186(.dina(w_n8209_0[1]),.dinb(n8419),.dout(n8420),.clk(gclk));
	jor g08187(.dina(n8420),.dinb(n8296),.dout(n8421),.clk(gclk));
	jor g08188(.dina(n8421),.dinb(w_asqrt57_28[0]),.dout(n8422),.clk(gclk));
	jnot g08189(.din(w_n8217_0[1]),.dout(n8423),.clk(gclk));
	jand g08190(.dina(n8423),.dinb(n8422),.dout(n8424),.clk(gclk));
	jor g08191(.dina(n8424),.dinb(n8295),.dout(n8425),.clk(gclk));
	jor g08192(.dina(n8425),.dinb(w_asqrt58_28[2]),.dout(n8426),.clk(gclk));
	jand g08193(.dina(w_n8224_0[1]),.dinb(n8426),.dout(n8427),.clk(gclk));
	jor g08194(.dina(n8427),.dinb(n8294),.dout(n8428),.clk(gclk));
	jor g08195(.dina(n8428),.dinb(w_asqrt59_28[1]),.dout(n8429),.clk(gclk));
	jand g08196(.dina(w_n8232_0[1]),.dinb(n8429),.dout(n8430),.clk(gclk));
	jor g08197(.dina(n8430),.dinb(n8293),.dout(n8431),.clk(gclk));
	jor g08198(.dina(n8431),.dinb(w_asqrt60_28[2]),.dout(n8432),.clk(gclk));
	jnot g08199(.din(w_n8240_0[1]),.dout(n8433),.clk(gclk));
	jand g08200(.dina(n8433),.dinb(n8432),.dout(n8434),.clk(gclk));
	jor g08201(.dina(n8434),.dinb(n8292),.dout(n8435),.clk(gclk));
	jor g08202(.dina(n8435),.dinb(w_asqrt61_28[2]),.dout(n8436),.clk(gclk));
	jnot g08203(.din(w_n8247_0[1]),.dout(n8437),.clk(gclk));
	jand g08204(.dina(n8437),.dinb(n8436),.dout(n8438),.clk(gclk));
	jor g08205(.dina(n8438),.dinb(n8291),.dout(n8439),.clk(gclk));
	jor g08206(.dina(n8439),.dinb(w_asqrt62_28[2]),.dout(n8440),.clk(gclk));
	jand g08207(.dina(w_n8274_0[0]),.dinb(n8440),.dout(n8441),.clk(gclk));
	jor g08208(.dina(n8441),.dinb(n8290),.dout(n8442),.clk(gclk));
	jnot g08209(.din(w_n8259_0[0]),.dout(n8443),.clk(gclk));
	jand g08210(.dina(n8443),.dinb(n8442),.dout(n8444),.clk(gclk));
	jand g08211(.dina(w_n8444_0[1]),.dinb(w_n7820_0[1]),.dout(n8445),.clk(gclk));
	jand g08212(.dina(n8445),.dinb(n8289),.dout(n8446),.clk(gclk));
	jor g08213(.dina(n8446),.dinb(w_asqrt63_36[1]),.dout(n8447),.clk(gclk));
	jnot g08214(.din(w_n8272_0[0]),.dout(n8448),.clk(gclk));
	jand g08215(.dina(n8448),.dinb(n8447),.dout(n8449),.clk(gclk));
	jor g08216(.dina(w_n8449_35[1]),.dinb(n8288),.dout(n8450),.clk(gclk));
	jand g08217(.dina(w_n8450_0[1]),.dinb(n8287),.dout(n8451),.clk(gclk));
	jand g08218(.dina(n8451),.dinb(n8285),.dout(n8452),.clk(gclk));
	jor g08219(.dina(n8452),.dinb(w_n8284_0[1]),.dout(n8453),.clk(gclk));
	jand g08220(.dina(w_n8453_0[2]),.dinb(w_asqrt30_26[0]),.dout(n8454),.clk(gclk));
	jor g08221(.dina(w_n8453_0[1]),.dinb(w_asqrt30_25[2]),.dout(n8455),.clk(gclk));
	jor g08222(.dina(w_n8270_0[0]),.dinb(w_n8265_1[0]),.dout(n8456),.clk(gclk));
	jor g08223(.dina(n8456),.dinb(w_n8263_0[0]),.dout(n8457),.clk(gclk));
	jor g08224(.dina(n8457),.dinb(w_n8003_40[1]),.dout(n8458),.clk(gclk));
	jand g08225(.dina(n8458),.dinb(w_n8450_0[0]),.dout(n8459),.clk(gclk));
	jxor g08226(.dina(n8459),.dinb(w_n7421_0[1]),.dout(n8460),.clk(gclk));
	jnot g08227(.din(w_n8460_0[1]),.dout(n8461),.clk(gclk));
	jand g08228(.dina(w_n8461_0[1]),.dinb(n8455),.dout(n8462),.clk(gclk));
	jor g08229(.dina(n8462),.dinb(w_n8454_0[1]),.dout(n8463),.clk(gclk));
	jand g08230(.dina(w_n8463_0[2]),.dinb(w_asqrt31_21[0]),.dout(n8464),.clk(gclk));
	jor g08231(.dina(w_n8463_0[1]),.dinb(w_asqrt31_20[2]),.dout(n8465),.clk(gclk));
	jxor g08232(.dina(w_n8005_0[0]),.dinb(w_n7581_35[2]),.dout(n8466),.clk(gclk));
	jand g08233(.dina(n8466),.dinb(w_asqrt28_36[1]),.dout(n8467),.clk(gclk));
	jxor g08234(.dina(n8467),.dinb(w_n8328_0[0]),.dout(n8468),.clk(gclk));
	jand g08235(.dina(w_n8468_0[2]),.dinb(n8465),.dout(n8469),.clk(gclk));
	jor g08236(.dina(n8469),.dinb(w_n8464_0[1]),.dout(n8470),.clk(gclk));
	jand g08237(.dina(w_n8470_0[2]),.dinb(w_asqrt32_26[0]),.dout(n8471),.clk(gclk));
	jor g08238(.dina(w_n8470_0[1]),.dinb(w_asqrt32_25[2]),.dout(n8472),.clk(gclk));
	jxor g08239(.dina(w_n8013_0[0]),.dinb(w_n7154_40[2]),.dout(n8473),.clk(gclk));
	jand g08240(.dina(n8473),.dinb(w_asqrt28_36[0]),.dout(n8474),.clk(gclk));
	jxor g08241(.dina(n8474),.dinb(w_n8022_0[0]),.dout(n8475),.clk(gclk));
	jnot g08242(.din(w_n8475_0[1]),.dout(n8476),.clk(gclk));
	jand g08243(.dina(w_n8476_0[1]),.dinb(n8472),.dout(n8477),.clk(gclk));
	jor g08244(.dina(n8477),.dinb(w_n8471_0[1]),.dout(n8478),.clk(gclk));
	jand g08245(.dina(w_n8478_0[2]),.dinb(w_asqrt33_21[2]),.dout(n8479),.clk(gclk));
	jor g08246(.dina(w_n8478_0[1]),.dinb(w_asqrt33_21[1]),.dout(n8480),.clk(gclk));
	jxor g08247(.dina(w_n8024_0[0]),.dinb(w_n6758_36[1]),.dout(n8481),.clk(gclk));
	jand g08248(.dina(n8481),.dinb(w_asqrt28_35[2]),.dout(n8482),.clk(gclk));
	jxor g08249(.dina(n8482),.dinb(w_n8029_0[0]),.dout(n8483),.clk(gclk));
	jnot g08250(.din(w_n8483_0[1]),.dout(n8484),.clk(gclk));
	jand g08251(.dina(w_n8484_0[1]),.dinb(n8480),.dout(n8485),.clk(gclk));
	jor g08252(.dina(n8485),.dinb(w_n8479_0[1]),.dout(n8486),.clk(gclk));
	jand g08253(.dina(w_n8486_0[2]),.dinb(w_asqrt34_26[1]),.dout(n8487),.clk(gclk));
	jor g08254(.dina(w_n8486_0[1]),.dinb(w_asqrt34_26[0]),.dout(n8488),.clk(gclk));
	jxor g08255(.dina(w_n8031_0[0]),.dinb(w_n6357_41[0]),.dout(n8489),.clk(gclk));
	jand g08256(.dina(n8489),.dinb(w_asqrt28_35[1]),.dout(n8490),.clk(gclk));
	jxor g08257(.dina(n8490),.dinb(w_n8036_0[0]),.dout(n8491),.clk(gclk));
	jnot g08258(.din(w_n8491_0[1]),.dout(n8492),.clk(gclk));
	jand g08259(.dina(w_n8492_0[1]),.dinb(n8488),.dout(n8493),.clk(gclk));
	jor g08260(.dina(n8493),.dinb(w_n8487_0[1]),.dout(n8494),.clk(gclk));
	jand g08261(.dina(w_n8494_0[2]),.dinb(w_asqrt35_22[1]),.dout(n8495),.clk(gclk));
	jxor g08262(.dina(w_n8038_0[0]),.dinb(w_n5989_37[0]),.dout(n8496),.clk(gclk));
	jand g08263(.dina(n8496),.dinb(w_asqrt28_35[0]),.dout(n8497),.clk(gclk));
	jxor g08264(.dina(n8497),.dinb(w_n8042_0[0]),.dout(n8498),.clk(gclk));
	jor g08265(.dina(w_n8494_0[1]),.dinb(w_asqrt35_22[0]),.dout(n8499),.clk(gclk));
	jand g08266(.dina(n8499),.dinb(w_n8498_0[1]),.dout(n8500),.clk(gclk));
	jor g08267(.dina(n8500),.dinb(w_n8495_0[1]),.dout(n8501),.clk(gclk));
	jand g08268(.dina(w_n8501_0[2]),.dinb(w_asqrt36_26[1]),.dout(n8502),.clk(gclk));
	jor g08269(.dina(w_n8501_0[1]),.dinb(w_asqrt36_26[0]),.dout(n8503),.clk(gclk));
	jxor g08270(.dina(w_n8046_0[0]),.dinb(w_n5606_41[1]),.dout(n8504),.clk(gclk));
	jand g08271(.dina(n8504),.dinb(w_asqrt28_34[2]),.dout(n8505),.clk(gclk));
	jxor g08272(.dina(n8505),.dinb(w_n8051_0[0]),.dout(n8506),.clk(gclk));
	jnot g08273(.din(w_n8506_0[1]),.dout(n8507),.clk(gclk));
	jand g08274(.dina(w_n8507_0[1]),.dinb(n8503),.dout(n8508),.clk(gclk));
	jor g08275(.dina(n8508),.dinb(w_n8502_0[1]),.dout(n8509),.clk(gclk));
	jand g08276(.dina(w_n8509_0[2]),.dinb(w_asqrt37_22[2]),.dout(n8510),.clk(gclk));
	jor g08277(.dina(w_n8509_0[1]),.dinb(w_asqrt37_22[1]),.dout(n8511),.clk(gclk));
	jxor g08278(.dina(w_n8053_0[0]),.dinb(w_n5259_38[0]),.dout(n8512),.clk(gclk));
	jand g08279(.dina(n8512),.dinb(w_asqrt28_34[1]),.dout(n8513),.clk(gclk));
	jxor g08280(.dina(n8513),.dinb(w_n8058_0[0]),.dout(n8514),.clk(gclk));
	jand g08281(.dina(w_n8514_0[1]),.dinb(n8511),.dout(n8515),.clk(gclk));
	jor g08282(.dina(n8515),.dinb(w_n8510_0[1]),.dout(n8516),.clk(gclk));
	jand g08283(.dina(w_n8516_0[2]),.dinb(w_asqrt38_26[2]),.dout(n8517),.clk(gclk));
	jor g08284(.dina(w_n8516_0[1]),.dinb(w_asqrt38_26[1]),.dout(n8518),.clk(gclk));
	jxor g08285(.dina(w_n8061_0[0]),.dinb(w_n4902_42[0]),.dout(n8519),.clk(gclk));
	jand g08286(.dina(n8519),.dinb(w_asqrt28_34[0]),.dout(n8520),.clk(gclk));
	jxor g08287(.dina(n8520),.dinb(w_n8066_0[0]),.dout(n8521),.clk(gclk));
	jnot g08288(.din(w_n8521_0[1]),.dout(n8522),.clk(gclk));
	jand g08289(.dina(w_n8522_0[1]),.dinb(n8518),.dout(n8523),.clk(gclk));
	jor g08290(.dina(n8523),.dinb(w_n8517_0[1]),.dout(n8524),.clk(gclk));
	jand g08291(.dina(w_n8524_0[2]),.dinb(w_asqrt39_23[1]),.dout(n8525),.clk(gclk));
	jor g08292(.dina(w_n8524_0[1]),.dinb(w_asqrt39_23[0]),.dout(n8526),.clk(gclk));
	jxor g08293(.dina(w_n8068_0[0]),.dinb(w_n4582_39[0]),.dout(n8527),.clk(gclk));
	jand g08294(.dina(n8527),.dinb(w_asqrt28_33[2]),.dout(n8528),.clk(gclk));
	jxor g08295(.dina(n8528),.dinb(w_n8073_0[0]),.dout(n8529),.clk(gclk));
	jand g08296(.dina(w_n8529_0[1]),.dinb(n8526),.dout(n8530),.clk(gclk));
	jor g08297(.dina(n8530),.dinb(w_n8525_0[1]),.dout(n8531),.clk(gclk));
	jand g08298(.dina(w_n8531_0[2]),.dinb(w_asqrt40_26[2]),.dout(n8532),.clk(gclk));
	jor g08299(.dina(w_n8531_0[1]),.dinb(w_asqrt40_26[1]),.dout(n8533),.clk(gclk));
	jxor g08300(.dina(w_n8076_0[0]),.dinb(w_n4249_42[2]),.dout(n8534),.clk(gclk));
	jand g08301(.dina(n8534),.dinb(w_asqrt28_33[1]),.dout(n8535),.clk(gclk));
	jxor g08302(.dina(n8535),.dinb(w_n8081_0[0]),.dout(n8536),.clk(gclk));
	jand g08303(.dina(w_n8536_0[1]),.dinb(n8533),.dout(n8537),.clk(gclk));
	jor g08304(.dina(n8537),.dinb(w_n8532_0[1]),.dout(n8538),.clk(gclk));
	jand g08305(.dina(w_n8538_0[2]),.dinb(w_asqrt41_23[2]),.dout(n8539),.clk(gclk));
	jor g08306(.dina(w_n8538_0[1]),.dinb(w_asqrt41_23[1]),.dout(n8540),.clk(gclk));
	jxor g08307(.dina(w_n8084_0[0]),.dinb(w_n3955_39[2]),.dout(n8541),.clk(gclk));
	jand g08308(.dina(n8541),.dinb(w_asqrt28_33[0]),.dout(n8542),.clk(gclk));
	jxor g08309(.dina(n8542),.dinb(w_n8089_0[0]),.dout(n8543),.clk(gclk));
	jand g08310(.dina(w_n8543_0[1]),.dinb(n8540),.dout(n8544),.clk(gclk));
	jor g08311(.dina(n8544),.dinb(w_n8539_0[1]),.dout(n8545),.clk(gclk));
	jand g08312(.dina(w_n8545_0[2]),.dinb(w_asqrt42_27[0]),.dout(n8546),.clk(gclk));
	jor g08313(.dina(w_n8545_0[1]),.dinb(w_asqrt42_26[2]),.dout(n8547),.clk(gclk));
	jxor g08314(.dina(w_n8092_0[0]),.dinb(w_n3642_43[0]),.dout(n8548),.clk(gclk));
	jand g08315(.dina(n8548),.dinb(w_asqrt28_32[2]),.dout(n8549),.clk(gclk));
	jxor g08316(.dina(n8549),.dinb(w_n8097_0[0]),.dout(n8550),.clk(gclk));
	jnot g08317(.din(w_n8550_0[1]),.dout(n8551),.clk(gclk));
	jand g08318(.dina(w_n8551_0[1]),.dinb(n8547),.dout(n8552),.clk(gclk));
	jor g08319(.dina(n8552),.dinb(w_n8546_0[1]),.dout(n8553),.clk(gclk));
	jand g08320(.dina(w_n8553_0[2]),.dinb(w_asqrt43_24[0]),.dout(n8554),.clk(gclk));
	jor g08321(.dina(w_n8553_0[1]),.dinb(w_asqrt43_23[2]),.dout(n8555),.clk(gclk));
	jxor g08322(.dina(w_n8099_0[0]),.dinb(w_n3368_40[1]),.dout(n8556),.clk(gclk));
	jand g08323(.dina(n8556),.dinb(w_asqrt28_32[1]),.dout(n8557),.clk(gclk));
	jxor g08324(.dina(n8557),.dinb(w_n8104_0[0]),.dout(n8558),.clk(gclk));
	jand g08325(.dina(w_n8558_0[1]),.dinb(n8555),.dout(n8559),.clk(gclk));
	jor g08326(.dina(n8559),.dinb(w_n8554_0[1]),.dout(n8560),.clk(gclk));
	jand g08327(.dina(w_n8560_0[2]),.dinb(w_asqrt44_27[0]),.dout(n8561),.clk(gclk));
	jor g08328(.dina(w_n8560_0[1]),.dinb(w_asqrt44_26[2]),.dout(n8562),.clk(gclk));
	jxor g08329(.dina(w_n8107_0[0]),.dinb(w_n3089_43[2]),.dout(n8563),.clk(gclk));
	jand g08330(.dina(n8563),.dinb(w_asqrt28_32[0]),.dout(n8564),.clk(gclk));
	jxor g08331(.dina(n8564),.dinb(w_n8112_0[0]),.dout(n8565),.clk(gclk));
	jnot g08332(.din(w_n8565_0[1]),.dout(n8566),.clk(gclk));
	jand g08333(.dina(w_n8566_0[1]),.dinb(n8562),.dout(n8567),.clk(gclk));
	jor g08334(.dina(n8567),.dinb(w_n8561_0[1]),.dout(n8568),.clk(gclk));
	jand g08335(.dina(w_n8568_0[2]),.dinb(w_asqrt45_24[2]),.dout(n8569),.clk(gclk));
	jor g08336(.dina(w_n8568_0[1]),.dinb(w_asqrt45_24[1]),.dout(n8570),.clk(gclk));
	jxor g08337(.dina(w_n8114_0[0]),.dinb(w_n2833_41[1]),.dout(n8571),.clk(gclk));
	jand g08338(.dina(n8571),.dinb(w_asqrt28_31[2]),.dout(n8572),.clk(gclk));
	jxor g08339(.dina(n8572),.dinb(w_n8119_0[0]),.dout(n8573),.clk(gclk));
	jand g08340(.dina(w_n8573_0[1]),.dinb(n8570),.dout(n8574),.clk(gclk));
	jor g08341(.dina(n8574),.dinb(w_n8569_0[1]),.dout(n8575),.clk(gclk));
	jand g08342(.dina(w_n8575_0[2]),.dinb(w_asqrt46_27[0]),.dout(n8576),.clk(gclk));
	jor g08343(.dina(w_n8575_0[1]),.dinb(w_asqrt46_26[2]),.dout(n8577),.clk(gclk));
	jxor g08344(.dina(w_n8122_0[0]),.dinb(w_n2572_44[0]),.dout(n8578),.clk(gclk));
	jand g08345(.dina(n8578),.dinb(w_asqrt28_31[1]),.dout(n8579),.clk(gclk));
	jxor g08346(.dina(n8579),.dinb(w_n8127_0[0]),.dout(n8580),.clk(gclk));
	jnot g08347(.din(w_n8580_0[1]),.dout(n8581),.clk(gclk));
	jand g08348(.dina(w_n8581_0[1]),.dinb(n8577),.dout(n8582),.clk(gclk));
	jor g08349(.dina(n8582),.dinb(w_n8576_0[1]),.dout(n8583),.clk(gclk));
	jand g08350(.dina(w_n8583_0[2]),.dinb(w_asqrt47_25[1]),.dout(n8584),.clk(gclk));
	jor g08351(.dina(w_n8583_0[1]),.dinb(w_asqrt47_25[0]),.dout(n8585),.clk(gclk));
	jxor g08352(.dina(w_n8129_0[0]),.dinb(w_n2345_42[0]),.dout(n8586),.clk(gclk));
	jand g08353(.dina(n8586),.dinb(w_asqrt28_31[0]),.dout(n8587),.clk(gclk));
	jxor g08354(.dina(n8587),.dinb(w_n8134_0[0]),.dout(n8588),.clk(gclk));
	jand g08355(.dina(w_n8588_0[1]),.dinb(n8585),.dout(n8589),.clk(gclk));
	jor g08356(.dina(n8589),.dinb(w_n8584_0[1]),.dout(n8590),.clk(gclk));
	jand g08357(.dina(w_n8590_0[2]),.dinb(w_asqrt48_27[1]),.dout(n8591),.clk(gclk));
	jor g08358(.dina(w_n8590_0[1]),.dinb(w_asqrt48_27[0]),.dout(n8592),.clk(gclk));
	jxor g08359(.dina(w_n8137_0[0]),.dinb(w_n2108_44[2]),.dout(n8593),.clk(gclk));
	jand g08360(.dina(n8593),.dinb(w_asqrt28_30[2]),.dout(n8594),.clk(gclk));
	jxor g08361(.dina(n8594),.dinb(w_n8142_0[0]),.dout(n8595),.clk(gclk));
	jnot g08362(.din(w_n8595_0[1]),.dout(n8596),.clk(gclk));
	jand g08363(.dina(w_n8596_0[1]),.dinb(n8592),.dout(n8597),.clk(gclk));
	jor g08364(.dina(n8597),.dinb(w_n8591_0[1]),.dout(n8598),.clk(gclk));
	jand g08365(.dina(w_n8598_0[2]),.dinb(w_asqrt49_25[2]),.dout(n8599),.clk(gclk));
	jor g08366(.dina(w_n8598_0[1]),.dinb(w_asqrt49_25[1]),.dout(n8600),.clk(gclk));
	jxor g08367(.dina(w_n8144_0[0]),.dinb(w_n1912_43[0]),.dout(n8601),.clk(gclk));
	jand g08368(.dina(n8601),.dinb(w_asqrt28_30[1]),.dout(n8602),.clk(gclk));
	jxor g08369(.dina(n8602),.dinb(w_n8149_0[0]),.dout(n8603),.clk(gclk));
	jand g08370(.dina(w_n8603_0[1]),.dinb(n8600),.dout(n8604),.clk(gclk));
	jor g08371(.dina(n8604),.dinb(w_n8599_0[1]),.dout(n8605),.clk(gclk));
	jand g08372(.dina(w_n8605_0[2]),.dinb(w_asqrt50_27[2]),.dout(n8606),.clk(gclk));
	jor g08373(.dina(w_n8605_0[1]),.dinb(w_asqrt50_27[1]),.dout(n8607),.clk(gclk));
	jxor g08374(.dina(w_n8152_0[0]),.dinb(w_n1699_45[1]),.dout(n8608),.clk(gclk));
	jand g08375(.dina(n8608),.dinb(w_asqrt28_30[0]),.dout(n8609),.clk(gclk));
	jxor g08376(.dina(n8609),.dinb(w_n8157_0[0]),.dout(n8610),.clk(gclk));
	jand g08377(.dina(w_n8610_0[1]),.dinb(n8607),.dout(n8611),.clk(gclk));
	jor g08378(.dina(n8611),.dinb(w_n8606_0[1]),.dout(n8612),.clk(gclk));
	jand g08379(.dina(w_n8612_0[2]),.dinb(w_asqrt51_26[0]),.dout(n8613),.clk(gclk));
	jor g08380(.dina(w_n8612_0[1]),.dinb(w_asqrt51_25[2]),.dout(n8614),.clk(gclk));
	jxor g08381(.dina(w_n8160_0[0]),.dinb(w_n1516_43[2]),.dout(n8615),.clk(gclk));
	jand g08382(.dina(n8615),.dinb(w_asqrt28_29[2]),.dout(n8616),.clk(gclk));
	jxor g08383(.dina(n8616),.dinb(w_n8165_0[0]),.dout(n8617),.clk(gclk));
	jand g08384(.dina(w_n8617_0[1]),.dinb(n8614),.dout(n8618),.clk(gclk));
	jor g08385(.dina(n8618),.dinb(w_n8613_0[1]),.dout(n8619),.clk(gclk));
	jand g08386(.dina(w_n8619_0[2]),.dinb(w_asqrt52_27[2]),.dout(n8620),.clk(gclk));
	jor g08387(.dina(w_n8619_0[1]),.dinb(w_asqrt52_27[1]),.dout(n8621),.clk(gclk));
	jxor g08388(.dina(w_n8168_0[0]),.dinb(w_n1332_45[1]),.dout(n8622),.clk(gclk));
	jand g08389(.dina(n8622),.dinb(w_asqrt28_29[1]),.dout(n8623),.clk(gclk));
	jxor g08390(.dina(n8623),.dinb(w_n8173_0[0]),.dout(n8624),.clk(gclk));
	jnot g08391(.din(w_n8624_0[1]),.dout(n8625),.clk(gclk));
	jand g08392(.dina(w_n8625_0[1]),.dinb(n8621),.dout(n8626),.clk(gclk));
	jor g08393(.dina(n8626),.dinb(w_n8620_0[1]),.dout(n8627),.clk(gclk));
	jand g08394(.dina(w_n8627_0[2]),.dinb(w_asqrt53_26[2]),.dout(n8628),.clk(gclk));
	jor g08395(.dina(w_n8627_0[1]),.dinb(w_asqrt53_26[1]),.dout(n8629),.clk(gclk));
	jxor g08396(.dina(w_n8175_0[0]),.dinb(w_n1173_44[1]),.dout(n8630),.clk(gclk));
	jand g08397(.dina(n8630),.dinb(w_asqrt28_29[0]),.dout(n8631),.clk(gclk));
	jxor g08398(.dina(n8631),.dinb(w_n8180_0[0]),.dout(n8632),.clk(gclk));
	jnot g08399(.din(w_n8632_0[1]),.dout(n8633),.clk(gclk));
	jand g08400(.dina(w_n8633_0[1]),.dinb(n8629),.dout(n8634),.clk(gclk));
	jor g08401(.dina(n8634),.dinb(w_n8628_0[1]),.dout(n8635),.clk(gclk));
	jand g08402(.dina(w_n8635_0[2]),.dinb(w_asqrt54_27[2]),.dout(n8636),.clk(gclk));
	jor g08403(.dina(w_n8635_0[1]),.dinb(w_asqrt54_27[1]),.dout(n8637),.clk(gclk));
	jxor g08404(.dina(w_n8182_0[0]),.dinb(w_n1008_46[1]),.dout(n8638),.clk(gclk));
	jand g08405(.dina(n8638),.dinb(w_asqrt28_28[2]),.dout(n8639),.clk(gclk));
	jxor g08406(.dina(n8639),.dinb(w_n8187_0[0]),.dout(n8640),.clk(gclk));
	jnot g08407(.din(w_n8640_0[1]),.dout(n8641),.clk(gclk));
	jand g08408(.dina(w_n8641_0[1]),.dinb(n8637),.dout(n8642),.clk(gclk));
	jor g08409(.dina(n8642),.dinb(w_n8636_0[1]),.dout(n8643),.clk(gclk));
	jand g08410(.dina(w_n8643_0[2]),.dinb(w_asqrt55_27[0]),.dout(n8644),.clk(gclk));
	jor g08411(.dina(w_n8643_0[1]),.dinb(w_asqrt55_26[2]),.dout(n8645),.clk(gclk));
	jxor g08412(.dina(w_n8189_0[0]),.dinb(w_n884_45[1]),.dout(n8646),.clk(gclk));
	jand g08413(.dina(n8646),.dinb(w_asqrt28_28[1]),.dout(n8647),.clk(gclk));
	jxor g08414(.dina(n8647),.dinb(w_n8194_0[0]),.dout(n8648),.clk(gclk));
	jand g08415(.dina(w_n8648_0[1]),.dinb(n8645),.dout(n8649),.clk(gclk));
	jor g08416(.dina(n8649),.dinb(w_n8644_0[1]),.dout(n8650),.clk(gclk));
	jand g08417(.dina(w_n8650_0[2]),.dinb(w_asqrt56_28[0]),.dout(n8651),.clk(gclk));
	jor g08418(.dina(w_n8650_0[1]),.dinb(w_asqrt56_27[2]),.dout(n8652),.clk(gclk));
	jxor g08419(.dina(w_n8197_0[0]),.dinb(w_n743_46[1]),.dout(n8653),.clk(gclk));
	jand g08420(.dina(n8653),.dinb(w_asqrt28_28[0]),.dout(n8654),.clk(gclk));
	jxor g08421(.dina(n8654),.dinb(w_n8202_0[0]),.dout(n8655),.clk(gclk));
	jnot g08422(.din(w_n8655_0[1]),.dout(n8656),.clk(gclk));
	jand g08423(.dina(w_n8656_0[1]),.dinb(n8652),.dout(n8657),.clk(gclk));
	jor g08424(.dina(n8657),.dinb(w_n8651_0[1]),.dout(n8658),.clk(gclk));
	jand g08425(.dina(w_n8658_0[2]),.dinb(w_asqrt57_27[2]),.dout(n8659),.clk(gclk));
	jor g08426(.dina(w_n8658_0[1]),.dinb(w_asqrt57_27[1]),.dout(n8660),.clk(gclk));
	jxor g08427(.dina(w_n8204_0[0]),.dinb(w_n635_46[1]),.dout(n8661),.clk(gclk));
	jand g08428(.dina(n8661),.dinb(w_asqrt28_27[2]),.dout(n8662),.clk(gclk));
	jxor g08429(.dina(n8662),.dinb(w_n8209_0[0]),.dout(n8663),.clk(gclk));
	jand g08430(.dina(w_n8663_0[1]),.dinb(n8660),.dout(n8664),.clk(gclk));
	jor g08431(.dina(n8664),.dinb(w_n8659_0[1]),.dout(n8665),.clk(gclk));
	jand g08432(.dina(w_n8665_0[2]),.dinb(w_asqrt58_28[1]),.dout(n8666),.clk(gclk));
	jor g08433(.dina(w_n8665_0[1]),.dinb(w_asqrt58_28[0]),.dout(n8667),.clk(gclk));
	jxor g08434(.dina(w_n8212_0[0]),.dinb(w_n515_47[1]),.dout(n8668),.clk(gclk));
	jand g08435(.dina(n8668),.dinb(w_asqrt28_27[1]),.dout(n8669),.clk(gclk));
	jxor g08436(.dina(n8669),.dinb(w_n8217_0[0]),.dout(n8670),.clk(gclk));
	jnot g08437(.din(w_n8670_0[1]),.dout(n8671),.clk(gclk));
	jand g08438(.dina(w_n8671_0[1]),.dinb(n8667),.dout(n8672),.clk(gclk));
	jor g08439(.dina(n8672),.dinb(w_n8666_0[1]),.dout(n8673),.clk(gclk));
	jand g08440(.dina(w_n8673_0[2]),.dinb(w_asqrt59_28[0]),.dout(n8674),.clk(gclk));
	jor g08441(.dina(w_n8673_0[1]),.dinb(w_asqrt59_27[2]),.dout(n8675),.clk(gclk));
	jxor g08442(.dina(w_n8219_0[0]),.dinb(w_n443_47[1]),.dout(n8676),.clk(gclk));
	jand g08443(.dina(n8676),.dinb(w_asqrt28_27[0]),.dout(n8677),.clk(gclk));
	jxor g08444(.dina(n8677),.dinb(w_n8224_0[0]),.dout(n8678),.clk(gclk));
	jand g08445(.dina(w_n8678_0[1]),.dinb(n8675),.dout(n8679),.clk(gclk));
	jor g08446(.dina(n8679),.dinb(w_n8674_0[1]),.dout(n8680),.clk(gclk));
	jand g08447(.dina(w_n8680_0[2]),.dinb(w_asqrt60_28[1]),.dout(n8681),.clk(gclk));
	jor g08448(.dina(w_n8680_0[1]),.dinb(w_asqrt60_28[0]),.dout(n8682),.clk(gclk));
	jxor g08449(.dina(w_n8227_0[0]),.dinb(w_n352_47[2]),.dout(n8683),.clk(gclk));
	jand g08450(.dina(n8683),.dinb(w_asqrt28_26[2]),.dout(n8684),.clk(gclk));
	jxor g08451(.dina(n8684),.dinb(w_n8232_0[0]),.dout(n8685),.clk(gclk));
	jand g08452(.dina(w_n8685_0[1]),.dinb(n8682),.dout(n8686),.clk(gclk));
	jor g08453(.dina(n8686),.dinb(w_n8681_0[1]),.dout(n8687),.clk(gclk));
	jand g08454(.dina(w_n8687_0[2]),.dinb(w_asqrt61_28[1]),.dout(n8688),.clk(gclk));
	jor g08455(.dina(w_n8687_0[1]),.dinb(w_asqrt61_28[0]),.dout(n8689),.clk(gclk));
	jxor g08456(.dina(w_n8235_0[0]),.dinb(w_n294_48[0]),.dout(n8690),.clk(gclk));
	jand g08457(.dina(n8690),.dinb(w_asqrt28_26[1]),.dout(n8691),.clk(gclk));
	jxor g08458(.dina(n8691),.dinb(w_n8240_0[0]),.dout(n8692),.clk(gclk));
	jnot g08459(.din(w_n8692_0[1]),.dout(n8693),.clk(gclk));
	jand g08460(.dina(w_n8693_0[1]),.dinb(n8689),.dout(n8694),.clk(gclk));
	jor g08461(.dina(n8694),.dinb(w_n8688_0[1]),.dout(n8695),.clk(gclk));
	jand g08462(.dina(w_n8695_0[2]),.dinb(w_asqrt62_28[1]),.dout(n8696),.clk(gclk));
	jor g08463(.dina(w_n8695_0[1]),.dinb(w_asqrt62_28[0]),.dout(n8697),.clk(gclk));
	jxor g08464(.dina(w_n8242_0[0]),.dinb(w_n239_48[0]),.dout(n8698),.clk(gclk));
	jand g08465(.dina(n8698),.dinb(w_asqrt28_26[0]),.dout(n8699),.clk(gclk));
	jxor g08466(.dina(n8699),.dinb(w_n8247_0[0]),.dout(n8700),.clk(gclk));
	jnot g08467(.din(w_n8700_0[2]),.dout(n8701),.clk(gclk));
	jand g08468(.dina(n8701),.dinb(n8697),.dout(n8702),.clk(gclk));
	jor g08469(.dina(n8702),.dinb(w_n8696_0[1]),.dout(n8703),.clk(gclk));
	jor g08470(.dina(w_n8703_0[1]),.dinb(w_n8277_0[2]),.dout(n8704),.clk(gclk));
	jnot g08471(.din(w_n8704_0[2]),.dout(n8705),.clk(gclk));
	jnot g08472(.din(w_n8277_0[1]),.dout(n8707),.clk(gclk));
	jnot g08473(.din(w_n8696_0[0]),.dout(n8708),.clk(gclk));
	jnot g08474(.din(w_n8688_0[0]),.dout(n8709),.clk(gclk));
	jnot g08475(.din(w_n8681_0[0]),.dout(n8710),.clk(gclk));
	jnot g08476(.din(w_n8674_0[0]),.dout(n8711),.clk(gclk));
	jnot g08477(.din(w_n8666_0[0]),.dout(n8712),.clk(gclk));
	jnot g08478(.din(w_n8659_0[0]),.dout(n8713),.clk(gclk));
	jnot g08479(.din(w_n8651_0[0]),.dout(n8714),.clk(gclk));
	jnot g08480(.din(w_n8644_0[0]),.dout(n8715),.clk(gclk));
	jnot g08481(.din(w_n8636_0[0]),.dout(n8716),.clk(gclk));
	jnot g08482(.din(w_n8628_0[0]),.dout(n8717),.clk(gclk));
	jnot g08483(.din(w_n8620_0[0]),.dout(n8718),.clk(gclk));
	jnot g08484(.din(w_n8613_0[0]),.dout(n8719),.clk(gclk));
	jnot g08485(.din(w_n8606_0[0]),.dout(n8720),.clk(gclk));
	jnot g08486(.din(w_n8599_0[0]),.dout(n8721),.clk(gclk));
	jnot g08487(.din(w_n8591_0[0]),.dout(n8722),.clk(gclk));
	jnot g08488(.din(w_n8584_0[0]),.dout(n8723),.clk(gclk));
	jnot g08489(.din(w_n8576_0[0]),.dout(n8724),.clk(gclk));
	jnot g08490(.din(w_n8569_0[0]),.dout(n8725),.clk(gclk));
	jnot g08491(.din(w_n8561_0[0]),.dout(n8726),.clk(gclk));
	jnot g08492(.din(w_n8554_0[0]),.dout(n8727),.clk(gclk));
	jnot g08493(.din(w_n8546_0[0]),.dout(n8728),.clk(gclk));
	jnot g08494(.din(w_n8539_0[0]),.dout(n8729),.clk(gclk));
	jnot g08495(.din(w_n8532_0[0]),.dout(n8730),.clk(gclk));
	jnot g08496(.din(w_n8525_0[0]),.dout(n8731),.clk(gclk));
	jnot g08497(.din(w_n8517_0[0]),.dout(n8732),.clk(gclk));
	jnot g08498(.din(w_n8510_0[0]),.dout(n8733),.clk(gclk));
	jnot g08499(.din(w_n8502_0[0]),.dout(n8734),.clk(gclk));
	jnot g08500(.din(w_n8495_0[0]),.dout(n8735),.clk(gclk));
	jnot g08501(.din(w_n8498_0[0]),.dout(n8736),.clk(gclk));
	jnot g08502(.din(w_n8487_0[0]),.dout(n8737),.clk(gclk));
	jnot g08503(.din(w_n8479_0[0]),.dout(n8738),.clk(gclk));
	jnot g08504(.din(w_n8471_0[0]),.dout(n8739),.clk(gclk));
	jnot g08505(.din(w_n8464_0[0]),.dout(n8740),.clk(gclk));
	jnot g08506(.din(w_n8454_0[0]),.dout(n8741),.clk(gclk));
	jnot g08507(.din(w_n8284_0[0]),.dout(n8742),.clk(gclk));
	jor g08508(.dina(w_n8449_35[0]),.dinb(w_n7991_0[2]),.dout(n8743),.clk(gclk));
	jnot g08509(.din(w_n8282_0[0]),.dout(n8744),.clk(gclk));
	jand g08510(.dina(n8744),.dinb(n8743),.dout(n8745),.clk(gclk));
	jand g08511(.dina(n8745),.dinb(w_n8003_40[0]),.dout(n8746),.clk(gclk));
	jor g08512(.dina(w_n8449_34[2]),.dinb(w_a56_0[0]),.dout(n8747),.clk(gclk));
	jand g08513(.dina(n8747),.dinb(w_a57_0[0]),.dout(n8748),.clk(gclk));
	jand g08514(.dina(w_asqrt28_25[2]),.dinb(w_n7993_0[0]),.dout(n8749),.clk(gclk));
	jor g08515(.dina(n8749),.dinb(n8748),.dout(n8750),.clk(gclk));
	jor g08516(.dina(w_n8750_0[1]),.dinb(n8746),.dout(n8751),.clk(gclk));
	jand g08517(.dina(n8751),.dinb(n8742),.dout(n8752),.clk(gclk));
	jand g08518(.dina(n8752),.dinb(w_n7581_35[1]),.dout(n8753),.clk(gclk));
	jor g08519(.dina(w_n8460_0[0]),.dinb(n8753),.dout(n8754),.clk(gclk));
	jand g08520(.dina(n8754),.dinb(n8741),.dout(n8755),.clk(gclk));
	jand g08521(.dina(n8755),.dinb(w_n7154_40[1]),.dout(n8756),.clk(gclk));
	jnot g08522(.din(w_n8468_0[1]),.dout(n8757),.clk(gclk));
	jor g08523(.dina(n8757),.dinb(n8756),.dout(n8758),.clk(gclk));
	jand g08524(.dina(n8758),.dinb(n8740),.dout(n8759),.clk(gclk));
	jand g08525(.dina(n8759),.dinb(w_n6758_36[0]),.dout(n8760),.clk(gclk));
	jor g08526(.dina(w_n8475_0[0]),.dinb(n8760),.dout(n8761),.clk(gclk));
	jand g08527(.dina(n8761),.dinb(n8739),.dout(n8762),.clk(gclk));
	jand g08528(.dina(n8762),.dinb(w_n6357_40[2]),.dout(n8763),.clk(gclk));
	jor g08529(.dina(w_n8483_0[0]),.dinb(n8763),.dout(n8764),.clk(gclk));
	jand g08530(.dina(n8764),.dinb(n8738),.dout(n8765),.clk(gclk));
	jand g08531(.dina(n8765),.dinb(w_n5989_36[2]),.dout(n8766),.clk(gclk));
	jor g08532(.dina(w_n8491_0[0]),.dinb(n8766),.dout(n8767),.clk(gclk));
	jand g08533(.dina(n8767),.dinb(n8737),.dout(n8768),.clk(gclk));
	jand g08534(.dina(n8768),.dinb(w_n5606_41[0]),.dout(n8769),.clk(gclk));
	jor g08535(.dina(n8769),.dinb(w_n8736_0[1]),.dout(n8770),.clk(gclk));
	jand g08536(.dina(n8770),.dinb(n8735),.dout(n8771),.clk(gclk));
	jand g08537(.dina(n8771),.dinb(w_n5259_37[2]),.dout(n8772),.clk(gclk));
	jor g08538(.dina(w_n8506_0[0]),.dinb(n8772),.dout(n8773),.clk(gclk));
	jand g08539(.dina(n8773),.dinb(n8734),.dout(n8774),.clk(gclk));
	jand g08540(.dina(n8774),.dinb(w_n4902_41[2]),.dout(n8775),.clk(gclk));
	jnot g08541(.din(w_n8514_0[0]),.dout(n8776),.clk(gclk));
	jor g08542(.dina(w_n8776_0[1]),.dinb(n8775),.dout(n8777),.clk(gclk));
	jand g08543(.dina(n8777),.dinb(n8733),.dout(n8778),.clk(gclk));
	jand g08544(.dina(n8778),.dinb(w_n4582_38[2]),.dout(n8779),.clk(gclk));
	jor g08545(.dina(w_n8521_0[0]),.dinb(n8779),.dout(n8780),.clk(gclk));
	jand g08546(.dina(n8780),.dinb(n8732),.dout(n8781),.clk(gclk));
	jand g08547(.dina(n8781),.dinb(w_n4249_42[1]),.dout(n8782),.clk(gclk));
	jnot g08548(.din(w_n8529_0[0]),.dout(n8783),.clk(gclk));
	jor g08549(.dina(w_n8783_0[1]),.dinb(n8782),.dout(n8784),.clk(gclk));
	jand g08550(.dina(n8784),.dinb(n8731),.dout(n8785),.clk(gclk));
	jand g08551(.dina(n8785),.dinb(w_n3955_39[1]),.dout(n8786),.clk(gclk));
	jnot g08552(.din(w_n8536_0[0]),.dout(n8787),.clk(gclk));
	jor g08553(.dina(w_n8787_0[1]),.dinb(n8786),.dout(n8788),.clk(gclk));
	jand g08554(.dina(n8788),.dinb(n8730),.dout(n8789),.clk(gclk));
	jand g08555(.dina(n8789),.dinb(w_n3642_42[2]),.dout(n8790),.clk(gclk));
	jnot g08556(.din(w_n8543_0[0]),.dout(n8791),.clk(gclk));
	jor g08557(.dina(w_n8791_0[1]),.dinb(n8790),.dout(n8792),.clk(gclk));
	jand g08558(.dina(n8792),.dinb(n8729),.dout(n8793),.clk(gclk));
	jand g08559(.dina(n8793),.dinb(w_n3368_40[0]),.dout(n8794),.clk(gclk));
	jor g08560(.dina(w_n8550_0[0]),.dinb(n8794),.dout(n8795),.clk(gclk));
	jand g08561(.dina(n8795),.dinb(n8728),.dout(n8796),.clk(gclk));
	jand g08562(.dina(n8796),.dinb(w_n3089_43[1]),.dout(n8797),.clk(gclk));
	jnot g08563(.din(w_n8558_0[0]),.dout(n8798),.clk(gclk));
	jor g08564(.dina(w_n8798_0[1]),.dinb(n8797),.dout(n8799),.clk(gclk));
	jand g08565(.dina(n8799),.dinb(n8727),.dout(n8800),.clk(gclk));
	jand g08566(.dina(n8800),.dinb(w_n2833_41[0]),.dout(n8801),.clk(gclk));
	jor g08567(.dina(w_n8565_0[0]),.dinb(n8801),.dout(n8802),.clk(gclk));
	jand g08568(.dina(n8802),.dinb(n8726),.dout(n8803),.clk(gclk));
	jand g08569(.dina(n8803),.dinb(w_n2572_43[2]),.dout(n8804),.clk(gclk));
	jnot g08570(.din(w_n8573_0[0]),.dout(n8805),.clk(gclk));
	jor g08571(.dina(w_n8805_0[1]),.dinb(n8804),.dout(n8806),.clk(gclk));
	jand g08572(.dina(n8806),.dinb(n8725),.dout(n8807),.clk(gclk));
	jand g08573(.dina(n8807),.dinb(w_n2345_41[2]),.dout(n8808),.clk(gclk));
	jor g08574(.dina(w_n8580_0[0]),.dinb(n8808),.dout(n8809),.clk(gclk));
	jand g08575(.dina(n8809),.dinb(n8724),.dout(n8810),.clk(gclk));
	jand g08576(.dina(n8810),.dinb(w_n2108_44[1]),.dout(n8811),.clk(gclk));
	jnot g08577(.din(w_n8588_0[0]),.dout(n8812),.clk(gclk));
	jor g08578(.dina(w_n8812_0[1]),.dinb(n8811),.dout(n8813),.clk(gclk));
	jand g08579(.dina(n8813),.dinb(n8723),.dout(n8814),.clk(gclk));
	jand g08580(.dina(n8814),.dinb(w_n1912_42[2]),.dout(n8815),.clk(gclk));
	jor g08581(.dina(w_n8595_0[0]),.dinb(n8815),.dout(n8816),.clk(gclk));
	jand g08582(.dina(n8816),.dinb(n8722),.dout(n8817),.clk(gclk));
	jand g08583(.dina(n8817),.dinb(w_n1699_45[0]),.dout(n8818),.clk(gclk));
	jnot g08584(.din(w_n8603_0[0]),.dout(n8819),.clk(gclk));
	jor g08585(.dina(w_n8819_0[1]),.dinb(n8818),.dout(n8820),.clk(gclk));
	jand g08586(.dina(n8820),.dinb(n8721),.dout(n8821),.clk(gclk));
	jand g08587(.dina(n8821),.dinb(w_n1516_43[1]),.dout(n8822),.clk(gclk));
	jnot g08588(.din(w_n8610_0[0]),.dout(n8823),.clk(gclk));
	jor g08589(.dina(w_n8823_0[1]),.dinb(n8822),.dout(n8824),.clk(gclk));
	jand g08590(.dina(n8824),.dinb(n8720),.dout(n8825),.clk(gclk));
	jand g08591(.dina(n8825),.dinb(w_n1332_45[0]),.dout(n8826),.clk(gclk));
	jnot g08592(.din(w_n8617_0[0]),.dout(n8827),.clk(gclk));
	jor g08593(.dina(w_n8827_0[1]),.dinb(n8826),.dout(n8828),.clk(gclk));
	jand g08594(.dina(n8828),.dinb(n8719),.dout(n8829),.clk(gclk));
	jand g08595(.dina(n8829),.dinb(w_n1173_44[0]),.dout(n8830),.clk(gclk));
	jor g08596(.dina(w_n8624_0[0]),.dinb(n8830),.dout(n8831),.clk(gclk));
	jand g08597(.dina(n8831),.dinb(n8718),.dout(n8832),.clk(gclk));
	jand g08598(.dina(n8832),.dinb(w_n1008_46[0]),.dout(n8833),.clk(gclk));
	jor g08599(.dina(w_n8632_0[0]),.dinb(n8833),.dout(n8834),.clk(gclk));
	jand g08600(.dina(n8834),.dinb(n8717),.dout(n8835),.clk(gclk));
	jand g08601(.dina(n8835),.dinb(w_n884_45[0]),.dout(n8836),.clk(gclk));
	jor g08602(.dina(w_n8640_0[0]),.dinb(n8836),.dout(n8837),.clk(gclk));
	jand g08603(.dina(n8837),.dinb(n8716),.dout(n8838),.clk(gclk));
	jand g08604(.dina(n8838),.dinb(w_n743_46[0]),.dout(n8839),.clk(gclk));
	jnot g08605(.din(w_n8648_0[0]),.dout(n8840),.clk(gclk));
	jor g08606(.dina(w_n8840_0[1]),.dinb(n8839),.dout(n8841),.clk(gclk));
	jand g08607(.dina(n8841),.dinb(n8715),.dout(n8842),.clk(gclk));
	jand g08608(.dina(n8842),.dinb(w_n635_46[0]),.dout(n8843),.clk(gclk));
	jor g08609(.dina(w_n8655_0[0]),.dinb(n8843),.dout(n8844),.clk(gclk));
	jand g08610(.dina(n8844),.dinb(n8714),.dout(n8845),.clk(gclk));
	jand g08611(.dina(n8845),.dinb(w_n515_47[0]),.dout(n8846),.clk(gclk));
	jnot g08612(.din(w_n8663_0[0]),.dout(n8847),.clk(gclk));
	jor g08613(.dina(w_n8847_0[1]),.dinb(n8846),.dout(n8848),.clk(gclk));
	jand g08614(.dina(n8848),.dinb(n8713),.dout(n8849),.clk(gclk));
	jand g08615(.dina(n8849),.dinb(w_n443_47[0]),.dout(n8850),.clk(gclk));
	jor g08616(.dina(w_n8670_0[0]),.dinb(n8850),.dout(n8851),.clk(gclk));
	jand g08617(.dina(n8851),.dinb(n8712),.dout(n8852),.clk(gclk));
	jand g08618(.dina(n8852),.dinb(w_n352_47[1]),.dout(n8853),.clk(gclk));
	jnot g08619(.din(w_n8678_0[0]),.dout(n8854),.clk(gclk));
	jor g08620(.dina(w_n8854_0[1]),.dinb(n8853),.dout(n8855),.clk(gclk));
	jand g08621(.dina(n8855),.dinb(n8711),.dout(n8856),.clk(gclk));
	jand g08622(.dina(n8856),.dinb(w_n294_47[2]),.dout(n8857),.clk(gclk));
	jnot g08623(.din(w_n8685_0[0]),.dout(n8858),.clk(gclk));
	jor g08624(.dina(w_n8858_0[1]),.dinb(n8857),.dout(n8859),.clk(gclk));
	jand g08625(.dina(n8859),.dinb(n8710),.dout(n8860),.clk(gclk));
	jand g08626(.dina(n8860),.dinb(w_n239_47[2]),.dout(n8861),.clk(gclk));
	jor g08627(.dina(w_n8692_0[0]),.dinb(n8861),.dout(n8862),.clk(gclk));
	jand g08628(.dina(n8862),.dinb(n8709),.dout(n8863),.clk(gclk));
	jand g08629(.dina(n8863),.dinb(w_n221_48[0]),.dout(n8864),.clk(gclk));
	jor g08630(.dina(w_n8700_0[1]),.dinb(n8864),.dout(n8865),.clk(gclk));
	jand g08631(.dina(n8865),.dinb(n8708),.dout(n8866),.clk(gclk));
	jor g08632(.dina(w_n8866_0[1]),.dinb(w_n8707_0[1]),.dout(n8867),.clk(gclk));
	jand g08633(.dina(w_asqrt28_25[1]),.dinb(w_n8444_0[0]),.dout(n8868),.clk(gclk));
	jor g08634(.dina(w_n8868_0[1]),.dinb(w_n8867_0[1]),.dout(n8869),.clk(gclk));
	jor g08635(.dina(n8869),.dinb(w_n8265_0[2]),.dout(n8870),.clk(gclk));
	jand g08636(.dina(n8870),.dinb(w_n218_20[0]),.dout(n8871),.clk(gclk));
	jand g08637(.dina(w_n8449_34[1]),.dinb(w_n8256_0[0]),.dout(n8872),.clk(gclk));
	jnot g08638(.din(n8872),.dout(n8873),.clk(gclk));
	jnot g08639(.din(w_n8265_0[1]),.dout(n8874),.clk(gclk));
	jand g08640(.dina(w_n8260_0[0]),.dinb(w_asqrt63_36[0]),.dout(n8875),.clk(gclk));
	jand g08641(.dina(n8875),.dinb(w_n8874_0[1]),.dout(n8876),.clk(gclk));
	jand g08642(.dina(w_n8876_0[1]),.dinb(n8873),.dout(n8877),.clk(gclk));
	jor g08643(.dina(w_n8877_0[1]),.dinb(w_n8871_0[1]),.dout(n8878),.clk(gclk));
	jor g08644(.dina(w_n8878_0[1]),.dinb(w_n8705_0[2]),.dout(asqrt_fa_28),.clk(gclk));
	jand g08645(.dina(w_n8703_0[0]),.dinb(w_n8277_0[0]),.dout(n8882),.clk(gclk));
	jnot g08646(.din(w_n8868_0[0]),.dout(n8883),.clk(gclk));
	jand g08647(.dina(n8883),.dinb(w_n8882_0[1]),.dout(n8884),.clk(gclk));
	jand g08648(.dina(n8884),.dinb(w_n8874_0[0]),.dout(n8885),.clk(gclk));
	jor g08649(.dina(n8885),.dinb(w_asqrt63_35[2]),.dout(n8886),.clk(gclk));
	jnot g08650(.din(w_n8877_0[0]),.dout(n8887),.clk(gclk));
	jand g08651(.dina(n8887),.dinb(n8886),.dout(n8888),.clk(gclk));
	jand g08652(.dina(w_n8888_0[1]),.dinb(w_n8704_0[1]),.dout(n8890),.clk(gclk));
	jxor g08653(.dina(w_n8695_0[0]),.dinb(w_n221_47[2]),.dout(n8891),.clk(gclk));
	jor g08654(.dina(n8891),.dinb(w_n8890_50[1]),.dout(n8892),.clk(gclk));
	jxor g08655(.dina(n8892),.dinb(w_n8700_0[0]),.dout(n8893),.clk(gclk));
	jnot g08656(.din(w_n8893_0[1]),.dout(n8894),.clk(gclk));
	jnot g08657(.din(w_a52_0[2]),.dout(n8895),.clk(gclk));
	jnot g08658(.din(w_a53_0[1]),.dout(n8896),.clk(gclk));
	jand g08659(.dina(w_n8896_0[1]),.dinb(w_n8895_1[2]),.dout(n8897),.clk(gclk));
	jand g08660(.dina(w_n8897_0[2]),.dinb(w_n8279_1[0]),.dout(n8898),.clk(gclk));
	jnot g08661(.din(w_n8898_0[1]),.dout(n8899),.clk(gclk));
	jor g08662(.dina(w_n8890_50[0]),.dinb(w_n8279_0[2]),.dout(n8900),.clk(gclk));
	jand g08663(.dina(n8900),.dinb(n8899),.dout(n8901),.clk(gclk));
	jor g08664(.dina(w_n8901_0[2]),.dinb(w_n8449_34[0]),.dout(n8902),.clk(gclk));
	jand g08665(.dina(w_n8901_0[1]),.dinb(w_n8449_33[2]),.dout(n8903),.clk(gclk));
	jor g08666(.dina(w_n8890_49[2]),.dinb(w_a54_1[0]),.dout(n8904),.clk(gclk));
	jand g08667(.dina(n8904),.dinb(w_a55_0[0]),.dout(n8905),.clk(gclk));
	jand g08668(.dina(w_asqrt27_20[1]),.dinb(w_n8281_0[1]),.dout(n8906),.clk(gclk));
	jor g08669(.dina(n8906),.dinb(n8905),.dout(n8907),.clk(gclk));
	jor g08670(.dina(n8907),.dinb(n8903),.dout(n8908),.clk(gclk));
	jand g08671(.dina(n8908),.dinb(w_n8902_0[1]),.dout(n8909),.clk(gclk));
	jor g08672(.dina(w_n8909_0[2]),.dinb(w_n8003_39[2]),.dout(n8910),.clk(gclk));
	jand g08673(.dina(w_n8909_0[1]),.dinb(w_n8003_39[1]),.dout(n8911),.clk(gclk));
	jnot g08674(.din(w_n8281_0[0]),.dout(n8912),.clk(gclk));
	jor g08675(.dina(w_n8890_49[1]),.dinb(n8912),.dout(n8913),.clk(gclk));
	jor g08676(.dina(w_n8705_0[1]),.dinb(w_n8449_33[1]),.dout(n8914),.clk(gclk));
	jor g08677(.dina(n8914),.dinb(w_n8876_0[0]),.dout(n8915),.clk(gclk));
	jor g08678(.dina(n8915),.dinb(w_n8871_0[0]),.dout(n8916),.clk(gclk));
	jand g08679(.dina(n8916),.dinb(w_n8913_0[1]),.dout(n8917),.clk(gclk));
	jxor g08680(.dina(n8917),.dinb(w_n7991_0[1]),.dout(n8918),.clk(gclk));
	jor g08681(.dina(w_n8918_0[2]),.dinb(n8911),.dout(n8919),.clk(gclk));
	jand g08682(.dina(n8919),.dinb(w_n8910_0[1]),.dout(n8920),.clk(gclk));
	jor g08683(.dina(w_n8920_0[2]),.dinb(w_n7581_35[0]),.dout(n8921),.clk(gclk));
	jand g08684(.dina(w_n8920_0[1]),.dinb(w_n7581_34[2]),.dout(n8922),.clk(gclk));
	jxor g08685(.dina(w_n8283_0[0]),.dinb(w_n8003_39[0]),.dout(n8923),.clk(gclk));
	jor g08686(.dina(n8923),.dinb(w_n8890_49[0]),.dout(n8924),.clk(gclk));
	jxor g08687(.dina(n8924),.dinb(w_n8750_0[0]),.dout(n8925),.clk(gclk));
	jnot g08688(.din(w_n8925_0[2]),.dout(n8926),.clk(gclk));
	jor g08689(.dina(n8926),.dinb(n8922),.dout(n8927),.clk(gclk));
	jand g08690(.dina(n8927),.dinb(w_n8921_0[1]),.dout(n8928),.clk(gclk));
	jor g08691(.dina(w_n8928_0[2]),.dinb(w_n7154_40[0]),.dout(n8929),.clk(gclk));
	jand g08692(.dina(w_n8928_0[1]),.dinb(w_n7154_39[2]),.dout(n8930),.clk(gclk));
	jxor g08693(.dina(w_n8453_0[0]),.dinb(w_n7581_34[1]),.dout(n8931),.clk(gclk));
	jor g08694(.dina(n8931),.dinb(w_n8890_48[2]),.dout(n8932),.clk(gclk));
	jxor g08695(.dina(n8932),.dinb(w_n8461_0[0]),.dout(n8933),.clk(gclk));
	jor g08696(.dina(w_n8933_0[2]),.dinb(n8930),.dout(n8934),.clk(gclk));
	jand g08697(.dina(n8934),.dinb(w_n8929_0[1]),.dout(n8935),.clk(gclk));
	jor g08698(.dina(w_n8935_0[2]),.dinb(w_n6758_35[2]),.dout(n8936),.clk(gclk));
	jand g08699(.dina(w_n8935_0[1]),.dinb(w_n6758_35[1]),.dout(n8937),.clk(gclk));
	jxor g08700(.dina(w_n8463_0[0]),.dinb(w_n7154_39[1]),.dout(n8938),.clk(gclk));
	jor g08701(.dina(n8938),.dinb(w_n8890_48[1]),.dout(n8939),.clk(gclk));
	jxor g08702(.dina(n8939),.dinb(w_n8468_0[0]),.dout(n8940),.clk(gclk));
	jor g08703(.dina(w_n8940_0[2]),.dinb(n8937),.dout(n8941),.clk(gclk));
	jand g08704(.dina(n8941),.dinb(w_n8936_0[1]),.dout(n8942),.clk(gclk));
	jor g08705(.dina(w_n8942_0[2]),.dinb(w_n6357_40[1]),.dout(n8943),.clk(gclk));
	jand g08706(.dina(w_n8942_0[1]),.dinb(w_n6357_40[0]),.dout(n8944),.clk(gclk));
	jxor g08707(.dina(w_n8470_0[0]),.dinb(w_n6758_35[0]),.dout(n8945),.clk(gclk));
	jor g08708(.dina(n8945),.dinb(w_n8890_48[0]),.dout(n8946),.clk(gclk));
	jxor g08709(.dina(n8946),.dinb(w_n8476_0[0]),.dout(n8947),.clk(gclk));
	jor g08710(.dina(w_n8947_0[2]),.dinb(n8944),.dout(n8948),.clk(gclk));
	jand g08711(.dina(n8948),.dinb(w_n8943_0[1]),.dout(n8949),.clk(gclk));
	jor g08712(.dina(w_n8949_0[2]),.dinb(w_n5989_36[1]),.dout(n8950),.clk(gclk));
	jand g08713(.dina(w_n8949_0[1]),.dinb(w_n5989_36[0]),.dout(n8951),.clk(gclk));
	jxor g08714(.dina(w_n8478_0[0]),.dinb(w_n6357_39[2]),.dout(n8952),.clk(gclk));
	jor g08715(.dina(n8952),.dinb(w_n8890_47[2]),.dout(n8953),.clk(gclk));
	jxor g08716(.dina(n8953),.dinb(w_n8484_0[0]),.dout(n8954),.clk(gclk));
	jor g08717(.dina(w_n8954_0[2]),.dinb(n8951),.dout(n8955),.clk(gclk));
	jand g08718(.dina(n8955),.dinb(w_n8950_0[1]),.dout(n8956),.clk(gclk));
	jor g08719(.dina(w_n8956_0[2]),.dinb(w_n5606_40[2]),.dout(n8957),.clk(gclk));
	jand g08720(.dina(w_n8956_0[1]),.dinb(w_n5606_40[1]),.dout(n8958),.clk(gclk));
	jxor g08721(.dina(w_n8486_0[0]),.dinb(w_n5989_35[2]),.dout(n8959),.clk(gclk));
	jor g08722(.dina(n8959),.dinb(w_n8890_47[1]),.dout(n8960),.clk(gclk));
	jxor g08723(.dina(n8960),.dinb(w_n8492_0[0]),.dout(n8961),.clk(gclk));
	jor g08724(.dina(w_n8961_0[2]),.dinb(n8958),.dout(n8962),.clk(gclk));
	jand g08725(.dina(n8962),.dinb(w_n8957_0[1]),.dout(n8963),.clk(gclk));
	jor g08726(.dina(w_n8963_0[2]),.dinb(w_n5259_37[1]),.dout(n8964),.clk(gclk));
	jxor g08727(.dina(w_n8494_0[0]),.dinb(w_n5606_40[0]),.dout(n8965),.clk(gclk));
	jor g08728(.dina(n8965),.dinb(w_n8890_47[0]),.dout(n8966),.clk(gclk));
	jxor g08729(.dina(n8966),.dinb(w_n8736_0[0]),.dout(n8967),.clk(gclk));
	jnot g08730(.din(w_n8967_0[2]),.dout(n8968),.clk(gclk));
	jand g08731(.dina(w_n8963_0[1]),.dinb(w_n5259_37[0]),.dout(n8969),.clk(gclk));
	jor g08732(.dina(n8969),.dinb(n8968),.dout(n8970),.clk(gclk));
	jand g08733(.dina(n8970),.dinb(w_n8964_0[1]),.dout(n8971),.clk(gclk));
	jor g08734(.dina(w_n8971_0[2]),.dinb(w_n4902_41[1]),.dout(n8972),.clk(gclk));
	jand g08735(.dina(w_n8971_0[1]),.dinb(w_n4902_41[0]),.dout(n8973),.clk(gclk));
	jxor g08736(.dina(w_n8501_0[0]),.dinb(w_n5259_36[2]),.dout(n8974),.clk(gclk));
	jor g08737(.dina(n8974),.dinb(w_n8890_46[2]),.dout(n8975),.clk(gclk));
	jxor g08738(.dina(n8975),.dinb(w_n8507_0[0]),.dout(n8976),.clk(gclk));
	jor g08739(.dina(w_n8976_0[2]),.dinb(n8973),.dout(n8977),.clk(gclk));
	jand g08740(.dina(n8977),.dinb(w_n8972_0[1]),.dout(n8978),.clk(gclk));
	jor g08741(.dina(w_n8978_0[2]),.dinb(w_n4582_38[1]),.dout(n8979),.clk(gclk));
	jand g08742(.dina(w_n8978_0[1]),.dinb(w_n4582_38[0]),.dout(n8980),.clk(gclk));
	jxor g08743(.dina(w_n8509_0[0]),.dinb(w_n4902_40[2]),.dout(n8981),.clk(gclk));
	jor g08744(.dina(n8981),.dinb(w_n8890_46[1]),.dout(n8982),.clk(gclk));
	jxor g08745(.dina(n8982),.dinb(w_n8776_0[0]),.dout(n8983),.clk(gclk));
	jnot g08746(.din(w_n8983_0[2]),.dout(n8984),.clk(gclk));
	jor g08747(.dina(n8984),.dinb(n8980),.dout(n8985),.clk(gclk));
	jand g08748(.dina(n8985),.dinb(w_n8979_0[1]),.dout(n8986),.clk(gclk));
	jor g08749(.dina(w_n8986_0[2]),.dinb(w_n4249_42[0]),.dout(n8987),.clk(gclk));
	jand g08750(.dina(w_n8986_0[1]),.dinb(w_n4249_41[2]),.dout(n8988),.clk(gclk));
	jxor g08751(.dina(w_n8516_0[0]),.dinb(w_n4582_37[2]),.dout(n8989),.clk(gclk));
	jor g08752(.dina(n8989),.dinb(w_n8890_46[0]),.dout(n8990),.clk(gclk));
	jxor g08753(.dina(n8990),.dinb(w_n8522_0[0]),.dout(n8991),.clk(gclk));
	jor g08754(.dina(w_n8991_0[2]),.dinb(n8988),.dout(n8992),.clk(gclk));
	jand g08755(.dina(n8992),.dinb(w_n8987_0[1]),.dout(n8993),.clk(gclk));
	jor g08756(.dina(w_n8993_0[2]),.dinb(w_n3955_39[0]),.dout(n8994),.clk(gclk));
	jand g08757(.dina(w_n8993_0[1]),.dinb(w_n3955_38[2]),.dout(n8995),.clk(gclk));
	jxor g08758(.dina(w_n8524_0[0]),.dinb(w_n4249_41[1]),.dout(n8996),.clk(gclk));
	jor g08759(.dina(n8996),.dinb(w_n8890_45[2]),.dout(n8997),.clk(gclk));
	jxor g08760(.dina(n8997),.dinb(w_n8783_0[0]),.dout(n8998),.clk(gclk));
	jnot g08761(.din(w_n8998_0[2]),.dout(n8999),.clk(gclk));
	jor g08762(.dina(n8999),.dinb(n8995),.dout(n9000),.clk(gclk));
	jand g08763(.dina(n9000),.dinb(w_n8994_0[1]),.dout(n9001),.clk(gclk));
	jor g08764(.dina(w_n9001_0[2]),.dinb(w_n3642_42[1]),.dout(n9002),.clk(gclk));
	jand g08765(.dina(w_n9001_0[1]),.dinb(w_n3642_42[0]),.dout(n9003),.clk(gclk));
	jxor g08766(.dina(w_n8531_0[0]),.dinb(w_n3955_38[1]),.dout(n9004),.clk(gclk));
	jor g08767(.dina(n9004),.dinb(w_n8890_45[1]),.dout(n9005),.clk(gclk));
	jxor g08768(.dina(n9005),.dinb(w_n8787_0[0]),.dout(n9006),.clk(gclk));
	jnot g08769(.din(w_n9006_0[2]),.dout(n9007),.clk(gclk));
	jor g08770(.dina(n9007),.dinb(n9003),.dout(n9008),.clk(gclk));
	jand g08771(.dina(n9008),.dinb(w_n9002_0[1]),.dout(n9009),.clk(gclk));
	jor g08772(.dina(w_n9009_0[2]),.dinb(w_n3368_39[2]),.dout(n9010),.clk(gclk));
	jand g08773(.dina(w_n9009_0[1]),.dinb(w_n3368_39[1]),.dout(n9011),.clk(gclk));
	jxor g08774(.dina(w_n8538_0[0]),.dinb(w_n3642_41[2]),.dout(n9012),.clk(gclk));
	jor g08775(.dina(n9012),.dinb(w_n8890_45[0]),.dout(n9013),.clk(gclk));
	jxor g08776(.dina(n9013),.dinb(w_n8791_0[0]),.dout(n9014),.clk(gclk));
	jnot g08777(.din(w_n9014_0[1]),.dout(n9015),.clk(gclk));
	jor g08778(.dina(w_n9015_0[1]),.dinb(n9011),.dout(n9016),.clk(gclk));
	jand g08779(.dina(n9016),.dinb(w_n9010_0[1]),.dout(n9017),.clk(gclk));
	jor g08780(.dina(w_n9017_0[2]),.dinb(w_n3089_43[0]),.dout(n9018),.clk(gclk));
	jand g08781(.dina(w_n9017_0[1]),.dinb(w_n3089_42[2]),.dout(n9019),.clk(gclk));
	jxor g08782(.dina(w_n8545_0[0]),.dinb(w_n3368_39[0]),.dout(n9020),.clk(gclk));
	jor g08783(.dina(n9020),.dinb(w_n8890_44[2]),.dout(n9021),.clk(gclk));
	jxor g08784(.dina(n9021),.dinb(w_n8551_0[0]),.dout(n9022),.clk(gclk));
	jor g08785(.dina(w_n9022_0[2]),.dinb(n9019),.dout(n9023),.clk(gclk));
	jand g08786(.dina(n9023),.dinb(w_n9018_0[1]),.dout(n9024),.clk(gclk));
	jor g08787(.dina(w_n9024_0[2]),.dinb(w_n2833_40[2]),.dout(n9025),.clk(gclk));
	jand g08788(.dina(w_n9024_0[1]),.dinb(w_n2833_40[1]),.dout(n9026),.clk(gclk));
	jxor g08789(.dina(w_n8553_0[0]),.dinb(w_n3089_42[1]),.dout(n9027),.clk(gclk));
	jor g08790(.dina(n9027),.dinb(w_n8890_44[1]),.dout(n9028),.clk(gclk));
	jxor g08791(.dina(n9028),.dinb(w_n8798_0[0]),.dout(n9029),.clk(gclk));
	jnot g08792(.din(w_n9029_0[2]),.dout(n9030),.clk(gclk));
	jor g08793(.dina(n9030),.dinb(n9026),.dout(n9031),.clk(gclk));
	jand g08794(.dina(n9031),.dinb(w_n9025_0[1]),.dout(n9032),.clk(gclk));
	jor g08795(.dina(w_n9032_0[2]),.dinb(w_n2572_43[1]),.dout(n9033),.clk(gclk));
	jand g08796(.dina(w_n9032_0[1]),.dinb(w_n2572_43[0]),.dout(n9034),.clk(gclk));
	jxor g08797(.dina(w_n8560_0[0]),.dinb(w_n2833_40[0]),.dout(n9035),.clk(gclk));
	jor g08798(.dina(n9035),.dinb(w_n8890_44[0]),.dout(n9036),.clk(gclk));
	jxor g08799(.dina(n9036),.dinb(w_n8566_0[0]),.dout(n9037),.clk(gclk));
	jor g08800(.dina(w_n9037_0[2]),.dinb(n9034),.dout(n9038),.clk(gclk));
	jand g08801(.dina(n9038),.dinb(w_n9033_0[1]),.dout(n9039),.clk(gclk));
	jor g08802(.dina(w_n9039_0[2]),.dinb(w_n2345_41[1]),.dout(n9040),.clk(gclk));
	jand g08803(.dina(w_n9039_0[1]),.dinb(w_n2345_41[0]),.dout(n9041),.clk(gclk));
	jxor g08804(.dina(w_n8568_0[0]),.dinb(w_n2572_42[2]),.dout(n9042),.clk(gclk));
	jor g08805(.dina(n9042),.dinb(w_n8890_43[2]),.dout(n9043),.clk(gclk));
	jxor g08806(.dina(n9043),.dinb(w_n8805_0[0]),.dout(n9044),.clk(gclk));
	jnot g08807(.din(w_n9044_0[2]),.dout(n9045),.clk(gclk));
	jor g08808(.dina(n9045),.dinb(n9041),.dout(n9046),.clk(gclk));
	jand g08809(.dina(n9046),.dinb(w_n9040_0[1]),.dout(n9047),.clk(gclk));
	jor g08810(.dina(w_n9047_0[2]),.dinb(w_n2108_44[0]),.dout(n9048),.clk(gclk));
	jand g08811(.dina(w_n9047_0[1]),.dinb(w_n2108_43[2]),.dout(n9049),.clk(gclk));
	jxor g08812(.dina(w_n8575_0[0]),.dinb(w_n2345_40[2]),.dout(n9050),.clk(gclk));
	jor g08813(.dina(n9050),.dinb(w_n8890_43[1]),.dout(n9051),.clk(gclk));
	jxor g08814(.dina(n9051),.dinb(w_n8581_0[0]),.dout(n9052),.clk(gclk));
	jor g08815(.dina(w_n9052_0[2]),.dinb(n9049),.dout(n9053),.clk(gclk));
	jand g08816(.dina(n9053),.dinb(w_n9048_0[1]),.dout(n9054),.clk(gclk));
	jor g08817(.dina(w_n9054_0[2]),.dinb(w_n1912_42[1]),.dout(n9055),.clk(gclk));
	jand g08818(.dina(w_n9054_0[1]),.dinb(w_n1912_42[0]),.dout(n9056),.clk(gclk));
	jxor g08819(.dina(w_n8583_0[0]),.dinb(w_n2108_43[1]),.dout(n9057),.clk(gclk));
	jor g08820(.dina(n9057),.dinb(w_n8890_43[0]),.dout(n9058),.clk(gclk));
	jxor g08821(.dina(n9058),.dinb(w_n8812_0[0]),.dout(n9059),.clk(gclk));
	jnot g08822(.din(w_n9059_0[2]),.dout(n9060),.clk(gclk));
	jor g08823(.dina(n9060),.dinb(n9056),.dout(n9061),.clk(gclk));
	jand g08824(.dina(n9061),.dinb(w_n9055_0[1]),.dout(n9062),.clk(gclk));
	jor g08825(.dina(w_n9062_0[2]),.dinb(w_n1699_44[2]),.dout(n9063),.clk(gclk));
	jand g08826(.dina(w_n9062_0[1]),.dinb(w_n1699_44[1]),.dout(n9064),.clk(gclk));
	jxor g08827(.dina(w_n8590_0[0]),.dinb(w_n1912_41[2]),.dout(n9065),.clk(gclk));
	jor g08828(.dina(n9065),.dinb(w_n8890_42[2]),.dout(n9066),.clk(gclk));
	jxor g08829(.dina(n9066),.dinb(w_n8596_0[0]),.dout(n9067),.clk(gclk));
	jor g08830(.dina(w_n9067_0[2]),.dinb(n9064),.dout(n9068),.clk(gclk));
	jand g08831(.dina(n9068),.dinb(w_n9063_0[1]),.dout(n9069),.clk(gclk));
	jor g08832(.dina(w_n9069_0[2]),.dinb(w_n1516_43[0]),.dout(n9070),.clk(gclk));
	jand g08833(.dina(w_n9069_0[1]),.dinb(w_n1516_42[2]),.dout(n9071),.clk(gclk));
	jxor g08834(.dina(w_n8598_0[0]),.dinb(w_n1699_44[0]),.dout(n9072),.clk(gclk));
	jor g08835(.dina(n9072),.dinb(w_n8890_42[1]),.dout(n9073),.clk(gclk));
	jxor g08836(.dina(n9073),.dinb(w_n8819_0[0]),.dout(n9074),.clk(gclk));
	jnot g08837(.din(w_n9074_0[2]),.dout(n9075),.clk(gclk));
	jor g08838(.dina(n9075),.dinb(n9071),.dout(n9076),.clk(gclk));
	jand g08839(.dina(n9076),.dinb(w_n9070_0[1]),.dout(n9077),.clk(gclk));
	jor g08840(.dina(w_n9077_0[2]),.dinb(w_n1332_44[2]),.dout(n9078),.clk(gclk));
	jand g08841(.dina(w_n9077_0[1]),.dinb(w_n1332_44[1]),.dout(n9079),.clk(gclk));
	jxor g08842(.dina(w_n8605_0[0]),.dinb(w_n1516_42[1]),.dout(n9080),.clk(gclk));
	jor g08843(.dina(n9080),.dinb(w_n8890_42[0]),.dout(n9081),.clk(gclk));
	jxor g08844(.dina(n9081),.dinb(w_n8823_0[0]),.dout(n9082),.clk(gclk));
	jnot g08845(.din(w_n9082_0[2]),.dout(n9083),.clk(gclk));
	jor g08846(.dina(n9083),.dinb(n9079),.dout(n9084),.clk(gclk));
	jand g08847(.dina(n9084),.dinb(w_n9078_0[1]),.dout(n9085),.clk(gclk));
	jor g08848(.dina(w_n9085_0[2]),.dinb(w_n1173_43[2]),.dout(n9086),.clk(gclk));
	jand g08849(.dina(w_n9085_0[1]),.dinb(w_n1173_43[1]),.dout(n9087),.clk(gclk));
	jxor g08850(.dina(w_n8612_0[0]),.dinb(w_n1332_44[0]),.dout(n9088),.clk(gclk));
	jor g08851(.dina(n9088),.dinb(w_n8890_41[2]),.dout(n9089),.clk(gclk));
	jxor g08852(.dina(n9089),.dinb(w_n8827_0[0]),.dout(n9090),.clk(gclk));
	jnot g08853(.din(w_n9090_0[2]),.dout(n9091),.clk(gclk));
	jor g08854(.dina(n9091),.dinb(n9087),.dout(n9092),.clk(gclk));
	jand g08855(.dina(n9092),.dinb(w_n9086_0[1]),.dout(n9093),.clk(gclk));
	jor g08856(.dina(w_n9093_0[2]),.dinb(w_n1008_45[2]),.dout(n9094),.clk(gclk));
	jand g08857(.dina(w_n9093_0[1]),.dinb(w_n1008_45[1]),.dout(n9095),.clk(gclk));
	jxor g08858(.dina(w_n8619_0[0]),.dinb(w_n1173_43[0]),.dout(n9096),.clk(gclk));
	jor g08859(.dina(n9096),.dinb(w_n8890_41[1]),.dout(n9097),.clk(gclk));
	jxor g08860(.dina(n9097),.dinb(w_n8625_0[0]),.dout(n9098),.clk(gclk));
	jor g08861(.dina(w_n9098_0[2]),.dinb(n9095),.dout(n9099),.clk(gclk));
	jand g08862(.dina(n9099),.dinb(w_n9094_0[1]),.dout(n9100),.clk(gclk));
	jor g08863(.dina(w_n9100_0[2]),.dinb(w_n884_44[2]),.dout(n9101),.clk(gclk));
	jand g08864(.dina(w_n9100_0[1]),.dinb(w_n884_44[1]),.dout(n9102),.clk(gclk));
	jxor g08865(.dina(w_n8627_0[0]),.dinb(w_n1008_45[0]),.dout(n9103),.clk(gclk));
	jor g08866(.dina(n9103),.dinb(w_n8890_41[0]),.dout(n9104),.clk(gclk));
	jxor g08867(.dina(n9104),.dinb(w_n8633_0[0]),.dout(n9105),.clk(gclk));
	jor g08868(.dina(w_n9105_0[2]),.dinb(n9102),.dout(n9106),.clk(gclk));
	jand g08869(.dina(n9106),.dinb(w_n9101_0[1]),.dout(n9107),.clk(gclk));
	jor g08870(.dina(w_n9107_0[2]),.dinb(w_n743_45[2]),.dout(n9108),.clk(gclk));
	jand g08871(.dina(w_n9107_0[1]),.dinb(w_n743_45[1]),.dout(n9109),.clk(gclk));
	jxor g08872(.dina(w_n8635_0[0]),.dinb(w_n884_44[0]),.dout(n9110),.clk(gclk));
	jor g08873(.dina(n9110),.dinb(w_n8890_40[2]),.dout(n9111),.clk(gclk));
	jxor g08874(.dina(n9111),.dinb(w_n8641_0[0]),.dout(n9112),.clk(gclk));
	jor g08875(.dina(w_n9112_0[2]),.dinb(n9109),.dout(n9113),.clk(gclk));
	jand g08876(.dina(n9113),.dinb(w_n9108_0[1]),.dout(n9114),.clk(gclk));
	jor g08877(.dina(w_n9114_0[2]),.dinb(w_n635_45[2]),.dout(n9115),.clk(gclk));
	jand g08878(.dina(w_n9114_0[1]),.dinb(w_n635_45[1]),.dout(n9116),.clk(gclk));
	jxor g08879(.dina(w_n8643_0[0]),.dinb(w_n743_45[0]),.dout(n9117),.clk(gclk));
	jor g08880(.dina(n9117),.dinb(w_n8890_40[1]),.dout(n9118),.clk(gclk));
	jxor g08881(.dina(n9118),.dinb(w_n8840_0[0]),.dout(n9119),.clk(gclk));
	jnot g08882(.din(w_n9119_0[2]),.dout(n9120),.clk(gclk));
	jor g08883(.dina(n9120),.dinb(n9116),.dout(n9121),.clk(gclk));
	jand g08884(.dina(n9121),.dinb(w_n9115_0[1]),.dout(n9122),.clk(gclk));
	jor g08885(.dina(w_n9122_0[2]),.dinb(w_n515_46[2]),.dout(n9123),.clk(gclk));
	jand g08886(.dina(w_n9122_0[1]),.dinb(w_n515_46[1]),.dout(n9124),.clk(gclk));
	jxor g08887(.dina(w_n8650_0[0]),.dinb(w_n635_45[0]),.dout(n9125),.clk(gclk));
	jor g08888(.dina(n9125),.dinb(w_n8890_40[0]),.dout(n9126),.clk(gclk));
	jxor g08889(.dina(n9126),.dinb(w_n8656_0[0]),.dout(n9127),.clk(gclk));
	jor g08890(.dina(w_n9127_0[2]),.dinb(n9124),.dout(n9128),.clk(gclk));
	jand g08891(.dina(n9128),.dinb(w_n9123_0[1]),.dout(n9129),.clk(gclk));
	jor g08892(.dina(w_n9129_0[2]),.dinb(w_n443_46[2]),.dout(n9130),.clk(gclk));
	jand g08893(.dina(w_n9129_0[1]),.dinb(w_n443_46[1]),.dout(n9131),.clk(gclk));
	jxor g08894(.dina(w_n8658_0[0]),.dinb(w_n515_46[0]),.dout(n9132),.clk(gclk));
	jor g08895(.dina(n9132),.dinb(w_n8890_39[2]),.dout(n9133),.clk(gclk));
	jxor g08896(.dina(n9133),.dinb(w_n8847_0[0]),.dout(n9134),.clk(gclk));
	jnot g08897(.din(w_n9134_0[1]),.dout(n9135),.clk(gclk));
	jor g08898(.dina(w_n9135_0[1]),.dinb(n9131),.dout(n9136),.clk(gclk));
	jand g08899(.dina(n9136),.dinb(w_n9130_0[1]),.dout(n9137),.clk(gclk));
	jor g08900(.dina(w_n9137_0[2]),.dinb(w_n352_47[0]),.dout(n9138),.clk(gclk));
	jand g08901(.dina(w_n9137_0[1]),.dinb(w_n352_46[2]),.dout(n9139),.clk(gclk));
	jxor g08902(.dina(w_n8665_0[0]),.dinb(w_n443_46[0]),.dout(n9140),.clk(gclk));
	jor g08903(.dina(n9140),.dinb(w_n8890_39[1]),.dout(n9141),.clk(gclk));
	jxor g08904(.dina(n9141),.dinb(w_n8671_0[0]),.dout(n9142),.clk(gclk));
	jor g08905(.dina(w_n9142_0[2]),.dinb(n9139),.dout(n9143),.clk(gclk));
	jand g08906(.dina(n9143),.dinb(w_n9138_0[1]),.dout(n9144),.clk(gclk));
	jor g08907(.dina(w_n9144_0[2]),.dinb(w_n294_47[1]),.dout(n9145),.clk(gclk));
	jand g08908(.dina(w_n9144_0[1]),.dinb(w_n294_47[0]),.dout(n9146),.clk(gclk));
	jxor g08909(.dina(w_n8673_0[0]),.dinb(w_n352_46[1]),.dout(n9147),.clk(gclk));
	jor g08910(.dina(n9147),.dinb(w_n8890_39[0]),.dout(n9148),.clk(gclk));
	jxor g08911(.dina(n9148),.dinb(w_n8854_0[0]),.dout(n9149),.clk(gclk));
	jnot g08912(.din(w_n9149_0[2]),.dout(n9150),.clk(gclk));
	jor g08913(.dina(n9150),.dinb(n9146),.dout(n9151),.clk(gclk));
	jand g08914(.dina(n9151),.dinb(w_n9145_0[1]),.dout(n9152),.clk(gclk));
	jor g08915(.dina(w_n9152_0[2]),.dinb(w_n239_47[1]),.dout(n9153),.clk(gclk));
	jand g08916(.dina(w_n9152_0[1]),.dinb(w_n239_47[0]),.dout(n9154),.clk(gclk));
	jxor g08917(.dina(w_n8680_0[0]),.dinb(w_n294_46[2]),.dout(n9155),.clk(gclk));
	jor g08918(.dina(n9155),.dinb(w_n8890_38[2]),.dout(n9156),.clk(gclk));
	jxor g08919(.dina(n9156),.dinb(w_n8858_0[0]),.dout(n9157),.clk(gclk));
	jnot g08920(.din(w_n9157_0[2]),.dout(n9158),.clk(gclk));
	jor g08921(.dina(n9158),.dinb(n9154),.dout(n9159),.clk(gclk));
	jand g08922(.dina(n9159),.dinb(w_n9153_0[1]),.dout(n9160),.clk(gclk));
	jor g08923(.dina(w_n9160_0[2]),.dinb(w_n221_47[1]),.dout(n9161),.clk(gclk));
	jand g08924(.dina(w_n9160_0[1]),.dinb(w_n221_47[0]),.dout(n9162),.clk(gclk));
	jxor g08925(.dina(w_n8687_0[0]),.dinb(w_n239_46[2]),.dout(n9163),.clk(gclk));
	jor g08926(.dina(n9163),.dinb(w_n8890_38[1]),.dout(n9164),.clk(gclk));
	jxor g08927(.dina(n9164),.dinb(w_n8693_0[0]),.dout(n9165),.clk(gclk));
	jor g08928(.dina(w_n9165_0[1]),.dinb(n9162),.dout(n9166),.clk(gclk));
	jand g08929(.dina(n9166),.dinb(w_n9161_0[1]),.dout(n9167),.clk(gclk));
	jand g08930(.dina(w_n9167_1[1]),.dinb(w_n8894_1[1]),.dout(n9168),.clk(gclk));
	jand g08931(.dina(w_n8888_0[0]),.dinb(w_n8866_0[0]),.dout(n9169),.clk(gclk));
	jand g08932(.dina(w_n8867_0[0]),.dinb(w_asqrt63_35[1]),.dout(n9170),.clk(gclk));
	jand g08933(.dina(n9170),.dinb(w_n8704_0[0]),.dout(n9171),.clk(gclk));
	jnot g08934(.din(n9171),.dout(n9172),.clk(gclk));
	jor g08935(.dina(w_n9172_0[1]),.dinb(n9169),.dout(n9173),.clk(gclk));
	jnot g08936(.din(w_n9173_0[1]),.dout(n9174),.clk(gclk));
	jor g08937(.dina(w_n9167_1[0]),.dinb(w_n8894_1[0]),.dout(n9175),.clk(gclk));
	jand g08938(.dina(w_n8878_0[0]),.dinb(w_n8882_0[0]),.dout(n9176),.clk(gclk));
	jor g08939(.dina(n9176),.dinb(w_n8705_0[0]),.dout(n9177),.clk(gclk));
	jor g08940(.dina(w_n9177_0[1]),.dinb(n9175),.dout(n9178),.clk(gclk));
	jand g08941(.dina(n9178),.dinb(w_n218_19[2]),.dout(n9179),.clk(gclk));
	jand g08942(.dina(w_n8890_38[0]),.dinb(w_n8707_0[0]),.dout(n9180),.clk(gclk));
	jor g08943(.dina(w_n9180_0[1]),.dinb(n9179),.dout(n9181),.clk(gclk));
	jor g08944(.dina(n9181),.dinb(n9174),.dout(n9182),.clk(gclk));
	jor g08945(.dina(n9182),.dinb(w_n9168_0[1]),.dout(asqrt_fa_27),.clk(gclk));
	jnot g08946(.din(w_n9165_0[0]),.dout(n9184),.clk(gclk));
	jxor g08947(.dina(w_n9160_0[0]),.dinb(w_n221_46[2]),.dout(n9185),.clk(gclk));
	jand g08948(.dina(n9185),.dinb(w_asqrt26_36[1]),.dout(n9186),.clk(gclk));
	jxor g08949(.dina(n9186),.dinb(w_n9184_0[1]),.dout(n9187),.clk(gclk));
	jnot g08950(.din(w_a50_0[2]),.dout(n9188),.clk(gclk));
	jnot g08951(.din(w_a51_0[1]),.dout(n9189),.clk(gclk));
	jand g08952(.dina(w_n9189_0[1]),.dinb(w_n9188_1[2]),.dout(n9190),.clk(gclk));
	jand g08953(.dina(w_n9190_0[2]),.dinb(w_n8895_1[1]),.dout(n9191),.clk(gclk));
	jand g08954(.dina(w_asqrt26_36[0]),.dinb(w_a52_0[1]),.dout(n9192),.clk(gclk));
	jor g08955(.dina(n9192),.dinb(w_n9191_0[1]),.dout(n9193),.clk(gclk));
	jand g08956(.dina(w_n9193_0[2]),.dinb(w_asqrt27_20[0]),.dout(n9194),.clk(gclk));
	jor g08957(.dina(w_n9193_0[1]),.dinb(w_asqrt27_19[2]),.dout(n9195),.clk(gclk));
	jand g08958(.dina(w_asqrt26_35[2]),.dinb(w_n8895_1[0]),.dout(n9196),.clk(gclk));
	jor g08959(.dina(n9196),.dinb(w_n8896_0[0]),.dout(n9197),.clk(gclk));
	jnot g08960(.din(w_n8897_0[1]),.dout(n9198),.clk(gclk));
	jnot g08961(.din(w_n9168_0[0]),.dout(n9199),.clk(gclk));
	jnot g08962(.din(w_n9161_0[0]),.dout(n9200),.clk(gclk));
	jnot g08963(.din(w_n9153_0[0]),.dout(n9201),.clk(gclk));
	jnot g08964(.din(w_n9145_0[0]),.dout(n9202),.clk(gclk));
	jnot g08965(.din(w_n9138_0[0]),.dout(n9203),.clk(gclk));
	jnot g08966(.din(w_n9130_0[0]),.dout(n9204),.clk(gclk));
	jnot g08967(.din(w_n9123_0[0]),.dout(n9205),.clk(gclk));
	jnot g08968(.din(w_n9115_0[0]),.dout(n9206),.clk(gclk));
	jnot g08969(.din(w_n9108_0[0]),.dout(n9207),.clk(gclk));
	jnot g08970(.din(w_n9101_0[0]),.dout(n9208),.clk(gclk));
	jnot g08971(.din(w_n9094_0[0]),.dout(n9209),.clk(gclk));
	jnot g08972(.din(w_n9086_0[0]),.dout(n9210),.clk(gclk));
	jnot g08973(.din(w_n9078_0[0]),.dout(n9211),.clk(gclk));
	jnot g08974(.din(w_n9070_0[0]),.dout(n9212),.clk(gclk));
	jnot g08975(.din(w_n9063_0[0]),.dout(n9213),.clk(gclk));
	jnot g08976(.din(w_n9055_0[0]),.dout(n9214),.clk(gclk));
	jnot g08977(.din(w_n9048_0[0]),.dout(n9215),.clk(gclk));
	jnot g08978(.din(w_n9040_0[0]),.dout(n9216),.clk(gclk));
	jnot g08979(.din(w_n9033_0[0]),.dout(n9217),.clk(gclk));
	jnot g08980(.din(w_n9025_0[0]),.dout(n9218),.clk(gclk));
	jnot g08981(.din(w_n9018_0[0]),.dout(n9219),.clk(gclk));
	jnot g08982(.din(w_n9010_0[0]),.dout(n9220),.clk(gclk));
	jnot g08983(.din(w_n9002_0[0]),.dout(n9221),.clk(gclk));
	jnot g08984(.din(w_n8994_0[0]),.dout(n9222),.clk(gclk));
	jnot g08985(.din(w_n8987_0[0]),.dout(n9223),.clk(gclk));
	jnot g08986(.din(w_n8979_0[0]),.dout(n9224),.clk(gclk));
	jnot g08987(.din(w_n8972_0[0]),.dout(n9225),.clk(gclk));
	jnot g08988(.din(w_n8964_0[0]),.dout(n9226),.clk(gclk));
	jnot g08989(.din(w_n8957_0[0]),.dout(n9227),.clk(gclk));
	jnot g08990(.din(w_n8950_0[0]),.dout(n9228),.clk(gclk));
	jnot g08991(.din(w_n8943_0[0]),.dout(n9229),.clk(gclk));
	jnot g08992(.din(w_n8936_0[0]),.dout(n9230),.clk(gclk));
	jnot g08993(.din(w_n8929_0[0]),.dout(n9231),.clk(gclk));
	jnot g08994(.din(w_n8921_0[0]),.dout(n9232),.clk(gclk));
	jnot g08995(.din(w_n8910_0[0]),.dout(n9233),.clk(gclk));
	jnot g08996(.din(w_n8902_0[0]),.dout(n9234),.clk(gclk));
	jand g08997(.dina(w_asqrt27_19[1]),.dinb(w_a54_0[2]),.dout(n9235),.clk(gclk));
	jor g08998(.dina(n9235),.dinb(w_n8898_0[0]),.dout(n9236),.clk(gclk));
	jor g08999(.dina(n9236),.dinb(w_asqrt28_25[0]),.dout(n9237),.clk(gclk));
	jand g09000(.dina(w_asqrt27_19[0]),.dinb(w_n8279_0[1]),.dout(n9238),.clk(gclk));
	jor g09001(.dina(n9238),.dinb(w_n8280_0[0]),.dout(n9239),.clk(gclk));
	jand g09002(.dina(w_n8913_0[0]),.dinb(n9239),.dout(n9240),.clk(gclk));
	jand g09003(.dina(w_n9240_0[1]),.dinb(n9237),.dout(n9241),.clk(gclk));
	jor g09004(.dina(n9241),.dinb(n9234),.dout(n9242),.clk(gclk));
	jor g09005(.dina(n9242),.dinb(w_asqrt29_19[2]),.dout(n9243),.clk(gclk));
	jnot g09006(.din(w_n8918_0[1]),.dout(n9244),.clk(gclk));
	jand g09007(.dina(n9244),.dinb(n9243),.dout(n9245),.clk(gclk));
	jor g09008(.dina(n9245),.dinb(n9233),.dout(n9246),.clk(gclk));
	jor g09009(.dina(n9246),.dinb(w_asqrt30_25[1]),.dout(n9247),.clk(gclk));
	jand g09010(.dina(w_n8925_0[1]),.dinb(n9247),.dout(n9248),.clk(gclk));
	jor g09011(.dina(n9248),.dinb(n9232),.dout(n9249),.clk(gclk));
	jor g09012(.dina(n9249),.dinb(w_asqrt31_20[1]),.dout(n9250),.clk(gclk));
	jnot g09013(.din(w_n8933_0[1]),.dout(n9251),.clk(gclk));
	jand g09014(.dina(n9251),.dinb(n9250),.dout(n9252),.clk(gclk));
	jor g09015(.dina(n9252),.dinb(n9231),.dout(n9253),.clk(gclk));
	jor g09016(.dina(n9253),.dinb(w_asqrt32_25[1]),.dout(n9254),.clk(gclk));
	jnot g09017(.din(w_n8940_0[1]),.dout(n9255),.clk(gclk));
	jand g09018(.dina(n9255),.dinb(n9254),.dout(n9256),.clk(gclk));
	jor g09019(.dina(n9256),.dinb(n9230),.dout(n9257),.clk(gclk));
	jor g09020(.dina(n9257),.dinb(w_asqrt33_21[0]),.dout(n9258),.clk(gclk));
	jnot g09021(.din(w_n8947_0[1]),.dout(n9259),.clk(gclk));
	jand g09022(.dina(n9259),.dinb(n9258),.dout(n9260),.clk(gclk));
	jor g09023(.dina(n9260),.dinb(n9229),.dout(n9261),.clk(gclk));
	jor g09024(.dina(n9261),.dinb(w_asqrt34_25[2]),.dout(n9262),.clk(gclk));
	jnot g09025(.din(w_n8954_0[1]),.dout(n9263),.clk(gclk));
	jand g09026(.dina(n9263),.dinb(n9262),.dout(n9264),.clk(gclk));
	jor g09027(.dina(n9264),.dinb(n9228),.dout(n9265),.clk(gclk));
	jor g09028(.dina(n9265),.dinb(w_asqrt35_21[2]),.dout(n9266),.clk(gclk));
	jnot g09029(.din(w_n8961_0[1]),.dout(n9267),.clk(gclk));
	jand g09030(.dina(n9267),.dinb(n9266),.dout(n9268),.clk(gclk));
	jor g09031(.dina(n9268),.dinb(n9227),.dout(n9269),.clk(gclk));
	jor g09032(.dina(n9269),.dinb(w_asqrt36_25[2]),.dout(n9270),.clk(gclk));
	jand g09033(.dina(n9270),.dinb(w_n8967_0[1]),.dout(n9271),.clk(gclk));
	jor g09034(.dina(n9271),.dinb(n9226),.dout(n9272),.clk(gclk));
	jor g09035(.dina(n9272),.dinb(w_asqrt37_22[0]),.dout(n9273),.clk(gclk));
	jnot g09036(.din(w_n8976_0[1]),.dout(n9274),.clk(gclk));
	jand g09037(.dina(n9274),.dinb(n9273),.dout(n9275),.clk(gclk));
	jor g09038(.dina(n9275),.dinb(n9225),.dout(n9276),.clk(gclk));
	jor g09039(.dina(n9276),.dinb(w_asqrt38_26[0]),.dout(n9277),.clk(gclk));
	jand g09040(.dina(w_n8983_0[1]),.dinb(n9277),.dout(n9278),.clk(gclk));
	jor g09041(.dina(n9278),.dinb(n9224),.dout(n9279),.clk(gclk));
	jor g09042(.dina(n9279),.dinb(w_asqrt39_22[2]),.dout(n9280),.clk(gclk));
	jnot g09043(.din(w_n8991_0[1]),.dout(n9281),.clk(gclk));
	jand g09044(.dina(n9281),.dinb(n9280),.dout(n9282),.clk(gclk));
	jor g09045(.dina(n9282),.dinb(n9223),.dout(n9283),.clk(gclk));
	jor g09046(.dina(n9283),.dinb(w_asqrt40_26[0]),.dout(n9284),.clk(gclk));
	jand g09047(.dina(w_n8998_0[1]),.dinb(n9284),.dout(n9285),.clk(gclk));
	jor g09048(.dina(n9285),.dinb(n9222),.dout(n9286),.clk(gclk));
	jor g09049(.dina(n9286),.dinb(w_asqrt41_23[0]),.dout(n9287),.clk(gclk));
	jand g09050(.dina(w_n9006_0[1]),.dinb(n9287),.dout(n9288),.clk(gclk));
	jor g09051(.dina(n9288),.dinb(n9221),.dout(n9289),.clk(gclk));
	jor g09052(.dina(n9289),.dinb(w_asqrt42_26[1]),.dout(n9290),.clk(gclk));
	jand g09053(.dina(w_n9014_0[0]),.dinb(n9290),.dout(n9291),.clk(gclk));
	jor g09054(.dina(n9291),.dinb(n9220),.dout(n9292),.clk(gclk));
	jor g09055(.dina(n9292),.dinb(w_asqrt43_23[1]),.dout(n9293),.clk(gclk));
	jnot g09056(.din(w_n9022_0[1]),.dout(n9294),.clk(gclk));
	jand g09057(.dina(n9294),.dinb(n9293),.dout(n9295),.clk(gclk));
	jor g09058(.dina(n9295),.dinb(n9219),.dout(n9296),.clk(gclk));
	jor g09059(.dina(n9296),.dinb(w_asqrt44_26[1]),.dout(n9297),.clk(gclk));
	jand g09060(.dina(w_n9029_0[1]),.dinb(n9297),.dout(n9298),.clk(gclk));
	jor g09061(.dina(n9298),.dinb(n9218),.dout(n9299),.clk(gclk));
	jor g09062(.dina(n9299),.dinb(w_asqrt45_24[0]),.dout(n9300),.clk(gclk));
	jnot g09063(.din(w_n9037_0[1]),.dout(n9301),.clk(gclk));
	jand g09064(.dina(n9301),.dinb(n9300),.dout(n9302),.clk(gclk));
	jor g09065(.dina(n9302),.dinb(n9217),.dout(n9303),.clk(gclk));
	jor g09066(.dina(n9303),.dinb(w_asqrt46_26[1]),.dout(n9304),.clk(gclk));
	jand g09067(.dina(w_n9044_0[1]),.dinb(n9304),.dout(n9305),.clk(gclk));
	jor g09068(.dina(n9305),.dinb(n9216),.dout(n9306),.clk(gclk));
	jor g09069(.dina(n9306),.dinb(w_asqrt47_24[2]),.dout(n9307),.clk(gclk));
	jnot g09070(.din(w_n9052_0[1]),.dout(n9308),.clk(gclk));
	jand g09071(.dina(n9308),.dinb(n9307),.dout(n9309),.clk(gclk));
	jor g09072(.dina(n9309),.dinb(n9215),.dout(n9310),.clk(gclk));
	jor g09073(.dina(n9310),.dinb(w_asqrt48_26[2]),.dout(n9311),.clk(gclk));
	jand g09074(.dina(w_n9059_0[1]),.dinb(n9311),.dout(n9312),.clk(gclk));
	jor g09075(.dina(n9312),.dinb(n9214),.dout(n9313),.clk(gclk));
	jor g09076(.dina(n9313),.dinb(w_asqrt49_25[0]),.dout(n9314),.clk(gclk));
	jnot g09077(.din(w_n9067_0[1]),.dout(n9315),.clk(gclk));
	jand g09078(.dina(n9315),.dinb(n9314),.dout(n9316),.clk(gclk));
	jor g09079(.dina(n9316),.dinb(n9213),.dout(n9317),.clk(gclk));
	jor g09080(.dina(n9317),.dinb(w_asqrt50_27[0]),.dout(n9318),.clk(gclk));
	jand g09081(.dina(w_n9074_0[1]),.dinb(n9318),.dout(n9319),.clk(gclk));
	jor g09082(.dina(n9319),.dinb(n9212),.dout(n9320),.clk(gclk));
	jor g09083(.dina(n9320),.dinb(w_asqrt51_25[1]),.dout(n9321),.clk(gclk));
	jand g09084(.dina(w_n9082_0[1]),.dinb(n9321),.dout(n9322),.clk(gclk));
	jor g09085(.dina(n9322),.dinb(n9211),.dout(n9323),.clk(gclk));
	jor g09086(.dina(n9323),.dinb(w_asqrt52_27[0]),.dout(n9324),.clk(gclk));
	jand g09087(.dina(w_n9090_0[1]),.dinb(n9324),.dout(n9325),.clk(gclk));
	jor g09088(.dina(n9325),.dinb(n9210),.dout(n9326),.clk(gclk));
	jor g09089(.dina(n9326),.dinb(w_asqrt53_26[0]),.dout(n9327),.clk(gclk));
	jnot g09090(.din(w_n9098_0[1]),.dout(n9328),.clk(gclk));
	jand g09091(.dina(n9328),.dinb(n9327),.dout(n9329),.clk(gclk));
	jor g09092(.dina(n9329),.dinb(n9209),.dout(n9330),.clk(gclk));
	jor g09093(.dina(n9330),.dinb(w_asqrt54_27[0]),.dout(n9331),.clk(gclk));
	jnot g09094(.din(w_n9105_0[1]),.dout(n9332),.clk(gclk));
	jand g09095(.dina(n9332),.dinb(n9331),.dout(n9333),.clk(gclk));
	jor g09096(.dina(n9333),.dinb(n9208),.dout(n9334),.clk(gclk));
	jor g09097(.dina(n9334),.dinb(w_asqrt55_26[1]),.dout(n9335),.clk(gclk));
	jnot g09098(.din(w_n9112_0[1]),.dout(n9336),.clk(gclk));
	jand g09099(.dina(n9336),.dinb(n9335),.dout(n9337),.clk(gclk));
	jor g09100(.dina(n9337),.dinb(n9207),.dout(n9338),.clk(gclk));
	jor g09101(.dina(n9338),.dinb(w_asqrt56_27[1]),.dout(n9339),.clk(gclk));
	jand g09102(.dina(w_n9119_0[1]),.dinb(n9339),.dout(n9340),.clk(gclk));
	jor g09103(.dina(n9340),.dinb(n9206),.dout(n9341),.clk(gclk));
	jor g09104(.dina(n9341),.dinb(w_asqrt57_27[0]),.dout(n9342),.clk(gclk));
	jnot g09105(.din(w_n9127_0[1]),.dout(n9343),.clk(gclk));
	jand g09106(.dina(n9343),.dinb(n9342),.dout(n9344),.clk(gclk));
	jor g09107(.dina(n9344),.dinb(n9205),.dout(n9345),.clk(gclk));
	jor g09108(.dina(n9345),.dinb(w_asqrt58_27[2]),.dout(n9346),.clk(gclk));
	jand g09109(.dina(w_n9134_0[0]),.dinb(n9346),.dout(n9347),.clk(gclk));
	jor g09110(.dina(n9347),.dinb(n9204),.dout(n9348),.clk(gclk));
	jor g09111(.dina(n9348),.dinb(w_asqrt59_27[1]),.dout(n9349),.clk(gclk));
	jnot g09112(.din(w_n9142_0[1]),.dout(n9350),.clk(gclk));
	jand g09113(.dina(n9350),.dinb(n9349),.dout(n9351),.clk(gclk));
	jor g09114(.dina(n9351),.dinb(n9203),.dout(n9352),.clk(gclk));
	jor g09115(.dina(n9352),.dinb(w_asqrt60_27[2]),.dout(n9353),.clk(gclk));
	jand g09116(.dina(w_n9149_0[1]),.dinb(n9353),.dout(n9354),.clk(gclk));
	jor g09117(.dina(n9354),.dinb(n9202),.dout(n9355),.clk(gclk));
	jor g09118(.dina(n9355),.dinb(w_asqrt61_27[2]),.dout(n9356),.clk(gclk));
	jand g09119(.dina(w_n9157_0[1]),.dinb(n9356),.dout(n9357),.clk(gclk));
	jor g09120(.dina(n9357),.dinb(n9201),.dout(n9358),.clk(gclk));
	jor g09121(.dina(n9358),.dinb(w_asqrt62_27[2]),.dout(n9359),.clk(gclk));
	jand g09122(.dina(w_n9184_0[0]),.dinb(n9359),.dout(n9360),.clk(gclk));
	jor g09123(.dina(n9360),.dinb(n9200),.dout(n9361),.clk(gclk));
	jand g09124(.dina(n9361),.dinb(w_n8893_0[0]),.dout(n9362),.clk(gclk));
	jnot g09125(.din(w_n9177_0[0]),.dout(n9363),.clk(gclk));
	jand g09126(.dina(n9363),.dinb(n9362),.dout(n9364),.clk(gclk));
	jor g09127(.dina(n9364),.dinb(w_asqrt63_35[0]),.dout(n9365),.clk(gclk));
	jnot g09128(.din(w_n9180_0[0]),.dout(n9366),.clk(gclk));
	jand g09129(.dina(n9366),.dinb(w_n9365_0[1]),.dout(n9367),.clk(gclk));
	jand g09130(.dina(n9367),.dinb(w_n9173_0[0]),.dout(n9368),.clk(gclk));
	jand g09131(.dina(w_n9368_0[1]),.dinb(w_n9199_0[1]),.dout(n9369),.clk(gclk));
	jor g09132(.dina(w_n9369_33[1]),.dinb(n9198),.dout(n9370),.clk(gclk));
	jand g09133(.dina(n9370),.dinb(n9197),.dout(n9371),.clk(gclk));
	jand g09134(.dina(n9371),.dinb(n9195),.dout(n9372),.clk(gclk));
	jor g09135(.dina(n9372),.dinb(w_n9194_0[1]),.dout(n9373),.clk(gclk));
	jand g09136(.dina(w_n9373_0[2]),.dinb(w_asqrt28_24[2]),.dout(n9374),.clk(gclk));
	jor g09137(.dina(w_n9373_0[1]),.dinb(w_asqrt28_24[1]),.dout(n9375),.clk(gclk));
	jand g09138(.dina(w_asqrt26_35[1]),.dinb(w_n8897_0[0]),.dout(n9376),.clk(gclk));
	jand g09139(.dina(w_n9172_0[0]),.dinb(w_n9199_0[0]),.dout(n9377),.clk(gclk));
	jand g09140(.dina(n9377),.dinb(w_n9365_0[0]),.dout(n9378),.clk(gclk));
	jand g09141(.dina(n9378),.dinb(w_asqrt27_18[2]),.dout(n9379),.clk(gclk));
	jor g09142(.dina(n9379),.dinb(w_n9376_0[1]),.dout(n9380),.clk(gclk));
	jxor g09143(.dina(n9380),.dinb(w_a54_0[1]),.dout(n9381),.clk(gclk));
	jnot g09144(.din(w_n9381_0[1]),.dout(n9382),.clk(gclk));
	jand g09145(.dina(w_n9382_0[1]),.dinb(n9375),.dout(n9383),.clk(gclk));
	jor g09146(.dina(n9383),.dinb(w_n9374_0[1]),.dout(n9384),.clk(gclk));
	jand g09147(.dina(w_n9384_0[2]),.dinb(w_asqrt29_19[1]),.dout(n9385),.clk(gclk));
	jor g09148(.dina(w_n9384_0[1]),.dinb(w_asqrt29_19[0]),.dout(n9386),.clk(gclk));
	jxor g09149(.dina(w_n8901_0[0]),.dinb(w_n8449_33[0]),.dout(n9387),.clk(gclk));
	jand g09150(.dina(n9387),.dinb(w_asqrt26_35[0]),.dout(n9388),.clk(gclk));
	jxor g09151(.dina(n9388),.dinb(w_n9240_0[0]),.dout(n9389),.clk(gclk));
	jand g09152(.dina(w_n9389_0[2]),.dinb(n9386),.dout(n9390),.clk(gclk));
	jor g09153(.dina(n9390),.dinb(w_n9385_0[1]),.dout(n9391),.clk(gclk));
	jand g09154(.dina(w_n9391_0[2]),.dinb(w_asqrt30_25[0]),.dout(n9392),.clk(gclk));
	jor g09155(.dina(w_n9391_0[1]),.dinb(w_asqrt30_24[2]),.dout(n9393),.clk(gclk));
	jxor g09156(.dina(w_n8909_0[0]),.dinb(w_n8003_38[2]),.dout(n9394),.clk(gclk));
	jand g09157(.dina(n9394),.dinb(w_asqrt26_34[2]),.dout(n9395),.clk(gclk));
	jxor g09158(.dina(n9395),.dinb(w_n8918_0[0]),.dout(n9396),.clk(gclk));
	jnot g09159(.din(w_n9396_0[1]),.dout(n9397),.clk(gclk));
	jand g09160(.dina(w_n9397_0[1]),.dinb(n9393),.dout(n9398),.clk(gclk));
	jor g09161(.dina(n9398),.dinb(w_n9392_0[1]),.dout(n9399),.clk(gclk));
	jand g09162(.dina(w_n9399_0[2]),.dinb(w_asqrt31_20[0]),.dout(n9400),.clk(gclk));
	jor g09163(.dina(w_n9399_0[1]),.dinb(w_asqrt31_19[2]),.dout(n9401),.clk(gclk));
	jxor g09164(.dina(w_n8920_0[0]),.dinb(w_n7581_34[0]),.dout(n9402),.clk(gclk));
	jand g09165(.dina(n9402),.dinb(w_asqrt26_34[1]),.dout(n9403),.clk(gclk));
	jxor g09166(.dina(n9403),.dinb(w_n8925_0[0]),.dout(n9404),.clk(gclk));
	jand g09167(.dina(w_n9404_0[1]),.dinb(n9401),.dout(n9405),.clk(gclk));
	jor g09168(.dina(n9405),.dinb(w_n9400_0[1]),.dout(n9406),.clk(gclk));
	jand g09169(.dina(w_n9406_0[2]),.dinb(w_asqrt32_25[0]),.dout(n9407),.clk(gclk));
	jor g09170(.dina(w_n9406_0[1]),.dinb(w_asqrt32_24[2]),.dout(n9408),.clk(gclk));
	jxor g09171(.dina(w_n8928_0[0]),.dinb(w_n7154_39[0]),.dout(n9409),.clk(gclk));
	jand g09172(.dina(n9409),.dinb(w_asqrt26_34[0]),.dout(n9410),.clk(gclk));
	jxor g09173(.dina(n9410),.dinb(w_n8933_0[0]),.dout(n9411),.clk(gclk));
	jnot g09174(.din(w_n9411_0[1]),.dout(n9412),.clk(gclk));
	jand g09175(.dina(w_n9412_0[1]),.dinb(n9408),.dout(n9413),.clk(gclk));
	jor g09176(.dina(n9413),.dinb(w_n9407_0[1]),.dout(n9414),.clk(gclk));
	jand g09177(.dina(w_n9414_0[2]),.dinb(w_asqrt33_20[2]),.dout(n9415),.clk(gclk));
	jor g09178(.dina(w_n9414_0[1]),.dinb(w_asqrt33_20[1]),.dout(n9416),.clk(gclk));
	jxor g09179(.dina(w_n8935_0[0]),.dinb(w_n6758_34[2]),.dout(n9417),.clk(gclk));
	jand g09180(.dina(n9417),.dinb(w_asqrt26_33[2]),.dout(n9418),.clk(gclk));
	jxor g09181(.dina(n9418),.dinb(w_n8940_0[0]),.dout(n9419),.clk(gclk));
	jnot g09182(.din(w_n9419_0[1]),.dout(n9420),.clk(gclk));
	jand g09183(.dina(w_n9420_0[1]),.dinb(n9416),.dout(n9421),.clk(gclk));
	jor g09184(.dina(n9421),.dinb(w_n9415_0[1]),.dout(n9422),.clk(gclk));
	jand g09185(.dina(w_n9422_0[2]),.dinb(w_asqrt34_25[1]),.dout(n9423),.clk(gclk));
	jor g09186(.dina(w_n9422_0[1]),.dinb(w_asqrt34_25[0]),.dout(n9424),.clk(gclk));
	jxor g09187(.dina(w_n8942_0[0]),.dinb(w_n6357_39[1]),.dout(n9425),.clk(gclk));
	jand g09188(.dina(n9425),.dinb(w_asqrt26_33[1]),.dout(n9426),.clk(gclk));
	jxor g09189(.dina(n9426),.dinb(w_n8947_0[0]),.dout(n9427),.clk(gclk));
	jnot g09190(.din(w_n9427_0[1]),.dout(n9428),.clk(gclk));
	jand g09191(.dina(w_n9428_0[1]),.dinb(n9424),.dout(n9429),.clk(gclk));
	jor g09192(.dina(n9429),.dinb(w_n9423_0[1]),.dout(n9430),.clk(gclk));
	jand g09193(.dina(w_n9430_0[2]),.dinb(w_asqrt35_21[1]),.dout(n9431),.clk(gclk));
	jor g09194(.dina(w_n9430_0[1]),.dinb(w_asqrt35_21[0]),.dout(n9432),.clk(gclk));
	jxor g09195(.dina(w_n8949_0[0]),.dinb(w_n5989_35[1]),.dout(n9433),.clk(gclk));
	jand g09196(.dina(n9433),.dinb(w_asqrt26_33[0]),.dout(n9434),.clk(gclk));
	jxor g09197(.dina(n9434),.dinb(w_n8954_0[0]),.dout(n9435),.clk(gclk));
	jnot g09198(.din(w_n9435_0[1]),.dout(n9436),.clk(gclk));
	jand g09199(.dina(w_n9436_0[1]),.dinb(n9432),.dout(n9437),.clk(gclk));
	jor g09200(.dina(n9437),.dinb(w_n9431_0[1]),.dout(n9438),.clk(gclk));
	jand g09201(.dina(w_n9438_0[2]),.dinb(w_asqrt36_25[1]),.dout(n9439),.clk(gclk));
	jor g09202(.dina(w_n9438_0[1]),.dinb(w_asqrt36_25[0]),.dout(n9440),.clk(gclk));
	jxor g09203(.dina(w_n8956_0[0]),.dinb(w_n5606_39[2]),.dout(n9441),.clk(gclk));
	jand g09204(.dina(n9441),.dinb(w_asqrt26_32[2]),.dout(n9442),.clk(gclk));
	jxor g09205(.dina(n9442),.dinb(w_n8961_0[0]),.dout(n9443),.clk(gclk));
	jnot g09206(.din(w_n9443_0[1]),.dout(n9444),.clk(gclk));
	jand g09207(.dina(w_n9444_0[1]),.dinb(n9440),.dout(n9445),.clk(gclk));
	jor g09208(.dina(n9445),.dinb(w_n9439_0[1]),.dout(n9446),.clk(gclk));
	jand g09209(.dina(w_n9446_0[2]),.dinb(w_asqrt37_21[2]),.dout(n9447),.clk(gclk));
	jxor g09210(.dina(w_n8963_0[0]),.dinb(w_n5259_36[1]),.dout(n9448),.clk(gclk));
	jand g09211(.dina(n9448),.dinb(w_asqrt26_32[1]),.dout(n9449),.clk(gclk));
	jxor g09212(.dina(n9449),.dinb(w_n8967_0[0]),.dout(n9450),.clk(gclk));
	jor g09213(.dina(w_n9446_0[1]),.dinb(w_asqrt37_21[1]),.dout(n9451),.clk(gclk));
	jand g09214(.dina(n9451),.dinb(w_n9450_0[1]),.dout(n9452),.clk(gclk));
	jor g09215(.dina(n9452),.dinb(w_n9447_0[1]),.dout(n9453),.clk(gclk));
	jand g09216(.dina(w_n9453_0[2]),.dinb(w_asqrt38_25[2]),.dout(n9454),.clk(gclk));
	jor g09217(.dina(w_n9453_0[1]),.dinb(w_asqrt38_25[1]),.dout(n9455),.clk(gclk));
	jxor g09218(.dina(w_n8971_0[0]),.dinb(w_n4902_40[1]),.dout(n9456),.clk(gclk));
	jand g09219(.dina(n9456),.dinb(w_asqrt26_32[0]),.dout(n9457),.clk(gclk));
	jxor g09220(.dina(n9457),.dinb(w_n8976_0[0]),.dout(n9458),.clk(gclk));
	jnot g09221(.din(w_n9458_0[1]),.dout(n9459),.clk(gclk));
	jand g09222(.dina(w_n9459_0[1]),.dinb(n9455),.dout(n9460),.clk(gclk));
	jor g09223(.dina(n9460),.dinb(w_n9454_0[1]),.dout(n9461),.clk(gclk));
	jand g09224(.dina(w_n9461_0[2]),.dinb(w_asqrt39_22[1]),.dout(n9462),.clk(gclk));
	jor g09225(.dina(w_n9461_0[1]),.dinb(w_asqrt39_22[0]),.dout(n9463),.clk(gclk));
	jxor g09226(.dina(w_n8978_0[0]),.dinb(w_n4582_37[1]),.dout(n9464),.clk(gclk));
	jand g09227(.dina(n9464),.dinb(w_asqrt26_31[2]),.dout(n9465),.clk(gclk));
	jxor g09228(.dina(n9465),.dinb(w_n8983_0[0]),.dout(n9466),.clk(gclk));
	jand g09229(.dina(w_n9466_0[1]),.dinb(n9463),.dout(n9467),.clk(gclk));
	jor g09230(.dina(n9467),.dinb(w_n9462_0[1]),.dout(n9468),.clk(gclk));
	jand g09231(.dina(w_n9468_0[2]),.dinb(w_asqrt40_25[2]),.dout(n9469),.clk(gclk));
	jor g09232(.dina(w_n9468_0[1]),.dinb(w_asqrt40_25[1]),.dout(n9470),.clk(gclk));
	jxor g09233(.dina(w_n8986_0[0]),.dinb(w_n4249_41[0]),.dout(n9471),.clk(gclk));
	jand g09234(.dina(n9471),.dinb(w_asqrt26_31[1]),.dout(n9472),.clk(gclk));
	jxor g09235(.dina(n9472),.dinb(w_n8991_0[0]),.dout(n9473),.clk(gclk));
	jnot g09236(.din(w_n9473_0[1]),.dout(n9474),.clk(gclk));
	jand g09237(.dina(w_n9474_0[1]),.dinb(n9470),.dout(n9475),.clk(gclk));
	jor g09238(.dina(n9475),.dinb(w_n9469_0[1]),.dout(n9476),.clk(gclk));
	jand g09239(.dina(w_n9476_0[2]),.dinb(w_asqrt41_22[2]),.dout(n9477),.clk(gclk));
	jor g09240(.dina(w_n9476_0[1]),.dinb(w_asqrt41_22[1]),.dout(n9478),.clk(gclk));
	jxor g09241(.dina(w_n8993_0[0]),.dinb(w_n3955_38[0]),.dout(n9479),.clk(gclk));
	jand g09242(.dina(n9479),.dinb(w_asqrt26_31[0]),.dout(n9480),.clk(gclk));
	jxor g09243(.dina(n9480),.dinb(w_n8998_0[0]),.dout(n9481),.clk(gclk));
	jand g09244(.dina(w_n9481_0[1]),.dinb(n9478),.dout(n9482),.clk(gclk));
	jor g09245(.dina(n9482),.dinb(w_n9477_0[1]),.dout(n9483),.clk(gclk));
	jand g09246(.dina(w_n9483_0[2]),.dinb(w_asqrt42_26[0]),.dout(n9484),.clk(gclk));
	jor g09247(.dina(w_n9483_0[1]),.dinb(w_asqrt42_25[2]),.dout(n9485),.clk(gclk));
	jxor g09248(.dina(w_n9001_0[0]),.dinb(w_n3642_41[1]),.dout(n9486),.clk(gclk));
	jand g09249(.dina(n9486),.dinb(w_asqrt26_30[2]),.dout(n9487),.clk(gclk));
	jxor g09250(.dina(n9487),.dinb(w_n9006_0[0]),.dout(n9488),.clk(gclk));
	jand g09251(.dina(w_n9488_0[2]),.dinb(n9485),.dout(n9489),.clk(gclk));
	jor g09252(.dina(n9489),.dinb(w_n9484_0[1]),.dout(n9490),.clk(gclk));
	jand g09253(.dina(w_n9490_0[2]),.dinb(w_asqrt43_23[0]),.dout(n9491),.clk(gclk));
	jor g09254(.dina(w_n9490_0[1]),.dinb(w_asqrt43_22[2]),.dout(n9492),.clk(gclk));
	jxor g09255(.dina(w_n9009_0[0]),.dinb(w_n3368_38[2]),.dout(n9493),.clk(gclk));
	jand g09256(.dina(n9493),.dinb(w_asqrt26_30[1]),.dout(n9494),.clk(gclk));
	jxor g09257(.dina(n9494),.dinb(w_n9015_0[0]),.dout(n9495),.clk(gclk));
	jnot g09258(.din(w_n9495_0[1]),.dout(n9496),.clk(gclk));
	jand g09259(.dina(w_n9496_0[1]),.dinb(n9492),.dout(n9497),.clk(gclk));
	jor g09260(.dina(n9497),.dinb(w_n9491_0[1]),.dout(n9498),.clk(gclk));
	jand g09261(.dina(w_n9498_0[2]),.dinb(w_asqrt44_26[0]),.dout(n9499),.clk(gclk));
	jor g09262(.dina(w_n9498_0[1]),.dinb(w_asqrt44_25[2]),.dout(n9500),.clk(gclk));
	jxor g09263(.dina(w_n9017_0[0]),.dinb(w_n3089_42[0]),.dout(n9501),.clk(gclk));
	jand g09264(.dina(n9501),.dinb(w_asqrt26_30[0]),.dout(n9502),.clk(gclk));
	jxor g09265(.dina(n9502),.dinb(w_n9022_0[0]),.dout(n9503),.clk(gclk));
	jnot g09266(.din(w_n9503_0[1]),.dout(n9504),.clk(gclk));
	jand g09267(.dina(w_n9504_0[1]),.dinb(n9500),.dout(n9505),.clk(gclk));
	jor g09268(.dina(n9505),.dinb(w_n9499_0[1]),.dout(n9506),.clk(gclk));
	jand g09269(.dina(w_n9506_0[2]),.dinb(w_asqrt45_23[2]),.dout(n9507),.clk(gclk));
	jor g09270(.dina(w_n9506_0[1]),.dinb(w_asqrt45_23[1]),.dout(n9508),.clk(gclk));
	jxor g09271(.dina(w_n9024_0[0]),.dinb(w_n2833_39[2]),.dout(n9509),.clk(gclk));
	jand g09272(.dina(n9509),.dinb(w_asqrt26_29[2]),.dout(n9510),.clk(gclk));
	jxor g09273(.dina(n9510),.dinb(w_n9029_0[0]),.dout(n9511),.clk(gclk));
	jand g09274(.dina(w_n9511_0[1]),.dinb(n9508),.dout(n9512),.clk(gclk));
	jor g09275(.dina(n9512),.dinb(w_n9507_0[1]),.dout(n9513),.clk(gclk));
	jand g09276(.dina(w_n9513_0[2]),.dinb(w_asqrt46_26[0]),.dout(n9514),.clk(gclk));
	jor g09277(.dina(w_n9513_0[1]),.dinb(w_asqrt46_25[2]),.dout(n9515),.clk(gclk));
	jxor g09278(.dina(w_n9032_0[0]),.dinb(w_n2572_42[1]),.dout(n9516),.clk(gclk));
	jand g09279(.dina(n9516),.dinb(w_asqrt26_29[1]),.dout(n9517),.clk(gclk));
	jxor g09280(.dina(n9517),.dinb(w_n9037_0[0]),.dout(n9518),.clk(gclk));
	jnot g09281(.din(w_n9518_0[1]),.dout(n9519),.clk(gclk));
	jand g09282(.dina(w_n9519_0[1]),.dinb(n9515),.dout(n9520),.clk(gclk));
	jor g09283(.dina(n9520),.dinb(w_n9514_0[1]),.dout(n9521),.clk(gclk));
	jand g09284(.dina(w_n9521_0[2]),.dinb(w_asqrt47_24[1]),.dout(n9522),.clk(gclk));
	jor g09285(.dina(w_n9521_0[1]),.dinb(w_asqrt47_24[0]),.dout(n9523),.clk(gclk));
	jxor g09286(.dina(w_n9039_0[0]),.dinb(w_n2345_40[1]),.dout(n9524),.clk(gclk));
	jand g09287(.dina(n9524),.dinb(w_asqrt26_29[0]),.dout(n9525),.clk(gclk));
	jxor g09288(.dina(n9525),.dinb(w_n9044_0[0]),.dout(n9526),.clk(gclk));
	jand g09289(.dina(w_n9526_0[1]),.dinb(n9523),.dout(n9527),.clk(gclk));
	jor g09290(.dina(n9527),.dinb(w_n9522_0[1]),.dout(n9528),.clk(gclk));
	jand g09291(.dina(w_n9528_0[2]),.dinb(w_asqrt48_26[1]),.dout(n9529),.clk(gclk));
	jor g09292(.dina(w_n9528_0[1]),.dinb(w_asqrt48_26[0]),.dout(n9530),.clk(gclk));
	jxor g09293(.dina(w_n9047_0[0]),.dinb(w_n2108_43[0]),.dout(n9531),.clk(gclk));
	jand g09294(.dina(n9531),.dinb(w_asqrt26_28[2]),.dout(n9532),.clk(gclk));
	jxor g09295(.dina(n9532),.dinb(w_n9052_0[0]),.dout(n9533),.clk(gclk));
	jnot g09296(.din(w_n9533_0[1]),.dout(n9534),.clk(gclk));
	jand g09297(.dina(w_n9534_0[1]),.dinb(n9530),.dout(n9535),.clk(gclk));
	jor g09298(.dina(n9535),.dinb(w_n9529_0[1]),.dout(n9536),.clk(gclk));
	jand g09299(.dina(w_n9536_0[2]),.dinb(w_asqrt49_24[2]),.dout(n9537),.clk(gclk));
	jor g09300(.dina(w_n9536_0[1]),.dinb(w_asqrt49_24[1]),.dout(n9538),.clk(gclk));
	jxor g09301(.dina(w_n9054_0[0]),.dinb(w_n1912_41[1]),.dout(n9539),.clk(gclk));
	jand g09302(.dina(n9539),.dinb(w_asqrt26_28[1]),.dout(n9540),.clk(gclk));
	jxor g09303(.dina(n9540),.dinb(w_n9059_0[0]),.dout(n9541),.clk(gclk));
	jand g09304(.dina(w_n9541_0[1]),.dinb(n9538),.dout(n9542),.clk(gclk));
	jor g09305(.dina(n9542),.dinb(w_n9537_0[1]),.dout(n9543),.clk(gclk));
	jand g09306(.dina(w_n9543_0[2]),.dinb(w_asqrt50_26[2]),.dout(n9544),.clk(gclk));
	jor g09307(.dina(w_n9543_0[1]),.dinb(w_asqrt50_26[1]),.dout(n9545),.clk(gclk));
	jxor g09308(.dina(w_n9062_0[0]),.dinb(w_n1699_43[2]),.dout(n9546),.clk(gclk));
	jand g09309(.dina(n9546),.dinb(w_asqrt26_28[0]),.dout(n9547),.clk(gclk));
	jxor g09310(.dina(n9547),.dinb(w_n9067_0[0]),.dout(n9548),.clk(gclk));
	jnot g09311(.din(w_n9548_0[1]),.dout(n9549),.clk(gclk));
	jand g09312(.dina(w_n9549_0[1]),.dinb(n9545),.dout(n9550),.clk(gclk));
	jor g09313(.dina(n9550),.dinb(w_n9544_0[1]),.dout(n9551),.clk(gclk));
	jand g09314(.dina(w_n9551_0[2]),.dinb(w_asqrt51_25[0]),.dout(n9552),.clk(gclk));
	jor g09315(.dina(w_n9551_0[1]),.dinb(w_asqrt51_24[2]),.dout(n9553),.clk(gclk));
	jxor g09316(.dina(w_n9069_0[0]),.dinb(w_n1516_42[0]),.dout(n9554),.clk(gclk));
	jand g09317(.dina(n9554),.dinb(w_asqrt26_27[2]),.dout(n9555),.clk(gclk));
	jxor g09318(.dina(n9555),.dinb(w_n9074_0[0]),.dout(n9556),.clk(gclk));
	jand g09319(.dina(w_n9556_0[1]),.dinb(n9553),.dout(n9557),.clk(gclk));
	jor g09320(.dina(n9557),.dinb(w_n9552_0[1]),.dout(n9558),.clk(gclk));
	jand g09321(.dina(w_n9558_0[2]),.dinb(w_asqrt52_26[2]),.dout(n9559),.clk(gclk));
	jor g09322(.dina(w_n9558_0[1]),.dinb(w_asqrt52_26[1]),.dout(n9560),.clk(gclk));
	jxor g09323(.dina(w_n9077_0[0]),.dinb(w_n1332_43[2]),.dout(n9561),.clk(gclk));
	jand g09324(.dina(n9561),.dinb(w_asqrt26_27[1]),.dout(n9562),.clk(gclk));
	jxor g09325(.dina(n9562),.dinb(w_n9082_0[0]),.dout(n9563),.clk(gclk));
	jand g09326(.dina(w_n9563_0[1]),.dinb(n9560),.dout(n9564),.clk(gclk));
	jor g09327(.dina(n9564),.dinb(w_n9559_0[1]),.dout(n9565),.clk(gclk));
	jand g09328(.dina(w_n9565_0[2]),.dinb(w_asqrt53_25[2]),.dout(n9566),.clk(gclk));
	jor g09329(.dina(w_n9565_0[1]),.dinb(w_asqrt53_25[1]),.dout(n9567),.clk(gclk));
	jxor g09330(.dina(w_n9085_0[0]),.dinb(w_n1173_42[2]),.dout(n9568),.clk(gclk));
	jand g09331(.dina(n9568),.dinb(w_asqrt26_27[0]),.dout(n9569),.clk(gclk));
	jxor g09332(.dina(n9569),.dinb(w_n9090_0[0]),.dout(n9570),.clk(gclk));
	jand g09333(.dina(w_n9570_0[1]),.dinb(n9567),.dout(n9571),.clk(gclk));
	jor g09334(.dina(n9571),.dinb(w_n9566_0[1]),.dout(n9572),.clk(gclk));
	jand g09335(.dina(w_n9572_0[2]),.dinb(w_asqrt54_26[2]),.dout(n9573),.clk(gclk));
	jor g09336(.dina(w_n9572_0[1]),.dinb(w_asqrt54_26[1]),.dout(n9574),.clk(gclk));
	jxor g09337(.dina(w_n9093_0[0]),.dinb(w_n1008_44[2]),.dout(n9575),.clk(gclk));
	jand g09338(.dina(n9575),.dinb(w_asqrt26_26[2]),.dout(n9576),.clk(gclk));
	jxor g09339(.dina(n9576),.dinb(w_n9098_0[0]),.dout(n9577),.clk(gclk));
	jnot g09340(.din(w_n9577_0[1]),.dout(n9578),.clk(gclk));
	jand g09341(.dina(w_n9578_0[1]),.dinb(n9574),.dout(n9579),.clk(gclk));
	jor g09342(.dina(n9579),.dinb(w_n9573_0[1]),.dout(n9580),.clk(gclk));
	jand g09343(.dina(w_n9580_0[2]),.dinb(w_asqrt55_26[0]),.dout(n9581),.clk(gclk));
	jor g09344(.dina(w_n9580_0[1]),.dinb(w_asqrt55_25[2]),.dout(n9582),.clk(gclk));
	jxor g09345(.dina(w_n9100_0[0]),.dinb(w_n884_43[2]),.dout(n9583),.clk(gclk));
	jand g09346(.dina(n9583),.dinb(w_asqrt26_26[1]),.dout(n9584),.clk(gclk));
	jxor g09347(.dina(n9584),.dinb(w_n9105_0[0]),.dout(n9585),.clk(gclk));
	jnot g09348(.din(w_n9585_0[1]),.dout(n9586),.clk(gclk));
	jand g09349(.dina(w_n9586_0[1]),.dinb(n9582),.dout(n9587),.clk(gclk));
	jor g09350(.dina(n9587),.dinb(w_n9581_0[1]),.dout(n9588),.clk(gclk));
	jand g09351(.dina(w_n9588_0[2]),.dinb(w_asqrt56_27[0]),.dout(n9589),.clk(gclk));
	jor g09352(.dina(w_n9588_0[1]),.dinb(w_asqrt56_26[2]),.dout(n9590),.clk(gclk));
	jxor g09353(.dina(w_n9107_0[0]),.dinb(w_n743_44[2]),.dout(n9591),.clk(gclk));
	jand g09354(.dina(n9591),.dinb(w_asqrt26_26[0]),.dout(n9592),.clk(gclk));
	jxor g09355(.dina(n9592),.dinb(w_n9112_0[0]),.dout(n9593),.clk(gclk));
	jnot g09356(.din(w_n9593_0[1]),.dout(n9594),.clk(gclk));
	jand g09357(.dina(w_n9594_0[1]),.dinb(n9590),.dout(n9595),.clk(gclk));
	jor g09358(.dina(n9595),.dinb(w_n9589_0[1]),.dout(n9596),.clk(gclk));
	jand g09359(.dina(w_n9596_0[2]),.dinb(w_asqrt57_26[2]),.dout(n9597),.clk(gclk));
	jor g09360(.dina(w_n9596_0[1]),.dinb(w_asqrt57_26[1]),.dout(n9598),.clk(gclk));
	jxor g09361(.dina(w_n9114_0[0]),.dinb(w_n635_44[2]),.dout(n9599),.clk(gclk));
	jand g09362(.dina(n9599),.dinb(w_asqrt26_25[2]),.dout(n9600),.clk(gclk));
	jxor g09363(.dina(n9600),.dinb(w_n9119_0[0]),.dout(n9601),.clk(gclk));
	jand g09364(.dina(w_n9601_0[1]),.dinb(n9598),.dout(n9602),.clk(gclk));
	jor g09365(.dina(n9602),.dinb(w_n9597_0[1]),.dout(n9603),.clk(gclk));
	jand g09366(.dina(w_n9603_0[2]),.dinb(w_asqrt58_27[1]),.dout(n9604),.clk(gclk));
	jor g09367(.dina(w_n9603_0[1]),.dinb(w_asqrt58_27[0]),.dout(n9605),.clk(gclk));
	jxor g09368(.dina(w_n9122_0[0]),.dinb(w_n515_45[2]),.dout(n9606),.clk(gclk));
	jand g09369(.dina(n9606),.dinb(w_asqrt26_25[1]),.dout(n9607),.clk(gclk));
	jxor g09370(.dina(n9607),.dinb(w_n9127_0[0]),.dout(n9608),.clk(gclk));
	jnot g09371(.din(w_n9608_0[1]),.dout(n9609),.clk(gclk));
	jand g09372(.dina(w_n9609_0[1]),.dinb(n9605),.dout(n9610),.clk(gclk));
	jor g09373(.dina(n9610),.dinb(w_n9604_0[1]),.dout(n9611),.clk(gclk));
	jand g09374(.dina(w_n9611_0[2]),.dinb(w_asqrt59_27[0]),.dout(n9612),.clk(gclk));
	jor g09375(.dina(w_n9611_0[1]),.dinb(w_asqrt59_26[2]),.dout(n9613),.clk(gclk));
	jxor g09376(.dina(w_n9129_0[0]),.dinb(w_n443_45[2]),.dout(n9614),.clk(gclk));
	jand g09377(.dina(n9614),.dinb(w_asqrt26_25[0]),.dout(n9615),.clk(gclk));
	jxor g09378(.dina(n9615),.dinb(w_n9135_0[0]),.dout(n9616),.clk(gclk));
	jnot g09379(.din(w_n9616_0[1]),.dout(n9617),.clk(gclk));
	jand g09380(.dina(w_n9617_0[1]),.dinb(n9613),.dout(n9618),.clk(gclk));
	jor g09381(.dina(n9618),.dinb(w_n9612_0[1]),.dout(n9619),.clk(gclk));
	jand g09382(.dina(w_n9619_0[2]),.dinb(w_asqrt60_27[1]),.dout(n9620),.clk(gclk));
	jor g09383(.dina(w_n9619_0[1]),.dinb(w_asqrt60_27[0]),.dout(n9621),.clk(gclk));
	jxor g09384(.dina(w_n9137_0[0]),.dinb(w_n352_46[0]),.dout(n9622),.clk(gclk));
	jand g09385(.dina(n9622),.dinb(w_asqrt26_24[2]),.dout(n9623),.clk(gclk));
	jxor g09386(.dina(n9623),.dinb(w_n9142_0[0]),.dout(n9624),.clk(gclk));
	jnot g09387(.din(w_n9624_0[1]),.dout(n9625),.clk(gclk));
	jand g09388(.dina(w_n9625_0[1]),.dinb(n9621),.dout(n9626),.clk(gclk));
	jor g09389(.dina(n9626),.dinb(w_n9620_0[1]),.dout(n9627),.clk(gclk));
	jand g09390(.dina(w_n9627_0[2]),.dinb(w_asqrt61_27[1]),.dout(n9628),.clk(gclk));
	jor g09391(.dina(w_n9627_0[1]),.dinb(w_asqrt61_27[0]),.dout(n9629),.clk(gclk));
	jxor g09392(.dina(w_n9144_0[0]),.dinb(w_n294_46[1]),.dout(n9630),.clk(gclk));
	jand g09393(.dina(n9630),.dinb(w_asqrt26_24[1]),.dout(n9631),.clk(gclk));
	jxor g09394(.dina(n9631),.dinb(w_n9149_0[0]),.dout(n9632),.clk(gclk));
	jand g09395(.dina(w_n9632_0[1]),.dinb(n9629),.dout(n9633),.clk(gclk));
	jor g09396(.dina(n9633),.dinb(w_n9628_0[1]),.dout(n9634),.clk(gclk));
	jand g09397(.dina(w_n9634_0[2]),.dinb(w_asqrt62_27[1]),.dout(n9635),.clk(gclk));
	jor g09398(.dina(w_n9634_0[1]),.dinb(w_asqrt62_27[0]),.dout(n9636),.clk(gclk));
	jxor g09399(.dina(w_n9152_0[0]),.dinb(w_n239_46[1]),.dout(n9637),.clk(gclk));
	jand g09400(.dina(n9637),.dinb(w_asqrt26_24[0]),.dout(n9638),.clk(gclk));
	jxor g09401(.dina(n9638),.dinb(w_n9157_0[0]),.dout(n9639),.clk(gclk));
	jand g09402(.dina(w_n9639_0[2]),.dinb(n9636),.dout(n9640),.clk(gclk));
	jor g09403(.dina(n9640),.dinb(w_n9635_0[1]),.dout(n9641),.clk(gclk));
	jor g09404(.dina(w_n9641_0[1]),.dinb(w_n9187_0[2]),.dout(n9642),.clk(gclk));
	jnot g09405(.din(w_n9642_1[1]),.dout(n9643),.clk(gclk));
	jand g09406(.dina(w_n9368_0[0]),.dinb(w_n9167_0[2]),.dout(n9644),.clk(gclk));
	jnot g09407(.din(n9644),.dout(n9645),.clk(gclk));
	jxor g09408(.dina(w_n9167_0[1]),.dinb(w_n8894_0[2]),.dout(n9646),.clk(gclk));
	jand g09409(.dina(w_n9646_0[1]),.dinb(w_asqrt63_34[2]),.dout(n9647),.clk(gclk));
	jand g09410(.dina(w_n9647_0[1]),.dinb(n9645),.dout(n9648),.clk(gclk));
	jnot g09411(.din(w_n9187_0[1]),.dout(n9649),.clk(gclk));
	jnot g09412(.din(w_n9635_0[0]),.dout(n9650),.clk(gclk));
	jnot g09413(.din(w_n9628_0[0]),.dout(n9651),.clk(gclk));
	jnot g09414(.din(w_n9620_0[0]),.dout(n9652),.clk(gclk));
	jnot g09415(.din(w_n9612_0[0]),.dout(n9653),.clk(gclk));
	jnot g09416(.din(w_n9604_0[0]),.dout(n9654),.clk(gclk));
	jnot g09417(.din(w_n9597_0[0]),.dout(n9655),.clk(gclk));
	jnot g09418(.din(w_n9589_0[0]),.dout(n9656),.clk(gclk));
	jnot g09419(.din(w_n9581_0[0]),.dout(n9657),.clk(gclk));
	jnot g09420(.din(w_n9573_0[0]),.dout(n9658),.clk(gclk));
	jnot g09421(.din(w_n9566_0[0]),.dout(n9659),.clk(gclk));
	jnot g09422(.din(w_n9559_0[0]),.dout(n9660),.clk(gclk));
	jnot g09423(.din(w_n9552_0[0]),.dout(n9661),.clk(gclk));
	jnot g09424(.din(w_n9544_0[0]),.dout(n9662),.clk(gclk));
	jnot g09425(.din(w_n9537_0[0]),.dout(n9663),.clk(gclk));
	jnot g09426(.din(w_n9529_0[0]),.dout(n9664),.clk(gclk));
	jnot g09427(.din(w_n9522_0[0]),.dout(n9665),.clk(gclk));
	jnot g09428(.din(w_n9514_0[0]),.dout(n9666),.clk(gclk));
	jnot g09429(.din(w_n9507_0[0]),.dout(n9667),.clk(gclk));
	jnot g09430(.din(w_n9499_0[0]),.dout(n9668),.clk(gclk));
	jnot g09431(.din(w_n9491_0[0]),.dout(n9669),.clk(gclk));
	jnot g09432(.din(w_n9484_0[0]),.dout(n9670),.clk(gclk));
	jnot g09433(.din(w_n9477_0[0]),.dout(n9671),.clk(gclk));
	jnot g09434(.din(w_n9469_0[0]),.dout(n9672),.clk(gclk));
	jnot g09435(.din(w_n9462_0[0]),.dout(n9673),.clk(gclk));
	jnot g09436(.din(w_n9454_0[0]),.dout(n9674),.clk(gclk));
	jnot g09437(.din(w_n9447_0[0]),.dout(n9675),.clk(gclk));
	jnot g09438(.din(w_n9450_0[0]),.dout(n9676),.clk(gclk));
	jnot g09439(.din(w_n9439_0[0]),.dout(n9677),.clk(gclk));
	jnot g09440(.din(w_n9431_0[0]),.dout(n9678),.clk(gclk));
	jnot g09441(.din(w_n9423_0[0]),.dout(n9679),.clk(gclk));
	jnot g09442(.din(w_n9415_0[0]),.dout(n9680),.clk(gclk));
	jnot g09443(.din(w_n9407_0[0]),.dout(n9681),.clk(gclk));
	jnot g09444(.din(w_n9400_0[0]),.dout(n9682),.clk(gclk));
	jnot g09445(.din(w_n9392_0[0]),.dout(n9683),.clk(gclk));
	jnot g09446(.din(w_n9385_0[0]),.dout(n9684),.clk(gclk));
	jnot g09447(.din(w_n9374_0[0]),.dout(n9685),.clk(gclk));
	jnot g09448(.din(w_n9194_0[0]),.dout(n9686),.clk(gclk));
	jnot g09449(.din(w_n9191_0[0]),.dout(n9687),.clk(gclk));
	jor g09450(.dina(w_n9369_33[0]),.dinb(w_n8895_0[2]),.dout(n9688),.clk(gclk));
	jand g09451(.dina(n9688),.dinb(n9687),.dout(n9689),.clk(gclk));
	jand g09452(.dina(n9689),.dinb(w_n8890_37[2]),.dout(n9690),.clk(gclk));
	jor g09453(.dina(w_n9369_32[2]),.dinb(w_a52_0[0]),.dout(n9691),.clk(gclk));
	jand g09454(.dina(n9691),.dinb(w_a53_0[0]),.dout(n9692),.clk(gclk));
	jor g09455(.dina(w_n9376_0[0]),.dinb(n9692),.dout(n9693),.clk(gclk));
	jor g09456(.dina(w_n9693_0[1]),.dinb(n9690),.dout(n9694),.clk(gclk));
	jand g09457(.dina(n9694),.dinb(n9686),.dout(n9695),.clk(gclk));
	jand g09458(.dina(n9695),.dinb(w_n8449_32[2]),.dout(n9696),.clk(gclk));
	jor g09459(.dina(w_n9381_0[0]),.dinb(n9696),.dout(n9697),.clk(gclk));
	jand g09460(.dina(n9697),.dinb(n9685),.dout(n9698),.clk(gclk));
	jand g09461(.dina(n9698),.dinb(w_n8003_38[1]),.dout(n9699),.clk(gclk));
	jnot g09462(.din(w_n9389_0[1]),.dout(n9700),.clk(gclk));
	jor g09463(.dina(n9700),.dinb(n9699),.dout(n9701),.clk(gclk));
	jand g09464(.dina(n9701),.dinb(n9684),.dout(n9702),.clk(gclk));
	jand g09465(.dina(n9702),.dinb(w_n7581_33[2]),.dout(n9703),.clk(gclk));
	jor g09466(.dina(w_n9396_0[0]),.dinb(n9703),.dout(n9704),.clk(gclk));
	jand g09467(.dina(n9704),.dinb(n9683),.dout(n9705),.clk(gclk));
	jand g09468(.dina(n9705),.dinb(w_n7154_38[2]),.dout(n9706),.clk(gclk));
	jnot g09469(.din(w_n9404_0[0]),.dout(n9707),.clk(gclk));
	jor g09470(.dina(w_n9707_0[1]),.dinb(n9706),.dout(n9708),.clk(gclk));
	jand g09471(.dina(n9708),.dinb(n9682),.dout(n9709),.clk(gclk));
	jand g09472(.dina(n9709),.dinb(w_n6758_34[1]),.dout(n9710),.clk(gclk));
	jor g09473(.dina(w_n9411_0[0]),.dinb(n9710),.dout(n9711),.clk(gclk));
	jand g09474(.dina(n9711),.dinb(n9681),.dout(n9712),.clk(gclk));
	jand g09475(.dina(n9712),.dinb(w_n6357_39[0]),.dout(n9713),.clk(gclk));
	jor g09476(.dina(w_n9419_0[0]),.dinb(n9713),.dout(n9714),.clk(gclk));
	jand g09477(.dina(n9714),.dinb(n9680),.dout(n9715),.clk(gclk));
	jand g09478(.dina(n9715),.dinb(w_n5989_35[0]),.dout(n9716),.clk(gclk));
	jor g09479(.dina(w_n9427_0[0]),.dinb(n9716),.dout(n9717),.clk(gclk));
	jand g09480(.dina(n9717),.dinb(n9679),.dout(n9718),.clk(gclk));
	jand g09481(.dina(n9718),.dinb(w_n5606_39[1]),.dout(n9719),.clk(gclk));
	jor g09482(.dina(w_n9435_0[0]),.dinb(n9719),.dout(n9720),.clk(gclk));
	jand g09483(.dina(n9720),.dinb(n9678),.dout(n9721),.clk(gclk));
	jand g09484(.dina(n9721),.dinb(w_n5259_36[0]),.dout(n9722),.clk(gclk));
	jor g09485(.dina(w_n9443_0[0]),.dinb(n9722),.dout(n9723),.clk(gclk));
	jand g09486(.dina(n9723),.dinb(n9677),.dout(n9724),.clk(gclk));
	jand g09487(.dina(n9724),.dinb(w_n4902_40[0]),.dout(n9725),.clk(gclk));
	jor g09488(.dina(n9725),.dinb(w_n9676_0[1]),.dout(n9726),.clk(gclk));
	jand g09489(.dina(n9726),.dinb(n9675),.dout(n9727),.clk(gclk));
	jand g09490(.dina(n9727),.dinb(w_n4582_37[0]),.dout(n9728),.clk(gclk));
	jor g09491(.dina(w_n9458_0[0]),.dinb(n9728),.dout(n9729),.clk(gclk));
	jand g09492(.dina(n9729),.dinb(n9674),.dout(n9730),.clk(gclk));
	jand g09493(.dina(n9730),.dinb(w_n4249_40[2]),.dout(n9731),.clk(gclk));
	jnot g09494(.din(w_n9466_0[0]),.dout(n9732),.clk(gclk));
	jor g09495(.dina(w_n9732_0[1]),.dinb(n9731),.dout(n9733),.clk(gclk));
	jand g09496(.dina(n9733),.dinb(n9673),.dout(n9734),.clk(gclk));
	jand g09497(.dina(n9734),.dinb(w_n3955_37[2]),.dout(n9735),.clk(gclk));
	jor g09498(.dina(w_n9473_0[0]),.dinb(n9735),.dout(n9736),.clk(gclk));
	jand g09499(.dina(n9736),.dinb(n9672),.dout(n9737),.clk(gclk));
	jand g09500(.dina(n9737),.dinb(w_n3642_41[0]),.dout(n9738),.clk(gclk));
	jnot g09501(.din(w_n9481_0[0]),.dout(n9739),.clk(gclk));
	jor g09502(.dina(w_n9739_0[1]),.dinb(n9738),.dout(n9740),.clk(gclk));
	jand g09503(.dina(n9740),.dinb(n9671),.dout(n9741),.clk(gclk));
	jand g09504(.dina(n9741),.dinb(w_n3368_38[1]),.dout(n9742),.clk(gclk));
	jnot g09505(.din(w_n9488_0[1]),.dout(n9743),.clk(gclk));
	jor g09506(.dina(n9743),.dinb(n9742),.dout(n9744),.clk(gclk));
	jand g09507(.dina(n9744),.dinb(n9670),.dout(n9745),.clk(gclk));
	jand g09508(.dina(n9745),.dinb(w_n3089_41[2]),.dout(n9746),.clk(gclk));
	jor g09509(.dina(w_n9495_0[0]),.dinb(n9746),.dout(n9747),.clk(gclk));
	jand g09510(.dina(n9747),.dinb(n9669),.dout(n9748),.clk(gclk));
	jand g09511(.dina(n9748),.dinb(w_n2833_39[1]),.dout(n9749),.clk(gclk));
	jor g09512(.dina(w_n9503_0[0]),.dinb(n9749),.dout(n9750),.clk(gclk));
	jand g09513(.dina(n9750),.dinb(n9668),.dout(n9751),.clk(gclk));
	jand g09514(.dina(n9751),.dinb(w_n2572_42[0]),.dout(n9752),.clk(gclk));
	jnot g09515(.din(w_n9511_0[0]),.dout(n9753),.clk(gclk));
	jor g09516(.dina(w_n9753_0[1]),.dinb(n9752),.dout(n9754),.clk(gclk));
	jand g09517(.dina(n9754),.dinb(n9667),.dout(n9755),.clk(gclk));
	jand g09518(.dina(n9755),.dinb(w_n2345_40[0]),.dout(n9756),.clk(gclk));
	jor g09519(.dina(w_n9518_0[0]),.dinb(n9756),.dout(n9757),.clk(gclk));
	jand g09520(.dina(n9757),.dinb(n9666),.dout(n9758),.clk(gclk));
	jand g09521(.dina(n9758),.dinb(w_n2108_42[2]),.dout(n9759),.clk(gclk));
	jnot g09522(.din(w_n9526_0[0]),.dout(n9760),.clk(gclk));
	jor g09523(.dina(w_n9760_0[1]),.dinb(n9759),.dout(n9761),.clk(gclk));
	jand g09524(.dina(n9761),.dinb(n9665),.dout(n9762),.clk(gclk));
	jand g09525(.dina(n9762),.dinb(w_n1912_41[0]),.dout(n9763),.clk(gclk));
	jor g09526(.dina(w_n9533_0[0]),.dinb(n9763),.dout(n9764),.clk(gclk));
	jand g09527(.dina(n9764),.dinb(n9664),.dout(n9765),.clk(gclk));
	jand g09528(.dina(n9765),.dinb(w_n1699_43[1]),.dout(n9766),.clk(gclk));
	jnot g09529(.din(w_n9541_0[0]),.dout(n9767),.clk(gclk));
	jor g09530(.dina(w_n9767_0[1]),.dinb(n9766),.dout(n9768),.clk(gclk));
	jand g09531(.dina(n9768),.dinb(n9663),.dout(n9769),.clk(gclk));
	jand g09532(.dina(n9769),.dinb(w_n1516_41[2]),.dout(n9770),.clk(gclk));
	jor g09533(.dina(w_n9548_0[0]),.dinb(n9770),.dout(n9771),.clk(gclk));
	jand g09534(.dina(n9771),.dinb(n9662),.dout(n9772),.clk(gclk));
	jand g09535(.dina(n9772),.dinb(w_n1332_43[1]),.dout(n9773),.clk(gclk));
	jnot g09536(.din(w_n9556_0[0]),.dout(n9774),.clk(gclk));
	jor g09537(.dina(w_n9774_0[1]),.dinb(n9773),.dout(n9775),.clk(gclk));
	jand g09538(.dina(n9775),.dinb(n9661),.dout(n9776),.clk(gclk));
	jand g09539(.dina(n9776),.dinb(w_n1173_42[1]),.dout(n9777),.clk(gclk));
	jnot g09540(.din(w_n9563_0[0]),.dout(n9778),.clk(gclk));
	jor g09541(.dina(w_n9778_0[1]),.dinb(n9777),.dout(n9779),.clk(gclk));
	jand g09542(.dina(n9779),.dinb(n9660),.dout(n9780),.clk(gclk));
	jand g09543(.dina(n9780),.dinb(w_n1008_44[1]),.dout(n9781),.clk(gclk));
	jnot g09544(.din(w_n9570_0[0]),.dout(n9782),.clk(gclk));
	jor g09545(.dina(w_n9782_0[1]),.dinb(n9781),.dout(n9783),.clk(gclk));
	jand g09546(.dina(n9783),.dinb(n9659),.dout(n9784),.clk(gclk));
	jand g09547(.dina(n9784),.dinb(w_n884_43[1]),.dout(n9785),.clk(gclk));
	jor g09548(.dina(w_n9577_0[0]),.dinb(n9785),.dout(n9786),.clk(gclk));
	jand g09549(.dina(n9786),.dinb(n9658),.dout(n9787),.clk(gclk));
	jand g09550(.dina(n9787),.dinb(w_n743_44[1]),.dout(n9788),.clk(gclk));
	jor g09551(.dina(w_n9585_0[0]),.dinb(n9788),.dout(n9789),.clk(gclk));
	jand g09552(.dina(n9789),.dinb(n9657),.dout(n9790),.clk(gclk));
	jand g09553(.dina(n9790),.dinb(w_n635_44[1]),.dout(n9791),.clk(gclk));
	jor g09554(.dina(w_n9593_0[0]),.dinb(n9791),.dout(n9792),.clk(gclk));
	jand g09555(.dina(n9792),.dinb(n9656),.dout(n9793),.clk(gclk));
	jand g09556(.dina(n9793),.dinb(w_n515_45[1]),.dout(n9794),.clk(gclk));
	jnot g09557(.din(w_n9601_0[0]),.dout(n9795),.clk(gclk));
	jor g09558(.dina(w_n9795_0[1]),.dinb(n9794),.dout(n9796),.clk(gclk));
	jand g09559(.dina(n9796),.dinb(n9655),.dout(n9797),.clk(gclk));
	jand g09560(.dina(n9797),.dinb(w_n443_45[1]),.dout(n9798),.clk(gclk));
	jor g09561(.dina(w_n9608_0[0]),.dinb(n9798),.dout(n9799),.clk(gclk));
	jand g09562(.dina(n9799),.dinb(n9654),.dout(n9800),.clk(gclk));
	jand g09563(.dina(n9800),.dinb(w_n352_45[2]),.dout(n9801),.clk(gclk));
	jor g09564(.dina(w_n9616_0[0]),.dinb(n9801),.dout(n9802),.clk(gclk));
	jand g09565(.dina(n9802),.dinb(n9653),.dout(n9803),.clk(gclk));
	jand g09566(.dina(n9803),.dinb(w_n294_46[0]),.dout(n9804),.clk(gclk));
	jor g09567(.dina(w_n9624_0[0]),.dinb(n9804),.dout(n9805),.clk(gclk));
	jand g09568(.dina(n9805),.dinb(n9652),.dout(n9806),.clk(gclk));
	jand g09569(.dina(n9806),.dinb(w_n239_46[0]),.dout(n9807),.clk(gclk));
	jnot g09570(.din(w_n9632_0[0]),.dout(n9808),.clk(gclk));
	jor g09571(.dina(w_n9808_0[1]),.dinb(n9807),.dout(n9809),.clk(gclk));
	jand g09572(.dina(n9809),.dinb(n9651),.dout(n9810),.clk(gclk));
	jand g09573(.dina(n9810),.dinb(w_n221_46[1]),.dout(n9811),.clk(gclk));
	jnot g09574(.din(w_n9639_0[1]),.dout(n9812),.clk(gclk));
	jor g09575(.dina(n9812),.dinb(n9811),.dout(n9813),.clk(gclk));
	jand g09576(.dina(n9813),.dinb(n9650),.dout(n9814),.clk(gclk));
	jor g09577(.dina(w_n9814_0[1]),.dinb(w_n9649_0[1]),.dout(n9815),.clk(gclk));
	jor g09578(.dina(w_n9646_0[0]),.dinb(w_n9369_32[1]),.dout(n9816),.clk(gclk));
	jnot g09579(.din(w_n9816_0[1]),.dout(n9817),.clk(gclk));
	jor g09580(.dina(n9817),.dinb(w_n9815_0[1]),.dout(n9818),.clk(gclk));
	jand g09581(.dina(n9818),.dinb(w_n218_19[1]),.dout(n9819),.clk(gclk));
	jand g09582(.dina(w_n9369_32[0]),.dinb(w_n8894_0[1]),.dout(n9820),.clk(gclk));
	jor g09583(.dina(w_n9820_0[1]),.dinb(w_n9819_0[1]),.dout(n9821),.clk(gclk));
	jor g09584(.dina(n9821),.dinb(w_n9648_0[1]),.dout(n9822),.clk(gclk));
	jor g09585(.dina(w_n9822_0[1]),.dinb(w_n9643_0[2]),.dout(asqrt_fa_26),.clk(gclk));
	jand g09586(.dina(w_n9641_0[0]),.dinb(w_n9187_0[0]),.dout(n9824),.clk(gclk));
	jand g09587(.dina(w_n9822_0[0]),.dinb(w_n9824_0[1]),.dout(n9825),.clk(gclk));
	jnot g09588(.din(w_n9648_0[0]),.dout(n9826),.clk(gclk));
	jand g09589(.dina(w_n9816_0[0]),.dinb(w_n9824_0[0]),.dout(n9827),.clk(gclk));
	jor g09590(.dina(n9827),.dinb(w_asqrt63_34[1]),.dout(n9828),.clk(gclk));
	jnot g09591(.din(w_n9820_0[0]),.dout(n9829),.clk(gclk));
	jand g09592(.dina(n9829),.dinb(n9828),.dout(n9830),.clk(gclk));
	jand g09593(.dina(n9830),.dinb(n9826),.dout(n9831),.clk(gclk));
	jand g09594(.dina(w_n9831_0[1]),.dinb(w_n9642_1[0]),.dout(n9832),.clk(gclk));
	jor g09595(.dina(w_n9832_49[1]),.dinb(w_n9188_1[1]),.dout(n9833),.clk(gclk));
	jnot g09596(.din(w_a48_0[2]),.dout(n9834),.clk(gclk));
	jnot g09597(.din(w_a49_0[1]),.dout(n9835),.clk(gclk));
	jand g09598(.dina(w_n9835_0[1]),.dinb(w_n9834_1[2]),.dout(n9836),.clk(gclk));
	jand g09599(.dina(w_n9836_0[2]),.dinb(w_n9188_1[0]),.dout(n9837),.clk(gclk));
	jnot g09600(.din(w_n9837_0[1]),.dout(n9838),.clk(gclk));
	jand g09601(.dina(n9838),.dinb(n9833),.dout(n9839),.clk(gclk));
	jor g09602(.dina(w_n9839_0[2]),.dinb(w_n9369_31[2]),.dout(n9840),.clk(gclk));
	jand g09603(.dina(w_n9839_0[1]),.dinb(w_n9369_31[1]),.dout(n9841),.clk(gclk));
	jor g09604(.dina(w_n9832_49[0]),.dinb(w_a50_0[1]),.dout(n9842),.clk(gclk));
	jand g09605(.dina(n9842),.dinb(w_a51_0[0]),.dout(n9843),.clk(gclk));
	jand g09606(.dina(w_asqrt25_18[1]),.dinb(w_n9190_0[1]),.dout(n9844),.clk(gclk));
	jor g09607(.dina(n9844),.dinb(n9843),.dout(n9845),.clk(gclk));
	jor g09608(.dina(n9845),.dinb(n9841),.dout(n9846),.clk(gclk));
	jand g09609(.dina(n9846),.dinb(w_n9840_0[1]),.dout(n9847),.clk(gclk));
	jor g09610(.dina(w_n9847_0[2]),.dinb(w_n8890_37[1]),.dout(n9848),.clk(gclk));
	jand g09611(.dina(w_n9847_0[1]),.dinb(w_n8890_37[0]),.dout(n9849),.clk(gclk));
	jnot g09612(.din(w_n9190_0[0]),.dout(n9850),.clk(gclk));
	jor g09613(.dina(w_n9832_48[2]),.dinb(n9850),.dout(n9851),.clk(gclk));
	jor g09614(.dina(w_n9647_0[0]),.dinb(w_n9643_0[1]),.dout(n9852),.clk(gclk));
	jor g09615(.dina(n9852),.dinb(w_n9819_0[0]),.dout(n9853),.clk(gclk));
	jor g09616(.dina(n9853),.dinb(w_n9369_31[0]),.dout(n9854),.clk(gclk));
	jand g09617(.dina(n9854),.dinb(w_n9851_0[1]),.dout(n9855),.clk(gclk));
	jxor g09618(.dina(n9855),.dinb(w_n8895_0[1]),.dout(n9856),.clk(gclk));
	jor g09619(.dina(w_n9856_0[2]),.dinb(n9849),.dout(n9857),.clk(gclk));
	jand g09620(.dina(n9857),.dinb(w_n9848_0[1]),.dout(n9858),.clk(gclk));
	jor g09621(.dina(w_n9858_0[2]),.dinb(w_n8449_32[1]),.dout(n9859),.clk(gclk));
	jand g09622(.dina(w_n9858_0[1]),.dinb(w_n8449_32[0]),.dout(n9860),.clk(gclk));
	jxor g09623(.dina(w_n9193_0[0]),.dinb(w_n8890_36[2]),.dout(n9861),.clk(gclk));
	jor g09624(.dina(n9861),.dinb(w_n9832_48[1]),.dout(n9862),.clk(gclk));
	jxor g09625(.dina(n9862),.dinb(w_n9693_0[0]),.dout(n9863),.clk(gclk));
	jnot g09626(.din(w_n9863_0[2]),.dout(n9864),.clk(gclk));
	jor g09627(.dina(n9864),.dinb(n9860),.dout(n9865),.clk(gclk));
	jand g09628(.dina(n9865),.dinb(w_n9859_0[1]),.dout(n9866),.clk(gclk));
	jor g09629(.dina(w_n9866_0[2]),.dinb(w_n8003_38[0]),.dout(n9867),.clk(gclk));
	jand g09630(.dina(w_n9866_0[1]),.dinb(w_n8003_37[2]),.dout(n9868),.clk(gclk));
	jxor g09631(.dina(w_n9373_0[0]),.dinb(w_n8449_31[2]),.dout(n9869),.clk(gclk));
	jor g09632(.dina(n9869),.dinb(w_n9832_48[0]),.dout(n9870),.clk(gclk));
	jxor g09633(.dina(n9870),.dinb(w_n9382_0[0]),.dout(n9871),.clk(gclk));
	jor g09634(.dina(w_n9871_0[2]),.dinb(n9868),.dout(n9872),.clk(gclk));
	jand g09635(.dina(n9872),.dinb(w_n9867_0[1]),.dout(n9873),.clk(gclk));
	jor g09636(.dina(w_n9873_0[2]),.dinb(w_n7581_33[1]),.dout(n9874),.clk(gclk));
	jand g09637(.dina(w_n9873_0[1]),.dinb(w_n7581_33[0]),.dout(n9875),.clk(gclk));
	jxor g09638(.dina(w_n9384_0[0]),.dinb(w_n8003_37[1]),.dout(n9876),.clk(gclk));
	jor g09639(.dina(n9876),.dinb(w_n9832_47[2]),.dout(n9877),.clk(gclk));
	jxor g09640(.dina(n9877),.dinb(w_n9389_0[0]),.dout(n9878),.clk(gclk));
	jor g09641(.dina(w_n9878_0[2]),.dinb(n9875),.dout(n9879),.clk(gclk));
	jand g09642(.dina(n9879),.dinb(w_n9874_0[1]),.dout(n9880),.clk(gclk));
	jor g09643(.dina(w_n9880_0[2]),.dinb(w_n7154_38[1]),.dout(n9881),.clk(gclk));
	jand g09644(.dina(w_n9880_0[1]),.dinb(w_n7154_38[0]),.dout(n9882),.clk(gclk));
	jxor g09645(.dina(w_n9391_0[0]),.dinb(w_n7581_32[2]),.dout(n9883),.clk(gclk));
	jor g09646(.dina(n9883),.dinb(w_n9832_47[1]),.dout(n9884),.clk(gclk));
	jxor g09647(.dina(n9884),.dinb(w_n9397_0[0]),.dout(n9885),.clk(gclk));
	jor g09648(.dina(w_n9885_0[2]),.dinb(n9882),.dout(n9886),.clk(gclk));
	jand g09649(.dina(n9886),.dinb(w_n9881_0[1]),.dout(n9887),.clk(gclk));
	jor g09650(.dina(w_n9887_0[2]),.dinb(w_n6758_34[0]),.dout(n9888),.clk(gclk));
	jand g09651(.dina(w_n9887_0[1]),.dinb(w_n6758_33[2]),.dout(n9889),.clk(gclk));
	jxor g09652(.dina(w_n9399_0[0]),.dinb(w_n7154_37[2]),.dout(n9890),.clk(gclk));
	jor g09653(.dina(n9890),.dinb(w_n9832_47[0]),.dout(n9891),.clk(gclk));
	jxor g09654(.dina(n9891),.dinb(w_n9707_0[0]),.dout(n9892),.clk(gclk));
	jnot g09655(.din(w_n9892_0[2]),.dout(n9893),.clk(gclk));
	jor g09656(.dina(n9893),.dinb(n9889),.dout(n9894),.clk(gclk));
	jand g09657(.dina(n9894),.dinb(w_n9888_0[1]),.dout(n9895),.clk(gclk));
	jor g09658(.dina(w_n9895_0[2]),.dinb(w_n6357_38[2]),.dout(n9896),.clk(gclk));
	jand g09659(.dina(w_n9895_0[1]),.dinb(w_n6357_38[1]),.dout(n9897),.clk(gclk));
	jxor g09660(.dina(w_n9406_0[0]),.dinb(w_n6758_33[1]),.dout(n9898),.clk(gclk));
	jor g09661(.dina(n9898),.dinb(w_n9832_46[2]),.dout(n9899),.clk(gclk));
	jxor g09662(.dina(n9899),.dinb(w_n9412_0[0]),.dout(n9900),.clk(gclk));
	jor g09663(.dina(w_n9900_0[2]),.dinb(n9897),.dout(n9901),.clk(gclk));
	jand g09664(.dina(n9901),.dinb(w_n9896_0[1]),.dout(n9902),.clk(gclk));
	jor g09665(.dina(w_n9902_0[2]),.dinb(w_n5989_34[2]),.dout(n9903),.clk(gclk));
	jand g09666(.dina(w_n9902_0[1]),.dinb(w_n5989_34[1]),.dout(n9904),.clk(gclk));
	jxor g09667(.dina(w_n9414_0[0]),.dinb(w_n6357_38[0]),.dout(n9905),.clk(gclk));
	jor g09668(.dina(n9905),.dinb(w_n9832_46[1]),.dout(n9906),.clk(gclk));
	jxor g09669(.dina(n9906),.dinb(w_n9420_0[0]),.dout(n9907),.clk(gclk));
	jor g09670(.dina(w_n9907_0[2]),.dinb(n9904),.dout(n9908),.clk(gclk));
	jand g09671(.dina(n9908),.dinb(w_n9903_0[1]),.dout(n9909),.clk(gclk));
	jor g09672(.dina(w_n9909_0[2]),.dinb(w_n5606_39[0]),.dout(n9910),.clk(gclk));
	jand g09673(.dina(w_n9909_0[1]),.dinb(w_n5606_38[2]),.dout(n9911),.clk(gclk));
	jxor g09674(.dina(w_n9422_0[0]),.dinb(w_n5989_34[0]),.dout(n9912),.clk(gclk));
	jor g09675(.dina(n9912),.dinb(w_n9832_46[0]),.dout(n9913),.clk(gclk));
	jxor g09676(.dina(n9913),.dinb(w_n9428_0[0]),.dout(n9914),.clk(gclk));
	jor g09677(.dina(w_n9914_0[2]),.dinb(n9911),.dout(n9915),.clk(gclk));
	jand g09678(.dina(n9915),.dinb(w_n9910_0[1]),.dout(n9916),.clk(gclk));
	jor g09679(.dina(w_n9916_0[2]),.dinb(w_n5259_35[2]),.dout(n9917),.clk(gclk));
	jand g09680(.dina(w_n9916_0[1]),.dinb(w_n5259_35[1]),.dout(n9918),.clk(gclk));
	jxor g09681(.dina(w_n9430_0[0]),.dinb(w_n5606_38[1]),.dout(n9919),.clk(gclk));
	jor g09682(.dina(n9919),.dinb(w_n9832_45[2]),.dout(n9920),.clk(gclk));
	jxor g09683(.dina(n9920),.dinb(w_n9436_0[0]),.dout(n9921),.clk(gclk));
	jor g09684(.dina(w_n9921_0[2]),.dinb(n9918),.dout(n9922),.clk(gclk));
	jand g09685(.dina(n9922),.dinb(w_n9917_0[1]),.dout(n9923),.clk(gclk));
	jor g09686(.dina(w_n9923_0[2]),.dinb(w_n4902_39[2]),.dout(n9924),.clk(gclk));
	jand g09687(.dina(w_n9923_0[1]),.dinb(w_n4902_39[1]),.dout(n9925),.clk(gclk));
	jxor g09688(.dina(w_n9438_0[0]),.dinb(w_n5259_35[0]),.dout(n9926),.clk(gclk));
	jor g09689(.dina(n9926),.dinb(w_n9832_45[1]),.dout(n9927),.clk(gclk));
	jxor g09690(.dina(n9927),.dinb(w_n9444_0[0]),.dout(n9928),.clk(gclk));
	jor g09691(.dina(w_n9928_0[2]),.dinb(n9925),.dout(n9929),.clk(gclk));
	jand g09692(.dina(n9929),.dinb(w_n9924_0[1]),.dout(n9930),.clk(gclk));
	jor g09693(.dina(w_n9930_0[2]),.dinb(w_n4582_36[2]),.dout(n9931),.clk(gclk));
	jxor g09694(.dina(w_n9446_0[0]),.dinb(w_n4902_39[0]),.dout(n9932),.clk(gclk));
	jor g09695(.dina(n9932),.dinb(w_n9832_45[0]),.dout(n9933),.clk(gclk));
	jxor g09696(.dina(n9933),.dinb(w_n9676_0[0]),.dout(n9934),.clk(gclk));
	jnot g09697(.din(w_n9934_0[2]),.dout(n9935),.clk(gclk));
	jand g09698(.dina(w_n9930_0[1]),.dinb(w_n4582_36[1]),.dout(n9936),.clk(gclk));
	jor g09699(.dina(n9936),.dinb(n9935),.dout(n9937),.clk(gclk));
	jand g09700(.dina(n9937),.dinb(w_n9931_0[1]),.dout(n9938),.clk(gclk));
	jor g09701(.dina(w_n9938_0[2]),.dinb(w_n4249_40[1]),.dout(n9939),.clk(gclk));
	jand g09702(.dina(w_n9938_0[1]),.dinb(w_n4249_40[0]),.dout(n9940),.clk(gclk));
	jxor g09703(.dina(w_n9453_0[0]),.dinb(w_n4582_36[0]),.dout(n9941),.clk(gclk));
	jor g09704(.dina(n9941),.dinb(w_n9832_44[2]),.dout(n9942),.clk(gclk));
	jxor g09705(.dina(n9942),.dinb(w_n9459_0[0]),.dout(n9943),.clk(gclk));
	jor g09706(.dina(w_n9943_0[2]),.dinb(n9940),.dout(n9944),.clk(gclk));
	jand g09707(.dina(n9944),.dinb(w_n9939_0[1]),.dout(n9945),.clk(gclk));
	jor g09708(.dina(w_n9945_0[2]),.dinb(w_n3955_37[1]),.dout(n9946),.clk(gclk));
	jand g09709(.dina(w_n9945_0[1]),.dinb(w_n3955_37[0]),.dout(n9947),.clk(gclk));
	jxor g09710(.dina(w_n9461_0[0]),.dinb(w_n4249_39[2]),.dout(n9948),.clk(gclk));
	jor g09711(.dina(n9948),.dinb(w_n9832_44[1]),.dout(n9949),.clk(gclk));
	jxor g09712(.dina(n9949),.dinb(w_n9732_0[0]),.dout(n9950),.clk(gclk));
	jnot g09713(.din(w_n9950_0[2]),.dout(n9951),.clk(gclk));
	jor g09714(.dina(n9951),.dinb(n9947),.dout(n9952),.clk(gclk));
	jand g09715(.dina(n9952),.dinb(w_n9946_0[1]),.dout(n9953),.clk(gclk));
	jor g09716(.dina(w_n9953_0[2]),.dinb(w_n3642_40[2]),.dout(n9954),.clk(gclk));
	jand g09717(.dina(w_n9953_0[1]),.dinb(w_n3642_40[1]),.dout(n9955),.clk(gclk));
	jxor g09718(.dina(w_n9468_0[0]),.dinb(w_n3955_36[2]),.dout(n9956),.clk(gclk));
	jor g09719(.dina(n9956),.dinb(w_n9832_44[0]),.dout(n9957),.clk(gclk));
	jxor g09720(.dina(n9957),.dinb(w_n9474_0[0]),.dout(n9958),.clk(gclk));
	jor g09721(.dina(w_n9958_0[2]),.dinb(n9955),.dout(n9959),.clk(gclk));
	jand g09722(.dina(n9959),.dinb(w_n9954_0[1]),.dout(n9960),.clk(gclk));
	jor g09723(.dina(w_n9960_0[2]),.dinb(w_n3368_38[0]),.dout(n9961),.clk(gclk));
	jand g09724(.dina(w_n9960_0[1]),.dinb(w_n3368_37[2]),.dout(n9962),.clk(gclk));
	jxor g09725(.dina(w_n9476_0[0]),.dinb(w_n3642_40[0]),.dout(n9963),.clk(gclk));
	jor g09726(.dina(n9963),.dinb(w_n9832_43[2]),.dout(n9964),.clk(gclk));
	jxor g09727(.dina(n9964),.dinb(w_n9739_0[0]),.dout(n9965),.clk(gclk));
	jnot g09728(.din(w_n9965_0[2]),.dout(n9966),.clk(gclk));
	jor g09729(.dina(n9966),.dinb(n9962),.dout(n9967),.clk(gclk));
	jand g09730(.dina(n9967),.dinb(w_n9961_0[1]),.dout(n9968),.clk(gclk));
	jor g09731(.dina(w_n9968_0[2]),.dinb(w_n3089_41[1]),.dout(n9969),.clk(gclk));
	jand g09732(.dina(w_n9968_0[1]),.dinb(w_n3089_41[0]),.dout(n9970),.clk(gclk));
	jxor g09733(.dina(w_n9483_0[0]),.dinb(w_n3368_37[1]),.dout(n9971),.clk(gclk));
	jor g09734(.dina(n9971),.dinb(w_n9832_43[1]),.dout(n9972),.clk(gclk));
	jxor g09735(.dina(n9972),.dinb(w_n9488_0[0]),.dout(n9973),.clk(gclk));
	jor g09736(.dina(w_n9973_0[2]),.dinb(n9970),.dout(n9974),.clk(gclk));
	jand g09737(.dina(n9974),.dinb(w_n9969_0[1]),.dout(n9975),.clk(gclk));
	jor g09738(.dina(w_n9975_0[2]),.dinb(w_n2833_39[0]),.dout(n9976),.clk(gclk));
	jand g09739(.dina(w_n9975_0[1]),.dinb(w_n2833_38[2]),.dout(n9977),.clk(gclk));
	jxor g09740(.dina(w_n9490_0[0]),.dinb(w_n3089_40[2]),.dout(n9978),.clk(gclk));
	jor g09741(.dina(n9978),.dinb(w_n9832_43[0]),.dout(n9979),.clk(gclk));
	jxor g09742(.dina(n9979),.dinb(w_n9496_0[0]),.dout(n9980),.clk(gclk));
	jor g09743(.dina(w_n9980_0[2]),.dinb(n9977),.dout(n9981),.clk(gclk));
	jand g09744(.dina(n9981),.dinb(w_n9976_0[1]),.dout(n9982),.clk(gclk));
	jor g09745(.dina(w_n9982_0[2]),.dinb(w_n2572_41[2]),.dout(n9983),.clk(gclk));
	jand g09746(.dina(w_n9982_0[1]),.dinb(w_n2572_41[1]),.dout(n9984),.clk(gclk));
	jxor g09747(.dina(w_n9498_0[0]),.dinb(w_n2833_38[1]),.dout(n9985),.clk(gclk));
	jor g09748(.dina(n9985),.dinb(w_n9832_42[2]),.dout(n9986),.clk(gclk));
	jxor g09749(.dina(n9986),.dinb(w_n9504_0[0]),.dout(n9987),.clk(gclk));
	jor g09750(.dina(w_n9987_0[2]),.dinb(n9984),.dout(n9988),.clk(gclk));
	jand g09751(.dina(n9988),.dinb(w_n9983_0[1]),.dout(n9989),.clk(gclk));
	jor g09752(.dina(w_n9989_0[2]),.dinb(w_n2345_39[2]),.dout(n9990),.clk(gclk));
	jand g09753(.dina(w_n9989_0[1]),.dinb(w_n2345_39[1]),.dout(n9991),.clk(gclk));
	jxor g09754(.dina(w_n9506_0[0]),.dinb(w_n2572_41[0]),.dout(n9992),.clk(gclk));
	jor g09755(.dina(n9992),.dinb(w_n9832_42[1]),.dout(n9993),.clk(gclk));
	jxor g09756(.dina(n9993),.dinb(w_n9753_0[0]),.dout(n9994),.clk(gclk));
	jnot g09757(.din(w_n9994_0[2]),.dout(n9995),.clk(gclk));
	jor g09758(.dina(n9995),.dinb(n9991),.dout(n9996),.clk(gclk));
	jand g09759(.dina(n9996),.dinb(w_n9990_0[1]),.dout(n9997),.clk(gclk));
	jor g09760(.dina(w_n9997_0[2]),.dinb(w_n2108_42[1]),.dout(n9998),.clk(gclk));
	jand g09761(.dina(w_n9997_0[1]),.dinb(w_n2108_42[0]),.dout(n9999),.clk(gclk));
	jxor g09762(.dina(w_n9513_0[0]),.dinb(w_n2345_39[0]),.dout(n10000),.clk(gclk));
	jor g09763(.dina(n10000),.dinb(w_n9832_42[0]),.dout(n10001),.clk(gclk));
	jxor g09764(.dina(n10001),.dinb(w_n9519_0[0]),.dout(n10002),.clk(gclk));
	jor g09765(.dina(w_n10002_0[2]),.dinb(n9999),.dout(n10003),.clk(gclk));
	jand g09766(.dina(n10003),.dinb(w_n9998_0[1]),.dout(n10004),.clk(gclk));
	jor g09767(.dina(w_n10004_0[2]),.dinb(w_n1912_40[2]),.dout(n10005),.clk(gclk));
	jand g09768(.dina(w_n10004_0[1]),.dinb(w_n1912_40[1]),.dout(n10006),.clk(gclk));
	jxor g09769(.dina(w_n9521_0[0]),.dinb(w_n2108_41[2]),.dout(n10007),.clk(gclk));
	jor g09770(.dina(n10007),.dinb(w_n9832_41[2]),.dout(n10008),.clk(gclk));
	jxor g09771(.dina(n10008),.dinb(w_n9760_0[0]),.dout(n10009),.clk(gclk));
	jnot g09772(.din(w_n10009_0[2]),.dout(n10010),.clk(gclk));
	jor g09773(.dina(n10010),.dinb(n10006),.dout(n10011),.clk(gclk));
	jand g09774(.dina(n10011),.dinb(w_n10005_0[1]),.dout(n10012),.clk(gclk));
	jor g09775(.dina(w_n10012_0[2]),.dinb(w_n1699_43[0]),.dout(n10013),.clk(gclk));
	jand g09776(.dina(w_n10012_0[1]),.dinb(w_n1699_42[2]),.dout(n10014),.clk(gclk));
	jxor g09777(.dina(w_n9528_0[0]),.dinb(w_n1912_40[0]),.dout(n10015),.clk(gclk));
	jor g09778(.dina(n10015),.dinb(w_n9832_41[1]),.dout(n10016),.clk(gclk));
	jxor g09779(.dina(n10016),.dinb(w_n9534_0[0]),.dout(n10017),.clk(gclk));
	jor g09780(.dina(w_n10017_0[2]),.dinb(n10014),.dout(n10018),.clk(gclk));
	jand g09781(.dina(n10018),.dinb(w_n10013_0[1]),.dout(n10019),.clk(gclk));
	jor g09782(.dina(w_n10019_0[2]),.dinb(w_n1516_41[1]),.dout(n10020),.clk(gclk));
	jand g09783(.dina(w_n10019_0[1]),.dinb(w_n1516_41[0]),.dout(n10021),.clk(gclk));
	jxor g09784(.dina(w_n9536_0[0]),.dinb(w_n1699_42[1]),.dout(n10022),.clk(gclk));
	jor g09785(.dina(n10022),.dinb(w_n9832_41[0]),.dout(n10023),.clk(gclk));
	jxor g09786(.dina(n10023),.dinb(w_n9767_0[0]),.dout(n10024),.clk(gclk));
	jnot g09787(.din(w_n10024_0[2]),.dout(n10025),.clk(gclk));
	jor g09788(.dina(n10025),.dinb(n10021),.dout(n10026),.clk(gclk));
	jand g09789(.dina(n10026),.dinb(w_n10020_0[1]),.dout(n10027),.clk(gclk));
	jor g09790(.dina(w_n10027_0[2]),.dinb(w_n1332_43[0]),.dout(n10028),.clk(gclk));
	jand g09791(.dina(w_n10027_0[1]),.dinb(w_n1332_42[2]),.dout(n10029),.clk(gclk));
	jxor g09792(.dina(w_n9543_0[0]),.dinb(w_n1516_40[2]),.dout(n10030),.clk(gclk));
	jor g09793(.dina(n10030),.dinb(w_n9832_40[2]),.dout(n10031),.clk(gclk));
	jxor g09794(.dina(n10031),.dinb(w_n9549_0[0]),.dout(n10032),.clk(gclk));
	jor g09795(.dina(w_n10032_0[2]),.dinb(n10029),.dout(n10033),.clk(gclk));
	jand g09796(.dina(n10033),.dinb(w_n10028_0[1]),.dout(n10034),.clk(gclk));
	jor g09797(.dina(w_n10034_0[2]),.dinb(w_n1173_42[0]),.dout(n10035),.clk(gclk));
	jand g09798(.dina(w_n10034_0[1]),.dinb(w_n1173_41[2]),.dout(n10036),.clk(gclk));
	jxor g09799(.dina(w_n9551_0[0]),.dinb(w_n1332_42[1]),.dout(n10037),.clk(gclk));
	jor g09800(.dina(n10037),.dinb(w_n9832_40[1]),.dout(n10038),.clk(gclk));
	jxor g09801(.dina(n10038),.dinb(w_n9774_0[0]),.dout(n10039),.clk(gclk));
	jnot g09802(.din(w_n10039_0[2]),.dout(n10040),.clk(gclk));
	jor g09803(.dina(n10040),.dinb(n10036),.dout(n10041),.clk(gclk));
	jand g09804(.dina(n10041),.dinb(w_n10035_0[1]),.dout(n10042),.clk(gclk));
	jor g09805(.dina(w_n10042_0[2]),.dinb(w_n1008_44[0]),.dout(n10043),.clk(gclk));
	jand g09806(.dina(w_n10042_0[1]),.dinb(w_n1008_43[2]),.dout(n10044),.clk(gclk));
	jxor g09807(.dina(w_n9558_0[0]),.dinb(w_n1173_41[1]),.dout(n10045),.clk(gclk));
	jor g09808(.dina(n10045),.dinb(w_n9832_40[0]),.dout(n10046),.clk(gclk));
	jxor g09809(.dina(n10046),.dinb(w_n9778_0[0]),.dout(n10047),.clk(gclk));
	jnot g09810(.din(w_n10047_0[2]),.dout(n10048),.clk(gclk));
	jor g09811(.dina(n10048),.dinb(n10044),.dout(n10049),.clk(gclk));
	jand g09812(.dina(n10049),.dinb(w_n10043_0[1]),.dout(n10050),.clk(gclk));
	jor g09813(.dina(w_n10050_0[2]),.dinb(w_n884_43[0]),.dout(n10051),.clk(gclk));
	jand g09814(.dina(w_n10050_0[1]),.dinb(w_n884_42[2]),.dout(n10052),.clk(gclk));
	jxor g09815(.dina(w_n9565_0[0]),.dinb(w_n1008_43[1]),.dout(n10053),.clk(gclk));
	jor g09816(.dina(n10053),.dinb(w_n9832_39[2]),.dout(n10054),.clk(gclk));
	jxor g09817(.dina(n10054),.dinb(w_n9782_0[0]),.dout(n10055),.clk(gclk));
	jnot g09818(.din(w_n10055_0[2]),.dout(n10056),.clk(gclk));
	jor g09819(.dina(n10056),.dinb(n10052),.dout(n10057),.clk(gclk));
	jand g09820(.dina(n10057),.dinb(w_n10051_0[1]),.dout(n10058),.clk(gclk));
	jor g09821(.dina(w_n10058_0[2]),.dinb(w_n743_44[0]),.dout(n10059),.clk(gclk));
	jand g09822(.dina(w_n10058_0[1]),.dinb(w_n743_43[2]),.dout(n10060),.clk(gclk));
	jxor g09823(.dina(w_n9572_0[0]),.dinb(w_n884_42[1]),.dout(n10061),.clk(gclk));
	jor g09824(.dina(n10061),.dinb(w_n9832_39[1]),.dout(n10062),.clk(gclk));
	jxor g09825(.dina(n10062),.dinb(w_n9578_0[0]),.dout(n10063),.clk(gclk));
	jor g09826(.dina(w_n10063_0[2]),.dinb(n10060),.dout(n10064),.clk(gclk));
	jand g09827(.dina(n10064),.dinb(w_n10059_0[1]),.dout(n10065),.clk(gclk));
	jor g09828(.dina(w_n10065_0[2]),.dinb(w_n635_44[0]),.dout(n10066),.clk(gclk));
	jand g09829(.dina(w_n10065_0[1]),.dinb(w_n635_43[2]),.dout(n10067),.clk(gclk));
	jxor g09830(.dina(w_n9580_0[0]),.dinb(w_n743_43[1]),.dout(n10068),.clk(gclk));
	jor g09831(.dina(n10068),.dinb(w_n9832_39[0]),.dout(n10069),.clk(gclk));
	jxor g09832(.dina(n10069),.dinb(w_n9586_0[0]),.dout(n10070),.clk(gclk));
	jor g09833(.dina(w_n10070_0[2]),.dinb(n10067),.dout(n10071),.clk(gclk));
	jand g09834(.dina(n10071),.dinb(w_n10066_0[1]),.dout(n10072),.clk(gclk));
	jor g09835(.dina(w_n10072_0[2]),.dinb(w_n515_45[0]),.dout(n10073),.clk(gclk));
	jand g09836(.dina(w_n10072_0[1]),.dinb(w_n515_44[2]),.dout(n10074),.clk(gclk));
	jxor g09837(.dina(w_n9588_0[0]),.dinb(w_n635_43[1]),.dout(n10075),.clk(gclk));
	jor g09838(.dina(n10075),.dinb(w_n9832_38[2]),.dout(n10076),.clk(gclk));
	jxor g09839(.dina(n10076),.dinb(w_n9594_0[0]),.dout(n10077),.clk(gclk));
	jor g09840(.dina(w_n10077_0[2]),.dinb(n10074),.dout(n10078),.clk(gclk));
	jand g09841(.dina(n10078),.dinb(w_n10073_0[1]),.dout(n10079),.clk(gclk));
	jor g09842(.dina(w_n10079_0[2]),.dinb(w_n443_45[0]),.dout(n10080),.clk(gclk));
	jand g09843(.dina(w_n10079_0[1]),.dinb(w_n443_44[2]),.dout(n10081),.clk(gclk));
	jxor g09844(.dina(w_n9596_0[0]),.dinb(w_n515_44[1]),.dout(n10082),.clk(gclk));
	jor g09845(.dina(n10082),.dinb(w_n9832_38[1]),.dout(n10083),.clk(gclk));
	jxor g09846(.dina(n10083),.dinb(w_n9795_0[0]),.dout(n10084),.clk(gclk));
	jnot g09847(.din(w_n10084_0[2]),.dout(n10085),.clk(gclk));
	jor g09848(.dina(n10085),.dinb(n10081),.dout(n10086),.clk(gclk));
	jand g09849(.dina(n10086),.dinb(w_n10080_0[1]),.dout(n10087),.clk(gclk));
	jor g09850(.dina(w_n10087_0[2]),.dinb(w_n352_45[1]),.dout(n10088),.clk(gclk));
	jand g09851(.dina(w_n10087_0[1]),.dinb(w_n352_45[0]),.dout(n10089),.clk(gclk));
	jxor g09852(.dina(w_n9603_0[0]),.dinb(w_n443_44[1]),.dout(n10090),.clk(gclk));
	jor g09853(.dina(n10090),.dinb(w_n9832_38[0]),.dout(n10091),.clk(gclk));
	jxor g09854(.dina(n10091),.dinb(w_n9609_0[0]),.dout(n10092),.clk(gclk));
	jor g09855(.dina(w_n10092_0[2]),.dinb(n10089),.dout(n10093),.clk(gclk));
	jand g09856(.dina(n10093),.dinb(w_n10088_0[1]),.dout(n10094),.clk(gclk));
	jor g09857(.dina(w_n10094_0[2]),.dinb(w_n294_45[2]),.dout(n10095),.clk(gclk));
	jand g09858(.dina(w_n10094_0[1]),.dinb(w_n294_45[1]),.dout(n10096),.clk(gclk));
	jxor g09859(.dina(w_n9611_0[0]),.dinb(w_n352_44[2]),.dout(n10097),.clk(gclk));
	jor g09860(.dina(n10097),.dinb(w_n9832_37[2]),.dout(n10098),.clk(gclk));
	jxor g09861(.dina(n10098),.dinb(w_n9617_0[0]),.dout(n10099),.clk(gclk));
	jor g09862(.dina(w_n10099_0[2]),.dinb(n10096),.dout(n10100),.clk(gclk));
	jand g09863(.dina(n10100),.dinb(w_n10095_0[1]),.dout(n10101),.clk(gclk));
	jor g09864(.dina(w_n10101_0[2]),.dinb(w_n239_45[2]),.dout(n10102),.clk(gclk));
	jand g09865(.dina(w_n10101_0[1]),.dinb(w_n239_45[1]),.dout(n10103),.clk(gclk));
	jxor g09866(.dina(w_n9619_0[0]),.dinb(w_n294_45[0]),.dout(n10104),.clk(gclk));
	jor g09867(.dina(n10104),.dinb(w_n9832_37[1]),.dout(n10105),.clk(gclk));
	jxor g09868(.dina(n10105),.dinb(w_n9625_0[0]),.dout(n10106),.clk(gclk));
	jor g09869(.dina(w_n10106_0[2]),.dinb(n10103),.dout(n10107),.clk(gclk));
	jand g09870(.dina(n10107),.dinb(w_n10102_0[1]),.dout(n10108),.clk(gclk));
	jor g09871(.dina(w_n10108_0[2]),.dinb(w_n221_46[0]),.dout(n10109),.clk(gclk));
	jand g09872(.dina(w_n10108_0[1]),.dinb(w_n221_45[2]),.dout(n10110),.clk(gclk));
	jxor g09873(.dina(w_n9627_0[0]),.dinb(w_n239_45[0]),.dout(n10111),.clk(gclk));
	jor g09874(.dina(n10111),.dinb(w_n9832_37[0]),.dout(n10112),.clk(gclk));
	jxor g09875(.dina(n10112),.dinb(w_n9808_0[0]),.dout(n10113),.clk(gclk));
	jnot g09876(.din(w_n10113_0[1]),.dout(n10114),.clk(gclk));
	jor g09877(.dina(w_n10114_0[1]),.dinb(n10110),.dout(n10115),.clk(gclk));
	jand g09878(.dina(n10115),.dinb(w_n10109_0[1]),.dout(n10116),.clk(gclk));
	jxor g09879(.dina(w_n9634_0[0]),.dinb(w_n221_45[1]),.dout(n10117),.clk(gclk));
	jor g09880(.dina(n10117),.dinb(w_n9832_36[2]),.dout(n10118),.clk(gclk));
	jxor g09881(.dina(n10118),.dinb(w_n9639_0[0]),.dout(n10119),.clk(gclk));
	jor g09882(.dina(w_n10119_1[1]),.dinb(w_n10116_0[2]),.dout(n10120),.clk(gclk));
	jor g09883(.dina(w_n10120_0[1]),.dinb(w_n9643_0[0]),.dout(n10121),.clk(gclk));
	jor g09884(.dina(n10121),.dinb(w_n9825_0[1]),.dout(n10122),.clk(gclk));
	jand g09885(.dina(n10122),.dinb(w_n218_19[0]),.dout(n10123),.clk(gclk));
	jand g09886(.dina(w_n9832_36[1]),.dinb(w_n9649_0[0]),.dout(n10124),.clk(gclk));
	jand g09887(.dina(w_n10119_1[0]),.dinb(w_n10116_0[1]),.dout(n10125),.clk(gclk));
	jor g09888(.dina(w_n10125_1[1]),.dinb(n10124),.dout(n10126),.clk(gclk));
	jand g09889(.dina(w_n9831_0[0]),.dinb(w_n9814_0[0]),.dout(n10127),.clk(gclk));
	jnot g09890(.din(n10127),.dout(n10128),.clk(gclk));
	jand g09891(.dina(w_n9815_0[0]),.dinb(w_asqrt63_34[0]),.dout(n10129),.clk(gclk));
	jand g09892(.dina(n10129),.dinb(w_n9642_0[2]),.dout(n10130),.clk(gclk));
	jand g09893(.dina(w_n10130_0[1]),.dinb(n10128),.dout(n10131),.clk(gclk));
	jor g09894(.dina(n10131),.dinb(n10126),.dout(n10132),.clk(gclk));
	jor g09895(.dina(w_n10132_0[1]),.dinb(w_n10123_0[1]),.dout(asqrt_fa_25),.clk(gclk));
	jnot g09896(.din(w_a46_1[1]),.dout(n10134),.clk(gclk));
	jnot g09897(.din(w_a47_0[1]),.dout(n10135),.clk(gclk));
	jand g09898(.dina(w_n10135_0[1]),.dinb(w_n10134_1[1]),.dout(n10136),.clk(gclk));
	jand g09899(.dina(w_n10136_0[2]),.dinb(w_n9834_1[1]),.dout(n10137),.clk(gclk));
	jand g09900(.dina(w_asqrt24_36[1]),.dinb(w_a48_0[1]),.dout(n10138),.clk(gclk));
	jor g09901(.dina(n10138),.dinb(w_n10137_0[1]),.dout(n10139),.clk(gclk));
	jand g09902(.dina(w_n10139_0[2]),.dinb(w_asqrt25_18[0]),.dout(n10140),.clk(gclk));
	jor g09903(.dina(w_n10139_0[1]),.dinb(w_asqrt25_17[2]),.dout(n10141),.clk(gclk));
	jand g09904(.dina(w_asqrt24_36[0]),.dinb(w_n9834_1[0]),.dout(n10142),.clk(gclk));
	jor g09905(.dina(n10142),.dinb(w_n9835_0[0]),.dout(n10143),.clk(gclk));
	jnot g09906(.din(w_n9836_0[1]),.dout(n10144),.clk(gclk));
	jnot g09907(.din(w_n9825_0[0]),.dout(n10145),.clk(gclk));
	jnot g09908(.din(w_n10109_0[0]),.dout(n10146),.clk(gclk));
	jnot g09909(.din(w_n10102_0[0]),.dout(n10147),.clk(gclk));
	jnot g09910(.din(w_n10095_0[0]),.dout(n10148),.clk(gclk));
	jnot g09911(.din(w_n10088_0[0]),.dout(n10149),.clk(gclk));
	jnot g09912(.din(w_n10080_0[0]),.dout(n10150),.clk(gclk));
	jnot g09913(.din(w_n10073_0[0]),.dout(n10151),.clk(gclk));
	jnot g09914(.din(w_n10066_0[0]),.dout(n10152),.clk(gclk));
	jnot g09915(.din(w_n10059_0[0]),.dout(n10153),.clk(gclk));
	jnot g09916(.din(w_n10051_0[0]),.dout(n10154),.clk(gclk));
	jnot g09917(.din(w_n10043_0[0]),.dout(n10155),.clk(gclk));
	jnot g09918(.din(w_n10035_0[0]),.dout(n10156),.clk(gclk));
	jnot g09919(.din(w_n10028_0[0]),.dout(n10157),.clk(gclk));
	jnot g09920(.din(w_n10020_0[0]),.dout(n10158),.clk(gclk));
	jnot g09921(.din(w_n10013_0[0]),.dout(n10159),.clk(gclk));
	jnot g09922(.din(w_n10005_0[0]),.dout(n10160),.clk(gclk));
	jnot g09923(.din(w_n9998_0[0]),.dout(n10161),.clk(gclk));
	jnot g09924(.din(w_n9990_0[0]),.dout(n10162),.clk(gclk));
	jnot g09925(.din(w_n9983_0[0]),.dout(n10163),.clk(gclk));
	jnot g09926(.din(w_n9976_0[0]),.dout(n10164),.clk(gclk));
	jnot g09927(.din(w_n9969_0[0]),.dout(n10165),.clk(gclk));
	jnot g09928(.din(w_n9961_0[0]),.dout(n10166),.clk(gclk));
	jnot g09929(.din(w_n9954_0[0]),.dout(n10167),.clk(gclk));
	jnot g09930(.din(w_n9946_0[0]),.dout(n10168),.clk(gclk));
	jnot g09931(.din(w_n9939_0[0]),.dout(n10169),.clk(gclk));
	jnot g09932(.din(w_n9931_0[0]),.dout(n10170),.clk(gclk));
	jnot g09933(.din(w_n9924_0[0]),.dout(n10171),.clk(gclk));
	jnot g09934(.din(w_n9917_0[0]),.dout(n10172),.clk(gclk));
	jnot g09935(.din(w_n9910_0[0]),.dout(n10173),.clk(gclk));
	jnot g09936(.din(w_n9903_0[0]),.dout(n10174),.clk(gclk));
	jnot g09937(.din(w_n9896_0[0]),.dout(n10175),.clk(gclk));
	jnot g09938(.din(w_n9888_0[0]),.dout(n10176),.clk(gclk));
	jnot g09939(.din(w_n9881_0[0]),.dout(n10177),.clk(gclk));
	jnot g09940(.din(w_n9874_0[0]),.dout(n10178),.clk(gclk));
	jnot g09941(.din(w_n9867_0[0]),.dout(n10179),.clk(gclk));
	jnot g09942(.din(w_n9859_0[0]),.dout(n10180),.clk(gclk));
	jnot g09943(.din(w_n9848_0[0]),.dout(n10181),.clk(gclk));
	jnot g09944(.din(w_n9840_0[0]),.dout(n10182),.clk(gclk));
	jand g09945(.dina(w_asqrt25_17[1]),.dinb(w_a50_0[0]),.dout(n10183),.clk(gclk));
	jor g09946(.dina(w_n9837_0[0]),.dinb(n10183),.dout(n10184),.clk(gclk));
	jor g09947(.dina(n10184),.dinb(w_asqrt26_23[2]),.dout(n10185),.clk(gclk));
	jand g09948(.dina(w_asqrt25_17[0]),.dinb(w_n9188_0[2]),.dout(n10186),.clk(gclk));
	jor g09949(.dina(n10186),.dinb(w_n9189_0[0]),.dout(n10187),.clk(gclk));
	jand g09950(.dina(w_n9851_0[0]),.dinb(n10187),.dout(n10188),.clk(gclk));
	jand g09951(.dina(w_n10188_0[1]),.dinb(n10185),.dout(n10189),.clk(gclk));
	jor g09952(.dina(n10189),.dinb(n10182),.dout(n10190),.clk(gclk));
	jor g09953(.dina(n10190),.dinb(w_asqrt27_18[1]),.dout(n10191),.clk(gclk));
	jnot g09954(.din(w_n9856_0[1]),.dout(n10192),.clk(gclk));
	jand g09955(.dina(n10192),.dinb(n10191),.dout(n10193),.clk(gclk));
	jor g09956(.dina(n10193),.dinb(n10181),.dout(n10194),.clk(gclk));
	jor g09957(.dina(n10194),.dinb(w_asqrt28_24[0]),.dout(n10195),.clk(gclk));
	jand g09958(.dina(w_n9863_0[1]),.dinb(n10195),.dout(n10196),.clk(gclk));
	jor g09959(.dina(n10196),.dinb(n10180),.dout(n10197),.clk(gclk));
	jor g09960(.dina(n10197),.dinb(w_asqrt29_18[2]),.dout(n10198),.clk(gclk));
	jnot g09961(.din(w_n9871_0[1]),.dout(n10199),.clk(gclk));
	jand g09962(.dina(n10199),.dinb(n10198),.dout(n10200),.clk(gclk));
	jor g09963(.dina(n10200),.dinb(n10179),.dout(n10201),.clk(gclk));
	jor g09964(.dina(n10201),.dinb(w_asqrt30_24[1]),.dout(n10202),.clk(gclk));
	jnot g09965(.din(w_n9878_0[1]),.dout(n10203),.clk(gclk));
	jand g09966(.dina(n10203),.dinb(n10202),.dout(n10204),.clk(gclk));
	jor g09967(.dina(n10204),.dinb(n10178),.dout(n10205),.clk(gclk));
	jor g09968(.dina(n10205),.dinb(w_asqrt31_19[1]),.dout(n10206),.clk(gclk));
	jnot g09969(.din(w_n9885_0[1]),.dout(n10207),.clk(gclk));
	jand g09970(.dina(n10207),.dinb(n10206),.dout(n10208),.clk(gclk));
	jor g09971(.dina(n10208),.dinb(n10177),.dout(n10209),.clk(gclk));
	jor g09972(.dina(n10209),.dinb(w_asqrt32_24[1]),.dout(n10210),.clk(gclk));
	jand g09973(.dina(w_n9892_0[1]),.dinb(n10210),.dout(n10211),.clk(gclk));
	jor g09974(.dina(n10211),.dinb(n10176),.dout(n10212),.clk(gclk));
	jor g09975(.dina(n10212),.dinb(w_asqrt33_20[0]),.dout(n10213),.clk(gclk));
	jnot g09976(.din(w_n9900_0[1]),.dout(n10214),.clk(gclk));
	jand g09977(.dina(n10214),.dinb(n10213),.dout(n10215),.clk(gclk));
	jor g09978(.dina(n10215),.dinb(n10175),.dout(n10216),.clk(gclk));
	jor g09979(.dina(n10216),.dinb(w_asqrt34_24[2]),.dout(n10217),.clk(gclk));
	jnot g09980(.din(w_n9907_0[1]),.dout(n10218),.clk(gclk));
	jand g09981(.dina(n10218),.dinb(n10217),.dout(n10219),.clk(gclk));
	jor g09982(.dina(n10219),.dinb(n10174),.dout(n10220),.clk(gclk));
	jor g09983(.dina(n10220),.dinb(w_asqrt35_20[2]),.dout(n10221),.clk(gclk));
	jnot g09984(.din(w_n9914_0[1]),.dout(n10222),.clk(gclk));
	jand g09985(.dina(n10222),.dinb(n10221),.dout(n10223),.clk(gclk));
	jor g09986(.dina(n10223),.dinb(n10173),.dout(n10224),.clk(gclk));
	jor g09987(.dina(n10224),.dinb(w_asqrt36_24[2]),.dout(n10225),.clk(gclk));
	jnot g09988(.din(w_n9921_0[1]),.dout(n10226),.clk(gclk));
	jand g09989(.dina(n10226),.dinb(n10225),.dout(n10227),.clk(gclk));
	jor g09990(.dina(n10227),.dinb(n10172),.dout(n10228),.clk(gclk));
	jor g09991(.dina(n10228),.dinb(w_asqrt37_21[0]),.dout(n10229),.clk(gclk));
	jnot g09992(.din(w_n9928_0[1]),.dout(n10230),.clk(gclk));
	jand g09993(.dina(n10230),.dinb(n10229),.dout(n10231),.clk(gclk));
	jor g09994(.dina(n10231),.dinb(n10171),.dout(n10232),.clk(gclk));
	jor g09995(.dina(n10232),.dinb(w_asqrt38_25[0]),.dout(n10233),.clk(gclk));
	jand g09996(.dina(n10233),.dinb(w_n9934_0[1]),.dout(n10234),.clk(gclk));
	jor g09997(.dina(n10234),.dinb(n10170),.dout(n10235),.clk(gclk));
	jor g09998(.dina(n10235),.dinb(w_asqrt39_21[2]),.dout(n10236),.clk(gclk));
	jnot g09999(.din(w_n9943_0[1]),.dout(n10237),.clk(gclk));
	jand g10000(.dina(n10237),.dinb(n10236),.dout(n10238),.clk(gclk));
	jor g10001(.dina(n10238),.dinb(n10169),.dout(n10239),.clk(gclk));
	jor g10002(.dina(n10239),.dinb(w_asqrt40_25[0]),.dout(n10240),.clk(gclk));
	jand g10003(.dina(w_n9950_0[1]),.dinb(n10240),.dout(n10241),.clk(gclk));
	jor g10004(.dina(n10241),.dinb(n10168),.dout(n10242),.clk(gclk));
	jor g10005(.dina(n10242),.dinb(w_asqrt41_22[0]),.dout(n10243),.clk(gclk));
	jnot g10006(.din(w_n9958_0[1]),.dout(n10244),.clk(gclk));
	jand g10007(.dina(n10244),.dinb(n10243),.dout(n10245),.clk(gclk));
	jor g10008(.dina(n10245),.dinb(n10167),.dout(n10246),.clk(gclk));
	jor g10009(.dina(n10246),.dinb(w_asqrt42_25[1]),.dout(n10247),.clk(gclk));
	jand g10010(.dina(w_n9965_0[1]),.dinb(n10247),.dout(n10248),.clk(gclk));
	jor g10011(.dina(n10248),.dinb(n10166),.dout(n10249),.clk(gclk));
	jor g10012(.dina(n10249),.dinb(w_asqrt43_22[1]),.dout(n10250),.clk(gclk));
	jnot g10013(.din(w_n9973_0[1]),.dout(n10251),.clk(gclk));
	jand g10014(.dina(n10251),.dinb(n10250),.dout(n10252),.clk(gclk));
	jor g10015(.dina(n10252),.dinb(n10165),.dout(n10253),.clk(gclk));
	jor g10016(.dina(n10253),.dinb(w_asqrt44_25[1]),.dout(n10254),.clk(gclk));
	jnot g10017(.din(w_n9980_0[1]),.dout(n10255),.clk(gclk));
	jand g10018(.dina(n10255),.dinb(n10254),.dout(n10256),.clk(gclk));
	jor g10019(.dina(n10256),.dinb(n10164),.dout(n10257),.clk(gclk));
	jor g10020(.dina(n10257),.dinb(w_asqrt45_23[0]),.dout(n10258),.clk(gclk));
	jnot g10021(.din(w_n9987_0[1]),.dout(n10259),.clk(gclk));
	jand g10022(.dina(n10259),.dinb(n10258),.dout(n10260),.clk(gclk));
	jor g10023(.dina(n10260),.dinb(n10163),.dout(n10261),.clk(gclk));
	jor g10024(.dina(n10261),.dinb(w_asqrt46_25[1]),.dout(n10262),.clk(gclk));
	jand g10025(.dina(w_n9994_0[1]),.dinb(n10262),.dout(n10263),.clk(gclk));
	jor g10026(.dina(n10263),.dinb(n10162),.dout(n10264),.clk(gclk));
	jor g10027(.dina(n10264),.dinb(w_asqrt47_23[2]),.dout(n10265),.clk(gclk));
	jnot g10028(.din(w_n10002_0[1]),.dout(n10266),.clk(gclk));
	jand g10029(.dina(n10266),.dinb(n10265),.dout(n10267),.clk(gclk));
	jor g10030(.dina(n10267),.dinb(n10161),.dout(n10268),.clk(gclk));
	jor g10031(.dina(n10268),.dinb(w_asqrt48_25[2]),.dout(n10269),.clk(gclk));
	jand g10032(.dina(w_n10009_0[1]),.dinb(n10269),.dout(n10270),.clk(gclk));
	jor g10033(.dina(n10270),.dinb(n10160),.dout(n10271),.clk(gclk));
	jor g10034(.dina(n10271),.dinb(w_asqrt49_24[0]),.dout(n10272),.clk(gclk));
	jnot g10035(.din(w_n10017_0[1]),.dout(n10273),.clk(gclk));
	jand g10036(.dina(n10273),.dinb(n10272),.dout(n10274),.clk(gclk));
	jor g10037(.dina(n10274),.dinb(n10159),.dout(n10275),.clk(gclk));
	jor g10038(.dina(n10275),.dinb(w_asqrt50_26[0]),.dout(n10276),.clk(gclk));
	jand g10039(.dina(w_n10024_0[1]),.dinb(n10276),.dout(n10277),.clk(gclk));
	jor g10040(.dina(n10277),.dinb(n10158),.dout(n10278),.clk(gclk));
	jor g10041(.dina(n10278),.dinb(w_asqrt51_24[1]),.dout(n10279),.clk(gclk));
	jnot g10042(.din(w_n10032_0[1]),.dout(n10280),.clk(gclk));
	jand g10043(.dina(n10280),.dinb(n10279),.dout(n10281),.clk(gclk));
	jor g10044(.dina(n10281),.dinb(n10157),.dout(n10282),.clk(gclk));
	jor g10045(.dina(n10282),.dinb(w_asqrt52_26[0]),.dout(n10283),.clk(gclk));
	jand g10046(.dina(w_n10039_0[1]),.dinb(n10283),.dout(n10284),.clk(gclk));
	jor g10047(.dina(n10284),.dinb(n10156),.dout(n10285),.clk(gclk));
	jor g10048(.dina(n10285),.dinb(w_asqrt53_25[0]),.dout(n10286),.clk(gclk));
	jand g10049(.dina(w_n10047_0[1]),.dinb(n10286),.dout(n10287),.clk(gclk));
	jor g10050(.dina(n10287),.dinb(n10155),.dout(n10288),.clk(gclk));
	jor g10051(.dina(n10288),.dinb(w_asqrt54_26[0]),.dout(n10289),.clk(gclk));
	jand g10052(.dina(w_n10055_0[1]),.dinb(n10289),.dout(n10290),.clk(gclk));
	jor g10053(.dina(n10290),.dinb(n10154),.dout(n10291),.clk(gclk));
	jor g10054(.dina(n10291),.dinb(w_asqrt55_25[1]),.dout(n10292),.clk(gclk));
	jnot g10055(.din(w_n10063_0[1]),.dout(n10293),.clk(gclk));
	jand g10056(.dina(n10293),.dinb(n10292),.dout(n10294),.clk(gclk));
	jor g10057(.dina(n10294),.dinb(n10153),.dout(n10295),.clk(gclk));
	jor g10058(.dina(n10295),.dinb(w_asqrt56_26[1]),.dout(n10296),.clk(gclk));
	jnot g10059(.din(w_n10070_0[1]),.dout(n10297),.clk(gclk));
	jand g10060(.dina(n10297),.dinb(n10296),.dout(n10298),.clk(gclk));
	jor g10061(.dina(n10298),.dinb(n10152),.dout(n10299),.clk(gclk));
	jor g10062(.dina(n10299),.dinb(w_asqrt57_26[0]),.dout(n10300),.clk(gclk));
	jnot g10063(.din(w_n10077_0[1]),.dout(n10301),.clk(gclk));
	jand g10064(.dina(n10301),.dinb(n10300),.dout(n10302),.clk(gclk));
	jor g10065(.dina(n10302),.dinb(n10151),.dout(n10303),.clk(gclk));
	jor g10066(.dina(n10303),.dinb(w_asqrt58_26[2]),.dout(n10304),.clk(gclk));
	jand g10067(.dina(w_n10084_0[1]),.dinb(n10304),.dout(n10305),.clk(gclk));
	jor g10068(.dina(n10305),.dinb(n10150),.dout(n10306),.clk(gclk));
	jor g10069(.dina(n10306),.dinb(w_asqrt59_26[1]),.dout(n10307),.clk(gclk));
	jnot g10070(.din(w_n10092_0[1]),.dout(n10308),.clk(gclk));
	jand g10071(.dina(n10308),.dinb(n10307),.dout(n10309),.clk(gclk));
	jor g10072(.dina(n10309),.dinb(n10149),.dout(n10310),.clk(gclk));
	jor g10073(.dina(n10310),.dinb(w_asqrt60_26[2]),.dout(n10311),.clk(gclk));
	jnot g10074(.din(w_n10099_0[1]),.dout(n10312),.clk(gclk));
	jand g10075(.dina(n10312),.dinb(n10311),.dout(n10313),.clk(gclk));
	jor g10076(.dina(n10313),.dinb(n10148),.dout(n10314),.clk(gclk));
	jor g10077(.dina(n10314),.dinb(w_asqrt61_26[2]),.dout(n10315),.clk(gclk));
	jnot g10078(.din(w_n10106_0[1]),.dout(n10316),.clk(gclk));
	jand g10079(.dina(n10316),.dinb(n10315),.dout(n10317),.clk(gclk));
	jor g10080(.dina(n10317),.dinb(n10147),.dout(n10318),.clk(gclk));
	jor g10081(.dina(n10318),.dinb(w_asqrt62_26[2]),.dout(n10319),.clk(gclk));
	jand g10082(.dina(w_n10113_0[0]),.dinb(n10319),.dout(n10320),.clk(gclk));
	jor g10083(.dina(n10320),.dinb(n10146),.dout(n10321),.clk(gclk));
	jnot g10084(.din(w_n10119_0[2]),.dout(n10322),.clk(gclk));
	jand g10085(.dina(n10322),.dinb(n10321),.dout(n10323),.clk(gclk));
	jand g10086(.dina(w_n10323_0[1]),.dinb(w_n9642_0[1]),.dout(n10324),.clk(gclk));
	jand g10087(.dina(n10324),.dinb(n10145),.dout(n10325),.clk(gclk));
	jor g10088(.dina(n10325),.dinb(w_asqrt63_33[2]),.dout(n10326),.clk(gclk));
	jnot g10089(.din(w_n10132_0[0]),.dout(n10327),.clk(gclk));
	jand g10090(.dina(n10327),.dinb(n10326),.dout(n10328),.clk(gclk));
	jor g10091(.dina(w_n10328_30[2]),.dinb(n10144),.dout(n10329),.clk(gclk));
	jand g10092(.dina(w_n10329_0[1]),.dinb(n10143),.dout(n10330),.clk(gclk));
	jand g10093(.dina(w_n10330_0[1]),.dinb(n10141),.dout(n10331),.clk(gclk));
	jor g10094(.dina(n10331),.dinb(w_n10140_0[1]),.dout(n10332),.clk(gclk));
	jand g10095(.dina(w_n10332_0[2]),.dinb(w_asqrt26_23[1]),.dout(n10333),.clk(gclk));
	jor g10096(.dina(w_n10332_0[1]),.dinb(w_asqrt26_23[0]),.dout(n10334),.clk(gclk));
	jor g10097(.dina(w_n10130_0[0]),.dinb(w_n10125_1[0]),.dout(n10335),.clk(gclk));
	jor g10098(.dina(n10335),.dinb(w_n10123_0[0]),.dout(n10336),.clk(gclk));
	jor g10099(.dina(n10336),.dinb(w_n9832_36[0]),.dout(n10337),.clk(gclk));
	jand g10100(.dina(n10337),.dinb(w_n10329_0[0]),.dout(n10338),.clk(gclk));
	jxor g10101(.dina(n10338),.dinb(w_n9188_0[1]),.dout(n10339),.clk(gclk));
	jnot g10102(.din(w_n10339_0[1]),.dout(n10340),.clk(gclk));
	jand g10103(.dina(w_n10340_0[1]),.dinb(n10334),.dout(n10341),.clk(gclk));
	jor g10104(.dina(n10341),.dinb(w_n10333_0[1]),.dout(n10342),.clk(gclk));
	jand g10105(.dina(w_n10342_0[2]),.dinb(w_asqrt27_18[0]),.dout(n10343),.clk(gclk));
	jor g10106(.dina(w_n10342_0[1]),.dinb(w_asqrt27_17[2]),.dout(n10344),.clk(gclk));
	jxor g10107(.dina(w_n9839_0[0]),.dinb(w_n9369_30[2]),.dout(n10345),.clk(gclk));
	jand g10108(.dina(n10345),.dinb(w_asqrt24_35[2]),.dout(n10346),.clk(gclk));
	jxor g10109(.dina(n10346),.dinb(w_n10188_0[0]),.dout(n10347),.clk(gclk));
	jand g10110(.dina(w_n10347_0[1]),.dinb(n10344),.dout(n10348),.clk(gclk));
	jor g10111(.dina(n10348),.dinb(w_n10343_0[1]),.dout(n10349),.clk(gclk));
	jand g10112(.dina(w_n10349_0[2]),.dinb(w_asqrt28_23[2]),.dout(n10350),.clk(gclk));
	jor g10113(.dina(w_n10349_0[1]),.dinb(w_asqrt28_23[1]),.dout(n10351),.clk(gclk));
	jxor g10114(.dina(w_n9847_0[0]),.dinb(w_n8890_36[1]),.dout(n10352),.clk(gclk));
	jand g10115(.dina(n10352),.dinb(w_asqrt24_35[1]),.dout(n10353),.clk(gclk));
	jxor g10116(.dina(n10353),.dinb(w_n9856_0[0]),.dout(n10354),.clk(gclk));
	jnot g10117(.din(w_n10354_0[1]),.dout(n10355),.clk(gclk));
	jand g10118(.dina(w_n10355_0[1]),.dinb(n10351),.dout(n10356),.clk(gclk));
	jor g10119(.dina(n10356),.dinb(w_n10350_0[1]),.dout(n10357),.clk(gclk));
	jand g10120(.dina(w_n10357_0[2]),.dinb(w_asqrt29_18[1]),.dout(n10358),.clk(gclk));
	jor g10121(.dina(w_n10357_0[1]),.dinb(w_asqrt29_18[0]),.dout(n10359),.clk(gclk));
	jxor g10122(.dina(w_n9858_0[0]),.dinb(w_n8449_31[1]),.dout(n10360),.clk(gclk));
	jand g10123(.dina(n10360),.dinb(w_asqrt24_35[0]),.dout(n10361),.clk(gclk));
	jxor g10124(.dina(n10361),.dinb(w_n9863_0[0]),.dout(n10362),.clk(gclk));
	jand g10125(.dina(w_n10362_0[1]),.dinb(n10359),.dout(n10363),.clk(gclk));
	jor g10126(.dina(n10363),.dinb(w_n10358_0[1]),.dout(n10364),.clk(gclk));
	jand g10127(.dina(w_n10364_0[2]),.dinb(w_asqrt30_24[0]),.dout(n10365),.clk(gclk));
	jor g10128(.dina(w_n10364_0[1]),.dinb(w_asqrt30_23[2]),.dout(n10366),.clk(gclk));
	jxor g10129(.dina(w_n9866_0[0]),.dinb(w_n8003_37[0]),.dout(n10367),.clk(gclk));
	jand g10130(.dina(n10367),.dinb(w_asqrt24_34[2]),.dout(n10368),.clk(gclk));
	jxor g10131(.dina(n10368),.dinb(w_n9871_0[0]),.dout(n10369),.clk(gclk));
	jnot g10132(.din(w_n10369_0[1]),.dout(n10370),.clk(gclk));
	jand g10133(.dina(w_n10370_0[1]),.dinb(n10366),.dout(n10371),.clk(gclk));
	jor g10134(.dina(n10371),.dinb(w_n10365_0[1]),.dout(n10372),.clk(gclk));
	jand g10135(.dina(w_n10372_0[2]),.dinb(w_asqrt31_19[0]),.dout(n10373),.clk(gclk));
	jor g10136(.dina(w_n10372_0[1]),.dinb(w_asqrt31_18[2]),.dout(n10374),.clk(gclk));
	jxor g10137(.dina(w_n9873_0[0]),.dinb(w_n7581_32[1]),.dout(n10375),.clk(gclk));
	jand g10138(.dina(n10375),.dinb(w_asqrt24_34[1]),.dout(n10376),.clk(gclk));
	jxor g10139(.dina(n10376),.dinb(w_n9878_0[0]),.dout(n10377),.clk(gclk));
	jnot g10140(.din(w_n10377_0[1]),.dout(n10378),.clk(gclk));
	jand g10141(.dina(w_n10378_0[1]),.dinb(n10374),.dout(n10379),.clk(gclk));
	jor g10142(.dina(n10379),.dinb(w_n10373_0[1]),.dout(n10380),.clk(gclk));
	jand g10143(.dina(w_n10380_0[2]),.dinb(w_asqrt32_24[0]),.dout(n10381),.clk(gclk));
	jor g10144(.dina(w_n10380_0[1]),.dinb(w_asqrt32_23[2]),.dout(n10382),.clk(gclk));
	jxor g10145(.dina(w_n9880_0[0]),.dinb(w_n7154_37[1]),.dout(n10383),.clk(gclk));
	jand g10146(.dina(n10383),.dinb(w_asqrt24_34[0]),.dout(n10384),.clk(gclk));
	jxor g10147(.dina(n10384),.dinb(w_n9885_0[0]),.dout(n10385),.clk(gclk));
	jnot g10148(.din(w_n10385_0[1]),.dout(n10386),.clk(gclk));
	jand g10149(.dina(w_n10386_0[1]),.dinb(n10382),.dout(n10387),.clk(gclk));
	jor g10150(.dina(n10387),.dinb(w_n10381_0[1]),.dout(n10388),.clk(gclk));
	jand g10151(.dina(w_n10388_0[2]),.dinb(w_asqrt33_19[2]),.dout(n10389),.clk(gclk));
	jor g10152(.dina(w_n10388_0[1]),.dinb(w_asqrt33_19[1]),.dout(n10390),.clk(gclk));
	jxor g10153(.dina(w_n9887_0[0]),.dinb(w_n6758_33[0]),.dout(n10391),.clk(gclk));
	jand g10154(.dina(n10391),.dinb(w_asqrt24_33[2]),.dout(n10392),.clk(gclk));
	jxor g10155(.dina(n10392),.dinb(w_n9892_0[0]),.dout(n10393),.clk(gclk));
	jand g10156(.dina(w_n10393_0[1]),.dinb(n10390),.dout(n10394),.clk(gclk));
	jor g10157(.dina(n10394),.dinb(w_n10389_0[1]),.dout(n10395),.clk(gclk));
	jand g10158(.dina(w_n10395_0[2]),.dinb(w_asqrt34_24[1]),.dout(n10396),.clk(gclk));
	jor g10159(.dina(w_n10395_0[1]),.dinb(w_asqrt34_24[0]),.dout(n10397),.clk(gclk));
	jxor g10160(.dina(w_n9895_0[0]),.dinb(w_n6357_37[2]),.dout(n10398),.clk(gclk));
	jand g10161(.dina(n10398),.dinb(w_asqrt24_33[1]),.dout(n10399),.clk(gclk));
	jxor g10162(.dina(n10399),.dinb(w_n9900_0[0]),.dout(n10400),.clk(gclk));
	jnot g10163(.din(w_n10400_0[1]),.dout(n10401),.clk(gclk));
	jand g10164(.dina(w_n10401_0[1]),.dinb(n10397),.dout(n10402),.clk(gclk));
	jor g10165(.dina(n10402),.dinb(w_n10396_0[1]),.dout(n10403),.clk(gclk));
	jand g10166(.dina(w_n10403_0[2]),.dinb(w_asqrt35_20[1]),.dout(n10404),.clk(gclk));
	jor g10167(.dina(w_n10403_0[1]),.dinb(w_asqrt35_20[0]),.dout(n10405),.clk(gclk));
	jxor g10168(.dina(w_n9902_0[0]),.dinb(w_n5989_33[2]),.dout(n10406),.clk(gclk));
	jand g10169(.dina(n10406),.dinb(w_asqrt24_33[0]),.dout(n10407),.clk(gclk));
	jxor g10170(.dina(n10407),.dinb(w_n9907_0[0]),.dout(n10408),.clk(gclk));
	jnot g10171(.din(w_n10408_0[1]),.dout(n10409),.clk(gclk));
	jand g10172(.dina(w_n10409_0[1]),.dinb(n10405),.dout(n10410),.clk(gclk));
	jor g10173(.dina(n10410),.dinb(w_n10404_0[1]),.dout(n10411),.clk(gclk));
	jand g10174(.dina(w_n10411_0[2]),.dinb(w_asqrt36_24[1]),.dout(n10412),.clk(gclk));
	jor g10175(.dina(w_n10411_0[1]),.dinb(w_asqrt36_24[0]),.dout(n10413),.clk(gclk));
	jxor g10176(.dina(w_n9909_0[0]),.dinb(w_n5606_38[0]),.dout(n10414),.clk(gclk));
	jand g10177(.dina(n10414),.dinb(w_asqrt24_32[2]),.dout(n10415),.clk(gclk));
	jxor g10178(.dina(n10415),.dinb(w_n9914_0[0]),.dout(n10416),.clk(gclk));
	jnot g10179(.din(w_n10416_0[1]),.dout(n10417),.clk(gclk));
	jand g10180(.dina(w_n10417_0[1]),.dinb(n10413),.dout(n10418),.clk(gclk));
	jor g10181(.dina(n10418),.dinb(w_n10412_0[1]),.dout(n10419),.clk(gclk));
	jand g10182(.dina(w_n10419_0[2]),.dinb(w_asqrt37_20[2]),.dout(n10420),.clk(gclk));
	jor g10183(.dina(w_n10419_0[1]),.dinb(w_asqrt37_20[1]),.dout(n10421),.clk(gclk));
	jxor g10184(.dina(w_n9916_0[0]),.dinb(w_n5259_34[2]),.dout(n10422),.clk(gclk));
	jand g10185(.dina(n10422),.dinb(w_asqrt24_32[1]),.dout(n10423),.clk(gclk));
	jxor g10186(.dina(n10423),.dinb(w_n9921_0[0]),.dout(n10424),.clk(gclk));
	jnot g10187(.din(w_n10424_0[1]),.dout(n10425),.clk(gclk));
	jand g10188(.dina(w_n10425_0[1]),.dinb(n10421),.dout(n10426),.clk(gclk));
	jor g10189(.dina(n10426),.dinb(w_n10420_0[1]),.dout(n10427),.clk(gclk));
	jand g10190(.dina(w_n10427_0[2]),.dinb(w_asqrt38_24[2]),.dout(n10428),.clk(gclk));
	jor g10191(.dina(w_n10427_0[1]),.dinb(w_asqrt38_24[1]),.dout(n10429),.clk(gclk));
	jxor g10192(.dina(w_n9923_0[0]),.dinb(w_n4902_38[2]),.dout(n10430),.clk(gclk));
	jand g10193(.dina(n10430),.dinb(w_asqrt24_32[0]),.dout(n10431),.clk(gclk));
	jxor g10194(.dina(n10431),.dinb(w_n9928_0[0]),.dout(n10432),.clk(gclk));
	jnot g10195(.din(w_n10432_0[1]),.dout(n10433),.clk(gclk));
	jand g10196(.dina(w_n10433_0[1]),.dinb(n10429),.dout(n10434),.clk(gclk));
	jor g10197(.dina(n10434),.dinb(w_n10428_0[1]),.dout(n10435),.clk(gclk));
	jand g10198(.dina(w_n10435_0[2]),.dinb(w_asqrt39_21[1]),.dout(n10436),.clk(gclk));
	jxor g10199(.dina(w_n9930_0[0]),.dinb(w_n4582_35[2]),.dout(n10437),.clk(gclk));
	jand g10200(.dina(n10437),.dinb(w_asqrt24_31[2]),.dout(n10438),.clk(gclk));
	jxor g10201(.dina(n10438),.dinb(w_n9934_0[0]),.dout(n10439),.clk(gclk));
	jor g10202(.dina(w_n10435_0[1]),.dinb(w_asqrt39_21[0]),.dout(n10440),.clk(gclk));
	jand g10203(.dina(n10440),.dinb(w_n10439_0[1]),.dout(n10441),.clk(gclk));
	jor g10204(.dina(n10441),.dinb(w_n10436_0[1]),.dout(n10442),.clk(gclk));
	jand g10205(.dina(w_n10442_0[2]),.dinb(w_asqrt40_24[2]),.dout(n10443),.clk(gclk));
	jor g10206(.dina(w_n10442_0[1]),.dinb(w_asqrt40_24[1]),.dout(n10444),.clk(gclk));
	jxor g10207(.dina(w_n9938_0[0]),.dinb(w_n4249_39[1]),.dout(n10445),.clk(gclk));
	jand g10208(.dina(n10445),.dinb(w_asqrt24_31[1]),.dout(n10446),.clk(gclk));
	jxor g10209(.dina(n10446),.dinb(w_n9943_0[0]),.dout(n10447),.clk(gclk));
	jnot g10210(.din(w_n10447_0[1]),.dout(n10448),.clk(gclk));
	jand g10211(.dina(w_n10448_0[1]),.dinb(n10444),.dout(n10449),.clk(gclk));
	jor g10212(.dina(n10449),.dinb(w_n10443_0[1]),.dout(n10450),.clk(gclk));
	jand g10213(.dina(w_n10450_0[2]),.dinb(w_asqrt41_21[2]),.dout(n10451),.clk(gclk));
	jor g10214(.dina(w_n10450_0[1]),.dinb(w_asqrt41_21[1]),.dout(n10452),.clk(gclk));
	jxor g10215(.dina(w_n9945_0[0]),.dinb(w_n3955_36[1]),.dout(n10453),.clk(gclk));
	jand g10216(.dina(n10453),.dinb(w_asqrt24_31[0]),.dout(n10454),.clk(gclk));
	jxor g10217(.dina(n10454),.dinb(w_n9950_0[0]),.dout(n10455),.clk(gclk));
	jand g10218(.dina(w_n10455_0[1]),.dinb(n10452),.dout(n10456),.clk(gclk));
	jor g10219(.dina(n10456),.dinb(w_n10451_0[1]),.dout(n10457),.clk(gclk));
	jand g10220(.dina(w_n10457_0[2]),.dinb(w_asqrt42_25[0]),.dout(n10458),.clk(gclk));
	jor g10221(.dina(w_n10457_0[1]),.dinb(w_asqrt42_24[2]),.dout(n10459),.clk(gclk));
	jxor g10222(.dina(w_n9953_0[0]),.dinb(w_n3642_39[2]),.dout(n10460),.clk(gclk));
	jand g10223(.dina(n10460),.dinb(w_asqrt24_30[2]),.dout(n10461),.clk(gclk));
	jxor g10224(.dina(n10461),.dinb(w_n9958_0[0]),.dout(n10462),.clk(gclk));
	jnot g10225(.din(w_n10462_0[1]),.dout(n10463),.clk(gclk));
	jand g10226(.dina(w_n10463_0[1]),.dinb(n10459),.dout(n10464),.clk(gclk));
	jor g10227(.dina(n10464),.dinb(w_n10458_0[1]),.dout(n10465),.clk(gclk));
	jand g10228(.dina(w_n10465_0[2]),.dinb(w_asqrt43_22[0]),.dout(n10466),.clk(gclk));
	jor g10229(.dina(w_n10465_0[1]),.dinb(w_asqrt43_21[2]),.dout(n10467),.clk(gclk));
	jxor g10230(.dina(w_n9960_0[0]),.dinb(w_n3368_37[0]),.dout(n10468),.clk(gclk));
	jand g10231(.dina(n10468),.dinb(w_asqrt24_30[1]),.dout(n10469),.clk(gclk));
	jxor g10232(.dina(n10469),.dinb(w_n9965_0[0]),.dout(n10470),.clk(gclk));
	jand g10233(.dina(w_n10470_0[1]),.dinb(n10467),.dout(n10471),.clk(gclk));
	jor g10234(.dina(n10471),.dinb(w_n10466_0[1]),.dout(n10472),.clk(gclk));
	jand g10235(.dina(w_n10472_0[2]),.dinb(w_asqrt44_25[0]),.dout(n10473),.clk(gclk));
	jor g10236(.dina(w_n10472_0[1]),.dinb(w_asqrt44_24[2]),.dout(n10474),.clk(gclk));
	jxor g10237(.dina(w_n9968_0[0]),.dinb(w_n3089_40[1]),.dout(n10475),.clk(gclk));
	jand g10238(.dina(n10475),.dinb(w_asqrt24_30[0]),.dout(n10476),.clk(gclk));
	jxor g10239(.dina(n10476),.dinb(w_n9973_0[0]),.dout(n10477),.clk(gclk));
	jnot g10240(.din(w_n10477_0[1]),.dout(n10478),.clk(gclk));
	jand g10241(.dina(w_n10478_0[1]),.dinb(n10474),.dout(n10479),.clk(gclk));
	jor g10242(.dina(n10479),.dinb(w_n10473_0[1]),.dout(n10480),.clk(gclk));
	jand g10243(.dina(w_n10480_0[2]),.dinb(w_asqrt45_22[2]),.dout(n10481),.clk(gclk));
	jor g10244(.dina(w_n10480_0[1]),.dinb(w_asqrt45_22[1]),.dout(n10482),.clk(gclk));
	jxor g10245(.dina(w_n9975_0[0]),.dinb(w_n2833_38[0]),.dout(n10483),.clk(gclk));
	jand g10246(.dina(n10483),.dinb(w_asqrt24_29[2]),.dout(n10484),.clk(gclk));
	jxor g10247(.dina(n10484),.dinb(w_n9980_0[0]),.dout(n10485),.clk(gclk));
	jnot g10248(.din(w_n10485_0[1]),.dout(n10486),.clk(gclk));
	jand g10249(.dina(w_n10486_0[1]),.dinb(n10482),.dout(n10487),.clk(gclk));
	jor g10250(.dina(n10487),.dinb(w_n10481_0[1]),.dout(n10488),.clk(gclk));
	jand g10251(.dina(w_n10488_0[2]),.dinb(w_asqrt46_25[0]),.dout(n10489),.clk(gclk));
	jor g10252(.dina(w_n10488_0[1]),.dinb(w_asqrt46_24[2]),.dout(n10490),.clk(gclk));
	jxor g10253(.dina(w_n9982_0[0]),.dinb(w_n2572_40[2]),.dout(n10491),.clk(gclk));
	jand g10254(.dina(n10491),.dinb(w_asqrt24_29[1]),.dout(n10492),.clk(gclk));
	jxor g10255(.dina(n10492),.dinb(w_n9987_0[0]),.dout(n10493),.clk(gclk));
	jnot g10256(.din(w_n10493_0[1]),.dout(n10494),.clk(gclk));
	jand g10257(.dina(w_n10494_0[1]),.dinb(n10490),.dout(n10495),.clk(gclk));
	jor g10258(.dina(n10495),.dinb(w_n10489_0[1]),.dout(n10496),.clk(gclk));
	jand g10259(.dina(w_n10496_0[2]),.dinb(w_asqrt47_23[1]),.dout(n10497),.clk(gclk));
	jor g10260(.dina(w_n10496_0[1]),.dinb(w_asqrt47_23[0]),.dout(n10498),.clk(gclk));
	jxor g10261(.dina(w_n9989_0[0]),.dinb(w_n2345_38[2]),.dout(n10499),.clk(gclk));
	jand g10262(.dina(n10499),.dinb(w_asqrt24_29[0]),.dout(n10500),.clk(gclk));
	jxor g10263(.dina(n10500),.dinb(w_n9994_0[0]),.dout(n10501),.clk(gclk));
	jand g10264(.dina(w_n10501_0[1]),.dinb(n10498),.dout(n10502),.clk(gclk));
	jor g10265(.dina(n10502),.dinb(w_n10497_0[1]),.dout(n10503),.clk(gclk));
	jand g10266(.dina(w_n10503_0[2]),.dinb(w_asqrt48_25[1]),.dout(n10504),.clk(gclk));
	jor g10267(.dina(w_n10503_0[1]),.dinb(w_asqrt48_25[0]),.dout(n10505),.clk(gclk));
	jxor g10268(.dina(w_n9997_0[0]),.dinb(w_n2108_41[1]),.dout(n10506),.clk(gclk));
	jand g10269(.dina(n10506),.dinb(w_asqrt24_28[2]),.dout(n10507),.clk(gclk));
	jxor g10270(.dina(n10507),.dinb(w_n10002_0[0]),.dout(n10508),.clk(gclk));
	jnot g10271(.din(w_n10508_0[1]),.dout(n10509),.clk(gclk));
	jand g10272(.dina(w_n10509_0[1]),.dinb(n10505),.dout(n10510),.clk(gclk));
	jor g10273(.dina(n10510),.dinb(w_n10504_0[1]),.dout(n10511),.clk(gclk));
	jand g10274(.dina(w_n10511_0[2]),.dinb(w_asqrt49_23[2]),.dout(n10512),.clk(gclk));
	jor g10275(.dina(w_n10511_0[1]),.dinb(w_asqrt49_23[1]),.dout(n10513),.clk(gclk));
	jxor g10276(.dina(w_n10004_0[0]),.dinb(w_n1912_39[2]),.dout(n10514),.clk(gclk));
	jand g10277(.dina(n10514),.dinb(w_asqrt24_28[1]),.dout(n10515),.clk(gclk));
	jxor g10278(.dina(n10515),.dinb(w_n10009_0[0]),.dout(n10516),.clk(gclk));
	jand g10279(.dina(w_n10516_0[1]),.dinb(n10513),.dout(n10517),.clk(gclk));
	jor g10280(.dina(n10517),.dinb(w_n10512_0[1]),.dout(n10518),.clk(gclk));
	jand g10281(.dina(w_n10518_0[2]),.dinb(w_asqrt50_25[2]),.dout(n10519),.clk(gclk));
	jor g10282(.dina(w_n10518_0[1]),.dinb(w_asqrt50_25[1]),.dout(n10520),.clk(gclk));
	jxor g10283(.dina(w_n10012_0[0]),.dinb(w_n1699_42[0]),.dout(n10521),.clk(gclk));
	jand g10284(.dina(n10521),.dinb(w_asqrt24_28[0]),.dout(n10522),.clk(gclk));
	jxor g10285(.dina(n10522),.dinb(w_n10017_0[0]),.dout(n10523),.clk(gclk));
	jnot g10286(.din(w_n10523_0[1]),.dout(n10524),.clk(gclk));
	jand g10287(.dina(w_n10524_0[1]),.dinb(n10520),.dout(n10525),.clk(gclk));
	jor g10288(.dina(n10525),.dinb(w_n10519_0[1]),.dout(n10526),.clk(gclk));
	jand g10289(.dina(w_n10526_0[2]),.dinb(w_asqrt51_24[0]),.dout(n10527),.clk(gclk));
	jor g10290(.dina(w_n10526_0[1]),.dinb(w_asqrt51_23[2]),.dout(n10528),.clk(gclk));
	jxor g10291(.dina(w_n10019_0[0]),.dinb(w_n1516_40[1]),.dout(n10529),.clk(gclk));
	jand g10292(.dina(n10529),.dinb(w_asqrt24_27[2]),.dout(n10530),.clk(gclk));
	jxor g10293(.dina(n10530),.dinb(w_n10024_0[0]),.dout(n10531),.clk(gclk));
	jand g10294(.dina(w_n10531_0[1]),.dinb(n10528),.dout(n10532),.clk(gclk));
	jor g10295(.dina(n10532),.dinb(w_n10527_0[1]),.dout(n10533),.clk(gclk));
	jand g10296(.dina(w_n10533_0[2]),.dinb(w_asqrt52_25[2]),.dout(n10534),.clk(gclk));
	jor g10297(.dina(w_n10533_0[1]),.dinb(w_asqrt52_25[1]),.dout(n10535),.clk(gclk));
	jxor g10298(.dina(w_n10027_0[0]),.dinb(w_n1332_42[0]),.dout(n10536),.clk(gclk));
	jand g10299(.dina(n10536),.dinb(w_asqrt24_27[1]),.dout(n10537),.clk(gclk));
	jxor g10300(.dina(n10537),.dinb(w_n10032_0[0]),.dout(n10538),.clk(gclk));
	jnot g10301(.din(w_n10538_0[1]),.dout(n10539),.clk(gclk));
	jand g10302(.dina(w_n10539_0[1]),.dinb(n10535),.dout(n10540),.clk(gclk));
	jor g10303(.dina(n10540),.dinb(w_n10534_0[1]),.dout(n10541),.clk(gclk));
	jand g10304(.dina(w_n10541_0[2]),.dinb(w_asqrt53_24[2]),.dout(n10542),.clk(gclk));
	jor g10305(.dina(w_n10541_0[1]),.dinb(w_asqrt53_24[1]),.dout(n10543),.clk(gclk));
	jxor g10306(.dina(w_n10034_0[0]),.dinb(w_n1173_41[0]),.dout(n10544),.clk(gclk));
	jand g10307(.dina(n10544),.dinb(w_asqrt24_27[0]),.dout(n10545),.clk(gclk));
	jxor g10308(.dina(n10545),.dinb(w_n10039_0[0]),.dout(n10546),.clk(gclk));
	jand g10309(.dina(w_n10546_0[1]),.dinb(n10543),.dout(n10547),.clk(gclk));
	jor g10310(.dina(n10547),.dinb(w_n10542_0[1]),.dout(n10548),.clk(gclk));
	jand g10311(.dina(w_n10548_0[2]),.dinb(w_asqrt54_25[2]),.dout(n10549),.clk(gclk));
	jor g10312(.dina(w_n10548_0[1]),.dinb(w_asqrt54_25[1]),.dout(n10550),.clk(gclk));
	jxor g10313(.dina(w_n10042_0[0]),.dinb(w_n1008_43[0]),.dout(n10551),.clk(gclk));
	jand g10314(.dina(n10551),.dinb(w_asqrt24_26[2]),.dout(n10552),.clk(gclk));
	jxor g10315(.dina(n10552),.dinb(w_n10047_0[0]),.dout(n10553),.clk(gclk));
	jand g10316(.dina(w_n10553_0[1]),.dinb(n10550),.dout(n10554),.clk(gclk));
	jor g10317(.dina(n10554),.dinb(w_n10549_0[1]),.dout(n10555),.clk(gclk));
	jand g10318(.dina(w_n10555_0[2]),.dinb(w_asqrt55_25[0]),.dout(n10556),.clk(gclk));
	jor g10319(.dina(w_n10555_0[1]),.dinb(w_asqrt55_24[2]),.dout(n10557),.clk(gclk));
	jxor g10320(.dina(w_n10050_0[0]),.dinb(w_n884_42[0]),.dout(n10558),.clk(gclk));
	jand g10321(.dina(n10558),.dinb(w_asqrt24_26[1]),.dout(n10559),.clk(gclk));
	jxor g10322(.dina(n10559),.dinb(w_n10055_0[0]),.dout(n10560),.clk(gclk));
	jand g10323(.dina(w_n10560_0[1]),.dinb(n10557),.dout(n10561),.clk(gclk));
	jor g10324(.dina(n10561),.dinb(w_n10556_0[1]),.dout(n10562),.clk(gclk));
	jand g10325(.dina(w_n10562_0[2]),.dinb(w_asqrt56_26[0]),.dout(n10563),.clk(gclk));
	jor g10326(.dina(w_n10562_0[1]),.dinb(w_asqrt56_25[2]),.dout(n10564),.clk(gclk));
	jxor g10327(.dina(w_n10058_0[0]),.dinb(w_n743_43[0]),.dout(n10565),.clk(gclk));
	jand g10328(.dina(n10565),.dinb(w_asqrt24_26[0]),.dout(n10566),.clk(gclk));
	jxor g10329(.dina(n10566),.dinb(w_n10063_0[0]),.dout(n10567),.clk(gclk));
	jnot g10330(.din(w_n10567_0[1]),.dout(n10568),.clk(gclk));
	jand g10331(.dina(w_n10568_0[1]),.dinb(n10564),.dout(n10569),.clk(gclk));
	jor g10332(.dina(n10569),.dinb(w_n10563_0[1]),.dout(n10570),.clk(gclk));
	jand g10333(.dina(w_n10570_0[2]),.dinb(w_asqrt57_25[2]),.dout(n10571),.clk(gclk));
	jor g10334(.dina(w_n10570_0[1]),.dinb(w_asqrt57_25[1]),.dout(n10572),.clk(gclk));
	jxor g10335(.dina(w_n10065_0[0]),.dinb(w_n635_43[0]),.dout(n10573),.clk(gclk));
	jand g10336(.dina(n10573),.dinb(w_asqrt24_25[2]),.dout(n10574),.clk(gclk));
	jxor g10337(.dina(n10574),.dinb(w_n10070_0[0]),.dout(n10575),.clk(gclk));
	jnot g10338(.din(w_n10575_0[1]),.dout(n10576),.clk(gclk));
	jand g10339(.dina(w_n10576_0[1]),.dinb(n10572),.dout(n10577),.clk(gclk));
	jor g10340(.dina(n10577),.dinb(w_n10571_0[1]),.dout(n10578),.clk(gclk));
	jand g10341(.dina(w_n10578_0[2]),.dinb(w_asqrt58_26[1]),.dout(n10579),.clk(gclk));
	jor g10342(.dina(w_n10578_0[1]),.dinb(w_asqrt58_26[0]),.dout(n10580),.clk(gclk));
	jxor g10343(.dina(w_n10072_0[0]),.dinb(w_n515_44[0]),.dout(n10581),.clk(gclk));
	jand g10344(.dina(n10581),.dinb(w_asqrt24_25[1]),.dout(n10582),.clk(gclk));
	jxor g10345(.dina(n10582),.dinb(w_n10077_0[0]),.dout(n10583),.clk(gclk));
	jnot g10346(.din(w_n10583_0[1]),.dout(n10584),.clk(gclk));
	jand g10347(.dina(w_n10584_0[1]),.dinb(n10580),.dout(n10585),.clk(gclk));
	jor g10348(.dina(n10585),.dinb(w_n10579_0[1]),.dout(n10586),.clk(gclk));
	jand g10349(.dina(w_n10586_0[2]),.dinb(w_asqrt59_26[0]),.dout(n10587),.clk(gclk));
	jor g10350(.dina(w_n10586_0[1]),.dinb(w_asqrt59_25[2]),.dout(n10588),.clk(gclk));
	jxor g10351(.dina(w_n10079_0[0]),.dinb(w_n443_44[0]),.dout(n10589),.clk(gclk));
	jand g10352(.dina(n10589),.dinb(w_asqrt24_25[0]),.dout(n10590),.clk(gclk));
	jxor g10353(.dina(n10590),.dinb(w_n10084_0[0]),.dout(n10591),.clk(gclk));
	jand g10354(.dina(w_n10591_0[1]),.dinb(n10588),.dout(n10592),.clk(gclk));
	jor g10355(.dina(n10592),.dinb(w_n10587_0[1]),.dout(n10593),.clk(gclk));
	jand g10356(.dina(w_n10593_0[2]),.dinb(w_asqrt60_26[1]),.dout(n10594),.clk(gclk));
	jor g10357(.dina(w_n10593_0[1]),.dinb(w_asqrt60_26[0]),.dout(n10595),.clk(gclk));
	jxor g10358(.dina(w_n10087_0[0]),.dinb(w_n352_44[1]),.dout(n10596),.clk(gclk));
	jand g10359(.dina(n10596),.dinb(w_asqrt24_24[2]),.dout(n10597),.clk(gclk));
	jxor g10360(.dina(n10597),.dinb(w_n10092_0[0]),.dout(n10598),.clk(gclk));
	jnot g10361(.din(w_n10598_0[1]),.dout(n10599),.clk(gclk));
	jand g10362(.dina(w_n10599_0[1]),.dinb(n10595),.dout(n10600),.clk(gclk));
	jor g10363(.dina(n10600),.dinb(w_n10594_0[1]),.dout(n10601),.clk(gclk));
	jand g10364(.dina(w_n10601_0[2]),.dinb(w_asqrt61_26[1]),.dout(n10602),.clk(gclk));
	jor g10365(.dina(w_n10601_0[1]),.dinb(w_asqrt61_26[0]),.dout(n10603),.clk(gclk));
	jxor g10366(.dina(w_n10094_0[0]),.dinb(w_n294_44[2]),.dout(n10604),.clk(gclk));
	jand g10367(.dina(n10604),.dinb(w_asqrt24_24[1]),.dout(n10605),.clk(gclk));
	jxor g10368(.dina(n10605),.dinb(w_n10099_0[0]),.dout(n10606),.clk(gclk));
	jnot g10369(.din(w_n10606_0[1]),.dout(n10607),.clk(gclk));
	jand g10370(.dina(w_n10607_0[1]),.dinb(n10603),.dout(n10608),.clk(gclk));
	jor g10371(.dina(n10608),.dinb(w_n10602_0[1]),.dout(n10609),.clk(gclk));
	jand g10372(.dina(w_n10609_0[2]),.dinb(w_asqrt62_26[1]),.dout(n10610),.clk(gclk));
	jnot g10373(.din(w_n10610_0[1]),.dout(n10611),.clk(gclk));
	jnot g10374(.din(w_n10602_0[0]),.dout(n10612),.clk(gclk));
	jnot g10375(.din(w_n10594_0[0]),.dout(n10613),.clk(gclk));
	jnot g10376(.din(w_n10587_0[0]),.dout(n10614),.clk(gclk));
	jnot g10377(.din(w_n10579_0[0]),.dout(n10615),.clk(gclk));
	jnot g10378(.din(w_n10571_0[0]),.dout(n10616),.clk(gclk));
	jnot g10379(.din(w_n10563_0[0]),.dout(n10617),.clk(gclk));
	jnot g10380(.din(w_n10556_0[0]),.dout(n10618),.clk(gclk));
	jnot g10381(.din(w_n10549_0[0]),.dout(n10619),.clk(gclk));
	jnot g10382(.din(w_n10542_0[0]),.dout(n10620),.clk(gclk));
	jnot g10383(.din(w_n10534_0[0]),.dout(n10621),.clk(gclk));
	jnot g10384(.din(w_n10527_0[0]),.dout(n10622),.clk(gclk));
	jnot g10385(.din(w_n10519_0[0]),.dout(n10623),.clk(gclk));
	jnot g10386(.din(w_n10512_0[0]),.dout(n10624),.clk(gclk));
	jnot g10387(.din(w_n10504_0[0]),.dout(n10625),.clk(gclk));
	jnot g10388(.din(w_n10497_0[0]),.dout(n10626),.clk(gclk));
	jnot g10389(.din(w_n10489_0[0]),.dout(n10627),.clk(gclk));
	jnot g10390(.din(w_n10481_0[0]),.dout(n10628),.clk(gclk));
	jnot g10391(.din(w_n10473_0[0]),.dout(n10629),.clk(gclk));
	jnot g10392(.din(w_n10466_0[0]),.dout(n10630),.clk(gclk));
	jnot g10393(.din(w_n10458_0[0]),.dout(n10631),.clk(gclk));
	jnot g10394(.din(w_n10451_0[0]),.dout(n10632),.clk(gclk));
	jnot g10395(.din(w_n10443_0[0]),.dout(n10633),.clk(gclk));
	jnot g10396(.din(w_n10436_0[0]),.dout(n10634),.clk(gclk));
	jnot g10397(.din(w_n10439_0[0]),.dout(n10635),.clk(gclk));
	jnot g10398(.din(w_n10428_0[0]),.dout(n10636),.clk(gclk));
	jnot g10399(.din(w_n10420_0[0]),.dout(n10637),.clk(gclk));
	jnot g10400(.din(w_n10412_0[0]),.dout(n10638),.clk(gclk));
	jnot g10401(.din(w_n10404_0[0]),.dout(n10639),.clk(gclk));
	jnot g10402(.din(w_n10396_0[0]),.dout(n10640),.clk(gclk));
	jnot g10403(.din(w_n10389_0[0]),.dout(n10641),.clk(gclk));
	jnot g10404(.din(w_n10381_0[0]),.dout(n10642),.clk(gclk));
	jnot g10405(.din(w_n10373_0[0]),.dout(n10643),.clk(gclk));
	jnot g10406(.din(w_n10365_0[0]),.dout(n10644),.clk(gclk));
	jnot g10407(.din(w_n10358_0[0]),.dout(n10645),.clk(gclk));
	jnot g10408(.din(w_n10350_0[0]),.dout(n10646),.clk(gclk));
	jnot g10409(.din(w_n10343_0[0]),.dout(n10647),.clk(gclk));
	jnot g10410(.din(w_n10333_0[0]),.dout(n10648),.clk(gclk));
	jnot g10411(.din(w_n10140_0[0]),.dout(n10649),.clk(gclk));
	jnot g10412(.din(w_n10137_0[0]),.dout(n10650),.clk(gclk));
	jor g10413(.dina(w_n10328_30[1]),.dinb(w_n9834_0[2]),.dout(n10651),.clk(gclk));
	jand g10414(.dina(n10651),.dinb(n10650),.dout(n10652),.clk(gclk));
	jand g10415(.dina(n10652),.dinb(w_n9832_35[2]),.dout(n10653),.clk(gclk));
	jor g10416(.dina(w_n10328_30[0]),.dinb(w_a48_0[0]),.dout(n10654),.clk(gclk));
	jand g10417(.dina(n10654),.dinb(w_a49_0[0]),.dout(n10655),.clk(gclk));
	jand g10418(.dina(w_asqrt24_24[0]),.dinb(w_n9836_0[0]),.dout(n10656),.clk(gclk));
	jor g10419(.dina(n10656),.dinb(n10655),.dout(n10657),.clk(gclk));
	jor g10420(.dina(n10657),.dinb(n10653),.dout(n10658),.clk(gclk));
	jand g10421(.dina(n10658),.dinb(n10649),.dout(n10659),.clk(gclk));
	jand g10422(.dina(n10659),.dinb(w_n9369_30[1]),.dout(n10660),.clk(gclk));
	jor g10423(.dina(w_n10339_0[0]),.dinb(n10660),.dout(n10661),.clk(gclk));
	jand g10424(.dina(n10661),.dinb(n10648),.dout(n10662),.clk(gclk));
	jand g10425(.dina(n10662),.dinb(w_n8890_36[0]),.dout(n10663),.clk(gclk));
	jnot g10426(.din(w_n10347_0[0]),.dout(n10664),.clk(gclk));
	jor g10427(.dina(w_n10664_0[1]),.dinb(n10663),.dout(n10665),.clk(gclk));
	jand g10428(.dina(n10665),.dinb(n10647),.dout(n10666),.clk(gclk));
	jand g10429(.dina(n10666),.dinb(w_n8449_31[0]),.dout(n10667),.clk(gclk));
	jor g10430(.dina(w_n10354_0[0]),.dinb(n10667),.dout(n10668),.clk(gclk));
	jand g10431(.dina(n10668),.dinb(n10646),.dout(n10669),.clk(gclk));
	jand g10432(.dina(n10669),.dinb(w_n8003_36[2]),.dout(n10670),.clk(gclk));
	jnot g10433(.din(w_n10362_0[0]),.dout(n10671),.clk(gclk));
	jor g10434(.dina(w_n10671_0[1]),.dinb(n10670),.dout(n10672),.clk(gclk));
	jand g10435(.dina(n10672),.dinb(n10645),.dout(n10673),.clk(gclk));
	jand g10436(.dina(n10673),.dinb(w_n7581_32[0]),.dout(n10674),.clk(gclk));
	jor g10437(.dina(w_n10369_0[0]),.dinb(n10674),.dout(n10675),.clk(gclk));
	jand g10438(.dina(n10675),.dinb(n10644),.dout(n10676),.clk(gclk));
	jand g10439(.dina(n10676),.dinb(w_n7154_37[0]),.dout(n10677),.clk(gclk));
	jor g10440(.dina(w_n10377_0[0]),.dinb(n10677),.dout(n10678),.clk(gclk));
	jand g10441(.dina(n10678),.dinb(n10643),.dout(n10679),.clk(gclk));
	jand g10442(.dina(n10679),.dinb(w_n6758_32[2]),.dout(n10680),.clk(gclk));
	jor g10443(.dina(w_n10385_0[0]),.dinb(n10680),.dout(n10681),.clk(gclk));
	jand g10444(.dina(n10681),.dinb(n10642),.dout(n10682),.clk(gclk));
	jand g10445(.dina(n10682),.dinb(w_n6357_37[1]),.dout(n10683),.clk(gclk));
	jnot g10446(.din(w_n10393_0[0]),.dout(n10684),.clk(gclk));
	jor g10447(.dina(w_n10684_0[1]),.dinb(n10683),.dout(n10685),.clk(gclk));
	jand g10448(.dina(n10685),.dinb(n10641),.dout(n10686),.clk(gclk));
	jand g10449(.dina(n10686),.dinb(w_n5989_33[1]),.dout(n10687),.clk(gclk));
	jor g10450(.dina(w_n10400_0[0]),.dinb(n10687),.dout(n10688),.clk(gclk));
	jand g10451(.dina(n10688),.dinb(n10640),.dout(n10689),.clk(gclk));
	jand g10452(.dina(n10689),.dinb(w_n5606_37[2]),.dout(n10690),.clk(gclk));
	jor g10453(.dina(w_n10408_0[0]),.dinb(n10690),.dout(n10691),.clk(gclk));
	jand g10454(.dina(n10691),.dinb(n10639),.dout(n10692),.clk(gclk));
	jand g10455(.dina(n10692),.dinb(w_n5259_34[1]),.dout(n10693),.clk(gclk));
	jor g10456(.dina(w_n10416_0[0]),.dinb(n10693),.dout(n10694),.clk(gclk));
	jand g10457(.dina(n10694),.dinb(n10638),.dout(n10695),.clk(gclk));
	jand g10458(.dina(n10695),.dinb(w_n4902_38[1]),.dout(n10696),.clk(gclk));
	jor g10459(.dina(w_n10424_0[0]),.dinb(n10696),.dout(n10697),.clk(gclk));
	jand g10460(.dina(n10697),.dinb(n10637),.dout(n10698),.clk(gclk));
	jand g10461(.dina(n10698),.dinb(w_n4582_35[1]),.dout(n10699),.clk(gclk));
	jor g10462(.dina(w_n10432_0[0]),.dinb(n10699),.dout(n10700),.clk(gclk));
	jand g10463(.dina(n10700),.dinb(n10636),.dout(n10701),.clk(gclk));
	jand g10464(.dina(n10701),.dinb(w_n4249_39[0]),.dout(n10702),.clk(gclk));
	jor g10465(.dina(n10702),.dinb(w_n10635_0[1]),.dout(n10703),.clk(gclk));
	jand g10466(.dina(n10703),.dinb(n10634),.dout(n10704),.clk(gclk));
	jand g10467(.dina(n10704),.dinb(w_n3955_36[0]),.dout(n10705),.clk(gclk));
	jor g10468(.dina(w_n10447_0[0]),.dinb(n10705),.dout(n10706),.clk(gclk));
	jand g10469(.dina(n10706),.dinb(n10633),.dout(n10707),.clk(gclk));
	jand g10470(.dina(n10707),.dinb(w_n3642_39[1]),.dout(n10708),.clk(gclk));
	jnot g10471(.din(w_n10455_0[0]),.dout(n10709),.clk(gclk));
	jor g10472(.dina(w_n10709_0[1]),.dinb(n10708),.dout(n10710),.clk(gclk));
	jand g10473(.dina(n10710),.dinb(n10632),.dout(n10711),.clk(gclk));
	jand g10474(.dina(n10711),.dinb(w_n3368_36[2]),.dout(n10712),.clk(gclk));
	jor g10475(.dina(w_n10462_0[0]),.dinb(n10712),.dout(n10713),.clk(gclk));
	jand g10476(.dina(n10713),.dinb(n10631),.dout(n10714),.clk(gclk));
	jand g10477(.dina(n10714),.dinb(w_n3089_40[0]),.dout(n10715),.clk(gclk));
	jnot g10478(.din(w_n10470_0[0]),.dout(n10716),.clk(gclk));
	jor g10479(.dina(w_n10716_0[1]),.dinb(n10715),.dout(n10717),.clk(gclk));
	jand g10480(.dina(n10717),.dinb(n10630),.dout(n10718),.clk(gclk));
	jand g10481(.dina(n10718),.dinb(w_n2833_37[2]),.dout(n10719),.clk(gclk));
	jor g10482(.dina(w_n10477_0[0]),.dinb(n10719),.dout(n10720),.clk(gclk));
	jand g10483(.dina(n10720),.dinb(n10629),.dout(n10721),.clk(gclk));
	jand g10484(.dina(n10721),.dinb(w_n2572_40[1]),.dout(n10722),.clk(gclk));
	jor g10485(.dina(w_n10485_0[0]),.dinb(n10722),.dout(n10723),.clk(gclk));
	jand g10486(.dina(n10723),.dinb(n10628),.dout(n10724),.clk(gclk));
	jand g10487(.dina(n10724),.dinb(w_n2345_38[1]),.dout(n10725),.clk(gclk));
	jor g10488(.dina(w_n10493_0[0]),.dinb(n10725),.dout(n10726),.clk(gclk));
	jand g10489(.dina(n10726),.dinb(n10627),.dout(n10727),.clk(gclk));
	jand g10490(.dina(n10727),.dinb(w_n2108_41[0]),.dout(n10728),.clk(gclk));
	jnot g10491(.din(w_n10501_0[0]),.dout(n10729),.clk(gclk));
	jor g10492(.dina(w_n10729_0[1]),.dinb(n10728),.dout(n10730),.clk(gclk));
	jand g10493(.dina(n10730),.dinb(n10626),.dout(n10731),.clk(gclk));
	jand g10494(.dina(n10731),.dinb(w_n1912_39[1]),.dout(n10732),.clk(gclk));
	jor g10495(.dina(w_n10508_0[0]),.dinb(n10732),.dout(n10733),.clk(gclk));
	jand g10496(.dina(n10733),.dinb(n10625),.dout(n10734),.clk(gclk));
	jand g10497(.dina(n10734),.dinb(w_n1699_41[2]),.dout(n10735),.clk(gclk));
	jnot g10498(.din(w_n10516_0[0]),.dout(n10736),.clk(gclk));
	jor g10499(.dina(w_n10736_0[1]),.dinb(n10735),.dout(n10737),.clk(gclk));
	jand g10500(.dina(n10737),.dinb(n10624),.dout(n10738),.clk(gclk));
	jand g10501(.dina(n10738),.dinb(w_n1516_40[0]),.dout(n10739),.clk(gclk));
	jor g10502(.dina(w_n10523_0[0]),.dinb(n10739),.dout(n10740),.clk(gclk));
	jand g10503(.dina(n10740),.dinb(n10623),.dout(n10741),.clk(gclk));
	jand g10504(.dina(n10741),.dinb(w_n1332_41[2]),.dout(n10742),.clk(gclk));
	jnot g10505(.din(w_n10531_0[0]),.dout(n10743),.clk(gclk));
	jor g10506(.dina(w_n10743_0[1]),.dinb(n10742),.dout(n10744),.clk(gclk));
	jand g10507(.dina(n10744),.dinb(n10622),.dout(n10745),.clk(gclk));
	jand g10508(.dina(n10745),.dinb(w_n1173_40[2]),.dout(n10746),.clk(gclk));
	jor g10509(.dina(w_n10538_0[0]),.dinb(n10746),.dout(n10747),.clk(gclk));
	jand g10510(.dina(n10747),.dinb(n10621),.dout(n10748),.clk(gclk));
	jand g10511(.dina(n10748),.dinb(w_n1008_42[2]),.dout(n10749),.clk(gclk));
	jnot g10512(.din(w_n10546_0[0]),.dout(n10750),.clk(gclk));
	jor g10513(.dina(w_n10750_0[1]),.dinb(n10749),.dout(n10751),.clk(gclk));
	jand g10514(.dina(n10751),.dinb(n10620),.dout(n10752),.clk(gclk));
	jand g10515(.dina(n10752),.dinb(w_n884_41[2]),.dout(n10753),.clk(gclk));
	jnot g10516(.din(w_n10553_0[0]),.dout(n10754),.clk(gclk));
	jor g10517(.dina(w_n10754_0[1]),.dinb(n10753),.dout(n10755),.clk(gclk));
	jand g10518(.dina(n10755),.dinb(n10619),.dout(n10756),.clk(gclk));
	jand g10519(.dina(n10756),.dinb(w_n743_42[2]),.dout(n10757),.clk(gclk));
	jnot g10520(.din(w_n10560_0[0]),.dout(n10758),.clk(gclk));
	jor g10521(.dina(w_n10758_0[1]),.dinb(n10757),.dout(n10759),.clk(gclk));
	jand g10522(.dina(n10759),.dinb(n10618),.dout(n10760),.clk(gclk));
	jand g10523(.dina(n10760),.dinb(w_n635_42[2]),.dout(n10761),.clk(gclk));
	jor g10524(.dina(w_n10567_0[0]),.dinb(n10761),.dout(n10762),.clk(gclk));
	jand g10525(.dina(n10762),.dinb(n10617),.dout(n10763),.clk(gclk));
	jand g10526(.dina(n10763),.dinb(w_n515_43[2]),.dout(n10764),.clk(gclk));
	jor g10527(.dina(w_n10575_0[0]),.dinb(n10764),.dout(n10765),.clk(gclk));
	jand g10528(.dina(n10765),.dinb(n10616),.dout(n10766),.clk(gclk));
	jand g10529(.dina(n10766),.dinb(w_n443_43[2]),.dout(n10767),.clk(gclk));
	jor g10530(.dina(w_n10583_0[0]),.dinb(n10767),.dout(n10768),.clk(gclk));
	jand g10531(.dina(n10768),.dinb(n10615),.dout(n10769),.clk(gclk));
	jand g10532(.dina(n10769),.dinb(w_n352_44[0]),.dout(n10770),.clk(gclk));
	jnot g10533(.din(w_n10591_0[0]),.dout(n10771),.clk(gclk));
	jor g10534(.dina(w_n10771_0[1]),.dinb(n10770),.dout(n10772),.clk(gclk));
	jand g10535(.dina(n10772),.dinb(n10614),.dout(n10773),.clk(gclk));
	jand g10536(.dina(n10773),.dinb(w_n294_44[1]),.dout(n10774),.clk(gclk));
	jor g10537(.dina(w_n10598_0[0]),.dinb(n10774),.dout(n10775),.clk(gclk));
	jand g10538(.dina(n10775),.dinb(n10613),.dout(n10776),.clk(gclk));
	jand g10539(.dina(n10776),.dinb(w_n239_44[2]),.dout(n10777),.clk(gclk));
	jor g10540(.dina(w_n10606_0[0]),.dinb(n10777),.dout(n10778),.clk(gclk));
	jand g10541(.dina(n10778),.dinb(n10612),.dout(n10779),.clk(gclk));
	jand g10542(.dina(n10779),.dinb(w_n221_45[0]),.dout(n10780),.clk(gclk));
	jxor g10543(.dina(w_n10101_0[0]),.dinb(w_n239_44[1]),.dout(n10781),.clk(gclk));
	jand g10544(.dina(n10781),.dinb(w_asqrt24_23[2]),.dout(n10782),.clk(gclk));
	jxor g10545(.dina(n10782),.dinb(w_n10106_0[0]),.dout(n10783),.clk(gclk));
	jor g10546(.dina(w_n10783_0[1]),.dinb(n10780),.dout(n10784),.clk(gclk));
	jand g10547(.dina(n10784),.dinb(n10611),.dout(n10785),.clk(gclk));
	jxor g10548(.dina(w_n10108_0[0]),.dinb(w_n221_44[2]),.dout(n10786),.clk(gclk));
	jand g10549(.dina(n10786),.dinb(w_asqrt24_23[1]),.dout(n10787),.clk(gclk));
	jxor g10550(.dina(n10787),.dinb(w_n10114_0[0]),.dout(n10788),.clk(gclk));
	jor g10551(.dina(w_n10788_1[1]),.dinb(w_n10785_0[2]),.dout(n10789),.clk(gclk));
	jand g10552(.dina(w_asqrt24_23[0]),.dinb(w_n10323_0[0]),.dout(n10790),.clk(gclk));
	jor g10553(.dina(n10790),.dinb(w_n10125_0[2]),.dout(n10791),.clk(gclk));
	jor g10554(.dina(w_n10791_0[1]),.dinb(w_n10789_0[1]),.dout(n10792),.clk(gclk));
	jand g10555(.dina(n10792),.dinb(w_n218_18[2]),.dout(n10793),.clk(gclk));
	jand g10556(.dina(w_n10328_29[2]),.dinb(w_n10119_0[1]),.dout(n10794),.clk(gclk));
	jand g10557(.dina(w_n10788_1[0]),.dinb(w_n10785_0[1]),.dout(n10795),.clk(gclk));
	jor g10558(.dina(w_n10795_0[2]),.dinb(w_n10794_0[1]),.dout(n10796),.clk(gclk));
	jand g10559(.dina(w_n10328_29[1]),.dinb(w_n10116_0[0]),.dout(n10797),.clk(gclk));
	jnot g10560(.din(n10797),.dout(n10798),.clk(gclk));
	jnot g10561(.din(w_n10125_0[1]),.dout(n10799),.clk(gclk));
	jand g10562(.dina(w_n10120_0[0]),.dinb(w_asqrt63_33[1]),.dout(n10800),.clk(gclk));
	jand g10563(.dina(n10800),.dinb(n10799),.dout(n10801),.clk(gclk));
	jand g10564(.dina(w_n10801_0[1]),.dinb(n10798),.dout(n10802),.clk(gclk));
	jor g10565(.dina(w_n10802_0[1]),.dinb(n10796),.dout(n10803),.clk(gclk));
	jor g10566(.dina(n10803),.dinb(w_n10793_0[1]),.dout(asqrt_fa_24),.clk(gclk));
	jnot g10567(.din(w_a44_0[2]),.dout(n10805),.clk(gclk));
	jnot g10568(.din(w_a45_0[1]),.dout(n10806),.clk(gclk));
	jand g10569(.dina(w_n10806_0[1]),.dinb(w_n10805_1[2]),.dout(n10807),.clk(gclk));
	jand g10570(.dina(w_n10807_0[2]),.dinb(w_n10134_1[0]),.dout(n10808),.clk(gclk));
	jnot g10571(.din(w_n10808_0[1]),.dout(n10809),.clk(gclk));
	jor g10572(.dina(w_n10609_0[1]),.dinb(w_asqrt62_26[0]),.dout(n10810),.clk(gclk));
	jnot g10573(.din(w_n10783_0[0]),.dout(n10811),.clk(gclk));
	jand g10574(.dina(w_n10811_0[1]),.dinb(n10810),.dout(n10812),.clk(gclk));
	jor g10575(.dina(n10812),.dinb(w_n10610_0[0]),.dout(n10813),.clk(gclk));
	jnot g10576(.din(w_n10788_0[2]),.dout(n10814),.clk(gclk));
	jand g10577(.dina(w_n10814_0[1]),.dinb(w_n10813_0[1]),.dout(n10815),.clk(gclk));
	jnot g10578(.din(w_n10791_0[0]),.dout(n10816),.clk(gclk));
	jand g10579(.dina(n10816),.dinb(w_n10815_0[1]),.dout(n10817),.clk(gclk));
	jor g10580(.dina(n10817),.dinb(w_asqrt63_33[0]),.dout(n10818),.clk(gclk));
	jnot g10581(.din(w_n10794_0[0]),.dout(n10819),.clk(gclk));
	jor g10582(.dina(w_n10814_0[0]),.dinb(w_n10813_0[0]),.dout(n10820),.clk(gclk));
	jand g10583(.dina(w_n10820_0[2]),.dinb(n10819),.dout(n10821),.clk(gclk));
	jnot g10584(.din(w_n10802_0[0]),.dout(n10822),.clk(gclk));
	jand g10585(.dina(n10822),.dinb(n10821),.dout(n10823),.clk(gclk));
	jand g10586(.dina(n10823),.dinb(n10818),.dout(n10824),.clk(gclk));
	jor g10587(.dina(w_n10824_47[2]),.dinb(w_n10134_0[2]),.dout(n10825),.clk(gclk));
	jand g10588(.dina(n10825),.dinb(n10809),.dout(n10826),.clk(gclk));
	jor g10589(.dina(w_n10826_0[2]),.dinb(w_n10328_29[0]),.dout(n10827),.clk(gclk));
	jand g10590(.dina(w_n10826_0[1]),.dinb(w_n10328_28[2]),.dout(n10828),.clk(gclk));
	jor g10591(.dina(w_n10824_47[1]),.dinb(w_a46_1[0]),.dout(n10829),.clk(gclk));
	jand g10592(.dina(n10829),.dinb(w_a47_0[0]),.dout(n10830),.clk(gclk));
	jand g10593(.dina(w_asqrt23_18),.dinb(w_n10136_0[1]),.dout(n10831),.clk(gclk));
	jor g10594(.dina(n10831),.dinb(n10830),.dout(n10832),.clk(gclk));
	jor g10595(.dina(n10832),.dinb(n10828),.dout(n10833),.clk(gclk));
	jand g10596(.dina(n10833),.dinb(w_n10827_0[1]),.dout(n10834),.clk(gclk));
	jor g10597(.dina(w_n10834_0[2]),.dinb(w_n9832_35[1]),.dout(n10835),.clk(gclk));
	jand g10598(.dina(w_n10834_0[1]),.dinb(w_n9832_35[0]),.dout(n10836),.clk(gclk));
	jnot g10599(.din(w_n10136_0[0]),.dout(n10837),.clk(gclk));
	jor g10600(.dina(w_n10824_47[0]),.dinb(n10837),.dout(n10838),.clk(gclk));
	jor g10601(.dina(w_n10801_0[0]),.dinb(w_n10328_28[1]),.dout(n10839),.clk(gclk));
	jor g10602(.dina(n10839),.dinb(w_n10795_0[1]),.dout(n10840),.clk(gclk));
	jor g10603(.dina(n10840),.dinb(w_n10793_0[0]),.dout(n10841),.clk(gclk));
	jand g10604(.dina(n10841),.dinb(w_n10838_0[1]),.dout(n10842),.clk(gclk));
	jxor g10605(.dina(n10842),.dinb(w_n9834_0[1]),.dout(n10843),.clk(gclk));
	jor g10606(.dina(w_n10843_0[2]),.dinb(n10836),.dout(n10844),.clk(gclk));
	jand g10607(.dina(n10844),.dinb(w_n10835_0[1]),.dout(n10845),.clk(gclk));
	jor g10608(.dina(w_n10845_0[2]),.dinb(w_n9369_30[0]),.dout(n10846),.clk(gclk));
	jand g10609(.dina(w_n10845_0[1]),.dinb(w_n9369_29[2]),.dout(n10847),.clk(gclk));
	jxor g10610(.dina(w_n10139_0[0]),.dinb(w_n9832_34[2]),.dout(n10848),.clk(gclk));
	jor g10611(.dina(n10848),.dinb(w_n10824_46[2]),.dout(n10849),.clk(gclk));
	jxor g10612(.dina(n10849),.dinb(w_n10330_0[0]),.dout(n10850),.clk(gclk));
	jor g10613(.dina(w_n10850_0[2]),.dinb(n10847),.dout(n10851),.clk(gclk));
	jand g10614(.dina(n10851),.dinb(w_n10846_0[1]),.dout(n10852),.clk(gclk));
	jor g10615(.dina(w_n10852_0[2]),.dinb(w_n8890_35[2]),.dout(n10853),.clk(gclk));
	jand g10616(.dina(w_n10852_0[1]),.dinb(w_n8890_35[1]),.dout(n10854),.clk(gclk));
	jxor g10617(.dina(w_n10332_0[0]),.dinb(w_n9369_29[1]),.dout(n10855),.clk(gclk));
	jor g10618(.dina(n10855),.dinb(w_n10824_46[1]),.dout(n10856),.clk(gclk));
	jxor g10619(.dina(n10856),.dinb(w_n10340_0[0]),.dout(n10857),.clk(gclk));
	jor g10620(.dina(w_n10857_0[2]),.dinb(n10854),.dout(n10858),.clk(gclk));
	jand g10621(.dina(n10858),.dinb(w_n10853_0[1]),.dout(n10859),.clk(gclk));
	jor g10622(.dina(w_n10859_0[2]),.dinb(w_n8449_30[2]),.dout(n10860),.clk(gclk));
	jand g10623(.dina(w_n10859_0[1]),.dinb(w_n8449_30[1]),.dout(n10861),.clk(gclk));
	jxor g10624(.dina(w_n10342_0[0]),.dinb(w_n8890_35[0]),.dout(n10862),.clk(gclk));
	jor g10625(.dina(n10862),.dinb(w_n10824_46[0]),.dout(n10863),.clk(gclk));
	jxor g10626(.dina(n10863),.dinb(w_n10664_0[0]),.dout(n10864),.clk(gclk));
	jnot g10627(.din(w_n10864_0[2]),.dout(n10865),.clk(gclk));
	jor g10628(.dina(n10865),.dinb(n10861),.dout(n10866),.clk(gclk));
	jand g10629(.dina(n10866),.dinb(w_n10860_0[1]),.dout(n10867),.clk(gclk));
	jor g10630(.dina(w_n10867_0[2]),.dinb(w_n8003_36[1]),.dout(n10868),.clk(gclk));
	jand g10631(.dina(w_n10867_0[1]),.dinb(w_n8003_36[0]),.dout(n10869),.clk(gclk));
	jxor g10632(.dina(w_n10349_0[0]),.dinb(w_n8449_30[0]),.dout(n10870),.clk(gclk));
	jor g10633(.dina(n10870),.dinb(w_n10824_45[2]),.dout(n10871),.clk(gclk));
	jxor g10634(.dina(n10871),.dinb(w_n10355_0[0]),.dout(n10872),.clk(gclk));
	jor g10635(.dina(w_n10872_0[2]),.dinb(n10869),.dout(n10873),.clk(gclk));
	jand g10636(.dina(n10873),.dinb(w_n10868_0[1]),.dout(n10874),.clk(gclk));
	jor g10637(.dina(w_n10874_0[2]),.dinb(w_n7581_31[2]),.dout(n10875),.clk(gclk));
	jand g10638(.dina(w_n10874_0[1]),.dinb(w_n7581_31[1]),.dout(n10876),.clk(gclk));
	jxor g10639(.dina(w_n10357_0[0]),.dinb(w_n8003_35[2]),.dout(n10877),.clk(gclk));
	jor g10640(.dina(n10877),.dinb(w_n10824_45[1]),.dout(n10878),.clk(gclk));
	jxor g10641(.dina(n10878),.dinb(w_n10671_0[0]),.dout(n10879),.clk(gclk));
	jnot g10642(.din(w_n10879_0[2]),.dout(n10880),.clk(gclk));
	jor g10643(.dina(n10880),.dinb(n10876),.dout(n10881),.clk(gclk));
	jand g10644(.dina(n10881),.dinb(w_n10875_0[1]),.dout(n10882),.clk(gclk));
	jor g10645(.dina(w_n10882_0[2]),.dinb(w_n7154_36[2]),.dout(n10883),.clk(gclk));
	jand g10646(.dina(w_n10882_0[1]),.dinb(w_n7154_36[1]),.dout(n10884),.clk(gclk));
	jxor g10647(.dina(w_n10364_0[0]),.dinb(w_n7581_31[0]),.dout(n10885),.clk(gclk));
	jor g10648(.dina(n10885),.dinb(w_n10824_45[0]),.dout(n10886),.clk(gclk));
	jxor g10649(.dina(n10886),.dinb(w_n10370_0[0]),.dout(n10887),.clk(gclk));
	jor g10650(.dina(w_n10887_0[2]),.dinb(n10884),.dout(n10888),.clk(gclk));
	jand g10651(.dina(n10888),.dinb(w_n10883_0[1]),.dout(n10889),.clk(gclk));
	jor g10652(.dina(w_n10889_0[2]),.dinb(w_n6758_32[1]),.dout(n10890),.clk(gclk));
	jand g10653(.dina(w_n10889_0[1]),.dinb(w_n6758_32[0]),.dout(n10891),.clk(gclk));
	jxor g10654(.dina(w_n10372_0[0]),.dinb(w_n7154_36[0]),.dout(n10892),.clk(gclk));
	jor g10655(.dina(n10892),.dinb(w_n10824_44[2]),.dout(n10893),.clk(gclk));
	jxor g10656(.dina(n10893),.dinb(w_n10378_0[0]),.dout(n10894),.clk(gclk));
	jor g10657(.dina(w_n10894_0[2]),.dinb(n10891),.dout(n10895),.clk(gclk));
	jand g10658(.dina(n10895),.dinb(w_n10890_0[1]),.dout(n10896),.clk(gclk));
	jor g10659(.dina(w_n10896_0[2]),.dinb(w_n6357_37[0]),.dout(n10897),.clk(gclk));
	jand g10660(.dina(w_n10896_0[1]),.dinb(w_n6357_36[2]),.dout(n10898),.clk(gclk));
	jxor g10661(.dina(w_n10380_0[0]),.dinb(w_n6758_31[2]),.dout(n10899),.clk(gclk));
	jor g10662(.dina(n10899),.dinb(w_n10824_44[1]),.dout(n10900),.clk(gclk));
	jxor g10663(.dina(n10900),.dinb(w_n10386_0[0]),.dout(n10901),.clk(gclk));
	jor g10664(.dina(w_n10901_0[2]),.dinb(n10898),.dout(n10902),.clk(gclk));
	jand g10665(.dina(n10902),.dinb(w_n10897_0[1]),.dout(n10903),.clk(gclk));
	jor g10666(.dina(w_n10903_0[2]),.dinb(w_n5989_33[0]),.dout(n10904),.clk(gclk));
	jand g10667(.dina(w_n10903_0[1]),.dinb(w_n5989_32[2]),.dout(n10905),.clk(gclk));
	jxor g10668(.dina(w_n10388_0[0]),.dinb(w_n6357_36[1]),.dout(n10906),.clk(gclk));
	jor g10669(.dina(n10906),.dinb(w_n10824_44[0]),.dout(n10907),.clk(gclk));
	jxor g10670(.dina(n10907),.dinb(w_n10684_0[0]),.dout(n10908),.clk(gclk));
	jnot g10671(.din(w_n10908_0[2]),.dout(n10909),.clk(gclk));
	jor g10672(.dina(n10909),.dinb(n10905),.dout(n10910),.clk(gclk));
	jand g10673(.dina(n10910),.dinb(w_n10904_0[1]),.dout(n10911),.clk(gclk));
	jor g10674(.dina(w_n10911_0[2]),.dinb(w_n5606_37[1]),.dout(n10912),.clk(gclk));
	jand g10675(.dina(w_n10911_0[1]),.dinb(w_n5606_37[0]),.dout(n10913),.clk(gclk));
	jxor g10676(.dina(w_n10395_0[0]),.dinb(w_n5989_32[1]),.dout(n10914),.clk(gclk));
	jor g10677(.dina(n10914),.dinb(w_n10824_43[2]),.dout(n10915),.clk(gclk));
	jxor g10678(.dina(n10915),.dinb(w_n10401_0[0]),.dout(n10916),.clk(gclk));
	jor g10679(.dina(w_n10916_0[2]),.dinb(n10913),.dout(n10917),.clk(gclk));
	jand g10680(.dina(n10917),.dinb(w_n10912_0[1]),.dout(n10918),.clk(gclk));
	jor g10681(.dina(w_n10918_0[2]),.dinb(w_n5259_34[0]),.dout(n10919),.clk(gclk));
	jand g10682(.dina(w_n10918_0[1]),.dinb(w_n5259_33[2]),.dout(n10920),.clk(gclk));
	jxor g10683(.dina(w_n10403_0[0]),.dinb(w_n5606_36[2]),.dout(n10921),.clk(gclk));
	jor g10684(.dina(n10921),.dinb(w_n10824_43[1]),.dout(n10922),.clk(gclk));
	jxor g10685(.dina(n10922),.dinb(w_n10409_0[0]),.dout(n10923),.clk(gclk));
	jor g10686(.dina(w_n10923_0[2]),.dinb(n10920),.dout(n10924),.clk(gclk));
	jand g10687(.dina(n10924),.dinb(w_n10919_0[1]),.dout(n10925),.clk(gclk));
	jor g10688(.dina(w_n10925_0[2]),.dinb(w_n4902_38[0]),.dout(n10926),.clk(gclk));
	jand g10689(.dina(w_n10925_0[1]),.dinb(w_n4902_37[2]),.dout(n10927),.clk(gclk));
	jxor g10690(.dina(w_n10411_0[0]),.dinb(w_n5259_33[1]),.dout(n10928),.clk(gclk));
	jor g10691(.dina(n10928),.dinb(w_n10824_43[0]),.dout(n10929),.clk(gclk));
	jxor g10692(.dina(n10929),.dinb(w_n10417_0[0]),.dout(n10930),.clk(gclk));
	jor g10693(.dina(w_n10930_0[2]),.dinb(n10927),.dout(n10931),.clk(gclk));
	jand g10694(.dina(n10931),.dinb(w_n10926_0[1]),.dout(n10932),.clk(gclk));
	jor g10695(.dina(w_n10932_0[2]),.dinb(w_n4582_35[0]),.dout(n10933),.clk(gclk));
	jand g10696(.dina(w_n10932_0[1]),.dinb(w_n4582_34[2]),.dout(n10934),.clk(gclk));
	jxor g10697(.dina(w_n10419_0[0]),.dinb(w_n4902_37[1]),.dout(n10935),.clk(gclk));
	jor g10698(.dina(n10935),.dinb(w_n10824_42[2]),.dout(n10936),.clk(gclk));
	jxor g10699(.dina(n10936),.dinb(w_n10425_0[0]),.dout(n10937),.clk(gclk));
	jor g10700(.dina(w_n10937_0[2]),.dinb(n10934),.dout(n10938),.clk(gclk));
	jand g10701(.dina(n10938),.dinb(w_n10933_0[1]),.dout(n10939),.clk(gclk));
	jor g10702(.dina(w_n10939_0[2]),.dinb(w_n4249_38[2]),.dout(n10940),.clk(gclk));
	jand g10703(.dina(w_n10939_0[1]),.dinb(w_n4249_38[1]),.dout(n10941),.clk(gclk));
	jxor g10704(.dina(w_n10427_0[0]),.dinb(w_n4582_34[1]),.dout(n10942),.clk(gclk));
	jor g10705(.dina(n10942),.dinb(w_n10824_42[1]),.dout(n10943),.clk(gclk));
	jxor g10706(.dina(n10943),.dinb(w_n10433_0[0]),.dout(n10944),.clk(gclk));
	jor g10707(.dina(w_n10944_0[2]),.dinb(n10941),.dout(n10945),.clk(gclk));
	jand g10708(.dina(n10945),.dinb(w_n10940_0[1]),.dout(n10946),.clk(gclk));
	jor g10709(.dina(w_n10946_0[2]),.dinb(w_n3955_35[2]),.dout(n10947),.clk(gclk));
	jxor g10710(.dina(w_n10435_0[0]),.dinb(w_n4249_38[0]),.dout(n10948),.clk(gclk));
	jor g10711(.dina(n10948),.dinb(w_n10824_42[0]),.dout(n10949),.clk(gclk));
	jxor g10712(.dina(n10949),.dinb(w_n10635_0[0]),.dout(n10950),.clk(gclk));
	jnot g10713(.din(w_n10950_0[2]),.dout(n10951),.clk(gclk));
	jand g10714(.dina(w_n10946_0[1]),.dinb(w_n3955_35[1]),.dout(n10952),.clk(gclk));
	jor g10715(.dina(n10952),.dinb(n10951),.dout(n10953),.clk(gclk));
	jand g10716(.dina(n10953),.dinb(w_n10947_0[1]),.dout(n10954),.clk(gclk));
	jor g10717(.dina(w_n10954_0[2]),.dinb(w_n3642_39[0]),.dout(n10955),.clk(gclk));
	jand g10718(.dina(w_n10954_0[1]),.dinb(w_n3642_38[2]),.dout(n10956),.clk(gclk));
	jxor g10719(.dina(w_n10442_0[0]),.dinb(w_n3955_35[0]),.dout(n10957),.clk(gclk));
	jor g10720(.dina(n10957),.dinb(w_n10824_41[2]),.dout(n10958),.clk(gclk));
	jxor g10721(.dina(n10958),.dinb(w_n10448_0[0]),.dout(n10959),.clk(gclk));
	jor g10722(.dina(w_n10959_0[2]),.dinb(n10956),.dout(n10960),.clk(gclk));
	jand g10723(.dina(n10960),.dinb(w_n10955_0[1]),.dout(n10961),.clk(gclk));
	jor g10724(.dina(w_n10961_0[2]),.dinb(w_n3368_36[1]),.dout(n10962),.clk(gclk));
	jand g10725(.dina(w_n10961_0[1]),.dinb(w_n3368_36[0]),.dout(n10963),.clk(gclk));
	jxor g10726(.dina(w_n10450_0[0]),.dinb(w_n3642_38[1]),.dout(n10964),.clk(gclk));
	jor g10727(.dina(n10964),.dinb(w_n10824_41[1]),.dout(n10965),.clk(gclk));
	jxor g10728(.dina(n10965),.dinb(w_n10709_0[0]),.dout(n10966),.clk(gclk));
	jnot g10729(.din(w_n10966_0[2]),.dout(n10967),.clk(gclk));
	jor g10730(.dina(n10967),.dinb(n10963),.dout(n10968),.clk(gclk));
	jand g10731(.dina(n10968),.dinb(w_n10962_0[1]),.dout(n10969),.clk(gclk));
	jor g10732(.dina(w_n10969_0[2]),.dinb(w_n3089_39[2]),.dout(n10970),.clk(gclk));
	jand g10733(.dina(w_n10969_0[1]),.dinb(w_n3089_39[1]),.dout(n10971),.clk(gclk));
	jxor g10734(.dina(w_n10457_0[0]),.dinb(w_n3368_35[2]),.dout(n10972),.clk(gclk));
	jor g10735(.dina(n10972),.dinb(w_n10824_41[0]),.dout(n10973),.clk(gclk));
	jxor g10736(.dina(n10973),.dinb(w_n10463_0[0]),.dout(n10974),.clk(gclk));
	jor g10737(.dina(w_n10974_0[2]),.dinb(n10971),.dout(n10975),.clk(gclk));
	jand g10738(.dina(n10975),.dinb(w_n10970_0[1]),.dout(n10976),.clk(gclk));
	jor g10739(.dina(w_n10976_0[2]),.dinb(w_n2833_37[1]),.dout(n10977),.clk(gclk));
	jand g10740(.dina(w_n10976_0[1]),.dinb(w_n2833_37[0]),.dout(n10978),.clk(gclk));
	jxor g10741(.dina(w_n10465_0[0]),.dinb(w_n3089_39[0]),.dout(n10979),.clk(gclk));
	jor g10742(.dina(n10979),.dinb(w_n10824_40[2]),.dout(n10980),.clk(gclk));
	jxor g10743(.dina(n10980),.dinb(w_n10716_0[0]),.dout(n10981),.clk(gclk));
	jnot g10744(.din(w_n10981_0[2]),.dout(n10982),.clk(gclk));
	jor g10745(.dina(n10982),.dinb(n10978),.dout(n10983),.clk(gclk));
	jand g10746(.dina(n10983),.dinb(w_n10977_0[1]),.dout(n10984),.clk(gclk));
	jor g10747(.dina(w_n10984_0[2]),.dinb(w_n2572_40[0]),.dout(n10985),.clk(gclk));
	jand g10748(.dina(w_n10984_0[1]),.dinb(w_n2572_39[2]),.dout(n10986),.clk(gclk));
	jxor g10749(.dina(w_n10472_0[0]),.dinb(w_n2833_36[2]),.dout(n10987),.clk(gclk));
	jor g10750(.dina(n10987),.dinb(w_n10824_40[1]),.dout(n10988),.clk(gclk));
	jxor g10751(.dina(n10988),.dinb(w_n10478_0[0]),.dout(n10989),.clk(gclk));
	jor g10752(.dina(w_n10989_0[2]),.dinb(n10986),.dout(n10990),.clk(gclk));
	jand g10753(.dina(n10990),.dinb(w_n10985_0[1]),.dout(n10991),.clk(gclk));
	jor g10754(.dina(w_n10991_0[2]),.dinb(w_n2345_38[0]),.dout(n10992),.clk(gclk));
	jand g10755(.dina(w_n10991_0[1]),.dinb(w_n2345_37[2]),.dout(n10993),.clk(gclk));
	jxor g10756(.dina(w_n10480_0[0]),.dinb(w_n2572_39[1]),.dout(n10994),.clk(gclk));
	jor g10757(.dina(n10994),.dinb(w_n10824_40[0]),.dout(n10995),.clk(gclk));
	jxor g10758(.dina(n10995),.dinb(w_n10486_0[0]),.dout(n10996),.clk(gclk));
	jor g10759(.dina(w_n10996_0[2]),.dinb(n10993),.dout(n10997),.clk(gclk));
	jand g10760(.dina(n10997),.dinb(w_n10992_0[1]),.dout(n10998),.clk(gclk));
	jor g10761(.dina(w_n10998_0[2]),.dinb(w_n2108_40[2]),.dout(n10999),.clk(gclk));
	jand g10762(.dina(w_n10998_0[1]),.dinb(w_n2108_40[1]),.dout(n11000),.clk(gclk));
	jxor g10763(.dina(w_n10488_0[0]),.dinb(w_n2345_37[1]),.dout(n11001),.clk(gclk));
	jor g10764(.dina(n11001),.dinb(w_n10824_39[2]),.dout(n11002),.clk(gclk));
	jxor g10765(.dina(n11002),.dinb(w_n10494_0[0]),.dout(n11003),.clk(gclk));
	jor g10766(.dina(w_n11003_0[2]),.dinb(n11000),.dout(n11004),.clk(gclk));
	jand g10767(.dina(n11004),.dinb(w_n10999_0[1]),.dout(n11005),.clk(gclk));
	jor g10768(.dina(w_n11005_0[2]),.dinb(w_n1912_39[0]),.dout(n11006),.clk(gclk));
	jand g10769(.dina(w_n11005_0[1]),.dinb(w_n1912_38[2]),.dout(n11007),.clk(gclk));
	jxor g10770(.dina(w_n10496_0[0]),.dinb(w_n2108_40[0]),.dout(n11008),.clk(gclk));
	jor g10771(.dina(n11008),.dinb(w_n10824_39[1]),.dout(n11009),.clk(gclk));
	jxor g10772(.dina(n11009),.dinb(w_n10729_0[0]),.dout(n11010),.clk(gclk));
	jnot g10773(.din(w_n11010_0[2]),.dout(n11011),.clk(gclk));
	jor g10774(.dina(n11011),.dinb(n11007),.dout(n11012),.clk(gclk));
	jand g10775(.dina(n11012),.dinb(w_n11006_0[1]),.dout(n11013),.clk(gclk));
	jor g10776(.dina(w_n11013_0[2]),.dinb(w_n1699_41[1]),.dout(n11014),.clk(gclk));
	jand g10777(.dina(w_n11013_0[1]),.dinb(w_n1699_41[0]),.dout(n11015),.clk(gclk));
	jxor g10778(.dina(w_n10503_0[0]),.dinb(w_n1912_38[1]),.dout(n11016),.clk(gclk));
	jor g10779(.dina(n11016),.dinb(w_n10824_39[0]),.dout(n11017),.clk(gclk));
	jxor g10780(.dina(n11017),.dinb(w_n10509_0[0]),.dout(n11018),.clk(gclk));
	jor g10781(.dina(w_n11018_0[2]),.dinb(n11015),.dout(n11019),.clk(gclk));
	jand g10782(.dina(n11019),.dinb(w_n11014_0[1]),.dout(n11020),.clk(gclk));
	jor g10783(.dina(w_n11020_0[2]),.dinb(w_n1516_39[2]),.dout(n11021),.clk(gclk));
	jand g10784(.dina(w_n11020_0[1]),.dinb(w_n1516_39[1]),.dout(n11022),.clk(gclk));
	jxor g10785(.dina(w_n10511_0[0]),.dinb(w_n1699_40[2]),.dout(n11023),.clk(gclk));
	jor g10786(.dina(n11023),.dinb(w_n10824_38[2]),.dout(n11024),.clk(gclk));
	jxor g10787(.dina(n11024),.dinb(w_n10736_0[0]),.dout(n11025),.clk(gclk));
	jnot g10788(.din(w_n11025_0[2]),.dout(n11026),.clk(gclk));
	jor g10789(.dina(n11026),.dinb(n11022),.dout(n11027),.clk(gclk));
	jand g10790(.dina(n11027),.dinb(w_n11021_0[1]),.dout(n11028),.clk(gclk));
	jor g10791(.dina(w_n11028_0[2]),.dinb(w_n1332_41[1]),.dout(n11029),.clk(gclk));
	jand g10792(.dina(w_n11028_0[1]),.dinb(w_n1332_41[0]),.dout(n11030),.clk(gclk));
	jxor g10793(.dina(w_n10518_0[0]),.dinb(w_n1516_39[0]),.dout(n11031),.clk(gclk));
	jor g10794(.dina(n11031),.dinb(w_n10824_38[1]),.dout(n11032),.clk(gclk));
	jxor g10795(.dina(n11032),.dinb(w_n10524_0[0]),.dout(n11033),.clk(gclk));
	jor g10796(.dina(w_n11033_0[2]),.dinb(n11030),.dout(n11034),.clk(gclk));
	jand g10797(.dina(n11034),.dinb(w_n11029_0[1]),.dout(n11035),.clk(gclk));
	jor g10798(.dina(w_n11035_0[2]),.dinb(w_n1173_40[1]),.dout(n11036),.clk(gclk));
	jand g10799(.dina(w_n11035_0[1]),.dinb(w_n1173_40[0]),.dout(n11037),.clk(gclk));
	jxor g10800(.dina(w_n10526_0[0]),.dinb(w_n1332_40[2]),.dout(n11038),.clk(gclk));
	jor g10801(.dina(n11038),.dinb(w_n10824_38[0]),.dout(n11039),.clk(gclk));
	jxor g10802(.dina(n11039),.dinb(w_n10743_0[0]),.dout(n11040),.clk(gclk));
	jnot g10803(.din(w_n11040_0[2]),.dout(n11041),.clk(gclk));
	jor g10804(.dina(n11041),.dinb(n11037),.dout(n11042),.clk(gclk));
	jand g10805(.dina(n11042),.dinb(w_n11036_0[1]),.dout(n11043),.clk(gclk));
	jor g10806(.dina(w_n11043_0[2]),.dinb(w_n1008_42[1]),.dout(n11044),.clk(gclk));
	jand g10807(.dina(w_n11043_0[1]),.dinb(w_n1008_42[0]),.dout(n11045),.clk(gclk));
	jxor g10808(.dina(w_n10533_0[0]),.dinb(w_n1173_39[2]),.dout(n11046),.clk(gclk));
	jor g10809(.dina(n11046),.dinb(w_n10824_37[2]),.dout(n11047),.clk(gclk));
	jxor g10810(.dina(n11047),.dinb(w_n10539_0[0]),.dout(n11048),.clk(gclk));
	jor g10811(.dina(w_n11048_0[2]),.dinb(n11045),.dout(n11049),.clk(gclk));
	jand g10812(.dina(n11049),.dinb(w_n11044_0[1]),.dout(n11050),.clk(gclk));
	jor g10813(.dina(w_n11050_0[2]),.dinb(w_n884_41[1]),.dout(n11051),.clk(gclk));
	jand g10814(.dina(w_n11050_0[1]),.dinb(w_n884_41[0]),.dout(n11052),.clk(gclk));
	jxor g10815(.dina(w_n10541_0[0]),.dinb(w_n1008_41[2]),.dout(n11053),.clk(gclk));
	jor g10816(.dina(n11053),.dinb(w_n10824_37[1]),.dout(n11054),.clk(gclk));
	jxor g10817(.dina(n11054),.dinb(w_n10750_0[0]),.dout(n11055),.clk(gclk));
	jnot g10818(.din(w_n11055_0[2]),.dout(n11056),.clk(gclk));
	jor g10819(.dina(n11056),.dinb(n11052),.dout(n11057),.clk(gclk));
	jand g10820(.dina(n11057),.dinb(w_n11051_0[1]),.dout(n11058),.clk(gclk));
	jor g10821(.dina(w_n11058_0[2]),.dinb(w_n743_42[1]),.dout(n11059),.clk(gclk));
	jand g10822(.dina(w_n11058_0[1]),.dinb(w_n743_42[0]),.dout(n11060),.clk(gclk));
	jxor g10823(.dina(w_n10548_0[0]),.dinb(w_n884_40[2]),.dout(n11061),.clk(gclk));
	jor g10824(.dina(n11061),.dinb(w_n10824_37[0]),.dout(n11062),.clk(gclk));
	jxor g10825(.dina(n11062),.dinb(w_n10754_0[0]),.dout(n11063),.clk(gclk));
	jnot g10826(.din(w_n11063_0[2]),.dout(n11064),.clk(gclk));
	jor g10827(.dina(n11064),.dinb(n11060),.dout(n11065),.clk(gclk));
	jand g10828(.dina(n11065),.dinb(w_n11059_0[1]),.dout(n11066),.clk(gclk));
	jor g10829(.dina(w_n11066_0[2]),.dinb(w_n635_42[1]),.dout(n11067),.clk(gclk));
	jand g10830(.dina(w_n11066_0[1]),.dinb(w_n635_42[0]),.dout(n11068),.clk(gclk));
	jxor g10831(.dina(w_n10555_0[0]),.dinb(w_n743_41[2]),.dout(n11069),.clk(gclk));
	jor g10832(.dina(n11069),.dinb(w_n10824_36[2]),.dout(n11070),.clk(gclk));
	jxor g10833(.dina(n11070),.dinb(w_n10758_0[0]),.dout(n11071),.clk(gclk));
	jnot g10834(.din(w_n11071_0[2]),.dout(n11072),.clk(gclk));
	jor g10835(.dina(n11072),.dinb(n11068),.dout(n11073),.clk(gclk));
	jand g10836(.dina(n11073),.dinb(w_n11067_0[1]),.dout(n11074),.clk(gclk));
	jor g10837(.dina(w_n11074_0[2]),.dinb(w_n515_43[1]),.dout(n11075),.clk(gclk));
	jand g10838(.dina(w_n11074_0[1]),.dinb(w_n515_43[0]),.dout(n11076),.clk(gclk));
	jxor g10839(.dina(w_n10562_0[0]),.dinb(w_n635_41[2]),.dout(n11077),.clk(gclk));
	jor g10840(.dina(n11077),.dinb(w_n10824_36[1]),.dout(n11078),.clk(gclk));
	jxor g10841(.dina(n11078),.dinb(w_n10568_0[0]),.dout(n11079),.clk(gclk));
	jor g10842(.dina(w_n11079_0[2]),.dinb(n11076),.dout(n11080),.clk(gclk));
	jand g10843(.dina(n11080),.dinb(w_n11075_0[1]),.dout(n11081),.clk(gclk));
	jor g10844(.dina(w_n11081_0[2]),.dinb(w_n443_43[1]),.dout(n11082),.clk(gclk));
	jand g10845(.dina(w_n11081_0[1]),.dinb(w_n443_43[0]),.dout(n11083),.clk(gclk));
	jxor g10846(.dina(w_n10570_0[0]),.dinb(w_n515_42[2]),.dout(n11084),.clk(gclk));
	jor g10847(.dina(n11084),.dinb(w_n10824_36[0]),.dout(n11085),.clk(gclk));
	jxor g10848(.dina(n11085),.dinb(w_n10576_0[0]),.dout(n11086),.clk(gclk));
	jor g10849(.dina(w_n11086_0[2]),.dinb(n11083),.dout(n11087),.clk(gclk));
	jand g10850(.dina(n11087),.dinb(w_n11082_0[1]),.dout(n11088),.clk(gclk));
	jor g10851(.dina(w_n11088_0[2]),.dinb(w_n352_43[2]),.dout(n11089),.clk(gclk));
	jand g10852(.dina(w_n11088_0[1]),.dinb(w_n352_43[1]),.dout(n11090),.clk(gclk));
	jxor g10853(.dina(w_n10578_0[0]),.dinb(w_n443_42[2]),.dout(n11091),.clk(gclk));
	jor g10854(.dina(n11091),.dinb(w_n10824_35[2]),.dout(n11092),.clk(gclk));
	jxor g10855(.dina(n11092),.dinb(w_n10584_0[0]),.dout(n11093),.clk(gclk));
	jor g10856(.dina(w_n11093_0[2]),.dinb(n11090),.dout(n11094),.clk(gclk));
	jand g10857(.dina(n11094),.dinb(w_n11089_0[1]),.dout(n11095),.clk(gclk));
	jor g10858(.dina(w_n11095_0[2]),.dinb(w_n294_44[0]),.dout(n11096),.clk(gclk));
	jand g10859(.dina(w_n11095_0[1]),.dinb(w_n294_43[2]),.dout(n11097),.clk(gclk));
	jxor g10860(.dina(w_n10586_0[0]),.dinb(w_n352_43[0]),.dout(n11098),.clk(gclk));
	jor g10861(.dina(n11098),.dinb(w_n10824_35[1]),.dout(n11099),.clk(gclk));
	jxor g10862(.dina(n11099),.dinb(w_n10771_0[0]),.dout(n11100),.clk(gclk));
	jnot g10863(.din(w_n11100_0[2]),.dout(n11101),.clk(gclk));
	jor g10864(.dina(n11101),.dinb(n11097),.dout(n11102),.clk(gclk));
	jand g10865(.dina(n11102),.dinb(w_n11096_0[1]),.dout(n11103),.clk(gclk));
	jor g10866(.dina(w_n11103_0[2]),.dinb(w_n239_44[0]),.dout(n11104),.clk(gclk));
	jand g10867(.dina(w_n11103_0[1]),.dinb(w_n239_43[2]),.dout(n11105),.clk(gclk));
	jxor g10868(.dina(w_n10593_0[0]),.dinb(w_n294_43[1]),.dout(n11106),.clk(gclk));
	jor g10869(.dina(n11106),.dinb(w_n10824_35[0]),.dout(n11107),.clk(gclk));
	jxor g10870(.dina(n11107),.dinb(w_n10599_0[0]),.dout(n11108),.clk(gclk));
	jor g10871(.dina(w_n11108_0[2]),.dinb(n11105),.dout(n11109),.clk(gclk));
	jand g10872(.dina(n11109),.dinb(w_n11104_0[1]),.dout(n11110),.clk(gclk));
	jor g10873(.dina(w_n11110_0[2]),.dinb(w_n221_44[1]),.dout(n11111),.clk(gclk));
	jand g10874(.dina(w_n11110_0[1]),.dinb(w_n221_44[0]),.dout(n11112),.clk(gclk));
	jxor g10875(.dina(w_n10601_0[0]),.dinb(w_n239_43[1]),.dout(n11113),.clk(gclk));
	jor g10876(.dina(n11113),.dinb(w_n10824_34[2]),.dout(n11114),.clk(gclk));
	jxor g10877(.dina(n11114),.dinb(w_n10607_0[0]),.dout(n11115),.clk(gclk));
	jor g10878(.dina(w_n11115_0[1]),.dinb(n11112),.dout(n11116),.clk(gclk));
	jand g10879(.dina(n11116),.dinb(w_n11111_0[1]),.dout(n11117),.clk(gclk));
	jxor g10880(.dina(w_n10609_0[0]),.dinb(w_n221_43[2]),.dout(n11118),.clk(gclk));
	jor g10881(.dina(n11118),.dinb(w_n10824_34[1]),.dout(n11119),.clk(gclk));
	jxor g10882(.dina(n11119),.dinb(w_n10811_0[0]),.dout(n11120),.clk(gclk));
	jand g10883(.dina(w_n11120_1[1]),.dinb(w_n11117_1[1]),.dout(n11121),.clk(gclk));
	jand g10884(.dina(w_n10824_34[0]),.dinb(w_n10785_0[0]),.dout(n11122),.clk(gclk));
	jand g10885(.dina(w_n10789_0[0]),.dinb(w_asqrt63_32[2]),.dout(n11123),.clk(gclk));
	jand g10886(.dina(n11123),.dinb(w_n10820_0[1]),.dout(n11124),.clk(gclk));
	jnot g10887(.din(n11124),.dout(n11125),.clk(gclk));
	jor g10888(.dina(w_n11125_0[1]),.dinb(n11122),.dout(n11126),.clk(gclk));
	jnot g10889(.din(w_n11126_0[1]),.dout(n11127),.clk(gclk));
	jand g10890(.dina(w_asqrt23_17[2]),.dinb(w_n10815_0[0]),.dout(n11128),.clk(gclk));
	jor g10891(.dina(w_n11120_1[0]),.dinb(w_n11117_1[0]),.dout(n11129),.clk(gclk));
	jor g10892(.dina(n11129),.dinb(w_n10795_0[0]),.dout(n11130),.clk(gclk));
	jor g10893(.dina(n11130),.dinb(w_n11128_0[1]),.dout(n11131),.clk(gclk));
	jand g10894(.dina(n11131),.dinb(w_n218_18[1]),.dout(n11132),.clk(gclk));
	jand g10895(.dina(w_n10824_33[2]),.dinb(w_n10788_0[1]),.dout(n11133),.clk(gclk));
	jor g10896(.dina(w_n11133_0[1]),.dinb(n11132),.dout(n11134),.clk(gclk));
	jor g10897(.dina(n11134),.dinb(n11127),.dout(n11135),.clk(gclk));
	jor g10898(.dina(n11135),.dinb(w_n11121_0[1]),.dout(asqrt_fa_23),.clk(gclk));
	jnot g10899(.din(w_n11115_0[0]),.dout(n11137),.clk(gclk));
	jxor g10900(.dina(w_n11110_0[0]),.dinb(w_n221_43[1]),.dout(n11138),.clk(gclk));
	jand g10901(.dina(n11138),.dinb(w_asqrt22_36),.dout(n11139),.clk(gclk));
	jxor g10902(.dina(n11139),.dinb(w_n11137_0[1]),.dout(n11140),.clk(gclk));
	jand g10903(.dina(w_asqrt22_35[2]),.dinb(w_a44_0[1]),.dout(n11141),.clk(gclk));
	jnot g10904(.din(w_a42_1[1]),.dout(n11142),.clk(gclk));
	jnot g10905(.din(w_a43_0[1]),.dout(n11143),.clk(gclk));
	jand g10906(.dina(w_n11143_0[1]),.dinb(w_n11142_1[1]),.dout(n11144),.clk(gclk));
	jand g10907(.dina(w_n11144_0[2]),.dinb(w_n10805_1[1]),.dout(n11145),.clk(gclk));
	jor g10908(.dina(w_n11145_0[1]),.dinb(n11141),.dout(n11146),.clk(gclk));
	jand g10909(.dina(w_n11146_0[2]),.dinb(w_asqrt23_17[1]),.dout(n11147),.clk(gclk));
	jor g10910(.dina(w_n11146_0[1]),.dinb(w_asqrt23_17[0]),.dout(n11148),.clk(gclk));
	jand g10911(.dina(w_asqrt22_35[1]),.dinb(w_n10805_1[0]),.dout(n11149),.clk(gclk));
	jor g10912(.dina(n11149),.dinb(w_n10806_0[0]),.dout(n11150),.clk(gclk));
	jnot g10913(.din(w_n10807_0[1]),.dout(n11151),.clk(gclk));
	jnot g10914(.din(w_n11121_0[0]),.dout(n11152),.clk(gclk));
	jnot g10915(.din(w_n11128_0[0]),.dout(n11153),.clk(gclk));
	jnot g10916(.din(w_n11111_0[0]),.dout(n11154),.clk(gclk));
	jnot g10917(.din(w_n11104_0[0]),.dout(n11155),.clk(gclk));
	jnot g10918(.din(w_n11096_0[0]),.dout(n11156),.clk(gclk));
	jnot g10919(.din(w_n11089_0[0]),.dout(n11157),.clk(gclk));
	jnot g10920(.din(w_n11082_0[0]),.dout(n11158),.clk(gclk));
	jnot g10921(.din(w_n11075_0[0]),.dout(n11159),.clk(gclk));
	jnot g10922(.din(w_n11067_0[0]),.dout(n11160),.clk(gclk));
	jnot g10923(.din(w_n11059_0[0]),.dout(n11161),.clk(gclk));
	jnot g10924(.din(w_n11051_0[0]),.dout(n11162),.clk(gclk));
	jnot g10925(.din(w_n11044_0[0]),.dout(n11163),.clk(gclk));
	jnot g10926(.din(w_n11036_0[0]),.dout(n11164),.clk(gclk));
	jnot g10927(.din(w_n11029_0[0]),.dout(n11165),.clk(gclk));
	jnot g10928(.din(w_n11021_0[0]),.dout(n11166),.clk(gclk));
	jnot g10929(.din(w_n11014_0[0]),.dout(n11167),.clk(gclk));
	jnot g10930(.din(w_n11006_0[0]),.dout(n11168),.clk(gclk));
	jnot g10931(.din(w_n10999_0[0]),.dout(n11169),.clk(gclk));
	jnot g10932(.din(w_n10992_0[0]),.dout(n11170),.clk(gclk));
	jnot g10933(.din(w_n10985_0[0]),.dout(n11171),.clk(gclk));
	jnot g10934(.din(w_n10977_0[0]),.dout(n11172),.clk(gclk));
	jnot g10935(.din(w_n10970_0[0]),.dout(n11173),.clk(gclk));
	jnot g10936(.din(w_n10962_0[0]),.dout(n11174),.clk(gclk));
	jnot g10937(.din(w_n10955_0[0]),.dout(n11175),.clk(gclk));
	jnot g10938(.din(w_n10947_0[0]),.dout(n11176),.clk(gclk));
	jnot g10939(.din(w_n10940_0[0]),.dout(n11177),.clk(gclk));
	jnot g10940(.din(w_n10933_0[0]),.dout(n11178),.clk(gclk));
	jnot g10941(.din(w_n10926_0[0]),.dout(n11179),.clk(gclk));
	jnot g10942(.din(w_n10919_0[0]),.dout(n11180),.clk(gclk));
	jnot g10943(.din(w_n10912_0[0]),.dout(n11181),.clk(gclk));
	jnot g10944(.din(w_n10904_0[0]),.dout(n11182),.clk(gclk));
	jnot g10945(.din(w_n10897_0[0]),.dout(n11183),.clk(gclk));
	jnot g10946(.din(w_n10890_0[0]),.dout(n11184),.clk(gclk));
	jnot g10947(.din(w_n10883_0[0]),.dout(n11185),.clk(gclk));
	jnot g10948(.din(w_n10875_0[0]),.dout(n11186),.clk(gclk));
	jnot g10949(.din(w_n10868_0[0]),.dout(n11187),.clk(gclk));
	jnot g10950(.din(w_n10860_0[0]),.dout(n11188),.clk(gclk));
	jnot g10951(.din(w_n10853_0[0]),.dout(n11189),.clk(gclk));
	jnot g10952(.din(w_n10846_0[0]),.dout(n11190),.clk(gclk));
	jnot g10953(.din(w_n10835_0[0]),.dout(n11191),.clk(gclk));
	jnot g10954(.din(w_n10827_0[0]),.dout(n11192),.clk(gclk));
	jand g10955(.dina(w_asqrt23_16[2]),.dinb(w_a46_0[2]),.dout(n11193),.clk(gclk));
	jor g10956(.dina(n11193),.dinb(w_n10808_0[0]),.dout(n11194),.clk(gclk));
	jor g10957(.dina(n11194),.dinb(w_asqrt24_22[2]),.dout(n11195),.clk(gclk));
	jand g10958(.dina(w_asqrt23_16[1]),.dinb(w_n10134_0[1]),.dout(n11196),.clk(gclk));
	jor g10959(.dina(n11196),.dinb(w_n10135_0[0]),.dout(n11197),.clk(gclk));
	jand g10960(.dina(w_n10838_0[0]),.dinb(n11197),.dout(n11198),.clk(gclk));
	jand g10961(.dina(w_n11198_0[1]),.dinb(n11195),.dout(n11199),.clk(gclk));
	jor g10962(.dina(n11199),.dinb(n11192),.dout(n11200),.clk(gclk));
	jor g10963(.dina(n11200),.dinb(w_asqrt25_16[2]),.dout(n11201),.clk(gclk));
	jnot g10964(.din(w_n10843_0[1]),.dout(n11202),.clk(gclk));
	jand g10965(.dina(n11202),.dinb(n11201),.dout(n11203),.clk(gclk));
	jor g10966(.dina(n11203),.dinb(n11191),.dout(n11204),.clk(gclk));
	jor g10967(.dina(n11204),.dinb(w_asqrt26_22[2]),.dout(n11205),.clk(gclk));
	jnot g10968(.din(w_n10850_0[1]),.dout(n11206),.clk(gclk));
	jand g10969(.dina(n11206),.dinb(n11205),.dout(n11207),.clk(gclk));
	jor g10970(.dina(n11207),.dinb(n11190),.dout(n11208),.clk(gclk));
	jor g10971(.dina(n11208),.dinb(w_asqrt27_17[1]),.dout(n11209),.clk(gclk));
	jnot g10972(.din(w_n10857_0[1]),.dout(n11210),.clk(gclk));
	jand g10973(.dina(n11210),.dinb(n11209),.dout(n11211),.clk(gclk));
	jor g10974(.dina(n11211),.dinb(n11189),.dout(n11212),.clk(gclk));
	jor g10975(.dina(n11212),.dinb(w_asqrt28_23[0]),.dout(n11213),.clk(gclk));
	jand g10976(.dina(w_n10864_0[1]),.dinb(n11213),.dout(n11214),.clk(gclk));
	jor g10977(.dina(n11214),.dinb(n11188),.dout(n11215),.clk(gclk));
	jor g10978(.dina(n11215),.dinb(w_asqrt29_17[2]),.dout(n11216),.clk(gclk));
	jnot g10979(.din(w_n10872_0[1]),.dout(n11217),.clk(gclk));
	jand g10980(.dina(n11217),.dinb(n11216),.dout(n11218),.clk(gclk));
	jor g10981(.dina(n11218),.dinb(n11187),.dout(n11219),.clk(gclk));
	jor g10982(.dina(n11219),.dinb(w_asqrt30_23[1]),.dout(n11220),.clk(gclk));
	jand g10983(.dina(w_n10879_0[1]),.dinb(n11220),.dout(n11221),.clk(gclk));
	jor g10984(.dina(n11221),.dinb(n11186),.dout(n11222),.clk(gclk));
	jor g10985(.dina(n11222),.dinb(w_asqrt31_18[1]),.dout(n11223),.clk(gclk));
	jnot g10986(.din(w_n10887_0[1]),.dout(n11224),.clk(gclk));
	jand g10987(.dina(n11224),.dinb(n11223),.dout(n11225),.clk(gclk));
	jor g10988(.dina(n11225),.dinb(n11185),.dout(n11226),.clk(gclk));
	jor g10989(.dina(n11226),.dinb(w_asqrt32_23[1]),.dout(n11227),.clk(gclk));
	jnot g10990(.din(w_n10894_0[1]),.dout(n11228),.clk(gclk));
	jand g10991(.dina(n11228),.dinb(n11227),.dout(n11229),.clk(gclk));
	jor g10992(.dina(n11229),.dinb(n11184),.dout(n11230),.clk(gclk));
	jor g10993(.dina(n11230),.dinb(w_asqrt33_19[0]),.dout(n11231),.clk(gclk));
	jnot g10994(.din(w_n10901_0[1]),.dout(n11232),.clk(gclk));
	jand g10995(.dina(n11232),.dinb(n11231),.dout(n11233),.clk(gclk));
	jor g10996(.dina(n11233),.dinb(n11183),.dout(n11234),.clk(gclk));
	jor g10997(.dina(n11234),.dinb(w_asqrt34_23[2]),.dout(n11235),.clk(gclk));
	jand g10998(.dina(w_n10908_0[1]),.dinb(n11235),.dout(n11236),.clk(gclk));
	jor g10999(.dina(n11236),.dinb(n11182),.dout(n11237),.clk(gclk));
	jor g11000(.dina(n11237),.dinb(w_asqrt35_19[2]),.dout(n11238),.clk(gclk));
	jnot g11001(.din(w_n10916_0[1]),.dout(n11239),.clk(gclk));
	jand g11002(.dina(n11239),.dinb(n11238),.dout(n11240),.clk(gclk));
	jor g11003(.dina(n11240),.dinb(n11181),.dout(n11241),.clk(gclk));
	jor g11004(.dina(n11241),.dinb(w_asqrt36_23[2]),.dout(n11242),.clk(gclk));
	jnot g11005(.din(w_n10923_0[1]),.dout(n11243),.clk(gclk));
	jand g11006(.dina(n11243),.dinb(n11242),.dout(n11244),.clk(gclk));
	jor g11007(.dina(n11244),.dinb(n11180),.dout(n11245),.clk(gclk));
	jor g11008(.dina(n11245),.dinb(w_asqrt37_20[0]),.dout(n11246),.clk(gclk));
	jnot g11009(.din(w_n10930_0[1]),.dout(n11247),.clk(gclk));
	jand g11010(.dina(n11247),.dinb(n11246),.dout(n11248),.clk(gclk));
	jor g11011(.dina(n11248),.dinb(n11179),.dout(n11249),.clk(gclk));
	jor g11012(.dina(n11249),.dinb(w_asqrt38_24[0]),.dout(n11250),.clk(gclk));
	jnot g11013(.din(w_n10937_0[1]),.dout(n11251),.clk(gclk));
	jand g11014(.dina(n11251),.dinb(n11250),.dout(n11252),.clk(gclk));
	jor g11015(.dina(n11252),.dinb(n11178),.dout(n11253),.clk(gclk));
	jor g11016(.dina(n11253),.dinb(w_asqrt39_20[2]),.dout(n11254),.clk(gclk));
	jnot g11017(.din(w_n10944_0[1]),.dout(n11255),.clk(gclk));
	jand g11018(.dina(n11255),.dinb(n11254),.dout(n11256),.clk(gclk));
	jor g11019(.dina(n11256),.dinb(n11177),.dout(n11257),.clk(gclk));
	jor g11020(.dina(n11257),.dinb(w_asqrt40_24[0]),.dout(n11258),.clk(gclk));
	jand g11021(.dina(n11258),.dinb(w_n10950_0[1]),.dout(n11259),.clk(gclk));
	jor g11022(.dina(n11259),.dinb(n11176),.dout(n11260),.clk(gclk));
	jor g11023(.dina(n11260),.dinb(w_asqrt41_21[0]),.dout(n11261),.clk(gclk));
	jnot g11024(.din(w_n10959_0[1]),.dout(n11262),.clk(gclk));
	jand g11025(.dina(n11262),.dinb(n11261),.dout(n11263),.clk(gclk));
	jor g11026(.dina(n11263),.dinb(n11175),.dout(n11264),.clk(gclk));
	jor g11027(.dina(n11264),.dinb(w_asqrt42_24[1]),.dout(n11265),.clk(gclk));
	jand g11028(.dina(w_n10966_0[1]),.dinb(n11265),.dout(n11266),.clk(gclk));
	jor g11029(.dina(n11266),.dinb(n11174),.dout(n11267),.clk(gclk));
	jor g11030(.dina(n11267),.dinb(w_asqrt43_21[1]),.dout(n11268),.clk(gclk));
	jnot g11031(.din(w_n10974_0[1]),.dout(n11269),.clk(gclk));
	jand g11032(.dina(n11269),.dinb(n11268),.dout(n11270),.clk(gclk));
	jor g11033(.dina(n11270),.dinb(n11173),.dout(n11271),.clk(gclk));
	jor g11034(.dina(n11271),.dinb(w_asqrt44_24[1]),.dout(n11272),.clk(gclk));
	jand g11035(.dina(w_n10981_0[1]),.dinb(n11272),.dout(n11273),.clk(gclk));
	jor g11036(.dina(n11273),.dinb(n11172),.dout(n11274),.clk(gclk));
	jor g11037(.dina(n11274),.dinb(w_asqrt45_22[0]),.dout(n11275),.clk(gclk));
	jnot g11038(.din(w_n10989_0[1]),.dout(n11276),.clk(gclk));
	jand g11039(.dina(n11276),.dinb(n11275),.dout(n11277),.clk(gclk));
	jor g11040(.dina(n11277),.dinb(n11171),.dout(n11278),.clk(gclk));
	jor g11041(.dina(n11278),.dinb(w_asqrt46_24[1]),.dout(n11279),.clk(gclk));
	jnot g11042(.din(w_n10996_0[1]),.dout(n11280),.clk(gclk));
	jand g11043(.dina(n11280),.dinb(n11279),.dout(n11281),.clk(gclk));
	jor g11044(.dina(n11281),.dinb(n11170),.dout(n11282),.clk(gclk));
	jor g11045(.dina(n11282),.dinb(w_asqrt47_22[2]),.dout(n11283),.clk(gclk));
	jnot g11046(.din(w_n11003_0[1]),.dout(n11284),.clk(gclk));
	jand g11047(.dina(n11284),.dinb(n11283),.dout(n11285),.clk(gclk));
	jor g11048(.dina(n11285),.dinb(n11169),.dout(n11286),.clk(gclk));
	jor g11049(.dina(n11286),.dinb(w_asqrt48_24[2]),.dout(n11287),.clk(gclk));
	jand g11050(.dina(w_n11010_0[1]),.dinb(n11287),.dout(n11288),.clk(gclk));
	jor g11051(.dina(n11288),.dinb(n11168),.dout(n11289),.clk(gclk));
	jor g11052(.dina(n11289),.dinb(w_asqrt49_23[0]),.dout(n11290),.clk(gclk));
	jnot g11053(.din(w_n11018_0[1]),.dout(n11291),.clk(gclk));
	jand g11054(.dina(n11291),.dinb(n11290),.dout(n11292),.clk(gclk));
	jor g11055(.dina(n11292),.dinb(n11167),.dout(n11293),.clk(gclk));
	jor g11056(.dina(n11293),.dinb(w_asqrt50_25[0]),.dout(n11294),.clk(gclk));
	jand g11057(.dina(w_n11025_0[1]),.dinb(n11294),.dout(n11295),.clk(gclk));
	jor g11058(.dina(n11295),.dinb(n11166),.dout(n11296),.clk(gclk));
	jor g11059(.dina(n11296),.dinb(w_asqrt51_23[1]),.dout(n11297),.clk(gclk));
	jnot g11060(.din(w_n11033_0[1]),.dout(n11298),.clk(gclk));
	jand g11061(.dina(n11298),.dinb(n11297),.dout(n11299),.clk(gclk));
	jor g11062(.dina(n11299),.dinb(n11165),.dout(n11300),.clk(gclk));
	jor g11063(.dina(n11300),.dinb(w_asqrt52_25[0]),.dout(n11301),.clk(gclk));
	jand g11064(.dina(w_n11040_0[1]),.dinb(n11301),.dout(n11302),.clk(gclk));
	jor g11065(.dina(n11302),.dinb(n11164),.dout(n11303),.clk(gclk));
	jor g11066(.dina(n11303),.dinb(w_asqrt53_24[0]),.dout(n11304),.clk(gclk));
	jnot g11067(.din(w_n11048_0[1]),.dout(n11305),.clk(gclk));
	jand g11068(.dina(n11305),.dinb(n11304),.dout(n11306),.clk(gclk));
	jor g11069(.dina(n11306),.dinb(n11163),.dout(n11307),.clk(gclk));
	jor g11070(.dina(n11307),.dinb(w_asqrt54_25[0]),.dout(n11308),.clk(gclk));
	jand g11071(.dina(w_n11055_0[1]),.dinb(n11308),.dout(n11309),.clk(gclk));
	jor g11072(.dina(n11309),.dinb(n11162),.dout(n11310),.clk(gclk));
	jor g11073(.dina(n11310),.dinb(w_asqrt55_24[1]),.dout(n11311),.clk(gclk));
	jand g11074(.dina(w_n11063_0[1]),.dinb(n11311),.dout(n11312),.clk(gclk));
	jor g11075(.dina(n11312),.dinb(n11161),.dout(n11313),.clk(gclk));
	jor g11076(.dina(n11313),.dinb(w_asqrt56_25[1]),.dout(n11314),.clk(gclk));
	jand g11077(.dina(w_n11071_0[1]),.dinb(n11314),.dout(n11315),.clk(gclk));
	jor g11078(.dina(n11315),.dinb(n11160),.dout(n11316),.clk(gclk));
	jor g11079(.dina(n11316),.dinb(w_asqrt57_25[0]),.dout(n11317),.clk(gclk));
	jnot g11080(.din(w_n11079_0[1]),.dout(n11318),.clk(gclk));
	jand g11081(.dina(n11318),.dinb(n11317),.dout(n11319),.clk(gclk));
	jor g11082(.dina(n11319),.dinb(n11159),.dout(n11320),.clk(gclk));
	jor g11083(.dina(n11320),.dinb(w_asqrt58_25[2]),.dout(n11321),.clk(gclk));
	jnot g11084(.din(w_n11086_0[1]),.dout(n11322),.clk(gclk));
	jand g11085(.dina(n11322),.dinb(n11321),.dout(n11323),.clk(gclk));
	jor g11086(.dina(n11323),.dinb(n11158),.dout(n11324),.clk(gclk));
	jor g11087(.dina(n11324),.dinb(w_asqrt59_25[1]),.dout(n11325),.clk(gclk));
	jnot g11088(.din(w_n11093_0[1]),.dout(n11326),.clk(gclk));
	jand g11089(.dina(n11326),.dinb(n11325),.dout(n11327),.clk(gclk));
	jor g11090(.dina(n11327),.dinb(n11157),.dout(n11328),.clk(gclk));
	jor g11091(.dina(n11328),.dinb(w_asqrt60_25[2]),.dout(n11329),.clk(gclk));
	jand g11092(.dina(w_n11100_0[1]),.dinb(n11329),.dout(n11330),.clk(gclk));
	jor g11093(.dina(n11330),.dinb(n11156),.dout(n11331),.clk(gclk));
	jor g11094(.dina(n11331),.dinb(w_asqrt61_25[2]),.dout(n11332),.clk(gclk));
	jnot g11095(.din(w_n11108_0[1]),.dout(n11333),.clk(gclk));
	jand g11096(.dina(n11333),.dinb(n11332),.dout(n11334),.clk(gclk));
	jor g11097(.dina(n11334),.dinb(n11155),.dout(n11335),.clk(gclk));
	jor g11098(.dina(n11335),.dinb(w_asqrt62_25[2]),.dout(n11336),.clk(gclk));
	jand g11099(.dina(w_n11137_0[0]),.dinb(n11336),.dout(n11337),.clk(gclk));
	jor g11100(.dina(n11337),.dinb(n11154),.dout(n11338),.clk(gclk));
	jnot g11101(.din(w_n11120_0[2]),.dout(n11339),.clk(gclk));
	jand g11102(.dina(n11339),.dinb(n11338),.dout(n11340),.clk(gclk));
	jand g11103(.dina(n11340),.dinb(w_n10820_0[0]),.dout(n11341),.clk(gclk));
	jand g11104(.dina(n11341),.dinb(n11153),.dout(n11342),.clk(gclk));
	jor g11105(.dina(n11342),.dinb(w_asqrt63_32[1]),.dout(n11343),.clk(gclk));
	jnot g11106(.din(w_n11133_0[0]),.dout(n11344),.clk(gclk));
	jand g11107(.dina(n11344),.dinb(w_n11343_0[1]),.dout(n11345),.clk(gclk));
	jand g11108(.dina(n11345),.dinb(w_n11126_0[0]),.dout(n11346),.clk(gclk));
	jand g11109(.dina(w_n11346_0[1]),.dinb(w_n11152_0[1]),.dout(n11347),.clk(gclk));
	jor g11110(.dina(w_n11347_27[1]),.dinb(n11151),.dout(n11348),.clk(gclk));
	jand g11111(.dina(n11348),.dinb(n11150),.dout(n11349),.clk(gclk));
	jand g11112(.dina(n11349),.dinb(n11148),.dout(n11350),.clk(gclk));
	jor g11113(.dina(n11350),.dinb(w_n11147_0[1]),.dout(n11351),.clk(gclk));
	jand g11114(.dina(w_n11351_0[2]),.dinb(w_asqrt24_22[1]),.dout(n11352),.clk(gclk));
	jor g11115(.dina(w_n11351_0[1]),.dinb(w_asqrt24_22[0]),.dout(n11353),.clk(gclk));
	jand g11116(.dina(w_asqrt22_35[0]),.dinb(w_n10807_0[0]),.dout(n11354),.clk(gclk));
	jand g11117(.dina(w_n11152_0[0]),.dinb(w_asqrt23_16[0]),.dout(n11355),.clk(gclk));
	jand g11118(.dina(n11355),.dinb(w_n11125_0[0]),.dout(n11356),.clk(gclk));
	jand g11119(.dina(n11356),.dinb(w_n11343_0[0]),.dout(n11357),.clk(gclk));
	jor g11120(.dina(n11357),.dinb(w_n11354_0[1]),.dout(n11358),.clk(gclk));
	jxor g11121(.dina(n11358),.dinb(w_a46_0[1]),.dout(n11359),.clk(gclk));
	jnot g11122(.din(w_n11359_0[1]),.dout(n11360),.clk(gclk));
	jand g11123(.dina(w_n11360_0[1]),.dinb(n11353),.dout(n11361),.clk(gclk));
	jor g11124(.dina(n11361),.dinb(w_n11352_0[1]),.dout(n11362),.clk(gclk));
	jand g11125(.dina(w_n11362_0[2]),.dinb(w_asqrt25_16[1]),.dout(n11363),.clk(gclk));
	jor g11126(.dina(w_n11362_0[1]),.dinb(w_asqrt25_16[0]),.dout(n11364),.clk(gclk));
	jxor g11127(.dina(w_n10826_0[0]),.dinb(w_n10328_28[0]),.dout(n11365),.clk(gclk));
	jand g11128(.dina(n11365),.dinb(w_asqrt22_34[2]),.dout(n11366),.clk(gclk));
	jxor g11129(.dina(n11366),.dinb(w_n11198_0[0]),.dout(n11367),.clk(gclk));
	jand g11130(.dina(w_n11367_0[1]),.dinb(n11364),.dout(n11368),.clk(gclk));
	jor g11131(.dina(n11368),.dinb(w_n11363_0[1]),.dout(n11369),.clk(gclk));
	jand g11132(.dina(w_n11369_0[2]),.dinb(w_asqrt26_22[1]),.dout(n11370),.clk(gclk));
	jor g11133(.dina(w_n11369_0[1]),.dinb(w_asqrt26_22[0]),.dout(n11371),.clk(gclk));
	jxor g11134(.dina(w_n10834_0[0]),.dinb(w_n9832_34[1]),.dout(n11372),.clk(gclk));
	jand g11135(.dina(n11372),.dinb(w_asqrt22_34[1]),.dout(n11373),.clk(gclk));
	jxor g11136(.dina(n11373),.dinb(w_n10843_0[0]),.dout(n11374),.clk(gclk));
	jnot g11137(.din(w_n11374_0[1]),.dout(n11375),.clk(gclk));
	jand g11138(.dina(w_n11375_0[1]),.dinb(n11371),.dout(n11376),.clk(gclk));
	jor g11139(.dina(n11376),.dinb(w_n11370_0[1]),.dout(n11377),.clk(gclk));
	jand g11140(.dina(w_n11377_0[2]),.dinb(w_asqrt27_17[0]),.dout(n11378),.clk(gclk));
	jor g11141(.dina(w_n11377_0[1]),.dinb(w_asqrt27_16[2]),.dout(n11379),.clk(gclk));
	jxor g11142(.dina(w_n10845_0[0]),.dinb(w_n9369_29[0]),.dout(n11380),.clk(gclk));
	jand g11143(.dina(n11380),.dinb(w_asqrt22_34[0]),.dout(n11381),.clk(gclk));
	jxor g11144(.dina(n11381),.dinb(w_n10850_0[0]),.dout(n11382),.clk(gclk));
	jnot g11145(.din(w_n11382_0[1]),.dout(n11383),.clk(gclk));
	jand g11146(.dina(w_n11383_0[1]),.dinb(n11379),.dout(n11384),.clk(gclk));
	jor g11147(.dina(n11384),.dinb(w_n11378_0[1]),.dout(n11385),.clk(gclk));
	jand g11148(.dina(w_n11385_0[2]),.dinb(w_asqrt28_22[2]),.dout(n11386),.clk(gclk));
	jor g11149(.dina(w_n11385_0[1]),.dinb(w_asqrt28_22[1]),.dout(n11387),.clk(gclk));
	jxor g11150(.dina(w_n10852_0[0]),.dinb(w_n8890_34[2]),.dout(n11388),.clk(gclk));
	jand g11151(.dina(n11388),.dinb(w_asqrt22_33[2]),.dout(n11389),.clk(gclk));
	jxor g11152(.dina(n11389),.dinb(w_n10857_0[0]),.dout(n11390),.clk(gclk));
	jnot g11153(.din(w_n11390_0[1]),.dout(n11391),.clk(gclk));
	jand g11154(.dina(w_n11391_0[1]),.dinb(n11387),.dout(n11392),.clk(gclk));
	jor g11155(.dina(n11392),.dinb(w_n11386_0[1]),.dout(n11393),.clk(gclk));
	jand g11156(.dina(w_n11393_0[2]),.dinb(w_asqrt29_17[1]),.dout(n11394),.clk(gclk));
	jor g11157(.dina(w_n11393_0[1]),.dinb(w_asqrt29_17[0]),.dout(n11395),.clk(gclk));
	jxor g11158(.dina(w_n10859_0[0]),.dinb(w_n8449_29[2]),.dout(n11396),.clk(gclk));
	jand g11159(.dina(n11396),.dinb(w_asqrt22_33[1]),.dout(n11397),.clk(gclk));
	jxor g11160(.dina(n11397),.dinb(w_n10864_0[0]),.dout(n11398),.clk(gclk));
	jand g11161(.dina(w_n11398_0[1]),.dinb(n11395),.dout(n11399),.clk(gclk));
	jor g11162(.dina(n11399),.dinb(w_n11394_0[1]),.dout(n11400),.clk(gclk));
	jand g11163(.dina(w_n11400_0[2]),.dinb(w_asqrt30_23[0]),.dout(n11401),.clk(gclk));
	jor g11164(.dina(w_n11400_0[1]),.dinb(w_asqrt30_22[2]),.dout(n11402),.clk(gclk));
	jxor g11165(.dina(w_n10867_0[0]),.dinb(w_n8003_35[1]),.dout(n11403),.clk(gclk));
	jand g11166(.dina(n11403),.dinb(w_asqrt22_33[0]),.dout(n11404),.clk(gclk));
	jxor g11167(.dina(n11404),.dinb(w_n10872_0[0]),.dout(n11405),.clk(gclk));
	jnot g11168(.din(w_n11405_0[1]),.dout(n11406),.clk(gclk));
	jand g11169(.dina(w_n11406_0[1]),.dinb(n11402),.dout(n11407),.clk(gclk));
	jor g11170(.dina(n11407),.dinb(w_n11401_0[1]),.dout(n11408),.clk(gclk));
	jand g11171(.dina(w_n11408_0[2]),.dinb(w_asqrt31_18[0]),.dout(n11409),.clk(gclk));
	jor g11172(.dina(w_n11408_0[1]),.dinb(w_asqrt31_17[2]),.dout(n11410),.clk(gclk));
	jxor g11173(.dina(w_n10874_0[0]),.dinb(w_n7581_30[2]),.dout(n11411),.clk(gclk));
	jand g11174(.dina(n11411),.dinb(w_asqrt22_32[2]),.dout(n11412),.clk(gclk));
	jxor g11175(.dina(n11412),.dinb(w_n10879_0[0]),.dout(n11413),.clk(gclk));
	jand g11176(.dina(w_n11413_0[1]),.dinb(n11410),.dout(n11414),.clk(gclk));
	jor g11177(.dina(n11414),.dinb(w_n11409_0[1]),.dout(n11415),.clk(gclk));
	jand g11178(.dina(w_n11415_0[2]),.dinb(w_asqrt32_23[0]),.dout(n11416),.clk(gclk));
	jor g11179(.dina(w_n11415_0[1]),.dinb(w_asqrt32_22[2]),.dout(n11417),.clk(gclk));
	jxor g11180(.dina(w_n10882_0[0]),.dinb(w_n7154_35[2]),.dout(n11418),.clk(gclk));
	jand g11181(.dina(n11418),.dinb(w_asqrt22_32[1]),.dout(n11419),.clk(gclk));
	jxor g11182(.dina(n11419),.dinb(w_n10887_0[0]),.dout(n11420),.clk(gclk));
	jnot g11183(.din(w_n11420_0[1]),.dout(n11421),.clk(gclk));
	jand g11184(.dina(w_n11421_0[1]),.dinb(n11417),.dout(n11422),.clk(gclk));
	jor g11185(.dina(n11422),.dinb(w_n11416_0[1]),.dout(n11423),.clk(gclk));
	jand g11186(.dina(w_n11423_0[2]),.dinb(w_asqrt33_18[2]),.dout(n11424),.clk(gclk));
	jor g11187(.dina(w_n11423_0[1]),.dinb(w_asqrt33_18[1]),.dout(n11425),.clk(gclk));
	jxor g11188(.dina(w_n10889_0[0]),.dinb(w_n6758_31[1]),.dout(n11426),.clk(gclk));
	jand g11189(.dina(n11426),.dinb(w_asqrt22_32[0]),.dout(n11427),.clk(gclk));
	jxor g11190(.dina(n11427),.dinb(w_n10894_0[0]),.dout(n11428),.clk(gclk));
	jnot g11191(.din(w_n11428_0[1]),.dout(n11429),.clk(gclk));
	jand g11192(.dina(w_n11429_0[1]),.dinb(n11425),.dout(n11430),.clk(gclk));
	jor g11193(.dina(n11430),.dinb(w_n11424_0[1]),.dout(n11431),.clk(gclk));
	jand g11194(.dina(w_n11431_0[2]),.dinb(w_asqrt34_23[1]),.dout(n11432),.clk(gclk));
	jor g11195(.dina(w_n11431_0[1]),.dinb(w_asqrt34_23[0]),.dout(n11433),.clk(gclk));
	jxor g11196(.dina(w_n10896_0[0]),.dinb(w_n6357_36[0]),.dout(n11434),.clk(gclk));
	jand g11197(.dina(n11434),.dinb(w_asqrt22_31[2]),.dout(n11435),.clk(gclk));
	jxor g11198(.dina(n11435),.dinb(w_n10901_0[0]),.dout(n11436),.clk(gclk));
	jnot g11199(.din(w_n11436_0[1]),.dout(n11437),.clk(gclk));
	jand g11200(.dina(w_n11437_0[1]),.dinb(n11433),.dout(n11438),.clk(gclk));
	jor g11201(.dina(n11438),.dinb(w_n11432_0[1]),.dout(n11439),.clk(gclk));
	jand g11202(.dina(w_n11439_0[2]),.dinb(w_asqrt35_19[1]),.dout(n11440),.clk(gclk));
	jor g11203(.dina(w_n11439_0[1]),.dinb(w_asqrt35_19[0]),.dout(n11441),.clk(gclk));
	jxor g11204(.dina(w_n10903_0[0]),.dinb(w_n5989_32[0]),.dout(n11442),.clk(gclk));
	jand g11205(.dina(n11442),.dinb(w_asqrt22_31[1]),.dout(n11443),.clk(gclk));
	jxor g11206(.dina(n11443),.dinb(w_n10908_0[0]),.dout(n11444),.clk(gclk));
	jand g11207(.dina(w_n11444_0[1]),.dinb(n11441),.dout(n11445),.clk(gclk));
	jor g11208(.dina(n11445),.dinb(w_n11440_0[1]),.dout(n11446),.clk(gclk));
	jand g11209(.dina(w_n11446_0[2]),.dinb(w_asqrt36_23[1]),.dout(n11447),.clk(gclk));
	jor g11210(.dina(w_n11446_0[1]),.dinb(w_asqrt36_23[0]),.dout(n11448),.clk(gclk));
	jxor g11211(.dina(w_n10911_0[0]),.dinb(w_n5606_36[1]),.dout(n11449),.clk(gclk));
	jand g11212(.dina(n11449),.dinb(w_asqrt22_31[0]),.dout(n11450),.clk(gclk));
	jxor g11213(.dina(n11450),.dinb(w_n10916_0[0]),.dout(n11451),.clk(gclk));
	jnot g11214(.din(w_n11451_0[1]),.dout(n11452),.clk(gclk));
	jand g11215(.dina(w_n11452_0[1]),.dinb(n11448),.dout(n11453),.clk(gclk));
	jor g11216(.dina(n11453),.dinb(w_n11447_0[1]),.dout(n11454),.clk(gclk));
	jand g11217(.dina(w_n11454_0[2]),.dinb(w_asqrt37_19[2]),.dout(n11455),.clk(gclk));
	jor g11218(.dina(w_n11454_0[1]),.dinb(w_asqrt37_19[1]),.dout(n11456),.clk(gclk));
	jxor g11219(.dina(w_n10918_0[0]),.dinb(w_n5259_33[0]),.dout(n11457),.clk(gclk));
	jand g11220(.dina(n11457),.dinb(w_asqrt22_30[2]),.dout(n11458),.clk(gclk));
	jxor g11221(.dina(n11458),.dinb(w_n10923_0[0]),.dout(n11459),.clk(gclk));
	jnot g11222(.din(w_n11459_0[1]),.dout(n11460),.clk(gclk));
	jand g11223(.dina(w_n11460_0[1]),.dinb(n11456),.dout(n11461),.clk(gclk));
	jor g11224(.dina(n11461),.dinb(w_n11455_0[1]),.dout(n11462),.clk(gclk));
	jand g11225(.dina(w_n11462_0[2]),.dinb(w_asqrt38_23[2]),.dout(n11463),.clk(gclk));
	jor g11226(.dina(w_n11462_0[1]),.dinb(w_asqrt38_23[1]),.dout(n11464),.clk(gclk));
	jxor g11227(.dina(w_n10925_0[0]),.dinb(w_n4902_37[0]),.dout(n11465),.clk(gclk));
	jand g11228(.dina(n11465),.dinb(w_asqrt22_30[1]),.dout(n11466),.clk(gclk));
	jxor g11229(.dina(n11466),.dinb(w_n10930_0[0]),.dout(n11467),.clk(gclk));
	jnot g11230(.din(w_n11467_0[1]),.dout(n11468),.clk(gclk));
	jand g11231(.dina(w_n11468_0[1]),.dinb(n11464),.dout(n11469),.clk(gclk));
	jor g11232(.dina(n11469),.dinb(w_n11463_0[1]),.dout(n11470),.clk(gclk));
	jand g11233(.dina(w_n11470_0[2]),.dinb(w_asqrt39_20[1]),.dout(n11471),.clk(gclk));
	jor g11234(.dina(w_n11470_0[1]),.dinb(w_asqrt39_20[0]),.dout(n11472),.clk(gclk));
	jxor g11235(.dina(w_n10932_0[0]),.dinb(w_n4582_34[0]),.dout(n11473),.clk(gclk));
	jand g11236(.dina(n11473),.dinb(w_asqrt22_30[0]),.dout(n11474),.clk(gclk));
	jxor g11237(.dina(n11474),.dinb(w_n10937_0[0]),.dout(n11475),.clk(gclk));
	jnot g11238(.din(w_n11475_0[1]),.dout(n11476),.clk(gclk));
	jand g11239(.dina(w_n11476_0[1]),.dinb(n11472),.dout(n11477),.clk(gclk));
	jor g11240(.dina(n11477),.dinb(w_n11471_0[1]),.dout(n11478),.clk(gclk));
	jand g11241(.dina(w_n11478_0[2]),.dinb(w_asqrt40_23[2]),.dout(n11479),.clk(gclk));
	jor g11242(.dina(w_n11478_0[1]),.dinb(w_asqrt40_23[1]),.dout(n11480),.clk(gclk));
	jxor g11243(.dina(w_n10939_0[0]),.dinb(w_n4249_37[2]),.dout(n11481),.clk(gclk));
	jand g11244(.dina(n11481),.dinb(w_asqrt22_29[2]),.dout(n11482),.clk(gclk));
	jxor g11245(.dina(n11482),.dinb(w_n10944_0[0]),.dout(n11483),.clk(gclk));
	jnot g11246(.din(w_n11483_0[1]),.dout(n11484),.clk(gclk));
	jand g11247(.dina(w_n11484_0[1]),.dinb(n11480),.dout(n11485),.clk(gclk));
	jor g11248(.dina(n11485),.dinb(w_n11479_0[1]),.dout(n11486),.clk(gclk));
	jand g11249(.dina(w_n11486_0[2]),.dinb(w_asqrt41_20[2]),.dout(n11487),.clk(gclk));
	jxor g11250(.dina(w_n10946_0[0]),.dinb(w_n3955_34[2]),.dout(n11488),.clk(gclk));
	jand g11251(.dina(n11488),.dinb(w_asqrt22_29[1]),.dout(n11489),.clk(gclk));
	jxor g11252(.dina(n11489),.dinb(w_n10950_0[0]),.dout(n11490),.clk(gclk));
	jor g11253(.dina(w_n11486_0[1]),.dinb(w_asqrt41_20[1]),.dout(n11491),.clk(gclk));
	jand g11254(.dina(n11491),.dinb(w_n11490_0[1]),.dout(n11492),.clk(gclk));
	jor g11255(.dina(n11492),.dinb(w_n11487_0[1]),.dout(n11493),.clk(gclk));
	jand g11256(.dina(w_n11493_0[2]),.dinb(w_asqrt42_24[0]),.dout(n11494),.clk(gclk));
	jor g11257(.dina(w_n11493_0[1]),.dinb(w_asqrt42_23[2]),.dout(n11495),.clk(gclk));
	jxor g11258(.dina(w_n10954_0[0]),.dinb(w_n3642_38[0]),.dout(n11496),.clk(gclk));
	jand g11259(.dina(n11496),.dinb(w_asqrt22_29[0]),.dout(n11497),.clk(gclk));
	jxor g11260(.dina(n11497),.dinb(w_n10959_0[0]),.dout(n11498),.clk(gclk));
	jnot g11261(.din(w_n11498_0[1]),.dout(n11499),.clk(gclk));
	jand g11262(.dina(w_n11499_0[1]),.dinb(n11495),.dout(n11500),.clk(gclk));
	jor g11263(.dina(n11500),.dinb(w_n11494_0[1]),.dout(n11501),.clk(gclk));
	jand g11264(.dina(w_n11501_0[2]),.dinb(w_asqrt43_21[0]),.dout(n11502),.clk(gclk));
	jor g11265(.dina(w_n11501_0[1]),.dinb(w_asqrt43_20[2]),.dout(n11503),.clk(gclk));
	jxor g11266(.dina(w_n10961_0[0]),.dinb(w_n3368_35[1]),.dout(n11504),.clk(gclk));
	jand g11267(.dina(n11504),.dinb(w_asqrt22_28[2]),.dout(n11505),.clk(gclk));
	jxor g11268(.dina(n11505),.dinb(w_n10966_0[0]),.dout(n11506),.clk(gclk));
	jand g11269(.dina(w_n11506_0[1]),.dinb(n11503),.dout(n11507),.clk(gclk));
	jor g11270(.dina(n11507),.dinb(w_n11502_0[1]),.dout(n11508),.clk(gclk));
	jand g11271(.dina(w_n11508_0[2]),.dinb(w_asqrt44_24[0]),.dout(n11509),.clk(gclk));
	jor g11272(.dina(w_n11508_0[1]),.dinb(w_asqrt44_23[2]),.dout(n11510),.clk(gclk));
	jxor g11273(.dina(w_n10969_0[0]),.dinb(w_n3089_38[2]),.dout(n11511),.clk(gclk));
	jand g11274(.dina(n11511),.dinb(w_asqrt22_28[1]),.dout(n11512),.clk(gclk));
	jxor g11275(.dina(n11512),.dinb(w_n10974_0[0]),.dout(n11513),.clk(gclk));
	jnot g11276(.din(w_n11513_0[1]),.dout(n11514),.clk(gclk));
	jand g11277(.dina(w_n11514_0[1]),.dinb(n11510),.dout(n11515),.clk(gclk));
	jor g11278(.dina(n11515),.dinb(w_n11509_0[1]),.dout(n11516),.clk(gclk));
	jand g11279(.dina(w_n11516_0[2]),.dinb(w_asqrt45_21[2]),.dout(n11517),.clk(gclk));
	jor g11280(.dina(w_n11516_0[1]),.dinb(w_asqrt45_21[1]),.dout(n11518),.clk(gclk));
	jxor g11281(.dina(w_n10976_0[0]),.dinb(w_n2833_36[1]),.dout(n11519),.clk(gclk));
	jand g11282(.dina(n11519),.dinb(w_asqrt22_28[0]),.dout(n11520),.clk(gclk));
	jxor g11283(.dina(n11520),.dinb(w_n10981_0[0]),.dout(n11521),.clk(gclk));
	jand g11284(.dina(w_n11521_0[1]),.dinb(n11518),.dout(n11522),.clk(gclk));
	jor g11285(.dina(n11522),.dinb(w_n11517_0[1]),.dout(n11523),.clk(gclk));
	jand g11286(.dina(w_n11523_0[2]),.dinb(w_asqrt46_24[0]),.dout(n11524),.clk(gclk));
	jor g11287(.dina(w_n11523_0[1]),.dinb(w_asqrt46_23[2]),.dout(n11525),.clk(gclk));
	jxor g11288(.dina(w_n10984_0[0]),.dinb(w_n2572_39[0]),.dout(n11526),.clk(gclk));
	jand g11289(.dina(n11526),.dinb(w_asqrt22_27[2]),.dout(n11527),.clk(gclk));
	jxor g11290(.dina(n11527),.dinb(w_n10989_0[0]),.dout(n11528),.clk(gclk));
	jnot g11291(.din(w_n11528_0[1]),.dout(n11529),.clk(gclk));
	jand g11292(.dina(w_n11529_0[1]),.dinb(n11525),.dout(n11530),.clk(gclk));
	jor g11293(.dina(n11530),.dinb(w_n11524_0[1]),.dout(n11531),.clk(gclk));
	jand g11294(.dina(w_n11531_0[2]),.dinb(w_asqrt47_22[1]),.dout(n11532),.clk(gclk));
	jor g11295(.dina(w_n11531_0[1]),.dinb(w_asqrt47_22[0]),.dout(n11533),.clk(gclk));
	jxor g11296(.dina(w_n10991_0[0]),.dinb(w_n2345_37[0]),.dout(n11534),.clk(gclk));
	jand g11297(.dina(n11534),.dinb(w_asqrt22_27[1]),.dout(n11535),.clk(gclk));
	jxor g11298(.dina(n11535),.dinb(w_n10996_0[0]),.dout(n11536),.clk(gclk));
	jnot g11299(.din(w_n11536_0[1]),.dout(n11537),.clk(gclk));
	jand g11300(.dina(w_n11537_0[1]),.dinb(n11533),.dout(n11538),.clk(gclk));
	jor g11301(.dina(n11538),.dinb(w_n11532_0[1]),.dout(n11539),.clk(gclk));
	jand g11302(.dina(w_n11539_0[2]),.dinb(w_asqrt48_24[1]),.dout(n11540),.clk(gclk));
	jor g11303(.dina(w_n11539_0[1]),.dinb(w_asqrt48_24[0]),.dout(n11541),.clk(gclk));
	jxor g11304(.dina(w_n10998_0[0]),.dinb(w_n2108_39[2]),.dout(n11542),.clk(gclk));
	jand g11305(.dina(n11542),.dinb(w_asqrt22_27[0]),.dout(n11543),.clk(gclk));
	jxor g11306(.dina(n11543),.dinb(w_n11003_0[0]),.dout(n11544),.clk(gclk));
	jnot g11307(.din(w_n11544_0[1]),.dout(n11545),.clk(gclk));
	jand g11308(.dina(w_n11545_0[1]),.dinb(n11541),.dout(n11546),.clk(gclk));
	jor g11309(.dina(n11546),.dinb(w_n11540_0[1]),.dout(n11547),.clk(gclk));
	jand g11310(.dina(w_n11547_0[2]),.dinb(w_asqrt49_22[2]),.dout(n11548),.clk(gclk));
	jor g11311(.dina(w_n11547_0[1]),.dinb(w_asqrt49_22[1]),.dout(n11549),.clk(gclk));
	jxor g11312(.dina(w_n11005_0[0]),.dinb(w_n1912_38[0]),.dout(n11550),.clk(gclk));
	jand g11313(.dina(n11550),.dinb(w_asqrt22_26[2]),.dout(n11551),.clk(gclk));
	jxor g11314(.dina(n11551),.dinb(w_n11010_0[0]),.dout(n11552),.clk(gclk));
	jand g11315(.dina(w_n11552_0[1]),.dinb(n11549),.dout(n11553),.clk(gclk));
	jor g11316(.dina(n11553),.dinb(w_n11548_0[1]),.dout(n11554),.clk(gclk));
	jand g11317(.dina(w_n11554_0[2]),.dinb(w_asqrt50_24[2]),.dout(n11555),.clk(gclk));
	jor g11318(.dina(w_n11554_0[1]),.dinb(w_asqrt50_24[1]),.dout(n11556),.clk(gclk));
	jxor g11319(.dina(w_n11013_0[0]),.dinb(w_n1699_40[1]),.dout(n11557),.clk(gclk));
	jand g11320(.dina(n11557),.dinb(w_asqrt22_26[1]),.dout(n11558),.clk(gclk));
	jxor g11321(.dina(n11558),.dinb(w_n11018_0[0]),.dout(n11559),.clk(gclk));
	jnot g11322(.din(w_n11559_0[1]),.dout(n11560),.clk(gclk));
	jand g11323(.dina(w_n11560_0[1]),.dinb(n11556),.dout(n11561),.clk(gclk));
	jor g11324(.dina(n11561),.dinb(w_n11555_0[1]),.dout(n11562),.clk(gclk));
	jand g11325(.dina(w_n11562_0[2]),.dinb(w_asqrt51_23[0]),.dout(n11563),.clk(gclk));
	jor g11326(.dina(w_n11562_0[1]),.dinb(w_asqrt51_22[2]),.dout(n11564),.clk(gclk));
	jxor g11327(.dina(w_n11020_0[0]),.dinb(w_n1516_38[2]),.dout(n11565),.clk(gclk));
	jand g11328(.dina(n11565),.dinb(w_asqrt22_26[0]),.dout(n11566),.clk(gclk));
	jxor g11329(.dina(n11566),.dinb(w_n11025_0[0]),.dout(n11567),.clk(gclk));
	jand g11330(.dina(w_n11567_0[1]),.dinb(n11564),.dout(n11568),.clk(gclk));
	jor g11331(.dina(n11568),.dinb(w_n11563_0[1]),.dout(n11569),.clk(gclk));
	jand g11332(.dina(w_n11569_0[2]),.dinb(w_asqrt52_24[2]),.dout(n11570),.clk(gclk));
	jor g11333(.dina(w_n11569_0[1]),.dinb(w_asqrt52_24[1]),.dout(n11571),.clk(gclk));
	jxor g11334(.dina(w_n11028_0[0]),.dinb(w_n1332_40[1]),.dout(n11572),.clk(gclk));
	jand g11335(.dina(n11572),.dinb(w_asqrt22_25[2]),.dout(n11573),.clk(gclk));
	jxor g11336(.dina(n11573),.dinb(w_n11033_0[0]),.dout(n11574),.clk(gclk));
	jnot g11337(.din(w_n11574_0[1]),.dout(n11575),.clk(gclk));
	jand g11338(.dina(w_n11575_0[1]),.dinb(n11571),.dout(n11576),.clk(gclk));
	jor g11339(.dina(n11576),.dinb(w_n11570_0[1]),.dout(n11577),.clk(gclk));
	jand g11340(.dina(w_n11577_0[2]),.dinb(w_asqrt53_23[2]),.dout(n11578),.clk(gclk));
	jor g11341(.dina(w_n11577_0[1]),.dinb(w_asqrt53_23[1]),.dout(n11579),.clk(gclk));
	jxor g11342(.dina(w_n11035_0[0]),.dinb(w_n1173_39[1]),.dout(n11580),.clk(gclk));
	jand g11343(.dina(n11580),.dinb(w_asqrt22_25[1]),.dout(n11581),.clk(gclk));
	jxor g11344(.dina(n11581),.dinb(w_n11040_0[0]),.dout(n11582),.clk(gclk));
	jand g11345(.dina(w_n11582_0[1]),.dinb(n11579),.dout(n11583),.clk(gclk));
	jor g11346(.dina(n11583),.dinb(w_n11578_0[1]),.dout(n11584),.clk(gclk));
	jand g11347(.dina(w_n11584_0[2]),.dinb(w_asqrt54_24[2]),.dout(n11585),.clk(gclk));
	jor g11348(.dina(w_n11584_0[1]),.dinb(w_asqrt54_24[1]),.dout(n11586),.clk(gclk));
	jxor g11349(.dina(w_n11043_0[0]),.dinb(w_n1008_41[1]),.dout(n11587),.clk(gclk));
	jand g11350(.dina(n11587),.dinb(w_asqrt22_25[0]),.dout(n11588),.clk(gclk));
	jxor g11351(.dina(n11588),.dinb(w_n11048_0[0]),.dout(n11589),.clk(gclk));
	jnot g11352(.din(w_n11589_0[1]),.dout(n11590),.clk(gclk));
	jand g11353(.dina(w_n11590_0[1]),.dinb(n11586),.dout(n11591),.clk(gclk));
	jor g11354(.dina(n11591),.dinb(w_n11585_0[1]),.dout(n11592),.clk(gclk));
	jand g11355(.dina(w_n11592_0[2]),.dinb(w_asqrt55_24[0]),.dout(n11593),.clk(gclk));
	jor g11356(.dina(w_n11592_0[1]),.dinb(w_asqrt55_23[2]),.dout(n11594),.clk(gclk));
	jxor g11357(.dina(w_n11050_0[0]),.dinb(w_n884_40[1]),.dout(n11595),.clk(gclk));
	jand g11358(.dina(n11595),.dinb(w_asqrt22_24[2]),.dout(n11596),.clk(gclk));
	jxor g11359(.dina(n11596),.dinb(w_n11055_0[0]),.dout(n11597),.clk(gclk));
	jand g11360(.dina(w_n11597_0[1]),.dinb(n11594),.dout(n11598),.clk(gclk));
	jor g11361(.dina(n11598),.dinb(w_n11593_0[1]),.dout(n11599),.clk(gclk));
	jand g11362(.dina(w_n11599_0[2]),.dinb(w_asqrt56_25[0]),.dout(n11600),.clk(gclk));
	jor g11363(.dina(w_n11599_0[1]),.dinb(w_asqrt56_24[2]),.dout(n11601),.clk(gclk));
	jxor g11364(.dina(w_n11058_0[0]),.dinb(w_n743_41[1]),.dout(n11602),.clk(gclk));
	jand g11365(.dina(n11602),.dinb(w_asqrt22_24[1]),.dout(n11603),.clk(gclk));
	jxor g11366(.dina(n11603),.dinb(w_n11063_0[0]),.dout(n11604),.clk(gclk));
	jand g11367(.dina(w_n11604_0[1]),.dinb(n11601),.dout(n11605),.clk(gclk));
	jor g11368(.dina(n11605),.dinb(w_n11600_0[1]),.dout(n11606),.clk(gclk));
	jand g11369(.dina(w_n11606_0[2]),.dinb(w_asqrt57_24[2]),.dout(n11607),.clk(gclk));
	jor g11370(.dina(w_n11606_0[1]),.dinb(w_asqrt57_24[1]),.dout(n11608),.clk(gclk));
	jxor g11371(.dina(w_n11066_0[0]),.dinb(w_n635_41[1]),.dout(n11609),.clk(gclk));
	jand g11372(.dina(n11609),.dinb(w_asqrt22_24[0]),.dout(n11610),.clk(gclk));
	jxor g11373(.dina(n11610),.dinb(w_n11071_0[0]),.dout(n11611),.clk(gclk));
	jand g11374(.dina(w_n11611_0[1]),.dinb(n11608),.dout(n11612),.clk(gclk));
	jor g11375(.dina(n11612),.dinb(w_n11607_0[1]),.dout(n11613),.clk(gclk));
	jand g11376(.dina(w_n11613_0[2]),.dinb(w_asqrt58_25[1]),.dout(n11614),.clk(gclk));
	jor g11377(.dina(w_n11613_0[1]),.dinb(w_asqrt58_25[0]),.dout(n11615),.clk(gclk));
	jxor g11378(.dina(w_n11074_0[0]),.dinb(w_n515_42[1]),.dout(n11616),.clk(gclk));
	jand g11379(.dina(n11616),.dinb(w_asqrt22_23[2]),.dout(n11617),.clk(gclk));
	jxor g11380(.dina(n11617),.dinb(w_n11079_0[0]),.dout(n11618),.clk(gclk));
	jnot g11381(.din(w_n11618_0[1]),.dout(n11619),.clk(gclk));
	jand g11382(.dina(w_n11619_0[1]),.dinb(n11615),.dout(n11620),.clk(gclk));
	jor g11383(.dina(n11620),.dinb(w_n11614_0[1]),.dout(n11621),.clk(gclk));
	jand g11384(.dina(w_n11621_0[2]),.dinb(w_asqrt59_25[0]),.dout(n11622),.clk(gclk));
	jor g11385(.dina(w_n11621_0[1]),.dinb(w_asqrt59_24[2]),.dout(n11623),.clk(gclk));
	jxor g11386(.dina(w_n11081_0[0]),.dinb(w_n443_42[1]),.dout(n11624),.clk(gclk));
	jand g11387(.dina(n11624),.dinb(w_asqrt22_23[1]),.dout(n11625),.clk(gclk));
	jxor g11388(.dina(n11625),.dinb(w_n11086_0[0]),.dout(n11626),.clk(gclk));
	jnot g11389(.din(w_n11626_0[1]),.dout(n11627),.clk(gclk));
	jand g11390(.dina(w_n11627_0[1]),.dinb(n11623),.dout(n11628),.clk(gclk));
	jor g11391(.dina(n11628),.dinb(w_n11622_0[1]),.dout(n11629),.clk(gclk));
	jand g11392(.dina(w_n11629_0[2]),.dinb(w_asqrt60_25[1]),.dout(n11630),.clk(gclk));
	jor g11393(.dina(w_n11629_0[1]),.dinb(w_asqrt60_25[0]),.dout(n11631),.clk(gclk));
	jxor g11394(.dina(w_n11088_0[0]),.dinb(w_n352_42[2]),.dout(n11632),.clk(gclk));
	jand g11395(.dina(n11632),.dinb(w_asqrt22_23[0]),.dout(n11633),.clk(gclk));
	jxor g11396(.dina(n11633),.dinb(w_n11093_0[0]),.dout(n11634),.clk(gclk));
	jnot g11397(.din(w_n11634_0[1]),.dout(n11635),.clk(gclk));
	jand g11398(.dina(w_n11635_0[1]),.dinb(n11631),.dout(n11636),.clk(gclk));
	jor g11399(.dina(n11636),.dinb(w_n11630_0[1]),.dout(n11637),.clk(gclk));
	jand g11400(.dina(w_n11637_0[2]),.dinb(w_asqrt61_25[1]),.dout(n11638),.clk(gclk));
	jor g11401(.dina(w_n11637_0[1]),.dinb(w_asqrt61_25[0]),.dout(n11639),.clk(gclk));
	jxor g11402(.dina(w_n11095_0[0]),.dinb(w_n294_43[0]),.dout(n11640),.clk(gclk));
	jand g11403(.dina(n11640),.dinb(w_asqrt22_22[2]),.dout(n11641),.clk(gclk));
	jxor g11404(.dina(n11641),.dinb(w_n11100_0[0]),.dout(n11642),.clk(gclk));
	jand g11405(.dina(w_n11642_0[1]),.dinb(n11639),.dout(n11643),.clk(gclk));
	jor g11406(.dina(n11643),.dinb(w_n11638_0[1]),.dout(n11644),.clk(gclk));
	jand g11407(.dina(w_n11644_0[2]),.dinb(w_asqrt62_25[1]),.dout(n11645),.clk(gclk));
	jor g11408(.dina(w_n11644_0[1]),.dinb(w_asqrt62_25[0]),.dout(n11646),.clk(gclk));
	jxor g11409(.dina(w_n11103_0[0]),.dinb(w_n239_43[0]),.dout(n11647),.clk(gclk));
	jand g11410(.dina(n11647),.dinb(w_asqrt22_22[1]),.dout(n11648),.clk(gclk));
	jxor g11411(.dina(n11648),.dinb(w_n11108_0[0]),.dout(n11649),.clk(gclk));
	jnot g11412(.din(w_n11649_0[2]),.dout(n11650),.clk(gclk));
	jand g11413(.dina(n11650),.dinb(n11646),.dout(n11651),.clk(gclk));
	jor g11414(.dina(n11651),.dinb(w_n11645_0[1]),.dout(n11652),.clk(gclk));
	jor g11415(.dina(w_n11652_0[1]),.dinb(w_n11140_0[2]),.dout(n11653),.clk(gclk));
	jnot g11416(.din(w_n11653_1[1]),.dout(n11654),.clk(gclk));
	jnot g11417(.din(w_n11140_0[1]),.dout(n11656),.clk(gclk));
	jnot g11418(.din(w_n11645_0[0]),.dout(n11657),.clk(gclk));
	jnot g11419(.din(w_n11638_0[0]),.dout(n11658),.clk(gclk));
	jnot g11420(.din(w_n11630_0[0]),.dout(n11659),.clk(gclk));
	jnot g11421(.din(w_n11622_0[0]),.dout(n11660),.clk(gclk));
	jnot g11422(.din(w_n11614_0[0]),.dout(n11661),.clk(gclk));
	jnot g11423(.din(w_n11607_0[0]),.dout(n11662),.clk(gclk));
	jnot g11424(.din(w_n11600_0[0]),.dout(n11663),.clk(gclk));
	jnot g11425(.din(w_n11593_0[0]),.dout(n11664),.clk(gclk));
	jnot g11426(.din(w_n11585_0[0]),.dout(n11665),.clk(gclk));
	jnot g11427(.din(w_n11578_0[0]),.dout(n11666),.clk(gclk));
	jnot g11428(.din(w_n11570_0[0]),.dout(n11667),.clk(gclk));
	jnot g11429(.din(w_n11563_0[0]),.dout(n11668),.clk(gclk));
	jnot g11430(.din(w_n11555_0[0]),.dout(n11669),.clk(gclk));
	jnot g11431(.din(w_n11548_0[0]),.dout(n11670),.clk(gclk));
	jnot g11432(.din(w_n11540_0[0]),.dout(n11671),.clk(gclk));
	jnot g11433(.din(w_n11532_0[0]),.dout(n11672),.clk(gclk));
	jnot g11434(.din(w_n11524_0[0]),.dout(n11673),.clk(gclk));
	jnot g11435(.din(w_n11517_0[0]),.dout(n11674),.clk(gclk));
	jnot g11436(.din(w_n11509_0[0]),.dout(n11675),.clk(gclk));
	jnot g11437(.din(w_n11502_0[0]),.dout(n11676),.clk(gclk));
	jnot g11438(.din(w_n11494_0[0]),.dout(n11677),.clk(gclk));
	jnot g11439(.din(w_n11487_0[0]),.dout(n11678),.clk(gclk));
	jnot g11440(.din(w_n11490_0[0]),.dout(n11679),.clk(gclk));
	jnot g11441(.din(w_n11479_0[0]),.dout(n11680),.clk(gclk));
	jnot g11442(.din(w_n11471_0[0]),.dout(n11681),.clk(gclk));
	jnot g11443(.din(w_n11463_0[0]),.dout(n11682),.clk(gclk));
	jnot g11444(.din(w_n11455_0[0]),.dout(n11683),.clk(gclk));
	jnot g11445(.din(w_n11447_0[0]),.dout(n11684),.clk(gclk));
	jnot g11446(.din(w_n11440_0[0]),.dout(n11685),.clk(gclk));
	jnot g11447(.din(w_n11432_0[0]),.dout(n11686),.clk(gclk));
	jnot g11448(.din(w_n11424_0[0]),.dout(n11687),.clk(gclk));
	jnot g11449(.din(w_n11416_0[0]),.dout(n11688),.clk(gclk));
	jnot g11450(.din(w_n11409_0[0]),.dout(n11689),.clk(gclk));
	jnot g11451(.din(w_n11401_0[0]),.dout(n11690),.clk(gclk));
	jnot g11452(.din(w_n11394_0[0]),.dout(n11691),.clk(gclk));
	jnot g11453(.din(w_n11386_0[0]),.dout(n11692),.clk(gclk));
	jnot g11454(.din(w_n11378_0[0]),.dout(n11693),.clk(gclk));
	jnot g11455(.din(w_n11370_0[0]),.dout(n11694),.clk(gclk));
	jnot g11456(.din(w_n11363_0[0]),.dout(n11695),.clk(gclk));
	jnot g11457(.din(w_n11352_0[0]),.dout(n11696),.clk(gclk));
	jnot g11458(.din(w_n11147_0[0]),.dout(n11697),.clk(gclk));
	jor g11459(.dina(w_n11347_27[0]),.dinb(w_n10805_0[2]),.dout(n11698),.clk(gclk));
	jnot g11460(.din(w_n11145_0[0]),.dout(n11699),.clk(gclk));
	jand g11461(.dina(n11699),.dinb(n11698),.dout(n11700),.clk(gclk));
	jand g11462(.dina(n11700),.dinb(w_n10824_33[1]),.dout(n11701),.clk(gclk));
	jor g11463(.dina(w_n11347_26[2]),.dinb(w_a44_0[0]),.dout(n11702),.clk(gclk));
	jand g11464(.dina(n11702),.dinb(w_a45_0[0]),.dout(n11703),.clk(gclk));
	jor g11465(.dina(w_n11354_0[0]),.dinb(n11703),.dout(n11704),.clk(gclk));
	jor g11466(.dina(w_n11704_0[1]),.dinb(n11701),.dout(n11705),.clk(gclk));
	jand g11467(.dina(n11705),.dinb(n11697),.dout(n11706),.clk(gclk));
	jand g11468(.dina(n11706),.dinb(w_n10328_27[2]),.dout(n11707),.clk(gclk));
	jor g11469(.dina(w_n11359_0[0]),.dinb(n11707),.dout(n11708),.clk(gclk));
	jand g11470(.dina(n11708),.dinb(n11696),.dout(n11709),.clk(gclk));
	jand g11471(.dina(n11709),.dinb(w_n9832_34[0]),.dout(n11710),.clk(gclk));
	jnot g11472(.din(w_n11367_0[0]),.dout(n11711),.clk(gclk));
	jor g11473(.dina(w_n11711_0[1]),.dinb(n11710),.dout(n11712),.clk(gclk));
	jand g11474(.dina(n11712),.dinb(n11695),.dout(n11713),.clk(gclk));
	jand g11475(.dina(n11713),.dinb(w_n9369_28[2]),.dout(n11714),.clk(gclk));
	jor g11476(.dina(w_n11374_0[0]),.dinb(n11714),.dout(n11715),.clk(gclk));
	jand g11477(.dina(n11715),.dinb(n11694),.dout(n11716),.clk(gclk));
	jand g11478(.dina(n11716),.dinb(w_n8890_34[1]),.dout(n11717),.clk(gclk));
	jor g11479(.dina(w_n11382_0[0]),.dinb(n11717),.dout(n11718),.clk(gclk));
	jand g11480(.dina(n11718),.dinb(n11693),.dout(n11719),.clk(gclk));
	jand g11481(.dina(n11719),.dinb(w_n8449_29[1]),.dout(n11720),.clk(gclk));
	jor g11482(.dina(w_n11390_0[0]),.dinb(n11720),.dout(n11721),.clk(gclk));
	jand g11483(.dina(n11721),.dinb(n11692),.dout(n11722),.clk(gclk));
	jand g11484(.dina(n11722),.dinb(w_n8003_35[0]),.dout(n11723),.clk(gclk));
	jnot g11485(.din(w_n11398_0[0]),.dout(n11724),.clk(gclk));
	jor g11486(.dina(w_n11724_0[1]),.dinb(n11723),.dout(n11725),.clk(gclk));
	jand g11487(.dina(n11725),.dinb(n11691),.dout(n11726),.clk(gclk));
	jand g11488(.dina(n11726),.dinb(w_n7581_30[1]),.dout(n11727),.clk(gclk));
	jor g11489(.dina(w_n11405_0[0]),.dinb(n11727),.dout(n11728),.clk(gclk));
	jand g11490(.dina(n11728),.dinb(n11690),.dout(n11729),.clk(gclk));
	jand g11491(.dina(n11729),.dinb(w_n7154_35[1]),.dout(n11730),.clk(gclk));
	jnot g11492(.din(w_n11413_0[0]),.dout(n11731),.clk(gclk));
	jor g11493(.dina(w_n11731_0[1]),.dinb(n11730),.dout(n11732),.clk(gclk));
	jand g11494(.dina(n11732),.dinb(n11689),.dout(n11733),.clk(gclk));
	jand g11495(.dina(n11733),.dinb(w_n6758_31[0]),.dout(n11734),.clk(gclk));
	jor g11496(.dina(w_n11420_0[0]),.dinb(n11734),.dout(n11735),.clk(gclk));
	jand g11497(.dina(n11735),.dinb(n11688),.dout(n11736),.clk(gclk));
	jand g11498(.dina(n11736),.dinb(w_n6357_35[2]),.dout(n11737),.clk(gclk));
	jor g11499(.dina(w_n11428_0[0]),.dinb(n11737),.dout(n11738),.clk(gclk));
	jand g11500(.dina(n11738),.dinb(n11687),.dout(n11739),.clk(gclk));
	jand g11501(.dina(n11739),.dinb(w_n5989_31[2]),.dout(n11740),.clk(gclk));
	jor g11502(.dina(w_n11436_0[0]),.dinb(n11740),.dout(n11741),.clk(gclk));
	jand g11503(.dina(n11741),.dinb(n11686),.dout(n11742),.clk(gclk));
	jand g11504(.dina(n11742),.dinb(w_n5606_36[0]),.dout(n11743),.clk(gclk));
	jnot g11505(.din(w_n11444_0[0]),.dout(n11744),.clk(gclk));
	jor g11506(.dina(w_n11744_0[1]),.dinb(n11743),.dout(n11745),.clk(gclk));
	jand g11507(.dina(n11745),.dinb(n11685),.dout(n11746),.clk(gclk));
	jand g11508(.dina(n11746),.dinb(w_n5259_32[2]),.dout(n11747),.clk(gclk));
	jor g11509(.dina(w_n11451_0[0]),.dinb(n11747),.dout(n11748),.clk(gclk));
	jand g11510(.dina(n11748),.dinb(n11684),.dout(n11749),.clk(gclk));
	jand g11511(.dina(n11749),.dinb(w_n4902_36[2]),.dout(n11750),.clk(gclk));
	jor g11512(.dina(w_n11459_0[0]),.dinb(n11750),.dout(n11751),.clk(gclk));
	jand g11513(.dina(n11751),.dinb(n11683),.dout(n11752),.clk(gclk));
	jand g11514(.dina(n11752),.dinb(w_n4582_33[2]),.dout(n11753),.clk(gclk));
	jor g11515(.dina(w_n11467_0[0]),.dinb(n11753),.dout(n11754),.clk(gclk));
	jand g11516(.dina(n11754),.dinb(n11682),.dout(n11755),.clk(gclk));
	jand g11517(.dina(n11755),.dinb(w_n4249_37[1]),.dout(n11756),.clk(gclk));
	jor g11518(.dina(w_n11475_0[0]),.dinb(n11756),.dout(n11757),.clk(gclk));
	jand g11519(.dina(n11757),.dinb(n11681),.dout(n11758),.clk(gclk));
	jand g11520(.dina(n11758),.dinb(w_n3955_34[1]),.dout(n11759),.clk(gclk));
	jor g11521(.dina(w_n11483_0[0]),.dinb(n11759),.dout(n11760),.clk(gclk));
	jand g11522(.dina(n11760),.dinb(n11680),.dout(n11761),.clk(gclk));
	jand g11523(.dina(n11761),.dinb(w_n3642_37[2]),.dout(n11762),.clk(gclk));
	jor g11524(.dina(n11762),.dinb(w_n11679_0[1]),.dout(n11763),.clk(gclk));
	jand g11525(.dina(n11763),.dinb(n11678),.dout(n11764),.clk(gclk));
	jand g11526(.dina(n11764),.dinb(w_n3368_35[0]),.dout(n11765),.clk(gclk));
	jor g11527(.dina(w_n11498_0[0]),.dinb(n11765),.dout(n11766),.clk(gclk));
	jand g11528(.dina(n11766),.dinb(n11677),.dout(n11767),.clk(gclk));
	jand g11529(.dina(n11767),.dinb(w_n3089_38[1]),.dout(n11768),.clk(gclk));
	jnot g11530(.din(w_n11506_0[0]),.dout(n11769),.clk(gclk));
	jor g11531(.dina(w_n11769_0[1]),.dinb(n11768),.dout(n11770),.clk(gclk));
	jand g11532(.dina(n11770),.dinb(n11676),.dout(n11771),.clk(gclk));
	jand g11533(.dina(n11771),.dinb(w_n2833_36[0]),.dout(n11772),.clk(gclk));
	jor g11534(.dina(w_n11513_0[0]),.dinb(n11772),.dout(n11773),.clk(gclk));
	jand g11535(.dina(n11773),.dinb(n11675),.dout(n11774),.clk(gclk));
	jand g11536(.dina(n11774),.dinb(w_n2572_38[2]),.dout(n11775),.clk(gclk));
	jnot g11537(.din(w_n11521_0[0]),.dout(n11776),.clk(gclk));
	jor g11538(.dina(w_n11776_0[1]),.dinb(n11775),.dout(n11777),.clk(gclk));
	jand g11539(.dina(n11777),.dinb(n11674),.dout(n11778),.clk(gclk));
	jand g11540(.dina(n11778),.dinb(w_n2345_36[2]),.dout(n11779),.clk(gclk));
	jor g11541(.dina(w_n11528_0[0]),.dinb(n11779),.dout(n11780),.clk(gclk));
	jand g11542(.dina(n11780),.dinb(n11673),.dout(n11781),.clk(gclk));
	jand g11543(.dina(n11781),.dinb(w_n2108_39[1]),.dout(n11782),.clk(gclk));
	jor g11544(.dina(w_n11536_0[0]),.dinb(n11782),.dout(n11783),.clk(gclk));
	jand g11545(.dina(n11783),.dinb(n11672),.dout(n11784),.clk(gclk));
	jand g11546(.dina(n11784),.dinb(w_n1912_37[2]),.dout(n11785),.clk(gclk));
	jor g11547(.dina(w_n11544_0[0]),.dinb(n11785),.dout(n11786),.clk(gclk));
	jand g11548(.dina(n11786),.dinb(n11671),.dout(n11787),.clk(gclk));
	jand g11549(.dina(n11787),.dinb(w_n1699_40[0]),.dout(n11788),.clk(gclk));
	jnot g11550(.din(w_n11552_0[0]),.dout(n11789),.clk(gclk));
	jor g11551(.dina(w_n11789_0[1]),.dinb(n11788),.dout(n11790),.clk(gclk));
	jand g11552(.dina(n11790),.dinb(n11670),.dout(n11791),.clk(gclk));
	jand g11553(.dina(n11791),.dinb(w_n1516_38[1]),.dout(n11792),.clk(gclk));
	jor g11554(.dina(w_n11559_0[0]),.dinb(n11792),.dout(n11793),.clk(gclk));
	jand g11555(.dina(n11793),.dinb(n11669),.dout(n11794),.clk(gclk));
	jand g11556(.dina(n11794),.dinb(w_n1332_40[0]),.dout(n11795),.clk(gclk));
	jnot g11557(.din(w_n11567_0[0]),.dout(n11796),.clk(gclk));
	jor g11558(.dina(w_n11796_0[1]),.dinb(n11795),.dout(n11797),.clk(gclk));
	jand g11559(.dina(n11797),.dinb(n11668),.dout(n11798),.clk(gclk));
	jand g11560(.dina(n11798),.dinb(w_n1173_39[0]),.dout(n11799),.clk(gclk));
	jor g11561(.dina(w_n11574_0[0]),.dinb(n11799),.dout(n11800),.clk(gclk));
	jand g11562(.dina(n11800),.dinb(n11667),.dout(n11801),.clk(gclk));
	jand g11563(.dina(n11801),.dinb(w_n1008_41[0]),.dout(n11802),.clk(gclk));
	jnot g11564(.din(w_n11582_0[0]),.dout(n11803),.clk(gclk));
	jor g11565(.dina(w_n11803_0[1]),.dinb(n11802),.dout(n11804),.clk(gclk));
	jand g11566(.dina(n11804),.dinb(n11666),.dout(n11805),.clk(gclk));
	jand g11567(.dina(n11805),.dinb(w_n884_40[0]),.dout(n11806),.clk(gclk));
	jor g11568(.dina(w_n11589_0[0]),.dinb(n11806),.dout(n11807),.clk(gclk));
	jand g11569(.dina(n11807),.dinb(n11665),.dout(n11808),.clk(gclk));
	jand g11570(.dina(n11808),.dinb(w_n743_41[0]),.dout(n11809),.clk(gclk));
	jnot g11571(.din(w_n11597_0[0]),.dout(n11810),.clk(gclk));
	jor g11572(.dina(w_n11810_0[1]),.dinb(n11809),.dout(n11811),.clk(gclk));
	jand g11573(.dina(n11811),.dinb(n11664),.dout(n11812),.clk(gclk));
	jand g11574(.dina(n11812),.dinb(w_n635_41[0]),.dout(n11813),.clk(gclk));
	jnot g11575(.din(w_n11604_0[0]),.dout(n11814),.clk(gclk));
	jor g11576(.dina(w_n11814_0[1]),.dinb(n11813),.dout(n11815),.clk(gclk));
	jand g11577(.dina(n11815),.dinb(n11663),.dout(n11816),.clk(gclk));
	jand g11578(.dina(n11816),.dinb(w_n515_42[0]),.dout(n11817),.clk(gclk));
	jnot g11579(.din(w_n11611_0[0]),.dout(n11818),.clk(gclk));
	jor g11580(.dina(w_n11818_0[1]),.dinb(n11817),.dout(n11819),.clk(gclk));
	jand g11581(.dina(n11819),.dinb(n11662),.dout(n11820),.clk(gclk));
	jand g11582(.dina(n11820),.dinb(w_n443_42[0]),.dout(n11821),.clk(gclk));
	jor g11583(.dina(w_n11618_0[0]),.dinb(n11821),.dout(n11822),.clk(gclk));
	jand g11584(.dina(n11822),.dinb(n11661),.dout(n11823),.clk(gclk));
	jand g11585(.dina(n11823),.dinb(w_n352_42[1]),.dout(n11824),.clk(gclk));
	jor g11586(.dina(w_n11626_0[0]),.dinb(n11824),.dout(n11825),.clk(gclk));
	jand g11587(.dina(n11825),.dinb(n11660),.dout(n11826),.clk(gclk));
	jand g11588(.dina(n11826),.dinb(w_n294_42[2]),.dout(n11827),.clk(gclk));
	jor g11589(.dina(w_n11634_0[0]),.dinb(n11827),.dout(n11828),.clk(gclk));
	jand g11590(.dina(n11828),.dinb(n11659),.dout(n11829),.clk(gclk));
	jand g11591(.dina(n11829),.dinb(w_n239_42[2]),.dout(n11830),.clk(gclk));
	jnot g11592(.din(w_n11642_0[0]),.dout(n11831),.clk(gclk));
	jor g11593(.dina(w_n11831_0[1]),.dinb(n11830),.dout(n11832),.clk(gclk));
	jand g11594(.dina(n11832),.dinb(n11658),.dout(n11833),.clk(gclk));
	jand g11595(.dina(n11833),.dinb(w_n221_43[0]),.dout(n11834),.clk(gclk));
	jor g11596(.dina(w_n11649_0[1]),.dinb(n11834),.dout(n11835),.clk(gclk));
	jand g11597(.dina(n11835),.dinb(n11657),.dout(n11836),.clk(gclk));
	jor g11598(.dina(w_n11836_0[1]),.dinb(n11656),.dout(n11837),.clk(gclk));
	jxor g11599(.dina(w_n11120_0[1]),.dinb(w_n11117_0[2]),.dout(n11838),.clk(gclk));
	jnot g11600(.din(w_n11838_0[1]),.dout(n11839),.clk(gclk));
	jand g11601(.dina(n11839),.dinb(w_asqrt22_22[0]),.dout(n11840),.clk(gclk));
	jor g11602(.dina(w_n11840_0[1]),.dinb(w_n11837_0[1]),.dout(n11841),.clk(gclk));
	jand g11603(.dina(n11841),.dinb(w_n218_18[0]),.dout(n11842),.clk(gclk));
	jand g11604(.dina(w_n11346_0[0]),.dinb(w_n11117_0[1]),.dout(n11843),.clk(gclk));
	jnot g11605(.din(n11843),.dout(n11844),.clk(gclk));
	jand g11606(.dina(w_n11838_0[0]),.dinb(w_asqrt63_32[0]),.dout(n11845),.clk(gclk));
	jand g11607(.dina(w_n11845_0[1]),.dinb(n11844),.dout(n11846),.clk(gclk));
	jor g11608(.dina(w_n11846_0[1]),.dinb(w_n11842_0[1]),.dout(n11847),.clk(gclk));
	jor g11609(.dina(w_n11847_0[1]),.dinb(w_n11654_0[2]),.dout(asqrt_fa_22),.clk(gclk));
	jand g11610(.dina(w_n11652_0[0]),.dinb(w_n11140_0[0]),.dout(n11851),.clk(gclk));
	jnot g11611(.din(w_n11840_0[0]),.dout(n11852),.clk(gclk));
	jand g11612(.dina(n11852),.dinb(w_n11851_0[1]),.dout(n11853),.clk(gclk));
	jor g11613(.dina(n11853),.dinb(w_asqrt63_31[2]),.dout(n11854),.clk(gclk));
	jnot g11614(.din(w_n11846_0[0]),.dout(n11855),.clk(gclk));
	jand g11615(.dina(n11855),.dinb(n11854),.dout(n11856),.clk(gclk));
	jand g11616(.dina(w_n11856_0[1]),.dinb(w_n11653_1[0]),.dout(n11858),.clk(gclk));
	jxor g11617(.dina(w_n11644_0[0]),.dinb(w_n221_42[2]),.dout(n11859),.clk(gclk));
	jor g11618(.dina(n11859),.dinb(w_n11858_45[1]),.dout(n11860),.clk(gclk));
	jxor g11619(.dina(n11860),.dinb(w_n11649_0[0]),.dout(n11861),.clk(gclk));
	jnot g11620(.din(w_n11861_0[1]),.dout(n11862),.clk(gclk));
	jor g11621(.dina(w_n11858_45[0]),.dinb(w_n11142_1[0]),.dout(n11863),.clk(gclk));
	jnot g11622(.din(w_a40_0[2]),.dout(n11864),.clk(gclk));
	jnot g11623(.din(w_a41_0[1]),.dout(n11865),.clk(gclk));
	jand g11624(.dina(w_n11865_0[1]),.dinb(w_n11864_1[2]),.dout(n11866),.clk(gclk));
	jand g11625(.dina(w_n11866_0[2]),.dinb(w_n11142_0[2]),.dout(n11867),.clk(gclk));
	jnot g11626(.din(w_n11867_0[1]),.dout(n11868),.clk(gclk));
	jand g11627(.dina(n11868),.dinb(n11863),.dout(n11869),.clk(gclk));
	jor g11628(.dina(w_n11869_0[2]),.dinb(w_n11347_26[1]),.dout(n11870),.clk(gclk));
	jand g11629(.dina(w_n11869_0[1]),.dinb(w_n11347_26[0]),.dout(n11871),.clk(gclk));
	jor g11630(.dina(w_n11858_44[2]),.dinb(w_a42_1[0]),.dout(n11872),.clk(gclk));
	jand g11631(.dina(n11872),.dinb(w_a43_0[0]),.dout(n11873),.clk(gclk));
	jand g11632(.dina(w_asqrt21_16),.dinb(w_n11144_0[1]),.dout(n11874),.clk(gclk));
	jor g11633(.dina(n11874),.dinb(n11873),.dout(n11875),.clk(gclk));
	jor g11634(.dina(n11875),.dinb(n11871),.dout(n11876),.clk(gclk));
	jand g11635(.dina(n11876),.dinb(w_n11870_0[1]),.dout(n11877),.clk(gclk));
	jor g11636(.dina(w_n11877_0[2]),.dinb(w_n10824_33[0]),.dout(n11878),.clk(gclk));
	jand g11637(.dina(w_n11877_0[1]),.dinb(w_n10824_32[2]),.dout(n11879),.clk(gclk));
	jnot g11638(.din(w_n11144_0[0]),.dout(n11880),.clk(gclk));
	jor g11639(.dina(w_n11858_44[1]),.dinb(n11880),.dout(n11881),.clk(gclk));
	jor g11640(.dina(w_n11845_0[0]),.dinb(w_n11654_0[1]),.dout(n11882),.clk(gclk));
	jor g11641(.dina(n11882),.dinb(w_n11842_0[0]),.dout(n11883),.clk(gclk));
	jor g11642(.dina(n11883),.dinb(w_n11347_25[2]),.dout(n11884),.clk(gclk));
	jand g11643(.dina(n11884),.dinb(w_n11881_0[1]),.dout(n11885),.clk(gclk));
	jxor g11644(.dina(n11885),.dinb(w_n10805_0[1]),.dout(n11886),.clk(gclk));
	jor g11645(.dina(w_n11886_0[2]),.dinb(n11879),.dout(n11887),.clk(gclk));
	jand g11646(.dina(n11887),.dinb(w_n11878_0[1]),.dout(n11888),.clk(gclk));
	jor g11647(.dina(w_n11888_0[2]),.dinb(w_n10328_27[1]),.dout(n11889),.clk(gclk));
	jand g11648(.dina(w_n11888_0[1]),.dinb(w_n10328_27[0]),.dout(n11890),.clk(gclk));
	jxor g11649(.dina(w_n11146_0[0]),.dinb(w_n10824_32[1]),.dout(n11891),.clk(gclk));
	jor g11650(.dina(n11891),.dinb(w_n11858_44[0]),.dout(n11892),.clk(gclk));
	jxor g11651(.dina(n11892),.dinb(w_n11704_0[0]),.dout(n11893),.clk(gclk));
	jnot g11652(.din(w_n11893_0[2]),.dout(n11894),.clk(gclk));
	jor g11653(.dina(n11894),.dinb(n11890),.dout(n11895),.clk(gclk));
	jand g11654(.dina(n11895),.dinb(w_n11889_0[1]),.dout(n11896),.clk(gclk));
	jor g11655(.dina(w_n11896_0[2]),.dinb(w_n9832_33[2]),.dout(n11897),.clk(gclk));
	jand g11656(.dina(w_n11896_0[1]),.dinb(w_n9832_33[1]),.dout(n11898),.clk(gclk));
	jxor g11657(.dina(w_n11351_0[0]),.dinb(w_n10328_26[2]),.dout(n11899),.clk(gclk));
	jor g11658(.dina(n11899),.dinb(w_n11858_43[2]),.dout(n11900),.clk(gclk));
	jxor g11659(.dina(n11900),.dinb(w_n11360_0[0]),.dout(n11901),.clk(gclk));
	jor g11660(.dina(w_n11901_0[2]),.dinb(n11898),.dout(n11902),.clk(gclk));
	jand g11661(.dina(n11902),.dinb(w_n11897_0[1]),.dout(n11903),.clk(gclk));
	jor g11662(.dina(w_n11903_0[2]),.dinb(w_n9369_28[1]),.dout(n11904),.clk(gclk));
	jand g11663(.dina(w_n11903_0[1]),.dinb(w_n9369_28[0]),.dout(n11905),.clk(gclk));
	jxor g11664(.dina(w_n11362_0[0]),.dinb(w_n9832_33[0]),.dout(n11906),.clk(gclk));
	jor g11665(.dina(n11906),.dinb(w_n11858_43[1]),.dout(n11907),.clk(gclk));
	jxor g11666(.dina(n11907),.dinb(w_n11711_0[0]),.dout(n11908),.clk(gclk));
	jnot g11667(.din(w_n11908_0[2]),.dout(n11909),.clk(gclk));
	jor g11668(.dina(n11909),.dinb(n11905),.dout(n11910),.clk(gclk));
	jand g11669(.dina(n11910),.dinb(w_n11904_0[1]),.dout(n11911),.clk(gclk));
	jor g11670(.dina(w_n11911_0[2]),.dinb(w_n8890_34[0]),.dout(n11912),.clk(gclk));
	jand g11671(.dina(w_n11911_0[1]),.dinb(w_n8890_33[2]),.dout(n11913),.clk(gclk));
	jxor g11672(.dina(w_n11369_0[0]),.dinb(w_n9369_27[2]),.dout(n11914),.clk(gclk));
	jor g11673(.dina(n11914),.dinb(w_n11858_43[0]),.dout(n11915),.clk(gclk));
	jxor g11674(.dina(n11915),.dinb(w_n11375_0[0]),.dout(n11916),.clk(gclk));
	jor g11675(.dina(w_n11916_0[2]),.dinb(n11913),.dout(n11917),.clk(gclk));
	jand g11676(.dina(n11917),.dinb(w_n11912_0[1]),.dout(n11918),.clk(gclk));
	jor g11677(.dina(w_n11918_0[2]),.dinb(w_n8449_29[0]),.dout(n11919),.clk(gclk));
	jand g11678(.dina(w_n11918_0[1]),.dinb(w_n8449_28[2]),.dout(n11920),.clk(gclk));
	jxor g11679(.dina(w_n11377_0[0]),.dinb(w_n8890_33[1]),.dout(n11921),.clk(gclk));
	jor g11680(.dina(n11921),.dinb(w_n11858_42[2]),.dout(n11922),.clk(gclk));
	jxor g11681(.dina(n11922),.dinb(w_n11383_0[0]),.dout(n11923),.clk(gclk));
	jor g11682(.dina(w_n11923_0[2]),.dinb(n11920),.dout(n11924),.clk(gclk));
	jand g11683(.dina(n11924),.dinb(w_n11919_0[1]),.dout(n11925),.clk(gclk));
	jor g11684(.dina(w_n11925_0[2]),.dinb(w_n8003_34[2]),.dout(n11926),.clk(gclk));
	jand g11685(.dina(w_n11925_0[1]),.dinb(w_n8003_34[1]),.dout(n11927),.clk(gclk));
	jxor g11686(.dina(w_n11385_0[0]),.dinb(w_n8449_28[1]),.dout(n11928),.clk(gclk));
	jor g11687(.dina(n11928),.dinb(w_n11858_42[1]),.dout(n11929),.clk(gclk));
	jxor g11688(.dina(n11929),.dinb(w_n11391_0[0]),.dout(n11930),.clk(gclk));
	jor g11689(.dina(w_n11930_0[2]),.dinb(n11927),.dout(n11931),.clk(gclk));
	jand g11690(.dina(n11931),.dinb(w_n11926_0[1]),.dout(n11932),.clk(gclk));
	jor g11691(.dina(w_n11932_0[2]),.dinb(w_n7581_30[0]),.dout(n11933),.clk(gclk));
	jand g11692(.dina(w_n11932_0[1]),.dinb(w_n7581_29[2]),.dout(n11934),.clk(gclk));
	jxor g11693(.dina(w_n11393_0[0]),.dinb(w_n8003_34[0]),.dout(n11935),.clk(gclk));
	jor g11694(.dina(n11935),.dinb(w_n11858_42[0]),.dout(n11936),.clk(gclk));
	jxor g11695(.dina(n11936),.dinb(w_n11724_0[0]),.dout(n11937),.clk(gclk));
	jnot g11696(.din(w_n11937_0[2]),.dout(n11938),.clk(gclk));
	jor g11697(.dina(n11938),.dinb(n11934),.dout(n11939),.clk(gclk));
	jand g11698(.dina(n11939),.dinb(w_n11933_0[1]),.dout(n11940),.clk(gclk));
	jor g11699(.dina(w_n11940_0[2]),.dinb(w_n7154_35[0]),.dout(n11941),.clk(gclk));
	jand g11700(.dina(w_n11940_0[1]),.dinb(w_n7154_34[2]),.dout(n11942),.clk(gclk));
	jxor g11701(.dina(w_n11400_0[0]),.dinb(w_n7581_29[1]),.dout(n11943),.clk(gclk));
	jor g11702(.dina(n11943),.dinb(w_n11858_41[2]),.dout(n11944),.clk(gclk));
	jxor g11703(.dina(n11944),.dinb(w_n11406_0[0]),.dout(n11945),.clk(gclk));
	jor g11704(.dina(w_n11945_0[2]),.dinb(n11942),.dout(n11946),.clk(gclk));
	jand g11705(.dina(n11946),.dinb(w_n11941_0[1]),.dout(n11947),.clk(gclk));
	jor g11706(.dina(w_n11947_0[2]),.dinb(w_n6758_30[2]),.dout(n11948),.clk(gclk));
	jand g11707(.dina(w_n11947_0[1]),.dinb(w_n6758_30[1]),.dout(n11949),.clk(gclk));
	jxor g11708(.dina(w_n11408_0[0]),.dinb(w_n7154_34[1]),.dout(n11950),.clk(gclk));
	jor g11709(.dina(n11950),.dinb(w_n11858_41[1]),.dout(n11951),.clk(gclk));
	jxor g11710(.dina(n11951),.dinb(w_n11731_0[0]),.dout(n11952),.clk(gclk));
	jnot g11711(.din(w_n11952_0[2]),.dout(n11953),.clk(gclk));
	jor g11712(.dina(n11953),.dinb(n11949),.dout(n11954),.clk(gclk));
	jand g11713(.dina(n11954),.dinb(w_n11948_0[1]),.dout(n11955),.clk(gclk));
	jor g11714(.dina(w_n11955_0[2]),.dinb(w_n6357_35[1]),.dout(n11956),.clk(gclk));
	jand g11715(.dina(w_n11955_0[1]),.dinb(w_n6357_35[0]),.dout(n11957),.clk(gclk));
	jxor g11716(.dina(w_n11415_0[0]),.dinb(w_n6758_30[0]),.dout(n11958),.clk(gclk));
	jor g11717(.dina(n11958),.dinb(w_n11858_41[0]),.dout(n11959),.clk(gclk));
	jxor g11718(.dina(n11959),.dinb(w_n11421_0[0]),.dout(n11960),.clk(gclk));
	jor g11719(.dina(w_n11960_0[2]),.dinb(n11957),.dout(n11961),.clk(gclk));
	jand g11720(.dina(n11961),.dinb(w_n11956_0[1]),.dout(n11962),.clk(gclk));
	jor g11721(.dina(w_n11962_0[2]),.dinb(w_n5989_31[1]),.dout(n11963),.clk(gclk));
	jand g11722(.dina(w_n11962_0[1]),.dinb(w_n5989_31[0]),.dout(n11964),.clk(gclk));
	jxor g11723(.dina(w_n11423_0[0]),.dinb(w_n6357_34[2]),.dout(n11965),.clk(gclk));
	jor g11724(.dina(n11965),.dinb(w_n11858_40[2]),.dout(n11966),.clk(gclk));
	jxor g11725(.dina(n11966),.dinb(w_n11429_0[0]),.dout(n11967),.clk(gclk));
	jor g11726(.dina(w_n11967_0[2]),.dinb(n11964),.dout(n11968),.clk(gclk));
	jand g11727(.dina(n11968),.dinb(w_n11963_0[1]),.dout(n11969),.clk(gclk));
	jor g11728(.dina(w_n11969_0[2]),.dinb(w_n5606_35[2]),.dout(n11970),.clk(gclk));
	jand g11729(.dina(w_n11969_0[1]),.dinb(w_n5606_35[1]),.dout(n11971),.clk(gclk));
	jxor g11730(.dina(w_n11431_0[0]),.dinb(w_n5989_30[2]),.dout(n11972),.clk(gclk));
	jor g11731(.dina(n11972),.dinb(w_n11858_40[1]),.dout(n11973),.clk(gclk));
	jxor g11732(.dina(n11973),.dinb(w_n11437_0[0]),.dout(n11974),.clk(gclk));
	jor g11733(.dina(w_n11974_0[2]),.dinb(n11971),.dout(n11975),.clk(gclk));
	jand g11734(.dina(n11975),.dinb(w_n11970_0[1]),.dout(n11976),.clk(gclk));
	jor g11735(.dina(w_n11976_0[2]),.dinb(w_n5259_32[1]),.dout(n11977),.clk(gclk));
	jand g11736(.dina(w_n11976_0[1]),.dinb(w_n5259_32[0]),.dout(n11978),.clk(gclk));
	jxor g11737(.dina(w_n11439_0[0]),.dinb(w_n5606_35[0]),.dout(n11979),.clk(gclk));
	jor g11738(.dina(n11979),.dinb(w_n11858_40[0]),.dout(n11980),.clk(gclk));
	jxor g11739(.dina(n11980),.dinb(w_n11744_0[0]),.dout(n11981),.clk(gclk));
	jnot g11740(.din(w_n11981_0[2]),.dout(n11982),.clk(gclk));
	jor g11741(.dina(n11982),.dinb(n11978),.dout(n11983),.clk(gclk));
	jand g11742(.dina(n11983),.dinb(w_n11977_0[1]),.dout(n11984),.clk(gclk));
	jor g11743(.dina(w_n11984_0[2]),.dinb(w_n4902_36[1]),.dout(n11985),.clk(gclk));
	jand g11744(.dina(w_n11984_0[1]),.dinb(w_n4902_36[0]),.dout(n11986),.clk(gclk));
	jxor g11745(.dina(w_n11446_0[0]),.dinb(w_n5259_31[2]),.dout(n11987),.clk(gclk));
	jor g11746(.dina(n11987),.dinb(w_n11858_39[2]),.dout(n11988),.clk(gclk));
	jxor g11747(.dina(n11988),.dinb(w_n11452_0[0]),.dout(n11989),.clk(gclk));
	jor g11748(.dina(w_n11989_0[2]),.dinb(n11986),.dout(n11990),.clk(gclk));
	jand g11749(.dina(n11990),.dinb(w_n11985_0[1]),.dout(n11991),.clk(gclk));
	jor g11750(.dina(w_n11991_0[2]),.dinb(w_n4582_33[1]),.dout(n11992),.clk(gclk));
	jand g11751(.dina(w_n11991_0[1]),.dinb(w_n4582_33[0]),.dout(n11993),.clk(gclk));
	jxor g11752(.dina(w_n11454_0[0]),.dinb(w_n4902_35[2]),.dout(n11994),.clk(gclk));
	jor g11753(.dina(n11994),.dinb(w_n11858_39[1]),.dout(n11995),.clk(gclk));
	jxor g11754(.dina(n11995),.dinb(w_n11460_0[0]),.dout(n11996),.clk(gclk));
	jor g11755(.dina(w_n11996_0[2]),.dinb(n11993),.dout(n11997),.clk(gclk));
	jand g11756(.dina(n11997),.dinb(w_n11992_0[1]),.dout(n11998),.clk(gclk));
	jor g11757(.dina(w_n11998_0[2]),.dinb(w_n4249_37[0]),.dout(n11999),.clk(gclk));
	jand g11758(.dina(w_n11998_0[1]),.dinb(w_n4249_36[2]),.dout(n12000),.clk(gclk));
	jxor g11759(.dina(w_n11462_0[0]),.dinb(w_n4582_32[2]),.dout(n12001),.clk(gclk));
	jor g11760(.dina(n12001),.dinb(w_n11858_39[0]),.dout(n12002),.clk(gclk));
	jxor g11761(.dina(n12002),.dinb(w_n11468_0[0]),.dout(n12003),.clk(gclk));
	jor g11762(.dina(w_n12003_0[2]),.dinb(n12000),.dout(n12004),.clk(gclk));
	jand g11763(.dina(n12004),.dinb(w_n11999_0[1]),.dout(n12005),.clk(gclk));
	jor g11764(.dina(w_n12005_0[2]),.dinb(w_n3955_34[0]),.dout(n12006),.clk(gclk));
	jand g11765(.dina(w_n12005_0[1]),.dinb(w_n3955_33[2]),.dout(n12007),.clk(gclk));
	jxor g11766(.dina(w_n11470_0[0]),.dinb(w_n4249_36[1]),.dout(n12008),.clk(gclk));
	jor g11767(.dina(n12008),.dinb(w_n11858_38[2]),.dout(n12009),.clk(gclk));
	jxor g11768(.dina(n12009),.dinb(w_n11476_0[0]),.dout(n12010),.clk(gclk));
	jor g11769(.dina(w_n12010_0[2]),.dinb(n12007),.dout(n12011),.clk(gclk));
	jand g11770(.dina(n12011),.dinb(w_n12006_0[1]),.dout(n12012),.clk(gclk));
	jor g11771(.dina(w_n12012_0[2]),.dinb(w_n3642_37[1]),.dout(n12013),.clk(gclk));
	jand g11772(.dina(w_n12012_0[1]),.dinb(w_n3642_37[0]),.dout(n12014),.clk(gclk));
	jxor g11773(.dina(w_n11478_0[0]),.dinb(w_n3955_33[1]),.dout(n12015),.clk(gclk));
	jor g11774(.dina(n12015),.dinb(w_n11858_38[1]),.dout(n12016),.clk(gclk));
	jxor g11775(.dina(n12016),.dinb(w_n11484_0[0]),.dout(n12017),.clk(gclk));
	jor g11776(.dina(w_n12017_0[2]),.dinb(n12014),.dout(n12018),.clk(gclk));
	jand g11777(.dina(n12018),.dinb(w_n12013_0[1]),.dout(n12019),.clk(gclk));
	jor g11778(.dina(w_n12019_0[2]),.dinb(w_n3368_34[2]),.dout(n12020),.clk(gclk));
	jxor g11779(.dina(w_n11486_0[0]),.dinb(w_n3642_36[2]),.dout(n12021),.clk(gclk));
	jor g11780(.dina(n12021),.dinb(w_n11858_38[0]),.dout(n12022),.clk(gclk));
	jxor g11781(.dina(n12022),.dinb(w_n11679_0[0]),.dout(n12023),.clk(gclk));
	jnot g11782(.din(w_n12023_0[2]),.dout(n12024),.clk(gclk));
	jand g11783(.dina(w_n12019_0[1]),.dinb(w_n3368_34[1]),.dout(n12025),.clk(gclk));
	jor g11784(.dina(n12025),.dinb(n12024),.dout(n12026),.clk(gclk));
	jand g11785(.dina(n12026),.dinb(w_n12020_0[1]),.dout(n12027),.clk(gclk));
	jor g11786(.dina(w_n12027_0[2]),.dinb(w_n3089_38[0]),.dout(n12028),.clk(gclk));
	jand g11787(.dina(w_n12027_0[1]),.dinb(w_n3089_37[2]),.dout(n12029),.clk(gclk));
	jxor g11788(.dina(w_n11493_0[0]),.dinb(w_n3368_34[0]),.dout(n12030),.clk(gclk));
	jor g11789(.dina(n12030),.dinb(w_n11858_37[2]),.dout(n12031),.clk(gclk));
	jxor g11790(.dina(n12031),.dinb(w_n11499_0[0]),.dout(n12032),.clk(gclk));
	jor g11791(.dina(w_n12032_0[2]),.dinb(n12029),.dout(n12033),.clk(gclk));
	jand g11792(.dina(n12033),.dinb(w_n12028_0[1]),.dout(n12034),.clk(gclk));
	jor g11793(.dina(w_n12034_0[2]),.dinb(w_n2833_35[2]),.dout(n12035),.clk(gclk));
	jand g11794(.dina(w_n12034_0[1]),.dinb(w_n2833_35[1]),.dout(n12036),.clk(gclk));
	jxor g11795(.dina(w_n11501_0[0]),.dinb(w_n3089_37[1]),.dout(n12037),.clk(gclk));
	jor g11796(.dina(n12037),.dinb(w_n11858_37[1]),.dout(n12038),.clk(gclk));
	jxor g11797(.dina(n12038),.dinb(w_n11769_0[0]),.dout(n12039),.clk(gclk));
	jnot g11798(.din(w_n12039_0[2]),.dout(n12040),.clk(gclk));
	jor g11799(.dina(n12040),.dinb(n12036),.dout(n12041),.clk(gclk));
	jand g11800(.dina(n12041),.dinb(w_n12035_0[1]),.dout(n12042),.clk(gclk));
	jor g11801(.dina(w_n12042_0[2]),.dinb(w_n2572_38[1]),.dout(n12043),.clk(gclk));
	jand g11802(.dina(w_n12042_0[1]),.dinb(w_n2572_38[0]),.dout(n12044),.clk(gclk));
	jxor g11803(.dina(w_n11508_0[0]),.dinb(w_n2833_35[0]),.dout(n12045),.clk(gclk));
	jor g11804(.dina(n12045),.dinb(w_n11858_37[0]),.dout(n12046),.clk(gclk));
	jxor g11805(.dina(n12046),.dinb(w_n11514_0[0]),.dout(n12047),.clk(gclk));
	jor g11806(.dina(w_n12047_0[2]),.dinb(n12044),.dout(n12048),.clk(gclk));
	jand g11807(.dina(n12048),.dinb(w_n12043_0[1]),.dout(n12049),.clk(gclk));
	jor g11808(.dina(w_n12049_0[2]),.dinb(w_n2345_36[1]),.dout(n12050),.clk(gclk));
	jand g11809(.dina(w_n12049_0[1]),.dinb(w_n2345_36[0]),.dout(n12051),.clk(gclk));
	jxor g11810(.dina(w_n11516_0[0]),.dinb(w_n2572_37[2]),.dout(n12052),.clk(gclk));
	jor g11811(.dina(n12052),.dinb(w_n11858_36[2]),.dout(n12053),.clk(gclk));
	jxor g11812(.dina(n12053),.dinb(w_n11776_0[0]),.dout(n12054),.clk(gclk));
	jnot g11813(.din(w_n12054_0[2]),.dout(n12055),.clk(gclk));
	jor g11814(.dina(n12055),.dinb(n12051),.dout(n12056),.clk(gclk));
	jand g11815(.dina(n12056),.dinb(w_n12050_0[1]),.dout(n12057),.clk(gclk));
	jor g11816(.dina(w_n12057_0[2]),.dinb(w_n2108_39[0]),.dout(n12058),.clk(gclk));
	jand g11817(.dina(w_n12057_0[1]),.dinb(w_n2108_38[2]),.dout(n12059),.clk(gclk));
	jxor g11818(.dina(w_n11523_0[0]),.dinb(w_n2345_35[2]),.dout(n12060),.clk(gclk));
	jor g11819(.dina(n12060),.dinb(w_n11858_36[1]),.dout(n12061),.clk(gclk));
	jxor g11820(.dina(n12061),.dinb(w_n11529_0[0]),.dout(n12062),.clk(gclk));
	jor g11821(.dina(w_n12062_0[2]),.dinb(n12059),.dout(n12063),.clk(gclk));
	jand g11822(.dina(n12063),.dinb(w_n12058_0[1]),.dout(n12064),.clk(gclk));
	jor g11823(.dina(w_n12064_0[2]),.dinb(w_n1912_37[1]),.dout(n12065),.clk(gclk));
	jand g11824(.dina(w_n12064_0[1]),.dinb(w_n1912_37[0]),.dout(n12066),.clk(gclk));
	jxor g11825(.dina(w_n11531_0[0]),.dinb(w_n2108_38[1]),.dout(n12067),.clk(gclk));
	jor g11826(.dina(n12067),.dinb(w_n11858_36[0]),.dout(n12068),.clk(gclk));
	jxor g11827(.dina(n12068),.dinb(w_n11537_0[0]),.dout(n12069),.clk(gclk));
	jor g11828(.dina(w_n12069_0[2]),.dinb(n12066),.dout(n12070),.clk(gclk));
	jand g11829(.dina(n12070),.dinb(w_n12065_0[1]),.dout(n12071),.clk(gclk));
	jor g11830(.dina(w_n12071_0[2]),.dinb(w_n1699_39[2]),.dout(n12072),.clk(gclk));
	jand g11831(.dina(w_n12071_0[1]),.dinb(w_n1699_39[1]),.dout(n12073),.clk(gclk));
	jxor g11832(.dina(w_n11539_0[0]),.dinb(w_n1912_36[2]),.dout(n12074),.clk(gclk));
	jor g11833(.dina(n12074),.dinb(w_n11858_35[2]),.dout(n12075),.clk(gclk));
	jxor g11834(.dina(n12075),.dinb(w_n11545_0[0]),.dout(n12076),.clk(gclk));
	jor g11835(.dina(w_n12076_0[2]),.dinb(n12073),.dout(n12077),.clk(gclk));
	jand g11836(.dina(n12077),.dinb(w_n12072_0[1]),.dout(n12078),.clk(gclk));
	jor g11837(.dina(w_n12078_0[2]),.dinb(w_n1516_38[0]),.dout(n12079),.clk(gclk));
	jand g11838(.dina(w_n12078_0[1]),.dinb(w_n1516_37[2]),.dout(n12080),.clk(gclk));
	jxor g11839(.dina(w_n11547_0[0]),.dinb(w_n1699_39[0]),.dout(n12081),.clk(gclk));
	jor g11840(.dina(n12081),.dinb(w_n11858_35[1]),.dout(n12082),.clk(gclk));
	jxor g11841(.dina(n12082),.dinb(w_n11789_0[0]),.dout(n12083),.clk(gclk));
	jnot g11842(.din(w_n12083_0[2]),.dout(n12084),.clk(gclk));
	jor g11843(.dina(n12084),.dinb(n12080),.dout(n12085),.clk(gclk));
	jand g11844(.dina(n12085),.dinb(w_n12079_0[1]),.dout(n12086),.clk(gclk));
	jor g11845(.dina(w_n12086_0[2]),.dinb(w_n1332_39[2]),.dout(n12087),.clk(gclk));
	jand g11846(.dina(w_n12086_0[1]),.dinb(w_n1332_39[1]),.dout(n12088),.clk(gclk));
	jxor g11847(.dina(w_n11554_0[0]),.dinb(w_n1516_37[1]),.dout(n12089),.clk(gclk));
	jor g11848(.dina(n12089),.dinb(w_n11858_35[0]),.dout(n12090),.clk(gclk));
	jxor g11849(.dina(n12090),.dinb(w_n11560_0[0]),.dout(n12091),.clk(gclk));
	jor g11850(.dina(w_n12091_0[2]),.dinb(n12088),.dout(n12092),.clk(gclk));
	jand g11851(.dina(n12092),.dinb(w_n12087_0[1]),.dout(n12093),.clk(gclk));
	jor g11852(.dina(w_n12093_0[2]),.dinb(w_n1173_38[2]),.dout(n12094),.clk(gclk));
	jand g11853(.dina(w_n12093_0[1]),.dinb(w_n1173_38[1]),.dout(n12095),.clk(gclk));
	jxor g11854(.dina(w_n11562_0[0]),.dinb(w_n1332_39[0]),.dout(n12096),.clk(gclk));
	jor g11855(.dina(n12096),.dinb(w_n11858_34[2]),.dout(n12097),.clk(gclk));
	jxor g11856(.dina(n12097),.dinb(w_n11796_0[0]),.dout(n12098),.clk(gclk));
	jnot g11857(.din(w_n12098_0[2]),.dout(n12099),.clk(gclk));
	jor g11858(.dina(n12099),.dinb(n12095),.dout(n12100),.clk(gclk));
	jand g11859(.dina(n12100),.dinb(w_n12094_0[1]),.dout(n12101),.clk(gclk));
	jor g11860(.dina(w_n12101_0[2]),.dinb(w_n1008_40[2]),.dout(n12102),.clk(gclk));
	jand g11861(.dina(w_n12101_0[1]),.dinb(w_n1008_40[1]),.dout(n12103),.clk(gclk));
	jxor g11862(.dina(w_n11569_0[0]),.dinb(w_n1173_38[0]),.dout(n12104),.clk(gclk));
	jor g11863(.dina(n12104),.dinb(w_n11858_34[1]),.dout(n12105),.clk(gclk));
	jxor g11864(.dina(n12105),.dinb(w_n11575_0[0]),.dout(n12106),.clk(gclk));
	jor g11865(.dina(w_n12106_0[2]),.dinb(n12103),.dout(n12107),.clk(gclk));
	jand g11866(.dina(n12107),.dinb(w_n12102_0[1]),.dout(n12108),.clk(gclk));
	jor g11867(.dina(w_n12108_0[2]),.dinb(w_n884_39[2]),.dout(n12109),.clk(gclk));
	jand g11868(.dina(w_n12108_0[1]),.dinb(w_n884_39[1]),.dout(n12110),.clk(gclk));
	jxor g11869(.dina(w_n11577_0[0]),.dinb(w_n1008_40[0]),.dout(n12111),.clk(gclk));
	jor g11870(.dina(n12111),.dinb(w_n11858_34[0]),.dout(n12112),.clk(gclk));
	jxor g11871(.dina(n12112),.dinb(w_n11803_0[0]),.dout(n12113),.clk(gclk));
	jnot g11872(.din(w_n12113_0[2]),.dout(n12114),.clk(gclk));
	jor g11873(.dina(n12114),.dinb(n12110),.dout(n12115),.clk(gclk));
	jand g11874(.dina(n12115),.dinb(w_n12109_0[1]),.dout(n12116),.clk(gclk));
	jor g11875(.dina(w_n12116_0[2]),.dinb(w_n743_40[2]),.dout(n12117),.clk(gclk));
	jand g11876(.dina(w_n12116_0[1]),.dinb(w_n743_40[1]),.dout(n12118),.clk(gclk));
	jxor g11877(.dina(w_n11584_0[0]),.dinb(w_n884_39[0]),.dout(n12119),.clk(gclk));
	jor g11878(.dina(n12119),.dinb(w_n11858_33[2]),.dout(n12120),.clk(gclk));
	jxor g11879(.dina(n12120),.dinb(w_n11590_0[0]),.dout(n12121),.clk(gclk));
	jor g11880(.dina(w_n12121_0[2]),.dinb(n12118),.dout(n12122),.clk(gclk));
	jand g11881(.dina(n12122),.dinb(w_n12117_0[1]),.dout(n12123),.clk(gclk));
	jor g11882(.dina(w_n12123_0[2]),.dinb(w_n635_40[2]),.dout(n12124),.clk(gclk));
	jand g11883(.dina(w_n12123_0[1]),.dinb(w_n635_40[1]),.dout(n12125),.clk(gclk));
	jxor g11884(.dina(w_n11592_0[0]),.dinb(w_n743_40[0]),.dout(n12126),.clk(gclk));
	jor g11885(.dina(n12126),.dinb(w_n11858_33[1]),.dout(n12127),.clk(gclk));
	jxor g11886(.dina(n12127),.dinb(w_n11810_0[0]),.dout(n12128),.clk(gclk));
	jnot g11887(.din(w_n12128_0[2]),.dout(n12129),.clk(gclk));
	jor g11888(.dina(n12129),.dinb(n12125),.dout(n12130),.clk(gclk));
	jand g11889(.dina(n12130),.dinb(w_n12124_0[1]),.dout(n12131),.clk(gclk));
	jor g11890(.dina(w_n12131_0[2]),.dinb(w_n515_41[2]),.dout(n12132),.clk(gclk));
	jand g11891(.dina(w_n12131_0[1]),.dinb(w_n515_41[1]),.dout(n12133),.clk(gclk));
	jxor g11892(.dina(w_n11599_0[0]),.dinb(w_n635_40[0]),.dout(n12134),.clk(gclk));
	jor g11893(.dina(n12134),.dinb(w_n11858_33[0]),.dout(n12135),.clk(gclk));
	jxor g11894(.dina(n12135),.dinb(w_n11814_0[0]),.dout(n12136),.clk(gclk));
	jnot g11895(.din(w_n12136_0[2]),.dout(n12137),.clk(gclk));
	jor g11896(.dina(n12137),.dinb(n12133),.dout(n12138),.clk(gclk));
	jand g11897(.dina(n12138),.dinb(w_n12132_0[1]),.dout(n12139),.clk(gclk));
	jor g11898(.dina(w_n12139_0[2]),.dinb(w_n443_41[2]),.dout(n12140),.clk(gclk));
	jand g11899(.dina(w_n12139_0[1]),.dinb(w_n443_41[1]),.dout(n12141),.clk(gclk));
	jxor g11900(.dina(w_n11606_0[0]),.dinb(w_n515_41[0]),.dout(n12142),.clk(gclk));
	jor g11901(.dina(n12142),.dinb(w_n11858_32[2]),.dout(n12143),.clk(gclk));
	jxor g11902(.dina(n12143),.dinb(w_n11818_0[0]),.dout(n12144),.clk(gclk));
	jnot g11903(.din(w_n12144_0[2]),.dout(n12145),.clk(gclk));
	jor g11904(.dina(n12145),.dinb(n12141),.dout(n12146),.clk(gclk));
	jand g11905(.dina(n12146),.dinb(w_n12140_0[1]),.dout(n12147),.clk(gclk));
	jor g11906(.dina(w_n12147_0[2]),.dinb(w_n352_42[0]),.dout(n12148),.clk(gclk));
	jand g11907(.dina(w_n12147_0[1]),.dinb(w_n352_41[2]),.dout(n12149),.clk(gclk));
	jxor g11908(.dina(w_n11613_0[0]),.dinb(w_n443_41[0]),.dout(n12150),.clk(gclk));
	jor g11909(.dina(n12150),.dinb(w_n11858_32[1]),.dout(n12151),.clk(gclk));
	jxor g11910(.dina(n12151),.dinb(w_n11619_0[0]),.dout(n12152),.clk(gclk));
	jor g11911(.dina(w_n12152_0[2]),.dinb(n12149),.dout(n12153),.clk(gclk));
	jand g11912(.dina(n12153),.dinb(w_n12148_0[1]),.dout(n12154),.clk(gclk));
	jor g11913(.dina(w_n12154_0[2]),.dinb(w_n294_42[1]),.dout(n12155),.clk(gclk));
	jand g11914(.dina(w_n12154_0[1]),.dinb(w_n294_42[0]),.dout(n12156),.clk(gclk));
	jxor g11915(.dina(w_n11621_0[0]),.dinb(w_n352_41[1]),.dout(n12157),.clk(gclk));
	jor g11916(.dina(n12157),.dinb(w_n11858_32[0]),.dout(n12158),.clk(gclk));
	jxor g11917(.dina(n12158),.dinb(w_n11627_0[0]),.dout(n12159),.clk(gclk));
	jor g11918(.dina(w_n12159_0[2]),.dinb(n12156),.dout(n12160),.clk(gclk));
	jand g11919(.dina(n12160),.dinb(w_n12155_0[1]),.dout(n12161),.clk(gclk));
	jor g11920(.dina(w_n12161_0[2]),.dinb(w_n239_42[1]),.dout(n12162),.clk(gclk));
	jand g11921(.dina(w_n12161_0[1]),.dinb(w_n239_42[0]),.dout(n12163),.clk(gclk));
	jxor g11922(.dina(w_n11629_0[0]),.dinb(w_n294_41[2]),.dout(n12164),.clk(gclk));
	jor g11923(.dina(n12164),.dinb(w_n11858_31[2]),.dout(n12165),.clk(gclk));
	jxor g11924(.dina(n12165),.dinb(w_n11635_0[0]),.dout(n12166),.clk(gclk));
	jor g11925(.dina(w_n12166_0[2]),.dinb(n12163),.dout(n12167),.clk(gclk));
	jand g11926(.dina(n12167),.dinb(w_n12162_0[1]),.dout(n12168),.clk(gclk));
	jor g11927(.dina(w_n12168_0[2]),.dinb(w_n221_42[1]),.dout(n12169),.clk(gclk));
	jand g11928(.dina(w_n12168_0[1]),.dinb(w_n221_42[0]),.dout(n12170),.clk(gclk));
	jxor g11929(.dina(w_n11637_0[0]),.dinb(w_n239_41[2]),.dout(n12171),.clk(gclk));
	jor g11930(.dina(n12171),.dinb(w_n11858_31[1]),.dout(n12172),.clk(gclk));
	jxor g11931(.dina(n12172),.dinb(w_n11831_0[0]),.dout(n12173),.clk(gclk));
	jnot g11932(.din(w_n12173_0[2]),.dout(n12174),.clk(gclk));
	jor g11933(.dina(n12174),.dinb(n12170),.dout(n12175),.clk(gclk));
	jand g11934(.dina(n12175),.dinb(w_n12169_0[1]),.dout(n12176),.clk(gclk));
	jand g11935(.dina(w_n12176_0[2]),.dinb(w_n11862_0[2]),.dout(n12177),.clk(gclk));
	jand g11936(.dina(w_n11847_0[0]),.dinb(w_n11851_0[0]),.dout(n12179),.clk(gclk));
	jor g11937(.dina(w_n12176_0[1]),.dinb(w_n11862_0[1]),.dout(n12180),.clk(gclk));
	jor g11938(.dina(w_n12180_0[1]),.dinb(w_n11654_0[0]),.dout(n12181),.clk(gclk));
	jor g11939(.dina(n12181),.dinb(w_n12179_0[1]),.dout(n12182),.clk(gclk));
	jand g11940(.dina(n12182),.dinb(w_n218_17[2]),.dout(n12183),.clk(gclk));
	jand g11941(.dina(w_n11856_0[0]),.dinb(w_n11836_0[0]),.dout(n12184),.clk(gclk));
	jand g11942(.dina(w_n11837_0[0]),.dinb(w_asqrt63_31[1]),.dout(n12185),.clk(gclk));
	jand g11943(.dina(n12185),.dinb(w_n11653_0[2]),.dout(n12186),.clk(gclk));
	jnot g11944(.din(n12186),.dout(n12187),.clk(gclk));
	jor g11945(.dina(w_n12187_0[1]),.dinb(n12184),.dout(n12188),.clk(gclk));
	jnot g11946(.din(w_n12188_0[1]),.dout(n12189),.clk(gclk));
	jor g11947(.dina(n12189),.dinb(n12183),.dout(n12190),.clk(gclk));
	jor g11948(.dina(w_n12190_0[1]),.dinb(w_n12177_0[2]),.dout(asqrt_fa_21),.clk(gclk));
	jxor g11949(.dina(w_n12168_0[0]),.dinb(w_n221_41[2]),.dout(n12193),.clk(gclk));
	jand g11950(.dina(n12193),.dinb(w_asqrt20_35),.dout(n12194),.clk(gclk));
	jxor g11951(.dina(n12194),.dinb(w_n12173_0[1]),.dout(n12195),.clk(gclk));
	jnot g11952(.din(w_a38_0[2]),.dout(n12196),.clk(gclk));
	jnot g11953(.din(w_a39_0[1]),.dout(n12197),.clk(gclk));
	jand g11954(.dina(w_n12197_0[1]),.dinb(w_n12196_1[2]),.dout(n12198),.clk(gclk));
	jand g11955(.dina(w_n12198_0[2]),.dinb(w_n11864_1[1]),.dout(n12199),.clk(gclk));
	jand g11956(.dina(w_asqrt20_34[2]),.dinb(w_a40_0[1]),.dout(n12200),.clk(gclk));
	jor g11957(.dina(n12200),.dinb(w_n12199_0[1]),.dout(n12201),.clk(gclk));
	jand g11958(.dina(w_n12201_0[2]),.dinb(w_asqrt21_15[2]),.dout(n12202),.clk(gclk));
	jor g11959(.dina(w_n12201_0[1]),.dinb(w_asqrt21_15[1]),.dout(n12203),.clk(gclk));
	jand g11960(.dina(w_asqrt20_34[1]),.dinb(w_n11864_1[0]),.dout(n12204),.clk(gclk));
	jor g11961(.dina(n12204),.dinb(w_n11865_0[0]),.dout(n12205),.clk(gclk));
	jnot g11962(.din(w_n11866_0[1]),.dout(n12206),.clk(gclk));
	jnot g11963(.din(w_n12177_0[1]),.dout(n12207),.clk(gclk));
	jnot g11964(.din(w_n12179_0[0]),.dout(n12209),.clk(gclk));
	jnot g11965(.din(w_n12169_0[0]),.dout(n12210),.clk(gclk));
	jnot g11966(.din(w_n12162_0[0]),.dout(n12211),.clk(gclk));
	jnot g11967(.din(w_n12155_0[0]),.dout(n12212),.clk(gclk));
	jnot g11968(.din(w_n12148_0[0]),.dout(n12213),.clk(gclk));
	jnot g11969(.din(w_n12140_0[0]),.dout(n12214),.clk(gclk));
	jnot g11970(.din(w_n12132_0[0]),.dout(n12215),.clk(gclk));
	jnot g11971(.din(w_n12124_0[0]),.dout(n12216),.clk(gclk));
	jnot g11972(.din(w_n12117_0[0]),.dout(n12217),.clk(gclk));
	jnot g11973(.din(w_n12109_0[0]),.dout(n12218),.clk(gclk));
	jnot g11974(.din(w_n12102_0[0]),.dout(n12219),.clk(gclk));
	jnot g11975(.din(w_n12094_0[0]),.dout(n12220),.clk(gclk));
	jnot g11976(.din(w_n12087_0[0]),.dout(n12221),.clk(gclk));
	jnot g11977(.din(w_n12079_0[0]),.dout(n12222),.clk(gclk));
	jnot g11978(.din(w_n12072_0[0]),.dout(n12223),.clk(gclk));
	jnot g11979(.din(w_n12065_0[0]),.dout(n12224),.clk(gclk));
	jnot g11980(.din(w_n12058_0[0]),.dout(n12225),.clk(gclk));
	jnot g11981(.din(w_n12050_0[0]),.dout(n12226),.clk(gclk));
	jnot g11982(.din(w_n12043_0[0]),.dout(n12227),.clk(gclk));
	jnot g11983(.din(w_n12035_0[0]),.dout(n12228),.clk(gclk));
	jnot g11984(.din(w_n12028_0[0]),.dout(n12229),.clk(gclk));
	jnot g11985(.din(w_n12020_0[0]),.dout(n12230),.clk(gclk));
	jnot g11986(.din(w_n12013_0[0]),.dout(n12231),.clk(gclk));
	jnot g11987(.din(w_n12006_0[0]),.dout(n12232),.clk(gclk));
	jnot g11988(.din(w_n11999_0[0]),.dout(n12233),.clk(gclk));
	jnot g11989(.din(w_n11992_0[0]),.dout(n12234),.clk(gclk));
	jnot g11990(.din(w_n11985_0[0]),.dout(n12235),.clk(gclk));
	jnot g11991(.din(w_n11977_0[0]),.dout(n12236),.clk(gclk));
	jnot g11992(.din(w_n11970_0[0]),.dout(n12237),.clk(gclk));
	jnot g11993(.din(w_n11963_0[0]),.dout(n12238),.clk(gclk));
	jnot g11994(.din(w_n11956_0[0]),.dout(n12239),.clk(gclk));
	jnot g11995(.din(w_n11948_0[0]),.dout(n12240),.clk(gclk));
	jnot g11996(.din(w_n11941_0[0]),.dout(n12241),.clk(gclk));
	jnot g11997(.din(w_n11933_0[0]),.dout(n12242),.clk(gclk));
	jnot g11998(.din(w_n11926_0[0]),.dout(n12243),.clk(gclk));
	jnot g11999(.din(w_n11919_0[0]),.dout(n12244),.clk(gclk));
	jnot g12000(.din(w_n11912_0[0]),.dout(n12245),.clk(gclk));
	jnot g12001(.din(w_n11904_0[0]),.dout(n12246),.clk(gclk));
	jnot g12002(.din(w_n11897_0[0]),.dout(n12247),.clk(gclk));
	jnot g12003(.din(w_n11889_0[0]),.dout(n12248),.clk(gclk));
	jnot g12004(.din(w_n11878_0[0]),.dout(n12249),.clk(gclk));
	jnot g12005(.din(w_n11870_0[0]),.dout(n12250),.clk(gclk));
	jand g12006(.dina(w_asqrt21_15[0]),.dinb(w_a42_0[2]),.dout(n12251),.clk(gclk));
	jor g12007(.dina(w_n11867_0[0]),.dinb(n12251),.dout(n12252),.clk(gclk));
	jor g12008(.dina(n12252),.dinb(w_asqrt22_21[2]),.dout(n12253),.clk(gclk));
	jand g12009(.dina(w_asqrt21_14[2]),.dinb(w_n11142_0[1]),.dout(n12254),.clk(gclk));
	jor g12010(.dina(n12254),.dinb(w_n11143_0[0]),.dout(n12255),.clk(gclk));
	jand g12011(.dina(w_n11881_0[0]),.dinb(n12255),.dout(n12256),.clk(gclk));
	jand g12012(.dina(w_n12256_0[1]),.dinb(n12253),.dout(n12257),.clk(gclk));
	jor g12013(.dina(n12257),.dinb(n12250),.dout(n12258),.clk(gclk));
	jor g12014(.dina(n12258),.dinb(w_asqrt23_15[2]),.dout(n12259),.clk(gclk));
	jnot g12015(.din(w_n11886_0[1]),.dout(n12260),.clk(gclk));
	jand g12016(.dina(n12260),.dinb(n12259),.dout(n12261),.clk(gclk));
	jor g12017(.dina(n12261),.dinb(n12249),.dout(n12262),.clk(gclk));
	jor g12018(.dina(n12262),.dinb(w_asqrt24_21[2]),.dout(n12263),.clk(gclk));
	jand g12019(.dina(w_n11893_0[1]),.dinb(n12263),.dout(n12264),.clk(gclk));
	jor g12020(.dina(n12264),.dinb(n12248),.dout(n12265),.clk(gclk));
	jor g12021(.dina(n12265),.dinb(w_asqrt25_15[2]),.dout(n12266),.clk(gclk));
	jnot g12022(.din(w_n11901_0[1]),.dout(n12267),.clk(gclk));
	jand g12023(.dina(n12267),.dinb(n12266),.dout(n12268),.clk(gclk));
	jor g12024(.dina(n12268),.dinb(n12247),.dout(n12269),.clk(gclk));
	jor g12025(.dina(n12269),.dinb(w_asqrt26_21[2]),.dout(n12270),.clk(gclk));
	jand g12026(.dina(w_n11908_0[1]),.dinb(n12270),.dout(n12271),.clk(gclk));
	jor g12027(.dina(n12271),.dinb(n12246),.dout(n12272),.clk(gclk));
	jor g12028(.dina(n12272),.dinb(w_asqrt27_16[1]),.dout(n12273),.clk(gclk));
	jnot g12029(.din(w_n11916_0[1]),.dout(n12274),.clk(gclk));
	jand g12030(.dina(n12274),.dinb(n12273),.dout(n12275),.clk(gclk));
	jor g12031(.dina(n12275),.dinb(n12245),.dout(n12276),.clk(gclk));
	jor g12032(.dina(n12276),.dinb(w_asqrt28_22[0]),.dout(n12277),.clk(gclk));
	jnot g12033(.din(w_n11923_0[1]),.dout(n12278),.clk(gclk));
	jand g12034(.dina(n12278),.dinb(n12277),.dout(n12279),.clk(gclk));
	jor g12035(.dina(n12279),.dinb(n12244),.dout(n12280),.clk(gclk));
	jor g12036(.dina(n12280),.dinb(w_asqrt29_16[2]),.dout(n12281),.clk(gclk));
	jnot g12037(.din(w_n11930_0[1]),.dout(n12282),.clk(gclk));
	jand g12038(.dina(n12282),.dinb(n12281),.dout(n12283),.clk(gclk));
	jor g12039(.dina(n12283),.dinb(n12243),.dout(n12284),.clk(gclk));
	jor g12040(.dina(n12284),.dinb(w_asqrt30_22[1]),.dout(n12285),.clk(gclk));
	jand g12041(.dina(w_n11937_0[1]),.dinb(n12285),.dout(n12286),.clk(gclk));
	jor g12042(.dina(n12286),.dinb(n12242),.dout(n12287),.clk(gclk));
	jor g12043(.dina(n12287),.dinb(w_asqrt31_17[1]),.dout(n12288),.clk(gclk));
	jnot g12044(.din(w_n11945_0[1]),.dout(n12289),.clk(gclk));
	jand g12045(.dina(n12289),.dinb(n12288),.dout(n12290),.clk(gclk));
	jor g12046(.dina(n12290),.dinb(n12241),.dout(n12291),.clk(gclk));
	jor g12047(.dina(n12291),.dinb(w_asqrt32_22[1]),.dout(n12292),.clk(gclk));
	jand g12048(.dina(w_n11952_0[1]),.dinb(n12292),.dout(n12293),.clk(gclk));
	jor g12049(.dina(n12293),.dinb(n12240),.dout(n12294),.clk(gclk));
	jor g12050(.dina(n12294),.dinb(w_asqrt33_18[0]),.dout(n12295),.clk(gclk));
	jnot g12051(.din(w_n11960_0[1]),.dout(n12296),.clk(gclk));
	jand g12052(.dina(n12296),.dinb(n12295),.dout(n12297),.clk(gclk));
	jor g12053(.dina(n12297),.dinb(n12239),.dout(n12298),.clk(gclk));
	jor g12054(.dina(n12298),.dinb(w_asqrt34_22[2]),.dout(n12299),.clk(gclk));
	jnot g12055(.din(w_n11967_0[1]),.dout(n12300),.clk(gclk));
	jand g12056(.dina(n12300),.dinb(n12299),.dout(n12301),.clk(gclk));
	jor g12057(.dina(n12301),.dinb(n12238),.dout(n12302),.clk(gclk));
	jor g12058(.dina(n12302),.dinb(w_asqrt35_18[2]),.dout(n12303),.clk(gclk));
	jnot g12059(.din(w_n11974_0[1]),.dout(n12304),.clk(gclk));
	jand g12060(.dina(n12304),.dinb(n12303),.dout(n12305),.clk(gclk));
	jor g12061(.dina(n12305),.dinb(n12237),.dout(n12306),.clk(gclk));
	jor g12062(.dina(n12306),.dinb(w_asqrt36_22[2]),.dout(n12307),.clk(gclk));
	jand g12063(.dina(w_n11981_0[1]),.dinb(n12307),.dout(n12308),.clk(gclk));
	jor g12064(.dina(n12308),.dinb(n12236),.dout(n12309),.clk(gclk));
	jor g12065(.dina(n12309),.dinb(w_asqrt37_19[0]),.dout(n12310),.clk(gclk));
	jnot g12066(.din(w_n11989_0[1]),.dout(n12311),.clk(gclk));
	jand g12067(.dina(n12311),.dinb(n12310),.dout(n12312),.clk(gclk));
	jor g12068(.dina(n12312),.dinb(n12235),.dout(n12313),.clk(gclk));
	jor g12069(.dina(n12313),.dinb(w_asqrt38_23[0]),.dout(n12314),.clk(gclk));
	jnot g12070(.din(w_n11996_0[1]),.dout(n12315),.clk(gclk));
	jand g12071(.dina(n12315),.dinb(n12314),.dout(n12316),.clk(gclk));
	jor g12072(.dina(n12316),.dinb(n12234),.dout(n12317),.clk(gclk));
	jor g12073(.dina(n12317),.dinb(w_asqrt39_19[2]),.dout(n12318),.clk(gclk));
	jnot g12074(.din(w_n12003_0[1]),.dout(n12319),.clk(gclk));
	jand g12075(.dina(n12319),.dinb(n12318),.dout(n12320),.clk(gclk));
	jor g12076(.dina(n12320),.dinb(n12233),.dout(n12321),.clk(gclk));
	jor g12077(.dina(n12321),.dinb(w_asqrt40_23[0]),.dout(n12322),.clk(gclk));
	jnot g12078(.din(w_n12010_0[1]),.dout(n12323),.clk(gclk));
	jand g12079(.dina(n12323),.dinb(n12322),.dout(n12324),.clk(gclk));
	jor g12080(.dina(n12324),.dinb(n12232),.dout(n12325),.clk(gclk));
	jor g12081(.dina(n12325),.dinb(w_asqrt41_20[0]),.dout(n12326),.clk(gclk));
	jnot g12082(.din(w_n12017_0[1]),.dout(n12327),.clk(gclk));
	jand g12083(.dina(n12327),.dinb(n12326),.dout(n12328),.clk(gclk));
	jor g12084(.dina(n12328),.dinb(n12231),.dout(n12329),.clk(gclk));
	jor g12085(.dina(n12329),.dinb(w_asqrt42_23[1]),.dout(n12330),.clk(gclk));
	jand g12086(.dina(n12330),.dinb(w_n12023_0[1]),.dout(n12331),.clk(gclk));
	jor g12087(.dina(n12331),.dinb(n12230),.dout(n12332),.clk(gclk));
	jor g12088(.dina(n12332),.dinb(w_asqrt43_20[1]),.dout(n12333),.clk(gclk));
	jnot g12089(.din(w_n12032_0[1]),.dout(n12334),.clk(gclk));
	jand g12090(.dina(n12334),.dinb(n12333),.dout(n12335),.clk(gclk));
	jor g12091(.dina(n12335),.dinb(n12229),.dout(n12336),.clk(gclk));
	jor g12092(.dina(n12336),.dinb(w_asqrt44_23[1]),.dout(n12337),.clk(gclk));
	jand g12093(.dina(w_n12039_0[1]),.dinb(n12337),.dout(n12338),.clk(gclk));
	jor g12094(.dina(n12338),.dinb(n12228),.dout(n12339),.clk(gclk));
	jor g12095(.dina(n12339),.dinb(w_asqrt45_21[0]),.dout(n12340),.clk(gclk));
	jnot g12096(.din(w_n12047_0[1]),.dout(n12341),.clk(gclk));
	jand g12097(.dina(n12341),.dinb(n12340),.dout(n12342),.clk(gclk));
	jor g12098(.dina(n12342),.dinb(n12227),.dout(n12343),.clk(gclk));
	jor g12099(.dina(n12343),.dinb(w_asqrt46_23[1]),.dout(n12344),.clk(gclk));
	jand g12100(.dina(w_n12054_0[1]),.dinb(n12344),.dout(n12345),.clk(gclk));
	jor g12101(.dina(n12345),.dinb(n12226),.dout(n12346),.clk(gclk));
	jor g12102(.dina(n12346),.dinb(w_asqrt47_21[2]),.dout(n12347),.clk(gclk));
	jnot g12103(.din(w_n12062_0[1]),.dout(n12348),.clk(gclk));
	jand g12104(.dina(n12348),.dinb(n12347),.dout(n12349),.clk(gclk));
	jor g12105(.dina(n12349),.dinb(n12225),.dout(n12350),.clk(gclk));
	jor g12106(.dina(n12350),.dinb(w_asqrt48_23[2]),.dout(n12351),.clk(gclk));
	jnot g12107(.din(w_n12069_0[1]),.dout(n12352),.clk(gclk));
	jand g12108(.dina(n12352),.dinb(n12351),.dout(n12353),.clk(gclk));
	jor g12109(.dina(n12353),.dinb(n12224),.dout(n12354),.clk(gclk));
	jor g12110(.dina(n12354),.dinb(w_asqrt49_22[0]),.dout(n12355),.clk(gclk));
	jnot g12111(.din(w_n12076_0[1]),.dout(n12356),.clk(gclk));
	jand g12112(.dina(n12356),.dinb(n12355),.dout(n12357),.clk(gclk));
	jor g12113(.dina(n12357),.dinb(n12223),.dout(n12358),.clk(gclk));
	jor g12114(.dina(n12358),.dinb(w_asqrt50_24[0]),.dout(n12359),.clk(gclk));
	jand g12115(.dina(w_n12083_0[1]),.dinb(n12359),.dout(n12360),.clk(gclk));
	jor g12116(.dina(n12360),.dinb(n12222),.dout(n12361),.clk(gclk));
	jor g12117(.dina(n12361),.dinb(w_asqrt51_22[1]),.dout(n12362),.clk(gclk));
	jnot g12118(.din(w_n12091_0[1]),.dout(n12363),.clk(gclk));
	jand g12119(.dina(n12363),.dinb(n12362),.dout(n12364),.clk(gclk));
	jor g12120(.dina(n12364),.dinb(n12221),.dout(n12365),.clk(gclk));
	jor g12121(.dina(n12365),.dinb(w_asqrt52_24[0]),.dout(n12366),.clk(gclk));
	jand g12122(.dina(w_n12098_0[1]),.dinb(n12366),.dout(n12367),.clk(gclk));
	jor g12123(.dina(n12367),.dinb(n12220),.dout(n12368),.clk(gclk));
	jor g12124(.dina(n12368),.dinb(w_asqrt53_23[0]),.dout(n12369),.clk(gclk));
	jnot g12125(.din(w_n12106_0[1]),.dout(n12370),.clk(gclk));
	jand g12126(.dina(n12370),.dinb(n12369),.dout(n12371),.clk(gclk));
	jor g12127(.dina(n12371),.dinb(n12219),.dout(n12372),.clk(gclk));
	jor g12128(.dina(n12372),.dinb(w_asqrt54_24[0]),.dout(n12373),.clk(gclk));
	jand g12129(.dina(w_n12113_0[1]),.dinb(n12373),.dout(n12374),.clk(gclk));
	jor g12130(.dina(n12374),.dinb(n12218),.dout(n12375),.clk(gclk));
	jor g12131(.dina(n12375),.dinb(w_asqrt55_23[1]),.dout(n12376),.clk(gclk));
	jnot g12132(.din(w_n12121_0[1]),.dout(n12377),.clk(gclk));
	jand g12133(.dina(n12377),.dinb(n12376),.dout(n12378),.clk(gclk));
	jor g12134(.dina(n12378),.dinb(n12217),.dout(n12379),.clk(gclk));
	jor g12135(.dina(n12379),.dinb(w_asqrt56_24[1]),.dout(n12380),.clk(gclk));
	jand g12136(.dina(w_n12128_0[1]),.dinb(n12380),.dout(n12381),.clk(gclk));
	jor g12137(.dina(n12381),.dinb(n12216),.dout(n12382),.clk(gclk));
	jor g12138(.dina(n12382),.dinb(w_asqrt57_24[0]),.dout(n12383),.clk(gclk));
	jand g12139(.dina(w_n12136_0[1]),.dinb(n12383),.dout(n12384),.clk(gclk));
	jor g12140(.dina(n12384),.dinb(n12215),.dout(n12385),.clk(gclk));
	jor g12141(.dina(n12385),.dinb(w_asqrt58_24[2]),.dout(n12386),.clk(gclk));
	jand g12142(.dina(w_n12144_0[1]),.dinb(n12386),.dout(n12387),.clk(gclk));
	jor g12143(.dina(n12387),.dinb(n12214),.dout(n12388),.clk(gclk));
	jor g12144(.dina(n12388),.dinb(w_asqrt59_24[1]),.dout(n12389),.clk(gclk));
	jnot g12145(.din(w_n12152_0[1]),.dout(n12390),.clk(gclk));
	jand g12146(.dina(n12390),.dinb(n12389),.dout(n12391),.clk(gclk));
	jor g12147(.dina(n12391),.dinb(n12213),.dout(n12392),.clk(gclk));
	jor g12148(.dina(n12392),.dinb(w_asqrt60_24[2]),.dout(n12393),.clk(gclk));
	jnot g12149(.din(w_n12159_0[1]),.dout(n12394),.clk(gclk));
	jand g12150(.dina(n12394),.dinb(n12393),.dout(n12395),.clk(gclk));
	jor g12151(.dina(n12395),.dinb(n12212),.dout(n12396),.clk(gclk));
	jor g12152(.dina(n12396),.dinb(w_asqrt61_24[2]),.dout(n12397),.clk(gclk));
	jnot g12153(.din(w_n12166_0[1]),.dout(n12398),.clk(gclk));
	jand g12154(.dina(n12398),.dinb(n12397),.dout(n12399),.clk(gclk));
	jor g12155(.dina(n12399),.dinb(n12211),.dout(n12400),.clk(gclk));
	jor g12156(.dina(n12400),.dinb(w_asqrt62_24[2]),.dout(n12401),.clk(gclk));
	jand g12157(.dina(w_n12173_0[0]),.dinb(n12401),.dout(n12402),.clk(gclk));
	jor g12158(.dina(n12402),.dinb(n12210),.dout(n12403),.clk(gclk));
	jand g12159(.dina(n12403),.dinb(w_n11861_0[0]),.dout(n12404),.clk(gclk));
	jand g12160(.dina(w_n12404_0[1]),.dinb(w_n11653_0[1]),.dout(n12405),.clk(gclk));
	jand g12161(.dina(n12405),.dinb(n12209),.dout(n12406),.clk(gclk));
	jor g12162(.dina(n12406),.dinb(w_asqrt63_31[0]),.dout(n12407),.clk(gclk));
	jand g12163(.dina(w_n12188_0[0]),.dinb(w_n12407_0[1]),.dout(n12408),.clk(gclk));
	jand g12164(.dina(w_n12408_0[1]),.dinb(w_n12207_1[1]),.dout(n12410),.clk(gclk));
	jor g12165(.dina(w_n12410_25[1]),.dinb(n12206),.dout(n12411),.clk(gclk));
	jand g12166(.dina(n12411),.dinb(n12205),.dout(n12412),.clk(gclk));
	jand g12167(.dina(n12412),.dinb(n12203),.dout(n12413),.clk(gclk));
	jor g12168(.dina(n12413),.dinb(w_n12202_0[1]),.dout(n12414),.clk(gclk));
	jand g12169(.dina(w_n12414_0[2]),.dinb(w_asqrt22_21[1]),.dout(n12415),.clk(gclk));
	jor g12170(.dina(w_n12414_0[1]),.dinb(w_asqrt22_21[0]),.dout(n12416),.clk(gclk));
	jand g12171(.dina(w_asqrt20_34[0]),.dinb(w_n11866_0[0]),.dout(n12417),.clk(gclk));
	jand g12172(.dina(w_n12187_0[0]),.dinb(w_n12207_1[0]),.dout(n12418),.clk(gclk));
	jand g12173(.dina(n12418),.dinb(w_n12407_0[0]),.dout(n12419),.clk(gclk));
	jand g12174(.dina(n12419),.dinb(w_asqrt21_14[1]),.dout(n12420),.clk(gclk));
	jor g12175(.dina(n12420),.dinb(w_n12417_0[1]),.dout(n12421),.clk(gclk));
	jxor g12176(.dina(n12421),.dinb(w_a42_0[1]),.dout(n12422),.clk(gclk));
	jnot g12177(.din(w_n12422_0[1]),.dout(n12423),.clk(gclk));
	jand g12178(.dina(w_n12423_0[1]),.dinb(n12416),.dout(n12424),.clk(gclk));
	jor g12179(.dina(n12424),.dinb(w_n12415_0[1]),.dout(n12425),.clk(gclk));
	jand g12180(.dina(w_n12425_0[2]),.dinb(w_asqrt23_15[1]),.dout(n12426),.clk(gclk));
	jor g12181(.dina(w_n12425_0[1]),.dinb(w_asqrt23_15[0]),.dout(n12427),.clk(gclk));
	jxor g12182(.dina(w_n11869_0[0]),.dinb(w_n11347_25[1]),.dout(n12428),.clk(gclk));
	jand g12183(.dina(n12428),.dinb(w_asqrt20_33[2]),.dout(n12429),.clk(gclk));
	jxor g12184(.dina(n12429),.dinb(w_n12256_0[0]),.dout(n12430),.clk(gclk));
	jand g12185(.dina(w_n12430_0[1]),.dinb(n12427),.dout(n12431),.clk(gclk));
	jor g12186(.dina(n12431),.dinb(w_n12426_0[1]),.dout(n12432),.clk(gclk));
	jand g12187(.dina(w_n12432_0[2]),.dinb(w_asqrt24_21[1]),.dout(n12433),.clk(gclk));
	jor g12188(.dina(w_n12432_0[1]),.dinb(w_asqrt24_21[0]),.dout(n12434),.clk(gclk));
	jxor g12189(.dina(w_n11877_0[0]),.dinb(w_n10824_32[0]),.dout(n12435),.clk(gclk));
	jand g12190(.dina(n12435),.dinb(w_asqrt20_33[1]),.dout(n12436),.clk(gclk));
	jxor g12191(.dina(n12436),.dinb(w_n11886_0[0]),.dout(n12437),.clk(gclk));
	jnot g12192(.din(w_n12437_0[1]),.dout(n12438),.clk(gclk));
	jand g12193(.dina(w_n12438_0[1]),.dinb(n12434),.dout(n12439),.clk(gclk));
	jor g12194(.dina(n12439),.dinb(w_n12433_0[1]),.dout(n12440),.clk(gclk));
	jand g12195(.dina(w_n12440_0[2]),.dinb(w_asqrt25_15[1]),.dout(n12441),.clk(gclk));
	jor g12196(.dina(w_n12440_0[1]),.dinb(w_asqrt25_15[0]),.dout(n12442),.clk(gclk));
	jxor g12197(.dina(w_n11888_0[0]),.dinb(w_n10328_26[1]),.dout(n12443),.clk(gclk));
	jand g12198(.dina(n12443),.dinb(w_asqrt20_33[0]),.dout(n12444),.clk(gclk));
	jxor g12199(.dina(n12444),.dinb(w_n11893_0[0]),.dout(n12445),.clk(gclk));
	jand g12200(.dina(w_n12445_0[1]),.dinb(n12442),.dout(n12446),.clk(gclk));
	jor g12201(.dina(n12446),.dinb(w_n12441_0[1]),.dout(n12447),.clk(gclk));
	jand g12202(.dina(w_n12447_0[2]),.dinb(w_asqrt26_21[1]),.dout(n12448),.clk(gclk));
	jor g12203(.dina(w_n12447_0[1]),.dinb(w_asqrt26_21[0]),.dout(n12449),.clk(gclk));
	jxor g12204(.dina(w_n11896_0[0]),.dinb(w_n9832_32[2]),.dout(n12450),.clk(gclk));
	jand g12205(.dina(n12450),.dinb(w_asqrt20_32[2]),.dout(n12451),.clk(gclk));
	jxor g12206(.dina(n12451),.dinb(w_n11901_0[0]),.dout(n12452),.clk(gclk));
	jnot g12207(.din(w_n12452_0[1]),.dout(n12453),.clk(gclk));
	jand g12208(.dina(w_n12453_0[1]),.dinb(n12449),.dout(n12454),.clk(gclk));
	jor g12209(.dina(n12454),.dinb(w_n12448_0[1]),.dout(n12455),.clk(gclk));
	jand g12210(.dina(w_n12455_0[2]),.dinb(w_asqrt27_16[0]),.dout(n12456),.clk(gclk));
	jor g12211(.dina(w_n12455_0[1]),.dinb(w_asqrt27_15[2]),.dout(n12457),.clk(gclk));
	jxor g12212(.dina(w_n11903_0[0]),.dinb(w_n9369_27[1]),.dout(n12458),.clk(gclk));
	jand g12213(.dina(n12458),.dinb(w_asqrt20_32[1]),.dout(n12459),.clk(gclk));
	jxor g12214(.dina(n12459),.dinb(w_n11908_0[0]),.dout(n12460),.clk(gclk));
	jand g12215(.dina(w_n12460_0[1]),.dinb(n12457),.dout(n12461),.clk(gclk));
	jor g12216(.dina(n12461),.dinb(w_n12456_0[1]),.dout(n12462),.clk(gclk));
	jand g12217(.dina(w_n12462_0[2]),.dinb(w_asqrt28_21[2]),.dout(n12463),.clk(gclk));
	jor g12218(.dina(w_n12462_0[1]),.dinb(w_asqrt28_21[1]),.dout(n12464),.clk(gclk));
	jxor g12219(.dina(w_n11911_0[0]),.dinb(w_n8890_33[0]),.dout(n12465),.clk(gclk));
	jand g12220(.dina(n12465),.dinb(w_asqrt20_32[0]),.dout(n12466),.clk(gclk));
	jxor g12221(.dina(n12466),.dinb(w_n11916_0[0]),.dout(n12467),.clk(gclk));
	jnot g12222(.din(w_n12467_0[1]),.dout(n12468),.clk(gclk));
	jand g12223(.dina(w_n12468_0[1]),.dinb(n12464),.dout(n12469),.clk(gclk));
	jor g12224(.dina(n12469),.dinb(w_n12463_0[1]),.dout(n12470),.clk(gclk));
	jand g12225(.dina(w_n12470_0[2]),.dinb(w_asqrt29_16[1]),.dout(n12471),.clk(gclk));
	jor g12226(.dina(w_n12470_0[1]),.dinb(w_asqrt29_16[0]),.dout(n12472),.clk(gclk));
	jxor g12227(.dina(w_n11918_0[0]),.dinb(w_n8449_28[0]),.dout(n12473),.clk(gclk));
	jand g12228(.dina(n12473),.dinb(w_asqrt20_31[2]),.dout(n12474),.clk(gclk));
	jxor g12229(.dina(n12474),.dinb(w_n11923_0[0]),.dout(n12475),.clk(gclk));
	jnot g12230(.din(w_n12475_0[1]),.dout(n12476),.clk(gclk));
	jand g12231(.dina(w_n12476_0[1]),.dinb(n12472),.dout(n12477),.clk(gclk));
	jor g12232(.dina(n12477),.dinb(w_n12471_0[1]),.dout(n12478),.clk(gclk));
	jand g12233(.dina(w_n12478_0[2]),.dinb(w_asqrt30_22[0]),.dout(n12479),.clk(gclk));
	jor g12234(.dina(w_n12478_0[1]),.dinb(w_asqrt30_21[2]),.dout(n12480),.clk(gclk));
	jxor g12235(.dina(w_n11925_0[0]),.dinb(w_n8003_33[2]),.dout(n12481),.clk(gclk));
	jand g12236(.dina(n12481),.dinb(w_asqrt20_31[1]),.dout(n12482),.clk(gclk));
	jxor g12237(.dina(n12482),.dinb(w_n11930_0[0]),.dout(n12483),.clk(gclk));
	jnot g12238(.din(w_n12483_0[1]),.dout(n12484),.clk(gclk));
	jand g12239(.dina(w_n12484_0[1]),.dinb(n12480),.dout(n12485),.clk(gclk));
	jor g12240(.dina(n12485),.dinb(w_n12479_0[1]),.dout(n12486),.clk(gclk));
	jand g12241(.dina(w_n12486_0[2]),.dinb(w_asqrt31_17[0]),.dout(n12487),.clk(gclk));
	jor g12242(.dina(w_n12486_0[1]),.dinb(w_asqrt31_16[2]),.dout(n12488),.clk(gclk));
	jxor g12243(.dina(w_n11932_0[0]),.dinb(w_n7581_29[0]),.dout(n12489),.clk(gclk));
	jand g12244(.dina(n12489),.dinb(w_asqrt20_31[0]),.dout(n12490),.clk(gclk));
	jxor g12245(.dina(n12490),.dinb(w_n11937_0[0]),.dout(n12491),.clk(gclk));
	jand g12246(.dina(w_n12491_0[1]),.dinb(n12488),.dout(n12492),.clk(gclk));
	jor g12247(.dina(n12492),.dinb(w_n12487_0[1]),.dout(n12493),.clk(gclk));
	jand g12248(.dina(w_n12493_0[2]),.dinb(w_asqrt32_22[0]),.dout(n12494),.clk(gclk));
	jor g12249(.dina(w_n12493_0[1]),.dinb(w_asqrt32_21[2]),.dout(n12495),.clk(gclk));
	jxor g12250(.dina(w_n11940_0[0]),.dinb(w_n7154_34[0]),.dout(n12496),.clk(gclk));
	jand g12251(.dina(n12496),.dinb(w_asqrt20_30[2]),.dout(n12497),.clk(gclk));
	jxor g12252(.dina(n12497),.dinb(w_n11945_0[0]),.dout(n12498),.clk(gclk));
	jnot g12253(.din(w_n12498_0[1]),.dout(n12499),.clk(gclk));
	jand g12254(.dina(w_n12499_0[1]),.dinb(n12495),.dout(n12500),.clk(gclk));
	jor g12255(.dina(n12500),.dinb(w_n12494_0[1]),.dout(n12501),.clk(gclk));
	jand g12256(.dina(w_n12501_0[2]),.dinb(w_asqrt33_17[2]),.dout(n12502),.clk(gclk));
	jor g12257(.dina(w_n12501_0[1]),.dinb(w_asqrt33_17[1]),.dout(n12503),.clk(gclk));
	jxor g12258(.dina(w_n11947_0[0]),.dinb(w_n6758_29[2]),.dout(n12504),.clk(gclk));
	jand g12259(.dina(n12504),.dinb(w_asqrt20_30[1]),.dout(n12505),.clk(gclk));
	jxor g12260(.dina(n12505),.dinb(w_n11952_0[0]),.dout(n12506),.clk(gclk));
	jand g12261(.dina(w_n12506_0[1]),.dinb(n12503),.dout(n12507),.clk(gclk));
	jor g12262(.dina(n12507),.dinb(w_n12502_0[1]),.dout(n12508),.clk(gclk));
	jand g12263(.dina(w_n12508_0[2]),.dinb(w_asqrt34_22[1]),.dout(n12509),.clk(gclk));
	jor g12264(.dina(w_n12508_0[1]),.dinb(w_asqrt34_22[0]),.dout(n12510),.clk(gclk));
	jxor g12265(.dina(w_n11955_0[0]),.dinb(w_n6357_34[1]),.dout(n12511),.clk(gclk));
	jand g12266(.dina(n12511),.dinb(w_asqrt20_30[0]),.dout(n12512),.clk(gclk));
	jxor g12267(.dina(n12512),.dinb(w_n11960_0[0]),.dout(n12513),.clk(gclk));
	jnot g12268(.din(w_n12513_0[1]),.dout(n12514),.clk(gclk));
	jand g12269(.dina(w_n12514_0[1]),.dinb(n12510),.dout(n12515),.clk(gclk));
	jor g12270(.dina(n12515),.dinb(w_n12509_0[1]),.dout(n12516),.clk(gclk));
	jand g12271(.dina(w_n12516_0[2]),.dinb(w_asqrt35_18[1]),.dout(n12517),.clk(gclk));
	jor g12272(.dina(w_n12516_0[1]),.dinb(w_asqrt35_18[0]),.dout(n12518),.clk(gclk));
	jxor g12273(.dina(w_n11962_0[0]),.dinb(w_n5989_30[1]),.dout(n12519),.clk(gclk));
	jand g12274(.dina(n12519),.dinb(w_asqrt20_29[2]),.dout(n12520),.clk(gclk));
	jxor g12275(.dina(n12520),.dinb(w_n11967_0[0]),.dout(n12521),.clk(gclk));
	jnot g12276(.din(w_n12521_0[1]),.dout(n12522),.clk(gclk));
	jand g12277(.dina(w_n12522_0[1]),.dinb(n12518),.dout(n12523),.clk(gclk));
	jor g12278(.dina(n12523),.dinb(w_n12517_0[1]),.dout(n12524),.clk(gclk));
	jand g12279(.dina(w_n12524_0[2]),.dinb(w_asqrt36_22[1]),.dout(n12525),.clk(gclk));
	jor g12280(.dina(w_n12524_0[1]),.dinb(w_asqrt36_22[0]),.dout(n12526),.clk(gclk));
	jxor g12281(.dina(w_n11969_0[0]),.dinb(w_n5606_34[2]),.dout(n12527),.clk(gclk));
	jand g12282(.dina(n12527),.dinb(w_asqrt20_29[1]),.dout(n12528),.clk(gclk));
	jxor g12283(.dina(n12528),.dinb(w_n11974_0[0]),.dout(n12529),.clk(gclk));
	jnot g12284(.din(w_n12529_0[1]),.dout(n12530),.clk(gclk));
	jand g12285(.dina(w_n12530_0[1]),.dinb(n12526),.dout(n12531),.clk(gclk));
	jor g12286(.dina(n12531),.dinb(w_n12525_0[1]),.dout(n12532),.clk(gclk));
	jand g12287(.dina(w_n12532_0[2]),.dinb(w_asqrt37_18[2]),.dout(n12533),.clk(gclk));
	jor g12288(.dina(w_n12532_0[1]),.dinb(w_asqrt37_18[1]),.dout(n12534),.clk(gclk));
	jxor g12289(.dina(w_n11976_0[0]),.dinb(w_n5259_31[1]),.dout(n12535),.clk(gclk));
	jand g12290(.dina(n12535),.dinb(w_asqrt20_29[0]),.dout(n12536),.clk(gclk));
	jxor g12291(.dina(n12536),.dinb(w_n11981_0[0]),.dout(n12537),.clk(gclk));
	jand g12292(.dina(w_n12537_0[1]),.dinb(n12534),.dout(n12538),.clk(gclk));
	jor g12293(.dina(n12538),.dinb(w_n12533_0[1]),.dout(n12539),.clk(gclk));
	jand g12294(.dina(w_n12539_0[2]),.dinb(w_asqrt38_22[2]),.dout(n12540),.clk(gclk));
	jor g12295(.dina(w_n12539_0[1]),.dinb(w_asqrt38_22[1]),.dout(n12541),.clk(gclk));
	jxor g12296(.dina(w_n11984_0[0]),.dinb(w_n4902_35[1]),.dout(n12542),.clk(gclk));
	jand g12297(.dina(n12542),.dinb(w_asqrt20_28[2]),.dout(n12543),.clk(gclk));
	jxor g12298(.dina(n12543),.dinb(w_n11989_0[0]),.dout(n12544),.clk(gclk));
	jnot g12299(.din(w_n12544_0[1]),.dout(n12545),.clk(gclk));
	jand g12300(.dina(w_n12545_0[1]),.dinb(n12541),.dout(n12546),.clk(gclk));
	jor g12301(.dina(n12546),.dinb(w_n12540_0[1]),.dout(n12547),.clk(gclk));
	jand g12302(.dina(w_n12547_0[2]),.dinb(w_asqrt39_19[1]),.dout(n12548),.clk(gclk));
	jor g12303(.dina(w_n12547_0[1]),.dinb(w_asqrt39_19[0]),.dout(n12549),.clk(gclk));
	jxor g12304(.dina(w_n11991_0[0]),.dinb(w_n4582_32[1]),.dout(n12550),.clk(gclk));
	jand g12305(.dina(n12550),.dinb(w_asqrt20_28[1]),.dout(n12551),.clk(gclk));
	jxor g12306(.dina(n12551),.dinb(w_n11996_0[0]),.dout(n12552),.clk(gclk));
	jnot g12307(.din(w_n12552_0[1]),.dout(n12553),.clk(gclk));
	jand g12308(.dina(w_n12553_0[1]),.dinb(n12549),.dout(n12554),.clk(gclk));
	jor g12309(.dina(n12554),.dinb(w_n12548_0[1]),.dout(n12555),.clk(gclk));
	jand g12310(.dina(w_n12555_0[2]),.dinb(w_asqrt40_22[2]),.dout(n12556),.clk(gclk));
	jor g12311(.dina(w_n12555_0[1]),.dinb(w_asqrt40_22[1]),.dout(n12557),.clk(gclk));
	jxor g12312(.dina(w_n11998_0[0]),.dinb(w_n4249_36[0]),.dout(n12558),.clk(gclk));
	jand g12313(.dina(n12558),.dinb(w_asqrt20_28[0]),.dout(n12559),.clk(gclk));
	jxor g12314(.dina(n12559),.dinb(w_n12003_0[0]),.dout(n12560),.clk(gclk));
	jnot g12315(.din(w_n12560_0[1]),.dout(n12561),.clk(gclk));
	jand g12316(.dina(w_n12561_0[1]),.dinb(n12557),.dout(n12562),.clk(gclk));
	jor g12317(.dina(n12562),.dinb(w_n12556_0[1]),.dout(n12563),.clk(gclk));
	jand g12318(.dina(w_n12563_0[2]),.dinb(w_asqrt41_19[2]),.dout(n12564),.clk(gclk));
	jor g12319(.dina(w_n12563_0[1]),.dinb(w_asqrt41_19[1]),.dout(n12565),.clk(gclk));
	jxor g12320(.dina(w_n12005_0[0]),.dinb(w_n3955_33[0]),.dout(n12566),.clk(gclk));
	jand g12321(.dina(n12566),.dinb(w_asqrt20_27[2]),.dout(n12567),.clk(gclk));
	jxor g12322(.dina(n12567),.dinb(w_n12010_0[0]),.dout(n12568),.clk(gclk));
	jnot g12323(.din(w_n12568_0[1]),.dout(n12569),.clk(gclk));
	jand g12324(.dina(w_n12569_0[1]),.dinb(n12565),.dout(n12570),.clk(gclk));
	jor g12325(.dina(n12570),.dinb(w_n12564_0[1]),.dout(n12571),.clk(gclk));
	jand g12326(.dina(w_n12571_0[2]),.dinb(w_asqrt42_23[0]),.dout(n12572),.clk(gclk));
	jor g12327(.dina(w_n12571_0[1]),.dinb(w_asqrt42_22[2]),.dout(n12573),.clk(gclk));
	jxor g12328(.dina(w_n12012_0[0]),.dinb(w_n3642_36[1]),.dout(n12574),.clk(gclk));
	jand g12329(.dina(n12574),.dinb(w_asqrt20_27[1]),.dout(n12575),.clk(gclk));
	jxor g12330(.dina(n12575),.dinb(w_n12017_0[0]),.dout(n12576),.clk(gclk));
	jnot g12331(.din(w_n12576_0[2]),.dout(n12577),.clk(gclk));
	jand g12332(.dina(n12577),.dinb(n12573),.dout(n12578),.clk(gclk));
	jor g12333(.dina(n12578),.dinb(w_n12572_0[1]),.dout(n12579),.clk(gclk));
	jand g12334(.dina(w_n12579_0[2]),.dinb(w_asqrt43_20[0]),.dout(n12580),.clk(gclk));
	jxor g12335(.dina(w_n12019_0[0]),.dinb(w_n3368_33[2]),.dout(n12581),.clk(gclk));
	jand g12336(.dina(n12581),.dinb(w_asqrt20_27[0]),.dout(n12582),.clk(gclk));
	jxor g12337(.dina(n12582),.dinb(w_n12023_0[0]),.dout(n12583),.clk(gclk));
	jor g12338(.dina(w_n12579_0[1]),.dinb(w_asqrt43_19[2]),.dout(n12584),.clk(gclk));
	jand g12339(.dina(n12584),.dinb(w_n12583_0[1]),.dout(n12585),.clk(gclk));
	jor g12340(.dina(n12585),.dinb(w_n12580_0[1]),.dout(n12586),.clk(gclk));
	jand g12341(.dina(w_n12586_0[2]),.dinb(w_asqrt44_23[0]),.dout(n12587),.clk(gclk));
	jor g12342(.dina(w_n12586_0[1]),.dinb(w_asqrt44_22[2]),.dout(n12588),.clk(gclk));
	jxor g12343(.dina(w_n12027_0[0]),.dinb(w_n3089_37[0]),.dout(n12589),.clk(gclk));
	jand g12344(.dina(n12589),.dinb(w_asqrt20_26[2]),.dout(n12590),.clk(gclk));
	jxor g12345(.dina(n12590),.dinb(w_n12032_0[0]),.dout(n12591),.clk(gclk));
	jnot g12346(.din(w_n12591_0[1]),.dout(n12592),.clk(gclk));
	jand g12347(.dina(w_n12592_0[1]),.dinb(n12588),.dout(n12593),.clk(gclk));
	jor g12348(.dina(n12593),.dinb(w_n12587_0[1]),.dout(n12594),.clk(gclk));
	jand g12349(.dina(w_n12594_0[2]),.dinb(w_asqrt45_20[2]),.dout(n12595),.clk(gclk));
	jor g12350(.dina(w_n12594_0[1]),.dinb(w_asqrt45_20[1]),.dout(n12596),.clk(gclk));
	jxor g12351(.dina(w_n12034_0[0]),.dinb(w_n2833_34[2]),.dout(n12597),.clk(gclk));
	jand g12352(.dina(n12597),.dinb(w_asqrt20_26[1]),.dout(n12598),.clk(gclk));
	jxor g12353(.dina(n12598),.dinb(w_n12039_0[0]),.dout(n12599),.clk(gclk));
	jand g12354(.dina(w_n12599_0[1]),.dinb(n12596),.dout(n12600),.clk(gclk));
	jor g12355(.dina(n12600),.dinb(w_n12595_0[1]),.dout(n12601),.clk(gclk));
	jand g12356(.dina(w_n12601_0[2]),.dinb(w_asqrt46_23[0]),.dout(n12602),.clk(gclk));
	jor g12357(.dina(w_n12601_0[1]),.dinb(w_asqrt46_22[2]),.dout(n12603),.clk(gclk));
	jxor g12358(.dina(w_n12042_0[0]),.dinb(w_n2572_37[1]),.dout(n12604),.clk(gclk));
	jand g12359(.dina(n12604),.dinb(w_asqrt20_26[0]),.dout(n12605),.clk(gclk));
	jxor g12360(.dina(n12605),.dinb(w_n12047_0[0]),.dout(n12606),.clk(gclk));
	jnot g12361(.din(w_n12606_0[1]),.dout(n12607),.clk(gclk));
	jand g12362(.dina(w_n12607_0[1]),.dinb(n12603),.dout(n12608),.clk(gclk));
	jor g12363(.dina(n12608),.dinb(w_n12602_0[1]),.dout(n12609),.clk(gclk));
	jand g12364(.dina(w_n12609_0[2]),.dinb(w_asqrt47_21[1]),.dout(n12610),.clk(gclk));
	jor g12365(.dina(w_n12609_0[1]),.dinb(w_asqrt47_21[0]),.dout(n12611),.clk(gclk));
	jxor g12366(.dina(w_n12049_0[0]),.dinb(w_n2345_35[1]),.dout(n12612),.clk(gclk));
	jand g12367(.dina(n12612),.dinb(w_asqrt20_25[2]),.dout(n12613),.clk(gclk));
	jxor g12368(.dina(n12613),.dinb(w_n12054_0[0]),.dout(n12614),.clk(gclk));
	jand g12369(.dina(w_n12614_0[1]),.dinb(n12611),.dout(n12615),.clk(gclk));
	jor g12370(.dina(n12615),.dinb(w_n12610_0[1]),.dout(n12616),.clk(gclk));
	jand g12371(.dina(w_n12616_0[2]),.dinb(w_asqrt48_23[1]),.dout(n12617),.clk(gclk));
	jor g12372(.dina(w_n12616_0[1]),.dinb(w_asqrt48_23[0]),.dout(n12618),.clk(gclk));
	jxor g12373(.dina(w_n12057_0[0]),.dinb(w_n2108_38[0]),.dout(n12619),.clk(gclk));
	jand g12374(.dina(n12619),.dinb(w_asqrt20_25[1]),.dout(n12620),.clk(gclk));
	jxor g12375(.dina(n12620),.dinb(w_n12062_0[0]),.dout(n12621),.clk(gclk));
	jnot g12376(.din(w_n12621_0[1]),.dout(n12622),.clk(gclk));
	jand g12377(.dina(w_n12622_0[1]),.dinb(n12618),.dout(n12623),.clk(gclk));
	jor g12378(.dina(n12623),.dinb(w_n12617_0[1]),.dout(n12624),.clk(gclk));
	jand g12379(.dina(w_n12624_0[2]),.dinb(w_asqrt49_21[2]),.dout(n12625),.clk(gclk));
	jor g12380(.dina(w_n12624_0[1]),.dinb(w_asqrt49_21[1]),.dout(n12626),.clk(gclk));
	jxor g12381(.dina(w_n12064_0[0]),.dinb(w_n1912_36[1]),.dout(n12627),.clk(gclk));
	jand g12382(.dina(n12627),.dinb(w_asqrt20_25[0]),.dout(n12628),.clk(gclk));
	jxor g12383(.dina(n12628),.dinb(w_n12069_0[0]),.dout(n12629),.clk(gclk));
	jnot g12384(.din(w_n12629_0[1]),.dout(n12630),.clk(gclk));
	jand g12385(.dina(w_n12630_0[1]),.dinb(n12626),.dout(n12631),.clk(gclk));
	jor g12386(.dina(n12631),.dinb(w_n12625_0[1]),.dout(n12632),.clk(gclk));
	jand g12387(.dina(w_n12632_0[2]),.dinb(w_asqrt50_23[2]),.dout(n12633),.clk(gclk));
	jor g12388(.dina(w_n12632_0[1]),.dinb(w_asqrt50_23[1]),.dout(n12634),.clk(gclk));
	jxor g12389(.dina(w_n12071_0[0]),.dinb(w_n1699_38[2]),.dout(n12635),.clk(gclk));
	jand g12390(.dina(n12635),.dinb(w_asqrt20_24[2]),.dout(n12636),.clk(gclk));
	jxor g12391(.dina(n12636),.dinb(w_n12076_0[0]),.dout(n12637),.clk(gclk));
	jnot g12392(.din(w_n12637_0[1]),.dout(n12638),.clk(gclk));
	jand g12393(.dina(w_n12638_0[1]),.dinb(n12634),.dout(n12639),.clk(gclk));
	jor g12394(.dina(n12639),.dinb(w_n12633_0[1]),.dout(n12640),.clk(gclk));
	jand g12395(.dina(w_n12640_0[2]),.dinb(w_asqrt51_22[0]),.dout(n12641),.clk(gclk));
	jor g12396(.dina(w_n12640_0[1]),.dinb(w_asqrt51_21[2]),.dout(n12642),.clk(gclk));
	jxor g12397(.dina(w_n12078_0[0]),.dinb(w_n1516_37[0]),.dout(n12643),.clk(gclk));
	jand g12398(.dina(n12643),.dinb(w_asqrt20_24[1]),.dout(n12644),.clk(gclk));
	jxor g12399(.dina(n12644),.dinb(w_n12083_0[0]),.dout(n12645),.clk(gclk));
	jand g12400(.dina(w_n12645_0[1]),.dinb(n12642),.dout(n12646),.clk(gclk));
	jor g12401(.dina(n12646),.dinb(w_n12641_0[1]),.dout(n12647),.clk(gclk));
	jand g12402(.dina(w_n12647_0[2]),.dinb(w_asqrt52_23[2]),.dout(n12648),.clk(gclk));
	jor g12403(.dina(w_n12647_0[1]),.dinb(w_asqrt52_23[1]),.dout(n12649),.clk(gclk));
	jxor g12404(.dina(w_n12086_0[0]),.dinb(w_n1332_38[2]),.dout(n12650),.clk(gclk));
	jand g12405(.dina(n12650),.dinb(w_asqrt20_24[0]),.dout(n12651),.clk(gclk));
	jxor g12406(.dina(n12651),.dinb(w_n12091_0[0]),.dout(n12652),.clk(gclk));
	jnot g12407(.din(w_n12652_0[1]),.dout(n12653),.clk(gclk));
	jand g12408(.dina(w_n12653_0[1]),.dinb(n12649),.dout(n12654),.clk(gclk));
	jor g12409(.dina(n12654),.dinb(w_n12648_0[1]),.dout(n12655),.clk(gclk));
	jand g12410(.dina(w_n12655_0[2]),.dinb(w_asqrt53_22[2]),.dout(n12656),.clk(gclk));
	jor g12411(.dina(w_n12655_0[1]),.dinb(w_asqrt53_22[1]),.dout(n12657),.clk(gclk));
	jxor g12412(.dina(w_n12093_0[0]),.dinb(w_n1173_37[2]),.dout(n12658),.clk(gclk));
	jand g12413(.dina(n12658),.dinb(w_asqrt20_23[2]),.dout(n12659),.clk(gclk));
	jxor g12414(.dina(n12659),.dinb(w_n12098_0[0]),.dout(n12660),.clk(gclk));
	jand g12415(.dina(w_n12660_0[1]),.dinb(n12657),.dout(n12661),.clk(gclk));
	jor g12416(.dina(n12661),.dinb(w_n12656_0[1]),.dout(n12662),.clk(gclk));
	jand g12417(.dina(w_n12662_0[2]),.dinb(w_asqrt54_23[2]),.dout(n12663),.clk(gclk));
	jor g12418(.dina(w_n12662_0[1]),.dinb(w_asqrt54_23[1]),.dout(n12664),.clk(gclk));
	jxor g12419(.dina(w_n12101_0[0]),.dinb(w_n1008_39[2]),.dout(n12665),.clk(gclk));
	jand g12420(.dina(n12665),.dinb(w_asqrt20_23[1]),.dout(n12666),.clk(gclk));
	jxor g12421(.dina(n12666),.dinb(w_n12106_0[0]),.dout(n12667),.clk(gclk));
	jnot g12422(.din(w_n12667_0[1]),.dout(n12668),.clk(gclk));
	jand g12423(.dina(w_n12668_0[1]),.dinb(n12664),.dout(n12669),.clk(gclk));
	jor g12424(.dina(n12669),.dinb(w_n12663_0[1]),.dout(n12670),.clk(gclk));
	jand g12425(.dina(w_n12670_0[2]),.dinb(w_asqrt55_23[0]),.dout(n12671),.clk(gclk));
	jor g12426(.dina(w_n12670_0[1]),.dinb(w_asqrt55_22[2]),.dout(n12672),.clk(gclk));
	jxor g12427(.dina(w_n12108_0[0]),.dinb(w_n884_38[2]),.dout(n12673),.clk(gclk));
	jand g12428(.dina(n12673),.dinb(w_asqrt20_23[0]),.dout(n12674),.clk(gclk));
	jxor g12429(.dina(n12674),.dinb(w_n12113_0[0]),.dout(n12675),.clk(gclk));
	jand g12430(.dina(w_n12675_0[1]),.dinb(n12672),.dout(n12676),.clk(gclk));
	jor g12431(.dina(n12676),.dinb(w_n12671_0[1]),.dout(n12677),.clk(gclk));
	jand g12432(.dina(w_n12677_0[2]),.dinb(w_asqrt56_24[0]),.dout(n12678),.clk(gclk));
	jor g12433(.dina(w_n12677_0[1]),.dinb(w_asqrt56_23[2]),.dout(n12679),.clk(gclk));
	jxor g12434(.dina(w_n12116_0[0]),.dinb(w_n743_39[2]),.dout(n12680),.clk(gclk));
	jand g12435(.dina(n12680),.dinb(w_asqrt20_22[2]),.dout(n12681),.clk(gclk));
	jxor g12436(.dina(n12681),.dinb(w_n12121_0[0]),.dout(n12682),.clk(gclk));
	jnot g12437(.din(w_n12682_0[1]),.dout(n12683),.clk(gclk));
	jand g12438(.dina(w_n12683_0[1]),.dinb(n12679),.dout(n12684),.clk(gclk));
	jor g12439(.dina(n12684),.dinb(w_n12678_0[1]),.dout(n12685),.clk(gclk));
	jand g12440(.dina(w_n12685_0[2]),.dinb(w_asqrt57_23[2]),.dout(n12686),.clk(gclk));
	jor g12441(.dina(w_n12685_0[1]),.dinb(w_asqrt57_23[1]),.dout(n12687),.clk(gclk));
	jxor g12442(.dina(w_n12123_0[0]),.dinb(w_n635_39[2]),.dout(n12688),.clk(gclk));
	jand g12443(.dina(n12688),.dinb(w_asqrt20_22[1]),.dout(n12689),.clk(gclk));
	jxor g12444(.dina(n12689),.dinb(w_n12128_0[0]),.dout(n12690),.clk(gclk));
	jand g12445(.dina(w_n12690_0[1]),.dinb(n12687),.dout(n12691),.clk(gclk));
	jor g12446(.dina(n12691),.dinb(w_n12686_0[1]),.dout(n12692),.clk(gclk));
	jand g12447(.dina(w_n12692_0[2]),.dinb(w_asqrt58_24[1]),.dout(n12693),.clk(gclk));
	jor g12448(.dina(w_n12692_0[1]),.dinb(w_asqrt58_24[0]),.dout(n12694),.clk(gclk));
	jxor g12449(.dina(w_n12131_0[0]),.dinb(w_n515_40[2]),.dout(n12695),.clk(gclk));
	jand g12450(.dina(n12695),.dinb(w_asqrt20_22[0]),.dout(n12696),.clk(gclk));
	jxor g12451(.dina(n12696),.dinb(w_n12136_0[0]),.dout(n12697),.clk(gclk));
	jand g12452(.dina(w_n12697_0[1]),.dinb(n12694),.dout(n12698),.clk(gclk));
	jor g12453(.dina(n12698),.dinb(w_n12693_0[1]),.dout(n12699),.clk(gclk));
	jand g12454(.dina(w_n12699_0[2]),.dinb(w_asqrt59_24[0]),.dout(n12700),.clk(gclk));
	jor g12455(.dina(w_n12699_0[1]),.dinb(w_asqrt59_23[2]),.dout(n12701),.clk(gclk));
	jxor g12456(.dina(w_n12139_0[0]),.dinb(w_n443_40[2]),.dout(n12702),.clk(gclk));
	jand g12457(.dina(n12702),.dinb(w_asqrt20_21[2]),.dout(n12703),.clk(gclk));
	jxor g12458(.dina(n12703),.dinb(w_n12144_0[0]),.dout(n12704),.clk(gclk));
	jand g12459(.dina(w_n12704_0[1]),.dinb(n12701),.dout(n12705),.clk(gclk));
	jor g12460(.dina(n12705),.dinb(w_n12700_0[1]),.dout(n12706),.clk(gclk));
	jand g12461(.dina(w_n12706_0[2]),.dinb(w_asqrt60_24[1]),.dout(n12707),.clk(gclk));
	jor g12462(.dina(w_n12706_0[1]),.dinb(w_asqrt60_24[0]),.dout(n12708),.clk(gclk));
	jxor g12463(.dina(w_n12147_0[0]),.dinb(w_n352_41[0]),.dout(n12709),.clk(gclk));
	jand g12464(.dina(n12709),.dinb(w_asqrt20_21[1]),.dout(n12710),.clk(gclk));
	jxor g12465(.dina(n12710),.dinb(w_n12152_0[0]),.dout(n12711),.clk(gclk));
	jnot g12466(.din(w_n12711_0[1]),.dout(n12712),.clk(gclk));
	jand g12467(.dina(w_n12712_0[1]),.dinb(n12708),.dout(n12713),.clk(gclk));
	jor g12468(.dina(n12713),.dinb(w_n12707_0[1]),.dout(n12714),.clk(gclk));
	jand g12469(.dina(w_n12714_0[2]),.dinb(w_asqrt61_24[1]),.dout(n12715),.clk(gclk));
	jor g12470(.dina(w_n12714_0[1]),.dinb(w_asqrt61_24[0]),.dout(n12716),.clk(gclk));
	jxor g12471(.dina(w_n12154_0[0]),.dinb(w_n294_41[1]),.dout(n12717),.clk(gclk));
	jand g12472(.dina(n12717),.dinb(w_asqrt20_21[0]),.dout(n12718),.clk(gclk));
	jxor g12473(.dina(n12718),.dinb(w_n12159_0[0]),.dout(n12719),.clk(gclk));
	jnot g12474(.din(w_n12719_0[1]),.dout(n12720),.clk(gclk));
	jand g12475(.dina(w_n12720_0[1]),.dinb(n12716),.dout(n12721),.clk(gclk));
	jor g12476(.dina(n12721),.dinb(w_n12715_0[1]),.dout(n12722),.clk(gclk));
	jand g12477(.dina(w_n12722_0[2]),.dinb(w_asqrt62_24[1]),.dout(n12723),.clk(gclk));
	jor g12478(.dina(w_n12722_0[1]),.dinb(w_asqrt62_24[0]),.dout(n12724),.clk(gclk));
	jxor g12479(.dina(w_n12161_0[0]),.dinb(w_n239_41[1]),.dout(n12725),.clk(gclk));
	jand g12480(.dina(n12725),.dinb(w_asqrt20_20[2]),.dout(n12726),.clk(gclk));
	jxor g12481(.dina(n12726),.dinb(w_n12166_0[0]),.dout(n12727),.clk(gclk));
	jnot g12482(.din(w_n12727_0[2]),.dout(n12728),.clk(gclk));
	jand g12483(.dina(n12728),.dinb(n12724),.dout(n12729),.clk(gclk));
	jor g12484(.dina(n12729),.dinb(w_n12723_0[1]),.dout(n12730),.clk(gclk));
	jor g12485(.dina(w_n12730_0[1]),.dinb(w_n12195_0[2]),.dout(n12731),.clk(gclk));
	jnot g12486(.din(w_n12731_1[1]),.dout(n12732),.clk(gclk));
	jand g12487(.dina(w_n12408_0[0]),.dinb(w_n12176_0[0]),.dout(n12733),.clk(gclk));
	jnot g12488(.din(n12733),.dout(n12734),.clk(gclk));
	jand g12489(.dina(w_n12180_0[0]),.dinb(w_asqrt63_30[2]),.dout(n12735),.clk(gclk));
	jand g12490(.dina(n12735),.dinb(w_n12207_0[2]),.dout(n12736),.clk(gclk));
	jand g12491(.dina(w_n12736_0[1]),.dinb(n12734),.dout(n12737),.clk(gclk));
	jand g12492(.dina(w_n12190_0[0]),.dinb(w_n12404_0[0]),.dout(n12738),.clk(gclk));
	jnot g12493(.din(w_n12195_0[1]),.dout(n12739),.clk(gclk));
	jnot g12494(.din(w_n12723_0[0]),.dout(n12740),.clk(gclk));
	jnot g12495(.din(w_n12715_0[0]),.dout(n12741),.clk(gclk));
	jnot g12496(.din(w_n12707_0[0]),.dout(n12742),.clk(gclk));
	jnot g12497(.din(w_n12700_0[0]),.dout(n12743),.clk(gclk));
	jnot g12498(.din(w_n12693_0[0]),.dout(n12744),.clk(gclk));
	jnot g12499(.din(w_n12686_0[0]),.dout(n12745),.clk(gclk));
	jnot g12500(.din(w_n12678_0[0]),.dout(n12746),.clk(gclk));
	jnot g12501(.din(w_n12671_0[0]),.dout(n12747),.clk(gclk));
	jnot g12502(.din(w_n12663_0[0]),.dout(n12748),.clk(gclk));
	jnot g12503(.din(w_n12656_0[0]),.dout(n12749),.clk(gclk));
	jnot g12504(.din(w_n12648_0[0]),.dout(n12750),.clk(gclk));
	jnot g12505(.din(w_n12641_0[0]),.dout(n12751),.clk(gclk));
	jnot g12506(.din(w_n12633_0[0]),.dout(n12752),.clk(gclk));
	jnot g12507(.din(w_n12625_0[0]),.dout(n12753),.clk(gclk));
	jnot g12508(.din(w_n12617_0[0]),.dout(n12754),.clk(gclk));
	jnot g12509(.din(w_n12610_0[0]),.dout(n12755),.clk(gclk));
	jnot g12510(.din(w_n12602_0[0]),.dout(n12756),.clk(gclk));
	jnot g12511(.din(w_n12595_0[0]),.dout(n12757),.clk(gclk));
	jnot g12512(.din(w_n12587_0[0]),.dout(n12758),.clk(gclk));
	jnot g12513(.din(w_n12580_0[0]),.dout(n12759),.clk(gclk));
	jnot g12514(.din(w_n12583_0[0]),.dout(n12760),.clk(gclk));
	jnot g12515(.din(w_n12572_0[0]),.dout(n12761),.clk(gclk));
	jnot g12516(.din(w_n12564_0[0]),.dout(n12762),.clk(gclk));
	jnot g12517(.din(w_n12556_0[0]),.dout(n12763),.clk(gclk));
	jnot g12518(.din(w_n12548_0[0]),.dout(n12764),.clk(gclk));
	jnot g12519(.din(w_n12540_0[0]),.dout(n12765),.clk(gclk));
	jnot g12520(.din(w_n12533_0[0]),.dout(n12766),.clk(gclk));
	jnot g12521(.din(w_n12525_0[0]),.dout(n12767),.clk(gclk));
	jnot g12522(.din(w_n12517_0[0]),.dout(n12768),.clk(gclk));
	jnot g12523(.din(w_n12509_0[0]),.dout(n12769),.clk(gclk));
	jnot g12524(.din(w_n12502_0[0]),.dout(n12770),.clk(gclk));
	jnot g12525(.din(w_n12494_0[0]),.dout(n12771),.clk(gclk));
	jnot g12526(.din(w_n12487_0[0]),.dout(n12772),.clk(gclk));
	jnot g12527(.din(w_n12479_0[0]),.dout(n12773),.clk(gclk));
	jnot g12528(.din(w_n12471_0[0]),.dout(n12774),.clk(gclk));
	jnot g12529(.din(w_n12463_0[0]),.dout(n12775),.clk(gclk));
	jnot g12530(.din(w_n12456_0[0]),.dout(n12776),.clk(gclk));
	jnot g12531(.din(w_n12448_0[0]),.dout(n12777),.clk(gclk));
	jnot g12532(.din(w_n12441_0[0]),.dout(n12778),.clk(gclk));
	jnot g12533(.din(w_n12433_0[0]),.dout(n12779),.clk(gclk));
	jnot g12534(.din(w_n12426_0[0]),.dout(n12780),.clk(gclk));
	jnot g12535(.din(w_n12415_0[0]),.dout(n12781),.clk(gclk));
	jnot g12536(.din(w_n12202_0[0]),.dout(n12782),.clk(gclk));
	jnot g12537(.din(w_n12199_0[0]),.dout(n12783),.clk(gclk));
	jor g12538(.dina(w_n12410_25[0]),.dinb(w_n11864_0[2]),.dout(n12784),.clk(gclk));
	jand g12539(.dina(n12784),.dinb(n12783),.dout(n12785),.clk(gclk));
	jand g12540(.dina(n12785),.dinb(w_n11858_31[0]),.dout(n12786),.clk(gclk));
	jor g12541(.dina(w_n12410_24[2]),.dinb(w_a40_0[0]),.dout(n12787),.clk(gclk));
	jand g12542(.dina(n12787),.dinb(w_a41_0[0]),.dout(n12788),.clk(gclk));
	jor g12543(.dina(w_n12417_0[0]),.dinb(n12788),.dout(n12789),.clk(gclk));
	jor g12544(.dina(w_n12789_0[1]),.dinb(n12786),.dout(n12790),.clk(gclk));
	jand g12545(.dina(n12790),.dinb(n12782),.dout(n12791),.clk(gclk));
	jand g12546(.dina(n12791),.dinb(w_n11347_25[0]),.dout(n12792),.clk(gclk));
	jor g12547(.dina(w_n12422_0[0]),.dinb(n12792),.dout(n12793),.clk(gclk));
	jand g12548(.dina(n12793),.dinb(n12781),.dout(n12794),.clk(gclk));
	jand g12549(.dina(n12794),.dinb(w_n10824_31[2]),.dout(n12795),.clk(gclk));
	jnot g12550(.din(w_n12430_0[0]),.dout(n12796),.clk(gclk));
	jor g12551(.dina(w_n12796_0[1]),.dinb(n12795),.dout(n12797),.clk(gclk));
	jand g12552(.dina(n12797),.dinb(n12780),.dout(n12798),.clk(gclk));
	jand g12553(.dina(n12798),.dinb(w_n10328_26[0]),.dout(n12799),.clk(gclk));
	jor g12554(.dina(w_n12437_0[0]),.dinb(n12799),.dout(n12800),.clk(gclk));
	jand g12555(.dina(n12800),.dinb(n12779),.dout(n12801),.clk(gclk));
	jand g12556(.dina(n12801),.dinb(w_n9832_32[1]),.dout(n12802),.clk(gclk));
	jnot g12557(.din(w_n12445_0[0]),.dout(n12803),.clk(gclk));
	jor g12558(.dina(w_n12803_0[1]),.dinb(n12802),.dout(n12804),.clk(gclk));
	jand g12559(.dina(n12804),.dinb(n12778),.dout(n12805),.clk(gclk));
	jand g12560(.dina(n12805),.dinb(w_n9369_27[0]),.dout(n12806),.clk(gclk));
	jor g12561(.dina(w_n12452_0[0]),.dinb(n12806),.dout(n12807),.clk(gclk));
	jand g12562(.dina(n12807),.dinb(n12777),.dout(n12808),.clk(gclk));
	jand g12563(.dina(n12808),.dinb(w_n8890_32[2]),.dout(n12809),.clk(gclk));
	jnot g12564(.din(w_n12460_0[0]),.dout(n12810),.clk(gclk));
	jor g12565(.dina(w_n12810_0[1]),.dinb(n12809),.dout(n12811),.clk(gclk));
	jand g12566(.dina(n12811),.dinb(n12776),.dout(n12812),.clk(gclk));
	jand g12567(.dina(n12812),.dinb(w_n8449_27[2]),.dout(n12813),.clk(gclk));
	jor g12568(.dina(w_n12467_0[0]),.dinb(n12813),.dout(n12814),.clk(gclk));
	jand g12569(.dina(n12814),.dinb(n12775),.dout(n12815),.clk(gclk));
	jand g12570(.dina(n12815),.dinb(w_n8003_33[1]),.dout(n12816),.clk(gclk));
	jor g12571(.dina(w_n12475_0[0]),.dinb(n12816),.dout(n12817),.clk(gclk));
	jand g12572(.dina(n12817),.dinb(n12774),.dout(n12818),.clk(gclk));
	jand g12573(.dina(n12818),.dinb(w_n7581_28[2]),.dout(n12819),.clk(gclk));
	jor g12574(.dina(w_n12483_0[0]),.dinb(n12819),.dout(n12820),.clk(gclk));
	jand g12575(.dina(n12820),.dinb(n12773),.dout(n12821),.clk(gclk));
	jand g12576(.dina(n12821),.dinb(w_n7154_33[2]),.dout(n12822),.clk(gclk));
	jnot g12577(.din(w_n12491_0[0]),.dout(n12823),.clk(gclk));
	jor g12578(.dina(w_n12823_0[1]),.dinb(n12822),.dout(n12824),.clk(gclk));
	jand g12579(.dina(n12824),.dinb(n12772),.dout(n12825),.clk(gclk));
	jand g12580(.dina(n12825),.dinb(w_n6758_29[1]),.dout(n12826),.clk(gclk));
	jor g12581(.dina(w_n12498_0[0]),.dinb(n12826),.dout(n12827),.clk(gclk));
	jand g12582(.dina(n12827),.dinb(n12771),.dout(n12828),.clk(gclk));
	jand g12583(.dina(n12828),.dinb(w_n6357_34[0]),.dout(n12829),.clk(gclk));
	jnot g12584(.din(w_n12506_0[0]),.dout(n12830),.clk(gclk));
	jor g12585(.dina(w_n12830_0[1]),.dinb(n12829),.dout(n12831),.clk(gclk));
	jand g12586(.dina(n12831),.dinb(n12770),.dout(n12832),.clk(gclk));
	jand g12587(.dina(n12832),.dinb(w_n5989_30[0]),.dout(n12833),.clk(gclk));
	jor g12588(.dina(w_n12513_0[0]),.dinb(n12833),.dout(n12834),.clk(gclk));
	jand g12589(.dina(n12834),.dinb(n12769),.dout(n12835),.clk(gclk));
	jand g12590(.dina(n12835),.dinb(w_n5606_34[1]),.dout(n12836),.clk(gclk));
	jor g12591(.dina(w_n12521_0[0]),.dinb(n12836),.dout(n12837),.clk(gclk));
	jand g12592(.dina(n12837),.dinb(n12768),.dout(n12838),.clk(gclk));
	jand g12593(.dina(n12838),.dinb(w_n5259_31[0]),.dout(n12839),.clk(gclk));
	jor g12594(.dina(w_n12529_0[0]),.dinb(n12839),.dout(n12840),.clk(gclk));
	jand g12595(.dina(n12840),.dinb(n12767),.dout(n12841),.clk(gclk));
	jand g12596(.dina(n12841),.dinb(w_n4902_35[0]),.dout(n12842),.clk(gclk));
	jnot g12597(.din(w_n12537_0[0]),.dout(n12843),.clk(gclk));
	jor g12598(.dina(w_n12843_0[1]),.dinb(n12842),.dout(n12844),.clk(gclk));
	jand g12599(.dina(n12844),.dinb(n12766),.dout(n12845),.clk(gclk));
	jand g12600(.dina(n12845),.dinb(w_n4582_32[0]),.dout(n12846),.clk(gclk));
	jor g12601(.dina(w_n12544_0[0]),.dinb(n12846),.dout(n12847),.clk(gclk));
	jand g12602(.dina(n12847),.dinb(n12765),.dout(n12848),.clk(gclk));
	jand g12603(.dina(n12848),.dinb(w_n4249_35[2]),.dout(n12849),.clk(gclk));
	jor g12604(.dina(w_n12552_0[0]),.dinb(n12849),.dout(n12850),.clk(gclk));
	jand g12605(.dina(n12850),.dinb(n12764),.dout(n12851),.clk(gclk));
	jand g12606(.dina(n12851),.dinb(w_n3955_32[2]),.dout(n12852),.clk(gclk));
	jor g12607(.dina(w_n12560_0[0]),.dinb(n12852),.dout(n12853),.clk(gclk));
	jand g12608(.dina(n12853),.dinb(n12763),.dout(n12854),.clk(gclk));
	jand g12609(.dina(n12854),.dinb(w_n3642_36[0]),.dout(n12855),.clk(gclk));
	jor g12610(.dina(w_n12568_0[0]),.dinb(n12855),.dout(n12856),.clk(gclk));
	jand g12611(.dina(n12856),.dinb(n12762),.dout(n12857),.clk(gclk));
	jand g12612(.dina(n12857),.dinb(w_n3368_33[1]),.dout(n12858),.clk(gclk));
	jor g12613(.dina(w_n12576_0[1]),.dinb(n12858),.dout(n12859),.clk(gclk));
	jand g12614(.dina(n12859),.dinb(n12761),.dout(n12860),.clk(gclk));
	jand g12615(.dina(n12860),.dinb(w_n3089_36[2]),.dout(n12861),.clk(gclk));
	jor g12616(.dina(n12861),.dinb(w_n12760_0[1]),.dout(n12862),.clk(gclk));
	jand g12617(.dina(n12862),.dinb(n12759),.dout(n12863),.clk(gclk));
	jand g12618(.dina(n12863),.dinb(w_n2833_34[1]),.dout(n12864),.clk(gclk));
	jor g12619(.dina(w_n12591_0[0]),.dinb(n12864),.dout(n12865),.clk(gclk));
	jand g12620(.dina(n12865),.dinb(n12758),.dout(n12866),.clk(gclk));
	jand g12621(.dina(n12866),.dinb(w_n2572_37[0]),.dout(n12867),.clk(gclk));
	jnot g12622(.din(w_n12599_0[0]),.dout(n12868),.clk(gclk));
	jor g12623(.dina(w_n12868_0[1]),.dinb(n12867),.dout(n12869),.clk(gclk));
	jand g12624(.dina(n12869),.dinb(n12757),.dout(n12870),.clk(gclk));
	jand g12625(.dina(n12870),.dinb(w_n2345_35[0]),.dout(n12871),.clk(gclk));
	jor g12626(.dina(w_n12606_0[0]),.dinb(n12871),.dout(n12872),.clk(gclk));
	jand g12627(.dina(n12872),.dinb(n12756),.dout(n12873),.clk(gclk));
	jand g12628(.dina(n12873),.dinb(w_n2108_37[2]),.dout(n12874),.clk(gclk));
	jnot g12629(.din(w_n12614_0[0]),.dout(n12875),.clk(gclk));
	jor g12630(.dina(w_n12875_0[1]),.dinb(n12874),.dout(n12876),.clk(gclk));
	jand g12631(.dina(n12876),.dinb(n12755),.dout(n12877),.clk(gclk));
	jand g12632(.dina(n12877),.dinb(w_n1912_36[0]),.dout(n12878),.clk(gclk));
	jor g12633(.dina(w_n12621_0[0]),.dinb(n12878),.dout(n12879),.clk(gclk));
	jand g12634(.dina(n12879),.dinb(n12754),.dout(n12880),.clk(gclk));
	jand g12635(.dina(n12880),.dinb(w_n1699_38[1]),.dout(n12881),.clk(gclk));
	jor g12636(.dina(w_n12629_0[0]),.dinb(n12881),.dout(n12882),.clk(gclk));
	jand g12637(.dina(n12882),.dinb(n12753),.dout(n12883),.clk(gclk));
	jand g12638(.dina(n12883),.dinb(w_n1516_36[2]),.dout(n12884),.clk(gclk));
	jor g12639(.dina(w_n12637_0[0]),.dinb(n12884),.dout(n12885),.clk(gclk));
	jand g12640(.dina(n12885),.dinb(n12752),.dout(n12886),.clk(gclk));
	jand g12641(.dina(n12886),.dinb(w_n1332_38[1]),.dout(n12887),.clk(gclk));
	jnot g12642(.din(w_n12645_0[0]),.dout(n12888),.clk(gclk));
	jor g12643(.dina(w_n12888_0[1]),.dinb(n12887),.dout(n12889),.clk(gclk));
	jand g12644(.dina(n12889),.dinb(n12751),.dout(n12890),.clk(gclk));
	jand g12645(.dina(n12890),.dinb(w_n1173_37[1]),.dout(n12891),.clk(gclk));
	jor g12646(.dina(w_n12652_0[0]),.dinb(n12891),.dout(n12892),.clk(gclk));
	jand g12647(.dina(n12892),.dinb(n12750),.dout(n12893),.clk(gclk));
	jand g12648(.dina(n12893),.dinb(w_n1008_39[1]),.dout(n12894),.clk(gclk));
	jnot g12649(.din(w_n12660_0[0]),.dout(n12895),.clk(gclk));
	jor g12650(.dina(w_n12895_0[1]),.dinb(n12894),.dout(n12896),.clk(gclk));
	jand g12651(.dina(n12896),.dinb(n12749),.dout(n12897),.clk(gclk));
	jand g12652(.dina(n12897),.dinb(w_n884_38[1]),.dout(n12898),.clk(gclk));
	jor g12653(.dina(w_n12667_0[0]),.dinb(n12898),.dout(n12899),.clk(gclk));
	jand g12654(.dina(n12899),.dinb(n12748),.dout(n12900),.clk(gclk));
	jand g12655(.dina(n12900),.dinb(w_n743_39[1]),.dout(n12901),.clk(gclk));
	jnot g12656(.din(w_n12675_0[0]),.dout(n12902),.clk(gclk));
	jor g12657(.dina(w_n12902_0[1]),.dinb(n12901),.dout(n12903),.clk(gclk));
	jand g12658(.dina(n12903),.dinb(n12747),.dout(n12904),.clk(gclk));
	jand g12659(.dina(n12904),.dinb(w_n635_39[1]),.dout(n12905),.clk(gclk));
	jor g12660(.dina(w_n12682_0[0]),.dinb(n12905),.dout(n12906),.clk(gclk));
	jand g12661(.dina(n12906),.dinb(n12746),.dout(n12907),.clk(gclk));
	jand g12662(.dina(n12907),.dinb(w_n515_40[1]),.dout(n12908),.clk(gclk));
	jnot g12663(.din(w_n12690_0[0]),.dout(n12909),.clk(gclk));
	jor g12664(.dina(w_n12909_0[1]),.dinb(n12908),.dout(n12910),.clk(gclk));
	jand g12665(.dina(n12910),.dinb(n12745),.dout(n12911),.clk(gclk));
	jand g12666(.dina(n12911),.dinb(w_n443_40[1]),.dout(n12912),.clk(gclk));
	jnot g12667(.din(w_n12697_0[0]),.dout(n12913),.clk(gclk));
	jor g12668(.dina(w_n12913_0[1]),.dinb(n12912),.dout(n12914),.clk(gclk));
	jand g12669(.dina(n12914),.dinb(n12744),.dout(n12915),.clk(gclk));
	jand g12670(.dina(n12915),.dinb(w_n352_40[2]),.dout(n12916),.clk(gclk));
	jnot g12671(.din(w_n12704_0[0]),.dout(n12917),.clk(gclk));
	jor g12672(.dina(w_n12917_0[1]),.dinb(n12916),.dout(n12918),.clk(gclk));
	jand g12673(.dina(n12918),.dinb(n12743),.dout(n12919),.clk(gclk));
	jand g12674(.dina(n12919),.dinb(w_n294_41[0]),.dout(n12920),.clk(gclk));
	jor g12675(.dina(w_n12711_0[0]),.dinb(n12920),.dout(n12921),.clk(gclk));
	jand g12676(.dina(n12921),.dinb(n12742),.dout(n12922),.clk(gclk));
	jand g12677(.dina(n12922),.dinb(w_n239_41[0]),.dout(n12923),.clk(gclk));
	jor g12678(.dina(w_n12719_0[0]),.dinb(n12923),.dout(n12924),.clk(gclk));
	jand g12679(.dina(n12924),.dinb(n12741),.dout(n12925),.clk(gclk));
	jand g12680(.dina(n12925),.dinb(w_n221_41[1]),.dout(n12926),.clk(gclk));
	jor g12681(.dina(w_n12727_0[1]),.dinb(n12926),.dout(n12927),.clk(gclk));
	jand g12682(.dina(n12927),.dinb(n12740),.dout(n12928),.clk(gclk));
	jor g12683(.dina(w_n12928_0[1]),.dinb(w_n12739_0[1]),.dout(n12929),.clk(gclk));
	jor g12684(.dina(w_n12929_0[1]),.dinb(w_n12177_0[0]),.dout(n12930),.clk(gclk));
	jor g12685(.dina(n12930),.dinb(w_n12738_0[1]),.dout(n12931),.clk(gclk));
	jand g12686(.dina(n12931),.dinb(w_n218_17[1]),.dout(n12932),.clk(gclk));
	jand g12687(.dina(w_n12410_24[1]),.dinb(w_n11862_0[0]),.dout(n12933),.clk(gclk));
	jor g12688(.dina(w_n12933_0[1]),.dinb(w_n12932_0[1]),.dout(n12934),.clk(gclk));
	jor g12689(.dina(n12934),.dinb(w_n12737_0[1]),.dout(n12935),.clk(gclk));
	jor g12690(.dina(w_n12935_0[1]),.dinb(w_n12732_0[2]),.dout(asqrt_fa_20),.clk(gclk));
	jand g12691(.dina(w_n12730_0[0]),.dinb(w_n12195_0[0]),.dout(n12937),.clk(gclk));
	jand g12692(.dina(w_n12935_0[0]),.dinb(w_n12937_0[1]),.dout(n12938),.clk(gclk));
	jnot g12693(.din(w_n12737_0[0]),.dout(n12939),.clk(gclk));
	jnot g12694(.din(w_n12738_0[0]),.dout(n12940),.clk(gclk));
	jand g12695(.dina(w_n12937_0[0]),.dinb(w_n12207_0[1]),.dout(n12941),.clk(gclk));
	jand g12696(.dina(n12941),.dinb(n12940),.dout(n12942),.clk(gclk));
	jor g12697(.dina(n12942),.dinb(w_asqrt63_30[1]),.dout(n12943),.clk(gclk));
	jnot g12698(.din(w_n12933_0[0]),.dout(n12944),.clk(gclk));
	jand g12699(.dina(n12944),.dinb(n12943),.dout(n12945),.clk(gclk));
	jand g12700(.dina(n12945),.dinb(n12939),.dout(n12946),.clk(gclk));
	jand g12701(.dina(w_n12946_0[1]),.dinb(w_n12731_1[0]),.dout(n12947),.clk(gclk));
	jxor g12702(.dina(w_n12722_0[0]),.dinb(w_n221_41[0]),.dout(n12948),.clk(gclk));
	jor g12703(.dina(n12948),.dinb(w_n12947_44[2]),.dout(n12949),.clk(gclk));
	jxor g12704(.dina(n12949),.dinb(w_n12727_0[0]),.dout(n12950),.clk(gclk));
	jnot g12705(.din(w_n12950_0[1]),.dout(n12951),.clk(gclk));
	jor g12706(.dina(w_n12947_44[1]),.dinb(w_n12196_1[1]),.dout(n12952),.clk(gclk));
	jnot g12707(.din(w_a36_0[2]),.dout(n12953),.clk(gclk));
	jnot g12708(.din(w_a37_0[1]),.dout(n12954),.clk(gclk));
	jand g12709(.dina(w_n12954_0[1]),.dinb(w_n12953_1[2]),.dout(n12955),.clk(gclk));
	jand g12710(.dina(w_n12955_0[2]),.dinb(w_n12196_1[0]),.dout(n12956),.clk(gclk));
	jnot g12711(.din(w_n12956_0[1]),.dout(n12957),.clk(gclk));
	jand g12712(.dina(n12957),.dinb(n12952),.dout(n12958),.clk(gclk));
	jor g12713(.dina(w_n12958_0[2]),.dinb(w_n12410_24[0]),.dout(n12959),.clk(gclk));
	jand g12714(.dina(w_n12958_0[1]),.dinb(w_n12410_23[2]),.dout(n12960),.clk(gclk));
	jor g12715(.dina(w_n12947_44[0]),.dinb(w_a38_0[1]),.dout(n12961),.clk(gclk));
	jand g12716(.dina(n12961),.dinb(w_a39_0[0]),.dout(n12962),.clk(gclk));
	jand g12717(.dina(w_asqrt19_14),.dinb(w_n12198_0[1]),.dout(n12963),.clk(gclk));
	jor g12718(.dina(n12963),.dinb(n12962),.dout(n12964),.clk(gclk));
	jor g12719(.dina(w_n12964_0[1]),.dinb(n12960),.dout(n12965),.clk(gclk));
	jand g12720(.dina(n12965),.dinb(w_n12959_0[1]),.dout(n12966),.clk(gclk));
	jor g12721(.dina(w_n12966_0[2]),.dinb(w_n11858_30[2]),.dout(n12967),.clk(gclk));
	jand g12722(.dina(w_n12966_0[1]),.dinb(w_n11858_30[1]),.dout(n12968),.clk(gclk));
	jnot g12723(.din(w_n12198_0[0]),.dout(n12969),.clk(gclk));
	jor g12724(.dina(w_n12947_43[2]),.dinb(n12969),.dout(n12970),.clk(gclk));
	jor g12725(.dina(w_n12732_0[1]),.dinb(w_n12410_23[1]),.dout(n12971),.clk(gclk));
	jor g12726(.dina(n12971),.dinb(w_n12736_0[0]),.dout(n12972),.clk(gclk));
	jor g12727(.dina(n12972),.dinb(w_n12932_0[0]),.dout(n12973),.clk(gclk));
	jand g12728(.dina(n12973),.dinb(w_n12970_0[1]),.dout(n12974),.clk(gclk));
	jxor g12729(.dina(n12974),.dinb(w_n11864_0[1]),.dout(n12975),.clk(gclk));
	jor g12730(.dina(w_n12975_0[2]),.dinb(n12968),.dout(n12976),.clk(gclk));
	jand g12731(.dina(n12976),.dinb(w_n12967_0[1]),.dout(n12977),.clk(gclk));
	jor g12732(.dina(w_n12977_0[2]),.dinb(w_n11347_24[2]),.dout(n12978),.clk(gclk));
	jand g12733(.dina(w_n12977_0[1]),.dinb(w_n11347_24[1]),.dout(n12979),.clk(gclk));
	jxor g12734(.dina(w_n12201_0[0]),.dinb(w_n11858_30[0]),.dout(n12980),.clk(gclk));
	jor g12735(.dina(n12980),.dinb(w_n12947_43[1]),.dout(n12981),.clk(gclk));
	jxor g12736(.dina(n12981),.dinb(w_n12789_0[0]),.dout(n12982),.clk(gclk));
	jnot g12737(.din(w_n12982_0[2]),.dout(n12983),.clk(gclk));
	jor g12738(.dina(n12983),.dinb(n12979),.dout(n12984),.clk(gclk));
	jand g12739(.dina(n12984),.dinb(w_n12978_0[1]),.dout(n12985),.clk(gclk));
	jor g12740(.dina(w_n12985_0[2]),.dinb(w_n10824_31[1]),.dout(n12986),.clk(gclk));
	jand g12741(.dina(w_n12985_0[1]),.dinb(w_n10824_31[0]),.dout(n12987),.clk(gclk));
	jxor g12742(.dina(w_n12414_0[0]),.dinb(w_n11347_24[0]),.dout(n12988),.clk(gclk));
	jor g12743(.dina(n12988),.dinb(w_n12947_43[0]),.dout(n12989),.clk(gclk));
	jxor g12744(.dina(n12989),.dinb(w_n12423_0[0]),.dout(n12990),.clk(gclk));
	jor g12745(.dina(w_n12990_0[2]),.dinb(n12987),.dout(n12991),.clk(gclk));
	jand g12746(.dina(n12991),.dinb(w_n12986_0[1]),.dout(n12992),.clk(gclk));
	jor g12747(.dina(w_n12992_0[2]),.dinb(w_n10328_25[2]),.dout(n12993),.clk(gclk));
	jand g12748(.dina(w_n12992_0[1]),.dinb(w_n10328_25[1]),.dout(n12994),.clk(gclk));
	jxor g12749(.dina(w_n12425_0[0]),.dinb(w_n10824_30[2]),.dout(n12995),.clk(gclk));
	jor g12750(.dina(n12995),.dinb(w_n12947_42[2]),.dout(n12996),.clk(gclk));
	jxor g12751(.dina(n12996),.dinb(w_n12796_0[0]),.dout(n12997),.clk(gclk));
	jnot g12752(.din(w_n12997_0[2]),.dout(n12998),.clk(gclk));
	jor g12753(.dina(n12998),.dinb(n12994),.dout(n12999),.clk(gclk));
	jand g12754(.dina(n12999),.dinb(w_n12993_0[1]),.dout(n13000),.clk(gclk));
	jor g12755(.dina(w_n13000_0[2]),.dinb(w_n9832_32[0]),.dout(n13001),.clk(gclk));
	jand g12756(.dina(w_n13000_0[1]),.dinb(w_n9832_31[2]),.dout(n13002),.clk(gclk));
	jxor g12757(.dina(w_n12432_0[0]),.dinb(w_n10328_25[0]),.dout(n13003),.clk(gclk));
	jor g12758(.dina(n13003),.dinb(w_n12947_42[1]),.dout(n13004),.clk(gclk));
	jxor g12759(.dina(n13004),.dinb(w_n12438_0[0]),.dout(n13005),.clk(gclk));
	jor g12760(.dina(w_n13005_0[2]),.dinb(n13002),.dout(n13006),.clk(gclk));
	jand g12761(.dina(n13006),.dinb(w_n13001_0[1]),.dout(n13007),.clk(gclk));
	jor g12762(.dina(w_n13007_0[2]),.dinb(w_n9369_26[2]),.dout(n13008),.clk(gclk));
	jand g12763(.dina(w_n13007_0[1]),.dinb(w_n9369_26[1]),.dout(n13009),.clk(gclk));
	jxor g12764(.dina(w_n12440_0[0]),.dinb(w_n9832_31[1]),.dout(n13010),.clk(gclk));
	jor g12765(.dina(n13010),.dinb(w_n12947_42[0]),.dout(n13011),.clk(gclk));
	jxor g12766(.dina(n13011),.dinb(w_n12803_0[0]),.dout(n13012),.clk(gclk));
	jnot g12767(.din(w_n13012_0[2]),.dout(n13013),.clk(gclk));
	jor g12768(.dina(n13013),.dinb(n13009),.dout(n13014),.clk(gclk));
	jand g12769(.dina(n13014),.dinb(w_n13008_0[1]),.dout(n13015),.clk(gclk));
	jor g12770(.dina(w_n13015_0[2]),.dinb(w_n8890_32[1]),.dout(n13016),.clk(gclk));
	jand g12771(.dina(w_n13015_0[1]),.dinb(w_n8890_32[0]),.dout(n13017),.clk(gclk));
	jxor g12772(.dina(w_n12447_0[0]),.dinb(w_n9369_26[0]),.dout(n13018),.clk(gclk));
	jor g12773(.dina(n13018),.dinb(w_n12947_41[2]),.dout(n13019),.clk(gclk));
	jxor g12774(.dina(n13019),.dinb(w_n12453_0[0]),.dout(n13020),.clk(gclk));
	jor g12775(.dina(w_n13020_0[2]),.dinb(n13017),.dout(n13021),.clk(gclk));
	jand g12776(.dina(n13021),.dinb(w_n13016_0[1]),.dout(n13022),.clk(gclk));
	jor g12777(.dina(w_n13022_0[2]),.dinb(w_n8449_27[1]),.dout(n13023),.clk(gclk));
	jand g12778(.dina(w_n13022_0[1]),.dinb(w_n8449_27[0]),.dout(n13024),.clk(gclk));
	jxor g12779(.dina(w_n12455_0[0]),.dinb(w_n8890_31[2]),.dout(n13025),.clk(gclk));
	jor g12780(.dina(n13025),.dinb(w_n12947_41[1]),.dout(n13026),.clk(gclk));
	jxor g12781(.dina(n13026),.dinb(w_n12810_0[0]),.dout(n13027),.clk(gclk));
	jnot g12782(.din(w_n13027_0[2]),.dout(n13028),.clk(gclk));
	jor g12783(.dina(n13028),.dinb(n13024),.dout(n13029),.clk(gclk));
	jand g12784(.dina(n13029),.dinb(w_n13023_0[1]),.dout(n13030),.clk(gclk));
	jor g12785(.dina(w_n13030_0[2]),.dinb(w_n8003_33[0]),.dout(n13031),.clk(gclk));
	jand g12786(.dina(w_n13030_0[1]),.dinb(w_n8003_32[2]),.dout(n13032),.clk(gclk));
	jxor g12787(.dina(w_n12462_0[0]),.dinb(w_n8449_26[2]),.dout(n13033),.clk(gclk));
	jor g12788(.dina(n13033),.dinb(w_n12947_41[0]),.dout(n13034),.clk(gclk));
	jxor g12789(.dina(n13034),.dinb(w_n12468_0[0]),.dout(n13035),.clk(gclk));
	jor g12790(.dina(w_n13035_0[2]),.dinb(n13032),.dout(n13036),.clk(gclk));
	jand g12791(.dina(n13036),.dinb(w_n13031_0[1]),.dout(n13037),.clk(gclk));
	jor g12792(.dina(w_n13037_0[2]),.dinb(w_n7581_28[1]),.dout(n13038),.clk(gclk));
	jand g12793(.dina(w_n13037_0[1]),.dinb(w_n7581_28[0]),.dout(n13039),.clk(gclk));
	jxor g12794(.dina(w_n12470_0[0]),.dinb(w_n8003_32[1]),.dout(n13040),.clk(gclk));
	jor g12795(.dina(n13040),.dinb(w_n12947_40[2]),.dout(n13041),.clk(gclk));
	jxor g12796(.dina(n13041),.dinb(w_n12476_0[0]),.dout(n13042),.clk(gclk));
	jor g12797(.dina(w_n13042_0[2]),.dinb(n13039),.dout(n13043),.clk(gclk));
	jand g12798(.dina(n13043),.dinb(w_n13038_0[1]),.dout(n13044),.clk(gclk));
	jor g12799(.dina(w_n13044_0[2]),.dinb(w_n7154_33[1]),.dout(n13045),.clk(gclk));
	jand g12800(.dina(w_n13044_0[1]),.dinb(w_n7154_33[0]),.dout(n13046),.clk(gclk));
	jxor g12801(.dina(w_n12478_0[0]),.dinb(w_n7581_27[2]),.dout(n13047),.clk(gclk));
	jor g12802(.dina(n13047),.dinb(w_n12947_40[1]),.dout(n13048),.clk(gclk));
	jxor g12803(.dina(n13048),.dinb(w_n12484_0[0]),.dout(n13049),.clk(gclk));
	jor g12804(.dina(w_n13049_0[2]),.dinb(n13046),.dout(n13050),.clk(gclk));
	jand g12805(.dina(n13050),.dinb(w_n13045_0[1]),.dout(n13051),.clk(gclk));
	jor g12806(.dina(w_n13051_0[2]),.dinb(w_n6758_29[0]),.dout(n13052),.clk(gclk));
	jand g12807(.dina(w_n13051_0[1]),.dinb(w_n6758_28[2]),.dout(n13053),.clk(gclk));
	jxor g12808(.dina(w_n12486_0[0]),.dinb(w_n7154_32[2]),.dout(n13054),.clk(gclk));
	jor g12809(.dina(n13054),.dinb(w_n12947_40[0]),.dout(n13055),.clk(gclk));
	jxor g12810(.dina(n13055),.dinb(w_n12823_0[0]),.dout(n13056),.clk(gclk));
	jnot g12811(.din(w_n13056_0[2]),.dout(n13057),.clk(gclk));
	jor g12812(.dina(n13057),.dinb(n13053),.dout(n13058),.clk(gclk));
	jand g12813(.dina(n13058),.dinb(w_n13052_0[1]),.dout(n13059),.clk(gclk));
	jor g12814(.dina(w_n13059_0[2]),.dinb(w_n6357_33[2]),.dout(n13060),.clk(gclk));
	jand g12815(.dina(w_n13059_0[1]),.dinb(w_n6357_33[1]),.dout(n13061),.clk(gclk));
	jxor g12816(.dina(w_n12493_0[0]),.dinb(w_n6758_28[1]),.dout(n13062),.clk(gclk));
	jor g12817(.dina(n13062),.dinb(w_n12947_39[2]),.dout(n13063),.clk(gclk));
	jxor g12818(.dina(n13063),.dinb(w_n12499_0[0]),.dout(n13064),.clk(gclk));
	jor g12819(.dina(w_n13064_0[2]),.dinb(n13061),.dout(n13065),.clk(gclk));
	jand g12820(.dina(n13065),.dinb(w_n13060_0[1]),.dout(n13066),.clk(gclk));
	jor g12821(.dina(w_n13066_0[2]),.dinb(w_n5989_29[2]),.dout(n13067),.clk(gclk));
	jand g12822(.dina(w_n13066_0[1]),.dinb(w_n5989_29[1]),.dout(n13068),.clk(gclk));
	jxor g12823(.dina(w_n12501_0[0]),.dinb(w_n6357_33[0]),.dout(n13069),.clk(gclk));
	jor g12824(.dina(n13069),.dinb(w_n12947_39[1]),.dout(n13070),.clk(gclk));
	jxor g12825(.dina(n13070),.dinb(w_n12830_0[0]),.dout(n13071),.clk(gclk));
	jnot g12826(.din(w_n13071_0[2]),.dout(n13072),.clk(gclk));
	jor g12827(.dina(n13072),.dinb(n13068),.dout(n13073),.clk(gclk));
	jand g12828(.dina(n13073),.dinb(w_n13067_0[1]),.dout(n13074),.clk(gclk));
	jor g12829(.dina(w_n13074_0[2]),.dinb(w_n5606_34[0]),.dout(n13075),.clk(gclk));
	jand g12830(.dina(w_n13074_0[1]),.dinb(w_n5606_33[2]),.dout(n13076),.clk(gclk));
	jxor g12831(.dina(w_n12508_0[0]),.dinb(w_n5989_29[0]),.dout(n13077),.clk(gclk));
	jor g12832(.dina(n13077),.dinb(w_n12947_39[0]),.dout(n13078),.clk(gclk));
	jxor g12833(.dina(n13078),.dinb(w_n12514_0[0]),.dout(n13079),.clk(gclk));
	jor g12834(.dina(w_n13079_0[2]),.dinb(n13076),.dout(n13080),.clk(gclk));
	jand g12835(.dina(n13080),.dinb(w_n13075_0[1]),.dout(n13081),.clk(gclk));
	jor g12836(.dina(w_n13081_0[2]),.dinb(w_n5259_30[2]),.dout(n13082),.clk(gclk));
	jand g12837(.dina(w_n13081_0[1]),.dinb(w_n5259_30[1]),.dout(n13083),.clk(gclk));
	jxor g12838(.dina(w_n12516_0[0]),.dinb(w_n5606_33[1]),.dout(n13084),.clk(gclk));
	jor g12839(.dina(n13084),.dinb(w_n12947_38[2]),.dout(n13085),.clk(gclk));
	jxor g12840(.dina(n13085),.dinb(w_n12522_0[0]),.dout(n13086),.clk(gclk));
	jor g12841(.dina(w_n13086_0[2]),.dinb(n13083),.dout(n13087),.clk(gclk));
	jand g12842(.dina(n13087),.dinb(w_n13082_0[1]),.dout(n13088),.clk(gclk));
	jor g12843(.dina(w_n13088_0[2]),.dinb(w_n4902_34[2]),.dout(n13089),.clk(gclk));
	jand g12844(.dina(w_n13088_0[1]),.dinb(w_n4902_34[1]),.dout(n13090),.clk(gclk));
	jxor g12845(.dina(w_n12524_0[0]),.dinb(w_n5259_30[0]),.dout(n13091),.clk(gclk));
	jor g12846(.dina(n13091),.dinb(w_n12947_38[1]),.dout(n13092),.clk(gclk));
	jxor g12847(.dina(n13092),.dinb(w_n12530_0[0]),.dout(n13093),.clk(gclk));
	jor g12848(.dina(w_n13093_0[2]),.dinb(n13090),.dout(n13094),.clk(gclk));
	jand g12849(.dina(n13094),.dinb(w_n13089_0[1]),.dout(n13095),.clk(gclk));
	jor g12850(.dina(w_n13095_0[2]),.dinb(w_n4582_31[2]),.dout(n13096),.clk(gclk));
	jand g12851(.dina(w_n13095_0[1]),.dinb(w_n4582_31[1]),.dout(n13097),.clk(gclk));
	jxor g12852(.dina(w_n12532_0[0]),.dinb(w_n4902_34[0]),.dout(n13098),.clk(gclk));
	jor g12853(.dina(n13098),.dinb(w_n12947_38[0]),.dout(n13099),.clk(gclk));
	jxor g12854(.dina(n13099),.dinb(w_n12843_0[0]),.dout(n13100),.clk(gclk));
	jnot g12855(.din(w_n13100_0[2]),.dout(n13101),.clk(gclk));
	jor g12856(.dina(n13101),.dinb(n13097),.dout(n13102),.clk(gclk));
	jand g12857(.dina(n13102),.dinb(w_n13096_0[1]),.dout(n13103),.clk(gclk));
	jor g12858(.dina(w_n13103_0[2]),.dinb(w_n4249_35[1]),.dout(n13104),.clk(gclk));
	jand g12859(.dina(w_n13103_0[1]),.dinb(w_n4249_35[0]),.dout(n13105),.clk(gclk));
	jxor g12860(.dina(w_n12539_0[0]),.dinb(w_n4582_31[0]),.dout(n13106),.clk(gclk));
	jor g12861(.dina(n13106),.dinb(w_n12947_37[2]),.dout(n13107),.clk(gclk));
	jxor g12862(.dina(n13107),.dinb(w_n12545_0[0]),.dout(n13108),.clk(gclk));
	jor g12863(.dina(w_n13108_0[2]),.dinb(n13105),.dout(n13109),.clk(gclk));
	jand g12864(.dina(n13109),.dinb(w_n13104_0[1]),.dout(n13110),.clk(gclk));
	jor g12865(.dina(w_n13110_0[2]),.dinb(w_n3955_32[1]),.dout(n13111),.clk(gclk));
	jand g12866(.dina(w_n13110_0[1]),.dinb(w_n3955_32[0]),.dout(n13112),.clk(gclk));
	jxor g12867(.dina(w_n12547_0[0]),.dinb(w_n4249_34[2]),.dout(n13113),.clk(gclk));
	jor g12868(.dina(n13113),.dinb(w_n12947_37[1]),.dout(n13114),.clk(gclk));
	jxor g12869(.dina(n13114),.dinb(w_n12553_0[0]),.dout(n13115),.clk(gclk));
	jor g12870(.dina(w_n13115_0[2]),.dinb(n13112),.dout(n13116),.clk(gclk));
	jand g12871(.dina(n13116),.dinb(w_n13111_0[1]),.dout(n13117),.clk(gclk));
	jor g12872(.dina(w_n13117_0[2]),.dinb(w_n3642_35[2]),.dout(n13118),.clk(gclk));
	jand g12873(.dina(w_n13117_0[1]),.dinb(w_n3642_35[1]),.dout(n13119),.clk(gclk));
	jxor g12874(.dina(w_n12555_0[0]),.dinb(w_n3955_31[2]),.dout(n13120),.clk(gclk));
	jor g12875(.dina(n13120),.dinb(w_n12947_37[0]),.dout(n13121),.clk(gclk));
	jxor g12876(.dina(n13121),.dinb(w_n12561_0[0]),.dout(n13122),.clk(gclk));
	jor g12877(.dina(w_n13122_0[2]),.dinb(n13119),.dout(n13123),.clk(gclk));
	jand g12878(.dina(n13123),.dinb(w_n13118_0[1]),.dout(n13124),.clk(gclk));
	jor g12879(.dina(w_n13124_0[2]),.dinb(w_n3368_33[0]),.dout(n13125),.clk(gclk));
	jand g12880(.dina(w_n13124_0[1]),.dinb(w_n3368_32[2]),.dout(n13126),.clk(gclk));
	jxor g12881(.dina(w_n12563_0[0]),.dinb(w_n3642_35[0]),.dout(n13127),.clk(gclk));
	jor g12882(.dina(n13127),.dinb(w_n12947_36[2]),.dout(n13128),.clk(gclk));
	jxor g12883(.dina(n13128),.dinb(w_n12569_0[0]),.dout(n13129),.clk(gclk));
	jor g12884(.dina(w_n13129_0[2]),.dinb(n13126),.dout(n13130),.clk(gclk));
	jand g12885(.dina(n13130),.dinb(w_n13125_0[1]),.dout(n13131),.clk(gclk));
	jor g12886(.dina(w_n13131_0[2]),.dinb(w_n3089_36[1]),.dout(n13132),.clk(gclk));
	jand g12887(.dina(w_n13131_0[1]),.dinb(w_n3089_36[0]),.dout(n13133),.clk(gclk));
	jxor g12888(.dina(w_n12571_0[0]),.dinb(w_n3368_32[1]),.dout(n13134),.clk(gclk));
	jor g12889(.dina(n13134),.dinb(w_n12947_36[1]),.dout(n13135),.clk(gclk));
	jxor g12890(.dina(n13135),.dinb(w_n12576_0[0]),.dout(n13136),.clk(gclk));
	jnot g12891(.din(w_n13136_0[2]),.dout(n13137),.clk(gclk));
	jor g12892(.dina(n13137),.dinb(n13133),.dout(n13138),.clk(gclk));
	jand g12893(.dina(n13138),.dinb(w_n13132_0[1]),.dout(n13139),.clk(gclk));
	jor g12894(.dina(w_n13139_0[2]),.dinb(w_n2833_34[0]),.dout(n13140),.clk(gclk));
	jxor g12895(.dina(w_n12579_0[0]),.dinb(w_n3089_35[2]),.dout(n13141),.clk(gclk));
	jor g12896(.dina(n13141),.dinb(w_n12947_36[0]),.dout(n13142),.clk(gclk));
	jxor g12897(.dina(n13142),.dinb(w_n12760_0[0]),.dout(n13143),.clk(gclk));
	jnot g12898(.din(w_n13143_0[2]),.dout(n13144),.clk(gclk));
	jand g12899(.dina(w_n13139_0[1]),.dinb(w_n2833_33[2]),.dout(n13145),.clk(gclk));
	jor g12900(.dina(n13145),.dinb(n13144),.dout(n13146),.clk(gclk));
	jand g12901(.dina(n13146),.dinb(w_n13140_0[1]),.dout(n13147),.clk(gclk));
	jor g12902(.dina(w_n13147_0[2]),.dinb(w_n2572_36[2]),.dout(n13148),.clk(gclk));
	jand g12903(.dina(w_n13147_0[1]),.dinb(w_n2572_36[1]),.dout(n13149),.clk(gclk));
	jxor g12904(.dina(w_n12586_0[0]),.dinb(w_n2833_33[1]),.dout(n13150),.clk(gclk));
	jor g12905(.dina(n13150),.dinb(w_n12947_35[2]),.dout(n13151),.clk(gclk));
	jxor g12906(.dina(n13151),.dinb(w_n12592_0[0]),.dout(n13152),.clk(gclk));
	jor g12907(.dina(w_n13152_0[2]),.dinb(n13149),.dout(n13153),.clk(gclk));
	jand g12908(.dina(n13153),.dinb(w_n13148_0[1]),.dout(n13154),.clk(gclk));
	jor g12909(.dina(w_n13154_0[2]),.dinb(w_n2345_34[2]),.dout(n13155),.clk(gclk));
	jand g12910(.dina(w_n13154_0[1]),.dinb(w_n2345_34[1]),.dout(n13156),.clk(gclk));
	jxor g12911(.dina(w_n12594_0[0]),.dinb(w_n2572_36[0]),.dout(n13157),.clk(gclk));
	jor g12912(.dina(n13157),.dinb(w_n12947_35[1]),.dout(n13158),.clk(gclk));
	jxor g12913(.dina(n13158),.dinb(w_n12868_0[0]),.dout(n13159),.clk(gclk));
	jnot g12914(.din(w_n13159_0[2]),.dout(n13160),.clk(gclk));
	jor g12915(.dina(n13160),.dinb(n13156),.dout(n13161),.clk(gclk));
	jand g12916(.dina(n13161),.dinb(w_n13155_0[1]),.dout(n13162),.clk(gclk));
	jor g12917(.dina(w_n13162_0[2]),.dinb(w_n2108_37[1]),.dout(n13163),.clk(gclk));
	jand g12918(.dina(w_n13162_0[1]),.dinb(w_n2108_37[0]),.dout(n13164),.clk(gclk));
	jxor g12919(.dina(w_n12601_0[0]),.dinb(w_n2345_34[0]),.dout(n13165),.clk(gclk));
	jor g12920(.dina(n13165),.dinb(w_n12947_35[0]),.dout(n13166),.clk(gclk));
	jxor g12921(.dina(n13166),.dinb(w_n12607_0[0]),.dout(n13167),.clk(gclk));
	jor g12922(.dina(w_n13167_0[2]),.dinb(n13164),.dout(n13168),.clk(gclk));
	jand g12923(.dina(n13168),.dinb(w_n13163_0[1]),.dout(n13169),.clk(gclk));
	jor g12924(.dina(w_n13169_0[2]),.dinb(w_n1912_35[2]),.dout(n13170),.clk(gclk));
	jand g12925(.dina(w_n13169_0[1]),.dinb(w_n1912_35[1]),.dout(n13171),.clk(gclk));
	jxor g12926(.dina(w_n12609_0[0]),.dinb(w_n2108_36[2]),.dout(n13172),.clk(gclk));
	jor g12927(.dina(n13172),.dinb(w_n12947_34[2]),.dout(n13173),.clk(gclk));
	jxor g12928(.dina(n13173),.dinb(w_n12875_0[0]),.dout(n13174),.clk(gclk));
	jnot g12929(.din(w_n13174_0[2]),.dout(n13175),.clk(gclk));
	jor g12930(.dina(n13175),.dinb(n13171),.dout(n13176),.clk(gclk));
	jand g12931(.dina(n13176),.dinb(w_n13170_0[1]),.dout(n13177),.clk(gclk));
	jor g12932(.dina(w_n13177_0[2]),.dinb(w_n1699_38[0]),.dout(n13178),.clk(gclk));
	jand g12933(.dina(w_n13177_0[1]),.dinb(w_n1699_37[2]),.dout(n13179),.clk(gclk));
	jxor g12934(.dina(w_n12616_0[0]),.dinb(w_n1912_35[0]),.dout(n13180),.clk(gclk));
	jor g12935(.dina(n13180),.dinb(w_n12947_34[1]),.dout(n13181),.clk(gclk));
	jxor g12936(.dina(n13181),.dinb(w_n12622_0[0]),.dout(n13182),.clk(gclk));
	jor g12937(.dina(w_n13182_0[2]),.dinb(n13179),.dout(n13183),.clk(gclk));
	jand g12938(.dina(n13183),.dinb(w_n13178_0[1]),.dout(n13184),.clk(gclk));
	jor g12939(.dina(w_n13184_0[2]),.dinb(w_n1516_36[1]),.dout(n13185),.clk(gclk));
	jand g12940(.dina(w_n13184_0[1]),.dinb(w_n1516_36[0]),.dout(n13186),.clk(gclk));
	jxor g12941(.dina(w_n12624_0[0]),.dinb(w_n1699_37[1]),.dout(n13187),.clk(gclk));
	jor g12942(.dina(n13187),.dinb(w_n12947_34[0]),.dout(n13188),.clk(gclk));
	jxor g12943(.dina(n13188),.dinb(w_n12630_0[0]),.dout(n13189),.clk(gclk));
	jor g12944(.dina(w_n13189_0[2]),.dinb(n13186),.dout(n13190),.clk(gclk));
	jand g12945(.dina(n13190),.dinb(w_n13185_0[1]),.dout(n13191),.clk(gclk));
	jor g12946(.dina(w_n13191_0[2]),.dinb(w_n1332_38[0]),.dout(n13192),.clk(gclk));
	jand g12947(.dina(w_n13191_0[1]),.dinb(w_n1332_37[2]),.dout(n13193),.clk(gclk));
	jxor g12948(.dina(w_n12632_0[0]),.dinb(w_n1516_35[2]),.dout(n13194),.clk(gclk));
	jor g12949(.dina(n13194),.dinb(w_n12947_33[2]),.dout(n13195),.clk(gclk));
	jxor g12950(.dina(n13195),.dinb(w_n12638_0[0]),.dout(n13196),.clk(gclk));
	jor g12951(.dina(w_n13196_0[2]),.dinb(n13193),.dout(n13197),.clk(gclk));
	jand g12952(.dina(n13197),.dinb(w_n13192_0[1]),.dout(n13198),.clk(gclk));
	jor g12953(.dina(w_n13198_0[2]),.dinb(w_n1173_37[0]),.dout(n13199),.clk(gclk));
	jand g12954(.dina(w_n13198_0[1]),.dinb(w_n1173_36[2]),.dout(n13200),.clk(gclk));
	jxor g12955(.dina(w_n12640_0[0]),.dinb(w_n1332_37[1]),.dout(n13201),.clk(gclk));
	jor g12956(.dina(n13201),.dinb(w_n12947_33[1]),.dout(n13202),.clk(gclk));
	jxor g12957(.dina(n13202),.dinb(w_n12888_0[0]),.dout(n13203),.clk(gclk));
	jnot g12958(.din(w_n13203_0[2]),.dout(n13204),.clk(gclk));
	jor g12959(.dina(n13204),.dinb(n13200),.dout(n13205),.clk(gclk));
	jand g12960(.dina(n13205),.dinb(w_n13199_0[1]),.dout(n13206),.clk(gclk));
	jor g12961(.dina(w_n13206_0[2]),.dinb(w_n1008_39[0]),.dout(n13207),.clk(gclk));
	jand g12962(.dina(w_n13206_0[1]),.dinb(w_n1008_38[2]),.dout(n13208),.clk(gclk));
	jxor g12963(.dina(w_n12647_0[0]),.dinb(w_n1173_36[1]),.dout(n13209),.clk(gclk));
	jor g12964(.dina(n13209),.dinb(w_n12947_33[0]),.dout(n13210),.clk(gclk));
	jxor g12965(.dina(n13210),.dinb(w_n12653_0[0]),.dout(n13211),.clk(gclk));
	jor g12966(.dina(w_n13211_0[2]),.dinb(n13208),.dout(n13212),.clk(gclk));
	jand g12967(.dina(n13212),.dinb(w_n13207_0[1]),.dout(n13213),.clk(gclk));
	jor g12968(.dina(w_n13213_0[2]),.dinb(w_n884_38[0]),.dout(n13214),.clk(gclk));
	jand g12969(.dina(w_n13213_0[1]),.dinb(w_n884_37[2]),.dout(n13215),.clk(gclk));
	jxor g12970(.dina(w_n12655_0[0]),.dinb(w_n1008_38[1]),.dout(n13216),.clk(gclk));
	jor g12971(.dina(n13216),.dinb(w_n12947_32[2]),.dout(n13217),.clk(gclk));
	jxor g12972(.dina(n13217),.dinb(w_n12895_0[0]),.dout(n13218),.clk(gclk));
	jnot g12973(.din(w_n13218_0[2]),.dout(n13219),.clk(gclk));
	jor g12974(.dina(n13219),.dinb(n13215),.dout(n13220),.clk(gclk));
	jand g12975(.dina(n13220),.dinb(w_n13214_0[1]),.dout(n13221),.clk(gclk));
	jor g12976(.dina(w_n13221_0[2]),.dinb(w_n743_39[0]),.dout(n13222),.clk(gclk));
	jand g12977(.dina(w_n13221_0[1]),.dinb(w_n743_38[2]),.dout(n13223),.clk(gclk));
	jxor g12978(.dina(w_n12662_0[0]),.dinb(w_n884_37[1]),.dout(n13224),.clk(gclk));
	jor g12979(.dina(n13224),.dinb(w_n12947_32[1]),.dout(n13225),.clk(gclk));
	jxor g12980(.dina(n13225),.dinb(w_n12668_0[0]),.dout(n13226),.clk(gclk));
	jor g12981(.dina(w_n13226_0[2]),.dinb(n13223),.dout(n13227),.clk(gclk));
	jand g12982(.dina(n13227),.dinb(w_n13222_0[1]),.dout(n13228),.clk(gclk));
	jor g12983(.dina(w_n13228_0[2]),.dinb(w_n635_39[0]),.dout(n13229),.clk(gclk));
	jand g12984(.dina(w_n13228_0[1]),.dinb(w_n635_38[2]),.dout(n13230),.clk(gclk));
	jxor g12985(.dina(w_n12670_0[0]),.dinb(w_n743_38[1]),.dout(n13231),.clk(gclk));
	jor g12986(.dina(n13231),.dinb(w_n12947_32[0]),.dout(n13232),.clk(gclk));
	jxor g12987(.dina(n13232),.dinb(w_n12902_0[0]),.dout(n13233),.clk(gclk));
	jnot g12988(.din(w_n13233_0[2]),.dout(n13234),.clk(gclk));
	jor g12989(.dina(n13234),.dinb(n13230),.dout(n13235),.clk(gclk));
	jand g12990(.dina(n13235),.dinb(w_n13229_0[1]),.dout(n13236),.clk(gclk));
	jor g12991(.dina(w_n13236_0[2]),.dinb(w_n515_40[0]),.dout(n13237),.clk(gclk));
	jand g12992(.dina(w_n13236_0[1]),.dinb(w_n515_39[2]),.dout(n13238),.clk(gclk));
	jxor g12993(.dina(w_n12677_0[0]),.dinb(w_n635_38[1]),.dout(n13239),.clk(gclk));
	jor g12994(.dina(n13239),.dinb(w_n12947_31[2]),.dout(n13240),.clk(gclk));
	jxor g12995(.dina(n13240),.dinb(w_n12683_0[0]),.dout(n13241),.clk(gclk));
	jor g12996(.dina(w_n13241_0[2]),.dinb(n13238),.dout(n13242),.clk(gclk));
	jand g12997(.dina(n13242),.dinb(w_n13237_0[1]),.dout(n13243),.clk(gclk));
	jor g12998(.dina(w_n13243_0[2]),.dinb(w_n443_40[0]),.dout(n13244),.clk(gclk));
	jand g12999(.dina(w_n13243_0[1]),.dinb(w_n443_39[2]),.dout(n13245),.clk(gclk));
	jxor g13000(.dina(w_n12685_0[0]),.dinb(w_n515_39[1]),.dout(n13246),.clk(gclk));
	jor g13001(.dina(n13246),.dinb(w_n12947_31[1]),.dout(n13247),.clk(gclk));
	jxor g13002(.dina(n13247),.dinb(w_n12909_0[0]),.dout(n13248),.clk(gclk));
	jnot g13003(.din(w_n13248_0[2]),.dout(n13249),.clk(gclk));
	jor g13004(.dina(n13249),.dinb(n13245),.dout(n13250),.clk(gclk));
	jand g13005(.dina(n13250),.dinb(w_n13244_0[1]),.dout(n13251),.clk(gclk));
	jor g13006(.dina(w_n13251_0[2]),.dinb(w_n352_40[1]),.dout(n13252),.clk(gclk));
	jand g13007(.dina(w_n13251_0[1]),.dinb(w_n352_40[0]),.dout(n13253),.clk(gclk));
	jxor g13008(.dina(w_n12692_0[0]),.dinb(w_n443_39[1]),.dout(n13254),.clk(gclk));
	jor g13009(.dina(n13254),.dinb(w_n12947_31[0]),.dout(n13255),.clk(gclk));
	jxor g13010(.dina(n13255),.dinb(w_n12913_0[0]),.dout(n13256),.clk(gclk));
	jnot g13011(.din(w_n13256_0[2]),.dout(n13257),.clk(gclk));
	jor g13012(.dina(n13257),.dinb(n13253),.dout(n13258),.clk(gclk));
	jand g13013(.dina(n13258),.dinb(w_n13252_0[1]),.dout(n13259),.clk(gclk));
	jor g13014(.dina(w_n13259_0[2]),.dinb(w_n294_40[2]),.dout(n13260),.clk(gclk));
	jand g13015(.dina(w_n13259_0[1]),.dinb(w_n294_40[1]),.dout(n13261),.clk(gclk));
	jxor g13016(.dina(w_n12699_0[0]),.dinb(w_n352_39[2]),.dout(n13262),.clk(gclk));
	jor g13017(.dina(n13262),.dinb(w_n12947_30[2]),.dout(n13263),.clk(gclk));
	jxor g13018(.dina(n13263),.dinb(w_n12917_0[0]),.dout(n13264),.clk(gclk));
	jnot g13019(.din(w_n13264_0[2]),.dout(n13265),.clk(gclk));
	jor g13020(.dina(n13265),.dinb(n13261),.dout(n13266),.clk(gclk));
	jand g13021(.dina(n13266),.dinb(w_n13260_0[1]),.dout(n13267),.clk(gclk));
	jor g13022(.dina(w_n13267_0[2]),.dinb(w_n239_40[2]),.dout(n13268),.clk(gclk));
	jand g13023(.dina(w_n13267_0[1]),.dinb(w_n239_40[1]),.dout(n13269),.clk(gclk));
	jxor g13024(.dina(w_n12706_0[0]),.dinb(w_n294_40[0]),.dout(n13270),.clk(gclk));
	jor g13025(.dina(n13270),.dinb(w_n12947_30[1]),.dout(n13271),.clk(gclk));
	jxor g13026(.dina(n13271),.dinb(w_n12712_0[0]),.dout(n13272),.clk(gclk));
	jor g13027(.dina(w_n13272_0[2]),.dinb(n13269),.dout(n13273),.clk(gclk));
	jand g13028(.dina(n13273),.dinb(w_n13268_0[1]),.dout(n13274),.clk(gclk));
	jor g13029(.dina(w_n13274_0[2]),.dinb(w_n221_40[2]),.dout(n13275),.clk(gclk));
	jand g13030(.dina(w_n13274_0[1]),.dinb(w_n221_40[1]),.dout(n13276),.clk(gclk));
	jxor g13031(.dina(w_n12714_0[0]),.dinb(w_n239_40[0]),.dout(n13277),.clk(gclk));
	jor g13032(.dina(n13277),.dinb(w_n12947_30[0]),.dout(n13278),.clk(gclk));
	jxor g13033(.dina(n13278),.dinb(w_n12720_0[0]),.dout(n13279),.clk(gclk));
	jor g13034(.dina(w_n13279_0[2]),.dinb(n13276),.dout(n13280),.clk(gclk));
	jand g13035(.dina(n13280),.dinb(w_n13275_0[1]),.dout(n13281),.clk(gclk));
	jor g13036(.dina(w_n13281_0[2]),.dinb(w_n12951_0[2]),.dout(n13282),.clk(gclk));
	jor g13037(.dina(w_n13282_0[1]),.dinb(w_n12732_0[0]),.dout(n13283),.clk(gclk));
	jor g13038(.dina(n13283),.dinb(w_n12938_0[1]),.dout(n13284),.clk(gclk));
	jand g13039(.dina(n13284),.dinb(w_n218_17[0]),.dout(n13285),.clk(gclk));
	jand g13040(.dina(w_n12947_29[2]),.dinb(w_n12739_0[0]),.dout(n13286),.clk(gclk));
	jand g13041(.dina(w_n13281_0[1]),.dinb(w_n12951_0[1]),.dout(n13287),.clk(gclk));
	jor g13042(.dina(w_n13287_1[1]),.dinb(n13286),.dout(n13288),.clk(gclk));
	jand g13043(.dina(w_n12946_0[0]),.dinb(w_n12928_0[0]),.dout(n13289),.clk(gclk));
	jnot g13044(.din(n13289),.dout(n13290),.clk(gclk));
	jand g13045(.dina(w_n12929_0[0]),.dinb(w_asqrt63_30[0]),.dout(n13291),.clk(gclk));
	jand g13046(.dina(n13291),.dinb(w_n12731_0[2]),.dout(n13292),.clk(gclk));
	jand g13047(.dina(w_n13292_0[1]),.dinb(n13290),.dout(n13293),.clk(gclk));
	jor g13048(.dina(n13293),.dinb(n13288),.dout(n13294),.clk(gclk));
	jor g13049(.dina(w_n13294_0[1]),.dinb(w_n13285_0[1]),.dout(asqrt_fa_19),.clk(gclk));
	jnot g13050(.din(w_a34_1[1]),.dout(n13296),.clk(gclk));
	jnot g13051(.din(w_a35_0[1]),.dout(n13297),.clk(gclk));
	jand g13052(.dina(w_n13297_0[1]),.dinb(w_n13296_1[1]),.dout(n13298),.clk(gclk));
	jand g13053(.dina(w_n13298_0[2]),.dinb(w_n12953_1[1]),.dout(n13299),.clk(gclk));
	jand g13054(.dina(w_asqrt18_35),.dinb(w_a36_0[1]),.dout(n13300),.clk(gclk));
	jor g13055(.dina(n13300),.dinb(w_n13299_0[1]),.dout(n13301),.clk(gclk));
	jand g13056(.dina(w_n13301_0[2]),.dinb(w_asqrt19_13[2]),.dout(n13302),.clk(gclk));
	jor g13057(.dina(w_n13301_0[1]),.dinb(w_asqrt19_13[1]),.dout(n13303),.clk(gclk));
	jand g13058(.dina(w_asqrt18_34[2]),.dinb(w_n12953_1[0]),.dout(n13304),.clk(gclk));
	jor g13059(.dina(n13304),.dinb(w_n12954_0[0]),.dout(n13305),.clk(gclk));
	jnot g13060(.din(w_n12955_0[1]),.dout(n13306),.clk(gclk));
	jnot g13061(.din(w_n12938_0[0]),.dout(n13307),.clk(gclk));
	jnot g13062(.din(w_n13275_0[0]),.dout(n13308),.clk(gclk));
	jnot g13063(.din(w_n13268_0[0]),.dout(n13309),.clk(gclk));
	jnot g13064(.din(w_n13260_0[0]),.dout(n13310),.clk(gclk));
	jnot g13065(.din(w_n13252_0[0]),.dout(n13311),.clk(gclk));
	jnot g13066(.din(w_n13244_0[0]),.dout(n13312),.clk(gclk));
	jnot g13067(.din(w_n13237_0[0]),.dout(n13313),.clk(gclk));
	jnot g13068(.din(w_n13229_0[0]),.dout(n13314),.clk(gclk));
	jnot g13069(.din(w_n13222_0[0]),.dout(n13315),.clk(gclk));
	jnot g13070(.din(w_n13214_0[0]),.dout(n13316),.clk(gclk));
	jnot g13071(.din(w_n13207_0[0]),.dout(n13317),.clk(gclk));
	jnot g13072(.din(w_n13199_0[0]),.dout(n13318),.clk(gclk));
	jnot g13073(.din(w_n13192_0[0]),.dout(n13319),.clk(gclk));
	jnot g13074(.din(w_n13185_0[0]),.dout(n13320),.clk(gclk));
	jnot g13075(.din(w_n13178_0[0]),.dout(n13321),.clk(gclk));
	jnot g13076(.din(w_n13170_0[0]),.dout(n13322),.clk(gclk));
	jnot g13077(.din(w_n13163_0[0]),.dout(n13323),.clk(gclk));
	jnot g13078(.din(w_n13155_0[0]),.dout(n13324),.clk(gclk));
	jnot g13079(.din(w_n13148_0[0]),.dout(n13325),.clk(gclk));
	jnot g13080(.din(w_n13140_0[0]),.dout(n13326),.clk(gclk));
	jnot g13081(.din(w_n13132_0[0]),.dout(n13327),.clk(gclk));
	jnot g13082(.din(w_n13125_0[0]),.dout(n13328),.clk(gclk));
	jnot g13083(.din(w_n13118_0[0]),.dout(n13329),.clk(gclk));
	jnot g13084(.din(w_n13111_0[0]),.dout(n13330),.clk(gclk));
	jnot g13085(.din(w_n13104_0[0]),.dout(n13331),.clk(gclk));
	jnot g13086(.din(w_n13096_0[0]),.dout(n13332),.clk(gclk));
	jnot g13087(.din(w_n13089_0[0]),.dout(n13333),.clk(gclk));
	jnot g13088(.din(w_n13082_0[0]),.dout(n13334),.clk(gclk));
	jnot g13089(.din(w_n13075_0[0]),.dout(n13335),.clk(gclk));
	jnot g13090(.din(w_n13067_0[0]),.dout(n13336),.clk(gclk));
	jnot g13091(.din(w_n13060_0[0]),.dout(n13337),.clk(gclk));
	jnot g13092(.din(w_n13052_0[0]),.dout(n13338),.clk(gclk));
	jnot g13093(.din(w_n13045_0[0]),.dout(n13339),.clk(gclk));
	jnot g13094(.din(w_n13038_0[0]),.dout(n13340),.clk(gclk));
	jnot g13095(.din(w_n13031_0[0]),.dout(n13341),.clk(gclk));
	jnot g13096(.din(w_n13023_0[0]),.dout(n13342),.clk(gclk));
	jnot g13097(.din(w_n13016_0[0]),.dout(n13343),.clk(gclk));
	jnot g13098(.din(w_n13008_0[0]),.dout(n13344),.clk(gclk));
	jnot g13099(.din(w_n13001_0[0]),.dout(n13345),.clk(gclk));
	jnot g13100(.din(w_n12993_0[0]),.dout(n13346),.clk(gclk));
	jnot g13101(.din(w_n12986_0[0]),.dout(n13347),.clk(gclk));
	jnot g13102(.din(w_n12978_0[0]),.dout(n13348),.clk(gclk));
	jnot g13103(.din(w_n12967_0[0]),.dout(n13349),.clk(gclk));
	jnot g13104(.din(w_n12959_0[0]),.dout(n13350),.clk(gclk));
	jand g13105(.dina(w_asqrt19_13[0]),.dinb(w_a38_0[0]),.dout(n13351),.clk(gclk));
	jor g13106(.dina(w_n12956_0[0]),.dinb(n13351),.dout(n13352),.clk(gclk));
	jor g13107(.dina(n13352),.dinb(w_asqrt20_20[1]),.dout(n13353),.clk(gclk));
	jand g13108(.dina(w_asqrt19_12[2]),.dinb(w_n12196_0[2]),.dout(n13354),.clk(gclk));
	jor g13109(.dina(n13354),.dinb(w_n12197_0[0]),.dout(n13355),.clk(gclk));
	jand g13110(.dina(w_n12970_0[0]),.dinb(n13355),.dout(n13356),.clk(gclk));
	jand g13111(.dina(n13356),.dinb(n13353),.dout(n13357),.clk(gclk));
	jor g13112(.dina(n13357),.dinb(n13350),.dout(n13358),.clk(gclk));
	jor g13113(.dina(n13358),.dinb(w_asqrt21_14[0]),.dout(n13359),.clk(gclk));
	jnot g13114(.din(w_n12975_0[1]),.dout(n13360),.clk(gclk));
	jand g13115(.dina(n13360),.dinb(n13359),.dout(n13361),.clk(gclk));
	jor g13116(.dina(n13361),.dinb(n13349),.dout(n13362),.clk(gclk));
	jor g13117(.dina(n13362),.dinb(w_asqrt22_20[2]),.dout(n13363),.clk(gclk));
	jand g13118(.dina(w_n12982_0[1]),.dinb(n13363),.dout(n13364),.clk(gclk));
	jor g13119(.dina(n13364),.dinb(n13348),.dout(n13365),.clk(gclk));
	jor g13120(.dina(n13365),.dinb(w_asqrt23_14[2]),.dout(n13366),.clk(gclk));
	jnot g13121(.din(w_n12990_0[1]),.dout(n13367),.clk(gclk));
	jand g13122(.dina(n13367),.dinb(n13366),.dout(n13368),.clk(gclk));
	jor g13123(.dina(n13368),.dinb(n13347),.dout(n13369),.clk(gclk));
	jor g13124(.dina(n13369),.dinb(w_asqrt24_20[2]),.dout(n13370),.clk(gclk));
	jand g13125(.dina(w_n12997_0[1]),.dinb(n13370),.dout(n13371),.clk(gclk));
	jor g13126(.dina(n13371),.dinb(n13346),.dout(n13372),.clk(gclk));
	jor g13127(.dina(n13372),.dinb(w_asqrt25_14[2]),.dout(n13373),.clk(gclk));
	jnot g13128(.din(w_n13005_0[1]),.dout(n13374),.clk(gclk));
	jand g13129(.dina(n13374),.dinb(n13373),.dout(n13375),.clk(gclk));
	jor g13130(.dina(n13375),.dinb(n13345),.dout(n13376),.clk(gclk));
	jor g13131(.dina(n13376),.dinb(w_asqrt26_20[2]),.dout(n13377),.clk(gclk));
	jand g13132(.dina(w_n13012_0[1]),.dinb(n13377),.dout(n13378),.clk(gclk));
	jor g13133(.dina(n13378),.dinb(n13344),.dout(n13379),.clk(gclk));
	jor g13134(.dina(n13379),.dinb(w_asqrt27_15[1]),.dout(n13380),.clk(gclk));
	jnot g13135(.din(w_n13020_0[1]),.dout(n13381),.clk(gclk));
	jand g13136(.dina(n13381),.dinb(n13380),.dout(n13382),.clk(gclk));
	jor g13137(.dina(n13382),.dinb(n13343),.dout(n13383),.clk(gclk));
	jor g13138(.dina(n13383),.dinb(w_asqrt28_21[0]),.dout(n13384),.clk(gclk));
	jand g13139(.dina(w_n13027_0[1]),.dinb(n13384),.dout(n13385),.clk(gclk));
	jor g13140(.dina(n13385),.dinb(n13342),.dout(n13386),.clk(gclk));
	jor g13141(.dina(n13386),.dinb(w_asqrt29_15[2]),.dout(n13387),.clk(gclk));
	jnot g13142(.din(w_n13035_0[1]),.dout(n13388),.clk(gclk));
	jand g13143(.dina(n13388),.dinb(n13387),.dout(n13389),.clk(gclk));
	jor g13144(.dina(n13389),.dinb(n13341),.dout(n13390),.clk(gclk));
	jor g13145(.dina(n13390),.dinb(w_asqrt30_21[1]),.dout(n13391),.clk(gclk));
	jnot g13146(.din(w_n13042_0[1]),.dout(n13392),.clk(gclk));
	jand g13147(.dina(n13392),.dinb(n13391),.dout(n13393),.clk(gclk));
	jor g13148(.dina(n13393),.dinb(n13340),.dout(n13394),.clk(gclk));
	jor g13149(.dina(n13394),.dinb(w_asqrt31_16[1]),.dout(n13395),.clk(gclk));
	jnot g13150(.din(w_n13049_0[1]),.dout(n13396),.clk(gclk));
	jand g13151(.dina(n13396),.dinb(n13395),.dout(n13397),.clk(gclk));
	jor g13152(.dina(n13397),.dinb(n13339),.dout(n13398),.clk(gclk));
	jor g13153(.dina(n13398),.dinb(w_asqrt32_21[1]),.dout(n13399),.clk(gclk));
	jand g13154(.dina(w_n13056_0[1]),.dinb(n13399),.dout(n13400),.clk(gclk));
	jor g13155(.dina(n13400),.dinb(n13338),.dout(n13401),.clk(gclk));
	jor g13156(.dina(n13401),.dinb(w_asqrt33_17[0]),.dout(n13402),.clk(gclk));
	jnot g13157(.din(w_n13064_0[1]),.dout(n13403),.clk(gclk));
	jand g13158(.dina(n13403),.dinb(n13402),.dout(n13404),.clk(gclk));
	jor g13159(.dina(n13404),.dinb(n13337),.dout(n13405),.clk(gclk));
	jor g13160(.dina(n13405),.dinb(w_asqrt34_21[2]),.dout(n13406),.clk(gclk));
	jand g13161(.dina(w_n13071_0[1]),.dinb(n13406),.dout(n13407),.clk(gclk));
	jor g13162(.dina(n13407),.dinb(n13336),.dout(n13408),.clk(gclk));
	jor g13163(.dina(n13408),.dinb(w_asqrt35_17[2]),.dout(n13409),.clk(gclk));
	jnot g13164(.din(w_n13079_0[1]),.dout(n13410),.clk(gclk));
	jand g13165(.dina(n13410),.dinb(n13409),.dout(n13411),.clk(gclk));
	jor g13166(.dina(n13411),.dinb(n13335),.dout(n13412),.clk(gclk));
	jor g13167(.dina(n13412),.dinb(w_asqrt36_21[2]),.dout(n13413),.clk(gclk));
	jnot g13168(.din(w_n13086_0[1]),.dout(n13414),.clk(gclk));
	jand g13169(.dina(n13414),.dinb(n13413),.dout(n13415),.clk(gclk));
	jor g13170(.dina(n13415),.dinb(n13334),.dout(n13416),.clk(gclk));
	jor g13171(.dina(n13416),.dinb(w_asqrt37_18[0]),.dout(n13417),.clk(gclk));
	jnot g13172(.din(w_n13093_0[1]),.dout(n13418),.clk(gclk));
	jand g13173(.dina(n13418),.dinb(n13417),.dout(n13419),.clk(gclk));
	jor g13174(.dina(n13419),.dinb(n13333),.dout(n13420),.clk(gclk));
	jor g13175(.dina(n13420),.dinb(w_asqrt38_22[0]),.dout(n13421),.clk(gclk));
	jand g13176(.dina(w_n13100_0[1]),.dinb(n13421),.dout(n13422),.clk(gclk));
	jor g13177(.dina(n13422),.dinb(n13332),.dout(n13423),.clk(gclk));
	jor g13178(.dina(n13423),.dinb(w_asqrt39_18[2]),.dout(n13424),.clk(gclk));
	jnot g13179(.din(w_n13108_0[1]),.dout(n13425),.clk(gclk));
	jand g13180(.dina(n13425),.dinb(n13424),.dout(n13426),.clk(gclk));
	jor g13181(.dina(n13426),.dinb(n13331),.dout(n13427),.clk(gclk));
	jor g13182(.dina(n13427),.dinb(w_asqrt40_22[0]),.dout(n13428),.clk(gclk));
	jnot g13183(.din(w_n13115_0[1]),.dout(n13429),.clk(gclk));
	jand g13184(.dina(n13429),.dinb(n13428),.dout(n13430),.clk(gclk));
	jor g13185(.dina(n13430),.dinb(n13330),.dout(n13431),.clk(gclk));
	jor g13186(.dina(n13431),.dinb(w_asqrt41_19[0]),.dout(n13432),.clk(gclk));
	jnot g13187(.din(w_n13122_0[1]),.dout(n13433),.clk(gclk));
	jand g13188(.dina(n13433),.dinb(n13432),.dout(n13434),.clk(gclk));
	jor g13189(.dina(n13434),.dinb(n13329),.dout(n13435),.clk(gclk));
	jor g13190(.dina(n13435),.dinb(w_asqrt42_22[1]),.dout(n13436),.clk(gclk));
	jnot g13191(.din(w_n13129_0[1]),.dout(n13437),.clk(gclk));
	jand g13192(.dina(n13437),.dinb(n13436),.dout(n13438),.clk(gclk));
	jor g13193(.dina(n13438),.dinb(n13328),.dout(n13439),.clk(gclk));
	jor g13194(.dina(n13439),.dinb(w_asqrt43_19[1]),.dout(n13440),.clk(gclk));
	jand g13195(.dina(w_n13136_0[1]),.dinb(n13440),.dout(n13441),.clk(gclk));
	jor g13196(.dina(n13441),.dinb(n13327),.dout(n13442),.clk(gclk));
	jor g13197(.dina(n13442),.dinb(w_asqrt44_22[1]),.dout(n13443),.clk(gclk));
	jand g13198(.dina(n13443),.dinb(w_n13143_0[1]),.dout(n13444),.clk(gclk));
	jor g13199(.dina(n13444),.dinb(n13326),.dout(n13445),.clk(gclk));
	jor g13200(.dina(n13445),.dinb(w_asqrt45_20[0]),.dout(n13446),.clk(gclk));
	jnot g13201(.din(w_n13152_0[1]),.dout(n13447),.clk(gclk));
	jand g13202(.dina(n13447),.dinb(n13446),.dout(n13448),.clk(gclk));
	jor g13203(.dina(n13448),.dinb(n13325),.dout(n13449),.clk(gclk));
	jor g13204(.dina(n13449),.dinb(w_asqrt46_22[1]),.dout(n13450),.clk(gclk));
	jand g13205(.dina(w_n13159_0[1]),.dinb(n13450),.dout(n13451),.clk(gclk));
	jor g13206(.dina(n13451),.dinb(n13324),.dout(n13452),.clk(gclk));
	jor g13207(.dina(n13452),.dinb(w_asqrt47_20[2]),.dout(n13453),.clk(gclk));
	jnot g13208(.din(w_n13167_0[1]),.dout(n13454),.clk(gclk));
	jand g13209(.dina(n13454),.dinb(n13453),.dout(n13455),.clk(gclk));
	jor g13210(.dina(n13455),.dinb(n13323),.dout(n13456),.clk(gclk));
	jor g13211(.dina(n13456),.dinb(w_asqrt48_22[2]),.dout(n13457),.clk(gclk));
	jand g13212(.dina(w_n13174_0[1]),.dinb(n13457),.dout(n13458),.clk(gclk));
	jor g13213(.dina(n13458),.dinb(n13322),.dout(n13459),.clk(gclk));
	jor g13214(.dina(n13459),.dinb(w_asqrt49_21[0]),.dout(n13460),.clk(gclk));
	jnot g13215(.din(w_n13182_0[1]),.dout(n13461),.clk(gclk));
	jand g13216(.dina(n13461),.dinb(n13460),.dout(n13462),.clk(gclk));
	jor g13217(.dina(n13462),.dinb(n13321),.dout(n13463),.clk(gclk));
	jor g13218(.dina(n13463),.dinb(w_asqrt50_23[0]),.dout(n13464),.clk(gclk));
	jnot g13219(.din(w_n13189_0[1]),.dout(n13465),.clk(gclk));
	jand g13220(.dina(n13465),.dinb(n13464),.dout(n13466),.clk(gclk));
	jor g13221(.dina(n13466),.dinb(n13320),.dout(n13467),.clk(gclk));
	jor g13222(.dina(n13467),.dinb(w_asqrt51_21[1]),.dout(n13468),.clk(gclk));
	jnot g13223(.din(w_n13196_0[1]),.dout(n13469),.clk(gclk));
	jand g13224(.dina(n13469),.dinb(n13468),.dout(n13470),.clk(gclk));
	jor g13225(.dina(n13470),.dinb(n13319),.dout(n13471),.clk(gclk));
	jor g13226(.dina(n13471),.dinb(w_asqrt52_23[0]),.dout(n13472),.clk(gclk));
	jand g13227(.dina(w_n13203_0[1]),.dinb(n13472),.dout(n13473),.clk(gclk));
	jor g13228(.dina(n13473),.dinb(n13318),.dout(n13474),.clk(gclk));
	jor g13229(.dina(n13474),.dinb(w_asqrt53_22[0]),.dout(n13475),.clk(gclk));
	jnot g13230(.din(w_n13211_0[1]),.dout(n13476),.clk(gclk));
	jand g13231(.dina(n13476),.dinb(n13475),.dout(n13477),.clk(gclk));
	jor g13232(.dina(n13477),.dinb(n13317),.dout(n13478),.clk(gclk));
	jor g13233(.dina(n13478),.dinb(w_asqrt54_23[0]),.dout(n13479),.clk(gclk));
	jand g13234(.dina(w_n13218_0[1]),.dinb(n13479),.dout(n13480),.clk(gclk));
	jor g13235(.dina(n13480),.dinb(n13316),.dout(n13481),.clk(gclk));
	jor g13236(.dina(n13481),.dinb(w_asqrt55_22[1]),.dout(n13482),.clk(gclk));
	jnot g13237(.din(w_n13226_0[1]),.dout(n13483),.clk(gclk));
	jand g13238(.dina(n13483),.dinb(n13482),.dout(n13484),.clk(gclk));
	jor g13239(.dina(n13484),.dinb(n13315),.dout(n13485),.clk(gclk));
	jor g13240(.dina(n13485),.dinb(w_asqrt56_23[1]),.dout(n13486),.clk(gclk));
	jand g13241(.dina(w_n13233_0[1]),.dinb(n13486),.dout(n13487),.clk(gclk));
	jor g13242(.dina(n13487),.dinb(n13314),.dout(n13488),.clk(gclk));
	jor g13243(.dina(n13488),.dinb(w_asqrt57_23[0]),.dout(n13489),.clk(gclk));
	jnot g13244(.din(w_n13241_0[1]),.dout(n13490),.clk(gclk));
	jand g13245(.dina(n13490),.dinb(n13489),.dout(n13491),.clk(gclk));
	jor g13246(.dina(n13491),.dinb(n13313),.dout(n13492),.clk(gclk));
	jor g13247(.dina(n13492),.dinb(w_asqrt58_23[2]),.dout(n13493),.clk(gclk));
	jand g13248(.dina(w_n13248_0[1]),.dinb(n13493),.dout(n13494),.clk(gclk));
	jor g13249(.dina(n13494),.dinb(n13312),.dout(n13495),.clk(gclk));
	jor g13250(.dina(n13495),.dinb(w_asqrt59_23[1]),.dout(n13496),.clk(gclk));
	jand g13251(.dina(w_n13256_0[1]),.dinb(n13496),.dout(n13497),.clk(gclk));
	jor g13252(.dina(n13497),.dinb(n13311),.dout(n13498),.clk(gclk));
	jor g13253(.dina(n13498),.dinb(w_asqrt60_23[2]),.dout(n13499),.clk(gclk));
	jand g13254(.dina(w_n13264_0[1]),.dinb(n13499),.dout(n13500),.clk(gclk));
	jor g13255(.dina(n13500),.dinb(n13310),.dout(n13501),.clk(gclk));
	jor g13256(.dina(n13501),.dinb(w_asqrt61_23[2]),.dout(n13502),.clk(gclk));
	jnot g13257(.din(w_n13272_0[1]),.dout(n13503),.clk(gclk));
	jand g13258(.dina(n13503),.dinb(n13502),.dout(n13504),.clk(gclk));
	jor g13259(.dina(n13504),.dinb(n13309),.dout(n13505),.clk(gclk));
	jor g13260(.dina(n13505),.dinb(w_asqrt62_23[2]),.dout(n13506),.clk(gclk));
	jnot g13261(.din(w_n13279_0[1]),.dout(n13507),.clk(gclk));
	jand g13262(.dina(n13507),.dinb(n13506),.dout(n13508),.clk(gclk));
	jor g13263(.dina(n13508),.dinb(n13308),.dout(n13509),.clk(gclk));
	jand g13264(.dina(n13509),.dinb(w_n12950_0[0]),.dout(n13510),.clk(gclk));
	jand g13265(.dina(w_n13510_0[1]),.dinb(w_n12731_0[1]),.dout(n13511),.clk(gclk));
	jand g13266(.dina(n13511),.dinb(n13307),.dout(n13512),.clk(gclk));
	jor g13267(.dina(n13512),.dinb(w_asqrt63_29[2]),.dout(n13513),.clk(gclk));
	jnot g13268(.din(w_n13294_0[0]),.dout(n13514),.clk(gclk));
	jand g13269(.dina(n13514),.dinb(n13513),.dout(n13515),.clk(gclk));
	jor g13270(.dina(w_n13515_23[1]),.dinb(n13306),.dout(n13516),.clk(gclk));
	jand g13271(.dina(w_n13516_0[1]),.dinb(n13305),.dout(n13517),.clk(gclk));
	jand g13272(.dina(n13517),.dinb(n13303),.dout(n13518),.clk(gclk));
	jor g13273(.dina(n13518),.dinb(w_n13302_0[1]),.dout(n13519),.clk(gclk));
	jand g13274(.dina(w_n13519_0[2]),.dinb(w_asqrt20_20[0]),.dout(n13520),.clk(gclk));
	jor g13275(.dina(w_n13519_0[1]),.dinb(w_asqrt20_19[2]),.dout(n13521),.clk(gclk));
	jor g13276(.dina(w_n13292_0[0]),.dinb(w_n13287_1[0]),.dout(n13522),.clk(gclk));
	jor g13277(.dina(n13522),.dinb(w_n13285_0[0]),.dout(n13523),.clk(gclk));
	jor g13278(.dina(n13523),.dinb(w_n12947_29[1]),.dout(n13524),.clk(gclk));
	jand g13279(.dina(n13524),.dinb(w_n13516_0[0]),.dout(n13525),.clk(gclk));
	jxor g13280(.dina(n13525),.dinb(w_n12196_0[1]),.dout(n13526),.clk(gclk));
	jnot g13281(.din(w_n13526_0[1]),.dout(n13527),.clk(gclk));
	jand g13282(.dina(w_n13527_0[1]),.dinb(n13521),.dout(n13528),.clk(gclk));
	jor g13283(.dina(n13528),.dinb(w_n13520_0[1]),.dout(n13529),.clk(gclk));
	jand g13284(.dina(w_n13529_0[2]),.dinb(w_asqrt21_13[2]),.dout(n13530),.clk(gclk));
	jor g13285(.dina(w_n13529_0[1]),.dinb(w_asqrt21_13[1]),.dout(n13531),.clk(gclk));
	jxor g13286(.dina(w_n12958_0[0]),.dinb(w_n12410_23[0]),.dout(n13532),.clk(gclk));
	jand g13287(.dina(n13532),.dinb(w_asqrt18_34[1]),.dout(n13533),.clk(gclk));
	jxor g13288(.dina(n13533),.dinb(w_n12964_0[0]),.dout(n13534),.clk(gclk));
	jnot g13289(.din(w_n13534_0[1]),.dout(n13535),.clk(gclk));
	jand g13290(.dina(w_n13535_0[1]),.dinb(n13531),.dout(n13536),.clk(gclk));
	jor g13291(.dina(n13536),.dinb(w_n13530_0[1]),.dout(n13537),.clk(gclk));
	jand g13292(.dina(w_n13537_0[2]),.dinb(w_asqrt22_20[1]),.dout(n13538),.clk(gclk));
	jor g13293(.dina(w_n13537_0[1]),.dinb(w_asqrt22_20[0]),.dout(n13539),.clk(gclk));
	jxor g13294(.dina(w_n12966_0[0]),.dinb(w_n11858_29[2]),.dout(n13540),.clk(gclk));
	jand g13295(.dina(n13540),.dinb(w_asqrt18_34[0]),.dout(n13541),.clk(gclk));
	jxor g13296(.dina(n13541),.dinb(w_n12975_0[0]),.dout(n13542),.clk(gclk));
	jnot g13297(.din(w_n13542_0[1]),.dout(n13543),.clk(gclk));
	jand g13298(.dina(w_n13543_0[1]),.dinb(n13539),.dout(n13544),.clk(gclk));
	jor g13299(.dina(n13544),.dinb(w_n13538_0[1]),.dout(n13545),.clk(gclk));
	jand g13300(.dina(w_n13545_0[2]),.dinb(w_asqrt23_14[1]),.dout(n13546),.clk(gclk));
	jor g13301(.dina(w_n13545_0[1]),.dinb(w_asqrt23_14[0]),.dout(n13547),.clk(gclk));
	jxor g13302(.dina(w_n12977_0[0]),.dinb(w_n11347_23[2]),.dout(n13548),.clk(gclk));
	jand g13303(.dina(n13548),.dinb(w_asqrt18_33[2]),.dout(n13549),.clk(gclk));
	jxor g13304(.dina(n13549),.dinb(w_n12982_0[0]),.dout(n13550),.clk(gclk));
	jand g13305(.dina(w_n13550_0[1]),.dinb(n13547),.dout(n13551),.clk(gclk));
	jor g13306(.dina(n13551),.dinb(w_n13546_0[1]),.dout(n13552),.clk(gclk));
	jand g13307(.dina(w_n13552_0[2]),.dinb(w_asqrt24_20[1]),.dout(n13553),.clk(gclk));
	jor g13308(.dina(w_n13552_0[1]),.dinb(w_asqrt24_20[0]),.dout(n13554),.clk(gclk));
	jxor g13309(.dina(w_n12985_0[0]),.dinb(w_n10824_30[1]),.dout(n13555),.clk(gclk));
	jand g13310(.dina(n13555),.dinb(w_asqrt18_33[1]),.dout(n13556),.clk(gclk));
	jxor g13311(.dina(n13556),.dinb(w_n12990_0[0]),.dout(n13557),.clk(gclk));
	jnot g13312(.din(w_n13557_0[1]),.dout(n13558),.clk(gclk));
	jand g13313(.dina(w_n13558_0[1]),.dinb(n13554),.dout(n13559),.clk(gclk));
	jor g13314(.dina(n13559),.dinb(w_n13553_0[1]),.dout(n13560),.clk(gclk));
	jand g13315(.dina(w_n13560_0[2]),.dinb(w_asqrt25_14[1]),.dout(n13561),.clk(gclk));
	jor g13316(.dina(w_n13560_0[1]),.dinb(w_asqrt25_14[0]),.dout(n13562),.clk(gclk));
	jxor g13317(.dina(w_n12992_0[0]),.dinb(w_n10328_24[2]),.dout(n13563),.clk(gclk));
	jand g13318(.dina(n13563),.dinb(w_asqrt18_33[0]),.dout(n13564),.clk(gclk));
	jxor g13319(.dina(n13564),.dinb(w_n12997_0[0]),.dout(n13565),.clk(gclk));
	jand g13320(.dina(w_n13565_0[1]),.dinb(n13562),.dout(n13566),.clk(gclk));
	jor g13321(.dina(n13566),.dinb(w_n13561_0[1]),.dout(n13567),.clk(gclk));
	jand g13322(.dina(w_n13567_0[2]),.dinb(w_asqrt26_20[1]),.dout(n13568),.clk(gclk));
	jor g13323(.dina(w_n13567_0[1]),.dinb(w_asqrt26_20[0]),.dout(n13569),.clk(gclk));
	jxor g13324(.dina(w_n13000_0[0]),.dinb(w_n9832_31[0]),.dout(n13570),.clk(gclk));
	jand g13325(.dina(n13570),.dinb(w_asqrt18_32[2]),.dout(n13571),.clk(gclk));
	jxor g13326(.dina(n13571),.dinb(w_n13005_0[0]),.dout(n13572),.clk(gclk));
	jnot g13327(.din(w_n13572_0[1]),.dout(n13573),.clk(gclk));
	jand g13328(.dina(w_n13573_0[1]),.dinb(n13569),.dout(n13574),.clk(gclk));
	jor g13329(.dina(n13574),.dinb(w_n13568_0[1]),.dout(n13575),.clk(gclk));
	jand g13330(.dina(w_n13575_0[2]),.dinb(w_asqrt27_15[0]),.dout(n13576),.clk(gclk));
	jor g13331(.dina(w_n13575_0[1]),.dinb(w_asqrt27_14[2]),.dout(n13577),.clk(gclk));
	jxor g13332(.dina(w_n13007_0[0]),.dinb(w_n9369_25[2]),.dout(n13578),.clk(gclk));
	jand g13333(.dina(n13578),.dinb(w_asqrt18_32[1]),.dout(n13579),.clk(gclk));
	jxor g13334(.dina(n13579),.dinb(w_n13012_0[0]),.dout(n13580),.clk(gclk));
	jand g13335(.dina(w_n13580_0[1]),.dinb(n13577),.dout(n13581),.clk(gclk));
	jor g13336(.dina(n13581),.dinb(w_n13576_0[1]),.dout(n13582),.clk(gclk));
	jand g13337(.dina(w_n13582_0[2]),.dinb(w_asqrt28_20[2]),.dout(n13583),.clk(gclk));
	jor g13338(.dina(w_n13582_0[1]),.dinb(w_asqrt28_20[1]),.dout(n13584),.clk(gclk));
	jxor g13339(.dina(w_n13015_0[0]),.dinb(w_n8890_31[1]),.dout(n13585),.clk(gclk));
	jand g13340(.dina(n13585),.dinb(w_asqrt18_32[0]),.dout(n13586),.clk(gclk));
	jxor g13341(.dina(n13586),.dinb(w_n13020_0[0]),.dout(n13587),.clk(gclk));
	jnot g13342(.din(w_n13587_0[1]),.dout(n13588),.clk(gclk));
	jand g13343(.dina(w_n13588_0[1]),.dinb(n13584),.dout(n13589),.clk(gclk));
	jor g13344(.dina(n13589),.dinb(w_n13583_0[1]),.dout(n13590),.clk(gclk));
	jand g13345(.dina(w_n13590_0[2]),.dinb(w_asqrt29_15[1]),.dout(n13591),.clk(gclk));
	jor g13346(.dina(w_n13590_0[1]),.dinb(w_asqrt29_15[0]),.dout(n13592),.clk(gclk));
	jxor g13347(.dina(w_n13022_0[0]),.dinb(w_n8449_26[1]),.dout(n13593),.clk(gclk));
	jand g13348(.dina(n13593),.dinb(w_asqrt18_31[2]),.dout(n13594),.clk(gclk));
	jxor g13349(.dina(n13594),.dinb(w_n13027_0[0]),.dout(n13595),.clk(gclk));
	jand g13350(.dina(w_n13595_0[1]),.dinb(n13592),.dout(n13596),.clk(gclk));
	jor g13351(.dina(n13596),.dinb(w_n13591_0[1]),.dout(n13597),.clk(gclk));
	jand g13352(.dina(w_n13597_0[2]),.dinb(w_asqrt30_21[0]),.dout(n13598),.clk(gclk));
	jor g13353(.dina(w_n13597_0[1]),.dinb(w_asqrt30_20[2]),.dout(n13599),.clk(gclk));
	jxor g13354(.dina(w_n13030_0[0]),.dinb(w_n8003_32[0]),.dout(n13600),.clk(gclk));
	jand g13355(.dina(n13600),.dinb(w_asqrt18_31[1]),.dout(n13601),.clk(gclk));
	jxor g13356(.dina(n13601),.dinb(w_n13035_0[0]),.dout(n13602),.clk(gclk));
	jnot g13357(.din(w_n13602_0[1]),.dout(n13603),.clk(gclk));
	jand g13358(.dina(w_n13603_0[1]),.dinb(n13599),.dout(n13604),.clk(gclk));
	jor g13359(.dina(n13604),.dinb(w_n13598_0[1]),.dout(n13605),.clk(gclk));
	jand g13360(.dina(w_n13605_0[2]),.dinb(w_asqrt31_16[0]),.dout(n13606),.clk(gclk));
	jor g13361(.dina(w_n13605_0[1]),.dinb(w_asqrt31_15[2]),.dout(n13607),.clk(gclk));
	jxor g13362(.dina(w_n13037_0[0]),.dinb(w_n7581_27[1]),.dout(n13608),.clk(gclk));
	jand g13363(.dina(n13608),.dinb(w_asqrt18_31[0]),.dout(n13609),.clk(gclk));
	jxor g13364(.dina(n13609),.dinb(w_n13042_0[0]),.dout(n13610),.clk(gclk));
	jnot g13365(.din(w_n13610_0[1]),.dout(n13611),.clk(gclk));
	jand g13366(.dina(w_n13611_0[1]),.dinb(n13607),.dout(n13612),.clk(gclk));
	jor g13367(.dina(n13612),.dinb(w_n13606_0[1]),.dout(n13613),.clk(gclk));
	jand g13368(.dina(w_n13613_0[2]),.dinb(w_asqrt32_21[0]),.dout(n13614),.clk(gclk));
	jor g13369(.dina(w_n13613_0[1]),.dinb(w_asqrt32_20[2]),.dout(n13615),.clk(gclk));
	jxor g13370(.dina(w_n13044_0[0]),.dinb(w_n7154_32[1]),.dout(n13616),.clk(gclk));
	jand g13371(.dina(n13616),.dinb(w_asqrt18_30[2]),.dout(n13617),.clk(gclk));
	jxor g13372(.dina(n13617),.dinb(w_n13049_0[0]),.dout(n13618),.clk(gclk));
	jnot g13373(.din(w_n13618_0[1]),.dout(n13619),.clk(gclk));
	jand g13374(.dina(w_n13619_0[1]),.dinb(n13615),.dout(n13620),.clk(gclk));
	jor g13375(.dina(n13620),.dinb(w_n13614_0[1]),.dout(n13621),.clk(gclk));
	jand g13376(.dina(w_n13621_0[2]),.dinb(w_asqrt33_16[2]),.dout(n13622),.clk(gclk));
	jor g13377(.dina(w_n13621_0[1]),.dinb(w_asqrt33_16[1]),.dout(n13623),.clk(gclk));
	jxor g13378(.dina(w_n13051_0[0]),.dinb(w_n6758_28[0]),.dout(n13624),.clk(gclk));
	jand g13379(.dina(n13624),.dinb(w_asqrt18_30[1]),.dout(n13625),.clk(gclk));
	jxor g13380(.dina(n13625),.dinb(w_n13056_0[0]),.dout(n13626),.clk(gclk));
	jand g13381(.dina(w_n13626_0[1]),.dinb(n13623),.dout(n13627),.clk(gclk));
	jor g13382(.dina(n13627),.dinb(w_n13622_0[1]),.dout(n13628),.clk(gclk));
	jand g13383(.dina(w_n13628_0[2]),.dinb(w_asqrt34_21[1]),.dout(n13629),.clk(gclk));
	jor g13384(.dina(w_n13628_0[1]),.dinb(w_asqrt34_21[0]),.dout(n13630),.clk(gclk));
	jxor g13385(.dina(w_n13059_0[0]),.dinb(w_n6357_32[2]),.dout(n13631),.clk(gclk));
	jand g13386(.dina(n13631),.dinb(w_asqrt18_30[0]),.dout(n13632),.clk(gclk));
	jxor g13387(.dina(n13632),.dinb(w_n13064_0[0]),.dout(n13633),.clk(gclk));
	jnot g13388(.din(w_n13633_0[1]),.dout(n13634),.clk(gclk));
	jand g13389(.dina(w_n13634_0[1]),.dinb(n13630),.dout(n13635),.clk(gclk));
	jor g13390(.dina(n13635),.dinb(w_n13629_0[1]),.dout(n13636),.clk(gclk));
	jand g13391(.dina(w_n13636_0[2]),.dinb(w_asqrt35_17[1]),.dout(n13637),.clk(gclk));
	jor g13392(.dina(w_n13636_0[1]),.dinb(w_asqrt35_17[0]),.dout(n13638),.clk(gclk));
	jxor g13393(.dina(w_n13066_0[0]),.dinb(w_n5989_28[2]),.dout(n13639),.clk(gclk));
	jand g13394(.dina(n13639),.dinb(w_asqrt18_29[2]),.dout(n13640),.clk(gclk));
	jxor g13395(.dina(n13640),.dinb(w_n13071_0[0]),.dout(n13641),.clk(gclk));
	jand g13396(.dina(w_n13641_0[1]),.dinb(n13638),.dout(n13642),.clk(gclk));
	jor g13397(.dina(n13642),.dinb(w_n13637_0[1]),.dout(n13643),.clk(gclk));
	jand g13398(.dina(w_n13643_0[2]),.dinb(w_asqrt36_21[1]),.dout(n13644),.clk(gclk));
	jor g13399(.dina(w_n13643_0[1]),.dinb(w_asqrt36_21[0]),.dout(n13645),.clk(gclk));
	jxor g13400(.dina(w_n13074_0[0]),.dinb(w_n5606_33[0]),.dout(n13646),.clk(gclk));
	jand g13401(.dina(n13646),.dinb(w_asqrt18_29[1]),.dout(n13647),.clk(gclk));
	jxor g13402(.dina(n13647),.dinb(w_n13079_0[0]),.dout(n13648),.clk(gclk));
	jnot g13403(.din(w_n13648_0[1]),.dout(n13649),.clk(gclk));
	jand g13404(.dina(w_n13649_0[1]),.dinb(n13645),.dout(n13650),.clk(gclk));
	jor g13405(.dina(n13650),.dinb(w_n13644_0[1]),.dout(n13651),.clk(gclk));
	jand g13406(.dina(w_n13651_0[2]),.dinb(w_asqrt37_17[2]),.dout(n13652),.clk(gclk));
	jor g13407(.dina(w_n13651_0[1]),.dinb(w_asqrt37_17[1]),.dout(n13653),.clk(gclk));
	jxor g13408(.dina(w_n13081_0[0]),.dinb(w_n5259_29[2]),.dout(n13654),.clk(gclk));
	jand g13409(.dina(n13654),.dinb(w_asqrt18_29[0]),.dout(n13655),.clk(gclk));
	jxor g13410(.dina(n13655),.dinb(w_n13086_0[0]),.dout(n13656),.clk(gclk));
	jnot g13411(.din(w_n13656_0[1]),.dout(n13657),.clk(gclk));
	jand g13412(.dina(w_n13657_0[1]),.dinb(n13653),.dout(n13658),.clk(gclk));
	jor g13413(.dina(n13658),.dinb(w_n13652_0[1]),.dout(n13659),.clk(gclk));
	jand g13414(.dina(w_n13659_0[2]),.dinb(w_asqrt38_21[2]),.dout(n13660),.clk(gclk));
	jor g13415(.dina(w_n13659_0[1]),.dinb(w_asqrt38_21[1]),.dout(n13661),.clk(gclk));
	jxor g13416(.dina(w_n13088_0[0]),.dinb(w_n4902_33[2]),.dout(n13662),.clk(gclk));
	jand g13417(.dina(n13662),.dinb(w_asqrt18_28[2]),.dout(n13663),.clk(gclk));
	jxor g13418(.dina(n13663),.dinb(w_n13093_0[0]),.dout(n13664),.clk(gclk));
	jnot g13419(.din(w_n13664_0[1]),.dout(n13665),.clk(gclk));
	jand g13420(.dina(w_n13665_0[1]),.dinb(n13661),.dout(n13666),.clk(gclk));
	jor g13421(.dina(n13666),.dinb(w_n13660_0[1]),.dout(n13667),.clk(gclk));
	jand g13422(.dina(w_n13667_0[2]),.dinb(w_asqrt39_18[1]),.dout(n13668),.clk(gclk));
	jor g13423(.dina(w_n13667_0[1]),.dinb(w_asqrt39_18[0]),.dout(n13669),.clk(gclk));
	jxor g13424(.dina(w_n13095_0[0]),.dinb(w_n4582_30[2]),.dout(n13670),.clk(gclk));
	jand g13425(.dina(n13670),.dinb(w_asqrt18_28[1]),.dout(n13671),.clk(gclk));
	jxor g13426(.dina(n13671),.dinb(w_n13100_0[0]),.dout(n13672),.clk(gclk));
	jand g13427(.dina(w_n13672_0[1]),.dinb(n13669),.dout(n13673),.clk(gclk));
	jor g13428(.dina(n13673),.dinb(w_n13668_0[1]),.dout(n13674),.clk(gclk));
	jand g13429(.dina(w_n13674_0[2]),.dinb(w_asqrt40_21[2]),.dout(n13675),.clk(gclk));
	jor g13430(.dina(w_n13674_0[1]),.dinb(w_asqrt40_21[1]),.dout(n13676),.clk(gclk));
	jxor g13431(.dina(w_n13103_0[0]),.dinb(w_n4249_34[1]),.dout(n13677),.clk(gclk));
	jand g13432(.dina(n13677),.dinb(w_asqrt18_28[0]),.dout(n13678),.clk(gclk));
	jxor g13433(.dina(n13678),.dinb(w_n13108_0[0]),.dout(n13679),.clk(gclk));
	jnot g13434(.din(w_n13679_0[1]),.dout(n13680),.clk(gclk));
	jand g13435(.dina(w_n13680_0[1]),.dinb(n13676),.dout(n13681),.clk(gclk));
	jor g13436(.dina(n13681),.dinb(w_n13675_0[1]),.dout(n13682),.clk(gclk));
	jand g13437(.dina(w_n13682_0[2]),.dinb(w_asqrt41_18[2]),.dout(n13683),.clk(gclk));
	jor g13438(.dina(w_n13682_0[1]),.dinb(w_asqrt41_18[1]),.dout(n13684),.clk(gclk));
	jxor g13439(.dina(w_n13110_0[0]),.dinb(w_n3955_31[1]),.dout(n13685),.clk(gclk));
	jand g13440(.dina(n13685),.dinb(w_asqrt18_27[2]),.dout(n13686),.clk(gclk));
	jxor g13441(.dina(n13686),.dinb(w_n13115_0[0]),.dout(n13687),.clk(gclk));
	jnot g13442(.din(w_n13687_0[1]),.dout(n13688),.clk(gclk));
	jand g13443(.dina(w_n13688_0[1]),.dinb(n13684),.dout(n13689),.clk(gclk));
	jor g13444(.dina(n13689),.dinb(w_n13683_0[1]),.dout(n13690),.clk(gclk));
	jand g13445(.dina(w_n13690_0[2]),.dinb(w_asqrt42_22[0]),.dout(n13691),.clk(gclk));
	jor g13446(.dina(w_n13690_0[1]),.dinb(w_asqrt42_21[2]),.dout(n13692),.clk(gclk));
	jxor g13447(.dina(w_n13117_0[0]),.dinb(w_n3642_34[2]),.dout(n13693),.clk(gclk));
	jand g13448(.dina(n13693),.dinb(w_asqrt18_27[1]),.dout(n13694),.clk(gclk));
	jxor g13449(.dina(n13694),.dinb(w_n13122_0[0]),.dout(n13695),.clk(gclk));
	jnot g13450(.din(w_n13695_0[1]),.dout(n13696),.clk(gclk));
	jand g13451(.dina(w_n13696_0[1]),.dinb(n13692),.dout(n13697),.clk(gclk));
	jor g13452(.dina(n13697),.dinb(w_n13691_0[1]),.dout(n13698),.clk(gclk));
	jand g13453(.dina(w_n13698_0[2]),.dinb(w_asqrt43_19[0]),.dout(n13699),.clk(gclk));
	jor g13454(.dina(w_n13698_0[1]),.dinb(w_asqrt43_18[2]),.dout(n13700),.clk(gclk));
	jxor g13455(.dina(w_n13124_0[0]),.dinb(w_n3368_32[0]),.dout(n13701),.clk(gclk));
	jand g13456(.dina(n13701),.dinb(w_asqrt18_27[0]),.dout(n13702),.clk(gclk));
	jxor g13457(.dina(n13702),.dinb(w_n13129_0[0]),.dout(n13703),.clk(gclk));
	jnot g13458(.din(w_n13703_0[1]),.dout(n13704),.clk(gclk));
	jand g13459(.dina(w_n13704_0[1]),.dinb(n13700),.dout(n13705),.clk(gclk));
	jor g13460(.dina(n13705),.dinb(w_n13699_0[1]),.dout(n13706),.clk(gclk));
	jand g13461(.dina(w_n13706_0[2]),.dinb(w_asqrt44_22[0]),.dout(n13707),.clk(gclk));
	jor g13462(.dina(w_n13706_0[1]),.dinb(w_asqrt44_21[2]),.dout(n13708),.clk(gclk));
	jxor g13463(.dina(w_n13131_0[0]),.dinb(w_n3089_35[1]),.dout(n13709),.clk(gclk));
	jand g13464(.dina(n13709),.dinb(w_asqrt18_26[2]),.dout(n13710),.clk(gclk));
	jxor g13465(.dina(n13710),.dinb(w_n13136_0[0]),.dout(n13711),.clk(gclk));
	jand g13466(.dina(w_n13711_0[1]),.dinb(n13708),.dout(n13712),.clk(gclk));
	jor g13467(.dina(n13712),.dinb(w_n13707_0[1]),.dout(n13713),.clk(gclk));
	jand g13468(.dina(w_n13713_0[2]),.dinb(w_asqrt45_19[2]),.dout(n13714),.clk(gclk));
	jxor g13469(.dina(w_n13139_0[0]),.dinb(w_n2833_33[0]),.dout(n13715),.clk(gclk));
	jand g13470(.dina(n13715),.dinb(w_asqrt18_26[1]),.dout(n13716),.clk(gclk));
	jxor g13471(.dina(n13716),.dinb(w_n13143_0[0]),.dout(n13717),.clk(gclk));
	jor g13472(.dina(w_n13713_0[1]),.dinb(w_asqrt45_19[1]),.dout(n13718),.clk(gclk));
	jand g13473(.dina(n13718),.dinb(w_n13717_0[1]),.dout(n13719),.clk(gclk));
	jor g13474(.dina(n13719),.dinb(w_n13714_0[1]),.dout(n13720),.clk(gclk));
	jand g13475(.dina(w_n13720_0[2]),.dinb(w_asqrt46_22[0]),.dout(n13721),.clk(gclk));
	jor g13476(.dina(w_n13720_0[1]),.dinb(w_asqrt46_21[2]),.dout(n13722),.clk(gclk));
	jxor g13477(.dina(w_n13147_0[0]),.dinb(w_n2572_35[2]),.dout(n13723),.clk(gclk));
	jand g13478(.dina(n13723),.dinb(w_asqrt18_26[0]),.dout(n13724),.clk(gclk));
	jxor g13479(.dina(n13724),.dinb(w_n13152_0[0]),.dout(n13725),.clk(gclk));
	jnot g13480(.din(w_n13725_0[1]),.dout(n13726),.clk(gclk));
	jand g13481(.dina(w_n13726_0[1]),.dinb(n13722),.dout(n13727),.clk(gclk));
	jor g13482(.dina(n13727),.dinb(w_n13721_0[1]),.dout(n13728),.clk(gclk));
	jand g13483(.dina(w_n13728_0[2]),.dinb(w_asqrt47_20[1]),.dout(n13729),.clk(gclk));
	jor g13484(.dina(w_n13728_0[1]),.dinb(w_asqrt47_20[0]),.dout(n13730),.clk(gclk));
	jxor g13485(.dina(w_n13154_0[0]),.dinb(w_n2345_33[2]),.dout(n13731),.clk(gclk));
	jand g13486(.dina(n13731),.dinb(w_asqrt18_25[2]),.dout(n13732),.clk(gclk));
	jxor g13487(.dina(n13732),.dinb(w_n13159_0[0]),.dout(n13733),.clk(gclk));
	jand g13488(.dina(w_n13733_0[1]),.dinb(n13730),.dout(n13734),.clk(gclk));
	jor g13489(.dina(n13734),.dinb(w_n13729_0[1]),.dout(n13735),.clk(gclk));
	jand g13490(.dina(w_n13735_0[2]),.dinb(w_asqrt48_22[1]),.dout(n13736),.clk(gclk));
	jor g13491(.dina(w_n13735_0[1]),.dinb(w_asqrt48_22[0]),.dout(n13737),.clk(gclk));
	jxor g13492(.dina(w_n13162_0[0]),.dinb(w_n2108_36[1]),.dout(n13738),.clk(gclk));
	jand g13493(.dina(n13738),.dinb(w_asqrt18_25[1]),.dout(n13739),.clk(gclk));
	jxor g13494(.dina(n13739),.dinb(w_n13167_0[0]),.dout(n13740),.clk(gclk));
	jnot g13495(.din(w_n13740_0[1]),.dout(n13741),.clk(gclk));
	jand g13496(.dina(w_n13741_0[1]),.dinb(n13737),.dout(n13742),.clk(gclk));
	jor g13497(.dina(n13742),.dinb(w_n13736_0[1]),.dout(n13743),.clk(gclk));
	jand g13498(.dina(w_n13743_0[2]),.dinb(w_asqrt49_20[2]),.dout(n13744),.clk(gclk));
	jor g13499(.dina(w_n13743_0[1]),.dinb(w_asqrt49_20[1]),.dout(n13745),.clk(gclk));
	jxor g13500(.dina(w_n13169_0[0]),.dinb(w_n1912_34[2]),.dout(n13746),.clk(gclk));
	jand g13501(.dina(n13746),.dinb(w_asqrt18_25[0]),.dout(n13747),.clk(gclk));
	jxor g13502(.dina(n13747),.dinb(w_n13174_0[0]),.dout(n13748),.clk(gclk));
	jand g13503(.dina(w_n13748_0[1]),.dinb(n13745),.dout(n13749),.clk(gclk));
	jor g13504(.dina(n13749),.dinb(w_n13744_0[1]),.dout(n13750),.clk(gclk));
	jand g13505(.dina(w_n13750_0[2]),.dinb(w_asqrt50_22[2]),.dout(n13751),.clk(gclk));
	jor g13506(.dina(w_n13750_0[1]),.dinb(w_asqrt50_22[1]),.dout(n13752),.clk(gclk));
	jxor g13507(.dina(w_n13177_0[0]),.dinb(w_n1699_37[0]),.dout(n13753),.clk(gclk));
	jand g13508(.dina(n13753),.dinb(w_asqrt18_24[2]),.dout(n13754),.clk(gclk));
	jxor g13509(.dina(n13754),.dinb(w_n13182_0[0]),.dout(n13755),.clk(gclk));
	jnot g13510(.din(w_n13755_0[1]),.dout(n13756),.clk(gclk));
	jand g13511(.dina(w_n13756_0[1]),.dinb(n13752),.dout(n13757),.clk(gclk));
	jor g13512(.dina(n13757),.dinb(w_n13751_0[1]),.dout(n13758),.clk(gclk));
	jand g13513(.dina(w_n13758_0[2]),.dinb(w_asqrt51_21[0]),.dout(n13759),.clk(gclk));
	jor g13514(.dina(w_n13758_0[1]),.dinb(w_asqrt51_20[2]),.dout(n13760),.clk(gclk));
	jxor g13515(.dina(w_n13184_0[0]),.dinb(w_n1516_35[1]),.dout(n13761),.clk(gclk));
	jand g13516(.dina(n13761),.dinb(w_asqrt18_24[1]),.dout(n13762),.clk(gclk));
	jxor g13517(.dina(n13762),.dinb(w_n13189_0[0]),.dout(n13763),.clk(gclk));
	jnot g13518(.din(w_n13763_0[1]),.dout(n13764),.clk(gclk));
	jand g13519(.dina(w_n13764_0[1]),.dinb(n13760),.dout(n13765),.clk(gclk));
	jor g13520(.dina(n13765),.dinb(w_n13759_0[1]),.dout(n13766),.clk(gclk));
	jand g13521(.dina(w_n13766_0[2]),.dinb(w_asqrt52_22[2]),.dout(n13767),.clk(gclk));
	jor g13522(.dina(w_n13766_0[1]),.dinb(w_asqrt52_22[1]),.dout(n13768),.clk(gclk));
	jxor g13523(.dina(w_n13191_0[0]),.dinb(w_n1332_37[0]),.dout(n13769),.clk(gclk));
	jand g13524(.dina(n13769),.dinb(w_asqrt18_24[0]),.dout(n13770),.clk(gclk));
	jxor g13525(.dina(n13770),.dinb(w_n13196_0[0]),.dout(n13771),.clk(gclk));
	jnot g13526(.din(w_n13771_0[1]),.dout(n13772),.clk(gclk));
	jand g13527(.dina(w_n13772_0[1]),.dinb(n13768),.dout(n13773),.clk(gclk));
	jor g13528(.dina(n13773),.dinb(w_n13767_0[1]),.dout(n13774),.clk(gclk));
	jand g13529(.dina(w_n13774_0[2]),.dinb(w_asqrt53_21[2]),.dout(n13775),.clk(gclk));
	jor g13530(.dina(w_n13774_0[1]),.dinb(w_asqrt53_21[1]),.dout(n13776),.clk(gclk));
	jxor g13531(.dina(w_n13198_0[0]),.dinb(w_n1173_36[0]),.dout(n13777),.clk(gclk));
	jand g13532(.dina(n13777),.dinb(w_asqrt18_23[2]),.dout(n13778),.clk(gclk));
	jxor g13533(.dina(n13778),.dinb(w_n13203_0[0]),.dout(n13779),.clk(gclk));
	jand g13534(.dina(w_n13779_0[1]),.dinb(n13776),.dout(n13780),.clk(gclk));
	jor g13535(.dina(n13780),.dinb(w_n13775_0[1]),.dout(n13781),.clk(gclk));
	jand g13536(.dina(w_n13781_0[2]),.dinb(w_asqrt54_22[2]),.dout(n13782),.clk(gclk));
	jor g13537(.dina(w_n13781_0[1]),.dinb(w_asqrt54_22[1]),.dout(n13783),.clk(gclk));
	jxor g13538(.dina(w_n13206_0[0]),.dinb(w_n1008_38[0]),.dout(n13784),.clk(gclk));
	jand g13539(.dina(n13784),.dinb(w_asqrt18_23[1]),.dout(n13785),.clk(gclk));
	jxor g13540(.dina(n13785),.dinb(w_n13211_0[0]),.dout(n13786),.clk(gclk));
	jnot g13541(.din(w_n13786_0[1]),.dout(n13787),.clk(gclk));
	jand g13542(.dina(w_n13787_0[1]),.dinb(n13783),.dout(n13788),.clk(gclk));
	jor g13543(.dina(n13788),.dinb(w_n13782_0[1]),.dout(n13789),.clk(gclk));
	jand g13544(.dina(w_n13789_0[2]),.dinb(w_asqrt55_22[0]),.dout(n13790),.clk(gclk));
	jor g13545(.dina(w_n13789_0[1]),.dinb(w_asqrt55_21[2]),.dout(n13791),.clk(gclk));
	jxor g13546(.dina(w_n13213_0[0]),.dinb(w_n884_37[0]),.dout(n13792),.clk(gclk));
	jand g13547(.dina(n13792),.dinb(w_asqrt18_23[0]),.dout(n13793),.clk(gclk));
	jxor g13548(.dina(n13793),.dinb(w_n13218_0[0]),.dout(n13794),.clk(gclk));
	jand g13549(.dina(w_n13794_0[1]),.dinb(n13791),.dout(n13795),.clk(gclk));
	jor g13550(.dina(n13795),.dinb(w_n13790_0[1]),.dout(n13796),.clk(gclk));
	jand g13551(.dina(w_n13796_0[2]),.dinb(w_asqrt56_23[0]),.dout(n13797),.clk(gclk));
	jor g13552(.dina(w_n13796_0[1]),.dinb(w_asqrt56_22[2]),.dout(n13798),.clk(gclk));
	jxor g13553(.dina(w_n13221_0[0]),.dinb(w_n743_38[0]),.dout(n13799),.clk(gclk));
	jand g13554(.dina(n13799),.dinb(w_asqrt18_22[2]),.dout(n13800),.clk(gclk));
	jxor g13555(.dina(n13800),.dinb(w_n13226_0[0]),.dout(n13801),.clk(gclk));
	jnot g13556(.din(w_n13801_0[1]),.dout(n13802),.clk(gclk));
	jand g13557(.dina(w_n13802_0[1]),.dinb(n13798),.dout(n13803),.clk(gclk));
	jor g13558(.dina(n13803),.dinb(w_n13797_0[1]),.dout(n13804),.clk(gclk));
	jand g13559(.dina(w_n13804_0[2]),.dinb(w_asqrt57_22[2]),.dout(n13805),.clk(gclk));
	jor g13560(.dina(w_n13804_0[1]),.dinb(w_asqrt57_22[1]),.dout(n13806),.clk(gclk));
	jxor g13561(.dina(w_n13228_0[0]),.dinb(w_n635_38[0]),.dout(n13807),.clk(gclk));
	jand g13562(.dina(n13807),.dinb(w_asqrt18_22[1]),.dout(n13808),.clk(gclk));
	jxor g13563(.dina(n13808),.dinb(w_n13233_0[0]),.dout(n13809),.clk(gclk));
	jand g13564(.dina(w_n13809_0[1]),.dinb(n13806),.dout(n13810),.clk(gclk));
	jor g13565(.dina(n13810),.dinb(w_n13805_0[1]),.dout(n13811),.clk(gclk));
	jand g13566(.dina(w_n13811_0[2]),.dinb(w_asqrt58_23[1]),.dout(n13812),.clk(gclk));
	jor g13567(.dina(w_n13811_0[1]),.dinb(w_asqrt58_23[0]),.dout(n13813),.clk(gclk));
	jxor g13568(.dina(w_n13236_0[0]),.dinb(w_n515_39[0]),.dout(n13814),.clk(gclk));
	jand g13569(.dina(n13814),.dinb(w_asqrt18_22[0]),.dout(n13815),.clk(gclk));
	jxor g13570(.dina(n13815),.dinb(w_n13241_0[0]),.dout(n13816),.clk(gclk));
	jnot g13571(.din(w_n13816_0[1]),.dout(n13817),.clk(gclk));
	jand g13572(.dina(w_n13817_0[1]),.dinb(n13813),.dout(n13818),.clk(gclk));
	jor g13573(.dina(n13818),.dinb(w_n13812_0[1]),.dout(n13819),.clk(gclk));
	jand g13574(.dina(w_n13819_0[2]),.dinb(w_asqrt59_23[0]),.dout(n13820),.clk(gclk));
	jor g13575(.dina(w_n13819_0[1]),.dinb(w_asqrt59_22[2]),.dout(n13821),.clk(gclk));
	jxor g13576(.dina(w_n13243_0[0]),.dinb(w_n443_39[0]),.dout(n13822),.clk(gclk));
	jand g13577(.dina(n13822),.dinb(w_asqrt18_21[2]),.dout(n13823),.clk(gclk));
	jxor g13578(.dina(n13823),.dinb(w_n13248_0[0]),.dout(n13824),.clk(gclk));
	jand g13579(.dina(w_n13824_0[1]),.dinb(n13821),.dout(n13825),.clk(gclk));
	jor g13580(.dina(n13825),.dinb(w_n13820_0[1]),.dout(n13826),.clk(gclk));
	jand g13581(.dina(w_n13826_0[2]),.dinb(w_asqrt60_23[1]),.dout(n13827),.clk(gclk));
	jor g13582(.dina(w_n13826_0[1]),.dinb(w_asqrt60_23[0]),.dout(n13828),.clk(gclk));
	jxor g13583(.dina(w_n13251_0[0]),.dinb(w_n352_39[1]),.dout(n13829),.clk(gclk));
	jand g13584(.dina(n13829),.dinb(w_asqrt18_21[1]),.dout(n13830),.clk(gclk));
	jxor g13585(.dina(n13830),.dinb(w_n13256_0[0]),.dout(n13831),.clk(gclk));
	jand g13586(.dina(w_n13831_0[1]),.dinb(n13828),.dout(n13832),.clk(gclk));
	jor g13587(.dina(n13832),.dinb(w_n13827_0[1]),.dout(n13833),.clk(gclk));
	jand g13588(.dina(w_n13833_0[2]),.dinb(w_asqrt61_23[1]),.dout(n13834),.clk(gclk));
	jor g13589(.dina(w_n13833_0[1]),.dinb(w_asqrt61_23[0]),.dout(n13835),.clk(gclk));
	jxor g13590(.dina(w_n13259_0[0]),.dinb(w_n294_39[2]),.dout(n13836),.clk(gclk));
	jand g13591(.dina(n13836),.dinb(w_asqrt18_21[0]),.dout(n13837),.clk(gclk));
	jxor g13592(.dina(n13837),.dinb(w_n13264_0[0]),.dout(n13838),.clk(gclk));
	jand g13593(.dina(w_n13838_0[1]),.dinb(n13835),.dout(n13839),.clk(gclk));
	jor g13594(.dina(n13839),.dinb(w_n13834_0[1]),.dout(n13840),.clk(gclk));
	jand g13595(.dina(w_n13840_0[2]),.dinb(w_asqrt62_23[1]),.dout(n13841),.clk(gclk));
	jor g13596(.dina(w_n13840_0[1]),.dinb(w_asqrt62_23[0]),.dout(n13842),.clk(gclk));
	jxor g13597(.dina(w_n13267_0[0]),.dinb(w_n239_39[2]),.dout(n13843),.clk(gclk));
	jand g13598(.dina(n13843),.dinb(w_asqrt18_20[2]),.dout(n13844),.clk(gclk));
	jxor g13599(.dina(n13844),.dinb(w_n13272_0[0]),.dout(n13845),.clk(gclk));
	jnot g13600(.din(w_n13845_0[1]),.dout(n13846),.clk(gclk));
	jand g13601(.dina(w_n13846_0[1]),.dinb(n13842),.dout(n13847),.clk(gclk));
	jor g13602(.dina(n13847),.dinb(w_n13841_0[1]),.dout(n13848),.clk(gclk));
	jxor g13603(.dina(w_n13274_0[0]),.dinb(w_n221_40[0]),.dout(n13849),.clk(gclk));
	jand g13604(.dina(n13849),.dinb(w_asqrt18_20[1]),.dout(n13850),.clk(gclk));
	jxor g13605(.dina(n13850),.dinb(w_n13279_0[0]),.dout(n13851),.clk(gclk));
	jnot g13606(.din(w_n13851_0[1]),.dout(n13852),.clk(gclk));
	jor g13607(.dina(w_n13852_0[2]),.dinb(w_n13848_0[2]),.dout(n13853),.clk(gclk));
	jnot g13608(.din(w_n13853_0[1]),.dout(n13854),.clk(gclk));
	jand g13609(.dina(w_n13515_23[0]),.dinb(w_n13281_0[0]),.dout(n13855),.clk(gclk));
	jnot g13610(.din(n13855),.dout(n13856),.clk(gclk));
	jnot g13611(.din(w_n13287_0[2]),.dout(n13857),.clk(gclk));
	jand g13612(.dina(w_n13282_0[0]),.dinb(w_asqrt63_29[1]),.dout(n13858),.clk(gclk));
	jand g13613(.dina(n13858),.dinb(n13857),.dout(n13859),.clk(gclk));
	jand g13614(.dina(w_n13859_0[1]),.dinb(n13856),.dout(n13860),.clk(gclk));
	jnot g13615(.din(w_n13841_0[0]),.dout(n13861),.clk(gclk));
	jnot g13616(.din(w_n13834_0[0]),.dout(n13862),.clk(gclk));
	jnot g13617(.din(w_n13827_0[0]),.dout(n13863),.clk(gclk));
	jnot g13618(.din(w_n13820_0[0]),.dout(n13864),.clk(gclk));
	jnot g13619(.din(w_n13812_0[0]),.dout(n13865),.clk(gclk));
	jnot g13620(.din(w_n13805_0[0]),.dout(n13866),.clk(gclk));
	jnot g13621(.din(w_n13797_0[0]),.dout(n13867),.clk(gclk));
	jnot g13622(.din(w_n13790_0[0]),.dout(n13868),.clk(gclk));
	jnot g13623(.din(w_n13782_0[0]),.dout(n13869),.clk(gclk));
	jnot g13624(.din(w_n13775_0[0]),.dout(n13870),.clk(gclk));
	jnot g13625(.din(w_n13767_0[0]),.dout(n13871),.clk(gclk));
	jnot g13626(.din(w_n13759_0[0]),.dout(n13872),.clk(gclk));
	jnot g13627(.din(w_n13751_0[0]),.dout(n13873),.clk(gclk));
	jnot g13628(.din(w_n13744_0[0]),.dout(n13874),.clk(gclk));
	jnot g13629(.din(w_n13736_0[0]),.dout(n13875),.clk(gclk));
	jnot g13630(.din(w_n13729_0[0]),.dout(n13876),.clk(gclk));
	jnot g13631(.din(w_n13721_0[0]),.dout(n13877),.clk(gclk));
	jnot g13632(.din(w_n13714_0[0]),.dout(n13878),.clk(gclk));
	jnot g13633(.din(w_n13717_0[0]),.dout(n13879),.clk(gclk));
	jnot g13634(.din(w_n13707_0[0]),.dout(n13880),.clk(gclk));
	jnot g13635(.din(w_n13699_0[0]),.dout(n13881),.clk(gclk));
	jnot g13636(.din(w_n13691_0[0]),.dout(n13882),.clk(gclk));
	jnot g13637(.din(w_n13683_0[0]),.dout(n13883),.clk(gclk));
	jnot g13638(.din(w_n13675_0[0]),.dout(n13884),.clk(gclk));
	jnot g13639(.din(w_n13668_0[0]),.dout(n13885),.clk(gclk));
	jnot g13640(.din(w_n13660_0[0]),.dout(n13886),.clk(gclk));
	jnot g13641(.din(w_n13652_0[0]),.dout(n13887),.clk(gclk));
	jnot g13642(.din(w_n13644_0[0]),.dout(n13888),.clk(gclk));
	jnot g13643(.din(w_n13637_0[0]),.dout(n13889),.clk(gclk));
	jnot g13644(.din(w_n13629_0[0]),.dout(n13890),.clk(gclk));
	jnot g13645(.din(w_n13622_0[0]),.dout(n13891),.clk(gclk));
	jnot g13646(.din(w_n13614_0[0]),.dout(n13892),.clk(gclk));
	jnot g13647(.din(w_n13606_0[0]),.dout(n13893),.clk(gclk));
	jnot g13648(.din(w_n13598_0[0]),.dout(n13894),.clk(gclk));
	jnot g13649(.din(w_n13591_0[0]),.dout(n13895),.clk(gclk));
	jnot g13650(.din(w_n13583_0[0]),.dout(n13896),.clk(gclk));
	jnot g13651(.din(w_n13576_0[0]),.dout(n13897),.clk(gclk));
	jnot g13652(.din(w_n13568_0[0]),.dout(n13898),.clk(gclk));
	jnot g13653(.din(w_n13561_0[0]),.dout(n13899),.clk(gclk));
	jnot g13654(.din(w_n13553_0[0]),.dout(n13900),.clk(gclk));
	jnot g13655(.din(w_n13546_0[0]),.dout(n13901),.clk(gclk));
	jnot g13656(.din(w_n13538_0[0]),.dout(n13902),.clk(gclk));
	jnot g13657(.din(w_n13530_0[0]),.dout(n13903),.clk(gclk));
	jnot g13658(.din(w_n13520_0[0]),.dout(n13904),.clk(gclk));
	jnot g13659(.din(w_n13302_0[0]),.dout(n13905),.clk(gclk));
	jnot g13660(.din(w_n13299_0[0]),.dout(n13906),.clk(gclk));
	jor g13661(.dina(w_n13515_22[2]),.dinb(w_n12953_0[2]),.dout(n13907),.clk(gclk));
	jand g13662(.dina(n13907),.dinb(n13906),.dout(n13908),.clk(gclk));
	jand g13663(.dina(n13908),.dinb(w_n12947_29[0]),.dout(n13909),.clk(gclk));
	jor g13664(.dina(w_n13515_22[1]),.dinb(w_a36_0[0]),.dout(n13910),.clk(gclk));
	jand g13665(.dina(n13910),.dinb(w_a37_0[0]),.dout(n13911),.clk(gclk));
	jand g13666(.dina(w_asqrt18_20[0]),.dinb(w_n12955_0[0]),.dout(n13912),.clk(gclk));
	jor g13667(.dina(n13912),.dinb(n13911),.dout(n13913),.clk(gclk));
	jor g13668(.dina(w_n13913_0[1]),.dinb(n13909),.dout(n13914),.clk(gclk));
	jand g13669(.dina(n13914),.dinb(n13905),.dout(n13915),.clk(gclk));
	jand g13670(.dina(n13915),.dinb(w_n12410_22[2]),.dout(n13916),.clk(gclk));
	jor g13671(.dina(w_n13526_0[0]),.dinb(n13916),.dout(n13917),.clk(gclk));
	jand g13672(.dina(n13917),.dinb(n13904),.dout(n13918),.clk(gclk));
	jand g13673(.dina(n13918),.dinb(w_n11858_29[1]),.dout(n13919),.clk(gclk));
	jor g13674(.dina(w_n13534_0[0]),.dinb(n13919),.dout(n13920),.clk(gclk));
	jand g13675(.dina(n13920),.dinb(n13903),.dout(n13921),.clk(gclk));
	jand g13676(.dina(n13921),.dinb(w_n11347_23[1]),.dout(n13922),.clk(gclk));
	jor g13677(.dina(w_n13542_0[0]),.dinb(n13922),.dout(n13923),.clk(gclk));
	jand g13678(.dina(n13923),.dinb(n13902),.dout(n13924),.clk(gclk));
	jand g13679(.dina(n13924),.dinb(w_n10824_30[0]),.dout(n13925),.clk(gclk));
	jnot g13680(.din(w_n13550_0[0]),.dout(n13926),.clk(gclk));
	jor g13681(.dina(w_n13926_0[1]),.dinb(n13925),.dout(n13927),.clk(gclk));
	jand g13682(.dina(n13927),.dinb(n13901),.dout(n13928),.clk(gclk));
	jand g13683(.dina(n13928),.dinb(w_n10328_24[1]),.dout(n13929),.clk(gclk));
	jor g13684(.dina(w_n13557_0[0]),.dinb(n13929),.dout(n13930),.clk(gclk));
	jand g13685(.dina(n13930),.dinb(n13900),.dout(n13931),.clk(gclk));
	jand g13686(.dina(n13931),.dinb(w_n9832_30[2]),.dout(n13932),.clk(gclk));
	jnot g13687(.din(w_n13565_0[0]),.dout(n13933),.clk(gclk));
	jor g13688(.dina(w_n13933_0[1]),.dinb(n13932),.dout(n13934),.clk(gclk));
	jand g13689(.dina(n13934),.dinb(n13899),.dout(n13935),.clk(gclk));
	jand g13690(.dina(n13935),.dinb(w_n9369_25[1]),.dout(n13936),.clk(gclk));
	jor g13691(.dina(w_n13572_0[0]),.dinb(n13936),.dout(n13937),.clk(gclk));
	jand g13692(.dina(n13937),.dinb(n13898),.dout(n13938),.clk(gclk));
	jand g13693(.dina(n13938),.dinb(w_n8890_31[0]),.dout(n13939),.clk(gclk));
	jnot g13694(.din(w_n13580_0[0]),.dout(n13940),.clk(gclk));
	jor g13695(.dina(w_n13940_0[1]),.dinb(n13939),.dout(n13941),.clk(gclk));
	jand g13696(.dina(n13941),.dinb(n13897),.dout(n13942),.clk(gclk));
	jand g13697(.dina(n13942),.dinb(w_n8449_26[0]),.dout(n13943),.clk(gclk));
	jor g13698(.dina(w_n13587_0[0]),.dinb(n13943),.dout(n13944),.clk(gclk));
	jand g13699(.dina(n13944),.dinb(n13896),.dout(n13945),.clk(gclk));
	jand g13700(.dina(n13945),.dinb(w_n8003_31[2]),.dout(n13946),.clk(gclk));
	jnot g13701(.din(w_n13595_0[0]),.dout(n13947),.clk(gclk));
	jor g13702(.dina(w_n13947_0[1]),.dinb(n13946),.dout(n13948),.clk(gclk));
	jand g13703(.dina(n13948),.dinb(n13895),.dout(n13949),.clk(gclk));
	jand g13704(.dina(n13949),.dinb(w_n7581_27[0]),.dout(n13950),.clk(gclk));
	jor g13705(.dina(w_n13602_0[0]),.dinb(n13950),.dout(n13951),.clk(gclk));
	jand g13706(.dina(n13951),.dinb(n13894),.dout(n13952),.clk(gclk));
	jand g13707(.dina(n13952),.dinb(w_n7154_32[0]),.dout(n13953),.clk(gclk));
	jor g13708(.dina(w_n13610_0[0]),.dinb(n13953),.dout(n13954),.clk(gclk));
	jand g13709(.dina(n13954),.dinb(n13893),.dout(n13955),.clk(gclk));
	jand g13710(.dina(n13955),.dinb(w_n6758_27[2]),.dout(n13956),.clk(gclk));
	jor g13711(.dina(w_n13618_0[0]),.dinb(n13956),.dout(n13957),.clk(gclk));
	jand g13712(.dina(n13957),.dinb(n13892),.dout(n13958),.clk(gclk));
	jand g13713(.dina(n13958),.dinb(w_n6357_32[1]),.dout(n13959),.clk(gclk));
	jnot g13714(.din(w_n13626_0[0]),.dout(n13960),.clk(gclk));
	jor g13715(.dina(w_n13960_0[1]),.dinb(n13959),.dout(n13961),.clk(gclk));
	jand g13716(.dina(n13961),.dinb(n13891),.dout(n13962),.clk(gclk));
	jand g13717(.dina(n13962),.dinb(w_n5989_28[1]),.dout(n13963),.clk(gclk));
	jor g13718(.dina(w_n13633_0[0]),.dinb(n13963),.dout(n13964),.clk(gclk));
	jand g13719(.dina(n13964),.dinb(n13890),.dout(n13965),.clk(gclk));
	jand g13720(.dina(n13965),.dinb(w_n5606_32[2]),.dout(n13966),.clk(gclk));
	jnot g13721(.din(w_n13641_0[0]),.dout(n13967),.clk(gclk));
	jor g13722(.dina(w_n13967_0[1]),.dinb(n13966),.dout(n13968),.clk(gclk));
	jand g13723(.dina(n13968),.dinb(n13889),.dout(n13969),.clk(gclk));
	jand g13724(.dina(n13969),.dinb(w_n5259_29[1]),.dout(n13970),.clk(gclk));
	jor g13725(.dina(w_n13648_0[0]),.dinb(n13970),.dout(n13971),.clk(gclk));
	jand g13726(.dina(n13971),.dinb(n13888),.dout(n13972),.clk(gclk));
	jand g13727(.dina(n13972),.dinb(w_n4902_33[1]),.dout(n13973),.clk(gclk));
	jor g13728(.dina(w_n13656_0[0]),.dinb(n13973),.dout(n13974),.clk(gclk));
	jand g13729(.dina(n13974),.dinb(n13887),.dout(n13975),.clk(gclk));
	jand g13730(.dina(n13975),.dinb(w_n4582_30[1]),.dout(n13976),.clk(gclk));
	jor g13731(.dina(w_n13664_0[0]),.dinb(n13976),.dout(n13977),.clk(gclk));
	jand g13732(.dina(n13977),.dinb(n13886),.dout(n13978),.clk(gclk));
	jand g13733(.dina(n13978),.dinb(w_n4249_34[0]),.dout(n13979),.clk(gclk));
	jnot g13734(.din(w_n13672_0[0]),.dout(n13980),.clk(gclk));
	jor g13735(.dina(w_n13980_0[1]),.dinb(n13979),.dout(n13981),.clk(gclk));
	jand g13736(.dina(n13981),.dinb(n13885),.dout(n13982),.clk(gclk));
	jand g13737(.dina(n13982),.dinb(w_n3955_31[0]),.dout(n13983),.clk(gclk));
	jor g13738(.dina(w_n13679_0[0]),.dinb(n13983),.dout(n13984),.clk(gclk));
	jand g13739(.dina(n13984),.dinb(n13884),.dout(n13985),.clk(gclk));
	jand g13740(.dina(n13985),.dinb(w_n3642_34[1]),.dout(n13986),.clk(gclk));
	jor g13741(.dina(w_n13687_0[0]),.dinb(n13986),.dout(n13987),.clk(gclk));
	jand g13742(.dina(n13987),.dinb(n13883),.dout(n13988),.clk(gclk));
	jand g13743(.dina(n13988),.dinb(w_n3368_31[2]),.dout(n13989),.clk(gclk));
	jor g13744(.dina(w_n13695_0[0]),.dinb(n13989),.dout(n13990),.clk(gclk));
	jand g13745(.dina(n13990),.dinb(n13882),.dout(n13991),.clk(gclk));
	jand g13746(.dina(n13991),.dinb(w_n3089_35[0]),.dout(n13992),.clk(gclk));
	jor g13747(.dina(w_n13703_0[0]),.dinb(n13992),.dout(n13993),.clk(gclk));
	jand g13748(.dina(n13993),.dinb(n13881),.dout(n13994),.clk(gclk));
	jand g13749(.dina(n13994),.dinb(w_n2833_32[2]),.dout(n13995),.clk(gclk));
	jnot g13750(.din(w_n13711_0[0]),.dout(n13996),.clk(gclk));
	jor g13751(.dina(w_n13996_0[1]),.dinb(n13995),.dout(n13997),.clk(gclk));
	jand g13752(.dina(n13997),.dinb(n13880),.dout(n13998),.clk(gclk));
	jand g13753(.dina(n13998),.dinb(w_n2572_35[1]),.dout(n13999),.clk(gclk));
	jor g13754(.dina(n13999),.dinb(w_n13879_0[1]),.dout(n14000),.clk(gclk));
	jand g13755(.dina(n14000),.dinb(n13878),.dout(n14001),.clk(gclk));
	jand g13756(.dina(n14001),.dinb(w_n2345_33[1]),.dout(n14002),.clk(gclk));
	jor g13757(.dina(w_n13725_0[0]),.dinb(n14002),.dout(n14003),.clk(gclk));
	jand g13758(.dina(n14003),.dinb(n13877),.dout(n14004),.clk(gclk));
	jand g13759(.dina(n14004),.dinb(w_n2108_36[0]),.dout(n14005),.clk(gclk));
	jnot g13760(.din(w_n13733_0[0]),.dout(n14006),.clk(gclk));
	jor g13761(.dina(w_n14006_0[1]),.dinb(n14005),.dout(n14007),.clk(gclk));
	jand g13762(.dina(n14007),.dinb(n13876),.dout(n14008),.clk(gclk));
	jand g13763(.dina(n14008),.dinb(w_n1912_34[1]),.dout(n14009),.clk(gclk));
	jor g13764(.dina(w_n13740_0[0]),.dinb(n14009),.dout(n14010),.clk(gclk));
	jand g13765(.dina(n14010),.dinb(n13875),.dout(n14011),.clk(gclk));
	jand g13766(.dina(n14011),.dinb(w_n1699_36[2]),.dout(n14012),.clk(gclk));
	jnot g13767(.din(w_n13748_0[0]),.dout(n14013),.clk(gclk));
	jor g13768(.dina(w_n14013_0[1]),.dinb(n14012),.dout(n14014),.clk(gclk));
	jand g13769(.dina(n14014),.dinb(n13874),.dout(n14015),.clk(gclk));
	jand g13770(.dina(n14015),.dinb(w_n1516_35[0]),.dout(n14016),.clk(gclk));
	jor g13771(.dina(w_n13755_0[0]),.dinb(n14016),.dout(n14017),.clk(gclk));
	jand g13772(.dina(n14017),.dinb(n13873),.dout(n14018),.clk(gclk));
	jand g13773(.dina(n14018),.dinb(w_n1332_36[2]),.dout(n14019),.clk(gclk));
	jor g13774(.dina(w_n13763_0[0]),.dinb(n14019),.dout(n14020),.clk(gclk));
	jand g13775(.dina(n14020),.dinb(n13872),.dout(n14021),.clk(gclk));
	jand g13776(.dina(n14021),.dinb(w_n1173_35[2]),.dout(n14022),.clk(gclk));
	jor g13777(.dina(w_n13771_0[0]),.dinb(n14022),.dout(n14023),.clk(gclk));
	jand g13778(.dina(n14023),.dinb(n13871),.dout(n14024),.clk(gclk));
	jand g13779(.dina(n14024),.dinb(w_n1008_37[2]),.dout(n14025),.clk(gclk));
	jnot g13780(.din(w_n13779_0[0]),.dout(n14026),.clk(gclk));
	jor g13781(.dina(w_n14026_0[1]),.dinb(n14025),.dout(n14027),.clk(gclk));
	jand g13782(.dina(n14027),.dinb(n13870),.dout(n14028),.clk(gclk));
	jand g13783(.dina(n14028),.dinb(w_n884_36[2]),.dout(n14029),.clk(gclk));
	jor g13784(.dina(w_n13786_0[0]),.dinb(n14029),.dout(n14030),.clk(gclk));
	jand g13785(.dina(n14030),.dinb(n13869),.dout(n14031),.clk(gclk));
	jand g13786(.dina(n14031),.dinb(w_n743_37[2]),.dout(n14032),.clk(gclk));
	jnot g13787(.din(w_n13794_0[0]),.dout(n14033),.clk(gclk));
	jor g13788(.dina(w_n14033_0[1]),.dinb(n14032),.dout(n14034),.clk(gclk));
	jand g13789(.dina(n14034),.dinb(n13868),.dout(n14035),.clk(gclk));
	jand g13790(.dina(n14035),.dinb(w_n635_37[2]),.dout(n14036),.clk(gclk));
	jor g13791(.dina(w_n13801_0[0]),.dinb(n14036),.dout(n14037),.clk(gclk));
	jand g13792(.dina(n14037),.dinb(n13867),.dout(n14038),.clk(gclk));
	jand g13793(.dina(n14038),.dinb(w_n515_38[2]),.dout(n14039),.clk(gclk));
	jnot g13794(.din(w_n13809_0[0]),.dout(n14040),.clk(gclk));
	jor g13795(.dina(w_n14040_0[1]),.dinb(n14039),.dout(n14041),.clk(gclk));
	jand g13796(.dina(n14041),.dinb(n13866),.dout(n14042),.clk(gclk));
	jand g13797(.dina(n14042),.dinb(w_n443_38[2]),.dout(n14043),.clk(gclk));
	jor g13798(.dina(w_n13816_0[0]),.dinb(n14043),.dout(n14044),.clk(gclk));
	jand g13799(.dina(n14044),.dinb(n13865),.dout(n14045),.clk(gclk));
	jand g13800(.dina(n14045),.dinb(w_n352_39[0]),.dout(n14046),.clk(gclk));
	jnot g13801(.din(w_n13824_0[0]),.dout(n14047),.clk(gclk));
	jor g13802(.dina(w_n14047_0[1]),.dinb(n14046),.dout(n14048),.clk(gclk));
	jand g13803(.dina(n14048),.dinb(n13864),.dout(n14049),.clk(gclk));
	jand g13804(.dina(n14049),.dinb(w_n294_39[1]),.dout(n14050),.clk(gclk));
	jnot g13805(.din(w_n13831_0[0]),.dout(n14051),.clk(gclk));
	jor g13806(.dina(w_n14051_0[1]),.dinb(n14050),.dout(n14052),.clk(gclk));
	jand g13807(.dina(n14052),.dinb(n13863),.dout(n14053),.clk(gclk));
	jand g13808(.dina(n14053),.dinb(w_n239_39[1]),.dout(n14054),.clk(gclk));
	jnot g13809(.din(w_n13838_0[0]),.dout(n14055),.clk(gclk));
	jor g13810(.dina(w_n14055_0[1]),.dinb(n14054),.dout(n14056),.clk(gclk));
	jand g13811(.dina(n14056),.dinb(n13862),.dout(n14057),.clk(gclk));
	jand g13812(.dina(n14057),.dinb(w_n221_39[2]),.dout(n14058),.clk(gclk));
	jor g13813(.dina(w_n13845_0[0]),.dinb(n14058),.dout(n14059),.clk(gclk));
	jand g13814(.dina(n14059),.dinb(n13861),.dout(n14060),.clk(gclk));
	jor g13815(.dina(w_n13851_0[0]),.dinb(w_n14060_0[1]),.dout(n14061),.clk(gclk));
	jand g13816(.dina(w_asqrt18_19[2]),.dinb(w_n13510_0[0]),.dout(n14062),.clk(gclk));
	jor g13817(.dina(n14062),.dinb(w_n13287_0[1]),.dout(n14063),.clk(gclk));
	jor g13818(.dina(w_n14063_0[1]),.dinb(n14061),.dout(n14064),.clk(gclk));
	jand g13819(.dina(n14064),.dinb(w_n218_16[2]),.dout(n14065),.clk(gclk));
	jand g13820(.dina(w_n13515_22[0]),.dinb(w_n12951_0[0]),.dout(n14066),.clk(gclk));
	jor g13821(.dina(w_n14066_0[1]),.dinb(w_n14065_0[1]),.dout(n14067),.clk(gclk));
	jor g13822(.dina(n14067),.dinb(w_n13860_0[1]),.dout(n14068),.clk(gclk));
	jor g13823(.dina(n14068),.dinb(w_n13854_0[1]),.dout(asqrt_fa_18),.clk(gclk));
	jnot g13824(.din(w_n13860_0[0]),.dout(n14070),.clk(gclk));
	jand g13825(.dina(w_n13852_0[1]),.dinb(w_n13848_0[1]),.dout(n14071),.clk(gclk));
	jnot g13826(.din(w_n14063_0[0]),.dout(n14072),.clk(gclk));
	jand g13827(.dina(n14072),.dinb(n14071),.dout(n14073),.clk(gclk));
	jor g13828(.dina(n14073),.dinb(w_asqrt63_29[0]),.dout(n14074),.clk(gclk));
	jnot g13829(.din(w_n14066_0[0]),.dout(n14075),.clk(gclk));
	jand g13830(.dina(n14075),.dinb(n14074),.dout(n14076),.clk(gclk));
	jand g13831(.dina(n14076),.dinb(n14070),.dout(n14077),.clk(gclk));
	jand g13832(.dina(w_n14077_0[1]),.dinb(w_n13853_0[0]),.dout(n14078),.clk(gclk));
	jor g13833(.dina(w_n14078_42[1]),.dinb(w_n13296_1[0]),.dout(n14079),.clk(gclk));
	jnot g13834(.din(w_a32_0[2]),.dout(n14080),.clk(gclk));
	jnot g13835(.din(w_a33_0[1]),.dout(n14081),.clk(gclk));
	jand g13836(.dina(w_n14081_0[1]),.dinb(w_n14080_1[2]),.dout(n14082),.clk(gclk));
	jand g13837(.dina(w_n14082_0[2]),.dinb(w_n13296_0[2]),.dout(n14083),.clk(gclk));
	jnot g13838(.din(w_n14083_0[1]),.dout(n14084),.clk(gclk));
	jand g13839(.dina(n14084),.dinb(n14079),.dout(n14085),.clk(gclk));
	jor g13840(.dina(w_n14085_0[2]),.dinb(w_n13515_21[2]),.dout(n14086),.clk(gclk));
	jand g13841(.dina(w_n14085_0[1]),.dinb(w_n13515_21[1]),.dout(n14087),.clk(gclk));
	jor g13842(.dina(w_n14078_42[0]),.dinb(w_a34_1[0]),.dout(n14088),.clk(gclk));
	jand g13843(.dina(n14088),.dinb(w_a35_0[0]),.dout(n14089),.clk(gclk));
	jand g13844(.dina(w_asqrt17_13[1]),.dinb(w_n13298_0[1]),.dout(n14090),.clk(gclk));
	jor g13845(.dina(n14090),.dinb(n14089),.dout(n14091),.clk(gclk));
	jor g13846(.dina(n14091),.dinb(n14087),.dout(n14092),.clk(gclk));
	jand g13847(.dina(n14092),.dinb(w_n14086_0[1]),.dout(n14093),.clk(gclk));
	jor g13848(.dina(w_n14093_0[2]),.dinb(w_n12947_28[2]),.dout(n14094),.clk(gclk));
	jand g13849(.dina(w_n14093_0[1]),.dinb(w_n12947_28[1]),.dout(n14095),.clk(gclk));
	jnot g13850(.din(w_n13298_0[0]),.dout(n14096),.clk(gclk));
	jor g13851(.dina(w_n14078_41[2]),.dinb(n14096),.dout(n14097),.clk(gclk));
	jor g13852(.dina(w_n13854_0[0]),.dinb(w_n13515_21[0]),.dout(n14098),.clk(gclk));
	jor g13853(.dina(n14098),.dinb(w_n14065_0[0]),.dout(n14099),.clk(gclk));
	jor g13854(.dina(n14099),.dinb(w_n13859_0[0]),.dout(n14100),.clk(gclk));
	jand g13855(.dina(n14100),.dinb(w_n14097_0[1]),.dout(n14101),.clk(gclk));
	jxor g13856(.dina(n14101),.dinb(w_n12953_0[1]),.dout(n14102),.clk(gclk));
	jor g13857(.dina(w_n14102_0[2]),.dinb(n14095),.dout(n14103),.clk(gclk));
	jand g13858(.dina(n14103),.dinb(w_n14094_0[1]),.dout(n14104),.clk(gclk));
	jor g13859(.dina(w_n14104_0[2]),.dinb(w_n12410_22[1]),.dout(n14105),.clk(gclk));
	jand g13860(.dina(w_n14104_0[1]),.dinb(w_n12410_22[0]),.dout(n14106),.clk(gclk));
	jxor g13861(.dina(w_n13301_0[0]),.dinb(w_n12947_28[0]),.dout(n14107),.clk(gclk));
	jor g13862(.dina(n14107),.dinb(w_n14078_41[1]),.dout(n14108),.clk(gclk));
	jxor g13863(.dina(n14108),.dinb(w_n13913_0[0]),.dout(n14109),.clk(gclk));
	jnot g13864(.din(w_n14109_0[2]),.dout(n14110),.clk(gclk));
	jor g13865(.dina(n14110),.dinb(n14106),.dout(n14111),.clk(gclk));
	jand g13866(.dina(n14111),.dinb(w_n14105_0[1]),.dout(n14112),.clk(gclk));
	jor g13867(.dina(w_n14112_0[2]),.dinb(w_n11858_29[0]),.dout(n14113),.clk(gclk));
	jand g13868(.dina(w_n14112_0[1]),.dinb(w_n11858_28[2]),.dout(n14114),.clk(gclk));
	jxor g13869(.dina(w_n13519_0[0]),.dinb(w_n12410_21[2]),.dout(n14115),.clk(gclk));
	jor g13870(.dina(n14115),.dinb(w_n14078_41[0]),.dout(n14116),.clk(gclk));
	jxor g13871(.dina(n14116),.dinb(w_n13527_0[0]),.dout(n14117),.clk(gclk));
	jor g13872(.dina(w_n14117_0[2]),.dinb(n14114),.dout(n14118),.clk(gclk));
	jand g13873(.dina(n14118),.dinb(w_n14113_0[1]),.dout(n14119),.clk(gclk));
	jor g13874(.dina(w_n14119_0[2]),.dinb(w_n11347_23[0]),.dout(n14120),.clk(gclk));
	jand g13875(.dina(w_n14119_0[1]),.dinb(w_n11347_22[2]),.dout(n14121),.clk(gclk));
	jxor g13876(.dina(w_n13529_0[0]),.dinb(w_n11858_28[1]),.dout(n14122),.clk(gclk));
	jor g13877(.dina(n14122),.dinb(w_n14078_40[2]),.dout(n14123),.clk(gclk));
	jxor g13878(.dina(n14123),.dinb(w_n13535_0[0]),.dout(n14124),.clk(gclk));
	jor g13879(.dina(w_n14124_0[2]),.dinb(n14121),.dout(n14125),.clk(gclk));
	jand g13880(.dina(n14125),.dinb(w_n14120_0[1]),.dout(n14126),.clk(gclk));
	jor g13881(.dina(w_n14126_0[2]),.dinb(w_n10824_29[2]),.dout(n14127),.clk(gclk));
	jand g13882(.dina(w_n14126_0[1]),.dinb(w_n10824_29[1]),.dout(n14128),.clk(gclk));
	jxor g13883(.dina(w_n13537_0[0]),.dinb(w_n11347_22[1]),.dout(n14129),.clk(gclk));
	jor g13884(.dina(n14129),.dinb(w_n14078_40[1]),.dout(n14130),.clk(gclk));
	jxor g13885(.dina(n14130),.dinb(w_n13543_0[0]),.dout(n14131),.clk(gclk));
	jor g13886(.dina(w_n14131_0[2]),.dinb(n14128),.dout(n14132),.clk(gclk));
	jand g13887(.dina(n14132),.dinb(w_n14127_0[1]),.dout(n14133),.clk(gclk));
	jor g13888(.dina(w_n14133_0[2]),.dinb(w_n10328_24[0]),.dout(n14134),.clk(gclk));
	jand g13889(.dina(w_n14133_0[1]),.dinb(w_n10328_23[2]),.dout(n14135),.clk(gclk));
	jxor g13890(.dina(w_n13545_0[0]),.dinb(w_n10824_29[0]),.dout(n14136),.clk(gclk));
	jor g13891(.dina(n14136),.dinb(w_n14078_40[0]),.dout(n14137),.clk(gclk));
	jxor g13892(.dina(n14137),.dinb(w_n13926_0[0]),.dout(n14138),.clk(gclk));
	jnot g13893(.din(w_n14138_0[2]),.dout(n14139),.clk(gclk));
	jor g13894(.dina(n14139),.dinb(n14135),.dout(n14140),.clk(gclk));
	jand g13895(.dina(n14140),.dinb(w_n14134_0[1]),.dout(n14141),.clk(gclk));
	jor g13896(.dina(w_n14141_0[2]),.dinb(w_n9832_30[1]),.dout(n14142),.clk(gclk));
	jand g13897(.dina(w_n14141_0[1]),.dinb(w_n9832_30[0]),.dout(n14143),.clk(gclk));
	jxor g13898(.dina(w_n13552_0[0]),.dinb(w_n10328_23[1]),.dout(n14144),.clk(gclk));
	jor g13899(.dina(n14144),.dinb(w_n14078_39[2]),.dout(n14145),.clk(gclk));
	jxor g13900(.dina(n14145),.dinb(w_n13558_0[0]),.dout(n14146),.clk(gclk));
	jor g13901(.dina(w_n14146_0[2]),.dinb(n14143),.dout(n14147),.clk(gclk));
	jand g13902(.dina(n14147),.dinb(w_n14142_0[1]),.dout(n14148),.clk(gclk));
	jor g13903(.dina(w_n14148_0[2]),.dinb(w_n9369_25[0]),.dout(n14149),.clk(gclk));
	jand g13904(.dina(w_n14148_0[1]),.dinb(w_n9369_24[2]),.dout(n14150),.clk(gclk));
	jxor g13905(.dina(w_n13560_0[0]),.dinb(w_n9832_29[2]),.dout(n14151),.clk(gclk));
	jor g13906(.dina(n14151),.dinb(w_n14078_39[1]),.dout(n14152),.clk(gclk));
	jxor g13907(.dina(n14152),.dinb(w_n13933_0[0]),.dout(n14153),.clk(gclk));
	jnot g13908(.din(w_n14153_0[2]),.dout(n14154),.clk(gclk));
	jor g13909(.dina(n14154),.dinb(n14150),.dout(n14155),.clk(gclk));
	jand g13910(.dina(n14155),.dinb(w_n14149_0[1]),.dout(n14156),.clk(gclk));
	jor g13911(.dina(w_n14156_0[2]),.dinb(w_n8890_30[2]),.dout(n14157),.clk(gclk));
	jand g13912(.dina(w_n14156_0[1]),.dinb(w_n8890_30[1]),.dout(n14158),.clk(gclk));
	jxor g13913(.dina(w_n13567_0[0]),.dinb(w_n9369_24[1]),.dout(n14159),.clk(gclk));
	jor g13914(.dina(n14159),.dinb(w_n14078_39[0]),.dout(n14160),.clk(gclk));
	jxor g13915(.dina(n14160),.dinb(w_n13573_0[0]),.dout(n14161),.clk(gclk));
	jor g13916(.dina(w_n14161_0[2]),.dinb(n14158),.dout(n14162),.clk(gclk));
	jand g13917(.dina(n14162),.dinb(w_n14157_0[1]),.dout(n14163),.clk(gclk));
	jor g13918(.dina(w_n14163_0[2]),.dinb(w_n8449_25[2]),.dout(n14164),.clk(gclk));
	jand g13919(.dina(w_n14163_0[1]),.dinb(w_n8449_25[1]),.dout(n14165),.clk(gclk));
	jxor g13920(.dina(w_n13575_0[0]),.dinb(w_n8890_30[0]),.dout(n14166),.clk(gclk));
	jor g13921(.dina(n14166),.dinb(w_n14078_38[2]),.dout(n14167),.clk(gclk));
	jxor g13922(.dina(n14167),.dinb(w_n13940_0[0]),.dout(n14168),.clk(gclk));
	jnot g13923(.din(w_n14168_0[2]),.dout(n14169),.clk(gclk));
	jor g13924(.dina(n14169),.dinb(n14165),.dout(n14170),.clk(gclk));
	jand g13925(.dina(n14170),.dinb(w_n14164_0[1]),.dout(n14171),.clk(gclk));
	jor g13926(.dina(w_n14171_0[2]),.dinb(w_n8003_31[1]),.dout(n14172),.clk(gclk));
	jand g13927(.dina(w_n14171_0[1]),.dinb(w_n8003_31[0]),.dout(n14173),.clk(gclk));
	jxor g13928(.dina(w_n13582_0[0]),.dinb(w_n8449_25[0]),.dout(n14174),.clk(gclk));
	jor g13929(.dina(n14174),.dinb(w_n14078_38[1]),.dout(n14175),.clk(gclk));
	jxor g13930(.dina(n14175),.dinb(w_n13588_0[0]),.dout(n14176),.clk(gclk));
	jor g13931(.dina(w_n14176_0[2]),.dinb(n14173),.dout(n14177),.clk(gclk));
	jand g13932(.dina(n14177),.dinb(w_n14172_0[1]),.dout(n14178),.clk(gclk));
	jor g13933(.dina(w_n14178_0[2]),.dinb(w_n7581_26[2]),.dout(n14179),.clk(gclk));
	jand g13934(.dina(w_n14178_0[1]),.dinb(w_n7581_26[1]),.dout(n14180),.clk(gclk));
	jxor g13935(.dina(w_n13590_0[0]),.dinb(w_n8003_30[2]),.dout(n14181),.clk(gclk));
	jor g13936(.dina(n14181),.dinb(w_n14078_38[0]),.dout(n14182),.clk(gclk));
	jxor g13937(.dina(n14182),.dinb(w_n13947_0[0]),.dout(n14183),.clk(gclk));
	jnot g13938(.din(w_n14183_0[2]),.dout(n14184),.clk(gclk));
	jor g13939(.dina(n14184),.dinb(n14180),.dout(n14185),.clk(gclk));
	jand g13940(.dina(n14185),.dinb(w_n14179_0[1]),.dout(n14186),.clk(gclk));
	jor g13941(.dina(w_n14186_0[2]),.dinb(w_n7154_31[2]),.dout(n14187),.clk(gclk));
	jand g13942(.dina(w_n14186_0[1]),.dinb(w_n7154_31[1]),.dout(n14188),.clk(gclk));
	jxor g13943(.dina(w_n13597_0[0]),.dinb(w_n7581_26[0]),.dout(n14189),.clk(gclk));
	jor g13944(.dina(n14189),.dinb(w_n14078_37[2]),.dout(n14190),.clk(gclk));
	jxor g13945(.dina(n14190),.dinb(w_n13603_0[0]),.dout(n14191),.clk(gclk));
	jor g13946(.dina(w_n14191_0[2]),.dinb(n14188),.dout(n14192),.clk(gclk));
	jand g13947(.dina(n14192),.dinb(w_n14187_0[1]),.dout(n14193),.clk(gclk));
	jor g13948(.dina(w_n14193_0[2]),.dinb(w_n6758_27[1]),.dout(n14194),.clk(gclk));
	jand g13949(.dina(w_n14193_0[1]),.dinb(w_n6758_27[0]),.dout(n14195),.clk(gclk));
	jxor g13950(.dina(w_n13605_0[0]),.dinb(w_n7154_31[0]),.dout(n14196),.clk(gclk));
	jor g13951(.dina(n14196),.dinb(w_n14078_37[1]),.dout(n14197),.clk(gclk));
	jxor g13952(.dina(n14197),.dinb(w_n13611_0[0]),.dout(n14198),.clk(gclk));
	jor g13953(.dina(w_n14198_0[2]),.dinb(n14195),.dout(n14199),.clk(gclk));
	jand g13954(.dina(n14199),.dinb(w_n14194_0[1]),.dout(n14200),.clk(gclk));
	jor g13955(.dina(w_n14200_0[2]),.dinb(w_n6357_32[0]),.dout(n14201),.clk(gclk));
	jand g13956(.dina(w_n14200_0[1]),.dinb(w_n6357_31[2]),.dout(n14202),.clk(gclk));
	jxor g13957(.dina(w_n13613_0[0]),.dinb(w_n6758_26[2]),.dout(n14203),.clk(gclk));
	jor g13958(.dina(n14203),.dinb(w_n14078_37[0]),.dout(n14204),.clk(gclk));
	jxor g13959(.dina(n14204),.dinb(w_n13619_0[0]),.dout(n14205),.clk(gclk));
	jor g13960(.dina(w_n14205_0[2]),.dinb(n14202),.dout(n14206),.clk(gclk));
	jand g13961(.dina(n14206),.dinb(w_n14201_0[1]),.dout(n14207),.clk(gclk));
	jor g13962(.dina(w_n14207_0[2]),.dinb(w_n5989_28[0]),.dout(n14208),.clk(gclk));
	jand g13963(.dina(w_n14207_0[1]),.dinb(w_n5989_27[2]),.dout(n14209),.clk(gclk));
	jxor g13964(.dina(w_n13621_0[0]),.dinb(w_n6357_31[1]),.dout(n14210),.clk(gclk));
	jor g13965(.dina(n14210),.dinb(w_n14078_36[2]),.dout(n14211),.clk(gclk));
	jxor g13966(.dina(n14211),.dinb(w_n13960_0[0]),.dout(n14212),.clk(gclk));
	jnot g13967(.din(w_n14212_0[2]),.dout(n14213),.clk(gclk));
	jor g13968(.dina(n14213),.dinb(n14209),.dout(n14214),.clk(gclk));
	jand g13969(.dina(n14214),.dinb(w_n14208_0[1]),.dout(n14215),.clk(gclk));
	jor g13970(.dina(w_n14215_0[2]),.dinb(w_n5606_32[1]),.dout(n14216),.clk(gclk));
	jand g13971(.dina(w_n14215_0[1]),.dinb(w_n5606_32[0]),.dout(n14217),.clk(gclk));
	jxor g13972(.dina(w_n13628_0[0]),.dinb(w_n5989_27[1]),.dout(n14218),.clk(gclk));
	jor g13973(.dina(n14218),.dinb(w_n14078_36[1]),.dout(n14219),.clk(gclk));
	jxor g13974(.dina(n14219),.dinb(w_n13634_0[0]),.dout(n14220),.clk(gclk));
	jor g13975(.dina(w_n14220_0[2]),.dinb(n14217),.dout(n14221),.clk(gclk));
	jand g13976(.dina(n14221),.dinb(w_n14216_0[1]),.dout(n14222),.clk(gclk));
	jor g13977(.dina(w_n14222_0[2]),.dinb(w_n5259_29[0]),.dout(n14223),.clk(gclk));
	jand g13978(.dina(w_n14222_0[1]),.dinb(w_n5259_28[2]),.dout(n14224),.clk(gclk));
	jxor g13979(.dina(w_n13636_0[0]),.dinb(w_n5606_31[2]),.dout(n14225),.clk(gclk));
	jor g13980(.dina(n14225),.dinb(w_n14078_36[0]),.dout(n14226),.clk(gclk));
	jxor g13981(.dina(n14226),.dinb(w_n13967_0[0]),.dout(n14227),.clk(gclk));
	jnot g13982(.din(w_n14227_0[2]),.dout(n14228),.clk(gclk));
	jor g13983(.dina(n14228),.dinb(n14224),.dout(n14229),.clk(gclk));
	jand g13984(.dina(n14229),.dinb(w_n14223_0[1]),.dout(n14230),.clk(gclk));
	jor g13985(.dina(w_n14230_0[2]),.dinb(w_n4902_33[0]),.dout(n14231),.clk(gclk));
	jand g13986(.dina(w_n14230_0[1]),.dinb(w_n4902_32[2]),.dout(n14232),.clk(gclk));
	jxor g13987(.dina(w_n13643_0[0]),.dinb(w_n5259_28[1]),.dout(n14233),.clk(gclk));
	jor g13988(.dina(n14233),.dinb(w_n14078_35[2]),.dout(n14234),.clk(gclk));
	jxor g13989(.dina(n14234),.dinb(w_n13649_0[0]),.dout(n14235),.clk(gclk));
	jor g13990(.dina(w_n14235_0[2]),.dinb(n14232),.dout(n14236),.clk(gclk));
	jand g13991(.dina(n14236),.dinb(w_n14231_0[1]),.dout(n14237),.clk(gclk));
	jor g13992(.dina(w_n14237_0[2]),.dinb(w_n4582_30[0]),.dout(n14238),.clk(gclk));
	jand g13993(.dina(w_n14237_0[1]),.dinb(w_n4582_29[2]),.dout(n14239),.clk(gclk));
	jxor g13994(.dina(w_n13651_0[0]),.dinb(w_n4902_32[1]),.dout(n14240),.clk(gclk));
	jor g13995(.dina(n14240),.dinb(w_n14078_35[1]),.dout(n14241),.clk(gclk));
	jxor g13996(.dina(n14241),.dinb(w_n13657_0[0]),.dout(n14242),.clk(gclk));
	jor g13997(.dina(w_n14242_0[2]),.dinb(n14239),.dout(n14243),.clk(gclk));
	jand g13998(.dina(n14243),.dinb(w_n14238_0[1]),.dout(n14244),.clk(gclk));
	jor g13999(.dina(w_n14244_0[2]),.dinb(w_n4249_33[2]),.dout(n14245),.clk(gclk));
	jand g14000(.dina(w_n14244_0[1]),.dinb(w_n4249_33[1]),.dout(n14246),.clk(gclk));
	jxor g14001(.dina(w_n13659_0[0]),.dinb(w_n4582_29[1]),.dout(n14247),.clk(gclk));
	jor g14002(.dina(n14247),.dinb(w_n14078_35[0]),.dout(n14248),.clk(gclk));
	jxor g14003(.dina(n14248),.dinb(w_n13665_0[0]),.dout(n14249),.clk(gclk));
	jor g14004(.dina(w_n14249_0[2]),.dinb(n14246),.dout(n14250),.clk(gclk));
	jand g14005(.dina(n14250),.dinb(w_n14245_0[1]),.dout(n14251),.clk(gclk));
	jor g14006(.dina(w_n14251_0[2]),.dinb(w_n3955_30[2]),.dout(n14252),.clk(gclk));
	jand g14007(.dina(w_n14251_0[1]),.dinb(w_n3955_30[1]),.dout(n14253),.clk(gclk));
	jxor g14008(.dina(w_n13667_0[0]),.dinb(w_n4249_33[0]),.dout(n14254),.clk(gclk));
	jor g14009(.dina(n14254),.dinb(w_n14078_34[2]),.dout(n14255),.clk(gclk));
	jxor g14010(.dina(n14255),.dinb(w_n13980_0[0]),.dout(n14256),.clk(gclk));
	jnot g14011(.din(w_n14256_0[2]),.dout(n14257),.clk(gclk));
	jor g14012(.dina(n14257),.dinb(n14253),.dout(n14258),.clk(gclk));
	jand g14013(.dina(n14258),.dinb(w_n14252_0[1]),.dout(n14259),.clk(gclk));
	jor g14014(.dina(w_n14259_0[2]),.dinb(w_n3642_34[0]),.dout(n14260),.clk(gclk));
	jand g14015(.dina(w_n14259_0[1]),.dinb(w_n3642_33[2]),.dout(n14261),.clk(gclk));
	jxor g14016(.dina(w_n13674_0[0]),.dinb(w_n3955_30[0]),.dout(n14262),.clk(gclk));
	jor g14017(.dina(n14262),.dinb(w_n14078_34[1]),.dout(n14263),.clk(gclk));
	jxor g14018(.dina(n14263),.dinb(w_n13680_0[0]),.dout(n14264),.clk(gclk));
	jor g14019(.dina(w_n14264_0[2]),.dinb(n14261),.dout(n14265),.clk(gclk));
	jand g14020(.dina(n14265),.dinb(w_n14260_0[1]),.dout(n14266),.clk(gclk));
	jor g14021(.dina(w_n14266_0[2]),.dinb(w_n3368_31[1]),.dout(n14267),.clk(gclk));
	jand g14022(.dina(w_n14266_0[1]),.dinb(w_n3368_31[0]),.dout(n14268),.clk(gclk));
	jxor g14023(.dina(w_n13682_0[0]),.dinb(w_n3642_33[1]),.dout(n14269),.clk(gclk));
	jor g14024(.dina(n14269),.dinb(w_n14078_34[0]),.dout(n14270),.clk(gclk));
	jxor g14025(.dina(n14270),.dinb(w_n13688_0[0]),.dout(n14271),.clk(gclk));
	jor g14026(.dina(w_n14271_0[1]),.dinb(n14268),.dout(n14272),.clk(gclk));
	jand g14027(.dina(n14272),.dinb(w_n14267_0[1]),.dout(n14273),.clk(gclk));
	jor g14028(.dina(w_n14273_0[2]),.dinb(w_n3089_34[2]),.dout(n14274),.clk(gclk));
	jand g14029(.dina(w_n14273_0[1]),.dinb(w_n3089_34[1]),.dout(n14275),.clk(gclk));
	jxor g14030(.dina(w_n13690_0[0]),.dinb(w_n3368_30[2]),.dout(n14276),.clk(gclk));
	jor g14031(.dina(n14276),.dinb(w_n14078_33[2]),.dout(n14277),.clk(gclk));
	jxor g14032(.dina(n14277),.dinb(w_n13696_0[0]),.dout(n14278),.clk(gclk));
	jor g14033(.dina(w_n14278_0[2]),.dinb(n14275),.dout(n14279),.clk(gclk));
	jand g14034(.dina(n14279),.dinb(w_n14274_0[1]),.dout(n14280),.clk(gclk));
	jor g14035(.dina(w_n14280_0[2]),.dinb(w_n2833_32[1]),.dout(n14281),.clk(gclk));
	jand g14036(.dina(w_n14280_0[1]),.dinb(w_n2833_32[0]),.dout(n14282),.clk(gclk));
	jxor g14037(.dina(w_n13698_0[0]),.dinb(w_n3089_34[0]),.dout(n14283),.clk(gclk));
	jor g14038(.dina(n14283),.dinb(w_n14078_33[1]),.dout(n14284),.clk(gclk));
	jxor g14039(.dina(n14284),.dinb(w_n13704_0[0]),.dout(n14285),.clk(gclk));
	jor g14040(.dina(w_n14285_0[2]),.dinb(n14282),.dout(n14286),.clk(gclk));
	jand g14041(.dina(n14286),.dinb(w_n14281_0[1]),.dout(n14287),.clk(gclk));
	jor g14042(.dina(w_n14287_0[2]),.dinb(w_n2572_35[0]),.dout(n14288),.clk(gclk));
	jand g14043(.dina(w_n14287_0[1]),.dinb(w_n2572_34[2]),.dout(n14289),.clk(gclk));
	jxor g14044(.dina(w_n13706_0[0]),.dinb(w_n2833_31[2]),.dout(n14290),.clk(gclk));
	jor g14045(.dina(n14290),.dinb(w_n14078_33[0]),.dout(n14291),.clk(gclk));
	jxor g14046(.dina(n14291),.dinb(w_n13996_0[0]),.dout(n14292),.clk(gclk));
	jnot g14047(.din(w_n14292_0[2]),.dout(n14293),.clk(gclk));
	jor g14048(.dina(n14293),.dinb(n14289),.dout(n14294),.clk(gclk));
	jand g14049(.dina(n14294),.dinb(w_n14288_0[1]),.dout(n14295),.clk(gclk));
	jor g14050(.dina(w_n14295_0[2]),.dinb(w_n2345_33[0]),.dout(n14296),.clk(gclk));
	jxor g14051(.dina(w_n13713_0[0]),.dinb(w_n2572_34[1]),.dout(n14297),.clk(gclk));
	jor g14052(.dina(n14297),.dinb(w_n14078_32[2]),.dout(n14298),.clk(gclk));
	jxor g14053(.dina(n14298),.dinb(w_n13879_0[0]),.dout(n14299),.clk(gclk));
	jnot g14054(.din(w_n14299_0[2]),.dout(n14300),.clk(gclk));
	jand g14055(.dina(w_n14295_0[1]),.dinb(w_n2345_32[2]),.dout(n14301),.clk(gclk));
	jor g14056(.dina(n14301),.dinb(n14300),.dout(n14302),.clk(gclk));
	jand g14057(.dina(n14302),.dinb(w_n14296_0[1]),.dout(n14303),.clk(gclk));
	jor g14058(.dina(w_n14303_0[2]),.dinb(w_n2108_35[2]),.dout(n14304),.clk(gclk));
	jand g14059(.dina(w_n14303_0[1]),.dinb(w_n2108_35[1]),.dout(n14305),.clk(gclk));
	jxor g14060(.dina(w_n13720_0[0]),.dinb(w_n2345_32[1]),.dout(n14306),.clk(gclk));
	jor g14061(.dina(n14306),.dinb(w_n14078_32[1]),.dout(n14307),.clk(gclk));
	jxor g14062(.dina(n14307),.dinb(w_n13726_0[0]),.dout(n14308),.clk(gclk));
	jor g14063(.dina(w_n14308_0[2]),.dinb(n14305),.dout(n14309),.clk(gclk));
	jand g14064(.dina(n14309),.dinb(w_n14304_0[1]),.dout(n14310),.clk(gclk));
	jor g14065(.dina(w_n14310_0[2]),.dinb(w_n1912_34[0]),.dout(n14311),.clk(gclk));
	jand g14066(.dina(w_n14310_0[1]),.dinb(w_n1912_33[2]),.dout(n14312),.clk(gclk));
	jxor g14067(.dina(w_n13728_0[0]),.dinb(w_n2108_35[0]),.dout(n14313),.clk(gclk));
	jor g14068(.dina(n14313),.dinb(w_n14078_32[0]),.dout(n14314),.clk(gclk));
	jxor g14069(.dina(n14314),.dinb(w_n14006_0[0]),.dout(n14315),.clk(gclk));
	jnot g14070(.din(w_n14315_0[2]),.dout(n14316),.clk(gclk));
	jor g14071(.dina(n14316),.dinb(n14312),.dout(n14317),.clk(gclk));
	jand g14072(.dina(n14317),.dinb(w_n14311_0[1]),.dout(n14318),.clk(gclk));
	jor g14073(.dina(w_n14318_0[2]),.dinb(w_n1699_36[1]),.dout(n14319),.clk(gclk));
	jand g14074(.dina(w_n14318_0[1]),.dinb(w_n1699_36[0]),.dout(n14320),.clk(gclk));
	jxor g14075(.dina(w_n13735_0[0]),.dinb(w_n1912_33[1]),.dout(n14321),.clk(gclk));
	jor g14076(.dina(n14321),.dinb(w_n14078_31[2]),.dout(n14322),.clk(gclk));
	jxor g14077(.dina(n14322),.dinb(w_n13741_0[0]),.dout(n14323),.clk(gclk));
	jor g14078(.dina(w_n14323_0[2]),.dinb(n14320),.dout(n14324),.clk(gclk));
	jand g14079(.dina(n14324),.dinb(w_n14319_0[1]),.dout(n14325),.clk(gclk));
	jor g14080(.dina(w_n14325_0[2]),.dinb(w_n1516_34[2]),.dout(n14326),.clk(gclk));
	jand g14081(.dina(w_n14325_0[1]),.dinb(w_n1516_34[1]),.dout(n14327),.clk(gclk));
	jxor g14082(.dina(w_n13743_0[0]),.dinb(w_n1699_35[2]),.dout(n14328),.clk(gclk));
	jor g14083(.dina(n14328),.dinb(w_n14078_31[1]),.dout(n14329),.clk(gclk));
	jxor g14084(.dina(n14329),.dinb(w_n14013_0[0]),.dout(n14330),.clk(gclk));
	jnot g14085(.din(w_n14330_0[2]),.dout(n14331),.clk(gclk));
	jor g14086(.dina(n14331),.dinb(n14327),.dout(n14332),.clk(gclk));
	jand g14087(.dina(n14332),.dinb(w_n14326_0[1]),.dout(n14333),.clk(gclk));
	jor g14088(.dina(w_n14333_0[2]),.dinb(w_n1332_36[1]),.dout(n14334),.clk(gclk));
	jand g14089(.dina(w_n14333_0[1]),.dinb(w_n1332_36[0]),.dout(n14335),.clk(gclk));
	jxor g14090(.dina(w_n13750_0[0]),.dinb(w_n1516_34[0]),.dout(n14336),.clk(gclk));
	jor g14091(.dina(n14336),.dinb(w_n14078_31[0]),.dout(n14337),.clk(gclk));
	jxor g14092(.dina(n14337),.dinb(w_n13756_0[0]),.dout(n14338),.clk(gclk));
	jor g14093(.dina(w_n14338_0[2]),.dinb(n14335),.dout(n14339),.clk(gclk));
	jand g14094(.dina(n14339),.dinb(w_n14334_0[1]),.dout(n14340),.clk(gclk));
	jor g14095(.dina(w_n14340_0[2]),.dinb(w_n1173_35[1]),.dout(n14341),.clk(gclk));
	jand g14096(.dina(w_n14340_0[1]),.dinb(w_n1173_35[0]),.dout(n14342),.clk(gclk));
	jxor g14097(.dina(w_n13758_0[0]),.dinb(w_n1332_35[2]),.dout(n14343),.clk(gclk));
	jor g14098(.dina(n14343),.dinb(w_n14078_30[2]),.dout(n14344),.clk(gclk));
	jxor g14099(.dina(n14344),.dinb(w_n13764_0[0]),.dout(n14345),.clk(gclk));
	jor g14100(.dina(w_n14345_0[2]),.dinb(n14342),.dout(n14346),.clk(gclk));
	jand g14101(.dina(n14346),.dinb(w_n14341_0[1]),.dout(n14347),.clk(gclk));
	jor g14102(.dina(w_n14347_0[2]),.dinb(w_n1008_37[1]),.dout(n14348),.clk(gclk));
	jand g14103(.dina(w_n14347_0[1]),.dinb(w_n1008_37[0]),.dout(n14349),.clk(gclk));
	jxor g14104(.dina(w_n13766_0[0]),.dinb(w_n1173_34[2]),.dout(n14350),.clk(gclk));
	jor g14105(.dina(n14350),.dinb(w_n14078_30[1]),.dout(n14351),.clk(gclk));
	jxor g14106(.dina(n14351),.dinb(w_n13772_0[0]),.dout(n14352),.clk(gclk));
	jor g14107(.dina(w_n14352_0[2]),.dinb(n14349),.dout(n14353),.clk(gclk));
	jand g14108(.dina(n14353),.dinb(w_n14348_0[1]),.dout(n14354),.clk(gclk));
	jor g14109(.dina(w_n14354_0[2]),.dinb(w_n884_36[1]),.dout(n14355),.clk(gclk));
	jand g14110(.dina(w_n14354_0[1]),.dinb(w_n884_36[0]),.dout(n14356),.clk(gclk));
	jxor g14111(.dina(w_n13774_0[0]),.dinb(w_n1008_36[2]),.dout(n14357),.clk(gclk));
	jor g14112(.dina(n14357),.dinb(w_n14078_30[0]),.dout(n14358),.clk(gclk));
	jxor g14113(.dina(n14358),.dinb(w_n14026_0[0]),.dout(n14359),.clk(gclk));
	jnot g14114(.din(w_n14359_0[2]),.dout(n14360),.clk(gclk));
	jor g14115(.dina(n14360),.dinb(n14356),.dout(n14361),.clk(gclk));
	jand g14116(.dina(n14361),.dinb(w_n14355_0[1]),.dout(n14362),.clk(gclk));
	jor g14117(.dina(w_n14362_0[2]),.dinb(w_n743_37[1]),.dout(n14363),.clk(gclk));
	jand g14118(.dina(w_n14362_0[1]),.dinb(w_n743_37[0]),.dout(n14364),.clk(gclk));
	jxor g14119(.dina(w_n13781_0[0]),.dinb(w_n884_35[2]),.dout(n14365),.clk(gclk));
	jor g14120(.dina(n14365),.dinb(w_n14078_29[2]),.dout(n14366),.clk(gclk));
	jxor g14121(.dina(n14366),.dinb(w_n13787_0[0]),.dout(n14367),.clk(gclk));
	jor g14122(.dina(w_n14367_0[2]),.dinb(n14364),.dout(n14368),.clk(gclk));
	jand g14123(.dina(n14368),.dinb(w_n14363_0[1]),.dout(n14369),.clk(gclk));
	jor g14124(.dina(w_n14369_0[2]),.dinb(w_n635_37[1]),.dout(n14370),.clk(gclk));
	jand g14125(.dina(w_n14369_0[1]),.dinb(w_n635_37[0]),.dout(n14371),.clk(gclk));
	jxor g14126(.dina(w_n13789_0[0]),.dinb(w_n743_36[2]),.dout(n14372),.clk(gclk));
	jor g14127(.dina(n14372),.dinb(w_n14078_29[1]),.dout(n14373),.clk(gclk));
	jxor g14128(.dina(n14373),.dinb(w_n14033_0[0]),.dout(n14374),.clk(gclk));
	jnot g14129(.din(w_n14374_0[2]),.dout(n14375),.clk(gclk));
	jor g14130(.dina(n14375),.dinb(n14371),.dout(n14376),.clk(gclk));
	jand g14131(.dina(n14376),.dinb(w_n14370_0[1]),.dout(n14377),.clk(gclk));
	jor g14132(.dina(w_n14377_0[2]),.dinb(w_n515_38[1]),.dout(n14378),.clk(gclk));
	jand g14133(.dina(w_n14377_0[1]),.dinb(w_n515_38[0]),.dout(n14379),.clk(gclk));
	jxor g14134(.dina(w_n13796_0[0]),.dinb(w_n635_36[2]),.dout(n14380),.clk(gclk));
	jor g14135(.dina(n14380),.dinb(w_n14078_29[0]),.dout(n14381),.clk(gclk));
	jxor g14136(.dina(n14381),.dinb(w_n13802_0[0]),.dout(n14382),.clk(gclk));
	jor g14137(.dina(w_n14382_0[2]),.dinb(n14379),.dout(n14383),.clk(gclk));
	jand g14138(.dina(n14383),.dinb(w_n14378_0[1]),.dout(n14384),.clk(gclk));
	jor g14139(.dina(w_n14384_0[2]),.dinb(w_n443_38[1]),.dout(n14385),.clk(gclk));
	jand g14140(.dina(w_n14384_0[1]),.dinb(w_n443_38[0]),.dout(n14386),.clk(gclk));
	jxor g14141(.dina(w_n13804_0[0]),.dinb(w_n515_37[2]),.dout(n14387),.clk(gclk));
	jor g14142(.dina(n14387),.dinb(w_n14078_28[2]),.dout(n14388),.clk(gclk));
	jxor g14143(.dina(n14388),.dinb(w_n14040_0[0]),.dout(n14389),.clk(gclk));
	jnot g14144(.din(w_n14389_0[2]),.dout(n14390),.clk(gclk));
	jor g14145(.dina(n14390),.dinb(n14386),.dout(n14391),.clk(gclk));
	jand g14146(.dina(n14391),.dinb(w_n14385_0[1]),.dout(n14392),.clk(gclk));
	jor g14147(.dina(w_n14392_0[2]),.dinb(w_n352_38[2]),.dout(n14393),.clk(gclk));
	jand g14148(.dina(w_n14392_0[1]),.dinb(w_n352_38[1]),.dout(n14394),.clk(gclk));
	jxor g14149(.dina(w_n13811_0[0]),.dinb(w_n443_37[2]),.dout(n14395),.clk(gclk));
	jor g14150(.dina(n14395),.dinb(w_n14078_28[1]),.dout(n14396),.clk(gclk));
	jxor g14151(.dina(n14396),.dinb(w_n13817_0[0]),.dout(n14397),.clk(gclk));
	jor g14152(.dina(w_n14397_0[2]),.dinb(n14394),.dout(n14398),.clk(gclk));
	jand g14153(.dina(n14398),.dinb(w_n14393_0[1]),.dout(n14399),.clk(gclk));
	jor g14154(.dina(w_n14399_0[2]),.dinb(w_n294_39[0]),.dout(n14400),.clk(gclk));
	jand g14155(.dina(w_n14399_0[1]),.dinb(w_n294_38[2]),.dout(n14401),.clk(gclk));
	jxor g14156(.dina(w_n13819_0[0]),.dinb(w_n352_38[0]),.dout(n14402),.clk(gclk));
	jor g14157(.dina(n14402),.dinb(w_n14078_28[0]),.dout(n14403),.clk(gclk));
	jxor g14158(.dina(n14403),.dinb(w_n14047_0[0]),.dout(n14404),.clk(gclk));
	jnot g14159(.din(w_n14404_0[2]),.dout(n14405),.clk(gclk));
	jor g14160(.dina(n14405),.dinb(n14401),.dout(n14406),.clk(gclk));
	jand g14161(.dina(n14406),.dinb(w_n14400_0[1]),.dout(n14407),.clk(gclk));
	jor g14162(.dina(w_n14407_0[2]),.dinb(w_n239_39[0]),.dout(n14408),.clk(gclk));
	jand g14163(.dina(w_n14407_0[1]),.dinb(w_n239_38[2]),.dout(n14409),.clk(gclk));
	jxor g14164(.dina(w_n13826_0[0]),.dinb(w_n294_38[1]),.dout(n14410),.clk(gclk));
	jor g14165(.dina(n14410),.dinb(w_n14078_27[2]),.dout(n14411),.clk(gclk));
	jxor g14166(.dina(n14411),.dinb(w_n14051_0[0]),.dout(n14412),.clk(gclk));
	jnot g14167(.din(w_n14412_0[2]),.dout(n14413),.clk(gclk));
	jor g14168(.dina(n14413),.dinb(n14409),.dout(n14414),.clk(gclk));
	jand g14169(.dina(n14414),.dinb(w_n14408_0[1]),.dout(n14415),.clk(gclk));
	jor g14170(.dina(w_n14415_0[2]),.dinb(w_n221_39[1]),.dout(n14416),.clk(gclk));
	jand g14171(.dina(w_n14415_0[1]),.dinb(w_n221_39[0]),.dout(n14417),.clk(gclk));
	jxor g14172(.dina(w_n13833_0[0]),.dinb(w_n239_38[1]),.dout(n14418),.clk(gclk));
	jor g14173(.dina(n14418),.dinb(w_n14078_27[1]),.dout(n14419),.clk(gclk));
	jxor g14174(.dina(n14419),.dinb(w_n14055_0[0]),.dout(n14420),.clk(gclk));
	jnot g14175(.din(w_n14420_0[1]),.dout(n14421),.clk(gclk));
	jor g14176(.dina(w_n14421_0[1]),.dinb(n14417),.dout(n14422),.clk(gclk));
	jand g14177(.dina(n14422),.dinb(w_n14416_0[1]),.dout(n14423),.clk(gclk));
	jxor g14178(.dina(w_n13840_0[0]),.dinb(w_n221_38[2]),.dout(n14424),.clk(gclk));
	jor g14179(.dina(n14424),.dinb(w_n14078_27[0]),.dout(n14425),.clk(gclk));
	jxor g14180(.dina(n14425),.dinb(w_n13846_0[0]),.dout(n14426),.clk(gclk));
	jand g14181(.dina(w_n14426_1[2]),.dinb(w_n14423_1[1]),.dout(n14427),.clk(gclk));
	jor g14182(.dina(w_n14426_1[1]),.dinb(w_n14423_1[0]),.dout(n14429),.clk(gclk));
	jxor g14183(.dina(w_n13852_0[0]),.dinb(w_n13848_0[0]),.dout(n14430),.clk(gclk));
	jnot g14184(.din(w_n14430_0[1]),.dout(n14431),.clk(gclk));
	jand g14185(.dina(n14431),.dinb(w_asqrt17_13[0]),.dout(n14432),.clk(gclk));
	jor g14186(.dina(w_n14432_0[1]),.dinb(n14429),.dout(n14433),.clk(gclk));
	jand g14187(.dina(n14433),.dinb(w_n218_16[1]),.dout(n14434),.clk(gclk));
	jand g14188(.dina(w_n14077_0[0]),.dinb(w_n14060_0[0]),.dout(n14435),.clk(gclk));
	jand g14189(.dina(w_n14430_0[0]),.dinb(w_asqrt63_28[2]),.dout(n14436),.clk(gclk));
	jnot g14190(.din(n14436),.dout(n14437),.clk(gclk));
	jor g14191(.dina(w_n14437_0[1]),.dinb(n14435),.dout(n14438),.clk(gclk));
	jnot g14192(.din(w_n14438_0[1]),.dout(n14439),.clk(gclk));
	jor g14193(.dina(n14439),.dinb(n14434),.dout(n14440),.clk(gclk));
	jor g14194(.dina(n14440),.dinb(w_n14427_0[1]),.dout(asqrt_fa_17),.clk(gclk));
	jnot g14195(.din(w_a30_1[1]),.dout(n14443),.clk(gclk));
	jnot g14196(.din(w_a31_0[1]),.dout(n14444),.clk(gclk));
	jand g14197(.dina(w_n14444_0[1]),.dinb(w_n14443_1[1]),.dout(n14445),.clk(gclk));
	jand g14198(.dina(w_n14445_0[2]),.dinb(w_n14080_1[1]),.dout(n14446),.clk(gclk));
	jand g14199(.dina(w_asqrt16_34[1]),.dinb(w_a32_0[1]),.dout(n14447),.clk(gclk));
	jor g14200(.dina(n14447),.dinb(w_n14446_0[1]),.dout(n14448),.clk(gclk));
	jand g14201(.dina(w_n14448_0[2]),.dinb(w_asqrt17_12[2]),.dout(n14449),.clk(gclk));
	jor g14202(.dina(w_n14448_0[1]),.dinb(w_asqrt17_12[1]),.dout(n14450),.clk(gclk));
	jand g14203(.dina(w_asqrt16_34[0]),.dinb(w_n14080_1[0]),.dout(n14451),.clk(gclk));
	jor g14204(.dina(n14451),.dinb(w_n14081_0[0]),.dout(n14452),.clk(gclk));
	jnot g14205(.din(w_n14082_0[1]),.dout(n14453),.clk(gclk));
	jnot g14206(.din(w_n14427_0[0]),.dout(n14454),.clk(gclk));
	jnot g14207(.din(w_n14416_0[0]),.dout(n14456),.clk(gclk));
	jnot g14208(.din(w_n14408_0[0]),.dout(n14457),.clk(gclk));
	jnot g14209(.din(w_n14400_0[0]),.dout(n14458),.clk(gclk));
	jnot g14210(.din(w_n14393_0[0]),.dout(n14459),.clk(gclk));
	jnot g14211(.din(w_n14385_0[0]),.dout(n14460),.clk(gclk));
	jnot g14212(.din(w_n14378_0[0]),.dout(n14461),.clk(gclk));
	jnot g14213(.din(w_n14370_0[0]),.dout(n14462),.clk(gclk));
	jnot g14214(.din(w_n14363_0[0]),.dout(n14463),.clk(gclk));
	jnot g14215(.din(w_n14355_0[0]),.dout(n14464),.clk(gclk));
	jnot g14216(.din(w_n14348_0[0]),.dout(n14465),.clk(gclk));
	jnot g14217(.din(w_n14341_0[0]),.dout(n14466),.clk(gclk));
	jnot g14218(.din(w_n14334_0[0]),.dout(n14467),.clk(gclk));
	jnot g14219(.din(w_n14326_0[0]),.dout(n14468),.clk(gclk));
	jnot g14220(.din(w_n14319_0[0]),.dout(n14469),.clk(gclk));
	jnot g14221(.din(w_n14311_0[0]),.dout(n14470),.clk(gclk));
	jnot g14222(.din(w_n14304_0[0]),.dout(n14471),.clk(gclk));
	jnot g14223(.din(w_n14296_0[0]),.dout(n14472),.clk(gclk));
	jnot g14224(.din(w_n14288_0[0]),.dout(n14473),.clk(gclk));
	jnot g14225(.din(w_n14281_0[0]),.dout(n14474),.clk(gclk));
	jnot g14226(.din(w_n14274_0[0]),.dout(n14475),.clk(gclk));
	jnot g14227(.din(w_n14267_0[0]),.dout(n14476),.clk(gclk));
	jnot g14228(.din(w_n14260_0[0]),.dout(n14477),.clk(gclk));
	jnot g14229(.din(w_n14252_0[0]),.dout(n14478),.clk(gclk));
	jnot g14230(.din(w_n14245_0[0]),.dout(n14479),.clk(gclk));
	jnot g14231(.din(w_n14238_0[0]),.dout(n14480),.clk(gclk));
	jnot g14232(.din(w_n14231_0[0]),.dout(n14481),.clk(gclk));
	jnot g14233(.din(w_n14223_0[0]),.dout(n14482),.clk(gclk));
	jnot g14234(.din(w_n14216_0[0]),.dout(n14483),.clk(gclk));
	jnot g14235(.din(w_n14208_0[0]),.dout(n14484),.clk(gclk));
	jnot g14236(.din(w_n14201_0[0]),.dout(n14485),.clk(gclk));
	jnot g14237(.din(w_n14194_0[0]),.dout(n14486),.clk(gclk));
	jnot g14238(.din(w_n14187_0[0]),.dout(n14487),.clk(gclk));
	jnot g14239(.din(w_n14179_0[0]),.dout(n14488),.clk(gclk));
	jnot g14240(.din(w_n14172_0[0]),.dout(n14489),.clk(gclk));
	jnot g14241(.din(w_n14164_0[0]),.dout(n14490),.clk(gclk));
	jnot g14242(.din(w_n14157_0[0]),.dout(n14491),.clk(gclk));
	jnot g14243(.din(w_n14149_0[0]),.dout(n14492),.clk(gclk));
	jnot g14244(.din(w_n14142_0[0]),.dout(n14493),.clk(gclk));
	jnot g14245(.din(w_n14134_0[0]),.dout(n14494),.clk(gclk));
	jnot g14246(.din(w_n14127_0[0]),.dout(n14495),.clk(gclk));
	jnot g14247(.din(w_n14120_0[0]),.dout(n14496),.clk(gclk));
	jnot g14248(.din(w_n14113_0[0]),.dout(n14497),.clk(gclk));
	jnot g14249(.din(w_n14105_0[0]),.dout(n14498),.clk(gclk));
	jnot g14250(.din(w_n14094_0[0]),.dout(n14499),.clk(gclk));
	jnot g14251(.din(w_n14086_0[0]),.dout(n14500),.clk(gclk));
	jand g14252(.dina(w_asqrt17_12[0]),.dinb(w_a34_0[2]),.dout(n14501),.clk(gclk));
	jor g14253(.dina(w_n14083_0[0]),.dinb(n14501),.dout(n14502),.clk(gclk));
	jor g14254(.dina(n14502),.dinb(w_asqrt18_19[1]),.dout(n14503),.clk(gclk));
	jand g14255(.dina(w_asqrt17_11[2]),.dinb(w_n13296_0[1]),.dout(n14504),.clk(gclk));
	jor g14256(.dina(n14504),.dinb(w_n13297_0[0]),.dout(n14505),.clk(gclk));
	jand g14257(.dina(w_n14097_0[0]),.dinb(n14505),.dout(n14506),.clk(gclk));
	jand g14258(.dina(w_n14506_0[1]),.dinb(n14503),.dout(n14507),.clk(gclk));
	jor g14259(.dina(n14507),.dinb(n14500),.dout(n14508),.clk(gclk));
	jor g14260(.dina(n14508),.dinb(w_asqrt19_12[1]),.dout(n14509),.clk(gclk));
	jnot g14261(.din(w_n14102_0[1]),.dout(n14510),.clk(gclk));
	jand g14262(.dina(n14510),.dinb(n14509),.dout(n14511),.clk(gclk));
	jor g14263(.dina(n14511),.dinb(n14499),.dout(n14512),.clk(gclk));
	jor g14264(.dina(n14512),.dinb(w_asqrt20_19[1]),.dout(n14513),.clk(gclk));
	jand g14265(.dina(w_n14109_0[1]),.dinb(n14513),.dout(n14514),.clk(gclk));
	jor g14266(.dina(n14514),.dinb(n14498),.dout(n14515),.clk(gclk));
	jor g14267(.dina(n14515),.dinb(w_asqrt21_13[0]),.dout(n14516),.clk(gclk));
	jnot g14268(.din(w_n14117_0[1]),.dout(n14517),.clk(gclk));
	jand g14269(.dina(n14517),.dinb(n14516),.dout(n14518),.clk(gclk));
	jor g14270(.dina(n14518),.dinb(n14497),.dout(n14519),.clk(gclk));
	jor g14271(.dina(n14519),.dinb(w_asqrt22_19[2]),.dout(n14520),.clk(gclk));
	jnot g14272(.din(w_n14124_0[1]),.dout(n14521),.clk(gclk));
	jand g14273(.dina(n14521),.dinb(n14520),.dout(n14522),.clk(gclk));
	jor g14274(.dina(n14522),.dinb(n14496),.dout(n14523),.clk(gclk));
	jor g14275(.dina(n14523),.dinb(w_asqrt23_13[2]),.dout(n14524),.clk(gclk));
	jnot g14276(.din(w_n14131_0[1]),.dout(n14525),.clk(gclk));
	jand g14277(.dina(n14525),.dinb(n14524),.dout(n14526),.clk(gclk));
	jor g14278(.dina(n14526),.dinb(n14495),.dout(n14527),.clk(gclk));
	jor g14279(.dina(n14527),.dinb(w_asqrt24_19[2]),.dout(n14528),.clk(gclk));
	jand g14280(.dina(w_n14138_0[1]),.dinb(n14528),.dout(n14529),.clk(gclk));
	jor g14281(.dina(n14529),.dinb(n14494),.dout(n14530),.clk(gclk));
	jor g14282(.dina(n14530),.dinb(w_asqrt25_13[2]),.dout(n14531),.clk(gclk));
	jnot g14283(.din(w_n14146_0[1]),.dout(n14532),.clk(gclk));
	jand g14284(.dina(n14532),.dinb(n14531),.dout(n14533),.clk(gclk));
	jor g14285(.dina(n14533),.dinb(n14493),.dout(n14534),.clk(gclk));
	jor g14286(.dina(n14534),.dinb(w_asqrt26_19[2]),.dout(n14535),.clk(gclk));
	jand g14287(.dina(w_n14153_0[1]),.dinb(n14535),.dout(n14536),.clk(gclk));
	jor g14288(.dina(n14536),.dinb(n14492),.dout(n14537),.clk(gclk));
	jor g14289(.dina(n14537),.dinb(w_asqrt27_14[1]),.dout(n14538),.clk(gclk));
	jnot g14290(.din(w_n14161_0[1]),.dout(n14539),.clk(gclk));
	jand g14291(.dina(n14539),.dinb(n14538),.dout(n14540),.clk(gclk));
	jor g14292(.dina(n14540),.dinb(n14491),.dout(n14541),.clk(gclk));
	jor g14293(.dina(n14541),.dinb(w_asqrt28_20[0]),.dout(n14542),.clk(gclk));
	jand g14294(.dina(w_n14168_0[1]),.dinb(n14542),.dout(n14543),.clk(gclk));
	jor g14295(.dina(n14543),.dinb(n14490),.dout(n14544),.clk(gclk));
	jor g14296(.dina(n14544),.dinb(w_asqrt29_14[2]),.dout(n14545),.clk(gclk));
	jnot g14297(.din(w_n14176_0[1]),.dout(n14546),.clk(gclk));
	jand g14298(.dina(n14546),.dinb(n14545),.dout(n14547),.clk(gclk));
	jor g14299(.dina(n14547),.dinb(n14489),.dout(n14548),.clk(gclk));
	jor g14300(.dina(n14548),.dinb(w_asqrt30_20[1]),.dout(n14549),.clk(gclk));
	jand g14301(.dina(w_n14183_0[1]),.dinb(n14549),.dout(n14550),.clk(gclk));
	jor g14302(.dina(n14550),.dinb(n14488),.dout(n14551),.clk(gclk));
	jor g14303(.dina(n14551),.dinb(w_asqrt31_15[1]),.dout(n14552),.clk(gclk));
	jnot g14304(.din(w_n14191_0[1]),.dout(n14553),.clk(gclk));
	jand g14305(.dina(n14553),.dinb(n14552),.dout(n14554),.clk(gclk));
	jor g14306(.dina(n14554),.dinb(n14487),.dout(n14555),.clk(gclk));
	jor g14307(.dina(n14555),.dinb(w_asqrt32_20[1]),.dout(n14556),.clk(gclk));
	jnot g14308(.din(w_n14198_0[1]),.dout(n14557),.clk(gclk));
	jand g14309(.dina(n14557),.dinb(n14556),.dout(n14558),.clk(gclk));
	jor g14310(.dina(n14558),.dinb(n14486),.dout(n14559),.clk(gclk));
	jor g14311(.dina(n14559),.dinb(w_asqrt33_16[0]),.dout(n14560),.clk(gclk));
	jnot g14312(.din(w_n14205_0[1]),.dout(n14561),.clk(gclk));
	jand g14313(.dina(n14561),.dinb(n14560),.dout(n14562),.clk(gclk));
	jor g14314(.dina(n14562),.dinb(n14485),.dout(n14563),.clk(gclk));
	jor g14315(.dina(n14563),.dinb(w_asqrt34_20[2]),.dout(n14564),.clk(gclk));
	jand g14316(.dina(w_n14212_0[1]),.dinb(n14564),.dout(n14565),.clk(gclk));
	jor g14317(.dina(n14565),.dinb(n14484),.dout(n14566),.clk(gclk));
	jor g14318(.dina(n14566),.dinb(w_asqrt35_16[2]),.dout(n14567),.clk(gclk));
	jnot g14319(.din(w_n14220_0[1]),.dout(n14568),.clk(gclk));
	jand g14320(.dina(n14568),.dinb(n14567),.dout(n14569),.clk(gclk));
	jor g14321(.dina(n14569),.dinb(n14483),.dout(n14570),.clk(gclk));
	jor g14322(.dina(n14570),.dinb(w_asqrt36_20[2]),.dout(n14571),.clk(gclk));
	jand g14323(.dina(w_n14227_0[1]),.dinb(n14571),.dout(n14572),.clk(gclk));
	jor g14324(.dina(n14572),.dinb(n14482),.dout(n14573),.clk(gclk));
	jor g14325(.dina(n14573),.dinb(w_asqrt37_17[0]),.dout(n14574),.clk(gclk));
	jnot g14326(.din(w_n14235_0[1]),.dout(n14575),.clk(gclk));
	jand g14327(.dina(n14575),.dinb(n14574),.dout(n14576),.clk(gclk));
	jor g14328(.dina(n14576),.dinb(n14481),.dout(n14577),.clk(gclk));
	jor g14329(.dina(n14577),.dinb(w_asqrt38_21[0]),.dout(n14578),.clk(gclk));
	jnot g14330(.din(w_n14242_0[1]),.dout(n14579),.clk(gclk));
	jand g14331(.dina(n14579),.dinb(n14578),.dout(n14580),.clk(gclk));
	jor g14332(.dina(n14580),.dinb(n14480),.dout(n14581),.clk(gclk));
	jor g14333(.dina(n14581),.dinb(w_asqrt39_17[2]),.dout(n14582),.clk(gclk));
	jnot g14334(.din(w_n14249_0[1]),.dout(n14583),.clk(gclk));
	jand g14335(.dina(n14583),.dinb(n14582),.dout(n14584),.clk(gclk));
	jor g14336(.dina(n14584),.dinb(n14479),.dout(n14585),.clk(gclk));
	jor g14337(.dina(n14585),.dinb(w_asqrt40_21[0]),.dout(n14586),.clk(gclk));
	jand g14338(.dina(w_n14256_0[1]),.dinb(n14586),.dout(n14587),.clk(gclk));
	jor g14339(.dina(n14587),.dinb(n14478),.dout(n14588),.clk(gclk));
	jor g14340(.dina(n14588),.dinb(w_asqrt41_18[0]),.dout(n14589),.clk(gclk));
	jnot g14341(.din(w_n14264_0[1]),.dout(n14590),.clk(gclk));
	jand g14342(.dina(n14590),.dinb(n14589),.dout(n14591),.clk(gclk));
	jor g14343(.dina(n14591),.dinb(n14477),.dout(n14592),.clk(gclk));
	jor g14344(.dina(n14592),.dinb(w_asqrt42_21[1]),.dout(n14593),.clk(gclk));
	jnot g14345(.din(w_n14271_0[0]),.dout(n14594),.clk(gclk));
	jand g14346(.dina(w_n14594_0[1]),.dinb(n14593),.dout(n14595),.clk(gclk));
	jor g14347(.dina(n14595),.dinb(n14476),.dout(n14596),.clk(gclk));
	jor g14348(.dina(n14596),.dinb(w_asqrt43_18[1]),.dout(n14597),.clk(gclk));
	jnot g14349(.din(w_n14278_0[1]),.dout(n14598),.clk(gclk));
	jand g14350(.dina(n14598),.dinb(n14597),.dout(n14599),.clk(gclk));
	jor g14351(.dina(n14599),.dinb(n14475),.dout(n14600),.clk(gclk));
	jor g14352(.dina(n14600),.dinb(w_asqrt44_21[1]),.dout(n14601),.clk(gclk));
	jnot g14353(.din(w_n14285_0[1]),.dout(n14602),.clk(gclk));
	jand g14354(.dina(n14602),.dinb(n14601),.dout(n14603),.clk(gclk));
	jor g14355(.dina(n14603),.dinb(n14474),.dout(n14604),.clk(gclk));
	jor g14356(.dina(n14604),.dinb(w_asqrt45_19[0]),.dout(n14605),.clk(gclk));
	jand g14357(.dina(w_n14292_0[1]),.dinb(n14605),.dout(n14606),.clk(gclk));
	jor g14358(.dina(n14606),.dinb(n14473),.dout(n14607),.clk(gclk));
	jor g14359(.dina(n14607),.dinb(w_asqrt46_21[1]),.dout(n14608),.clk(gclk));
	jand g14360(.dina(n14608),.dinb(w_n14299_0[1]),.dout(n14609),.clk(gclk));
	jor g14361(.dina(n14609),.dinb(n14472),.dout(n14610),.clk(gclk));
	jor g14362(.dina(n14610),.dinb(w_asqrt47_19[2]),.dout(n14611),.clk(gclk));
	jnot g14363(.din(w_n14308_0[1]),.dout(n14612),.clk(gclk));
	jand g14364(.dina(n14612),.dinb(n14611),.dout(n14613),.clk(gclk));
	jor g14365(.dina(n14613),.dinb(n14471),.dout(n14614),.clk(gclk));
	jor g14366(.dina(n14614),.dinb(w_asqrt48_21[2]),.dout(n14615),.clk(gclk));
	jand g14367(.dina(w_n14315_0[1]),.dinb(n14615),.dout(n14616),.clk(gclk));
	jor g14368(.dina(n14616),.dinb(n14470),.dout(n14617),.clk(gclk));
	jor g14369(.dina(n14617),.dinb(w_asqrt49_20[0]),.dout(n14618),.clk(gclk));
	jnot g14370(.din(w_n14323_0[1]),.dout(n14619),.clk(gclk));
	jand g14371(.dina(n14619),.dinb(n14618),.dout(n14620),.clk(gclk));
	jor g14372(.dina(n14620),.dinb(n14469),.dout(n14621),.clk(gclk));
	jor g14373(.dina(n14621),.dinb(w_asqrt50_22[0]),.dout(n14622),.clk(gclk));
	jand g14374(.dina(w_n14330_0[1]),.dinb(n14622),.dout(n14623),.clk(gclk));
	jor g14375(.dina(n14623),.dinb(n14468),.dout(n14624),.clk(gclk));
	jor g14376(.dina(n14624),.dinb(w_asqrt51_20[1]),.dout(n14625),.clk(gclk));
	jnot g14377(.din(w_n14338_0[1]),.dout(n14626),.clk(gclk));
	jand g14378(.dina(n14626),.dinb(n14625),.dout(n14627),.clk(gclk));
	jor g14379(.dina(n14627),.dinb(n14467),.dout(n14628),.clk(gclk));
	jor g14380(.dina(n14628),.dinb(w_asqrt52_22[0]),.dout(n14629),.clk(gclk));
	jnot g14381(.din(w_n14345_0[1]),.dout(n14630),.clk(gclk));
	jand g14382(.dina(n14630),.dinb(n14629),.dout(n14631),.clk(gclk));
	jor g14383(.dina(n14631),.dinb(n14466),.dout(n14632),.clk(gclk));
	jor g14384(.dina(n14632),.dinb(w_asqrt53_21[0]),.dout(n14633),.clk(gclk));
	jnot g14385(.din(w_n14352_0[1]),.dout(n14634),.clk(gclk));
	jand g14386(.dina(n14634),.dinb(n14633),.dout(n14635),.clk(gclk));
	jor g14387(.dina(n14635),.dinb(n14465),.dout(n14636),.clk(gclk));
	jor g14388(.dina(n14636),.dinb(w_asqrt54_22[0]),.dout(n14637),.clk(gclk));
	jand g14389(.dina(w_n14359_0[1]),.dinb(n14637),.dout(n14638),.clk(gclk));
	jor g14390(.dina(n14638),.dinb(n14464),.dout(n14639),.clk(gclk));
	jor g14391(.dina(n14639),.dinb(w_asqrt55_21[1]),.dout(n14640),.clk(gclk));
	jnot g14392(.din(w_n14367_0[1]),.dout(n14641),.clk(gclk));
	jand g14393(.dina(n14641),.dinb(n14640),.dout(n14642),.clk(gclk));
	jor g14394(.dina(n14642),.dinb(n14463),.dout(n14643),.clk(gclk));
	jor g14395(.dina(n14643),.dinb(w_asqrt56_22[1]),.dout(n14644),.clk(gclk));
	jand g14396(.dina(w_n14374_0[1]),.dinb(n14644),.dout(n14645),.clk(gclk));
	jor g14397(.dina(n14645),.dinb(n14462),.dout(n14646),.clk(gclk));
	jor g14398(.dina(n14646),.dinb(w_asqrt57_22[0]),.dout(n14647),.clk(gclk));
	jnot g14399(.din(w_n14382_0[1]),.dout(n14648),.clk(gclk));
	jand g14400(.dina(n14648),.dinb(n14647),.dout(n14649),.clk(gclk));
	jor g14401(.dina(n14649),.dinb(n14461),.dout(n14650),.clk(gclk));
	jor g14402(.dina(n14650),.dinb(w_asqrt58_22[2]),.dout(n14651),.clk(gclk));
	jand g14403(.dina(w_n14389_0[1]),.dinb(n14651),.dout(n14652),.clk(gclk));
	jor g14404(.dina(n14652),.dinb(n14460),.dout(n14653),.clk(gclk));
	jor g14405(.dina(n14653),.dinb(w_asqrt59_22[1]),.dout(n14654),.clk(gclk));
	jnot g14406(.din(w_n14397_0[1]),.dout(n14655),.clk(gclk));
	jand g14407(.dina(n14655),.dinb(n14654),.dout(n14656),.clk(gclk));
	jor g14408(.dina(n14656),.dinb(n14459),.dout(n14657),.clk(gclk));
	jor g14409(.dina(n14657),.dinb(w_asqrt60_22[2]),.dout(n14658),.clk(gclk));
	jand g14410(.dina(w_n14404_0[1]),.dinb(n14658),.dout(n14659),.clk(gclk));
	jor g14411(.dina(n14659),.dinb(n14458),.dout(n14660),.clk(gclk));
	jor g14412(.dina(n14660),.dinb(w_asqrt61_22[2]),.dout(n14661),.clk(gclk));
	jand g14413(.dina(w_n14412_0[1]),.dinb(n14661),.dout(n14662),.clk(gclk));
	jor g14414(.dina(n14662),.dinb(n14457),.dout(n14663),.clk(gclk));
	jor g14415(.dina(n14663),.dinb(w_asqrt62_22[2]),.dout(n14664),.clk(gclk));
	jand g14416(.dina(w_n14420_0[0]),.dinb(n14664),.dout(n14665),.clk(gclk));
	jor g14417(.dina(n14665),.dinb(n14456),.dout(n14666),.clk(gclk));
	jnot g14418(.din(w_n14426_1[0]),.dout(n14667),.clk(gclk));
	jand g14419(.dina(n14667),.dinb(n14666),.dout(n14668),.clk(gclk));
	jnot g14420(.din(w_n14432_0[0]),.dout(n14669),.clk(gclk));
	jand g14421(.dina(n14669),.dinb(n14668),.dout(n14670),.clk(gclk));
	jor g14422(.dina(n14670),.dinb(w_asqrt63_28[1]),.dout(n14671),.clk(gclk));
	jand g14423(.dina(w_n14438_0[0]),.dinb(w_n14671_0[1]),.dout(n14672),.clk(gclk));
	jand g14424(.dina(w_n14672_0[1]),.dinb(w_n14454_0[1]),.dout(n14674),.clk(gclk));
	jor g14425(.dina(w_n14674_20[1]),.dinb(n14453),.dout(n14675),.clk(gclk));
	jand g14426(.dina(n14675),.dinb(n14452),.dout(n14676),.clk(gclk));
	jand g14427(.dina(n14676),.dinb(n14450),.dout(n14677),.clk(gclk));
	jor g14428(.dina(n14677),.dinb(w_n14449_0[1]),.dout(n14678),.clk(gclk));
	jand g14429(.dina(w_n14678_0[2]),.dinb(w_asqrt18_19[0]),.dout(n14679),.clk(gclk));
	jor g14430(.dina(w_n14678_0[1]),.dinb(w_asqrt18_18[2]),.dout(n14680),.clk(gclk));
	jand g14431(.dina(w_asqrt16_33[2]),.dinb(w_n14082_0[0]),.dout(n14681),.clk(gclk));
	jand g14432(.dina(w_n14437_0[0]),.dinb(w_n14454_0[0]),.dout(n14682),.clk(gclk));
	jand g14433(.dina(n14682),.dinb(w_n14671_0[0]),.dout(n14683),.clk(gclk));
	jand g14434(.dina(n14683),.dinb(w_asqrt17_11[1]),.dout(n14684),.clk(gclk));
	jor g14435(.dina(n14684),.dinb(w_n14681_0[1]),.dout(n14685),.clk(gclk));
	jxor g14436(.dina(n14685),.dinb(w_a34_0[1]),.dout(n14686),.clk(gclk));
	jnot g14437(.din(w_n14686_0[1]),.dout(n14687),.clk(gclk));
	jand g14438(.dina(w_n14687_0[1]),.dinb(n14680),.dout(n14688),.clk(gclk));
	jor g14439(.dina(n14688),.dinb(w_n14679_0[1]),.dout(n14689),.clk(gclk));
	jand g14440(.dina(w_n14689_0[2]),.dinb(w_asqrt19_12[0]),.dout(n14690),.clk(gclk));
	jor g14441(.dina(w_n14689_0[1]),.dinb(w_asqrt19_11[2]),.dout(n14691),.clk(gclk));
	jxor g14442(.dina(w_n14085_0[0]),.dinb(w_n13515_20[2]),.dout(n14692),.clk(gclk));
	jand g14443(.dina(n14692),.dinb(w_asqrt16_33[1]),.dout(n14693),.clk(gclk));
	jxor g14444(.dina(n14693),.dinb(w_n14506_0[0]),.dout(n14694),.clk(gclk));
	jand g14445(.dina(w_n14694_0[1]),.dinb(n14691),.dout(n14695),.clk(gclk));
	jor g14446(.dina(n14695),.dinb(w_n14690_0[1]),.dout(n14696),.clk(gclk));
	jand g14447(.dina(w_n14696_0[2]),.dinb(w_asqrt20_19[0]),.dout(n14697),.clk(gclk));
	jor g14448(.dina(w_n14696_0[1]),.dinb(w_asqrt20_18[2]),.dout(n14698),.clk(gclk));
	jxor g14449(.dina(w_n14093_0[0]),.dinb(w_n12947_27[2]),.dout(n14699),.clk(gclk));
	jand g14450(.dina(n14699),.dinb(w_asqrt16_33[0]),.dout(n14700),.clk(gclk));
	jxor g14451(.dina(n14700),.dinb(w_n14102_0[0]),.dout(n14701),.clk(gclk));
	jnot g14452(.din(w_n14701_0[1]),.dout(n14702),.clk(gclk));
	jand g14453(.dina(w_n14702_0[1]),.dinb(n14698),.dout(n14703),.clk(gclk));
	jor g14454(.dina(n14703),.dinb(w_n14697_0[1]),.dout(n14704),.clk(gclk));
	jand g14455(.dina(w_n14704_0[2]),.dinb(w_asqrt21_12[2]),.dout(n14705),.clk(gclk));
	jor g14456(.dina(w_n14704_0[1]),.dinb(w_asqrt21_12[1]),.dout(n14706),.clk(gclk));
	jxor g14457(.dina(w_n14104_0[0]),.dinb(w_n12410_21[1]),.dout(n14707),.clk(gclk));
	jand g14458(.dina(n14707),.dinb(w_asqrt16_32[2]),.dout(n14708),.clk(gclk));
	jxor g14459(.dina(n14708),.dinb(w_n14109_0[0]),.dout(n14709),.clk(gclk));
	jand g14460(.dina(w_n14709_0[1]),.dinb(n14706),.dout(n14710),.clk(gclk));
	jor g14461(.dina(n14710),.dinb(w_n14705_0[1]),.dout(n14711),.clk(gclk));
	jand g14462(.dina(w_n14711_0[2]),.dinb(w_asqrt22_19[1]),.dout(n14712),.clk(gclk));
	jor g14463(.dina(w_n14711_0[1]),.dinb(w_asqrt22_19[0]),.dout(n14713),.clk(gclk));
	jxor g14464(.dina(w_n14112_0[0]),.dinb(w_n11858_28[0]),.dout(n14714),.clk(gclk));
	jand g14465(.dina(n14714),.dinb(w_asqrt16_32[1]),.dout(n14715),.clk(gclk));
	jxor g14466(.dina(n14715),.dinb(w_n14117_0[0]),.dout(n14716),.clk(gclk));
	jnot g14467(.din(w_n14716_0[1]),.dout(n14717),.clk(gclk));
	jand g14468(.dina(w_n14717_0[1]),.dinb(n14713),.dout(n14718),.clk(gclk));
	jor g14469(.dina(n14718),.dinb(w_n14712_0[1]),.dout(n14719),.clk(gclk));
	jand g14470(.dina(w_n14719_0[2]),.dinb(w_asqrt23_13[1]),.dout(n14720),.clk(gclk));
	jor g14471(.dina(w_n14719_0[1]),.dinb(w_asqrt23_13[0]),.dout(n14721),.clk(gclk));
	jxor g14472(.dina(w_n14119_0[0]),.dinb(w_n11347_22[0]),.dout(n14722),.clk(gclk));
	jand g14473(.dina(n14722),.dinb(w_asqrt16_32[0]),.dout(n14723),.clk(gclk));
	jxor g14474(.dina(n14723),.dinb(w_n14124_0[0]),.dout(n14724),.clk(gclk));
	jnot g14475(.din(w_n14724_0[1]),.dout(n14725),.clk(gclk));
	jand g14476(.dina(w_n14725_0[1]),.dinb(n14721),.dout(n14726),.clk(gclk));
	jor g14477(.dina(n14726),.dinb(w_n14720_0[1]),.dout(n14727),.clk(gclk));
	jand g14478(.dina(w_n14727_0[2]),.dinb(w_asqrt24_19[1]),.dout(n14728),.clk(gclk));
	jor g14479(.dina(w_n14727_0[1]),.dinb(w_asqrt24_19[0]),.dout(n14729),.clk(gclk));
	jxor g14480(.dina(w_n14126_0[0]),.dinb(w_n10824_28[2]),.dout(n14730),.clk(gclk));
	jand g14481(.dina(n14730),.dinb(w_asqrt16_31[2]),.dout(n14731),.clk(gclk));
	jxor g14482(.dina(n14731),.dinb(w_n14131_0[0]),.dout(n14732),.clk(gclk));
	jnot g14483(.din(w_n14732_0[1]),.dout(n14733),.clk(gclk));
	jand g14484(.dina(w_n14733_0[1]),.dinb(n14729),.dout(n14734),.clk(gclk));
	jor g14485(.dina(n14734),.dinb(w_n14728_0[1]),.dout(n14735),.clk(gclk));
	jand g14486(.dina(w_n14735_0[2]),.dinb(w_asqrt25_13[1]),.dout(n14736),.clk(gclk));
	jor g14487(.dina(w_n14735_0[1]),.dinb(w_asqrt25_13[0]),.dout(n14737),.clk(gclk));
	jxor g14488(.dina(w_n14133_0[0]),.dinb(w_n10328_23[0]),.dout(n14738),.clk(gclk));
	jand g14489(.dina(n14738),.dinb(w_asqrt16_31[1]),.dout(n14739),.clk(gclk));
	jxor g14490(.dina(n14739),.dinb(w_n14138_0[0]),.dout(n14740),.clk(gclk));
	jand g14491(.dina(w_n14740_0[1]),.dinb(n14737),.dout(n14741),.clk(gclk));
	jor g14492(.dina(n14741),.dinb(w_n14736_0[1]),.dout(n14742),.clk(gclk));
	jand g14493(.dina(w_n14742_0[2]),.dinb(w_asqrt26_19[1]),.dout(n14743),.clk(gclk));
	jor g14494(.dina(w_n14742_0[1]),.dinb(w_asqrt26_19[0]),.dout(n14744),.clk(gclk));
	jxor g14495(.dina(w_n14141_0[0]),.dinb(w_n9832_29[1]),.dout(n14745),.clk(gclk));
	jand g14496(.dina(n14745),.dinb(w_asqrt16_31[0]),.dout(n14746),.clk(gclk));
	jxor g14497(.dina(n14746),.dinb(w_n14146_0[0]),.dout(n14747),.clk(gclk));
	jnot g14498(.din(w_n14747_0[1]),.dout(n14748),.clk(gclk));
	jand g14499(.dina(w_n14748_0[1]),.dinb(n14744),.dout(n14749),.clk(gclk));
	jor g14500(.dina(n14749),.dinb(w_n14743_0[1]),.dout(n14750),.clk(gclk));
	jand g14501(.dina(w_n14750_0[2]),.dinb(w_asqrt27_14[0]),.dout(n14751),.clk(gclk));
	jor g14502(.dina(w_n14750_0[1]),.dinb(w_asqrt27_13[2]),.dout(n14752),.clk(gclk));
	jxor g14503(.dina(w_n14148_0[0]),.dinb(w_n9369_24[0]),.dout(n14753),.clk(gclk));
	jand g14504(.dina(n14753),.dinb(w_asqrt16_30[2]),.dout(n14754),.clk(gclk));
	jxor g14505(.dina(n14754),.dinb(w_n14153_0[0]),.dout(n14755),.clk(gclk));
	jand g14506(.dina(w_n14755_0[1]),.dinb(n14752),.dout(n14756),.clk(gclk));
	jor g14507(.dina(n14756),.dinb(w_n14751_0[1]),.dout(n14757),.clk(gclk));
	jand g14508(.dina(w_n14757_0[2]),.dinb(w_asqrt28_19[2]),.dout(n14758),.clk(gclk));
	jor g14509(.dina(w_n14757_0[1]),.dinb(w_asqrt28_19[1]),.dout(n14759),.clk(gclk));
	jxor g14510(.dina(w_n14156_0[0]),.dinb(w_n8890_29[2]),.dout(n14760),.clk(gclk));
	jand g14511(.dina(n14760),.dinb(w_asqrt16_30[1]),.dout(n14761),.clk(gclk));
	jxor g14512(.dina(n14761),.dinb(w_n14161_0[0]),.dout(n14762),.clk(gclk));
	jnot g14513(.din(w_n14762_0[1]),.dout(n14763),.clk(gclk));
	jand g14514(.dina(w_n14763_0[1]),.dinb(n14759),.dout(n14764),.clk(gclk));
	jor g14515(.dina(n14764),.dinb(w_n14758_0[1]),.dout(n14765),.clk(gclk));
	jand g14516(.dina(w_n14765_0[2]),.dinb(w_asqrt29_14[1]),.dout(n14766),.clk(gclk));
	jor g14517(.dina(w_n14765_0[1]),.dinb(w_asqrt29_14[0]),.dout(n14767),.clk(gclk));
	jxor g14518(.dina(w_n14163_0[0]),.dinb(w_n8449_24[2]),.dout(n14768),.clk(gclk));
	jand g14519(.dina(n14768),.dinb(w_asqrt16_30[0]),.dout(n14769),.clk(gclk));
	jxor g14520(.dina(n14769),.dinb(w_n14168_0[0]),.dout(n14770),.clk(gclk));
	jand g14521(.dina(w_n14770_0[1]),.dinb(n14767),.dout(n14771),.clk(gclk));
	jor g14522(.dina(n14771),.dinb(w_n14766_0[1]),.dout(n14772),.clk(gclk));
	jand g14523(.dina(w_n14772_0[2]),.dinb(w_asqrt30_20[0]),.dout(n14773),.clk(gclk));
	jor g14524(.dina(w_n14772_0[1]),.dinb(w_asqrt30_19[2]),.dout(n14774),.clk(gclk));
	jxor g14525(.dina(w_n14171_0[0]),.dinb(w_n8003_30[1]),.dout(n14775),.clk(gclk));
	jand g14526(.dina(n14775),.dinb(w_asqrt16_29[2]),.dout(n14776),.clk(gclk));
	jxor g14527(.dina(n14776),.dinb(w_n14176_0[0]),.dout(n14777),.clk(gclk));
	jnot g14528(.din(w_n14777_0[1]),.dout(n14778),.clk(gclk));
	jand g14529(.dina(w_n14778_0[1]),.dinb(n14774),.dout(n14779),.clk(gclk));
	jor g14530(.dina(n14779),.dinb(w_n14773_0[1]),.dout(n14780),.clk(gclk));
	jand g14531(.dina(w_n14780_0[2]),.dinb(w_asqrt31_15[0]),.dout(n14781),.clk(gclk));
	jor g14532(.dina(w_n14780_0[1]),.dinb(w_asqrt31_14[2]),.dout(n14782),.clk(gclk));
	jxor g14533(.dina(w_n14178_0[0]),.dinb(w_n7581_25[2]),.dout(n14783),.clk(gclk));
	jand g14534(.dina(n14783),.dinb(w_asqrt16_29[1]),.dout(n14784),.clk(gclk));
	jxor g14535(.dina(n14784),.dinb(w_n14183_0[0]),.dout(n14785),.clk(gclk));
	jand g14536(.dina(w_n14785_0[1]),.dinb(n14782),.dout(n14786),.clk(gclk));
	jor g14537(.dina(n14786),.dinb(w_n14781_0[1]),.dout(n14787),.clk(gclk));
	jand g14538(.dina(w_n14787_0[2]),.dinb(w_asqrt32_20[0]),.dout(n14788),.clk(gclk));
	jor g14539(.dina(w_n14787_0[1]),.dinb(w_asqrt32_19[2]),.dout(n14789),.clk(gclk));
	jxor g14540(.dina(w_n14186_0[0]),.dinb(w_n7154_30[2]),.dout(n14790),.clk(gclk));
	jand g14541(.dina(n14790),.dinb(w_asqrt16_29[0]),.dout(n14791),.clk(gclk));
	jxor g14542(.dina(n14791),.dinb(w_n14191_0[0]),.dout(n14792),.clk(gclk));
	jnot g14543(.din(w_n14792_0[1]),.dout(n14793),.clk(gclk));
	jand g14544(.dina(w_n14793_0[1]),.dinb(n14789),.dout(n14794),.clk(gclk));
	jor g14545(.dina(n14794),.dinb(w_n14788_0[1]),.dout(n14795),.clk(gclk));
	jand g14546(.dina(w_n14795_0[2]),.dinb(w_asqrt33_15[2]),.dout(n14796),.clk(gclk));
	jor g14547(.dina(w_n14795_0[1]),.dinb(w_asqrt33_15[1]),.dout(n14797),.clk(gclk));
	jxor g14548(.dina(w_n14193_0[0]),.dinb(w_n6758_26[1]),.dout(n14798),.clk(gclk));
	jand g14549(.dina(n14798),.dinb(w_asqrt16_28[2]),.dout(n14799),.clk(gclk));
	jxor g14550(.dina(n14799),.dinb(w_n14198_0[0]),.dout(n14800),.clk(gclk));
	jnot g14551(.din(w_n14800_0[1]),.dout(n14801),.clk(gclk));
	jand g14552(.dina(w_n14801_0[1]),.dinb(n14797),.dout(n14802),.clk(gclk));
	jor g14553(.dina(n14802),.dinb(w_n14796_0[1]),.dout(n14803),.clk(gclk));
	jand g14554(.dina(w_n14803_0[2]),.dinb(w_asqrt34_20[1]),.dout(n14804),.clk(gclk));
	jor g14555(.dina(w_n14803_0[1]),.dinb(w_asqrt34_20[0]),.dout(n14805),.clk(gclk));
	jxor g14556(.dina(w_n14200_0[0]),.dinb(w_n6357_31[0]),.dout(n14806),.clk(gclk));
	jand g14557(.dina(n14806),.dinb(w_asqrt16_28[1]),.dout(n14807),.clk(gclk));
	jxor g14558(.dina(n14807),.dinb(w_n14205_0[0]),.dout(n14808),.clk(gclk));
	jnot g14559(.din(w_n14808_0[1]),.dout(n14809),.clk(gclk));
	jand g14560(.dina(w_n14809_0[1]),.dinb(n14805),.dout(n14810),.clk(gclk));
	jor g14561(.dina(n14810),.dinb(w_n14804_0[1]),.dout(n14811),.clk(gclk));
	jand g14562(.dina(w_n14811_0[2]),.dinb(w_asqrt35_16[1]),.dout(n14812),.clk(gclk));
	jor g14563(.dina(w_n14811_0[1]),.dinb(w_asqrt35_16[0]),.dout(n14813),.clk(gclk));
	jxor g14564(.dina(w_n14207_0[0]),.dinb(w_n5989_27[0]),.dout(n14814),.clk(gclk));
	jand g14565(.dina(n14814),.dinb(w_asqrt16_28[0]),.dout(n14815),.clk(gclk));
	jxor g14566(.dina(n14815),.dinb(w_n14212_0[0]),.dout(n14816),.clk(gclk));
	jand g14567(.dina(w_n14816_0[1]),.dinb(n14813),.dout(n14817),.clk(gclk));
	jor g14568(.dina(n14817),.dinb(w_n14812_0[1]),.dout(n14818),.clk(gclk));
	jand g14569(.dina(w_n14818_0[2]),.dinb(w_asqrt36_20[1]),.dout(n14819),.clk(gclk));
	jor g14570(.dina(w_n14818_0[1]),.dinb(w_asqrt36_20[0]),.dout(n14820),.clk(gclk));
	jxor g14571(.dina(w_n14215_0[0]),.dinb(w_n5606_31[1]),.dout(n14821),.clk(gclk));
	jand g14572(.dina(n14821),.dinb(w_asqrt16_27[2]),.dout(n14822),.clk(gclk));
	jxor g14573(.dina(n14822),.dinb(w_n14220_0[0]),.dout(n14823),.clk(gclk));
	jnot g14574(.din(w_n14823_0[1]),.dout(n14824),.clk(gclk));
	jand g14575(.dina(w_n14824_0[1]),.dinb(n14820),.dout(n14825),.clk(gclk));
	jor g14576(.dina(n14825),.dinb(w_n14819_0[1]),.dout(n14826),.clk(gclk));
	jand g14577(.dina(w_n14826_0[2]),.dinb(w_asqrt37_16[2]),.dout(n14827),.clk(gclk));
	jor g14578(.dina(w_n14826_0[1]),.dinb(w_asqrt37_16[1]),.dout(n14828),.clk(gclk));
	jxor g14579(.dina(w_n14222_0[0]),.dinb(w_n5259_28[0]),.dout(n14829),.clk(gclk));
	jand g14580(.dina(n14829),.dinb(w_asqrt16_27[1]),.dout(n14830),.clk(gclk));
	jxor g14581(.dina(n14830),.dinb(w_n14227_0[0]),.dout(n14831),.clk(gclk));
	jand g14582(.dina(w_n14831_0[1]),.dinb(n14828),.dout(n14832),.clk(gclk));
	jor g14583(.dina(n14832),.dinb(w_n14827_0[1]),.dout(n14833),.clk(gclk));
	jand g14584(.dina(w_n14833_0[2]),.dinb(w_asqrt38_20[2]),.dout(n14834),.clk(gclk));
	jor g14585(.dina(w_n14833_0[1]),.dinb(w_asqrt38_20[1]),.dout(n14835),.clk(gclk));
	jxor g14586(.dina(w_n14230_0[0]),.dinb(w_n4902_32[0]),.dout(n14836),.clk(gclk));
	jand g14587(.dina(n14836),.dinb(w_asqrt16_27[0]),.dout(n14837),.clk(gclk));
	jxor g14588(.dina(n14837),.dinb(w_n14235_0[0]),.dout(n14838),.clk(gclk));
	jnot g14589(.din(w_n14838_0[1]),.dout(n14839),.clk(gclk));
	jand g14590(.dina(w_n14839_0[1]),.dinb(n14835),.dout(n14840),.clk(gclk));
	jor g14591(.dina(n14840),.dinb(w_n14834_0[1]),.dout(n14841),.clk(gclk));
	jand g14592(.dina(w_n14841_0[2]),.dinb(w_asqrt39_17[1]),.dout(n14842),.clk(gclk));
	jor g14593(.dina(w_n14841_0[1]),.dinb(w_asqrt39_17[0]),.dout(n14843),.clk(gclk));
	jxor g14594(.dina(w_n14237_0[0]),.dinb(w_n4582_29[0]),.dout(n14844),.clk(gclk));
	jand g14595(.dina(n14844),.dinb(w_asqrt16_26[2]),.dout(n14845),.clk(gclk));
	jxor g14596(.dina(n14845),.dinb(w_n14242_0[0]),.dout(n14846),.clk(gclk));
	jnot g14597(.din(w_n14846_0[1]),.dout(n14847),.clk(gclk));
	jand g14598(.dina(w_n14847_0[1]),.dinb(n14843),.dout(n14848),.clk(gclk));
	jor g14599(.dina(n14848),.dinb(w_n14842_0[1]),.dout(n14849),.clk(gclk));
	jand g14600(.dina(w_n14849_0[2]),.dinb(w_asqrt40_20[2]),.dout(n14850),.clk(gclk));
	jor g14601(.dina(w_n14849_0[1]),.dinb(w_asqrt40_20[1]),.dout(n14851),.clk(gclk));
	jxor g14602(.dina(w_n14244_0[0]),.dinb(w_n4249_32[2]),.dout(n14852),.clk(gclk));
	jand g14603(.dina(n14852),.dinb(w_asqrt16_26[1]),.dout(n14853),.clk(gclk));
	jxor g14604(.dina(n14853),.dinb(w_n14249_0[0]),.dout(n14854),.clk(gclk));
	jnot g14605(.din(w_n14854_0[1]),.dout(n14855),.clk(gclk));
	jand g14606(.dina(w_n14855_0[1]),.dinb(n14851),.dout(n14856),.clk(gclk));
	jor g14607(.dina(n14856),.dinb(w_n14850_0[1]),.dout(n14857),.clk(gclk));
	jand g14608(.dina(w_n14857_0[2]),.dinb(w_asqrt41_17[2]),.dout(n14858),.clk(gclk));
	jor g14609(.dina(w_n14857_0[1]),.dinb(w_asqrt41_17[1]),.dout(n14859),.clk(gclk));
	jxor g14610(.dina(w_n14251_0[0]),.dinb(w_n3955_29[2]),.dout(n14860),.clk(gclk));
	jand g14611(.dina(n14860),.dinb(w_asqrt16_26[0]),.dout(n14861),.clk(gclk));
	jxor g14612(.dina(n14861),.dinb(w_n14256_0[0]),.dout(n14862),.clk(gclk));
	jand g14613(.dina(w_n14862_0[1]),.dinb(n14859),.dout(n14863),.clk(gclk));
	jor g14614(.dina(n14863),.dinb(w_n14858_0[1]),.dout(n14864),.clk(gclk));
	jand g14615(.dina(w_n14864_0[2]),.dinb(w_asqrt42_21[0]),.dout(n14865),.clk(gclk));
	jor g14616(.dina(w_n14864_0[1]),.dinb(w_asqrt42_20[2]),.dout(n14866),.clk(gclk));
	jxor g14617(.dina(w_n14259_0[0]),.dinb(w_n3642_33[0]),.dout(n14867),.clk(gclk));
	jand g14618(.dina(n14867),.dinb(w_asqrt16_25[2]),.dout(n14868),.clk(gclk));
	jxor g14619(.dina(n14868),.dinb(w_n14264_0[0]),.dout(n14869),.clk(gclk));
	jnot g14620(.din(w_n14869_0[1]),.dout(n14870),.clk(gclk));
	jand g14621(.dina(w_n14870_0[1]),.dinb(n14866),.dout(n14871),.clk(gclk));
	jor g14622(.dina(n14871),.dinb(w_n14865_0[1]),.dout(n14872),.clk(gclk));
	jand g14623(.dina(w_n14872_0[2]),.dinb(w_asqrt43_18[0]),.dout(n14873),.clk(gclk));
	jor g14624(.dina(w_n14872_0[1]),.dinb(w_asqrt43_17[2]),.dout(n14874),.clk(gclk));
	jxor g14625(.dina(w_n14266_0[0]),.dinb(w_n3368_30[1]),.dout(n14875),.clk(gclk));
	jand g14626(.dina(n14875),.dinb(w_asqrt16_25[1]),.dout(n14876),.clk(gclk));
	jxor g14627(.dina(n14876),.dinb(w_n14594_0[0]),.dout(n14877),.clk(gclk));
	jand g14628(.dina(w_n14877_0[1]),.dinb(n14874),.dout(n14878),.clk(gclk));
	jor g14629(.dina(n14878),.dinb(w_n14873_0[1]),.dout(n14879),.clk(gclk));
	jand g14630(.dina(w_n14879_0[2]),.dinb(w_asqrt44_21[0]),.dout(n14880),.clk(gclk));
	jor g14631(.dina(w_n14879_0[1]),.dinb(w_asqrt44_20[2]),.dout(n14881),.clk(gclk));
	jxor g14632(.dina(w_n14273_0[0]),.dinb(w_n3089_33[2]),.dout(n14882),.clk(gclk));
	jand g14633(.dina(n14882),.dinb(w_asqrt16_25[0]),.dout(n14883),.clk(gclk));
	jxor g14634(.dina(n14883),.dinb(w_n14278_0[0]),.dout(n14884),.clk(gclk));
	jnot g14635(.din(w_n14884_0[1]),.dout(n14885),.clk(gclk));
	jand g14636(.dina(w_n14885_0[1]),.dinb(n14881),.dout(n14886),.clk(gclk));
	jor g14637(.dina(n14886),.dinb(w_n14880_0[1]),.dout(n14887),.clk(gclk));
	jand g14638(.dina(w_n14887_0[2]),.dinb(w_asqrt45_18[2]),.dout(n14888),.clk(gclk));
	jor g14639(.dina(w_n14887_0[1]),.dinb(w_asqrt45_18[1]),.dout(n14889),.clk(gclk));
	jxor g14640(.dina(w_n14280_0[0]),.dinb(w_n2833_31[1]),.dout(n14890),.clk(gclk));
	jand g14641(.dina(n14890),.dinb(w_asqrt16_24[2]),.dout(n14891),.clk(gclk));
	jxor g14642(.dina(n14891),.dinb(w_n14285_0[0]),.dout(n14892),.clk(gclk));
	jnot g14643(.din(w_n14892_0[1]),.dout(n14893),.clk(gclk));
	jand g14644(.dina(w_n14893_0[1]),.dinb(n14889),.dout(n14894),.clk(gclk));
	jor g14645(.dina(n14894),.dinb(w_n14888_0[1]),.dout(n14895),.clk(gclk));
	jand g14646(.dina(w_n14895_0[2]),.dinb(w_asqrt46_21[0]),.dout(n14896),.clk(gclk));
	jor g14647(.dina(w_n14895_0[1]),.dinb(w_asqrt46_20[2]),.dout(n14897),.clk(gclk));
	jxor g14648(.dina(w_n14287_0[0]),.dinb(w_n2572_34[0]),.dout(n14898),.clk(gclk));
	jand g14649(.dina(n14898),.dinb(w_asqrt16_24[1]),.dout(n14899),.clk(gclk));
	jxor g14650(.dina(n14899),.dinb(w_n14292_0[0]),.dout(n14900),.clk(gclk));
	jand g14651(.dina(w_n14900_0[1]),.dinb(n14897),.dout(n14901),.clk(gclk));
	jor g14652(.dina(n14901),.dinb(w_n14896_0[1]),.dout(n14902),.clk(gclk));
	jand g14653(.dina(w_n14902_0[2]),.dinb(w_asqrt47_19[1]),.dout(n14903),.clk(gclk));
	jxor g14654(.dina(w_n14295_0[0]),.dinb(w_n2345_32[0]),.dout(n14904),.clk(gclk));
	jand g14655(.dina(n14904),.dinb(w_asqrt16_24[0]),.dout(n14905),.clk(gclk));
	jxor g14656(.dina(n14905),.dinb(w_n14299_0[0]),.dout(n14906),.clk(gclk));
	jor g14657(.dina(w_n14902_0[1]),.dinb(w_asqrt47_19[0]),.dout(n14907),.clk(gclk));
	jand g14658(.dina(n14907),.dinb(w_n14906_0[1]),.dout(n14908),.clk(gclk));
	jor g14659(.dina(n14908),.dinb(w_n14903_0[1]),.dout(n14909),.clk(gclk));
	jand g14660(.dina(w_n14909_0[2]),.dinb(w_asqrt48_21[1]),.dout(n14910),.clk(gclk));
	jor g14661(.dina(w_n14909_0[1]),.dinb(w_asqrt48_21[0]),.dout(n14911),.clk(gclk));
	jxor g14662(.dina(w_n14303_0[0]),.dinb(w_n2108_34[2]),.dout(n14912),.clk(gclk));
	jand g14663(.dina(n14912),.dinb(w_asqrt16_23[2]),.dout(n14913),.clk(gclk));
	jxor g14664(.dina(n14913),.dinb(w_n14308_0[0]),.dout(n14914),.clk(gclk));
	jnot g14665(.din(w_n14914_0[1]),.dout(n14915),.clk(gclk));
	jand g14666(.dina(w_n14915_0[1]),.dinb(n14911),.dout(n14916),.clk(gclk));
	jor g14667(.dina(n14916),.dinb(w_n14910_0[1]),.dout(n14917),.clk(gclk));
	jand g14668(.dina(w_n14917_0[2]),.dinb(w_asqrt49_19[2]),.dout(n14918),.clk(gclk));
	jor g14669(.dina(w_n14917_0[1]),.dinb(w_asqrt49_19[1]),.dout(n14919),.clk(gclk));
	jxor g14670(.dina(w_n14310_0[0]),.dinb(w_n1912_33[0]),.dout(n14920),.clk(gclk));
	jand g14671(.dina(n14920),.dinb(w_asqrt16_23[1]),.dout(n14921),.clk(gclk));
	jxor g14672(.dina(n14921),.dinb(w_n14315_0[0]),.dout(n14922),.clk(gclk));
	jand g14673(.dina(w_n14922_0[1]),.dinb(n14919),.dout(n14923),.clk(gclk));
	jor g14674(.dina(n14923),.dinb(w_n14918_0[1]),.dout(n14924),.clk(gclk));
	jand g14675(.dina(w_n14924_0[2]),.dinb(w_asqrt50_21[2]),.dout(n14925),.clk(gclk));
	jor g14676(.dina(w_n14924_0[1]),.dinb(w_asqrt50_21[1]),.dout(n14926),.clk(gclk));
	jxor g14677(.dina(w_n14318_0[0]),.dinb(w_n1699_35[1]),.dout(n14927),.clk(gclk));
	jand g14678(.dina(n14927),.dinb(w_asqrt16_23[0]),.dout(n14928),.clk(gclk));
	jxor g14679(.dina(n14928),.dinb(w_n14323_0[0]),.dout(n14929),.clk(gclk));
	jnot g14680(.din(w_n14929_0[1]),.dout(n14930),.clk(gclk));
	jand g14681(.dina(w_n14930_0[1]),.dinb(n14926),.dout(n14931),.clk(gclk));
	jor g14682(.dina(n14931),.dinb(w_n14925_0[1]),.dout(n14932),.clk(gclk));
	jand g14683(.dina(w_n14932_0[2]),.dinb(w_asqrt51_20[0]),.dout(n14933),.clk(gclk));
	jor g14684(.dina(w_n14932_0[1]),.dinb(w_asqrt51_19[2]),.dout(n14934),.clk(gclk));
	jxor g14685(.dina(w_n14325_0[0]),.dinb(w_n1516_33[2]),.dout(n14935),.clk(gclk));
	jand g14686(.dina(n14935),.dinb(w_asqrt16_22[2]),.dout(n14936),.clk(gclk));
	jxor g14687(.dina(n14936),.dinb(w_n14330_0[0]),.dout(n14937),.clk(gclk));
	jand g14688(.dina(w_n14937_0[1]),.dinb(n14934),.dout(n14938),.clk(gclk));
	jor g14689(.dina(n14938),.dinb(w_n14933_0[1]),.dout(n14939),.clk(gclk));
	jand g14690(.dina(w_n14939_0[2]),.dinb(w_asqrt52_21[2]),.dout(n14940),.clk(gclk));
	jor g14691(.dina(w_n14939_0[1]),.dinb(w_asqrt52_21[1]),.dout(n14941),.clk(gclk));
	jxor g14692(.dina(w_n14333_0[0]),.dinb(w_n1332_35[1]),.dout(n14942),.clk(gclk));
	jand g14693(.dina(n14942),.dinb(w_asqrt16_22[1]),.dout(n14943),.clk(gclk));
	jxor g14694(.dina(n14943),.dinb(w_n14338_0[0]),.dout(n14944),.clk(gclk));
	jnot g14695(.din(w_n14944_0[1]),.dout(n14945),.clk(gclk));
	jand g14696(.dina(w_n14945_0[1]),.dinb(n14941),.dout(n14946),.clk(gclk));
	jor g14697(.dina(n14946),.dinb(w_n14940_0[1]),.dout(n14947),.clk(gclk));
	jand g14698(.dina(w_n14947_0[2]),.dinb(w_asqrt53_20[2]),.dout(n14948),.clk(gclk));
	jor g14699(.dina(w_n14947_0[1]),.dinb(w_asqrt53_20[1]),.dout(n14949),.clk(gclk));
	jxor g14700(.dina(w_n14340_0[0]),.dinb(w_n1173_34[1]),.dout(n14950),.clk(gclk));
	jand g14701(.dina(n14950),.dinb(w_asqrt16_22[0]),.dout(n14951),.clk(gclk));
	jxor g14702(.dina(n14951),.dinb(w_n14345_0[0]),.dout(n14952),.clk(gclk));
	jnot g14703(.din(w_n14952_0[1]),.dout(n14953),.clk(gclk));
	jand g14704(.dina(w_n14953_0[1]),.dinb(n14949),.dout(n14954),.clk(gclk));
	jor g14705(.dina(n14954),.dinb(w_n14948_0[1]),.dout(n14955),.clk(gclk));
	jand g14706(.dina(w_n14955_0[2]),.dinb(w_asqrt54_21[2]),.dout(n14956),.clk(gclk));
	jor g14707(.dina(w_n14955_0[1]),.dinb(w_asqrt54_21[1]),.dout(n14957),.clk(gclk));
	jxor g14708(.dina(w_n14347_0[0]),.dinb(w_n1008_36[1]),.dout(n14958),.clk(gclk));
	jand g14709(.dina(n14958),.dinb(w_asqrt16_21[2]),.dout(n14959),.clk(gclk));
	jxor g14710(.dina(n14959),.dinb(w_n14352_0[0]),.dout(n14960),.clk(gclk));
	jnot g14711(.din(w_n14960_0[1]),.dout(n14961),.clk(gclk));
	jand g14712(.dina(w_n14961_0[1]),.dinb(n14957),.dout(n14962),.clk(gclk));
	jor g14713(.dina(n14962),.dinb(w_n14956_0[1]),.dout(n14963),.clk(gclk));
	jand g14714(.dina(w_n14963_0[2]),.dinb(w_asqrt55_21[0]),.dout(n14964),.clk(gclk));
	jor g14715(.dina(w_n14963_0[1]),.dinb(w_asqrt55_20[2]),.dout(n14965),.clk(gclk));
	jxor g14716(.dina(w_n14354_0[0]),.dinb(w_n884_35[1]),.dout(n14966),.clk(gclk));
	jand g14717(.dina(n14966),.dinb(w_asqrt16_21[1]),.dout(n14967),.clk(gclk));
	jxor g14718(.dina(n14967),.dinb(w_n14359_0[0]),.dout(n14968),.clk(gclk));
	jand g14719(.dina(w_n14968_0[1]),.dinb(n14965),.dout(n14969),.clk(gclk));
	jor g14720(.dina(n14969),.dinb(w_n14964_0[1]),.dout(n14970),.clk(gclk));
	jand g14721(.dina(w_n14970_0[2]),.dinb(w_asqrt56_22[0]),.dout(n14971),.clk(gclk));
	jor g14722(.dina(w_n14970_0[1]),.dinb(w_asqrt56_21[2]),.dout(n14972),.clk(gclk));
	jxor g14723(.dina(w_n14362_0[0]),.dinb(w_n743_36[1]),.dout(n14973),.clk(gclk));
	jand g14724(.dina(n14973),.dinb(w_asqrt16_21[0]),.dout(n14974),.clk(gclk));
	jxor g14725(.dina(n14974),.dinb(w_n14367_0[0]),.dout(n14975),.clk(gclk));
	jnot g14726(.din(w_n14975_0[1]),.dout(n14976),.clk(gclk));
	jand g14727(.dina(w_n14976_0[1]),.dinb(n14972),.dout(n14977),.clk(gclk));
	jor g14728(.dina(n14977),.dinb(w_n14971_0[1]),.dout(n14978),.clk(gclk));
	jand g14729(.dina(w_n14978_0[2]),.dinb(w_asqrt57_21[2]),.dout(n14979),.clk(gclk));
	jor g14730(.dina(w_n14978_0[1]),.dinb(w_asqrt57_21[1]),.dout(n14980),.clk(gclk));
	jxor g14731(.dina(w_n14369_0[0]),.dinb(w_n635_36[1]),.dout(n14981),.clk(gclk));
	jand g14732(.dina(n14981),.dinb(w_asqrt16_20[2]),.dout(n14982),.clk(gclk));
	jxor g14733(.dina(n14982),.dinb(w_n14374_0[0]),.dout(n14983),.clk(gclk));
	jand g14734(.dina(w_n14983_0[1]),.dinb(n14980),.dout(n14984),.clk(gclk));
	jor g14735(.dina(n14984),.dinb(w_n14979_0[1]),.dout(n14985),.clk(gclk));
	jand g14736(.dina(w_n14985_0[2]),.dinb(w_asqrt58_22[1]),.dout(n14986),.clk(gclk));
	jor g14737(.dina(w_n14985_0[1]),.dinb(w_asqrt58_22[0]),.dout(n14987),.clk(gclk));
	jxor g14738(.dina(w_n14377_0[0]),.dinb(w_n515_37[1]),.dout(n14988),.clk(gclk));
	jand g14739(.dina(n14988),.dinb(w_asqrt16_20[1]),.dout(n14989),.clk(gclk));
	jxor g14740(.dina(n14989),.dinb(w_n14382_0[0]),.dout(n14990),.clk(gclk));
	jnot g14741(.din(w_n14990_0[1]),.dout(n14991),.clk(gclk));
	jand g14742(.dina(w_n14991_0[1]),.dinb(n14987),.dout(n14992),.clk(gclk));
	jor g14743(.dina(n14992),.dinb(w_n14986_0[1]),.dout(n14993),.clk(gclk));
	jand g14744(.dina(w_n14993_0[2]),.dinb(w_asqrt59_22[0]),.dout(n14994),.clk(gclk));
	jor g14745(.dina(w_n14993_0[1]),.dinb(w_asqrt59_21[2]),.dout(n14995),.clk(gclk));
	jxor g14746(.dina(w_n14384_0[0]),.dinb(w_n443_37[1]),.dout(n14996),.clk(gclk));
	jand g14747(.dina(n14996),.dinb(w_asqrt16_20[0]),.dout(n14997),.clk(gclk));
	jxor g14748(.dina(n14997),.dinb(w_n14389_0[0]),.dout(n14998),.clk(gclk));
	jand g14749(.dina(w_n14998_0[1]),.dinb(n14995),.dout(n14999),.clk(gclk));
	jor g14750(.dina(n14999),.dinb(w_n14994_0[1]),.dout(n15000),.clk(gclk));
	jand g14751(.dina(w_n15000_0[2]),.dinb(w_asqrt60_22[1]),.dout(n15001),.clk(gclk));
	jor g14752(.dina(w_n15000_0[1]),.dinb(w_asqrt60_22[0]),.dout(n15002),.clk(gclk));
	jxor g14753(.dina(w_n14392_0[0]),.dinb(w_n352_37[2]),.dout(n15003),.clk(gclk));
	jand g14754(.dina(n15003),.dinb(w_asqrt16_19[2]),.dout(n15004),.clk(gclk));
	jxor g14755(.dina(n15004),.dinb(w_n14397_0[0]),.dout(n15005),.clk(gclk));
	jnot g14756(.din(w_n15005_0[1]),.dout(n15006),.clk(gclk));
	jand g14757(.dina(w_n15006_0[1]),.dinb(n15002),.dout(n15007),.clk(gclk));
	jor g14758(.dina(n15007),.dinb(w_n15001_0[1]),.dout(n15008),.clk(gclk));
	jand g14759(.dina(w_n15008_0[2]),.dinb(w_asqrt61_22[1]),.dout(n15009),.clk(gclk));
	jor g14760(.dina(w_n15008_0[1]),.dinb(w_asqrt61_22[0]),.dout(n15010),.clk(gclk));
	jxor g14761(.dina(w_n14399_0[0]),.dinb(w_n294_38[0]),.dout(n15011),.clk(gclk));
	jand g14762(.dina(n15011),.dinb(w_asqrt16_19[1]),.dout(n15012),.clk(gclk));
	jxor g14763(.dina(n15012),.dinb(w_n14404_0[0]),.dout(n15013),.clk(gclk));
	jand g14764(.dina(w_n15013_0[1]),.dinb(n15010),.dout(n15014),.clk(gclk));
	jor g14765(.dina(n15014),.dinb(w_n15009_0[1]),.dout(n15015),.clk(gclk));
	jand g14766(.dina(w_n15015_0[2]),.dinb(w_asqrt62_22[1]),.dout(n15016),.clk(gclk));
	jnot g14767(.din(w_n15016_0[1]),.dout(n15017),.clk(gclk));
	jnot g14768(.din(w_n15009_0[0]),.dout(n15018),.clk(gclk));
	jnot g14769(.din(w_n15001_0[0]),.dout(n15019),.clk(gclk));
	jnot g14770(.din(w_n14994_0[0]),.dout(n15020),.clk(gclk));
	jnot g14771(.din(w_n14986_0[0]),.dout(n15021),.clk(gclk));
	jnot g14772(.din(w_n14979_0[0]),.dout(n15022),.clk(gclk));
	jnot g14773(.din(w_n14971_0[0]),.dout(n15023),.clk(gclk));
	jnot g14774(.din(w_n14964_0[0]),.dout(n15024),.clk(gclk));
	jnot g14775(.din(w_n14956_0[0]),.dout(n15025),.clk(gclk));
	jnot g14776(.din(w_n14948_0[0]),.dout(n15026),.clk(gclk));
	jnot g14777(.din(w_n14940_0[0]),.dout(n15027),.clk(gclk));
	jnot g14778(.din(w_n14933_0[0]),.dout(n15028),.clk(gclk));
	jnot g14779(.din(w_n14925_0[0]),.dout(n15029),.clk(gclk));
	jnot g14780(.din(w_n14918_0[0]),.dout(n15030),.clk(gclk));
	jnot g14781(.din(w_n14910_0[0]),.dout(n15031),.clk(gclk));
	jnot g14782(.din(w_n14903_0[0]),.dout(n15032),.clk(gclk));
	jnot g14783(.din(w_n14906_0[0]),.dout(n15033),.clk(gclk));
	jnot g14784(.din(w_n14896_0[0]),.dout(n15034),.clk(gclk));
	jnot g14785(.din(w_n14888_0[0]),.dout(n15035),.clk(gclk));
	jnot g14786(.din(w_n14880_0[0]),.dout(n15036),.clk(gclk));
	jnot g14787(.din(w_n14873_0[0]),.dout(n15037),.clk(gclk));
	jnot g14788(.din(w_n14865_0[0]),.dout(n15038),.clk(gclk));
	jnot g14789(.din(w_n14858_0[0]),.dout(n15039),.clk(gclk));
	jnot g14790(.din(w_n14850_0[0]),.dout(n15040),.clk(gclk));
	jnot g14791(.din(w_n14842_0[0]),.dout(n15041),.clk(gclk));
	jnot g14792(.din(w_n14834_0[0]),.dout(n15042),.clk(gclk));
	jnot g14793(.din(w_n14827_0[0]),.dout(n15043),.clk(gclk));
	jnot g14794(.din(w_n14819_0[0]),.dout(n15044),.clk(gclk));
	jnot g14795(.din(w_n14812_0[0]),.dout(n15045),.clk(gclk));
	jnot g14796(.din(w_n14804_0[0]),.dout(n15046),.clk(gclk));
	jnot g14797(.din(w_n14796_0[0]),.dout(n15047),.clk(gclk));
	jnot g14798(.din(w_n14788_0[0]),.dout(n15048),.clk(gclk));
	jnot g14799(.din(w_n14781_0[0]),.dout(n15049),.clk(gclk));
	jnot g14800(.din(w_n14773_0[0]),.dout(n15050),.clk(gclk));
	jnot g14801(.din(w_n14766_0[0]),.dout(n15051),.clk(gclk));
	jnot g14802(.din(w_n14758_0[0]),.dout(n15052),.clk(gclk));
	jnot g14803(.din(w_n14751_0[0]),.dout(n15053),.clk(gclk));
	jnot g14804(.din(w_n14743_0[0]),.dout(n15054),.clk(gclk));
	jnot g14805(.din(w_n14736_0[0]),.dout(n15055),.clk(gclk));
	jnot g14806(.din(w_n14728_0[0]),.dout(n15056),.clk(gclk));
	jnot g14807(.din(w_n14720_0[0]),.dout(n15057),.clk(gclk));
	jnot g14808(.din(w_n14712_0[0]),.dout(n15058),.clk(gclk));
	jnot g14809(.din(w_n14705_0[0]),.dout(n15059),.clk(gclk));
	jnot g14810(.din(w_n14697_0[0]),.dout(n15060),.clk(gclk));
	jnot g14811(.din(w_n14690_0[0]),.dout(n15061),.clk(gclk));
	jnot g14812(.din(w_n14679_0[0]),.dout(n15062),.clk(gclk));
	jnot g14813(.din(w_n14449_0[0]),.dout(n15063),.clk(gclk));
	jnot g14814(.din(w_n14446_0[0]),.dout(n15064),.clk(gclk));
	jor g14815(.dina(w_n14674_20[0]),.dinb(w_n14080_0[2]),.dout(n15065),.clk(gclk));
	jand g14816(.dina(n15065),.dinb(n15064),.dout(n15066),.clk(gclk));
	jand g14817(.dina(n15066),.dinb(w_n14078_26[2]),.dout(n15067),.clk(gclk));
	jor g14818(.dina(w_n14674_19[2]),.dinb(w_a32_0[0]),.dout(n15068),.clk(gclk));
	jand g14819(.dina(n15068),.dinb(w_a33_0[0]),.dout(n15069),.clk(gclk));
	jor g14820(.dina(w_n14681_0[0]),.dinb(n15069),.dout(n15070),.clk(gclk));
	jor g14821(.dina(w_n15070_0[1]),.dinb(n15067),.dout(n15071),.clk(gclk));
	jand g14822(.dina(n15071),.dinb(n15063),.dout(n15072),.clk(gclk));
	jand g14823(.dina(n15072),.dinb(w_n13515_20[1]),.dout(n15073),.clk(gclk));
	jor g14824(.dina(w_n14686_0[0]),.dinb(n15073),.dout(n15074),.clk(gclk));
	jand g14825(.dina(n15074),.dinb(n15062),.dout(n15075),.clk(gclk));
	jand g14826(.dina(n15075),.dinb(w_n12947_27[1]),.dout(n15076),.clk(gclk));
	jnot g14827(.din(w_n14694_0[0]),.dout(n15077),.clk(gclk));
	jor g14828(.dina(w_n15077_0[1]),.dinb(n15076),.dout(n15078),.clk(gclk));
	jand g14829(.dina(n15078),.dinb(n15061),.dout(n15079),.clk(gclk));
	jand g14830(.dina(n15079),.dinb(w_n12410_21[0]),.dout(n15080),.clk(gclk));
	jor g14831(.dina(w_n14701_0[0]),.dinb(n15080),.dout(n15081),.clk(gclk));
	jand g14832(.dina(n15081),.dinb(n15060),.dout(n15082),.clk(gclk));
	jand g14833(.dina(n15082),.dinb(w_n11858_27[2]),.dout(n15083),.clk(gclk));
	jnot g14834(.din(w_n14709_0[0]),.dout(n15084),.clk(gclk));
	jor g14835(.dina(w_n15084_0[1]),.dinb(n15083),.dout(n15085),.clk(gclk));
	jand g14836(.dina(n15085),.dinb(n15059),.dout(n15086),.clk(gclk));
	jand g14837(.dina(n15086),.dinb(w_n11347_21[2]),.dout(n15087),.clk(gclk));
	jor g14838(.dina(w_n14716_0[0]),.dinb(n15087),.dout(n15088),.clk(gclk));
	jand g14839(.dina(n15088),.dinb(n15058),.dout(n15089),.clk(gclk));
	jand g14840(.dina(n15089),.dinb(w_n10824_28[1]),.dout(n15090),.clk(gclk));
	jor g14841(.dina(w_n14724_0[0]),.dinb(n15090),.dout(n15091),.clk(gclk));
	jand g14842(.dina(n15091),.dinb(n15057),.dout(n15092),.clk(gclk));
	jand g14843(.dina(n15092),.dinb(w_n10328_22[2]),.dout(n15093),.clk(gclk));
	jor g14844(.dina(w_n14732_0[0]),.dinb(n15093),.dout(n15094),.clk(gclk));
	jand g14845(.dina(n15094),.dinb(n15056),.dout(n15095),.clk(gclk));
	jand g14846(.dina(n15095),.dinb(w_n9832_29[0]),.dout(n15096),.clk(gclk));
	jnot g14847(.din(w_n14740_0[0]),.dout(n15097),.clk(gclk));
	jor g14848(.dina(w_n15097_0[1]),.dinb(n15096),.dout(n15098),.clk(gclk));
	jand g14849(.dina(n15098),.dinb(n15055),.dout(n15099),.clk(gclk));
	jand g14850(.dina(n15099),.dinb(w_n9369_23[2]),.dout(n15100),.clk(gclk));
	jor g14851(.dina(w_n14747_0[0]),.dinb(n15100),.dout(n15101),.clk(gclk));
	jand g14852(.dina(n15101),.dinb(n15054),.dout(n15102),.clk(gclk));
	jand g14853(.dina(n15102),.dinb(w_n8890_29[1]),.dout(n15103),.clk(gclk));
	jnot g14854(.din(w_n14755_0[0]),.dout(n15104),.clk(gclk));
	jor g14855(.dina(w_n15104_0[1]),.dinb(n15103),.dout(n15105),.clk(gclk));
	jand g14856(.dina(n15105),.dinb(n15053),.dout(n15106),.clk(gclk));
	jand g14857(.dina(n15106),.dinb(w_n8449_24[1]),.dout(n15107),.clk(gclk));
	jor g14858(.dina(w_n14762_0[0]),.dinb(n15107),.dout(n15108),.clk(gclk));
	jand g14859(.dina(n15108),.dinb(n15052),.dout(n15109),.clk(gclk));
	jand g14860(.dina(n15109),.dinb(w_n8003_30[0]),.dout(n15110),.clk(gclk));
	jnot g14861(.din(w_n14770_0[0]),.dout(n15111),.clk(gclk));
	jor g14862(.dina(w_n15111_0[1]),.dinb(n15110),.dout(n15112),.clk(gclk));
	jand g14863(.dina(n15112),.dinb(n15051),.dout(n15113),.clk(gclk));
	jand g14864(.dina(n15113),.dinb(w_n7581_25[1]),.dout(n15114),.clk(gclk));
	jor g14865(.dina(w_n14777_0[0]),.dinb(n15114),.dout(n15115),.clk(gclk));
	jand g14866(.dina(n15115),.dinb(n15050),.dout(n15116),.clk(gclk));
	jand g14867(.dina(n15116),.dinb(w_n7154_30[1]),.dout(n15117),.clk(gclk));
	jnot g14868(.din(w_n14785_0[0]),.dout(n15118),.clk(gclk));
	jor g14869(.dina(w_n15118_0[1]),.dinb(n15117),.dout(n15119),.clk(gclk));
	jand g14870(.dina(n15119),.dinb(n15049),.dout(n15120),.clk(gclk));
	jand g14871(.dina(n15120),.dinb(w_n6758_26[0]),.dout(n15121),.clk(gclk));
	jor g14872(.dina(w_n14792_0[0]),.dinb(n15121),.dout(n15122),.clk(gclk));
	jand g14873(.dina(n15122),.dinb(n15048),.dout(n15123),.clk(gclk));
	jand g14874(.dina(n15123),.dinb(w_n6357_30[2]),.dout(n15124),.clk(gclk));
	jor g14875(.dina(w_n14800_0[0]),.dinb(n15124),.dout(n15125),.clk(gclk));
	jand g14876(.dina(n15125),.dinb(n15047),.dout(n15126),.clk(gclk));
	jand g14877(.dina(n15126),.dinb(w_n5989_26[2]),.dout(n15127),.clk(gclk));
	jor g14878(.dina(w_n14808_0[0]),.dinb(n15127),.dout(n15128),.clk(gclk));
	jand g14879(.dina(n15128),.dinb(n15046),.dout(n15129),.clk(gclk));
	jand g14880(.dina(n15129),.dinb(w_n5606_31[0]),.dout(n15130),.clk(gclk));
	jnot g14881(.din(w_n14816_0[0]),.dout(n15131),.clk(gclk));
	jor g14882(.dina(w_n15131_0[1]),.dinb(n15130),.dout(n15132),.clk(gclk));
	jand g14883(.dina(n15132),.dinb(n15045),.dout(n15133),.clk(gclk));
	jand g14884(.dina(n15133),.dinb(w_n5259_27[2]),.dout(n15134),.clk(gclk));
	jor g14885(.dina(w_n14823_0[0]),.dinb(n15134),.dout(n15135),.clk(gclk));
	jand g14886(.dina(n15135),.dinb(n15044),.dout(n15136),.clk(gclk));
	jand g14887(.dina(n15136),.dinb(w_n4902_31[2]),.dout(n15137),.clk(gclk));
	jnot g14888(.din(w_n14831_0[0]),.dout(n15138),.clk(gclk));
	jor g14889(.dina(w_n15138_0[1]),.dinb(n15137),.dout(n15139),.clk(gclk));
	jand g14890(.dina(n15139),.dinb(n15043),.dout(n15140),.clk(gclk));
	jand g14891(.dina(n15140),.dinb(w_n4582_28[2]),.dout(n15141),.clk(gclk));
	jor g14892(.dina(w_n14838_0[0]),.dinb(n15141),.dout(n15142),.clk(gclk));
	jand g14893(.dina(n15142),.dinb(n15042),.dout(n15143),.clk(gclk));
	jand g14894(.dina(n15143),.dinb(w_n4249_32[1]),.dout(n15144),.clk(gclk));
	jor g14895(.dina(w_n14846_0[0]),.dinb(n15144),.dout(n15145),.clk(gclk));
	jand g14896(.dina(n15145),.dinb(n15041),.dout(n15146),.clk(gclk));
	jand g14897(.dina(n15146),.dinb(w_n3955_29[1]),.dout(n15147),.clk(gclk));
	jor g14898(.dina(w_n14854_0[0]),.dinb(n15147),.dout(n15148),.clk(gclk));
	jand g14899(.dina(n15148),.dinb(n15040),.dout(n15149),.clk(gclk));
	jand g14900(.dina(n15149),.dinb(w_n3642_32[2]),.dout(n15150),.clk(gclk));
	jnot g14901(.din(w_n14862_0[0]),.dout(n15151),.clk(gclk));
	jor g14902(.dina(w_n15151_0[1]),.dinb(n15150),.dout(n15152),.clk(gclk));
	jand g14903(.dina(n15152),.dinb(n15039),.dout(n15153),.clk(gclk));
	jand g14904(.dina(n15153),.dinb(w_n3368_30[0]),.dout(n15154),.clk(gclk));
	jor g14905(.dina(w_n14869_0[0]),.dinb(n15154),.dout(n15155),.clk(gclk));
	jand g14906(.dina(n15155),.dinb(n15038),.dout(n15156),.clk(gclk));
	jand g14907(.dina(n15156),.dinb(w_n3089_33[1]),.dout(n15157),.clk(gclk));
	jnot g14908(.din(w_n14877_0[0]),.dout(n15158),.clk(gclk));
	jor g14909(.dina(w_n15158_0[1]),.dinb(n15157),.dout(n15159),.clk(gclk));
	jand g14910(.dina(n15159),.dinb(n15037),.dout(n15160),.clk(gclk));
	jand g14911(.dina(n15160),.dinb(w_n2833_31[0]),.dout(n15161),.clk(gclk));
	jor g14912(.dina(w_n14884_0[0]),.dinb(n15161),.dout(n15162),.clk(gclk));
	jand g14913(.dina(n15162),.dinb(n15036),.dout(n15163),.clk(gclk));
	jand g14914(.dina(n15163),.dinb(w_n2572_33[2]),.dout(n15164),.clk(gclk));
	jor g14915(.dina(w_n14892_0[0]),.dinb(n15164),.dout(n15165),.clk(gclk));
	jand g14916(.dina(n15165),.dinb(n15035),.dout(n15166),.clk(gclk));
	jand g14917(.dina(n15166),.dinb(w_n2345_31[2]),.dout(n15167),.clk(gclk));
	jnot g14918(.din(w_n14900_0[0]),.dout(n15168),.clk(gclk));
	jor g14919(.dina(w_n15168_0[1]),.dinb(n15167),.dout(n15169),.clk(gclk));
	jand g14920(.dina(n15169),.dinb(n15034),.dout(n15170),.clk(gclk));
	jand g14921(.dina(n15170),.dinb(w_n2108_34[1]),.dout(n15171),.clk(gclk));
	jor g14922(.dina(n15171),.dinb(w_n15033_0[1]),.dout(n15172),.clk(gclk));
	jand g14923(.dina(n15172),.dinb(n15032),.dout(n15173),.clk(gclk));
	jand g14924(.dina(n15173),.dinb(w_n1912_32[2]),.dout(n15174),.clk(gclk));
	jor g14925(.dina(w_n14914_0[0]),.dinb(n15174),.dout(n15175),.clk(gclk));
	jand g14926(.dina(n15175),.dinb(n15031),.dout(n15176),.clk(gclk));
	jand g14927(.dina(n15176),.dinb(w_n1699_35[0]),.dout(n15177),.clk(gclk));
	jnot g14928(.din(w_n14922_0[0]),.dout(n15178),.clk(gclk));
	jor g14929(.dina(w_n15178_0[1]),.dinb(n15177),.dout(n15179),.clk(gclk));
	jand g14930(.dina(n15179),.dinb(n15030),.dout(n15180),.clk(gclk));
	jand g14931(.dina(n15180),.dinb(w_n1516_33[1]),.dout(n15181),.clk(gclk));
	jor g14932(.dina(w_n14929_0[0]),.dinb(n15181),.dout(n15182),.clk(gclk));
	jand g14933(.dina(n15182),.dinb(n15029),.dout(n15183),.clk(gclk));
	jand g14934(.dina(n15183),.dinb(w_n1332_35[0]),.dout(n15184),.clk(gclk));
	jnot g14935(.din(w_n14937_0[0]),.dout(n15185),.clk(gclk));
	jor g14936(.dina(w_n15185_0[1]),.dinb(n15184),.dout(n15186),.clk(gclk));
	jand g14937(.dina(n15186),.dinb(n15028),.dout(n15187),.clk(gclk));
	jand g14938(.dina(n15187),.dinb(w_n1173_34[0]),.dout(n15188),.clk(gclk));
	jor g14939(.dina(w_n14944_0[0]),.dinb(n15188),.dout(n15189),.clk(gclk));
	jand g14940(.dina(n15189),.dinb(n15027),.dout(n15190),.clk(gclk));
	jand g14941(.dina(n15190),.dinb(w_n1008_36[0]),.dout(n15191),.clk(gclk));
	jor g14942(.dina(w_n14952_0[0]),.dinb(n15191),.dout(n15192),.clk(gclk));
	jand g14943(.dina(n15192),.dinb(n15026),.dout(n15193),.clk(gclk));
	jand g14944(.dina(n15193),.dinb(w_n884_35[0]),.dout(n15194),.clk(gclk));
	jor g14945(.dina(w_n14960_0[0]),.dinb(n15194),.dout(n15195),.clk(gclk));
	jand g14946(.dina(n15195),.dinb(n15025),.dout(n15196),.clk(gclk));
	jand g14947(.dina(n15196),.dinb(w_n743_36[0]),.dout(n15197),.clk(gclk));
	jnot g14948(.din(w_n14968_0[0]),.dout(n15198),.clk(gclk));
	jor g14949(.dina(w_n15198_0[1]),.dinb(n15197),.dout(n15199),.clk(gclk));
	jand g14950(.dina(n15199),.dinb(n15024),.dout(n15200),.clk(gclk));
	jand g14951(.dina(n15200),.dinb(w_n635_36[0]),.dout(n15201),.clk(gclk));
	jor g14952(.dina(w_n14975_0[0]),.dinb(n15201),.dout(n15202),.clk(gclk));
	jand g14953(.dina(n15202),.dinb(n15023),.dout(n15203),.clk(gclk));
	jand g14954(.dina(n15203),.dinb(w_n515_37[0]),.dout(n15204),.clk(gclk));
	jnot g14955(.din(w_n14983_0[0]),.dout(n15205),.clk(gclk));
	jor g14956(.dina(w_n15205_0[1]),.dinb(n15204),.dout(n15206),.clk(gclk));
	jand g14957(.dina(n15206),.dinb(n15022),.dout(n15207),.clk(gclk));
	jand g14958(.dina(n15207),.dinb(w_n443_37[0]),.dout(n15208),.clk(gclk));
	jor g14959(.dina(w_n14990_0[0]),.dinb(n15208),.dout(n15209),.clk(gclk));
	jand g14960(.dina(n15209),.dinb(n15021),.dout(n15210),.clk(gclk));
	jand g14961(.dina(n15210),.dinb(w_n352_37[1]),.dout(n15211),.clk(gclk));
	jnot g14962(.din(w_n14998_0[0]),.dout(n15212),.clk(gclk));
	jor g14963(.dina(w_n15212_0[1]),.dinb(n15211),.dout(n15213),.clk(gclk));
	jand g14964(.dina(n15213),.dinb(n15020),.dout(n15214),.clk(gclk));
	jand g14965(.dina(n15214),.dinb(w_n294_37[2]),.dout(n15215),.clk(gclk));
	jor g14966(.dina(w_n15005_0[0]),.dinb(n15215),.dout(n15216),.clk(gclk));
	jand g14967(.dina(n15216),.dinb(n15019),.dout(n15217),.clk(gclk));
	jand g14968(.dina(n15217),.dinb(w_n239_38[0]),.dout(n15218),.clk(gclk));
	jnot g14969(.din(w_n15013_0[0]),.dout(n15219),.clk(gclk));
	jor g14970(.dina(w_n15219_0[1]),.dinb(n15218),.dout(n15220),.clk(gclk));
	jand g14971(.dina(n15220),.dinb(n15018),.dout(n15221),.clk(gclk));
	jand g14972(.dina(n15221),.dinb(w_n221_38[1]),.dout(n15222),.clk(gclk));
	jxor g14973(.dina(w_n14407_0[0]),.dinb(w_n239_37[2]),.dout(n15223),.clk(gclk));
	jand g14974(.dina(n15223),.dinb(w_asqrt16_19[0]),.dout(n15224),.clk(gclk));
	jxor g14975(.dina(n15224),.dinb(w_n14412_0[0]),.dout(n15225),.clk(gclk));
	jnot g14976(.din(w_n15225_0[1]),.dout(n15226),.clk(gclk));
	jor g14977(.dina(w_n15226_0[1]),.dinb(n15222),.dout(n15227),.clk(gclk));
	jand g14978(.dina(n15227),.dinb(n15017),.dout(n15228),.clk(gclk));
	jxor g14979(.dina(w_n14415_0[0]),.dinb(w_n221_38[0]),.dout(n15229),.clk(gclk));
	jand g14980(.dina(n15229),.dinb(w_asqrt16_18[2]),.dout(n15230),.clk(gclk));
	jxor g14981(.dina(n15230),.dinb(w_n14421_0[0]),.dout(n15231),.clk(gclk));
	jor g14982(.dina(w_n15231_1[1]),.dinb(w_n15228_0[2]),.dout(n15232),.clk(gclk));
	jxor g14983(.dina(w_n14426_0[2]),.dinb(w_n14423_0[2]),.dout(n15233),.clk(gclk));
	jnot g14984(.din(w_n15233_0[1]),.dout(n15234),.clk(gclk));
	jand g14985(.dina(n15234),.dinb(w_asqrt16_18[1]),.dout(n15235),.clk(gclk));
	jor g14986(.dina(w_n15235_0[1]),.dinb(w_n15232_0[1]),.dout(n15236),.clk(gclk));
	jand g14987(.dina(n15236),.dinb(w_n218_16[0]),.dout(n15237),.clk(gclk));
	jand g14988(.dina(w_n14674_19[1]),.dinb(w_n14426_0[1]),.dout(n15238),.clk(gclk));
	jand g14989(.dina(w_n15231_1[0]),.dinb(w_n15228_0[1]),.dout(n15239),.clk(gclk));
	jor g14990(.dina(w_n15239_0[2]),.dinb(w_n15238_0[1]),.dout(n15240),.clk(gclk));
	jand g14991(.dina(w_n14672_0[0]),.dinb(w_n14423_0[1]),.dout(n15241),.clk(gclk));
	jnot g14992(.din(n15241),.dout(n15242),.clk(gclk));
	jand g14993(.dina(w_n15233_0[0]),.dinb(w_asqrt63_28[0]),.dout(n15243),.clk(gclk));
	jand g14994(.dina(w_n15243_0[1]),.dinb(n15242),.dout(n15244),.clk(gclk));
	jor g14995(.dina(w_n15244_0[1]),.dinb(n15240),.dout(n15245),.clk(gclk));
	jor g14996(.dina(n15245),.dinb(w_n15237_0[1]),.dout(asqrt_fa_16),.clk(gclk));
	jor g14997(.dina(w_n15015_0[1]),.dinb(w_asqrt62_22[0]),.dout(n15247),.clk(gclk));
	jand g14998(.dina(w_n15225_0[0]),.dinb(n15247),.dout(n15248),.clk(gclk));
	jor g14999(.dina(n15248),.dinb(w_n15016_0[0]),.dout(n15249),.clk(gclk));
	jnot g15000(.din(w_n15231_0[2]),.dout(n15250),.clk(gclk));
	jand g15001(.dina(w_n15250_0[1]),.dinb(w_n15249_0[1]),.dout(n15251),.clk(gclk));
	jnot g15002(.din(w_n15235_0[0]),.dout(n15252),.clk(gclk));
	jand g15003(.dina(n15252),.dinb(w_n15251_0[1]),.dout(n15253),.clk(gclk));
	jor g15004(.dina(n15253),.dinb(w_asqrt63_27[2]),.dout(n15254),.clk(gclk));
	jnot g15005(.din(w_n15238_0[0]),.dout(n15255),.clk(gclk));
	jor g15006(.dina(w_n15250_0[0]),.dinb(w_n15249_0[0]),.dout(n15256),.clk(gclk));
	jand g15007(.dina(w_n15256_0[2]),.dinb(n15255),.dout(n15257),.clk(gclk));
	jnot g15008(.din(w_n15244_0[0]),.dout(n15258),.clk(gclk));
	jand g15009(.dina(n15258),.dinb(n15257),.dout(n15259),.clk(gclk));
	jand g15010(.dina(n15259),.dinb(n15254),.dout(n15260),.clk(gclk));
	jxor g15011(.dina(w_n15015_0[0]),.dinb(w_n221_37[2]),.dout(n15261),.clk(gclk));
	jor g15012(.dina(n15261),.dinb(w_n15260_41[2]),.dout(n15262),.clk(gclk));
	jxor g15013(.dina(n15262),.dinb(w_n15226_0[0]),.dout(n15263),.clk(gclk));
	jnot g15014(.din(w_n15263_0[1]),.dout(n15264),.clk(gclk));
	jnot g15015(.din(w_a28_0[2]),.dout(n15265),.clk(gclk));
	jnot g15016(.din(w_a29_0[1]),.dout(n15266),.clk(gclk));
	jand g15017(.dina(w_n15266_0[1]),.dinb(w_n15265_1[2]),.dout(n15267),.clk(gclk));
	jand g15018(.dina(w_n15267_0[2]),.dinb(w_n14443_1[0]),.dout(n15268),.clk(gclk));
	jnot g15019(.din(w_n15268_0[1]),.dout(n15269),.clk(gclk));
	jor g15020(.dina(w_n15260_41[1]),.dinb(w_n14443_0[2]),.dout(n15270),.clk(gclk));
	jand g15021(.dina(n15270),.dinb(n15269),.dout(n15271),.clk(gclk));
	jor g15022(.dina(w_n15271_0[2]),.dinb(w_n14674_19[0]),.dout(n15272),.clk(gclk));
	jand g15023(.dina(w_n15271_0[1]),.dinb(w_n14674_18[2]),.dout(n15273),.clk(gclk));
	jor g15024(.dina(w_n15260_41[0]),.dinb(w_a30_1[0]),.dout(n15274),.clk(gclk));
	jand g15025(.dina(n15274),.dinb(w_a31_0[0]),.dout(n15275),.clk(gclk));
	jand g15026(.dina(w_asqrt15_12),.dinb(w_n14445_0[1]),.dout(n15276),.clk(gclk));
	jor g15027(.dina(n15276),.dinb(n15275),.dout(n15277),.clk(gclk));
	jor g15028(.dina(n15277),.dinb(n15273),.dout(n15278),.clk(gclk));
	jand g15029(.dina(n15278),.dinb(w_n15272_0[1]),.dout(n15279),.clk(gclk));
	jor g15030(.dina(w_n15279_0[2]),.dinb(w_n14078_26[1]),.dout(n15280),.clk(gclk));
	jand g15031(.dina(w_n15279_0[1]),.dinb(w_n14078_26[0]),.dout(n15281),.clk(gclk));
	jnot g15032(.din(w_n14445_0[0]),.dout(n15282),.clk(gclk));
	jor g15033(.dina(w_n15260_40[2]),.dinb(n15282),.dout(n15283),.clk(gclk));
	jor g15034(.dina(w_n15239_0[1]),.dinb(w_n14674_18[1]),.dout(n15284),.clk(gclk));
	jor g15035(.dina(n15284),.dinb(w_n15237_0[0]),.dout(n15285),.clk(gclk));
	jor g15036(.dina(n15285),.dinb(w_n15243_0[0]),.dout(n15286),.clk(gclk));
	jand g15037(.dina(n15286),.dinb(w_n15283_0[1]),.dout(n15287),.clk(gclk));
	jxor g15038(.dina(n15287),.dinb(w_n14080_0[1]),.dout(n15288),.clk(gclk));
	jor g15039(.dina(w_n15288_0[1]),.dinb(n15281),.dout(n15289),.clk(gclk));
	jand g15040(.dina(n15289),.dinb(w_n15280_0[1]),.dout(n15290),.clk(gclk));
	jor g15041(.dina(w_n15290_0[2]),.dinb(w_n13515_20[0]),.dout(n15291),.clk(gclk));
	jand g15042(.dina(w_n15290_0[1]),.dinb(w_n13515_19[2]),.dout(n15292),.clk(gclk));
	jxor g15043(.dina(w_n14448_0[0]),.dinb(w_n14078_25[2]),.dout(n15293),.clk(gclk));
	jor g15044(.dina(n15293),.dinb(w_n15260_40[1]),.dout(n15294),.clk(gclk));
	jxor g15045(.dina(n15294),.dinb(w_n15070_0[0]),.dout(n15295),.clk(gclk));
	jnot g15046(.din(w_n15295_0[2]),.dout(n15296),.clk(gclk));
	jor g15047(.dina(n15296),.dinb(n15292),.dout(n15297),.clk(gclk));
	jand g15048(.dina(n15297),.dinb(w_n15291_0[1]),.dout(n15298),.clk(gclk));
	jor g15049(.dina(w_n15298_0[2]),.dinb(w_n12947_27[0]),.dout(n15299),.clk(gclk));
	jand g15050(.dina(w_n15298_0[1]),.dinb(w_n12947_26[2]),.dout(n15300),.clk(gclk));
	jxor g15051(.dina(w_n14678_0[0]),.dinb(w_n13515_19[1]),.dout(n15301),.clk(gclk));
	jor g15052(.dina(n15301),.dinb(w_n15260_40[0]),.dout(n15302),.clk(gclk));
	jxor g15053(.dina(n15302),.dinb(w_n14687_0[0]),.dout(n15303),.clk(gclk));
	jor g15054(.dina(w_n15303_0[2]),.dinb(n15300),.dout(n15304),.clk(gclk));
	jand g15055(.dina(n15304),.dinb(w_n15299_0[1]),.dout(n15305),.clk(gclk));
	jor g15056(.dina(w_n15305_0[2]),.dinb(w_n12410_20[2]),.dout(n15306),.clk(gclk));
	jand g15057(.dina(w_n15305_0[1]),.dinb(w_n12410_20[1]),.dout(n15307),.clk(gclk));
	jxor g15058(.dina(w_n14689_0[0]),.dinb(w_n12947_26[1]),.dout(n15308),.clk(gclk));
	jor g15059(.dina(n15308),.dinb(w_n15260_39[2]),.dout(n15309),.clk(gclk));
	jxor g15060(.dina(n15309),.dinb(w_n15077_0[0]),.dout(n15310),.clk(gclk));
	jnot g15061(.din(w_n15310_0[2]),.dout(n15311),.clk(gclk));
	jor g15062(.dina(n15311),.dinb(n15307),.dout(n15312),.clk(gclk));
	jand g15063(.dina(n15312),.dinb(w_n15306_0[1]),.dout(n15313),.clk(gclk));
	jor g15064(.dina(w_n15313_0[2]),.dinb(w_n11858_27[1]),.dout(n15314),.clk(gclk));
	jand g15065(.dina(w_n15313_0[1]),.dinb(w_n11858_27[0]),.dout(n15315),.clk(gclk));
	jxor g15066(.dina(w_n14696_0[0]),.dinb(w_n12410_20[0]),.dout(n15316),.clk(gclk));
	jor g15067(.dina(n15316),.dinb(w_n15260_39[1]),.dout(n15317),.clk(gclk));
	jxor g15068(.dina(n15317),.dinb(w_n14702_0[0]),.dout(n15318),.clk(gclk));
	jor g15069(.dina(w_n15318_0[2]),.dinb(n15315),.dout(n15319),.clk(gclk));
	jand g15070(.dina(n15319),.dinb(w_n15314_0[1]),.dout(n15320),.clk(gclk));
	jor g15071(.dina(w_n15320_0[2]),.dinb(w_n11347_21[1]),.dout(n15321),.clk(gclk));
	jand g15072(.dina(w_n15320_0[1]),.dinb(w_n11347_21[0]),.dout(n15322),.clk(gclk));
	jxor g15073(.dina(w_n14704_0[0]),.dinb(w_n11858_26[2]),.dout(n15323),.clk(gclk));
	jor g15074(.dina(n15323),.dinb(w_n15260_39[0]),.dout(n15324),.clk(gclk));
	jxor g15075(.dina(n15324),.dinb(w_n15084_0[0]),.dout(n15325),.clk(gclk));
	jnot g15076(.din(w_n15325_0[2]),.dout(n15326),.clk(gclk));
	jor g15077(.dina(n15326),.dinb(n15322),.dout(n15327),.clk(gclk));
	jand g15078(.dina(n15327),.dinb(w_n15321_0[1]),.dout(n15328),.clk(gclk));
	jor g15079(.dina(w_n15328_0[2]),.dinb(w_n10824_28[0]),.dout(n15329),.clk(gclk));
	jand g15080(.dina(w_n15328_0[1]),.dinb(w_n10824_27[2]),.dout(n15330),.clk(gclk));
	jxor g15081(.dina(w_n14711_0[0]),.dinb(w_n11347_20[2]),.dout(n15331),.clk(gclk));
	jor g15082(.dina(n15331),.dinb(w_n15260_38[2]),.dout(n15332),.clk(gclk));
	jxor g15083(.dina(n15332),.dinb(w_n14717_0[0]),.dout(n15333),.clk(gclk));
	jor g15084(.dina(w_n15333_0[2]),.dinb(n15330),.dout(n15334),.clk(gclk));
	jand g15085(.dina(n15334),.dinb(w_n15329_0[1]),.dout(n15335),.clk(gclk));
	jor g15086(.dina(w_n15335_0[2]),.dinb(w_n10328_22[1]),.dout(n15336),.clk(gclk));
	jand g15087(.dina(w_n15335_0[1]),.dinb(w_n10328_22[0]),.dout(n15337),.clk(gclk));
	jxor g15088(.dina(w_n14719_0[0]),.dinb(w_n10824_27[1]),.dout(n15338),.clk(gclk));
	jor g15089(.dina(n15338),.dinb(w_n15260_38[1]),.dout(n15339),.clk(gclk));
	jxor g15090(.dina(n15339),.dinb(w_n14725_0[0]),.dout(n15340),.clk(gclk));
	jor g15091(.dina(w_n15340_0[2]),.dinb(n15337),.dout(n15341),.clk(gclk));
	jand g15092(.dina(n15341),.dinb(w_n15336_0[1]),.dout(n15342),.clk(gclk));
	jor g15093(.dina(w_n15342_0[2]),.dinb(w_n9832_28[2]),.dout(n15343),.clk(gclk));
	jand g15094(.dina(w_n15342_0[1]),.dinb(w_n9832_28[1]),.dout(n15344),.clk(gclk));
	jxor g15095(.dina(w_n14727_0[0]),.dinb(w_n10328_21[2]),.dout(n15345),.clk(gclk));
	jor g15096(.dina(n15345),.dinb(w_n15260_38[0]),.dout(n15346),.clk(gclk));
	jxor g15097(.dina(n15346),.dinb(w_n14733_0[0]),.dout(n15347),.clk(gclk));
	jor g15098(.dina(w_n15347_0[2]),.dinb(n15344),.dout(n15348),.clk(gclk));
	jand g15099(.dina(n15348),.dinb(w_n15343_0[1]),.dout(n15349),.clk(gclk));
	jor g15100(.dina(w_n15349_0[2]),.dinb(w_n9369_23[1]),.dout(n15350),.clk(gclk));
	jand g15101(.dina(w_n15349_0[1]),.dinb(w_n9369_23[0]),.dout(n15351),.clk(gclk));
	jxor g15102(.dina(w_n14735_0[0]),.dinb(w_n9832_28[0]),.dout(n15352),.clk(gclk));
	jor g15103(.dina(n15352),.dinb(w_n15260_37[2]),.dout(n15353),.clk(gclk));
	jxor g15104(.dina(n15353),.dinb(w_n15097_0[0]),.dout(n15354),.clk(gclk));
	jnot g15105(.din(w_n15354_0[2]),.dout(n15355),.clk(gclk));
	jor g15106(.dina(n15355),.dinb(n15351),.dout(n15356),.clk(gclk));
	jand g15107(.dina(n15356),.dinb(w_n15350_0[1]),.dout(n15357),.clk(gclk));
	jor g15108(.dina(w_n15357_0[2]),.dinb(w_n8890_29[0]),.dout(n15358),.clk(gclk));
	jand g15109(.dina(w_n15357_0[1]),.dinb(w_n8890_28[2]),.dout(n15359),.clk(gclk));
	jxor g15110(.dina(w_n14742_0[0]),.dinb(w_n9369_22[2]),.dout(n15360),.clk(gclk));
	jor g15111(.dina(n15360),.dinb(w_n15260_37[1]),.dout(n15361),.clk(gclk));
	jxor g15112(.dina(n15361),.dinb(w_n14748_0[0]),.dout(n15362),.clk(gclk));
	jor g15113(.dina(w_n15362_0[2]),.dinb(n15359),.dout(n15363),.clk(gclk));
	jand g15114(.dina(n15363),.dinb(w_n15358_0[1]),.dout(n15364),.clk(gclk));
	jor g15115(.dina(w_n15364_0[2]),.dinb(w_n8449_24[0]),.dout(n15365),.clk(gclk));
	jand g15116(.dina(w_n15364_0[1]),.dinb(w_n8449_23[2]),.dout(n15366),.clk(gclk));
	jxor g15117(.dina(w_n14750_0[0]),.dinb(w_n8890_28[1]),.dout(n15367),.clk(gclk));
	jor g15118(.dina(n15367),.dinb(w_n15260_37[0]),.dout(n15368),.clk(gclk));
	jxor g15119(.dina(n15368),.dinb(w_n15104_0[0]),.dout(n15369),.clk(gclk));
	jnot g15120(.din(w_n15369_0[2]),.dout(n15370),.clk(gclk));
	jor g15121(.dina(n15370),.dinb(n15366),.dout(n15371),.clk(gclk));
	jand g15122(.dina(n15371),.dinb(w_n15365_0[1]),.dout(n15372),.clk(gclk));
	jor g15123(.dina(w_n15372_0[2]),.dinb(w_n8003_29[2]),.dout(n15373),.clk(gclk));
	jand g15124(.dina(w_n15372_0[1]),.dinb(w_n8003_29[1]),.dout(n15374),.clk(gclk));
	jxor g15125(.dina(w_n14757_0[0]),.dinb(w_n8449_23[1]),.dout(n15375),.clk(gclk));
	jor g15126(.dina(n15375),.dinb(w_n15260_36[2]),.dout(n15376),.clk(gclk));
	jxor g15127(.dina(n15376),.dinb(w_n14763_0[0]),.dout(n15377),.clk(gclk));
	jor g15128(.dina(w_n15377_0[2]),.dinb(n15374),.dout(n15378),.clk(gclk));
	jand g15129(.dina(n15378),.dinb(w_n15373_0[1]),.dout(n15379),.clk(gclk));
	jor g15130(.dina(w_n15379_0[2]),.dinb(w_n7581_25[0]),.dout(n15380),.clk(gclk));
	jand g15131(.dina(w_n15379_0[1]),.dinb(w_n7581_24[2]),.dout(n15381),.clk(gclk));
	jxor g15132(.dina(w_n14765_0[0]),.dinb(w_n8003_29[0]),.dout(n15382),.clk(gclk));
	jor g15133(.dina(n15382),.dinb(w_n15260_36[1]),.dout(n15383),.clk(gclk));
	jxor g15134(.dina(n15383),.dinb(w_n15111_0[0]),.dout(n15384),.clk(gclk));
	jnot g15135(.din(w_n15384_0[2]),.dout(n15385),.clk(gclk));
	jor g15136(.dina(n15385),.dinb(n15381),.dout(n15386),.clk(gclk));
	jand g15137(.dina(n15386),.dinb(w_n15380_0[1]),.dout(n15387),.clk(gclk));
	jor g15138(.dina(w_n15387_0[2]),.dinb(w_n7154_30[0]),.dout(n15388),.clk(gclk));
	jand g15139(.dina(w_n15387_0[1]),.dinb(w_n7154_29[2]),.dout(n15389),.clk(gclk));
	jxor g15140(.dina(w_n14772_0[0]),.dinb(w_n7581_24[1]),.dout(n15390),.clk(gclk));
	jor g15141(.dina(n15390),.dinb(w_n15260_36[0]),.dout(n15391),.clk(gclk));
	jxor g15142(.dina(n15391),.dinb(w_n14778_0[0]),.dout(n15392),.clk(gclk));
	jor g15143(.dina(w_n15392_0[2]),.dinb(n15389),.dout(n15393),.clk(gclk));
	jand g15144(.dina(n15393),.dinb(w_n15388_0[1]),.dout(n15394),.clk(gclk));
	jor g15145(.dina(w_n15394_0[2]),.dinb(w_n6758_25[2]),.dout(n15395),.clk(gclk));
	jand g15146(.dina(w_n15394_0[1]),.dinb(w_n6758_25[1]),.dout(n15396),.clk(gclk));
	jxor g15147(.dina(w_n14780_0[0]),.dinb(w_n7154_29[1]),.dout(n15397),.clk(gclk));
	jor g15148(.dina(n15397),.dinb(w_n15260_35[2]),.dout(n15398),.clk(gclk));
	jxor g15149(.dina(n15398),.dinb(w_n15118_0[0]),.dout(n15399),.clk(gclk));
	jnot g15150(.din(w_n15399_0[2]),.dout(n15400),.clk(gclk));
	jor g15151(.dina(n15400),.dinb(n15396),.dout(n15401),.clk(gclk));
	jand g15152(.dina(n15401),.dinb(w_n15395_0[1]),.dout(n15402),.clk(gclk));
	jor g15153(.dina(w_n15402_0[2]),.dinb(w_n6357_30[1]),.dout(n15403),.clk(gclk));
	jand g15154(.dina(w_n15402_0[1]),.dinb(w_n6357_30[0]),.dout(n15404),.clk(gclk));
	jxor g15155(.dina(w_n14787_0[0]),.dinb(w_n6758_25[0]),.dout(n15405),.clk(gclk));
	jor g15156(.dina(n15405),.dinb(w_n15260_35[1]),.dout(n15406),.clk(gclk));
	jxor g15157(.dina(n15406),.dinb(w_n14793_0[0]),.dout(n15407),.clk(gclk));
	jor g15158(.dina(w_n15407_0[2]),.dinb(n15404),.dout(n15408),.clk(gclk));
	jand g15159(.dina(n15408),.dinb(w_n15403_0[1]),.dout(n15409),.clk(gclk));
	jor g15160(.dina(w_n15409_0[2]),.dinb(w_n5989_26[1]),.dout(n15410),.clk(gclk));
	jand g15161(.dina(w_n15409_0[1]),.dinb(w_n5989_26[0]),.dout(n15411),.clk(gclk));
	jxor g15162(.dina(w_n14795_0[0]),.dinb(w_n6357_29[2]),.dout(n15412),.clk(gclk));
	jor g15163(.dina(n15412),.dinb(w_n15260_35[0]),.dout(n15413),.clk(gclk));
	jxor g15164(.dina(n15413),.dinb(w_n14801_0[0]),.dout(n15414),.clk(gclk));
	jor g15165(.dina(w_n15414_0[2]),.dinb(n15411),.dout(n15415),.clk(gclk));
	jand g15166(.dina(n15415),.dinb(w_n15410_0[1]),.dout(n15416),.clk(gclk));
	jor g15167(.dina(w_n15416_0[2]),.dinb(w_n5606_30[2]),.dout(n15417),.clk(gclk));
	jand g15168(.dina(w_n15416_0[1]),.dinb(w_n5606_30[1]),.dout(n15418),.clk(gclk));
	jxor g15169(.dina(w_n14803_0[0]),.dinb(w_n5989_25[2]),.dout(n15419),.clk(gclk));
	jor g15170(.dina(n15419),.dinb(w_n15260_34[2]),.dout(n15420),.clk(gclk));
	jxor g15171(.dina(n15420),.dinb(w_n14809_0[0]),.dout(n15421),.clk(gclk));
	jor g15172(.dina(w_n15421_0[2]),.dinb(n15418),.dout(n15422),.clk(gclk));
	jand g15173(.dina(n15422),.dinb(w_n15417_0[1]),.dout(n15423),.clk(gclk));
	jor g15174(.dina(w_n15423_0[2]),.dinb(w_n5259_27[1]),.dout(n15424),.clk(gclk));
	jand g15175(.dina(w_n15423_0[1]),.dinb(w_n5259_27[0]),.dout(n15425),.clk(gclk));
	jxor g15176(.dina(w_n14811_0[0]),.dinb(w_n5606_30[0]),.dout(n15426),.clk(gclk));
	jor g15177(.dina(n15426),.dinb(w_n15260_34[1]),.dout(n15427),.clk(gclk));
	jxor g15178(.dina(n15427),.dinb(w_n15131_0[0]),.dout(n15428),.clk(gclk));
	jnot g15179(.din(w_n15428_0[2]),.dout(n15429),.clk(gclk));
	jor g15180(.dina(n15429),.dinb(n15425),.dout(n15430),.clk(gclk));
	jand g15181(.dina(n15430),.dinb(w_n15424_0[1]),.dout(n15431),.clk(gclk));
	jor g15182(.dina(w_n15431_0[2]),.dinb(w_n4902_31[1]),.dout(n15432),.clk(gclk));
	jand g15183(.dina(w_n15431_0[1]),.dinb(w_n4902_31[0]),.dout(n15433),.clk(gclk));
	jxor g15184(.dina(w_n14818_0[0]),.dinb(w_n5259_26[2]),.dout(n15434),.clk(gclk));
	jor g15185(.dina(n15434),.dinb(w_n15260_34[0]),.dout(n15435),.clk(gclk));
	jxor g15186(.dina(n15435),.dinb(w_n14824_0[0]),.dout(n15436),.clk(gclk));
	jor g15187(.dina(w_n15436_0[2]),.dinb(n15433),.dout(n15437),.clk(gclk));
	jand g15188(.dina(n15437),.dinb(w_n15432_0[1]),.dout(n15438),.clk(gclk));
	jor g15189(.dina(w_n15438_0[2]),.dinb(w_n4582_28[1]),.dout(n15439),.clk(gclk));
	jand g15190(.dina(w_n15438_0[1]),.dinb(w_n4582_28[0]),.dout(n15440),.clk(gclk));
	jxor g15191(.dina(w_n14826_0[0]),.dinb(w_n4902_30[2]),.dout(n15441),.clk(gclk));
	jor g15192(.dina(n15441),.dinb(w_n15260_33[2]),.dout(n15442),.clk(gclk));
	jxor g15193(.dina(n15442),.dinb(w_n15138_0[0]),.dout(n15443),.clk(gclk));
	jnot g15194(.din(w_n15443_0[2]),.dout(n15444),.clk(gclk));
	jor g15195(.dina(n15444),.dinb(n15440),.dout(n15445),.clk(gclk));
	jand g15196(.dina(n15445),.dinb(w_n15439_0[1]),.dout(n15446),.clk(gclk));
	jor g15197(.dina(w_n15446_0[2]),.dinb(w_n4249_32[0]),.dout(n15447),.clk(gclk));
	jand g15198(.dina(w_n15446_0[1]),.dinb(w_n4249_31[2]),.dout(n15448),.clk(gclk));
	jxor g15199(.dina(w_n14833_0[0]),.dinb(w_n4582_27[2]),.dout(n15449),.clk(gclk));
	jor g15200(.dina(n15449),.dinb(w_n15260_33[1]),.dout(n15450),.clk(gclk));
	jxor g15201(.dina(n15450),.dinb(w_n14839_0[0]),.dout(n15451),.clk(gclk));
	jor g15202(.dina(w_n15451_0[2]),.dinb(n15448),.dout(n15452),.clk(gclk));
	jand g15203(.dina(n15452),.dinb(w_n15447_0[1]),.dout(n15453),.clk(gclk));
	jor g15204(.dina(w_n15453_0[2]),.dinb(w_n3955_29[0]),.dout(n15454),.clk(gclk));
	jand g15205(.dina(w_n15453_0[1]),.dinb(w_n3955_28[2]),.dout(n15455),.clk(gclk));
	jxor g15206(.dina(w_n14841_0[0]),.dinb(w_n4249_31[1]),.dout(n15456),.clk(gclk));
	jor g15207(.dina(n15456),.dinb(w_n15260_33[0]),.dout(n15457),.clk(gclk));
	jxor g15208(.dina(n15457),.dinb(w_n14847_0[0]),.dout(n15458),.clk(gclk));
	jor g15209(.dina(w_n15458_0[2]),.dinb(n15455),.dout(n15459),.clk(gclk));
	jand g15210(.dina(n15459),.dinb(w_n15454_0[1]),.dout(n15460),.clk(gclk));
	jor g15211(.dina(w_n15460_0[2]),.dinb(w_n3642_32[1]),.dout(n15461),.clk(gclk));
	jand g15212(.dina(w_n15460_0[1]),.dinb(w_n3642_32[0]),.dout(n15462),.clk(gclk));
	jxor g15213(.dina(w_n14849_0[0]),.dinb(w_n3955_28[1]),.dout(n15463),.clk(gclk));
	jor g15214(.dina(n15463),.dinb(w_n15260_32[2]),.dout(n15464),.clk(gclk));
	jxor g15215(.dina(n15464),.dinb(w_n14855_0[0]),.dout(n15465),.clk(gclk));
	jor g15216(.dina(w_n15465_0[2]),.dinb(n15462),.dout(n15466),.clk(gclk));
	jand g15217(.dina(n15466),.dinb(w_n15461_0[1]),.dout(n15467),.clk(gclk));
	jor g15218(.dina(w_n15467_0[2]),.dinb(w_n3368_29[2]),.dout(n15468),.clk(gclk));
	jand g15219(.dina(w_n15467_0[1]),.dinb(w_n3368_29[1]),.dout(n15469),.clk(gclk));
	jxor g15220(.dina(w_n14857_0[0]),.dinb(w_n3642_31[2]),.dout(n15470),.clk(gclk));
	jor g15221(.dina(n15470),.dinb(w_n15260_32[1]),.dout(n15471),.clk(gclk));
	jxor g15222(.dina(n15471),.dinb(w_n15151_0[0]),.dout(n15472),.clk(gclk));
	jnot g15223(.din(w_n15472_0[2]),.dout(n15473),.clk(gclk));
	jor g15224(.dina(n15473),.dinb(n15469),.dout(n15474),.clk(gclk));
	jand g15225(.dina(n15474),.dinb(w_n15468_0[1]),.dout(n15475),.clk(gclk));
	jor g15226(.dina(w_n15475_0[2]),.dinb(w_n3089_33[0]),.dout(n15476),.clk(gclk));
	jand g15227(.dina(w_n15475_0[1]),.dinb(w_n3089_32[2]),.dout(n15477),.clk(gclk));
	jxor g15228(.dina(w_n14864_0[0]),.dinb(w_n3368_29[0]),.dout(n15478),.clk(gclk));
	jor g15229(.dina(n15478),.dinb(w_n15260_32[0]),.dout(n15479),.clk(gclk));
	jxor g15230(.dina(n15479),.dinb(w_n14870_0[0]),.dout(n15480),.clk(gclk));
	jor g15231(.dina(w_n15480_0[2]),.dinb(n15477),.dout(n15481),.clk(gclk));
	jand g15232(.dina(n15481),.dinb(w_n15476_0[1]),.dout(n15482),.clk(gclk));
	jor g15233(.dina(w_n15482_0[2]),.dinb(w_n2833_30[2]),.dout(n15483),.clk(gclk));
	jand g15234(.dina(w_n15482_0[1]),.dinb(w_n2833_30[1]),.dout(n15484),.clk(gclk));
	jxor g15235(.dina(w_n14872_0[0]),.dinb(w_n3089_32[1]),.dout(n15485),.clk(gclk));
	jor g15236(.dina(n15485),.dinb(w_n15260_31[2]),.dout(n15486),.clk(gclk));
	jxor g15237(.dina(n15486),.dinb(w_n15158_0[0]),.dout(n15487),.clk(gclk));
	jnot g15238(.din(w_n15487_0[2]),.dout(n15488),.clk(gclk));
	jor g15239(.dina(n15488),.dinb(n15484),.dout(n15489),.clk(gclk));
	jand g15240(.dina(n15489),.dinb(w_n15483_0[1]),.dout(n15490),.clk(gclk));
	jor g15241(.dina(w_n15490_0[2]),.dinb(w_n2572_33[1]),.dout(n15491),.clk(gclk));
	jand g15242(.dina(w_n15490_0[1]),.dinb(w_n2572_33[0]),.dout(n15492),.clk(gclk));
	jxor g15243(.dina(w_n14879_0[0]),.dinb(w_n2833_30[0]),.dout(n15493),.clk(gclk));
	jor g15244(.dina(n15493),.dinb(w_n15260_31[1]),.dout(n15494),.clk(gclk));
	jxor g15245(.dina(n15494),.dinb(w_n14885_0[0]),.dout(n15495),.clk(gclk));
	jor g15246(.dina(w_n15495_0[2]),.dinb(n15492),.dout(n15496),.clk(gclk));
	jand g15247(.dina(n15496),.dinb(w_n15491_0[1]),.dout(n15497),.clk(gclk));
	jor g15248(.dina(w_n15497_0[2]),.dinb(w_n2345_31[1]),.dout(n15498),.clk(gclk));
	jand g15249(.dina(w_n15497_0[1]),.dinb(w_n2345_31[0]),.dout(n15499),.clk(gclk));
	jxor g15250(.dina(w_n14887_0[0]),.dinb(w_n2572_32[2]),.dout(n15500),.clk(gclk));
	jor g15251(.dina(n15500),.dinb(w_n15260_31[0]),.dout(n15501),.clk(gclk));
	jxor g15252(.dina(n15501),.dinb(w_n14893_0[0]),.dout(n15502),.clk(gclk));
	jor g15253(.dina(w_n15502_0[2]),.dinb(n15499),.dout(n15503),.clk(gclk));
	jand g15254(.dina(n15503),.dinb(w_n15498_0[1]),.dout(n15504),.clk(gclk));
	jor g15255(.dina(w_n15504_0[2]),.dinb(w_n2108_34[0]),.dout(n15505),.clk(gclk));
	jand g15256(.dina(w_n15504_0[1]),.dinb(w_n2108_33[2]),.dout(n15506),.clk(gclk));
	jxor g15257(.dina(w_n14895_0[0]),.dinb(w_n2345_30[2]),.dout(n15507),.clk(gclk));
	jor g15258(.dina(n15507),.dinb(w_n15260_30[2]),.dout(n15508),.clk(gclk));
	jxor g15259(.dina(n15508),.dinb(w_n15168_0[0]),.dout(n15509),.clk(gclk));
	jnot g15260(.din(w_n15509_0[2]),.dout(n15510),.clk(gclk));
	jor g15261(.dina(n15510),.dinb(n15506),.dout(n15511),.clk(gclk));
	jand g15262(.dina(n15511),.dinb(w_n15505_0[1]),.dout(n15512),.clk(gclk));
	jor g15263(.dina(w_n15512_0[2]),.dinb(w_n1912_32[1]),.dout(n15513),.clk(gclk));
	jxor g15264(.dina(w_n14902_0[0]),.dinb(w_n2108_33[1]),.dout(n15514),.clk(gclk));
	jor g15265(.dina(n15514),.dinb(w_n15260_30[1]),.dout(n15515),.clk(gclk));
	jxor g15266(.dina(n15515),.dinb(w_n15033_0[0]),.dout(n15516),.clk(gclk));
	jnot g15267(.din(w_n15516_0[2]),.dout(n15517),.clk(gclk));
	jand g15268(.dina(w_n15512_0[1]),.dinb(w_n1912_32[0]),.dout(n15518),.clk(gclk));
	jor g15269(.dina(n15518),.dinb(n15517),.dout(n15519),.clk(gclk));
	jand g15270(.dina(n15519),.dinb(w_n15513_0[1]),.dout(n15520),.clk(gclk));
	jor g15271(.dina(w_n15520_0[2]),.dinb(w_n1699_34[2]),.dout(n15521),.clk(gclk));
	jand g15272(.dina(w_n15520_0[1]),.dinb(w_n1699_34[1]),.dout(n15522),.clk(gclk));
	jxor g15273(.dina(w_n14909_0[0]),.dinb(w_n1912_31[2]),.dout(n15523),.clk(gclk));
	jor g15274(.dina(n15523),.dinb(w_n15260_30[0]),.dout(n15524),.clk(gclk));
	jxor g15275(.dina(n15524),.dinb(w_n14915_0[0]),.dout(n15525),.clk(gclk));
	jor g15276(.dina(w_n15525_0[2]),.dinb(n15522),.dout(n15526),.clk(gclk));
	jand g15277(.dina(n15526),.dinb(w_n15521_0[1]),.dout(n15527),.clk(gclk));
	jor g15278(.dina(w_n15527_0[2]),.dinb(w_n1516_33[0]),.dout(n15528),.clk(gclk));
	jand g15279(.dina(w_n15527_0[1]),.dinb(w_n1516_32[2]),.dout(n15529),.clk(gclk));
	jxor g15280(.dina(w_n14917_0[0]),.dinb(w_n1699_34[0]),.dout(n15530),.clk(gclk));
	jor g15281(.dina(n15530),.dinb(w_n15260_29[2]),.dout(n15531),.clk(gclk));
	jxor g15282(.dina(n15531),.dinb(w_n15178_0[0]),.dout(n15532),.clk(gclk));
	jnot g15283(.din(w_n15532_0[2]),.dout(n15533),.clk(gclk));
	jor g15284(.dina(n15533),.dinb(n15529),.dout(n15534),.clk(gclk));
	jand g15285(.dina(n15534),.dinb(w_n15528_0[1]),.dout(n15535),.clk(gclk));
	jor g15286(.dina(w_n15535_0[2]),.dinb(w_n1332_34[2]),.dout(n15536),.clk(gclk));
	jand g15287(.dina(w_n15535_0[1]),.dinb(w_n1332_34[1]),.dout(n15537),.clk(gclk));
	jxor g15288(.dina(w_n14924_0[0]),.dinb(w_n1516_32[1]),.dout(n15538),.clk(gclk));
	jor g15289(.dina(n15538),.dinb(w_n15260_29[1]),.dout(n15539),.clk(gclk));
	jxor g15290(.dina(n15539),.dinb(w_n14930_0[0]),.dout(n15540),.clk(gclk));
	jor g15291(.dina(w_n15540_0[2]),.dinb(n15537),.dout(n15541),.clk(gclk));
	jand g15292(.dina(n15541),.dinb(w_n15536_0[1]),.dout(n15542),.clk(gclk));
	jor g15293(.dina(w_n15542_0[2]),.dinb(w_n1173_33[2]),.dout(n15543),.clk(gclk));
	jand g15294(.dina(w_n15542_0[1]),.dinb(w_n1173_33[1]),.dout(n15544),.clk(gclk));
	jxor g15295(.dina(w_n14932_0[0]),.dinb(w_n1332_34[0]),.dout(n15545),.clk(gclk));
	jor g15296(.dina(n15545),.dinb(w_n15260_29[0]),.dout(n15546),.clk(gclk));
	jxor g15297(.dina(n15546),.dinb(w_n15185_0[0]),.dout(n15547),.clk(gclk));
	jnot g15298(.din(w_n15547_0[2]),.dout(n15548),.clk(gclk));
	jor g15299(.dina(n15548),.dinb(n15544),.dout(n15549),.clk(gclk));
	jand g15300(.dina(n15549),.dinb(w_n15543_0[1]),.dout(n15550),.clk(gclk));
	jor g15301(.dina(w_n15550_0[2]),.dinb(w_n1008_35[2]),.dout(n15551),.clk(gclk));
	jand g15302(.dina(w_n15550_0[1]),.dinb(w_n1008_35[1]),.dout(n15552),.clk(gclk));
	jxor g15303(.dina(w_n14939_0[0]),.dinb(w_n1173_33[0]),.dout(n15553),.clk(gclk));
	jor g15304(.dina(n15553),.dinb(w_n15260_28[2]),.dout(n15554),.clk(gclk));
	jxor g15305(.dina(n15554),.dinb(w_n14945_0[0]),.dout(n15555),.clk(gclk));
	jor g15306(.dina(w_n15555_0[2]),.dinb(n15552),.dout(n15556),.clk(gclk));
	jand g15307(.dina(n15556),.dinb(w_n15551_0[1]),.dout(n15557),.clk(gclk));
	jor g15308(.dina(w_n15557_0[2]),.dinb(w_n884_34[2]),.dout(n15558),.clk(gclk));
	jand g15309(.dina(w_n15557_0[1]),.dinb(w_n884_34[1]),.dout(n15559),.clk(gclk));
	jxor g15310(.dina(w_n14947_0[0]),.dinb(w_n1008_35[0]),.dout(n15560),.clk(gclk));
	jor g15311(.dina(n15560),.dinb(w_n15260_28[1]),.dout(n15561),.clk(gclk));
	jxor g15312(.dina(n15561),.dinb(w_n14953_0[0]),.dout(n15562),.clk(gclk));
	jor g15313(.dina(w_n15562_0[2]),.dinb(n15559),.dout(n15563),.clk(gclk));
	jand g15314(.dina(n15563),.dinb(w_n15558_0[1]),.dout(n15564),.clk(gclk));
	jor g15315(.dina(w_n15564_0[2]),.dinb(w_n743_35[2]),.dout(n15565),.clk(gclk));
	jand g15316(.dina(w_n15564_0[1]),.dinb(w_n743_35[1]),.dout(n15566),.clk(gclk));
	jxor g15317(.dina(w_n14955_0[0]),.dinb(w_n884_34[0]),.dout(n15567),.clk(gclk));
	jor g15318(.dina(n15567),.dinb(w_n15260_28[0]),.dout(n15568),.clk(gclk));
	jxor g15319(.dina(n15568),.dinb(w_n14961_0[0]),.dout(n15569),.clk(gclk));
	jor g15320(.dina(w_n15569_0[2]),.dinb(n15566),.dout(n15570),.clk(gclk));
	jand g15321(.dina(n15570),.dinb(w_n15565_0[1]),.dout(n15571),.clk(gclk));
	jor g15322(.dina(w_n15571_0[2]),.dinb(w_n635_35[2]),.dout(n15572),.clk(gclk));
	jand g15323(.dina(w_n15571_0[1]),.dinb(w_n635_35[1]),.dout(n15573),.clk(gclk));
	jxor g15324(.dina(w_n14963_0[0]),.dinb(w_n743_35[0]),.dout(n15574),.clk(gclk));
	jor g15325(.dina(n15574),.dinb(w_n15260_27[2]),.dout(n15575),.clk(gclk));
	jxor g15326(.dina(n15575),.dinb(w_n15198_0[0]),.dout(n15576),.clk(gclk));
	jnot g15327(.din(w_n15576_0[2]),.dout(n15577),.clk(gclk));
	jor g15328(.dina(n15577),.dinb(n15573),.dout(n15578),.clk(gclk));
	jand g15329(.dina(n15578),.dinb(w_n15572_0[1]),.dout(n15579),.clk(gclk));
	jor g15330(.dina(w_n15579_0[2]),.dinb(w_n515_36[2]),.dout(n15580),.clk(gclk));
	jand g15331(.dina(w_n15579_0[1]),.dinb(w_n515_36[1]),.dout(n15581),.clk(gclk));
	jxor g15332(.dina(w_n14970_0[0]),.dinb(w_n635_35[0]),.dout(n15582),.clk(gclk));
	jor g15333(.dina(n15582),.dinb(w_n15260_27[1]),.dout(n15583),.clk(gclk));
	jxor g15334(.dina(n15583),.dinb(w_n14976_0[0]),.dout(n15584),.clk(gclk));
	jor g15335(.dina(w_n15584_0[2]),.dinb(n15581),.dout(n15585),.clk(gclk));
	jand g15336(.dina(n15585),.dinb(w_n15580_0[1]),.dout(n15586),.clk(gclk));
	jor g15337(.dina(w_n15586_0[2]),.dinb(w_n443_36[2]),.dout(n15587),.clk(gclk));
	jand g15338(.dina(w_n15586_0[1]),.dinb(w_n443_36[1]),.dout(n15588),.clk(gclk));
	jxor g15339(.dina(w_n14978_0[0]),.dinb(w_n515_36[0]),.dout(n15589),.clk(gclk));
	jor g15340(.dina(n15589),.dinb(w_n15260_27[0]),.dout(n15590),.clk(gclk));
	jxor g15341(.dina(n15590),.dinb(w_n15205_0[0]),.dout(n15591),.clk(gclk));
	jnot g15342(.din(w_n15591_0[2]),.dout(n15592),.clk(gclk));
	jor g15343(.dina(n15592),.dinb(n15588),.dout(n15593),.clk(gclk));
	jand g15344(.dina(n15593),.dinb(w_n15587_0[1]),.dout(n15594),.clk(gclk));
	jor g15345(.dina(w_n15594_0[2]),.dinb(w_n352_37[0]),.dout(n15595),.clk(gclk));
	jand g15346(.dina(w_n15594_0[1]),.dinb(w_n352_36[2]),.dout(n15596),.clk(gclk));
	jxor g15347(.dina(w_n14985_0[0]),.dinb(w_n443_36[0]),.dout(n15597),.clk(gclk));
	jor g15348(.dina(n15597),.dinb(w_n15260_26[2]),.dout(n15598),.clk(gclk));
	jxor g15349(.dina(n15598),.dinb(w_n14991_0[0]),.dout(n15599),.clk(gclk));
	jor g15350(.dina(w_n15599_0[2]),.dinb(n15596),.dout(n15600),.clk(gclk));
	jand g15351(.dina(n15600),.dinb(w_n15595_0[1]),.dout(n15601),.clk(gclk));
	jor g15352(.dina(w_n15601_0[2]),.dinb(w_n294_37[1]),.dout(n15602),.clk(gclk));
	jand g15353(.dina(w_n15601_0[1]),.dinb(w_n294_37[0]),.dout(n15603),.clk(gclk));
	jxor g15354(.dina(w_n14993_0[0]),.dinb(w_n352_36[1]),.dout(n15604),.clk(gclk));
	jor g15355(.dina(n15604),.dinb(w_n15260_26[1]),.dout(n15605),.clk(gclk));
	jxor g15356(.dina(n15605),.dinb(w_n15212_0[0]),.dout(n15606),.clk(gclk));
	jnot g15357(.din(w_n15606_0[2]),.dout(n15607),.clk(gclk));
	jor g15358(.dina(n15607),.dinb(n15603),.dout(n15608),.clk(gclk));
	jand g15359(.dina(n15608),.dinb(w_n15602_0[1]),.dout(n15609),.clk(gclk));
	jor g15360(.dina(w_n15609_0[2]),.dinb(w_n239_37[1]),.dout(n15610),.clk(gclk));
	jand g15361(.dina(w_n15609_0[1]),.dinb(w_n239_37[0]),.dout(n15611),.clk(gclk));
	jxor g15362(.dina(w_n15000_0[0]),.dinb(w_n294_36[2]),.dout(n15612),.clk(gclk));
	jor g15363(.dina(n15612),.dinb(w_n15260_26[0]),.dout(n15613),.clk(gclk));
	jxor g15364(.dina(n15613),.dinb(w_n15006_0[0]),.dout(n15614),.clk(gclk));
	jor g15365(.dina(w_n15614_0[2]),.dinb(n15611),.dout(n15615),.clk(gclk));
	jand g15366(.dina(n15615),.dinb(w_n15610_0[1]),.dout(n15616),.clk(gclk));
	jor g15367(.dina(w_n15616_0[2]),.dinb(w_n221_37[1]),.dout(n15617),.clk(gclk));
	jand g15368(.dina(w_n15616_0[1]),.dinb(w_n221_37[0]),.dout(n15618),.clk(gclk));
	jxor g15369(.dina(w_n15008_0[0]),.dinb(w_n239_36[2]),.dout(n15619),.clk(gclk));
	jor g15370(.dina(n15619),.dinb(w_n15260_25[2]),.dout(n15620),.clk(gclk));
	jxor g15371(.dina(n15620),.dinb(w_n15219_0[0]),.dout(n15621),.clk(gclk));
	jnot g15372(.din(w_n15621_0[1]),.dout(n15622),.clk(gclk));
	jor g15373(.dina(w_n15622_0[1]),.dinb(n15618),.dout(n15623),.clk(gclk));
	jand g15374(.dina(n15623),.dinb(w_n15617_0[1]),.dout(n15624),.clk(gclk));
	jor g15375(.dina(w_n15624_0[2]),.dinb(w_n15264_0[2]),.dout(n15625),.clk(gclk));
	jand g15376(.dina(w_asqrt15_11[2]),.dinb(w_n15251_0[0]),.dout(n15626),.clk(gclk));
	jor g15377(.dina(w_n15626_0[1]),.dinb(w_n15625_0[1]),.dout(n15627),.clk(gclk));
	jor g15378(.dina(n15627),.dinb(w_n15239_0[0]),.dout(n15628),.clk(gclk));
	jand g15379(.dina(n15628),.dinb(w_n218_15[2]),.dout(n15629),.clk(gclk));
	jand g15380(.dina(w_n15260_25[1]),.dinb(w_n15231_0[1]),.dout(n15630),.clk(gclk));
	jand g15381(.dina(w_n15624_0[1]),.dinb(w_n15264_0[1]),.dout(n15631),.clk(gclk));
	jor g15382(.dina(w_n15631_0[2]),.dinb(n15630),.dout(n15632),.clk(gclk));
	jand g15383(.dina(w_n15260_25[0]),.dinb(w_n15228_0[0]),.dout(n15633),.clk(gclk));
	jand g15384(.dina(w_n15232_0[0]),.dinb(w_asqrt63_27[1]),.dout(n15634),.clk(gclk));
	jand g15385(.dina(n15634),.dinb(w_n15256_0[1]),.dout(n15635),.clk(gclk));
	jnot g15386(.din(n15635),.dout(n15636),.clk(gclk));
	jor g15387(.dina(w_n15636_0[1]),.dinb(n15633),.dout(n15637),.clk(gclk));
	jnot g15388(.din(n15637),.dout(n15638),.clk(gclk));
	jor g15389(.dina(n15638),.dinb(n15632),.dout(n15639),.clk(gclk));
	jor g15390(.dina(w_n15639_0[1]),.dinb(n15629),.dout(asqrt_fa_15),.clk(gclk));
	jand g15391(.dina(w_asqrt14_34),.dinb(w_a28_0[1]),.dout(n15641),.clk(gclk));
	jnot g15392(.din(w_a26_1[1]),.dout(n15642),.clk(gclk));
	jnot g15393(.din(w_a27_0[1]),.dout(n15643),.clk(gclk));
	jand g15394(.dina(w_n15643_0[1]),.dinb(w_n15642_1[1]),.dout(n15644),.clk(gclk));
	jand g15395(.dina(w_n15644_0[2]),.dinb(w_n15265_1[1]),.dout(n15645),.clk(gclk));
	jor g15396(.dina(w_n15645_0[1]),.dinb(n15641),.dout(n15646),.clk(gclk));
	jand g15397(.dina(w_n15646_0[2]),.dinb(w_asqrt15_11[1]),.dout(n15647),.clk(gclk));
	jor g15398(.dina(w_n15646_0[1]),.dinb(w_asqrt15_11[0]),.dout(n15648),.clk(gclk));
	jand g15399(.dina(w_asqrt14_33[2]),.dinb(w_n15265_1[0]),.dout(n15649),.clk(gclk));
	jor g15400(.dina(n15649),.dinb(w_n15266_0[0]),.dout(n15650),.clk(gclk));
	jnot g15401(.din(w_n15267_0[1]),.dout(n15651),.clk(gclk));
	jnot g15402(.din(w_n15617_0[0]),.dout(n15652),.clk(gclk));
	jnot g15403(.din(w_n15610_0[0]),.dout(n15653),.clk(gclk));
	jnot g15404(.din(w_n15602_0[0]),.dout(n15654),.clk(gclk));
	jnot g15405(.din(w_n15595_0[0]),.dout(n15655),.clk(gclk));
	jnot g15406(.din(w_n15587_0[0]),.dout(n15656),.clk(gclk));
	jnot g15407(.din(w_n15580_0[0]),.dout(n15657),.clk(gclk));
	jnot g15408(.din(w_n15572_0[0]),.dout(n15658),.clk(gclk));
	jnot g15409(.din(w_n15565_0[0]),.dout(n15659),.clk(gclk));
	jnot g15410(.din(w_n15558_0[0]),.dout(n15660),.clk(gclk));
	jnot g15411(.din(w_n15551_0[0]),.dout(n15661),.clk(gclk));
	jnot g15412(.din(w_n15543_0[0]),.dout(n15662),.clk(gclk));
	jnot g15413(.din(w_n15536_0[0]),.dout(n15663),.clk(gclk));
	jnot g15414(.din(w_n15528_0[0]),.dout(n15664),.clk(gclk));
	jnot g15415(.din(w_n15521_0[0]),.dout(n15665),.clk(gclk));
	jnot g15416(.din(w_n15513_0[0]),.dout(n15666),.clk(gclk));
	jnot g15417(.din(w_n15505_0[0]),.dout(n15667),.clk(gclk));
	jnot g15418(.din(w_n15498_0[0]),.dout(n15668),.clk(gclk));
	jnot g15419(.din(w_n15491_0[0]),.dout(n15669),.clk(gclk));
	jnot g15420(.din(w_n15483_0[0]),.dout(n15670),.clk(gclk));
	jnot g15421(.din(w_n15476_0[0]),.dout(n15671),.clk(gclk));
	jnot g15422(.din(w_n15468_0[0]),.dout(n15672),.clk(gclk));
	jnot g15423(.din(w_n15461_0[0]),.dout(n15673),.clk(gclk));
	jnot g15424(.din(w_n15454_0[0]),.dout(n15674),.clk(gclk));
	jnot g15425(.din(w_n15447_0[0]),.dout(n15675),.clk(gclk));
	jnot g15426(.din(w_n15439_0[0]),.dout(n15676),.clk(gclk));
	jnot g15427(.din(w_n15432_0[0]),.dout(n15677),.clk(gclk));
	jnot g15428(.din(w_n15424_0[0]),.dout(n15678),.clk(gclk));
	jnot g15429(.din(w_n15417_0[0]),.dout(n15679),.clk(gclk));
	jnot g15430(.din(w_n15410_0[0]),.dout(n15680),.clk(gclk));
	jnot g15431(.din(w_n15403_0[0]),.dout(n15681),.clk(gclk));
	jnot g15432(.din(w_n15395_0[0]),.dout(n15682),.clk(gclk));
	jnot g15433(.din(w_n15388_0[0]),.dout(n15683),.clk(gclk));
	jnot g15434(.din(w_n15380_0[0]),.dout(n15684),.clk(gclk));
	jnot g15435(.din(w_n15373_0[0]),.dout(n15685),.clk(gclk));
	jnot g15436(.din(w_n15365_0[0]),.dout(n15686),.clk(gclk));
	jnot g15437(.din(w_n15358_0[0]),.dout(n15687),.clk(gclk));
	jnot g15438(.din(w_n15350_0[0]),.dout(n15688),.clk(gclk));
	jnot g15439(.din(w_n15343_0[0]),.dout(n15689),.clk(gclk));
	jnot g15440(.din(w_n15336_0[0]),.dout(n15690),.clk(gclk));
	jnot g15441(.din(w_n15329_0[0]),.dout(n15691),.clk(gclk));
	jnot g15442(.din(w_n15321_0[0]),.dout(n15692),.clk(gclk));
	jnot g15443(.din(w_n15314_0[0]),.dout(n15693),.clk(gclk));
	jnot g15444(.din(w_n15306_0[0]),.dout(n15694),.clk(gclk));
	jnot g15445(.din(w_n15299_0[0]),.dout(n15695),.clk(gclk));
	jnot g15446(.din(w_n15291_0[0]),.dout(n15696),.clk(gclk));
	jnot g15447(.din(w_n15280_0[0]),.dout(n15697),.clk(gclk));
	jnot g15448(.din(w_n15272_0[0]),.dout(n15698),.clk(gclk));
	jand g15449(.dina(w_asqrt15_10[2]),.dinb(w_a30_0[2]),.dout(n15699),.clk(gclk));
	jor g15450(.dina(n15699),.dinb(w_n15268_0[0]),.dout(n15700),.clk(gclk));
	jor g15451(.dina(n15700),.dinb(w_asqrt16_18[0]),.dout(n15701),.clk(gclk));
	jand g15452(.dina(w_asqrt15_10[1]),.dinb(w_n14443_0[1]),.dout(n15702),.clk(gclk));
	jor g15453(.dina(n15702),.dinb(w_n14444_0[0]),.dout(n15703),.clk(gclk));
	jand g15454(.dina(w_n15283_0[0]),.dinb(n15703),.dout(n15704),.clk(gclk));
	jand g15455(.dina(w_n15704_0[1]),.dinb(n15701),.dout(n15705),.clk(gclk));
	jor g15456(.dina(n15705),.dinb(n15698),.dout(n15706),.clk(gclk));
	jor g15457(.dina(n15706),.dinb(w_asqrt17_11[0]),.dout(n15707),.clk(gclk));
	jnot g15458(.din(w_n15288_0[0]),.dout(n15708),.clk(gclk));
	jand g15459(.dina(w_n15708_0[1]),.dinb(n15707),.dout(n15709),.clk(gclk));
	jor g15460(.dina(n15709),.dinb(n15697),.dout(n15710),.clk(gclk));
	jor g15461(.dina(n15710),.dinb(w_asqrt18_18[1]),.dout(n15711),.clk(gclk));
	jand g15462(.dina(w_n15295_0[1]),.dinb(n15711),.dout(n15712),.clk(gclk));
	jor g15463(.dina(n15712),.dinb(n15696),.dout(n15713),.clk(gclk));
	jor g15464(.dina(n15713),.dinb(w_asqrt19_11[1]),.dout(n15714),.clk(gclk));
	jnot g15465(.din(w_n15303_0[1]),.dout(n15715),.clk(gclk));
	jand g15466(.dina(n15715),.dinb(n15714),.dout(n15716),.clk(gclk));
	jor g15467(.dina(n15716),.dinb(n15695),.dout(n15717),.clk(gclk));
	jor g15468(.dina(n15717),.dinb(w_asqrt20_18[1]),.dout(n15718),.clk(gclk));
	jand g15469(.dina(w_n15310_0[1]),.dinb(n15718),.dout(n15719),.clk(gclk));
	jor g15470(.dina(n15719),.dinb(n15694),.dout(n15720),.clk(gclk));
	jor g15471(.dina(n15720),.dinb(w_asqrt21_12[0]),.dout(n15721),.clk(gclk));
	jnot g15472(.din(w_n15318_0[1]),.dout(n15722),.clk(gclk));
	jand g15473(.dina(n15722),.dinb(n15721),.dout(n15723),.clk(gclk));
	jor g15474(.dina(n15723),.dinb(n15693),.dout(n15724),.clk(gclk));
	jor g15475(.dina(n15724),.dinb(w_asqrt22_18[2]),.dout(n15725),.clk(gclk));
	jand g15476(.dina(w_n15325_0[1]),.dinb(n15725),.dout(n15726),.clk(gclk));
	jor g15477(.dina(n15726),.dinb(n15692),.dout(n15727),.clk(gclk));
	jor g15478(.dina(n15727),.dinb(w_asqrt23_12[2]),.dout(n15728),.clk(gclk));
	jnot g15479(.din(w_n15333_0[1]),.dout(n15729),.clk(gclk));
	jand g15480(.dina(n15729),.dinb(n15728),.dout(n15730),.clk(gclk));
	jor g15481(.dina(n15730),.dinb(n15691),.dout(n15731),.clk(gclk));
	jor g15482(.dina(n15731),.dinb(w_asqrt24_18[2]),.dout(n15732),.clk(gclk));
	jnot g15483(.din(w_n15340_0[1]),.dout(n15733),.clk(gclk));
	jand g15484(.dina(n15733),.dinb(n15732),.dout(n15734),.clk(gclk));
	jor g15485(.dina(n15734),.dinb(n15690),.dout(n15735),.clk(gclk));
	jor g15486(.dina(n15735),.dinb(w_asqrt25_12[2]),.dout(n15736),.clk(gclk));
	jnot g15487(.din(w_n15347_0[1]),.dout(n15737),.clk(gclk));
	jand g15488(.dina(n15737),.dinb(n15736),.dout(n15738),.clk(gclk));
	jor g15489(.dina(n15738),.dinb(n15689),.dout(n15739),.clk(gclk));
	jor g15490(.dina(n15739),.dinb(w_asqrt26_18[2]),.dout(n15740),.clk(gclk));
	jand g15491(.dina(w_n15354_0[1]),.dinb(n15740),.dout(n15741),.clk(gclk));
	jor g15492(.dina(n15741),.dinb(n15688),.dout(n15742),.clk(gclk));
	jor g15493(.dina(n15742),.dinb(w_asqrt27_13[1]),.dout(n15743),.clk(gclk));
	jnot g15494(.din(w_n15362_0[1]),.dout(n15744),.clk(gclk));
	jand g15495(.dina(n15744),.dinb(n15743),.dout(n15745),.clk(gclk));
	jor g15496(.dina(n15745),.dinb(n15687),.dout(n15746),.clk(gclk));
	jor g15497(.dina(n15746),.dinb(w_asqrt28_19[0]),.dout(n15747),.clk(gclk));
	jand g15498(.dina(w_n15369_0[1]),.dinb(n15747),.dout(n15748),.clk(gclk));
	jor g15499(.dina(n15748),.dinb(n15686),.dout(n15749),.clk(gclk));
	jor g15500(.dina(n15749),.dinb(w_asqrt29_13[2]),.dout(n15750),.clk(gclk));
	jnot g15501(.din(w_n15377_0[1]),.dout(n15751),.clk(gclk));
	jand g15502(.dina(n15751),.dinb(n15750),.dout(n15752),.clk(gclk));
	jor g15503(.dina(n15752),.dinb(n15685),.dout(n15753),.clk(gclk));
	jor g15504(.dina(n15753),.dinb(w_asqrt30_19[1]),.dout(n15754),.clk(gclk));
	jand g15505(.dina(w_n15384_0[1]),.dinb(n15754),.dout(n15755),.clk(gclk));
	jor g15506(.dina(n15755),.dinb(n15684),.dout(n15756),.clk(gclk));
	jor g15507(.dina(n15756),.dinb(w_asqrt31_14[1]),.dout(n15757),.clk(gclk));
	jnot g15508(.din(w_n15392_0[1]),.dout(n15758),.clk(gclk));
	jand g15509(.dina(n15758),.dinb(n15757),.dout(n15759),.clk(gclk));
	jor g15510(.dina(n15759),.dinb(n15683),.dout(n15760),.clk(gclk));
	jor g15511(.dina(n15760),.dinb(w_asqrt32_19[1]),.dout(n15761),.clk(gclk));
	jand g15512(.dina(w_n15399_0[1]),.dinb(n15761),.dout(n15762),.clk(gclk));
	jor g15513(.dina(n15762),.dinb(n15682),.dout(n15763),.clk(gclk));
	jor g15514(.dina(n15763),.dinb(w_asqrt33_15[0]),.dout(n15764),.clk(gclk));
	jnot g15515(.din(w_n15407_0[1]),.dout(n15765),.clk(gclk));
	jand g15516(.dina(n15765),.dinb(n15764),.dout(n15766),.clk(gclk));
	jor g15517(.dina(n15766),.dinb(n15681),.dout(n15767),.clk(gclk));
	jor g15518(.dina(n15767),.dinb(w_asqrt34_19[2]),.dout(n15768),.clk(gclk));
	jnot g15519(.din(w_n15414_0[1]),.dout(n15769),.clk(gclk));
	jand g15520(.dina(n15769),.dinb(n15768),.dout(n15770),.clk(gclk));
	jor g15521(.dina(n15770),.dinb(n15680),.dout(n15771),.clk(gclk));
	jor g15522(.dina(n15771),.dinb(w_asqrt35_15[2]),.dout(n15772),.clk(gclk));
	jnot g15523(.din(w_n15421_0[1]),.dout(n15773),.clk(gclk));
	jand g15524(.dina(n15773),.dinb(n15772),.dout(n15774),.clk(gclk));
	jor g15525(.dina(n15774),.dinb(n15679),.dout(n15775),.clk(gclk));
	jor g15526(.dina(n15775),.dinb(w_asqrt36_19[2]),.dout(n15776),.clk(gclk));
	jand g15527(.dina(w_n15428_0[1]),.dinb(n15776),.dout(n15777),.clk(gclk));
	jor g15528(.dina(n15777),.dinb(n15678),.dout(n15778),.clk(gclk));
	jor g15529(.dina(n15778),.dinb(w_asqrt37_16[0]),.dout(n15779),.clk(gclk));
	jnot g15530(.din(w_n15436_0[1]),.dout(n15780),.clk(gclk));
	jand g15531(.dina(n15780),.dinb(n15779),.dout(n15781),.clk(gclk));
	jor g15532(.dina(n15781),.dinb(n15677),.dout(n15782),.clk(gclk));
	jor g15533(.dina(n15782),.dinb(w_asqrt38_20[0]),.dout(n15783),.clk(gclk));
	jand g15534(.dina(w_n15443_0[1]),.dinb(n15783),.dout(n15784),.clk(gclk));
	jor g15535(.dina(n15784),.dinb(n15676),.dout(n15785),.clk(gclk));
	jor g15536(.dina(n15785),.dinb(w_asqrt39_16[2]),.dout(n15786),.clk(gclk));
	jnot g15537(.din(w_n15451_0[1]),.dout(n15787),.clk(gclk));
	jand g15538(.dina(n15787),.dinb(n15786),.dout(n15788),.clk(gclk));
	jor g15539(.dina(n15788),.dinb(n15675),.dout(n15789),.clk(gclk));
	jor g15540(.dina(n15789),.dinb(w_asqrt40_20[0]),.dout(n15790),.clk(gclk));
	jnot g15541(.din(w_n15458_0[1]),.dout(n15791),.clk(gclk));
	jand g15542(.dina(n15791),.dinb(n15790),.dout(n15792),.clk(gclk));
	jor g15543(.dina(n15792),.dinb(n15674),.dout(n15793),.clk(gclk));
	jor g15544(.dina(n15793),.dinb(w_asqrt41_17[0]),.dout(n15794),.clk(gclk));
	jnot g15545(.din(w_n15465_0[1]),.dout(n15795),.clk(gclk));
	jand g15546(.dina(n15795),.dinb(n15794),.dout(n15796),.clk(gclk));
	jor g15547(.dina(n15796),.dinb(n15673),.dout(n15797),.clk(gclk));
	jor g15548(.dina(n15797),.dinb(w_asqrt42_20[1]),.dout(n15798),.clk(gclk));
	jand g15549(.dina(w_n15472_0[1]),.dinb(n15798),.dout(n15799),.clk(gclk));
	jor g15550(.dina(n15799),.dinb(n15672),.dout(n15800),.clk(gclk));
	jor g15551(.dina(n15800),.dinb(w_asqrt43_17[1]),.dout(n15801),.clk(gclk));
	jnot g15552(.din(w_n15480_0[1]),.dout(n15802),.clk(gclk));
	jand g15553(.dina(n15802),.dinb(n15801),.dout(n15803),.clk(gclk));
	jor g15554(.dina(n15803),.dinb(n15671),.dout(n15804),.clk(gclk));
	jor g15555(.dina(n15804),.dinb(w_asqrt44_20[1]),.dout(n15805),.clk(gclk));
	jand g15556(.dina(w_n15487_0[1]),.dinb(n15805),.dout(n15806),.clk(gclk));
	jor g15557(.dina(n15806),.dinb(n15670),.dout(n15807),.clk(gclk));
	jor g15558(.dina(n15807),.dinb(w_asqrt45_18[0]),.dout(n15808),.clk(gclk));
	jnot g15559(.din(w_n15495_0[1]),.dout(n15809),.clk(gclk));
	jand g15560(.dina(n15809),.dinb(n15808),.dout(n15810),.clk(gclk));
	jor g15561(.dina(n15810),.dinb(n15669),.dout(n15811),.clk(gclk));
	jor g15562(.dina(n15811),.dinb(w_asqrt46_20[1]),.dout(n15812),.clk(gclk));
	jnot g15563(.din(w_n15502_0[1]),.dout(n15813),.clk(gclk));
	jand g15564(.dina(n15813),.dinb(n15812),.dout(n15814),.clk(gclk));
	jor g15565(.dina(n15814),.dinb(n15668),.dout(n15815),.clk(gclk));
	jor g15566(.dina(n15815),.dinb(w_asqrt47_18[2]),.dout(n15816),.clk(gclk));
	jand g15567(.dina(w_n15509_0[1]),.dinb(n15816),.dout(n15817),.clk(gclk));
	jor g15568(.dina(n15817),.dinb(n15667),.dout(n15818),.clk(gclk));
	jor g15569(.dina(n15818),.dinb(w_asqrt48_20[2]),.dout(n15819),.clk(gclk));
	jand g15570(.dina(n15819),.dinb(w_n15516_0[1]),.dout(n15820),.clk(gclk));
	jor g15571(.dina(n15820),.dinb(n15666),.dout(n15821),.clk(gclk));
	jor g15572(.dina(n15821),.dinb(w_asqrt49_19[0]),.dout(n15822),.clk(gclk));
	jnot g15573(.din(w_n15525_0[1]),.dout(n15823),.clk(gclk));
	jand g15574(.dina(n15823),.dinb(n15822),.dout(n15824),.clk(gclk));
	jor g15575(.dina(n15824),.dinb(n15665),.dout(n15825),.clk(gclk));
	jor g15576(.dina(n15825),.dinb(w_asqrt50_21[0]),.dout(n15826),.clk(gclk));
	jand g15577(.dina(w_n15532_0[1]),.dinb(n15826),.dout(n15827),.clk(gclk));
	jor g15578(.dina(n15827),.dinb(n15664),.dout(n15828),.clk(gclk));
	jor g15579(.dina(n15828),.dinb(w_asqrt51_19[1]),.dout(n15829),.clk(gclk));
	jnot g15580(.din(w_n15540_0[1]),.dout(n15830),.clk(gclk));
	jand g15581(.dina(n15830),.dinb(n15829),.dout(n15831),.clk(gclk));
	jor g15582(.dina(n15831),.dinb(n15663),.dout(n15832),.clk(gclk));
	jor g15583(.dina(n15832),.dinb(w_asqrt52_21[0]),.dout(n15833),.clk(gclk));
	jand g15584(.dina(w_n15547_0[1]),.dinb(n15833),.dout(n15834),.clk(gclk));
	jor g15585(.dina(n15834),.dinb(n15662),.dout(n15835),.clk(gclk));
	jor g15586(.dina(n15835),.dinb(w_asqrt53_20[0]),.dout(n15836),.clk(gclk));
	jnot g15587(.din(w_n15555_0[1]),.dout(n15837),.clk(gclk));
	jand g15588(.dina(n15837),.dinb(n15836),.dout(n15838),.clk(gclk));
	jor g15589(.dina(n15838),.dinb(n15661),.dout(n15839),.clk(gclk));
	jor g15590(.dina(n15839),.dinb(w_asqrt54_21[0]),.dout(n15840),.clk(gclk));
	jnot g15591(.din(w_n15562_0[1]),.dout(n15841),.clk(gclk));
	jand g15592(.dina(n15841),.dinb(n15840),.dout(n15842),.clk(gclk));
	jor g15593(.dina(n15842),.dinb(n15660),.dout(n15843),.clk(gclk));
	jor g15594(.dina(n15843),.dinb(w_asqrt55_20[1]),.dout(n15844),.clk(gclk));
	jnot g15595(.din(w_n15569_0[1]),.dout(n15845),.clk(gclk));
	jand g15596(.dina(n15845),.dinb(n15844),.dout(n15846),.clk(gclk));
	jor g15597(.dina(n15846),.dinb(n15659),.dout(n15847),.clk(gclk));
	jor g15598(.dina(n15847),.dinb(w_asqrt56_21[1]),.dout(n15848),.clk(gclk));
	jand g15599(.dina(w_n15576_0[1]),.dinb(n15848),.dout(n15849),.clk(gclk));
	jor g15600(.dina(n15849),.dinb(n15658),.dout(n15850),.clk(gclk));
	jor g15601(.dina(n15850),.dinb(w_asqrt57_21[0]),.dout(n15851),.clk(gclk));
	jnot g15602(.din(w_n15584_0[1]),.dout(n15852),.clk(gclk));
	jand g15603(.dina(n15852),.dinb(n15851),.dout(n15853),.clk(gclk));
	jor g15604(.dina(n15853),.dinb(n15657),.dout(n15854),.clk(gclk));
	jor g15605(.dina(n15854),.dinb(w_asqrt58_21[2]),.dout(n15855),.clk(gclk));
	jand g15606(.dina(w_n15591_0[1]),.dinb(n15855),.dout(n15856),.clk(gclk));
	jor g15607(.dina(n15856),.dinb(n15656),.dout(n15857),.clk(gclk));
	jor g15608(.dina(n15857),.dinb(w_asqrt59_21[1]),.dout(n15858),.clk(gclk));
	jnot g15609(.din(w_n15599_0[1]),.dout(n15859),.clk(gclk));
	jand g15610(.dina(n15859),.dinb(n15858),.dout(n15860),.clk(gclk));
	jor g15611(.dina(n15860),.dinb(n15655),.dout(n15861),.clk(gclk));
	jor g15612(.dina(n15861),.dinb(w_asqrt60_21[2]),.dout(n15862),.clk(gclk));
	jand g15613(.dina(w_n15606_0[1]),.dinb(n15862),.dout(n15863),.clk(gclk));
	jor g15614(.dina(n15863),.dinb(n15654),.dout(n15864),.clk(gclk));
	jor g15615(.dina(n15864),.dinb(w_asqrt61_21[2]),.dout(n15865),.clk(gclk));
	jnot g15616(.din(w_n15614_0[1]),.dout(n15866),.clk(gclk));
	jand g15617(.dina(n15866),.dinb(n15865),.dout(n15867),.clk(gclk));
	jor g15618(.dina(n15867),.dinb(n15653),.dout(n15868),.clk(gclk));
	jor g15619(.dina(n15868),.dinb(w_asqrt62_21[2]),.dout(n15869),.clk(gclk));
	jand g15620(.dina(w_n15621_0[0]),.dinb(n15869),.dout(n15870),.clk(gclk));
	jor g15621(.dina(n15870),.dinb(n15652),.dout(n15871),.clk(gclk));
	jand g15622(.dina(n15871),.dinb(w_n15263_0[0]),.dout(n15872),.clk(gclk));
	jnot g15623(.din(w_n15626_0[0]),.dout(n15873),.clk(gclk));
	jand g15624(.dina(n15873),.dinb(w_n15872_0[1]),.dout(n15874),.clk(gclk));
	jand g15625(.dina(n15874),.dinb(w_n15256_0[0]),.dout(n15875),.clk(gclk));
	jor g15626(.dina(n15875),.dinb(w_asqrt63_27[0]),.dout(n15876),.clk(gclk));
	jnot g15627(.din(w_n15639_0[0]),.dout(n15877),.clk(gclk));
	jand g15628(.dina(n15877),.dinb(w_n15876_0[1]),.dout(n15878),.clk(gclk));
	jor g15629(.dina(w_n15878_18[1]),.dinb(n15651),.dout(n15879),.clk(gclk));
	jand g15630(.dina(n15879),.dinb(n15650),.dout(n15880),.clk(gclk));
	jand g15631(.dina(n15880),.dinb(n15648),.dout(n15881),.clk(gclk));
	jor g15632(.dina(n15881),.dinb(w_n15647_0[1]),.dout(n15882),.clk(gclk));
	jand g15633(.dina(w_n15882_0[2]),.dinb(w_asqrt16_17[2]),.dout(n15883),.clk(gclk));
	jor g15634(.dina(w_n15882_0[1]),.dinb(w_asqrt16_17[1]),.dout(n15884),.clk(gclk));
	jand g15635(.dina(w_asqrt14_33[1]),.dinb(w_n15267_0[0]),.dout(n15885),.clk(gclk));
	jnot g15636(.din(w_n15631_0[1]),.dout(n15886),.clk(gclk));
	jand g15637(.dina(w_n15636_0[0]),.dinb(w_asqrt15_10[0]),.dout(n15887),.clk(gclk));
	jand g15638(.dina(n15887),.dinb(w_n15886_0[1]),.dout(n15888),.clk(gclk));
	jand g15639(.dina(n15888),.dinb(w_n15876_0[0]),.dout(n15889),.clk(gclk));
	jor g15640(.dina(n15889),.dinb(w_n15885_0[1]),.dout(n15890),.clk(gclk));
	jxor g15641(.dina(n15890),.dinb(w_a30_0[1]),.dout(n15891),.clk(gclk));
	jnot g15642(.din(w_n15891_0[1]),.dout(n15892),.clk(gclk));
	jand g15643(.dina(w_n15892_0[1]),.dinb(n15884),.dout(n15893),.clk(gclk));
	jor g15644(.dina(n15893),.dinb(w_n15883_0[1]),.dout(n15894),.clk(gclk));
	jand g15645(.dina(w_n15894_0[2]),.dinb(w_asqrt17_10[2]),.dout(n15895),.clk(gclk));
	jor g15646(.dina(w_n15894_0[1]),.dinb(w_asqrt17_10[1]),.dout(n15896),.clk(gclk));
	jxor g15647(.dina(w_n15271_0[0]),.dinb(w_n14674_18[0]),.dout(n15897),.clk(gclk));
	jand g15648(.dina(n15897),.dinb(w_asqrt14_33[0]),.dout(n15898),.clk(gclk));
	jxor g15649(.dina(n15898),.dinb(w_n15704_0[0]),.dout(n15899),.clk(gclk));
	jand g15650(.dina(w_n15899_0[2]),.dinb(n15896),.dout(n15900),.clk(gclk));
	jor g15651(.dina(n15900),.dinb(w_n15895_0[1]),.dout(n15901),.clk(gclk));
	jand g15652(.dina(w_n15901_0[2]),.dinb(w_asqrt18_18[0]),.dout(n15902),.clk(gclk));
	jor g15653(.dina(w_n15901_0[1]),.dinb(w_asqrt18_17[2]),.dout(n15903),.clk(gclk));
	jxor g15654(.dina(w_n15279_0[0]),.dinb(w_n14078_25[1]),.dout(n15904),.clk(gclk));
	jand g15655(.dina(n15904),.dinb(w_asqrt14_32[2]),.dout(n15905),.clk(gclk));
	jxor g15656(.dina(n15905),.dinb(w_n15708_0[0]),.dout(n15906),.clk(gclk));
	jand g15657(.dina(w_n15906_0[1]),.dinb(n15903),.dout(n15907),.clk(gclk));
	jor g15658(.dina(n15907),.dinb(w_n15902_0[1]),.dout(n15908),.clk(gclk));
	jand g15659(.dina(w_n15908_0[2]),.dinb(w_asqrt19_11[0]),.dout(n15909),.clk(gclk));
	jor g15660(.dina(w_n15908_0[1]),.dinb(w_asqrt19_10[2]),.dout(n15910),.clk(gclk));
	jxor g15661(.dina(w_n15290_0[0]),.dinb(w_n13515_19[0]),.dout(n15911),.clk(gclk));
	jand g15662(.dina(n15911),.dinb(w_asqrt14_32[1]),.dout(n15912),.clk(gclk));
	jxor g15663(.dina(n15912),.dinb(w_n15295_0[0]),.dout(n15913),.clk(gclk));
	jand g15664(.dina(w_n15913_0[1]),.dinb(n15910),.dout(n15914),.clk(gclk));
	jor g15665(.dina(n15914),.dinb(w_n15909_0[1]),.dout(n15915),.clk(gclk));
	jand g15666(.dina(w_n15915_0[2]),.dinb(w_asqrt20_18[0]),.dout(n15916),.clk(gclk));
	jor g15667(.dina(w_n15915_0[1]),.dinb(w_asqrt20_17[2]),.dout(n15917),.clk(gclk));
	jxor g15668(.dina(w_n15298_0[0]),.dinb(w_n12947_26[0]),.dout(n15918),.clk(gclk));
	jand g15669(.dina(n15918),.dinb(w_asqrt14_32[0]),.dout(n15919),.clk(gclk));
	jxor g15670(.dina(n15919),.dinb(w_n15303_0[0]),.dout(n15920),.clk(gclk));
	jnot g15671(.din(w_n15920_0[1]),.dout(n15921),.clk(gclk));
	jand g15672(.dina(w_n15921_0[1]),.dinb(n15917),.dout(n15922),.clk(gclk));
	jor g15673(.dina(n15922),.dinb(w_n15916_0[1]),.dout(n15923),.clk(gclk));
	jand g15674(.dina(w_n15923_0[2]),.dinb(w_asqrt21_11[2]),.dout(n15924),.clk(gclk));
	jor g15675(.dina(w_n15923_0[1]),.dinb(w_asqrt21_11[1]),.dout(n15925),.clk(gclk));
	jxor g15676(.dina(w_n15305_0[0]),.dinb(w_n12410_19[2]),.dout(n15926),.clk(gclk));
	jand g15677(.dina(n15926),.dinb(w_asqrt14_31[2]),.dout(n15927),.clk(gclk));
	jxor g15678(.dina(n15927),.dinb(w_n15310_0[0]),.dout(n15928),.clk(gclk));
	jand g15679(.dina(w_n15928_0[1]),.dinb(n15925),.dout(n15929),.clk(gclk));
	jor g15680(.dina(n15929),.dinb(w_n15924_0[1]),.dout(n15930),.clk(gclk));
	jand g15681(.dina(w_n15930_0[2]),.dinb(w_asqrt22_18[1]),.dout(n15931),.clk(gclk));
	jor g15682(.dina(w_n15930_0[1]),.dinb(w_asqrt22_18[0]),.dout(n15932),.clk(gclk));
	jxor g15683(.dina(w_n15313_0[0]),.dinb(w_n11858_26[1]),.dout(n15933),.clk(gclk));
	jand g15684(.dina(n15933),.dinb(w_asqrt14_31[1]),.dout(n15934),.clk(gclk));
	jxor g15685(.dina(n15934),.dinb(w_n15318_0[0]),.dout(n15935),.clk(gclk));
	jnot g15686(.din(w_n15935_0[1]),.dout(n15936),.clk(gclk));
	jand g15687(.dina(w_n15936_0[1]),.dinb(n15932),.dout(n15937),.clk(gclk));
	jor g15688(.dina(n15937),.dinb(w_n15931_0[1]),.dout(n15938),.clk(gclk));
	jand g15689(.dina(w_n15938_0[2]),.dinb(w_asqrt23_12[1]),.dout(n15939),.clk(gclk));
	jor g15690(.dina(w_n15938_0[1]),.dinb(w_asqrt23_12[0]),.dout(n15940),.clk(gclk));
	jxor g15691(.dina(w_n15320_0[0]),.dinb(w_n11347_20[1]),.dout(n15941),.clk(gclk));
	jand g15692(.dina(n15941),.dinb(w_asqrt14_31[0]),.dout(n15942),.clk(gclk));
	jxor g15693(.dina(n15942),.dinb(w_n15325_0[0]),.dout(n15943),.clk(gclk));
	jand g15694(.dina(w_n15943_0[1]),.dinb(n15940),.dout(n15944),.clk(gclk));
	jor g15695(.dina(n15944),.dinb(w_n15939_0[1]),.dout(n15945),.clk(gclk));
	jand g15696(.dina(w_n15945_0[2]),.dinb(w_asqrt24_18[1]),.dout(n15946),.clk(gclk));
	jor g15697(.dina(w_n15945_0[1]),.dinb(w_asqrt24_18[0]),.dout(n15947),.clk(gclk));
	jxor g15698(.dina(w_n15328_0[0]),.dinb(w_n10824_27[0]),.dout(n15948),.clk(gclk));
	jand g15699(.dina(n15948),.dinb(w_asqrt14_30[2]),.dout(n15949),.clk(gclk));
	jxor g15700(.dina(n15949),.dinb(w_n15333_0[0]),.dout(n15950),.clk(gclk));
	jnot g15701(.din(w_n15950_0[1]),.dout(n15951),.clk(gclk));
	jand g15702(.dina(w_n15951_0[1]),.dinb(n15947),.dout(n15952),.clk(gclk));
	jor g15703(.dina(n15952),.dinb(w_n15946_0[1]),.dout(n15953),.clk(gclk));
	jand g15704(.dina(w_n15953_0[2]),.dinb(w_asqrt25_12[1]),.dout(n15954),.clk(gclk));
	jor g15705(.dina(w_n15953_0[1]),.dinb(w_asqrt25_12[0]),.dout(n15955),.clk(gclk));
	jxor g15706(.dina(w_n15335_0[0]),.dinb(w_n10328_21[1]),.dout(n15956),.clk(gclk));
	jand g15707(.dina(n15956),.dinb(w_asqrt14_30[1]),.dout(n15957),.clk(gclk));
	jxor g15708(.dina(n15957),.dinb(w_n15340_0[0]),.dout(n15958),.clk(gclk));
	jnot g15709(.din(w_n15958_0[1]),.dout(n15959),.clk(gclk));
	jand g15710(.dina(w_n15959_0[1]),.dinb(n15955),.dout(n15960),.clk(gclk));
	jor g15711(.dina(n15960),.dinb(w_n15954_0[1]),.dout(n15961),.clk(gclk));
	jand g15712(.dina(w_n15961_0[2]),.dinb(w_asqrt26_18[1]),.dout(n15962),.clk(gclk));
	jor g15713(.dina(w_n15961_0[1]),.dinb(w_asqrt26_18[0]),.dout(n15963),.clk(gclk));
	jxor g15714(.dina(w_n15342_0[0]),.dinb(w_n9832_27[2]),.dout(n15964),.clk(gclk));
	jand g15715(.dina(n15964),.dinb(w_asqrt14_30[0]),.dout(n15965),.clk(gclk));
	jxor g15716(.dina(n15965),.dinb(w_n15347_0[0]),.dout(n15966),.clk(gclk));
	jnot g15717(.din(w_n15966_0[1]),.dout(n15967),.clk(gclk));
	jand g15718(.dina(w_n15967_0[1]),.dinb(n15963),.dout(n15968),.clk(gclk));
	jor g15719(.dina(n15968),.dinb(w_n15962_0[1]),.dout(n15969),.clk(gclk));
	jand g15720(.dina(w_n15969_0[2]),.dinb(w_asqrt27_13[0]),.dout(n15970),.clk(gclk));
	jor g15721(.dina(w_n15969_0[1]),.dinb(w_asqrt27_12[2]),.dout(n15971),.clk(gclk));
	jxor g15722(.dina(w_n15349_0[0]),.dinb(w_n9369_22[1]),.dout(n15972),.clk(gclk));
	jand g15723(.dina(n15972),.dinb(w_asqrt14_29[2]),.dout(n15973),.clk(gclk));
	jxor g15724(.dina(n15973),.dinb(w_n15354_0[0]),.dout(n15974),.clk(gclk));
	jand g15725(.dina(w_n15974_0[1]),.dinb(n15971),.dout(n15975),.clk(gclk));
	jor g15726(.dina(n15975),.dinb(w_n15970_0[1]),.dout(n15976),.clk(gclk));
	jand g15727(.dina(w_n15976_0[2]),.dinb(w_asqrt28_18[2]),.dout(n15977),.clk(gclk));
	jor g15728(.dina(w_n15976_0[1]),.dinb(w_asqrt28_18[1]),.dout(n15978),.clk(gclk));
	jxor g15729(.dina(w_n15357_0[0]),.dinb(w_n8890_28[0]),.dout(n15979),.clk(gclk));
	jand g15730(.dina(n15979),.dinb(w_asqrt14_29[1]),.dout(n15980),.clk(gclk));
	jxor g15731(.dina(n15980),.dinb(w_n15362_0[0]),.dout(n15981),.clk(gclk));
	jnot g15732(.din(w_n15981_0[1]),.dout(n15982),.clk(gclk));
	jand g15733(.dina(w_n15982_0[1]),.dinb(n15978),.dout(n15983),.clk(gclk));
	jor g15734(.dina(n15983),.dinb(w_n15977_0[1]),.dout(n15984),.clk(gclk));
	jand g15735(.dina(w_n15984_0[2]),.dinb(w_asqrt29_13[1]),.dout(n15985),.clk(gclk));
	jor g15736(.dina(w_n15984_0[1]),.dinb(w_asqrt29_13[0]),.dout(n15986),.clk(gclk));
	jxor g15737(.dina(w_n15364_0[0]),.dinb(w_n8449_23[0]),.dout(n15987),.clk(gclk));
	jand g15738(.dina(n15987),.dinb(w_asqrt14_29[0]),.dout(n15988),.clk(gclk));
	jxor g15739(.dina(n15988),.dinb(w_n15369_0[0]),.dout(n15989),.clk(gclk));
	jand g15740(.dina(w_n15989_0[1]),.dinb(n15986),.dout(n15990),.clk(gclk));
	jor g15741(.dina(n15990),.dinb(w_n15985_0[1]),.dout(n15991),.clk(gclk));
	jand g15742(.dina(w_n15991_0[2]),.dinb(w_asqrt30_19[0]),.dout(n15992),.clk(gclk));
	jor g15743(.dina(w_n15991_0[1]),.dinb(w_asqrt30_18[2]),.dout(n15993),.clk(gclk));
	jxor g15744(.dina(w_n15372_0[0]),.dinb(w_n8003_28[2]),.dout(n15994),.clk(gclk));
	jand g15745(.dina(n15994),.dinb(w_asqrt14_28[2]),.dout(n15995),.clk(gclk));
	jxor g15746(.dina(n15995),.dinb(w_n15377_0[0]),.dout(n15996),.clk(gclk));
	jnot g15747(.din(w_n15996_0[1]),.dout(n15997),.clk(gclk));
	jand g15748(.dina(w_n15997_0[1]),.dinb(n15993),.dout(n15998),.clk(gclk));
	jor g15749(.dina(n15998),.dinb(w_n15992_0[1]),.dout(n15999),.clk(gclk));
	jand g15750(.dina(w_n15999_0[2]),.dinb(w_asqrt31_14[0]),.dout(n16000),.clk(gclk));
	jor g15751(.dina(w_n15999_0[1]),.dinb(w_asqrt31_13[2]),.dout(n16001),.clk(gclk));
	jxor g15752(.dina(w_n15379_0[0]),.dinb(w_n7581_24[0]),.dout(n16002),.clk(gclk));
	jand g15753(.dina(n16002),.dinb(w_asqrt14_28[1]),.dout(n16003),.clk(gclk));
	jxor g15754(.dina(n16003),.dinb(w_n15384_0[0]),.dout(n16004),.clk(gclk));
	jand g15755(.dina(w_n16004_0[1]),.dinb(n16001),.dout(n16005),.clk(gclk));
	jor g15756(.dina(n16005),.dinb(w_n16000_0[1]),.dout(n16006),.clk(gclk));
	jand g15757(.dina(w_n16006_0[2]),.dinb(w_asqrt32_19[0]),.dout(n16007),.clk(gclk));
	jor g15758(.dina(w_n16006_0[1]),.dinb(w_asqrt32_18[2]),.dout(n16008),.clk(gclk));
	jxor g15759(.dina(w_n15387_0[0]),.dinb(w_n7154_29[0]),.dout(n16009),.clk(gclk));
	jand g15760(.dina(n16009),.dinb(w_asqrt14_28[0]),.dout(n16010),.clk(gclk));
	jxor g15761(.dina(n16010),.dinb(w_n15392_0[0]),.dout(n16011),.clk(gclk));
	jnot g15762(.din(w_n16011_0[1]),.dout(n16012),.clk(gclk));
	jand g15763(.dina(w_n16012_0[1]),.dinb(n16008),.dout(n16013),.clk(gclk));
	jor g15764(.dina(n16013),.dinb(w_n16007_0[1]),.dout(n16014),.clk(gclk));
	jand g15765(.dina(w_n16014_0[2]),.dinb(w_asqrt33_14[2]),.dout(n16015),.clk(gclk));
	jor g15766(.dina(w_n16014_0[1]),.dinb(w_asqrt33_14[1]),.dout(n16016),.clk(gclk));
	jxor g15767(.dina(w_n15394_0[0]),.dinb(w_n6758_24[2]),.dout(n16017),.clk(gclk));
	jand g15768(.dina(n16017),.dinb(w_asqrt14_27[2]),.dout(n16018),.clk(gclk));
	jxor g15769(.dina(n16018),.dinb(w_n15399_0[0]),.dout(n16019),.clk(gclk));
	jand g15770(.dina(w_n16019_0[1]),.dinb(n16016),.dout(n16020),.clk(gclk));
	jor g15771(.dina(n16020),.dinb(w_n16015_0[1]),.dout(n16021),.clk(gclk));
	jand g15772(.dina(w_n16021_0[2]),.dinb(w_asqrt34_19[1]),.dout(n16022),.clk(gclk));
	jor g15773(.dina(w_n16021_0[1]),.dinb(w_asqrt34_19[0]),.dout(n16023),.clk(gclk));
	jxor g15774(.dina(w_n15402_0[0]),.dinb(w_n6357_29[1]),.dout(n16024),.clk(gclk));
	jand g15775(.dina(n16024),.dinb(w_asqrt14_27[1]),.dout(n16025),.clk(gclk));
	jxor g15776(.dina(n16025),.dinb(w_n15407_0[0]),.dout(n16026),.clk(gclk));
	jnot g15777(.din(w_n16026_0[1]),.dout(n16027),.clk(gclk));
	jand g15778(.dina(w_n16027_0[1]),.dinb(n16023),.dout(n16028),.clk(gclk));
	jor g15779(.dina(n16028),.dinb(w_n16022_0[1]),.dout(n16029),.clk(gclk));
	jand g15780(.dina(w_n16029_0[2]),.dinb(w_asqrt35_15[1]),.dout(n16030),.clk(gclk));
	jor g15781(.dina(w_n16029_0[1]),.dinb(w_asqrt35_15[0]),.dout(n16031),.clk(gclk));
	jxor g15782(.dina(w_n15409_0[0]),.dinb(w_n5989_25[1]),.dout(n16032),.clk(gclk));
	jand g15783(.dina(n16032),.dinb(w_asqrt14_27[0]),.dout(n16033),.clk(gclk));
	jxor g15784(.dina(n16033),.dinb(w_n15414_0[0]),.dout(n16034),.clk(gclk));
	jnot g15785(.din(w_n16034_0[1]),.dout(n16035),.clk(gclk));
	jand g15786(.dina(w_n16035_0[1]),.dinb(n16031),.dout(n16036),.clk(gclk));
	jor g15787(.dina(n16036),.dinb(w_n16030_0[1]),.dout(n16037),.clk(gclk));
	jand g15788(.dina(w_n16037_0[2]),.dinb(w_asqrt36_19[1]),.dout(n16038),.clk(gclk));
	jor g15789(.dina(w_n16037_0[1]),.dinb(w_asqrt36_19[0]),.dout(n16039),.clk(gclk));
	jxor g15790(.dina(w_n15416_0[0]),.dinb(w_n5606_29[2]),.dout(n16040),.clk(gclk));
	jand g15791(.dina(n16040),.dinb(w_asqrt14_26[2]),.dout(n16041),.clk(gclk));
	jxor g15792(.dina(n16041),.dinb(w_n15421_0[0]),.dout(n16042),.clk(gclk));
	jnot g15793(.din(w_n16042_0[1]),.dout(n16043),.clk(gclk));
	jand g15794(.dina(w_n16043_0[1]),.dinb(n16039),.dout(n16044),.clk(gclk));
	jor g15795(.dina(n16044),.dinb(w_n16038_0[1]),.dout(n16045),.clk(gclk));
	jand g15796(.dina(w_n16045_0[2]),.dinb(w_asqrt37_15[2]),.dout(n16046),.clk(gclk));
	jor g15797(.dina(w_n16045_0[1]),.dinb(w_asqrt37_15[1]),.dout(n16047),.clk(gclk));
	jxor g15798(.dina(w_n15423_0[0]),.dinb(w_n5259_26[1]),.dout(n16048),.clk(gclk));
	jand g15799(.dina(n16048),.dinb(w_asqrt14_26[1]),.dout(n16049),.clk(gclk));
	jxor g15800(.dina(n16049),.dinb(w_n15428_0[0]),.dout(n16050),.clk(gclk));
	jand g15801(.dina(w_n16050_0[1]),.dinb(n16047),.dout(n16051),.clk(gclk));
	jor g15802(.dina(n16051),.dinb(w_n16046_0[1]),.dout(n16052),.clk(gclk));
	jand g15803(.dina(w_n16052_0[2]),.dinb(w_asqrt38_19[2]),.dout(n16053),.clk(gclk));
	jor g15804(.dina(w_n16052_0[1]),.dinb(w_asqrt38_19[1]),.dout(n16054),.clk(gclk));
	jxor g15805(.dina(w_n15431_0[0]),.dinb(w_n4902_30[1]),.dout(n16055),.clk(gclk));
	jand g15806(.dina(n16055),.dinb(w_asqrt14_26[0]),.dout(n16056),.clk(gclk));
	jxor g15807(.dina(n16056),.dinb(w_n15436_0[0]),.dout(n16057),.clk(gclk));
	jnot g15808(.din(w_n16057_0[1]),.dout(n16058),.clk(gclk));
	jand g15809(.dina(w_n16058_0[1]),.dinb(n16054),.dout(n16059),.clk(gclk));
	jor g15810(.dina(n16059),.dinb(w_n16053_0[1]),.dout(n16060),.clk(gclk));
	jand g15811(.dina(w_n16060_0[2]),.dinb(w_asqrt39_16[1]),.dout(n16061),.clk(gclk));
	jor g15812(.dina(w_n16060_0[1]),.dinb(w_asqrt39_16[0]),.dout(n16062),.clk(gclk));
	jxor g15813(.dina(w_n15438_0[0]),.dinb(w_n4582_27[1]),.dout(n16063),.clk(gclk));
	jand g15814(.dina(n16063),.dinb(w_asqrt14_25[2]),.dout(n16064),.clk(gclk));
	jxor g15815(.dina(n16064),.dinb(w_n15443_0[0]),.dout(n16065),.clk(gclk));
	jand g15816(.dina(w_n16065_0[1]),.dinb(n16062),.dout(n16066),.clk(gclk));
	jor g15817(.dina(n16066),.dinb(w_n16061_0[1]),.dout(n16067),.clk(gclk));
	jand g15818(.dina(w_n16067_0[2]),.dinb(w_asqrt40_19[2]),.dout(n16068),.clk(gclk));
	jor g15819(.dina(w_n16067_0[1]),.dinb(w_asqrt40_19[1]),.dout(n16069),.clk(gclk));
	jxor g15820(.dina(w_n15446_0[0]),.dinb(w_n4249_31[0]),.dout(n16070),.clk(gclk));
	jand g15821(.dina(n16070),.dinb(w_asqrt14_25[1]),.dout(n16071),.clk(gclk));
	jxor g15822(.dina(n16071),.dinb(w_n15451_0[0]),.dout(n16072),.clk(gclk));
	jnot g15823(.din(w_n16072_0[1]),.dout(n16073),.clk(gclk));
	jand g15824(.dina(w_n16073_0[1]),.dinb(n16069),.dout(n16074),.clk(gclk));
	jor g15825(.dina(n16074),.dinb(w_n16068_0[1]),.dout(n16075),.clk(gclk));
	jand g15826(.dina(w_n16075_0[2]),.dinb(w_asqrt41_16[2]),.dout(n16076),.clk(gclk));
	jor g15827(.dina(w_n16075_0[1]),.dinb(w_asqrt41_16[1]),.dout(n16077),.clk(gclk));
	jxor g15828(.dina(w_n15453_0[0]),.dinb(w_n3955_28[0]),.dout(n16078),.clk(gclk));
	jand g15829(.dina(n16078),.dinb(w_asqrt14_25[0]),.dout(n16079),.clk(gclk));
	jxor g15830(.dina(n16079),.dinb(w_n15458_0[0]),.dout(n16080),.clk(gclk));
	jnot g15831(.din(w_n16080_0[1]),.dout(n16081),.clk(gclk));
	jand g15832(.dina(w_n16081_0[1]),.dinb(n16077),.dout(n16082),.clk(gclk));
	jor g15833(.dina(n16082),.dinb(w_n16076_0[1]),.dout(n16083),.clk(gclk));
	jand g15834(.dina(w_n16083_0[2]),.dinb(w_asqrt42_20[0]),.dout(n16084),.clk(gclk));
	jor g15835(.dina(w_n16083_0[1]),.dinb(w_asqrt42_19[2]),.dout(n16085),.clk(gclk));
	jxor g15836(.dina(w_n15460_0[0]),.dinb(w_n3642_31[1]),.dout(n16086),.clk(gclk));
	jand g15837(.dina(n16086),.dinb(w_asqrt14_24[2]),.dout(n16087),.clk(gclk));
	jxor g15838(.dina(n16087),.dinb(w_n15465_0[0]),.dout(n16088),.clk(gclk));
	jnot g15839(.din(w_n16088_0[1]),.dout(n16089),.clk(gclk));
	jand g15840(.dina(w_n16089_0[1]),.dinb(n16085),.dout(n16090),.clk(gclk));
	jor g15841(.dina(n16090),.dinb(w_n16084_0[1]),.dout(n16091),.clk(gclk));
	jand g15842(.dina(w_n16091_0[2]),.dinb(w_asqrt43_17[0]),.dout(n16092),.clk(gclk));
	jor g15843(.dina(w_n16091_0[1]),.dinb(w_asqrt43_16[2]),.dout(n16093),.clk(gclk));
	jxor g15844(.dina(w_n15467_0[0]),.dinb(w_n3368_28[2]),.dout(n16094),.clk(gclk));
	jand g15845(.dina(n16094),.dinb(w_asqrt14_24[1]),.dout(n16095),.clk(gclk));
	jxor g15846(.dina(n16095),.dinb(w_n15472_0[0]),.dout(n16096),.clk(gclk));
	jand g15847(.dina(w_n16096_0[1]),.dinb(n16093),.dout(n16097),.clk(gclk));
	jor g15848(.dina(n16097),.dinb(w_n16092_0[1]),.dout(n16098),.clk(gclk));
	jand g15849(.dina(w_n16098_0[2]),.dinb(w_asqrt44_20[0]),.dout(n16099),.clk(gclk));
	jor g15850(.dina(w_n16098_0[1]),.dinb(w_asqrt44_19[2]),.dout(n16100),.clk(gclk));
	jxor g15851(.dina(w_n15475_0[0]),.dinb(w_n3089_32[0]),.dout(n16101),.clk(gclk));
	jand g15852(.dina(n16101),.dinb(w_asqrt14_24[0]),.dout(n16102),.clk(gclk));
	jxor g15853(.dina(n16102),.dinb(w_n15480_0[0]),.dout(n16103),.clk(gclk));
	jnot g15854(.din(w_n16103_0[1]),.dout(n16104),.clk(gclk));
	jand g15855(.dina(w_n16104_0[1]),.dinb(n16100),.dout(n16105),.clk(gclk));
	jor g15856(.dina(n16105),.dinb(w_n16099_0[1]),.dout(n16106),.clk(gclk));
	jand g15857(.dina(w_n16106_0[2]),.dinb(w_asqrt45_17[2]),.dout(n16107),.clk(gclk));
	jor g15858(.dina(w_n16106_0[1]),.dinb(w_asqrt45_17[1]),.dout(n16108),.clk(gclk));
	jxor g15859(.dina(w_n15482_0[0]),.dinb(w_n2833_29[2]),.dout(n16109),.clk(gclk));
	jand g15860(.dina(n16109),.dinb(w_asqrt14_23[2]),.dout(n16110),.clk(gclk));
	jxor g15861(.dina(n16110),.dinb(w_n15487_0[0]),.dout(n16111),.clk(gclk));
	jand g15862(.dina(w_n16111_0[1]),.dinb(n16108),.dout(n16112),.clk(gclk));
	jor g15863(.dina(n16112),.dinb(w_n16107_0[1]),.dout(n16113),.clk(gclk));
	jand g15864(.dina(w_n16113_0[2]),.dinb(w_asqrt46_20[0]),.dout(n16114),.clk(gclk));
	jor g15865(.dina(w_n16113_0[1]),.dinb(w_asqrt46_19[2]),.dout(n16115),.clk(gclk));
	jxor g15866(.dina(w_n15490_0[0]),.dinb(w_n2572_32[1]),.dout(n16116),.clk(gclk));
	jand g15867(.dina(n16116),.dinb(w_asqrt14_23[1]),.dout(n16117),.clk(gclk));
	jxor g15868(.dina(n16117),.dinb(w_n15495_0[0]),.dout(n16118),.clk(gclk));
	jnot g15869(.din(w_n16118_0[1]),.dout(n16119),.clk(gclk));
	jand g15870(.dina(w_n16119_0[1]),.dinb(n16115),.dout(n16120),.clk(gclk));
	jor g15871(.dina(n16120),.dinb(w_n16114_0[1]),.dout(n16121),.clk(gclk));
	jand g15872(.dina(w_n16121_0[2]),.dinb(w_asqrt47_18[1]),.dout(n16122),.clk(gclk));
	jor g15873(.dina(w_n16121_0[1]),.dinb(w_asqrt47_18[0]),.dout(n16123),.clk(gclk));
	jxor g15874(.dina(w_n15497_0[0]),.dinb(w_n2345_30[1]),.dout(n16124),.clk(gclk));
	jand g15875(.dina(n16124),.dinb(w_asqrt14_23[0]),.dout(n16125),.clk(gclk));
	jxor g15876(.dina(n16125),.dinb(w_n15502_0[0]),.dout(n16126),.clk(gclk));
	jnot g15877(.din(w_n16126_0[1]),.dout(n16127),.clk(gclk));
	jand g15878(.dina(w_n16127_0[1]),.dinb(n16123),.dout(n16128),.clk(gclk));
	jor g15879(.dina(n16128),.dinb(w_n16122_0[1]),.dout(n16129),.clk(gclk));
	jand g15880(.dina(w_n16129_0[2]),.dinb(w_asqrt48_20[1]),.dout(n16130),.clk(gclk));
	jor g15881(.dina(w_n16129_0[1]),.dinb(w_asqrt48_20[0]),.dout(n16131),.clk(gclk));
	jxor g15882(.dina(w_n15504_0[0]),.dinb(w_n2108_33[0]),.dout(n16132),.clk(gclk));
	jand g15883(.dina(n16132),.dinb(w_asqrt14_22[2]),.dout(n16133),.clk(gclk));
	jxor g15884(.dina(n16133),.dinb(w_n15509_0[0]),.dout(n16134),.clk(gclk));
	jand g15885(.dina(w_n16134_0[1]),.dinb(n16131),.dout(n16135),.clk(gclk));
	jor g15886(.dina(n16135),.dinb(w_n16130_0[1]),.dout(n16136),.clk(gclk));
	jand g15887(.dina(w_n16136_0[2]),.dinb(w_asqrt49_18[2]),.dout(n16137),.clk(gclk));
	jxor g15888(.dina(w_n15512_0[0]),.dinb(w_n1912_31[1]),.dout(n16138),.clk(gclk));
	jand g15889(.dina(n16138),.dinb(w_asqrt14_22[1]),.dout(n16139),.clk(gclk));
	jxor g15890(.dina(n16139),.dinb(w_n15516_0[0]),.dout(n16140),.clk(gclk));
	jor g15891(.dina(w_n16136_0[1]),.dinb(w_asqrt49_18[1]),.dout(n16141),.clk(gclk));
	jand g15892(.dina(n16141),.dinb(w_n16140_0[1]),.dout(n16142),.clk(gclk));
	jor g15893(.dina(n16142),.dinb(w_n16137_0[1]),.dout(n16143),.clk(gclk));
	jand g15894(.dina(w_n16143_0[2]),.dinb(w_asqrt50_20[2]),.dout(n16144),.clk(gclk));
	jor g15895(.dina(w_n16143_0[1]),.dinb(w_asqrt50_20[1]),.dout(n16145),.clk(gclk));
	jxor g15896(.dina(w_n15520_0[0]),.dinb(w_n1699_33[2]),.dout(n16146),.clk(gclk));
	jand g15897(.dina(n16146),.dinb(w_asqrt14_22[0]),.dout(n16147),.clk(gclk));
	jxor g15898(.dina(n16147),.dinb(w_n15525_0[0]),.dout(n16148),.clk(gclk));
	jnot g15899(.din(w_n16148_0[1]),.dout(n16149),.clk(gclk));
	jand g15900(.dina(w_n16149_0[1]),.dinb(n16145),.dout(n16150),.clk(gclk));
	jor g15901(.dina(n16150),.dinb(w_n16144_0[1]),.dout(n16151),.clk(gclk));
	jand g15902(.dina(w_n16151_0[2]),.dinb(w_asqrt51_19[0]),.dout(n16152),.clk(gclk));
	jor g15903(.dina(w_n16151_0[1]),.dinb(w_asqrt51_18[2]),.dout(n16153),.clk(gclk));
	jxor g15904(.dina(w_n15527_0[0]),.dinb(w_n1516_32[0]),.dout(n16154),.clk(gclk));
	jand g15905(.dina(n16154),.dinb(w_asqrt14_21[2]),.dout(n16155),.clk(gclk));
	jxor g15906(.dina(n16155),.dinb(w_n15532_0[0]),.dout(n16156),.clk(gclk));
	jand g15907(.dina(w_n16156_0[1]),.dinb(n16153),.dout(n16157),.clk(gclk));
	jor g15908(.dina(n16157),.dinb(w_n16152_0[1]),.dout(n16158),.clk(gclk));
	jand g15909(.dina(w_n16158_0[2]),.dinb(w_asqrt52_20[2]),.dout(n16159),.clk(gclk));
	jor g15910(.dina(w_n16158_0[1]),.dinb(w_asqrt52_20[1]),.dout(n16160),.clk(gclk));
	jxor g15911(.dina(w_n15535_0[0]),.dinb(w_n1332_33[2]),.dout(n16161),.clk(gclk));
	jand g15912(.dina(n16161),.dinb(w_asqrt14_21[1]),.dout(n16162),.clk(gclk));
	jxor g15913(.dina(n16162),.dinb(w_n15540_0[0]),.dout(n16163),.clk(gclk));
	jnot g15914(.din(w_n16163_0[1]),.dout(n16164),.clk(gclk));
	jand g15915(.dina(w_n16164_0[1]),.dinb(n16160),.dout(n16165),.clk(gclk));
	jor g15916(.dina(n16165),.dinb(w_n16159_0[1]),.dout(n16166),.clk(gclk));
	jand g15917(.dina(w_n16166_0[2]),.dinb(w_asqrt53_19[2]),.dout(n16167),.clk(gclk));
	jor g15918(.dina(w_n16166_0[1]),.dinb(w_asqrt53_19[1]),.dout(n16168),.clk(gclk));
	jxor g15919(.dina(w_n15542_0[0]),.dinb(w_n1173_32[2]),.dout(n16169),.clk(gclk));
	jand g15920(.dina(n16169),.dinb(w_asqrt14_21[0]),.dout(n16170),.clk(gclk));
	jxor g15921(.dina(n16170),.dinb(w_n15547_0[0]),.dout(n16171),.clk(gclk));
	jand g15922(.dina(w_n16171_0[1]),.dinb(n16168),.dout(n16172),.clk(gclk));
	jor g15923(.dina(n16172),.dinb(w_n16167_0[1]),.dout(n16173),.clk(gclk));
	jand g15924(.dina(w_n16173_0[2]),.dinb(w_asqrt54_20[2]),.dout(n16174),.clk(gclk));
	jor g15925(.dina(w_n16173_0[1]),.dinb(w_asqrt54_20[1]),.dout(n16175),.clk(gclk));
	jxor g15926(.dina(w_n15550_0[0]),.dinb(w_n1008_34[2]),.dout(n16176),.clk(gclk));
	jand g15927(.dina(n16176),.dinb(w_asqrt14_20[2]),.dout(n16177),.clk(gclk));
	jxor g15928(.dina(n16177),.dinb(w_n15555_0[0]),.dout(n16178),.clk(gclk));
	jnot g15929(.din(w_n16178_0[1]),.dout(n16179),.clk(gclk));
	jand g15930(.dina(w_n16179_0[1]),.dinb(n16175),.dout(n16180),.clk(gclk));
	jor g15931(.dina(n16180),.dinb(w_n16174_0[1]),.dout(n16181),.clk(gclk));
	jand g15932(.dina(w_n16181_0[2]),.dinb(w_asqrt55_20[0]),.dout(n16182),.clk(gclk));
	jor g15933(.dina(w_n16181_0[1]),.dinb(w_asqrt55_19[2]),.dout(n16183),.clk(gclk));
	jxor g15934(.dina(w_n15557_0[0]),.dinb(w_n884_33[2]),.dout(n16184),.clk(gclk));
	jand g15935(.dina(n16184),.dinb(w_asqrt14_20[1]),.dout(n16185),.clk(gclk));
	jxor g15936(.dina(n16185),.dinb(w_n15562_0[0]),.dout(n16186),.clk(gclk));
	jnot g15937(.din(w_n16186_0[1]),.dout(n16187),.clk(gclk));
	jand g15938(.dina(w_n16187_0[1]),.dinb(n16183),.dout(n16188),.clk(gclk));
	jor g15939(.dina(n16188),.dinb(w_n16182_0[1]),.dout(n16189),.clk(gclk));
	jand g15940(.dina(w_n16189_0[2]),.dinb(w_asqrt56_21[0]),.dout(n16190),.clk(gclk));
	jor g15941(.dina(w_n16189_0[1]),.dinb(w_asqrt56_20[2]),.dout(n16191),.clk(gclk));
	jxor g15942(.dina(w_n15564_0[0]),.dinb(w_n743_34[2]),.dout(n16192),.clk(gclk));
	jand g15943(.dina(n16192),.dinb(w_asqrt14_20[0]),.dout(n16193),.clk(gclk));
	jxor g15944(.dina(n16193),.dinb(w_n15569_0[0]),.dout(n16194),.clk(gclk));
	jnot g15945(.din(w_n16194_0[1]),.dout(n16195),.clk(gclk));
	jand g15946(.dina(w_n16195_0[1]),.dinb(n16191),.dout(n16196),.clk(gclk));
	jor g15947(.dina(n16196),.dinb(w_n16190_0[1]),.dout(n16197),.clk(gclk));
	jand g15948(.dina(w_n16197_0[2]),.dinb(w_asqrt57_20[2]),.dout(n16198),.clk(gclk));
	jor g15949(.dina(w_n16197_0[1]),.dinb(w_asqrt57_20[1]),.dout(n16199),.clk(gclk));
	jxor g15950(.dina(w_n15571_0[0]),.dinb(w_n635_34[2]),.dout(n16200),.clk(gclk));
	jand g15951(.dina(n16200),.dinb(w_asqrt14_19[2]),.dout(n16201),.clk(gclk));
	jxor g15952(.dina(n16201),.dinb(w_n15576_0[0]),.dout(n16202),.clk(gclk));
	jand g15953(.dina(w_n16202_0[1]),.dinb(n16199),.dout(n16203),.clk(gclk));
	jor g15954(.dina(n16203),.dinb(w_n16198_0[1]),.dout(n16204),.clk(gclk));
	jand g15955(.dina(w_n16204_0[2]),.dinb(w_asqrt58_21[1]),.dout(n16205),.clk(gclk));
	jor g15956(.dina(w_n16204_0[1]),.dinb(w_asqrt58_21[0]),.dout(n16206),.clk(gclk));
	jxor g15957(.dina(w_n15579_0[0]),.dinb(w_n515_35[2]),.dout(n16207),.clk(gclk));
	jand g15958(.dina(n16207),.dinb(w_asqrt14_19[1]),.dout(n16208),.clk(gclk));
	jxor g15959(.dina(n16208),.dinb(w_n15584_0[0]),.dout(n16209),.clk(gclk));
	jnot g15960(.din(w_n16209_0[1]),.dout(n16210),.clk(gclk));
	jand g15961(.dina(w_n16210_0[1]),.dinb(n16206),.dout(n16211),.clk(gclk));
	jor g15962(.dina(n16211),.dinb(w_n16205_0[1]),.dout(n16212),.clk(gclk));
	jand g15963(.dina(w_n16212_0[2]),.dinb(w_asqrt59_21[0]),.dout(n16213),.clk(gclk));
	jor g15964(.dina(w_n16212_0[1]),.dinb(w_asqrt59_20[2]),.dout(n16214),.clk(gclk));
	jxor g15965(.dina(w_n15586_0[0]),.dinb(w_n443_35[2]),.dout(n16215),.clk(gclk));
	jand g15966(.dina(n16215),.dinb(w_asqrt14_19[0]),.dout(n16216),.clk(gclk));
	jxor g15967(.dina(n16216),.dinb(w_n15591_0[0]),.dout(n16217),.clk(gclk));
	jand g15968(.dina(w_n16217_0[1]),.dinb(n16214),.dout(n16218),.clk(gclk));
	jor g15969(.dina(n16218),.dinb(w_n16213_0[1]),.dout(n16219),.clk(gclk));
	jand g15970(.dina(w_n16219_0[2]),.dinb(w_asqrt60_21[1]),.dout(n16220),.clk(gclk));
	jor g15971(.dina(w_n16219_0[1]),.dinb(w_asqrt60_21[0]),.dout(n16221),.clk(gclk));
	jxor g15972(.dina(w_n15594_0[0]),.dinb(w_n352_36[0]),.dout(n16222),.clk(gclk));
	jand g15973(.dina(n16222),.dinb(w_asqrt14_18[2]),.dout(n16223),.clk(gclk));
	jxor g15974(.dina(n16223),.dinb(w_n15599_0[0]),.dout(n16224),.clk(gclk));
	jnot g15975(.din(w_n16224_0[1]),.dout(n16225),.clk(gclk));
	jand g15976(.dina(w_n16225_0[1]),.dinb(n16221),.dout(n16226),.clk(gclk));
	jor g15977(.dina(n16226),.dinb(w_n16220_0[1]),.dout(n16227),.clk(gclk));
	jand g15978(.dina(w_n16227_0[2]),.dinb(w_asqrt61_21[1]),.dout(n16228),.clk(gclk));
	jor g15979(.dina(w_n16227_0[1]),.dinb(w_asqrt61_21[0]),.dout(n16229),.clk(gclk));
	jxor g15980(.dina(w_n15601_0[0]),.dinb(w_n294_36[1]),.dout(n16230),.clk(gclk));
	jand g15981(.dina(n16230),.dinb(w_asqrt14_18[1]),.dout(n16231),.clk(gclk));
	jxor g15982(.dina(n16231),.dinb(w_n15606_0[0]),.dout(n16232),.clk(gclk));
	jand g15983(.dina(w_n16232_0[1]),.dinb(n16229),.dout(n16233),.clk(gclk));
	jor g15984(.dina(n16233),.dinb(w_n16228_0[1]),.dout(n16234),.clk(gclk));
	jand g15985(.dina(w_n16234_0[2]),.dinb(w_asqrt62_21[1]),.dout(n16235),.clk(gclk));
	jnot g15986(.din(w_n16235_0[1]),.dout(n16236),.clk(gclk));
	jnot g15987(.din(w_n16228_0[0]),.dout(n16237),.clk(gclk));
	jnot g15988(.din(w_n16220_0[0]),.dout(n16238),.clk(gclk));
	jnot g15989(.din(w_n16213_0[0]),.dout(n16239),.clk(gclk));
	jnot g15990(.din(w_n16205_0[0]),.dout(n16240),.clk(gclk));
	jnot g15991(.din(w_n16198_0[0]),.dout(n16241),.clk(gclk));
	jnot g15992(.din(w_n16190_0[0]),.dout(n16242),.clk(gclk));
	jnot g15993(.din(w_n16182_0[0]),.dout(n16243),.clk(gclk));
	jnot g15994(.din(w_n16174_0[0]),.dout(n16244),.clk(gclk));
	jnot g15995(.din(w_n16167_0[0]),.dout(n16245),.clk(gclk));
	jnot g15996(.din(w_n16159_0[0]),.dout(n16246),.clk(gclk));
	jnot g15997(.din(w_n16152_0[0]),.dout(n16247),.clk(gclk));
	jnot g15998(.din(w_n16144_0[0]),.dout(n16248),.clk(gclk));
	jnot g15999(.din(w_n16137_0[0]),.dout(n16249),.clk(gclk));
	jnot g16000(.din(w_n16140_0[0]),.dout(n16250),.clk(gclk));
	jnot g16001(.din(w_n16130_0[0]),.dout(n16251),.clk(gclk));
	jnot g16002(.din(w_n16122_0[0]),.dout(n16252),.clk(gclk));
	jnot g16003(.din(w_n16114_0[0]),.dout(n16253),.clk(gclk));
	jnot g16004(.din(w_n16107_0[0]),.dout(n16254),.clk(gclk));
	jnot g16005(.din(w_n16099_0[0]),.dout(n16255),.clk(gclk));
	jnot g16006(.din(w_n16092_0[0]),.dout(n16256),.clk(gclk));
	jnot g16007(.din(w_n16084_0[0]),.dout(n16257),.clk(gclk));
	jnot g16008(.din(w_n16076_0[0]),.dout(n16258),.clk(gclk));
	jnot g16009(.din(w_n16068_0[0]),.dout(n16259),.clk(gclk));
	jnot g16010(.din(w_n16061_0[0]),.dout(n16260),.clk(gclk));
	jnot g16011(.din(w_n16053_0[0]),.dout(n16261),.clk(gclk));
	jnot g16012(.din(w_n16046_0[0]),.dout(n16262),.clk(gclk));
	jnot g16013(.din(w_n16038_0[0]),.dout(n16263),.clk(gclk));
	jnot g16014(.din(w_n16030_0[0]),.dout(n16264),.clk(gclk));
	jnot g16015(.din(w_n16022_0[0]),.dout(n16265),.clk(gclk));
	jnot g16016(.din(w_n16015_0[0]),.dout(n16266),.clk(gclk));
	jnot g16017(.din(w_n16007_0[0]),.dout(n16267),.clk(gclk));
	jnot g16018(.din(w_n16000_0[0]),.dout(n16268),.clk(gclk));
	jnot g16019(.din(w_n15992_0[0]),.dout(n16269),.clk(gclk));
	jnot g16020(.din(w_n15985_0[0]),.dout(n16270),.clk(gclk));
	jnot g16021(.din(w_n15977_0[0]),.dout(n16271),.clk(gclk));
	jnot g16022(.din(w_n15970_0[0]),.dout(n16272),.clk(gclk));
	jnot g16023(.din(w_n15962_0[0]),.dout(n16273),.clk(gclk));
	jnot g16024(.din(w_n15954_0[0]),.dout(n16274),.clk(gclk));
	jnot g16025(.din(w_n15946_0[0]),.dout(n16275),.clk(gclk));
	jnot g16026(.din(w_n15939_0[0]),.dout(n16276),.clk(gclk));
	jnot g16027(.din(w_n15931_0[0]),.dout(n16277),.clk(gclk));
	jnot g16028(.din(w_n15924_0[0]),.dout(n16278),.clk(gclk));
	jnot g16029(.din(w_n15916_0[0]),.dout(n16279),.clk(gclk));
	jnot g16030(.din(w_n15909_0[0]),.dout(n16280),.clk(gclk));
	jnot g16031(.din(w_n15902_0[0]),.dout(n16281),.clk(gclk));
	jnot g16032(.din(w_n15895_0[0]),.dout(n16282),.clk(gclk));
	jnot g16033(.din(w_n15883_0[0]),.dout(n16283),.clk(gclk));
	jnot g16034(.din(w_n15647_0[0]),.dout(n16284),.clk(gclk));
	jor g16035(.dina(w_n15878_18[0]),.dinb(w_n15265_0[2]),.dout(n16285),.clk(gclk));
	jnot g16036(.din(w_n15645_0[0]),.dout(n16286),.clk(gclk));
	jand g16037(.dina(n16286),.dinb(n16285),.dout(n16287),.clk(gclk));
	jand g16038(.dina(n16287),.dinb(w_n15260_24[2]),.dout(n16288),.clk(gclk));
	jor g16039(.dina(w_n15878_17[2]),.dinb(w_a28_0[0]),.dout(n16289),.clk(gclk));
	jand g16040(.dina(n16289),.dinb(w_a29_0[0]),.dout(n16290),.clk(gclk));
	jor g16041(.dina(w_n15885_0[0]),.dinb(n16290),.dout(n16291),.clk(gclk));
	jor g16042(.dina(w_n16291_0[1]),.dinb(n16288),.dout(n16292),.clk(gclk));
	jand g16043(.dina(n16292),.dinb(n16284),.dout(n16293),.clk(gclk));
	jand g16044(.dina(n16293),.dinb(w_n14674_17[2]),.dout(n16294),.clk(gclk));
	jor g16045(.dina(w_n15891_0[0]),.dinb(n16294),.dout(n16295),.clk(gclk));
	jand g16046(.dina(n16295),.dinb(n16283),.dout(n16296),.clk(gclk));
	jand g16047(.dina(n16296),.dinb(w_n14078_25[0]),.dout(n16297),.clk(gclk));
	jnot g16048(.din(w_n15899_0[1]),.dout(n16298),.clk(gclk));
	jor g16049(.dina(n16298),.dinb(n16297),.dout(n16299),.clk(gclk));
	jand g16050(.dina(n16299),.dinb(n16282),.dout(n16300),.clk(gclk));
	jand g16051(.dina(n16300),.dinb(w_n13515_18[2]),.dout(n16301),.clk(gclk));
	jnot g16052(.din(w_n15906_0[0]),.dout(n16302),.clk(gclk));
	jor g16053(.dina(w_n16302_0[1]),.dinb(n16301),.dout(n16303),.clk(gclk));
	jand g16054(.dina(n16303),.dinb(n16281),.dout(n16304),.clk(gclk));
	jand g16055(.dina(n16304),.dinb(w_n12947_25[2]),.dout(n16305),.clk(gclk));
	jnot g16056(.din(w_n15913_0[0]),.dout(n16306),.clk(gclk));
	jor g16057(.dina(w_n16306_0[1]),.dinb(n16305),.dout(n16307),.clk(gclk));
	jand g16058(.dina(n16307),.dinb(n16280),.dout(n16308),.clk(gclk));
	jand g16059(.dina(n16308),.dinb(w_n12410_19[1]),.dout(n16309),.clk(gclk));
	jor g16060(.dina(w_n15920_0[0]),.dinb(n16309),.dout(n16310),.clk(gclk));
	jand g16061(.dina(n16310),.dinb(n16279),.dout(n16311),.clk(gclk));
	jand g16062(.dina(n16311),.dinb(w_n11858_26[0]),.dout(n16312),.clk(gclk));
	jnot g16063(.din(w_n15928_0[0]),.dout(n16313),.clk(gclk));
	jor g16064(.dina(w_n16313_0[1]),.dinb(n16312),.dout(n16314),.clk(gclk));
	jand g16065(.dina(n16314),.dinb(n16278),.dout(n16315),.clk(gclk));
	jand g16066(.dina(n16315),.dinb(w_n11347_20[0]),.dout(n16316),.clk(gclk));
	jor g16067(.dina(w_n15935_0[0]),.dinb(n16316),.dout(n16317),.clk(gclk));
	jand g16068(.dina(n16317),.dinb(n16277),.dout(n16318),.clk(gclk));
	jand g16069(.dina(n16318),.dinb(w_n10824_26[2]),.dout(n16319),.clk(gclk));
	jnot g16070(.din(w_n15943_0[0]),.dout(n16320),.clk(gclk));
	jor g16071(.dina(w_n16320_0[1]),.dinb(n16319),.dout(n16321),.clk(gclk));
	jand g16072(.dina(n16321),.dinb(n16276),.dout(n16322),.clk(gclk));
	jand g16073(.dina(n16322),.dinb(w_n10328_21[0]),.dout(n16323),.clk(gclk));
	jor g16074(.dina(w_n15950_0[0]),.dinb(n16323),.dout(n16324),.clk(gclk));
	jand g16075(.dina(n16324),.dinb(n16275),.dout(n16325),.clk(gclk));
	jand g16076(.dina(n16325),.dinb(w_n9832_27[1]),.dout(n16326),.clk(gclk));
	jor g16077(.dina(w_n15958_0[0]),.dinb(n16326),.dout(n16327),.clk(gclk));
	jand g16078(.dina(n16327),.dinb(n16274),.dout(n16328),.clk(gclk));
	jand g16079(.dina(n16328),.dinb(w_n9369_22[0]),.dout(n16329),.clk(gclk));
	jor g16080(.dina(w_n15966_0[0]),.dinb(n16329),.dout(n16330),.clk(gclk));
	jand g16081(.dina(n16330),.dinb(n16273),.dout(n16331),.clk(gclk));
	jand g16082(.dina(n16331),.dinb(w_n8890_27[2]),.dout(n16332),.clk(gclk));
	jnot g16083(.din(w_n15974_0[0]),.dout(n16333),.clk(gclk));
	jor g16084(.dina(w_n16333_0[1]),.dinb(n16332),.dout(n16334),.clk(gclk));
	jand g16085(.dina(n16334),.dinb(n16272),.dout(n16335),.clk(gclk));
	jand g16086(.dina(n16335),.dinb(w_n8449_22[2]),.dout(n16336),.clk(gclk));
	jor g16087(.dina(w_n15981_0[0]),.dinb(n16336),.dout(n16337),.clk(gclk));
	jand g16088(.dina(n16337),.dinb(n16271),.dout(n16338),.clk(gclk));
	jand g16089(.dina(n16338),.dinb(w_n8003_28[1]),.dout(n16339),.clk(gclk));
	jnot g16090(.din(w_n15989_0[0]),.dout(n16340),.clk(gclk));
	jor g16091(.dina(w_n16340_0[1]),.dinb(n16339),.dout(n16341),.clk(gclk));
	jand g16092(.dina(n16341),.dinb(n16270),.dout(n16342),.clk(gclk));
	jand g16093(.dina(n16342),.dinb(w_n7581_23[2]),.dout(n16343),.clk(gclk));
	jor g16094(.dina(w_n15996_0[0]),.dinb(n16343),.dout(n16344),.clk(gclk));
	jand g16095(.dina(n16344),.dinb(n16269),.dout(n16345),.clk(gclk));
	jand g16096(.dina(n16345),.dinb(w_n7154_28[2]),.dout(n16346),.clk(gclk));
	jnot g16097(.din(w_n16004_0[0]),.dout(n16347),.clk(gclk));
	jor g16098(.dina(w_n16347_0[1]),.dinb(n16346),.dout(n16348),.clk(gclk));
	jand g16099(.dina(n16348),.dinb(n16268),.dout(n16349),.clk(gclk));
	jand g16100(.dina(n16349),.dinb(w_n6758_24[1]),.dout(n16350),.clk(gclk));
	jor g16101(.dina(w_n16011_0[0]),.dinb(n16350),.dout(n16351),.clk(gclk));
	jand g16102(.dina(n16351),.dinb(n16267),.dout(n16352),.clk(gclk));
	jand g16103(.dina(n16352),.dinb(w_n6357_29[0]),.dout(n16353),.clk(gclk));
	jnot g16104(.din(w_n16019_0[0]),.dout(n16354),.clk(gclk));
	jor g16105(.dina(w_n16354_0[1]),.dinb(n16353),.dout(n16355),.clk(gclk));
	jand g16106(.dina(n16355),.dinb(n16266),.dout(n16356),.clk(gclk));
	jand g16107(.dina(n16356),.dinb(w_n5989_25[0]),.dout(n16357),.clk(gclk));
	jor g16108(.dina(w_n16026_0[0]),.dinb(n16357),.dout(n16358),.clk(gclk));
	jand g16109(.dina(n16358),.dinb(n16265),.dout(n16359),.clk(gclk));
	jand g16110(.dina(n16359),.dinb(w_n5606_29[1]),.dout(n16360),.clk(gclk));
	jor g16111(.dina(w_n16034_0[0]),.dinb(n16360),.dout(n16361),.clk(gclk));
	jand g16112(.dina(n16361),.dinb(n16264),.dout(n16362),.clk(gclk));
	jand g16113(.dina(n16362),.dinb(w_n5259_26[0]),.dout(n16363),.clk(gclk));
	jor g16114(.dina(w_n16042_0[0]),.dinb(n16363),.dout(n16364),.clk(gclk));
	jand g16115(.dina(n16364),.dinb(n16263),.dout(n16365),.clk(gclk));
	jand g16116(.dina(n16365),.dinb(w_n4902_30[0]),.dout(n16366),.clk(gclk));
	jnot g16117(.din(w_n16050_0[0]),.dout(n16367),.clk(gclk));
	jor g16118(.dina(w_n16367_0[1]),.dinb(n16366),.dout(n16368),.clk(gclk));
	jand g16119(.dina(n16368),.dinb(n16262),.dout(n16369),.clk(gclk));
	jand g16120(.dina(n16369),.dinb(w_n4582_27[0]),.dout(n16370),.clk(gclk));
	jor g16121(.dina(w_n16057_0[0]),.dinb(n16370),.dout(n16371),.clk(gclk));
	jand g16122(.dina(n16371),.dinb(n16261),.dout(n16372),.clk(gclk));
	jand g16123(.dina(n16372),.dinb(w_n4249_30[2]),.dout(n16373),.clk(gclk));
	jnot g16124(.din(w_n16065_0[0]),.dout(n16374),.clk(gclk));
	jor g16125(.dina(w_n16374_0[1]),.dinb(n16373),.dout(n16375),.clk(gclk));
	jand g16126(.dina(n16375),.dinb(n16260),.dout(n16376),.clk(gclk));
	jand g16127(.dina(n16376),.dinb(w_n3955_27[2]),.dout(n16377),.clk(gclk));
	jor g16128(.dina(w_n16072_0[0]),.dinb(n16377),.dout(n16378),.clk(gclk));
	jand g16129(.dina(n16378),.dinb(n16259),.dout(n16379),.clk(gclk));
	jand g16130(.dina(n16379),.dinb(w_n3642_31[0]),.dout(n16380),.clk(gclk));
	jor g16131(.dina(w_n16080_0[0]),.dinb(n16380),.dout(n16381),.clk(gclk));
	jand g16132(.dina(n16381),.dinb(n16258),.dout(n16382),.clk(gclk));
	jand g16133(.dina(n16382),.dinb(w_n3368_28[1]),.dout(n16383),.clk(gclk));
	jor g16134(.dina(w_n16088_0[0]),.dinb(n16383),.dout(n16384),.clk(gclk));
	jand g16135(.dina(n16384),.dinb(n16257),.dout(n16385),.clk(gclk));
	jand g16136(.dina(n16385),.dinb(w_n3089_31[2]),.dout(n16386),.clk(gclk));
	jnot g16137(.din(w_n16096_0[0]),.dout(n16387),.clk(gclk));
	jor g16138(.dina(w_n16387_0[1]),.dinb(n16386),.dout(n16388),.clk(gclk));
	jand g16139(.dina(n16388),.dinb(n16256),.dout(n16389),.clk(gclk));
	jand g16140(.dina(n16389),.dinb(w_n2833_29[1]),.dout(n16390),.clk(gclk));
	jor g16141(.dina(w_n16103_0[0]),.dinb(n16390),.dout(n16391),.clk(gclk));
	jand g16142(.dina(n16391),.dinb(n16255),.dout(n16392),.clk(gclk));
	jand g16143(.dina(n16392),.dinb(w_n2572_32[0]),.dout(n16393),.clk(gclk));
	jnot g16144(.din(w_n16111_0[0]),.dout(n16394),.clk(gclk));
	jor g16145(.dina(w_n16394_0[1]),.dinb(n16393),.dout(n16395),.clk(gclk));
	jand g16146(.dina(n16395),.dinb(n16254),.dout(n16396),.clk(gclk));
	jand g16147(.dina(n16396),.dinb(w_n2345_30[0]),.dout(n16397),.clk(gclk));
	jor g16148(.dina(w_n16118_0[0]),.dinb(n16397),.dout(n16398),.clk(gclk));
	jand g16149(.dina(n16398),.dinb(n16253),.dout(n16399),.clk(gclk));
	jand g16150(.dina(n16399),.dinb(w_n2108_32[2]),.dout(n16400),.clk(gclk));
	jor g16151(.dina(w_n16126_0[0]),.dinb(n16400),.dout(n16401),.clk(gclk));
	jand g16152(.dina(n16401),.dinb(n16252),.dout(n16402),.clk(gclk));
	jand g16153(.dina(n16402),.dinb(w_n1912_31[0]),.dout(n16403),.clk(gclk));
	jnot g16154(.din(w_n16134_0[0]),.dout(n16404),.clk(gclk));
	jor g16155(.dina(w_n16404_0[1]),.dinb(n16403),.dout(n16405),.clk(gclk));
	jand g16156(.dina(n16405),.dinb(n16251),.dout(n16406),.clk(gclk));
	jand g16157(.dina(n16406),.dinb(w_n1699_33[1]),.dout(n16407),.clk(gclk));
	jor g16158(.dina(n16407),.dinb(w_n16250_0[1]),.dout(n16408),.clk(gclk));
	jand g16159(.dina(n16408),.dinb(n16249),.dout(n16409),.clk(gclk));
	jand g16160(.dina(n16409),.dinb(w_n1516_31[2]),.dout(n16410),.clk(gclk));
	jor g16161(.dina(w_n16148_0[0]),.dinb(n16410),.dout(n16411),.clk(gclk));
	jand g16162(.dina(n16411),.dinb(n16248),.dout(n16412),.clk(gclk));
	jand g16163(.dina(n16412),.dinb(w_n1332_33[1]),.dout(n16413),.clk(gclk));
	jnot g16164(.din(w_n16156_0[0]),.dout(n16414),.clk(gclk));
	jor g16165(.dina(w_n16414_0[1]),.dinb(n16413),.dout(n16415),.clk(gclk));
	jand g16166(.dina(n16415),.dinb(n16247),.dout(n16416),.clk(gclk));
	jand g16167(.dina(n16416),.dinb(w_n1173_32[1]),.dout(n16417),.clk(gclk));
	jor g16168(.dina(w_n16163_0[0]),.dinb(n16417),.dout(n16418),.clk(gclk));
	jand g16169(.dina(n16418),.dinb(n16246),.dout(n16419),.clk(gclk));
	jand g16170(.dina(n16419),.dinb(w_n1008_34[1]),.dout(n16420),.clk(gclk));
	jnot g16171(.din(w_n16171_0[0]),.dout(n16421),.clk(gclk));
	jor g16172(.dina(w_n16421_0[1]),.dinb(n16420),.dout(n16422),.clk(gclk));
	jand g16173(.dina(n16422),.dinb(n16245),.dout(n16423),.clk(gclk));
	jand g16174(.dina(n16423),.dinb(w_n884_33[1]),.dout(n16424),.clk(gclk));
	jor g16175(.dina(w_n16178_0[0]),.dinb(n16424),.dout(n16425),.clk(gclk));
	jand g16176(.dina(n16425),.dinb(n16244),.dout(n16426),.clk(gclk));
	jand g16177(.dina(n16426),.dinb(w_n743_34[1]),.dout(n16427),.clk(gclk));
	jor g16178(.dina(w_n16186_0[0]),.dinb(n16427),.dout(n16428),.clk(gclk));
	jand g16179(.dina(n16428),.dinb(n16243),.dout(n16429),.clk(gclk));
	jand g16180(.dina(n16429),.dinb(w_n635_34[1]),.dout(n16430),.clk(gclk));
	jor g16181(.dina(w_n16194_0[0]),.dinb(n16430),.dout(n16431),.clk(gclk));
	jand g16182(.dina(n16431),.dinb(n16242),.dout(n16432),.clk(gclk));
	jand g16183(.dina(n16432),.dinb(w_n515_35[1]),.dout(n16433),.clk(gclk));
	jnot g16184(.din(w_n16202_0[0]),.dout(n16434),.clk(gclk));
	jor g16185(.dina(w_n16434_0[1]),.dinb(n16433),.dout(n16435),.clk(gclk));
	jand g16186(.dina(n16435),.dinb(n16241),.dout(n16436),.clk(gclk));
	jand g16187(.dina(n16436),.dinb(w_n443_35[1]),.dout(n16437),.clk(gclk));
	jor g16188(.dina(w_n16209_0[0]),.dinb(n16437),.dout(n16438),.clk(gclk));
	jand g16189(.dina(n16438),.dinb(n16240),.dout(n16439),.clk(gclk));
	jand g16190(.dina(n16439),.dinb(w_n352_35[2]),.dout(n16440),.clk(gclk));
	jnot g16191(.din(w_n16217_0[0]),.dout(n16441),.clk(gclk));
	jor g16192(.dina(w_n16441_0[1]),.dinb(n16440),.dout(n16442),.clk(gclk));
	jand g16193(.dina(n16442),.dinb(n16239),.dout(n16443),.clk(gclk));
	jand g16194(.dina(n16443),.dinb(w_n294_36[0]),.dout(n16444),.clk(gclk));
	jor g16195(.dina(w_n16224_0[0]),.dinb(n16444),.dout(n16445),.clk(gclk));
	jand g16196(.dina(n16445),.dinb(n16238),.dout(n16446),.clk(gclk));
	jand g16197(.dina(n16446),.dinb(w_n239_36[1]),.dout(n16447),.clk(gclk));
	jnot g16198(.din(w_n16232_0[0]),.dout(n16448),.clk(gclk));
	jor g16199(.dina(w_n16448_0[1]),.dinb(n16447),.dout(n16449),.clk(gclk));
	jand g16200(.dina(n16449),.dinb(n16237),.dout(n16450),.clk(gclk));
	jand g16201(.dina(n16450),.dinb(w_n221_36[2]),.dout(n16451),.clk(gclk));
	jxor g16202(.dina(w_n15609_0[0]),.dinb(w_n239_36[0]),.dout(n16452),.clk(gclk));
	jand g16203(.dina(n16452),.dinb(w_asqrt14_18[0]),.dout(n16453),.clk(gclk));
	jxor g16204(.dina(n16453),.dinb(w_n15614_0[0]),.dout(n16454),.clk(gclk));
	jor g16205(.dina(w_n16454_0[2]),.dinb(n16451),.dout(n16455),.clk(gclk));
	jand g16206(.dina(n16455),.dinb(n16236),.dout(n16456),.clk(gclk));
	jxor g16207(.dina(w_n15616_0[0]),.dinb(w_n221_36[1]),.dout(n16457),.clk(gclk));
	jand g16208(.dina(n16457),.dinb(w_asqrt14_17[2]),.dout(n16458),.clk(gclk));
	jxor g16209(.dina(n16458),.dinb(w_n15622_0[0]),.dout(n16459),.clk(gclk));
	jor g16210(.dina(w_n16459_0[2]),.dinb(w_n16456_0[2]),.dout(n16460),.clk(gclk));
	jand g16211(.dina(w_asqrt14_17[1]),.dinb(w_n15872_0[0]),.dout(n16461),.clk(gclk));
	jor g16212(.dina(n16461),.dinb(w_n15631_0[0]),.dout(n16462),.clk(gclk));
	jor g16213(.dina(w_n16462_0[1]),.dinb(w_n16460_0[1]),.dout(n16463),.clk(gclk));
	jand g16214(.dina(n16463),.dinb(w_n218_15[1]),.dout(n16464),.clk(gclk));
	jand g16215(.dina(w_n15878_17[1]),.dinb(w_n15264_0[0]),.dout(n16465),.clk(gclk));
	jand g16216(.dina(w_n16459_0[1]),.dinb(w_n16456_0[1]),.dout(n16466),.clk(gclk));
	jor g16217(.dina(w_n16466_0[2]),.dinb(w_n16465_0[1]),.dout(n16467),.clk(gclk));
	jand g16218(.dina(w_n15878_17[0]),.dinb(w_n15624_0[0]),.dout(n16468),.clk(gclk));
	jnot g16219(.din(n16468),.dout(n16469),.clk(gclk));
	jand g16220(.dina(w_n15625_0[0]),.dinb(w_asqrt63_26[2]),.dout(n16470),.clk(gclk));
	jand g16221(.dina(n16470),.dinb(w_n15886_0[0]),.dout(n16471),.clk(gclk));
	jand g16222(.dina(w_n16471_0[1]),.dinb(n16469),.dout(n16472),.clk(gclk));
	jor g16223(.dina(w_n16472_0[1]),.dinb(n16467),.dout(n16473),.clk(gclk));
	jor g16224(.dina(n16473),.dinb(w_n16464_0[1]),.dout(asqrt_fa_14),.clk(gclk));
	jor g16225(.dina(w_n16234_0[1]),.dinb(w_asqrt62_21[0]),.dout(n16475),.clk(gclk));
	jnot g16226(.din(w_n16454_0[1]),.dout(n16476),.clk(gclk));
	jand g16227(.dina(n16476),.dinb(n16475),.dout(n16477),.clk(gclk));
	jor g16228(.dina(n16477),.dinb(w_n16235_0[0]),.dout(n16478),.clk(gclk));
	jnot g16229(.din(w_n16459_0[0]),.dout(n16479),.clk(gclk));
	jand g16230(.dina(w_n16479_0[1]),.dinb(w_n16478_0[1]),.dout(n16480),.clk(gclk));
	jnot g16231(.din(w_n16462_0[0]),.dout(n16481),.clk(gclk));
	jand g16232(.dina(n16481),.dinb(w_n16480_0[1]),.dout(n16482),.clk(gclk));
	jor g16233(.dina(n16482),.dinb(w_asqrt63_26[1]),.dout(n16483),.clk(gclk));
	jnot g16234(.din(w_n16465_0[0]),.dout(n16484),.clk(gclk));
	jor g16235(.dina(w_n16479_0[0]),.dinb(w_n16478_0[0]),.dout(n16485),.clk(gclk));
	jand g16236(.dina(w_n16485_0[2]),.dinb(n16484),.dout(n16486),.clk(gclk));
	jnot g16237(.din(w_n16472_0[0]),.dout(n16487),.clk(gclk));
	jand g16238(.dina(n16487),.dinb(n16486),.dout(n16488),.clk(gclk));
	jand g16239(.dina(n16488),.dinb(n16483),.dout(n16489),.clk(gclk));
	jxor g16240(.dina(w_n16234_0[0]),.dinb(w_n221_36[0]),.dout(n16490),.clk(gclk));
	jor g16241(.dina(n16490),.dinb(w_n16489_39[2]),.dout(n16491),.clk(gclk));
	jxor g16242(.dina(n16491),.dinb(w_n16454_0[0]),.dout(n16492),.clk(gclk));
	jnot g16243(.din(w_n16492_0[1]),.dout(n16493),.clk(gclk));
	jnot g16244(.din(w_a24_0[2]),.dout(n16494),.clk(gclk));
	jnot g16245(.din(w_a25_0[1]),.dout(n16495),.clk(gclk));
	jand g16246(.dina(w_n16495_0[1]),.dinb(w_n16494_1[2]),.dout(n16496),.clk(gclk));
	jand g16247(.dina(w_n16496_0[2]),.dinb(w_n15642_1[0]),.dout(n16497),.clk(gclk));
	jnot g16248(.din(w_n16497_0[1]),.dout(n16498),.clk(gclk));
	jor g16249(.dina(w_n16489_39[1]),.dinb(w_n15642_0[2]),.dout(n16499),.clk(gclk));
	jand g16250(.dina(n16499),.dinb(n16498),.dout(n16500),.clk(gclk));
	jor g16251(.dina(w_n16500_0[2]),.dinb(w_n15878_16[2]),.dout(n16501),.clk(gclk));
	jand g16252(.dina(w_n16500_0[1]),.dinb(w_n15878_16[1]),.dout(n16502),.clk(gclk));
	jor g16253(.dina(w_n16489_39[0]),.dinb(w_a26_1[0]),.dout(n16503),.clk(gclk));
	jand g16254(.dina(n16503),.dinb(w_a27_0[0]),.dout(n16504),.clk(gclk));
	jand g16255(.dina(w_asqrt13_10[1]),.dinb(w_n15644_0[1]),.dout(n16505),.clk(gclk));
	jor g16256(.dina(n16505),.dinb(n16504),.dout(n16506),.clk(gclk));
	jor g16257(.dina(n16506),.dinb(n16502),.dout(n16507),.clk(gclk));
	jand g16258(.dina(n16507),.dinb(w_n16501_0[1]),.dout(n16508),.clk(gclk));
	jor g16259(.dina(w_n16508_0[2]),.dinb(w_n15260_24[1]),.dout(n16509),.clk(gclk));
	jand g16260(.dina(w_n16508_0[1]),.dinb(w_n15260_24[0]),.dout(n16510),.clk(gclk));
	jnot g16261(.din(w_n15644_0[0]),.dout(n16511),.clk(gclk));
	jor g16262(.dina(w_n16489_38[2]),.dinb(n16511),.dout(n16512),.clk(gclk));
	jor g16263(.dina(w_n16471_0[0]),.dinb(w_n15878_16[0]),.dout(n16513),.clk(gclk));
	jor g16264(.dina(n16513),.dinb(w_n16464_0[0]),.dout(n16514),.clk(gclk));
	jor g16265(.dina(n16514),.dinb(w_n16466_0[1]),.dout(n16515),.clk(gclk));
	jand g16266(.dina(n16515),.dinb(w_n16512_0[1]),.dout(n16516),.clk(gclk));
	jxor g16267(.dina(n16516),.dinb(w_n15265_0[1]),.dout(n16517),.clk(gclk));
	jor g16268(.dina(w_n16517_0[2]),.dinb(n16510),.dout(n16518),.clk(gclk));
	jand g16269(.dina(n16518),.dinb(w_n16509_0[1]),.dout(n16519),.clk(gclk));
	jor g16270(.dina(w_n16519_0[2]),.dinb(w_n14674_17[1]),.dout(n16520),.clk(gclk));
	jand g16271(.dina(w_n16519_0[1]),.dinb(w_n14674_17[0]),.dout(n16521),.clk(gclk));
	jxor g16272(.dina(w_n15646_0[0]),.dinb(w_n15260_23[2]),.dout(n16522),.clk(gclk));
	jor g16273(.dina(n16522),.dinb(w_n16489_38[1]),.dout(n16523),.clk(gclk));
	jxor g16274(.dina(n16523),.dinb(w_n16291_0[0]),.dout(n16524),.clk(gclk));
	jnot g16275(.din(w_n16524_0[2]),.dout(n16525),.clk(gclk));
	jor g16276(.dina(n16525),.dinb(n16521),.dout(n16526),.clk(gclk));
	jand g16277(.dina(n16526),.dinb(w_n16520_0[1]),.dout(n16527),.clk(gclk));
	jor g16278(.dina(w_n16527_0[2]),.dinb(w_n14078_24[2]),.dout(n16528),.clk(gclk));
	jand g16279(.dina(w_n16527_0[1]),.dinb(w_n14078_24[1]),.dout(n16529),.clk(gclk));
	jxor g16280(.dina(w_n15882_0[0]),.dinb(w_n14674_16[2]),.dout(n16530),.clk(gclk));
	jor g16281(.dina(n16530),.dinb(w_n16489_38[0]),.dout(n16531),.clk(gclk));
	jxor g16282(.dina(n16531),.dinb(w_n15892_0[0]),.dout(n16532),.clk(gclk));
	jor g16283(.dina(w_n16532_0[2]),.dinb(n16529),.dout(n16533),.clk(gclk));
	jand g16284(.dina(n16533),.dinb(w_n16528_0[1]),.dout(n16534),.clk(gclk));
	jor g16285(.dina(w_n16534_0[2]),.dinb(w_n13515_18[1]),.dout(n16535),.clk(gclk));
	jand g16286(.dina(w_n16534_0[1]),.dinb(w_n13515_18[0]),.dout(n16536),.clk(gclk));
	jxor g16287(.dina(w_n15894_0[0]),.dinb(w_n14078_24[0]),.dout(n16537),.clk(gclk));
	jor g16288(.dina(n16537),.dinb(w_n16489_37[2]),.dout(n16538),.clk(gclk));
	jxor g16289(.dina(n16538),.dinb(w_n15899_0[0]),.dout(n16539),.clk(gclk));
	jor g16290(.dina(w_n16539_0[2]),.dinb(n16536),.dout(n16540),.clk(gclk));
	jand g16291(.dina(n16540),.dinb(w_n16535_0[1]),.dout(n16541),.clk(gclk));
	jor g16292(.dina(w_n16541_0[2]),.dinb(w_n12947_25[1]),.dout(n16542),.clk(gclk));
	jand g16293(.dina(w_n16541_0[1]),.dinb(w_n12947_25[0]),.dout(n16543),.clk(gclk));
	jxor g16294(.dina(w_n15901_0[0]),.dinb(w_n13515_17[2]),.dout(n16544),.clk(gclk));
	jor g16295(.dina(n16544),.dinb(w_n16489_37[1]),.dout(n16545),.clk(gclk));
	jxor g16296(.dina(n16545),.dinb(w_n16302_0[0]),.dout(n16546),.clk(gclk));
	jnot g16297(.din(w_n16546_0[2]),.dout(n16547),.clk(gclk));
	jor g16298(.dina(n16547),.dinb(n16543),.dout(n16548),.clk(gclk));
	jand g16299(.dina(n16548),.dinb(w_n16542_0[1]),.dout(n16549),.clk(gclk));
	jor g16300(.dina(w_n16549_0[2]),.dinb(w_n12410_19[0]),.dout(n16550),.clk(gclk));
	jand g16301(.dina(w_n16549_0[1]),.dinb(w_n12410_18[2]),.dout(n16551),.clk(gclk));
	jxor g16302(.dina(w_n15908_0[0]),.dinb(w_n12947_24[2]),.dout(n16552),.clk(gclk));
	jor g16303(.dina(n16552),.dinb(w_n16489_37[0]),.dout(n16553),.clk(gclk));
	jxor g16304(.dina(n16553),.dinb(w_n16306_0[0]),.dout(n16554),.clk(gclk));
	jnot g16305(.din(w_n16554_0[2]),.dout(n16555),.clk(gclk));
	jor g16306(.dina(n16555),.dinb(n16551),.dout(n16556),.clk(gclk));
	jand g16307(.dina(n16556),.dinb(w_n16550_0[1]),.dout(n16557),.clk(gclk));
	jor g16308(.dina(w_n16557_0[2]),.dinb(w_n11858_25[2]),.dout(n16558),.clk(gclk));
	jand g16309(.dina(w_n16557_0[1]),.dinb(w_n11858_25[1]),.dout(n16559),.clk(gclk));
	jxor g16310(.dina(w_n15915_0[0]),.dinb(w_n12410_18[1]),.dout(n16560),.clk(gclk));
	jor g16311(.dina(n16560),.dinb(w_n16489_36[2]),.dout(n16561),.clk(gclk));
	jxor g16312(.dina(n16561),.dinb(w_n15921_0[0]),.dout(n16562),.clk(gclk));
	jor g16313(.dina(w_n16562_0[2]),.dinb(n16559),.dout(n16563),.clk(gclk));
	jand g16314(.dina(n16563),.dinb(w_n16558_0[1]),.dout(n16564),.clk(gclk));
	jor g16315(.dina(w_n16564_0[2]),.dinb(w_n11347_19[2]),.dout(n16565),.clk(gclk));
	jand g16316(.dina(w_n16564_0[1]),.dinb(w_n11347_19[1]),.dout(n16566),.clk(gclk));
	jxor g16317(.dina(w_n15923_0[0]),.dinb(w_n11858_25[0]),.dout(n16567),.clk(gclk));
	jor g16318(.dina(n16567),.dinb(w_n16489_36[1]),.dout(n16568),.clk(gclk));
	jxor g16319(.dina(n16568),.dinb(w_n16313_0[0]),.dout(n16569),.clk(gclk));
	jnot g16320(.din(w_n16569_0[2]),.dout(n16570),.clk(gclk));
	jor g16321(.dina(n16570),.dinb(n16566),.dout(n16571),.clk(gclk));
	jand g16322(.dina(n16571),.dinb(w_n16565_0[1]),.dout(n16572),.clk(gclk));
	jor g16323(.dina(w_n16572_0[2]),.dinb(w_n10824_26[1]),.dout(n16573),.clk(gclk));
	jand g16324(.dina(w_n16572_0[1]),.dinb(w_n10824_26[0]),.dout(n16574),.clk(gclk));
	jxor g16325(.dina(w_n15930_0[0]),.dinb(w_n11347_19[0]),.dout(n16575),.clk(gclk));
	jor g16326(.dina(n16575),.dinb(w_n16489_36[0]),.dout(n16576),.clk(gclk));
	jxor g16327(.dina(n16576),.dinb(w_n15936_0[0]),.dout(n16577),.clk(gclk));
	jor g16328(.dina(w_n16577_0[2]),.dinb(n16574),.dout(n16578),.clk(gclk));
	jand g16329(.dina(n16578),.dinb(w_n16573_0[1]),.dout(n16579),.clk(gclk));
	jor g16330(.dina(w_n16579_0[2]),.dinb(w_n10328_20[2]),.dout(n16580),.clk(gclk));
	jand g16331(.dina(w_n16579_0[1]),.dinb(w_n10328_20[1]),.dout(n16581),.clk(gclk));
	jxor g16332(.dina(w_n15938_0[0]),.dinb(w_n10824_25[2]),.dout(n16582),.clk(gclk));
	jor g16333(.dina(n16582),.dinb(w_n16489_35[2]),.dout(n16583),.clk(gclk));
	jxor g16334(.dina(n16583),.dinb(w_n16320_0[0]),.dout(n16584),.clk(gclk));
	jnot g16335(.din(w_n16584_0[2]),.dout(n16585),.clk(gclk));
	jor g16336(.dina(n16585),.dinb(n16581),.dout(n16586),.clk(gclk));
	jand g16337(.dina(n16586),.dinb(w_n16580_0[1]),.dout(n16587),.clk(gclk));
	jor g16338(.dina(w_n16587_0[2]),.dinb(w_n9832_27[0]),.dout(n16588),.clk(gclk));
	jand g16339(.dina(w_n16587_0[1]),.dinb(w_n9832_26[2]),.dout(n16589),.clk(gclk));
	jxor g16340(.dina(w_n15945_0[0]),.dinb(w_n10328_20[0]),.dout(n16590),.clk(gclk));
	jor g16341(.dina(n16590),.dinb(w_n16489_35[1]),.dout(n16591),.clk(gclk));
	jxor g16342(.dina(n16591),.dinb(w_n15951_0[0]),.dout(n16592),.clk(gclk));
	jor g16343(.dina(w_n16592_0[2]),.dinb(n16589),.dout(n16593),.clk(gclk));
	jand g16344(.dina(n16593),.dinb(w_n16588_0[1]),.dout(n16594),.clk(gclk));
	jor g16345(.dina(w_n16594_0[2]),.dinb(w_n9369_21[2]),.dout(n16595),.clk(gclk));
	jand g16346(.dina(w_n16594_0[1]),.dinb(w_n9369_21[1]),.dout(n16596),.clk(gclk));
	jxor g16347(.dina(w_n15953_0[0]),.dinb(w_n9832_26[1]),.dout(n16597),.clk(gclk));
	jor g16348(.dina(n16597),.dinb(w_n16489_35[0]),.dout(n16598),.clk(gclk));
	jxor g16349(.dina(n16598),.dinb(w_n15959_0[0]),.dout(n16599),.clk(gclk));
	jor g16350(.dina(w_n16599_0[2]),.dinb(n16596),.dout(n16600),.clk(gclk));
	jand g16351(.dina(n16600),.dinb(w_n16595_0[1]),.dout(n16601),.clk(gclk));
	jor g16352(.dina(w_n16601_0[2]),.dinb(w_n8890_27[1]),.dout(n16602),.clk(gclk));
	jand g16353(.dina(w_n16601_0[1]),.dinb(w_n8890_27[0]),.dout(n16603),.clk(gclk));
	jxor g16354(.dina(w_n15961_0[0]),.dinb(w_n9369_21[0]),.dout(n16604),.clk(gclk));
	jor g16355(.dina(n16604),.dinb(w_n16489_34[2]),.dout(n16605),.clk(gclk));
	jxor g16356(.dina(n16605),.dinb(w_n15967_0[0]),.dout(n16606),.clk(gclk));
	jor g16357(.dina(w_n16606_0[2]),.dinb(n16603),.dout(n16607),.clk(gclk));
	jand g16358(.dina(n16607),.dinb(w_n16602_0[1]),.dout(n16608),.clk(gclk));
	jor g16359(.dina(w_n16608_0[2]),.dinb(w_n8449_22[1]),.dout(n16609),.clk(gclk));
	jand g16360(.dina(w_n16608_0[1]),.dinb(w_n8449_22[0]),.dout(n16610),.clk(gclk));
	jxor g16361(.dina(w_n15969_0[0]),.dinb(w_n8890_26[2]),.dout(n16611),.clk(gclk));
	jor g16362(.dina(n16611),.dinb(w_n16489_34[1]),.dout(n16612),.clk(gclk));
	jxor g16363(.dina(n16612),.dinb(w_n16333_0[0]),.dout(n16613),.clk(gclk));
	jnot g16364(.din(w_n16613_0[2]),.dout(n16614),.clk(gclk));
	jor g16365(.dina(n16614),.dinb(n16610),.dout(n16615),.clk(gclk));
	jand g16366(.dina(n16615),.dinb(w_n16609_0[1]),.dout(n16616),.clk(gclk));
	jor g16367(.dina(w_n16616_0[2]),.dinb(w_n8003_28[0]),.dout(n16617),.clk(gclk));
	jand g16368(.dina(w_n16616_0[1]),.dinb(w_n8003_27[2]),.dout(n16618),.clk(gclk));
	jxor g16369(.dina(w_n15976_0[0]),.dinb(w_n8449_21[2]),.dout(n16619),.clk(gclk));
	jor g16370(.dina(n16619),.dinb(w_n16489_34[0]),.dout(n16620),.clk(gclk));
	jxor g16371(.dina(n16620),.dinb(w_n15982_0[0]),.dout(n16621),.clk(gclk));
	jor g16372(.dina(w_n16621_0[2]),.dinb(n16618),.dout(n16622),.clk(gclk));
	jand g16373(.dina(n16622),.dinb(w_n16617_0[1]),.dout(n16623),.clk(gclk));
	jor g16374(.dina(w_n16623_0[2]),.dinb(w_n7581_23[1]),.dout(n16624),.clk(gclk));
	jand g16375(.dina(w_n16623_0[1]),.dinb(w_n7581_23[0]),.dout(n16625),.clk(gclk));
	jxor g16376(.dina(w_n15984_0[0]),.dinb(w_n8003_27[1]),.dout(n16626),.clk(gclk));
	jor g16377(.dina(n16626),.dinb(w_n16489_33[2]),.dout(n16627),.clk(gclk));
	jxor g16378(.dina(n16627),.dinb(w_n16340_0[0]),.dout(n16628),.clk(gclk));
	jnot g16379(.din(w_n16628_0[2]),.dout(n16629),.clk(gclk));
	jor g16380(.dina(n16629),.dinb(n16625),.dout(n16630),.clk(gclk));
	jand g16381(.dina(n16630),.dinb(w_n16624_0[1]),.dout(n16631),.clk(gclk));
	jor g16382(.dina(w_n16631_0[2]),.dinb(w_n7154_28[1]),.dout(n16632),.clk(gclk));
	jand g16383(.dina(w_n16631_0[1]),.dinb(w_n7154_28[0]),.dout(n16633),.clk(gclk));
	jxor g16384(.dina(w_n15991_0[0]),.dinb(w_n7581_22[2]),.dout(n16634),.clk(gclk));
	jor g16385(.dina(n16634),.dinb(w_n16489_33[1]),.dout(n16635),.clk(gclk));
	jxor g16386(.dina(n16635),.dinb(w_n15997_0[0]),.dout(n16636),.clk(gclk));
	jor g16387(.dina(w_n16636_0[2]),.dinb(n16633),.dout(n16637),.clk(gclk));
	jand g16388(.dina(n16637),.dinb(w_n16632_0[1]),.dout(n16638),.clk(gclk));
	jor g16389(.dina(w_n16638_0[2]),.dinb(w_n6758_24[0]),.dout(n16639),.clk(gclk));
	jand g16390(.dina(w_n16638_0[1]),.dinb(w_n6758_23[2]),.dout(n16640),.clk(gclk));
	jxor g16391(.dina(w_n15999_0[0]),.dinb(w_n7154_27[2]),.dout(n16641),.clk(gclk));
	jor g16392(.dina(n16641),.dinb(w_n16489_33[0]),.dout(n16642),.clk(gclk));
	jxor g16393(.dina(n16642),.dinb(w_n16347_0[0]),.dout(n16643),.clk(gclk));
	jnot g16394(.din(w_n16643_0[2]),.dout(n16644),.clk(gclk));
	jor g16395(.dina(n16644),.dinb(n16640),.dout(n16645),.clk(gclk));
	jand g16396(.dina(n16645),.dinb(w_n16639_0[1]),.dout(n16646),.clk(gclk));
	jor g16397(.dina(w_n16646_0[2]),.dinb(w_n6357_28[2]),.dout(n16647),.clk(gclk));
	jand g16398(.dina(w_n16646_0[1]),.dinb(w_n6357_28[1]),.dout(n16648),.clk(gclk));
	jxor g16399(.dina(w_n16006_0[0]),.dinb(w_n6758_23[1]),.dout(n16649),.clk(gclk));
	jor g16400(.dina(n16649),.dinb(w_n16489_32[2]),.dout(n16650),.clk(gclk));
	jxor g16401(.dina(n16650),.dinb(w_n16012_0[0]),.dout(n16651),.clk(gclk));
	jor g16402(.dina(w_n16651_0[2]),.dinb(n16648),.dout(n16652),.clk(gclk));
	jand g16403(.dina(n16652),.dinb(w_n16647_0[1]),.dout(n16653),.clk(gclk));
	jor g16404(.dina(w_n16653_0[2]),.dinb(w_n5989_24[2]),.dout(n16654),.clk(gclk));
	jand g16405(.dina(w_n16653_0[1]),.dinb(w_n5989_24[1]),.dout(n16655),.clk(gclk));
	jxor g16406(.dina(w_n16014_0[0]),.dinb(w_n6357_28[0]),.dout(n16656),.clk(gclk));
	jor g16407(.dina(n16656),.dinb(w_n16489_32[1]),.dout(n16657),.clk(gclk));
	jxor g16408(.dina(n16657),.dinb(w_n16354_0[0]),.dout(n16658),.clk(gclk));
	jnot g16409(.din(w_n16658_0[2]),.dout(n16659),.clk(gclk));
	jor g16410(.dina(n16659),.dinb(n16655),.dout(n16660),.clk(gclk));
	jand g16411(.dina(n16660),.dinb(w_n16654_0[1]),.dout(n16661),.clk(gclk));
	jor g16412(.dina(w_n16661_0[2]),.dinb(w_n5606_29[0]),.dout(n16662),.clk(gclk));
	jand g16413(.dina(w_n16661_0[1]),.dinb(w_n5606_28[2]),.dout(n16663),.clk(gclk));
	jxor g16414(.dina(w_n16021_0[0]),.dinb(w_n5989_24[0]),.dout(n16664),.clk(gclk));
	jor g16415(.dina(n16664),.dinb(w_n16489_32[0]),.dout(n16665),.clk(gclk));
	jxor g16416(.dina(n16665),.dinb(w_n16027_0[0]),.dout(n16666),.clk(gclk));
	jor g16417(.dina(w_n16666_0[2]),.dinb(n16663),.dout(n16667),.clk(gclk));
	jand g16418(.dina(n16667),.dinb(w_n16662_0[1]),.dout(n16668),.clk(gclk));
	jor g16419(.dina(w_n16668_0[2]),.dinb(w_n5259_25[2]),.dout(n16669),.clk(gclk));
	jand g16420(.dina(w_n16668_0[1]),.dinb(w_n5259_25[1]),.dout(n16670),.clk(gclk));
	jxor g16421(.dina(w_n16029_0[0]),.dinb(w_n5606_28[1]),.dout(n16671),.clk(gclk));
	jor g16422(.dina(n16671),.dinb(w_n16489_31[2]),.dout(n16672),.clk(gclk));
	jxor g16423(.dina(n16672),.dinb(w_n16035_0[0]),.dout(n16673),.clk(gclk));
	jor g16424(.dina(w_n16673_0[2]),.dinb(n16670),.dout(n16674),.clk(gclk));
	jand g16425(.dina(n16674),.dinb(w_n16669_0[1]),.dout(n16675),.clk(gclk));
	jor g16426(.dina(w_n16675_0[2]),.dinb(w_n4902_29[2]),.dout(n16676),.clk(gclk));
	jand g16427(.dina(w_n16675_0[1]),.dinb(w_n4902_29[1]),.dout(n16677),.clk(gclk));
	jxor g16428(.dina(w_n16037_0[0]),.dinb(w_n5259_25[0]),.dout(n16678),.clk(gclk));
	jor g16429(.dina(n16678),.dinb(w_n16489_31[1]),.dout(n16679),.clk(gclk));
	jxor g16430(.dina(n16679),.dinb(w_n16043_0[0]),.dout(n16680),.clk(gclk));
	jor g16431(.dina(w_n16680_0[2]),.dinb(n16677),.dout(n16681),.clk(gclk));
	jand g16432(.dina(n16681),.dinb(w_n16676_0[1]),.dout(n16682),.clk(gclk));
	jor g16433(.dina(w_n16682_0[2]),.dinb(w_n4582_26[2]),.dout(n16683),.clk(gclk));
	jand g16434(.dina(w_n16682_0[1]),.dinb(w_n4582_26[1]),.dout(n16684),.clk(gclk));
	jxor g16435(.dina(w_n16045_0[0]),.dinb(w_n4902_29[0]),.dout(n16685),.clk(gclk));
	jor g16436(.dina(n16685),.dinb(w_n16489_31[0]),.dout(n16686),.clk(gclk));
	jxor g16437(.dina(n16686),.dinb(w_n16367_0[0]),.dout(n16687),.clk(gclk));
	jnot g16438(.din(w_n16687_0[2]),.dout(n16688),.clk(gclk));
	jor g16439(.dina(n16688),.dinb(n16684),.dout(n16689),.clk(gclk));
	jand g16440(.dina(n16689),.dinb(w_n16683_0[1]),.dout(n16690),.clk(gclk));
	jor g16441(.dina(w_n16690_0[2]),.dinb(w_n4249_30[1]),.dout(n16691),.clk(gclk));
	jand g16442(.dina(w_n16690_0[1]),.dinb(w_n4249_30[0]),.dout(n16692),.clk(gclk));
	jxor g16443(.dina(w_n16052_0[0]),.dinb(w_n4582_26[0]),.dout(n16693),.clk(gclk));
	jor g16444(.dina(n16693),.dinb(w_n16489_30[2]),.dout(n16694),.clk(gclk));
	jxor g16445(.dina(n16694),.dinb(w_n16058_0[0]),.dout(n16695),.clk(gclk));
	jor g16446(.dina(w_n16695_0[2]),.dinb(n16692),.dout(n16696),.clk(gclk));
	jand g16447(.dina(n16696),.dinb(w_n16691_0[1]),.dout(n16697),.clk(gclk));
	jor g16448(.dina(w_n16697_0[2]),.dinb(w_n3955_27[1]),.dout(n16698),.clk(gclk));
	jand g16449(.dina(w_n16697_0[1]),.dinb(w_n3955_27[0]),.dout(n16699),.clk(gclk));
	jxor g16450(.dina(w_n16060_0[0]),.dinb(w_n4249_29[2]),.dout(n16700),.clk(gclk));
	jor g16451(.dina(n16700),.dinb(w_n16489_30[1]),.dout(n16701),.clk(gclk));
	jxor g16452(.dina(n16701),.dinb(w_n16374_0[0]),.dout(n16702),.clk(gclk));
	jnot g16453(.din(w_n16702_0[2]),.dout(n16703),.clk(gclk));
	jor g16454(.dina(n16703),.dinb(n16699),.dout(n16704),.clk(gclk));
	jand g16455(.dina(n16704),.dinb(w_n16698_0[1]),.dout(n16705),.clk(gclk));
	jor g16456(.dina(w_n16705_0[2]),.dinb(w_n3642_30[2]),.dout(n16706),.clk(gclk));
	jand g16457(.dina(w_n16705_0[1]),.dinb(w_n3642_30[1]),.dout(n16707),.clk(gclk));
	jxor g16458(.dina(w_n16067_0[0]),.dinb(w_n3955_26[2]),.dout(n16708),.clk(gclk));
	jor g16459(.dina(n16708),.dinb(w_n16489_30[0]),.dout(n16709),.clk(gclk));
	jxor g16460(.dina(n16709),.dinb(w_n16073_0[0]),.dout(n16710),.clk(gclk));
	jor g16461(.dina(w_n16710_0[2]),.dinb(n16707),.dout(n16711),.clk(gclk));
	jand g16462(.dina(n16711),.dinb(w_n16706_0[1]),.dout(n16712),.clk(gclk));
	jor g16463(.dina(w_n16712_0[2]),.dinb(w_n3368_28[0]),.dout(n16713),.clk(gclk));
	jand g16464(.dina(w_n16712_0[1]),.dinb(w_n3368_27[2]),.dout(n16714),.clk(gclk));
	jxor g16465(.dina(w_n16075_0[0]),.dinb(w_n3642_30[0]),.dout(n16715),.clk(gclk));
	jor g16466(.dina(n16715),.dinb(w_n16489_29[2]),.dout(n16716),.clk(gclk));
	jxor g16467(.dina(n16716),.dinb(w_n16081_0[0]),.dout(n16717),.clk(gclk));
	jor g16468(.dina(w_n16717_0[2]),.dinb(n16714),.dout(n16718),.clk(gclk));
	jand g16469(.dina(n16718),.dinb(w_n16713_0[1]),.dout(n16719),.clk(gclk));
	jor g16470(.dina(w_n16719_0[2]),.dinb(w_n3089_31[1]),.dout(n16720),.clk(gclk));
	jand g16471(.dina(w_n16719_0[1]),.dinb(w_n3089_31[0]),.dout(n16721),.clk(gclk));
	jxor g16472(.dina(w_n16083_0[0]),.dinb(w_n3368_27[1]),.dout(n16722),.clk(gclk));
	jor g16473(.dina(n16722),.dinb(w_n16489_29[1]),.dout(n16723),.clk(gclk));
	jxor g16474(.dina(n16723),.dinb(w_n16089_0[0]),.dout(n16724),.clk(gclk));
	jor g16475(.dina(w_n16724_0[2]),.dinb(n16721),.dout(n16725),.clk(gclk));
	jand g16476(.dina(n16725),.dinb(w_n16720_0[1]),.dout(n16726),.clk(gclk));
	jor g16477(.dina(w_n16726_0[2]),.dinb(w_n2833_29[0]),.dout(n16727),.clk(gclk));
	jand g16478(.dina(w_n16726_0[1]),.dinb(w_n2833_28[2]),.dout(n16728),.clk(gclk));
	jxor g16479(.dina(w_n16091_0[0]),.dinb(w_n3089_30[2]),.dout(n16729),.clk(gclk));
	jor g16480(.dina(n16729),.dinb(w_n16489_29[0]),.dout(n16730),.clk(gclk));
	jxor g16481(.dina(n16730),.dinb(w_n16387_0[0]),.dout(n16731),.clk(gclk));
	jnot g16482(.din(w_n16731_0[2]),.dout(n16732),.clk(gclk));
	jor g16483(.dina(n16732),.dinb(n16728),.dout(n16733),.clk(gclk));
	jand g16484(.dina(n16733),.dinb(w_n16727_0[1]),.dout(n16734),.clk(gclk));
	jor g16485(.dina(w_n16734_0[2]),.dinb(w_n2572_31[2]),.dout(n16735),.clk(gclk));
	jand g16486(.dina(w_n16734_0[1]),.dinb(w_n2572_31[1]),.dout(n16736),.clk(gclk));
	jxor g16487(.dina(w_n16098_0[0]),.dinb(w_n2833_28[1]),.dout(n16737),.clk(gclk));
	jor g16488(.dina(n16737),.dinb(w_n16489_28[2]),.dout(n16738),.clk(gclk));
	jxor g16489(.dina(n16738),.dinb(w_n16104_0[0]),.dout(n16739),.clk(gclk));
	jor g16490(.dina(w_n16739_0[2]),.dinb(n16736),.dout(n16740),.clk(gclk));
	jand g16491(.dina(n16740),.dinb(w_n16735_0[1]),.dout(n16741),.clk(gclk));
	jor g16492(.dina(w_n16741_0[2]),.dinb(w_n2345_29[2]),.dout(n16742),.clk(gclk));
	jand g16493(.dina(w_n16741_0[1]),.dinb(w_n2345_29[1]),.dout(n16743),.clk(gclk));
	jxor g16494(.dina(w_n16106_0[0]),.dinb(w_n2572_31[0]),.dout(n16744),.clk(gclk));
	jor g16495(.dina(n16744),.dinb(w_n16489_28[1]),.dout(n16745),.clk(gclk));
	jxor g16496(.dina(n16745),.dinb(w_n16394_0[0]),.dout(n16746),.clk(gclk));
	jnot g16497(.din(w_n16746_0[2]),.dout(n16747),.clk(gclk));
	jor g16498(.dina(n16747),.dinb(n16743),.dout(n16748),.clk(gclk));
	jand g16499(.dina(n16748),.dinb(w_n16742_0[1]),.dout(n16749),.clk(gclk));
	jor g16500(.dina(w_n16749_0[2]),.dinb(w_n2108_32[1]),.dout(n16750),.clk(gclk));
	jand g16501(.dina(w_n16749_0[1]),.dinb(w_n2108_32[0]),.dout(n16751),.clk(gclk));
	jxor g16502(.dina(w_n16113_0[0]),.dinb(w_n2345_29[0]),.dout(n16752),.clk(gclk));
	jor g16503(.dina(n16752),.dinb(w_n16489_28[0]),.dout(n16753),.clk(gclk));
	jxor g16504(.dina(n16753),.dinb(w_n16119_0[0]),.dout(n16754),.clk(gclk));
	jor g16505(.dina(w_n16754_0[2]),.dinb(n16751),.dout(n16755),.clk(gclk));
	jand g16506(.dina(n16755),.dinb(w_n16750_0[1]),.dout(n16756),.clk(gclk));
	jor g16507(.dina(w_n16756_0[2]),.dinb(w_n1912_30[2]),.dout(n16757),.clk(gclk));
	jand g16508(.dina(w_n16756_0[1]),.dinb(w_n1912_30[1]),.dout(n16758),.clk(gclk));
	jxor g16509(.dina(w_n16121_0[0]),.dinb(w_n2108_31[2]),.dout(n16759),.clk(gclk));
	jor g16510(.dina(n16759),.dinb(w_n16489_27[2]),.dout(n16760),.clk(gclk));
	jxor g16511(.dina(n16760),.dinb(w_n16127_0[0]),.dout(n16761),.clk(gclk));
	jor g16512(.dina(w_n16761_0[2]),.dinb(n16758),.dout(n16762),.clk(gclk));
	jand g16513(.dina(n16762),.dinb(w_n16757_0[1]),.dout(n16763),.clk(gclk));
	jor g16514(.dina(w_n16763_0[2]),.dinb(w_n1699_33[0]),.dout(n16764),.clk(gclk));
	jand g16515(.dina(w_n16763_0[1]),.dinb(w_n1699_32[2]),.dout(n16765),.clk(gclk));
	jxor g16516(.dina(w_n16129_0[0]),.dinb(w_n1912_30[0]),.dout(n16766),.clk(gclk));
	jor g16517(.dina(n16766),.dinb(w_n16489_27[1]),.dout(n16767),.clk(gclk));
	jxor g16518(.dina(n16767),.dinb(w_n16404_0[0]),.dout(n16768),.clk(gclk));
	jnot g16519(.din(w_n16768_0[2]),.dout(n16769),.clk(gclk));
	jor g16520(.dina(n16769),.dinb(n16765),.dout(n16770),.clk(gclk));
	jand g16521(.dina(n16770),.dinb(w_n16764_0[1]),.dout(n16771),.clk(gclk));
	jor g16522(.dina(w_n16771_0[2]),.dinb(w_n1516_31[1]),.dout(n16772),.clk(gclk));
	jxor g16523(.dina(w_n16136_0[0]),.dinb(w_n1699_32[1]),.dout(n16773),.clk(gclk));
	jor g16524(.dina(n16773),.dinb(w_n16489_27[0]),.dout(n16774),.clk(gclk));
	jxor g16525(.dina(n16774),.dinb(w_n16250_0[0]),.dout(n16775),.clk(gclk));
	jnot g16526(.din(w_n16775_0[2]),.dout(n16776),.clk(gclk));
	jand g16527(.dina(w_n16771_0[1]),.dinb(w_n1516_31[0]),.dout(n16777),.clk(gclk));
	jor g16528(.dina(n16777),.dinb(n16776),.dout(n16778),.clk(gclk));
	jand g16529(.dina(n16778),.dinb(w_n16772_0[1]),.dout(n16779),.clk(gclk));
	jor g16530(.dina(w_n16779_0[2]),.dinb(w_n1332_33[0]),.dout(n16780),.clk(gclk));
	jand g16531(.dina(w_n16779_0[1]),.dinb(w_n1332_32[2]),.dout(n16781),.clk(gclk));
	jxor g16532(.dina(w_n16143_0[0]),.dinb(w_n1516_30[2]),.dout(n16782),.clk(gclk));
	jor g16533(.dina(n16782),.dinb(w_n16489_26[2]),.dout(n16783),.clk(gclk));
	jxor g16534(.dina(n16783),.dinb(w_n16149_0[0]),.dout(n16784),.clk(gclk));
	jor g16535(.dina(w_n16784_0[2]),.dinb(n16781),.dout(n16785),.clk(gclk));
	jand g16536(.dina(n16785),.dinb(w_n16780_0[1]),.dout(n16786),.clk(gclk));
	jor g16537(.dina(w_n16786_0[2]),.dinb(w_n1173_32[0]),.dout(n16787),.clk(gclk));
	jand g16538(.dina(w_n16786_0[1]),.dinb(w_n1173_31[2]),.dout(n16788),.clk(gclk));
	jxor g16539(.dina(w_n16151_0[0]),.dinb(w_n1332_32[1]),.dout(n16789),.clk(gclk));
	jor g16540(.dina(n16789),.dinb(w_n16489_26[1]),.dout(n16790),.clk(gclk));
	jxor g16541(.dina(n16790),.dinb(w_n16414_0[0]),.dout(n16791),.clk(gclk));
	jnot g16542(.din(w_n16791_0[2]),.dout(n16792),.clk(gclk));
	jor g16543(.dina(n16792),.dinb(n16788),.dout(n16793),.clk(gclk));
	jand g16544(.dina(n16793),.dinb(w_n16787_0[1]),.dout(n16794),.clk(gclk));
	jor g16545(.dina(w_n16794_0[2]),.dinb(w_n1008_34[0]),.dout(n16795),.clk(gclk));
	jand g16546(.dina(w_n16794_0[1]),.dinb(w_n1008_33[2]),.dout(n16796),.clk(gclk));
	jxor g16547(.dina(w_n16158_0[0]),.dinb(w_n1173_31[1]),.dout(n16797),.clk(gclk));
	jor g16548(.dina(n16797),.dinb(w_n16489_26[0]),.dout(n16798),.clk(gclk));
	jxor g16549(.dina(n16798),.dinb(w_n16164_0[0]),.dout(n16799),.clk(gclk));
	jor g16550(.dina(w_n16799_0[2]),.dinb(n16796),.dout(n16800),.clk(gclk));
	jand g16551(.dina(n16800),.dinb(w_n16795_0[1]),.dout(n16801),.clk(gclk));
	jor g16552(.dina(w_n16801_0[2]),.dinb(w_n884_33[0]),.dout(n16802),.clk(gclk));
	jand g16553(.dina(w_n16801_0[1]),.dinb(w_n884_32[2]),.dout(n16803),.clk(gclk));
	jxor g16554(.dina(w_n16166_0[0]),.dinb(w_n1008_33[1]),.dout(n16804),.clk(gclk));
	jor g16555(.dina(n16804),.dinb(w_n16489_25[2]),.dout(n16805),.clk(gclk));
	jxor g16556(.dina(n16805),.dinb(w_n16421_0[0]),.dout(n16806),.clk(gclk));
	jnot g16557(.din(w_n16806_0[2]),.dout(n16807),.clk(gclk));
	jor g16558(.dina(n16807),.dinb(n16803),.dout(n16808),.clk(gclk));
	jand g16559(.dina(n16808),.dinb(w_n16802_0[1]),.dout(n16809),.clk(gclk));
	jor g16560(.dina(w_n16809_0[2]),.dinb(w_n743_34[0]),.dout(n16810),.clk(gclk));
	jand g16561(.dina(w_n16809_0[1]),.dinb(w_n743_33[2]),.dout(n16811),.clk(gclk));
	jxor g16562(.dina(w_n16173_0[0]),.dinb(w_n884_32[1]),.dout(n16812),.clk(gclk));
	jor g16563(.dina(n16812),.dinb(w_n16489_25[1]),.dout(n16813),.clk(gclk));
	jxor g16564(.dina(n16813),.dinb(w_n16179_0[0]),.dout(n16814),.clk(gclk));
	jor g16565(.dina(w_n16814_0[2]),.dinb(n16811),.dout(n16815),.clk(gclk));
	jand g16566(.dina(n16815),.dinb(w_n16810_0[1]),.dout(n16816),.clk(gclk));
	jor g16567(.dina(w_n16816_0[2]),.dinb(w_n635_34[0]),.dout(n16817),.clk(gclk));
	jand g16568(.dina(w_n16816_0[1]),.dinb(w_n635_33[2]),.dout(n16818),.clk(gclk));
	jxor g16569(.dina(w_n16181_0[0]),.dinb(w_n743_33[1]),.dout(n16819),.clk(gclk));
	jor g16570(.dina(n16819),.dinb(w_n16489_25[0]),.dout(n16820),.clk(gclk));
	jxor g16571(.dina(n16820),.dinb(w_n16187_0[0]),.dout(n16821),.clk(gclk));
	jor g16572(.dina(w_n16821_0[2]),.dinb(n16818),.dout(n16822),.clk(gclk));
	jand g16573(.dina(n16822),.dinb(w_n16817_0[1]),.dout(n16823),.clk(gclk));
	jor g16574(.dina(w_n16823_0[2]),.dinb(w_n515_35[0]),.dout(n16824),.clk(gclk));
	jand g16575(.dina(w_n16823_0[1]),.dinb(w_n515_34[2]),.dout(n16825),.clk(gclk));
	jxor g16576(.dina(w_n16189_0[0]),.dinb(w_n635_33[1]),.dout(n16826),.clk(gclk));
	jor g16577(.dina(n16826),.dinb(w_n16489_24[2]),.dout(n16827),.clk(gclk));
	jxor g16578(.dina(n16827),.dinb(w_n16195_0[0]),.dout(n16828),.clk(gclk));
	jor g16579(.dina(w_n16828_0[2]),.dinb(n16825),.dout(n16829),.clk(gclk));
	jand g16580(.dina(n16829),.dinb(w_n16824_0[1]),.dout(n16830),.clk(gclk));
	jor g16581(.dina(w_n16830_0[2]),.dinb(w_n443_35[0]),.dout(n16831),.clk(gclk));
	jand g16582(.dina(w_n16830_0[1]),.dinb(w_n443_34[2]),.dout(n16832),.clk(gclk));
	jxor g16583(.dina(w_n16197_0[0]),.dinb(w_n515_34[1]),.dout(n16833),.clk(gclk));
	jor g16584(.dina(n16833),.dinb(w_n16489_24[1]),.dout(n16834),.clk(gclk));
	jxor g16585(.dina(n16834),.dinb(w_n16434_0[0]),.dout(n16835),.clk(gclk));
	jnot g16586(.din(w_n16835_0[2]),.dout(n16836),.clk(gclk));
	jor g16587(.dina(n16836),.dinb(n16832),.dout(n16837),.clk(gclk));
	jand g16588(.dina(n16837),.dinb(w_n16831_0[1]),.dout(n16838),.clk(gclk));
	jor g16589(.dina(w_n16838_0[2]),.dinb(w_n352_35[1]),.dout(n16839),.clk(gclk));
	jand g16590(.dina(w_n16838_0[1]),.dinb(w_n352_35[0]),.dout(n16840),.clk(gclk));
	jxor g16591(.dina(w_n16204_0[0]),.dinb(w_n443_34[1]),.dout(n16841),.clk(gclk));
	jor g16592(.dina(n16841),.dinb(w_n16489_24[0]),.dout(n16842),.clk(gclk));
	jxor g16593(.dina(n16842),.dinb(w_n16210_0[0]),.dout(n16843),.clk(gclk));
	jor g16594(.dina(w_n16843_0[2]),.dinb(n16840),.dout(n16844),.clk(gclk));
	jand g16595(.dina(n16844),.dinb(w_n16839_0[1]),.dout(n16845),.clk(gclk));
	jor g16596(.dina(w_n16845_0[2]),.dinb(w_n294_35[2]),.dout(n16846),.clk(gclk));
	jand g16597(.dina(w_n16845_0[1]),.dinb(w_n294_35[1]),.dout(n16847),.clk(gclk));
	jxor g16598(.dina(w_n16212_0[0]),.dinb(w_n352_34[2]),.dout(n16848),.clk(gclk));
	jor g16599(.dina(n16848),.dinb(w_n16489_23[2]),.dout(n16849),.clk(gclk));
	jxor g16600(.dina(n16849),.dinb(w_n16441_0[0]),.dout(n16850),.clk(gclk));
	jnot g16601(.din(w_n16850_0[2]),.dout(n16851),.clk(gclk));
	jor g16602(.dina(n16851),.dinb(n16847),.dout(n16852),.clk(gclk));
	jand g16603(.dina(n16852),.dinb(w_n16846_0[1]),.dout(n16853),.clk(gclk));
	jor g16604(.dina(w_n16853_0[2]),.dinb(w_n239_35[2]),.dout(n16854),.clk(gclk));
	jand g16605(.dina(w_n16853_0[1]),.dinb(w_n239_35[1]),.dout(n16855),.clk(gclk));
	jxor g16606(.dina(w_n16219_0[0]),.dinb(w_n294_35[0]),.dout(n16856),.clk(gclk));
	jor g16607(.dina(n16856),.dinb(w_n16489_23[1]),.dout(n16857),.clk(gclk));
	jxor g16608(.dina(n16857),.dinb(w_n16225_0[0]),.dout(n16858),.clk(gclk));
	jor g16609(.dina(w_n16858_0[2]),.dinb(n16855),.dout(n16859),.clk(gclk));
	jand g16610(.dina(n16859),.dinb(w_n16854_0[1]),.dout(n16860),.clk(gclk));
	jor g16611(.dina(w_n16860_0[2]),.dinb(w_n221_35[2]),.dout(n16861),.clk(gclk));
	jand g16612(.dina(w_n16860_0[1]),.dinb(w_n221_35[1]),.dout(n16862),.clk(gclk));
	jxor g16613(.dina(w_n16227_0[0]),.dinb(w_n239_35[0]),.dout(n16863),.clk(gclk));
	jor g16614(.dina(n16863),.dinb(w_n16489_23[0]),.dout(n16864),.clk(gclk));
	jxor g16615(.dina(n16864),.dinb(w_n16448_0[0]),.dout(n16865),.clk(gclk));
	jnot g16616(.din(w_n16865_0[1]),.dout(n16866),.clk(gclk));
	jor g16617(.dina(w_n16866_0[1]),.dinb(n16862),.dout(n16867),.clk(gclk));
	jand g16618(.dina(n16867),.dinb(w_n16861_0[1]),.dout(n16868),.clk(gclk));
	jand g16619(.dina(w_n16868_0[2]),.dinb(w_n16493_0[2]),.dout(n16869),.clk(gclk));
	jor g16620(.dina(w_n16868_0[1]),.dinb(w_n16493_0[1]),.dout(n16871),.clk(gclk));
	jand g16621(.dina(w_asqrt13_10[0]),.dinb(w_n16480_0[0]),.dout(n16872),.clk(gclk));
	jor g16622(.dina(w_n16872_0[1]),.dinb(w_n16871_0[1]),.dout(n16873),.clk(gclk));
	jor g16623(.dina(n16873),.dinb(w_n16466_0[0]),.dout(n16874),.clk(gclk));
	jand g16624(.dina(n16874),.dinb(w_n218_15[0]),.dout(n16875),.clk(gclk));
	jand g16625(.dina(w_n16489_22[2]),.dinb(w_n16456_0[0]),.dout(n16876),.clk(gclk));
	jand g16626(.dina(w_n16460_0[0]),.dinb(w_asqrt63_26[0]),.dout(n16877),.clk(gclk));
	jand g16627(.dina(n16877),.dinb(w_n16485_0[1]),.dout(n16878),.clk(gclk));
	jnot g16628(.din(n16878),.dout(n16879),.clk(gclk));
	jor g16629(.dina(w_n16879_0[1]),.dinb(n16876),.dout(n16880),.clk(gclk));
	jnot g16630(.din(w_n16880_0[1]),.dout(n16881),.clk(gclk));
	jor g16631(.dina(n16881),.dinb(n16875),.dout(n16882),.clk(gclk));
	jor g16632(.dina(w_n16882_0[1]),.dinb(w_n16869_0[2]),.dout(asqrt_fa_13),.clk(gclk));
	jnot g16633(.din(w_a22_1[1]),.dout(n16885),.clk(gclk));
	jnot g16634(.din(w_a23_0[1]),.dout(n16886),.clk(gclk));
	jand g16635(.dina(w_n16886_0[1]),.dinb(w_n16885_1[1]),.dout(n16887),.clk(gclk));
	jand g16636(.dina(w_n16887_0[2]),.dinb(w_n16494_1[1]),.dout(n16888),.clk(gclk));
	jand g16637(.dina(w_asqrt12_33),.dinb(w_a24_0[1]),.dout(n16889),.clk(gclk));
	jor g16638(.dina(n16889),.dinb(w_n16888_0[1]),.dout(n16890),.clk(gclk));
	jand g16639(.dina(w_n16890_0[2]),.dinb(w_asqrt13_9[2]),.dout(n16891),.clk(gclk));
	jor g16640(.dina(w_n16890_0[1]),.dinb(w_asqrt13_9[1]),.dout(n16892),.clk(gclk));
	jand g16641(.dina(w_asqrt12_32[2]),.dinb(w_n16494_1[0]),.dout(n16893),.clk(gclk));
	jor g16642(.dina(n16893),.dinb(w_n16495_0[0]),.dout(n16894),.clk(gclk));
	jnot g16643(.din(w_n16496_0[1]),.dout(n16895),.clk(gclk));
	jnot g16644(.din(w_n16869_0[1]),.dout(n16896),.clk(gclk));
	jnot g16645(.din(w_n16861_0[0]),.dout(n16898),.clk(gclk));
	jnot g16646(.din(w_n16854_0[0]),.dout(n16899),.clk(gclk));
	jnot g16647(.din(w_n16846_0[0]),.dout(n16900),.clk(gclk));
	jnot g16648(.din(w_n16839_0[0]),.dout(n16901),.clk(gclk));
	jnot g16649(.din(w_n16831_0[0]),.dout(n16902),.clk(gclk));
	jnot g16650(.din(w_n16824_0[0]),.dout(n16903),.clk(gclk));
	jnot g16651(.din(w_n16817_0[0]),.dout(n16904),.clk(gclk));
	jnot g16652(.din(w_n16810_0[0]),.dout(n16905),.clk(gclk));
	jnot g16653(.din(w_n16802_0[0]),.dout(n16906),.clk(gclk));
	jnot g16654(.din(w_n16795_0[0]),.dout(n16907),.clk(gclk));
	jnot g16655(.din(w_n16787_0[0]),.dout(n16908),.clk(gclk));
	jnot g16656(.din(w_n16780_0[0]),.dout(n16909),.clk(gclk));
	jnot g16657(.din(w_n16772_0[0]),.dout(n16910),.clk(gclk));
	jnot g16658(.din(w_n16764_0[0]),.dout(n16911),.clk(gclk));
	jnot g16659(.din(w_n16757_0[0]),.dout(n16912),.clk(gclk));
	jnot g16660(.din(w_n16750_0[0]),.dout(n16913),.clk(gclk));
	jnot g16661(.din(w_n16742_0[0]),.dout(n16914),.clk(gclk));
	jnot g16662(.din(w_n16735_0[0]),.dout(n16915),.clk(gclk));
	jnot g16663(.din(w_n16727_0[0]),.dout(n16916),.clk(gclk));
	jnot g16664(.din(w_n16720_0[0]),.dout(n16917),.clk(gclk));
	jnot g16665(.din(w_n16713_0[0]),.dout(n16918),.clk(gclk));
	jnot g16666(.din(w_n16706_0[0]),.dout(n16919),.clk(gclk));
	jnot g16667(.din(w_n16698_0[0]),.dout(n16920),.clk(gclk));
	jnot g16668(.din(w_n16691_0[0]),.dout(n16921),.clk(gclk));
	jnot g16669(.din(w_n16683_0[0]),.dout(n16922),.clk(gclk));
	jnot g16670(.din(w_n16676_0[0]),.dout(n16923),.clk(gclk));
	jnot g16671(.din(w_n16669_0[0]),.dout(n16924),.clk(gclk));
	jnot g16672(.din(w_n16662_0[0]),.dout(n16925),.clk(gclk));
	jnot g16673(.din(w_n16654_0[0]),.dout(n16926),.clk(gclk));
	jnot g16674(.din(w_n16647_0[0]),.dout(n16927),.clk(gclk));
	jnot g16675(.din(w_n16639_0[0]),.dout(n16928),.clk(gclk));
	jnot g16676(.din(w_n16632_0[0]),.dout(n16929),.clk(gclk));
	jnot g16677(.din(w_n16624_0[0]),.dout(n16930),.clk(gclk));
	jnot g16678(.din(w_n16617_0[0]),.dout(n16931),.clk(gclk));
	jnot g16679(.din(w_n16609_0[0]),.dout(n16932),.clk(gclk));
	jnot g16680(.din(w_n16602_0[0]),.dout(n16933),.clk(gclk));
	jnot g16681(.din(w_n16595_0[0]),.dout(n16934),.clk(gclk));
	jnot g16682(.din(w_n16588_0[0]),.dout(n16935),.clk(gclk));
	jnot g16683(.din(w_n16580_0[0]),.dout(n16936),.clk(gclk));
	jnot g16684(.din(w_n16573_0[0]),.dout(n16937),.clk(gclk));
	jnot g16685(.din(w_n16565_0[0]),.dout(n16938),.clk(gclk));
	jnot g16686(.din(w_n16558_0[0]),.dout(n16939),.clk(gclk));
	jnot g16687(.din(w_n16550_0[0]),.dout(n16940),.clk(gclk));
	jnot g16688(.din(w_n16542_0[0]),.dout(n16941),.clk(gclk));
	jnot g16689(.din(w_n16535_0[0]),.dout(n16942),.clk(gclk));
	jnot g16690(.din(w_n16528_0[0]),.dout(n16943),.clk(gclk));
	jnot g16691(.din(w_n16520_0[0]),.dout(n16944),.clk(gclk));
	jnot g16692(.din(w_n16509_0[0]),.dout(n16945),.clk(gclk));
	jnot g16693(.din(w_n16501_0[0]),.dout(n16946),.clk(gclk));
	jand g16694(.dina(w_asqrt13_9[0]),.dinb(w_a26_0[2]),.dout(n16947),.clk(gclk));
	jor g16695(.dina(n16947),.dinb(w_n16497_0[0]),.dout(n16948),.clk(gclk));
	jor g16696(.dina(n16948),.dinb(w_asqrt14_17[0]),.dout(n16949),.clk(gclk));
	jand g16697(.dina(w_asqrt13_8[2]),.dinb(w_n15642_0[1]),.dout(n16950),.clk(gclk));
	jor g16698(.dina(n16950),.dinb(w_n15643_0[0]),.dout(n16951),.clk(gclk));
	jand g16699(.dina(w_n16512_0[0]),.dinb(n16951),.dout(n16952),.clk(gclk));
	jand g16700(.dina(w_n16952_0[1]),.dinb(n16949),.dout(n16953),.clk(gclk));
	jor g16701(.dina(n16953),.dinb(n16946),.dout(n16954),.clk(gclk));
	jor g16702(.dina(n16954),.dinb(w_asqrt15_9[2]),.dout(n16955),.clk(gclk));
	jnot g16703(.din(w_n16517_0[1]),.dout(n16956),.clk(gclk));
	jand g16704(.dina(n16956),.dinb(n16955),.dout(n16957),.clk(gclk));
	jor g16705(.dina(n16957),.dinb(n16945),.dout(n16958),.clk(gclk));
	jor g16706(.dina(n16958),.dinb(w_asqrt16_17[0]),.dout(n16959),.clk(gclk));
	jand g16707(.dina(w_n16524_0[1]),.dinb(n16959),.dout(n16960),.clk(gclk));
	jor g16708(.dina(n16960),.dinb(n16944),.dout(n16961),.clk(gclk));
	jor g16709(.dina(n16961),.dinb(w_asqrt17_10[0]),.dout(n16962),.clk(gclk));
	jnot g16710(.din(w_n16532_0[1]),.dout(n16963),.clk(gclk));
	jand g16711(.dina(n16963),.dinb(n16962),.dout(n16964),.clk(gclk));
	jor g16712(.dina(n16964),.dinb(n16943),.dout(n16965),.clk(gclk));
	jor g16713(.dina(n16965),.dinb(w_asqrt18_17[1]),.dout(n16966),.clk(gclk));
	jnot g16714(.din(w_n16539_0[1]),.dout(n16967),.clk(gclk));
	jand g16715(.dina(n16967),.dinb(n16966),.dout(n16968),.clk(gclk));
	jor g16716(.dina(n16968),.dinb(n16942),.dout(n16969),.clk(gclk));
	jor g16717(.dina(n16969),.dinb(w_asqrt19_10[1]),.dout(n16970),.clk(gclk));
	jand g16718(.dina(w_n16546_0[1]),.dinb(n16970),.dout(n16971),.clk(gclk));
	jor g16719(.dina(n16971),.dinb(n16941),.dout(n16972),.clk(gclk));
	jor g16720(.dina(n16972),.dinb(w_asqrt20_17[1]),.dout(n16973),.clk(gclk));
	jand g16721(.dina(w_n16554_0[1]),.dinb(n16973),.dout(n16974),.clk(gclk));
	jor g16722(.dina(n16974),.dinb(n16940),.dout(n16975),.clk(gclk));
	jor g16723(.dina(n16975),.dinb(w_asqrt21_11[0]),.dout(n16976),.clk(gclk));
	jnot g16724(.din(w_n16562_0[1]),.dout(n16977),.clk(gclk));
	jand g16725(.dina(n16977),.dinb(n16976),.dout(n16978),.clk(gclk));
	jor g16726(.dina(n16978),.dinb(n16939),.dout(n16979),.clk(gclk));
	jor g16727(.dina(n16979),.dinb(w_asqrt22_17[2]),.dout(n16980),.clk(gclk));
	jand g16728(.dina(w_n16569_0[1]),.dinb(n16980),.dout(n16981),.clk(gclk));
	jor g16729(.dina(n16981),.dinb(n16938),.dout(n16982),.clk(gclk));
	jor g16730(.dina(n16982),.dinb(w_asqrt23_11[2]),.dout(n16983),.clk(gclk));
	jnot g16731(.din(w_n16577_0[1]),.dout(n16984),.clk(gclk));
	jand g16732(.dina(n16984),.dinb(n16983),.dout(n16985),.clk(gclk));
	jor g16733(.dina(n16985),.dinb(n16937),.dout(n16986),.clk(gclk));
	jor g16734(.dina(n16986),.dinb(w_asqrt24_17[2]),.dout(n16987),.clk(gclk));
	jand g16735(.dina(w_n16584_0[1]),.dinb(n16987),.dout(n16988),.clk(gclk));
	jor g16736(.dina(n16988),.dinb(n16936),.dout(n16989),.clk(gclk));
	jor g16737(.dina(n16989),.dinb(w_asqrt25_11[2]),.dout(n16990),.clk(gclk));
	jnot g16738(.din(w_n16592_0[1]),.dout(n16991),.clk(gclk));
	jand g16739(.dina(n16991),.dinb(n16990),.dout(n16992),.clk(gclk));
	jor g16740(.dina(n16992),.dinb(n16935),.dout(n16993),.clk(gclk));
	jor g16741(.dina(n16993),.dinb(w_asqrt26_17[2]),.dout(n16994),.clk(gclk));
	jnot g16742(.din(w_n16599_0[1]),.dout(n16995),.clk(gclk));
	jand g16743(.dina(n16995),.dinb(n16994),.dout(n16996),.clk(gclk));
	jor g16744(.dina(n16996),.dinb(n16934),.dout(n16997),.clk(gclk));
	jor g16745(.dina(n16997),.dinb(w_asqrt27_12[1]),.dout(n16998),.clk(gclk));
	jnot g16746(.din(w_n16606_0[1]),.dout(n16999),.clk(gclk));
	jand g16747(.dina(n16999),.dinb(n16998),.dout(n17000),.clk(gclk));
	jor g16748(.dina(n17000),.dinb(n16933),.dout(n17001),.clk(gclk));
	jor g16749(.dina(n17001),.dinb(w_asqrt28_18[0]),.dout(n17002),.clk(gclk));
	jand g16750(.dina(w_n16613_0[1]),.dinb(n17002),.dout(n17003),.clk(gclk));
	jor g16751(.dina(n17003),.dinb(n16932),.dout(n17004),.clk(gclk));
	jor g16752(.dina(n17004),.dinb(w_asqrt29_12[2]),.dout(n17005),.clk(gclk));
	jnot g16753(.din(w_n16621_0[1]),.dout(n17006),.clk(gclk));
	jand g16754(.dina(n17006),.dinb(n17005),.dout(n17007),.clk(gclk));
	jor g16755(.dina(n17007),.dinb(n16931),.dout(n17008),.clk(gclk));
	jor g16756(.dina(n17008),.dinb(w_asqrt30_18[1]),.dout(n17009),.clk(gclk));
	jand g16757(.dina(w_n16628_0[1]),.dinb(n17009),.dout(n17010),.clk(gclk));
	jor g16758(.dina(n17010),.dinb(n16930),.dout(n17011),.clk(gclk));
	jor g16759(.dina(n17011),.dinb(w_asqrt31_13[1]),.dout(n17012),.clk(gclk));
	jnot g16760(.din(w_n16636_0[1]),.dout(n17013),.clk(gclk));
	jand g16761(.dina(n17013),.dinb(n17012),.dout(n17014),.clk(gclk));
	jor g16762(.dina(n17014),.dinb(n16929),.dout(n17015),.clk(gclk));
	jor g16763(.dina(n17015),.dinb(w_asqrt32_18[1]),.dout(n17016),.clk(gclk));
	jand g16764(.dina(w_n16643_0[1]),.dinb(n17016),.dout(n17017),.clk(gclk));
	jor g16765(.dina(n17017),.dinb(n16928),.dout(n17018),.clk(gclk));
	jor g16766(.dina(n17018),.dinb(w_asqrt33_14[0]),.dout(n17019),.clk(gclk));
	jnot g16767(.din(w_n16651_0[1]),.dout(n17020),.clk(gclk));
	jand g16768(.dina(n17020),.dinb(n17019),.dout(n17021),.clk(gclk));
	jor g16769(.dina(n17021),.dinb(n16927),.dout(n17022),.clk(gclk));
	jor g16770(.dina(n17022),.dinb(w_asqrt34_18[2]),.dout(n17023),.clk(gclk));
	jand g16771(.dina(w_n16658_0[1]),.dinb(n17023),.dout(n17024),.clk(gclk));
	jor g16772(.dina(n17024),.dinb(n16926),.dout(n17025),.clk(gclk));
	jor g16773(.dina(n17025),.dinb(w_asqrt35_14[2]),.dout(n17026),.clk(gclk));
	jnot g16774(.din(w_n16666_0[1]),.dout(n17027),.clk(gclk));
	jand g16775(.dina(n17027),.dinb(n17026),.dout(n17028),.clk(gclk));
	jor g16776(.dina(n17028),.dinb(n16925),.dout(n17029),.clk(gclk));
	jor g16777(.dina(n17029),.dinb(w_asqrt36_18[2]),.dout(n17030),.clk(gclk));
	jnot g16778(.din(w_n16673_0[1]),.dout(n17031),.clk(gclk));
	jand g16779(.dina(n17031),.dinb(n17030),.dout(n17032),.clk(gclk));
	jor g16780(.dina(n17032),.dinb(n16924),.dout(n17033),.clk(gclk));
	jor g16781(.dina(n17033),.dinb(w_asqrt37_15[0]),.dout(n17034),.clk(gclk));
	jnot g16782(.din(w_n16680_0[1]),.dout(n17035),.clk(gclk));
	jand g16783(.dina(n17035),.dinb(n17034),.dout(n17036),.clk(gclk));
	jor g16784(.dina(n17036),.dinb(n16923),.dout(n17037),.clk(gclk));
	jor g16785(.dina(n17037),.dinb(w_asqrt38_19[0]),.dout(n17038),.clk(gclk));
	jand g16786(.dina(w_n16687_0[1]),.dinb(n17038),.dout(n17039),.clk(gclk));
	jor g16787(.dina(n17039),.dinb(n16922),.dout(n17040),.clk(gclk));
	jor g16788(.dina(n17040),.dinb(w_asqrt39_15[2]),.dout(n17041),.clk(gclk));
	jnot g16789(.din(w_n16695_0[1]),.dout(n17042),.clk(gclk));
	jand g16790(.dina(n17042),.dinb(n17041),.dout(n17043),.clk(gclk));
	jor g16791(.dina(n17043),.dinb(n16921),.dout(n17044),.clk(gclk));
	jor g16792(.dina(n17044),.dinb(w_asqrt40_19[0]),.dout(n17045),.clk(gclk));
	jand g16793(.dina(w_n16702_0[1]),.dinb(n17045),.dout(n17046),.clk(gclk));
	jor g16794(.dina(n17046),.dinb(n16920),.dout(n17047),.clk(gclk));
	jor g16795(.dina(n17047),.dinb(w_asqrt41_16[0]),.dout(n17048),.clk(gclk));
	jnot g16796(.din(w_n16710_0[1]),.dout(n17049),.clk(gclk));
	jand g16797(.dina(n17049),.dinb(n17048),.dout(n17050),.clk(gclk));
	jor g16798(.dina(n17050),.dinb(n16919),.dout(n17051),.clk(gclk));
	jor g16799(.dina(n17051),.dinb(w_asqrt42_19[1]),.dout(n17052),.clk(gclk));
	jnot g16800(.din(w_n16717_0[1]),.dout(n17053),.clk(gclk));
	jand g16801(.dina(n17053),.dinb(n17052),.dout(n17054),.clk(gclk));
	jor g16802(.dina(n17054),.dinb(n16918),.dout(n17055),.clk(gclk));
	jor g16803(.dina(n17055),.dinb(w_asqrt43_16[1]),.dout(n17056),.clk(gclk));
	jnot g16804(.din(w_n16724_0[1]),.dout(n17057),.clk(gclk));
	jand g16805(.dina(n17057),.dinb(n17056),.dout(n17058),.clk(gclk));
	jor g16806(.dina(n17058),.dinb(n16917),.dout(n17059),.clk(gclk));
	jor g16807(.dina(n17059),.dinb(w_asqrt44_19[1]),.dout(n17060),.clk(gclk));
	jand g16808(.dina(w_n16731_0[1]),.dinb(n17060),.dout(n17061),.clk(gclk));
	jor g16809(.dina(n17061),.dinb(n16916),.dout(n17062),.clk(gclk));
	jor g16810(.dina(n17062),.dinb(w_asqrt45_17[0]),.dout(n17063),.clk(gclk));
	jnot g16811(.din(w_n16739_0[1]),.dout(n17064),.clk(gclk));
	jand g16812(.dina(n17064),.dinb(n17063),.dout(n17065),.clk(gclk));
	jor g16813(.dina(n17065),.dinb(n16915),.dout(n17066),.clk(gclk));
	jor g16814(.dina(n17066),.dinb(w_asqrt46_19[1]),.dout(n17067),.clk(gclk));
	jand g16815(.dina(w_n16746_0[1]),.dinb(n17067),.dout(n17068),.clk(gclk));
	jor g16816(.dina(n17068),.dinb(n16914),.dout(n17069),.clk(gclk));
	jor g16817(.dina(n17069),.dinb(w_asqrt47_17[2]),.dout(n17070),.clk(gclk));
	jnot g16818(.din(w_n16754_0[1]),.dout(n17071),.clk(gclk));
	jand g16819(.dina(n17071),.dinb(n17070),.dout(n17072),.clk(gclk));
	jor g16820(.dina(n17072),.dinb(n16913),.dout(n17073),.clk(gclk));
	jor g16821(.dina(n17073),.dinb(w_asqrt48_19[2]),.dout(n17074),.clk(gclk));
	jnot g16822(.din(w_n16761_0[1]),.dout(n17075),.clk(gclk));
	jand g16823(.dina(n17075),.dinb(n17074),.dout(n17076),.clk(gclk));
	jor g16824(.dina(n17076),.dinb(n16912),.dout(n17077),.clk(gclk));
	jor g16825(.dina(n17077),.dinb(w_asqrt49_18[0]),.dout(n17078),.clk(gclk));
	jand g16826(.dina(w_n16768_0[1]),.dinb(n17078),.dout(n17079),.clk(gclk));
	jor g16827(.dina(n17079),.dinb(n16911),.dout(n17080),.clk(gclk));
	jor g16828(.dina(n17080),.dinb(w_asqrt50_20[0]),.dout(n17081),.clk(gclk));
	jand g16829(.dina(n17081),.dinb(w_n16775_0[1]),.dout(n17082),.clk(gclk));
	jor g16830(.dina(n17082),.dinb(n16910),.dout(n17083),.clk(gclk));
	jor g16831(.dina(n17083),.dinb(w_asqrt51_18[1]),.dout(n17084),.clk(gclk));
	jnot g16832(.din(w_n16784_0[1]),.dout(n17085),.clk(gclk));
	jand g16833(.dina(n17085),.dinb(n17084),.dout(n17086),.clk(gclk));
	jor g16834(.dina(n17086),.dinb(n16909),.dout(n17087),.clk(gclk));
	jor g16835(.dina(n17087),.dinb(w_asqrt52_20[0]),.dout(n17088),.clk(gclk));
	jand g16836(.dina(w_n16791_0[1]),.dinb(n17088),.dout(n17089),.clk(gclk));
	jor g16837(.dina(n17089),.dinb(n16908),.dout(n17090),.clk(gclk));
	jor g16838(.dina(n17090),.dinb(w_asqrt53_19[0]),.dout(n17091),.clk(gclk));
	jnot g16839(.din(w_n16799_0[1]),.dout(n17092),.clk(gclk));
	jand g16840(.dina(n17092),.dinb(n17091),.dout(n17093),.clk(gclk));
	jor g16841(.dina(n17093),.dinb(n16907),.dout(n17094),.clk(gclk));
	jor g16842(.dina(n17094),.dinb(w_asqrt54_20[0]),.dout(n17095),.clk(gclk));
	jand g16843(.dina(w_n16806_0[1]),.dinb(n17095),.dout(n17096),.clk(gclk));
	jor g16844(.dina(n17096),.dinb(n16906),.dout(n17097),.clk(gclk));
	jor g16845(.dina(n17097),.dinb(w_asqrt55_19[1]),.dout(n17098),.clk(gclk));
	jnot g16846(.din(w_n16814_0[1]),.dout(n17099),.clk(gclk));
	jand g16847(.dina(n17099),.dinb(n17098),.dout(n17100),.clk(gclk));
	jor g16848(.dina(n17100),.dinb(n16905),.dout(n17101),.clk(gclk));
	jor g16849(.dina(n17101),.dinb(w_asqrt56_20[1]),.dout(n17102),.clk(gclk));
	jnot g16850(.din(w_n16821_0[1]),.dout(n17103),.clk(gclk));
	jand g16851(.dina(n17103),.dinb(n17102),.dout(n17104),.clk(gclk));
	jor g16852(.dina(n17104),.dinb(n16904),.dout(n17105),.clk(gclk));
	jor g16853(.dina(n17105),.dinb(w_asqrt57_20[0]),.dout(n17106),.clk(gclk));
	jnot g16854(.din(w_n16828_0[1]),.dout(n17107),.clk(gclk));
	jand g16855(.dina(n17107),.dinb(n17106),.dout(n17108),.clk(gclk));
	jor g16856(.dina(n17108),.dinb(n16903),.dout(n17109),.clk(gclk));
	jor g16857(.dina(n17109),.dinb(w_asqrt58_20[2]),.dout(n17110),.clk(gclk));
	jand g16858(.dina(w_n16835_0[1]),.dinb(n17110),.dout(n17111),.clk(gclk));
	jor g16859(.dina(n17111),.dinb(n16902),.dout(n17112),.clk(gclk));
	jor g16860(.dina(n17112),.dinb(w_asqrt59_20[1]),.dout(n17113),.clk(gclk));
	jnot g16861(.din(w_n16843_0[1]),.dout(n17114),.clk(gclk));
	jand g16862(.dina(n17114),.dinb(n17113),.dout(n17115),.clk(gclk));
	jor g16863(.dina(n17115),.dinb(n16901),.dout(n17116),.clk(gclk));
	jor g16864(.dina(n17116),.dinb(w_asqrt60_20[2]),.dout(n17117),.clk(gclk));
	jand g16865(.dina(w_n16850_0[1]),.dinb(n17117),.dout(n17118),.clk(gclk));
	jor g16866(.dina(n17118),.dinb(n16900),.dout(n17119),.clk(gclk));
	jor g16867(.dina(n17119),.dinb(w_asqrt61_20[2]),.dout(n17120),.clk(gclk));
	jnot g16868(.din(w_n16858_0[1]),.dout(n17121),.clk(gclk));
	jand g16869(.dina(n17121),.dinb(n17120),.dout(n17122),.clk(gclk));
	jor g16870(.dina(n17122),.dinb(n16899),.dout(n17123),.clk(gclk));
	jor g16871(.dina(n17123),.dinb(w_asqrt62_20[2]),.dout(n17124),.clk(gclk));
	jand g16872(.dina(w_n16865_0[0]),.dinb(n17124),.dout(n17125),.clk(gclk));
	jor g16873(.dina(n17125),.dinb(n16898),.dout(n17126),.clk(gclk));
	jand g16874(.dina(n17126),.dinb(w_n16492_0[0]),.dout(n17127),.clk(gclk));
	jnot g16875(.din(w_n16872_0[0]),.dout(n17128),.clk(gclk));
	jand g16876(.dina(n17128),.dinb(w_n17127_0[1]),.dout(n17129),.clk(gclk));
	jand g16877(.dina(n17129),.dinb(w_n16485_0[0]),.dout(n17130),.clk(gclk));
	jor g16878(.dina(n17130),.dinb(w_asqrt63_25[2]),.dout(n17131),.clk(gclk));
	jand g16879(.dina(w_n16880_0[0]),.dinb(w_n17131_0[1]),.dout(n17132),.clk(gclk));
	jand g16880(.dina(w_n17132_0[1]),.dinb(w_n16896_1[1]),.dout(n17134),.clk(gclk));
	jor g16881(.dina(w_n17134_15[1]),.dinb(n16895),.dout(n17135),.clk(gclk));
	jand g16882(.dina(n17135),.dinb(n16894),.dout(n17136),.clk(gclk));
	jand g16883(.dina(n17136),.dinb(n16892),.dout(n17137),.clk(gclk));
	jor g16884(.dina(n17137),.dinb(w_n16891_0[1]),.dout(n17138),.clk(gclk));
	jand g16885(.dina(w_n17138_0[2]),.dinb(w_asqrt14_16[2]),.dout(n17139),.clk(gclk));
	jor g16886(.dina(w_n17138_0[1]),.dinb(w_asqrt14_16[1]),.dout(n17140),.clk(gclk));
	jand g16887(.dina(w_asqrt12_32[1]),.dinb(w_n16496_0[0]),.dout(n17141),.clk(gclk));
	jand g16888(.dina(w_n16896_1[0]),.dinb(w_asqrt13_8[1]),.dout(n17142),.clk(gclk));
	jand g16889(.dina(n17142),.dinb(w_n17131_0[0]),.dout(n17143),.clk(gclk));
	jand g16890(.dina(n17143),.dinb(w_n16879_0[0]),.dout(n17144),.clk(gclk));
	jor g16891(.dina(n17144),.dinb(w_n17141_0[1]),.dout(n17145),.clk(gclk));
	jxor g16892(.dina(n17145),.dinb(w_a26_0[1]),.dout(n17146),.clk(gclk));
	jnot g16893(.din(w_n17146_0[1]),.dout(n17147),.clk(gclk));
	jand g16894(.dina(w_n17147_0[1]),.dinb(n17140),.dout(n17148),.clk(gclk));
	jor g16895(.dina(n17148),.dinb(w_n17139_0[1]),.dout(n17149),.clk(gclk));
	jand g16896(.dina(w_n17149_0[2]),.dinb(w_asqrt15_9[1]),.dout(n17150),.clk(gclk));
	jor g16897(.dina(w_n17149_0[1]),.dinb(w_asqrt15_9[0]),.dout(n17151),.clk(gclk));
	jxor g16898(.dina(w_n16500_0[0]),.dinb(w_n15878_15[2]),.dout(n17152),.clk(gclk));
	jand g16899(.dina(n17152),.dinb(w_asqrt12_32[0]),.dout(n17153),.clk(gclk));
	jxor g16900(.dina(n17153),.dinb(w_n16952_0[0]),.dout(n17154),.clk(gclk));
	jand g16901(.dina(w_n17154_0[1]),.dinb(n17151),.dout(n17155),.clk(gclk));
	jor g16902(.dina(n17155),.dinb(w_n17150_0[1]),.dout(n17156),.clk(gclk));
	jand g16903(.dina(w_n17156_0[2]),.dinb(w_asqrt16_16[2]),.dout(n17157),.clk(gclk));
	jor g16904(.dina(w_n17156_0[1]),.dinb(w_asqrt16_16[1]),.dout(n17158),.clk(gclk));
	jxor g16905(.dina(w_n16508_0[0]),.dinb(w_n15260_23[1]),.dout(n17159),.clk(gclk));
	jand g16906(.dina(n17159),.dinb(w_asqrt12_31[2]),.dout(n17160),.clk(gclk));
	jxor g16907(.dina(n17160),.dinb(w_n16517_0[0]),.dout(n17161),.clk(gclk));
	jnot g16908(.din(w_n17161_0[1]),.dout(n17162),.clk(gclk));
	jand g16909(.dina(w_n17162_0[1]),.dinb(n17158),.dout(n17163),.clk(gclk));
	jor g16910(.dina(n17163),.dinb(w_n17157_0[1]),.dout(n17164),.clk(gclk));
	jand g16911(.dina(w_n17164_0[2]),.dinb(w_asqrt17_9[2]),.dout(n17165),.clk(gclk));
	jor g16912(.dina(w_n17164_0[1]),.dinb(w_asqrt17_9[1]),.dout(n17166),.clk(gclk));
	jxor g16913(.dina(w_n16519_0[0]),.dinb(w_n14674_16[1]),.dout(n17167),.clk(gclk));
	jand g16914(.dina(n17167),.dinb(w_asqrt12_31[1]),.dout(n17168),.clk(gclk));
	jxor g16915(.dina(n17168),.dinb(w_n16524_0[0]),.dout(n17169),.clk(gclk));
	jand g16916(.dina(w_n17169_0[1]),.dinb(n17166),.dout(n17170),.clk(gclk));
	jor g16917(.dina(n17170),.dinb(w_n17165_0[1]),.dout(n17171),.clk(gclk));
	jand g16918(.dina(w_n17171_0[2]),.dinb(w_asqrt18_17[0]),.dout(n17172),.clk(gclk));
	jor g16919(.dina(w_n17171_0[1]),.dinb(w_asqrt18_16[2]),.dout(n17173),.clk(gclk));
	jxor g16920(.dina(w_n16527_0[0]),.dinb(w_n14078_23[2]),.dout(n17174),.clk(gclk));
	jand g16921(.dina(n17174),.dinb(w_asqrt12_31[0]),.dout(n17175),.clk(gclk));
	jxor g16922(.dina(n17175),.dinb(w_n16532_0[0]),.dout(n17176),.clk(gclk));
	jnot g16923(.din(w_n17176_0[1]),.dout(n17177),.clk(gclk));
	jand g16924(.dina(w_n17177_0[1]),.dinb(n17173),.dout(n17178),.clk(gclk));
	jor g16925(.dina(n17178),.dinb(w_n17172_0[1]),.dout(n17179),.clk(gclk));
	jand g16926(.dina(w_n17179_0[2]),.dinb(w_asqrt19_10[0]),.dout(n17180),.clk(gclk));
	jor g16927(.dina(w_n17179_0[1]),.dinb(w_asqrt19_9[2]),.dout(n17181),.clk(gclk));
	jxor g16928(.dina(w_n16534_0[0]),.dinb(w_n13515_17[1]),.dout(n17182),.clk(gclk));
	jand g16929(.dina(n17182),.dinb(w_asqrt12_30[2]),.dout(n17183),.clk(gclk));
	jxor g16930(.dina(n17183),.dinb(w_n16539_0[0]),.dout(n17184),.clk(gclk));
	jnot g16931(.din(w_n17184_0[1]),.dout(n17185),.clk(gclk));
	jand g16932(.dina(w_n17185_0[1]),.dinb(n17181),.dout(n17186),.clk(gclk));
	jor g16933(.dina(n17186),.dinb(w_n17180_0[1]),.dout(n17187),.clk(gclk));
	jand g16934(.dina(w_n17187_0[2]),.dinb(w_asqrt20_17[0]),.dout(n17188),.clk(gclk));
	jor g16935(.dina(w_n17187_0[1]),.dinb(w_asqrt20_16[2]),.dout(n17189),.clk(gclk));
	jxor g16936(.dina(w_n16541_0[0]),.dinb(w_n12947_24[1]),.dout(n17190),.clk(gclk));
	jand g16937(.dina(n17190),.dinb(w_asqrt12_30[1]),.dout(n17191),.clk(gclk));
	jxor g16938(.dina(n17191),.dinb(w_n16546_0[0]),.dout(n17192),.clk(gclk));
	jand g16939(.dina(w_n17192_0[1]),.dinb(n17189),.dout(n17193),.clk(gclk));
	jor g16940(.dina(n17193),.dinb(w_n17188_0[1]),.dout(n17194),.clk(gclk));
	jand g16941(.dina(w_n17194_0[2]),.dinb(w_asqrt21_10[2]),.dout(n17195),.clk(gclk));
	jor g16942(.dina(w_n17194_0[1]),.dinb(w_asqrt21_10[1]),.dout(n17196),.clk(gclk));
	jxor g16943(.dina(w_n16549_0[0]),.dinb(w_n12410_18[0]),.dout(n17197),.clk(gclk));
	jand g16944(.dina(n17197),.dinb(w_asqrt12_30[0]),.dout(n17198),.clk(gclk));
	jxor g16945(.dina(n17198),.dinb(w_n16554_0[0]),.dout(n17199),.clk(gclk));
	jand g16946(.dina(w_n17199_0[1]),.dinb(n17196),.dout(n17200),.clk(gclk));
	jor g16947(.dina(n17200),.dinb(w_n17195_0[1]),.dout(n17201),.clk(gclk));
	jand g16948(.dina(w_n17201_0[2]),.dinb(w_asqrt22_17[1]),.dout(n17202),.clk(gclk));
	jor g16949(.dina(w_n17201_0[1]),.dinb(w_asqrt22_17[0]),.dout(n17203),.clk(gclk));
	jxor g16950(.dina(w_n16557_0[0]),.dinb(w_n11858_24[2]),.dout(n17204),.clk(gclk));
	jand g16951(.dina(n17204),.dinb(w_asqrt12_29[2]),.dout(n17205),.clk(gclk));
	jxor g16952(.dina(n17205),.dinb(w_n16562_0[0]),.dout(n17206),.clk(gclk));
	jnot g16953(.din(w_n17206_0[1]),.dout(n17207),.clk(gclk));
	jand g16954(.dina(w_n17207_0[1]),.dinb(n17203),.dout(n17208),.clk(gclk));
	jor g16955(.dina(n17208),.dinb(w_n17202_0[1]),.dout(n17209),.clk(gclk));
	jand g16956(.dina(w_n17209_0[2]),.dinb(w_asqrt23_11[1]),.dout(n17210),.clk(gclk));
	jor g16957(.dina(w_n17209_0[1]),.dinb(w_asqrt23_11[0]),.dout(n17211),.clk(gclk));
	jxor g16958(.dina(w_n16564_0[0]),.dinb(w_n11347_18[2]),.dout(n17212),.clk(gclk));
	jand g16959(.dina(n17212),.dinb(w_asqrt12_29[1]),.dout(n17213),.clk(gclk));
	jxor g16960(.dina(n17213),.dinb(w_n16569_0[0]),.dout(n17214),.clk(gclk));
	jand g16961(.dina(w_n17214_0[1]),.dinb(n17211),.dout(n17215),.clk(gclk));
	jor g16962(.dina(n17215),.dinb(w_n17210_0[1]),.dout(n17216),.clk(gclk));
	jand g16963(.dina(w_n17216_0[2]),.dinb(w_asqrt24_17[1]),.dout(n17217),.clk(gclk));
	jor g16964(.dina(w_n17216_0[1]),.dinb(w_asqrt24_17[0]),.dout(n17218),.clk(gclk));
	jxor g16965(.dina(w_n16572_0[0]),.dinb(w_n10824_25[1]),.dout(n17219),.clk(gclk));
	jand g16966(.dina(n17219),.dinb(w_asqrt12_29[0]),.dout(n17220),.clk(gclk));
	jxor g16967(.dina(n17220),.dinb(w_n16577_0[0]),.dout(n17221),.clk(gclk));
	jnot g16968(.din(w_n17221_0[1]),.dout(n17222),.clk(gclk));
	jand g16969(.dina(w_n17222_0[1]),.dinb(n17218),.dout(n17223),.clk(gclk));
	jor g16970(.dina(n17223),.dinb(w_n17217_0[1]),.dout(n17224),.clk(gclk));
	jand g16971(.dina(w_n17224_0[2]),.dinb(w_asqrt25_11[1]),.dout(n17225),.clk(gclk));
	jor g16972(.dina(w_n17224_0[1]),.dinb(w_asqrt25_11[0]),.dout(n17226),.clk(gclk));
	jxor g16973(.dina(w_n16579_0[0]),.dinb(w_n10328_19[2]),.dout(n17227),.clk(gclk));
	jand g16974(.dina(n17227),.dinb(w_asqrt12_28[2]),.dout(n17228),.clk(gclk));
	jxor g16975(.dina(n17228),.dinb(w_n16584_0[0]),.dout(n17229),.clk(gclk));
	jand g16976(.dina(w_n17229_0[1]),.dinb(n17226),.dout(n17230),.clk(gclk));
	jor g16977(.dina(n17230),.dinb(w_n17225_0[1]),.dout(n17231),.clk(gclk));
	jand g16978(.dina(w_n17231_0[2]),.dinb(w_asqrt26_17[1]),.dout(n17232),.clk(gclk));
	jor g16979(.dina(w_n17231_0[1]),.dinb(w_asqrt26_17[0]),.dout(n17233),.clk(gclk));
	jxor g16980(.dina(w_n16587_0[0]),.dinb(w_n9832_26[0]),.dout(n17234),.clk(gclk));
	jand g16981(.dina(n17234),.dinb(w_asqrt12_28[1]),.dout(n17235),.clk(gclk));
	jxor g16982(.dina(n17235),.dinb(w_n16592_0[0]),.dout(n17236),.clk(gclk));
	jnot g16983(.din(w_n17236_0[1]),.dout(n17237),.clk(gclk));
	jand g16984(.dina(w_n17237_0[1]),.dinb(n17233),.dout(n17238),.clk(gclk));
	jor g16985(.dina(n17238),.dinb(w_n17232_0[1]),.dout(n17239),.clk(gclk));
	jand g16986(.dina(w_n17239_0[2]),.dinb(w_asqrt27_12[0]),.dout(n17240),.clk(gclk));
	jor g16987(.dina(w_n17239_0[1]),.dinb(w_asqrt27_11[2]),.dout(n17241),.clk(gclk));
	jxor g16988(.dina(w_n16594_0[0]),.dinb(w_n9369_20[2]),.dout(n17242),.clk(gclk));
	jand g16989(.dina(n17242),.dinb(w_asqrt12_28[0]),.dout(n17243),.clk(gclk));
	jxor g16990(.dina(n17243),.dinb(w_n16599_0[0]),.dout(n17244),.clk(gclk));
	jnot g16991(.din(w_n17244_0[1]),.dout(n17245),.clk(gclk));
	jand g16992(.dina(w_n17245_0[1]),.dinb(n17241),.dout(n17246),.clk(gclk));
	jor g16993(.dina(n17246),.dinb(w_n17240_0[1]),.dout(n17247),.clk(gclk));
	jand g16994(.dina(w_n17247_0[2]),.dinb(w_asqrt28_17[2]),.dout(n17248),.clk(gclk));
	jor g16995(.dina(w_n17247_0[1]),.dinb(w_asqrt28_17[1]),.dout(n17249),.clk(gclk));
	jxor g16996(.dina(w_n16601_0[0]),.dinb(w_n8890_26[1]),.dout(n17250),.clk(gclk));
	jand g16997(.dina(n17250),.dinb(w_asqrt12_27[2]),.dout(n17251),.clk(gclk));
	jxor g16998(.dina(n17251),.dinb(w_n16606_0[0]),.dout(n17252),.clk(gclk));
	jnot g16999(.din(w_n17252_0[1]),.dout(n17253),.clk(gclk));
	jand g17000(.dina(w_n17253_0[1]),.dinb(n17249),.dout(n17254),.clk(gclk));
	jor g17001(.dina(n17254),.dinb(w_n17248_0[1]),.dout(n17255),.clk(gclk));
	jand g17002(.dina(w_n17255_0[2]),.dinb(w_asqrt29_12[1]),.dout(n17256),.clk(gclk));
	jor g17003(.dina(w_n17255_0[1]),.dinb(w_asqrt29_12[0]),.dout(n17257),.clk(gclk));
	jxor g17004(.dina(w_n16608_0[0]),.dinb(w_n8449_21[1]),.dout(n17258),.clk(gclk));
	jand g17005(.dina(n17258),.dinb(w_asqrt12_27[1]),.dout(n17259),.clk(gclk));
	jxor g17006(.dina(n17259),.dinb(w_n16613_0[0]),.dout(n17260),.clk(gclk));
	jand g17007(.dina(w_n17260_0[1]),.dinb(n17257),.dout(n17261),.clk(gclk));
	jor g17008(.dina(n17261),.dinb(w_n17256_0[1]),.dout(n17262),.clk(gclk));
	jand g17009(.dina(w_n17262_0[2]),.dinb(w_asqrt30_18[0]),.dout(n17263),.clk(gclk));
	jor g17010(.dina(w_n17262_0[1]),.dinb(w_asqrt30_17[2]),.dout(n17264),.clk(gclk));
	jxor g17011(.dina(w_n16616_0[0]),.dinb(w_n8003_27[0]),.dout(n17265),.clk(gclk));
	jand g17012(.dina(n17265),.dinb(w_asqrt12_27[0]),.dout(n17266),.clk(gclk));
	jxor g17013(.dina(n17266),.dinb(w_n16621_0[0]),.dout(n17267),.clk(gclk));
	jnot g17014(.din(w_n17267_0[1]),.dout(n17268),.clk(gclk));
	jand g17015(.dina(w_n17268_0[1]),.dinb(n17264),.dout(n17269),.clk(gclk));
	jor g17016(.dina(n17269),.dinb(w_n17263_0[1]),.dout(n17270),.clk(gclk));
	jand g17017(.dina(w_n17270_0[2]),.dinb(w_asqrt31_13[0]),.dout(n17271),.clk(gclk));
	jor g17018(.dina(w_n17270_0[1]),.dinb(w_asqrt31_12[2]),.dout(n17272),.clk(gclk));
	jxor g17019(.dina(w_n16623_0[0]),.dinb(w_n7581_22[1]),.dout(n17273),.clk(gclk));
	jand g17020(.dina(n17273),.dinb(w_asqrt12_26[2]),.dout(n17274),.clk(gclk));
	jxor g17021(.dina(n17274),.dinb(w_n16628_0[0]),.dout(n17275),.clk(gclk));
	jand g17022(.dina(w_n17275_0[1]),.dinb(n17272),.dout(n17276),.clk(gclk));
	jor g17023(.dina(n17276),.dinb(w_n17271_0[1]),.dout(n17277),.clk(gclk));
	jand g17024(.dina(w_n17277_0[2]),.dinb(w_asqrt32_18[0]),.dout(n17278),.clk(gclk));
	jor g17025(.dina(w_n17277_0[1]),.dinb(w_asqrt32_17[2]),.dout(n17279),.clk(gclk));
	jxor g17026(.dina(w_n16631_0[0]),.dinb(w_n7154_27[1]),.dout(n17280),.clk(gclk));
	jand g17027(.dina(n17280),.dinb(w_asqrt12_26[1]),.dout(n17281),.clk(gclk));
	jxor g17028(.dina(n17281),.dinb(w_n16636_0[0]),.dout(n17282),.clk(gclk));
	jnot g17029(.din(w_n17282_0[1]),.dout(n17283),.clk(gclk));
	jand g17030(.dina(w_n17283_0[1]),.dinb(n17279),.dout(n17284),.clk(gclk));
	jor g17031(.dina(n17284),.dinb(w_n17278_0[1]),.dout(n17285),.clk(gclk));
	jand g17032(.dina(w_n17285_0[2]),.dinb(w_asqrt33_13[2]),.dout(n17286),.clk(gclk));
	jor g17033(.dina(w_n17285_0[1]),.dinb(w_asqrt33_13[1]),.dout(n17287),.clk(gclk));
	jxor g17034(.dina(w_n16638_0[0]),.dinb(w_n6758_23[0]),.dout(n17288),.clk(gclk));
	jand g17035(.dina(n17288),.dinb(w_asqrt12_26[0]),.dout(n17289),.clk(gclk));
	jxor g17036(.dina(n17289),.dinb(w_n16643_0[0]),.dout(n17290),.clk(gclk));
	jand g17037(.dina(w_n17290_0[1]),.dinb(n17287),.dout(n17291),.clk(gclk));
	jor g17038(.dina(n17291),.dinb(w_n17286_0[1]),.dout(n17292),.clk(gclk));
	jand g17039(.dina(w_n17292_0[2]),.dinb(w_asqrt34_18[1]),.dout(n17293),.clk(gclk));
	jor g17040(.dina(w_n17292_0[1]),.dinb(w_asqrt34_18[0]),.dout(n17294),.clk(gclk));
	jxor g17041(.dina(w_n16646_0[0]),.dinb(w_n6357_27[2]),.dout(n17295),.clk(gclk));
	jand g17042(.dina(n17295),.dinb(w_asqrt12_25[2]),.dout(n17296),.clk(gclk));
	jxor g17043(.dina(n17296),.dinb(w_n16651_0[0]),.dout(n17297),.clk(gclk));
	jnot g17044(.din(w_n17297_0[1]),.dout(n17298),.clk(gclk));
	jand g17045(.dina(w_n17298_0[1]),.dinb(n17294),.dout(n17299),.clk(gclk));
	jor g17046(.dina(n17299),.dinb(w_n17293_0[1]),.dout(n17300),.clk(gclk));
	jand g17047(.dina(w_n17300_0[2]),.dinb(w_asqrt35_14[1]),.dout(n17301),.clk(gclk));
	jor g17048(.dina(w_n17300_0[1]),.dinb(w_asqrt35_14[0]),.dout(n17302),.clk(gclk));
	jxor g17049(.dina(w_n16653_0[0]),.dinb(w_n5989_23[2]),.dout(n17303),.clk(gclk));
	jand g17050(.dina(n17303),.dinb(w_asqrt12_25[1]),.dout(n17304),.clk(gclk));
	jxor g17051(.dina(n17304),.dinb(w_n16658_0[0]),.dout(n17305),.clk(gclk));
	jand g17052(.dina(w_n17305_0[1]),.dinb(n17302),.dout(n17306),.clk(gclk));
	jor g17053(.dina(n17306),.dinb(w_n17301_0[1]),.dout(n17307),.clk(gclk));
	jand g17054(.dina(w_n17307_0[2]),.dinb(w_asqrt36_18[1]),.dout(n17308),.clk(gclk));
	jor g17055(.dina(w_n17307_0[1]),.dinb(w_asqrt36_18[0]),.dout(n17309),.clk(gclk));
	jxor g17056(.dina(w_n16661_0[0]),.dinb(w_n5606_28[0]),.dout(n17310),.clk(gclk));
	jand g17057(.dina(n17310),.dinb(w_asqrt12_25[0]),.dout(n17311),.clk(gclk));
	jxor g17058(.dina(n17311),.dinb(w_n16666_0[0]),.dout(n17312),.clk(gclk));
	jnot g17059(.din(w_n17312_0[1]),.dout(n17313),.clk(gclk));
	jand g17060(.dina(w_n17313_0[1]),.dinb(n17309),.dout(n17314),.clk(gclk));
	jor g17061(.dina(n17314),.dinb(w_n17308_0[1]),.dout(n17315),.clk(gclk));
	jand g17062(.dina(w_n17315_0[2]),.dinb(w_asqrt37_14[2]),.dout(n17316),.clk(gclk));
	jor g17063(.dina(w_n17315_0[1]),.dinb(w_asqrt37_14[1]),.dout(n17317),.clk(gclk));
	jxor g17064(.dina(w_n16668_0[0]),.dinb(w_n5259_24[2]),.dout(n17318),.clk(gclk));
	jand g17065(.dina(n17318),.dinb(w_asqrt12_24[2]),.dout(n17319),.clk(gclk));
	jxor g17066(.dina(n17319),.dinb(w_n16673_0[0]),.dout(n17320),.clk(gclk));
	jnot g17067(.din(w_n17320_0[1]),.dout(n17321),.clk(gclk));
	jand g17068(.dina(w_n17321_0[1]),.dinb(n17317),.dout(n17322),.clk(gclk));
	jor g17069(.dina(n17322),.dinb(w_n17316_0[1]),.dout(n17323),.clk(gclk));
	jand g17070(.dina(w_n17323_0[2]),.dinb(w_asqrt38_18[2]),.dout(n17324),.clk(gclk));
	jor g17071(.dina(w_n17323_0[1]),.dinb(w_asqrt38_18[1]),.dout(n17325),.clk(gclk));
	jxor g17072(.dina(w_n16675_0[0]),.dinb(w_n4902_28[2]),.dout(n17326),.clk(gclk));
	jand g17073(.dina(n17326),.dinb(w_asqrt12_24[1]),.dout(n17327),.clk(gclk));
	jxor g17074(.dina(n17327),.dinb(w_n16680_0[0]),.dout(n17328),.clk(gclk));
	jnot g17075(.din(w_n17328_0[1]),.dout(n17329),.clk(gclk));
	jand g17076(.dina(w_n17329_0[1]),.dinb(n17325),.dout(n17330),.clk(gclk));
	jor g17077(.dina(n17330),.dinb(w_n17324_0[1]),.dout(n17331),.clk(gclk));
	jand g17078(.dina(w_n17331_0[2]),.dinb(w_asqrt39_15[1]),.dout(n17332),.clk(gclk));
	jor g17079(.dina(w_n17331_0[1]),.dinb(w_asqrt39_15[0]),.dout(n17333),.clk(gclk));
	jxor g17080(.dina(w_n16682_0[0]),.dinb(w_n4582_25[2]),.dout(n17334),.clk(gclk));
	jand g17081(.dina(n17334),.dinb(w_asqrt12_24[0]),.dout(n17335),.clk(gclk));
	jxor g17082(.dina(n17335),.dinb(w_n16687_0[0]),.dout(n17336),.clk(gclk));
	jand g17083(.dina(w_n17336_0[1]),.dinb(n17333),.dout(n17337),.clk(gclk));
	jor g17084(.dina(n17337),.dinb(w_n17332_0[1]),.dout(n17338),.clk(gclk));
	jand g17085(.dina(w_n17338_0[2]),.dinb(w_asqrt40_18[2]),.dout(n17339),.clk(gclk));
	jor g17086(.dina(w_n17338_0[1]),.dinb(w_asqrt40_18[1]),.dout(n17340),.clk(gclk));
	jxor g17087(.dina(w_n16690_0[0]),.dinb(w_n4249_29[1]),.dout(n17341),.clk(gclk));
	jand g17088(.dina(n17341),.dinb(w_asqrt12_23[2]),.dout(n17342),.clk(gclk));
	jxor g17089(.dina(n17342),.dinb(w_n16695_0[0]),.dout(n17343),.clk(gclk));
	jnot g17090(.din(w_n17343_0[1]),.dout(n17344),.clk(gclk));
	jand g17091(.dina(w_n17344_0[1]),.dinb(n17340),.dout(n17345),.clk(gclk));
	jor g17092(.dina(n17345),.dinb(w_n17339_0[1]),.dout(n17346),.clk(gclk));
	jand g17093(.dina(w_n17346_0[2]),.dinb(w_asqrt41_15[2]),.dout(n17347),.clk(gclk));
	jor g17094(.dina(w_n17346_0[1]),.dinb(w_asqrt41_15[1]),.dout(n17348),.clk(gclk));
	jxor g17095(.dina(w_n16697_0[0]),.dinb(w_n3955_26[1]),.dout(n17349),.clk(gclk));
	jand g17096(.dina(n17349),.dinb(w_asqrt12_23[1]),.dout(n17350),.clk(gclk));
	jxor g17097(.dina(n17350),.dinb(w_n16702_0[0]),.dout(n17351),.clk(gclk));
	jand g17098(.dina(w_n17351_0[1]),.dinb(n17348),.dout(n17352),.clk(gclk));
	jor g17099(.dina(n17352),.dinb(w_n17347_0[1]),.dout(n17353),.clk(gclk));
	jand g17100(.dina(w_n17353_0[2]),.dinb(w_asqrt42_19[0]),.dout(n17354),.clk(gclk));
	jor g17101(.dina(w_n17353_0[1]),.dinb(w_asqrt42_18[2]),.dout(n17355),.clk(gclk));
	jxor g17102(.dina(w_n16705_0[0]),.dinb(w_n3642_29[2]),.dout(n17356),.clk(gclk));
	jand g17103(.dina(n17356),.dinb(w_asqrt12_23[0]),.dout(n17357),.clk(gclk));
	jxor g17104(.dina(n17357),.dinb(w_n16710_0[0]),.dout(n17358),.clk(gclk));
	jnot g17105(.din(w_n17358_0[1]),.dout(n17359),.clk(gclk));
	jand g17106(.dina(w_n17359_0[1]),.dinb(n17355),.dout(n17360),.clk(gclk));
	jor g17107(.dina(n17360),.dinb(w_n17354_0[1]),.dout(n17361),.clk(gclk));
	jand g17108(.dina(w_n17361_0[2]),.dinb(w_asqrt43_16[0]),.dout(n17362),.clk(gclk));
	jor g17109(.dina(w_n17361_0[1]),.dinb(w_asqrt43_15[2]),.dout(n17363),.clk(gclk));
	jxor g17110(.dina(w_n16712_0[0]),.dinb(w_n3368_27[0]),.dout(n17364),.clk(gclk));
	jand g17111(.dina(n17364),.dinb(w_asqrt12_22[2]),.dout(n17365),.clk(gclk));
	jxor g17112(.dina(n17365),.dinb(w_n16717_0[0]),.dout(n17366),.clk(gclk));
	jnot g17113(.din(w_n17366_0[1]),.dout(n17367),.clk(gclk));
	jand g17114(.dina(w_n17367_0[1]),.dinb(n17363),.dout(n17368),.clk(gclk));
	jor g17115(.dina(n17368),.dinb(w_n17362_0[1]),.dout(n17369),.clk(gclk));
	jand g17116(.dina(w_n17369_0[2]),.dinb(w_asqrt44_19[0]),.dout(n17370),.clk(gclk));
	jor g17117(.dina(w_n17369_0[1]),.dinb(w_asqrt44_18[2]),.dout(n17371),.clk(gclk));
	jxor g17118(.dina(w_n16719_0[0]),.dinb(w_n3089_30[1]),.dout(n17372),.clk(gclk));
	jand g17119(.dina(n17372),.dinb(w_asqrt12_22[1]),.dout(n17373),.clk(gclk));
	jxor g17120(.dina(n17373),.dinb(w_n16724_0[0]),.dout(n17374),.clk(gclk));
	jnot g17121(.din(w_n17374_0[1]),.dout(n17375),.clk(gclk));
	jand g17122(.dina(w_n17375_0[1]),.dinb(n17371),.dout(n17376),.clk(gclk));
	jor g17123(.dina(n17376),.dinb(w_n17370_0[1]),.dout(n17377),.clk(gclk));
	jand g17124(.dina(w_n17377_0[2]),.dinb(w_asqrt45_16[2]),.dout(n17378),.clk(gclk));
	jor g17125(.dina(w_n17377_0[1]),.dinb(w_asqrt45_16[1]),.dout(n17379),.clk(gclk));
	jxor g17126(.dina(w_n16726_0[0]),.dinb(w_n2833_28[0]),.dout(n17380),.clk(gclk));
	jand g17127(.dina(n17380),.dinb(w_asqrt12_22[0]),.dout(n17381),.clk(gclk));
	jxor g17128(.dina(n17381),.dinb(w_n16731_0[0]),.dout(n17382),.clk(gclk));
	jand g17129(.dina(w_n17382_0[1]),.dinb(n17379),.dout(n17383),.clk(gclk));
	jor g17130(.dina(n17383),.dinb(w_n17378_0[1]),.dout(n17384),.clk(gclk));
	jand g17131(.dina(w_n17384_0[2]),.dinb(w_asqrt46_19[0]),.dout(n17385),.clk(gclk));
	jor g17132(.dina(w_n17384_0[1]),.dinb(w_asqrt46_18[2]),.dout(n17386),.clk(gclk));
	jxor g17133(.dina(w_n16734_0[0]),.dinb(w_n2572_30[2]),.dout(n17387),.clk(gclk));
	jand g17134(.dina(n17387),.dinb(w_asqrt12_21[2]),.dout(n17388),.clk(gclk));
	jxor g17135(.dina(n17388),.dinb(w_n16739_0[0]),.dout(n17389),.clk(gclk));
	jnot g17136(.din(w_n17389_0[1]),.dout(n17390),.clk(gclk));
	jand g17137(.dina(w_n17390_0[1]),.dinb(n17386),.dout(n17391),.clk(gclk));
	jor g17138(.dina(n17391),.dinb(w_n17385_0[1]),.dout(n17392),.clk(gclk));
	jand g17139(.dina(w_n17392_0[2]),.dinb(w_asqrt47_17[1]),.dout(n17393),.clk(gclk));
	jor g17140(.dina(w_n17392_0[1]),.dinb(w_asqrt47_17[0]),.dout(n17394),.clk(gclk));
	jxor g17141(.dina(w_n16741_0[0]),.dinb(w_n2345_28[2]),.dout(n17395),.clk(gclk));
	jand g17142(.dina(n17395),.dinb(w_asqrt12_21[1]),.dout(n17396),.clk(gclk));
	jxor g17143(.dina(n17396),.dinb(w_n16746_0[0]),.dout(n17397),.clk(gclk));
	jand g17144(.dina(w_n17397_0[1]),.dinb(n17394),.dout(n17398),.clk(gclk));
	jor g17145(.dina(n17398),.dinb(w_n17393_0[1]),.dout(n17399),.clk(gclk));
	jand g17146(.dina(w_n17399_0[2]),.dinb(w_asqrt48_19[1]),.dout(n17400),.clk(gclk));
	jor g17147(.dina(w_n17399_0[1]),.dinb(w_asqrt48_19[0]),.dout(n17401),.clk(gclk));
	jxor g17148(.dina(w_n16749_0[0]),.dinb(w_n2108_31[1]),.dout(n17402),.clk(gclk));
	jand g17149(.dina(n17402),.dinb(w_asqrt12_21[0]),.dout(n17403),.clk(gclk));
	jxor g17150(.dina(n17403),.dinb(w_n16754_0[0]),.dout(n17404),.clk(gclk));
	jnot g17151(.din(w_n17404_0[1]),.dout(n17405),.clk(gclk));
	jand g17152(.dina(w_n17405_0[1]),.dinb(n17401),.dout(n17406),.clk(gclk));
	jor g17153(.dina(n17406),.dinb(w_n17400_0[1]),.dout(n17407),.clk(gclk));
	jand g17154(.dina(w_n17407_0[2]),.dinb(w_asqrt49_17[2]),.dout(n17408),.clk(gclk));
	jor g17155(.dina(w_n17407_0[1]),.dinb(w_asqrt49_17[1]),.dout(n17409),.clk(gclk));
	jxor g17156(.dina(w_n16756_0[0]),.dinb(w_n1912_29[2]),.dout(n17410),.clk(gclk));
	jand g17157(.dina(n17410),.dinb(w_asqrt12_20[2]),.dout(n17411),.clk(gclk));
	jxor g17158(.dina(n17411),.dinb(w_n16761_0[0]),.dout(n17412),.clk(gclk));
	jnot g17159(.din(w_n17412_0[1]),.dout(n17413),.clk(gclk));
	jand g17160(.dina(w_n17413_0[1]),.dinb(n17409),.dout(n17414),.clk(gclk));
	jor g17161(.dina(n17414),.dinb(w_n17408_0[1]),.dout(n17415),.clk(gclk));
	jand g17162(.dina(w_n17415_0[2]),.dinb(w_asqrt50_19[2]),.dout(n17416),.clk(gclk));
	jor g17163(.dina(w_n17415_0[1]),.dinb(w_asqrt50_19[1]),.dout(n17417),.clk(gclk));
	jxor g17164(.dina(w_n16763_0[0]),.dinb(w_n1699_32[0]),.dout(n17418),.clk(gclk));
	jand g17165(.dina(n17418),.dinb(w_asqrt12_20[1]),.dout(n17419),.clk(gclk));
	jxor g17166(.dina(n17419),.dinb(w_n16768_0[0]),.dout(n17420),.clk(gclk));
	jand g17167(.dina(w_n17420_0[1]),.dinb(n17417),.dout(n17421),.clk(gclk));
	jor g17168(.dina(n17421),.dinb(w_n17416_0[1]),.dout(n17422),.clk(gclk));
	jand g17169(.dina(w_n17422_0[2]),.dinb(w_asqrt51_18[0]),.dout(n17423),.clk(gclk));
	jxor g17170(.dina(w_n16771_0[0]),.dinb(w_n1516_30[1]),.dout(n17424),.clk(gclk));
	jand g17171(.dina(n17424),.dinb(w_asqrt12_20[0]),.dout(n17425),.clk(gclk));
	jxor g17172(.dina(n17425),.dinb(w_n16775_0[0]),.dout(n17426),.clk(gclk));
	jor g17173(.dina(w_n17422_0[1]),.dinb(w_asqrt51_17[2]),.dout(n17427),.clk(gclk));
	jand g17174(.dina(n17427),.dinb(w_n17426_0[1]),.dout(n17428),.clk(gclk));
	jor g17175(.dina(n17428),.dinb(w_n17423_0[1]),.dout(n17429),.clk(gclk));
	jand g17176(.dina(w_n17429_0[2]),.dinb(w_asqrt52_19[2]),.dout(n17430),.clk(gclk));
	jor g17177(.dina(w_n17429_0[1]),.dinb(w_asqrt52_19[1]),.dout(n17431),.clk(gclk));
	jxor g17178(.dina(w_n16779_0[0]),.dinb(w_n1332_32[0]),.dout(n17432),.clk(gclk));
	jand g17179(.dina(n17432),.dinb(w_asqrt12_19[2]),.dout(n17433),.clk(gclk));
	jxor g17180(.dina(n17433),.dinb(w_n16784_0[0]),.dout(n17434),.clk(gclk));
	jnot g17181(.din(w_n17434_0[1]),.dout(n17435),.clk(gclk));
	jand g17182(.dina(w_n17435_0[1]),.dinb(n17431),.dout(n17436),.clk(gclk));
	jor g17183(.dina(n17436),.dinb(w_n17430_0[1]),.dout(n17437),.clk(gclk));
	jand g17184(.dina(w_n17437_0[2]),.dinb(w_asqrt53_18[2]),.dout(n17438),.clk(gclk));
	jor g17185(.dina(w_n17437_0[1]),.dinb(w_asqrt53_18[1]),.dout(n17439),.clk(gclk));
	jxor g17186(.dina(w_n16786_0[0]),.dinb(w_n1173_31[0]),.dout(n17440),.clk(gclk));
	jand g17187(.dina(n17440),.dinb(w_asqrt12_19[1]),.dout(n17441),.clk(gclk));
	jxor g17188(.dina(n17441),.dinb(w_n16791_0[0]),.dout(n17442),.clk(gclk));
	jand g17189(.dina(w_n17442_0[1]),.dinb(n17439),.dout(n17443),.clk(gclk));
	jor g17190(.dina(n17443),.dinb(w_n17438_0[1]),.dout(n17444),.clk(gclk));
	jand g17191(.dina(w_n17444_0[2]),.dinb(w_asqrt54_19[2]),.dout(n17445),.clk(gclk));
	jor g17192(.dina(w_n17444_0[1]),.dinb(w_asqrt54_19[1]),.dout(n17446),.clk(gclk));
	jxor g17193(.dina(w_n16794_0[0]),.dinb(w_n1008_33[0]),.dout(n17447),.clk(gclk));
	jand g17194(.dina(n17447),.dinb(w_asqrt12_19[0]),.dout(n17448),.clk(gclk));
	jxor g17195(.dina(n17448),.dinb(w_n16799_0[0]),.dout(n17449),.clk(gclk));
	jnot g17196(.din(w_n17449_0[1]),.dout(n17450),.clk(gclk));
	jand g17197(.dina(w_n17450_0[1]),.dinb(n17446),.dout(n17451),.clk(gclk));
	jor g17198(.dina(n17451),.dinb(w_n17445_0[1]),.dout(n17452),.clk(gclk));
	jand g17199(.dina(w_n17452_0[2]),.dinb(w_asqrt55_19[0]),.dout(n17453),.clk(gclk));
	jor g17200(.dina(w_n17452_0[1]),.dinb(w_asqrt55_18[2]),.dout(n17454),.clk(gclk));
	jxor g17201(.dina(w_n16801_0[0]),.dinb(w_n884_32[0]),.dout(n17455),.clk(gclk));
	jand g17202(.dina(n17455),.dinb(w_asqrt12_18[2]),.dout(n17456),.clk(gclk));
	jxor g17203(.dina(n17456),.dinb(w_n16806_0[0]),.dout(n17457),.clk(gclk));
	jand g17204(.dina(w_n17457_0[1]),.dinb(n17454),.dout(n17458),.clk(gclk));
	jor g17205(.dina(n17458),.dinb(w_n17453_0[1]),.dout(n17459),.clk(gclk));
	jand g17206(.dina(w_n17459_0[2]),.dinb(w_asqrt56_20[0]),.dout(n17460),.clk(gclk));
	jor g17207(.dina(w_n17459_0[1]),.dinb(w_asqrt56_19[2]),.dout(n17461),.clk(gclk));
	jxor g17208(.dina(w_n16809_0[0]),.dinb(w_n743_33[0]),.dout(n17462),.clk(gclk));
	jand g17209(.dina(n17462),.dinb(w_asqrt12_18[1]),.dout(n17463),.clk(gclk));
	jxor g17210(.dina(n17463),.dinb(w_n16814_0[0]),.dout(n17464),.clk(gclk));
	jnot g17211(.din(w_n17464_0[1]),.dout(n17465),.clk(gclk));
	jand g17212(.dina(w_n17465_0[1]),.dinb(n17461),.dout(n17466),.clk(gclk));
	jor g17213(.dina(n17466),.dinb(w_n17460_0[1]),.dout(n17467),.clk(gclk));
	jand g17214(.dina(w_n17467_0[2]),.dinb(w_asqrt57_19[2]),.dout(n17468),.clk(gclk));
	jor g17215(.dina(w_n17467_0[1]),.dinb(w_asqrt57_19[1]),.dout(n17469),.clk(gclk));
	jxor g17216(.dina(w_n16816_0[0]),.dinb(w_n635_33[0]),.dout(n17470),.clk(gclk));
	jand g17217(.dina(n17470),.dinb(w_asqrt12_18[0]),.dout(n17471),.clk(gclk));
	jxor g17218(.dina(n17471),.dinb(w_n16821_0[0]),.dout(n17472),.clk(gclk));
	jnot g17219(.din(w_n17472_0[1]),.dout(n17473),.clk(gclk));
	jand g17220(.dina(w_n17473_0[1]),.dinb(n17469),.dout(n17474),.clk(gclk));
	jor g17221(.dina(n17474),.dinb(w_n17468_0[1]),.dout(n17475),.clk(gclk));
	jand g17222(.dina(w_n17475_0[2]),.dinb(w_asqrt58_20[1]),.dout(n17476),.clk(gclk));
	jor g17223(.dina(w_n17475_0[1]),.dinb(w_asqrt58_20[0]),.dout(n17477),.clk(gclk));
	jxor g17224(.dina(w_n16823_0[0]),.dinb(w_n515_34[0]),.dout(n17478),.clk(gclk));
	jand g17225(.dina(n17478),.dinb(w_asqrt12_17[2]),.dout(n17479),.clk(gclk));
	jxor g17226(.dina(n17479),.dinb(w_n16828_0[0]),.dout(n17480),.clk(gclk));
	jnot g17227(.din(w_n17480_0[1]),.dout(n17481),.clk(gclk));
	jand g17228(.dina(w_n17481_0[1]),.dinb(n17477),.dout(n17482),.clk(gclk));
	jor g17229(.dina(n17482),.dinb(w_n17476_0[1]),.dout(n17483),.clk(gclk));
	jand g17230(.dina(w_n17483_0[2]),.dinb(w_asqrt59_20[0]),.dout(n17484),.clk(gclk));
	jor g17231(.dina(w_n17483_0[1]),.dinb(w_asqrt59_19[2]),.dout(n17485),.clk(gclk));
	jxor g17232(.dina(w_n16830_0[0]),.dinb(w_n443_34[0]),.dout(n17486),.clk(gclk));
	jand g17233(.dina(n17486),.dinb(w_asqrt12_17[1]),.dout(n17487),.clk(gclk));
	jxor g17234(.dina(n17487),.dinb(w_n16835_0[0]),.dout(n17488),.clk(gclk));
	jand g17235(.dina(w_n17488_0[1]),.dinb(n17485),.dout(n17489),.clk(gclk));
	jor g17236(.dina(n17489),.dinb(w_n17484_0[1]),.dout(n17490),.clk(gclk));
	jand g17237(.dina(w_n17490_0[2]),.dinb(w_asqrt60_20[1]),.dout(n17491),.clk(gclk));
	jor g17238(.dina(w_n17490_0[1]),.dinb(w_asqrt60_20[0]),.dout(n17492),.clk(gclk));
	jxor g17239(.dina(w_n16838_0[0]),.dinb(w_n352_34[1]),.dout(n17493),.clk(gclk));
	jand g17240(.dina(n17493),.dinb(w_asqrt12_17[0]),.dout(n17494),.clk(gclk));
	jxor g17241(.dina(n17494),.dinb(w_n16843_0[0]),.dout(n17495),.clk(gclk));
	jnot g17242(.din(w_n17495_0[1]),.dout(n17496),.clk(gclk));
	jand g17243(.dina(w_n17496_0[1]),.dinb(n17492),.dout(n17497),.clk(gclk));
	jor g17244(.dina(n17497),.dinb(w_n17491_0[1]),.dout(n17498),.clk(gclk));
	jand g17245(.dina(w_n17498_0[2]),.dinb(w_asqrt61_20[1]),.dout(n17499),.clk(gclk));
	jor g17246(.dina(w_n17498_0[1]),.dinb(w_asqrt61_20[0]),.dout(n17500),.clk(gclk));
	jxor g17247(.dina(w_n16845_0[0]),.dinb(w_n294_34[2]),.dout(n17501),.clk(gclk));
	jand g17248(.dina(n17501),.dinb(w_asqrt12_16[2]),.dout(n17502),.clk(gclk));
	jxor g17249(.dina(n17502),.dinb(w_n16850_0[0]),.dout(n17503),.clk(gclk));
	jand g17250(.dina(w_n17503_0[1]),.dinb(n17500),.dout(n17504),.clk(gclk));
	jor g17251(.dina(n17504),.dinb(w_n17499_0[1]),.dout(n17505),.clk(gclk));
	jand g17252(.dina(w_n17505_0[2]),.dinb(w_asqrt62_20[1]),.dout(n17506),.clk(gclk));
	jor g17253(.dina(w_n17505_0[1]),.dinb(w_asqrt62_20[0]),.dout(n17507),.clk(gclk));
	jxor g17254(.dina(w_n16853_0[0]),.dinb(w_n239_34[2]),.dout(n17508),.clk(gclk));
	jand g17255(.dina(n17508),.dinb(w_asqrt12_16[1]),.dout(n17509),.clk(gclk));
	jxor g17256(.dina(n17509),.dinb(w_n16858_0[0]),.dout(n17510),.clk(gclk));
	jnot g17257(.din(w_n17510_0[2]),.dout(n17511),.clk(gclk));
	jand g17258(.dina(n17511),.dinb(n17507),.dout(n17512),.clk(gclk));
	jor g17259(.dina(n17512),.dinb(w_n17506_0[1]),.dout(n17513),.clk(gclk));
	jxor g17260(.dina(w_n16860_0[0]),.dinb(w_n221_35[0]),.dout(n17514),.clk(gclk));
	jand g17261(.dina(n17514),.dinb(w_asqrt12_16[0]),.dout(n17515),.clk(gclk));
	jxor g17262(.dina(n17515),.dinb(w_n16866_0[0]),.dout(n17516),.clk(gclk));
	jnot g17263(.din(w_n17516_0[2]),.dout(n17517),.clk(gclk));
	jor g17264(.dina(w_n17517_0[1]),.dinb(w_n17513_0[1]),.dout(n17518),.clk(gclk));
	jnot g17265(.din(w_n17518_1[1]),.dout(n17519),.clk(gclk));
	jand g17266(.dina(w_n17132_0[0]),.dinb(w_n16868_0[0]),.dout(n17520),.clk(gclk));
	jnot g17267(.din(n17520),.dout(n17521),.clk(gclk));
	jand g17268(.dina(w_n16871_0[0]),.dinb(w_asqrt63_25[1]),.dout(n17522),.clk(gclk));
	jand g17269(.dina(n17522),.dinb(w_n16896_0[2]),.dout(n17523),.clk(gclk));
	jand g17270(.dina(w_n17523_0[1]),.dinb(n17521),.dout(n17524),.clk(gclk));
	jand g17271(.dina(w_n16882_0[0]),.dinb(w_n17127_0[0]),.dout(n17525),.clk(gclk));
	jnot g17272(.din(w_n17506_0[0]),.dout(n17526),.clk(gclk));
	jnot g17273(.din(w_n17499_0[0]),.dout(n17527),.clk(gclk));
	jnot g17274(.din(w_n17491_0[0]),.dout(n17528),.clk(gclk));
	jnot g17275(.din(w_n17484_0[0]),.dout(n17529),.clk(gclk));
	jnot g17276(.din(w_n17476_0[0]),.dout(n17530),.clk(gclk));
	jnot g17277(.din(w_n17468_0[0]),.dout(n17531),.clk(gclk));
	jnot g17278(.din(w_n17460_0[0]),.dout(n17532),.clk(gclk));
	jnot g17279(.din(w_n17453_0[0]),.dout(n17533),.clk(gclk));
	jnot g17280(.din(w_n17445_0[0]),.dout(n17534),.clk(gclk));
	jnot g17281(.din(w_n17438_0[0]),.dout(n17535),.clk(gclk));
	jnot g17282(.din(w_n17430_0[0]),.dout(n17536),.clk(gclk));
	jnot g17283(.din(w_n17423_0[0]),.dout(n17537),.clk(gclk));
	jnot g17284(.din(w_n17426_0[0]),.dout(n17538),.clk(gclk));
	jnot g17285(.din(w_n17416_0[0]),.dout(n17539),.clk(gclk));
	jnot g17286(.din(w_n17408_0[0]),.dout(n17540),.clk(gclk));
	jnot g17287(.din(w_n17400_0[0]),.dout(n17541),.clk(gclk));
	jnot g17288(.din(w_n17393_0[0]),.dout(n17542),.clk(gclk));
	jnot g17289(.din(w_n17385_0[0]),.dout(n17543),.clk(gclk));
	jnot g17290(.din(w_n17378_0[0]),.dout(n17544),.clk(gclk));
	jnot g17291(.din(w_n17370_0[0]),.dout(n17545),.clk(gclk));
	jnot g17292(.din(w_n17362_0[0]),.dout(n17546),.clk(gclk));
	jnot g17293(.din(w_n17354_0[0]),.dout(n17547),.clk(gclk));
	jnot g17294(.din(w_n17347_0[0]),.dout(n17548),.clk(gclk));
	jnot g17295(.din(w_n17339_0[0]),.dout(n17549),.clk(gclk));
	jnot g17296(.din(w_n17332_0[0]),.dout(n17550),.clk(gclk));
	jnot g17297(.din(w_n17324_0[0]),.dout(n17551),.clk(gclk));
	jnot g17298(.din(w_n17316_0[0]),.dout(n17552),.clk(gclk));
	jnot g17299(.din(w_n17308_0[0]),.dout(n17553),.clk(gclk));
	jnot g17300(.din(w_n17301_0[0]),.dout(n17554),.clk(gclk));
	jnot g17301(.din(w_n17293_0[0]),.dout(n17555),.clk(gclk));
	jnot g17302(.din(w_n17286_0[0]),.dout(n17556),.clk(gclk));
	jnot g17303(.din(w_n17278_0[0]),.dout(n17557),.clk(gclk));
	jnot g17304(.din(w_n17271_0[0]),.dout(n17558),.clk(gclk));
	jnot g17305(.din(w_n17263_0[0]),.dout(n17559),.clk(gclk));
	jnot g17306(.din(w_n17256_0[0]),.dout(n17560),.clk(gclk));
	jnot g17307(.din(w_n17248_0[0]),.dout(n17561),.clk(gclk));
	jnot g17308(.din(w_n17240_0[0]),.dout(n17562),.clk(gclk));
	jnot g17309(.din(w_n17232_0[0]),.dout(n17563),.clk(gclk));
	jnot g17310(.din(w_n17225_0[0]),.dout(n17564),.clk(gclk));
	jnot g17311(.din(w_n17217_0[0]),.dout(n17565),.clk(gclk));
	jnot g17312(.din(w_n17210_0[0]),.dout(n17566),.clk(gclk));
	jnot g17313(.din(w_n17202_0[0]),.dout(n17567),.clk(gclk));
	jnot g17314(.din(w_n17195_0[0]),.dout(n17568),.clk(gclk));
	jnot g17315(.din(w_n17188_0[0]),.dout(n17569),.clk(gclk));
	jnot g17316(.din(w_n17180_0[0]),.dout(n17570),.clk(gclk));
	jnot g17317(.din(w_n17172_0[0]),.dout(n17571),.clk(gclk));
	jnot g17318(.din(w_n17165_0[0]),.dout(n17572),.clk(gclk));
	jnot g17319(.din(w_n17157_0[0]),.dout(n17573),.clk(gclk));
	jnot g17320(.din(w_n17150_0[0]),.dout(n17574),.clk(gclk));
	jnot g17321(.din(w_n17139_0[0]),.dout(n17575),.clk(gclk));
	jnot g17322(.din(w_n16891_0[0]),.dout(n17576),.clk(gclk));
	jnot g17323(.din(w_n16888_0[0]),.dout(n17577),.clk(gclk));
	jor g17324(.dina(w_n17134_15[0]),.dinb(w_n16494_0[2]),.dout(n17578),.clk(gclk));
	jand g17325(.dina(n17578),.dinb(n17577),.dout(n17579),.clk(gclk));
	jand g17326(.dina(n17579),.dinb(w_n16489_22[1]),.dout(n17580),.clk(gclk));
	jor g17327(.dina(w_n17134_14[2]),.dinb(w_a24_0[0]),.dout(n17581),.clk(gclk));
	jand g17328(.dina(n17581),.dinb(w_a25_0[0]),.dout(n17582),.clk(gclk));
	jor g17329(.dina(w_n17141_0[0]),.dinb(n17582),.dout(n17583),.clk(gclk));
	jor g17330(.dina(w_n17583_0[1]),.dinb(n17580),.dout(n17584),.clk(gclk));
	jand g17331(.dina(n17584),.dinb(n17576),.dout(n17585),.clk(gclk));
	jand g17332(.dina(n17585),.dinb(w_n15878_15[1]),.dout(n17586),.clk(gclk));
	jor g17333(.dina(w_n17146_0[0]),.dinb(n17586),.dout(n17587),.clk(gclk));
	jand g17334(.dina(n17587),.dinb(n17575),.dout(n17588),.clk(gclk));
	jand g17335(.dina(n17588),.dinb(w_n15260_23[0]),.dout(n17589),.clk(gclk));
	jnot g17336(.din(w_n17154_0[0]),.dout(n17590),.clk(gclk));
	jor g17337(.dina(w_n17590_0[1]),.dinb(n17589),.dout(n17591),.clk(gclk));
	jand g17338(.dina(n17591),.dinb(n17574),.dout(n17592),.clk(gclk));
	jand g17339(.dina(n17592),.dinb(w_n14674_16[0]),.dout(n17593),.clk(gclk));
	jor g17340(.dina(w_n17161_0[0]),.dinb(n17593),.dout(n17594),.clk(gclk));
	jand g17341(.dina(n17594),.dinb(n17573),.dout(n17595),.clk(gclk));
	jand g17342(.dina(n17595),.dinb(w_n14078_23[1]),.dout(n17596),.clk(gclk));
	jnot g17343(.din(w_n17169_0[0]),.dout(n17597),.clk(gclk));
	jor g17344(.dina(w_n17597_0[1]),.dinb(n17596),.dout(n17598),.clk(gclk));
	jand g17345(.dina(n17598),.dinb(n17572),.dout(n17599),.clk(gclk));
	jand g17346(.dina(n17599),.dinb(w_n13515_17[0]),.dout(n17600),.clk(gclk));
	jor g17347(.dina(w_n17176_0[0]),.dinb(n17600),.dout(n17601),.clk(gclk));
	jand g17348(.dina(n17601),.dinb(n17571),.dout(n17602),.clk(gclk));
	jand g17349(.dina(n17602),.dinb(w_n12947_24[0]),.dout(n17603),.clk(gclk));
	jor g17350(.dina(w_n17184_0[0]),.dinb(n17603),.dout(n17604),.clk(gclk));
	jand g17351(.dina(n17604),.dinb(n17570),.dout(n17605),.clk(gclk));
	jand g17352(.dina(n17605),.dinb(w_n12410_17[2]),.dout(n17606),.clk(gclk));
	jnot g17353(.din(w_n17192_0[0]),.dout(n17607),.clk(gclk));
	jor g17354(.dina(w_n17607_0[1]),.dinb(n17606),.dout(n17608),.clk(gclk));
	jand g17355(.dina(n17608),.dinb(n17569),.dout(n17609),.clk(gclk));
	jand g17356(.dina(n17609),.dinb(w_n11858_24[1]),.dout(n17610),.clk(gclk));
	jnot g17357(.din(w_n17199_0[0]),.dout(n17611),.clk(gclk));
	jor g17358(.dina(w_n17611_0[1]),.dinb(n17610),.dout(n17612),.clk(gclk));
	jand g17359(.dina(n17612),.dinb(n17568),.dout(n17613),.clk(gclk));
	jand g17360(.dina(n17613),.dinb(w_n11347_18[1]),.dout(n17614),.clk(gclk));
	jor g17361(.dina(w_n17206_0[0]),.dinb(n17614),.dout(n17615),.clk(gclk));
	jand g17362(.dina(n17615),.dinb(n17567),.dout(n17616),.clk(gclk));
	jand g17363(.dina(n17616),.dinb(w_n10824_25[0]),.dout(n17617),.clk(gclk));
	jnot g17364(.din(w_n17214_0[0]),.dout(n17618),.clk(gclk));
	jor g17365(.dina(w_n17618_0[1]),.dinb(n17617),.dout(n17619),.clk(gclk));
	jand g17366(.dina(n17619),.dinb(n17566),.dout(n17620),.clk(gclk));
	jand g17367(.dina(n17620),.dinb(w_n10328_19[1]),.dout(n17621),.clk(gclk));
	jor g17368(.dina(w_n17221_0[0]),.dinb(n17621),.dout(n17622),.clk(gclk));
	jand g17369(.dina(n17622),.dinb(n17565),.dout(n17623),.clk(gclk));
	jand g17370(.dina(n17623),.dinb(w_n9832_25[2]),.dout(n17624),.clk(gclk));
	jnot g17371(.din(w_n17229_0[0]),.dout(n17625),.clk(gclk));
	jor g17372(.dina(w_n17625_0[1]),.dinb(n17624),.dout(n17626),.clk(gclk));
	jand g17373(.dina(n17626),.dinb(n17564),.dout(n17627),.clk(gclk));
	jand g17374(.dina(n17627),.dinb(w_n9369_20[1]),.dout(n17628),.clk(gclk));
	jor g17375(.dina(w_n17236_0[0]),.dinb(n17628),.dout(n17629),.clk(gclk));
	jand g17376(.dina(n17629),.dinb(n17563),.dout(n17630),.clk(gclk));
	jand g17377(.dina(n17630),.dinb(w_n8890_26[0]),.dout(n17631),.clk(gclk));
	jor g17378(.dina(w_n17244_0[0]),.dinb(n17631),.dout(n17632),.clk(gclk));
	jand g17379(.dina(n17632),.dinb(n17562),.dout(n17633),.clk(gclk));
	jand g17380(.dina(n17633),.dinb(w_n8449_21[0]),.dout(n17634),.clk(gclk));
	jor g17381(.dina(w_n17252_0[0]),.dinb(n17634),.dout(n17635),.clk(gclk));
	jand g17382(.dina(n17635),.dinb(n17561),.dout(n17636),.clk(gclk));
	jand g17383(.dina(n17636),.dinb(w_n8003_26[2]),.dout(n17637),.clk(gclk));
	jnot g17384(.din(w_n17260_0[0]),.dout(n17638),.clk(gclk));
	jor g17385(.dina(w_n17638_0[1]),.dinb(n17637),.dout(n17639),.clk(gclk));
	jand g17386(.dina(n17639),.dinb(n17560),.dout(n17640),.clk(gclk));
	jand g17387(.dina(n17640),.dinb(w_n7581_22[0]),.dout(n17641),.clk(gclk));
	jor g17388(.dina(w_n17267_0[0]),.dinb(n17641),.dout(n17642),.clk(gclk));
	jand g17389(.dina(n17642),.dinb(n17559),.dout(n17643),.clk(gclk));
	jand g17390(.dina(n17643),.dinb(w_n7154_27[0]),.dout(n17644),.clk(gclk));
	jnot g17391(.din(w_n17275_0[0]),.dout(n17645),.clk(gclk));
	jor g17392(.dina(w_n17645_0[1]),.dinb(n17644),.dout(n17646),.clk(gclk));
	jand g17393(.dina(n17646),.dinb(n17558),.dout(n17647),.clk(gclk));
	jand g17394(.dina(n17647),.dinb(w_n6758_22[2]),.dout(n17648),.clk(gclk));
	jor g17395(.dina(w_n17282_0[0]),.dinb(n17648),.dout(n17649),.clk(gclk));
	jand g17396(.dina(n17649),.dinb(n17557),.dout(n17650),.clk(gclk));
	jand g17397(.dina(n17650),.dinb(w_n6357_27[1]),.dout(n17651),.clk(gclk));
	jnot g17398(.din(w_n17290_0[0]),.dout(n17652),.clk(gclk));
	jor g17399(.dina(w_n17652_0[1]),.dinb(n17651),.dout(n17653),.clk(gclk));
	jand g17400(.dina(n17653),.dinb(n17556),.dout(n17654),.clk(gclk));
	jand g17401(.dina(n17654),.dinb(w_n5989_23[1]),.dout(n17655),.clk(gclk));
	jor g17402(.dina(w_n17297_0[0]),.dinb(n17655),.dout(n17656),.clk(gclk));
	jand g17403(.dina(n17656),.dinb(n17555),.dout(n17657),.clk(gclk));
	jand g17404(.dina(n17657),.dinb(w_n5606_27[2]),.dout(n17658),.clk(gclk));
	jnot g17405(.din(w_n17305_0[0]),.dout(n17659),.clk(gclk));
	jor g17406(.dina(w_n17659_0[1]),.dinb(n17658),.dout(n17660),.clk(gclk));
	jand g17407(.dina(n17660),.dinb(n17554),.dout(n17661),.clk(gclk));
	jand g17408(.dina(n17661),.dinb(w_n5259_24[1]),.dout(n17662),.clk(gclk));
	jor g17409(.dina(w_n17312_0[0]),.dinb(n17662),.dout(n17663),.clk(gclk));
	jand g17410(.dina(n17663),.dinb(n17553),.dout(n17664),.clk(gclk));
	jand g17411(.dina(n17664),.dinb(w_n4902_28[1]),.dout(n17665),.clk(gclk));
	jor g17412(.dina(w_n17320_0[0]),.dinb(n17665),.dout(n17666),.clk(gclk));
	jand g17413(.dina(n17666),.dinb(n17552),.dout(n17667),.clk(gclk));
	jand g17414(.dina(n17667),.dinb(w_n4582_25[1]),.dout(n17668),.clk(gclk));
	jor g17415(.dina(w_n17328_0[0]),.dinb(n17668),.dout(n17669),.clk(gclk));
	jand g17416(.dina(n17669),.dinb(n17551),.dout(n17670),.clk(gclk));
	jand g17417(.dina(n17670),.dinb(w_n4249_29[0]),.dout(n17671),.clk(gclk));
	jnot g17418(.din(w_n17336_0[0]),.dout(n17672),.clk(gclk));
	jor g17419(.dina(w_n17672_0[1]),.dinb(n17671),.dout(n17673),.clk(gclk));
	jand g17420(.dina(n17673),.dinb(n17550),.dout(n17674),.clk(gclk));
	jand g17421(.dina(n17674),.dinb(w_n3955_26[0]),.dout(n17675),.clk(gclk));
	jor g17422(.dina(w_n17343_0[0]),.dinb(n17675),.dout(n17676),.clk(gclk));
	jand g17423(.dina(n17676),.dinb(n17549),.dout(n17677),.clk(gclk));
	jand g17424(.dina(n17677),.dinb(w_n3642_29[1]),.dout(n17678),.clk(gclk));
	jnot g17425(.din(w_n17351_0[0]),.dout(n17679),.clk(gclk));
	jor g17426(.dina(w_n17679_0[1]),.dinb(n17678),.dout(n17680),.clk(gclk));
	jand g17427(.dina(n17680),.dinb(n17548),.dout(n17681),.clk(gclk));
	jand g17428(.dina(n17681),.dinb(w_n3368_26[2]),.dout(n17682),.clk(gclk));
	jor g17429(.dina(w_n17358_0[0]),.dinb(n17682),.dout(n17683),.clk(gclk));
	jand g17430(.dina(n17683),.dinb(n17547),.dout(n17684),.clk(gclk));
	jand g17431(.dina(n17684),.dinb(w_n3089_30[0]),.dout(n17685),.clk(gclk));
	jor g17432(.dina(w_n17366_0[0]),.dinb(n17685),.dout(n17686),.clk(gclk));
	jand g17433(.dina(n17686),.dinb(n17546),.dout(n17687),.clk(gclk));
	jand g17434(.dina(n17687),.dinb(w_n2833_27[2]),.dout(n17688),.clk(gclk));
	jor g17435(.dina(w_n17374_0[0]),.dinb(n17688),.dout(n17689),.clk(gclk));
	jand g17436(.dina(n17689),.dinb(n17545),.dout(n17690),.clk(gclk));
	jand g17437(.dina(n17690),.dinb(w_n2572_30[1]),.dout(n17691),.clk(gclk));
	jnot g17438(.din(w_n17382_0[0]),.dout(n17692),.clk(gclk));
	jor g17439(.dina(w_n17692_0[1]),.dinb(n17691),.dout(n17693),.clk(gclk));
	jand g17440(.dina(n17693),.dinb(n17544),.dout(n17694),.clk(gclk));
	jand g17441(.dina(n17694),.dinb(w_n2345_28[1]),.dout(n17695),.clk(gclk));
	jor g17442(.dina(w_n17389_0[0]),.dinb(n17695),.dout(n17696),.clk(gclk));
	jand g17443(.dina(n17696),.dinb(n17543),.dout(n17697),.clk(gclk));
	jand g17444(.dina(n17697),.dinb(w_n2108_31[0]),.dout(n17698),.clk(gclk));
	jnot g17445(.din(w_n17397_0[0]),.dout(n17699),.clk(gclk));
	jor g17446(.dina(w_n17699_0[1]),.dinb(n17698),.dout(n17700),.clk(gclk));
	jand g17447(.dina(n17700),.dinb(n17542),.dout(n17701),.clk(gclk));
	jand g17448(.dina(n17701),.dinb(w_n1912_29[1]),.dout(n17702),.clk(gclk));
	jor g17449(.dina(w_n17404_0[0]),.dinb(n17702),.dout(n17703),.clk(gclk));
	jand g17450(.dina(n17703),.dinb(n17541),.dout(n17704),.clk(gclk));
	jand g17451(.dina(n17704),.dinb(w_n1699_31[2]),.dout(n17705),.clk(gclk));
	jor g17452(.dina(w_n17412_0[0]),.dinb(n17705),.dout(n17706),.clk(gclk));
	jand g17453(.dina(n17706),.dinb(n17540),.dout(n17707),.clk(gclk));
	jand g17454(.dina(n17707),.dinb(w_n1516_30[0]),.dout(n17708),.clk(gclk));
	jnot g17455(.din(w_n17420_0[0]),.dout(n17709),.clk(gclk));
	jor g17456(.dina(w_n17709_0[1]),.dinb(n17708),.dout(n17710),.clk(gclk));
	jand g17457(.dina(n17710),.dinb(n17539),.dout(n17711),.clk(gclk));
	jand g17458(.dina(n17711),.dinb(w_n1332_31[2]),.dout(n17712),.clk(gclk));
	jor g17459(.dina(n17712),.dinb(w_n17538_0[1]),.dout(n17713),.clk(gclk));
	jand g17460(.dina(n17713),.dinb(n17537),.dout(n17714),.clk(gclk));
	jand g17461(.dina(n17714),.dinb(w_n1173_30[2]),.dout(n17715),.clk(gclk));
	jor g17462(.dina(w_n17434_0[0]),.dinb(n17715),.dout(n17716),.clk(gclk));
	jand g17463(.dina(n17716),.dinb(n17536),.dout(n17717),.clk(gclk));
	jand g17464(.dina(n17717),.dinb(w_n1008_32[2]),.dout(n17718),.clk(gclk));
	jnot g17465(.din(w_n17442_0[0]),.dout(n17719),.clk(gclk));
	jor g17466(.dina(w_n17719_0[1]),.dinb(n17718),.dout(n17720),.clk(gclk));
	jand g17467(.dina(n17720),.dinb(n17535),.dout(n17721),.clk(gclk));
	jand g17468(.dina(n17721),.dinb(w_n884_31[2]),.dout(n17722),.clk(gclk));
	jor g17469(.dina(w_n17449_0[0]),.dinb(n17722),.dout(n17723),.clk(gclk));
	jand g17470(.dina(n17723),.dinb(n17534),.dout(n17724),.clk(gclk));
	jand g17471(.dina(n17724),.dinb(w_n743_32[2]),.dout(n17725),.clk(gclk));
	jnot g17472(.din(w_n17457_0[0]),.dout(n17726),.clk(gclk));
	jor g17473(.dina(w_n17726_0[1]),.dinb(n17725),.dout(n17727),.clk(gclk));
	jand g17474(.dina(n17727),.dinb(n17533),.dout(n17728),.clk(gclk));
	jand g17475(.dina(n17728),.dinb(w_n635_32[2]),.dout(n17729),.clk(gclk));
	jor g17476(.dina(w_n17464_0[0]),.dinb(n17729),.dout(n17730),.clk(gclk));
	jand g17477(.dina(n17730),.dinb(n17532),.dout(n17731),.clk(gclk));
	jand g17478(.dina(n17731),.dinb(w_n515_33[2]),.dout(n17732),.clk(gclk));
	jor g17479(.dina(w_n17472_0[0]),.dinb(n17732),.dout(n17733),.clk(gclk));
	jand g17480(.dina(n17733),.dinb(n17531),.dout(n17734),.clk(gclk));
	jand g17481(.dina(n17734),.dinb(w_n443_33[2]),.dout(n17735),.clk(gclk));
	jor g17482(.dina(w_n17480_0[0]),.dinb(n17735),.dout(n17736),.clk(gclk));
	jand g17483(.dina(n17736),.dinb(n17530),.dout(n17737),.clk(gclk));
	jand g17484(.dina(n17737),.dinb(w_n352_34[0]),.dout(n17738),.clk(gclk));
	jnot g17485(.din(w_n17488_0[0]),.dout(n17739),.clk(gclk));
	jor g17486(.dina(w_n17739_0[1]),.dinb(n17738),.dout(n17740),.clk(gclk));
	jand g17487(.dina(n17740),.dinb(n17529),.dout(n17741),.clk(gclk));
	jand g17488(.dina(n17741),.dinb(w_n294_34[1]),.dout(n17742),.clk(gclk));
	jor g17489(.dina(w_n17495_0[0]),.dinb(n17742),.dout(n17743),.clk(gclk));
	jand g17490(.dina(n17743),.dinb(n17528),.dout(n17744),.clk(gclk));
	jand g17491(.dina(n17744),.dinb(w_n239_34[1]),.dout(n17745),.clk(gclk));
	jnot g17492(.din(w_n17503_0[0]),.dout(n17746),.clk(gclk));
	jor g17493(.dina(w_n17746_0[1]),.dinb(n17745),.dout(n17747),.clk(gclk));
	jand g17494(.dina(n17747),.dinb(n17527),.dout(n17748),.clk(gclk));
	jand g17495(.dina(n17748),.dinb(w_n221_34[2]),.dout(n17749),.clk(gclk));
	jor g17496(.dina(w_n17510_0[1]),.dinb(n17749),.dout(n17750),.clk(gclk));
	jand g17497(.dina(n17750),.dinb(n17526),.dout(n17751),.clk(gclk));
	jor g17498(.dina(w_n17516_0[1]),.dinb(w_n17751_0[1]),.dout(n17752),.clk(gclk));
	jor g17499(.dina(w_n17752_0[1]),.dinb(w_n16869_0[0]),.dout(n17753),.clk(gclk));
	jor g17500(.dina(n17753),.dinb(w_n17525_0[1]),.dout(n17754),.clk(gclk));
	jand g17501(.dina(n17754),.dinb(w_n218_14[2]),.dout(n17755),.clk(gclk));
	jand g17502(.dina(w_n17134_14[1]),.dinb(w_n16493_0[0]),.dout(n17756),.clk(gclk));
	jor g17503(.dina(w_n17756_0[1]),.dinb(w_n17755_0[1]),.dout(n17757),.clk(gclk));
	jor g17504(.dina(n17757),.dinb(w_n17524_0[1]),.dout(n17758),.clk(gclk));
	jor g17505(.dina(w_n17758_0[1]),.dinb(w_n17519_0[2]),.dout(asqrt_fa_12),.clk(gclk));
	jnot g17506(.din(w_n17524_0[0]),.dout(n17760),.clk(gclk));
	jnot g17507(.din(w_n17525_0[0]),.dout(n17761),.clk(gclk));
	jand g17508(.dina(w_n17517_0[0]),.dinb(w_n17513_0[0]),.dout(n17762),.clk(gclk));
	jand g17509(.dina(w_n17762_0[1]),.dinb(w_n16896_0[1]),.dout(n17763),.clk(gclk));
	jand g17510(.dina(n17763),.dinb(n17761),.dout(n17764),.clk(gclk));
	jor g17511(.dina(n17764),.dinb(w_asqrt63_25[0]),.dout(n17765),.clk(gclk));
	jnot g17512(.din(w_n17756_0[0]),.dout(n17766),.clk(gclk));
	jand g17513(.dina(n17766),.dinb(n17765),.dout(n17767),.clk(gclk));
	jand g17514(.dina(n17767),.dinb(n17760),.dout(n17768),.clk(gclk));
	jand g17515(.dina(w_n17768_0[1]),.dinb(w_n17518_1[0]),.dout(n17769),.clk(gclk));
	jxor g17516(.dina(w_n17505_0[0]),.dinb(w_n221_34[1]),.dout(n17770),.clk(gclk));
	jor g17517(.dina(n17770),.dinb(w_n17769_38[1]),.dout(n17771),.clk(gclk));
	jxor g17518(.dina(n17771),.dinb(w_n17510_0[0]),.dout(n17772),.clk(gclk));
	jnot g17519(.din(w_n17772_0[1]),.dout(n17773),.clk(gclk));
	jnot g17520(.din(w_a20_0[2]),.dout(n17774),.clk(gclk));
	jnot g17521(.din(w_a21_0[1]),.dout(n17775),.clk(gclk));
	jand g17522(.dina(w_n17775_0[1]),.dinb(w_n17774_1[2]),.dout(n17776),.clk(gclk));
	jand g17523(.dina(w_n17776_0[2]),.dinb(w_n16885_1[0]),.dout(n17777),.clk(gclk));
	jnot g17524(.din(w_n17777_0[1]),.dout(n17778),.clk(gclk));
	jor g17525(.dina(w_n17769_38[0]),.dinb(w_n16885_0[2]),.dout(n17779),.clk(gclk));
	jand g17526(.dina(n17779),.dinb(n17778),.dout(n17780),.clk(gclk));
	jor g17527(.dina(w_n17780_0[2]),.dinb(w_n17134_14[0]),.dout(n17781),.clk(gclk));
	jand g17528(.dina(w_n17780_0[1]),.dinb(w_n17134_13[2]),.dout(n17782),.clk(gclk));
	jor g17529(.dina(w_n17769_37[2]),.dinb(w_a22_1[0]),.dout(n17783),.clk(gclk));
	jand g17530(.dina(n17783),.dinb(w_a23_0[0]),.dout(n17784),.clk(gclk));
	jand g17531(.dina(w_asqrt11_8[1]),.dinb(w_n16887_0[1]),.dout(n17785),.clk(gclk));
	jor g17532(.dina(n17785),.dinb(n17784),.dout(n17786),.clk(gclk));
	jor g17533(.dina(n17786),.dinb(n17782),.dout(n17787),.clk(gclk));
	jand g17534(.dina(n17787),.dinb(w_n17781_0[1]),.dout(n17788),.clk(gclk));
	jor g17535(.dina(w_n17788_0[2]),.dinb(w_n16489_22[0]),.dout(n17789),.clk(gclk));
	jand g17536(.dina(w_n17788_0[1]),.dinb(w_n16489_21[2]),.dout(n17790),.clk(gclk));
	jnot g17537(.din(w_n16887_0[0]),.dout(n17791),.clk(gclk));
	jor g17538(.dina(w_n17769_37[1]),.dinb(n17791),.dout(n17792),.clk(gclk));
	jor g17539(.dina(w_n17519_0[1]),.dinb(w_n17134_13[1]),.dout(n17793),.clk(gclk));
	jor g17540(.dina(n17793),.dinb(w_n17523_0[0]),.dout(n17794),.clk(gclk));
	jor g17541(.dina(n17794),.dinb(w_n17755_0[0]),.dout(n17795),.clk(gclk));
	jand g17542(.dina(n17795),.dinb(w_n17792_0[1]),.dout(n17796),.clk(gclk));
	jxor g17543(.dina(n17796),.dinb(w_n16494_0[1]),.dout(n17797),.clk(gclk));
	jor g17544(.dina(w_n17797_0[2]),.dinb(n17790),.dout(n17798),.clk(gclk));
	jand g17545(.dina(n17798),.dinb(w_n17789_0[1]),.dout(n17799),.clk(gclk));
	jor g17546(.dina(w_n17799_0[2]),.dinb(w_n15878_15[0]),.dout(n17800),.clk(gclk));
	jand g17547(.dina(w_n17799_0[1]),.dinb(w_n15878_14[2]),.dout(n17801),.clk(gclk));
	jxor g17548(.dina(w_n16890_0[0]),.dinb(w_n16489_21[1]),.dout(n17802),.clk(gclk));
	jor g17549(.dina(n17802),.dinb(w_n17769_37[0]),.dout(n17803),.clk(gclk));
	jxor g17550(.dina(n17803),.dinb(w_n17583_0[0]),.dout(n17804),.clk(gclk));
	jnot g17551(.din(w_n17804_0[2]),.dout(n17805),.clk(gclk));
	jor g17552(.dina(n17805),.dinb(n17801),.dout(n17806),.clk(gclk));
	jand g17553(.dina(n17806),.dinb(w_n17800_0[1]),.dout(n17807),.clk(gclk));
	jor g17554(.dina(w_n17807_0[2]),.dinb(w_n15260_22[2]),.dout(n17808),.clk(gclk));
	jand g17555(.dina(w_n17807_0[1]),.dinb(w_n15260_22[1]),.dout(n17809),.clk(gclk));
	jxor g17556(.dina(w_n17138_0[0]),.dinb(w_n15878_14[1]),.dout(n17810),.clk(gclk));
	jor g17557(.dina(n17810),.dinb(w_n17769_36[2]),.dout(n17811),.clk(gclk));
	jxor g17558(.dina(n17811),.dinb(w_n17147_0[0]),.dout(n17812),.clk(gclk));
	jor g17559(.dina(w_n17812_0[2]),.dinb(n17809),.dout(n17813),.clk(gclk));
	jand g17560(.dina(n17813),.dinb(w_n17808_0[1]),.dout(n17814),.clk(gclk));
	jor g17561(.dina(w_n17814_0[2]),.dinb(w_n14674_15[2]),.dout(n17815),.clk(gclk));
	jand g17562(.dina(w_n17814_0[1]),.dinb(w_n14674_15[1]),.dout(n17816),.clk(gclk));
	jxor g17563(.dina(w_n17149_0[0]),.dinb(w_n15260_22[0]),.dout(n17817),.clk(gclk));
	jor g17564(.dina(n17817),.dinb(w_n17769_36[1]),.dout(n17818),.clk(gclk));
	jxor g17565(.dina(n17818),.dinb(w_n17590_0[0]),.dout(n17819),.clk(gclk));
	jnot g17566(.din(w_n17819_0[2]),.dout(n17820),.clk(gclk));
	jor g17567(.dina(n17820),.dinb(n17816),.dout(n17821),.clk(gclk));
	jand g17568(.dina(n17821),.dinb(w_n17815_0[1]),.dout(n17822),.clk(gclk));
	jor g17569(.dina(w_n17822_0[2]),.dinb(w_n14078_23[0]),.dout(n17823),.clk(gclk));
	jand g17570(.dina(w_n17822_0[1]),.dinb(w_n14078_22[2]),.dout(n17824),.clk(gclk));
	jxor g17571(.dina(w_n17156_0[0]),.dinb(w_n14674_15[0]),.dout(n17825),.clk(gclk));
	jor g17572(.dina(n17825),.dinb(w_n17769_36[0]),.dout(n17826),.clk(gclk));
	jxor g17573(.dina(n17826),.dinb(w_n17162_0[0]),.dout(n17827),.clk(gclk));
	jor g17574(.dina(w_n17827_0[2]),.dinb(n17824),.dout(n17828),.clk(gclk));
	jand g17575(.dina(n17828),.dinb(w_n17823_0[1]),.dout(n17829),.clk(gclk));
	jor g17576(.dina(w_n17829_0[2]),.dinb(w_n13515_16[2]),.dout(n17830),.clk(gclk));
	jand g17577(.dina(w_n17829_0[1]),.dinb(w_n13515_16[1]),.dout(n17831),.clk(gclk));
	jxor g17578(.dina(w_n17164_0[0]),.dinb(w_n14078_22[1]),.dout(n17832),.clk(gclk));
	jor g17579(.dina(n17832),.dinb(w_n17769_35[2]),.dout(n17833),.clk(gclk));
	jxor g17580(.dina(n17833),.dinb(w_n17597_0[0]),.dout(n17834),.clk(gclk));
	jnot g17581(.din(w_n17834_0[2]),.dout(n17835),.clk(gclk));
	jor g17582(.dina(n17835),.dinb(n17831),.dout(n17836),.clk(gclk));
	jand g17583(.dina(n17836),.dinb(w_n17830_0[1]),.dout(n17837),.clk(gclk));
	jor g17584(.dina(w_n17837_0[2]),.dinb(w_n12947_23[2]),.dout(n17838),.clk(gclk));
	jand g17585(.dina(w_n17837_0[1]),.dinb(w_n12947_23[1]),.dout(n17839),.clk(gclk));
	jxor g17586(.dina(w_n17171_0[0]),.dinb(w_n13515_16[0]),.dout(n17840),.clk(gclk));
	jor g17587(.dina(n17840),.dinb(w_n17769_35[1]),.dout(n17841),.clk(gclk));
	jxor g17588(.dina(n17841),.dinb(w_n17177_0[0]),.dout(n17842),.clk(gclk));
	jor g17589(.dina(w_n17842_0[2]),.dinb(n17839),.dout(n17843),.clk(gclk));
	jand g17590(.dina(n17843),.dinb(w_n17838_0[1]),.dout(n17844),.clk(gclk));
	jor g17591(.dina(w_n17844_0[2]),.dinb(w_n12410_17[1]),.dout(n17845),.clk(gclk));
	jand g17592(.dina(w_n17844_0[1]),.dinb(w_n12410_17[0]),.dout(n17846),.clk(gclk));
	jxor g17593(.dina(w_n17179_0[0]),.dinb(w_n12947_23[0]),.dout(n17847),.clk(gclk));
	jor g17594(.dina(n17847),.dinb(w_n17769_35[0]),.dout(n17848),.clk(gclk));
	jxor g17595(.dina(n17848),.dinb(w_n17185_0[0]),.dout(n17849),.clk(gclk));
	jor g17596(.dina(w_n17849_0[2]),.dinb(n17846),.dout(n17850),.clk(gclk));
	jand g17597(.dina(n17850),.dinb(w_n17845_0[1]),.dout(n17851),.clk(gclk));
	jor g17598(.dina(w_n17851_0[2]),.dinb(w_n11858_24[0]),.dout(n17852),.clk(gclk));
	jand g17599(.dina(w_n17851_0[1]),.dinb(w_n11858_23[2]),.dout(n17853),.clk(gclk));
	jxor g17600(.dina(w_n17187_0[0]),.dinb(w_n12410_16[2]),.dout(n17854),.clk(gclk));
	jor g17601(.dina(n17854),.dinb(w_n17769_34[2]),.dout(n17855),.clk(gclk));
	jxor g17602(.dina(n17855),.dinb(w_n17607_0[0]),.dout(n17856),.clk(gclk));
	jnot g17603(.din(w_n17856_0[2]),.dout(n17857),.clk(gclk));
	jor g17604(.dina(n17857),.dinb(n17853),.dout(n17858),.clk(gclk));
	jand g17605(.dina(n17858),.dinb(w_n17852_0[1]),.dout(n17859),.clk(gclk));
	jor g17606(.dina(w_n17859_0[2]),.dinb(w_n11347_18[0]),.dout(n17860),.clk(gclk));
	jand g17607(.dina(w_n17859_0[1]),.dinb(w_n11347_17[2]),.dout(n17861),.clk(gclk));
	jxor g17608(.dina(w_n17194_0[0]),.dinb(w_n11858_23[1]),.dout(n17862),.clk(gclk));
	jor g17609(.dina(n17862),.dinb(w_n17769_34[1]),.dout(n17863),.clk(gclk));
	jxor g17610(.dina(n17863),.dinb(w_n17611_0[0]),.dout(n17864),.clk(gclk));
	jnot g17611(.din(w_n17864_0[2]),.dout(n17865),.clk(gclk));
	jor g17612(.dina(n17865),.dinb(n17861),.dout(n17866),.clk(gclk));
	jand g17613(.dina(n17866),.dinb(w_n17860_0[1]),.dout(n17867),.clk(gclk));
	jor g17614(.dina(w_n17867_0[2]),.dinb(w_n10824_24[2]),.dout(n17868),.clk(gclk));
	jand g17615(.dina(w_n17867_0[1]),.dinb(w_n10824_24[1]),.dout(n17869),.clk(gclk));
	jxor g17616(.dina(w_n17201_0[0]),.dinb(w_n11347_17[1]),.dout(n17870),.clk(gclk));
	jor g17617(.dina(n17870),.dinb(w_n17769_34[0]),.dout(n17871),.clk(gclk));
	jxor g17618(.dina(n17871),.dinb(w_n17207_0[0]),.dout(n17872),.clk(gclk));
	jor g17619(.dina(w_n17872_0[2]),.dinb(n17869),.dout(n17873),.clk(gclk));
	jand g17620(.dina(n17873),.dinb(w_n17868_0[1]),.dout(n17874),.clk(gclk));
	jor g17621(.dina(w_n17874_0[2]),.dinb(w_n10328_19[0]),.dout(n17875),.clk(gclk));
	jand g17622(.dina(w_n17874_0[1]),.dinb(w_n10328_18[2]),.dout(n17876),.clk(gclk));
	jxor g17623(.dina(w_n17209_0[0]),.dinb(w_n10824_24[0]),.dout(n17877),.clk(gclk));
	jor g17624(.dina(n17877),.dinb(w_n17769_33[2]),.dout(n17878),.clk(gclk));
	jxor g17625(.dina(n17878),.dinb(w_n17618_0[0]),.dout(n17879),.clk(gclk));
	jnot g17626(.din(w_n17879_0[2]),.dout(n17880),.clk(gclk));
	jor g17627(.dina(n17880),.dinb(n17876),.dout(n17881),.clk(gclk));
	jand g17628(.dina(n17881),.dinb(w_n17875_0[1]),.dout(n17882),.clk(gclk));
	jor g17629(.dina(w_n17882_0[2]),.dinb(w_n9832_25[1]),.dout(n17883),.clk(gclk));
	jand g17630(.dina(w_n17882_0[1]),.dinb(w_n9832_25[0]),.dout(n17884),.clk(gclk));
	jxor g17631(.dina(w_n17216_0[0]),.dinb(w_n10328_18[1]),.dout(n17885),.clk(gclk));
	jor g17632(.dina(n17885),.dinb(w_n17769_33[1]),.dout(n17886),.clk(gclk));
	jxor g17633(.dina(n17886),.dinb(w_n17222_0[0]),.dout(n17887),.clk(gclk));
	jor g17634(.dina(w_n17887_0[2]),.dinb(n17884),.dout(n17888),.clk(gclk));
	jand g17635(.dina(n17888),.dinb(w_n17883_0[1]),.dout(n17889),.clk(gclk));
	jor g17636(.dina(w_n17889_0[2]),.dinb(w_n9369_20[0]),.dout(n17890),.clk(gclk));
	jand g17637(.dina(w_n17889_0[1]),.dinb(w_n9369_19[2]),.dout(n17891),.clk(gclk));
	jxor g17638(.dina(w_n17224_0[0]),.dinb(w_n9832_24[2]),.dout(n17892),.clk(gclk));
	jor g17639(.dina(n17892),.dinb(w_n17769_33[0]),.dout(n17893),.clk(gclk));
	jxor g17640(.dina(n17893),.dinb(w_n17625_0[0]),.dout(n17894),.clk(gclk));
	jnot g17641(.din(w_n17894_0[2]),.dout(n17895),.clk(gclk));
	jor g17642(.dina(n17895),.dinb(n17891),.dout(n17896),.clk(gclk));
	jand g17643(.dina(n17896),.dinb(w_n17890_0[1]),.dout(n17897),.clk(gclk));
	jor g17644(.dina(w_n17897_0[2]),.dinb(w_n8890_25[2]),.dout(n17898),.clk(gclk));
	jand g17645(.dina(w_n17897_0[1]),.dinb(w_n8890_25[1]),.dout(n17899),.clk(gclk));
	jxor g17646(.dina(w_n17231_0[0]),.dinb(w_n9369_19[1]),.dout(n17900),.clk(gclk));
	jor g17647(.dina(n17900),.dinb(w_n17769_32[2]),.dout(n17901),.clk(gclk));
	jxor g17648(.dina(n17901),.dinb(w_n17237_0[0]),.dout(n17902),.clk(gclk));
	jor g17649(.dina(w_n17902_0[2]),.dinb(n17899),.dout(n17903),.clk(gclk));
	jand g17650(.dina(n17903),.dinb(w_n17898_0[1]),.dout(n17904),.clk(gclk));
	jor g17651(.dina(w_n17904_0[2]),.dinb(w_n8449_20[2]),.dout(n17905),.clk(gclk));
	jand g17652(.dina(w_n17904_0[1]),.dinb(w_n8449_20[1]),.dout(n17906),.clk(gclk));
	jxor g17653(.dina(w_n17239_0[0]),.dinb(w_n8890_25[0]),.dout(n17907),.clk(gclk));
	jor g17654(.dina(n17907),.dinb(w_n17769_32[1]),.dout(n17908),.clk(gclk));
	jxor g17655(.dina(n17908),.dinb(w_n17245_0[0]),.dout(n17909),.clk(gclk));
	jor g17656(.dina(w_n17909_0[2]),.dinb(n17906),.dout(n17910),.clk(gclk));
	jand g17657(.dina(n17910),.dinb(w_n17905_0[1]),.dout(n17911),.clk(gclk));
	jor g17658(.dina(w_n17911_0[2]),.dinb(w_n8003_26[1]),.dout(n17912),.clk(gclk));
	jand g17659(.dina(w_n17911_0[1]),.dinb(w_n8003_26[0]),.dout(n17913),.clk(gclk));
	jxor g17660(.dina(w_n17247_0[0]),.dinb(w_n8449_20[0]),.dout(n17914),.clk(gclk));
	jor g17661(.dina(n17914),.dinb(w_n17769_32[0]),.dout(n17915),.clk(gclk));
	jxor g17662(.dina(n17915),.dinb(w_n17253_0[0]),.dout(n17916),.clk(gclk));
	jor g17663(.dina(w_n17916_0[2]),.dinb(n17913),.dout(n17917),.clk(gclk));
	jand g17664(.dina(n17917),.dinb(w_n17912_0[1]),.dout(n17918),.clk(gclk));
	jor g17665(.dina(w_n17918_0[2]),.dinb(w_n7581_21[2]),.dout(n17919),.clk(gclk));
	jand g17666(.dina(w_n17918_0[1]),.dinb(w_n7581_21[1]),.dout(n17920),.clk(gclk));
	jxor g17667(.dina(w_n17255_0[0]),.dinb(w_n8003_25[2]),.dout(n17921),.clk(gclk));
	jor g17668(.dina(n17921),.dinb(w_n17769_31[2]),.dout(n17922),.clk(gclk));
	jxor g17669(.dina(n17922),.dinb(w_n17638_0[0]),.dout(n17923),.clk(gclk));
	jnot g17670(.din(w_n17923_0[2]),.dout(n17924),.clk(gclk));
	jor g17671(.dina(n17924),.dinb(n17920),.dout(n17925),.clk(gclk));
	jand g17672(.dina(n17925),.dinb(w_n17919_0[1]),.dout(n17926),.clk(gclk));
	jor g17673(.dina(w_n17926_0[2]),.dinb(w_n7154_26[2]),.dout(n17927),.clk(gclk));
	jand g17674(.dina(w_n17926_0[1]),.dinb(w_n7154_26[1]),.dout(n17928),.clk(gclk));
	jxor g17675(.dina(w_n17262_0[0]),.dinb(w_n7581_21[0]),.dout(n17929),.clk(gclk));
	jor g17676(.dina(n17929),.dinb(w_n17769_31[1]),.dout(n17930),.clk(gclk));
	jxor g17677(.dina(n17930),.dinb(w_n17268_0[0]),.dout(n17931),.clk(gclk));
	jor g17678(.dina(w_n17931_0[2]),.dinb(n17928),.dout(n17932),.clk(gclk));
	jand g17679(.dina(n17932),.dinb(w_n17927_0[1]),.dout(n17933),.clk(gclk));
	jor g17680(.dina(w_n17933_0[2]),.dinb(w_n6758_22[1]),.dout(n17934),.clk(gclk));
	jand g17681(.dina(w_n17933_0[1]),.dinb(w_n6758_22[0]),.dout(n17935),.clk(gclk));
	jxor g17682(.dina(w_n17270_0[0]),.dinb(w_n7154_26[0]),.dout(n17936),.clk(gclk));
	jor g17683(.dina(n17936),.dinb(w_n17769_31[0]),.dout(n17937),.clk(gclk));
	jxor g17684(.dina(n17937),.dinb(w_n17645_0[0]),.dout(n17938),.clk(gclk));
	jnot g17685(.din(w_n17938_0[2]),.dout(n17939),.clk(gclk));
	jor g17686(.dina(n17939),.dinb(n17935),.dout(n17940),.clk(gclk));
	jand g17687(.dina(n17940),.dinb(w_n17934_0[1]),.dout(n17941),.clk(gclk));
	jor g17688(.dina(w_n17941_0[2]),.dinb(w_n6357_27[0]),.dout(n17942),.clk(gclk));
	jand g17689(.dina(w_n17941_0[1]),.dinb(w_n6357_26[2]),.dout(n17943),.clk(gclk));
	jxor g17690(.dina(w_n17277_0[0]),.dinb(w_n6758_21[2]),.dout(n17944),.clk(gclk));
	jor g17691(.dina(n17944),.dinb(w_n17769_30[2]),.dout(n17945),.clk(gclk));
	jxor g17692(.dina(n17945),.dinb(w_n17283_0[0]),.dout(n17946),.clk(gclk));
	jor g17693(.dina(w_n17946_0[2]),.dinb(n17943),.dout(n17947),.clk(gclk));
	jand g17694(.dina(n17947),.dinb(w_n17942_0[1]),.dout(n17948),.clk(gclk));
	jor g17695(.dina(w_n17948_0[2]),.dinb(w_n5989_23[0]),.dout(n17949),.clk(gclk));
	jand g17696(.dina(w_n17948_0[1]),.dinb(w_n5989_22[2]),.dout(n17950),.clk(gclk));
	jxor g17697(.dina(w_n17285_0[0]),.dinb(w_n6357_26[1]),.dout(n17951),.clk(gclk));
	jor g17698(.dina(n17951),.dinb(w_n17769_30[1]),.dout(n17952),.clk(gclk));
	jxor g17699(.dina(n17952),.dinb(w_n17652_0[0]),.dout(n17953),.clk(gclk));
	jnot g17700(.din(w_n17953_0[2]),.dout(n17954),.clk(gclk));
	jor g17701(.dina(n17954),.dinb(n17950),.dout(n17955),.clk(gclk));
	jand g17702(.dina(n17955),.dinb(w_n17949_0[1]),.dout(n17956),.clk(gclk));
	jor g17703(.dina(w_n17956_0[2]),.dinb(w_n5606_27[1]),.dout(n17957),.clk(gclk));
	jand g17704(.dina(w_n17956_0[1]),.dinb(w_n5606_27[0]),.dout(n17958),.clk(gclk));
	jxor g17705(.dina(w_n17292_0[0]),.dinb(w_n5989_22[1]),.dout(n17959),.clk(gclk));
	jor g17706(.dina(n17959),.dinb(w_n17769_30[0]),.dout(n17960),.clk(gclk));
	jxor g17707(.dina(n17960),.dinb(w_n17298_0[0]),.dout(n17961),.clk(gclk));
	jor g17708(.dina(w_n17961_0[2]),.dinb(n17958),.dout(n17962),.clk(gclk));
	jand g17709(.dina(n17962),.dinb(w_n17957_0[1]),.dout(n17963),.clk(gclk));
	jor g17710(.dina(w_n17963_0[2]),.dinb(w_n5259_24[0]),.dout(n17964),.clk(gclk));
	jand g17711(.dina(w_n17963_0[1]),.dinb(w_n5259_23[2]),.dout(n17965),.clk(gclk));
	jxor g17712(.dina(w_n17300_0[0]),.dinb(w_n5606_26[2]),.dout(n17966),.clk(gclk));
	jor g17713(.dina(n17966),.dinb(w_n17769_29[2]),.dout(n17967),.clk(gclk));
	jxor g17714(.dina(n17967),.dinb(w_n17659_0[0]),.dout(n17968),.clk(gclk));
	jnot g17715(.din(w_n17968_0[2]),.dout(n17969),.clk(gclk));
	jor g17716(.dina(n17969),.dinb(n17965),.dout(n17970),.clk(gclk));
	jand g17717(.dina(n17970),.dinb(w_n17964_0[1]),.dout(n17971),.clk(gclk));
	jor g17718(.dina(w_n17971_0[2]),.dinb(w_n4902_28[0]),.dout(n17972),.clk(gclk));
	jand g17719(.dina(w_n17971_0[1]),.dinb(w_n4902_27[2]),.dout(n17973),.clk(gclk));
	jxor g17720(.dina(w_n17307_0[0]),.dinb(w_n5259_23[1]),.dout(n17974),.clk(gclk));
	jor g17721(.dina(n17974),.dinb(w_n17769_29[1]),.dout(n17975),.clk(gclk));
	jxor g17722(.dina(n17975),.dinb(w_n17313_0[0]),.dout(n17976),.clk(gclk));
	jor g17723(.dina(w_n17976_0[2]),.dinb(n17973),.dout(n17977),.clk(gclk));
	jand g17724(.dina(n17977),.dinb(w_n17972_0[1]),.dout(n17978),.clk(gclk));
	jor g17725(.dina(w_n17978_0[2]),.dinb(w_n4582_25[0]),.dout(n17979),.clk(gclk));
	jand g17726(.dina(w_n17978_0[1]),.dinb(w_n4582_24[2]),.dout(n17980),.clk(gclk));
	jxor g17727(.dina(w_n17315_0[0]),.dinb(w_n4902_27[1]),.dout(n17981),.clk(gclk));
	jor g17728(.dina(n17981),.dinb(w_n17769_29[0]),.dout(n17982),.clk(gclk));
	jxor g17729(.dina(n17982),.dinb(w_n17321_0[0]),.dout(n17983),.clk(gclk));
	jor g17730(.dina(w_n17983_0[2]),.dinb(n17980),.dout(n17984),.clk(gclk));
	jand g17731(.dina(n17984),.dinb(w_n17979_0[1]),.dout(n17985),.clk(gclk));
	jor g17732(.dina(w_n17985_0[2]),.dinb(w_n4249_28[2]),.dout(n17986),.clk(gclk));
	jand g17733(.dina(w_n17985_0[1]),.dinb(w_n4249_28[1]),.dout(n17987),.clk(gclk));
	jxor g17734(.dina(w_n17323_0[0]),.dinb(w_n4582_24[1]),.dout(n17988),.clk(gclk));
	jor g17735(.dina(n17988),.dinb(w_n17769_28[2]),.dout(n17989),.clk(gclk));
	jxor g17736(.dina(n17989),.dinb(w_n17329_0[0]),.dout(n17990),.clk(gclk));
	jor g17737(.dina(w_n17990_0[2]),.dinb(n17987),.dout(n17991),.clk(gclk));
	jand g17738(.dina(n17991),.dinb(w_n17986_0[1]),.dout(n17992),.clk(gclk));
	jor g17739(.dina(w_n17992_0[2]),.dinb(w_n3955_25[2]),.dout(n17993),.clk(gclk));
	jand g17740(.dina(w_n17992_0[1]),.dinb(w_n3955_25[1]),.dout(n17994),.clk(gclk));
	jxor g17741(.dina(w_n17331_0[0]),.dinb(w_n4249_28[0]),.dout(n17995),.clk(gclk));
	jor g17742(.dina(n17995),.dinb(w_n17769_28[1]),.dout(n17996),.clk(gclk));
	jxor g17743(.dina(n17996),.dinb(w_n17672_0[0]),.dout(n17997),.clk(gclk));
	jnot g17744(.din(w_n17997_0[2]),.dout(n17998),.clk(gclk));
	jor g17745(.dina(n17998),.dinb(n17994),.dout(n17999),.clk(gclk));
	jand g17746(.dina(n17999),.dinb(w_n17993_0[1]),.dout(n18000),.clk(gclk));
	jor g17747(.dina(w_n18000_0[2]),.dinb(w_n3642_29[0]),.dout(n18001),.clk(gclk));
	jand g17748(.dina(w_n18000_0[1]),.dinb(w_n3642_28[2]),.dout(n18002),.clk(gclk));
	jxor g17749(.dina(w_n17338_0[0]),.dinb(w_n3955_25[0]),.dout(n18003),.clk(gclk));
	jor g17750(.dina(n18003),.dinb(w_n17769_28[0]),.dout(n18004),.clk(gclk));
	jxor g17751(.dina(n18004),.dinb(w_n17344_0[0]),.dout(n18005),.clk(gclk));
	jor g17752(.dina(w_n18005_0[2]),.dinb(n18002),.dout(n18006),.clk(gclk));
	jand g17753(.dina(n18006),.dinb(w_n18001_0[1]),.dout(n18007),.clk(gclk));
	jor g17754(.dina(w_n18007_0[2]),.dinb(w_n3368_26[1]),.dout(n18008),.clk(gclk));
	jand g17755(.dina(w_n18007_0[1]),.dinb(w_n3368_26[0]),.dout(n18009),.clk(gclk));
	jxor g17756(.dina(w_n17346_0[0]),.dinb(w_n3642_28[1]),.dout(n18010),.clk(gclk));
	jor g17757(.dina(n18010),.dinb(w_n17769_27[2]),.dout(n18011),.clk(gclk));
	jxor g17758(.dina(n18011),.dinb(w_n17679_0[0]),.dout(n18012),.clk(gclk));
	jnot g17759(.din(w_n18012_0[1]),.dout(n18013),.clk(gclk));
	jor g17760(.dina(w_n18013_0[1]),.dinb(n18009),.dout(n18014),.clk(gclk));
	jand g17761(.dina(n18014),.dinb(w_n18008_0[1]),.dout(n18015),.clk(gclk));
	jor g17762(.dina(w_n18015_0[2]),.dinb(w_n3089_29[2]),.dout(n18016),.clk(gclk));
	jand g17763(.dina(w_n18015_0[1]),.dinb(w_n3089_29[1]),.dout(n18017),.clk(gclk));
	jxor g17764(.dina(w_n17353_0[0]),.dinb(w_n3368_25[2]),.dout(n18018),.clk(gclk));
	jor g17765(.dina(n18018),.dinb(w_n17769_27[1]),.dout(n18019),.clk(gclk));
	jxor g17766(.dina(n18019),.dinb(w_n17359_0[0]),.dout(n18020),.clk(gclk));
	jor g17767(.dina(w_n18020_0[2]),.dinb(n18017),.dout(n18021),.clk(gclk));
	jand g17768(.dina(n18021),.dinb(w_n18016_0[1]),.dout(n18022),.clk(gclk));
	jor g17769(.dina(w_n18022_0[2]),.dinb(w_n2833_27[1]),.dout(n18023),.clk(gclk));
	jand g17770(.dina(w_n18022_0[1]),.dinb(w_n2833_27[0]),.dout(n18024),.clk(gclk));
	jxor g17771(.dina(w_n17361_0[0]),.dinb(w_n3089_29[0]),.dout(n18025),.clk(gclk));
	jor g17772(.dina(n18025),.dinb(w_n17769_27[0]),.dout(n18026),.clk(gclk));
	jxor g17773(.dina(n18026),.dinb(w_n17367_0[0]),.dout(n18027),.clk(gclk));
	jor g17774(.dina(w_n18027_0[2]),.dinb(n18024),.dout(n18028),.clk(gclk));
	jand g17775(.dina(n18028),.dinb(w_n18023_0[1]),.dout(n18029),.clk(gclk));
	jor g17776(.dina(w_n18029_0[2]),.dinb(w_n2572_30[0]),.dout(n18030),.clk(gclk));
	jand g17777(.dina(w_n18029_0[1]),.dinb(w_n2572_29[2]),.dout(n18031),.clk(gclk));
	jxor g17778(.dina(w_n17369_0[0]),.dinb(w_n2833_26[2]),.dout(n18032),.clk(gclk));
	jor g17779(.dina(n18032),.dinb(w_n17769_26[2]),.dout(n18033),.clk(gclk));
	jxor g17780(.dina(n18033),.dinb(w_n17375_0[0]),.dout(n18034),.clk(gclk));
	jor g17781(.dina(w_n18034_0[2]),.dinb(n18031),.dout(n18035),.clk(gclk));
	jand g17782(.dina(n18035),.dinb(w_n18030_0[1]),.dout(n18036),.clk(gclk));
	jor g17783(.dina(w_n18036_0[2]),.dinb(w_n2345_28[0]),.dout(n18037),.clk(gclk));
	jand g17784(.dina(w_n18036_0[1]),.dinb(w_n2345_27[2]),.dout(n18038),.clk(gclk));
	jxor g17785(.dina(w_n17377_0[0]),.dinb(w_n2572_29[1]),.dout(n18039),.clk(gclk));
	jor g17786(.dina(n18039),.dinb(w_n17769_26[1]),.dout(n18040),.clk(gclk));
	jxor g17787(.dina(n18040),.dinb(w_n17692_0[0]),.dout(n18041),.clk(gclk));
	jnot g17788(.din(w_n18041_0[2]),.dout(n18042),.clk(gclk));
	jor g17789(.dina(n18042),.dinb(n18038),.dout(n18043),.clk(gclk));
	jand g17790(.dina(n18043),.dinb(w_n18037_0[1]),.dout(n18044),.clk(gclk));
	jor g17791(.dina(w_n18044_0[2]),.dinb(w_n2108_30[2]),.dout(n18045),.clk(gclk));
	jand g17792(.dina(w_n18044_0[1]),.dinb(w_n2108_30[1]),.dout(n18046),.clk(gclk));
	jxor g17793(.dina(w_n17384_0[0]),.dinb(w_n2345_27[1]),.dout(n18047),.clk(gclk));
	jor g17794(.dina(n18047),.dinb(w_n17769_26[0]),.dout(n18048),.clk(gclk));
	jxor g17795(.dina(n18048),.dinb(w_n17390_0[0]),.dout(n18049),.clk(gclk));
	jor g17796(.dina(w_n18049_0[2]),.dinb(n18046),.dout(n18050),.clk(gclk));
	jand g17797(.dina(n18050),.dinb(w_n18045_0[1]),.dout(n18051),.clk(gclk));
	jor g17798(.dina(w_n18051_0[2]),.dinb(w_n1912_29[0]),.dout(n18052),.clk(gclk));
	jand g17799(.dina(w_n18051_0[1]),.dinb(w_n1912_28[2]),.dout(n18053),.clk(gclk));
	jxor g17800(.dina(w_n17392_0[0]),.dinb(w_n2108_30[0]),.dout(n18054),.clk(gclk));
	jor g17801(.dina(n18054),.dinb(w_n17769_25[2]),.dout(n18055),.clk(gclk));
	jxor g17802(.dina(n18055),.dinb(w_n17699_0[0]),.dout(n18056),.clk(gclk));
	jnot g17803(.din(w_n18056_0[2]),.dout(n18057),.clk(gclk));
	jor g17804(.dina(n18057),.dinb(n18053),.dout(n18058),.clk(gclk));
	jand g17805(.dina(n18058),.dinb(w_n18052_0[1]),.dout(n18059),.clk(gclk));
	jor g17806(.dina(w_n18059_0[2]),.dinb(w_n1699_31[1]),.dout(n18060),.clk(gclk));
	jand g17807(.dina(w_n18059_0[1]),.dinb(w_n1699_31[0]),.dout(n18061),.clk(gclk));
	jxor g17808(.dina(w_n17399_0[0]),.dinb(w_n1912_28[1]),.dout(n18062),.clk(gclk));
	jor g17809(.dina(n18062),.dinb(w_n17769_25[1]),.dout(n18063),.clk(gclk));
	jxor g17810(.dina(n18063),.dinb(w_n17405_0[0]),.dout(n18064),.clk(gclk));
	jor g17811(.dina(w_n18064_0[2]),.dinb(n18061),.dout(n18065),.clk(gclk));
	jand g17812(.dina(n18065),.dinb(w_n18060_0[1]),.dout(n18066),.clk(gclk));
	jor g17813(.dina(w_n18066_0[2]),.dinb(w_n1516_29[2]),.dout(n18067),.clk(gclk));
	jand g17814(.dina(w_n18066_0[1]),.dinb(w_n1516_29[1]),.dout(n18068),.clk(gclk));
	jxor g17815(.dina(w_n17407_0[0]),.dinb(w_n1699_30[2]),.dout(n18069),.clk(gclk));
	jor g17816(.dina(n18069),.dinb(w_n17769_25[0]),.dout(n18070),.clk(gclk));
	jxor g17817(.dina(n18070),.dinb(w_n17413_0[0]),.dout(n18071),.clk(gclk));
	jor g17818(.dina(w_n18071_0[2]),.dinb(n18068),.dout(n18072),.clk(gclk));
	jand g17819(.dina(n18072),.dinb(w_n18067_0[1]),.dout(n18073),.clk(gclk));
	jor g17820(.dina(w_n18073_0[2]),.dinb(w_n1332_31[1]),.dout(n18074),.clk(gclk));
	jand g17821(.dina(w_n18073_0[1]),.dinb(w_n1332_31[0]),.dout(n18075),.clk(gclk));
	jxor g17822(.dina(w_n17415_0[0]),.dinb(w_n1516_29[0]),.dout(n18076),.clk(gclk));
	jor g17823(.dina(n18076),.dinb(w_n17769_24[2]),.dout(n18077),.clk(gclk));
	jxor g17824(.dina(n18077),.dinb(w_n17709_0[0]),.dout(n18078),.clk(gclk));
	jnot g17825(.din(w_n18078_0[2]),.dout(n18079),.clk(gclk));
	jor g17826(.dina(n18079),.dinb(n18075),.dout(n18080),.clk(gclk));
	jand g17827(.dina(n18080),.dinb(w_n18074_0[1]),.dout(n18081),.clk(gclk));
	jor g17828(.dina(w_n18081_0[2]),.dinb(w_n1173_30[1]),.dout(n18082),.clk(gclk));
	jxor g17829(.dina(w_n17422_0[0]),.dinb(w_n1332_30[2]),.dout(n18083),.clk(gclk));
	jor g17830(.dina(n18083),.dinb(w_n17769_24[1]),.dout(n18084),.clk(gclk));
	jxor g17831(.dina(n18084),.dinb(w_n17538_0[0]),.dout(n18085),.clk(gclk));
	jnot g17832(.din(w_n18085_0[2]),.dout(n18086),.clk(gclk));
	jand g17833(.dina(w_n18081_0[1]),.dinb(w_n1173_30[0]),.dout(n18087),.clk(gclk));
	jor g17834(.dina(n18087),.dinb(n18086),.dout(n18088),.clk(gclk));
	jand g17835(.dina(n18088),.dinb(w_n18082_0[1]),.dout(n18089),.clk(gclk));
	jor g17836(.dina(w_n18089_0[2]),.dinb(w_n1008_32[1]),.dout(n18090),.clk(gclk));
	jand g17837(.dina(w_n18089_0[1]),.dinb(w_n1008_32[0]),.dout(n18091),.clk(gclk));
	jxor g17838(.dina(w_n17429_0[0]),.dinb(w_n1173_29[2]),.dout(n18092),.clk(gclk));
	jor g17839(.dina(n18092),.dinb(w_n17769_24[0]),.dout(n18093),.clk(gclk));
	jxor g17840(.dina(n18093),.dinb(w_n17435_0[0]),.dout(n18094),.clk(gclk));
	jor g17841(.dina(w_n18094_0[2]),.dinb(n18091),.dout(n18095),.clk(gclk));
	jand g17842(.dina(n18095),.dinb(w_n18090_0[1]),.dout(n18096),.clk(gclk));
	jor g17843(.dina(w_n18096_0[2]),.dinb(w_n884_31[1]),.dout(n18097),.clk(gclk));
	jand g17844(.dina(w_n18096_0[1]),.dinb(w_n884_31[0]),.dout(n18098),.clk(gclk));
	jxor g17845(.dina(w_n17437_0[0]),.dinb(w_n1008_31[2]),.dout(n18099),.clk(gclk));
	jor g17846(.dina(n18099),.dinb(w_n17769_23[2]),.dout(n18100),.clk(gclk));
	jxor g17847(.dina(n18100),.dinb(w_n17719_0[0]),.dout(n18101),.clk(gclk));
	jnot g17848(.din(w_n18101_0[2]),.dout(n18102),.clk(gclk));
	jor g17849(.dina(n18102),.dinb(n18098),.dout(n18103),.clk(gclk));
	jand g17850(.dina(n18103),.dinb(w_n18097_0[1]),.dout(n18104),.clk(gclk));
	jor g17851(.dina(w_n18104_0[2]),.dinb(w_n743_32[1]),.dout(n18105),.clk(gclk));
	jand g17852(.dina(w_n18104_0[1]),.dinb(w_n743_32[0]),.dout(n18106),.clk(gclk));
	jxor g17853(.dina(w_n17444_0[0]),.dinb(w_n884_30[2]),.dout(n18107),.clk(gclk));
	jor g17854(.dina(n18107),.dinb(w_n17769_23[1]),.dout(n18108),.clk(gclk));
	jxor g17855(.dina(n18108),.dinb(w_n17450_0[0]),.dout(n18109),.clk(gclk));
	jor g17856(.dina(w_n18109_0[2]),.dinb(n18106),.dout(n18110),.clk(gclk));
	jand g17857(.dina(n18110),.dinb(w_n18105_0[1]),.dout(n18111),.clk(gclk));
	jor g17858(.dina(w_n18111_0[2]),.dinb(w_n635_32[1]),.dout(n18112),.clk(gclk));
	jand g17859(.dina(w_n18111_0[1]),.dinb(w_n635_32[0]),.dout(n18113),.clk(gclk));
	jxor g17860(.dina(w_n17452_0[0]),.dinb(w_n743_31[2]),.dout(n18114),.clk(gclk));
	jor g17861(.dina(n18114),.dinb(w_n17769_23[0]),.dout(n18115),.clk(gclk));
	jxor g17862(.dina(n18115),.dinb(w_n17726_0[0]),.dout(n18116),.clk(gclk));
	jnot g17863(.din(w_n18116_0[2]),.dout(n18117),.clk(gclk));
	jor g17864(.dina(n18117),.dinb(n18113),.dout(n18118),.clk(gclk));
	jand g17865(.dina(n18118),.dinb(w_n18112_0[1]),.dout(n18119),.clk(gclk));
	jor g17866(.dina(w_n18119_0[2]),.dinb(w_n515_33[1]),.dout(n18120),.clk(gclk));
	jand g17867(.dina(w_n18119_0[1]),.dinb(w_n515_33[0]),.dout(n18121),.clk(gclk));
	jxor g17868(.dina(w_n17459_0[0]),.dinb(w_n635_31[2]),.dout(n18122),.clk(gclk));
	jor g17869(.dina(n18122),.dinb(w_n17769_22[2]),.dout(n18123),.clk(gclk));
	jxor g17870(.dina(n18123),.dinb(w_n17465_0[0]),.dout(n18124),.clk(gclk));
	jor g17871(.dina(w_n18124_0[2]),.dinb(n18121),.dout(n18125),.clk(gclk));
	jand g17872(.dina(n18125),.dinb(w_n18120_0[1]),.dout(n18126),.clk(gclk));
	jor g17873(.dina(w_n18126_0[2]),.dinb(w_n443_33[1]),.dout(n18127),.clk(gclk));
	jand g17874(.dina(w_n18126_0[1]),.dinb(w_n443_33[0]),.dout(n18128),.clk(gclk));
	jxor g17875(.dina(w_n17467_0[0]),.dinb(w_n515_32[2]),.dout(n18129),.clk(gclk));
	jor g17876(.dina(n18129),.dinb(w_n17769_22[1]),.dout(n18130),.clk(gclk));
	jxor g17877(.dina(n18130),.dinb(w_n17473_0[0]),.dout(n18131),.clk(gclk));
	jor g17878(.dina(w_n18131_0[2]),.dinb(n18128),.dout(n18132),.clk(gclk));
	jand g17879(.dina(n18132),.dinb(w_n18127_0[1]),.dout(n18133),.clk(gclk));
	jor g17880(.dina(w_n18133_0[2]),.dinb(w_n352_33[2]),.dout(n18134),.clk(gclk));
	jand g17881(.dina(w_n18133_0[1]),.dinb(w_n352_33[1]),.dout(n18135),.clk(gclk));
	jxor g17882(.dina(w_n17475_0[0]),.dinb(w_n443_32[2]),.dout(n18136),.clk(gclk));
	jor g17883(.dina(n18136),.dinb(w_n17769_22[0]),.dout(n18137),.clk(gclk));
	jxor g17884(.dina(n18137),.dinb(w_n17481_0[0]),.dout(n18138),.clk(gclk));
	jor g17885(.dina(w_n18138_0[2]),.dinb(n18135),.dout(n18139),.clk(gclk));
	jand g17886(.dina(n18139),.dinb(w_n18134_0[1]),.dout(n18140),.clk(gclk));
	jor g17887(.dina(w_n18140_0[2]),.dinb(w_n294_34[0]),.dout(n18141),.clk(gclk));
	jand g17888(.dina(w_n18140_0[1]),.dinb(w_n294_33[2]),.dout(n18142),.clk(gclk));
	jxor g17889(.dina(w_n17483_0[0]),.dinb(w_n352_33[0]),.dout(n18143),.clk(gclk));
	jor g17890(.dina(n18143),.dinb(w_n17769_21[2]),.dout(n18144),.clk(gclk));
	jxor g17891(.dina(n18144),.dinb(w_n17739_0[0]),.dout(n18145),.clk(gclk));
	jnot g17892(.din(w_n18145_0[2]),.dout(n18146),.clk(gclk));
	jor g17893(.dina(n18146),.dinb(n18142),.dout(n18147),.clk(gclk));
	jand g17894(.dina(n18147),.dinb(w_n18141_0[1]),.dout(n18148),.clk(gclk));
	jor g17895(.dina(w_n18148_0[2]),.dinb(w_n239_34[0]),.dout(n18149),.clk(gclk));
	jand g17896(.dina(w_n18148_0[1]),.dinb(w_n239_33[2]),.dout(n18150),.clk(gclk));
	jxor g17897(.dina(w_n17490_0[0]),.dinb(w_n294_33[1]),.dout(n18151),.clk(gclk));
	jor g17898(.dina(n18151),.dinb(w_n17769_21[1]),.dout(n18152),.clk(gclk));
	jxor g17899(.dina(n18152),.dinb(w_n17496_0[0]),.dout(n18153),.clk(gclk));
	jor g17900(.dina(w_n18153_0[2]),.dinb(n18150),.dout(n18154),.clk(gclk));
	jand g17901(.dina(n18154),.dinb(w_n18149_0[1]),.dout(n18155),.clk(gclk));
	jor g17902(.dina(w_n18155_0[2]),.dinb(w_n221_34[0]),.dout(n18156),.clk(gclk));
	jand g17903(.dina(w_n18155_0[1]),.dinb(w_n221_33[2]),.dout(n18157),.clk(gclk));
	jxor g17904(.dina(w_n17498_0[0]),.dinb(w_n239_33[1]),.dout(n18158),.clk(gclk));
	jor g17905(.dina(n18158),.dinb(w_n17769_21[0]),.dout(n18159),.clk(gclk));
	jxor g17906(.dina(n18159),.dinb(w_n17746_0[0]),.dout(n18160),.clk(gclk));
	jnot g17907(.din(w_n18160_0[2]),.dout(n18161),.clk(gclk));
	jor g17908(.dina(n18161),.dinb(n18157),.dout(n18162),.clk(gclk));
	jand g17909(.dina(n18162),.dinb(w_n18156_0[1]),.dout(n18163),.clk(gclk));
	jand g17910(.dina(w_n18163_0[2]),.dinb(w_n17773_0[2]),.dout(n18164),.clk(gclk));
	jand g17911(.dina(w_n17768_0[0]),.dinb(w_n17751_0[0]),.dout(n18165),.clk(gclk));
	jand g17912(.dina(w_n17752_0[0]),.dinb(w_asqrt63_24[2]),.dout(n18166),.clk(gclk));
	jand g17913(.dina(n18166),.dinb(w_n17518_0[2]),.dout(n18167),.clk(gclk));
	jnot g17914(.din(n18167),.dout(n18168),.clk(gclk));
	jor g17915(.dina(w_n18168_0[1]),.dinb(n18165),.dout(n18169),.clk(gclk));
	jnot g17916(.din(w_n18169_0[1]),.dout(n18170),.clk(gclk));
	jand g17917(.dina(w_n17758_0[0]),.dinb(w_n17762_0[0]),.dout(n18171),.clk(gclk));
	jor g17918(.dina(w_n18163_0[1]),.dinb(w_n17773_0[1]),.dout(n18172),.clk(gclk));
	jor g17919(.dina(w_n18172_0[1]),.dinb(w_n17519_0[0]),.dout(n18173),.clk(gclk));
	jor g17920(.dina(n18173),.dinb(w_n18171_0[1]),.dout(n18174),.clk(gclk));
	jand g17921(.dina(n18174),.dinb(w_n218_14[1]),.dout(n18175),.clk(gclk));
	jand g17922(.dina(w_n17769_20[2]),.dinb(w_n17516_0[0]),.dout(n18176),.clk(gclk));
	jor g17923(.dina(w_n18176_0[1]),.dinb(n18175),.dout(n18177),.clk(gclk));
	jor g17924(.dina(n18177),.dinb(n18170),.dout(n18178),.clk(gclk));
	jor g17925(.dina(w_n18178_0[1]),.dinb(w_n18164_0[2]),.dout(asqrt_fa_11),.clk(gclk));
	jxor g17926(.dina(w_n18155_0[0]),.dinb(w_n221_33[1]),.dout(n18180),.clk(gclk));
	jand g17927(.dina(n18180),.dinb(w_asqrt10_32[1]),.dout(n18181),.clk(gclk));
	jxor g17928(.dina(n18181),.dinb(w_n18160_0[1]),.dout(n18182),.clk(gclk));
	jnot g17929(.din(w_n18182_1[1]),.dout(n18183),.clk(gclk));
	jand g17930(.dina(w_asqrt10_32[0]),.dinb(w_a20_0[1]),.dout(n18184),.clk(gclk));
	jnot g17931(.din(w_a18_1[1]),.dout(n18185),.clk(gclk));
	jnot g17932(.din(w_a19_0[1]),.dout(n18186),.clk(gclk));
	jand g17933(.dina(w_n18186_0[1]),.dinb(w_n18185_1[1]),.dout(n18187),.clk(gclk));
	jand g17934(.dina(w_n18187_0[2]),.dinb(w_n17774_1[1]),.dout(n18188),.clk(gclk));
	jor g17935(.dina(w_n18188_0[1]),.dinb(n18184),.dout(n18189),.clk(gclk));
	jand g17936(.dina(w_n18189_0[2]),.dinb(w_asqrt11_8[0]),.dout(n18190),.clk(gclk));
	jor g17937(.dina(w_n18189_0[1]),.dinb(w_asqrt11_7[2]),.dout(n18191),.clk(gclk));
	jand g17938(.dina(w_asqrt10_31[2]),.dinb(w_n17774_1[0]),.dout(n18192),.clk(gclk));
	jor g17939(.dina(n18192),.dinb(w_n17775_0[0]),.dout(n18193),.clk(gclk));
	jnot g17940(.din(w_n17776_0[1]),.dout(n18194),.clk(gclk));
	jnot g17941(.din(w_n18164_0[1]),.dout(n18195),.clk(gclk));
	jnot g17942(.din(w_n18171_0[0]),.dout(n18196),.clk(gclk));
	jnot g17943(.din(w_n18156_0[0]),.dout(n18197),.clk(gclk));
	jnot g17944(.din(w_n18149_0[0]),.dout(n18198),.clk(gclk));
	jnot g17945(.din(w_n18141_0[0]),.dout(n18199),.clk(gclk));
	jnot g17946(.din(w_n18134_0[0]),.dout(n18200),.clk(gclk));
	jnot g17947(.din(w_n18127_0[0]),.dout(n18201),.clk(gclk));
	jnot g17948(.din(w_n18120_0[0]),.dout(n18202),.clk(gclk));
	jnot g17949(.din(w_n18112_0[0]),.dout(n18203),.clk(gclk));
	jnot g17950(.din(w_n18105_0[0]),.dout(n18204),.clk(gclk));
	jnot g17951(.din(w_n18097_0[0]),.dout(n18205),.clk(gclk));
	jnot g17952(.din(w_n18090_0[0]),.dout(n18206),.clk(gclk));
	jnot g17953(.din(w_n18082_0[0]),.dout(n18207),.clk(gclk));
	jnot g17954(.din(w_n18074_0[0]),.dout(n18208),.clk(gclk));
	jnot g17955(.din(w_n18067_0[0]),.dout(n18209),.clk(gclk));
	jnot g17956(.din(w_n18060_0[0]),.dout(n18210),.clk(gclk));
	jnot g17957(.din(w_n18052_0[0]),.dout(n18211),.clk(gclk));
	jnot g17958(.din(w_n18045_0[0]),.dout(n18212),.clk(gclk));
	jnot g17959(.din(w_n18037_0[0]),.dout(n18213),.clk(gclk));
	jnot g17960(.din(w_n18030_0[0]),.dout(n18214),.clk(gclk));
	jnot g17961(.din(w_n18023_0[0]),.dout(n18215),.clk(gclk));
	jnot g17962(.din(w_n18016_0[0]),.dout(n18216),.clk(gclk));
	jnot g17963(.din(w_n18008_0[0]),.dout(n18217),.clk(gclk));
	jnot g17964(.din(w_n18001_0[0]),.dout(n18218),.clk(gclk));
	jnot g17965(.din(w_n17993_0[0]),.dout(n18219),.clk(gclk));
	jnot g17966(.din(w_n17986_0[0]),.dout(n18220),.clk(gclk));
	jnot g17967(.din(w_n17979_0[0]),.dout(n18221),.clk(gclk));
	jnot g17968(.din(w_n17972_0[0]),.dout(n18222),.clk(gclk));
	jnot g17969(.din(w_n17964_0[0]),.dout(n18223),.clk(gclk));
	jnot g17970(.din(w_n17957_0[0]),.dout(n18224),.clk(gclk));
	jnot g17971(.din(w_n17949_0[0]),.dout(n18225),.clk(gclk));
	jnot g17972(.din(w_n17942_0[0]),.dout(n18226),.clk(gclk));
	jnot g17973(.din(w_n17934_0[0]),.dout(n18227),.clk(gclk));
	jnot g17974(.din(w_n17927_0[0]),.dout(n18228),.clk(gclk));
	jnot g17975(.din(w_n17919_0[0]),.dout(n18229),.clk(gclk));
	jnot g17976(.din(w_n17912_0[0]),.dout(n18230),.clk(gclk));
	jnot g17977(.din(w_n17905_0[0]),.dout(n18231),.clk(gclk));
	jnot g17978(.din(w_n17898_0[0]),.dout(n18232),.clk(gclk));
	jnot g17979(.din(w_n17890_0[0]),.dout(n18233),.clk(gclk));
	jnot g17980(.din(w_n17883_0[0]),.dout(n18234),.clk(gclk));
	jnot g17981(.din(w_n17875_0[0]),.dout(n18235),.clk(gclk));
	jnot g17982(.din(w_n17868_0[0]),.dout(n18236),.clk(gclk));
	jnot g17983(.din(w_n17860_0[0]),.dout(n18237),.clk(gclk));
	jnot g17984(.din(w_n17852_0[0]),.dout(n18238),.clk(gclk));
	jnot g17985(.din(w_n17845_0[0]),.dout(n18239),.clk(gclk));
	jnot g17986(.din(w_n17838_0[0]),.dout(n18240),.clk(gclk));
	jnot g17987(.din(w_n17830_0[0]),.dout(n18241),.clk(gclk));
	jnot g17988(.din(w_n17823_0[0]),.dout(n18242),.clk(gclk));
	jnot g17989(.din(w_n17815_0[0]),.dout(n18243),.clk(gclk));
	jnot g17990(.din(w_n17808_0[0]),.dout(n18244),.clk(gclk));
	jnot g17991(.din(w_n17800_0[0]),.dout(n18245),.clk(gclk));
	jnot g17992(.din(w_n17789_0[0]),.dout(n18246),.clk(gclk));
	jnot g17993(.din(w_n17781_0[0]),.dout(n18247),.clk(gclk));
	jand g17994(.dina(w_asqrt11_7[1]),.dinb(w_a22_0[2]),.dout(n18248),.clk(gclk));
	jor g17995(.dina(n18248),.dinb(w_n17777_0[0]),.dout(n18249),.clk(gclk));
	jor g17996(.dina(n18249),.dinb(w_asqrt12_15[2]),.dout(n18250),.clk(gclk));
	jand g17997(.dina(w_asqrt11_7[0]),.dinb(w_n16885_0[1]),.dout(n18251),.clk(gclk));
	jor g17998(.dina(n18251),.dinb(w_n16886_0[0]),.dout(n18252),.clk(gclk));
	jand g17999(.dina(w_n17792_0[0]),.dinb(n18252),.dout(n18253),.clk(gclk));
	jand g18000(.dina(w_n18253_0[1]),.dinb(n18250),.dout(n18254),.clk(gclk));
	jor g18001(.dina(n18254),.dinb(n18247),.dout(n18255),.clk(gclk));
	jor g18002(.dina(n18255),.dinb(w_asqrt13_8[0]),.dout(n18256),.clk(gclk));
	jnot g18003(.din(w_n17797_0[1]),.dout(n18257),.clk(gclk));
	jand g18004(.dina(n18257),.dinb(n18256),.dout(n18258),.clk(gclk));
	jor g18005(.dina(n18258),.dinb(n18246),.dout(n18259),.clk(gclk));
	jor g18006(.dina(n18259),.dinb(w_asqrt14_16[0]),.dout(n18260),.clk(gclk));
	jand g18007(.dina(w_n17804_0[1]),.dinb(n18260),.dout(n18261),.clk(gclk));
	jor g18008(.dina(n18261),.dinb(n18245),.dout(n18262),.clk(gclk));
	jor g18009(.dina(n18262),.dinb(w_asqrt15_8[2]),.dout(n18263),.clk(gclk));
	jnot g18010(.din(w_n17812_0[1]),.dout(n18264),.clk(gclk));
	jand g18011(.dina(n18264),.dinb(n18263),.dout(n18265),.clk(gclk));
	jor g18012(.dina(n18265),.dinb(n18244),.dout(n18266),.clk(gclk));
	jor g18013(.dina(n18266),.dinb(w_asqrt16_16[0]),.dout(n18267),.clk(gclk));
	jand g18014(.dina(w_n17819_0[1]),.dinb(n18267),.dout(n18268),.clk(gclk));
	jor g18015(.dina(n18268),.dinb(n18243),.dout(n18269),.clk(gclk));
	jor g18016(.dina(n18269),.dinb(w_asqrt17_9[0]),.dout(n18270),.clk(gclk));
	jnot g18017(.din(w_n17827_0[1]),.dout(n18271),.clk(gclk));
	jand g18018(.dina(n18271),.dinb(n18270),.dout(n18272),.clk(gclk));
	jor g18019(.dina(n18272),.dinb(n18242),.dout(n18273),.clk(gclk));
	jor g18020(.dina(n18273),.dinb(w_asqrt18_16[1]),.dout(n18274),.clk(gclk));
	jand g18021(.dina(w_n17834_0[1]),.dinb(n18274),.dout(n18275),.clk(gclk));
	jor g18022(.dina(n18275),.dinb(n18241),.dout(n18276),.clk(gclk));
	jor g18023(.dina(n18276),.dinb(w_asqrt19_9[1]),.dout(n18277),.clk(gclk));
	jnot g18024(.din(w_n17842_0[1]),.dout(n18278),.clk(gclk));
	jand g18025(.dina(n18278),.dinb(n18277),.dout(n18279),.clk(gclk));
	jor g18026(.dina(n18279),.dinb(n18240),.dout(n18280),.clk(gclk));
	jor g18027(.dina(n18280),.dinb(w_asqrt20_16[1]),.dout(n18281),.clk(gclk));
	jnot g18028(.din(w_n17849_0[1]),.dout(n18282),.clk(gclk));
	jand g18029(.dina(n18282),.dinb(n18281),.dout(n18283),.clk(gclk));
	jor g18030(.dina(n18283),.dinb(n18239),.dout(n18284),.clk(gclk));
	jor g18031(.dina(n18284),.dinb(w_asqrt21_10[0]),.dout(n18285),.clk(gclk));
	jand g18032(.dina(w_n17856_0[1]),.dinb(n18285),.dout(n18286),.clk(gclk));
	jor g18033(.dina(n18286),.dinb(n18238),.dout(n18287),.clk(gclk));
	jor g18034(.dina(n18287),.dinb(w_asqrt22_16[2]),.dout(n18288),.clk(gclk));
	jand g18035(.dina(w_n17864_0[1]),.dinb(n18288),.dout(n18289),.clk(gclk));
	jor g18036(.dina(n18289),.dinb(n18237),.dout(n18290),.clk(gclk));
	jor g18037(.dina(n18290),.dinb(w_asqrt23_10[2]),.dout(n18291),.clk(gclk));
	jnot g18038(.din(w_n17872_0[1]),.dout(n18292),.clk(gclk));
	jand g18039(.dina(n18292),.dinb(n18291),.dout(n18293),.clk(gclk));
	jor g18040(.dina(n18293),.dinb(n18236),.dout(n18294),.clk(gclk));
	jor g18041(.dina(n18294),.dinb(w_asqrt24_16[2]),.dout(n18295),.clk(gclk));
	jand g18042(.dina(w_n17879_0[1]),.dinb(n18295),.dout(n18296),.clk(gclk));
	jor g18043(.dina(n18296),.dinb(n18235),.dout(n18297),.clk(gclk));
	jor g18044(.dina(n18297),.dinb(w_asqrt25_10[2]),.dout(n18298),.clk(gclk));
	jnot g18045(.din(w_n17887_0[1]),.dout(n18299),.clk(gclk));
	jand g18046(.dina(n18299),.dinb(n18298),.dout(n18300),.clk(gclk));
	jor g18047(.dina(n18300),.dinb(n18234),.dout(n18301),.clk(gclk));
	jor g18048(.dina(n18301),.dinb(w_asqrt26_16[2]),.dout(n18302),.clk(gclk));
	jand g18049(.dina(w_n17894_0[1]),.dinb(n18302),.dout(n18303),.clk(gclk));
	jor g18050(.dina(n18303),.dinb(n18233),.dout(n18304),.clk(gclk));
	jor g18051(.dina(n18304),.dinb(w_asqrt27_11[1]),.dout(n18305),.clk(gclk));
	jnot g18052(.din(w_n17902_0[1]),.dout(n18306),.clk(gclk));
	jand g18053(.dina(n18306),.dinb(n18305),.dout(n18307),.clk(gclk));
	jor g18054(.dina(n18307),.dinb(n18232),.dout(n18308),.clk(gclk));
	jor g18055(.dina(n18308),.dinb(w_asqrt28_17[0]),.dout(n18309),.clk(gclk));
	jnot g18056(.din(w_n17909_0[1]),.dout(n18310),.clk(gclk));
	jand g18057(.dina(n18310),.dinb(n18309),.dout(n18311),.clk(gclk));
	jor g18058(.dina(n18311),.dinb(n18231),.dout(n18312),.clk(gclk));
	jor g18059(.dina(n18312),.dinb(w_asqrt29_11[2]),.dout(n18313),.clk(gclk));
	jnot g18060(.din(w_n17916_0[1]),.dout(n18314),.clk(gclk));
	jand g18061(.dina(n18314),.dinb(n18313),.dout(n18315),.clk(gclk));
	jor g18062(.dina(n18315),.dinb(n18230),.dout(n18316),.clk(gclk));
	jor g18063(.dina(n18316),.dinb(w_asqrt30_17[1]),.dout(n18317),.clk(gclk));
	jand g18064(.dina(w_n17923_0[1]),.dinb(n18317),.dout(n18318),.clk(gclk));
	jor g18065(.dina(n18318),.dinb(n18229),.dout(n18319),.clk(gclk));
	jor g18066(.dina(n18319),.dinb(w_asqrt31_12[1]),.dout(n18320),.clk(gclk));
	jnot g18067(.din(w_n17931_0[1]),.dout(n18321),.clk(gclk));
	jand g18068(.dina(n18321),.dinb(n18320),.dout(n18322),.clk(gclk));
	jor g18069(.dina(n18322),.dinb(n18228),.dout(n18323),.clk(gclk));
	jor g18070(.dina(n18323),.dinb(w_asqrt32_17[1]),.dout(n18324),.clk(gclk));
	jand g18071(.dina(w_n17938_0[1]),.dinb(n18324),.dout(n18325),.clk(gclk));
	jor g18072(.dina(n18325),.dinb(n18227),.dout(n18326),.clk(gclk));
	jor g18073(.dina(n18326),.dinb(w_asqrt33_13[0]),.dout(n18327),.clk(gclk));
	jnot g18074(.din(w_n17946_0[1]),.dout(n18328),.clk(gclk));
	jand g18075(.dina(n18328),.dinb(n18327),.dout(n18329),.clk(gclk));
	jor g18076(.dina(n18329),.dinb(n18226),.dout(n18330),.clk(gclk));
	jor g18077(.dina(n18330),.dinb(w_asqrt34_17[2]),.dout(n18331),.clk(gclk));
	jand g18078(.dina(w_n17953_0[1]),.dinb(n18331),.dout(n18332),.clk(gclk));
	jor g18079(.dina(n18332),.dinb(n18225),.dout(n18333),.clk(gclk));
	jor g18080(.dina(n18333),.dinb(w_asqrt35_13[2]),.dout(n18334),.clk(gclk));
	jnot g18081(.din(w_n17961_0[1]),.dout(n18335),.clk(gclk));
	jand g18082(.dina(n18335),.dinb(n18334),.dout(n18336),.clk(gclk));
	jor g18083(.dina(n18336),.dinb(n18224),.dout(n18337),.clk(gclk));
	jor g18084(.dina(n18337),.dinb(w_asqrt36_17[2]),.dout(n18338),.clk(gclk));
	jand g18085(.dina(w_n17968_0[1]),.dinb(n18338),.dout(n18339),.clk(gclk));
	jor g18086(.dina(n18339),.dinb(n18223),.dout(n18340),.clk(gclk));
	jor g18087(.dina(n18340),.dinb(w_asqrt37_14[0]),.dout(n18341),.clk(gclk));
	jnot g18088(.din(w_n17976_0[1]),.dout(n18342),.clk(gclk));
	jand g18089(.dina(n18342),.dinb(n18341),.dout(n18343),.clk(gclk));
	jor g18090(.dina(n18343),.dinb(n18222),.dout(n18344),.clk(gclk));
	jor g18091(.dina(n18344),.dinb(w_asqrt38_18[0]),.dout(n18345),.clk(gclk));
	jnot g18092(.din(w_n17983_0[1]),.dout(n18346),.clk(gclk));
	jand g18093(.dina(n18346),.dinb(n18345),.dout(n18347),.clk(gclk));
	jor g18094(.dina(n18347),.dinb(n18221),.dout(n18348),.clk(gclk));
	jor g18095(.dina(n18348),.dinb(w_asqrt39_14[2]),.dout(n18349),.clk(gclk));
	jnot g18096(.din(w_n17990_0[1]),.dout(n18350),.clk(gclk));
	jand g18097(.dina(n18350),.dinb(n18349),.dout(n18351),.clk(gclk));
	jor g18098(.dina(n18351),.dinb(n18220),.dout(n18352),.clk(gclk));
	jor g18099(.dina(n18352),.dinb(w_asqrt40_18[0]),.dout(n18353),.clk(gclk));
	jand g18100(.dina(w_n17997_0[1]),.dinb(n18353),.dout(n18354),.clk(gclk));
	jor g18101(.dina(n18354),.dinb(n18219),.dout(n18355),.clk(gclk));
	jor g18102(.dina(n18355),.dinb(w_asqrt41_15[0]),.dout(n18356),.clk(gclk));
	jnot g18103(.din(w_n18005_0[1]),.dout(n18357),.clk(gclk));
	jand g18104(.dina(n18357),.dinb(n18356),.dout(n18358),.clk(gclk));
	jor g18105(.dina(n18358),.dinb(n18218),.dout(n18359),.clk(gclk));
	jor g18106(.dina(n18359),.dinb(w_asqrt42_18[1]),.dout(n18360),.clk(gclk));
	jand g18107(.dina(w_n18012_0[0]),.dinb(n18360),.dout(n18361),.clk(gclk));
	jor g18108(.dina(n18361),.dinb(n18217),.dout(n18362),.clk(gclk));
	jor g18109(.dina(n18362),.dinb(w_asqrt43_15[1]),.dout(n18363),.clk(gclk));
	jnot g18110(.din(w_n18020_0[1]),.dout(n18364),.clk(gclk));
	jand g18111(.dina(n18364),.dinb(n18363),.dout(n18365),.clk(gclk));
	jor g18112(.dina(n18365),.dinb(n18216),.dout(n18366),.clk(gclk));
	jor g18113(.dina(n18366),.dinb(w_asqrt44_18[1]),.dout(n18367),.clk(gclk));
	jnot g18114(.din(w_n18027_0[1]),.dout(n18368),.clk(gclk));
	jand g18115(.dina(n18368),.dinb(n18367),.dout(n18369),.clk(gclk));
	jor g18116(.dina(n18369),.dinb(n18215),.dout(n18370),.clk(gclk));
	jor g18117(.dina(n18370),.dinb(w_asqrt45_16[0]),.dout(n18371),.clk(gclk));
	jnot g18118(.din(w_n18034_0[1]),.dout(n18372),.clk(gclk));
	jand g18119(.dina(n18372),.dinb(n18371),.dout(n18373),.clk(gclk));
	jor g18120(.dina(n18373),.dinb(n18214),.dout(n18374),.clk(gclk));
	jor g18121(.dina(n18374),.dinb(w_asqrt46_18[1]),.dout(n18375),.clk(gclk));
	jand g18122(.dina(w_n18041_0[1]),.dinb(n18375),.dout(n18376),.clk(gclk));
	jor g18123(.dina(n18376),.dinb(n18213),.dout(n18377),.clk(gclk));
	jor g18124(.dina(n18377),.dinb(w_asqrt47_16[2]),.dout(n18378),.clk(gclk));
	jnot g18125(.din(w_n18049_0[1]),.dout(n18379),.clk(gclk));
	jand g18126(.dina(n18379),.dinb(n18378),.dout(n18380),.clk(gclk));
	jor g18127(.dina(n18380),.dinb(n18212),.dout(n18381),.clk(gclk));
	jor g18128(.dina(n18381),.dinb(w_asqrt48_18[2]),.dout(n18382),.clk(gclk));
	jand g18129(.dina(w_n18056_0[1]),.dinb(n18382),.dout(n18383),.clk(gclk));
	jor g18130(.dina(n18383),.dinb(n18211),.dout(n18384),.clk(gclk));
	jor g18131(.dina(n18384),.dinb(w_asqrt49_17[0]),.dout(n18385),.clk(gclk));
	jnot g18132(.din(w_n18064_0[1]),.dout(n18386),.clk(gclk));
	jand g18133(.dina(n18386),.dinb(n18385),.dout(n18387),.clk(gclk));
	jor g18134(.dina(n18387),.dinb(n18210),.dout(n18388),.clk(gclk));
	jor g18135(.dina(n18388),.dinb(w_asqrt50_19[0]),.dout(n18389),.clk(gclk));
	jnot g18136(.din(w_n18071_0[1]),.dout(n18390),.clk(gclk));
	jand g18137(.dina(n18390),.dinb(n18389),.dout(n18391),.clk(gclk));
	jor g18138(.dina(n18391),.dinb(n18209),.dout(n18392),.clk(gclk));
	jor g18139(.dina(n18392),.dinb(w_asqrt51_17[1]),.dout(n18393),.clk(gclk));
	jand g18140(.dina(w_n18078_0[1]),.dinb(n18393),.dout(n18394),.clk(gclk));
	jor g18141(.dina(n18394),.dinb(n18208),.dout(n18395),.clk(gclk));
	jor g18142(.dina(n18395),.dinb(w_asqrt52_19[0]),.dout(n18396),.clk(gclk));
	jand g18143(.dina(n18396),.dinb(w_n18085_0[1]),.dout(n18397),.clk(gclk));
	jor g18144(.dina(n18397),.dinb(n18207),.dout(n18398),.clk(gclk));
	jor g18145(.dina(n18398),.dinb(w_asqrt53_18[0]),.dout(n18399),.clk(gclk));
	jnot g18146(.din(w_n18094_0[1]),.dout(n18400),.clk(gclk));
	jand g18147(.dina(n18400),.dinb(n18399),.dout(n18401),.clk(gclk));
	jor g18148(.dina(n18401),.dinb(n18206),.dout(n18402),.clk(gclk));
	jor g18149(.dina(n18402),.dinb(w_asqrt54_19[0]),.dout(n18403),.clk(gclk));
	jand g18150(.dina(w_n18101_0[1]),.dinb(n18403),.dout(n18404),.clk(gclk));
	jor g18151(.dina(n18404),.dinb(n18205),.dout(n18405),.clk(gclk));
	jor g18152(.dina(n18405),.dinb(w_asqrt55_18[1]),.dout(n18406),.clk(gclk));
	jnot g18153(.din(w_n18109_0[1]),.dout(n18407),.clk(gclk));
	jand g18154(.dina(n18407),.dinb(n18406),.dout(n18408),.clk(gclk));
	jor g18155(.dina(n18408),.dinb(n18204),.dout(n18409),.clk(gclk));
	jor g18156(.dina(n18409),.dinb(w_asqrt56_19[1]),.dout(n18410),.clk(gclk));
	jand g18157(.dina(w_n18116_0[1]),.dinb(n18410),.dout(n18411),.clk(gclk));
	jor g18158(.dina(n18411),.dinb(n18203),.dout(n18412),.clk(gclk));
	jor g18159(.dina(n18412),.dinb(w_asqrt57_19[0]),.dout(n18413),.clk(gclk));
	jnot g18160(.din(w_n18124_0[1]),.dout(n18414),.clk(gclk));
	jand g18161(.dina(n18414),.dinb(n18413),.dout(n18415),.clk(gclk));
	jor g18162(.dina(n18415),.dinb(n18202),.dout(n18416),.clk(gclk));
	jor g18163(.dina(n18416),.dinb(w_asqrt58_19[2]),.dout(n18417),.clk(gclk));
	jnot g18164(.din(w_n18131_0[1]),.dout(n18418),.clk(gclk));
	jand g18165(.dina(n18418),.dinb(n18417),.dout(n18419),.clk(gclk));
	jor g18166(.dina(n18419),.dinb(n18201),.dout(n18420),.clk(gclk));
	jor g18167(.dina(n18420),.dinb(w_asqrt59_19[1]),.dout(n18421),.clk(gclk));
	jnot g18168(.din(w_n18138_0[1]),.dout(n18422),.clk(gclk));
	jand g18169(.dina(n18422),.dinb(n18421),.dout(n18423),.clk(gclk));
	jor g18170(.dina(n18423),.dinb(n18200),.dout(n18424),.clk(gclk));
	jor g18171(.dina(n18424),.dinb(w_asqrt60_19[2]),.dout(n18425),.clk(gclk));
	jand g18172(.dina(w_n18145_0[1]),.dinb(n18425),.dout(n18426),.clk(gclk));
	jor g18173(.dina(n18426),.dinb(n18199),.dout(n18427),.clk(gclk));
	jor g18174(.dina(n18427),.dinb(w_asqrt61_19[2]),.dout(n18428),.clk(gclk));
	jnot g18175(.din(w_n18153_0[1]),.dout(n18429),.clk(gclk));
	jand g18176(.dina(n18429),.dinb(n18428),.dout(n18430),.clk(gclk));
	jor g18177(.dina(n18430),.dinb(n18198),.dout(n18431),.clk(gclk));
	jor g18178(.dina(n18431),.dinb(w_asqrt62_19[2]),.dout(n18432),.clk(gclk));
	jand g18179(.dina(w_n18160_0[0]),.dinb(n18432),.dout(n18433),.clk(gclk));
	jor g18180(.dina(n18433),.dinb(n18197),.dout(n18434),.clk(gclk));
	jand g18181(.dina(n18434),.dinb(w_n17772_0[0]),.dout(n18435),.clk(gclk));
	jand g18182(.dina(w_n18435_0[1]),.dinb(w_n17518_0[1]),.dout(n18436),.clk(gclk));
	jand g18183(.dina(n18436),.dinb(n18196),.dout(n18437),.clk(gclk));
	jor g18184(.dina(n18437),.dinb(w_asqrt63_24[1]),.dout(n18438),.clk(gclk));
	jnot g18185(.din(w_n18176_0[0]),.dout(n18439),.clk(gclk));
	jand g18186(.dina(n18439),.dinb(w_n18438_0[1]),.dout(n18440),.clk(gclk));
	jand g18187(.dina(n18440),.dinb(w_n18169_0[0]),.dout(n18441),.clk(gclk));
	jand g18188(.dina(w_n18441_0[1]),.dinb(w_n18195_0[2]),.dout(n18442),.clk(gclk));
	jor g18189(.dina(w_n18442_12[2]),.dinb(n18194),.dout(n18443),.clk(gclk));
	jand g18190(.dina(n18443),.dinb(n18193),.dout(n18444),.clk(gclk));
	jand g18191(.dina(n18444),.dinb(n18191),.dout(n18445),.clk(gclk));
	jor g18192(.dina(n18445),.dinb(w_n18190_0[1]),.dout(n18446),.clk(gclk));
	jand g18193(.dina(w_n18446_0[2]),.dinb(w_asqrt12_15[1]),.dout(n18447),.clk(gclk));
	jor g18194(.dina(w_n18446_0[1]),.dinb(w_asqrt12_15[0]),.dout(n18448),.clk(gclk));
	jand g18195(.dina(w_asqrt10_31[1]),.dinb(w_n17776_0[0]),.dout(n18449),.clk(gclk));
	jand g18196(.dina(w_n18195_0[1]),.dinb(w_asqrt11_6[2]),.dout(n18450),.clk(gclk));
	jand g18197(.dina(n18450),.dinb(w_n18438_0[0]),.dout(n18451),.clk(gclk));
	jand g18198(.dina(n18451),.dinb(w_n18168_0[0]),.dout(n18452),.clk(gclk));
	jor g18199(.dina(n18452),.dinb(w_n18449_0[1]),.dout(n18453),.clk(gclk));
	jxor g18200(.dina(n18453),.dinb(w_a22_0[1]),.dout(n18454),.clk(gclk));
	jnot g18201(.din(w_n18454_0[1]),.dout(n18455),.clk(gclk));
	jand g18202(.dina(w_n18455_0[1]),.dinb(n18448),.dout(n18456),.clk(gclk));
	jor g18203(.dina(n18456),.dinb(w_n18447_0[1]),.dout(n18457),.clk(gclk));
	jand g18204(.dina(w_n18457_0[2]),.dinb(w_asqrt13_7[2]),.dout(n18458),.clk(gclk));
	jor g18205(.dina(w_n18457_0[1]),.dinb(w_asqrt13_7[1]),.dout(n18459),.clk(gclk));
	jxor g18206(.dina(w_n17780_0[0]),.dinb(w_n17134_13[0]),.dout(n18460),.clk(gclk));
	jand g18207(.dina(n18460),.dinb(w_asqrt10_31[0]),.dout(n18461),.clk(gclk));
	jxor g18208(.dina(n18461),.dinb(w_n18253_0[0]),.dout(n18462),.clk(gclk));
	jand g18209(.dina(w_n18462_0[1]),.dinb(n18459),.dout(n18463),.clk(gclk));
	jor g18210(.dina(n18463),.dinb(w_n18458_0[1]),.dout(n18464),.clk(gclk));
	jand g18211(.dina(w_n18464_0[2]),.dinb(w_asqrt14_15[2]),.dout(n18465),.clk(gclk));
	jor g18212(.dina(w_n18464_0[1]),.dinb(w_asqrt14_15[1]),.dout(n18466),.clk(gclk));
	jxor g18213(.dina(w_n17788_0[0]),.dinb(w_n16489_21[0]),.dout(n18467),.clk(gclk));
	jand g18214(.dina(n18467),.dinb(w_asqrt10_30[2]),.dout(n18468),.clk(gclk));
	jxor g18215(.dina(n18468),.dinb(w_n17797_0[0]),.dout(n18469),.clk(gclk));
	jnot g18216(.din(w_n18469_0[1]),.dout(n18470),.clk(gclk));
	jand g18217(.dina(w_n18470_0[1]),.dinb(n18466),.dout(n18471),.clk(gclk));
	jor g18218(.dina(n18471),.dinb(w_n18465_0[1]),.dout(n18472),.clk(gclk));
	jand g18219(.dina(w_n18472_0[2]),.dinb(w_asqrt15_8[1]),.dout(n18473),.clk(gclk));
	jor g18220(.dina(w_n18472_0[1]),.dinb(w_asqrt15_8[0]),.dout(n18474),.clk(gclk));
	jxor g18221(.dina(w_n17799_0[0]),.dinb(w_n15878_14[0]),.dout(n18475),.clk(gclk));
	jand g18222(.dina(n18475),.dinb(w_asqrt10_30[1]),.dout(n18476),.clk(gclk));
	jxor g18223(.dina(n18476),.dinb(w_n17804_0[0]),.dout(n18477),.clk(gclk));
	jand g18224(.dina(w_n18477_0[1]),.dinb(n18474),.dout(n18478),.clk(gclk));
	jor g18225(.dina(n18478),.dinb(w_n18473_0[1]),.dout(n18479),.clk(gclk));
	jand g18226(.dina(w_n18479_0[2]),.dinb(w_asqrt16_15[2]),.dout(n18480),.clk(gclk));
	jor g18227(.dina(w_n18479_0[1]),.dinb(w_asqrt16_15[1]),.dout(n18481),.clk(gclk));
	jxor g18228(.dina(w_n17807_0[0]),.dinb(w_n15260_21[2]),.dout(n18482),.clk(gclk));
	jand g18229(.dina(n18482),.dinb(w_asqrt10_30[0]),.dout(n18483),.clk(gclk));
	jxor g18230(.dina(n18483),.dinb(w_n17812_0[0]),.dout(n18484),.clk(gclk));
	jnot g18231(.din(w_n18484_0[1]),.dout(n18485),.clk(gclk));
	jand g18232(.dina(w_n18485_0[1]),.dinb(n18481),.dout(n18486),.clk(gclk));
	jor g18233(.dina(n18486),.dinb(w_n18480_0[1]),.dout(n18487),.clk(gclk));
	jand g18234(.dina(w_n18487_0[2]),.dinb(w_asqrt17_8[2]),.dout(n18488),.clk(gclk));
	jor g18235(.dina(w_n18487_0[1]),.dinb(w_asqrt17_8[1]),.dout(n18489),.clk(gclk));
	jxor g18236(.dina(w_n17814_0[0]),.dinb(w_n14674_14[2]),.dout(n18490),.clk(gclk));
	jand g18237(.dina(n18490),.dinb(w_asqrt10_29[2]),.dout(n18491),.clk(gclk));
	jxor g18238(.dina(n18491),.dinb(w_n17819_0[0]),.dout(n18492),.clk(gclk));
	jand g18239(.dina(w_n18492_0[1]),.dinb(n18489),.dout(n18493),.clk(gclk));
	jor g18240(.dina(n18493),.dinb(w_n18488_0[1]),.dout(n18494),.clk(gclk));
	jand g18241(.dina(w_n18494_0[2]),.dinb(w_asqrt18_16[0]),.dout(n18495),.clk(gclk));
	jor g18242(.dina(w_n18494_0[1]),.dinb(w_asqrt18_15[2]),.dout(n18496),.clk(gclk));
	jxor g18243(.dina(w_n17822_0[0]),.dinb(w_n14078_22[0]),.dout(n18497),.clk(gclk));
	jand g18244(.dina(n18497),.dinb(w_asqrt10_29[1]),.dout(n18498),.clk(gclk));
	jxor g18245(.dina(n18498),.dinb(w_n17827_0[0]),.dout(n18499),.clk(gclk));
	jnot g18246(.din(w_n18499_0[1]),.dout(n18500),.clk(gclk));
	jand g18247(.dina(w_n18500_0[1]),.dinb(n18496),.dout(n18501),.clk(gclk));
	jor g18248(.dina(n18501),.dinb(w_n18495_0[1]),.dout(n18502),.clk(gclk));
	jand g18249(.dina(w_n18502_0[2]),.dinb(w_asqrt19_9[0]),.dout(n18503),.clk(gclk));
	jor g18250(.dina(w_n18502_0[1]),.dinb(w_asqrt19_8[2]),.dout(n18504),.clk(gclk));
	jxor g18251(.dina(w_n17829_0[0]),.dinb(w_n13515_15[2]),.dout(n18505),.clk(gclk));
	jand g18252(.dina(n18505),.dinb(w_asqrt10_29[0]),.dout(n18506),.clk(gclk));
	jxor g18253(.dina(n18506),.dinb(w_n17834_0[0]),.dout(n18507),.clk(gclk));
	jand g18254(.dina(w_n18507_0[1]),.dinb(n18504),.dout(n18508),.clk(gclk));
	jor g18255(.dina(n18508),.dinb(w_n18503_0[1]),.dout(n18509),.clk(gclk));
	jand g18256(.dina(w_n18509_0[2]),.dinb(w_asqrt20_16[0]),.dout(n18510),.clk(gclk));
	jor g18257(.dina(w_n18509_0[1]),.dinb(w_asqrt20_15[2]),.dout(n18511),.clk(gclk));
	jxor g18258(.dina(w_n17837_0[0]),.dinb(w_n12947_22[2]),.dout(n18512),.clk(gclk));
	jand g18259(.dina(n18512),.dinb(w_asqrt10_28[2]),.dout(n18513),.clk(gclk));
	jxor g18260(.dina(n18513),.dinb(w_n17842_0[0]),.dout(n18514),.clk(gclk));
	jnot g18261(.din(w_n18514_0[1]),.dout(n18515),.clk(gclk));
	jand g18262(.dina(w_n18515_0[1]),.dinb(n18511),.dout(n18516),.clk(gclk));
	jor g18263(.dina(n18516),.dinb(w_n18510_0[1]),.dout(n18517),.clk(gclk));
	jand g18264(.dina(w_n18517_0[2]),.dinb(w_asqrt21_9[2]),.dout(n18518),.clk(gclk));
	jor g18265(.dina(w_n18517_0[1]),.dinb(w_asqrt21_9[1]),.dout(n18519),.clk(gclk));
	jxor g18266(.dina(w_n17844_0[0]),.dinb(w_n12410_16[1]),.dout(n18520),.clk(gclk));
	jand g18267(.dina(n18520),.dinb(w_asqrt10_28[1]),.dout(n18521),.clk(gclk));
	jxor g18268(.dina(n18521),.dinb(w_n17849_0[0]),.dout(n18522),.clk(gclk));
	jnot g18269(.din(w_n18522_0[1]),.dout(n18523),.clk(gclk));
	jand g18270(.dina(w_n18523_0[1]),.dinb(n18519),.dout(n18524),.clk(gclk));
	jor g18271(.dina(n18524),.dinb(w_n18518_0[1]),.dout(n18525),.clk(gclk));
	jand g18272(.dina(w_n18525_0[2]),.dinb(w_asqrt22_16[1]),.dout(n18526),.clk(gclk));
	jor g18273(.dina(w_n18525_0[1]),.dinb(w_asqrt22_16[0]),.dout(n18527),.clk(gclk));
	jxor g18274(.dina(w_n17851_0[0]),.dinb(w_n11858_23[0]),.dout(n18528),.clk(gclk));
	jand g18275(.dina(n18528),.dinb(w_asqrt10_28[0]),.dout(n18529),.clk(gclk));
	jxor g18276(.dina(n18529),.dinb(w_n17856_0[0]),.dout(n18530),.clk(gclk));
	jand g18277(.dina(w_n18530_0[1]),.dinb(n18527),.dout(n18531),.clk(gclk));
	jor g18278(.dina(n18531),.dinb(w_n18526_0[1]),.dout(n18532),.clk(gclk));
	jand g18279(.dina(w_n18532_0[2]),.dinb(w_asqrt23_10[1]),.dout(n18533),.clk(gclk));
	jor g18280(.dina(w_n18532_0[1]),.dinb(w_asqrt23_10[0]),.dout(n18534),.clk(gclk));
	jxor g18281(.dina(w_n17859_0[0]),.dinb(w_n11347_17[0]),.dout(n18535),.clk(gclk));
	jand g18282(.dina(n18535),.dinb(w_asqrt10_27[2]),.dout(n18536),.clk(gclk));
	jxor g18283(.dina(n18536),.dinb(w_n17864_0[0]),.dout(n18537),.clk(gclk));
	jand g18284(.dina(w_n18537_0[1]),.dinb(n18534),.dout(n18538),.clk(gclk));
	jor g18285(.dina(n18538),.dinb(w_n18533_0[1]),.dout(n18539),.clk(gclk));
	jand g18286(.dina(w_n18539_0[2]),.dinb(w_asqrt24_16[1]),.dout(n18540),.clk(gclk));
	jor g18287(.dina(w_n18539_0[1]),.dinb(w_asqrt24_16[0]),.dout(n18541),.clk(gclk));
	jxor g18288(.dina(w_n17867_0[0]),.dinb(w_n10824_23[2]),.dout(n18542),.clk(gclk));
	jand g18289(.dina(n18542),.dinb(w_asqrt10_27[1]),.dout(n18543),.clk(gclk));
	jxor g18290(.dina(n18543),.dinb(w_n17872_0[0]),.dout(n18544),.clk(gclk));
	jnot g18291(.din(w_n18544_0[1]),.dout(n18545),.clk(gclk));
	jand g18292(.dina(w_n18545_0[1]),.dinb(n18541),.dout(n18546),.clk(gclk));
	jor g18293(.dina(n18546),.dinb(w_n18540_0[1]),.dout(n18547),.clk(gclk));
	jand g18294(.dina(w_n18547_0[2]),.dinb(w_asqrt25_10[1]),.dout(n18548),.clk(gclk));
	jor g18295(.dina(w_n18547_0[1]),.dinb(w_asqrt25_10[0]),.dout(n18549),.clk(gclk));
	jxor g18296(.dina(w_n17874_0[0]),.dinb(w_n10328_18[0]),.dout(n18550),.clk(gclk));
	jand g18297(.dina(n18550),.dinb(w_asqrt10_27[0]),.dout(n18551),.clk(gclk));
	jxor g18298(.dina(n18551),.dinb(w_n17879_0[0]),.dout(n18552),.clk(gclk));
	jand g18299(.dina(w_n18552_0[1]),.dinb(n18549),.dout(n18553),.clk(gclk));
	jor g18300(.dina(n18553),.dinb(w_n18548_0[1]),.dout(n18554),.clk(gclk));
	jand g18301(.dina(w_n18554_0[2]),.dinb(w_asqrt26_16[1]),.dout(n18555),.clk(gclk));
	jor g18302(.dina(w_n18554_0[1]),.dinb(w_asqrt26_16[0]),.dout(n18556),.clk(gclk));
	jxor g18303(.dina(w_n17882_0[0]),.dinb(w_n9832_24[1]),.dout(n18557),.clk(gclk));
	jand g18304(.dina(n18557),.dinb(w_asqrt10_26[2]),.dout(n18558),.clk(gclk));
	jxor g18305(.dina(n18558),.dinb(w_n17887_0[0]),.dout(n18559),.clk(gclk));
	jnot g18306(.din(w_n18559_0[1]),.dout(n18560),.clk(gclk));
	jand g18307(.dina(w_n18560_0[1]),.dinb(n18556),.dout(n18561),.clk(gclk));
	jor g18308(.dina(n18561),.dinb(w_n18555_0[1]),.dout(n18562),.clk(gclk));
	jand g18309(.dina(w_n18562_0[2]),.dinb(w_asqrt27_11[0]),.dout(n18563),.clk(gclk));
	jor g18310(.dina(w_n18562_0[1]),.dinb(w_asqrt27_10[2]),.dout(n18564),.clk(gclk));
	jxor g18311(.dina(w_n17889_0[0]),.dinb(w_n9369_19[0]),.dout(n18565),.clk(gclk));
	jand g18312(.dina(n18565),.dinb(w_asqrt10_26[1]),.dout(n18566),.clk(gclk));
	jxor g18313(.dina(n18566),.dinb(w_n17894_0[0]),.dout(n18567),.clk(gclk));
	jand g18314(.dina(w_n18567_0[1]),.dinb(n18564),.dout(n18568),.clk(gclk));
	jor g18315(.dina(n18568),.dinb(w_n18563_0[1]),.dout(n18569),.clk(gclk));
	jand g18316(.dina(w_n18569_0[2]),.dinb(w_asqrt28_16[2]),.dout(n18570),.clk(gclk));
	jor g18317(.dina(w_n18569_0[1]),.dinb(w_asqrt28_16[1]),.dout(n18571),.clk(gclk));
	jxor g18318(.dina(w_n17897_0[0]),.dinb(w_n8890_24[2]),.dout(n18572),.clk(gclk));
	jand g18319(.dina(n18572),.dinb(w_asqrt10_26[0]),.dout(n18573),.clk(gclk));
	jxor g18320(.dina(n18573),.dinb(w_n17902_0[0]),.dout(n18574),.clk(gclk));
	jnot g18321(.din(w_n18574_0[1]),.dout(n18575),.clk(gclk));
	jand g18322(.dina(w_n18575_0[1]),.dinb(n18571),.dout(n18576),.clk(gclk));
	jor g18323(.dina(n18576),.dinb(w_n18570_0[1]),.dout(n18577),.clk(gclk));
	jand g18324(.dina(w_n18577_0[2]),.dinb(w_asqrt29_11[1]),.dout(n18578),.clk(gclk));
	jor g18325(.dina(w_n18577_0[1]),.dinb(w_asqrt29_11[0]),.dout(n18579),.clk(gclk));
	jxor g18326(.dina(w_n17904_0[0]),.dinb(w_n8449_19[2]),.dout(n18580),.clk(gclk));
	jand g18327(.dina(n18580),.dinb(w_asqrt10_25[2]),.dout(n18581),.clk(gclk));
	jxor g18328(.dina(n18581),.dinb(w_n17909_0[0]),.dout(n18582),.clk(gclk));
	jnot g18329(.din(w_n18582_0[1]),.dout(n18583),.clk(gclk));
	jand g18330(.dina(w_n18583_0[1]),.dinb(n18579),.dout(n18584),.clk(gclk));
	jor g18331(.dina(n18584),.dinb(w_n18578_0[1]),.dout(n18585),.clk(gclk));
	jand g18332(.dina(w_n18585_0[2]),.dinb(w_asqrt30_17[0]),.dout(n18586),.clk(gclk));
	jor g18333(.dina(w_n18585_0[1]),.dinb(w_asqrt30_16[2]),.dout(n18587),.clk(gclk));
	jxor g18334(.dina(w_n17911_0[0]),.dinb(w_n8003_25[1]),.dout(n18588),.clk(gclk));
	jand g18335(.dina(n18588),.dinb(w_asqrt10_25[1]),.dout(n18589),.clk(gclk));
	jxor g18336(.dina(n18589),.dinb(w_n17916_0[0]),.dout(n18590),.clk(gclk));
	jnot g18337(.din(w_n18590_0[1]),.dout(n18591),.clk(gclk));
	jand g18338(.dina(w_n18591_0[1]),.dinb(n18587),.dout(n18592),.clk(gclk));
	jor g18339(.dina(n18592),.dinb(w_n18586_0[1]),.dout(n18593),.clk(gclk));
	jand g18340(.dina(w_n18593_0[2]),.dinb(w_asqrt31_12[0]),.dout(n18594),.clk(gclk));
	jor g18341(.dina(w_n18593_0[1]),.dinb(w_asqrt31_11[2]),.dout(n18595),.clk(gclk));
	jxor g18342(.dina(w_n17918_0[0]),.dinb(w_n7581_20[2]),.dout(n18596),.clk(gclk));
	jand g18343(.dina(n18596),.dinb(w_asqrt10_25[0]),.dout(n18597),.clk(gclk));
	jxor g18344(.dina(n18597),.dinb(w_n17923_0[0]),.dout(n18598),.clk(gclk));
	jand g18345(.dina(w_n18598_0[1]),.dinb(n18595),.dout(n18599),.clk(gclk));
	jor g18346(.dina(n18599),.dinb(w_n18594_0[1]),.dout(n18600),.clk(gclk));
	jand g18347(.dina(w_n18600_0[2]),.dinb(w_asqrt32_17[0]),.dout(n18601),.clk(gclk));
	jor g18348(.dina(w_n18600_0[1]),.dinb(w_asqrt32_16[2]),.dout(n18602),.clk(gclk));
	jxor g18349(.dina(w_n17926_0[0]),.dinb(w_n7154_25[2]),.dout(n18603),.clk(gclk));
	jand g18350(.dina(n18603),.dinb(w_asqrt10_24[2]),.dout(n18604),.clk(gclk));
	jxor g18351(.dina(n18604),.dinb(w_n17931_0[0]),.dout(n18605),.clk(gclk));
	jnot g18352(.din(w_n18605_0[1]),.dout(n18606),.clk(gclk));
	jand g18353(.dina(w_n18606_0[1]),.dinb(n18602),.dout(n18607),.clk(gclk));
	jor g18354(.dina(n18607),.dinb(w_n18601_0[1]),.dout(n18608),.clk(gclk));
	jand g18355(.dina(w_n18608_0[2]),.dinb(w_asqrt33_12[2]),.dout(n18609),.clk(gclk));
	jor g18356(.dina(w_n18608_0[1]),.dinb(w_asqrt33_12[1]),.dout(n18610),.clk(gclk));
	jxor g18357(.dina(w_n17933_0[0]),.dinb(w_n6758_21[1]),.dout(n18611),.clk(gclk));
	jand g18358(.dina(n18611),.dinb(w_asqrt10_24[1]),.dout(n18612),.clk(gclk));
	jxor g18359(.dina(n18612),.dinb(w_n17938_0[0]),.dout(n18613),.clk(gclk));
	jand g18360(.dina(w_n18613_0[1]),.dinb(n18610),.dout(n18614),.clk(gclk));
	jor g18361(.dina(n18614),.dinb(w_n18609_0[1]),.dout(n18615),.clk(gclk));
	jand g18362(.dina(w_n18615_0[2]),.dinb(w_asqrt34_17[1]),.dout(n18616),.clk(gclk));
	jor g18363(.dina(w_n18615_0[1]),.dinb(w_asqrt34_17[0]),.dout(n18617),.clk(gclk));
	jxor g18364(.dina(w_n17941_0[0]),.dinb(w_n6357_26[0]),.dout(n18618),.clk(gclk));
	jand g18365(.dina(n18618),.dinb(w_asqrt10_24[0]),.dout(n18619),.clk(gclk));
	jxor g18366(.dina(n18619),.dinb(w_n17946_0[0]),.dout(n18620),.clk(gclk));
	jnot g18367(.din(w_n18620_0[1]),.dout(n18621),.clk(gclk));
	jand g18368(.dina(w_n18621_0[1]),.dinb(n18617),.dout(n18622),.clk(gclk));
	jor g18369(.dina(n18622),.dinb(w_n18616_0[1]),.dout(n18623),.clk(gclk));
	jand g18370(.dina(w_n18623_0[2]),.dinb(w_asqrt35_13[1]),.dout(n18624),.clk(gclk));
	jor g18371(.dina(w_n18623_0[1]),.dinb(w_asqrt35_13[0]),.dout(n18625),.clk(gclk));
	jxor g18372(.dina(w_n17948_0[0]),.dinb(w_n5989_22[0]),.dout(n18626),.clk(gclk));
	jand g18373(.dina(n18626),.dinb(w_asqrt10_23[2]),.dout(n18627),.clk(gclk));
	jxor g18374(.dina(n18627),.dinb(w_n17953_0[0]),.dout(n18628),.clk(gclk));
	jand g18375(.dina(w_n18628_0[1]),.dinb(n18625),.dout(n18629),.clk(gclk));
	jor g18376(.dina(n18629),.dinb(w_n18624_0[1]),.dout(n18630),.clk(gclk));
	jand g18377(.dina(w_n18630_0[2]),.dinb(w_asqrt36_17[1]),.dout(n18631),.clk(gclk));
	jor g18378(.dina(w_n18630_0[1]),.dinb(w_asqrt36_17[0]),.dout(n18632),.clk(gclk));
	jxor g18379(.dina(w_n17956_0[0]),.dinb(w_n5606_26[1]),.dout(n18633),.clk(gclk));
	jand g18380(.dina(n18633),.dinb(w_asqrt10_23[1]),.dout(n18634),.clk(gclk));
	jxor g18381(.dina(n18634),.dinb(w_n17961_0[0]),.dout(n18635),.clk(gclk));
	jnot g18382(.din(w_n18635_0[1]),.dout(n18636),.clk(gclk));
	jand g18383(.dina(w_n18636_0[1]),.dinb(n18632),.dout(n18637),.clk(gclk));
	jor g18384(.dina(n18637),.dinb(w_n18631_0[1]),.dout(n18638),.clk(gclk));
	jand g18385(.dina(w_n18638_0[2]),.dinb(w_asqrt37_13[2]),.dout(n18639),.clk(gclk));
	jor g18386(.dina(w_n18638_0[1]),.dinb(w_asqrt37_13[1]),.dout(n18640),.clk(gclk));
	jxor g18387(.dina(w_n17963_0[0]),.dinb(w_n5259_23[0]),.dout(n18641),.clk(gclk));
	jand g18388(.dina(n18641),.dinb(w_asqrt10_23[0]),.dout(n18642),.clk(gclk));
	jxor g18389(.dina(n18642),.dinb(w_n17968_0[0]),.dout(n18643),.clk(gclk));
	jand g18390(.dina(w_n18643_0[1]),.dinb(n18640),.dout(n18644),.clk(gclk));
	jor g18391(.dina(n18644),.dinb(w_n18639_0[1]),.dout(n18645),.clk(gclk));
	jand g18392(.dina(w_n18645_0[2]),.dinb(w_asqrt38_17[2]),.dout(n18646),.clk(gclk));
	jor g18393(.dina(w_n18645_0[1]),.dinb(w_asqrt38_17[1]),.dout(n18647),.clk(gclk));
	jxor g18394(.dina(w_n17971_0[0]),.dinb(w_n4902_27[0]),.dout(n18648),.clk(gclk));
	jand g18395(.dina(n18648),.dinb(w_asqrt10_22[2]),.dout(n18649),.clk(gclk));
	jxor g18396(.dina(n18649),.dinb(w_n17976_0[0]),.dout(n18650),.clk(gclk));
	jnot g18397(.din(w_n18650_0[1]),.dout(n18651),.clk(gclk));
	jand g18398(.dina(w_n18651_0[1]),.dinb(n18647),.dout(n18652),.clk(gclk));
	jor g18399(.dina(n18652),.dinb(w_n18646_0[1]),.dout(n18653),.clk(gclk));
	jand g18400(.dina(w_n18653_0[2]),.dinb(w_asqrt39_14[1]),.dout(n18654),.clk(gclk));
	jor g18401(.dina(w_n18653_0[1]),.dinb(w_asqrt39_14[0]),.dout(n18655),.clk(gclk));
	jxor g18402(.dina(w_n17978_0[0]),.dinb(w_n4582_24[0]),.dout(n18656),.clk(gclk));
	jand g18403(.dina(n18656),.dinb(w_asqrt10_22[1]),.dout(n18657),.clk(gclk));
	jxor g18404(.dina(n18657),.dinb(w_n17983_0[0]),.dout(n18658),.clk(gclk));
	jnot g18405(.din(w_n18658_0[1]),.dout(n18659),.clk(gclk));
	jand g18406(.dina(w_n18659_0[1]),.dinb(n18655),.dout(n18660),.clk(gclk));
	jor g18407(.dina(n18660),.dinb(w_n18654_0[1]),.dout(n18661),.clk(gclk));
	jand g18408(.dina(w_n18661_0[2]),.dinb(w_asqrt40_17[2]),.dout(n18662),.clk(gclk));
	jor g18409(.dina(w_n18661_0[1]),.dinb(w_asqrt40_17[1]),.dout(n18663),.clk(gclk));
	jxor g18410(.dina(w_n17985_0[0]),.dinb(w_n4249_27[2]),.dout(n18664),.clk(gclk));
	jand g18411(.dina(n18664),.dinb(w_asqrt10_22[0]),.dout(n18665),.clk(gclk));
	jxor g18412(.dina(n18665),.dinb(w_n17990_0[0]),.dout(n18666),.clk(gclk));
	jnot g18413(.din(w_n18666_0[1]),.dout(n18667),.clk(gclk));
	jand g18414(.dina(w_n18667_0[1]),.dinb(n18663),.dout(n18668),.clk(gclk));
	jor g18415(.dina(n18668),.dinb(w_n18662_0[1]),.dout(n18669),.clk(gclk));
	jand g18416(.dina(w_n18669_0[2]),.dinb(w_asqrt41_14[2]),.dout(n18670),.clk(gclk));
	jor g18417(.dina(w_n18669_0[1]),.dinb(w_asqrt41_14[1]),.dout(n18671),.clk(gclk));
	jxor g18418(.dina(w_n17992_0[0]),.dinb(w_n3955_24[2]),.dout(n18672),.clk(gclk));
	jand g18419(.dina(n18672),.dinb(w_asqrt10_21[2]),.dout(n18673),.clk(gclk));
	jxor g18420(.dina(n18673),.dinb(w_n17997_0[0]),.dout(n18674),.clk(gclk));
	jand g18421(.dina(w_n18674_0[1]),.dinb(n18671),.dout(n18675),.clk(gclk));
	jor g18422(.dina(n18675),.dinb(w_n18670_0[1]),.dout(n18676),.clk(gclk));
	jand g18423(.dina(w_n18676_0[2]),.dinb(w_asqrt42_18[0]),.dout(n18677),.clk(gclk));
	jor g18424(.dina(w_n18676_0[1]),.dinb(w_asqrt42_17[2]),.dout(n18678),.clk(gclk));
	jxor g18425(.dina(w_n18000_0[0]),.dinb(w_n3642_28[0]),.dout(n18679),.clk(gclk));
	jand g18426(.dina(n18679),.dinb(w_asqrt10_21[1]),.dout(n18680),.clk(gclk));
	jxor g18427(.dina(n18680),.dinb(w_n18005_0[0]),.dout(n18681),.clk(gclk));
	jnot g18428(.din(w_n18681_0[1]),.dout(n18682),.clk(gclk));
	jand g18429(.dina(w_n18682_0[1]),.dinb(n18678),.dout(n18683),.clk(gclk));
	jor g18430(.dina(n18683),.dinb(w_n18677_0[1]),.dout(n18684),.clk(gclk));
	jand g18431(.dina(w_n18684_0[2]),.dinb(w_asqrt43_15[0]),.dout(n18685),.clk(gclk));
	jor g18432(.dina(w_n18684_0[1]),.dinb(w_asqrt43_14[2]),.dout(n18686),.clk(gclk));
	jxor g18433(.dina(w_n18007_0[0]),.dinb(w_n3368_25[1]),.dout(n18687),.clk(gclk));
	jand g18434(.dina(n18687),.dinb(w_asqrt10_21[0]),.dout(n18688),.clk(gclk));
	jxor g18435(.dina(n18688),.dinb(w_n18013_0[0]),.dout(n18689),.clk(gclk));
	jnot g18436(.din(w_n18689_0[1]),.dout(n18690),.clk(gclk));
	jand g18437(.dina(w_n18690_0[1]),.dinb(n18686),.dout(n18691),.clk(gclk));
	jor g18438(.dina(n18691),.dinb(w_n18685_0[1]),.dout(n18692),.clk(gclk));
	jand g18439(.dina(w_n18692_0[2]),.dinb(w_asqrt44_18[0]),.dout(n18693),.clk(gclk));
	jor g18440(.dina(w_n18692_0[1]),.dinb(w_asqrt44_17[2]),.dout(n18694),.clk(gclk));
	jxor g18441(.dina(w_n18015_0[0]),.dinb(w_n3089_28[2]),.dout(n18695),.clk(gclk));
	jand g18442(.dina(n18695),.dinb(w_asqrt10_20[2]),.dout(n18696),.clk(gclk));
	jxor g18443(.dina(n18696),.dinb(w_n18020_0[0]),.dout(n18697),.clk(gclk));
	jnot g18444(.din(w_n18697_0[1]),.dout(n18698),.clk(gclk));
	jand g18445(.dina(w_n18698_0[1]),.dinb(n18694),.dout(n18699),.clk(gclk));
	jor g18446(.dina(n18699),.dinb(w_n18693_0[1]),.dout(n18700),.clk(gclk));
	jand g18447(.dina(w_n18700_0[2]),.dinb(w_asqrt45_15[2]),.dout(n18701),.clk(gclk));
	jor g18448(.dina(w_n18700_0[1]),.dinb(w_asqrt45_15[1]),.dout(n18702),.clk(gclk));
	jxor g18449(.dina(w_n18022_0[0]),.dinb(w_n2833_26[1]),.dout(n18703),.clk(gclk));
	jand g18450(.dina(n18703),.dinb(w_asqrt10_20[1]),.dout(n18704),.clk(gclk));
	jxor g18451(.dina(n18704),.dinb(w_n18027_0[0]),.dout(n18705),.clk(gclk));
	jnot g18452(.din(w_n18705_0[1]),.dout(n18706),.clk(gclk));
	jand g18453(.dina(w_n18706_0[1]),.dinb(n18702),.dout(n18707),.clk(gclk));
	jor g18454(.dina(n18707),.dinb(w_n18701_0[1]),.dout(n18708),.clk(gclk));
	jand g18455(.dina(w_n18708_0[2]),.dinb(w_asqrt46_18[0]),.dout(n18709),.clk(gclk));
	jor g18456(.dina(w_n18708_0[1]),.dinb(w_asqrt46_17[2]),.dout(n18710),.clk(gclk));
	jxor g18457(.dina(w_n18029_0[0]),.dinb(w_n2572_29[0]),.dout(n18711),.clk(gclk));
	jand g18458(.dina(n18711),.dinb(w_asqrt10_20[0]),.dout(n18712),.clk(gclk));
	jxor g18459(.dina(n18712),.dinb(w_n18034_0[0]),.dout(n18713),.clk(gclk));
	jnot g18460(.din(w_n18713_0[1]),.dout(n18714),.clk(gclk));
	jand g18461(.dina(w_n18714_0[1]),.dinb(n18710),.dout(n18715),.clk(gclk));
	jor g18462(.dina(n18715),.dinb(w_n18709_0[1]),.dout(n18716),.clk(gclk));
	jand g18463(.dina(w_n18716_0[2]),.dinb(w_asqrt47_16[1]),.dout(n18717),.clk(gclk));
	jor g18464(.dina(w_n18716_0[1]),.dinb(w_asqrt47_16[0]),.dout(n18718),.clk(gclk));
	jxor g18465(.dina(w_n18036_0[0]),.dinb(w_n2345_27[0]),.dout(n18719),.clk(gclk));
	jand g18466(.dina(n18719),.dinb(w_asqrt10_19[2]),.dout(n18720),.clk(gclk));
	jxor g18467(.dina(n18720),.dinb(w_n18041_0[0]),.dout(n18721),.clk(gclk));
	jand g18468(.dina(w_n18721_0[1]),.dinb(n18718),.dout(n18722),.clk(gclk));
	jor g18469(.dina(n18722),.dinb(w_n18717_0[1]),.dout(n18723),.clk(gclk));
	jand g18470(.dina(w_n18723_0[2]),.dinb(w_asqrt48_18[1]),.dout(n18724),.clk(gclk));
	jor g18471(.dina(w_n18723_0[1]),.dinb(w_asqrt48_18[0]),.dout(n18725),.clk(gclk));
	jxor g18472(.dina(w_n18044_0[0]),.dinb(w_n2108_29[2]),.dout(n18726),.clk(gclk));
	jand g18473(.dina(n18726),.dinb(w_asqrt10_19[1]),.dout(n18727),.clk(gclk));
	jxor g18474(.dina(n18727),.dinb(w_n18049_0[0]),.dout(n18728),.clk(gclk));
	jnot g18475(.din(w_n18728_0[1]),.dout(n18729),.clk(gclk));
	jand g18476(.dina(w_n18729_0[1]),.dinb(n18725),.dout(n18730),.clk(gclk));
	jor g18477(.dina(n18730),.dinb(w_n18724_0[1]),.dout(n18731),.clk(gclk));
	jand g18478(.dina(w_n18731_0[2]),.dinb(w_asqrt49_16[2]),.dout(n18732),.clk(gclk));
	jor g18479(.dina(w_n18731_0[1]),.dinb(w_asqrt49_16[1]),.dout(n18733),.clk(gclk));
	jxor g18480(.dina(w_n18051_0[0]),.dinb(w_n1912_28[0]),.dout(n18734),.clk(gclk));
	jand g18481(.dina(n18734),.dinb(w_asqrt10_19[0]),.dout(n18735),.clk(gclk));
	jxor g18482(.dina(n18735),.dinb(w_n18056_0[0]),.dout(n18736),.clk(gclk));
	jand g18483(.dina(w_n18736_0[1]),.dinb(n18733),.dout(n18737),.clk(gclk));
	jor g18484(.dina(n18737),.dinb(w_n18732_0[1]),.dout(n18738),.clk(gclk));
	jand g18485(.dina(w_n18738_0[2]),.dinb(w_asqrt50_18[2]),.dout(n18739),.clk(gclk));
	jor g18486(.dina(w_n18738_0[1]),.dinb(w_asqrt50_18[1]),.dout(n18740),.clk(gclk));
	jxor g18487(.dina(w_n18059_0[0]),.dinb(w_n1699_30[1]),.dout(n18741),.clk(gclk));
	jand g18488(.dina(n18741),.dinb(w_asqrt10_18[2]),.dout(n18742),.clk(gclk));
	jxor g18489(.dina(n18742),.dinb(w_n18064_0[0]),.dout(n18743),.clk(gclk));
	jnot g18490(.din(w_n18743_0[1]),.dout(n18744),.clk(gclk));
	jand g18491(.dina(w_n18744_0[1]),.dinb(n18740),.dout(n18745),.clk(gclk));
	jor g18492(.dina(n18745),.dinb(w_n18739_0[1]),.dout(n18746),.clk(gclk));
	jand g18493(.dina(w_n18746_0[2]),.dinb(w_asqrt51_17[0]),.dout(n18747),.clk(gclk));
	jor g18494(.dina(w_n18746_0[1]),.dinb(w_asqrt51_16[2]),.dout(n18748),.clk(gclk));
	jxor g18495(.dina(w_n18066_0[0]),.dinb(w_n1516_28[2]),.dout(n18749),.clk(gclk));
	jand g18496(.dina(n18749),.dinb(w_asqrt10_18[1]),.dout(n18750),.clk(gclk));
	jxor g18497(.dina(n18750),.dinb(w_n18071_0[0]),.dout(n18751),.clk(gclk));
	jnot g18498(.din(w_n18751_0[1]),.dout(n18752),.clk(gclk));
	jand g18499(.dina(w_n18752_0[1]),.dinb(n18748),.dout(n18753),.clk(gclk));
	jor g18500(.dina(n18753),.dinb(w_n18747_0[1]),.dout(n18754),.clk(gclk));
	jand g18501(.dina(w_n18754_0[2]),.dinb(w_asqrt52_18[2]),.dout(n18755),.clk(gclk));
	jor g18502(.dina(w_n18754_0[1]),.dinb(w_asqrt52_18[1]),.dout(n18756),.clk(gclk));
	jxor g18503(.dina(w_n18073_0[0]),.dinb(w_n1332_30[1]),.dout(n18757),.clk(gclk));
	jand g18504(.dina(n18757),.dinb(w_asqrt10_18[0]),.dout(n18758),.clk(gclk));
	jxor g18505(.dina(n18758),.dinb(w_n18078_0[0]),.dout(n18759),.clk(gclk));
	jand g18506(.dina(w_n18759_0[1]),.dinb(n18756),.dout(n18760),.clk(gclk));
	jor g18507(.dina(n18760),.dinb(w_n18755_0[1]),.dout(n18761),.clk(gclk));
	jand g18508(.dina(w_n18761_0[2]),.dinb(w_asqrt53_17[2]),.dout(n18762),.clk(gclk));
	jxor g18509(.dina(w_n18081_0[0]),.dinb(w_n1173_29[1]),.dout(n18763),.clk(gclk));
	jand g18510(.dina(n18763),.dinb(w_asqrt10_17[2]),.dout(n18764),.clk(gclk));
	jxor g18511(.dina(n18764),.dinb(w_n18085_0[0]),.dout(n18765),.clk(gclk));
	jor g18512(.dina(w_n18761_0[1]),.dinb(w_asqrt53_17[1]),.dout(n18766),.clk(gclk));
	jand g18513(.dina(n18766),.dinb(w_n18765_0[1]),.dout(n18767),.clk(gclk));
	jor g18514(.dina(n18767),.dinb(w_n18762_0[1]),.dout(n18768),.clk(gclk));
	jand g18515(.dina(w_n18768_0[2]),.dinb(w_asqrt54_18[2]),.dout(n18769),.clk(gclk));
	jor g18516(.dina(w_n18768_0[1]),.dinb(w_asqrt54_18[1]),.dout(n18770),.clk(gclk));
	jxor g18517(.dina(w_n18089_0[0]),.dinb(w_n1008_31[1]),.dout(n18771),.clk(gclk));
	jand g18518(.dina(n18771),.dinb(w_asqrt10_17[1]),.dout(n18772),.clk(gclk));
	jxor g18519(.dina(n18772),.dinb(w_n18094_0[0]),.dout(n18773),.clk(gclk));
	jnot g18520(.din(w_n18773_0[1]),.dout(n18774),.clk(gclk));
	jand g18521(.dina(w_n18774_0[1]),.dinb(n18770),.dout(n18775),.clk(gclk));
	jor g18522(.dina(n18775),.dinb(w_n18769_0[1]),.dout(n18776),.clk(gclk));
	jand g18523(.dina(w_n18776_0[2]),.dinb(w_asqrt55_18[0]),.dout(n18777),.clk(gclk));
	jor g18524(.dina(w_n18776_0[1]),.dinb(w_asqrt55_17[2]),.dout(n18778),.clk(gclk));
	jxor g18525(.dina(w_n18096_0[0]),.dinb(w_n884_30[1]),.dout(n18779),.clk(gclk));
	jand g18526(.dina(n18779),.dinb(w_asqrt10_17[0]),.dout(n18780),.clk(gclk));
	jxor g18527(.dina(n18780),.dinb(w_n18101_0[0]),.dout(n18781),.clk(gclk));
	jand g18528(.dina(w_n18781_0[1]),.dinb(n18778),.dout(n18782),.clk(gclk));
	jor g18529(.dina(n18782),.dinb(w_n18777_0[1]),.dout(n18783),.clk(gclk));
	jand g18530(.dina(w_n18783_0[2]),.dinb(w_asqrt56_19[0]),.dout(n18784),.clk(gclk));
	jor g18531(.dina(w_n18783_0[1]),.dinb(w_asqrt56_18[2]),.dout(n18785),.clk(gclk));
	jxor g18532(.dina(w_n18104_0[0]),.dinb(w_n743_31[1]),.dout(n18786),.clk(gclk));
	jand g18533(.dina(n18786),.dinb(w_asqrt10_16[2]),.dout(n18787),.clk(gclk));
	jxor g18534(.dina(n18787),.dinb(w_n18109_0[0]),.dout(n18788),.clk(gclk));
	jnot g18535(.din(w_n18788_0[1]),.dout(n18789),.clk(gclk));
	jand g18536(.dina(w_n18789_0[1]),.dinb(n18785),.dout(n18790),.clk(gclk));
	jor g18537(.dina(n18790),.dinb(w_n18784_0[1]),.dout(n18791),.clk(gclk));
	jand g18538(.dina(w_n18791_0[2]),.dinb(w_asqrt57_18[2]),.dout(n18792),.clk(gclk));
	jor g18539(.dina(w_n18791_0[1]),.dinb(w_asqrt57_18[1]),.dout(n18793),.clk(gclk));
	jxor g18540(.dina(w_n18111_0[0]),.dinb(w_n635_31[1]),.dout(n18794),.clk(gclk));
	jand g18541(.dina(n18794),.dinb(w_asqrt10_16[1]),.dout(n18795),.clk(gclk));
	jxor g18542(.dina(n18795),.dinb(w_n18116_0[0]),.dout(n18796),.clk(gclk));
	jand g18543(.dina(w_n18796_0[1]),.dinb(n18793),.dout(n18797),.clk(gclk));
	jor g18544(.dina(n18797),.dinb(w_n18792_0[1]),.dout(n18798),.clk(gclk));
	jand g18545(.dina(w_n18798_0[2]),.dinb(w_asqrt58_19[1]),.dout(n18799),.clk(gclk));
	jor g18546(.dina(w_n18798_0[1]),.dinb(w_asqrt58_19[0]),.dout(n18800),.clk(gclk));
	jxor g18547(.dina(w_n18119_0[0]),.dinb(w_n515_32[1]),.dout(n18801),.clk(gclk));
	jand g18548(.dina(n18801),.dinb(w_asqrt10_16[0]),.dout(n18802),.clk(gclk));
	jxor g18549(.dina(n18802),.dinb(w_n18124_0[0]),.dout(n18803),.clk(gclk));
	jnot g18550(.din(w_n18803_0[2]),.dout(n18804),.clk(gclk));
	jand g18551(.dina(n18804),.dinb(n18800),.dout(n18805),.clk(gclk));
	jor g18552(.dina(n18805),.dinb(w_n18799_0[1]),.dout(n18806),.clk(gclk));
	jand g18553(.dina(w_n18806_0[2]),.dinb(w_asqrt59_19[0]),.dout(n18807),.clk(gclk));
	jor g18554(.dina(w_n18806_0[1]),.dinb(w_asqrt59_18[2]),.dout(n18808),.clk(gclk));
	jxor g18555(.dina(w_n18126_0[0]),.dinb(w_n443_32[1]),.dout(n18809),.clk(gclk));
	jand g18556(.dina(n18809),.dinb(w_asqrt10_15[2]),.dout(n18810),.clk(gclk));
	jxor g18557(.dina(n18810),.dinb(w_n18131_0[0]),.dout(n18811),.clk(gclk));
	jnot g18558(.din(w_n18811_0[1]),.dout(n18812),.clk(gclk));
	jand g18559(.dina(w_n18812_0[1]),.dinb(n18808),.dout(n18813),.clk(gclk));
	jor g18560(.dina(n18813),.dinb(w_n18807_0[1]),.dout(n18814),.clk(gclk));
	jand g18561(.dina(w_n18814_0[2]),.dinb(w_asqrt60_19[1]),.dout(n18815),.clk(gclk));
	jor g18562(.dina(w_n18814_0[1]),.dinb(w_asqrt60_19[0]),.dout(n18816),.clk(gclk));
	jxor g18563(.dina(w_n18133_0[0]),.dinb(w_n352_32[2]),.dout(n18817),.clk(gclk));
	jand g18564(.dina(n18817),.dinb(w_asqrt10_15[1]),.dout(n18818),.clk(gclk));
	jxor g18565(.dina(n18818),.dinb(w_n18138_0[0]),.dout(n18819),.clk(gclk));
	jnot g18566(.din(w_n18819_0[1]),.dout(n18820),.clk(gclk));
	jand g18567(.dina(w_n18820_0[1]),.dinb(n18816),.dout(n18821),.clk(gclk));
	jor g18568(.dina(n18821),.dinb(w_n18815_0[1]),.dout(n18822),.clk(gclk));
	jand g18569(.dina(w_n18822_0[2]),.dinb(w_asqrt61_19[1]),.dout(n18823),.clk(gclk));
	jor g18570(.dina(w_n18822_0[1]),.dinb(w_asqrt61_19[0]),.dout(n18824),.clk(gclk));
	jxor g18571(.dina(w_n18140_0[0]),.dinb(w_n294_33[0]),.dout(n18825),.clk(gclk));
	jand g18572(.dina(n18825),.dinb(w_asqrt10_15[0]),.dout(n18826),.clk(gclk));
	jxor g18573(.dina(n18826),.dinb(w_n18145_0[0]),.dout(n18827),.clk(gclk));
	jand g18574(.dina(w_n18827_0[1]),.dinb(n18824),.dout(n18828),.clk(gclk));
	jor g18575(.dina(n18828),.dinb(w_n18823_0[1]),.dout(n18829),.clk(gclk));
	jand g18576(.dina(w_n18829_0[2]),.dinb(w_asqrt62_19[1]),.dout(n18830),.clk(gclk));
	jnot g18577(.din(w_n18830_0[1]),.dout(n18831),.clk(gclk));
	jnot g18578(.din(w_n18823_0[0]),.dout(n18832),.clk(gclk));
	jnot g18579(.din(w_n18815_0[0]),.dout(n18833),.clk(gclk));
	jnot g18580(.din(w_n18807_0[0]),.dout(n18834),.clk(gclk));
	jnot g18581(.din(w_n18799_0[0]),.dout(n18835),.clk(gclk));
	jnot g18582(.din(w_n18792_0[0]),.dout(n18836),.clk(gclk));
	jnot g18583(.din(w_n18784_0[0]),.dout(n18837),.clk(gclk));
	jnot g18584(.din(w_n18777_0[0]),.dout(n18838),.clk(gclk));
	jnot g18585(.din(w_n18769_0[0]),.dout(n18839),.clk(gclk));
	jnot g18586(.din(w_n18762_0[0]),.dout(n18840),.clk(gclk));
	jnot g18587(.din(w_n18765_0[0]),.dout(n18841),.clk(gclk));
	jnot g18588(.din(w_n18755_0[0]),.dout(n18842),.clk(gclk));
	jnot g18589(.din(w_n18747_0[0]),.dout(n18843),.clk(gclk));
	jnot g18590(.din(w_n18739_0[0]),.dout(n18844),.clk(gclk));
	jnot g18591(.din(w_n18732_0[0]),.dout(n18845),.clk(gclk));
	jnot g18592(.din(w_n18724_0[0]),.dout(n18846),.clk(gclk));
	jnot g18593(.din(w_n18717_0[0]),.dout(n18847),.clk(gclk));
	jnot g18594(.din(w_n18709_0[0]),.dout(n18848),.clk(gclk));
	jnot g18595(.din(w_n18701_0[0]),.dout(n18849),.clk(gclk));
	jnot g18596(.din(w_n18693_0[0]),.dout(n18850),.clk(gclk));
	jnot g18597(.din(w_n18685_0[0]),.dout(n18851),.clk(gclk));
	jnot g18598(.din(w_n18677_0[0]),.dout(n18852),.clk(gclk));
	jnot g18599(.din(w_n18670_0[0]),.dout(n18853),.clk(gclk));
	jnot g18600(.din(w_n18662_0[0]),.dout(n18854),.clk(gclk));
	jnot g18601(.din(w_n18654_0[0]),.dout(n18855),.clk(gclk));
	jnot g18602(.din(w_n18646_0[0]),.dout(n18856),.clk(gclk));
	jnot g18603(.din(w_n18639_0[0]),.dout(n18857),.clk(gclk));
	jnot g18604(.din(w_n18631_0[0]),.dout(n18858),.clk(gclk));
	jnot g18605(.din(w_n18624_0[0]),.dout(n18859),.clk(gclk));
	jnot g18606(.din(w_n18616_0[0]),.dout(n18860),.clk(gclk));
	jnot g18607(.din(w_n18609_0[0]),.dout(n18861),.clk(gclk));
	jnot g18608(.din(w_n18601_0[0]),.dout(n18862),.clk(gclk));
	jnot g18609(.din(w_n18594_0[0]),.dout(n18863),.clk(gclk));
	jnot g18610(.din(w_n18586_0[0]),.dout(n18864),.clk(gclk));
	jnot g18611(.din(w_n18578_0[0]),.dout(n18865),.clk(gclk));
	jnot g18612(.din(w_n18570_0[0]),.dout(n18866),.clk(gclk));
	jnot g18613(.din(w_n18563_0[0]),.dout(n18867),.clk(gclk));
	jnot g18614(.din(w_n18555_0[0]),.dout(n18868),.clk(gclk));
	jnot g18615(.din(w_n18548_0[0]),.dout(n18869),.clk(gclk));
	jnot g18616(.din(w_n18540_0[0]),.dout(n18870),.clk(gclk));
	jnot g18617(.din(w_n18533_0[0]),.dout(n18871),.clk(gclk));
	jnot g18618(.din(w_n18526_0[0]),.dout(n18872),.clk(gclk));
	jnot g18619(.din(w_n18518_0[0]),.dout(n18873),.clk(gclk));
	jnot g18620(.din(w_n18510_0[0]),.dout(n18874),.clk(gclk));
	jnot g18621(.din(w_n18503_0[0]),.dout(n18875),.clk(gclk));
	jnot g18622(.din(w_n18495_0[0]),.dout(n18876),.clk(gclk));
	jnot g18623(.din(w_n18488_0[0]),.dout(n18877),.clk(gclk));
	jnot g18624(.din(w_n18480_0[0]),.dout(n18878),.clk(gclk));
	jnot g18625(.din(w_n18473_0[0]),.dout(n18879),.clk(gclk));
	jnot g18626(.din(w_n18465_0[0]),.dout(n18880),.clk(gclk));
	jnot g18627(.din(w_n18458_0[0]),.dout(n18881),.clk(gclk));
	jnot g18628(.din(w_n18447_0[0]),.dout(n18882),.clk(gclk));
	jnot g18629(.din(w_n18190_0[0]),.dout(n18883),.clk(gclk));
	jor g18630(.dina(w_n18442_12[1]),.dinb(w_n17774_0[2]),.dout(n18884),.clk(gclk));
	jnot g18631(.din(w_n18188_0[0]),.dout(n18885),.clk(gclk));
	jand g18632(.dina(n18885),.dinb(n18884),.dout(n18886),.clk(gclk));
	jand g18633(.dina(n18886),.dinb(w_n17769_20[1]),.dout(n18887),.clk(gclk));
	jor g18634(.dina(w_n18442_12[0]),.dinb(w_a20_0[0]),.dout(n18888),.clk(gclk));
	jand g18635(.dina(n18888),.dinb(w_a21_0[0]),.dout(n18889),.clk(gclk));
	jor g18636(.dina(w_n18449_0[0]),.dinb(n18889),.dout(n18890),.clk(gclk));
	jor g18637(.dina(w_n18890_0[1]),.dinb(n18887),.dout(n18891),.clk(gclk));
	jand g18638(.dina(n18891),.dinb(n18883),.dout(n18892),.clk(gclk));
	jand g18639(.dina(n18892),.dinb(w_n17134_12[2]),.dout(n18893),.clk(gclk));
	jor g18640(.dina(w_n18454_0[0]),.dinb(n18893),.dout(n18894),.clk(gclk));
	jand g18641(.dina(n18894),.dinb(n18882),.dout(n18895),.clk(gclk));
	jand g18642(.dina(n18895),.dinb(w_n16489_20[2]),.dout(n18896),.clk(gclk));
	jnot g18643(.din(w_n18462_0[0]),.dout(n18897),.clk(gclk));
	jor g18644(.dina(w_n18897_0[1]),.dinb(n18896),.dout(n18898),.clk(gclk));
	jand g18645(.dina(n18898),.dinb(n18881),.dout(n18899),.clk(gclk));
	jand g18646(.dina(n18899),.dinb(w_n15878_13[2]),.dout(n18900),.clk(gclk));
	jor g18647(.dina(w_n18469_0[0]),.dinb(n18900),.dout(n18901),.clk(gclk));
	jand g18648(.dina(n18901),.dinb(n18880),.dout(n18902),.clk(gclk));
	jand g18649(.dina(n18902),.dinb(w_n15260_21[1]),.dout(n18903),.clk(gclk));
	jnot g18650(.din(w_n18477_0[0]),.dout(n18904),.clk(gclk));
	jor g18651(.dina(w_n18904_0[1]),.dinb(n18903),.dout(n18905),.clk(gclk));
	jand g18652(.dina(n18905),.dinb(n18879),.dout(n18906),.clk(gclk));
	jand g18653(.dina(n18906),.dinb(w_n14674_14[1]),.dout(n18907),.clk(gclk));
	jor g18654(.dina(w_n18484_0[0]),.dinb(n18907),.dout(n18908),.clk(gclk));
	jand g18655(.dina(n18908),.dinb(n18878),.dout(n18909),.clk(gclk));
	jand g18656(.dina(n18909),.dinb(w_n14078_21[2]),.dout(n18910),.clk(gclk));
	jnot g18657(.din(w_n18492_0[0]),.dout(n18911),.clk(gclk));
	jor g18658(.dina(w_n18911_0[1]),.dinb(n18910),.dout(n18912),.clk(gclk));
	jand g18659(.dina(n18912),.dinb(n18877),.dout(n18913),.clk(gclk));
	jand g18660(.dina(n18913),.dinb(w_n13515_15[1]),.dout(n18914),.clk(gclk));
	jor g18661(.dina(w_n18499_0[0]),.dinb(n18914),.dout(n18915),.clk(gclk));
	jand g18662(.dina(n18915),.dinb(n18876),.dout(n18916),.clk(gclk));
	jand g18663(.dina(n18916),.dinb(w_n12947_22[1]),.dout(n18917),.clk(gclk));
	jnot g18664(.din(w_n18507_0[0]),.dout(n18918),.clk(gclk));
	jor g18665(.dina(w_n18918_0[1]),.dinb(n18917),.dout(n18919),.clk(gclk));
	jand g18666(.dina(n18919),.dinb(n18875),.dout(n18920),.clk(gclk));
	jand g18667(.dina(n18920),.dinb(w_n12410_16[0]),.dout(n18921),.clk(gclk));
	jor g18668(.dina(w_n18514_0[0]),.dinb(n18921),.dout(n18922),.clk(gclk));
	jand g18669(.dina(n18922),.dinb(n18874),.dout(n18923),.clk(gclk));
	jand g18670(.dina(n18923),.dinb(w_n11858_22[2]),.dout(n18924),.clk(gclk));
	jor g18671(.dina(w_n18522_0[0]),.dinb(n18924),.dout(n18925),.clk(gclk));
	jand g18672(.dina(n18925),.dinb(n18873),.dout(n18926),.clk(gclk));
	jand g18673(.dina(n18926),.dinb(w_n11347_16[2]),.dout(n18927),.clk(gclk));
	jnot g18674(.din(w_n18530_0[0]),.dout(n18928),.clk(gclk));
	jor g18675(.dina(w_n18928_0[1]),.dinb(n18927),.dout(n18929),.clk(gclk));
	jand g18676(.dina(n18929),.dinb(n18872),.dout(n18930),.clk(gclk));
	jand g18677(.dina(n18930),.dinb(w_n10824_23[1]),.dout(n18931),.clk(gclk));
	jnot g18678(.din(w_n18537_0[0]),.dout(n18932),.clk(gclk));
	jor g18679(.dina(w_n18932_0[1]),.dinb(n18931),.dout(n18933),.clk(gclk));
	jand g18680(.dina(n18933),.dinb(n18871),.dout(n18934),.clk(gclk));
	jand g18681(.dina(n18934),.dinb(w_n10328_17[2]),.dout(n18935),.clk(gclk));
	jor g18682(.dina(w_n18544_0[0]),.dinb(n18935),.dout(n18936),.clk(gclk));
	jand g18683(.dina(n18936),.dinb(n18870),.dout(n18937),.clk(gclk));
	jand g18684(.dina(n18937),.dinb(w_n9832_24[0]),.dout(n18938),.clk(gclk));
	jnot g18685(.din(w_n18552_0[0]),.dout(n18939),.clk(gclk));
	jor g18686(.dina(w_n18939_0[1]),.dinb(n18938),.dout(n18940),.clk(gclk));
	jand g18687(.dina(n18940),.dinb(n18869),.dout(n18941),.clk(gclk));
	jand g18688(.dina(n18941),.dinb(w_n9369_18[2]),.dout(n18942),.clk(gclk));
	jor g18689(.dina(w_n18559_0[0]),.dinb(n18942),.dout(n18943),.clk(gclk));
	jand g18690(.dina(n18943),.dinb(n18868),.dout(n18944),.clk(gclk));
	jand g18691(.dina(n18944),.dinb(w_n8890_24[1]),.dout(n18945),.clk(gclk));
	jnot g18692(.din(w_n18567_0[0]),.dout(n18946),.clk(gclk));
	jor g18693(.dina(w_n18946_0[1]),.dinb(n18945),.dout(n18947),.clk(gclk));
	jand g18694(.dina(n18947),.dinb(n18867),.dout(n18948),.clk(gclk));
	jand g18695(.dina(n18948),.dinb(w_n8449_19[1]),.dout(n18949),.clk(gclk));
	jor g18696(.dina(w_n18574_0[0]),.dinb(n18949),.dout(n18950),.clk(gclk));
	jand g18697(.dina(n18950),.dinb(n18866),.dout(n18951),.clk(gclk));
	jand g18698(.dina(n18951),.dinb(w_n8003_25[0]),.dout(n18952),.clk(gclk));
	jor g18699(.dina(w_n18582_0[0]),.dinb(n18952),.dout(n18953),.clk(gclk));
	jand g18700(.dina(n18953),.dinb(n18865),.dout(n18954),.clk(gclk));
	jand g18701(.dina(n18954),.dinb(w_n7581_20[1]),.dout(n18955),.clk(gclk));
	jor g18702(.dina(w_n18590_0[0]),.dinb(n18955),.dout(n18956),.clk(gclk));
	jand g18703(.dina(n18956),.dinb(n18864),.dout(n18957),.clk(gclk));
	jand g18704(.dina(n18957),.dinb(w_n7154_25[1]),.dout(n18958),.clk(gclk));
	jnot g18705(.din(w_n18598_0[0]),.dout(n18959),.clk(gclk));
	jor g18706(.dina(w_n18959_0[1]),.dinb(n18958),.dout(n18960),.clk(gclk));
	jand g18707(.dina(n18960),.dinb(n18863),.dout(n18961),.clk(gclk));
	jand g18708(.dina(n18961),.dinb(w_n6758_21[0]),.dout(n18962),.clk(gclk));
	jor g18709(.dina(w_n18605_0[0]),.dinb(n18962),.dout(n18963),.clk(gclk));
	jand g18710(.dina(n18963),.dinb(n18862),.dout(n18964),.clk(gclk));
	jand g18711(.dina(n18964),.dinb(w_n6357_25[2]),.dout(n18965),.clk(gclk));
	jnot g18712(.din(w_n18613_0[0]),.dout(n18966),.clk(gclk));
	jor g18713(.dina(w_n18966_0[1]),.dinb(n18965),.dout(n18967),.clk(gclk));
	jand g18714(.dina(n18967),.dinb(n18861),.dout(n18968),.clk(gclk));
	jand g18715(.dina(n18968),.dinb(w_n5989_21[2]),.dout(n18969),.clk(gclk));
	jor g18716(.dina(w_n18620_0[0]),.dinb(n18969),.dout(n18970),.clk(gclk));
	jand g18717(.dina(n18970),.dinb(n18860),.dout(n18971),.clk(gclk));
	jand g18718(.dina(n18971),.dinb(w_n5606_26[0]),.dout(n18972),.clk(gclk));
	jnot g18719(.din(w_n18628_0[0]),.dout(n18973),.clk(gclk));
	jor g18720(.dina(w_n18973_0[1]),.dinb(n18972),.dout(n18974),.clk(gclk));
	jand g18721(.dina(n18974),.dinb(n18859),.dout(n18975),.clk(gclk));
	jand g18722(.dina(n18975),.dinb(w_n5259_22[2]),.dout(n18976),.clk(gclk));
	jor g18723(.dina(w_n18635_0[0]),.dinb(n18976),.dout(n18977),.clk(gclk));
	jand g18724(.dina(n18977),.dinb(n18858),.dout(n18978),.clk(gclk));
	jand g18725(.dina(n18978),.dinb(w_n4902_26[2]),.dout(n18979),.clk(gclk));
	jnot g18726(.din(w_n18643_0[0]),.dout(n18980),.clk(gclk));
	jor g18727(.dina(w_n18980_0[1]),.dinb(n18979),.dout(n18981),.clk(gclk));
	jand g18728(.dina(n18981),.dinb(n18857),.dout(n18982),.clk(gclk));
	jand g18729(.dina(n18982),.dinb(w_n4582_23[2]),.dout(n18983),.clk(gclk));
	jor g18730(.dina(w_n18650_0[0]),.dinb(n18983),.dout(n18984),.clk(gclk));
	jand g18731(.dina(n18984),.dinb(n18856),.dout(n18985),.clk(gclk));
	jand g18732(.dina(n18985),.dinb(w_n4249_27[1]),.dout(n18986),.clk(gclk));
	jor g18733(.dina(w_n18658_0[0]),.dinb(n18986),.dout(n18987),.clk(gclk));
	jand g18734(.dina(n18987),.dinb(n18855),.dout(n18988),.clk(gclk));
	jand g18735(.dina(n18988),.dinb(w_n3955_24[1]),.dout(n18989),.clk(gclk));
	jor g18736(.dina(w_n18666_0[0]),.dinb(n18989),.dout(n18990),.clk(gclk));
	jand g18737(.dina(n18990),.dinb(n18854),.dout(n18991),.clk(gclk));
	jand g18738(.dina(n18991),.dinb(w_n3642_27[2]),.dout(n18992),.clk(gclk));
	jnot g18739(.din(w_n18674_0[0]),.dout(n18993),.clk(gclk));
	jor g18740(.dina(w_n18993_0[1]),.dinb(n18992),.dout(n18994),.clk(gclk));
	jand g18741(.dina(n18994),.dinb(n18853),.dout(n18995),.clk(gclk));
	jand g18742(.dina(n18995),.dinb(w_n3368_25[0]),.dout(n18996),.clk(gclk));
	jor g18743(.dina(w_n18681_0[0]),.dinb(n18996),.dout(n18997),.clk(gclk));
	jand g18744(.dina(n18997),.dinb(n18852),.dout(n18998),.clk(gclk));
	jand g18745(.dina(n18998),.dinb(w_n3089_28[1]),.dout(n18999),.clk(gclk));
	jor g18746(.dina(w_n18689_0[0]),.dinb(n18999),.dout(n19000),.clk(gclk));
	jand g18747(.dina(n19000),.dinb(n18851),.dout(n19001),.clk(gclk));
	jand g18748(.dina(n19001),.dinb(w_n2833_26[0]),.dout(n19002),.clk(gclk));
	jor g18749(.dina(w_n18697_0[0]),.dinb(n19002),.dout(n19003),.clk(gclk));
	jand g18750(.dina(n19003),.dinb(n18850),.dout(n19004),.clk(gclk));
	jand g18751(.dina(n19004),.dinb(w_n2572_28[2]),.dout(n19005),.clk(gclk));
	jor g18752(.dina(w_n18705_0[0]),.dinb(n19005),.dout(n19006),.clk(gclk));
	jand g18753(.dina(n19006),.dinb(n18849),.dout(n19007),.clk(gclk));
	jand g18754(.dina(n19007),.dinb(w_n2345_26[2]),.dout(n19008),.clk(gclk));
	jor g18755(.dina(w_n18713_0[0]),.dinb(n19008),.dout(n19009),.clk(gclk));
	jand g18756(.dina(n19009),.dinb(n18848),.dout(n19010),.clk(gclk));
	jand g18757(.dina(n19010),.dinb(w_n2108_29[1]),.dout(n19011),.clk(gclk));
	jnot g18758(.din(w_n18721_0[0]),.dout(n19012),.clk(gclk));
	jor g18759(.dina(w_n19012_0[1]),.dinb(n19011),.dout(n19013),.clk(gclk));
	jand g18760(.dina(n19013),.dinb(n18847),.dout(n19014),.clk(gclk));
	jand g18761(.dina(n19014),.dinb(w_n1912_27[2]),.dout(n19015),.clk(gclk));
	jor g18762(.dina(w_n18728_0[0]),.dinb(n19015),.dout(n19016),.clk(gclk));
	jand g18763(.dina(n19016),.dinb(n18846),.dout(n19017),.clk(gclk));
	jand g18764(.dina(n19017),.dinb(w_n1699_30[0]),.dout(n19018),.clk(gclk));
	jnot g18765(.din(w_n18736_0[0]),.dout(n19019),.clk(gclk));
	jor g18766(.dina(w_n19019_0[1]),.dinb(n19018),.dout(n19020),.clk(gclk));
	jand g18767(.dina(n19020),.dinb(n18845),.dout(n19021),.clk(gclk));
	jand g18768(.dina(n19021),.dinb(w_n1516_28[1]),.dout(n19022),.clk(gclk));
	jor g18769(.dina(w_n18743_0[0]),.dinb(n19022),.dout(n19023),.clk(gclk));
	jand g18770(.dina(n19023),.dinb(n18844),.dout(n19024),.clk(gclk));
	jand g18771(.dina(n19024),.dinb(w_n1332_30[0]),.dout(n19025),.clk(gclk));
	jor g18772(.dina(w_n18751_0[0]),.dinb(n19025),.dout(n19026),.clk(gclk));
	jand g18773(.dina(n19026),.dinb(n18843),.dout(n19027),.clk(gclk));
	jand g18774(.dina(n19027),.dinb(w_n1173_29[0]),.dout(n19028),.clk(gclk));
	jnot g18775(.din(w_n18759_0[0]),.dout(n19029),.clk(gclk));
	jor g18776(.dina(w_n19029_0[1]),.dinb(n19028),.dout(n19030),.clk(gclk));
	jand g18777(.dina(n19030),.dinb(n18842),.dout(n19031),.clk(gclk));
	jand g18778(.dina(n19031),.dinb(w_n1008_31[0]),.dout(n19032),.clk(gclk));
	jor g18779(.dina(n19032),.dinb(w_n18841_0[1]),.dout(n19033),.clk(gclk));
	jand g18780(.dina(n19033),.dinb(n18840),.dout(n19034),.clk(gclk));
	jand g18781(.dina(n19034),.dinb(w_n884_30[0]),.dout(n19035),.clk(gclk));
	jor g18782(.dina(w_n18773_0[0]),.dinb(n19035),.dout(n19036),.clk(gclk));
	jand g18783(.dina(n19036),.dinb(n18839),.dout(n19037),.clk(gclk));
	jand g18784(.dina(n19037),.dinb(w_n743_31[0]),.dout(n19038),.clk(gclk));
	jnot g18785(.din(w_n18781_0[0]),.dout(n19039),.clk(gclk));
	jor g18786(.dina(w_n19039_0[1]),.dinb(n19038),.dout(n19040),.clk(gclk));
	jand g18787(.dina(n19040),.dinb(n18838),.dout(n19041),.clk(gclk));
	jand g18788(.dina(n19041),.dinb(w_n635_31[0]),.dout(n19042),.clk(gclk));
	jor g18789(.dina(w_n18788_0[0]),.dinb(n19042),.dout(n19043),.clk(gclk));
	jand g18790(.dina(n19043),.dinb(n18837),.dout(n19044),.clk(gclk));
	jand g18791(.dina(n19044),.dinb(w_n515_32[0]),.dout(n19045),.clk(gclk));
	jnot g18792(.din(w_n18796_0[0]),.dout(n19046),.clk(gclk));
	jor g18793(.dina(w_n19046_0[1]),.dinb(n19045),.dout(n19047),.clk(gclk));
	jand g18794(.dina(n19047),.dinb(n18836),.dout(n19048),.clk(gclk));
	jand g18795(.dina(n19048),.dinb(w_n443_32[0]),.dout(n19049),.clk(gclk));
	jor g18796(.dina(w_n18803_0[1]),.dinb(n19049),.dout(n19050),.clk(gclk));
	jand g18797(.dina(n19050),.dinb(n18835),.dout(n19051),.clk(gclk));
	jand g18798(.dina(n19051),.dinb(w_n352_32[1]),.dout(n19052),.clk(gclk));
	jor g18799(.dina(w_n18811_0[0]),.dinb(n19052),.dout(n19053),.clk(gclk));
	jand g18800(.dina(n19053),.dinb(n18834),.dout(n19054),.clk(gclk));
	jand g18801(.dina(n19054),.dinb(w_n294_32[2]),.dout(n19055),.clk(gclk));
	jor g18802(.dina(w_n18819_0[0]),.dinb(n19055),.dout(n19056),.clk(gclk));
	jand g18803(.dina(n19056),.dinb(n18833),.dout(n19057),.clk(gclk));
	jand g18804(.dina(n19057),.dinb(w_n239_33[0]),.dout(n19058),.clk(gclk));
	jnot g18805(.din(w_n18827_0[0]),.dout(n19059),.clk(gclk));
	jor g18806(.dina(w_n19059_0[1]),.dinb(n19058),.dout(n19060),.clk(gclk));
	jand g18807(.dina(n19060),.dinb(n18832),.dout(n19061),.clk(gclk));
	jand g18808(.dina(n19061),.dinb(w_n221_33[0]),.dout(n19062),.clk(gclk));
	jxor g18809(.dina(w_n18148_0[0]),.dinb(w_n239_32[2]),.dout(n19063),.clk(gclk));
	jand g18810(.dina(n19063),.dinb(w_asqrt10_14[2]),.dout(n19064),.clk(gclk));
	jxor g18811(.dina(n19064),.dinb(w_n18153_0[0]),.dout(n19065),.clk(gclk));
	jor g18812(.dina(w_n19065_0[2]),.dinb(n19062),.dout(n19066),.clk(gclk));
	jand g18813(.dina(n19066),.dinb(n18831),.dout(n19067),.clk(gclk));
	jor g18814(.dina(w_n19067_0[1]),.dinb(w_n18183_0[1]),.dout(n19068),.clk(gclk));
	jand g18815(.dina(w_n18178_0[0]),.dinb(w_n18435_0[0]),.dout(n19069),.clk(gclk));
	jor g18816(.dina(n19069),.dinb(w_n18164_0[0]),.dout(n19070),.clk(gclk));
	jor g18817(.dina(w_n19070_0[1]),.dinb(w_n19068_0[1]),.dout(n19071),.clk(gclk));
	jand g18818(.dina(n19071),.dinb(w_n218_14[0]),.dout(n19072),.clk(gclk));
	jand g18819(.dina(w_n18442_11[2]),.dinb(w_n17773_0[0]),.dout(n19073),.clk(gclk));
	jand g18820(.dina(w_n19067_0[0]),.dinb(w_n18183_0[0]),.dout(n19074),.clk(gclk));
	jor g18821(.dina(w_n19074_0[2]),.dinb(w_n19073_0[1]),.dout(n19075),.clk(gclk));
	jand g18822(.dina(w_n18441_0[0]),.dinb(w_n18163_0[0]),.dout(n19076),.clk(gclk));
	jnot g18823(.din(n19076),.dout(n19077),.clk(gclk));
	jand g18824(.dina(w_n18172_0[0]),.dinb(w_asqrt63_24[0]),.dout(n19078),.clk(gclk));
	jand g18825(.dina(n19078),.dinb(w_n18195_0[0]),.dout(n19079),.clk(gclk));
	jand g18826(.dina(w_n19079_0[1]),.dinb(n19077),.dout(n19080),.clk(gclk));
	jor g18827(.dina(w_n19080_0[1]),.dinb(n19075),.dout(n19081),.clk(gclk));
	jor g18828(.dina(n19081),.dinb(w_n19072_0[1]),.dout(asqrt_fa_10),.clk(gclk));
	jor g18829(.dina(w_n18829_0[1]),.dinb(w_asqrt62_19[0]),.dout(n19083),.clk(gclk));
	jnot g18830(.din(w_n19065_0[1]),.dout(n19084),.clk(gclk));
	jand g18831(.dina(n19084),.dinb(n19083),.dout(n19085),.clk(gclk));
	jor g18832(.dina(n19085),.dinb(w_n18830_0[0]),.dout(n19086),.clk(gclk));
	jand g18833(.dina(w_n19086_0[2]),.dinb(w_n18182_1[0]),.dout(n19087),.clk(gclk));
	jnot g18834(.din(w_n19070_0[0]),.dout(n19088),.clk(gclk));
	jand g18835(.dina(n19088),.dinb(w_n19087_0[1]),.dout(n19089),.clk(gclk));
	jor g18836(.dina(n19089),.dinb(w_asqrt63_23[2]),.dout(n19090),.clk(gclk));
	jnot g18837(.din(w_n19073_0[0]),.dout(n19091),.clk(gclk));
	jor g18838(.dina(w_n19086_0[1]),.dinb(w_n18182_0[2]),.dout(n19092),.clk(gclk));
	jand g18839(.dina(n19092),.dinb(n19091),.dout(n19093),.clk(gclk));
	jnot g18840(.din(w_n19080_0[0]),.dout(n19094),.clk(gclk));
	jand g18841(.dina(n19094),.dinb(n19093),.dout(n19095),.clk(gclk));
	jand g18842(.dina(n19095),.dinb(n19090),.dout(n19096),.clk(gclk));
	jxor g18843(.dina(w_n18829_0[0]),.dinb(w_n221_32[2]),.dout(n19097),.clk(gclk));
	jor g18844(.dina(n19097),.dinb(w_n19096_36[1]),.dout(n19098),.clk(gclk));
	jxor g18845(.dina(n19098),.dinb(w_n19065_0[0]),.dout(n19099),.clk(gclk));
	jnot g18846(.din(w_n19099_0[2]),.dout(n19100),.clk(gclk));
	jnot g18847(.din(w_a16_0[2]),.dout(n19101),.clk(gclk));
	jnot g18848(.din(w_a17_0[1]),.dout(n19102),.clk(gclk));
	jand g18849(.dina(w_n19102_0[1]),.dinb(w_n19101_1[2]),.dout(n19103),.clk(gclk));
	jand g18850(.dina(w_n19103_0[2]),.dinb(w_n18185_1[0]),.dout(n19104),.clk(gclk));
	jnot g18851(.din(w_n19104_0[1]),.dout(n19105),.clk(gclk));
	jor g18852(.dina(w_n19096_36[0]),.dinb(w_n18185_0[2]),.dout(n19106),.clk(gclk));
	jand g18853(.dina(n19106),.dinb(n19105),.dout(n19107),.clk(gclk));
	jor g18854(.dina(w_n19107_0[2]),.dinb(w_n18442_11[1]),.dout(n19108),.clk(gclk));
	jand g18855(.dina(w_n19107_0[1]),.dinb(w_n18442_11[0]),.dout(n19109),.clk(gclk));
	jor g18856(.dina(w_n19096_35[2]),.dinb(w_a18_1[0]),.dout(n19110),.clk(gclk));
	jand g18857(.dina(n19110),.dinb(w_a19_0[0]),.dout(n19111),.clk(gclk));
	jand g18858(.dina(w_asqrt9_8),.dinb(w_n18187_0[1]),.dout(n19112),.clk(gclk));
	jor g18859(.dina(n19112),.dinb(n19111),.dout(n19113),.clk(gclk));
	jor g18860(.dina(w_n19113_0[1]),.dinb(n19109),.dout(n19114),.clk(gclk));
	jand g18861(.dina(n19114),.dinb(w_n19108_0[1]),.dout(n19115),.clk(gclk));
	jor g18862(.dina(w_n19115_0[2]),.dinb(w_n17769_20[0]),.dout(n19116),.clk(gclk));
	jand g18863(.dina(w_n19115_0[1]),.dinb(w_n17769_19[2]),.dout(n19117),.clk(gclk));
	jnot g18864(.din(w_n18187_0[0]),.dout(n19118),.clk(gclk));
	jor g18865(.dina(w_n19096_35[1]),.dinb(n19118),.dout(n19119),.clk(gclk));
	jor g18866(.dina(w_n19079_0[0]),.dinb(w_n18442_10[2]),.dout(n19120),.clk(gclk));
	jor g18867(.dina(n19120),.dinb(w_n19074_0[1]),.dout(n19121),.clk(gclk));
	jor g18868(.dina(n19121),.dinb(w_n19072_0[0]),.dout(n19122),.clk(gclk));
	jand g18869(.dina(n19122),.dinb(w_n19119_0[1]),.dout(n19123),.clk(gclk));
	jxor g18870(.dina(n19123),.dinb(w_n17774_0[1]),.dout(n19124),.clk(gclk));
	jor g18871(.dina(w_n19124_0[2]),.dinb(n19117),.dout(n19125),.clk(gclk));
	jand g18872(.dina(n19125),.dinb(w_n19116_0[1]),.dout(n19126),.clk(gclk));
	jor g18873(.dina(w_n19126_0[2]),.dinb(w_n17134_12[1]),.dout(n19127),.clk(gclk));
	jand g18874(.dina(w_n19126_0[1]),.dinb(w_n17134_12[0]),.dout(n19128),.clk(gclk));
	jxor g18875(.dina(w_n18189_0[0]),.dinb(w_n17769_19[1]),.dout(n19129),.clk(gclk));
	jor g18876(.dina(n19129),.dinb(w_n19096_35[0]),.dout(n19130),.clk(gclk));
	jxor g18877(.dina(n19130),.dinb(w_n18890_0[0]),.dout(n19131),.clk(gclk));
	jnot g18878(.din(w_n19131_0[2]),.dout(n19132),.clk(gclk));
	jor g18879(.dina(n19132),.dinb(n19128),.dout(n19133),.clk(gclk));
	jand g18880(.dina(n19133),.dinb(w_n19127_0[1]),.dout(n19134),.clk(gclk));
	jor g18881(.dina(w_n19134_0[2]),.dinb(w_n16489_20[1]),.dout(n19135),.clk(gclk));
	jand g18882(.dina(w_n19134_0[1]),.dinb(w_n16489_20[0]),.dout(n19136),.clk(gclk));
	jxor g18883(.dina(w_n18446_0[0]),.dinb(w_n17134_11[2]),.dout(n19137),.clk(gclk));
	jor g18884(.dina(n19137),.dinb(w_n19096_34[2]),.dout(n19138),.clk(gclk));
	jxor g18885(.dina(n19138),.dinb(w_n18455_0[0]),.dout(n19139),.clk(gclk));
	jor g18886(.dina(w_n19139_0[2]),.dinb(n19136),.dout(n19140),.clk(gclk));
	jand g18887(.dina(n19140),.dinb(w_n19135_0[1]),.dout(n19141),.clk(gclk));
	jor g18888(.dina(w_n19141_0[2]),.dinb(w_n15878_13[1]),.dout(n19142),.clk(gclk));
	jand g18889(.dina(w_n19141_0[1]),.dinb(w_n15878_13[0]),.dout(n19143),.clk(gclk));
	jxor g18890(.dina(w_n18457_0[0]),.dinb(w_n16489_19[2]),.dout(n19144),.clk(gclk));
	jor g18891(.dina(n19144),.dinb(w_n19096_34[1]),.dout(n19145),.clk(gclk));
	jxor g18892(.dina(n19145),.dinb(w_n18897_0[0]),.dout(n19146),.clk(gclk));
	jnot g18893(.din(w_n19146_0[2]),.dout(n19147),.clk(gclk));
	jor g18894(.dina(n19147),.dinb(n19143),.dout(n19148),.clk(gclk));
	jand g18895(.dina(n19148),.dinb(w_n19142_0[1]),.dout(n19149),.clk(gclk));
	jor g18896(.dina(w_n19149_0[2]),.dinb(w_n15260_21[0]),.dout(n19150),.clk(gclk));
	jand g18897(.dina(w_n19149_0[1]),.dinb(w_n15260_20[2]),.dout(n19151),.clk(gclk));
	jxor g18898(.dina(w_n18464_0[0]),.dinb(w_n15878_12[2]),.dout(n19152),.clk(gclk));
	jor g18899(.dina(n19152),.dinb(w_n19096_34[0]),.dout(n19153),.clk(gclk));
	jxor g18900(.dina(n19153),.dinb(w_n18470_0[0]),.dout(n19154),.clk(gclk));
	jor g18901(.dina(w_n19154_0[2]),.dinb(n19151),.dout(n19155),.clk(gclk));
	jand g18902(.dina(n19155),.dinb(w_n19150_0[1]),.dout(n19156),.clk(gclk));
	jor g18903(.dina(w_n19156_0[2]),.dinb(w_n14674_14[0]),.dout(n19157),.clk(gclk));
	jand g18904(.dina(w_n19156_0[1]),.dinb(w_n14674_13[2]),.dout(n19158),.clk(gclk));
	jxor g18905(.dina(w_n18472_0[0]),.dinb(w_n15260_20[1]),.dout(n19159),.clk(gclk));
	jor g18906(.dina(n19159),.dinb(w_n19096_33[2]),.dout(n19160),.clk(gclk));
	jxor g18907(.dina(n19160),.dinb(w_n18904_0[0]),.dout(n19161),.clk(gclk));
	jnot g18908(.din(w_n19161_0[2]),.dout(n19162),.clk(gclk));
	jor g18909(.dina(n19162),.dinb(n19158),.dout(n19163),.clk(gclk));
	jand g18910(.dina(n19163),.dinb(w_n19157_0[1]),.dout(n19164),.clk(gclk));
	jor g18911(.dina(w_n19164_0[2]),.dinb(w_n14078_21[1]),.dout(n19165),.clk(gclk));
	jand g18912(.dina(w_n19164_0[1]),.dinb(w_n14078_21[0]),.dout(n19166),.clk(gclk));
	jxor g18913(.dina(w_n18479_0[0]),.dinb(w_n14674_13[1]),.dout(n19167),.clk(gclk));
	jor g18914(.dina(n19167),.dinb(w_n19096_33[1]),.dout(n19168),.clk(gclk));
	jxor g18915(.dina(n19168),.dinb(w_n18485_0[0]),.dout(n19169),.clk(gclk));
	jor g18916(.dina(w_n19169_0[2]),.dinb(n19166),.dout(n19170),.clk(gclk));
	jand g18917(.dina(n19170),.dinb(w_n19165_0[1]),.dout(n19171),.clk(gclk));
	jor g18918(.dina(w_n19171_0[2]),.dinb(w_n13515_15[0]),.dout(n19172),.clk(gclk));
	jand g18919(.dina(w_n19171_0[1]),.dinb(w_n13515_14[2]),.dout(n19173),.clk(gclk));
	jxor g18920(.dina(w_n18487_0[0]),.dinb(w_n14078_20[2]),.dout(n19174),.clk(gclk));
	jor g18921(.dina(n19174),.dinb(w_n19096_33[0]),.dout(n19175),.clk(gclk));
	jxor g18922(.dina(n19175),.dinb(w_n18911_0[0]),.dout(n19176),.clk(gclk));
	jnot g18923(.din(w_n19176_0[2]),.dout(n19177),.clk(gclk));
	jor g18924(.dina(n19177),.dinb(n19173),.dout(n19178),.clk(gclk));
	jand g18925(.dina(n19178),.dinb(w_n19172_0[1]),.dout(n19179),.clk(gclk));
	jor g18926(.dina(w_n19179_0[2]),.dinb(w_n12947_22[0]),.dout(n19180),.clk(gclk));
	jand g18927(.dina(w_n19179_0[1]),.dinb(w_n12947_21[2]),.dout(n19181),.clk(gclk));
	jxor g18928(.dina(w_n18494_0[0]),.dinb(w_n13515_14[1]),.dout(n19182),.clk(gclk));
	jor g18929(.dina(n19182),.dinb(w_n19096_32[2]),.dout(n19183),.clk(gclk));
	jxor g18930(.dina(n19183),.dinb(w_n18500_0[0]),.dout(n19184),.clk(gclk));
	jor g18931(.dina(w_n19184_0[2]),.dinb(n19181),.dout(n19185),.clk(gclk));
	jand g18932(.dina(n19185),.dinb(w_n19180_0[1]),.dout(n19186),.clk(gclk));
	jor g18933(.dina(w_n19186_0[2]),.dinb(w_n12410_15[2]),.dout(n19187),.clk(gclk));
	jand g18934(.dina(w_n19186_0[1]),.dinb(w_n12410_15[1]),.dout(n19188),.clk(gclk));
	jxor g18935(.dina(w_n18502_0[0]),.dinb(w_n12947_21[1]),.dout(n19189),.clk(gclk));
	jor g18936(.dina(n19189),.dinb(w_n19096_32[1]),.dout(n19190),.clk(gclk));
	jxor g18937(.dina(n19190),.dinb(w_n18918_0[0]),.dout(n19191),.clk(gclk));
	jnot g18938(.din(w_n19191_0[2]),.dout(n19192),.clk(gclk));
	jor g18939(.dina(n19192),.dinb(n19188),.dout(n19193),.clk(gclk));
	jand g18940(.dina(n19193),.dinb(w_n19187_0[1]),.dout(n19194),.clk(gclk));
	jor g18941(.dina(w_n19194_0[2]),.dinb(w_n11858_22[1]),.dout(n19195),.clk(gclk));
	jand g18942(.dina(w_n19194_0[1]),.dinb(w_n11858_22[0]),.dout(n19196),.clk(gclk));
	jxor g18943(.dina(w_n18509_0[0]),.dinb(w_n12410_15[0]),.dout(n19197),.clk(gclk));
	jor g18944(.dina(n19197),.dinb(w_n19096_32[0]),.dout(n19198),.clk(gclk));
	jxor g18945(.dina(n19198),.dinb(w_n18515_0[0]),.dout(n19199),.clk(gclk));
	jor g18946(.dina(w_n19199_0[2]),.dinb(n19196),.dout(n19200),.clk(gclk));
	jand g18947(.dina(n19200),.dinb(w_n19195_0[1]),.dout(n19201),.clk(gclk));
	jor g18948(.dina(w_n19201_0[2]),.dinb(w_n11347_16[1]),.dout(n19202),.clk(gclk));
	jand g18949(.dina(w_n19201_0[1]),.dinb(w_n11347_16[0]),.dout(n19203),.clk(gclk));
	jxor g18950(.dina(w_n18517_0[0]),.dinb(w_n11858_21[2]),.dout(n19204),.clk(gclk));
	jor g18951(.dina(n19204),.dinb(w_n19096_31[2]),.dout(n19205),.clk(gclk));
	jxor g18952(.dina(n19205),.dinb(w_n18523_0[0]),.dout(n19206),.clk(gclk));
	jor g18953(.dina(w_n19206_0[2]),.dinb(n19203),.dout(n19207),.clk(gclk));
	jand g18954(.dina(n19207),.dinb(w_n19202_0[1]),.dout(n19208),.clk(gclk));
	jor g18955(.dina(w_n19208_0[2]),.dinb(w_n10824_23[0]),.dout(n19209),.clk(gclk));
	jand g18956(.dina(w_n19208_0[1]),.dinb(w_n10824_22[2]),.dout(n19210),.clk(gclk));
	jxor g18957(.dina(w_n18525_0[0]),.dinb(w_n11347_15[2]),.dout(n19211),.clk(gclk));
	jor g18958(.dina(n19211),.dinb(w_n19096_31[1]),.dout(n19212),.clk(gclk));
	jxor g18959(.dina(n19212),.dinb(w_n18928_0[0]),.dout(n19213),.clk(gclk));
	jnot g18960(.din(w_n19213_0[2]),.dout(n19214),.clk(gclk));
	jor g18961(.dina(n19214),.dinb(n19210),.dout(n19215),.clk(gclk));
	jand g18962(.dina(n19215),.dinb(w_n19209_0[1]),.dout(n19216),.clk(gclk));
	jor g18963(.dina(w_n19216_0[2]),.dinb(w_n10328_17[1]),.dout(n19217),.clk(gclk));
	jand g18964(.dina(w_n19216_0[1]),.dinb(w_n10328_17[0]),.dout(n19218),.clk(gclk));
	jxor g18965(.dina(w_n18532_0[0]),.dinb(w_n10824_22[1]),.dout(n19219),.clk(gclk));
	jor g18966(.dina(n19219),.dinb(w_n19096_31[0]),.dout(n19220),.clk(gclk));
	jxor g18967(.dina(n19220),.dinb(w_n18932_0[0]),.dout(n19221),.clk(gclk));
	jnot g18968(.din(w_n19221_0[2]),.dout(n19222),.clk(gclk));
	jor g18969(.dina(n19222),.dinb(n19218),.dout(n19223),.clk(gclk));
	jand g18970(.dina(n19223),.dinb(w_n19217_0[1]),.dout(n19224),.clk(gclk));
	jor g18971(.dina(w_n19224_0[2]),.dinb(w_n9832_23[2]),.dout(n19225),.clk(gclk));
	jand g18972(.dina(w_n19224_0[1]),.dinb(w_n9832_23[1]),.dout(n19226),.clk(gclk));
	jxor g18973(.dina(w_n18539_0[0]),.dinb(w_n10328_16[2]),.dout(n19227),.clk(gclk));
	jor g18974(.dina(n19227),.dinb(w_n19096_30[2]),.dout(n19228),.clk(gclk));
	jxor g18975(.dina(n19228),.dinb(w_n18545_0[0]),.dout(n19229),.clk(gclk));
	jor g18976(.dina(w_n19229_0[2]),.dinb(n19226),.dout(n19230),.clk(gclk));
	jand g18977(.dina(n19230),.dinb(w_n19225_0[1]),.dout(n19231),.clk(gclk));
	jor g18978(.dina(w_n19231_0[2]),.dinb(w_n9369_18[1]),.dout(n19232),.clk(gclk));
	jand g18979(.dina(w_n19231_0[1]),.dinb(w_n9369_18[0]),.dout(n19233),.clk(gclk));
	jxor g18980(.dina(w_n18547_0[0]),.dinb(w_n9832_23[0]),.dout(n19234),.clk(gclk));
	jor g18981(.dina(n19234),.dinb(w_n19096_30[1]),.dout(n19235),.clk(gclk));
	jxor g18982(.dina(n19235),.dinb(w_n18939_0[0]),.dout(n19236),.clk(gclk));
	jnot g18983(.din(w_n19236_0[2]),.dout(n19237),.clk(gclk));
	jor g18984(.dina(n19237),.dinb(n19233),.dout(n19238),.clk(gclk));
	jand g18985(.dina(n19238),.dinb(w_n19232_0[1]),.dout(n19239),.clk(gclk));
	jor g18986(.dina(w_n19239_0[2]),.dinb(w_n8890_24[0]),.dout(n19240),.clk(gclk));
	jand g18987(.dina(w_n19239_0[1]),.dinb(w_n8890_23[2]),.dout(n19241),.clk(gclk));
	jxor g18988(.dina(w_n18554_0[0]),.dinb(w_n9369_17[2]),.dout(n19242),.clk(gclk));
	jor g18989(.dina(n19242),.dinb(w_n19096_30[0]),.dout(n19243),.clk(gclk));
	jxor g18990(.dina(n19243),.dinb(w_n18560_0[0]),.dout(n19244),.clk(gclk));
	jor g18991(.dina(w_n19244_0[2]),.dinb(n19241),.dout(n19245),.clk(gclk));
	jand g18992(.dina(n19245),.dinb(w_n19240_0[1]),.dout(n19246),.clk(gclk));
	jor g18993(.dina(w_n19246_0[2]),.dinb(w_n8449_19[0]),.dout(n19247),.clk(gclk));
	jand g18994(.dina(w_n19246_0[1]),.dinb(w_n8449_18[2]),.dout(n19248),.clk(gclk));
	jxor g18995(.dina(w_n18562_0[0]),.dinb(w_n8890_23[1]),.dout(n19249),.clk(gclk));
	jor g18996(.dina(n19249),.dinb(w_n19096_29[2]),.dout(n19250),.clk(gclk));
	jxor g18997(.dina(n19250),.dinb(w_n18946_0[0]),.dout(n19251),.clk(gclk));
	jnot g18998(.din(w_n19251_0[2]),.dout(n19252),.clk(gclk));
	jor g18999(.dina(n19252),.dinb(n19248),.dout(n19253),.clk(gclk));
	jand g19000(.dina(n19253),.dinb(w_n19247_0[1]),.dout(n19254),.clk(gclk));
	jor g19001(.dina(w_n19254_0[2]),.dinb(w_n8003_24[2]),.dout(n19255),.clk(gclk));
	jand g19002(.dina(w_n19254_0[1]),.dinb(w_n8003_24[1]),.dout(n19256),.clk(gclk));
	jxor g19003(.dina(w_n18569_0[0]),.dinb(w_n8449_18[1]),.dout(n19257),.clk(gclk));
	jor g19004(.dina(n19257),.dinb(w_n19096_29[1]),.dout(n19258),.clk(gclk));
	jxor g19005(.dina(n19258),.dinb(w_n18575_0[0]),.dout(n19259),.clk(gclk));
	jor g19006(.dina(w_n19259_0[2]),.dinb(n19256),.dout(n19260),.clk(gclk));
	jand g19007(.dina(n19260),.dinb(w_n19255_0[1]),.dout(n19261),.clk(gclk));
	jor g19008(.dina(w_n19261_0[2]),.dinb(w_n7581_20[0]),.dout(n19262),.clk(gclk));
	jand g19009(.dina(w_n19261_0[1]),.dinb(w_n7581_19[2]),.dout(n19263),.clk(gclk));
	jxor g19010(.dina(w_n18577_0[0]),.dinb(w_n8003_24[0]),.dout(n19264),.clk(gclk));
	jor g19011(.dina(n19264),.dinb(w_n19096_29[0]),.dout(n19265),.clk(gclk));
	jxor g19012(.dina(n19265),.dinb(w_n18583_0[0]),.dout(n19266),.clk(gclk));
	jor g19013(.dina(w_n19266_0[2]),.dinb(n19263),.dout(n19267),.clk(gclk));
	jand g19014(.dina(n19267),.dinb(w_n19262_0[1]),.dout(n19268),.clk(gclk));
	jor g19015(.dina(w_n19268_0[2]),.dinb(w_n7154_25[0]),.dout(n19269),.clk(gclk));
	jand g19016(.dina(w_n19268_0[1]),.dinb(w_n7154_24[2]),.dout(n19270),.clk(gclk));
	jxor g19017(.dina(w_n18585_0[0]),.dinb(w_n7581_19[1]),.dout(n19271),.clk(gclk));
	jor g19018(.dina(n19271),.dinb(w_n19096_28[2]),.dout(n19272),.clk(gclk));
	jxor g19019(.dina(n19272),.dinb(w_n18591_0[0]),.dout(n19273),.clk(gclk));
	jor g19020(.dina(w_n19273_0[2]),.dinb(n19270),.dout(n19274),.clk(gclk));
	jand g19021(.dina(n19274),.dinb(w_n19269_0[1]),.dout(n19275),.clk(gclk));
	jor g19022(.dina(w_n19275_0[2]),.dinb(w_n6758_20[2]),.dout(n19276),.clk(gclk));
	jand g19023(.dina(w_n19275_0[1]),.dinb(w_n6758_20[1]),.dout(n19277),.clk(gclk));
	jxor g19024(.dina(w_n18593_0[0]),.dinb(w_n7154_24[1]),.dout(n19278),.clk(gclk));
	jor g19025(.dina(n19278),.dinb(w_n19096_28[1]),.dout(n19279),.clk(gclk));
	jxor g19026(.dina(n19279),.dinb(w_n18959_0[0]),.dout(n19280),.clk(gclk));
	jnot g19027(.din(w_n19280_0[2]),.dout(n19281),.clk(gclk));
	jor g19028(.dina(n19281),.dinb(n19277),.dout(n19282),.clk(gclk));
	jand g19029(.dina(n19282),.dinb(w_n19276_0[1]),.dout(n19283),.clk(gclk));
	jor g19030(.dina(w_n19283_0[2]),.dinb(w_n6357_25[1]),.dout(n19284),.clk(gclk));
	jand g19031(.dina(w_n19283_0[1]),.dinb(w_n6357_25[0]),.dout(n19285),.clk(gclk));
	jxor g19032(.dina(w_n18600_0[0]),.dinb(w_n6758_20[0]),.dout(n19286),.clk(gclk));
	jor g19033(.dina(n19286),.dinb(w_n19096_28[0]),.dout(n19287),.clk(gclk));
	jxor g19034(.dina(n19287),.dinb(w_n18606_0[0]),.dout(n19288),.clk(gclk));
	jor g19035(.dina(w_n19288_0[2]),.dinb(n19285),.dout(n19289),.clk(gclk));
	jand g19036(.dina(n19289),.dinb(w_n19284_0[1]),.dout(n19290),.clk(gclk));
	jor g19037(.dina(w_n19290_0[2]),.dinb(w_n5989_21[1]),.dout(n19291),.clk(gclk));
	jand g19038(.dina(w_n19290_0[1]),.dinb(w_n5989_21[0]),.dout(n19292),.clk(gclk));
	jxor g19039(.dina(w_n18608_0[0]),.dinb(w_n6357_24[2]),.dout(n19293),.clk(gclk));
	jor g19040(.dina(n19293),.dinb(w_n19096_27[2]),.dout(n19294),.clk(gclk));
	jxor g19041(.dina(n19294),.dinb(w_n18966_0[0]),.dout(n19295),.clk(gclk));
	jnot g19042(.din(w_n19295_0[2]),.dout(n19296),.clk(gclk));
	jor g19043(.dina(n19296),.dinb(n19292),.dout(n19297),.clk(gclk));
	jand g19044(.dina(n19297),.dinb(w_n19291_0[1]),.dout(n19298),.clk(gclk));
	jor g19045(.dina(w_n19298_0[2]),.dinb(w_n5606_25[2]),.dout(n19299),.clk(gclk));
	jand g19046(.dina(w_n19298_0[1]),.dinb(w_n5606_25[1]),.dout(n19300),.clk(gclk));
	jxor g19047(.dina(w_n18615_0[0]),.dinb(w_n5989_20[2]),.dout(n19301),.clk(gclk));
	jor g19048(.dina(n19301),.dinb(w_n19096_27[1]),.dout(n19302),.clk(gclk));
	jxor g19049(.dina(n19302),.dinb(w_n18621_0[0]),.dout(n19303),.clk(gclk));
	jor g19050(.dina(w_n19303_0[2]),.dinb(n19300),.dout(n19304),.clk(gclk));
	jand g19051(.dina(n19304),.dinb(w_n19299_0[1]),.dout(n19305),.clk(gclk));
	jor g19052(.dina(w_n19305_0[2]),.dinb(w_n5259_22[1]),.dout(n19306),.clk(gclk));
	jand g19053(.dina(w_n19305_0[1]),.dinb(w_n5259_22[0]),.dout(n19307),.clk(gclk));
	jxor g19054(.dina(w_n18623_0[0]),.dinb(w_n5606_25[0]),.dout(n19308),.clk(gclk));
	jor g19055(.dina(n19308),.dinb(w_n19096_27[0]),.dout(n19309),.clk(gclk));
	jxor g19056(.dina(n19309),.dinb(w_n18973_0[0]),.dout(n19310),.clk(gclk));
	jnot g19057(.din(w_n19310_0[2]),.dout(n19311),.clk(gclk));
	jor g19058(.dina(n19311),.dinb(n19307),.dout(n19312),.clk(gclk));
	jand g19059(.dina(n19312),.dinb(w_n19306_0[1]),.dout(n19313),.clk(gclk));
	jor g19060(.dina(w_n19313_0[2]),.dinb(w_n4902_26[1]),.dout(n19314),.clk(gclk));
	jand g19061(.dina(w_n19313_0[1]),.dinb(w_n4902_26[0]),.dout(n19315),.clk(gclk));
	jxor g19062(.dina(w_n18630_0[0]),.dinb(w_n5259_21[2]),.dout(n19316),.clk(gclk));
	jor g19063(.dina(n19316),.dinb(w_n19096_26[2]),.dout(n19317),.clk(gclk));
	jxor g19064(.dina(n19317),.dinb(w_n18636_0[0]),.dout(n19318),.clk(gclk));
	jor g19065(.dina(w_n19318_0[2]),.dinb(n19315),.dout(n19319),.clk(gclk));
	jand g19066(.dina(n19319),.dinb(w_n19314_0[1]),.dout(n19320),.clk(gclk));
	jor g19067(.dina(w_n19320_0[2]),.dinb(w_n4582_23[1]),.dout(n19321),.clk(gclk));
	jand g19068(.dina(w_n19320_0[1]),.dinb(w_n4582_23[0]),.dout(n19322),.clk(gclk));
	jxor g19069(.dina(w_n18638_0[0]),.dinb(w_n4902_25[2]),.dout(n19323),.clk(gclk));
	jor g19070(.dina(n19323),.dinb(w_n19096_26[1]),.dout(n19324),.clk(gclk));
	jxor g19071(.dina(n19324),.dinb(w_n18980_0[0]),.dout(n19325),.clk(gclk));
	jnot g19072(.din(w_n19325_0[2]),.dout(n19326),.clk(gclk));
	jor g19073(.dina(n19326),.dinb(n19322),.dout(n19327),.clk(gclk));
	jand g19074(.dina(n19327),.dinb(w_n19321_0[1]),.dout(n19328),.clk(gclk));
	jor g19075(.dina(w_n19328_0[2]),.dinb(w_n4249_27[0]),.dout(n19329),.clk(gclk));
	jand g19076(.dina(w_n19328_0[1]),.dinb(w_n4249_26[2]),.dout(n19330),.clk(gclk));
	jxor g19077(.dina(w_n18645_0[0]),.dinb(w_n4582_22[2]),.dout(n19331),.clk(gclk));
	jor g19078(.dina(n19331),.dinb(w_n19096_26[0]),.dout(n19332),.clk(gclk));
	jxor g19079(.dina(n19332),.dinb(w_n18651_0[0]),.dout(n19333),.clk(gclk));
	jor g19080(.dina(w_n19333_0[2]),.dinb(n19330),.dout(n19334),.clk(gclk));
	jand g19081(.dina(n19334),.dinb(w_n19329_0[1]),.dout(n19335),.clk(gclk));
	jor g19082(.dina(w_n19335_0[2]),.dinb(w_n3955_24[0]),.dout(n19336),.clk(gclk));
	jand g19083(.dina(w_n19335_0[1]),.dinb(w_n3955_23[2]),.dout(n19337),.clk(gclk));
	jxor g19084(.dina(w_n18653_0[0]),.dinb(w_n4249_26[1]),.dout(n19338),.clk(gclk));
	jor g19085(.dina(n19338),.dinb(w_n19096_25[2]),.dout(n19339),.clk(gclk));
	jxor g19086(.dina(n19339),.dinb(w_n18659_0[0]),.dout(n19340),.clk(gclk));
	jor g19087(.dina(w_n19340_0[2]),.dinb(n19337),.dout(n19341),.clk(gclk));
	jand g19088(.dina(n19341),.dinb(w_n19336_0[1]),.dout(n19342),.clk(gclk));
	jor g19089(.dina(w_n19342_0[2]),.dinb(w_n3642_27[1]),.dout(n19343),.clk(gclk));
	jand g19090(.dina(w_n19342_0[1]),.dinb(w_n3642_27[0]),.dout(n19344),.clk(gclk));
	jxor g19091(.dina(w_n18661_0[0]),.dinb(w_n3955_23[1]),.dout(n19345),.clk(gclk));
	jor g19092(.dina(n19345),.dinb(w_n19096_25[1]),.dout(n19346),.clk(gclk));
	jxor g19093(.dina(n19346),.dinb(w_n18667_0[0]),.dout(n19347),.clk(gclk));
	jor g19094(.dina(w_n19347_0[2]),.dinb(n19344),.dout(n19348),.clk(gclk));
	jand g19095(.dina(n19348),.dinb(w_n19343_0[1]),.dout(n19349),.clk(gclk));
	jor g19096(.dina(w_n19349_0[2]),.dinb(w_n3368_24[2]),.dout(n19350),.clk(gclk));
	jand g19097(.dina(w_n19349_0[1]),.dinb(w_n3368_24[1]),.dout(n19351),.clk(gclk));
	jxor g19098(.dina(w_n18669_0[0]),.dinb(w_n3642_26[2]),.dout(n19352),.clk(gclk));
	jor g19099(.dina(n19352),.dinb(w_n19096_25[0]),.dout(n19353),.clk(gclk));
	jxor g19100(.dina(n19353),.dinb(w_n18993_0[0]),.dout(n19354),.clk(gclk));
	jnot g19101(.din(w_n19354_0[2]),.dout(n19355),.clk(gclk));
	jor g19102(.dina(n19355),.dinb(n19351),.dout(n19356),.clk(gclk));
	jand g19103(.dina(n19356),.dinb(w_n19350_0[1]),.dout(n19357),.clk(gclk));
	jor g19104(.dina(w_n19357_0[2]),.dinb(w_n3089_28[0]),.dout(n19358),.clk(gclk));
	jand g19105(.dina(w_n19357_0[1]),.dinb(w_n3089_27[2]),.dout(n19359),.clk(gclk));
	jxor g19106(.dina(w_n18676_0[0]),.dinb(w_n3368_24[0]),.dout(n19360),.clk(gclk));
	jor g19107(.dina(n19360),.dinb(w_n19096_24[2]),.dout(n19361),.clk(gclk));
	jxor g19108(.dina(n19361),.dinb(w_n18682_0[0]),.dout(n19362),.clk(gclk));
	jor g19109(.dina(w_n19362_0[2]),.dinb(n19359),.dout(n19363),.clk(gclk));
	jand g19110(.dina(n19363),.dinb(w_n19358_0[1]),.dout(n19364),.clk(gclk));
	jor g19111(.dina(w_n19364_0[2]),.dinb(w_n2833_25[2]),.dout(n19365),.clk(gclk));
	jand g19112(.dina(w_n19364_0[1]),.dinb(w_n2833_25[1]),.dout(n19366),.clk(gclk));
	jxor g19113(.dina(w_n18684_0[0]),.dinb(w_n3089_27[1]),.dout(n19367),.clk(gclk));
	jor g19114(.dina(n19367),.dinb(w_n19096_24[1]),.dout(n19368),.clk(gclk));
	jxor g19115(.dina(n19368),.dinb(w_n18690_0[0]),.dout(n19369),.clk(gclk));
	jor g19116(.dina(w_n19369_0[2]),.dinb(n19366),.dout(n19370),.clk(gclk));
	jand g19117(.dina(n19370),.dinb(w_n19365_0[1]),.dout(n19371),.clk(gclk));
	jor g19118(.dina(w_n19371_0[2]),.dinb(w_n2572_28[1]),.dout(n19372),.clk(gclk));
	jand g19119(.dina(w_n19371_0[1]),.dinb(w_n2572_28[0]),.dout(n19373),.clk(gclk));
	jxor g19120(.dina(w_n18692_0[0]),.dinb(w_n2833_25[0]),.dout(n19374),.clk(gclk));
	jor g19121(.dina(n19374),.dinb(w_n19096_24[0]),.dout(n19375),.clk(gclk));
	jxor g19122(.dina(n19375),.dinb(w_n18698_0[0]),.dout(n19376),.clk(gclk));
	jor g19123(.dina(w_n19376_0[2]),.dinb(n19373),.dout(n19377),.clk(gclk));
	jand g19124(.dina(n19377),.dinb(w_n19372_0[1]),.dout(n19378),.clk(gclk));
	jor g19125(.dina(w_n19378_0[2]),.dinb(w_n2345_26[1]),.dout(n19379),.clk(gclk));
	jand g19126(.dina(w_n19378_0[1]),.dinb(w_n2345_26[0]),.dout(n19380),.clk(gclk));
	jxor g19127(.dina(w_n18700_0[0]),.dinb(w_n2572_27[2]),.dout(n19381),.clk(gclk));
	jor g19128(.dina(n19381),.dinb(w_n19096_23[2]),.dout(n19382),.clk(gclk));
	jxor g19129(.dina(n19382),.dinb(w_n18706_0[0]),.dout(n19383),.clk(gclk));
	jor g19130(.dina(w_n19383_0[2]),.dinb(n19380),.dout(n19384),.clk(gclk));
	jand g19131(.dina(n19384),.dinb(w_n19379_0[1]),.dout(n19385),.clk(gclk));
	jor g19132(.dina(w_n19385_0[2]),.dinb(w_n2108_29[0]),.dout(n19386),.clk(gclk));
	jand g19133(.dina(w_n19385_0[1]),.dinb(w_n2108_28[2]),.dout(n19387),.clk(gclk));
	jxor g19134(.dina(w_n18708_0[0]),.dinb(w_n2345_25[2]),.dout(n19388),.clk(gclk));
	jor g19135(.dina(n19388),.dinb(w_n19096_23[1]),.dout(n19389),.clk(gclk));
	jxor g19136(.dina(n19389),.dinb(w_n18714_0[0]),.dout(n19390),.clk(gclk));
	jor g19137(.dina(w_n19390_0[2]),.dinb(n19387),.dout(n19391),.clk(gclk));
	jand g19138(.dina(n19391),.dinb(w_n19386_0[1]),.dout(n19392),.clk(gclk));
	jor g19139(.dina(w_n19392_0[2]),.dinb(w_n1912_27[1]),.dout(n19393),.clk(gclk));
	jand g19140(.dina(w_n19392_0[1]),.dinb(w_n1912_27[0]),.dout(n19394),.clk(gclk));
	jxor g19141(.dina(w_n18716_0[0]),.dinb(w_n2108_28[1]),.dout(n19395),.clk(gclk));
	jor g19142(.dina(n19395),.dinb(w_n19096_23[0]),.dout(n19396),.clk(gclk));
	jxor g19143(.dina(n19396),.dinb(w_n19012_0[0]),.dout(n19397),.clk(gclk));
	jnot g19144(.din(w_n19397_0[2]),.dout(n19398),.clk(gclk));
	jor g19145(.dina(n19398),.dinb(n19394),.dout(n19399),.clk(gclk));
	jand g19146(.dina(n19399),.dinb(w_n19393_0[1]),.dout(n19400),.clk(gclk));
	jor g19147(.dina(w_n19400_0[2]),.dinb(w_n1699_29[2]),.dout(n19401),.clk(gclk));
	jand g19148(.dina(w_n19400_0[1]),.dinb(w_n1699_29[1]),.dout(n19402),.clk(gclk));
	jxor g19149(.dina(w_n18723_0[0]),.dinb(w_n1912_26[2]),.dout(n19403),.clk(gclk));
	jor g19150(.dina(n19403),.dinb(w_n19096_22[2]),.dout(n19404),.clk(gclk));
	jxor g19151(.dina(n19404),.dinb(w_n18729_0[0]),.dout(n19405),.clk(gclk));
	jor g19152(.dina(w_n19405_0[2]),.dinb(n19402),.dout(n19406),.clk(gclk));
	jand g19153(.dina(n19406),.dinb(w_n19401_0[1]),.dout(n19407),.clk(gclk));
	jor g19154(.dina(w_n19407_0[2]),.dinb(w_n1516_28[0]),.dout(n19408),.clk(gclk));
	jand g19155(.dina(w_n19407_0[1]),.dinb(w_n1516_27[2]),.dout(n19409),.clk(gclk));
	jxor g19156(.dina(w_n18731_0[0]),.dinb(w_n1699_29[0]),.dout(n19410),.clk(gclk));
	jor g19157(.dina(n19410),.dinb(w_n19096_22[1]),.dout(n19411),.clk(gclk));
	jxor g19158(.dina(n19411),.dinb(w_n19019_0[0]),.dout(n19412),.clk(gclk));
	jnot g19159(.din(w_n19412_0[2]),.dout(n19413),.clk(gclk));
	jor g19160(.dina(n19413),.dinb(n19409),.dout(n19414),.clk(gclk));
	jand g19161(.dina(n19414),.dinb(w_n19408_0[1]),.dout(n19415),.clk(gclk));
	jor g19162(.dina(w_n19415_0[2]),.dinb(w_n1332_29[2]),.dout(n19416),.clk(gclk));
	jand g19163(.dina(w_n19415_0[1]),.dinb(w_n1332_29[1]),.dout(n19417),.clk(gclk));
	jxor g19164(.dina(w_n18738_0[0]),.dinb(w_n1516_27[1]),.dout(n19418),.clk(gclk));
	jor g19165(.dina(n19418),.dinb(w_n19096_22[0]),.dout(n19419),.clk(gclk));
	jxor g19166(.dina(n19419),.dinb(w_n18744_0[0]),.dout(n19420),.clk(gclk));
	jor g19167(.dina(w_n19420_0[2]),.dinb(n19417),.dout(n19421),.clk(gclk));
	jand g19168(.dina(n19421),.dinb(w_n19416_0[1]),.dout(n19422),.clk(gclk));
	jor g19169(.dina(w_n19422_0[2]),.dinb(w_n1173_28[2]),.dout(n19423),.clk(gclk));
	jand g19170(.dina(w_n19422_0[1]),.dinb(w_n1173_28[1]),.dout(n19424),.clk(gclk));
	jxor g19171(.dina(w_n18746_0[0]),.dinb(w_n1332_29[0]),.dout(n19425),.clk(gclk));
	jor g19172(.dina(n19425),.dinb(w_n19096_21[2]),.dout(n19426),.clk(gclk));
	jxor g19173(.dina(n19426),.dinb(w_n18752_0[0]),.dout(n19427),.clk(gclk));
	jor g19174(.dina(w_n19427_0[2]),.dinb(n19424),.dout(n19428),.clk(gclk));
	jand g19175(.dina(n19428),.dinb(w_n19423_0[1]),.dout(n19429),.clk(gclk));
	jor g19176(.dina(w_n19429_0[2]),.dinb(w_n1008_30[2]),.dout(n19430),.clk(gclk));
	jand g19177(.dina(w_n19429_0[1]),.dinb(w_n1008_30[1]),.dout(n19431),.clk(gclk));
	jxor g19178(.dina(w_n18754_0[0]),.dinb(w_n1173_28[0]),.dout(n19432),.clk(gclk));
	jor g19179(.dina(n19432),.dinb(w_n19096_21[1]),.dout(n19433),.clk(gclk));
	jxor g19180(.dina(n19433),.dinb(w_n19029_0[0]),.dout(n19434),.clk(gclk));
	jnot g19181(.din(w_n19434_0[2]),.dout(n19435),.clk(gclk));
	jor g19182(.dina(n19435),.dinb(n19431),.dout(n19436),.clk(gclk));
	jand g19183(.dina(n19436),.dinb(w_n19430_0[1]),.dout(n19437),.clk(gclk));
	jor g19184(.dina(w_n19437_0[2]),.dinb(w_n884_29[2]),.dout(n19438),.clk(gclk));
	jxor g19185(.dina(w_n18761_0[0]),.dinb(w_n1008_30[0]),.dout(n19439),.clk(gclk));
	jor g19186(.dina(n19439),.dinb(w_n19096_21[0]),.dout(n19440),.clk(gclk));
	jxor g19187(.dina(n19440),.dinb(w_n18841_0[0]),.dout(n19441),.clk(gclk));
	jnot g19188(.din(w_n19441_0[2]),.dout(n19442),.clk(gclk));
	jand g19189(.dina(w_n19437_0[1]),.dinb(w_n884_29[1]),.dout(n19443),.clk(gclk));
	jor g19190(.dina(n19443),.dinb(n19442),.dout(n19444),.clk(gclk));
	jand g19191(.dina(n19444),.dinb(w_n19438_0[1]),.dout(n19445),.clk(gclk));
	jor g19192(.dina(w_n19445_0[2]),.dinb(w_n743_30[2]),.dout(n19446),.clk(gclk));
	jand g19193(.dina(w_n19445_0[1]),.dinb(w_n743_30[1]),.dout(n19447),.clk(gclk));
	jxor g19194(.dina(w_n18768_0[0]),.dinb(w_n884_29[0]),.dout(n19448),.clk(gclk));
	jor g19195(.dina(n19448),.dinb(w_n19096_20[2]),.dout(n19449),.clk(gclk));
	jxor g19196(.dina(n19449),.dinb(w_n18774_0[0]),.dout(n19450),.clk(gclk));
	jor g19197(.dina(w_n19450_0[2]),.dinb(n19447),.dout(n19451),.clk(gclk));
	jand g19198(.dina(n19451),.dinb(w_n19446_0[1]),.dout(n19452),.clk(gclk));
	jor g19199(.dina(w_n19452_0[2]),.dinb(w_n635_30[2]),.dout(n19453),.clk(gclk));
	jand g19200(.dina(w_n19452_0[1]),.dinb(w_n635_30[1]),.dout(n19454),.clk(gclk));
	jxor g19201(.dina(w_n18776_0[0]),.dinb(w_n743_30[0]),.dout(n19455),.clk(gclk));
	jor g19202(.dina(n19455),.dinb(w_n19096_20[1]),.dout(n19456),.clk(gclk));
	jxor g19203(.dina(n19456),.dinb(w_n19039_0[0]),.dout(n19457),.clk(gclk));
	jnot g19204(.din(w_n19457_0[2]),.dout(n19458),.clk(gclk));
	jor g19205(.dina(n19458),.dinb(n19454),.dout(n19459),.clk(gclk));
	jand g19206(.dina(n19459),.dinb(w_n19453_0[1]),.dout(n19460),.clk(gclk));
	jor g19207(.dina(w_n19460_0[2]),.dinb(w_n515_31[2]),.dout(n19461),.clk(gclk));
	jand g19208(.dina(w_n19460_0[1]),.dinb(w_n515_31[1]),.dout(n19462),.clk(gclk));
	jxor g19209(.dina(w_n18783_0[0]),.dinb(w_n635_30[0]),.dout(n19463),.clk(gclk));
	jor g19210(.dina(n19463),.dinb(w_n19096_20[0]),.dout(n19464),.clk(gclk));
	jxor g19211(.dina(n19464),.dinb(w_n18789_0[0]),.dout(n19465),.clk(gclk));
	jor g19212(.dina(w_n19465_0[2]),.dinb(n19462),.dout(n19466),.clk(gclk));
	jand g19213(.dina(n19466),.dinb(w_n19461_0[1]),.dout(n19467),.clk(gclk));
	jor g19214(.dina(w_n19467_0[2]),.dinb(w_n443_31[2]),.dout(n19468),.clk(gclk));
	jand g19215(.dina(w_n19467_0[1]),.dinb(w_n443_31[1]),.dout(n19469),.clk(gclk));
	jxor g19216(.dina(w_n18791_0[0]),.dinb(w_n515_31[0]),.dout(n19470),.clk(gclk));
	jor g19217(.dina(n19470),.dinb(w_n19096_19[2]),.dout(n19471),.clk(gclk));
	jxor g19218(.dina(n19471),.dinb(w_n19046_0[0]),.dout(n19472),.clk(gclk));
	jnot g19219(.din(w_n19472_0[1]),.dout(n19473),.clk(gclk));
	jor g19220(.dina(w_n19473_0[1]),.dinb(n19469),.dout(n19474),.clk(gclk));
	jand g19221(.dina(n19474),.dinb(w_n19468_0[1]),.dout(n19475),.clk(gclk));
	jor g19222(.dina(w_n19475_0[2]),.dinb(w_n352_32[0]),.dout(n19476),.clk(gclk));
	jand g19223(.dina(w_n19475_0[1]),.dinb(w_n352_31[2]),.dout(n19477),.clk(gclk));
	jxor g19224(.dina(w_n18798_0[0]),.dinb(w_n443_31[0]),.dout(n19478),.clk(gclk));
	jor g19225(.dina(n19478),.dinb(w_n19096_19[1]),.dout(n19479),.clk(gclk));
	jxor g19226(.dina(n19479),.dinb(w_n18803_0[0]),.dout(n19480),.clk(gclk));
	jnot g19227(.din(w_n19480_0[2]),.dout(n19481),.clk(gclk));
	jor g19228(.dina(n19481),.dinb(n19477),.dout(n19482),.clk(gclk));
	jand g19229(.dina(n19482),.dinb(w_n19476_0[1]),.dout(n19483),.clk(gclk));
	jor g19230(.dina(w_n19483_0[2]),.dinb(w_n294_32[1]),.dout(n19484),.clk(gclk));
	jand g19231(.dina(w_n19483_0[1]),.dinb(w_n294_32[0]),.dout(n19485),.clk(gclk));
	jxor g19232(.dina(w_n18806_0[0]),.dinb(w_n352_31[1]),.dout(n19486),.clk(gclk));
	jor g19233(.dina(n19486),.dinb(w_n19096_19[0]),.dout(n19487),.clk(gclk));
	jxor g19234(.dina(n19487),.dinb(w_n18812_0[0]),.dout(n19488),.clk(gclk));
	jor g19235(.dina(w_n19488_0[2]),.dinb(n19485),.dout(n19489),.clk(gclk));
	jand g19236(.dina(n19489),.dinb(w_n19484_0[1]),.dout(n19490),.clk(gclk));
	jor g19237(.dina(w_n19490_0[2]),.dinb(w_n239_32[1]),.dout(n19491),.clk(gclk));
	jand g19238(.dina(w_n19490_0[1]),.dinb(w_n239_32[0]),.dout(n19492),.clk(gclk));
	jxor g19239(.dina(w_n18814_0[0]),.dinb(w_n294_31[2]),.dout(n19493),.clk(gclk));
	jor g19240(.dina(n19493),.dinb(w_n19096_18[2]),.dout(n19494),.clk(gclk));
	jxor g19241(.dina(n19494),.dinb(w_n18820_0[0]),.dout(n19495),.clk(gclk));
	jor g19242(.dina(w_n19495_0[2]),.dinb(n19492),.dout(n19496),.clk(gclk));
	jand g19243(.dina(n19496),.dinb(w_n19491_0[1]),.dout(n19497),.clk(gclk));
	jor g19244(.dina(w_n19497_0[2]),.dinb(w_n221_32[1]),.dout(n19498),.clk(gclk));
	jand g19245(.dina(w_n19497_0[1]),.dinb(w_n221_32[0]),.dout(n19499),.clk(gclk));
	jxor g19246(.dina(w_n18822_0[0]),.dinb(w_n239_31[2]),.dout(n19500),.clk(gclk));
	jor g19247(.dina(n19500),.dinb(w_n19096_18[1]),.dout(n19501),.clk(gclk));
	jxor g19248(.dina(n19501),.dinb(w_n19059_0[0]),.dout(n19502),.clk(gclk));
	jnot g19249(.din(w_n19502_0[2]),.dout(n19503),.clk(gclk));
	jor g19250(.dina(n19503),.dinb(n19499),.dout(n19504),.clk(gclk));
	jand g19251(.dina(n19504),.dinb(w_n19498_0[1]),.dout(n19505),.clk(gclk));
	jor g19252(.dina(w_n19505_0[2]),.dinb(w_n19100_0[2]),.dout(n19506),.clk(gclk));
	jand g19253(.dina(w_asqrt9_7[2]),.dinb(w_n19087_0[0]),.dout(n19507),.clk(gclk));
	jor g19254(.dina(n19507),.dinb(w_n19074_0[0]),.dout(n19508),.clk(gclk));
	jor g19255(.dina(w_n19508_0[1]),.dinb(w_n19506_0[1]),.dout(n19509),.clk(gclk));
	jand g19256(.dina(n19509),.dinb(w_n218_13[2]),.dout(n19510),.clk(gclk));
	jand g19257(.dina(w_n19505_0[1]),.dinb(w_n19100_0[1]),.dout(n19511),.clk(gclk));
	jand g19258(.dina(w_asqrt9_7[1]),.dinb(w_n18182_0[1]),.dout(n19512),.clk(gclk));
	jor g19259(.dina(n19512),.dinb(w_n19086_0[0]),.dout(n19513),.clk(gclk));
	jand g19260(.dina(n19513),.dinb(w_n19068_0[0]),.dout(n19514),.clk(gclk));
	jand g19261(.dina(n19514),.dinb(w_asqrt63_23[1]),.dout(n19515),.clk(gclk));
	jor g19262(.dina(w_n19515_0[1]),.dinb(w_n19511_0[1]),.dout(n19516),.clk(gclk));
	jor g19263(.dina(n19516),.dinb(n19510),.dout(asqrt_fa_9),.clk(gclk));
	jxor g19264(.dina(w_n19497_0[0]),.dinb(w_n221_31[2]),.dout(n19520),.clk(gclk));
	jand g19265(.dina(n19520),.dinb(w_asqrt8_32[1]),.dout(n19521),.clk(gclk));
	jxor g19266(.dina(n19521),.dinb(w_n19502_0[1]),.dout(n19522),.clk(gclk));
	jnot g19267(.din(w_n19522_0[2]),.dout(n19523),.clk(gclk));
	jnot g19268(.din(w_a14_1[1]),.dout(n19524),.clk(gclk));
	jnot g19269(.din(w_a15_0[1]),.dout(n19525),.clk(gclk));
	jand g19270(.dina(w_n19525_0[1]),.dinb(w_n19524_1[1]),.dout(n19526),.clk(gclk));
	jand g19271(.dina(w_n19526_0[2]),.dinb(w_n19101_1[1]),.dout(n19527),.clk(gclk));
	jand g19272(.dina(w_asqrt8_32[0]),.dinb(w_a16_0[1]),.dout(n19528),.clk(gclk));
	jor g19273(.dina(n19528),.dinb(w_n19527_0[1]),.dout(n19529),.clk(gclk));
	jand g19274(.dina(w_n19529_0[2]),.dinb(w_asqrt9_7[0]),.dout(n19530),.clk(gclk));
	jor g19275(.dina(w_n19529_0[1]),.dinb(w_asqrt9_6[2]),.dout(n19531),.clk(gclk));
	jand g19276(.dina(w_asqrt8_31[2]),.dinb(w_n19101_1[0]),.dout(n19532),.clk(gclk));
	jor g19277(.dina(n19532),.dinb(w_n19102_0[0]),.dout(n19533),.clk(gclk));
	jnot g19278(.din(w_n19103_0[1]),.dout(n19534),.clk(gclk));
	jnot g19279(.din(w_n19498_0[0]),.dout(n19535),.clk(gclk));
	jnot g19280(.din(w_n19491_0[0]),.dout(n19536),.clk(gclk));
	jnot g19281(.din(w_n19484_0[0]),.dout(n19537),.clk(gclk));
	jnot g19282(.din(w_n19476_0[0]),.dout(n19538),.clk(gclk));
	jnot g19283(.din(w_n19468_0[0]),.dout(n19539),.clk(gclk));
	jnot g19284(.din(w_n19461_0[0]),.dout(n19540),.clk(gclk));
	jnot g19285(.din(w_n19453_0[0]),.dout(n19541),.clk(gclk));
	jnot g19286(.din(w_n19446_0[0]),.dout(n19542),.clk(gclk));
	jnot g19287(.din(w_n19438_0[0]),.dout(n19543),.clk(gclk));
	jnot g19288(.din(w_n19430_0[0]),.dout(n19544),.clk(gclk));
	jnot g19289(.din(w_n19423_0[0]),.dout(n19545),.clk(gclk));
	jnot g19290(.din(w_n19416_0[0]),.dout(n19546),.clk(gclk));
	jnot g19291(.din(w_n19408_0[0]),.dout(n19547),.clk(gclk));
	jnot g19292(.din(w_n19401_0[0]),.dout(n19548),.clk(gclk));
	jnot g19293(.din(w_n19393_0[0]),.dout(n19549),.clk(gclk));
	jnot g19294(.din(w_n19386_0[0]),.dout(n19550),.clk(gclk));
	jnot g19295(.din(w_n19379_0[0]),.dout(n19551),.clk(gclk));
	jnot g19296(.din(w_n19372_0[0]),.dout(n19552),.clk(gclk));
	jnot g19297(.din(w_n19365_0[0]),.dout(n19553),.clk(gclk));
	jnot g19298(.din(w_n19358_0[0]),.dout(n19554),.clk(gclk));
	jnot g19299(.din(w_n19350_0[0]),.dout(n19555),.clk(gclk));
	jnot g19300(.din(w_n19343_0[0]),.dout(n19556),.clk(gclk));
	jnot g19301(.din(w_n19336_0[0]),.dout(n19557),.clk(gclk));
	jnot g19302(.din(w_n19329_0[0]),.dout(n19558),.clk(gclk));
	jnot g19303(.din(w_n19321_0[0]),.dout(n19559),.clk(gclk));
	jnot g19304(.din(w_n19314_0[0]),.dout(n19560),.clk(gclk));
	jnot g19305(.din(w_n19306_0[0]),.dout(n19561),.clk(gclk));
	jnot g19306(.din(w_n19299_0[0]),.dout(n19562),.clk(gclk));
	jnot g19307(.din(w_n19291_0[0]),.dout(n19563),.clk(gclk));
	jnot g19308(.din(w_n19284_0[0]),.dout(n19564),.clk(gclk));
	jnot g19309(.din(w_n19276_0[0]),.dout(n19565),.clk(gclk));
	jnot g19310(.din(w_n19269_0[0]),.dout(n19566),.clk(gclk));
	jnot g19311(.din(w_n19262_0[0]),.dout(n19567),.clk(gclk));
	jnot g19312(.din(w_n19255_0[0]),.dout(n19568),.clk(gclk));
	jnot g19313(.din(w_n19247_0[0]),.dout(n19569),.clk(gclk));
	jnot g19314(.din(w_n19240_0[0]),.dout(n19570),.clk(gclk));
	jnot g19315(.din(w_n19232_0[0]),.dout(n19571),.clk(gclk));
	jnot g19316(.din(w_n19225_0[0]),.dout(n19572),.clk(gclk));
	jnot g19317(.din(w_n19217_0[0]),.dout(n19573),.clk(gclk));
	jnot g19318(.din(w_n19209_0[0]),.dout(n19574),.clk(gclk));
	jnot g19319(.din(w_n19202_0[0]),.dout(n19575),.clk(gclk));
	jnot g19320(.din(w_n19195_0[0]),.dout(n19576),.clk(gclk));
	jnot g19321(.din(w_n19187_0[0]),.dout(n19577),.clk(gclk));
	jnot g19322(.din(w_n19180_0[0]),.dout(n19578),.clk(gclk));
	jnot g19323(.din(w_n19172_0[0]),.dout(n19579),.clk(gclk));
	jnot g19324(.din(w_n19165_0[0]),.dout(n19580),.clk(gclk));
	jnot g19325(.din(w_n19157_0[0]),.dout(n19581),.clk(gclk));
	jnot g19326(.din(w_n19150_0[0]),.dout(n19582),.clk(gclk));
	jnot g19327(.din(w_n19142_0[0]),.dout(n19583),.clk(gclk));
	jnot g19328(.din(w_n19135_0[0]),.dout(n19584),.clk(gclk));
	jnot g19329(.din(w_n19127_0[0]),.dout(n19585),.clk(gclk));
	jnot g19330(.din(w_n19116_0[0]),.dout(n19586),.clk(gclk));
	jnot g19331(.din(w_n19108_0[0]),.dout(n19587),.clk(gclk));
	jand g19332(.dina(w_asqrt9_6[1]),.dinb(w_a18_0[2]),.dout(n19588),.clk(gclk));
	jor g19333(.dina(n19588),.dinb(w_n19104_0[0]),.dout(n19589),.clk(gclk));
	jor g19334(.dina(n19589),.dinb(w_asqrt10_14[1]),.dout(n19590),.clk(gclk));
	jand g19335(.dina(w_asqrt9_6[0]),.dinb(w_n18185_0[1]),.dout(n19591),.clk(gclk));
	jor g19336(.dina(n19591),.dinb(w_n18186_0[0]),.dout(n19592),.clk(gclk));
	jand g19337(.dina(w_n19119_0[0]),.dinb(n19592),.dout(n19593),.clk(gclk));
	jand g19338(.dina(n19593),.dinb(n19590),.dout(n19594),.clk(gclk));
	jor g19339(.dina(n19594),.dinb(n19587),.dout(n19595),.clk(gclk));
	jor g19340(.dina(n19595),.dinb(w_asqrt11_6[1]),.dout(n19596),.clk(gclk));
	jnot g19341(.din(w_n19124_0[1]),.dout(n19597),.clk(gclk));
	jand g19342(.dina(n19597),.dinb(n19596),.dout(n19598),.clk(gclk));
	jor g19343(.dina(n19598),.dinb(n19586),.dout(n19599),.clk(gclk));
	jor g19344(.dina(n19599),.dinb(w_asqrt12_14[2]),.dout(n19600),.clk(gclk));
	jand g19345(.dina(w_n19131_0[1]),.dinb(n19600),.dout(n19601),.clk(gclk));
	jor g19346(.dina(n19601),.dinb(n19585),.dout(n19602),.clk(gclk));
	jor g19347(.dina(n19602),.dinb(w_asqrt13_7[0]),.dout(n19603),.clk(gclk));
	jnot g19348(.din(w_n19139_0[1]),.dout(n19604),.clk(gclk));
	jand g19349(.dina(n19604),.dinb(n19603),.dout(n19605),.clk(gclk));
	jor g19350(.dina(n19605),.dinb(n19584),.dout(n19606),.clk(gclk));
	jor g19351(.dina(n19606),.dinb(w_asqrt14_15[0]),.dout(n19607),.clk(gclk));
	jand g19352(.dina(w_n19146_0[1]),.dinb(n19607),.dout(n19608),.clk(gclk));
	jor g19353(.dina(n19608),.dinb(n19583),.dout(n19609),.clk(gclk));
	jor g19354(.dina(n19609),.dinb(w_asqrt15_7[2]),.dout(n19610),.clk(gclk));
	jnot g19355(.din(w_n19154_0[1]),.dout(n19611),.clk(gclk));
	jand g19356(.dina(n19611),.dinb(n19610),.dout(n19612),.clk(gclk));
	jor g19357(.dina(n19612),.dinb(n19582),.dout(n19613),.clk(gclk));
	jor g19358(.dina(n19613),.dinb(w_asqrt16_15[0]),.dout(n19614),.clk(gclk));
	jand g19359(.dina(w_n19161_0[1]),.dinb(n19614),.dout(n19615),.clk(gclk));
	jor g19360(.dina(n19615),.dinb(n19581),.dout(n19616),.clk(gclk));
	jor g19361(.dina(n19616),.dinb(w_asqrt17_8[0]),.dout(n19617),.clk(gclk));
	jnot g19362(.din(w_n19169_0[1]),.dout(n19618),.clk(gclk));
	jand g19363(.dina(n19618),.dinb(n19617),.dout(n19619),.clk(gclk));
	jor g19364(.dina(n19619),.dinb(n19580),.dout(n19620),.clk(gclk));
	jor g19365(.dina(n19620),.dinb(w_asqrt18_15[1]),.dout(n19621),.clk(gclk));
	jand g19366(.dina(w_n19176_0[1]),.dinb(n19621),.dout(n19622),.clk(gclk));
	jor g19367(.dina(n19622),.dinb(n19579),.dout(n19623),.clk(gclk));
	jor g19368(.dina(n19623),.dinb(w_asqrt19_8[1]),.dout(n19624),.clk(gclk));
	jnot g19369(.din(w_n19184_0[1]),.dout(n19625),.clk(gclk));
	jand g19370(.dina(n19625),.dinb(n19624),.dout(n19626),.clk(gclk));
	jor g19371(.dina(n19626),.dinb(n19578),.dout(n19627),.clk(gclk));
	jor g19372(.dina(n19627),.dinb(w_asqrt20_15[1]),.dout(n19628),.clk(gclk));
	jand g19373(.dina(w_n19191_0[1]),.dinb(n19628),.dout(n19629),.clk(gclk));
	jor g19374(.dina(n19629),.dinb(n19577),.dout(n19630),.clk(gclk));
	jor g19375(.dina(n19630),.dinb(w_asqrt21_9[0]),.dout(n19631),.clk(gclk));
	jnot g19376(.din(w_n19199_0[1]),.dout(n19632),.clk(gclk));
	jand g19377(.dina(n19632),.dinb(n19631),.dout(n19633),.clk(gclk));
	jor g19378(.dina(n19633),.dinb(n19576),.dout(n19634),.clk(gclk));
	jor g19379(.dina(n19634),.dinb(w_asqrt22_15[2]),.dout(n19635),.clk(gclk));
	jnot g19380(.din(w_n19206_0[1]),.dout(n19636),.clk(gclk));
	jand g19381(.dina(n19636),.dinb(n19635),.dout(n19637),.clk(gclk));
	jor g19382(.dina(n19637),.dinb(n19575),.dout(n19638),.clk(gclk));
	jor g19383(.dina(n19638),.dinb(w_asqrt23_9[2]),.dout(n19639),.clk(gclk));
	jand g19384(.dina(w_n19213_0[1]),.dinb(n19639),.dout(n19640),.clk(gclk));
	jor g19385(.dina(n19640),.dinb(n19574),.dout(n19641),.clk(gclk));
	jor g19386(.dina(n19641),.dinb(w_asqrt24_15[2]),.dout(n19642),.clk(gclk));
	jand g19387(.dina(w_n19221_0[1]),.dinb(n19642),.dout(n19643),.clk(gclk));
	jor g19388(.dina(n19643),.dinb(n19573),.dout(n19644),.clk(gclk));
	jor g19389(.dina(n19644),.dinb(w_asqrt25_9[2]),.dout(n19645),.clk(gclk));
	jnot g19390(.din(w_n19229_0[1]),.dout(n19646),.clk(gclk));
	jand g19391(.dina(n19646),.dinb(n19645),.dout(n19647),.clk(gclk));
	jor g19392(.dina(n19647),.dinb(n19572),.dout(n19648),.clk(gclk));
	jor g19393(.dina(n19648),.dinb(w_asqrt26_15[2]),.dout(n19649),.clk(gclk));
	jand g19394(.dina(w_n19236_0[1]),.dinb(n19649),.dout(n19650),.clk(gclk));
	jor g19395(.dina(n19650),.dinb(n19571),.dout(n19651),.clk(gclk));
	jor g19396(.dina(n19651),.dinb(w_asqrt27_10[1]),.dout(n19652),.clk(gclk));
	jnot g19397(.din(w_n19244_0[1]),.dout(n19653),.clk(gclk));
	jand g19398(.dina(n19653),.dinb(n19652),.dout(n19654),.clk(gclk));
	jor g19399(.dina(n19654),.dinb(n19570),.dout(n19655),.clk(gclk));
	jor g19400(.dina(n19655),.dinb(w_asqrt28_16[0]),.dout(n19656),.clk(gclk));
	jand g19401(.dina(w_n19251_0[1]),.dinb(n19656),.dout(n19657),.clk(gclk));
	jor g19402(.dina(n19657),.dinb(n19569),.dout(n19658),.clk(gclk));
	jor g19403(.dina(n19658),.dinb(w_asqrt29_10[2]),.dout(n19659),.clk(gclk));
	jnot g19404(.din(w_n19259_0[1]),.dout(n19660),.clk(gclk));
	jand g19405(.dina(n19660),.dinb(n19659),.dout(n19661),.clk(gclk));
	jor g19406(.dina(n19661),.dinb(n19568),.dout(n19662),.clk(gclk));
	jor g19407(.dina(n19662),.dinb(w_asqrt30_16[1]),.dout(n19663),.clk(gclk));
	jnot g19408(.din(w_n19266_0[1]),.dout(n19664),.clk(gclk));
	jand g19409(.dina(n19664),.dinb(n19663),.dout(n19665),.clk(gclk));
	jor g19410(.dina(n19665),.dinb(n19567),.dout(n19666),.clk(gclk));
	jor g19411(.dina(n19666),.dinb(w_asqrt31_11[1]),.dout(n19667),.clk(gclk));
	jnot g19412(.din(w_n19273_0[1]),.dout(n19668),.clk(gclk));
	jand g19413(.dina(n19668),.dinb(n19667),.dout(n19669),.clk(gclk));
	jor g19414(.dina(n19669),.dinb(n19566),.dout(n19670),.clk(gclk));
	jor g19415(.dina(n19670),.dinb(w_asqrt32_16[1]),.dout(n19671),.clk(gclk));
	jand g19416(.dina(w_n19280_0[1]),.dinb(n19671),.dout(n19672),.clk(gclk));
	jor g19417(.dina(n19672),.dinb(n19565),.dout(n19673),.clk(gclk));
	jor g19418(.dina(n19673),.dinb(w_asqrt33_12[0]),.dout(n19674),.clk(gclk));
	jnot g19419(.din(w_n19288_0[1]),.dout(n19675),.clk(gclk));
	jand g19420(.dina(n19675),.dinb(n19674),.dout(n19676),.clk(gclk));
	jor g19421(.dina(n19676),.dinb(n19564),.dout(n19677),.clk(gclk));
	jor g19422(.dina(n19677),.dinb(w_asqrt34_16[2]),.dout(n19678),.clk(gclk));
	jand g19423(.dina(w_n19295_0[1]),.dinb(n19678),.dout(n19679),.clk(gclk));
	jor g19424(.dina(n19679),.dinb(n19563),.dout(n19680),.clk(gclk));
	jor g19425(.dina(n19680),.dinb(w_asqrt35_12[2]),.dout(n19681),.clk(gclk));
	jnot g19426(.din(w_n19303_0[1]),.dout(n19682),.clk(gclk));
	jand g19427(.dina(n19682),.dinb(n19681),.dout(n19683),.clk(gclk));
	jor g19428(.dina(n19683),.dinb(n19562),.dout(n19684),.clk(gclk));
	jor g19429(.dina(n19684),.dinb(w_asqrt36_16[2]),.dout(n19685),.clk(gclk));
	jand g19430(.dina(w_n19310_0[1]),.dinb(n19685),.dout(n19686),.clk(gclk));
	jor g19431(.dina(n19686),.dinb(n19561),.dout(n19687),.clk(gclk));
	jor g19432(.dina(n19687),.dinb(w_asqrt37_13[0]),.dout(n19688),.clk(gclk));
	jnot g19433(.din(w_n19318_0[1]),.dout(n19689),.clk(gclk));
	jand g19434(.dina(n19689),.dinb(n19688),.dout(n19690),.clk(gclk));
	jor g19435(.dina(n19690),.dinb(n19560),.dout(n19691),.clk(gclk));
	jor g19436(.dina(n19691),.dinb(w_asqrt38_17[0]),.dout(n19692),.clk(gclk));
	jand g19437(.dina(w_n19325_0[1]),.dinb(n19692),.dout(n19693),.clk(gclk));
	jor g19438(.dina(n19693),.dinb(n19559),.dout(n19694),.clk(gclk));
	jor g19439(.dina(n19694),.dinb(w_asqrt39_13[2]),.dout(n19695),.clk(gclk));
	jnot g19440(.din(w_n19333_0[1]),.dout(n19696),.clk(gclk));
	jand g19441(.dina(n19696),.dinb(n19695),.dout(n19697),.clk(gclk));
	jor g19442(.dina(n19697),.dinb(n19558),.dout(n19698),.clk(gclk));
	jor g19443(.dina(n19698),.dinb(w_asqrt40_17[0]),.dout(n19699),.clk(gclk));
	jnot g19444(.din(w_n19340_0[1]),.dout(n19700),.clk(gclk));
	jand g19445(.dina(n19700),.dinb(n19699),.dout(n19701),.clk(gclk));
	jor g19446(.dina(n19701),.dinb(n19557),.dout(n19702),.clk(gclk));
	jor g19447(.dina(n19702),.dinb(w_asqrt41_14[0]),.dout(n19703),.clk(gclk));
	jnot g19448(.din(w_n19347_0[1]),.dout(n19704),.clk(gclk));
	jand g19449(.dina(n19704),.dinb(n19703),.dout(n19705),.clk(gclk));
	jor g19450(.dina(n19705),.dinb(n19556),.dout(n19706),.clk(gclk));
	jor g19451(.dina(n19706),.dinb(w_asqrt42_17[1]),.dout(n19707),.clk(gclk));
	jand g19452(.dina(w_n19354_0[1]),.dinb(n19707),.dout(n19708),.clk(gclk));
	jor g19453(.dina(n19708),.dinb(n19555),.dout(n19709),.clk(gclk));
	jor g19454(.dina(n19709),.dinb(w_asqrt43_14[1]),.dout(n19710),.clk(gclk));
	jnot g19455(.din(w_n19362_0[1]),.dout(n19711),.clk(gclk));
	jand g19456(.dina(n19711),.dinb(n19710),.dout(n19712),.clk(gclk));
	jor g19457(.dina(n19712),.dinb(n19554),.dout(n19713),.clk(gclk));
	jor g19458(.dina(n19713),.dinb(w_asqrt44_17[1]),.dout(n19714),.clk(gclk));
	jnot g19459(.din(w_n19369_0[1]),.dout(n19715),.clk(gclk));
	jand g19460(.dina(n19715),.dinb(n19714),.dout(n19716),.clk(gclk));
	jor g19461(.dina(n19716),.dinb(n19553),.dout(n19717),.clk(gclk));
	jor g19462(.dina(n19717),.dinb(w_asqrt45_15[0]),.dout(n19718),.clk(gclk));
	jnot g19463(.din(w_n19376_0[1]),.dout(n19719),.clk(gclk));
	jand g19464(.dina(n19719),.dinb(n19718),.dout(n19720),.clk(gclk));
	jor g19465(.dina(n19720),.dinb(n19552),.dout(n19721),.clk(gclk));
	jor g19466(.dina(n19721),.dinb(w_asqrt46_17[1]),.dout(n19722),.clk(gclk));
	jnot g19467(.din(w_n19383_0[1]),.dout(n19723),.clk(gclk));
	jand g19468(.dina(n19723),.dinb(n19722),.dout(n19724),.clk(gclk));
	jor g19469(.dina(n19724),.dinb(n19551),.dout(n19725),.clk(gclk));
	jor g19470(.dina(n19725),.dinb(w_asqrt47_15[2]),.dout(n19726),.clk(gclk));
	jnot g19471(.din(w_n19390_0[1]),.dout(n19727),.clk(gclk));
	jand g19472(.dina(n19727),.dinb(n19726),.dout(n19728),.clk(gclk));
	jor g19473(.dina(n19728),.dinb(n19550),.dout(n19729),.clk(gclk));
	jor g19474(.dina(n19729),.dinb(w_asqrt48_17[2]),.dout(n19730),.clk(gclk));
	jand g19475(.dina(w_n19397_0[1]),.dinb(n19730),.dout(n19731),.clk(gclk));
	jor g19476(.dina(n19731),.dinb(n19549),.dout(n19732),.clk(gclk));
	jor g19477(.dina(n19732),.dinb(w_asqrt49_16[0]),.dout(n19733),.clk(gclk));
	jnot g19478(.din(w_n19405_0[1]),.dout(n19734),.clk(gclk));
	jand g19479(.dina(n19734),.dinb(n19733),.dout(n19735),.clk(gclk));
	jor g19480(.dina(n19735),.dinb(n19548),.dout(n19736),.clk(gclk));
	jor g19481(.dina(n19736),.dinb(w_asqrt50_18[0]),.dout(n19737),.clk(gclk));
	jand g19482(.dina(w_n19412_0[1]),.dinb(n19737),.dout(n19738),.clk(gclk));
	jor g19483(.dina(n19738),.dinb(n19547),.dout(n19739),.clk(gclk));
	jor g19484(.dina(n19739),.dinb(w_asqrt51_16[1]),.dout(n19740),.clk(gclk));
	jnot g19485(.din(w_n19420_0[1]),.dout(n19741),.clk(gclk));
	jand g19486(.dina(n19741),.dinb(n19740),.dout(n19742),.clk(gclk));
	jor g19487(.dina(n19742),.dinb(n19546),.dout(n19743),.clk(gclk));
	jor g19488(.dina(n19743),.dinb(w_asqrt52_18[0]),.dout(n19744),.clk(gclk));
	jnot g19489(.din(w_n19427_0[1]),.dout(n19745),.clk(gclk));
	jand g19490(.dina(n19745),.dinb(n19744),.dout(n19746),.clk(gclk));
	jor g19491(.dina(n19746),.dinb(n19545),.dout(n19747),.clk(gclk));
	jor g19492(.dina(n19747),.dinb(w_asqrt53_17[0]),.dout(n19748),.clk(gclk));
	jand g19493(.dina(w_n19434_0[1]),.dinb(n19748),.dout(n19749),.clk(gclk));
	jor g19494(.dina(n19749),.dinb(n19544),.dout(n19750),.clk(gclk));
	jor g19495(.dina(n19750),.dinb(w_asqrt54_18[0]),.dout(n19751),.clk(gclk));
	jand g19496(.dina(n19751),.dinb(w_n19441_0[1]),.dout(n19752),.clk(gclk));
	jor g19497(.dina(n19752),.dinb(n19543),.dout(n19753),.clk(gclk));
	jor g19498(.dina(n19753),.dinb(w_asqrt55_17[1]),.dout(n19754),.clk(gclk));
	jnot g19499(.din(w_n19450_0[1]),.dout(n19755),.clk(gclk));
	jand g19500(.dina(n19755),.dinb(n19754),.dout(n19756),.clk(gclk));
	jor g19501(.dina(n19756),.dinb(n19542),.dout(n19757),.clk(gclk));
	jor g19502(.dina(n19757),.dinb(w_asqrt56_18[1]),.dout(n19758),.clk(gclk));
	jand g19503(.dina(w_n19457_0[1]),.dinb(n19758),.dout(n19759),.clk(gclk));
	jor g19504(.dina(n19759),.dinb(n19541),.dout(n19760),.clk(gclk));
	jor g19505(.dina(n19760),.dinb(w_asqrt57_18[0]),.dout(n19761),.clk(gclk));
	jnot g19506(.din(w_n19465_0[1]),.dout(n19762),.clk(gclk));
	jand g19507(.dina(n19762),.dinb(n19761),.dout(n19763),.clk(gclk));
	jor g19508(.dina(n19763),.dinb(n19540),.dout(n19764),.clk(gclk));
	jor g19509(.dina(n19764),.dinb(w_asqrt58_18[2]),.dout(n19765),.clk(gclk));
	jand g19510(.dina(w_n19472_0[0]),.dinb(n19765),.dout(n19766),.clk(gclk));
	jor g19511(.dina(n19766),.dinb(n19539),.dout(n19767),.clk(gclk));
	jor g19512(.dina(n19767),.dinb(w_asqrt59_18[1]),.dout(n19768),.clk(gclk));
	jand g19513(.dina(w_n19480_0[1]),.dinb(n19768),.dout(n19769),.clk(gclk));
	jor g19514(.dina(n19769),.dinb(n19538),.dout(n19770),.clk(gclk));
	jor g19515(.dina(n19770),.dinb(w_asqrt60_18[2]),.dout(n19771),.clk(gclk));
	jnot g19516(.din(w_n19488_0[1]),.dout(n19772),.clk(gclk));
	jand g19517(.dina(n19772),.dinb(n19771),.dout(n19773),.clk(gclk));
	jor g19518(.dina(n19773),.dinb(n19537),.dout(n19774),.clk(gclk));
	jor g19519(.dina(n19774),.dinb(w_asqrt61_18[2]),.dout(n19775),.clk(gclk));
	jnot g19520(.din(w_n19495_0[1]),.dout(n19776),.clk(gclk));
	jand g19521(.dina(n19776),.dinb(n19775),.dout(n19777),.clk(gclk));
	jor g19522(.dina(n19777),.dinb(n19536),.dout(n19778),.clk(gclk));
	jor g19523(.dina(n19778),.dinb(w_asqrt62_18[2]),.dout(n19779),.clk(gclk));
	jand g19524(.dina(w_n19502_0[0]),.dinb(n19779),.dout(n19780),.clk(gclk));
	jor g19525(.dina(n19780),.dinb(n19535),.dout(n19781),.clk(gclk));
	jand g19526(.dina(w_n19781_0[1]),.dinb(w_n19099_0[1]),.dout(n19782),.clk(gclk));
	jnot g19527(.din(w_n19508_0[0]),.dout(n19783),.clk(gclk));
	jand g19528(.dina(n19783),.dinb(w_n19782_0[1]),.dout(n19784),.clk(gclk));
	jor g19529(.dina(n19784),.dinb(w_asqrt63_23[0]),.dout(n19785),.clk(gclk));
	jor g19530(.dina(w_n19781_0[0]),.dinb(w_n19099_0[0]),.dout(n19786),.clk(gclk));
	jnot g19531(.din(w_n19515_0[0]),.dout(n19787),.clk(gclk));
	jand g19532(.dina(n19787),.dinb(w_n19786_0[1]),.dout(n19788),.clk(gclk));
	jand g19533(.dina(w_n19788_0[1]),.dinb(w_n19785_0[1]),.dout(n19791),.clk(gclk));
	jor g19534(.dina(w_n19791_10[2]),.dinb(n19534),.dout(n19792),.clk(gclk));
	jand g19535(.dina(n19792),.dinb(n19533),.dout(n19793),.clk(gclk));
	jand g19536(.dina(n19793),.dinb(n19531),.dout(n19794),.clk(gclk));
	jor g19537(.dina(n19794),.dinb(w_n19530_0[1]),.dout(n19795),.clk(gclk));
	jand g19538(.dina(w_n19795_0[2]),.dinb(w_asqrt10_14[0]),.dout(n19796),.clk(gclk));
	jor g19539(.dina(w_n19795_0[1]),.dinb(w_asqrt10_13[2]),.dout(n19797),.clk(gclk));
	jand g19540(.dina(w_asqrt8_31[1]),.dinb(w_n19103_0[0]),.dout(n19798),.clk(gclk));
	jand g19541(.dina(w_n19788_0[0]),.dinb(w_asqrt9_5[2]),.dout(n19799),.clk(gclk));
	jand g19542(.dina(n19799),.dinb(w_n19785_0[0]),.dout(n19800),.clk(gclk));
	jor g19543(.dina(n19800),.dinb(w_n19798_0[1]),.dout(n19801),.clk(gclk));
	jxor g19544(.dina(n19801),.dinb(w_a18_0[1]),.dout(n19802),.clk(gclk));
	jnot g19545(.din(w_n19802_0[1]),.dout(n19803),.clk(gclk));
	jand g19546(.dina(w_n19803_0[1]),.dinb(n19797),.dout(n19804),.clk(gclk));
	jor g19547(.dina(n19804),.dinb(w_n19796_0[1]),.dout(n19805),.clk(gclk));
	jand g19548(.dina(w_n19805_0[2]),.dinb(w_asqrt11_6[0]),.dout(n19806),.clk(gclk));
	jor g19549(.dina(w_n19805_0[1]),.dinb(w_asqrt11_5[2]),.dout(n19807),.clk(gclk));
	jxor g19550(.dina(w_n19107_0[0]),.dinb(w_n18442_10[1]),.dout(n19808),.clk(gclk));
	jand g19551(.dina(n19808),.dinb(w_asqrt8_31[0]),.dout(n19809),.clk(gclk));
	jxor g19552(.dina(n19809),.dinb(w_n19113_0[0]),.dout(n19810),.clk(gclk));
	jnot g19553(.din(w_n19810_0[1]),.dout(n19811),.clk(gclk));
	jand g19554(.dina(w_n19811_0[1]),.dinb(n19807),.dout(n19812),.clk(gclk));
	jor g19555(.dina(n19812),.dinb(w_n19806_0[1]),.dout(n19813),.clk(gclk));
	jand g19556(.dina(w_n19813_0[2]),.dinb(w_asqrt12_14[1]),.dout(n19814),.clk(gclk));
	jor g19557(.dina(w_n19813_0[1]),.dinb(w_asqrt12_14[0]),.dout(n19815),.clk(gclk));
	jxor g19558(.dina(w_n19115_0[0]),.dinb(w_n17769_19[0]),.dout(n19816),.clk(gclk));
	jand g19559(.dina(n19816),.dinb(w_asqrt8_30[2]),.dout(n19817),.clk(gclk));
	jxor g19560(.dina(n19817),.dinb(w_n19124_0[0]),.dout(n19818),.clk(gclk));
	jnot g19561(.din(w_n19818_0[1]),.dout(n19819),.clk(gclk));
	jand g19562(.dina(w_n19819_0[1]),.dinb(n19815),.dout(n19820),.clk(gclk));
	jor g19563(.dina(n19820),.dinb(w_n19814_0[1]),.dout(n19821),.clk(gclk));
	jand g19564(.dina(w_n19821_0[2]),.dinb(w_asqrt13_6[2]),.dout(n19822),.clk(gclk));
	jor g19565(.dina(w_n19821_0[1]),.dinb(w_asqrt13_6[1]),.dout(n19823),.clk(gclk));
	jxor g19566(.dina(w_n19126_0[0]),.dinb(w_n17134_11[1]),.dout(n19824),.clk(gclk));
	jand g19567(.dina(n19824),.dinb(w_asqrt8_30[1]),.dout(n19825),.clk(gclk));
	jxor g19568(.dina(n19825),.dinb(w_n19131_0[0]),.dout(n19826),.clk(gclk));
	jand g19569(.dina(w_n19826_0[1]),.dinb(n19823),.dout(n19827),.clk(gclk));
	jor g19570(.dina(n19827),.dinb(w_n19822_0[1]),.dout(n19828),.clk(gclk));
	jand g19571(.dina(w_n19828_0[2]),.dinb(w_asqrt14_14[2]),.dout(n19829),.clk(gclk));
	jor g19572(.dina(w_n19828_0[1]),.dinb(w_asqrt14_14[1]),.dout(n19830),.clk(gclk));
	jxor g19573(.dina(w_n19134_0[0]),.dinb(w_n16489_19[1]),.dout(n19831),.clk(gclk));
	jand g19574(.dina(n19831),.dinb(w_asqrt8_30[0]),.dout(n19832),.clk(gclk));
	jxor g19575(.dina(n19832),.dinb(w_n19139_0[0]),.dout(n19833),.clk(gclk));
	jnot g19576(.din(w_n19833_0[1]),.dout(n19834),.clk(gclk));
	jand g19577(.dina(w_n19834_0[1]),.dinb(n19830),.dout(n19835),.clk(gclk));
	jor g19578(.dina(n19835),.dinb(w_n19829_0[1]),.dout(n19836),.clk(gclk));
	jand g19579(.dina(w_n19836_0[2]),.dinb(w_asqrt15_7[1]),.dout(n19837),.clk(gclk));
	jor g19580(.dina(w_n19836_0[1]),.dinb(w_asqrt15_7[0]),.dout(n19838),.clk(gclk));
	jxor g19581(.dina(w_n19141_0[0]),.dinb(w_n15878_12[1]),.dout(n19839),.clk(gclk));
	jand g19582(.dina(n19839),.dinb(w_asqrt8_29[2]),.dout(n19840),.clk(gclk));
	jxor g19583(.dina(n19840),.dinb(w_n19146_0[0]),.dout(n19841),.clk(gclk));
	jand g19584(.dina(w_n19841_0[1]),.dinb(n19838),.dout(n19842),.clk(gclk));
	jor g19585(.dina(n19842),.dinb(w_n19837_0[1]),.dout(n19843),.clk(gclk));
	jand g19586(.dina(w_n19843_0[2]),.dinb(w_asqrt16_14[2]),.dout(n19844),.clk(gclk));
	jor g19587(.dina(w_n19843_0[1]),.dinb(w_asqrt16_14[1]),.dout(n19845),.clk(gclk));
	jxor g19588(.dina(w_n19149_0[0]),.dinb(w_n15260_20[0]),.dout(n19846),.clk(gclk));
	jand g19589(.dina(n19846),.dinb(w_asqrt8_29[1]),.dout(n19847),.clk(gclk));
	jxor g19590(.dina(n19847),.dinb(w_n19154_0[0]),.dout(n19848),.clk(gclk));
	jnot g19591(.din(w_n19848_0[1]),.dout(n19849),.clk(gclk));
	jand g19592(.dina(w_n19849_0[1]),.dinb(n19845),.dout(n19850),.clk(gclk));
	jor g19593(.dina(n19850),.dinb(w_n19844_0[1]),.dout(n19851),.clk(gclk));
	jand g19594(.dina(w_n19851_0[2]),.dinb(w_asqrt17_7[2]),.dout(n19852),.clk(gclk));
	jor g19595(.dina(w_n19851_0[1]),.dinb(w_asqrt17_7[1]),.dout(n19853),.clk(gclk));
	jxor g19596(.dina(w_n19156_0[0]),.dinb(w_n14674_13[0]),.dout(n19854),.clk(gclk));
	jand g19597(.dina(n19854),.dinb(w_asqrt8_29[0]),.dout(n19855),.clk(gclk));
	jxor g19598(.dina(n19855),.dinb(w_n19161_0[0]),.dout(n19856),.clk(gclk));
	jand g19599(.dina(w_n19856_0[1]),.dinb(n19853),.dout(n19857),.clk(gclk));
	jor g19600(.dina(n19857),.dinb(w_n19852_0[1]),.dout(n19858),.clk(gclk));
	jand g19601(.dina(w_n19858_0[2]),.dinb(w_asqrt18_15[0]),.dout(n19859),.clk(gclk));
	jor g19602(.dina(w_n19858_0[1]),.dinb(w_asqrt18_14[2]),.dout(n19860),.clk(gclk));
	jxor g19603(.dina(w_n19164_0[0]),.dinb(w_n14078_20[1]),.dout(n19861),.clk(gclk));
	jand g19604(.dina(n19861),.dinb(w_asqrt8_28[2]),.dout(n19862),.clk(gclk));
	jxor g19605(.dina(n19862),.dinb(w_n19169_0[0]),.dout(n19863),.clk(gclk));
	jnot g19606(.din(w_n19863_0[1]),.dout(n19864),.clk(gclk));
	jand g19607(.dina(w_n19864_0[1]),.dinb(n19860),.dout(n19865),.clk(gclk));
	jor g19608(.dina(n19865),.dinb(w_n19859_0[1]),.dout(n19866),.clk(gclk));
	jand g19609(.dina(w_n19866_0[2]),.dinb(w_asqrt19_8[0]),.dout(n19867),.clk(gclk));
	jor g19610(.dina(w_n19866_0[1]),.dinb(w_asqrt19_7[2]),.dout(n19868),.clk(gclk));
	jxor g19611(.dina(w_n19171_0[0]),.dinb(w_n13515_14[0]),.dout(n19869),.clk(gclk));
	jand g19612(.dina(n19869),.dinb(w_asqrt8_28[1]),.dout(n19870),.clk(gclk));
	jxor g19613(.dina(n19870),.dinb(w_n19176_0[0]),.dout(n19871),.clk(gclk));
	jand g19614(.dina(w_n19871_0[1]),.dinb(n19868),.dout(n19872),.clk(gclk));
	jor g19615(.dina(n19872),.dinb(w_n19867_0[1]),.dout(n19873),.clk(gclk));
	jand g19616(.dina(w_n19873_0[2]),.dinb(w_asqrt20_15[0]),.dout(n19874),.clk(gclk));
	jor g19617(.dina(w_n19873_0[1]),.dinb(w_asqrt20_14[2]),.dout(n19875),.clk(gclk));
	jxor g19618(.dina(w_n19179_0[0]),.dinb(w_n12947_21[0]),.dout(n19876),.clk(gclk));
	jand g19619(.dina(n19876),.dinb(w_asqrt8_28[0]),.dout(n19877),.clk(gclk));
	jxor g19620(.dina(n19877),.dinb(w_n19184_0[0]),.dout(n19878),.clk(gclk));
	jnot g19621(.din(w_n19878_0[1]),.dout(n19879),.clk(gclk));
	jand g19622(.dina(w_n19879_0[1]),.dinb(n19875),.dout(n19880),.clk(gclk));
	jor g19623(.dina(n19880),.dinb(w_n19874_0[1]),.dout(n19881),.clk(gclk));
	jand g19624(.dina(w_n19881_0[2]),.dinb(w_asqrt21_8[2]),.dout(n19882),.clk(gclk));
	jor g19625(.dina(w_n19881_0[1]),.dinb(w_asqrt21_8[1]),.dout(n19883),.clk(gclk));
	jxor g19626(.dina(w_n19186_0[0]),.dinb(w_n12410_14[2]),.dout(n19884),.clk(gclk));
	jand g19627(.dina(n19884),.dinb(w_asqrt8_27[2]),.dout(n19885),.clk(gclk));
	jxor g19628(.dina(n19885),.dinb(w_n19191_0[0]),.dout(n19886),.clk(gclk));
	jand g19629(.dina(w_n19886_0[1]),.dinb(n19883),.dout(n19887),.clk(gclk));
	jor g19630(.dina(n19887),.dinb(w_n19882_0[1]),.dout(n19888),.clk(gclk));
	jand g19631(.dina(w_n19888_0[2]),.dinb(w_asqrt22_15[1]),.dout(n19889),.clk(gclk));
	jor g19632(.dina(w_n19888_0[1]),.dinb(w_asqrt22_15[0]),.dout(n19890),.clk(gclk));
	jxor g19633(.dina(w_n19194_0[0]),.dinb(w_n11858_21[1]),.dout(n19891),.clk(gclk));
	jand g19634(.dina(n19891),.dinb(w_asqrt8_27[1]),.dout(n19892),.clk(gclk));
	jxor g19635(.dina(n19892),.dinb(w_n19199_0[0]),.dout(n19893),.clk(gclk));
	jnot g19636(.din(w_n19893_0[1]),.dout(n19894),.clk(gclk));
	jand g19637(.dina(w_n19894_0[1]),.dinb(n19890),.dout(n19895),.clk(gclk));
	jor g19638(.dina(n19895),.dinb(w_n19889_0[1]),.dout(n19896),.clk(gclk));
	jand g19639(.dina(w_n19896_0[2]),.dinb(w_asqrt23_9[1]),.dout(n19897),.clk(gclk));
	jor g19640(.dina(w_n19896_0[1]),.dinb(w_asqrt23_9[0]),.dout(n19898),.clk(gclk));
	jxor g19641(.dina(w_n19201_0[0]),.dinb(w_n11347_15[1]),.dout(n19899),.clk(gclk));
	jand g19642(.dina(n19899),.dinb(w_asqrt8_27[0]),.dout(n19900),.clk(gclk));
	jxor g19643(.dina(n19900),.dinb(w_n19206_0[0]),.dout(n19901),.clk(gclk));
	jnot g19644(.din(w_n19901_0[1]),.dout(n19902),.clk(gclk));
	jand g19645(.dina(w_n19902_0[1]),.dinb(n19898),.dout(n19903),.clk(gclk));
	jor g19646(.dina(n19903),.dinb(w_n19897_0[1]),.dout(n19904),.clk(gclk));
	jand g19647(.dina(w_n19904_0[2]),.dinb(w_asqrt24_15[1]),.dout(n19905),.clk(gclk));
	jor g19648(.dina(w_n19904_0[1]),.dinb(w_asqrt24_15[0]),.dout(n19906),.clk(gclk));
	jxor g19649(.dina(w_n19208_0[0]),.dinb(w_n10824_22[0]),.dout(n19907),.clk(gclk));
	jand g19650(.dina(n19907),.dinb(w_asqrt8_26[2]),.dout(n19908),.clk(gclk));
	jxor g19651(.dina(n19908),.dinb(w_n19213_0[0]),.dout(n19909),.clk(gclk));
	jand g19652(.dina(w_n19909_0[1]),.dinb(n19906),.dout(n19910),.clk(gclk));
	jor g19653(.dina(n19910),.dinb(w_n19905_0[1]),.dout(n19911),.clk(gclk));
	jand g19654(.dina(w_n19911_0[2]),.dinb(w_asqrt25_9[1]),.dout(n19912),.clk(gclk));
	jor g19655(.dina(w_n19911_0[1]),.dinb(w_asqrt25_9[0]),.dout(n19913),.clk(gclk));
	jxor g19656(.dina(w_n19216_0[0]),.dinb(w_n10328_16[1]),.dout(n19914),.clk(gclk));
	jand g19657(.dina(n19914),.dinb(w_asqrt8_26[1]),.dout(n19915),.clk(gclk));
	jxor g19658(.dina(n19915),.dinb(w_n19221_0[0]),.dout(n19916),.clk(gclk));
	jand g19659(.dina(w_n19916_0[1]),.dinb(n19913),.dout(n19917),.clk(gclk));
	jor g19660(.dina(n19917),.dinb(w_n19912_0[1]),.dout(n19918),.clk(gclk));
	jand g19661(.dina(w_n19918_0[2]),.dinb(w_asqrt26_15[1]),.dout(n19919),.clk(gclk));
	jor g19662(.dina(w_n19918_0[1]),.dinb(w_asqrt26_15[0]),.dout(n19920),.clk(gclk));
	jxor g19663(.dina(w_n19224_0[0]),.dinb(w_n9832_22[2]),.dout(n19921),.clk(gclk));
	jand g19664(.dina(n19921),.dinb(w_asqrt8_26[0]),.dout(n19922),.clk(gclk));
	jxor g19665(.dina(n19922),.dinb(w_n19229_0[0]),.dout(n19923),.clk(gclk));
	jnot g19666(.din(w_n19923_0[1]),.dout(n19924),.clk(gclk));
	jand g19667(.dina(w_n19924_0[1]),.dinb(n19920),.dout(n19925),.clk(gclk));
	jor g19668(.dina(n19925),.dinb(w_n19919_0[1]),.dout(n19926),.clk(gclk));
	jand g19669(.dina(w_n19926_0[2]),.dinb(w_asqrt27_10[0]),.dout(n19927),.clk(gclk));
	jor g19670(.dina(w_n19926_0[1]),.dinb(w_asqrt27_9[2]),.dout(n19928),.clk(gclk));
	jxor g19671(.dina(w_n19231_0[0]),.dinb(w_n9369_17[1]),.dout(n19929),.clk(gclk));
	jand g19672(.dina(n19929),.dinb(w_asqrt8_25[2]),.dout(n19930),.clk(gclk));
	jxor g19673(.dina(n19930),.dinb(w_n19236_0[0]),.dout(n19931),.clk(gclk));
	jand g19674(.dina(w_n19931_0[1]),.dinb(n19928),.dout(n19932),.clk(gclk));
	jor g19675(.dina(n19932),.dinb(w_n19927_0[1]),.dout(n19933),.clk(gclk));
	jand g19676(.dina(w_n19933_0[2]),.dinb(w_asqrt28_15[2]),.dout(n19934),.clk(gclk));
	jor g19677(.dina(w_n19933_0[1]),.dinb(w_asqrt28_15[1]),.dout(n19935),.clk(gclk));
	jxor g19678(.dina(w_n19239_0[0]),.dinb(w_n8890_23[0]),.dout(n19936),.clk(gclk));
	jand g19679(.dina(n19936),.dinb(w_asqrt8_25[1]),.dout(n19937),.clk(gclk));
	jxor g19680(.dina(n19937),.dinb(w_n19244_0[0]),.dout(n19938),.clk(gclk));
	jnot g19681(.din(w_n19938_0[1]),.dout(n19939),.clk(gclk));
	jand g19682(.dina(w_n19939_0[1]),.dinb(n19935),.dout(n19940),.clk(gclk));
	jor g19683(.dina(n19940),.dinb(w_n19934_0[1]),.dout(n19941),.clk(gclk));
	jand g19684(.dina(w_n19941_0[2]),.dinb(w_asqrt29_10[1]),.dout(n19942),.clk(gclk));
	jor g19685(.dina(w_n19941_0[1]),.dinb(w_asqrt29_10[0]),.dout(n19943),.clk(gclk));
	jxor g19686(.dina(w_n19246_0[0]),.dinb(w_n8449_18[0]),.dout(n19944),.clk(gclk));
	jand g19687(.dina(n19944),.dinb(w_asqrt8_25[0]),.dout(n19945),.clk(gclk));
	jxor g19688(.dina(n19945),.dinb(w_n19251_0[0]),.dout(n19946),.clk(gclk));
	jand g19689(.dina(w_n19946_0[1]),.dinb(n19943),.dout(n19947),.clk(gclk));
	jor g19690(.dina(n19947),.dinb(w_n19942_0[1]),.dout(n19948),.clk(gclk));
	jand g19691(.dina(w_n19948_0[2]),.dinb(w_asqrt30_16[0]),.dout(n19949),.clk(gclk));
	jor g19692(.dina(w_n19948_0[1]),.dinb(w_asqrt30_15[2]),.dout(n19950),.clk(gclk));
	jxor g19693(.dina(w_n19254_0[0]),.dinb(w_n8003_23[2]),.dout(n19951),.clk(gclk));
	jand g19694(.dina(n19951),.dinb(w_asqrt8_24[2]),.dout(n19952),.clk(gclk));
	jxor g19695(.dina(n19952),.dinb(w_n19259_0[0]),.dout(n19953),.clk(gclk));
	jnot g19696(.din(w_n19953_0[1]),.dout(n19954),.clk(gclk));
	jand g19697(.dina(w_n19954_0[1]),.dinb(n19950),.dout(n19955),.clk(gclk));
	jor g19698(.dina(n19955),.dinb(w_n19949_0[1]),.dout(n19956),.clk(gclk));
	jand g19699(.dina(w_n19956_0[2]),.dinb(w_asqrt31_11[0]),.dout(n19957),.clk(gclk));
	jor g19700(.dina(w_n19956_0[1]),.dinb(w_asqrt31_10[2]),.dout(n19958),.clk(gclk));
	jxor g19701(.dina(w_n19261_0[0]),.dinb(w_n7581_19[0]),.dout(n19959),.clk(gclk));
	jand g19702(.dina(n19959),.dinb(w_asqrt8_24[1]),.dout(n19960),.clk(gclk));
	jxor g19703(.dina(n19960),.dinb(w_n19266_0[0]),.dout(n19961),.clk(gclk));
	jnot g19704(.din(w_n19961_0[1]),.dout(n19962),.clk(gclk));
	jand g19705(.dina(w_n19962_0[1]),.dinb(n19958),.dout(n19963),.clk(gclk));
	jor g19706(.dina(n19963),.dinb(w_n19957_0[1]),.dout(n19964),.clk(gclk));
	jand g19707(.dina(w_n19964_0[2]),.dinb(w_asqrt32_16[0]),.dout(n19965),.clk(gclk));
	jor g19708(.dina(w_n19964_0[1]),.dinb(w_asqrt32_15[2]),.dout(n19966),.clk(gclk));
	jxor g19709(.dina(w_n19268_0[0]),.dinb(w_n7154_24[0]),.dout(n19967),.clk(gclk));
	jand g19710(.dina(n19967),.dinb(w_asqrt8_24[0]),.dout(n19968),.clk(gclk));
	jxor g19711(.dina(n19968),.dinb(w_n19273_0[0]),.dout(n19969),.clk(gclk));
	jnot g19712(.din(w_n19969_0[1]),.dout(n19970),.clk(gclk));
	jand g19713(.dina(w_n19970_0[1]),.dinb(n19966),.dout(n19971),.clk(gclk));
	jor g19714(.dina(n19971),.dinb(w_n19965_0[1]),.dout(n19972),.clk(gclk));
	jand g19715(.dina(w_n19972_0[2]),.dinb(w_asqrt33_11[2]),.dout(n19973),.clk(gclk));
	jor g19716(.dina(w_n19972_0[1]),.dinb(w_asqrt33_11[1]),.dout(n19974),.clk(gclk));
	jxor g19717(.dina(w_n19275_0[0]),.dinb(w_n6758_19[2]),.dout(n19975),.clk(gclk));
	jand g19718(.dina(n19975),.dinb(w_asqrt8_23[2]),.dout(n19976),.clk(gclk));
	jxor g19719(.dina(n19976),.dinb(w_n19280_0[0]),.dout(n19977),.clk(gclk));
	jand g19720(.dina(w_n19977_0[1]),.dinb(n19974),.dout(n19978),.clk(gclk));
	jor g19721(.dina(n19978),.dinb(w_n19973_0[1]),.dout(n19979),.clk(gclk));
	jand g19722(.dina(w_n19979_0[2]),.dinb(w_asqrt34_16[1]),.dout(n19980),.clk(gclk));
	jor g19723(.dina(w_n19979_0[1]),.dinb(w_asqrt34_16[0]),.dout(n19981),.clk(gclk));
	jxor g19724(.dina(w_n19283_0[0]),.dinb(w_n6357_24[1]),.dout(n19982),.clk(gclk));
	jand g19725(.dina(n19982),.dinb(w_asqrt8_23[1]),.dout(n19983),.clk(gclk));
	jxor g19726(.dina(n19983),.dinb(w_n19288_0[0]),.dout(n19984),.clk(gclk));
	jnot g19727(.din(w_n19984_0[1]),.dout(n19985),.clk(gclk));
	jand g19728(.dina(w_n19985_0[1]),.dinb(n19981),.dout(n19986),.clk(gclk));
	jor g19729(.dina(n19986),.dinb(w_n19980_0[1]),.dout(n19987),.clk(gclk));
	jand g19730(.dina(w_n19987_0[2]),.dinb(w_asqrt35_12[1]),.dout(n19988),.clk(gclk));
	jor g19731(.dina(w_n19987_0[1]),.dinb(w_asqrt35_12[0]),.dout(n19989),.clk(gclk));
	jxor g19732(.dina(w_n19290_0[0]),.dinb(w_n5989_20[1]),.dout(n19990),.clk(gclk));
	jand g19733(.dina(n19990),.dinb(w_asqrt8_23[0]),.dout(n19991),.clk(gclk));
	jxor g19734(.dina(n19991),.dinb(w_n19295_0[0]),.dout(n19992),.clk(gclk));
	jand g19735(.dina(w_n19992_0[1]),.dinb(n19989),.dout(n19993),.clk(gclk));
	jor g19736(.dina(n19993),.dinb(w_n19988_0[1]),.dout(n19994),.clk(gclk));
	jand g19737(.dina(w_n19994_0[2]),.dinb(w_asqrt36_16[1]),.dout(n19995),.clk(gclk));
	jor g19738(.dina(w_n19994_0[1]),.dinb(w_asqrt36_16[0]),.dout(n19996),.clk(gclk));
	jxor g19739(.dina(w_n19298_0[0]),.dinb(w_n5606_24[2]),.dout(n19997),.clk(gclk));
	jand g19740(.dina(n19997),.dinb(w_asqrt8_22[2]),.dout(n19998),.clk(gclk));
	jxor g19741(.dina(n19998),.dinb(w_n19303_0[0]),.dout(n19999),.clk(gclk));
	jnot g19742(.din(w_n19999_0[1]),.dout(n20000),.clk(gclk));
	jand g19743(.dina(w_n20000_0[1]),.dinb(n19996),.dout(n20001),.clk(gclk));
	jor g19744(.dina(n20001),.dinb(w_n19995_0[1]),.dout(n20002),.clk(gclk));
	jand g19745(.dina(w_n20002_0[2]),.dinb(w_asqrt37_12[2]),.dout(n20003),.clk(gclk));
	jor g19746(.dina(w_n20002_0[1]),.dinb(w_asqrt37_12[1]),.dout(n20004),.clk(gclk));
	jxor g19747(.dina(w_n19305_0[0]),.dinb(w_n5259_21[1]),.dout(n20005),.clk(gclk));
	jand g19748(.dina(n20005),.dinb(w_asqrt8_22[1]),.dout(n20006),.clk(gclk));
	jxor g19749(.dina(n20006),.dinb(w_n19310_0[0]),.dout(n20007),.clk(gclk));
	jand g19750(.dina(w_n20007_0[1]),.dinb(n20004),.dout(n20008),.clk(gclk));
	jor g19751(.dina(n20008),.dinb(w_n20003_0[1]),.dout(n20009),.clk(gclk));
	jand g19752(.dina(w_n20009_0[2]),.dinb(w_asqrt38_16[2]),.dout(n20010),.clk(gclk));
	jor g19753(.dina(w_n20009_0[1]),.dinb(w_asqrt38_16[1]),.dout(n20011),.clk(gclk));
	jxor g19754(.dina(w_n19313_0[0]),.dinb(w_n4902_25[1]),.dout(n20012),.clk(gclk));
	jand g19755(.dina(n20012),.dinb(w_asqrt8_22[0]),.dout(n20013),.clk(gclk));
	jxor g19756(.dina(n20013),.dinb(w_n19318_0[0]),.dout(n20014),.clk(gclk));
	jnot g19757(.din(w_n20014_0[1]),.dout(n20015),.clk(gclk));
	jand g19758(.dina(w_n20015_0[1]),.dinb(n20011),.dout(n20016),.clk(gclk));
	jor g19759(.dina(n20016),.dinb(w_n20010_0[1]),.dout(n20017),.clk(gclk));
	jand g19760(.dina(w_n20017_0[2]),.dinb(w_asqrt39_13[1]),.dout(n20018),.clk(gclk));
	jor g19761(.dina(w_n20017_0[1]),.dinb(w_asqrt39_13[0]),.dout(n20019),.clk(gclk));
	jxor g19762(.dina(w_n19320_0[0]),.dinb(w_n4582_22[1]),.dout(n20020),.clk(gclk));
	jand g19763(.dina(n20020),.dinb(w_asqrt8_21[2]),.dout(n20021),.clk(gclk));
	jxor g19764(.dina(n20021),.dinb(w_n19325_0[0]),.dout(n20022),.clk(gclk));
	jand g19765(.dina(w_n20022_0[1]),.dinb(n20019),.dout(n20023),.clk(gclk));
	jor g19766(.dina(n20023),.dinb(w_n20018_0[1]),.dout(n20024),.clk(gclk));
	jand g19767(.dina(w_n20024_0[2]),.dinb(w_asqrt40_16[2]),.dout(n20025),.clk(gclk));
	jor g19768(.dina(w_n20024_0[1]),.dinb(w_asqrt40_16[1]),.dout(n20026),.clk(gclk));
	jxor g19769(.dina(w_n19328_0[0]),.dinb(w_n4249_26[0]),.dout(n20027),.clk(gclk));
	jand g19770(.dina(n20027),.dinb(w_asqrt8_21[1]),.dout(n20028),.clk(gclk));
	jxor g19771(.dina(n20028),.dinb(w_n19333_0[0]),.dout(n20029),.clk(gclk));
	jnot g19772(.din(w_n20029_0[1]),.dout(n20030),.clk(gclk));
	jand g19773(.dina(w_n20030_0[1]),.dinb(n20026),.dout(n20031),.clk(gclk));
	jor g19774(.dina(n20031),.dinb(w_n20025_0[1]),.dout(n20032),.clk(gclk));
	jand g19775(.dina(w_n20032_0[2]),.dinb(w_asqrt41_13[2]),.dout(n20033),.clk(gclk));
	jor g19776(.dina(w_n20032_0[1]),.dinb(w_asqrt41_13[1]),.dout(n20034),.clk(gclk));
	jxor g19777(.dina(w_n19335_0[0]),.dinb(w_n3955_23[0]),.dout(n20035),.clk(gclk));
	jand g19778(.dina(n20035),.dinb(w_asqrt8_21[0]),.dout(n20036),.clk(gclk));
	jxor g19779(.dina(n20036),.dinb(w_n19340_0[0]),.dout(n20037),.clk(gclk));
	jnot g19780(.din(w_n20037_0[1]),.dout(n20038),.clk(gclk));
	jand g19781(.dina(w_n20038_0[1]),.dinb(n20034),.dout(n20039),.clk(gclk));
	jor g19782(.dina(n20039),.dinb(w_n20033_0[1]),.dout(n20040),.clk(gclk));
	jand g19783(.dina(w_n20040_0[2]),.dinb(w_asqrt42_17[0]),.dout(n20041),.clk(gclk));
	jor g19784(.dina(w_n20040_0[1]),.dinb(w_asqrt42_16[2]),.dout(n20042),.clk(gclk));
	jxor g19785(.dina(w_n19342_0[0]),.dinb(w_n3642_26[1]),.dout(n20043),.clk(gclk));
	jand g19786(.dina(n20043),.dinb(w_asqrt8_20[2]),.dout(n20044),.clk(gclk));
	jxor g19787(.dina(n20044),.dinb(w_n19347_0[0]),.dout(n20045),.clk(gclk));
	jnot g19788(.din(w_n20045_0[1]),.dout(n20046),.clk(gclk));
	jand g19789(.dina(w_n20046_0[1]),.dinb(n20042),.dout(n20047),.clk(gclk));
	jor g19790(.dina(n20047),.dinb(w_n20041_0[1]),.dout(n20048),.clk(gclk));
	jand g19791(.dina(w_n20048_0[2]),.dinb(w_asqrt43_14[0]),.dout(n20049),.clk(gclk));
	jor g19792(.dina(w_n20048_0[1]),.dinb(w_asqrt43_13[2]),.dout(n20050),.clk(gclk));
	jxor g19793(.dina(w_n19349_0[0]),.dinb(w_n3368_23[2]),.dout(n20051),.clk(gclk));
	jand g19794(.dina(n20051),.dinb(w_asqrt8_20[1]),.dout(n20052),.clk(gclk));
	jxor g19795(.dina(n20052),.dinb(w_n19354_0[0]),.dout(n20053),.clk(gclk));
	jand g19796(.dina(w_n20053_0[1]),.dinb(n20050),.dout(n20054),.clk(gclk));
	jor g19797(.dina(n20054),.dinb(w_n20049_0[1]),.dout(n20055),.clk(gclk));
	jand g19798(.dina(w_n20055_0[2]),.dinb(w_asqrt44_17[0]),.dout(n20056),.clk(gclk));
	jor g19799(.dina(w_n20055_0[1]),.dinb(w_asqrt44_16[2]),.dout(n20057),.clk(gclk));
	jxor g19800(.dina(w_n19357_0[0]),.dinb(w_n3089_27[0]),.dout(n20058),.clk(gclk));
	jand g19801(.dina(n20058),.dinb(w_asqrt8_20[0]),.dout(n20059),.clk(gclk));
	jxor g19802(.dina(n20059),.dinb(w_n19362_0[0]),.dout(n20060),.clk(gclk));
	jnot g19803(.din(w_n20060_0[1]),.dout(n20061),.clk(gclk));
	jand g19804(.dina(w_n20061_0[1]),.dinb(n20057),.dout(n20062),.clk(gclk));
	jor g19805(.dina(n20062),.dinb(w_n20056_0[1]),.dout(n20063),.clk(gclk));
	jand g19806(.dina(w_n20063_0[2]),.dinb(w_asqrt45_14[2]),.dout(n20064),.clk(gclk));
	jor g19807(.dina(w_n20063_0[1]),.dinb(w_asqrt45_14[1]),.dout(n20065),.clk(gclk));
	jxor g19808(.dina(w_n19364_0[0]),.dinb(w_n2833_24[2]),.dout(n20066),.clk(gclk));
	jand g19809(.dina(n20066),.dinb(w_asqrt8_19[2]),.dout(n20067),.clk(gclk));
	jxor g19810(.dina(n20067),.dinb(w_n19369_0[0]),.dout(n20068),.clk(gclk));
	jnot g19811(.din(w_n20068_0[1]),.dout(n20069),.clk(gclk));
	jand g19812(.dina(w_n20069_0[1]),.dinb(n20065),.dout(n20070),.clk(gclk));
	jor g19813(.dina(n20070),.dinb(w_n20064_0[1]),.dout(n20071),.clk(gclk));
	jand g19814(.dina(w_n20071_0[2]),.dinb(w_asqrt46_17[0]),.dout(n20072),.clk(gclk));
	jor g19815(.dina(w_n20071_0[1]),.dinb(w_asqrt46_16[2]),.dout(n20073),.clk(gclk));
	jxor g19816(.dina(w_n19371_0[0]),.dinb(w_n2572_27[1]),.dout(n20074),.clk(gclk));
	jand g19817(.dina(n20074),.dinb(w_asqrt8_19[1]),.dout(n20075),.clk(gclk));
	jxor g19818(.dina(n20075),.dinb(w_n19376_0[0]),.dout(n20076),.clk(gclk));
	jnot g19819(.din(w_n20076_0[1]),.dout(n20077),.clk(gclk));
	jand g19820(.dina(w_n20077_0[1]),.dinb(n20073),.dout(n20078),.clk(gclk));
	jor g19821(.dina(n20078),.dinb(w_n20072_0[1]),.dout(n20079),.clk(gclk));
	jand g19822(.dina(w_n20079_0[2]),.dinb(w_asqrt47_15[1]),.dout(n20080),.clk(gclk));
	jor g19823(.dina(w_n20079_0[1]),.dinb(w_asqrt47_15[0]),.dout(n20081),.clk(gclk));
	jxor g19824(.dina(w_n19378_0[0]),.dinb(w_n2345_25[1]),.dout(n20082),.clk(gclk));
	jand g19825(.dina(n20082),.dinb(w_asqrt8_19[0]),.dout(n20083),.clk(gclk));
	jxor g19826(.dina(n20083),.dinb(w_n19383_0[0]),.dout(n20084),.clk(gclk));
	jnot g19827(.din(w_n20084_0[1]),.dout(n20085),.clk(gclk));
	jand g19828(.dina(w_n20085_0[1]),.dinb(n20081),.dout(n20086),.clk(gclk));
	jor g19829(.dina(n20086),.dinb(w_n20080_0[1]),.dout(n20087),.clk(gclk));
	jand g19830(.dina(w_n20087_0[2]),.dinb(w_asqrt48_17[1]),.dout(n20088),.clk(gclk));
	jor g19831(.dina(w_n20087_0[1]),.dinb(w_asqrt48_17[0]),.dout(n20089),.clk(gclk));
	jxor g19832(.dina(w_n19385_0[0]),.dinb(w_n2108_28[0]),.dout(n20090),.clk(gclk));
	jand g19833(.dina(n20090),.dinb(w_asqrt8_18[2]),.dout(n20091),.clk(gclk));
	jxor g19834(.dina(n20091),.dinb(w_n19390_0[0]),.dout(n20092),.clk(gclk));
	jnot g19835(.din(w_n20092_0[1]),.dout(n20093),.clk(gclk));
	jand g19836(.dina(w_n20093_0[1]),.dinb(n20089),.dout(n20094),.clk(gclk));
	jor g19837(.dina(n20094),.dinb(w_n20088_0[1]),.dout(n20095),.clk(gclk));
	jand g19838(.dina(w_n20095_0[2]),.dinb(w_asqrt49_15[2]),.dout(n20096),.clk(gclk));
	jor g19839(.dina(w_n20095_0[1]),.dinb(w_asqrt49_15[1]),.dout(n20097),.clk(gclk));
	jxor g19840(.dina(w_n19392_0[0]),.dinb(w_n1912_26[1]),.dout(n20098),.clk(gclk));
	jand g19841(.dina(n20098),.dinb(w_asqrt8_18[1]),.dout(n20099),.clk(gclk));
	jxor g19842(.dina(n20099),.dinb(w_n19397_0[0]),.dout(n20100),.clk(gclk));
	jand g19843(.dina(w_n20100_0[1]),.dinb(n20097),.dout(n20101),.clk(gclk));
	jor g19844(.dina(n20101),.dinb(w_n20096_0[1]),.dout(n20102),.clk(gclk));
	jand g19845(.dina(w_n20102_0[2]),.dinb(w_asqrt50_17[2]),.dout(n20103),.clk(gclk));
	jor g19846(.dina(w_n20102_0[1]),.dinb(w_asqrt50_17[1]),.dout(n20104),.clk(gclk));
	jxor g19847(.dina(w_n19400_0[0]),.dinb(w_n1699_28[2]),.dout(n20105),.clk(gclk));
	jand g19848(.dina(n20105),.dinb(w_asqrt8_18[0]),.dout(n20106),.clk(gclk));
	jxor g19849(.dina(n20106),.dinb(w_n19405_0[0]),.dout(n20107),.clk(gclk));
	jnot g19850(.din(w_n20107_0[1]),.dout(n20108),.clk(gclk));
	jand g19851(.dina(w_n20108_0[1]),.dinb(n20104),.dout(n20109),.clk(gclk));
	jor g19852(.dina(n20109),.dinb(w_n20103_0[1]),.dout(n20110),.clk(gclk));
	jand g19853(.dina(w_n20110_0[2]),.dinb(w_asqrt51_16[0]),.dout(n20111),.clk(gclk));
	jor g19854(.dina(w_n20110_0[1]),.dinb(w_asqrt51_15[2]),.dout(n20112),.clk(gclk));
	jxor g19855(.dina(w_n19407_0[0]),.dinb(w_n1516_27[0]),.dout(n20113),.clk(gclk));
	jand g19856(.dina(n20113),.dinb(w_asqrt8_17[2]),.dout(n20114),.clk(gclk));
	jxor g19857(.dina(n20114),.dinb(w_n19412_0[0]),.dout(n20115),.clk(gclk));
	jand g19858(.dina(w_n20115_0[1]),.dinb(n20112),.dout(n20116),.clk(gclk));
	jor g19859(.dina(n20116),.dinb(w_n20111_0[1]),.dout(n20117),.clk(gclk));
	jand g19860(.dina(w_n20117_0[2]),.dinb(w_asqrt52_17[2]),.dout(n20118),.clk(gclk));
	jor g19861(.dina(w_n20117_0[1]),.dinb(w_asqrt52_17[1]),.dout(n20119),.clk(gclk));
	jxor g19862(.dina(w_n19415_0[0]),.dinb(w_n1332_28[2]),.dout(n20120),.clk(gclk));
	jand g19863(.dina(n20120),.dinb(w_asqrt8_17[1]),.dout(n20121),.clk(gclk));
	jxor g19864(.dina(n20121),.dinb(w_n19420_0[0]),.dout(n20122),.clk(gclk));
	jnot g19865(.din(w_n20122_0[1]),.dout(n20123),.clk(gclk));
	jand g19866(.dina(w_n20123_0[1]),.dinb(n20119),.dout(n20124),.clk(gclk));
	jor g19867(.dina(n20124),.dinb(w_n20118_0[1]),.dout(n20125),.clk(gclk));
	jand g19868(.dina(w_n20125_0[2]),.dinb(w_asqrt53_16[2]),.dout(n20126),.clk(gclk));
	jor g19869(.dina(w_n20125_0[1]),.dinb(w_asqrt53_16[1]),.dout(n20127),.clk(gclk));
	jxor g19870(.dina(w_n19422_0[0]),.dinb(w_n1173_27[2]),.dout(n20128),.clk(gclk));
	jand g19871(.dina(n20128),.dinb(w_asqrt8_17[0]),.dout(n20129),.clk(gclk));
	jxor g19872(.dina(n20129),.dinb(w_n19427_0[0]),.dout(n20130),.clk(gclk));
	jnot g19873(.din(w_n20130_0[1]),.dout(n20131),.clk(gclk));
	jand g19874(.dina(w_n20131_0[1]),.dinb(n20127),.dout(n20132),.clk(gclk));
	jor g19875(.dina(n20132),.dinb(w_n20126_0[1]),.dout(n20133),.clk(gclk));
	jand g19876(.dina(w_n20133_0[2]),.dinb(w_asqrt54_17[2]),.dout(n20134),.clk(gclk));
	jor g19877(.dina(w_n20133_0[1]),.dinb(w_asqrt54_17[1]),.dout(n20135),.clk(gclk));
	jxor g19878(.dina(w_n19429_0[0]),.dinb(w_n1008_29[2]),.dout(n20136),.clk(gclk));
	jand g19879(.dina(n20136),.dinb(w_asqrt8_16[2]),.dout(n20137),.clk(gclk));
	jxor g19880(.dina(n20137),.dinb(w_n19434_0[0]),.dout(n20138),.clk(gclk));
	jand g19881(.dina(w_n20138_0[1]),.dinb(n20135),.dout(n20139),.clk(gclk));
	jor g19882(.dina(n20139),.dinb(w_n20134_0[1]),.dout(n20140),.clk(gclk));
	jand g19883(.dina(w_n20140_0[2]),.dinb(w_asqrt55_17[0]),.dout(n20141),.clk(gclk));
	jxor g19884(.dina(w_n19437_0[0]),.dinb(w_n884_28[2]),.dout(n20142),.clk(gclk));
	jand g19885(.dina(n20142),.dinb(w_asqrt8_16[1]),.dout(n20143),.clk(gclk));
	jxor g19886(.dina(n20143),.dinb(w_n19441_0[0]),.dout(n20144),.clk(gclk));
	jor g19887(.dina(w_n20140_0[1]),.dinb(w_asqrt55_16[2]),.dout(n20145),.clk(gclk));
	jand g19888(.dina(n20145),.dinb(w_n20144_0[1]),.dout(n20146),.clk(gclk));
	jor g19889(.dina(n20146),.dinb(w_n20141_0[1]),.dout(n20147),.clk(gclk));
	jand g19890(.dina(w_n20147_0[2]),.dinb(w_asqrt56_18[0]),.dout(n20148),.clk(gclk));
	jor g19891(.dina(w_n20147_0[1]),.dinb(w_asqrt56_17[2]),.dout(n20149),.clk(gclk));
	jxor g19892(.dina(w_n19445_0[0]),.dinb(w_n743_29[2]),.dout(n20150),.clk(gclk));
	jand g19893(.dina(n20150),.dinb(w_asqrt8_16[0]),.dout(n20151),.clk(gclk));
	jxor g19894(.dina(n20151),.dinb(w_n19450_0[0]),.dout(n20152),.clk(gclk));
	jnot g19895(.din(w_n20152_0[1]),.dout(n20153),.clk(gclk));
	jand g19896(.dina(w_n20153_0[1]),.dinb(n20149),.dout(n20154),.clk(gclk));
	jor g19897(.dina(n20154),.dinb(w_n20148_0[1]),.dout(n20155),.clk(gclk));
	jand g19898(.dina(w_n20155_0[2]),.dinb(w_asqrt57_17[2]),.dout(n20156),.clk(gclk));
	jor g19899(.dina(w_n20155_0[1]),.dinb(w_asqrt57_17[1]),.dout(n20157),.clk(gclk));
	jxor g19900(.dina(w_n19452_0[0]),.dinb(w_n635_29[2]),.dout(n20158),.clk(gclk));
	jand g19901(.dina(n20158),.dinb(w_asqrt8_15[2]),.dout(n20159),.clk(gclk));
	jxor g19902(.dina(n20159),.dinb(w_n19457_0[0]),.dout(n20160),.clk(gclk));
	jand g19903(.dina(w_n20160_0[1]),.dinb(n20157),.dout(n20161),.clk(gclk));
	jor g19904(.dina(n20161),.dinb(w_n20156_0[1]),.dout(n20162),.clk(gclk));
	jand g19905(.dina(w_n20162_0[2]),.dinb(w_asqrt58_18[1]),.dout(n20163),.clk(gclk));
	jor g19906(.dina(w_n20162_0[1]),.dinb(w_asqrt58_18[0]),.dout(n20164),.clk(gclk));
	jxor g19907(.dina(w_n19460_0[0]),.dinb(w_n515_30[2]),.dout(n20165),.clk(gclk));
	jand g19908(.dina(n20165),.dinb(w_asqrt8_15[1]),.dout(n20166),.clk(gclk));
	jxor g19909(.dina(n20166),.dinb(w_n19465_0[0]),.dout(n20167),.clk(gclk));
	jnot g19910(.din(w_n20167_0[1]),.dout(n20168),.clk(gclk));
	jand g19911(.dina(w_n20168_0[1]),.dinb(n20164),.dout(n20169),.clk(gclk));
	jor g19912(.dina(n20169),.dinb(w_n20163_0[1]),.dout(n20170),.clk(gclk));
	jand g19913(.dina(w_n20170_0[2]),.dinb(w_asqrt59_18[0]),.dout(n20171),.clk(gclk));
	jor g19914(.dina(w_n20170_0[1]),.dinb(w_asqrt59_17[2]),.dout(n20172),.clk(gclk));
	jxor g19915(.dina(w_n19467_0[0]),.dinb(w_n443_30[2]),.dout(n20173),.clk(gclk));
	jand g19916(.dina(n20173),.dinb(w_asqrt8_15[0]),.dout(n20174),.clk(gclk));
	jxor g19917(.dina(n20174),.dinb(w_n19473_0[0]),.dout(n20175),.clk(gclk));
	jnot g19918(.din(w_n20175_0[1]),.dout(n20176),.clk(gclk));
	jand g19919(.dina(w_n20176_0[1]),.dinb(n20172),.dout(n20177),.clk(gclk));
	jor g19920(.dina(n20177),.dinb(w_n20171_0[1]),.dout(n20178),.clk(gclk));
	jand g19921(.dina(w_n20178_0[2]),.dinb(w_asqrt60_18[1]),.dout(n20179),.clk(gclk));
	jor g19922(.dina(w_n20178_0[1]),.dinb(w_asqrt60_18[0]),.dout(n20180),.clk(gclk));
	jxor g19923(.dina(w_n19475_0[0]),.dinb(w_n352_31[0]),.dout(n20181),.clk(gclk));
	jand g19924(.dina(n20181),.dinb(w_asqrt8_14[2]),.dout(n20182),.clk(gclk));
	jxor g19925(.dina(n20182),.dinb(w_n19480_0[0]),.dout(n20183),.clk(gclk));
	jand g19926(.dina(w_n20183_0[1]),.dinb(n20180),.dout(n20184),.clk(gclk));
	jor g19927(.dina(n20184),.dinb(w_n20179_0[1]),.dout(n20185),.clk(gclk));
	jand g19928(.dina(w_n20185_0[2]),.dinb(w_asqrt61_18[1]),.dout(n20186),.clk(gclk));
	jor g19929(.dina(w_n20185_0[1]),.dinb(w_asqrt61_18[0]),.dout(n20187),.clk(gclk));
	jxor g19930(.dina(w_n19483_0[0]),.dinb(w_n294_31[1]),.dout(n20188),.clk(gclk));
	jand g19931(.dina(n20188),.dinb(w_asqrt8_14[1]),.dout(n20189),.clk(gclk));
	jxor g19932(.dina(n20189),.dinb(w_n19488_0[0]),.dout(n20190),.clk(gclk));
	jnot g19933(.din(w_n20190_0[1]),.dout(n20191),.clk(gclk));
	jand g19934(.dina(w_n20191_0[1]),.dinb(n20187),.dout(n20192),.clk(gclk));
	jor g19935(.dina(n20192),.dinb(w_n20186_0[1]),.dout(n20193),.clk(gclk));
	jand g19936(.dina(w_n20193_0[2]),.dinb(w_asqrt62_18[1]),.dout(n20194),.clk(gclk));
	jnot g19937(.din(w_n20194_0[1]),.dout(n20195),.clk(gclk));
	jnot g19938(.din(w_n20186_0[0]),.dout(n20196),.clk(gclk));
	jnot g19939(.din(w_n20179_0[0]),.dout(n20197),.clk(gclk));
	jnot g19940(.din(w_n20171_0[0]),.dout(n20198),.clk(gclk));
	jnot g19941(.din(w_n20163_0[0]),.dout(n20199),.clk(gclk));
	jnot g19942(.din(w_n20156_0[0]),.dout(n20200),.clk(gclk));
	jnot g19943(.din(w_n20148_0[0]),.dout(n20201),.clk(gclk));
	jnot g19944(.din(w_n20141_0[0]),.dout(n20202),.clk(gclk));
	jnot g19945(.din(w_n20144_0[0]),.dout(n20203),.clk(gclk));
	jnot g19946(.din(w_n20134_0[0]),.dout(n20204),.clk(gclk));
	jnot g19947(.din(w_n20126_0[0]),.dout(n20205),.clk(gclk));
	jnot g19948(.din(w_n20118_0[0]),.dout(n20206),.clk(gclk));
	jnot g19949(.din(w_n20111_0[0]),.dout(n20207),.clk(gclk));
	jnot g19950(.din(w_n20103_0[0]),.dout(n20208),.clk(gclk));
	jnot g19951(.din(w_n20096_0[0]),.dout(n20209),.clk(gclk));
	jnot g19952(.din(w_n20088_0[0]),.dout(n20210),.clk(gclk));
	jnot g19953(.din(w_n20080_0[0]),.dout(n20211),.clk(gclk));
	jnot g19954(.din(w_n20072_0[0]),.dout(n20212),.clk(gclk));
	jnot g19955(.din(w_n20064_0[0]),.dout(n20213),.clk(gclk));
	jnot g19956(.din(w_n20056_0[0]),.dout(n20214),.clk(gclk));
	jnot g19957(.din(w_n20049_0[0]),.dout(n20215),.clk(gclk));
	jnot g19958(.din(w_n20041_0[0]),.dout(n20216),.clk(gclk));
	jnot g19959(.din(w_n20033_0[0]),.dout(n20217),.clk(gclk));
	jnot g19960(.din(w_n20025_0[0]),.dout(n20218),.clk(gclk));
	jnot g19961(.din(w_n20018_0[0]),.dout(n20219),.clk(gclk));
	jnot g19962(.din(w_n20010_0[0]),.dout(n20220),.clk(gclk));
	jnot g19963(.din(w_n20003_0[0]),.dout(n20221),.clk(gclk));
	jnot g19964(.din(w_n19995_0[0]),.dout(n20222),.clk(gclk));
	jnot g19965(.din(w_n19988_0[0]),.dout(n20223),.clk(gclk));
	jnot g19966(.din(w_n19980_0[0]),.dout(n20224),.clk(gclk));
	jnot g19967(.din(w_n19973_0[0]),.dout(n20225),.clk(gclk));
	jnot g19968(.din(w_n19965_0[0]),.dout(n20226),.clk(gclk));
	jnot g19969(.din(w_n19957_0[0]),.dout(n20227),.clk(gclk));
	jnot g19970(.din(w_n19949_0[0]),.dout(n20228),.clk(gclk));
	jnot g19971(.din(w_n19942_0[0]),.dout(n20229),.clk(gclk));
	jnot g19972(.din(w_n19934_0[0]),.dout(n20230),.clk(gclk));
	jnot g19973(.din(w_n19927_0[0]),.dout(n20231),.clk(gclk));
	jnot g19974(.din(w_n19919_0[0]),.dout(n20232),.clk(gclk));
	jnot g19975(.din(w_n19912_0[0]),.dout(n20233),.clk(gclk));
	jnot g19976(.din(w_n19905_0[0]),.dout(n20234),.clk(gclk));
	jnot g19977(.din(w_n19897_0[0]),.dout(n20235),.clk(gclk));
	jnot g19978(.din(w_n19889_0[0]),.dout(n20236),.clk(gclk));
	jnot g19979(.din(w_n19882_0[0]),.dout(n20237),.clk(gclk));
	jnot g19980(.din(w_n19874_0[0]),.dout(n20238),.clk(gclk));
	jnot g19981(.din(w_n19867_0[0]),.dout(n20239),.clk(gclk));
	jnot g19982(.din(w_n19859_0[0]),.dout(n20240),.clk(gclk));
	jnot g19983(.din(w_n19852_0[0]),.dout(n20241),.clk(gclk));
	jnot g19984(.din(w_n19844_0[0]),.dout(n20242),.clk(gclk));
	jnot g19985(.din(w_n19837_0[0]),.dout(n20243),.clk(gclk));
	jnot g19986(.din(w_n19829_0[0]),.dout(n20244),.clk(gclk));
	jnot g19987(.din(w_n19822_0[0]),.dout(n20245),.clk(gclk));
	jnot g19988(.din(w_n19814_0[0]),.dout(n20246),.clk(gclk));
	jnot g19989(.din(w_n19806_0[0]),.dout(n20247),.clk(gclk));
	jnot g19990(.din(w_n19796_0[0]),.dout(n20248),.clk(gclk));
	jnot g19991(.din(w_n19530_0[0]),.dout(n20249),.clk(gclk));
	jnot g19992(.din(w_n19527_0[0]),.dout(n20250),.clk(gclk));
	jor g19993(.dina(w_n19791_10[1]),.dinb(w_n19101_0[2]),.dout(n20251),.clk(gclk));
	jand g19994(.dina(n20251),.dinb(n20250),.dout(n20252),.clk(gclk));
	jand g19995(.dina(n20252),.dinb(w_n19096_18[0]),.dout(n20253),.clk(gclk));
	jor g19996(.dina(w_n19791_10[0]),.dinb(w_a16_0[0]),.dout(n20254),.clk(gclk));
	jand g19997(.dina(n20254),.dinb(w_a17_0[0]),.dout(n20255),.clk(gclk));
	jor g19998(.dina(w_n19798_0[0]),.dinb(n20255),.dout(n20256),.clk(gclk));
	jor g19999(.dina(w_n20256_0[1]),.dinb(n20253),.dout(n20257),.clk(gclk));
	jand g20000(.dina(n20257),.dinb(n20249),.dout(n20258),.clk(gclk));
	jand g20001(.dina(n20258),.dinb(w_n18442_10[0]),.dout(n20259),.clk(gclk));
	jor g20002(.dina(w_n19802_0[0]),.dinb(n20259),.dout(n20260),.clk(gclk));
	jand g20003(.dina(n20260),.dinb(n20248),.dout(n20261),.clk(gclk));
	jand g20004(.dina(n20261),.dinb(w_n17769_18[2]),.dout(n20262),.clk(gclk));
	jor g20005(.dina(w_n19810_0[0]),.dinb(n20262),.dout(n20263),.clk(gclk));
	jand g20006(.dina(n20263),.dinb(n20247),.dout(n20264),.clk(gclk));
	jand g20007(.dina(n20264),.dinb(w_n17134_11[0]),.dout(n20265),.clk(gclk));
	jor g20008(.dina(w_n19818_0[0]),.dinb(n20265),.dout(n20266),.clk(gclk));
	jand g20009(.dina(n20266),.dinb(n20246),.dout(n20267),.clk(gclk));
	jand g20010(.dina(n20267),.dinb(w_n16489_19[0]),.dout(n20268),.clk(gclk));
	jnot g20011(.din(w_n19826_0[0]),.dout(n20269),.clk(gclk));
	jor g20012(.dina(w_n20269_0[1]),.dinb(n20268),.dout(n20270),.clk(gclk));
	jand g20013(.dina(n20270),.dinb(n20245),.dout(n20271),.clk(gclk));
	jand g20014(.dina(n20271),.dinb(w_n15878_12[0]),.dout(n20272),.clk(gclk));
	jor g20015(.dina(w_n19833_0[0]),.dinb(n20272),.dout(n20273),.clk(gclk));
	jand g20016(.dina(n20273),.dinb(n20244),.dout(n20274),.clk(gclk));
	jand g20017(.dina(n20274),.dinb(w_n15260_19[2]),.dout(n20275),.clk(gclk));
	jnot g20018(.din(w_n19841_0[0]),.dout(n20276),.clk(gclk));
	jor g20019(.dina(w_n20276_0[1]),.dinb(n20275),.dout(n20277),.clk(gclk));
	jand g20020(.dina(n20277),.dinb(n20243),.dout(n20278),.clk(gclk));
	jand g20021(.dina(n20278),.dinb(w_n14674_12[2]),.dout(n20279),.clk(gclk));
	jor g20022(.dina(w_n19848_0[0]),.dinb(n20279),.dout(n20280),.clk(gclk));
	jand g20023(.dina(n20280),.dinb(n20242),.dout(n20281),.clk(gclk));
	jand g20024(.dina(n20281),.dinb(w_n14078_20[0]),.dout(n20282),.clk(gclk));
	jnot g20025(.din(w_n19856_0[0]),.dout(n20283),.clk(gclk));
	jor g20026(.dina(w_n20283_0[1]),.dinb(n20282),.dout(n20284),.clk(gclk));
	jand g20027(.dina(n20284),.dinb(n20241),.dout(n20285),.clk(gclk));
	jand g20028(.dina(n20285),.dinb(w_n13515_13[2]),.dout(n20286),.clk(gclk));
	jor g20029(.dina(w_n19863_0[0]),.dinb(n20286),.dout(n20287),.clk(gclk));
	jand g20030(.dina(n20287),.dinb(n20240),.dout(n20288),.clk(gclk));
	jand g20031(.dina(n20288),.dinb(w_n12947_20[2]),.dout(n20289),.clk(gclk));
	jnot g20032(.din(w_n19871_0[0]),.dout(n20290),.clk(gclk));
	jor g20033(.dina(w_n20290_0[1]),.dinb(n20289),.dout(n20291),.clk(gclk));
	jand g20034(.dina(n20291),.dinb(n20239),.dout(n20292),.clk(gclk));
	jand g20035(.dina(n20292),.dinb(w_n12410_14[1]),.dout(n20293),.clk(gclk));
	jor g20036(.dina(w_n19878_0[0]),.dinb(n20293),.dout(n20294),.clk(gclk));
	jand g20037(.dina(n20294),.dinb(n20238),.dout(n20295),.clk(gclk));
	jand g20038(.dina(n20295),.dinb(w_n11858_21[0]),.dout(n20296),.clk(gclk));
	jnot g20039(.din(w_n19886_0[0]),.dout(n20297),.clk(gclk));
	jor g20040(.dina(w_n20297_0[1]),.dinb(n20296),.dout(n20298),.clk(gclk));
	jand g20041(.dina(n20298),.dinb(n20237),.dout(n20299),.clk(gclk));
	jand g20042(.dina(n20299),.dinb(w_n11347_15[0]),.dout(n20300),.clk(gclk));
	jor g20043(.dina(w_n19893_0[0]),.dinb(n20300),.dout(n20301),.clk(gclk));
	jand g20044(.dina(n20301),.dinb(n20236),.dout(n20302),.clk(gclk));
	jand g20045(.dina(n20302),.dinb(w_n10824_21[2]),.dout(n20303),.clk(gclk));
	jor g20046(.dina(w_n19901_0[0]),.dinb(n20303),.dout(n20304),.clk(gclk));
	jand g20047(.dina(n20304),.dinb(n20235),.dout(n20305),.clk(gclk));
	jand g20048(.dina(n20305),.dinb(w_n10328_16[0]),.dout(n20306),.clk(gclk));
	jnot g20049(.din(w_n19909_0[0]),.dout(n20307),.clk(gclk));
	jor g20050(.dina(w_n20307_0[1]),.dinb(n20306),.dout(n20308),.clk(gclk));
	jand g20051(.dina(n20308),.dinb(n20234),.dout(n20309),.clk(gclk));
	jand g20052(.dina(n20309),.dinb(w_n9832_22[1]),.dout(n20310),.clk(gclk));
	jnot g20053(.din(w_n19916_0[0]),.dout(n20311),.clk(gclk));
	jor g20054(.dina(w_n20311_0[1]),.dinb(n20310),.dout(n20312),.clk(gclk));
	jand g20055(.dina(n20312),.dinb(n20233),.dout(n20313),.clk(gclk));
	jand g20056(.dina(n20313),.dinb(w_n9369_17[0]),.dout(n20314),.clk(gclk));
	jor g20057(.dina(w_n19923_0[0]),.dinb(n20314),.dout(n20315),.clk(gclk));
	jand g20058(.dina(n20315),.dinb(n20232),.dout(n20316),.clk(gclk));
	jand g20059(.dina(n20316),.dinb(w_n8890_22[2]),.dout(n20317),.clk(gclk));
	jnot g20060(.din(w_n19931_0[0]),.dout(n20318),.clk(gclk));
	jor g20061(.dina(w_n20318_0[1]),.dinb(n20317),.dout(n20319),.clk(gclk));
	jand g20062(.dina(n20319),.dinb(n20231),.dout(n20320),.clk(gclk));
	jand g20063(.dina(n20320),.dinb(w_n8449_17[2]),.dout(n20321),.clk(gclk));
	jor g20064(.dina(w_n19938_0[0]),.dinb(n20321),.dout(n20322),.clk(gclk));
	jand g20065(.dina(n20322),.dinb(n20230),.dout(n20323),.clk(gclk));
	jand g20066(.dina(n20323),.dinb(w_n8003_23[1]),.dout(n20324),.clk(gclk));
	jnot g20067(.din(w_n19946_0[0]),.dout(n20325),.clk(gclk));
	jor g20068(.dina(w_n20325_0[1]),.dinb(n20324),.dout(n20326),.clk(gclk));
	jand g20069(.dina(n20326),.dinb(n20229),.dout(n20327),.clk(gclk));
	jand g20070(.dina(n20327),.dinb(w_n7581_18[2]),.dout(n20328),.clk(gclk));
	jor g20071(.dina(w_n19953_0[0]),.dinb(n20328),.dout(n20329),.clk(gclk));
	jand g20072(.dina(n20329),.dinb(n20228),.dout(n20330),.clk(gclk));
	jand g20073(.dina(n20330),.dinb(w_n7154_23[2]),.dout(n20331),.clk(gclk));
	jor g20074(.dina(w_n19961_0[0]),.dinb(n20331),.dout(n20332),.clk(gclk));
	jand g20075(.dina(n20332),.dinb(n20227),.dout(n20333),.clk(gclk));
	jand g20076(.dina(n20333),.dinb(w_n6758_19[1]),.dout(n20334),.clk(gclk));
	jor g20077(.dina(w_n19969_0[0]),.dinb(n20334),.dout(n20335),.clk(gclk));
	jand g20078(.dina(n20335),.dinb(n20226),.dout(n20336),.clk(gclk));
	jand g20079(.dina(n20336),.dinb(w_n6357_24[0]),.dout(n20337),.clk(gclk));
	jnot g20080(.din(w_n19977_0[0]),.dout(n20338),.clk(gclk));
	jor g20081(.dina(w_n20338_0[1]),.dinb(n20337),.dout(n20339),.clk(gclk));
	jand g20082(.dina(n20339),.dinb(n20225),.dout(n20340),.clk(gclk));
	jand g20083(.dina(n20340),.dinb(w_n5989_20[0]),.dout(n20341),.clk(gclk));
	jor g20084(.dina(w_n19984_0[0]),.dinb(n20341),.dout(n20342),.clk(gclk));
	jand g20085(.dina(n20342),.dinb(n20224),.dout(n20343),.clk(gclk));
	jand g20086(.dina(n20343),.dinb(w_n5606_24[1]),.dout(n20344),.clk(gclk));
	jnot g20087(.din(w_n19992_0[0]),.dout(n20345),.clk(gclk));
	jor g20088(.dina(w_n20345_0[1]),.dinb(n20344),.dout(n20346),.clk(gclk));
	jand g20089(.dina(n20346),.dinb(n20223),.dout(n20347),.clk(gclk));
	jand g20090(.dina(n20347),.dinb(w_n5259_21[0]),.dout(n20348),.clk(gclk));
	jor g20091(.dina(w_n19999_0[0]),.dinb(n20348),.dout(n20349),.clk(gclk));
	jand g20092(.dina(n20349),.dinb(n20222),.dout(n20350),.clk(gclk));
	jand g20093(.dina(n20350),.dinb(w_n4902_25[0]),.dout(n20351),.clk(gclk));
	jnot g20094(.din(w_n20007_0[0]),.dout(n20352),.clk(gclk));
	jor g20095(.dina(w_n20352_0[1]),.dinb(n20351),.dout(n20353),.clk(gclk));
	jand g20096(.dina(n20353),.dinb(n20221),.dout(n20354),.clk(gclk));
	jand g20097(.dina(n20354),.dinb(w_n4582_22[0]),.dout(n20355),.clk(gclk));
	jor g20098(.dina(w_n20014_0[0]),.dinb(n20355),.dout(n20356),.clk(gclk));
	jand g20099(.dina(n20356),.dinb(n20220),.dout(n20357),.clk(gclk));
	jand g20100(.dina(n20357),.dinb(w_n4249_25[2]),.dout(n20358),.clk(gclk));
	jnot g20101(.din(w_n20022_0[0]),.dout(n20359),.clk(gclk));
	jor g20102(.dina(w_n20359_0[1]),.dinb(n20358),.dout(n20360),.clk(gclk));
	jand g20103(.dina(n20360),.dinb(n20219),.dout(n20361),.clk(gclk));
	jand g20104(.dina(n20361),.dinb(w_n3955_22[2]),.dout(n20362),.clk(gclk));
	jor g20105(.dina(w_n20029_0[0]),.dinb(n20362),.dout(n20363),.clk(gclk));
	jand g20106(.dina(n20363),.dinb(n20218),.dout(n20364),.clk(gclk));
	jand g20107(.dina(n20364),.dinb(w_n3642_26[0]),.dout(n20365),.clk(gclk));
	jor g20108(.dina(w_n20037_0[0]),.dinb(n20365),.dout(n20366),.clk(gclk));
	jand g20109(.dina(n20366),.dinb(n20217),.dout(n20367),.clk(gclk));
	jand g20110(.dina(n20367),.dinb(w_n3368_23[1]),.dout(n20368),.clk(gclk));
	jor g20111(.dina(w_n20045_0[0]),.dinb(n20368),.dout(n20369),.clk(gclk));
	jand g20112(.dina(n20369),.dinb(n20216),.dout(n20370),.clk(gclk));
	jand g20113(.dina(n20370),.dinb(w_n3089_26[2]),.dout(n20371),.clk(gclk));
	jnot g20114(.din(w_n20053_0[0]),.dout(n20372),.clk(gclk));
	jor g20115(.dina(w_n20372_0[1]),.dinb(n20371),.dout(n20373),.clk(gclk));
	jand g20116(.dina(n20373),.dinb(n20215),.dout(n20374),.clk(gclk));
	jand g20117(.dina(n20374),.dinb(w_n2833_24[1]),.dout(n20375),.clk(gclk));
	jor g20118(.dina(w_n20060_0[0]),.dinb(n20375),.dout(n20376),.clk(gclk));
	jand g20119(.dina(n20376),.dinb(n20214),.dout(n20377),.clk(gclk));
	jand g20120(.dina(n20377),.dinb(w_n2572_27[0]),.dout(n20378),.clk(gclk));
	jor g20121(.dina(w_n20068_0[0]),.dinb(n20378),.dout(n20379),.clk(gclk));
	jand g20122(.dina(n20379),.dinb(n20213),.dout(n20380),.clk(gclk));
	jand g20123(.dina(n20380),.dinb(w_n2345_25[0]),.dout(n20381),.clk(gclk));
	jor g20124(.dina(w_n20076_0[0]),.dinb(n20381),.dout(n20382),.clk(gclk));
	jand g20125(.dina(n20382),.dinb(n20212),.dout(n20383),.clk(gclk));
	jand g20126(.dina(n20383),.dinb(w_n2108_27[2]),.dout(n20384),.clk(gclk));
	jor g20127(.dina(w_n20084_0[0]),.dinb(n20384),.dout(n20385),.clk(gclk));
	jand g20128(.dina(n20385),.dinb(n20211),.dout(n20386),.clk(gclk));
	jand g20129(.dina(n20386),.dinb(w_n1912_26[0]),.dout(n20387),.clk(gclk));
	jor g20130(.dina(w_n20092_0[0]),.dinb(n20387),.dout(n20388),.clk(gclk));
	jand g20131(.dina(n20388),.dinb(n20210),.dout(n20389),.clk(gclk));
	jand g20132(.dina(n20389),.dinb(w_n1699_28[1]),.dout(n20390),.clk(gclk));
	jnot g20133(.din(w_n20100_0[0]),.dout(n20391),.clk(gclk));
	jor g20134(.dina(w_n20391_0[1]),.dinb(n20390),.dout(n20392),.clk(gclk));
	jand g20135(.dina(n20392),.dinb(n20209),.dout(n20393),.clk(gclk));
	jand g20136(.dina(n20393),.dinb(w_n1516_26[2]),.dout(n20394),.clk(gclk));
	jor g20137(.dina(w_n20107_0[0]),.dinb(n20394),.dout(n20395),.clk(gclk));
	jand g20138(.dina(n20395),.dinb(n20208),.dout(n20396),.clk(gclk));
	jand g20139(.dina(n20396),.dinb(w_n1332_28[1]),.dout(n20397),.clk(gclk));
	jnot g20140(.din(w_n20115_0[0]),.dout(n20398),.clk(gclk));
	jor g20141(.dina(w_n20398_0[1]),.dinb(n20397),.dout(n20399),.clk(gclk));
	jand g20142(.dina(n20399),.dinb(n20207),.dout(n20400),.clk(gclk));
	jand g20143(.dina(n20400),.dinb(w_n1173_27[1]),.dout(n20401),.clk(gclk));
	jor g20144(.dina(w_n20122_0[0]),.dinb(n20401),.dout(n20402),.clk(gclk));
	jand g20145(.dina(n20402),.dinb(n20206),.dout(n20403),.clk(gclk));
	jand g20146(.dina(n20403),.dinb(w_n1008_29[1]),.dout(n20404),.clk(gclk));
	jor g20147(.dina(w_n20130_0[0]),.dinb(n20404),.dout(n20405),.clk(gclk));
	jand g20148(.dina(n20405),.dinb(n20205),.dout(n20406),.clk(gclk));
	jand g20149(.dina(n20406),.dinb(w_n884_28[1]),.dout(n20407),.clk(gclk));
	jnot g20150(.din(w_n20138_0[0]),.dout(n20408),.clk(gclk));
	jor g20151(.dina(w_n20408_0[1]),.dinb(n20407),.dout(n20409),.clk(gclk));
	jand g20152(.dina(n20409),.dinb(n20204),.dout(n20410),.clk(gclk));
	jand g20153(.dina(n20410),.dinb(w_n743_29[1]),.dout(n20411),.clk(gclk));
	jor g20154(.dina(n20411),.dinb(w_n20203_0[1]),.dout(n20412),.clk(gclk));
	jand g20155(.dina(n20412),.dinb(n20202),.dout(n20413),.clk(gclk));
	jand g20156(.dina(n20413),.dinb(w_n635_29[1]),.dout(n20414),.clk(gclk));
	jor g20157(.dina(w_n20152_0[0]),.dinb(n20414),.dout(n20415),.clk(gclk));
	jand g20158(.dina(n20415),.dinb(n20201),.dout(n20416),.clk(gclk));
	jand g20159(.dina(n20416),.dinb(w_n515_30[1]),.dout(n20417),.clk(gclk));
	jnot g20160(.din(w_n20160_0[0]),.dout(n20418),.clk(gclk));
	jor g20161(.dina(w_n20418_0[1]),.dinb(n20417),.dout(n20419),.clk(gclk));
	jand g20162(.dina(n20419),.dinb(n20200),.dout(n20420),.clk(gclk));
	jand g20163(.dina(n20420),.dinb(w_n443_30[1]),.dout(n20421),.clk(gclk));
	jor g20164(.dina(w_n20167_0[0]),.dinb(n20421),.dout(n20422),.clk(gclk));
	jand g20165(.dina(n20422),.dinb(n20199),.dout(n20423),.clk(gclk));
	jand g20166(.dina(n20423),.dinb(w_n352_30[2]),.dout(n20424),.clk(gclk));
	jor g20167(.dina(w_n20175_0[0]),.dinb(n20424),.dout(n20425),.clk(gclk));
	jand g20168(.dina(n20425),.dinb(n20198),.dout(n20426),.clk(gclk));
	jand g20169(.dina(n20426),.dinb(w_n294_31[0]),.dout(n20427),.clk(gclk));
	jnot g20170(.din(w_n20183_0[0]),.dout(n20428),.clk(gclk));
	jor g20171(.dina(w_n20428_0[1]),.dinb(n20427),.dout(n20429),.clk(gclk));
	jand g20172(.dina(n20429),.dinb(n20197),.dout(n20430),.clk(gclk));
	jand g20173(.dina(n20430),.dinb(w_n239_31[1]),.dout(n20431),.clk(gclk));
	jor g20174(.dina(w_n20190_0[0]),.dinb(n20431),.dout(n20432),.clk(gclk));
	jand g20175(.dina(n20432),.dinb(n20196),.dout(n20433),.clk(gclk));
	jand g20176(.dina(n20433),.dinb(w_n221_31[1]),.dout(n20434),.clk(gclk));
	jxor g20177(.dina(w_n19490_0[0]),.dinb(w_n239_31[0]),.dout(n20435),.clk(gclk));
	jand g20178(.dina(n20435),.dinb(w_asqrt8_14[0]),.dout(n20436),.clk(gclk));
	jxor g20179(.dina(n20436),.dinb(w_n19495_0[0]),.dout(n20437),.clk(gclk));
	jor g20180(.dina(w_n20437_0[2]),.dinb(n20434),.dout(n20438),.clk(gclk));
	jand g20181(.dina(n20438),.dinb(n20195),.dout(n20439),.clk(gclk));
	jor g20182(.dina(w_n20439_0[2]),.dinb(w_n19523_0[2]),.dout(n20440),.clk(gclk));
	jand g20183(.dina(w_asqrt8_13[2]),.dinb(w_n19782_0[0]),.dout(n20441),.clk(gclk));
	jor g20184(.dina(n20441),.dinb(w_n19511_0[0]),.dout(n20442),.clk(gclk));
	jor g20185(.dina(w_n20442_0[1]),.dinb(w_n20440_0[1]),.dout(n20443),.clk(gclk));
	jand g20186(.dina(n20443),.dinb(w_n218_13[1]),.dout(n20444),.clk(gclk));
	jand g20187(.dina(w_n19791_9[2]),.dinb(w_n19100_0[0]),.dout(n20445),.clk(gclk));
	jand g20188(.dina(w_n20439_0[1]),.dinb(w_n19523_0[1]),.dout(n20446),.clk(gclk));
	jor g20189(.dina(w_n20446_0[2]),.dinb(w_n20445_0[1]),.dout(n20447),.clk(gclk));
	jand g20190(.dina(w_n19791_9[1]),.dinb(w_n19505_0[0]),.dout(n20448),.clk(gclk));
	jnot g20191(.din(n20448),.dout(n20449),.clk(gclk));
	jand g20192(.dina(w_n19786_0[0]),.dinb(w_asqrt63_22[2]),.dout(n20450),.clk(gclk));
	jand g20193(.dina(n20450),.dinb(w_n19506_0[0]),.dout(n20451),.clk(gclk));
	jand g20194(.dina(w_n20451_0[1]),.dinb(n20449),.dout(n20452),.clk(gclk));
	jor g20195(.dina(w_n20452_0[1]),.dinb(n20447),.dout(n20453),.clk(gclk));
	jor g20196(.dina(n20453),.dinb(w_n20444_0[1]),.dout(asqrt_fa_8),.clk(gclk));
	jor g20197(.dina(w_n20193_0[1]),.dinb(w_asqrt62_18[0]),.dout(n20455),.clk(gclk));
	jnot g20198(.din(w_n20437_0[1]),.dout(n20456),.clk(gclk));
	jand g20199(.dina(n20456),.dinb(n20455),.dout(n20457),.clk(gclk));
	jor g20200(.dina(n20457),.dinb(w_n20194_0[0]),.dout(n20458),.clk(gclk));
	jand g20201(.dina(w_n20458_0[1]),.dinb(w_n19522_0[1]),.dout(n20459),.clk(gclk));
	jnot g20202(.din(w_n20442_0[0]),.dout(n20460),.clk(gclk));
	jand g20203(.dina(n20460),.dinb(w_n20459_0[1]),.dout(n20461),.clk(gclk));
	jor g20204(.dina(n20461),.dinb(w_asqrt63_22[1]),.dout(n20462),.clk(gclk));
	jnot g20205(.din(w_n20445_0[0]),.dout(n20463),.clk(gclk));
	jor g20206(.dina(w_n20458_0[0]),.dinb(w_n19522_0[0]),.dout(n20464),.clk(gclk));
	jand g20207(.dina(w_n20464_0[1]),.dinb(n20463),.dout(n20465),.clk(gclk));
	jnot g20208(.din(w_n20452_0[0]),.dout(n20466),.clk(gclk));
	jand g20209(.dina(n20466),.dinb(n20465),.dout(n20467),.clk(gclk));
	jand g20210(.dina(n20467),.dinb(n20462),.dout(n20468),.clk(gclk));
	jxor g20211(.dina(w_n20193_0[0]),.dinb(w_n221_31[0]),.dout(n20469),.clk(gclk));
	jor g20212(.dina(n20469),.dinb(w_n20468_35[2]),.dout(n20470),.clk(gclk));
	jxor g20213(.dina(n20470),.dinb(w_n20437_0[0]),.dout(n20471),.clk(gclk));
	jnot g20214(.din(w_n20471_0[2]),.dout(n20472),.clk(gclk));
	jnot g20215(.din(w_a12_0[2]),.dout(n20473),.clk(gclk));
	jnot g20216(.din(w_a13_0[1]),.dout(n20474),.clk(gclk));
	jand g20217(.dina(w_n20474_0[1]),.dinb(w_n20473_1[2]),.dout(n20475),.clk(gclk));
	jand g20218(.dina(w_n20475_0[2]),.dinb(w_n19524_1[0]),.dout(n20476),.clk(gclk));
	jnot g20219(.din(w_n20476_0[1]),.dout(n20477),.clk(gclk));
	jor g20220(.dina(w_n20468_35[1]),.dinb(w_n19524_0[2]),.dout(n20478),.clk(gclk));
	jand g20221(.dina(n20478),.dinb(n20477),.dout(n20479),.clk(gclk));
	jor g20222(.dina(w_n20479_0[2]),.dinb(w_n19791_9[0]),.dout(n20480),.clk(gclk));
	jand g20223(.dina(w_n20479_0[1]),.dinb(w_n19791_8[2]),.dout(n20481),.clk(gclk));
	jor g20224(.dina(w_n20468_35[0]),.dinb(w_a14_1[0]),.dout(n20482),.clk(gclk));
	jand g20225(.dina(n20482),.dinb(w_a15_0[0]),.dout(n20483),.clk(gclk));
	jand g20226(.dina(w_asqrt7_6),.dinb(w_n19526_0[1]),.dout(n20484),.clk(gclk));
	jor g20227(.dina(n20484),.dinb(n20483),.dout(n20485),.clk(gclk));
	jor g20228(.dina(n20485),.dinb(n20481),.dout(n20486),.clk(gclk));
	jand g20229(.dina(n20486),.dinb(w_n20480_0[1]),.dout(n20487),.clk(gclk));
	jor g20230(.dina(w_n20487_0[2]),.dinb(w_n19096_17[2]),.dout(n20488),.clk(gclk));
	jand g20231(.dina(w_n20487_0[1]),.dinb(w_n19096_17[1]),.dout(n20489),.clk(gclk));
	jnot g20232(.din(w_n19526_0[0]),.dout(n20490),.clk(gclk));
	jor g20233(.dina(w_n20468_34[2]),.dinb(n20490),.dout(n20491),.clk(gclk));
	jor g20234(.dina(w_n20451_0[0]),.dinb(w_n20446_0[1]),.dout(n20492),.clk(gclk));
	jor g20235(.dina(n20492),.dinb(w_n20444_0[0]),.dout(n20493),.clk(gclk));
	jor g20236(.dina(n20493),.dinb(w_n19791_8[1]),.dout(n20494),.clk(gclk));
	jand g20237(.dina(n20494),.dinb(w_n20491_0[1]),.dout(n20495),.clk(gclk));
	jxor g20238(.dina(n20495),.dinb(w_n19101_0[1]),.dout(n20496),.clk(gclk));
	jor g20239(.dina(w_n20496_0[2]),.dinb(n20489),.dout(n20497),.clk(gclk));
	jand g20240(.dina(n20497),.dinb(w_n20488_0[1]),.dout(n20498),.clk(gclk));
	jor g20241(.dina(w_n20498_0[2]),.dinb(w_n18442_9[2]),.dout(n20499),.clk(gclk));
	jand g20242(.dina(w_n20498_0[1]),.dinb(w_n18442_9[1]),.dout(n20500),.clk(gclk));
	jxor g20243(.dina(w_n19529_0[0]),.dinb(w_n19096_17[0]),.dout(n20501),.clk(gclk));
	jor g20244(.dina(n20501),.dinb(w_n20468_34[1]),.dout(n20502),.clk(gclk));
	jxor g20245(.dina(n20502),.dinb(w_n20256_0[0]),.dout(n20503),.clk(gclk));
	jnot g20246(.din(w_n20503_0[2]),.dout(n20504),.clk(gclk));
	jor g20247(.dina(n20504),.dinb(n20500),.dout(n20505),.clk(gclk));
	jand g20248(.dina(n20505),.dinb(w_n20499_0[1]),.dout(n20506),.clk(gclk));
	jor g20249(.dina(w_n20506_0[2]),.dinb(w_n17769_18[1]),.dout(n20507),.clk(gclk));
	jand g20250(.dina(w_n20506_0[1]),.dinb(w_n17769_18[0]),.dout(n20508),.clk(gclk));
	jxor g20251(.dina(w_n19795_0[0]),.dinb(w_n18442_9[0]),.dout(n20509),.clk(gclk));
	jor g20252(.dina(n20509),.dinb(w_n20468_34[0]),.dout(n20510),.clk(gclk));
	jxor g20253(.dina(n20510),.dinb(w_n19803_0[0]),.dout(n20511),.clk(gclk));
	jor g20254(.dina(w_n20511_0[2]),.dinb(n20508),.dout(n20512),.clk(gclk));
	jand g20255(.dina(n20512),.dinb(w_n20507_0[1]),.dout(n20513),.clk(gclk));
	jor g20256(.dina(w_n20513_0[2]),.dinb(w_n17134_10[2]),.dout(n20514),.clk(gclk));
	jand g20257(.dina(w_n20513_0[1]),.dinb(w_n17134_10[1]),.dout(n20515),.clk(gclk));
	jxor g20258(.dina(w_n19805_0[0]),.dinb(w_n17769_17[2]),.dout(n20516),.clk(gclk));
	jor g20259(.dina(n20516),.dinb(w_n20468_33[2]),.dout(n20517),.clk(gclk));
	jxor g20260(.dina(n20517),.dinb(w_n19811_0[0]),.dout(n20518),.clk(gclk));
	jor g20261(.dina(w_n20518_0[2]),.dinb(n20515),.dout(n20519),.clk(gclk));
	jand g20262(.dina(n20519),.dinb(w_n20514_0[1]),.dout(n20520),.clk(gclk));
	jor g20263(.dina(w_n20520_0[2]),.dinb(w_n16489_18[2]),.dout(n20521),.clk(gclk));
	jand g20264(.dina(w_n20520_0[1]),.dinb(w_n16489_18[1]),.dout(n20522),.clk(gclk));
	jxor g20265(.dina(w_n19813_0[0]),.dinb(w_n17134_10[0]),.dout(n20523),.clk(gclk));
	jor g20266(.dina(n20523),.dinb(w_n20468_33[1]),.dout(n20524),.clk(gclk));
	jxor g20267(.dina(n20524),.dinb(w_n19819_0[0]),.dout(n20525),.clk(gclk));
	jor g20268(.dina(w_n20525_0[2]),.dinb(n20522),.dout(n20526),.clk(gclk));
	jand g20269(.dina(n20526),.dinb(w_n20521_0[1]),.dout(n20527),.clk(gclk));
	jor g20270(.dina(w_n20527_0[2]),.dinb(w_n15878_11[2]),.dout(n20528),.clk(gclk));
	jand g20271(.dina(w_n20527_0[1]),.dinb(w_n15878_11[1]),.dout(n20529),.clk(gclk));
	jxor g20272(.dina(w_n19821_0[0]),.dinb(w_n16489_18[0]),.dout(n20530),.clk(gclk));
	jor g20273(.dina(n20530),.dinb(w_n20468_33[0]),.dout(n20531),.clk(gclk));
	jxor g20274(.dina(n20531),.dinb(w_n20269_0[0]),.dout(n20532),.clk(gclk));
	jnot g20275(.din(w_n20532_0[2]),.dout(n20533),.clk(gclk));
	jor g20276(.dina(n20533),.dinb(n20529),.dout(n20534),.clk(gclk));
	jand g20277(.dina(n20534),.dinb(w_n20528_0[1]),.dout(n20535),.clk(gclk));
	jor g20278(.dina(w_n20535_0[2]),.dinb(w_n15260_19[1]),.dout(n20536),.clk(gclk));
	jand g20279(.dina(w_n20535_0[1]),.dinb(w_n15260_19[0]),.dout(n20537),.clk(gclk));
	jxor g20280(.dina(w_n19828_0[0]),.dinb(w_n15878_11[0]),.dout(n20538),.clk(gclk));
	jor g20281(.dina(n20538),.dinb(w_n20468_32[2]),.dout(n20539),.clk(gclk));
	jxor g20282(.dina(n20539),.dinb(w_n19834_0[0]),.dout(n20540),.clk(gclk));
	jor g20283(.dina(w_n20540_0[2]),.dinb(n20537),.dout(n20541),.clk(gclk));
	jand g20284(.dina(n20541),.dinb(w_n20536_0[1]),.dout(n20542),.clk(gclk));
	jor g20285(.dina(w_n20542_0[2]),.dinb(w_n14674_12[1]),.dout(n20543),.clk(gclk));
	jand g20286(.dina(w_n20542_0[1]),.dinb(w_n14674_12[0]),.dout(n20544),.clk(gclk));
	jxor g20287(.dina(w_n19836_0[0]),.dinb(w_n15260_18[2]),.dout(n20545),.clk(gclk));
	jor g20288(.dina(n20545),.dinb(w_n20468_32[1]),.dout(n20546),.clk(gclk));
	jxor g20289(.dina(n20546),.dinb(w_n20276_0[0]),.dout(n20547),.clk(gclk));
	jnot g20290(.din(w_n20547_0[1]),.dout(n20548),.clk(gclk));
	jor g20291(.dina(w_n20548_0[1]),.dinb(n20544),.dout(n20549),.clk(gclk));
	jand g20292(.dina(n20549),.dinb(w_n20543_0[1]),.dout(n20550),.clk(gclk));
	jor g20293(.dina(w_n20550_0[2]),.dinb(w_n14078_19[2]),.dout(n20551),.clk(gclk));
	jand g20294(.dina(w_n20550_0[1]),.dinb(w_n14078_19[1]),.dout(n20552),.clk(gclk));
	jxor g20295(.dina(w_n19843_0[0]),.dinb(w_n14674_11[2]),.dout(n20553),.clk(gclk));
	jor g20296(.dina(n20553),.dinb(w_n20468_32[0]),.dout(n20554),.clk(gclk));
	jxor g20297(.dina(n20554),.dinb(w_n19849_0[0]),.dout(n20555),.clk(gclk));
	jor g20298(.dina(w_n20555_0[2]),.dinb(n20552),.dout(n20556),.clk(gclk));
	jand g20299(.dina(n20556),.dinb(w_n20551_0[1]),.dout(n20557),.clk(gclk));
	jor g20300(.dina(w_n20557_0[2]),.dinb(w_n13515_13[1]),.dout(n20558),.clk(gclk));
	jand g20301(.dina(w_n20557_0[1]),.dinb(w_n13515_13[0]),.dout(n20559),.clk(gclk));
	jxor g20302(.dina(w_n19851_0[0]),.dinb(w_n14078_19[0]),.dout(n20560),.clk(gclk));
	jor g20303(.dina(n20560),.dinb(w_n20468_31[2]),.dout(n20561),.clk(gclk));
	jxor g20304(.dina(n20561),.dinb(w_n20283_0[0]),.dout(n20562),.clk(gclk));
	jnot g20305(.din(w_n20562_0[2]),.dout(n20563),.clk(gclk));
	jor g20306(.dina(n20563),.dinb(n20559),.dout(n20564),.clk(gclk));
	jand g20307(.dina(n20564),.dinb(w_n20558_0[1]),.dout(n20565),.clk(gclk));
	jor g20308(.dina(w_n20565_0[2]),.dinb(w_n12947_20[1]),.dout(n20566),.clk(gclk));
	jand g20309(.dina(w_n20565_0[1]),.dinb(w_n12947_20[0]),.dout(n20567),.clk(gclk));
	jxor g20310(.dina(w_n19858_0[0]),.dinb(w_n13515_12[2]),.dout(n20568),.clk(gclk));
	jor g20311(.dina(n20568),.dinb(w_n20468_31[1]),.dout(n20569),.clk(gclk));
	jxor g20312(.dina(n20569),.dinb(w_n19864_0[0]),.dout(n20570),.clk(gclk));
	jor g20313(.dina(w_n20570_0[2]),.dinb(n20567),.dout(n20571),.clk(gclk));
	jand g20314(.dina(n20571),.dinb(w_n20566_0[1]),.dout(n20572),.clk(gclk));
	jor g20315(.dina(w_n20572_0[2]),.dinb(w_n12410_14[0]),.dout(n20573),.clk(gclk));
	jand g20316(.dina(w_n20572_0[1]),.dinb(w_n12410_13[2]),.dout(n20574),.clk(gclk));
	jxor g20317(.dina(w_n19866_0[0]),.dinb(w_n12947_19[2]),.dout(n20575),.clk(gclk));
	jor g20318(.dina(n20575),.dinb(w_n20468_31[0]),.dout(n20576),.clk(gclk));
	jxor g20319(.dina(n20576),.dinb(w_n20290_0[0]),.dout(n20577),.clk(gclk));
	jnot g20320(.din(w_n20577_0[2]),.dout(n20578),.clk(gclk));
	jor g20321(.dina(n20578),.dinb(n20574),.dout(n20579),.clk(gclk));
	jand g20322(.dina(n20579),.dinb(w_n20573_0[1]),.dout(n20580),.clk(gclk));
	jor g20323(.dina(w_n20580_0[2]),.dinb(w_n11858_20[2]),.dout(n20581),.clk(gclk));
	jand g20324(.dina(w_n20580_0[1]),.dinb(w_n11858_20[1]),.dout(n20582),.clk(gclk));
	jxor g20325(.dina(w_n19873_0[0]),.dinb(w_n12410_13[1]),.dout(n20583),.clk(gclk));
	jor g20326(.dina(n20583),.dinb(w_n20468_30[2]),.dout(n20584),.clk(gclk));
	jxor g20327(.dina(n20584),.dinb(w_n19879_0[0]),.dout(n20585),.clk(gclk));
	jor g20328(.dina(w_n20585_0[2]),.dinb(n20582),.dout(n20586),.clk(gclk));
	jand g20329(.dina(n20586),.dinb(w_n20581_0[1]),.dout(n20587),.clk(gclk));
	jor g20330(.dina(w_n20587_0[2]),.dinb(w_n11347_14[2]),.dout(n20588),.clk(gclk));
	jand g20331(.dina(w_n20587_0[1]),.dinb(w_n11347_14[1]),.dout(n20589),.clk(gclk));
	jxor g20332(.dina(w_n19881_0[0]),.dinb(w_n11858_20[0]),.dout(n20590),.clk(gclk));
	jor g20333(.dina(n20590),.dinb(w_n20468_30[1]),.dout(n20591),.clk(gclk));
	jxor g20334(.dina(n20591),.dinb(w_n20297_0[0]),.dout(n20592),.clk(gclk));
	jnot g20335(.din(w_n20592_0[2]),.dout(n20593),.clk(gclk));
	jor g20336(.dina(n20593),.dinb(n20589),.dout(n20594),.clk(gclk));
	jand g20337(.dina(n20594),.dinb(w_n20588_0[1]),.dout(n20595),.clk(gclk));
	jor g20338(.dina(w_n20595_0[2]),.dinb(w_n10824_21[1]),.dout(n20596),.clk(gclk));
	jand g20339(.dina(w_n20595_0[1]),.dinb(w_n10824_21[0]),.dout(n20597),.clk(gclk));
	jxor g20340(.dina(w_n19888_0[0]),.dinb(w_n11347_14[0]),.dout(n20598),.clk(gclk));
	jor g20341(.dina(n20598),.dinb(w_n20468_30[0]),.dout(n20599),.clk(gclk));
	jxor g20342(.dina(n20599),.dinb(w_n19894_0[0]),.dout(n20600),.clk(gclk));
	jor g20343(.dina(w_n20600_0[2]),.dinb(n20597),.dout(n20601),.clk(gclk));
	jand g20344(.dina(n20601),.dinb(w_n20596_0[1]),.dout(n20602),.clk(gclk));
	jor g20345(.dina(w_n20602_0[2]),.dinb(w_n10328_15[2]),.dout(n20603),.clk(gclk));
	jand g20346(.dina(w_n20602_0[1]),.dinb(w_n10328_15[1]),.dout(n20604),.clk(gclk));
	jxor g20347(.dina(w_n19896_0[0]),.dinb(w_n10824_20[2]),.dout(n20605),.clk(gclk));
	jor g20348(.dina(n20605),.dinb(w_n20468_29[2]),.dout(n20606),.clk(gclk));
	jxor g20349(.dina(n20606),.dinb(w_n19902_0[0]),.dout(n20607),.clk(gclk));
	jor g20350(.dina(w_n20607_0[2]),.dinb(n20604),.dout(n20608),.clk(gclk));
	jand g20351(.dina(n20608),.dinb(w_n20603_0[1]),.dout(n20609),.clk(gclk));
	jor g20352(.dina(w_n20609_0[2]),.dinb(w_n9832_22[0]),.dout(n20610),.clk(gclk));
	jand g20353(.dina(w_n20609_0[1]),.dinb(w_n9832_21[2]),.dout(n20611),.clk(gclk));
	jxor g20354(.dina(w_n19904_0[0]),.dinb(w_n10328_15[0]),.dout(n20612),.clk(gclk));
	jor g20355(.dina(n20612),.dinb(w_n20468_29[1]),.dout(n20613),.clk(gclk));
	jxor g20356(.dina(n20613),.dinb(w_n20307_0[0]),.dout(n20614),.clk(gclk));
	jnot g20357(.din(w_n20614_0[2]),.dout(n20615),.clk(gclk));
	jor g20358(.dina(n20615),.dinb(n20611),.dout(n20616),.clk(gclk));
	jand g20359(.dina(n20616),.dinb(w_n20610_0[1]),.dout(n20617),.clk(gclk));
	jor g20360(.dina(w_n20617_0[2]),.dinb(w_n9369_16[2]),.dout(n20618),.clk(gclk));
	jand g20361(.dina(w_n20617_0[1]),.dinb(w_n9369_16[1]),.dout(n20619),.clk(gclk));
	jxor g20362(.dina(w_n19911_0[0]),.dinb(w_n9832_21[1]),.dout(n20620),.clk(gclk));
	jor g20363(.dina(n20620),.dinb(w_n20468_29[0]),.dout(n20621),.clk(gclk));
	jxor g20364(.dina(n20621),.dinb(w_n20311_0[0]),.dout(n20622),.clk(gclk));
	jnot g20365(.din(w_n20622_0[2]),.dout(n20623),.clk(gclk));
	jor g20366(.dina(n20623),.dinb(n20619),.dout(n20624),.clk(gclk));
	jand g20367(.dina(n20624),.dinb(w_n20618_0[1]),.dout(n20625),.clk(gclk));
	jor g20368(.dina(w_n20625_0[2]),.dinb(w_n8890_22[1]),.dout(n20626),.clk(gclk));
	jand g20369(.dina(w_n20625_0[1]),.dinb(w_n8890_22[0]),.dout(n20627),.clk(gclk));
	jxor g20370(.dina(w_n19918_0[0]),.dinb(w_n9369_16[0]),.dout(n20628),.clk(gclk));
	jor g20371(.dina(n20628),.dinb(w_n20468_28[2]),.dout(n20629),.clk(gclk));
	jxor g20372(.dina(n20629),.dinb(w_n19924_0[0]),.dout(n20630),.clk(gclk));
	jor g20373(.dina(w_n20630_0[2]),.dinb(n20627),.dout(n20631),.clk(gclk));
	jand g20374(.dina(n20631),.dinb(w_n20626_0[1]),.dout(n20632),.clk(gclk));
	jor g20375(.dina(w_n20632_0[2]),.dinb(w_n8449_17[1]),.dout(n20633),.clk(gclk));
	jand g20376(.dina(w_n20632_0[1]),.dinb(w_n8449_17[0]),.dout(n20634),.clk(gclk));
	jxor g20377(.dina(w_n19926_0[0]),.dinb(w_n8890_21[2]),.dout(n20635),.clk(gclk));
	jor g20378(.dina(n20635),.dinb(w_n20468_28[1]),.dout(n20636),.clk(gclk));
	jxor g20379(.dina(n20636),.dinb(w_n20318_0[0]),.dout(n20637),.clk(gclk));
	jnot g20380(.din(w_n20637_0[2]),.dout(n20638),.clk(gclk));
	jor g20381(.dina(n20638),.dinb(n20634),.dout(n20639),.clk(gclk));
	jand g20382(.dina(n20639),.dinb(w_n20633_0[1]),.dout(n20640),.clk(gclk));
	jor g20383(.dina(w_n20640_0[2]),.dinb(w_n8003_23[0]),.dout(n20641),.clk(gclk));
	jand g20384(.dina(w_n20640_0[1]),.dinb(w_n8003_22[2]),.dout(n20642),.clk(gclk));
	jxor g20385(.dina(w_n19933_0[0]),.dinb(w_n8449_16[2]),.dout(n20643),.clk(gclk));
	jor g20386(.dina(n20643),.dinb(w_n20468_28[0]),.dout(n20644),.clk(gclk));
	jxor g20387(.dina(n20644),.dinb(w_n19939_0[0]),.dout(n20645),.clk(gclk));
	jor g20388(.dina(w_n20645_0[2]),.dinb(n20642),.dout(n20646),.clk(gclk));
	jand g20389(.dina(n20646),.dinb(w_n20641_0[1]),.dout(n20647),.clk(gclk));
	jor g20390(.dina(w_n20647_0[2]),.dinb(w_n7581_18[1]),.dout(n20648),.clk(gclk));
	jand g20391(.dina(w_n20647_0[1]),.dinb(w_n7581_18[0]),.dout(n20649),.clk(gclk));
	jxor g20392(.dina(w_n19941_0[0]),.dinb(w_n8003_22[1]),.dout(n20650),.clk(gclk));
	jor g20393(.dina(n20650),.dinb(w_n20468_27[2]),.dout(n20651),.clk(gclk));
	jxor g20394(.dina(n20651),.dinb(w_n20325_0[0]),.dout(n20652),.clk(gclk));
	jnot g20395(.din(w_n20652_0[2]),.dout(n20653),.clk(gclk));
	jor g20396(.dina(n20653),.dinb(n20649),.dout(n20654),.clk(gclk));
	jand g20397(.dina(n20654),.dinb(w_n20648_0[1]),.dout(n20655),.clk(gclk));
	jor g20398(.dina(w_n20655_0[2]),.dinb(w_n7154_23[1]),.dout(n20656),.clk(gclk));
	jand g20399(.dina(w_n20655_0[1]),.dinb(w_n7154_23[0]),.dout(n20657),.clk(gclk));
	jxor g20400(.dina(w_n19948_0[0]),.dinb(w_n7581_17[2]),.dout(n20658),.clk(gclk));
	jor g20401(.dina(n20658),.dinb(w_n20468_27[1]),.dout(n20659),.clk(gclk));
	jxor g20402(.dina(n20659),.dinb(w_n19954_0[0]),.dout(n20660),.clk(gclk));
	jor g20403(.dina(w_n20660_0[2]),.dinb(n20657),.dout(n20661),.clk(gclk));
	jand g20404(.dina(n20661),.dinb(w_n20656_0[1]),.dout(n20662),.clk(gclk));
	jor g20405(.dina(w_n20662_0[2]),.dinb(w_n6758_19[0]),.dout(n20663),.clk(gclk));
	jand g20406(.dina(w_n20662_0[1]),.dinb(w_n6758_18[2]),.dout(n20664),.clk(gclk));
	jxor g20407(.dina(w_n19956_0[0]),.dinb(w_n7154_22[2]),.dout(n20665),.clk(gclk));
	jor g20408(.dina(n20665),.dinb(w_n20468_27[0]),.dout(n20666),.clk(gclk));
	jxor g20409(.dina(n20666),.dinb(w_n19962_0[0]),.dout(n20667),.clk(gclk));
	jor g20410(.dina(w_n20667_0[2]),.dinb(n20664),.dout(n20668),.clk(gclk));
	jand g20411(.dina(n20668),.dinb(w_n20663_0[1]),.dout(n20669),.clk(gclk));
	jor g20412(.dina(w_n20669_0[2]),.dinb(w_n6357_23[2]),.dout(n20670),.clk(gclk));
	jand g20413(.dina(w_n20669_0[1]),.dinb(w_n6357_23[1]),.dout(n20671),.clk(gclk));
	jxor g20414(.dina(w_n19964_0[0]),.dinb(w_n6758_18[1]),.dout(n20672),.clk(gclk));
	jor g20415(.dina(n20672),.dinb(w_n20468_26[2]),.dout(n20673),.clk(gclk));
	jxor g20416(.dina(n20673),.dinb(w_n19970_0[0]),.dout(n20674),.clk(gclk));
	jor g20417(.dina(w_n20674_0[2]),.dinb(n20671),.dout(n20675),.clk(gclk));
	jand g20418(.dina(n20675),.dinb(w_n20670_0[1]),.dout(n20676),.clk(gclk));
	jor g20419(.dina(w_n20676_0[2]),.dinb(w_n5989_19[2]),.dout(n20677),.clk(gclk));
	jand g20420(.dina(w_n20676_0[1]),.dinb(w_n5989_19[1]),.dout(n20678),.clk(gclk));
	jxor g20421(.dina(w_n19972_0[0]),.dinb(w_n6357_23[0]),.dout(n20679),.clk(gclk));
	jor g20422(.dina(n20679),.dinb(w_n20468_26[1]),.dout(n20680),.clk(gclk));
	jxor g20423(.dina(n20680),.dinb(w_n20338_0[0]),.dout(n20681),.clk(gclk));
	jnot g20424(.din(w_n20681_0[2]),.dout(n20682),.clk(gclk));
	jor g20425(.dina(n20682),.dinb(n20678),.dout(n20683),.clk(gclk));
	jand g20426(.dina(n20683),.dinb(w_n20677_0[1]),.dout(n20684),.clk(gclk));
	jor g20427(.dina(w_n20684_0[2]),.dinb(w_n5606_24[0]),.dout(n20685),.clk(gclk));
	jand g20428(.dina(w_n20684_0[1]),.dinb(w_n5606_23[2]),.dout(n20686),.clk(gclk));
	jxor g20429(.dina(w_n19979_0[0]),.dinb(w_n5989_19[0]),.dout(n20687),.clk(gclk));
	jor g20430(.dina(n20687),.dinb(w_n20468_26[0]),.dout(n20688),.clk(gclk));
	jxor g20431(.dina(n20688),.dinb(w_n19985_0[0]),.dout(n20689),.clk(gclk));
	jor g20432(.dina(w_n20689_0[2]),.dinb(n20686),.dout(n20690),.clk(gclk));
	jand g20433(.dina(n20690),.dinb(w_n20685_0[1]),.dout(n20691),.clk(gclk));
	jor g20434(.dina(w_n20691_0[2]),.dinb(w_n5259_20[2]),.dout(n20692),.clk(gclk));
	jand g20435(.dina(w_n20691_0[1]),.dinb(w_n5259_20[1]),.dout(n20693),.clk(gclk));
	jxor g20436(.dina(w_n19987_0[0]),.dinb(w_n5606_23[1]),.dout(n20694),.clk(gclk));
	jor g20437(.dina(n20694),.dinb(w_n20468_25[2]),.dout(n20695),.clk(gclk));
	jxor g20438(.dina(n20695),.dinb(w_n20345_0[0]),.dout(n20696),.clk(gclk));
	jnot g20439(.din(w_n20696_0[2]),.dout(n20697),.clk(gclk));
	jor g20440(.dina(n20697),.dinb(n20693),.dout(n20698),.clk(gclk));
	jand g20441(.dina(n20698),.dinb(w_n20692_0[1]),.dout(n20699),.clk(gclk));
	jor g20442(.dina(w_n20699_0[2]),.dinb(w_n4902_24[2]),.dout(n20700),.clk(gclk));
	jand g20443(.dina(w_n20699_0[1]),.dinb(w_n4902_24[1]),.dout(n20701),.clk(gclk));
	jxor g20444(.dina(w_n19994_0[0]),.dinb(w_n5259_20[0]),.dout(n20702),.clk(gclk));
	jor g20445(.dina(n20702),.dinb(w_n20468_25[1]),.dout(n20703),.clk(gclk));
	jxor g20446(.dina(n20703),.dinb(w_n20000_0[0]),.dout(n20704),.clk(gclk));
	jor g20447(.dina(w_n20704_0[2]),.dinb(n20701),.dout(n20705),.clk(gclk));
	jand g20448(.dina(n20705),.dinb(w_n20700_0[1]),.dout(n20706),.clk(gclk));
	jor g20449(.dina(w_n20706_0[2]),.dinb(w_n4582_21[2]),.dout(n20707),.clk(gclk));
	jand g20450(.dina(w_n20706_0[1]),.dinb(w_n4582_21[1]),.dout(n20708),.clk(gclk));
	jxor g20451(.dina(w_n20002_0[0]),.dinb(w_n4902_24[0]),.dout(n20709),.clk(gclk));
	jor g20452(.dina(n20709),.dinb(w_n20468_25[0]),.dout(n20710),.clk(gclk));
	jxor g20453(.dina(n20710),.dinb(w_n20352_0[0]),.dout(n20711),.clk(gclk));
	jnot g20454(.din(w_n20711_0[2]),.dout(n20712),.clk(gclk));
	jor g20455(.dina(n20712),.dinb(n20708),.dout(n20713),.clk(gclk));
	jand g20456(.dina(n20713),.dinb(w_n20707_0[1]),.dout(n20714),.clk(gclk));
	jor g20457(.dina(w_n20714_0[2]),.dinb(w_n4249_25[1]),.dout(n20715),.clk(gclk));
	jand g20458(.dina(w_n20714_0[1]),.dinb(w_n4249_25[0]),.dout(n20716),.clk(gclk));
	jxor g20459(.dina(w_n20009_0[0]),.dinb(w_n4582_21[0]),.dout(n20717),.clk(gclk));
	jor g20460(.dina(n20717),.dinb(w_n20468_24[2]),.dout(n20718),.clk(gclk));
	jxor g20461(.dina(n20718),.dinb(w_n20015_0[0]),.dout(n20719),.clk(gclk));
	jor g20462(.dina(w_n20719_0[2]),.dinb(n20716),.dout(n20720),.clk(gclk));
	jand g20463(.dina(n20720),.dinb(w_n20715_0[1]),.dout(n20721),.clk(gclk));
	jor g20464(.dina(w_n20721_0[2]),.dinb(w_n3955_22[1]),.dout(n20722),.clk(gclk));
	jand g20465(.dina(w_n20721_0[1]),.dinb(w_n3955_22[0]),.dout(n20723),.clk(gclk));
	jxor g20466(.dina(w_n20017_0[0]),.dinb(w_n4249_24[2]),.dout(n20724),.clk(gclk));
	jor g20467(.dina(n20724),.dinb(w_n20468_24[1]),.dout(n20725),.clk(gclk));
	jxor g20468(.dina(n20725),.dinb(w_n20359_0[0]),.dout(n20726),.clk(gclk));
	jnot g20469(.din(w_n20726_0[2]),.dout(n20727),.clk(gclk));
	jor g20470(.dina(n20727),.dinb(n20723),.dout(n20728),.clk(gclk));
	jand g20471(.dina(n20728),.dinb(w_n20722_0[1]),.dout(n20729),.clk(gclk));
	jor g20472(.dina(w_n20729_0[2]),.dinb(w_n3642_25[2]),.dout(n20730),.clk(gclk));
	jand g20473(.dina(w_n20729_0[1]),.dinb(w_n3642_25[1]),.dout(n20731),.clk(gclk));
	jxor g20474(.dina(w_n20024_0[0]),.dinb(w_n3955_21[2]),.dout(n20732),.clk(gclk));
	jor g20475(.dina(n20732),.dinb(w_n20468_24[0]),.dout(n20733),.clk(gclk));
	jxor g20476(.dina(n20733),.dinb(w_n20030_0[0]),.dout(n20734),.clk(gclk));
	jor g20477(.dina(w_n20734_0[2]),.dinb(n20731),.dout(n20735),.clk(gclk));
	jand g20478(.dina(n20735),.dinb(w_n20730_0[1]),.dout(n20736),.clk(gclk));
	jor g20479(.dina(w_n20736_0[2]),.dinb(w_n3368_23[0]),.dout(n20737),.clk(gclk));
	jand g20480(.dina(w_n20736_0[1]),.dinb(w_n3368_22[2]),.dout(n20738),.clk(gclk));
	jxor g20481(.dina(w_n20032_0[0]),.dinb(w_n3642_25[0]),.dout(n20739),.clk(gclk));
	jor g20482(.dina(n20739),.dinb(w_n20468_23[2]),.dout(n20740),.clk(gclk));
	jxor g20483(.dina(n20740),.dinb(w_n20038_0[0]),.dout(n20741),.clk(gclk));
	jor g20484(.dina(w_n20741_0[2]),.dinb(n20738),.dout(n20742),.clk(gclk));
	jand g20485(.dina(n20742),.dinb(w_n20737_0[1]),.dout(n20743),.clk(gclk));
	jor g20486(.dina(w_n20743_0[2]),.dinb(w_n3089_26[1]),.dout(n20744),.clk(gclk));
	jand g20487(.dina(w_n20743_0[1]),.dinb(w_n3089_26[0]),.dout(n20745),.clk(gclk));
	jxor g20488(.dina(w_n20040_0[0]),.dinb(w_n3368_22[1]),.dout(n20746),.clk(gclk));
	jor g20489(.dina(n20746),.dinb(w_n20468_23[1]),.dout(n20747),.clk(gclk));
	jxor g20490(.dina(n20747),.dinb(w_n20046_0[0]),.dout(n20748),.clk(gclk));
	jor g20491(.dina(w_n20748_0[2]),.dinb(n20745),.dout(n20749),.clk(gclk));
	jand g20492(.dina(n20749),.dinb(w_n20744_0[1]),.dout(n20750),.clk(gclk));
	jor g20493(.dina(w_n20750_0[2]),.dinb(w_n2833_24[0]),.dout(n20751),.clk(gclk));
	jand g20494(.dina(w_n20750_0[1]),.dinb(w_n2833_23[2]),.dout(n20752),.clk(gclk));
	jxor g20495(.dina(w_n20048_0[0]),.dinb(w_n3089_25[2]),.dout(n20753),.clk(gclk));
	jor g20496(.dina(n20753),.dinb(w_n20468_23[0]),.dout(n20754),.clk(gclk));
	jxor g20497(.dina(n20754),.dinb(w_n20372_0[0]),.dout(n20755),.clk(gclk));
	jnot g20498(.din(w_n20755_0[2]),.dout(n20756),.clk(gclk));
	jor g20499(.dina(n20756),.dinb(n20752),.dout(n20757),.clk(gclk));
	jand g20500(.dina(n20757),.dinb(w_n20751_0[1]),.dout(n20758),.clk(gclk));
	jor g20501(.dina(w_n20758_0[2]),.dinb(w_n2572_26[2]),.dout(n20759),.clk(gclk));
	jand g20502(.dina(w_n20758_0[1]),.dinb(w_n2572_26[1]),.dout(n20760),.clk(gclk));
	jxor g20503(.dina(w_n20055_0[0]),.dinb(w_n2833_23[1]),.dout(n20761),.clk(gclk));
	jor g20504(.dina(n20761),.dinb(w_n20468_22[2]),.dout(n20762),.clk(gclk));
	jxor g20505(.dina(n20762),.dinb(w_n20061_0[0]),.dout(n20763),.clk(gclk));
	jor g20506(.dina(w_n20763_0[2]),.dinb(n20760),.dout(n20764),.clk(gclk));
	jand g20507(.dina(n20764),.dinb(w_n20759_0[1]),.dout(n20765),.clk(gclk));
	jor g20508(.dina(w_n20765_0[2]),.dinb(w_n2345_24[2]),.dout(n20766),.clk(gclk));
	jand g20509(.dina(w_n20765_0[1]),.dinb(w_n2345_24[1]),.dout(n20767),.clk(gclk));
	jxor g20510(.dina(w_n20063_0[0]),.dinb(w_n2572_26[0]),.dout(n20768),.clk(gclk));
	jor g20511(.dina(n20768),.dinb(w_n20468_22[1]),.dout(n20769),.clk(gclk));
	jxor g20512(.dina(n20769),.dinb(w_n20069_0[0]),.dout(n20770),.clk(gclk));
	jor g20513(.dina(w_n20770_0[2]),.dinb(n20767),.dout(n20771),.clk(gclk));
	jand g20514(.dina(n20771),.dinb(w_n20766_0[1]),.dout(n20772),.clk(gclk));
	jor g20515(.dina(w_n20772_0[2]),.dinb(w_n2108_27[1]),.dout(n20773),.clk(gclk));
	jand g20516(.dina(w_n20772_0[1]),.dinb(w_n2108_27[0]),.dout(n20774),.clk(gclk));
	jxor g20517(.dina(w_n20071_0[0]),.dinb(w_n2345_24[0]),.dout(n20775),.clk(gclk));
	jor g20518(.dina(n20775),.dinb(w_n20468_22[0]),.dout(n20776),.clk(gclk));
	jxor g20519(.dina(n20776),.dinb(w_n20077_0[0]),.dout(n20777),.clk(gclk));
	jor g20520(.dina(w_n20777_0[2]),.dinb(n20774),.dout(n20778),.clk(gclk));
	jand g20521(.dina(n20778),.dinb(w_n20773_0[1]),.dout(n20779),.clk(gclk));
	jor g20522(.dina(w_n20779_0[2]),.dinb(w_n1912_25[2]),.dout(n20780),.clk(gclk));
	jand g20523(.dina(w_n20779_0[1]),.dinb(w_n1912_25[1]),.dout(n20781),.clk(gclk));
	jxor g20524(.dina(w_n20079_0[0]),.dinb(w_n2108_26[2]),.dout(n20782),.clk(gclk));
	jor g20525(.dina(n20782),.dinb(w_n20468_21[2]),.dout(n20783),.clk(gclk));
	jxor g20526(.dina(n20783),.dinb(w_n20085_0[0]),.dout(n20784),.clk(gclk));
	jor g20527(.dina(w_n20784_0[2]),.dinb(n20781),.dout(n20785),.clk(gclk));
	jand g20528(.dina(n20785),.dinb(w_n20780_0[1]),.dout(n20786),.clk(gclk));
	jor g20529(.dina(w_n20786_0[2]),.dinb(w_n1699_28[0]),.dout(n20787),.clk(gclk));
	jand g20530(.dina(w_n20786_0[1]),.dinb(w_n1699_27[2]),.dout(n20788),.clk(gclk));
	jxor g20531(.dina(w_n20087_0[0]),.dinb(w_n1912_25[0]),.dout(n20789),.clk(gclk));
	jor g20532(.dina(n20789),.dinb(w_n20468_21[1]),.dout(n20790),.clk(gclk));
	jxor g20533(.dina(n20790),.dinb(w_n20093_0[0]),.dout(n20791),.clk(gclk));
	jor g20534(.dina(w_n20791_0[2]),.dinb(n20788),.dout(n20792),.clk(gclk));
	jand g20535(.dina(n20792),.dinb(w_n20787_0[1]),.dout(n20793),.clk(gclk));
	jor g20536(.dina(w_n20793_0[2]),.dinb(w_n1516_26[1]),.dout(n20794),.clk(gclk));
	jand g20537(.dina(w_n20793_0[1]),.dinb(w_n1516_26[0]),.dout(n20795),.clk(gclk));
	jxor g20538(.dina(w_n20095_0[0]),.dinb(w_n1699_27[1]),.dout(n20796),.clk(gclk));
	jor g20539(.dina(n20796),.dinb(w_n20468_21[0]),.dout(n20797),.clk(gclk));
	jxor g20540(.dina(n20797),.dinb(w_n20391_0[0]),.dout(n20798),.clk(gclk));
	jnot g20541(.din(w_n20798_0[2]),.dout(n20799),.clk(gclk));
	jor g20542(.dina(n20799),.dinb(n20795),.dout(n20800),.clk(gclk));
	jand g20543(.dina(n20800),.dinb(w_n20794_0[1]),.dout(n20801),.clk(gclk));
	jor g20544(.dina(w_n20801_0[2]),.dinb(w_n1332_28[0]),.dout(n20802),.clk(gclk));
	jand g20545(.dina(w_n20801_0[1]),.dinb(w_n1332_27[2]),.dout(n20803),.clk(gclk));
	jxor g20546(.dina(w_n20102_0[0]),.dinb(w_n1516_25[2]),.dout(n20804),.clk(gclk));
	jor g20547(.dina(n20804),.dinb(w_n20468_20[2]),.dout(n20805),.clk(gclk));
	jxor g20548(.dina(n20805),.dinb(w_n20108_0[0]),.dout(n20806),.clk(gclk));
	jor g20549(.dina(w_n20806_0[2]),.dinb(n20803),.dout(n20807),.clk(gclk));
	jand g20550(.dina(n20807),.dinb(w_n20802_0[1]),.dout(n20808),.clk(gclk));
	jor g20551(.dina(w_n20808_0[2]),.dinb(w_n1173_27[0]),.dout(n20809),.clk(gclk));
	jand g20552(.dina(w_n20808_0[1]),.dinb(w_n1173_26[2]),.dout(n20810),.clk(gclk));
	jxor g20553(.dina(w_n20110_0[0]),.dinb(w_n1332_27[1]),.dout(n20811),.clk(gclk));
	jor g20554(.dina(n20811),.dinb(w_n20468_20[1]),.dout(n20812),.clk(gclk));
	jxor g20555(.dina(n20812),.dinb(w_n20398_0[0]),.dout(n20813),.clk(gclk));
	jnot g20556(.din(w_n20813_0[2]),.dout(n20814),.clk(gclk));
	jor g20557(.dina(n20814),.dinb(n20810),.dout(n20815),.clk(gclk));
	jand g20558(.dina(n20815),.dinb(w_n20809_0[1]),.dout(n20816),.clk(gclk));
	jor g20559(.dina(w_n20816_0[2]),.dinb(w_n1008_29[0]),.dout(n20817),.clk(gclk));
	jand g20560(.dina(w_n20816_0[1]),.dinb(w_n1008_28[2]),.dout(n20818),.clk(gclk));
	jxor g20561(.dina(w_n20117_0[0]),.dinb(w_n1173_26[1]),.dout(n20819),.clk(gclk));
	jor g20562(.dina(n20819),.dinb(w_n20468_20[0]),.dout(n20820),.clk(gclk));
	jxor g20563(.dina(n20820),.dinb(w_n20123_0[0]),.dout(n20821),.clk(gclk));
	jor g20564(.dina(w_n20821_0[2]),.dinb(n20818),.dout(n20822),.clk(gclk));
	jand g20565(.dina(n20822),.dinb(w_n20817_0[1]),.dout(n20823),.clk(gclk));
	jor g20566(.dina(w_n20823_0[2]),.dinb(w_n884_28[0]),.dout(n20824),.clk(gclk));
	jand g20567(.dina(w_n20823_0[1]),.dinb(w_n884_27[2]),.dout(n20825),.clk(gclk));
	jxor g20568(.dina(w_n20125_0[0]),.dinb(w_n1008_28[1]),.dout(n20826),.clk(gclk));
	jor g20569(.dina(n20826),.dinb(w_n20468_19[2]),.dout(n20827),.clk(gclk));
	jxor g20570(.dina(n20827),.dinb(w_n20131_0[0]),.dout(n20828),.clk(gclk));
	jor g20571(.dina(w_n20828_0[2]),.dinb(n20825),.dout(n20829),.clk(gclk));
	jand g20572(.dina(n20829),.dinb(w_n20824_0[1]),.dout(n20830),.clk(gclk));
	jor g20573(.dina(w_n20830_0[2]),.dinb(w_n743_29[0]),.dout(n20831),.clk(gclk));
	jand g20574(.dina(w_n20830_0[1]),.dinb(w_n743_28[2]),.dout(n20832),.clk(gclk));
	jxor g20575(.dina(w_n20133_0[0]),.dinb(w_n884_27[1]),.dout(n20833),.clk(gclk));
	jor g20576(.dina(n20833),.dinb(w_n20468_19[1]),.dout(n20834),.clk(gclk));
	jxor g20577(.dina(n20834),.dinb(w_n20408_0[0]),.dout(n20835),.clk(gclk));
	jnot g20578(.din(w_n20835_0[2]),.dout(n20836),.clk(gclk));
	jor g20579(.dina(n20836),.dinb(n20832),.dout(n20837),.clk(gclk));
	jand g20580(.dina(n20837),.dinb(w_n20831_0[1]),.dout(n20838),.clk(gclk));
	jor g20581(.dina(w_n20838_0[2]),.dinb(w_n635_29[0]),.dout(n20839),.clk(gclk));
	jxor g20582(.dina(w_n20140_0[0]),.dinb(w_n743_28[1]),.dout(n20840),.clk(gclk));
	jor g20583(.dina(n20840),.dinb(w_n20468_19[0]),.dout(n20841),.clk(gclk));
	jxor g20584(.dina(n20841),.dinb(w_n20203_0[0]),.dout(n20842),.clk(gclk));
	jnot g20585(.din(w_n20842_0[2]),.dout(n20843),.clk(gclk));
	jand g20586(.dina(w_n20838_0[1]),.dinb(w_n635_28[2]),.dout(n20844),.clk(gclk));
	jor g20587(.dina(n20844),.dinb(n20843),.dout(n20845),.clk(gclk));
	jand g20588(.dina(n20845),.dinb(w_n20839_0[1]),.dout(n20846),.clk(gclk));
	jor g20589(.dina(w_n20846_0[2]),.dinb(w_n515_30[0]),.dout(n20847),.clk(gclk));
	jand g20590(.dina(w_n20846_0[1]),.dinb(w_n515_29[2]),.dout(n20848),.clk(gclk));
	jxor g20591(.dina(w_n20147_0[0]),.dinb(w_n635_28[1]),.dout(n20849),.clk(gclk));
	jor g20592(.dina(n20849),.dinb(w_n20468_18[2]),.dout(n20850),.clk(gclk));
	jxor g20593(.dina(n20850),.dinb(w_n20153_0[0]),.dout(n20851),.clk(gclk));
	jor g20594(.dina(w_n20851_0[2]),.dinb(n20848),.dout(n20852),.clk(gclk));
	jand g20595(.dina(n20852),.dinb(w_n20847_0[1]),.dout(n20853),.clk(gclk));
	jor g20596(.dina(w_n20853_0[2]),.dinb(w_n443_30[0]),.dout(n20854),.clk(gclk));
	jand g20597(.dina(w_n20853_0[1]),.dinb(w_n443_29[2]),.dout(n20855),.clk(gclk));
	jxor g20598(.dina(w_n20155_0[0]),.dinb(w_n515_29[1]),.dout(n20856),.clk(gclk));
	jor g20599(.dina(n20856),.dinb(w_n20468_18[1]),.dout(n20857),.clk(gclk));
	jxor g20600(.dina(n20857),.dinb(w_n20418_0[0]),.dout(n20858),.clk(gclk));
	jnot g20601(.din(w_n20858_0[1]),.dout(n20859),.clk(gclk));
	jor g20602(.dina(w_n20859_0[1]),.dinb(n20855),.dout(n20860),.clk(gclk));
	jand g20603(.dina(n20860),.dinb(w_n20854_0[1]),.dout(n20861),.clk(gclk));
	jor g20604(.dina(w_n20861_0[2]),.dinb(w_n352_30[1]),.dout(n20862),.clk(gclk));
	jand g20605(.dina(w_n20861_0[1]),.dinb(w_n352_30[0]),.dout(n20863),.clk(gclk));
	jxor g20606(.dina(w_n20162_0[0]),.dinb(w_n443_29[1]),.dout(n20864),.clk(gclk));
	jor g20607(.dina(n20864),.dinb(w_n20468_18[0]),.dout(n20865),.clk(gclk));
	jxor g20608(.dina(n20865),.dinb(w_n20168_0[0]),.dout(n20866),.clk(gclk));
	jor g20609(.dina(w_n20866_0[2]),.dinb(n20863),.dout(n20867),.clk(gclk));
	jand g20610(.dina(n20867),.dinb(w_n20862_0[1]),.dout(n20868),.clk(gclk));
	jor g20611(.dina(w_n20868_0[2]),.dinb(w_n294_30[2]),.dout(n20869),.clk(gclk));
	jand g20612(.dina(w_n20868_0[1]),.dinb(w_n294_30[1]),.dout(n20870),.clk(gclk));
	jxor g20613(.dina(w_n20170_0[0]),.dinb(w_n352_29[2]),.dout(n20871),.clk(gclk));
	jor g20614(.dina(n20871),.dinb(w_n20468_17[2]),.dout(n20872),.clk(gclk));
	jxor g20615(.dina(n20872),.dinb(w_n20176_0[0]),.dout(n20873),.clk(gclk));
	jor g20616(.dina(w_n20873_0[2]),.dinb(n20870),.dout(n20874),.clk(gclk));
	jand g20617(.dina(n20874),.dinb(w_n20869_0[1]),.dout(n20875),.clk(gclk));
	jor g20618(.dina(w_n20875_0[2]),.dinb(w_n239_30[2]),.dout(n20876),.clk(gclk));
	jand g20619(.dina(w_n20875_0[1]),.dinb(w_n239_30[1]),.dout(n20877),.clk(gclk));
	jxor g20620(.dina(w_n20178_0[0]),.dinb(w_n294_30[0]),.dout(n20878),.clk(gclk));
	jor g20621(.dina(n20878),.dinb(w_n20468_17[1]),.dout(n20879),.clk(gclk));
	jxor g20622(.dina(n20879),.dinb(w_n20428_0[0]),.dout(n20880),.clk(gclk));
	jnot g20623(.din(w_n20880_0[2]),.dout(n20881),.clk(gclk));
	jor g20624(.dina(n20881),.dinb(n20877),.dout(n20882),.clk(gclk));
	jand g20625(.dina(n20882),.dinb(w_n20876_0[1]),.dout(n20883),.clk(gclk));
	jor g20626(.dina(w_n20883_0[2]),.dinb(w_n221_30[2]),.dout(n20884),.clk(gclk));
	jand g20627(.dina(w_n20883_0[1]),.dinb(w_n221_30[1]),.dout(n20885),.clk(gclk));
	jxor g20628(.dina(w_n20185_0[0]),.dinb(w_n239_30[0]),.dout(n20886),.clk(gclk));
	jor g20629(.dina(n20886),.dinb(w_n20468_17[0]),.dout(n20887),.clk(gclk));
	jxor g20630(.dina(n20887),.dinb(w_n20191_0[0]),.dout(n20888),.clk(gclk));
	jor g20631(.dina(w_n20888_0[2]),.dinb(n20885),.dout(n20889),.clk(gclk));
	jand g20632(.dina(n20889),.dinb(w_n20884_0[1]),.dout(n20890),.clk(gclk));
	jor g20633(.dina(w_n20890_0[2]),.dinb(w_n20472_0[1]),.dout(n20891),.clk(gclk));
	jand g20634(.dina(w_asqrt7_5[2]),.dinb(w_n20459_0[0]),.dout(n20892),.clk(gclk));
	jor g20635(.dina(n20892),.dinb(w_n20446_0[0]),.dout(n20893),.clk(gclk));
	jor g20636(.dina(w_n20893_0[1]),.dinb(w_n20891_0[1]),.dout(n20894),.clk(gclk));
	jand g20637(.dina(n20894),.dinb(w_n218_13[0]),.dout(n20895),.clk(gclk));
	jand g20638(.dina(w_n20468_16[2]),.dinb(w_n19523_0[0]),.dout(n20896),.clk(gclk));
	jand g20639(.dina(w_n20890_0[1]),.dinb(w_n20472_0[0]),.dout(n20897),.clk(gclk));
	jor g20640(.dina(w_n20897_0[1]),.dinb(w_n20896_0[1]),.dout(n20898),.clk(gclk));
	jand g20641(.dina(w_n20468_16[1]),.dinb(w_n20439_0[0]),.dout(n20899),.clk(gclk));
	jand g20642(.dina(w_n20440_0[0]),.dinb(w_asqrt63_22[0]),.dout(n20900),.clk(gclk));
	jand g20643(.dina(n20900),.dinb(w_n20464_0[0]),.dout(n20901),.clk(gclk));
	jnot g20644(.din(n20901),.dout(n20902),.clk(gclk));
	jor g20645(.dina(w_n20902_0[1]),.dinb(n20899),.dout(n20903),.clk(gclk));
	jnot g20646(.din(w_n20903_0[1]),.dout(n20904),.clk(gclk));
	jor g20647(.dina(n20904),.dinb(n20898),.dout(n20905),.clk(gclk));
	jor g20648(.dina(n20905),.dinb(n20895),.dout(asqrt_fa_7),.clk(gclk));
	jnot g20649(.din(w_a10_0[2]),.dout(n20907),.clk(gclk));
	jnot g20650(.din(w_a11_0[1]),.dout(n20908),.clk(gclk));
	jand g20651(.dina(w_n20908_0[1]),.dinb(w_n20907_1[2]),.dout(n20909),.clk(gclk));
	jand g20652(.dina(w_n20909_0[2]),.dinb(w_n20473_1[1]),.dout(n20910),.clk(gclk));
	jand g20653(.dina(w_asqrt6_32),.dinb(w_a12_0[1]),.dout(n20911),.clk(gclk));
	jor g20654(.dina(n20911),.dinb(w_n20910_0[1]),.dout(n20912),.clk(gclk));
	jand g20655(.dina(w_n20912_0[2]),.dinb(w_asqrt7_5[1]),.dout(n20913),.clk(gclk));
	jor g20656(.dina(w_n20912_0[1]),.dinb(w_asqrt7_5[0]),.dout(n20914),.clk(gclk));
	jand g20657(.dina(w_asqrt6_31[2]),.dinb(w_n20473_1[0]),.dout(n20915),.clk(gclk));
	jor g20658(.dina(n20915),.dinb(w_n20474_0[0]),.dout(n20916),.clk(gclk));
	jnot g20659(.din(w_n20475_0[1]),.dout(n20917),.clk(gclk));
	jnot g20660(.din(w_n20884_0[0]),.dout(n20918),.clk(gclk));
	jnot g20661(.din(w_n20876_0[0]),.dout(n20919),.clk(gclk));
	jnot g20662(.din(w_n20869_0[0]),.dout(n20920),.clk(gclk));
	jnot g20663(.din(w_n20862_0[0]),.dout(n20921),.clk(gclk));
	jnot g20664(.din(w_n20854_0[0]),.dout(n20922),.clk(gclk));
	jnot g20665(.din(w_n20847_0[0]),.dout(n20923),.clk(gclk));
	jnot g20666(.din(w_n20839_0[0]),.dout(n20924),.clk(gclk));
	jnot g20667(.din(w_n20831_0[0]),.dout(n20925),.clk(gclk));
	jnot g20668(.din(w_n20824_0[0]),.dout(n20926),.clk(gclk));
	jnot g20669(.din(w_n20817_0[0]),.dout(n20927),.clk(gclk));
	jnot g20670(.din(w_n20809_0[0]),.dout(n20928),.clk(gclk));
	jnot g20671(.din(w_n20802_0[0]),.dout(n20929),.clk(gclk));
	jnot g20672(.din(w_n20794_0[0]),.dout(n20930),.clk(gclk));
	jnot g20673(.din(w_n20787_0[0]),.dout(n20931),.clk(gclk));
	jnot g20674(.din(w_n20780_0[0]),.dout(n20932),.clk(gclk));
	jnot g20675(.din(w_n20773_0[0]),.dout(n20933),.clk(gclk));
	jnot g20676(.din(w_n20766_0[0]),.dout(n20934),.clk(gclk));
	jnot g20677(.din(w_n20759_0[0]),.dout(n20935),.clk(gclk));
	jnot g20678(.din(w_n20751_0[0]),.dout(n20936),.clk(gclk));
	jnot g20679(.din(w_n20744_0[0]),.dout(n20937),.clk(gclk));
	jnot g20680(.din(w_n20737_0[0]),.dout(n20938),.clk(gclk));
	jnot g20681(.din(w_n20730_0[0]),.dout(n20939),.clk(gclk));
	jnot g20682(.din(w_n20722_0[0]),.dout(n20940),.clk(gclk));
	jnot g20683(.din(w_n20715_0[0]),.dout(n20941),.clk(gclk));
	jnot g20684(.din(w_n20707_0[0]),.dout(n20942),.clk(gclk));
	jnot g20685(.din(w_n20700_0[0]),.dout(n20943),.clk(gclk));
	jnot g20686(.din(w_n20692_0[0]),.dout(n20944),.clk(gclk));
	jnot g20687(.din(w_n20685_0[0]),.dout(n20945),.clk(gclk));
	jnot g20688(.din(w_n20677_0[0]),.dout(n20946),.clk(gclk));
	jnot g20689(.din(w_n20670_0[0]),.dout(n20947),.clk(gclk));
	jnot g20690(.din(w_n20663_0[0]),.dout(n20948),.clk(gclk));
	jnot g20691(.din(w_n20656_0[0]),.dout(n20949),.clk(gclk));
	jnot g20692(.din(w_n20648_0[0]),.dout(n20950),.clk(gclk));
	jnot g20693(.din(w_n20641_0[0]),.dout(n20951),.clk(gclk));
	jnot g20694(.din(w_n20633_0[0]),.dout(n20952),.clk(gclk));
	jnot g20695(.din(w_n20626_0[0]),.dout(n20953),.clk(gclk));
	jnot g20696(.din(w_n20618_0[0]),.dout(n20954),.clk(gclk));
	jnot g20697(.din(w_n20610_0[0]),.dout(n20955),.clk(gclk));
	jnot g20698(.din(w_n20603_0[0]),.dout(n20956),.clk(gclk));
	jnot g20699(.din(w_n20596_0[0]),.dout(n20957),.clk(gclk));
	jnot g20700(.din(w_n20588_0[0]),.dout(n20958),.clk(gclk));
	jnot g20701(.din(w_n20581_0[0]),.dout(n20959),.clk(gclk));
	jnot g20702(.din(w_n20573_0[0]),.dout(n20960),.clk(gclk));
	jnot g20703(.din(w_n20566_0[0]),.dout(n20961),.clk(gclk));
	jnot g20704(.din(w_n20558_0[0]),.dout(n20962),.clk(gclk));
	jnot g20705(.din(w_n20551_0[0]),.dout(n20963),.clk(gclk));
	jnot g20706(.din(w_n20543_0[0]),.dout(n20964),.clk(gclk));
	jnot g20707(.din(w_n20536_0[0]),.dout(n20965),.clk(gclk));
	jnot g20708(.din(w_n20528_0[0]),.dout(n20966),.clk(gclk));
	jnot g20709(.din(w_n20521_0[0]),.dout(n20967),.clk(gclk));
	jnot g20710(.din(w_n20514_0[0]),.dout(n20968),.clk(gclk));
	jnot g20711(.din(w_n20507_0[0]),.dout(n20969),.clk(gclk));
	jnot g20712(.din(w_n20499_0[0]),.dout(n20970),.clk(gclk));
	jnot g20713(.din(w_n20488_0[0]),.dout(n20971),.clk(gclk));
	jnot g20714(.din(w_n20480_0[0]),.dout(n20972),.clk(gclk));
	jand g20715(.dina(w_asqrt7_4[2]),.dinb(w_a14_0[2]),.dout(n20973),.clk(gclk));
	jor g20716(.dina(n20973),.dinb(w_n20476_0[0]),.dout(n20974),.clk(gclk));
	jor g20717(.dina(n20974),.dinb(w_asqrt8_13[1]),.dout(n20975),.clk(gclk));
	jand g20718(.dina(w_asqrt7_4[1]),.dinb(w_n19524_0[1]),.dout(n20976),.clk(gclk));
	jor g20719(.dina(n20976),.dinb(w_n19525_0[0]),.dout(n20977),.clk(gclk));
	jand g20720(.dina(w_n20491_0[0]),.dinb(n20977),.dout(n20978),.clk(gclk));
	jand g20721(.dina(w_n20978_0[1]),.dinb(n20975),.dout(n20979),.clk(gclk));
	jor g20722(.dina(n20979),.dinb(n20972),.dout(n20980),.clk(gclk));
	jor g20723(.dina(n20980),.dinb(w_asqrt9_5[1]),.dout(n20981),.clk(gclk));
	jnot g20724(.din(w_n20496_0[1]),.dout(n20982),.clk(gclk));
	jand g20725(.dina(n20982),.dinb(n20981),.dout(n20983),.clk(gclk));
	jor g20726(.dina(n20983),.dinb(n20971),.dout(n20984),.clk(gclk));
	jor g20727(.dina(n20984),.dinb(w_asqrt10_13[1]),.dout(n20985),.clk(gclk));
	jand g20728(.dina(w_n20503_0[1]),.dinb(n20985),.dout(n20986),.clk(gclk));
	jor g20729(.dina(n20986),.dinb(n20970),.dout(n20987),.clk(gclk));
	jor g20730(.dina(n20987),.dinb(w_asqrt11_5[1]),.dout(n20988),.clk(gclk));
	jnot g20731(.din(w_n20511_0[1]),.dout(n20989),.clk(gclk));
	jand g20732(.dina(n20989),.dinb(n20988),.dout(n20990),.clk(gclk));
	jor g20733(.dina(n20990),.dinb(n20969),.dout(n20991),.clk(gclk));
	jor g20734(.dina(n20991),.dinb(w_asqrt12_13[2]),.dout(n20992),.clk(gclk));
	jnot g20735(.din(w_n20518_0[1]),.dout(n20993),.clk(gclk));
	jand g20736(.dina(n20993),.dinb(n20992),.dout(n20994),.clk(gclk));
	jor g20737(.dina(n20994),.dinb(n20968),.dout(n20995),.clk(gclk));
	jor g20738(.dina(n20995),.dinb(w_asqrt13_6[0]),.dout(n20996),.clk(gclk));
	jnot g20739(.din(w_n20525_0[1]),.dout(n20997),.clk(gclk));
	jand g20740(.dina(n20997),.dinb(n20996),.dout(n20998),.clk(gclk));
	jor g20741(.dina(n20998),.dinb(n20967),.dout(n20999),.clk(gclk));
	jor g20742(.dina(n20999),.dinb(w_asqrt14_14[0]),.dout(n21000),.clk(gclk));
	jand g20743(.dina(w_n20532_0[1]),.dinb(n21000),.dout(n21001),.clk(gclk));
	jor g20744(.dina(n21001),.dinb(n20966),.dout(n21002),.clk(gclk));
	jor g20745(.dina(n21002),.dinb(w_asqrt15_6[2]),.dout(n21003),.clk(gclk));
	jnot g20746(.din(w_n20540_0[1]),.dout(n21004),.clk(gclk));
	jand g20747(.dina(n21004),.dinb(n21003),.dout(n21005),.clk(gclk));
	jor g20748(.dina(n21005),.dinb(n20965),.dout(n21006),.clk(gclk));
	jor g20749(.dina(n21006),.dinb(w_asqrt16_14[0]),.dout(n21007),.clk(gclk));
	jand g20750(.dina(w_n20547_0[0]),.dinb(n21007),.dout(n21008),.clk(gclk));
	jor g20751(.dina(n21008),.dinb(n20964),.dout(n21009),.clk(gclk));
	jor g20752(.dina(n21009),.dinb(w_asqrt17_7[0]),.dout(n21010),.clk(gclk));
	jnot g20753(.din(w_n20555_0[1]),.dout(n21011),.clk(gclk));
	jand g20754(.dina(n21011),.dinb(n21010),.dout(n21012),.clk(gclk));
	jor g20755(.dina(n21012),.dinb(n20963),.dout(n21013),.clk(gclk));
	jor g20756(.dina(n21013),.dinb(w_asqrt18_14[1]),.dout(n21014),.clk(gclk));
	jand g20757(.dina(w_n20562_0[1]),.dinb(n21014),.dout(n21015),.clk(gclk));
	jor g20758(.dina(n21015),.dinb(n20962),.dout(n21016),.clk(gclk));
	jor g20759(.dina(n21016),.dinb(w_asqrt19_7[1]),.dout(n21017),.clk(gclk));
	jnot g20760(.din(w_n20570_0[1]),.dout(n21018),.clk(gclk));
	jand g20761(.dina(n21018),.dinb(n21017),.dout(n21019),.clk(gclk));
	jor g20762(.dina(n21019),.dinb(n20961),.dout(n21020),.clk(gclk));
	jor g20763(.dina(n21020),.dinb(w_asqrt20_14[1]),.dout(n21021),.clk(gclk));
	jand g20764(.dina(w_n20577_0[1]),.dinb(n21021),.dout(n21022),.clk(gclk));
	jor g20765(.dina(n21022),.dinb(n20960),.dout(n21023),.clk(gclk));
	jor g20766(.dina(n21023),.dinb(w_asqrt21_8[0]),.dout(n21024),.clk(gclk));
	jnot g20767(.din(w_n20585_0[1]),.dout(n21025),.clk(gclk));
	jand g20768(.dina(n21025),.dinb(n21024),.dout(n21026),.clk(gclk));
	jor g20769(.dina(n21026),.dinb(n20959),.dout(n21027),.clk(gclk));
	jor g20770(.dina(n21027),.dinb(w_asqrt22_14[2]),.dout(n21028),.clk(gclk));
	jand g20771(.dina(w_n20592_0[1]),.dinb(n21028),.dout(n21029),.clk(gclk));
	jor g20772(.dina(n21029),.dinb(n20958),.dout(n21030),.clk(gclk));
	jor g20773(.dina(n21030),.dinb(w_asqrt23_8[2]),.dout(n21031),.clk(gclk));
	jnot g20774(.din(w_n20600_0[1]),.dout(n21032),.clk(gclk));
	jand g20775(.dina(n21032),.dinb(n21031),.dout(n21033),.clk(gclk));
	jor g20776(.dina(n21033),.dinb(n20957),.dout(n21034),.clk(gclk));
	jor g20777(.dina(n21034),.dinb(w_asqrt24_14[2]),.dout(n21035),.clk(gclk));
	jnot g20778(.din(w_n20607_0[1]),.dout(n21036),.clk(gclk));
	jand g20779(.dina(n21036),.dinb(n21035),.dout(n21037),.clk(gclk));
	jor g20780(.dina(n21037),.dinb(n20956),.dout(n21038),.clk(gclk));
	jor g20781(.dina(n21038),.dinb(w_asqrt25_8[2]),.dout(n21039),.clk(gclk));
	jand g20782(.dina(w_n20614_0[1]),.dinb(n21039),.dout(n21040),.clk(gclk));
	jor g20783(.dina(n21040),.dinb(n20955),.dout(n21041),.clk(gclk));
	jor g20784(.dina(n21041),.dinb(w_asqrt26_14[2]),.dout(n21042),.clk(gclk));
	jand g20785(.dina(w_n20622_0[1]),.dinb(n21042),.dout(n21043),.clk(gclk));
	jor g20786(.dina(n21043),.dinb(n20954),.dout(n21044),.clk(gclk));
	jor g20787(.dina(n21044),.dinb(w_asqrt27_9[1]),.dout(n21045),.clk(gclk));
	jnot g20788(.din(w_n20630_0[1]),.dout(n21046),.clk(gclk));
	jand g20789(.dina(n21046),.dinb(n21045),.dout(n21047),.clk(gclk));
	jor g20790(.dina(n21047),.dinb(n20953),.dout(n21048),.clk(gclk));
	jor g20791(.dina(n21048),.dinb(w_asqrt28_15[0]),.dout(n21049),.clk(gclk));
	jand g20792(.dina(w_n20637_0[1]),.dinb(n21049),.dout(n21050),.clk(gclk));
	jor g20793(.dina(n21050),.dinb(n20952),.dout(n21051),.clk(gclk));
	jor g20794(.dina(n21051),.dinb(w_asqrt29_9[2]),.dout(n21052),.clk(gclk));
	jnot g20795(.din(w_n20645_0[1]),.dout(n21053),.clk(gclk));
	jand g20796(.dina(n21053),.dinb(n21052),.dout(n21054),.clk(gclk));
	jor g20797(.dina(n21054),.dinb(n20951),.dout(n21055),.clk(gclk));
	jor g20798(.dina(n21055),.dinb(w_asqrt30_15[1]),.dout(n21056),.clk(gclk));
	jand g20799(.dina(w_n20652_0[1]),.dinb(n21056),.dout(n21057),.clk(gclk));
	jor g20800(.dina(n21057),.dinb(n20950),.dout(n21058),.clk(gclk));
	jor g20801(.dina(n21058),.dinb(w_asqrt31_10[1]),.dout(n21059),.clk(gclk));
	jnot g20802(.din(w_n20660_0[1]),.dout(n21060),.clk(gclk));
	jand g20803(.dina(n21060),.dinb(n21059),.dout(n21061),.clk(gclk));
	jor g20804(.dina(n21061),.dinb(n20949),.dout(n21062),.clk(gclk));
	jor g20805(.dina(n21062),.dinb(w_asqrt32_15[1]),.dout(n21063),.clk(gclk));
	jnot g20806(.din(w_n20667_0[1]),.dout(n21064),.clk(gclk));
	jand g20807(.dina(n21064),.dinb(n21063),.dout(n21065),.clk(gclk));
	jor g20808(.dina(n21065),.dinb(n20948),.dout(n21066),.clk(gclk));
	jor g20809(.dina(n21066),.dinb(w_asqrt33_11[0]),.dout(n21067),.clk(gclk));
	jnot g20810(.din(w_n20674_0[1]),.dout(n21068),.clk(gclk));
	jand g20811(.dina(n21068),.dinb(n21067),.dout(n21069),.clk(gclk));
	jor g20812(.dina(n21069),.dinb(n20947),.dout(n21070),.clk(gclk));
	jor g20813(.dina(n21070),.dinb(w_asqrt34_15[2]),.dout(n21071),.clk(gclk));
	jand g20814(.dina(w_n20681_0[1]),.dinb(n21071),.dout(n21072),.clk(gclk));
	jor g20815(.dina(n21072),.dinb(n20946),.dout(n21073),.clk(gclk));
	jor g20816(.dina(n21073),.dinb(w_asqrt35_11[2]),.dout(n21074),.clk(gclk));
	jnot g20817(.din(w_n20689_0[1]),.dout(n21075),.clk(gclk));
	jand g20818(.dina(n21075),.dinb(n21074),.dout(n21076),.clk(gclk));
	jor g20819(.dina(n21076),.dinb(n20945),.dout(n21077),.clk(gclk));
	jor g20820(.dina(n21077),.dinb(w_asqrt36_15[2]),.dout(n21078),.clk(gclk));
	jand g20821(.dina(w_n20696_0[1]),.dinb(n21078),.dout(n21079),.clk(gclk));
	jor g20822(.dina(n21079),.dinb(n20944),.dout(n21080),.clk(gclk));
	jor g20823(.dina(n21080),.dinb(w_asqrt37_12[0]),.dout(n21081),.clk(gclk));
	jnot g20824(.din(w_n20704_0[1]),.dout(n21082),.clk(gclk));
	jand g20825(.dina(n21082),.dinb(n21081),.dout(n21083),.clk(gclk));
	jor g20826(.dina(n21083),.dinb(n20943),.dout(n21084),.clk(gclk));
	jor g20827(.dina(n21084),.dinb(w_asqrt38_16[0]),.dout(n21085),.clk(gclk));
	jand g20828(.dina(w_n20711_0[1]),.dinb(n21085),.dout(n21086),.clk(gclk));
	jor g20829(.dina(n21086),.dinb(n20942),.dout(n21087),.clk(gclk));
	jor g20830(.dina(n21087),.dinb(w_asqrt39_12[2]),.dout(n21088),.clk(gclk));
	jnot g20831(.din(w_n20719_0[1]),.dout(n21089),.clk(gclk));
	jand g20832(.dina(n21089),.dinb(n21088),.dout(n21090),.clk(gclk));
	jor g20833(.dina(n21090),.dinb(n20941),.dout(n21091),.clk(gclk));
	jor g20834(.dina(n21091),.dinb(w_asqrt40_16[0]),.dout(n21092),.clk(gclk));
	jand g20835(.dina(w_n20726_0[1]),.dinb(n21092),.dout(n21093),.clk(gclk));
	jor g20836(.dina(n21093),.dinb(n20940),.dout(n21094),.clk(gclk));
	jor g20837(.dina(n21094),.dinb(w_asqrt41_13[0]),.dout(n21095),.clk(gclk));
	jnot g20838(.din(w_n20734_0[1]),.dout(n21096),.clk(gclk));
	jand g20839(.dina(n21096),.dinb(n21095),.dout(n21097),.clk(gclk));
	jor g20840(.dina(n21097),.dinb(n20939),.dout(n21098),.clk(gclk));
	jor g20841(.dina(n21098),.dinb(w_asqrt42_16[1]),.dout(n21099),.clk(gclk));
	jnot g20842(.din(w_n20741_0[1]),.dout(n21100),.clk(gclk));
	jand g20843(.dina(n21100),.dinb(n21099),.dout(n21101),.clk(gclk));
	jor g20844(.dina(n21101),.dinb(n20938),.dout(n21102),.clk(gclk));
	jor g20845(.dina(n21102),.dinb(w_asqrt43_13[1]),.dout(n21103),.clk(gclk));
	jnot g20846(.din(w_n20748_0[1]),.dout(n21104),.clk(gclk));
	jand g20847(.dina(n21104),.dinb(n21103),.dout(n21105),.clk(gclk));
	jor g20848(.dina(n21105),.dinb(n20937),.dout(n21106),.clk(gclk));
	jor g20849(.dina(n21106),.dinb(w_asqrt44_16[1]),.dout(n21107),.clk(gclk));
	jand g20850(.dina(w_n20755_0[1]),.dinb(n21107),.dout(n21108),.clk(gclk));
	jor g20851(.dina(n21108),.dinb(n20936),.dout(n21109),.clk(gclk));
	jor g20852(.dina(n21109),.dinb(w_asqrt45_14[0]),.dout(n21110),.clk(gclk));
	jnot g20853(.din(w_n20763_0[1]),.dout(n21111),.clk(gclk));
	jand g20854(.dina(n21111),.dinb(n21110),.dout(n21112),.clk(gclk));
	jor g20855(.dina(n21112),.dinb(n20935),.dout(n21113),.clk(gclk));
	jor g20856(.dina(n21113),.dinb(w_asqrt46_16[1]),.dout(n21114),.clk(gclk));
	jnot g20857(.din(w_n20770_0[1]),.dout(n21115),.clk(gclk));
	jand g20858(.dina(n21115),.dinb(n21114),.dout(n21116),.clk(gclk));
	jor g20859(.dina(n21116),.dinb(n20934),.dout(n21117),.clk(gclk));
	jor g20860(.dina(n21117),.dinb(w_asqrt47_14[2]),.dout(n21118),.clk(gclk));
	jnot g20861(.din(w_n20777_0[1]),.dout(n21119),.clk(gclk));
	jand g20862(.dina(n21119),.dinb(n21118),.dout(n21120),.clk(gclk));
	jor g20863(.dina(n21120),.dinb(n20933),.dout(n21121),.clk(gclk));
	jor g20864(.dina(n21121),.dinb(w_asqrt48_16[2]),.dout(n21122),.clk(gclk));
	jnot g20865(.din(w_n20784_0[1]),.dout(n21123),.clk(gclk));
	jand g20866(.dina(n21123),.dinb(n21122),.dout(n21124),.clk(gclk));
	jor g20867(.dina(n21124),.dinb(n20932),.dout(n21125),.clk(gclk));
	jor g20868(.dina(n21125),.dinb(w_asqrt49_15[0]),.dout(n21126),.clk(gclk));
	jnot g20869(.din(w_n20791_0[1]),.dout(n21127),.clk(gclk));
	jand g20870(.dina(n21127),.dinb(n21126),.dout(n21128),.clk(gclk));
	jor g20871(.dina(n21128),.dinb(n20931),.dout(n21129),.clk(gclk));
	jor g20872(.dina(n21129),.dinb(w_asqrt50_17[0]),.dout(n21130),.clk(gclk));
	jand g20873(.dina(w_n20798_0[1]),.dinb(n21130),.dout(n21131),.clk(gclk));
	jor g20874(.dina(n21131),.dinb(n20930),.dout(n21132),.clk(gclk));
	jor g20875(.dina(n21132),.dinb(w_asqrt51_15[1]),.dout(n21133),.clk(gclk));
	jnot g20876(.din(w_n20806_0[1]),.dout(n21134),.clk(gclk));
	jand g20877(.dina(n21134),.dinb(n21133),.dout(n21135),.clk(gclk));
	jor g20878(.dina(n21135),.dinb(n20929),.dout(n21136),.clk(gclk));
	jor g20879(.dina(n21136),.dinb(w_asqrt52_17[0]),.dout(n21137),.clk(gclk));
	jand g20880(.dina(w_n20813_0[1]),.dinb(n21137),.dout(n21138),.clk(gclk));
	jor g20881(.dina(n21138),.dinb(n20928),.dout(n21139),.clk(gclk));
	jor g20882(.dina(n21139),.dinb(w_asqrt53_16[0]),.dout(n21140),.clk(gclk));
	jnot g20883(.din(w_n20821_0[1]),.dout(n21141),.clk(gclk));
	jand g20884(.dina(n21141),.dinb(n21140),.dout(n21142),.clk(gclk));
	jor g20885(.dina(n21142),.dinb(n20927),.dout(n21143),.clk(gclk));
	jor g20886(.dina(n21143),.dinb(w_asqrt54_17[0]),.dout(n21144),.clk(gclk));
	jnot g20887(.din(w_n20828_0[1]),.dout(n21145),.clk(gclk));
	jand g20888(.dina(n21145),.dinb(n21144),.dout(n21146),.clk(gclk));
	jor g20889(.dina(n21146),.dinb(n20926),.dout(n21147),.clk(gclk));
	jor g20890(.dina(n21147),.dinb(w_asqrt55_16[1]),.dout(n21148),.clk(gclk));
	jand g20891(.dina(w_n20835_0[1]),.dinb(n21148),.dout(n21149),.clk(gclk));
	jor g20892(.dina(n21149),.dinb(n20925),.dout(n21150),.clk(gclk));
	jor g20893(.dina(n21150),.dinb(w_asqrt56_17[1]),.dout(n21151),.clk(gclk));
	jand g20894(.dina(n21151),.dinb(w_n20842_0[1]),.dout(n21152),.clk(gclk));
	jor g20895(.dina(n21152),.dinb(n20924),.dout(n21153),.clk(gclk));
	jor g20896(.dina(n21153),.dinb(w_asqrt57_17[0]),.dout(n21154),.clk(gclk));
	jnot g20897(.din(w_n20851_0[1]),.dout(n21155),.clk(gclk));
	jand g20898(.dina(n21155),.dinb(n21154),.dout(n21156),.clk(gclk));
	jor g20899(.dina(n21156),.dinb(n20923),.dout(n21157),.clk(gclk));
	jor g20900(.dina(n21157),.dinb(w_asqrt58_17[2]),.dout(n21158),.clk(gclk));
	jand g20901(.dina(w_n20858_0[0]),.dinb(n21158),.dout(n21159),.clk(gclk));
	jor g20902(.dina(n21159),.dinb(n20922),.dout(n21160),.clk(gclk));
	jor g20903(.dina(n21160),.dinb(w_asqrt59_17[1]),.dout(n21161),.clk(gclk));
	jnot g20904(.din(w_n20866_0[1]),.dout(n21162),.clk(gclk));
	jand g20905(.dina(n21162),.dinb(n21161),.dout(n21163),.clk(gclk));
	jor g20906(.dina(n21163),.dinb(n20921),.dout(n21164),.clk(gclk));
	jor g20907(.dina(n21164),.dinb(w_asqrt60_17[2]),.dout(n21165),.clk(gclk));
	jnot g20908(.din(w_n20873_0[1]),.dout(n21166),.clk(gclk));
	jand g20909(.dina(n21166),.dinb(n21165),.dout(n21167),.clk(gclk));
	jor g20910(.dina(n21167),.dinb(n20920),.dout(n21168),.clk(gclk));
	jor g20911(.dina(n21168),.dinb(w_asqrt61_17[2]),.dout(n21169),.clk(gclk));
	jand g20912(.dina(w_n20880_0[1]),.dinb(n21169),.dout(n21170),.clk(gclk));
	jor g20913(.dina(n21170),.dinb(n20919),.dout(n21171),.clk(gclk));
	jor g20914(.dina(n21171),.dinb(w_asqrt62_17[2]),.dout(n21172),.clk(gclk));
	jnot g20915(.din(w_n20888_0[1]),.dout(n21173),.clk(gclk));
	jand g20916(.dina(n21173),.dinb(n21172),.dout(n21174),.clk(gclk));
	jor g20917(.dina(n21174),.dinb(n20918),.dout(n21175),.clk(gclk));
	jand g20918(.dina(w_n21175_0[1]),.dinb(w_n20471_0[1]),.dout(n21176),.clk(gclk));
	jnot g20919(.din(w_n20893_0[0]),.dout(n21177),.clk(gclk));
	jand g20920(.dina(n21177),.dinb(w_n21176_0[1]),.dout(n21178),.clk(gclk));
	jor g20921(.dina(n21178),.dinb(w_asqrt63_21[2]),.dout(n21179),.clk(gclk));
	jnot g20922(.din(w_n20896_0[0]),.dout(n21180),.clk(gclk));
	jor g20923(.dina(w_n21175_0[0]),.dinb(w_n20471_0[0]),.dout(n21181),.clk(gclk));
	jand g20924(.dina(w_n21181_1[1]),.dinb(n21180),.dout(n21182),.clk(gclk));
	jand g20925(.dina(w_n20903_0[0]),.dinb(n21182),.dout(n21183),.clk(gclk));
	jand g20926(.dina(n21183),.dinb(w_n21179_0[1]),.dout(n21184),.clk(gclk));
	jor g20927(.dina(w_n21184_7[2]),.dinb(n20917),.dout(n21185),.clk(gclk));
	jand g20928(.dina(n21185),.dinb(n20916),.dout(n21186),.clk(gclk));
	jand g20929(.dina(n21186),.dinb(n20914),.dout(n21187),.clk(gclk));
	jor g20930(.dina(n21187),.dinb(w_n20913_0[1]),.dout(n21188),.clk(gclk));
	jand g20931(.dina(w_n21188_0[2]),.dinb(w_asqrt8_13[0]),.dout(n21189),.clk(gclk));
	jor g20932(.dina(w_n21188_0[1]),.dinb(w_asqrt8_12[2]),.dout(n21190),.clk(gclk));
	jand g20933(.dina(w_asqrt6_31[1]),.dinb(w_n20475_0[0]),.dout(n21191),.clk(gclk));
	jand g20934(.dina(w_n20902_0[0]),.dinb(w_asqrt7_4[0]),.dout(n21192),.clk(gclk));
	jand g20935(.dina(n21192),.dinb(w_n21181_1[0]),.dout(n21193),.clk(gclk));
	jand g20936(.dina(n21193),.dinb(w_n21179_0[0]),.dout(n21194),.clk(gclk));
	jor g20937(.dina(n21194),.dinb(w_n21191_0[1]),.dout(n21195),.clk(gclk));
	jxor g20938(.dina(n21195),.dinb(w_a14_0[1]),.dout(n21196),.clk(gclk));
	jnot g20939(.din(w_n21196_0[1]),.dout(n21197),.clk(gclk));
	jand g20940(.dina(w_n21197_0[1]),.dinb(n21190),.dout(n21198),.clk(gclk));
	jor g20941(.dina(n21198),.dinb(w_n21189_0[1]),.dout(n21199),.clk(gclk));
	jand g20942(.dina(w_n21199_0[2]),.dinb(w_asqrt9_5[0]),.dout(n21200),.clk(gclk));
	jor g20943(.dina(w_n21199_0[1]),.dinb(w_asqrt9_4[2]),.dout(n21201),.clk(gclk));
	jxor g20944(.dina(w_n20479_0[0]),.dinb(w_n19791_8[0]),.dout(n21202),.clk(gclk));
	jand g20945(.dina(n21202),.dinb(w_asqrt6_31[0]),.dout(n21203),.clk(gclk));
	jxor g20946(.dina(n21203),.dinb(w_n20978_0[0]),.dout(n21204),.clk(gclk));
	jand g20947(.dina(w_n21204_0[1]),.dinb(n21201),.dout(n21205),.clk(gclk));
	jor g20948(.dina(n21205),.dinb(w_n21200_0[1]),.dout(n21206),.clk(gclk));
	jand g20949(.dina(w_n21206_0[2]),.dinb(w_asqrt10_13[0]),.dout(n21207),.clk(gclk));
	jor g20950(.dina(w_n21206_0[1]),.dinb(w_asqrt10_12[2]),.dout(n21208),.clk(gclk));
	jxor g20951(.dina(w_n20487_0[0]),.dinb(w_n19096_16[2]),.dout(n21209),.clk(gclk));
	jand g20952(.dina(n21209),.dinb(w_asqrt6_30[2]),.dout(n21210),.clk(gclk));
	jxor g20953(.dina(n21210),.dinb(w_n20496_0[0]),.dout(n21211),.clk(gclk));
	jnot g20954(.din(w_n21211_0[1]),.dout(n21212),.clk(gclk));
	jand g20955(.dina(w_n21212_0[1]),.dinb(n21208),.dout(n21213),.clk(gclk));
	jor g20956(.dina(n21213),.dinb(w_n21207_0[1]),.dout(n21214),.clk(gclk));
	jand g20957(.dina(w_n21214_0[2]),.dinb(w_asqrt11_5[0]),.dout(n21215),.clk(gclk));
	jor g20958(.dina(w_n21214_0[1]),.dinb(w_asqrt11_4[2]),.dout(n21216),.clk(gclk));
	jxor g20959(.dina(w_n20498_0[0]),.dinb(w_n18442_8[2]),.dout(n21217),.clk(gclk));
	jand g20960(.dina(n21217),.dinb(w_asqrt6_30[1]),.dout(n21218),.clk(gclk));
	jxor g20961(.dina(n21218),.dinb(w_n20503_0[0]),.dout(n21219),.clk(gclk));
	jand g20962(.dina(w_n21219_0[1]),.dinb(n21216),.dout(n21220),.clk(gclk));
	jor g20963(.dina(n21220),.dinb(w_n21215_0[1]),.dout(n21221),.clk(gclk));
	jand g20964(.dina(w_n21221_0[2]),.dinb(w_asqrt12_13[1]),.dout(n21222),.clk(gclk));
	jor g20965(.dina(w_n21221_0[1]),.dinb(w_asqrt12_13[0]),.dout(n21223),.clk(gclk));
	jxor g20966(.dina(w_n20506_0[0]),.dinb(w_n17769_17[1]),.dout(n21224),.clk(gclk));
	jand g20967(.dina(n21224),.dinb(w_asqrt6_30[0]),.dout(n21225),.clk(gclk));
	jxor g20968(.dina(n21225),.dinb(w_n20511_0[0]),.dout(n21226),.clk(gclk));
	jnot g20969(.din(w_n21226_0[1]),.dout(n21227),.clk(gclk));
	jand g20970(.dina(w_n21227_0[1]),.dinb(n21223),.dout(n21228),.clk(gclk));
	jor g20971(.dina(n21228),.dinb(w_n21222_0[1]),.dout(n21229),.clk(gclk));
	jand g20972(.dina(w_n21229_0[2]),.dinb(w_asqrt13_5[2]),.dout(n21230),.clk(gclk));
	jor g20973(.dina(w_n21229_0[1]),.dinb(w_asqrt13_5[1]),.dout(n21231),.clk(gclk));
	jxor g20974(.dina(w_n20513_0[0]),.dinb(w_n17134_9[2]),.dout(n21232),.clk(gclk));
	jand g20975(.dina(n21232),.dinb(w_asqrt6_29[2]),.dout(n21233),.clk(gclk));
	jxor g20976(.dina(n21233),.dinb(w_n20518_0[0]),.dout(n21234),.clk(gclk));
	jnot g20977(.din(w_n21234_0[1]),.dout(n21235),.clk(gclk));
	jand g20978(.dina(w_n21235_0[1]),.dinb(n21231),.dout(n21236),.clk(gclk));
	jor g20979(.dina(n21236),.dinb(w_n21230_0[1]),.dout(n21237),.clk(gclk));
	jand g20980(.dina(w_n21237_0[2]),.dinb(w_asqrt14_13[2]),.dout(n21238),.clk(gclk));
	jor g20981(.dina(w_n21237_0[1]),.dinb(w_asqrt14_13[1]),.dout(n21239),.clk(gclk));
	jxor g20982(.dina(w_n20520_0[0]),.dinb(w_n16489_17[2]),.dout(n21240),.clk(gclk));
	jand g20983(.dina(n21240),.dinb(w_asqrt6_29[1]),.dout(n21241),.clk(gclk));
	jxor g20984(.dina(n21241),.dinb(w_n20525_0[0]),.dout(n21242),.clk(gclk));
	jnot g20985(.din(w_n21242_0[1]),.dout(n21243),.clk(gclk));
	jand g20986(.dina(w_n21243_0[1]),.dinb(n21239),.dout(n21244),.clk(gclk));
	jor g20987(.dina(n21244),.dinb(w_n21238_0[1]),.dout(n21245),.clk(gclk));
	jand g20988(.dina(w_n21245_0[2]),.dinb(w_asqrt15_6[1]),.dout(n21246),.clk(gclk));
	jor g20989(.dina(w_n21245_0[1]),.dinb(w_asqrt15_6[0]),.dout(n21247),.clk(gclk));
	jxor g20990(.dina(w_n20527_0[0]),.dinb(w_n15878_10[2]),.dout(n21248),.clk(gclk));
	jand g20991(.dina(n21248),.dinb(w_asqrt6_29[0]),.dout(n21249),.clk(gclk));
	jxor g20992(.dina(n21249),.dinb(w_n20532_0[0]),.dout(n21250),.clk(gclk));
	jand g20993(.dina(w_n21250_0[1]),.dinb(n21247),.dout(n21251),.clk(gclk));
	jor g20994(.dina(n21251),.dinb(w_n21246_0[1]),.dout(n21252),.clk(gclk));
	jand g20995(.dina(w_n21252_0[2]),.dinb(w_asqrt16_13[2]),.dout(n21253),.clk(gclk));
	jor g20996(.dina(w_n21252_0[1]),.dinb(w_asqrt16_13[1]),.dout(n21254),.clk(gclk));
	jxor g20997(.dina(w_n20535_0[0]),.dinb(w_n15260_18[1]),.dout(n21255),.clk(gclk));
	jand g20998(.dina(n21255),.dinb(w_asqrt6_28[2]),.dout(n21256),.clk(gclk));
	jxor g20999(.dina(n21256),.dinb(w_n20540_0[0]),.dout(n21257),.clk(gclk));
	jnot g21000(.din(w_n21257_0[1]),.dout(n21258),.clk(gclk));
	jand g21001(.dina(w_n21258_0[1]),.dinb(n21254),.dout(n21259),.clk(gclk));
	jor g21002(.dina(n21259),.dinb(w_n21253_0[1]),.dout(n21260),.clk(gclk));
	jand g21003(.dina(w_n21260_0[2]),.dinb(w_asqrt17_6[2]),.dout(n21261),.clk(gclk));
	jor g21004(.dina(w_n21260_0[1]),.dinb(w_asqrt17_6[1]),.dout(n21262),.clk(gclk));
	jxor g21005(.dina(w_n20542_0[0]),.dinb(w_n14674_11[1]),.dout(n21263),.clk(gclk));
	jand g21006(.dina(n21263),.dinb(w_asqrt6_28[1]),.dout(n21264),.clk(gclk));
	jxor g21007(.dina(n21264),.dinb(w_n20548_0[0]),.dout(n21265),.clk(gclk));
	jnot g21008(.din(w_n21265_0[1]),.dout(n21266),.clk(gclk));
	jand g21009(.dina(w_n21266_0[1]),.dinb(n21262),.dout(n21267),.clk(gclk));
	jor g21010(.dina(n21267),.dinb(w_n21261_0[1]),.dout(n21268),.clk(gclk));
	jand g21011(.dina(w_n21268_0[2]),.dinb(w_asqrt18_14[0]),.dout(n21269),.clk(gclk));
	jor g21012(.dina(w_n21268_0[1]),.dinb(w_asqrt18_13[2]),.dout(n21270),.clk(gclk));
	jxor g21013(.dina(w_n20550_0[0]),.dinb(w_n14078_18[2]),.dout(n21271),.clk(gclk));
	jand g21014(.dina(n21271),.dinb(w_asqrt6_28[0]),.dout(n21272),.clk(gclk));
	jxor g21015(.dina(n21272),.dinb(w_n20555_0[0]),.dout(n21273),.clk(gclk));
	jnot g21016(.din(w_n21273_0[1]),.dout(n21274),.clk(gclk));
	jand g21017(.dina(w_n21274_0[1]),.dinb(n21270),.dout(n21275),.clk(gclk));
	jor g21018(.dina(n21275),.dinb(w_n21269_0[1]),.dout(n21276),.clk(gclk));
	jand g21019(.dina(w_n21276_0[2]),.dinb(w_asqrt19_7[0]),.dout(n21277),.clk(gclk));
	jor g21020(.dina(w_n21276_0[1]),.dinb(w_asqrt19_6[2]),.dout(n21278),.clk(gclk));
	jxor g21021(.dina(w_n20557_0[0]),.dinb(w_n13515_12[1]),.dout(n21279),.clk(gclk));
	jand g21022(.dina(n21279),.dinb(w_asqrt6_27[2]),.dout(n21280),.clk(gclk));
	jxor g21023(.dina(n21280),.dinb(w_n20562_0[0]),.dout(n21281),.clk(gclk));
	jand g21024(.dina(w_n21281_0[1]),.dinb(n21278),.dout(n21282),.clk(gclk));
	jor g21025(.dina(n21282),.dinb(w_n21277_0[1]),.dout(n21283),.clk(gclk));
	jand g21026(.dina(w_n21283_0[2]),.dinb(w_asqrt20_14[0]),.dout(n21284),.clk(gclk));
	jor g21027(.dina(w_n21283_0[1]),.dinb(w_asqrt20_13[2]),.dout(n21285),.clk(gclk));
	jxor g21028(.dina(w_n20565_0[0]),.dinb(w_n12947_19[1]),.dout(n21286),.clk(gclk));
	jand g21029(.dina(n21286),.dinb(w_asqrt6_27[1]),.dout(n21287),.clk(gclk));
	jxor g21030(.dina(n21287),.dinb(w_n20570_0[0]),.dout(n21288),.clk(gclk));
	jnot g21031(.din(w_n21288_0[1]),.dout(n21289),.clk(gclk));
	jand g21032(.dina(w_n21289_0[1]),.dinb(n21285),.dout(n21290),.clk(gclk));
	jor g21033(.dina(n21290),.dinb(w_n21284_0[1]),.dout(n21291),.clk(gclk));
	jand g21034(.dina(w_n21291_0[2]),.dinb(w_asqrt21_7[2]),.dout(n21292),.clk(gclk));
	jor g21035(.dina(w_n21291_0[1]),.dinb(w_asqrt21_7[1]),.dout(n21293),.clk(gclk));
	jxor g21036(.dina(w_n20572_0[0]),.dinb(w_n12410_13[0]),.dout(n21294),.clk(gclk));
	jand g21037(.dina(n21294),.dinb(w_asqrt6_27[0]),.dout(n21295),.clk(gclk));
	jxor g21038(.dina(n21295),.dinb(w_n20577_0[0]),.dout(n21296),.clk(gclk));
	jand g21039(.dina(w_n21296_0[1]),.dinb(n21293),.dout(n21297),.clk(gclk));
	jor g21040(.dina(n21297),.dinb(w_n21292_0[1]),.dout(n21298),.clk(gclk));
	jand g21041(.dina(w_n21298_0[2]),.dinb(w_asqrt22_14[1]),.dout(n21299),.clk(gclk));
	jor g21042(.dina(w_n21298_0[1]),.dinb(w_asqrt22_14[0]),.dout(n21300),.clk(gclk));
	jxor g21043(.dina(w_n20580_0[0]),.dinb(w_n11858_19[2]),.dout(n21301),.clk(gclk));
	jand g21044(.dina(n21301),.dinb(w_asqrt6_26[2]),.dout(n21302),.clk(gclk));
	jxor g21045(.dina(n21302),.dinb(w_n20585_0[0]),.dout(n21303),.clk(gclk));
	jnot g21046(.din(w_n21303_0[1]),.dout(n21304),.clk(gclk));
	jand g21047(.dina(w_n21304_0[1]),.dinb(n21300),.dout(n21305),.clk(gclk));
	jor g21048(.dina(n21305),.dinb(w_n21299_0[1]),.dout(n21306),.clk(gclk));
	jand g21049(.dina(w_n21306_0[2]),.dinb(w_asqrt23_8[1]),.dout(n21307),.clk(gclk));
	jor g21050(.dina(w_n21306_0[1]),.dinb(w_asqrt23_8[0]),.dout(n21308),.clk(gclk));
	jxor g21051(.dina(w_n20587_0[0]),.dinb(w_n11347_13[2]),.dout(n21309),.clk(gclk));
	jand g21052(.dina(n21309),.dinb(w_asqrt6_26[1]),.dout(n21310),.clk(gclk));
	jxor g21053(.dina(n21310),.dinb(w_n20592_0[0]),.dout(n21311),.clk(gclk));
	jand g21054(.dina(w_n21311_0[1]),.dinb(n21308),.dout(n21312),.clk(gclk));
	jor g21055(.dina(n21312),.dinb(w_n21307_0[1]),.dout(n21313),.clk(gclk));
	jand g21056(.dina(w_n21313_0[2]),.dinb(w_asqrt24_14[1]),.dout(n21314),.clk(gclk));
	jor g21057(.dina(w_n21313_0[1]),.dinb(w_asqrt24_14[0]),.dout(n21315),.clk(gclk));
	jxor g21058(.dina(w_n20595_0[0]),.dinb(w_n10824_20[1]),.dout(n21316),.clk(gclk));
	jand g21059(.dina(n21316),.dinb(w_asqrt6_26[0]),.dout(n21317),.clk(gclk));
	jxor g21060(.dina(n21317),.dinb(w_n20600_0[0]),.dout(n21318),.clk(gclk));
	jnot g21061(.din(w_n21318_0[1]),.dout(n21319),.clk(gclk));
	jand g21062(.dina(w_n21319_0[1]),.dinb(n21315),.dout(n21320),.clk(gclk));
	jor g21063(.dina(n21320),.dinb(w_n21314_0[1]),.dout(n21321),.clk(gclk));
	jand g21064(.dina(w_n21321_0[2]),.dinb(w_asqrt25_8[1]),.dout(n21322),.clk(gclk));
	jor g21065(.dina(w_n21321_0[1]),.dinb(w_asqrt25_8[0]),.dout(n21323),.clk(gclk));
	jxor g21066(.dina(w_n20602_0[0]),.dinb(w_n10328_14[2]),.dout(n21324),.clk(gclk));
	jand g21067(.dina(n21324),.dinb(w_asqrt6_25[2]),.dout(n21325),.clk(gclk));
	jxor g21068(.dina(n21325),.dinb(w_n20607_0[0]),.dout(n21326),.clk(gclk));
	jnot g21069(.din(w_n21326_0[1]),.dout(n21327),.clk(gclk));
	jand g21070(.dina(w_n21327_0[1]),.dinb(n21323),.dout(n21328),.clk(gclk));
	jor g21071(.dina(n21328),.dinb(w_n21322_0[1]),.dout(n21329),.clk(gclk));
	jand g21072(.dina(w_n21329_0[2]),.dinb(w_asqrt26_14[1]),.dout(n21330),.clk(gclk));
	jor g21073(.dina(w_n21329_0[1]),.dinb(w_asqrt26_14[0]),.dout(n21331),.clk(gclk));
	jxor g21074(.dina(w_n20609_0[0]),.dinb(w_n9832_21[0]),.dout(n21332),.clk(gclk));
	jand g21075(.dina(n21332),.dinb(w_asqrt6_25[1]),.dout(n21333),.clk(gclk));
	jxor g21076(.dina(n21333),.dinb(w_n20614_0[0]),.dout(n21334),.clk(gclk));
	jand g21077(.dina(w_n21334_0[1]),.dinb(n21331),.dout(n21335),.clk(gclk));
	jor g21078(.dina(n21335),.dinb(w_n21330_0[1]),.dout(n21336),.clk(gclk));
	jand g21079(.dina(w_n21336_0[2]),.dinb(w_asqrt27_9[0]),.dout(n21337),.clk(gclk));
	jor g21080(.dina(w_n21336_0[1]),.dinb(w_asqrt27_8[2]),.dout(n21338),.clk(gclk));
	jxor g21081(.dina(w_n20617_0[0]),.dinb(w_n9369_15[2]),.dout(n21339),.clk(gclk));
	jand g21082(.dina(n21339),.dinb(w_asqrt6_25[0]),.dout(n21340),.clk(gclk));
	jxor g21083(.dina(n21340),.dinb(w_n20622_0[0]),.dout(n21341),.clk(gclk));
	jand g21084(.dina(w_n21341_0[1]),.dinb(n21338),.dout(n21342),.clk(gclk));
	jor g21085(.dina(n21342),.dinb(w_n21337_0[1]),.dout(n21343),.clk(gclk));
	jand g21086(.dina(w_n21343_0[2]),.dinb(w_asqrt28_14[2]),.dout(n21344),.clk(gclk));
	jor g21087(.dina(w_n21343_0[1]),.dinb(w_asqrt28_14[1]),.dout(n21345),.clk(gclk));
	jxor g21088(.dina(w_n20625_0[0]),.dinb(w_n8890_21[1]),.dout(n21346),.clk(gclk));
	jand g21089(.dina(n21346),.dinb(w_asqrt6_24[2]),.dout(n21347),.clk(gclk));
	jxor g21090(.dina(n21347),.dinb(w_n20630_0[0]),.dout(n21348),.clk(gclk));
	jnot g21091(.din(w_n21348_0[1]),.dout(n21349),.clk(gclk));
	jand g21092(.dina(w_n21349_0[1]),.dinb(n21345),.dout(n21350),.clk(gclk));
	jor g21093(.dina(n21350),.dinb(w_n21344_0[1]),.dout(n21351),.clk(gclk));
	jand g21094(.dina(w_n21351_0[2]),.dinb(w_asqrt29_9[1]),.dout(n21352),.clk(gclk));
	jor g21095(.dina(w_n21351_0[1]),.dinb(w_asqrt29_9[0]),.dout(n21353),.clk(gclk));
	jxor g21096(.dina(w_n20632_0[0]),.dinb(w_n8449_16[1]),.dout(n21354),.clk(gclk));
	jand g21097(.dina(n21354),.dinb(w_asqrt6_24[1]),.dout(n21355),.clk(gclk));
	jxor g21098(.dina(n21355),.dinb(w_n20637_0[0]),.dout(n21356),.clk(gclk));
	jand g21099(.dina(w_n21356_0[1]),.dinb(n21353),.dout(n21357),.clk(gclk));
	jor g21100(.dina(n21357),.dinb(w_n21352_0[1]),.dout(n21358),.clk(gclk));
	jand g21101(.dina(w_n21358_0[2]),.dinb(w_asqrt30_15[0]),.dout(n21359),.clk(gclk));
	jor g21102(.dina(w_n21358_0[1]),.dinb(w_asqrt30_14[2]),.dout(n21360),.clk(gclk));
	jxor g21103(.dina(w_n20640_0[0]),.dinb(w_n8003_22[0]),.dout(n21361),.clk(gclk));
	jand g21104(.dina(n21361),.dinb(w_asqrt6_24[0]),.dout(n21362),.clk(gclk));
	jxor g21105(.dina(n21362),.dinb(w_n20645_0[0]),.dout(n21363),.clk(gclk));
	jnot g21106(.din(w_n21363_0[1]),.dout(n21364),.clk(gclk));
	jand g21107(.dina(w_n21364_0[1]),.dinb(n21360),.dout(n21365),.clk(gclk));
	jor g21108(.dina(n21365),.dinb(w_n21359_0[1]),.dout(n21366),.clk(gclk));
	jand g21109(.dina(w_n21366_0[2]),.dinb(w_asqrt31_10[0]),.dout(n21367),.clk(gclk));
	jor g21110(.dina(w_n21366_0[1]),.dinb(w_asqrt31_9[2]),.dout(n21368),.clk(gclk));
	jxor g21111(.dina(w_n20647_0[0]),.dinb(w_n7581_17[1]),.dout(n21369),.clk(gclk));
	jand g21112(.dina(n21369),.dinb(w_asqrt6_23[2]),.dout(n21370),.clk(gclk));
	jxor g21113(.dina(n21370),.dinb(w_n20652_0[0]),.dout(n21371),.clk(gclk));
	jand g21114(.dina(w_n21371_0[1]),.dinb(n21368),.dout(n21372),.clk(gclk));
	jor g21115(.dina(n21372),.dinb(w_n21367_0[1]),.dout(n21373),.clk(gclk));
	jand g21116(.dina(w_n21373_0[2]),.dinb(w_asqrt32_15[0]),.dout(n21374),.clk(gclk));
	jor g21117(.dina(w_n21373_0[1]),.dinb(w_asqrt32_14[2]),.dout(n21375),.clk(gclk));
	jxor g21118(.dina(w_n20655_0[0]),.dinb(w_n7154_22[1]),.dout(n21376),.clk(gclk));
	jand g21119(.dina(n21376),.dinb(w_asqrt6_23[1]),.dout(n21377),.clk(gclk));
	jxor g21120(.dina(n21377),.dinb(w_n20660_0[0]),.dout(n21378),.clk(gclk));
	jnot g21121(.din(w_n21378_0[1]),.dout(n21379),.clk(gclk));
	jand g21122(.dina(w_n21379_0[1]),.dinb(n21375),.dout(n21380),.clk(gclk));
	jor g21123(.dina(n21380),.dinb(w_n21374_0[1]),.dout(n21381),.clk(gclk));
	jand g21124(.dina(w_n21381_0[2]),.dinb(w_asqrt33_10[2]),.dout(n21382),.clk(gclk));
	jor g21125(.dina(w_n21381_0[1]),.dinb(w_asqrt33_10[1]),.dout(n21383),.clk(gclk));
	jxor g21126(.dina(w_n20662_0[0]),.dinb(w_n6758_18[0]),.dout(n21384),.clk(gclk));
	jand g21127(.dina(n21384),.dinb(w_asqrt6_23[0]),.dout(n21385),.clk(gclk));
	jxor g21128(.dina(n21385),.dinb(w_n20667_0[0]),.dout(n21386),.clk(gclk));
	jnot g21129(.din(w_n21386_0[1]),.dout(n21387),.clk(gclk));
	jand g21130(.dina(w_n21387_0[1]),.dinb(n21383),.dout(n21388),.clk(gclk));
	jor g21131(.dina(n21388),.dinb(w_n21382_0[1]),.dout(n21389),.clk(gclk));
	jand g21132(.dina(w_n21389_0[2]),.dinb(w_asqrt34_15[1]),.dout(n21390),.clk(gclk));
	jor g21133(.dina(w_n21389_0[1]),.dinb(w_asqrt34_15[0]),.dout(n21391),.clk(gclk));
	jxor g21134(.dina(w_n20669_0[0]),.dinb(w_n6357_22[2]),.dout(n21392),.clk(gclk));
	jand g21135(.dina(n21392),.dinb(w_asqrt6_22[2]),.dout(n21393),.clk(gclk));
	jxor g21136(.dina(n21393),.dinb(w_n20674_0[0]),.dout(n21394),.clk(gclk));
	jnot g21137(.din(w_n21394_0[1]),.dout(n21395),.clk(gclk));
	jand g21138(.dina(w_n21395_0[1]),.dinb(n21391),.dout(n21396),.clk(gclk));
	jor g21139(.dina(n21396),.dinb(w_n21390_0[1]),.dout(n21397),.clk(gclk));
	jand g21140(.dina(w_n21397_0[2]),.dinb(w_asqrt35_11[1]),.dout(n21398),.clk(gclk));
	jor g21141(.dina(w_n21397_0[1]),.dinb(w_asqrt35_11[0]),.dout(n21399),.clk(gclk));
	jxor g21142(.dina(w_n20676_0[0]),.dinb(w_n5989_18[2]),.dout(n21400),.clk(gclk));
	jand g21143(.dina(n21400),.dinb(w_asqrt6_22[1]),.dout(n21401),.clk(gclk));
	jxor g21144(.dina(n21401),.dinb(w_n20681_0[0]),.dout(n21402),.clk(gclk));
	jand g21145(.dina(w_n21402_0[1]),.dinb(n21399),.dout(n21403),.clk(gclk));
	jor g21146(.dina(n21403),.dinb(w_n21398_0[1]),.dout(n21404),.clk(gclk));
	jand g21147(.dina(w_n21404_0[2]),.dinb(w_asqrt36_15[1]),.dout(n21405),.clk(gclk));
	jor g21148(.dina(w_n21404_0[1]),.dinb(w_asqrt36_15[0]),.dout(n21406),.clk(gclk));
	jxor g21149(.dina(w_n20684_0[0]),.dinb(w_n5606_23[0]),.dout(n21407),.clk(gclk));
	jand g21150(.dina(n21407),.dinb(w_asqrt6_22[0]),.dout(n21408),.clk(gclk));
	jxor g21151(.dina(n21408),.dinb(w_n20689_0[0]),.dout(n21409),.clk(gclk));
	jnot g21152(.din(w_n21409_0[1]),.dout(n21410),.clk(gclk));
	jand g21153(.dina(w_n21410_0[1]),.dinb(n21406),.dout(n21411),.clk(gclk));
	jor g21154(.dina(n21411),.dinb(w_n21405_0[1]),.dout(n21412),.clk(gclk));
	jand g21155(.dina(w_n21412_0[2]),.dinb(w_asqrt37_11[2]),.dout(n21413),.clk(gclk));
	jor g21156(.dina(w_n21412_0[1]),.dinb(w_asqrt37_11[1]),.dout(n21414),.clk(gclk));
	jxor g21157(.dina(w_n20691_0[0]),.dinb(w_n5259_19[2]),.dout(n21415),.clk(gclk));
	jand g21158(.dina(n21415),.dinb(w_asqrt6_21[2]),.dout(n21416),.clk(gclk));
	jxor g21159(.dina(n21416),.dinb(w_n20696_0[0]),.dout(n21417),.clk(gclk));
	jand g21160(.dina(w_n21417_0[1]),.dinb(n21414),.dout(n21418),.clk(gclk));
	jor g21161(.dina(n21418),.dinb(w_n21413_0[1]),.dout(n21419),.clk(gclk));
	jand g21162(.dina(w_n21419_0[2]),.dinb(w_asqrt38_15[2]),.dout(n21420),.clk(gclk));
	jor g21163(.dina(w_n21419_0[1]),.dinb(w_asqrt38_15[1]),.dout(n21421),.clk(gclk));
	jxor g21164(.dina(w_n20699_0[0]),.dinb(w_n4902_23[2]),.dout(n21422),.clk(gclk));
	jand g21165(.dina(n21422),.dinb(w_asqrt6_21[1]),.dout(n21423),.clk(gclk));
	jxor g21166(.dina(n21423),.dinb(w_n20704_0[0]),.dout(n21424),.clk(gclk));
	jnot g21167(.din(w_n21424_0[1]),.dout(n21425),.clk(gclk));
	jand g21168(.dina(w_n21425_0[1]),.dinb(n21421),.dout(n21426),.clk(gclk));
	jor g21169(.dina(n21426),.dinb(w_n21420_0[1]),.dout(n21427),.clk(gclk));
	jand g21170(.dina(w_n21427_0[2]),.dinb(w_asqrt39_12[1]),.dout(n21428),.clk(gclk));
	jor g21171(.dina(w_n21427_0[1]),.dinb(w_asqrt39_12[0]),.dout(n21429),.clk(gclk));
	jxor g21172(.dina(w_n20706_0[0]),.dinb(w_n4582_20[2]),.dout(n21430),.clk(gclk));
	jand g21173(.dina(n21430),.dinb(w_asqrt6_21[0]),.dout(n21431),.clk(gclk));
	jxor g21174(.dina(n21431),.dinb(w_n20711_0[0]),.dout(n21432),.clk(gclk));
	jand g21175(.dina(w_n21432_0[1]),.dinb(n21429),.dout(n21433),.clk(gclk));
	jor g21176(.dina(n21433),.dinb(w_n21428_0[1]),.dout(n21434),.clk(gclk));
	jand g21177(.dina(w_n21434_0[2]),.dinb(w_asqrt40_15[2]),.dout(n21435),.clk(gclk));
	jor g21178(.dina(w_n21434_0[1]),.dinb(w_asqrt40_15[1]),.dout(n21436),.clk(gclk));
	jxor g21179(.dina(w_n20714_0[0]),.dinb(w_n4249_24[1]),.dout(n21437),.clk(gclk));
	jand g21180(.dina(n21437),.dinb(w_asqrt6_20[2]),.dout(n21438),.clk(gclk));
	jxor g21181(.dina(n21438),.dinb(w_n20719_0[0]),.dout(n21439),.clk(gclk));
	jnot g21182(.din(w_n21439_0[1]),.dout(n21440),.clk(gclk));
	jand g21183(.dina(w_n21440_0[1]),.dinb(n21436),.dout(n21441),.clk(gclk));
	jor g21184(.dina(n21441),.dinb(w_n21435_0[1]),.dout(n21442),.clk(gclk));
	jand g21185(.dina(w_n21442_0[2]),.dinb(w_asqrt41_12[2]),.dout(n21443),.clk(gclk));
	jor g21186(.dina(w_n21442_0[1]),.dinb(w_asqrt41_12[1]),.dout(n21444),.clk(gclk));
	jxor g21187(.dina(w_n20721_0[0]),.dinb(w_n3955_21[1]),.dout(n21445),.clk(gclk));
	jand g21188(.dina(n21445),.dinb(w_asqrt6_20[1]),.dout(n21446),.clk(gclk));
	jxor g21189(.dina(n21446),.dinb(w_n20726_0[0]),.dout(n21447),.clk(gclk));
	jand g21190(.dina(w_n21447_0[1]),.dinb(n21444),.dout(n21448),.clk(gclk));
	jor g21191(.dina(n21448),.dinb(w_n21443_0[1]),.dout(n21449),.clk(gclk));
	jand g21192(.dina(w_n21449_0[2]),.dinb(w_asqrt42_16[0]),.dout(n21450),.clk(gclk));
	jor g21193(.dina(w_n21449_0[1]),.dinb(w_asqrt42_15[2]),.dout(n21451),.clk(gclk));
	jxor g21194(.dina(w_n20729_0[0]),.dinb(w_n3642_24[2]),.dout(n21452),.clk(gclk));
	jand g21195(.dina(n21452),.dinb(w_asqrt6_20[0]),.dout(n21453),.clk(gclk));
	jxor g21196(.dina(n21453),.dinb(w_n20734_0[0]),.dout(n21454),.clk(gclk));
	jnot g21197(.din(w_n21454_0[1]),.dout(n21455),.clk(gclk));
	jand g21198(.dina(w_n21455_0[1]),.dinb(n21451),.dout(n21456),.clk(gclk));
	jor g21199(.dina(n21456),.dinb(w_n21450_0[1]),.dout(n21457),.clk(gclk));
	jand g21200(.dina(w_n21457_0[2]),.dinb(w_asqrt43_13[0]),.dout(n21458),.clk(gclk));
	jor g21201(.dina(w_n21457_0[1]),.dinb(w_asqrt43_12[2]),.dout(n21459),.clk(gclk));
	jxor g21202(.dina(w_n20736_0[0]),.dinb(w_n3368_22[0]),.dout(n21460),.clk(gclk));
	jand g21203(.dina(n21460),.dinb(w_asqrt6_19[2]),.dout(n21461),.clk(gclk));
	jxor g21204(.dina(n21461),.dinb(w_n20741_0[0]),.dout(n21462),.clk(gclk));
	jnot g21205(.din(w_n21462_0[1]),.dout(n21463),.clk(gclk));
	jand g21206(.dina(w_n21463_0[1]),.dinb(n21459),.dout(n21464),.clk(gclk));
	jor g21207(.dina(n21464),.dinb(w_n21458_0[1]),.dout(n21465),.clk(gclk));
	jand g21208(.dina(w_n21465_0[2]),.dinb(w_asqrt44_16[0]),.dout(n21466),.clk(gclk));
	jor g21209(.dina(w_n21465_0[1]),.dinb(w_asqrt44_15[2]),.dout(n21467),.clk(gclk));
	jxor g21210(.dina(w_n20743_0[0]),.dinb(w_n3089_25[1]),.dout(n21468),.clk(gclk));
	jand g21211(.dina(n21468),.dinb(w_asqrt6_19[1]),.dout(n21469),.clk(gclk));
	jxor g21212(.dina(n21469),.dinb(w_n20748_0[0]),.dout(n21470),.clk(gclk));
	jnot g21213(.din(w_n21470_0[1]),.dout(n21471),.clk(gclk));
	jand g21214(.dina(w_n21471_0[1]),.dinb(n21467),.dout(n21472),.clk(gclk));
	jor g21215(.dina(n21472),.dinb(w_n21466_0[1]),.dout(n21473),.clk(gclk));
	jand g21216(.dina(w_n21473_0[2]),.dinb(w_asqrt45_13[2]),.dout(n21474),.clk(gclk));
	jor g21217(.dina(w_n21473_0[1]),.dinb(w_asqrt45_13[1]),.dout(n21475),.clk(gclk));
	jxor g21218(.dina(w_n20750_0[0]),.dinb(w_n2833_23[0]),.dout(n21476),.clk(gclk));
	jand g21219(.dina(n21476),.dinb(w_asqrt6_19[0]),.dout(n21477),.clk(gclk));
	jxor g21220(.dina(n21477),.dinb(w_n20755_0[0]),.dout(n21478),.clk(gclk));
	jand g21221(.dina(w_n21478_0[1]),.dinb(n21475),.dout(n21479),.clk(gclk));
	jor g21222(.dina(n21479),.dinb(w_n21474_0[1]),.dout(n21480),.clk(gclk));
	jand g21223(.dina(w_n21480_0[2]),.dinb(w_asqrt46_16[0]),.dout(n21481),.clk(gclk));
	jor g21224(.dina(w_n21480_0[1]),.dinb(w_asqrt46_15[2]),.dout(n21482),.clk(gclk));
	jxor g21225(.dina(w_n20758_0[0]),.dinb(w_n2572_25[2]),.dout(n21483),.clk(gclk));
	jand g21226(.dina(n21483),.dinb(w_asqrt6_18[2]),.dout(n21484),.clk(gclk));
	jxor g21227(.dina(n21484),.dinb(w_n20763_0[0]),.dout(n21485),.clk(gclk));
	jnot g21228(.din(w_n21485_0[1]),.dout(n21486),.clk(gclk));
	jand g21229(.dina(w_n21486_0[1]),.dinb(n21482),.dout(n21487),.clk(gclk));
	jor g21230(.dina(n21487),.dinb(w_n21481_0[1]),.dout(n21488),.clk(gclk));
	jand g21231(.dina(w_n21488_0[2]),.dinb(w_asqrt47_14[1]),.dout(n21489),.clk(gclk));
	jor g21232(.dina(w_n21488_0[1]),.dinb(w_asqrt47_14[0]),.dout(n21490),.clk(gclk));
	jxor g21233(.dina(w_n20765_0[0]),.dinb(w_n2345_23[2]),.dout(n21491),.clk(gclk));
	jand g21234(.dina(n21491),.dinb(w_asqrt6_18[1]),.dout(n21492),.clk(gclk));
	jxor g21235(.dina(n21492),.dinb(w_n20770_0[0]),.dout(n21493),.clk(gclk));
	jnot g21236(.din(w_n21493_0[1]),.dout(n21494),.clk(gclk));
	jand g21237(.dina(w_n21494_0[1]),.dinb(n21490),.dout(n21495),.clk(gclk));
	jor g21238(.dina(n21495),.dinb(w_n21489_0[1]),.dout(n21496),.clk(gclk));
	jand g21239(.dina(w_n21496_0[2]),.dinb(w_asqrt48_16[1]),.dout(n21497),.clk(gclk));
	jor g21240(.dina(w_n21496_0[1]),.dinb(w_asqrt48_16[0]),.dout(n21498),.clk(gclk));
	jxor g21241(.dina(w_n20772_0[0]),.dinb(w_n2108_26[1]),.dout(n21499),.clk(gclk));
	jand g21242(.dina(n21499),.dinb(w_asqrt6_18[0]),.dout(n21500),.clk(gclk));
	jxor g21243(.dina(n21500),.dinb(w_n20777_0[0]),.dout(n21501),.clk(gclk));
	jnot g21244(.din(w_n21501_0[1]),.dout(n21502),.clk(gclk));
	jand g21245(.dina(w_n21502_0[1]),.dinb(n21498),.dout(n21503),.clk(gclk));
	jor g21246(.dina(n21503),.dinb(w_n21497_0[1]),.dout(n21504),.clk(gclk));
	jand g21247(.dina(w_n21504_0[2]),.dinb(w_asqrt49_14[2]),.dout(n21505),.clk(gclk));
	jor g21248(.dina(w_n21504_0[1]),.dinb(w_asqrt49_14[1]),.dout(n21506),.clk(gclk));
	jxor g21249(.dina(w_n20779_0[0]),.dinb(w_n1912_24[2]),.dout(n21507),.clk(gclk));
	jand g21250(.dina(n21507),.dinb(w_asqrt6_17[2]),.dout(n21508),.clk(gclk));
	jxor g21251(.dina(n21508),.dinb(w_n20784_0[0]),.dout(n21509),.clk(gclk));
	jnot g21252(.din(w_n21509_0[1]),.dout(n21510),.clk(gclk));
	jand g21253(.dina(w_n21510_0[1]),.dinb(n21506),.dout(n21511),.clk(gclk));
	jor g21254(.dina(n21511),.dinb(w_n21505_0[1]),.dout(n21512),.clk(gclk));
	jand g21255(.dina(w_n21512_0[2]),.dinb(w_asqrt50_16[2]),.dout(n21513),.clk(gclk));
	jor g21256(.dina(w_n21512_0[1]),.dinb(w_asqrt50_16[1]),.dout(n21514),.clk(gclk));
	jxor g21257(.dina(w_n20786_0[0]),.dinb(w_n1699_27[0]),.dout(n21515),.clk(gclk));
	jand g21258(.dina(n21515),.dinb(w_asqrt6_17[1]),.dout(n21516),.clk(gclk));
	jxor g21259(.dina(n21516),.dinb(w_n20791_0[0]),.dout(n21517),.clk(gclk));
	jnot g21260(.din(w_n21517_0[1]),.dout(n21518),.clk(gclk));
	jand g21261(.dina(w_n21518_0[1]),.dinb(n21514),.dout(n21519),.clk(gclk));
	jor g21262(.dina(n21519),.dinb(w_n21513_0[1]),.dout(n21520),.clk(gclk));
	jand g21263(.dina(w_n21520_0[2]),.dinb(w_asqrt51_15[0]),.dout(n21521),.clk(gclk));
	jor g21264(.dina(w_n21520_0[1]),.dinb(w_asqrt51_14[2]),.dout(n21522),.clk(gclk));
	jxor g21265(.dina(w_n20793_0[0]),.dinb(w_n1516_25[1]),.dout(n21523),.clk(gclk));
	jand g21266(.dina(n21523),.dinb(w_asqrt6_17[0]),.dout(n21524),.clk(gclk));
	jxor g21267(.dina(n21524),.dinb(w_n20798_0[0]),.dout(n21525),.clk(gclk));
	jand g21268(.dina(w_n21525_0[1]),.dinb(n21522),.dout(n21526),.clk(gclk));
	jor g21269(.dina(n21526),.dinb(w_n21521_0[1]),.dout(n21527),.clk(gclk));
	jand g21270(.dina(w_n21527_0[2]),.dinb(w_asqrt52_16[2]),.dout(n21528),.clk(gclk));
	jor g21271(.dina(w_n21527_0[1]),.dinb(w_asqrt52_16[1]),.dout(n21529),.clk(gclk));
	jxor g21272(.dina(w_n20801_0[0]),.dinb(w_n1332_27[0]),.dout(n21530),.clk(gclk));
	jand g21273(.dina(n21530),.dinb(w_asqrt6_16[2]),.dout(n21531),.clk(gclk));
	jxor g21274(.dina(n21531),.dinb(w_n20806_0[0]),.dout(n21532),.clk(gclk));
	jnot g21275(.din(w_n21532_0[1]),.dout(n21533),.clk(gclk));
	jand g21276(.dina(w_n21533_0[1]),.dinb(n21529),.dout(n21534),.clk(gclk));
	jor g21277(.dina(n21534),.dinb(w_n21528_0[1]),.dout(n21535),.clk(gclk));
	jand g21278(.dina(w_n21535_0[2]),.dinb(w_asqrt53_15[2]),.dout(n21536),.clk(gclk));
	jor g21279(.dina(w_n21535_0[1]),.dinb(w_asqrt53_15[1]),.dout(n21537),.clk(gclk));
	jxor g21280(.dina(w_n20808_0[0]),.dinb(w_n1173_26[0]),.dout(n21538),.clk(gclk));
	jand g21281(.dina(n21538),.dinb(w_asqrt6_16[1]),.dout(n21539),.clk(gclk));
	jxor g21282(.dina(n21539),.dinb(w_n20813_0[0]),.dout(n21540),.clk(gclk));
	jand g21283(.dina(w_n21540_0[1]),.dinb(n21537),.dout(n21541),.clk(gclk));
	jor g21284(.dina(n21541),.dinb(w_n21536_0[1]),.dout(n21542),.clk(gclk));
	jand g21285(.dina(w_n21542_0[2]),.dinb(w_asqrt54_16[2]),.dout(n21543),.clk(gclk));
	jor g21286(.dina(w_n21542_0[1]),.dinb(w_asqrt54_16[1]),.dout(n21544),.clk(gclk));
	jxor g21287(.dina(w_n20816_0[0]),.dinb(w_n1008_28[0]),.dout(n21545),.clk(gclk));
	jand g21288(.dina(n21545),.dinb(w_asqrt6_16[0]),.dout(n21546),.clk(gclk));
	jxor g21289(.dina(n21546),.dinb(w_n20821_0[0]),.dout(n21547),.clk(gclk));
	jnot g21290(.din(w_n21547_0[1]),.dout(n21548),.clk(gclk));
	jand g21291(.dina(w_n21548_0[1]),.dinb(n21544),.dout(n21549),.clk(gclk));
	jor g21292(.dina(n21549),.dinb(w_n21543_0[1]),.dout(n21550),.clk(gclk));
	jand g21293(.dina(w_n21550_0[2]),.dinb(w_asqrt55_16[0]),.dout(n21551),.clk(gclk));
	jor g21294(.dina(w_n21550_0[1]),.dinb(w_asqrt55_15[2]),.dout(n21552),.clk(gclk));
	jxor g21295(.dina(w_n20823_0[0]),.dinb(w_n884_27[0]),.dout(n21553),.clk(gclk));
	jand g21296(.dina(n21553),.dinb(w_asqrt6_15[2]),.dout(n21554),.clk(gclk));
	jxor g21297(.dina(n21554),.dinb(w_n20828_0[0]),.dout(n21555),.clk(gclk));
	jnot g21298(.din(w_n21555_0[1]),.dout(n21556),.clk(gclk));
	jand g21299(.dina(w_n21556_0[1]),.dinb(n21552),.dout(n21557),.clk(gclk));
	jor g21300(.dina(n21557),.dinb(w_n21551_0[1]),.dout(n21558),.clk(gclk));
	jand g21301(.dina(w_n21558_0[2]),.dinb(w_asqrt56_17[0]),.dout(n21559),.clk(gclk));
	jor g21302(.dina(w_n21558_0[1]),.dinb(w_asqrt56_16[2]),.dout(n21560),.clk(gclk));
	jxor g21303(.dina(w_n20830_0[0]),.dinb(w_n743_28[0]),.dout(n21561),.clk(gclk));
	jand g21304(.dina(n21561),.dinb(w_asqrt6_15[1]),.dout(n21562),.clk(gclk));
	jxor g21305(.dina(n21562),.dinb(w_n20835_0[0]),.dout(n21563),.clk(gclk));
	jand g21306(.dina(w_n21563_0[1]),.dinb(n21560),.dout(n21564),.clk(gclk));
	jor g21307(.dina(n21564),.dinb(w_n21559_0[1]),.dout(n21565),.clk(gclk));
	jand g21308(.dina(w_n21565_0[2]),.dinb(w_asqrt57_16[2]),.dout(n21566),.clk(gclk));
	jor g21309(.dina(w_n21565_0[1]),.dinb(w_asqrt57_16[1]),.dout(n21567),.clk(gclk));
	jxor g21310(.dina(w_n20838_0[0]),.dinb(w_n635_28[0]),.dout(n21568),.clk(gclk));
	jand g21311(.dina(n21568),.dinb(w_asqrt6_15[0]),.dout(n21569),.clk(gclk));
	jxor g21312(.dina(n21569),.dinb(w_n20842_0[0]),.dout(n21570),.clk(gclk));
	jand g21313(.dina(w_n21570_0[1]),.dinb(n21567),.dout(n21571),.clk(gclk));
	jor g21314(.dina(n21571),.dinb(w_n21566_0[1]),.dout(n21572),.clk(gclk));
	jand g21315(.dina(w_n21572_0[2]),.dinb(w_asqrt58_17[1]),.dout(n21573),.clk(gclk));
	jor g21316(.dina(w_n21572_0[1]),.dinb(w_asqrt58_17[0]),.dout(n21574),.clk(gclk));
	jxor g21317(.dina(w_n20846_0[0]),.dinb(w_n515_29[0]),.dout(n21575),.clk(gclk));
	jand g21318(.dina(n21575),.dinb(w_asqrt6_14[2]),.dout(n21576),.clk(gclk));
	jxor g21319(.dina(n21576),.dinb(w_n20851_0[0]),.dout(n21577),.clk(gclk));
	jnot g21320(.din(w_n21577_0[1]),.dout(n21578),.clk(gclk));
	jand g21321(.dina(w_n21578_0[1]),.dinb(n21574),.dout(n21579),.clk(gclk));
	jor g21322(.dina(n21579),.dinb(w_n21573_0[1]),.dout(n21580),.clk(gclk));
	jand g21323(.dina(w_n21580_0[2]),.dinb(w_asqrt59_17[0]),.dout(n21581),.clk(gclk));
	jor g21324(.dina(w_n21580_0[1]),.dinb(w_asqrt59_16[2]),.dout(n21582),.clk(gclk));
	jxor g21325(.dina(w_n20853_0[0]),.dinb(w_n443_29[0]),.dout(n21583),.clk(gclk));
	jand g21326(.dina(n21583),.dinb(w_asqrt6_14[1]),.dout(n21584),.clk(gclk));
	jxor g21327(.dina(n21584),.dinb(w_n20859_0[0]),.dout(n21585),.clk(gclk));
	jnot g21328(.din(w_n21585_0[1]),.dout(n21586),.clk(gclk));
	jand g21329(.dina(w_n21586_0[1]),.dinb(n21582),.dout(n21587),.clk(gclk));
	jor g21330(.dina(n21587),.dinb(w_n21581_0[1]),.dout(n21588),.clk(gclk));
	jand g21331(.dina(w_n21588_0[2]),.dinb(w_asqrt60_17[1]),.dout(n21589),.clk(gclk));
	jor g21332(.dina(w_n21588_0[1]),.dinb(w_asqrt60_17[0]),.dout(n21590),.clk(gclk));
	jxor g21333(.dina(w_n20861_0[0]),.dinb(w_n352_29[1]),.dout(n21591),.clk(gclk));
	jand g21334(.dina(n21591),.dinb(w_asqrt6_14[0]),.dout(n21592),.clk(gclk));
	jxor g21335(.dina(n21592),.dinb(w_n20866_0[0]),.dout(n21593),.clk(gclk));
	jnot g21336(.din(w_n21593_0[1]),.dout(n21594),.clk(gclk));
	jand g21337(.dina(w_n21594_0[1]),.dinb(n21590),.dout(n21595),.clk(gclk));
	jor g21338(.dina(n21595),.dinb(w_n21589_0[1]),.dout(n21596),.clk(gclk));
	jand g21339(.dina(w_n21596_0[2]),.dinb(w_asqrt61_17[1]),.dout(n21597),.clk(gclk));
	jor g21340(.dina(w_n21596_0[1]),.dinb(w_asqrt61_17[0]),.dout(n21598),.clk(gclk));
	jxor g21341(.dina(w_n20868_0[0]),.dinb(w_n294_29[2]),.dout(n21599),.clk(gclk));
	jand g21342(.dina(n21599),.dinb(w_asqrt6_13[2]),.dout(n21600),.clk(gclk));
	jxor g21343(.dina(n21600),.dinb(w_n20873_0[0]),.dout(n21601),.clk(gclk));
	jnot g21344(.din(w_n21601_0[2]),.dout(n21602),.clk(gclk));
	jand g21345(.dina(n21602),.dinb(n21598),.dout(n21603),.clk(gclk));
	jor g21346(.dina(n21603),.dinb(w_n21597_0[1]),.dout(n21604),.clk(gclk));
	jand g21347(.dina(w_n21604_0[2]),.dinb(w_asqrt62_17[1]),.dout(n21605),.clk(gclk));
	jor g21348(.dina(w_n21604_0[1]),.dinb(w_asqrt62_17[0]),.dout(n21606),.clk(gclk));
	jxor g21349(.dina(w_n20875_0[0]),.dinb(w_n239_29[2]),.dout(n21607),.clk(gclk));
	jand g21350(.dina(n21607),.dinb(w_asqrt6_13[1]),.dout(n21608),.clk(gclk));
	jxor g21351(.dina(n21608),.dinb(w_n20880_0[0]),.dout(n21609),.clk(gclk));
	jand g21352(.dina(w_n21609_0[2]),.dinb(n21606),.dout(n21610),.clk(gclk));
	jor g21353(.dina(n21610),.dinb(w_n21605_0[1]),.dout(n21611),.clk(gclk));
	jxor g21354(.dina(w_n20883_0[0]),.dinb(w_n221_30[0]),.dout(n21612),.clk(gclk));
	jand g21355(.dina(n21612),.dinb(w_asqrt6_13[0]),.dout(n21613),.clk(gclk));
	jxor g21356(.dina(n21613),.dinb(w_n20888_0[0]),.dout(n21614),.clk(gclk));
	jnot g21357(.din(w_n21614_0[1]),.dout(n21615),.clk(gclk));
	jor g21358(.dina(w_n21615_0[2]),.dinb(w_n21611_0[2]),.dout(n21616),.clk(gclk));
	jnot g21359(.din(w_n21616_0[1]),.dout(n21617),.clk(gclk));
	jand g21360(.dina(w_asqrt6_12[2]),.dinb(w_n21176_0[0]),.dout(n21618),.clk(gclk));
	jnot g21361(.din(w_n21605_0[0]),.dout(n21619),.clk(gclk));
	jnot g21362(.din(w_n21597_0[0]),.dout(n21620),.clk(gclk));
	jnot g21363(.din(w_n21589_0[0]),.dout(n21621),.clk(gclk));
	jnot g21364(.din(w_n21581_0[0]),.dout(n21622),.clk(gclk));
	jnot g21365(.din(w_n21573_0[0]),.dout(n21623),.clk(gclk));
	jnot g21366(.din(w_n21566_0[0]),.dout(n21624),.clk(gclk));
	jnot g21367(.din(w_n21559_0[0]),.dout(n21625),.clk(gclk));
	jnot g21368(.din(w_n21551_0[0]),.dout(n21626),.clk(gclk));
	jnot g21369(.din(w_n21543_0[0]),.dout(n21627),.clk(gclk));
	jnot g21370(.din(w_n21536_0[0]),.dout(n21628),.clk(gclk));
	jnot g21371(.din(w_n21528_0[0]),.dout(n21629),.clk(gclk));
	jnot g21372(.din(w_n21521_0[0]),.dout(n21630),.clk(gclk));
	jnot g21373(.din(w_n21513_0[0]),.dout(n21631),.clk(gclk));
	jnot g21374(.din(w_n21505_0[0]),.dout(n21632),.clk(gclk));
	jnot g21375(.din(w_n21497_0[0]),.dout(n21633),.clk(gclk));
	jnot g21376(.din(w_n21489_0[0]),.dout(n21634),.clk(gclk));
	jnot g21377(.din(w_n21481_0[0]),.dout(n21635),.clk(gclk));
	jnot g21378(.din(w_n21474_0[0]),.dout(n21636),.clk(gclk));
	jnot g21379(.din(w_n21466_0[0]),.dout(n21637),.clk(gclk));
	jnot g21380(.din(w_n21458_0[0]),.dout(n21638),.clk(gclk));
	jnot g21381(.din(w_n21450_0[0]),.dout(n21639),.clk(gclk));
	jnot g21382(.din(w_n21443_0[0]),.dout(n21640),.clk(gclk));
	jnot g21383(.din(w_n21435_0[0]),.dout(n21641),.clk(gclk));
	jnot g21384(.din(w_n21428_0[0]),.dout(n21642),.clk(gclk));
	jnot g21385(.din(w_n21420_0[0]),.dout(n21643),.clk(gclk));
	jnot g21386(.din(w_n21413_0[0]),.dout(n21644),.clk(gclk));
	jnot g21387(.din(w_n21405_0[0]),.dout(n21645),.clk(gclk));
	jnot g21388(.din(w_n21398_0[0]),.dout(n21646),.clk(gclk));
	jnot g21389(.din(w_n21390_0[0]),.dout(n21647),.clk(gclk));
	jnot g21390(.din(w_n21382_0[0]),.dout(n21648),.clk(gclk));
	jnot g21391(.din(w_n21374_0[0]),.dout(n21649),.clk(gclk));
	jnot g21392(.din(w_n21367_0[0]),.dout(n21650),.clk(gclk));
	jnot g21393(.din(w_n21359_0[0]),.dout(n21651),.clk(gclk));
	jnot g21394(.din(w_n21352_0[0]),.dout(n21652),.clk(gclk));
	jnot g21395(.din(w_n21344_0[0]),.dout(n21653),.clk(gclk));
	jnot g21396(.din(w_n21337_0[0]),.dout(n21654),.clk(gclk));
	jnot g21397(.din(w_n21330_0[0]),.dout(n21655),.clk(gclk));
	jnot g21398(.din(w_n21322_0[0]),.dout(n21656),.clk(gclk));
	jnot g21399(.din(w_n21314_0[0]),.dout(n21657),.clk(gclk));
	jnot g21400(.din(w_n21307_0[0]),.dout(n21658),.clk(gclk));
	jnot g21401(.din(w_n21299_0[0]),.dout(n21659),.clk(gclk));
	jnot g21402(.din(w_n21292_0[0]),.dout(n21660),.clk(gclk));
	jnot g21403(.din(w_n21284_0[0]),.dout(n21661),.clk(gclk));
	jnot g21404(.din(w_n21277_0[0]),.dout(n21662),.clk(gclk));
	jnot g21405(.din(w_n21269_0[0]),.dout(n21663),.clk(gclk));
	jnot g21406(.din(w_n21261_0[0]),.dout(n21664),.clk(gclk));
	jnot g21407(.din(w_n21253_0[0]),.dout(n21665),.clk(gclk));
	jnot g21408(.din(w_n21246_0[0]),.dout(n21666),.clk(gclk));
	jnot g21409(.din(w_n21238_0[0]),.dout(n21667),.clk(gclk));
	jnot g21410(.din(w_n21230_0[0]),.dout(n21668),.clk(gclk));
	jnot g21411(.din(w_n21222_0[0]),.dout(n21669),.clk(gclk));
	jnot g21412(.din(w_n21215_0[0]),.dout(n21670),.clk(gclk));
	jnot g21413(.din(w_n21207_0[0]),.dout(n21671),.clk(gclk));
	jnot g21414(.din(w_n21200_0[0]),.dout(n21672),.clk(gclk));
	jnot g21415(.din(w_n21189_0[0]),.dout(n21673),.clk(gclk));
	jnot g21416(.din(w_n20913_0[0]),.dout(n21674),.clk(gclk));
	jnot g21417(.din(w_n20910_0[0]),.dout(n21675),.clk(gclk));
	jor g21418(.dina(w_n21184_7[1]),.dinb(w_n20473_0[2]),.dout(n21676),.clk(gclk));
	jand g21419(.dina(n21676),.dinb(n21675),.dout(n21677),.clk(gclk));
	jand g21420(.dina(n21677),.dinb(w_n20468_16[0]),.dout(n21678),.clk(gclk));
	jor g21421(.dina(w_n21184_7[0]),.dinb(w_a12_0[0]),.dout(n21679),.clk(gclk));
	jand g21422(.dina(n21679),.dinb(w_a13_0[0]),.dout(n21680),.clk(gclk));
	jor g21423(.dina(w_n21191_0[0]),.dinb(n21680),.dout(n21681),.clk(gclk));
	jor g21424(.dina(w_n21681_0[1]),.dinb(n21678),.dout(n21682),.clk(gclk));
	jand g21425(.dina(n21682),.dinb(n21674),.dout(n21683),.clk(gclk));
	jand g21426(.dina(n21683),.dinb(w_n19791_7[2]),.dout(n21684),.clk(gclk));
	jor g21427(.dina(w_n21196_0[0]),.dinb(n21684),.dout(n21685),.clk(gclk));
	jand g21428(.dina(n21685),.dinb(n21673),.dout(n21686),.clk(gclk));
	jand g21429(.dina(n21686),.dinb(w_n19096_16[1]),.dout(n21687),.clk(gclk));
	jnot g21430(.din(w_n21204_0[0]),.dout(n21688),.clk(gclk));
	jor g21431(.dina(w_n21688_0[1]),.dinb(n21687),.dout(n21689),.clk(gclk));
	jand g21432(.dina(n21689),.dinb(n21672),.dout(n21690),.clk(gclk));
	jand g21433(.dina(n21690),.dinb(w_n18442_8[1]),.dout(n21691),.clk(gclk));
	jor g21434(.dina(w_n21211_0[0]),.dinb(n21691),.dout(n21692),.clk(gclk));
	jand g21435(.dina(n21692),.dinb(n21671),.dout(n21693),.clk(gclk));
	jand g21436(.dina(n21693),.dinb(w_n17769_17[0]),.dout(n21694),.clk(gclk));
	jnot g21437(.din(w_n21219_0[0]),.dout(n21695),.clk(gclk));
	jor g21438(.dina(w_n21695_0[1]),.dinb(n21694),.dout(n21696),.clk(gclk));
	jand g21439(.dina(n21696),.dinb(n21670),.dout(n21697),.clk(gclk));
	jand g21440(.dina(n21697),.dinb(w_n17134_9[1]),.dout(n21698),.clk(gclk));
	jor g21441(.dina(w_n21226_0[0]),.dinb(n21698),.dout(n21699),.clk(gclk));
	jand g21442(.dina(n21699),.dinb(n21669),.dout(n21700),.clk(gclk));
	jand g21443(.dina(n21700),.dinb(w_n16489_17[1]),.dout(n21701),.clk(gclk));
	jor g21444(.dina(w_n21234_0[0]),.dinb(n21701),.dout(n21702),.clk(gclk));
	jand g21445(.dina(n21702),.dinb(n21668),.dout(n21703),.clk(gclk));
	jand g21446(.dina(n21703),.dinb(w_n15878_10[1]),.dout(n21704),.clk(gclk));
	jor g21447(.dina(w_n21242_0[0]),.dinb(n21704),.dout(n21705),.clk(gclk));
	jand g21448(.dina(n21705),.dinb(n21667),.dout(n21706),.clk(gclk));
	jand g21449(.dina(n21706),.dinb(w_n15260_18[0]),.dout(n21707),.clk(gclk));
	jnot g21450(.din(w_n21250_0[0]),.dout(n21708),.clk(gclk));
	jor g21451(.dina(w_n21708_0[1]),.dinb(n21707),.dout(n21709),.clk(gclk));
	jand g21452(.dina(n21709),.dinb(n21666),.dout(n21710),.clk(gclk));
	jand g21453(.dina(n21710),.dinb(w_n14674_11[0]),.dout(n21711),.clk(gclk));
	jor g21454(.dina(w_n21257_0[0]),.dinb(n21711),.dout(n21712),.clk(gclk));
	jand g21455(.dina(n21712),.dinb(n21665),.dout(n21713),.clk(gclk));
	jand g21456(.dina(n21713),.dinb(w_n14078_18[1]),.dout(n21714),.clk(gclk));
	jor g21457(.dina(w_n21265_0[0]),.dinb(n21714),.dout(n21715),.clk(gclk));
	jand g21458(.dina(n21715),.dinb(n21664),.dout(n21716),.clk(gclk));
	jand g21459(.dina(n21716),.dinb(w_n13515_12[0]),.dout(n21717),.clk(gclk));
	jor g21460(.dina(w_n21273_0[0]),.dinb(n21717),.dout(n21718),.clk(gclk));
	jand g21461(.dina(n21718),.dinb(n21663),.dout(n21719),.clk(gclk));
	jand g21462(.dina(n21719),.dinb(w_n12947_19[0]),.dout(n21720),.clk(gclk));
	jnot g21463(.din(w_n21281_0[0]),.dout(n21721),.clk(gclk));
	jor g21464(.dina(w_n21721_0[1]),.dinb(n21720),.dout(n21722),.clk(gclk));
	jand g21465(.dina(n21722),.dinb(n21662),.dout(n21723),.clk(gclk));
	jand g21466(.dina(n21723),.dinb(w_n12410_12[2]),.dout(n21724),.clk(gclk));
	jor g21467(.dina(w_n21288_0[0]),.dinb(n21724),.dout(n21725),.clk(gclk));
	jand g21468(.dina(n21725),.dinb(n21661),.dout(n21726),.clk(gclk));
	jand g21469(.dina(n21726),.dinb(w_n11858_19[1]),.dout(n21727),.clk(gclk));
	jnot g21470(.din(w_n21296_0[0]),.dout(n21728),.clk(gclk));
	jor g21471(.dina(w_n21728_0[1]),.dinb(n21727),.dout(n21729),.clk(gclk));
	jand g21472(.dina(n21729),.dinb(n21660),.dout(n21730),.clk(gclk));
	jand g21473(.dina(n21730),.dinb(w_n11347_13[1]),.dout(n21731),.clk(gclk));
	jor g21474(.dina(w_n21303_0[0]),.dinb(n21731),.dout(n21732),.clk(gclk));
	jand g21475(.dina(n21732),.dinb(n21659),.dout(n21733),.clk(gclk));
	jand g21476(.dina(n21733),.dinb(w_n10824_20[0]),.dout(n21734),.clk(gclk));
	jnot g21477(.din(w_n21311_0[0]),.dout(n21735),.clk(gclk));
	jor g21478(.dina(w_n21735_0[1]),.dinb(n21734),.dout(n21736),.clk(gclk));
	jand g21479(.dina(n21736),.dinb(n21658),.dout(n21737),.clk(gclk));
	jand g21480(.dina(n21737),.dinb(w_n10328_14[1]),.dout(n21738),.clk(gclk));
	jor g21481(.dina(w_n21318_0[0]),.dinb(n21738),.dout(n21739),.clk(gclk));
	jand g21482(.dina(n21739),.dinb(n21657),.dout(n21740),.clk(gclk));
	jand g21483(.dina(n21740),.dinb(w_n9832_20[2]),.dout(n21741),.clk(gclk));
	jor g21484(.dina(w_n21326_0[0]),.dinb(n21741),.dout(n21742),.clk(gclk));
	jand g21485(.dina(n21742),.dinb(n21656),.dout(n21743),.clk(gclk));
	jand g21486(.dina(n21743),.dinb(w_n9369_15[1]),.dout(n21744),.clk(gclk));
	jnot g21487(.din(w_n21334_0[0]),.dout(n21745),.clk(gclk));
	jor g21488(.dina(w_n21745_0[1]),.dinb(n21744),.dout(n21746),.clk(gclk));
	jand g21489(.dina(n21746),.dinb(n21655),.dout(n21747),.clk(gclk));
	jand g21490(.dina(n21747),.dinb(w_n8890_21[0]),.dout(n21748),.clk(gclk));
	jnot g21491(.din(w_n21341_0[0]),.dout(n21749),.clk(gclk));
	jor g21492(.dina(w_n21749_0[1]),.dinb(n21748),.dout(n21750),.clk(gclk));
	jand g21493(.dina(n21750),.dinb(n21654),.dout(n21751),.clk(gclk));
	jand g21494(.dina(n21751),.dinb(w_n8449_16[0]),.dout(n21752),.clk(gclk));
	jor g21495(.dina(w_n21348_0[0]),.dinb(n21752),.dout(n21753),.clk(gclk));
	jand g21496(.dina(n21753),.dinb(n21653),.dout(n21754),.clk(gclk));
	jand g21497(.dina(n21754),.dinb(w_n8003_21[2]),.dout(n21755),.clk(gclk));
	jnot g21498(.din(w_n21356_0[0]),.dout(n21756),.clk(gclk));
	jor g21499(.dina(w_n21756_0[1]),.dinb(n21755),.dout(n21757),.clk(gclk));
	jand g21500(.dina(n21757),.dinb(n21652),.dout(n21758),.clk(gclk));
	jand g21501(.dina(n21758),.dinb(w_n7581_17[0]),.dout(n21759),.clk(gclk));
	jor g21502(.dina(w_n21363_0[0]),.dinb(n21759),.dout(n21760),.clk(gclk));
	jand g21503(.dina(n21760),.dinb(n21651),.dout(n21761),.clk(gclk));
	jand g21504(.dina(n21761),.dinb(w_n7154_22[0]),.dout(n21762),.clk(gclk));
	jnot g21505(.din(w_n21371_0[0]),.dout(n21763),.clk(gclk));
	jor g21506(.dina(w_n21763_0[1]),.dinb(n21762),.dout(n21764),.clk(gclk));
	jand g21507(.dina(n21764),.dinb(n21650),.dout(n21765),.clk(gclk));
	jand g21508(.dina(n21765),.dinb(w_n6758_17[2]),.dout(n21766),.clk(gclk));
	jor g21509(.dina(w_n21378_0[0]),.dinb(n21766),.dout(n21767),.clk(gclk));
	jand g21510(.dina(n21767),.dinb(n21649),.dout(n21768),.clk(gclk));
	jand g21511(.dina(n21768),.dinb(w_n6357_22[1]),.dout(n21769),.clk(gclk));
	jor g21512(.dina(w_n21386_0[0]),.dinb(n21769),.dout(n21770),.clk(gclk));
	jand g21513(.dina(n21770),.dinb(n21648),.dout(n21771),.clk(gclk));
	jand g21514(.dina(n21771),.dinb(w_n5989_18[1]),.dout(n21772),.clk(gclk));
	jor g21515(.dina(w_n21394_0[0]),.dinb(n21772),.dout(n21773),.clk(gclk));
	jand g21516(.dina(n21773),.dinb(n21647),.dout(n21774),.clk(gclk));
	jand g21517(.dina(n21774),.dinb(w_n5606_22[2]),.dout(n21775),.clk(gclk));
	jnot g21518(.din(w_n21402_0[0]),.dout(n21776),.clk(gclk));
	jor g21519(.dina(w_n21776_0[1]),.dinb(n21775),.dout(n21777),.clk(gclk));
	jand g21520(.dina(n21777),.dinb(n21646),.dout(n21778),.clk(gclk));
	jand g21521(.dina(n21778),.dinb(w_n5259_19[1]),.dout(n21779),.clk(gclk));
	jor g21522(.dina(w_n21409_0[0]),.dinb(n21779),.dout(n21780),.clk(gclk));
	jand g21523(.dina(n21780),.dinb(n21645),.dout(n21781),.clk(gclk));
	jand g21524(.dina(n21781),.dinb(w_n4902_23[1]),.dout(n21782),.clk(gclk));
	jnot g21525(.din(w_n21417_0[0]),.dout(n21783),.clk(gclk));
	jor g21526(.dina(w_n21783_0[1]),.dinb(n21782),.dout(n21784),.clk(gclk));
	jand g21527(.dina(n21784),.dinb(n21644),.dout(n21785),.clk(gclk));
	jand g21528(.dina(n21785),.dinb(w_n4582_20[1]),.dout(n21786),.clk(gclk));
	jor g21529(.dina(w_n21424_0[0]),.dinb(n21786),.dout(n21787),.clk(gclk));
	jand g21530(.dina(n21787),.dinb(n21643),.dout(n21788),.clk(gclk));
	jand g21531(.dina(n21788),.dinb(w_n4249_24[0]),.dout(n21789),.clk(gclk));
	jnot g21532(.din(w_n21432_0[0]),.dout(n21790),.clk(gclk));
	jor g21533(.dina(w_n21790_0[1]),.dinb(n21789),.dout(n21791),.clk(gclk));
	jand g21534(.dina(n21791),.dinb(n21642),.dout(n21792),.clk(gclk));
	jand g21535(.dina(n21792),.dinb(w_n3955_21[0]),.dout(n21793),.clk(gclk));
	jor g21536(.dina(w_n21439_0[0]),.dinb(n21793),.dout(n21794),.clk(gclk));
	jand g21537(.dina(n21794),.dinb(n21641),.dout(n21795),.clk(gclk));
	jand g21538(.dina(n21795),.dinb(w_n3642_24[1]),.dout(n21796),.clk(gclk));
	jnot g21539(.din(w_n21447_0[0]),.dout(n21797),.clk(gclk));
	jor g21540(.dina(w_n21797_0[1]),.dinb(n21796),.dout(n21798),.clk(gclk));
	jand g21541(.dina(n21798),.dinb(n21640),.dout(n21799),.clk(gclk));
	jand g21542(.dina(n21799),.dinb(w_n3368_21[2]),.dout(n21800),.clk(gclk));
	jor g21543(.dina(w_n21454_0[0]),.dinb(n21800),.dout(n21801),.clk(gclk));
	jand g21544(.dina(n21801),.dinb(n21639),.dout(n21802),.clk(gclk));
	jand g21545(.dina(n21802),.dinb(w_n3089_25[0]),.dout(n21803),.clk(gclk));
	jor g21546(.dina(w_n21462_0[0]),.dinb(n21803),.dout(n21804),.clk(gclk));
	jand g21547(.dina(n21804),.dinb(n21638),.dout(n21805),.clk(gclk));
	jand g21548(.dina(n21805),.dinb(w_n2833_22[2]),.dout(n21806),.clk(gclk));
	jor g21549(.dina(w_n21470_0[0]),.dinb(n21806),.dout(n21807),.clk(gclk));
	jand g21550(.dina(n21807),.dinb(n21637),.dout(n21808),.clk(gclk));
	jand g21551(.dina(n21808),.dinb(w_n2572_25[1]),.dout(n21809),.clk(gclk));
	jnot g21552(.din(w_n21478_0[0]),.dout(n21810),.clk(gclk));
	jor g21553(.dina(w_n21810_0[1]),.dinb(n21809),.dout(n21811),.clk(gclk));
	jand g21554(.dina(n21811),.dinb(n21636),.dout(n21812),.clk(gclk));
	jand g21555(.dina(n21812),.dinb(w_n2345_23[1]),.dout(n21813),.clk(gclk));
	jor g21556(.dina(w_n21485_0[0]),.dinb(n21813),.dout(n21814),.clk(gclk));
	jand g21557(.dina(n21814),.dinb(n21635),.dout(n21815),.clk(gclk));
	jand g21558(.dina(n21815),.dinb(w_n2108_26[0]),.dout(n21816),.clk(gclk));
	jor g21559(.dina(w_n21493_0[0]),.dinb(n21816),.dout(n21817),.clk(gclk));
	jand g21560(.dina(n21817),.dinb(n21634),.dout(n21818),.clk(gclk));
	jand g21561(.dina(n21818),.dinb(w_n1912_24[1]),.dout(n21819),.clk(gclk));
	jor g21562(.dina(w_n21501_0[0]),.dinb(n21819),.dout(n21820),.clk(gclk));
	jand g21563(.dina(n21820),.dinb(n21633),.dout(n21821),.clk(gclk));
	jand g21564(.dina(n21821),.dinb(w_n1699_26[2]),.dout(n21822),.clk(gclk));
	jor g21565(.dina(w_n21509_0[0]),.dinb(n21822),.dout(n21823),.clk(gclk));
	jand g21566(.dina(n21823),.dinb(n21632),.dout(n21824),.clk(gclk));
	jand g21567(.dina(n21824),.dinb(w_n1516_25[0]),.dout(n21825),.clk(gclk));
	jor g21568(.dina(w_n21517_0[0]),.dinb(n21825),.dout(n21826),.clk(gclk));
	jand g21569(.dina(n21826),.dinb(n21631),.dout(n21827),.clk(gclk));
	jand g21570(.dina(n21827),.dinb(w_n1332_26[2]),.dout(n21828),.clk(gclk));
	jnot g21571(.din(w_n21525_0[0]),.dout(n21829),.clk(gclk));
	jor g21572(.dina(w_n21829_0[1]),.dinb(n21828),.dout(n21830),.clk(gclk));
	jand g21573(.dina(n21830),.dinb(n21630),.dout(n21831),.clk(gclk));
	jand g21574(.dina(n21831),.dinb(w_n1173_25[2]),.dout(n21832),.clk(gclk));
	jor g21575(.dina(w_n21532_0[0]),.dinb(n21832),.dout(n21833),.clk(gclk));
	jand g21576(.dina(n21833),.dinb(n21629),.dout(n21834),.clk(gclk));
	jand g21577(.dina(n21834),.dinb(w_n1008_27[2]),.dout(n21835),.clk(gclk));
	jnot g21578(.din(w_n21540_0[0]),.dout(n21836),.clk(gclk));
	jor g21579(.dina(w_n21836_0[1]),.dinb(n21835),.dout(n21837),.clk(gclk));
	jand g21580(.dina(n21837),.dinb(n21628),.dout(n21838),.clk(gclk));
	jand g21581(.dina(n21838),.dinb(w_n884_26[2]),.dout(n21839),.clk(gclk));
	jor g21582(.dina(w_n21547_0[0]),.dinb(n21839),.dout(n21840),.clk(gclk));
	jand g21583(.dina(n21840),.dinb(n21627),.dout(n21841),.clk(gclk));
	jand g21584(.dina(n21841),.dinb(w_n743_27[2]),.dout(n21842),.clk(gclk));
	jor g21585(.dina(w_n21555_0[0]),.dinb(n21842),.dout(n21843),.clk(gclk));
	jand g21586(.dina(n21843),.dinb(n21626),.dout(n21844),.clk(gclk));
	jand g21587(.dina(n21844),.dinb(w_n635_27[2]),.dout(n21845),.clk(gclk));
	jnot g21588(.din(w_n21563_0[0]),.dout(n21846),.clk(gclk));
	jor g21589(.dina(w_n21846_0[1]),.dinb(n21845),.dout(n21847),.clk(gclk));
	jand g21590(.dina(n21847),.dinb(n21625),.dout(n21848),.clk(gclk));
	jand g21591(.dina(n21848),.dinb(w_n515_28[2]),.dout(n21849),.clk(gclk));
	jnot g21592(.din(w_n21570_0[0]),.dout(n21850),.clk(gclk));
	jor g21593(.dina(w_n21850_0[1]),.dinb(n21849),.dout(n21851),.clk(gclk));
	jand g21594(.dina(n21851),.dinb(n21624),.dout(n21852),.clk(gclk));
	jand g21595(.dina(n21852),.dinb(w_n443_28[2]),.dout(n21853),.clk(gclk));
	jor g21596(.dina(w_n21577_0[0]),.dinb(n21853),.dout(n21854),.clk(gclk));
	jand g21597(.dina(n21854),.dinb(n21623),.dout(n21855),.clk(gclk));
	jand g21598(.dina(n21855),.dinb(w_n352_29[0]),.dout(n21856),.clk(gclk));
	jor g21599(.dina(w_n21585_0[0]),.dinb(n21856),.dout(n21857),.clk(gclk));
	jand g21600(.dina(n21857),.dinb(n21622),.dout(n21858),.clk(gclk));
	jand g21601(.dina(n21858),.dinb(w_n294_29[1]),.dout(n21859),.clk(gclk));
	jor g21602(.dina(w_n21593_0[0]),.dinb(n21859),.dout(n21860),.clk(gclk));
	jand g21603(.dina(n21860),.dinb(n21621),.dout(n21861),.clk(gclk));
	jand g21604(.dina(n21861),.dinb(w_n239_29[1]),.dout(n21862),.clk(gclk));
	jor g21605(.dina(w_n21601_0[1]),.dinb(n21862),.dout(n21863),.clk(gclk));
	jand g21606(.dina(n21863),.dinb(n21620),.dout(n21864),.clk(gclk));
	jand g21607(.dina(n21864),.dinb(w_n221_29[2]),.dout(n21865),.clk(gclk));
	jnot g21608(.din(w_n21609_0[1]),.dout(n21866),.clk(gclk));
	jor g21609(.dina(n21866),.dinb(n21865),.dout(n21867),.clk(gclk));
	jand g21610(.dina(n21867),.dinb(n21619),.dout(n21868),.clk(gclk));
	jor g21611(.dina(w_n21614_0[0]),.dinb(w_n21868_0[1]),.dout(n21869),.clk(gclk));
	jor g21612(.dina(n21869),.dinb(w_n20897_0[0]),.dout(n21870),.clk(gclk));
	jor g21613(.dina(n21870),.dinb(w_n21618_0[1]),.dout(n21871),.clk(gclk));
	jand g21614(.dina(n21871),.dinb(w_n218_12[2]),.dout(n21872),.clk(gclk));
	jand g21615(.dina(w_n21184_6[2]),.dinb(w_n20890_0[0]),.dout(n21873),.clk(gclk));
	jnot g21616(.din(n21873),.dout(n21874),.clk(gclk));
	jand g21617(.dina(w_n20891_0[0]),.dinb(w_asqrt63_21[1]),.dout(n21875),.clk(gclk));
	jand g21618(.dina(n21875),.dinb(w_n21181_0[2]),.dout(n21876),.clk(gclk));
	jand g21619(.dina(n21876),.dinb(n21874),.dout(n21877),.clk(gclk));
	jor g21620(.dina(w_n21877_0[1]),.dinb(n21872),.dout(n21878),.clk(gclk));
	jor g21621(.dina(n21878),.dinb(n21617),.dout(asqrt_fa_6),.clk(gclk));
	jnot g21622(.din(w_n21618_0[0]),.dout(n21880),.clk(gclk));
	jand g21623(.dina(w_n21615_0[1]),.dinb(w_n21611_0[1]),.dout(n21881),.clk(gclk));
	jand g21624(.dina(n21881),.dinb(w_n21181_0[1]),.dout(n21882),.clk(gclk));
	jand g21625(.dina(n21882),.dinb(n21880),.dout(n21883),.clk(gclk));
	jor g21626(.dina(n21883),.dinb(w_asqrt63_21[0]),.dout(n21884),.clk(gclk));
	jnot g21627(.din(w_n21877_0[0]),.dout(n21885),.clk(gclk));
	jand g21628(.dina(n21885),.dinb(n21884),.dout(n21886),.clk(gclk));
	jand g21629(.dina(n21886),.dinb(w_n21616_0[0]),.dout(n21887),.clk(gclk));
	jor g21630(.dina(w_n21887_34[1]),.dinb(w_n20907_1[1]),.dout(n21888),.clk(gclk));
	jnot g21631(.din(w_a8_0[2]),.dout(n21889),.clk(gclk));
	jnot g21632(.din(w_a9_0[1]),.dout(n21890),.clk(gclk));
	jand g21633(.dina(w_n21890_0[1]),.dinb(w_n21889_1[2]),.dout(n21891),.clk(gclk));
	jand g21634(.dina(w_n21891_0[2]),.dinb(w_n20907_1[0]),.dout(n21892),.clk(gclk));
	jnot g21635(.din(w_n21892_0[1]),.dout(n21893),.clk(gclk));
	jand g21636(.dina(n21893),.dinb(n21888),.dout(n21894),.clk(gclk));
	jor g21637(.dina(w_n21894_0[2]),.dinb(w_n21184_6[1]),.dout(n21895),.clk(gclk));
	jand g21638(.dina(w_n21894_0[1]),.dinb(w_n21184_6[0]),.dout(n21896),.clk(gclk));
	jor g21639(.dina(w_n21887_34[0]),.dinb(w_a10_0[1]),.dout(n21897),.clk(gclk));
	jand g21640(.dina(n21897),.dinb(w_a11_0[0]),.dout(n21898),.clk(gclk));
	jand g21641(.dina(w_asqrt5_4[1]),.dinb(w_n20909_0[1]),.dout(n21899),.clk(gclk));
	jor g21642(.dina(n21899),.dinb(n21898),.dout(n21900),.clk(gclk));
	jor g21643(.dina(n21900),.dinb(n21896),.dout(n21901),.clk(gclk));
	jand g21644(.dina(n21901),.dinb(w_n21895_0[1]),.dout(n21902),.clk(gclk));
	jor g21645(.dina(w_n21902_0[2]),.dinb(w_n20468_15[2]),.dout(n21903),.clk(gclk));
	jand g21646(.dina(w_n21902_0[1]),.dinb(w_n20468_15[1]),.dout(n21904),.clk(gclk));
	jnot g21647(.din(w_n20909_0[0]),.dout(n21905),.clk(gclk));
	jor g21648(.dina(w_n21887_33[2]),.dinb(n21905),.dout(n21906),.clk(gclk));
	jor g21649(.dina(w_asqrt5_4[0]),.dinb(w_n21184_5[2]),.dout(n21907),.clk(gclk));
	jand g21650(.dina(n21907),.dinb(w_n21906_0[1]),.dout(n21908),.clk(gclk));
	jxor g21651(.dina(n21908),.dinb(w_n20473_0[1]),.dout(n21909),.clk(gclk));
	jor g21652(.dina(w_n21909_0[1]),.dinb(n21904),.dout(n21910),.clk(gclk));
	jand g21653(.dina(n21910),.dinb(w_n21903_0[1]),.dout(n21911),.clk(gclk));
	jor g21654(.dina(w_n21911_0[2]),.dinb(w_n19791_7[1]),.dout(n21912),.clk(gclk));
	jand g21655(.dina(w_n21911_0[1]),.dinb(w_n19791_7[0]),.dout(n21913),.clk(gclk));
	jxor g21656(.dina(w_n20912_0[0]),.dinb(w_n20468_15[0]),.dout(n21914),.clk(gclk));
	jor g21657(.dina(n21914),.dinb(w_n21887_33[1]),.dout(n21915),.clk(gclk));
	jxor g21658(.dina(n21915),.dinb(w_n21681_0[0]),.dout(n21916),.clk(gclk));
	jnot g21659(.din(w_n21916_0[2]),.dout(n21917),.clk(gclk));
	jor g21660(.dina(n21917),.dinb(n21913),.dout(n21918),.clk(gclk));
	jand g21661(.dina(n21918),.dinb(w_n21912_0[1]),.dout(n21919),.clk(gclk));
	jor g21662(.dina(w_n21919_0[2]),.dinb(w_n19096_16[0]),.dout(n21920),.clk(gclk));
	jand g21663(.dina(w_n21919_0[1]),.dinb(w_n19096_15[2]),.dout(n21921),.clk(gclk));
	jxor g21664(.dina(w_n21188_0[0]),.dinb(w_n19791_6[2]),.dout(n21922),.clk(gclk));
	jor g21665(.dina(n21922),.dinb(w_n21887_33[0]),.dout(n21923),.clk(gclk));
	jxor g21666(.dina(n21923),.dinb(w_n21197_0[0]),.dout(n21924),.clk(gclk));
	jor g21667(.dina(w_n21924_0[2]),.dinb(n21921),.dout(n21925),.clk(gclk));
	jand g21668(.dina(n21925),.dinb(w_n21920_0[1]),.dout(n21926),.clk(gclk));
	jor g21669(.dina(w_n21926_0[2]),.dinb(w_n18442_8[0]),.dout(n21927),.clk(gclk));
	jand g21670(.dina(w_n21926_0[1]),.dinb(w_n18442_7[2]),.dout(n21928),.clk(gclk));
	jxor g21671(.dina(w_n21199_0[0]),.dinb(w_n19096_15[1]),.dout(n21929),.clk(gclk));
	jor g21672(.dina(n21929),.dinb(w_n21887_32[2]),.dout(n21930),.clk(gclk));
	jxor g21673(.dina(n21930),.dinb(w_n21688_0[0]),.dout(n21931),.clk(gclk));
	jnot g21674(.din(w_n21931_0[2]),.dout(n21932),.clk(gclk));
	jor g21675(.dina(n21932),.dinb(n21928),.dout(n21933),.clk(gclk));
	jand g21676(.dina(n21933),.dinb(w_n21927_0[1]),.dout(n21934),.clk(gclk));
	jor g21677(.dina(w_n21934_0[2]),.dinb(w_n17769_16[2]),.dout(n21935),.clk(gclk));
	jand g21678(.dina(w_n21934_0[1]),.dinb(w_n17769_16[1]),.dout(n21936),.clk(gclk));
	jxor g21679(.dina(w_n21206_0[0]),.dinb(w_n18442_7[1]),.dout(n21937),.clk(gclk));
	jor g21680(.dina(n21937),.dinb(w_n21887_32[1]),.dout(n21938),.clk(gclk));
	jxor g21681(.dina(n21938),.dinb(w_n21212_0[0]),.dout(n21939),.clk(gclk));
	jor g21682(.dina(w_n21939_0[2]),.dinb(n21936),.dout(n21940),.clk(gclk));
	jand g21683(.dina(n21940),.dinb(w_n21935_0[1]),.dout(n21941),.clk(gclk));
	jor g21684(.dina(w_n21941_0[2]),.dinb(w_n17134_9[0]),.dout(n21942),.clk(gclk));
	jand g21685(.dina(w_n21941_0[1]),.dinb(w_n17134_8[2]),.dout(n21943),.clk(gclk));
	jxor g21686(.dina(w_n21214_0[0]),.dinb(w_n17769_16[0]),.dout(n21944),.clk(gclk));
	jor g21687(.dina(n21944),.dinb(w_n21887_32[0]),.dout(n21945),.clk(gclk));
	jxor g21688(.dina(n21945),.dinb(w_n21695_0[0]),.dout(n21946),.clk(gclk));
	jnot g21689(.din(w_n21946_0[2]),.dout(n21947),.clk(gclk));
	jor g21690(.dina(n21947),.dinb(n21943),.dout(n21948),.clk(gclk));
	jand g21691(.dina(n21948),.dinb(w_n21942_0[1]),.dout(n21949),.clk(gclk));
	jor g21692(.dina(w_n21949_0[2]),.dinb(w_n16489_17[0]),.dout(n21950),.clk(gclk));
	jand g21693(.dina(w_n21949_0[1]),.dinb(w_n16489_16[2]),.dout(n21951),.clk(gclk));
	jxor g21694(.dina(w_n21221_0[0]),.dinb(w_n17134_8[1]),.dout(n21952),.clk(gclk));
	jor g21695(.dina(n21952),.dinb(w_n21887_31[2]),.dout(n21953),.clk(gclk));
	jxor g21696(.dina(n21953),.dinb(w_n21227_0[0]),.dout(n21954),.clk(gclk));
	jor g21697(.dina(w_n21954_0[2]),.dinb(n21951),.dout(n21955),.clk(gclk));
	jand g21698(.dina(n21955),.dinb(w_n21950_0[1]),.dout(n21956),.clk(gclk));
	jor g21699(.dina(w_n21956_0[2]),.dinb(w_n15878_10[0]),.dout(n21957),.clk(gclk));
	jand g21700(.dina(w_n21956_0[1]),.dinb(w_n15878_9[2]),.dout(n21958),.clk(gclk));
	jxor g21701(.dina(w_n21229_0[0]),.dinb(w_n16489_16[1]),.dout(n21959),.clk(gclk));
	jor g21702(.dina(n21959),.dinb(w_n21887_31[1]),.dout(n21960),.clk(gclk));
	jxor g21703(.dina(n21960),.dinb(w_n21235_0[0]),.dout(n21961),.clk(gclk));
	jor g21704(.dina(w_n21961_0[2]),.dinb(n21958),.dout(n21962),.clk(gclk));
	jand g21705(.dina(n21962),.dinb(w_n21957_0[1]),.dout(n21963),.clk(gclk));
	jor g21706(.dina(w_n21963_0[2]),.dinb(w_n15260_17[2]),.dout(n21964),.clk(gclk));
	jand g21707(.dina(w_n21963_0[1]),.dinb(w_n15260_17[1]),.dout(n21965),.clk(gclk));
	jxor g21708(.dina(w_n21237_0[0]),.dinb(w_n15878_9[1]),.dout(n21966),.clk(gclk));
	jor g21709(.dina(n21966),.dinb(w_n21887_31[0]),.dout(n21967),.clk(gclk));
	jxor g21710(.dina(n21967),.dinb(w_n21243_0[0]),.dout(n21968),.clk(gclk));
	jor g21711(.dina(w_n21968_0[2]),.dinb(n21965),.dout(n21969),.clk(gclk));
	jand g21712(.dina(n21969),.dinb(w_n21964_0[1]),.dout(n21970),.clk(gclk));
	jor g21713(.dina(w_n21970_0[2]),.dinb(w_n14674_10[2]),.dout(n21971),.clk(gclk));
	jand g21714(.dina(w_n21970_0[1]),.dinb(w_n14674_10[1]),.dout(n21972),.clk(gclk));
	jxor g21715(.dina(w_n21245_0[0]),.dinb(w_n15260_17[0]),.dout(n21973),.clk(gclk));
	jor g21716(.dina(n21973),.dinb(w_n21887_30[2]),.dout(n21974),.clk(gclk));
	jxor g21717(.dina(n21974),.dinb(w_n21708_0[0]),.dout(n21975),.clk(gclk));
	jnot g21718(.din(w_n21975_0[2]),.dout(n21976),.clk(gclk));
	jor g21719(.dina(n21976),.dinb(n21972),.dout(n21977),.clk(gclk));
	jand g21720(.dina(n21977),.dinb(w_n21971_0[1]),.dout(n21978),.clk(gclk));
	jor g21721(.dina(w_n21978_0[2]),.dinb(w_n14078_18[0]),.dout(n21979),.clk(gclk));
	jand g21722(.dina(w_n21978_0[1]),.dinb(w_n14078_17[2]),.dout(n21980),.clk(gclk));
	jxor g21723(.dina(w_n21252_0[0]),.dinb(w_n14674_10[0]),.dout(n21981),.clk(gclk));
	jor g21724(.dina(n21981),.dinb(w_n21887_30[1]),.dout(n21982),.clk(gclk));
	jxor g21725(.dina(n21982),.dinb(w_n21258_0[0]),.dout(n21983),.clk(gclk));
	jor g21726(.dina(w_n21983_0[2]),.dinb(n21980),.dout(n21984),.clk(gclk));
	jand g21727(.dina(n21984),.dinb(w_n21979_0[1]),.dout(n21985),.clk(gclk));
	jor g21728(.dina(w_n21985_0[2]),.dinb(w_n13515_11[2]),.dout(n21986),.clk(gclk));
	jand g21729(.dina(w_n21985_0[1]),.dinb(w_n13515_11[1]),.dout(n21987),.clk(gclk));
	jxor g21730(.dina(w_n21260_0[0]),.dinb(w_n14078_17[1]),.dout(n21988),.clk(gclk));
	jor g21731(.dina(n21988),.dinb(w_n21887_30[0]),.dout(n21989),.clk(gclk));
	jxor g21732(.dina(n21989),.dinb(w_n21266_0[0]),.dout(n21990),.clk(gclk));
	jor g21733(.dina(w_n21990_0[2]),.dinb(n21987),.dout(n21991),.clk(gclk));
	jand g21734(.dina(n21991),.dinb(w_n21986_0[1]),.dout(n21992),.clk(gclk));
	jor g21735(.dina(w_n21992_0[2]),.dinb(w_n12947_18[2]),.dout(n21993),.clk(gclk));
	jand g21736(.dina(w_n21992_0[1]),.dinb(w_n12947_18[1]),.dout(n21994),.clk(gclk));
	jxor g21737(.dina(w_n21268_0[0]),.dinb(w_n13515_11[0]),.dout(n21995),.clk(gclk));
	jor g21738(.dina(n21995),.dinb(w_n21887_29[2]),.dout(n21996),.clk(gclk));
	jxor g21739(.dina(n21996),.dinb(w_n21274_0[0]),.dout(n21997),.clk(gclk));
	jor g21740(.dina(w_n21997_0[2]),.dinb(n21994),.dout(n21998),.clk(gclk));
	jand g21741(.dina(n21998),.dinb(w_n21993_0[1]),.dout(n21999),.clk(gclk));
	jor g21742(.dina(w_n21999_0[2]),.dinb(w_n12410_12[1]),.dout(n22000),.clk(gclk));
	jand g21743(.dina(w_n21999_0[1]),.dinb(w_n12410_12[0]),.dout(n22001),.clk(gclk));
	jxor g21744(.dina(w_n21276_0[0]),.dinb(w_n12947_18[0]),.dout(n22002),.clk(gclk));
	jor g21745(.dina(n22002),.dinb(w_n21887_29[1]),.dout(n22003),.clk(gclk));
	jxor g21746(.dina(n22003),.dinb(w_n21721_0[0]),.dout(n22004),.clk(gclk));
	jnot g21747(.din(w_n22004_0[2]),.dout(n22005),.clk(gclk));
	jor g21748(.dina(n22005),.dinb(n22001),.dout(n22006),.clk(gclk));
	jand g21749(.dina(n22006),.dinb(w_n22000_0[1]),.dout(n22007),.clk(gclk));
	jor g21750(.dina(w_n22007_0[2]),.dinb(w_n11858_19[0]),.dout(n22008),.clk(gclk));
	jand g21751(.dina(w_n22007_0[1]),.dinb(w_n11858_18[2]),.dout(n22009),.clk(gclk));
	jxor g21752(.dina(w_n21283_0[0]),.dinb(w_n12410_11[2]),.dout(n22010),.clk(gclk));
	jor g21753(.dina(n22010),.dinb(w_n21887_29[0]),.dout(n22011),.clk(gclk));
	jxor g21754(.dina(n22011),.dinb(w_n21289_0[0]),.dout(n22012),.clk(gclk));
	jor g21755(.dina(w_n22012_0[2]),.dinb(n22009),.dout(n22013),.clk(gclk));
	jand g21756(.dina(n22013),.dinb(w_n22008_0[1]),.dout(n22014),.clk(gclk));
	jor g21757(.dina(w_n22014_0[2]),.dinb(w_n11347_13[0]),.dout(n22015),.clk(gclk));
	jand g21758(.dina(w_n22014_0[1]),.dinb(w_n11347_12[2]),.dout(n22016),.clk(gclk));
	jxor g21759(.dina(w_n21291_0[0]),.dinb(w_n11858_18[1]),.dout(n22017),.clk(gclk));
	jor g21760(.dina(n22017),.dinb(w_n21887_28[2]),.dout(n22018),.clk(gclk));
	jxor g21761(.dina(n22018),.dinb(w_n21728_0[0]),.dout(n22019),.clk(gclk));
	jnot g21762(.din(w_n22019_0[2]),.dout(n22020),.clk(gclk));
	jor g21763(.dina(n22020),.dinb(n22016),.dout(n22021),.clk(gclk));
	jand g21764(.dina(n22021),.dinb(w_n22015_0[1]),.dout(n22022),.clk(gclk));
	jor g21765(.dina(w_n22022_0[2]),.dinb(w_n10824_19[2]),.dout(n22023),.clk(gclk));
	jand g21766(.dina(w_n22022_0[1]),.dinb(w_n10824_19[1]),.dout(n22024),.clk(gclk));
	jxor g21767(.dina(w_n21298_0[0]),.dinb(w_n11347_12[1]),.dout(n22025),.clk(gclk));
	jor g21768(.dina(n22025),.dinb(w_n21887_28[1]),.dout(n22026),.clk(gclk));
	jxor g21769(.dina(n22026),.dinb(w_n21304_0[0]),.dout(n22027),.clk(gclk));
	jor g21770(.dina(w_n22027_0[2]),.dinb(n22024),.dout(n22028),.clk(gclk));
	jand g21771(.dina(n22028),.dinb(w_n22023_0[1]),.dout(n22029),.clk(gclk));
	jor g21772(.dina(w_n22029_0[2]),.dinb(w_n10328_14[0]),.dout(n22030),.clk(gclk));
	jand g21773(.dina(w_n22029_0[1]),.dinb(w_n10328_13[2]),.dout(n22031),.clk(gclk));
	jxor g21774(.dina(w_n21306_0[0]),.dinb(w_n10824_19[0]),.dout(n22032),.clk(gclk));
	jor g21775(.dina(n22032),.dinb(w_n21887_28[0]),.dout(n22033),.clk(gclk));
	jxor g21776(.dina(n22033),.dinb(w_n21735_0[0]),.dout(n22034),.clk(gclk));
	jnot g21777(.din(w_n22034_0[2]),.dout(n22035),.clk(gclk));
	jor g21778(.dina(n22035),.dinb(n22031),.dout(n22036),.clk(gclk));
	jand g21779(.dina(n22036),.dinb(w_n22030_0[1]),.dout(n22037),.clk(gclk));
	jor g21780(.dina(w_n22037_0[2]),.dinb(w_n9832_20[1]),.dout(n22038),.clk(gclk));
	jand g21781(.dina(w_n22037_0[1]),.dinb(w_n9832_20[0]),.dout(n22039),.clk(gclk));
	jxor g21782(.dina(w_n21313_0[0]),.dinb(w_n10328_13[1]),.dout(n22040),.clk(gclk));
	jor g21783(.dina(n22040),.dinb(w_n21887_27[2]),.dout(n22041),.clk(gclk));
	jxor g21784(.dina(n22041),.dinb(w_n21319_0[0]),.dout(n22042),.clk(gclk));
	jor g21785(.dina(w_n22042_0[2]),.dinb(n22039),.dout(n22043),.clk(gclk));
	jand g21786(.dina(n22043),.dinb(w_n22038_0[1]),.dout(n22044),.clk(gclk));
	jor g21787(.dina(w_n22044_0[2]),.dinb(w_n9369_15[0]),.dout(n22045),.clk(gclk));
	jand g21788(.dina(w_n22044_0[1]),.dinb(w_n9369_14[2]),.dout(n22046),.clk(gclk));
	jxor g21789(.dina(w_n21321_0[0]),.dinb(w_n9832_19[2]),.dout(n22047),.clk(gclk));
	jor g21790(.dina(n22047),.dinb(w_n21887_27[1]),.dout(n22048),.clk(gclk));
	jxor g21791(.dina(n22048),.dinb(w_n21327_0[0]),.dout(n22049),.clk(gclk));
	jor g21792(.dina(w_n22049_0[2]),.dinb(n22046),.dout(n22050),.clk(gclk));
	jand g21793(.dina(n22050),.dinb(w_n22045_0[1]),.dout(n22051),.clk(gclk));
	jor g21794(.dina(w_n22051_0[2]),.dinb(w_n8890_20[2]),.dout(n22052),.clk(gclk));
	jand g21795(.dina(w_n22051_0[1]),.dinb(w_n8890_20[1]),.dout(n22053),.clk(gclk));
	jxor g21796(.dina(w_n21329_0[0]),.dinb(w_n9369_14[1]),.dout(n22054),.clk(gclk));
	jor g21797(.dina(n22054),.dinb(w_n21887_27[0]),.dout(n22055),.clk(gclk));
	jxor g21798(.dina(n22055),.dinb(w_n21745_0[0]),.dout(n22056),.clk(gclk));
	jnot g21799(.din(w_n22056_0[2]),.dout(n22057),.clk(gclk));
	jor g21800(.dina(n22057),.dinb(n22053),.dout(n22058),.clk(gclk));
	jand g21801(.dina(n22058),.dinb(w_n22052_0[1]),.dout(n22059),.clk(gclk));
	jor g21802(.dina(w_n22059_0[2]),.dinb(w_n8449_15[2]),.dout(n22060),.clk(gclk));
	jand g21803(.dina(w_n22059_0[1]),.dinb(w_n8449_15[1]),.dout(n22061),.clk(gclk));
	jxor g21804(.dina(w_n21336_0[0]),.dinb(w_n8890_20[0]),.dout(n22062),.clk(gclk));
	jor g21805(.dina(n22062),.dinb(w_n21887_26[2]),.dout(n22063),.clk(gclk));
	jxor g21806(.dina(n22063),.dinb(w_n21749_0[0]),.dout(n22064),.clk(gclk));
	jnot g21807(.din(w_n22064_0[2]),.dout(n22065),.clk(gclk));
	jor g21808(.dina(n22065),.dinb(n22061),.dout(n22066),.clk(gclk));
	jand g21809(.dina(n22066),.dinb(w_n22060_0[1]),.dout(n22067),.clk(gclk));
	jor g21810(.dina(w_n22067_0[2]),.dinb(w_n8003_21[1]),.dout(n22068),.clk(gclk));
	jand g21811(.dina(w_n22067_0[1]),.dinb(w_n8003_21[0]),.dout(n22069),.clk(gclk));
	jxor g21812(.dina(w_n21343_0[0]),.dinb(w_n8449_15[0]),.dout(n22070),.clk(gclk));
	jor g21813(.dina(n22070),.dinb(w_n21887_26[1]),.dout(n22071),.clk(gclk));
	jxor g21814(.dina(n22071),.dinb(w_n21349_0[0]),.dout(n22072),.clk(gclk));
	jor g21815(.dina(w_n22072_0[2]),.dinb(n22069),.dout(n22073),.clk(gclk));
	jand g21816(.dina(n22073),.dinb(w_n22068_0[1]),.dout(n22074),.clk(gclk));
	jor g21817(.dina(w_n22074_0[2]),.dinb(w_n7581_16[2]),.dout(n22075),.clk(gclk));
	jand g21818(.dina(w_n22074_0[1]),.dinb(w_n7581_16[1]),.dout(n22076),.clk(gclk));
	jxor g21819(.dina(w_n21351_0[0]),.dinb(w_n8003_20[2]),.dout(n22077),.clk(gclk));
	jor g21820(.dina(n22077),.dinb(w_n21887_26[0]),.dout(n22078),.clk(gclk));
	jxor g21821(.dina(n22078),.dinb(w_n21756_0[0]),.dout(n22079),.clk(gclk));
	jnot g21822(.din(w_n22079_0[2]),.dout(n22080),.clk(gclk));
	jor g21823(.dina(n22080),.dinb(n22076),.dout(n22081),.clk(gclk));
	jand g21824(.dina(n22081),.dinb(w_n22075_0[1]),.dout(n22082),.clk(gclk));
	jor g21825(.dina(w_n22082_0[2]),.dinb(w_n7154_21[2]),.dout(n22083),.clk(gclk));
	jand g21826(.dina(w_n22082_0[1]),.dinb(w_n7154_21[1]),.dout(n22084),.clk(gclk));
	jxor g21827(.dina(w_n21358_0[0]),.dinb(w_n7581_16[0]),.dout(n22085),.clk(gclk));
	jor g21828(.dina(n22085),.dinb(w_n21887_25[2]),.dout(n22086),.clk(gclk));
	jxor g21829(.dina(n22086),.dinb(w_n21364_0[0]),.dout(n22087),.clk(gclk));
	jor g21830(.dina(w_n22087_0[2]),.dinb(n22084),.dout(n22088),.clk(gclk));
	jand g21831(.dina(n22088),.dinb(w_n22083_0[1]),.dout(n22089),.clk(gclk));
	jor g21832(.dina(w_n22089_0[2]),.dinb(w_n6758_17[1]),.dout(n22090),.clk(gclk));
	jand g21833(.dina(w_n22089_0[1]),.dinb(w_n6758_17[0]),.dout(n22091),.clk(gclk));
	jxor g21834(.dina(w_n21366_0[0]),.dinb(w_n7154_21[0]),.dout(n22092),.clk(gclk));
	jor g21835(.dina(n22092),.dinb(w_n21887_25[1]),.dout(n22093),.clk(gclk));
	jxor g21836(.dina(n22093),.dinb(w_n21763_0[0]),.dout(n22094),.clk(gclk));
	jnot g21837(.din(w_n22094_0[2]),.dout(n22095),.clk(gclk));
	jor g21838(.dina(n22095),.dinb(n22091),.dout(n22096),.clk(gclk));
	jand g21839(.dina(n22096),.dinb(w_n22090_0[1]),.dout(n22097),.clk(gclk));
	jor g21840(.dina(w_n22097_0[2]),.dinb(w_n6357_22[0]),.dout(n22098),.clk(gclk));
	jand g21841(.dina(w_n22097_0[1]),.dinb(w_n6357_21[2]),.dout(n22099),.clk(gclk));
	jxor g21842(.dina(w_n21373_0[0]),.dinb(w_n6758_16[2]),.dout(n22100),.clk(gclk));
	jor g21843(.dina(n22100),.dinb(w_n21887_25[0]),.dout(n22101),.clk(gclk));
	jxor g21844(.dina(n22101),.dinb(w_n21379_0[0]),.dout(n22102),.clk(gclk));
	jor g21845(.dina(w_n22102_0[2]),.dinb(n22099),.dout(n22103),.clk(gclk));
	jand g21846(.dina(n22103),.dinb(w_n22098_0[1]),.dout(n22104),.clk(gclk));
	jor g21847(.dina(w_n22104_0[2]),.dinb(w_n5989_18[0]),.dout(n22105),.clk(gclk));
	jand g21848(.dina(w_n22104_0[1]),.dinb(w_n5989_17[2]),.dout(n22106),.clk(gclk));
	jxor g21849(.dina(w_n21381_0[0]),.dinb(w_n6357_21[1]),.dout(n22107),.clk(gclk));
	jor g21850(.dina(n22107),.dinb(w_n21887_24[2]),.dout(n22108),.clk(gclk));
	jxor g21851(.dina(n22108),.dinb(w_n21387_0[0]),.dout(n22109),.clk(gclk));
	jor g21852(.dina(w_n22109_0[2]),.dinb(n22106),.dout(n22110),.clk(gclk));
	jand g21853(.dina(n22110),.dinb(w_n22105_0[1]),.dout(n22111),.clk(gclk));
	jor g21854(.dina(w_n22111_0[2]),.dinb(w_n5606_22[1]),.dout(n22112),.clk(gclk));
	jand g21855(.dina(w_n22111_0[1]),.dinb(w_n5606_22[0]),.dout(n22113),.clk(gclk));
	jxor g21856(.dina(w_n21389_0[0]),.dinb(w_n5989_17[1]),.dout(n22114),.clk(gclk));
	jor g21857(.dina(n22114),.dinb(w_n21887_24[1]),.dout(n22115),.clk(gclk));
	jxor g21858(.dina(n22115),.dinb(w_n21395_0[0]),.dout(n22116),.clk(gclk));
	jor g21859(.dina(w_n22116_0[2]),.dinb(n22113),.dout(n22117),.clk(gclk));
	jand g21860(.dina(n22117),.dinb(w_n22112_0[1]),.dout(n22118),.clk(gclk));
	jor g21861(.dina(w_n22118_0[2]),.dinb(w_n5259_19[0]),.dout(n22119),.clk(gclk));
	jand g21862(.dina(w_n22118_0[1]),.dinb(w_n5259_18[2]),.dout(n22120),.clk(gclk));
	jxor g21863(.dina(w_n21397_0[0]),.dinb(w_n5606_21[2]),.dout(n22121),.clk(gclk));
	jor g21864(.dina(n22121),.dinb(w_n21887_24[0]),.dout(n22122),.clk(gclk));
	jxor g21865(.dina(n22122),.dinb(w_n21776_0[0]),.dout(n22123),.clk(gclk));
	jnot g21866(.din(w_n22123_0[2]),.dout(n22124),.clk(gclk));
	jor g21867(.dina(n22124),.dinb(n22120),.dout(n22125),.clk(gclk));
	jand g21868(.dina(n22125),.dinb(w_n22119_0[1]),.dout(n22126),.clk(gclk));
	jor g21869(.dina(w_n22126_0[2]),.dinb(w_n4902_23[0]),.dout(n22127),.clk(gclk));
	jand g21870(.dina(w_n22126_0[1]),.dinb(w_n4902_22[2]),.dout(n22128),.clk(gclk));
	jxor g21871(.dina(w_n21404_0[0]),.dinb(w_n5259_18[1]),.dout(n22129),.clk(gclk));
	jor g21872(.dina(n22129),.dinb(w_n21887_23[2]),.dout(n22130),.clk(gclk));
	jxor g21873(.dina(n22130),.dinb(w_n21410_0[0]),.dout(n22131),.clk(gclk));
	jor g21874(.dina(w_n22131_0[2]),.dinb(n22128),.dout(n22132),.clk(gclk));
	jand g21875(.dina(n22132),.dinb(w_n22127_0[1]),.dout(n22133),.clk(gclk));
	jor g21876(.dina(w_n22133_0[2]),.dinb(w_n4582_20[0]),.dout(n22134),.clk(gclk));
	jand g21877(.dina(w_n22133_0[1]),.dinb(w_n4582_19[2]),.dout(n22135),.clk(gclk));
	jxor g21878(.dina(w_n21412_0[0]),.dinb(w_n4902_22[1]),.dout(n22136),.clk(gclk));
	jor g21879(.dina(n22136),.dinb(w_n21887_23[1]),.dout(n22137),.clk(gclk));
	jxor g21880(.dina(n22137),.dinb(w_n21783_0[0]),.dout(n22138),.clk(gclk));
	jnot g21881(.din(w_n22138_0[2]),.dout(n22139),.clk(gclk));
	jor g21882(.dina(n22139),.dinb(n22135),.dout(n22140),.clk(gclk));
	jand g21883(.dina(n22140),.dinb(w_n22134_0[1]),.dout(n22141),.clk(gclk));
	jor g21884(.dina(w_n22141_0[2]),.dinb(w_n4249_23[2]),.dout(n22142),.clk(gclk));
	jand g21885(.dina(w_n22141_0[1]),.dinb(w_n4249_23[1]),.dout(n22143),.clk(gclk));
	jxor g21886(.dina(w_n21419_0[0]),.dinb(w_n4582_19[1]),.dout(n22144),.clk(gclk));
	jor g21887(.dina(n22144),.dinb(w_n21887_23[0]),.dout(n22145),.clk(gclk));
	jxor g21888(.dina(n22145),.dinb(w_n21425_0[0]),.dout(n22146),.clk(gclk));
	jor g21889(.dina(w_n22146_0[2]),.dinb(n22143),.dout(n22147),.clk(gclk));
	jand g21890(.dina(n22147),.dinb(w_n22142_0[1]),.dout(n22148),.clk(gclk));
	jor g21891(.dina(w_n22148_0[2]),.dinb(w_n3955_20[2]),.dout(n22149),.clk(gclk));
	jand g21892(.dina(w_n22148_0[1]),.dinb(w_n3955_20[1]),.dout(n22150),.clk(gclk));
	jxor g21893(.dina(w_n21427_0[0]),.dinb(w_n4249_23[0]),.dout(n22151),.clk(gclk));
	jor g21894(.dina(n22151),.dinb(w_n21887_22[2]),.dout(n22152),.clk(gclk));
	jxor g21895(.dina(n22152),.dinb(w_n21790_0[0]),.dout(n22153),.clk(gclk));
	jnot g21896(.din(w_n22153_0[2]),.dout(n22154),.clk(gclk));
	jor g21897(.dina(n22154),.dinb(n22150),.dout(n22155),.clk(gclk));
	jand g21898(.dina(n22155),.dinb(w_n22149_0[1]),.dout(n22156),.clk(gclk));
	jor g21899(.dina(w_n22156_0[2]),.dinb(w_n3642_24[0]),.dout(n22157),.clk(gclk));
	jand g21900(.dina(w_n22156_0[1]),.dinb(w_n3642_23[2]),.dout(n22158),.clk(gclk));
	jxor g21901(.dina(w_n21434_0[0]),.dinb(w_n3955_20[0]),.dout(n22159),.clk(gclk));
	jor g21902(.dina(n22159),.dinb(w_n21887_22[1]),.dout(n22160),.clk(gclk));
	jxor g21903(.dina(n22160),.dinb(w_n21440_0[0]),.dout(n22161),.clk(gclk));
	jor g21904(.dina(w_n22161_0[2]),.dinb(n22158),.dout(n22162),.clk(gclk));
	jand g21905(.dina(n22162),.dinb(w_n22157_0[1]),.dout(n22163),.clk(gclk));
	jor g21906(.dina(w_n22163_0[2]),.dinb(w_n3368_21[1]),.dout(n22164),.clk(gclk));
	jand g21907(.dina(w_n22163_0[1]),.dinb(w_n3368_21[0]),.dout(n22165),.clk(gclk));
	jxor g21908(.dina(w_n21442_0[0]),.dinb(w_n3642_23[1]),.dout(n22166),.clk(gclk));
	jor g21909(.dina(n22166),.dinb(w_n21887_22[0]),.dout(n22167),.clk(gclk));
	jxor g21910(.dina(n22167),.dinb(w_n21797_0[0]),.dout(n22168),.clk(gclk));
	jnot g21911(.din(w_n22168_0[2]),.dout(n22169),.clk(gclk));
	jor g21912(.dina(n22169),.dinb(n22165),.dout(n22170),.clk(gclk));
	jand g21913(.dina(n22170),.dinb(w_n22164_0[1]),.dout(n22171),.clk(gclk));
	jor g21914(.dina(w_n22171_0[2]),.dinb(w_n3089_24[2]),.dout(n22172),.clk(gclk));
	jand g21915(.dina(w_n22171_0[1]),.dinb(w_n3089_24[1]),.dout(n22173),.clk(gclk));
	jxor g21916(.dina(w_n21449_0[0]),.dinb(w_n3368_20[2]),.dout(n22174),.clk(gclk));
	jor g21917(.dina(n22174),.dinb(w_n21887_21[2]),.dout(n22175),.clk(gclk));
	jxor g21918(.dina(n22175),.dinb(w_n21455_0[0]),.dout(n22176),.clk(gclk));
	jor g21919(.dina(w_n22176_0[2]),.dinb(n22173),.dout(n22177),.clk(gclk));
	jand g21920(.dina(n22177),.dinb(w_n22172_0[1]),.dout(n22178),.clk(gclk));
	jor g21921(.dina(w_n22178_0[2]),.dinb(w_n2833_22[1]),.dout(n22179),.clk(gclk));
	jand g21922(.dina(w_n22178_0[1]),.dinb(w_n2833_22[0]),.dout(n22180),.clk(gclk));
	jxor g21923(.dina(w_n21457_0[0]),.dinb(w_n3089_24[0]),.dout(n22181),.clk(gclk));
	jor g21924(.dina(n22181),.dinb(w_n21887_21[1]),.dout(n22182),.clk(gclk));
	jxor g21925(.dina(n22182),.dinb(w_n21463_0[0]),.dout(n22183),.clk(gclk));
	jor g21926(.dina(w_n22183_0[2]),.dinb(n22180),.dout(n22184),.clk(gclk));
	jand g21927(.dina(n22184),.dinb(w_n22179_0[1]),.dout(n22185),.clk(gclk));
	jor g21928(.dina(w_n22185_0[2]),.dinb(w_n2572_25[0]),.dout(n22186),.clk(gclk));
	jand g21929(.dina(w_n22185_0[1]),.dinb(w_n2572_24[2]),.dout(n22187),.clk(gclk));
	jxor g21930(.dina(w_n21465_0[0]),.dinb(w_n2833_21[2]),.dout(n22188),.clk(gclk));
	jor g21931(.dina(n22188),.dinb(w_n21887_21[0]),.dout(n22189),.clk(gclk));
	jxor g21932(.dina(n22189),.dinb(w_n21471_0[0]),.dout(n22190),.clk(gclk));
	jor g21933(.dina(w_n22190_0[2]),.dinb(n22187),.dout(n22191),.clk(gclk));
	jand g21934(.dina(n22191),.dinb(w_n22186_0[1]),.dout(n22192),.clk(gclk));
	jor g21935(.dina(w_n22192_0[2]),.dinb(w_n2345_23[0]),.dout(n22193),.clk(gclk));
	jand g21936(.dina(w_n22192_0[1]),.dinb(w_n2345_22[2]),.dout(n22194),.clk(gclk));
	jxor g21937(.dina(w_n21473_0[0]),.dinb(w_n2572_24[1]),.dout(n22195),.clk(gclk));
	jor g21938(.dina(n22195),.dinb(w_n21887_20[2]),.dout(n22196),.clk(gclk));
	jxor g21939(.dina(n22196),.dinb(w_n21810_0[0]),.dout(n22197),.clk(gclk));
	jnot g21940(.din(w_n22197_0[2]),.dout(n22198),.clk(gclk));
	jor g21941(.dina(n22198),.dinb(n22194),.dout(n22199),.clk(gclk));
	jand g21942(.dina(n22199),.dinb(w_n22193_0[1]),.dout(n22200),.clk(gclk));
	jor g21943(.dina(w_n22200_0[2]),.dinb(w_n2108_25[2]),.dout(n22201),.clk(gclk));
	jand g21944(.dina(w_n22200_0[1]),.dinb(w_n2108_25[1]),.dout(n22202),.clk(gclk));
	jxor g21945(.dina(w_n21480_0[0]),.dinb(w_n2345_22[1]),.dout(n22203),.clk(gclk));
	jor g21946(.dina(n22203),.dinb(w_n21887_20[1]),.dout(n22204),.clk(gclk));
	jxor g21947(.dina(n22204),.dinb(w_n21486_0[0]),.dout(n22205),.clk(gclk));
	jor g21948(.dina(w_n22205_0[2]),.dinb(n22202),.dout(n22206),.clk(gclk));
	jand g21949(.dina(n22206),.dinb(w_n22201_0[1]),.dout(n22207),.clk(gclk));
	jor g21950(.dina(w_n22207_0[2]),.dinb(w_n1912_24[0]),.dout(n22208),.clk(gclk));
	jand g21951(.dina(w_n22207_0[1]),.dinb(w_n1912_23[2]),.dout(n22209),.clk(gclk));
	jxor g21952(.dina(w_n21488_0[0]),.dinb(w_n2108_25[0]),.dout(n22210),.clk(gclk));
	jor g21953(.dina(n22210),.dinb(w_n21887_20[0]),.dout(n22211),.clk(gclk));
	jxor g21954(.dina(n22211),.dinb(w_n21494_0[0]),.dout(n22212),.clk(gclk));
	jor g21955(.dina(w_n22212_0[2]),.dinb(n22209),.dout(n22213),.clk(gclk));
	jand g21956(.dina(n22213),.dinb(w_n22208_0[1]),.dout(n22214),.clk(gclk));
	jor g21957(.dina(w_n22214_0[2]),.dinb(w_n1699_26[1]),.dout(n22215),.clk(gclk));
	jand g21958(.dina(w_n22214_0[1]),.dinb(w_n1699_26[0]),.dout(n22216),.clk(gclk));
	jxor g21959(.dina(w_n21496_0[0]),.dinb(w_n1912_23[1]),.dout(n22217),.clk(gclk));
	jor g21960(.dina(n22217),.dinb(w_n21887_19[2]),.dout(n22218),.clk(gclk));
	jxor g21961(.dina(n22218),.dinb(w_n21502_0[0]),.dout(n22219),.clk(gclk));
	jor g21962(.dina(w_n22219_0[2]),.dinb(n22216),.dout(n22220),.clk(gclk));
	jand g21963(.dina(n22220),.dinb(w_n22215_0[1]),.dout(n22221),.clk(gclk));
	jor g21964(.dina(w_n22221_0[2]),.dinb(w_n1516_24[2]),.dout(n22222),.clk(gclk));
	jand g21965(.dina(w_n22221_0[1]),.dinb(w_n1516_24[1]),.dout(n22223),.clk(gclk));
	jxor g21966(.dina(w_n21504_0[0]),.dinb(w_n1699_25[2]),.dout(n22224),.clk(gclk));
	jor g21967(.dina(n22224),.dinb(w_n21887_19[1]),.dout(n22225),.clk(gclk));
	jxor g21968(.dina(n22225),.dinb(w_n21510_0[0]),.dout(n22226),.clk(gclk));
	jor g21969(.dina(w_n22226_0[2]),.dinb(n22223),.dout(n22227),.clk(gclk));
	jand g21970(.dina(n22227),.dinb(w_n22222_0[1]),.dout(n22228),.clk(gclk));
	jor g21971(.dina(w_n22228_0[2]),.dinb(w_n1332_26[1]),.dout(n22229),.clk(gclk));
	jand g21972(.dina(w_n22228_0[1]),.dinb(w_n1332_26[0]),.dout(n22230),.clk(gclk));
	jxor g21973(.dina(w_n21512_0[0]),.dinb(w_n1516_24[0]),.dout(n22231),.clk(gclk));
	jor g21974(.dina(n22231),.dinb(w_n21887_19[0]),.dout(n22232),.clk(gclk));
	jxor g21975(.dina(n22232),.dinb(w_n21518_0[0]),.dout(n22233),.clk(gclk));
	jor g21976(.dina(w_n22233_0[2]),.dinb(n22230),.dout(n22234),.clk(gclk));
	jand g21977(.dina(n22234),.dinb(w_n22229_0[1]),.dout(n22235),.clk(gclk));
	jor g21978(.dina(w_n22235_0[2]),.dinb(w_n1173_25[1]),.dout(n22236),.clk(gclk));
	jand g21979(.dina(w_n22235_0[1]),.dinb(w_n1173_25[0]),.dout(n22237),.clk(gclk));
	jxor g21980(.dina(w_n21520_0[0]),.dinb(w_n1332_25[2]),.dout(n22238),.clk(gclk));
	jor g21981(.dina(n22238),.dinb(w_n21887_18[2]),.dout(n22239),.clk(gclk));
	jxor g21982(.dina(n22239),.dinb(w_n21829_0[0]),.dout(n22240),.clk(gclk));
	jnot g21983(.din(w_n22240_0[2]),.dout(n22241),.clk(gclk));
	jor g21984(.dina(n22241),.dinb(n22237),.dout(n22242),.clk(gclk));
	jand g21985(.dina(n22242),.dinb(w_n22236_0[1]),.dout(n22243),.clk(gclk));
	jor g21986(.dina(w_n22243_0[2]),.dinb(w_n1008_27[1]),.dout(n22244),.clk(gclk));
	jand g21987(.dina(w_n22243_0[1]),.dinb(w_n1008_27[0]),.dout(n22245),.clk(gclk));
	jxor g21988(.dina(w_n21527_0[0]),.dinb(w_n1173_24[2]),.dout(n22246),.clk(gclk));
	jor g21989(.dina(n22246),.dinb(w_n21887_18[1]),.dout(n22247),.clk(gclk));
	jxor g21990(.dina(n22247),.dinb(w_n21533_0[0]),.dout(n22248),.clk(gclk));
	jor g21991(.dina(w_n22248_0[2]),.dinb(n22245),.dout(n22249),.clk(gclk));
	jand g21992(.dina(n22249),.dinb(w_n22244_0[1]),.dout(n22250),.clk(gclk));
	jor g21993(.dina(w_n22250_0[2]),.dinb(w_n884_26[1]),.dout(n22251),.clk(gclk));
	jand g21994(.dina(w_n22250_0[1]),.dinb(w_n884_26[0]),.dout(n22252),.clk(gclk));
	jxor g21995(.dina(w_n21535_0[0]),.dinb(w_n1008_26[2]),.dout(n22253),.clk(gclk));
	jor g21996(.dina(n22253),.dinb(w_n21887_18[0]),.dout(n22254),.clk(gclk));
	jxor g21997(.dina(n22254),.dinb(w_n21836_0[0]),.dout(n22255),.clk(gclk));
	jnot g21998(.din(w_n22255_0[2]),.dout(n22256),.clk(gclk));
	jor g21999(.dina(n22256),.dinb(n22252),.dout(n22257),.clk(gclk));
	jand g22000(.dina(n22257),.dinb(w_n22251_0[1]),.dout(n22258),.clk(gclk));
	jor g22001(.dina(w_n22258_0[2]),.dinb(w_n743_27[1]),.dout(n22259),.clk(gclk));
	jand g22002(.dina(w_n22258_0[1]),.dinb(w_n743_27[0]),.dout(n22260),.clk(gclk));
	jxor g22003(.dina(w_n21542_0[0]),.dinb(w_n884_25[2]),.dout(n22261),.clk(gclk));
	jor g22004(.dina(n22261),.dinb(w_n21887_17[2]),.dout(n22262),.clk(gclk));
	jxor g22005(.dina(n22262),.dinb(w_n21548_0[0]),.dout(n22263),.clk(gclk));
	jor g22006(.dina(w_n22263_0[2]),.dinb(n22260),.dout(n22264),.clk(gclk));
	jand g22007(.dina(n22264),.dinb(w_n22259_0[1]),.dout(n22265),.clk(gclk));
	jor g22008(.dina(w_n22265_0[2]),.dinb(w_n635_27[1]),.dout(n22266),.clk(gclk));
	jand g22009(.dina(w_n22265_0[1]),.dinb(w_n635_27[0]),.dout(n22267),.clk(gclk));
	jxor g22010(.dina(w_n21550_0[0]),.dinb(w_n743_26[2]),.dout(n22268),.clk(gclk));
	jor g22011(.dina(n22268),.dinb(w_n21887_17[1]),.dout(n22269),.clk(gclk));
	jxor g22012(.dina(n22269),.dinb(w_n21556_0[0]),.dout(n22270),.clk(gclk));
	jor g22013(.dina(w_n22270_0[2]),.dinb(n22267),.dout(n22271),.clk(gclk));
	jand g22014(.dina(n22271),.dinb(w_n22266_0[1]),.dout(n22272),.clk(gclk));
	jor g22015(.dina(w_n22272_0[2]),.dinb(w_n515_28[1]),.dout(n22273),.clk(gclk));
	jand g22016(.dina(w_n22272_0[1]),.dinb(w_n515_28[0]),.dout(n22274),.clk(gclk));
	jxor g22017(.dina(w_n21558_0[0]),.dinb(w_n635_26[2]),.dout(n22275),.clk(gclk));
	jor g22018(.dina(n22275),.dinb(w_n21887_17[0]),.dout(n22276),.clk(gclk));
	jxor g22019(.dina(n22276),.dinb(w_n21846_0[0]),.dout(n22277),.clk(gclk));
	jnot g22020(.din(w_n22277_0[2]),.dout(n22278),.clk(gclk));
	jor g22021(.dina(n22278),.dinb(n22274),.dout(n22279),.clk(gclk));
	jand g22022(.dina(n22279),.dinb(w_n22273_0[1]),.dout(n22280),.clk(gclk));
	jor g22023(.dina(w_n22280_0[2]),.dinb(w_n443_28[1]),.dout(n22281),.clk(gclk));
	jand g22024(.dina(w_n22280_0[1]),.dinb(w_n443_28[0]),.dout(n22282),.clk(gclk));
	jxor g22025(.dina(w_n21565_0[0]),.dinb(w_n515_27[2]),.dout(n22283),.clk(gclk));
	jor g22026(.dina(n22283),.dinb(w_n21887_16[2]),.dout(n22284),.clk(gclk));
	jxor g22027(.dina(n22284),.dinb(w_n21850_0[0]),.dout(n22285),.clk(gclk));
	jnot g22028(.din(w_n22285_0[2]),.dout(n22286),.clk(gclk));
	jor g22029(.dina(n22286),.dinb(n22282),.dout(n22287),.clk(gclk));
	jand g22030(.dina(n22287),.dinb(w_n22281_0[1]),.dout(n22288),.clk(gclk));
	jor g22031(.dina(w_n22288_0[2]),.dinb(w_n352_28[2]),.dout(n22289),.clk(gclk));
	jand g22032(.dina(w_n22288_0[1]),.dinb(w_n352_28[1]),.dout(n22290),.clk(gclk));
	jxor g22033(.dina(w_n21572_0[0]),.dinb(w_n443_27[2]),.dout(n22291),.clk(gclk));
	jor g22034(.dina(n22291),.dinb(w_n21887_16[1]),.dout(n22292),.clk(gclk));
	jxor g22035(.dina(n22292),.dinb(w_n21578_0[0]),.dout(n22293),.clk(gclk));
	jor g22036(.dina(w_n22293_0[2]),.dinb(n22290),.dout(n22294),.clk(gclk));
	jand g22037(.dina(n22294),.dinb(w_n22289_0[1]),.dout(n22295),.clk(gclk));
	jor g22038(.dina(w_n22295_0[2]),.dinb(w_n294_29[0]),.dout(n22296),.clk(gclk));
	jand g22039(.dina(w_n22295_0[1]),.dinb(w_n294_28[2]),.dout(n22297),.clk(gclk));
	jxor g22040(.dina(w_n21580_0[0]),.dinb(w_n352_28[0]),.dout(n22298),.clk(gclk));
	jor g22041(.dina(n22298),.dinb(w_n21887_16[0]),.dout(n22299),.clk(gclk));
	jxor g22042(.dina(n22299),.dinb(w_n21586_0[0]),.dout(n22300),.clk(gclk));
	jor g22043(.dina(w_n22300_0[2]),.dinb(n22297),.dout(n22301),.clk(gclk));
	jand g22044(.dina(n22301),.dinb(w_n22296_0[1]),.dout(n22302),.clk(gclk));
	jor g22045(.dina(w_n22302_0[2]),.dinb(w_n239_29[0]),.dout(n22303),.clk(gclk));
	jand g22046(.dina(w_n22302_0[1]),.dinb(w_n239_28[2]),.dout(n22304),.clk(gclk));
	jxor g22047(.dina(w_n21588_0[0]),.dinb(w_n294_28[1]),.dout(n22305),.clk(gclk));
	jor g22048(.dina(n22305),.dinb(w_n21887_15[2]),.dout(n22306),.clk(gclk));
	jxor g22049(.dina(n22306),.dinb(w_n21594_0[0]),.dout(n22307),.clk(gclk));
	jor g22050(.dina(w_n22307_0[2]),.dinb(n22304),.dout(n22308),.clk(gclk));
	jand g22051(.dina(n22308),.dinb(w_n22303_0[1]),.dout(n22309),.clk(gclk));
	jor g22052(.dina(w_n22309_0[2]),.dinb(w_n221_29[1]),.dout(n22310),.clk(gclk));
	jand g22053(.dina(w_n22309_0[1]),.dinb(w_n221_29[0]),.dout(n22311),.clk(gclk));
	jxor g22054(.dina(w_n21596_0[0]),.dinb(w_n239_28[1]),.dout(n22312),.clk(gclk));
	jor g22055(.dina(n22312),.dinb(w_n21887_15[1]),.dout(n22313),.clk(gclk));
	jxor g22056(.dina(n22313),.dinb(w_n21601_0[0]),.dout(n22314),.clk(gclk));
	jnot g22057(.din(w_n22314_0[1]),.dout(n22315),.clk(gclk));
	jor g22058(.dina(w_n22315_0[1]),.dinb(n22311),.dout(n22316),.clk(gclk));
	jand g22059(.dina(n22316),.dinb(w_n22310_0[1]),.dout(n22317),.clk(gclk));
	jxor g22060(.dina(w_n21604_0[0]),.dinb(w_n221_28[2]),.dout(n22318),.clk(gclk));
	jor g22061(.dina(n22318),.dinb(w_n21887_15[0]),.dout(n22319),.clk(gclk));
	jxor g22062(.dina(n22319),.dinb(w_n21609_0[0]),.dout(n22320),.clk(gclk));
	jand g22063(.dina(w_n22320_1[1]),.dinb(w_n22317_1[1]),.dout(n22321),.clk(gclk));
	jor g22064(.dina(w_n22320_1[0]),.dinb(w_n22317_1[0]),.dout(n22322),.clk(gclk));
	jxor g22065(.dina(w_n21615_0[0]),.dinb(w_n21611_0[0]),.dout(n22323),.clk(gclk));
	jnot g22066(.din(n22323),.dout(n22324),.clk(gclk));
	jand g22067(.dina(w_n22324_0[1]),.dinb(w_asqrt5_3[2]),.dout(n22325),.clk(gclk));
	jor g22068(.dina(w_n22325_0[1]),.dinb(n22322),.dout(n22326),.clk(gclk));
	jand g22069(.dina(n22326),.dinb(w_n218_12[1]),.dout(n22327),.clk(gclk));
	jand g22070(.dina(w_n21887_14[2]),.dinb(w_n21868_0[0]),.dout(n22328),.clk(gclk));
	jor g22071(.dina(n22328),.dinb(w_n22324_0[0]),.dout(n22329),.clk(gclk));
	jor g22072(.dina(n22329),.dinb(w_n218_12[0]),.dout(n22330),.clk(gclk));
	jnot g22073(.din(w_n22330_0[1]),.dout(n22331),.clk(gclk));
	jor g22074(.dina(n22331),.dinb(n22327),.dout(n22332),.clk(gclk));
	jor g22075(.dina(w_n22332_0[1]),.dinb(w_n22321_0[2]),.dout(asqrt_fa_5),.clk(gclk));
	jnot g22076(.din(w_a6_0[2]),.dout(n22334),.clk(gclk));
	jnot g22077(.din(w_a7_0[1]),.dout(n22335),.clk(gclk));
	jand g22078(.dina(w_n22335_0[1]),.dinb(w_n22334_1[2]),.dout(n22336),.clk(gclk));
	jand g22079(.dina(w_n22336_0[2]),.dinb(w_n21889_1[1]),.dout(n22337),.clk(gclk));
	jand g22080(.dina(w_asqrt4_31[1]),.dinb(w_a8_0[1]),.dout(n22338),.clk(gclk));
	jor g22081(.dina(n22338),.dinb(w_n22337_0[1]),.dout(n22339),.clk(gclk));
	jand g22082(.dina(w_n22339_0[2]),.dinb(w_asqrt5_3[1]),.dout(n22340),.clk(gclk));
	jor g22083(.dina(w_n22339_0[1]),.dinb(w_asqrt5_3[0]),.dout(n22341),.clk(gclk));
	jand g22084(.dina(w_asqrt4_31[0]),.dinb(w_n21889_1[0]),.dout(n22342),.clk(gclk));
	jor g22085(.dina(n22342),.dinb(w_n21890_0[0]),.dout(n22343),.clk(gclk));
	jnot g22086(.din(w_n21891_0[1]),.dout(n22344),.clk(gclk));
	jnot g22087(.din(w_n22321_0[1]),.dout(n22345),.clk(gclk));
	jnot g22088(.din(w_n22310_0[0]),.dout(n22346),.clk(gclk));
	jnot g22089(.din(w_n22303_0[0]),.dout(n22347),.clk(gclk));
	jnot g22090(.din(w_n22296_0[0]),.dout(n22348),.clk(gclk));
	jnot g22091(.din(w_n22289_0[0]),.dout(n22349),.clk(gclk));
	jnot g22092(.din(w_n22281_0[0]),.dout(n22350),.clk(gclk));
	jnot g22093(.din(w_n22273_0[0]),.dout(n22351),.clk(gclk));
	jnot g22094(.din(w_n22266_0[0]),.dout(n22352),.clk(gclk));
	jnot g22095(.din(w_n22259_0[0]),.dout(n22353),.clk(gclk));
	jnot g22096(.din(w_n22251_0[0]),.dout(n22354),.clk(gclk));
	jnot g22097(.din(w_n22244_0[0]),.dout(n22355),.clk(gclk));
	jnot g22098(.din(w_n22236_0[0]),.dout(n22356),.clk(gclk));
	jnot g22099(.din(w_n22229_0[0]),.dout(n22357),.clk(gclk));
	jnot g22100(.din(w_n22222_0[0]),.dout(n22358),.clk(gclk));
	jnot g22101(.din(w_n22215_0[0]),.dout(n22359),.clk(gclk));
	jnot g22102(.din(w_n22208_0[0]),.dout(n22360),.clk(gclk));
	jnot g22103(.din(w_n22201_0[0]),.dout(n22361),.clk(gclk));
	jnot g22104(.din(w_n22193_0[0]),.dout(n22362),.clk(gclk));
	jnot g22105(.din(w_n22186_0[0]),.dout(n22363),.clk(gclk));
	jnot g22106(.din(w_n22179_0[0]),.dout(n22364),.clk(gclk));
	jnot g22107(.din(w_n22172_0[0]),.dout(n22365),.clk(gclk));
	jnot g22108(.din(w_n22164_0[0]),.dout(n22366),.clk(gclk));
	jnot g22109(.din(w_n22157_0[0]),.dout(n22367),.clk(gclk));
	jnot g22110(.din(w_n22149_0[0]),.dout(n22368),.clk(gclk));
	jnot g22111(.din(w_n22142_0[0]),.dout(n22369),.clk(gclk));
	jnot g22112(.din(w_n22134_0[0]),.dout(n22370),.clk(gclk));
	jnot g22113(.din(w_n22127_0[0]),.dout(n22371),.clk(gclk));
	jnot g22114(.din(w_n22119_0[0]),.dout(n22372),.clk(gclk));
	jnot g22115(.din(w_n22112_0[0]),.dout(n22373),.clk(gclk));
	jnot g22116(.din(w_n22105_0[0]),.dout(n22374),.clk(gclk));
	jnot g22117(.din(w_n22098_0[0]),.dout(n22375),.clk(gclk));
	jnot g22118(.din(w_n22090_0[0]),.dout(n22376),.clk(gclk));
	jnot g22119(.din(w_n22083_0[0]),.dout(n22377),.clk(gclk));
	jnot g22120(.din(w_n22075_0[0]),.dout(n22378),.clk(gclk));
	jnot g22121(.din(w_n22068_0[0]),.dout(n22379),.clk(gclk));
	jnot g22122(.din(w_n22060_0[0]),.dout(n22380),.clk(gclk));
	jnot g22123(.din(w_n22052_0[0]),.dout(n22381),.clk(gclk));
	jnot g22124(.din(w_n22045_0[0]),.dout(n22382),.clk(gclk));
	jnot g22125(.din(w_n22038_0[0]),.dout(n22383),.clk(gclk));
	jnot g22126(.din(w_n22030_0[0]),.dout(n22384),.clk(gclk));
	jnot g22127(.din(w_n22023_0[0]),.dout(n22385),.clk(gclk));
	jnot g22128(.din(w_n22015_0[0]),.dout(n22386),.clk(gclk));
	jnot g22129(.din(w_n22008_0[0]),.dout(n22387),.clk(gclk));
	jnot g22130(.din(w_n22000_0[0]),.dout(n22388),.clk(gclk));
	jnot g22131(.din(w_n21993_0[0]),.dout(n22389),.clk(gclk));
	jnot g22132(.din(w_n21986_0[0]),.dout(n22390),.clk(gclk));
	jnot g22133(.din(w_n21979_0[0]),.dout(n22391),.clk(gclk));
	jnot g22134(.din(w_n21971_0[0]),.dout(n22392),.clk(gclk));
	jnot g22135(.din(w_n21964_0[0]),.dout(n22393),.clk(gclk));
	jnot g22136(.din(w_n21957_0[0]),.dout(n22394),.clk(gclk));
	jnot g22137(.din(w_n21950_0[0]),.dout(n22395),.clk(gclk));
	jnot g22138(.din(w_n21942_0[0]),.dout(n22396),.clk(gclk));
	jnot g22139(.din(w_n21935_0[0]),.dout(n22397),.clk(gclk));
	jnot g22140(.din(w_n21927_0[0]),.dout(n22398),.clk(gclk));
	jnot g22141(.din(w_n21920_0[0]),.dout(n22399),.clk(gclk));
	jnot g22142(.din(w_n21912_0[0]),.dout(n22400),.clk(gclk));
	jnot g22143(.din(w_n21903_0[0]),.dout(n22401),.clk(gclk));
	jnot g22144(.din(w_n21895_0[0]),.dout(n22402),.clk(gclk));
	jand g22145(.dina(w_asqrt5_2[2]),.dinb(w_a10_0[0]),.dout(n22403),.clk(gclk));
	jor g22146(.dina(w_n21892_0[0]),.dinb(n22403),.dout(n22404),.clk(gclk));
	jor g22147(.dina(n22404),.dinb(w_asqrt6_12[1]),.dout(n22405),.clk(gclk));
	jand g22148(.dina(w_asqrt5_2[1]),.dinb(w_n20907_0[2]),.dout(n22406),.clk(gclk));
	jor g22149(.dina(n22406),.dinb(w_n20908_0[0]),.dout(n22407),.clk(gclk));
	jand g22150(.dina(w_n21906_0[0]),.dinb(n22407),.dout(n22408),.clk(gclk));
	jand g22151(.dina(w_n22408_0[1]),.dinb(n22405),.dout(n22409),.clk(gclk));
	jor g22152(.dina(n22409),.dinb(n22402),.dout(n22410),.clk(gclk));
	jor g22153(.dina(n22410),.dinb(w_asqrt7_3[2]),.dout(n22411),.clk(gclk));
	jnot g22154(.din(w_n21909_0[0]),.dout(n22412),.clk(gclk));
	jand g22155(.dina(w_n22412_0[1]),.dinb(n22411),.dout(n22413),.clk(gclk));
	jor g22156(.dina(n22413),.dinb(n22401),.dout(n22414),.clk(gclk));
	jor g22157(.dina(n22414),.dinb(w_asqrt8_12[1]),.dout(n22415),.clk(gclk));
	jand g22158(.dina(w_n21916_0[1]),.dinb(n22415),.dout(n22416),.clk(gclk));
	jor g22159(.dina(n22416),.dinb(n22400),.dout(n22417),.clk(gclk));
	jor g22160(.dina(n22417),.dinb(w_asqrt9_4[1]),.dout(n22418),.clk(gclk));
	jnot g22161(.din(w_n21924_0[1]),.dout(n22419),.clk(gclk));
	jand g22162(.dina(n22419),.dinb(n22418),.dout(n22420),.clk(gclk));
	jor g22163(.dina(n22420),.dinb(n22399),.dout(n22421),.clk(gclk));
	jor g22164(.dina(n22421),.dinb(w_asqrt10_12[1]),.dout(n22422),.clk(gclk));
	jand g22165(.dina(w_n21931_0[1]),.dinb(n22422),.dout(n22423),.clk(gclk));
	jor g22166(.dina(n22423),.dinb(n22398),.dout(n22424),.clk(gclk));
	jor g22167(.dina(n22424),.dinb(w_asqrt11_4[1]),.dout(n22425),.clk(gclk));
	jnot g22168(.din(w_n21939_0[1]),.dout(n22426),.clk(gclk));
	jand g22169(.dina(n22426),.dinb(n22425),.dout(n22427),.clk(gclk));
	jor g22170(.dina(n22427),.dinb(n22397),.dout(n22428),.clk(gclk));
	jor g22171(.dina(n22428),.dinb(w_asqrt12_12[2]),.dout(n22429),.clk(gclk));
	jand g22172(.dina(w_n21946_0[1]),.dinb(n22429),.dout(n22430),.clk(gclk));
	jor g22173(.dina(n22430),.dinb(n22396),.dout(n22431),.clk(gclk));
	jor g22174(.dina(n22431),.dinb(w_asqrt13_5[0]),.dout(n22432),.clk(gclk));
	jnot g22175(.din(w_n21954_0[1]),.dout(n22433),.clk(gclk));
	jand g22176(.dina(n22433),.dinb(n22432),.dout(n22434),.clk(gclk));
	jor g22177(.dina(n22434),.dinb(n22395),.dout(n22435),.clk(gclk));
	jor g22178(.dina(n22435),.dinb(w_asqrt14_13[0]),.dout(n22436),.clk(gclk));
	jnot g22179(.din(w_n21961_0[1]),.dout(n22437),.clk(gclk));
	jand g22180(.dina(n22437),.dinb(n22436),.dout(n22438),.clk(gclk));
	jor g22181(.dina(n22438),.dinb(n22394),.dout(n22439),.clk(gclk));
	jor g22182(.dina(n22439),.dinb(w_asqrt15_5[2]),.dout(n22440),.clk(gclk));
	jnot g22183(.din(w_n21968_0[1]),.dout(n22441),.clk(gclk));
	jand g22184(.dina(n22441),.dinb(n22440),.dout(n22442),.clk(gclk));
	jor g22185(.dina(n22442),.dinb(n22393),.dout(n22443),.clk(gclk));
	jor g22186(.dina(n22443),.dinb(w_asqrt16_13[0]),.dout(n22444),.clk(gclk));
	jand g22187(.dina(w_n21975_0[1]),.dinb(n22444),.dout(n22445),.clk(gclk));
	jor g22188(.dina(n22445),.dinb(n22392),.dout(n22446),.clk(gclk));
	jor g22189(.dina(n22446),.dinb(w_asqrt17_6[0]),.dout(n22447),.clk(gclk));
	jnot g22190(.din(w_n21983_0[1]),.dout(n22448),.clk(gclk));
	jand g22191(.dina(n22448),.dinb(n22447),.dout(n22449),.clk(gclk));
	jor g22192(.dina(n22449),.dinb(n22391),.dout(n22450),.clk(gclk));
	jor g22193(.dina(n22450),.dinb(w_asqrt18_13[1]),.dout(n22451),.clk(gclk));
	jnot g22194(.din(w_n21990_0[1]),.dout(n22452),.clk(gclk));
	jand g22195(.dina(n22452),.dinb(n22451),.dout(n22453),.clk(gclk));
	jor g22196(.dina(n22453),.dinb(n22390),.dout(n22454),.clk(gclk));
	jor g22197(.dina(n22454),.dinb(w_asqrt19_6[1]),.dout(n22455),.clk(gclk));
	jnot g22198(.din(w_n21997_0[1]),.dout(n22456),.clk(gclk));
	jand g22199(.dina(n22456),.dinb(n22455),.dout(n22457),.clk(gclk));
	jor g22200(.dina(n22457),.dinb(n22389),.dout(n22458),.clk(gclk));
	jor g22201(.dina(n22458),.dinb(w_asqrt20_13[1]),.dout(n22459),.clk(gclk));
	jand g22202(.dina(w_n22004_0[1]),.dinb(n22459),.dout(n22460),.clk(gclk));
	jor g22203(.dina(n22460),.dinb(n22388),.dout(n22461),.clk(gclk));
	jor g22204(.dina(n22461),.dinb(w_asqrt21_7[0]),.dout(n22462),.clk(gclk));
	jnot g22205(.din(w_n22012_0[1]),.dout(n22463),.clk(gclk));
	jand g22206(.dina(n22463),.dinb(n22462),.dout(n22464),.clk(gclk));
	jor g22207(.dina(n22464),.dinb(n22387),.dout(n22465),.clk(gclk));
	jor g22208(.dina(n22465),.dinb(w_asqrt22_13[2]),.dout(n22466),.clk(gclk));
	jand g22209(.dina(w_n22019_0[1]),.dinb(n22466),.dout(n22467),.clk(gclk));
	jor g22210(.dina(n22467),.dinb(n22386),.dout(n22468),.clk(gclk));
	jor g22211(.dina(n22468),.dinb(w_asqrt23_7[2]),.dout(n22469),.clk(gclk));
	jnot g22212(.din(w_n22027_0[1]),.dout(n22470),.clk(gclk));
	jand g22213(.dina(n22470),.dinb(n22469),.dout(n22471),.clk(gclk));
	jor g22214(.dina(n22471),.dinb(n22385),.dout(n22472),.clk(gclk));
	jor g22215(.dina(n22472),.dinb(w_asqrt24_13[2]),.dout(n22473),.clk(gclk));
	jand g22216(.dina(w_n22034_0[1]),.dinb(n22473),.dout(n22474),.clk(gclk));
	jor g22217(.dina(n22474),.dinb(n22384),.dout(n22475),.clk(gclk));
	jor g22218(.dina(n22475),.dinb(w_asqrt25_7[2]),.dout(n22476),.clk(gclk));
	jnot g22219(.din(w_n22042_0[1]),.dout(n22477),.clk(gclk));
	jand g22220(.dina(n22477),.dinb(n22476),.dout(n22478),.clk(gclk));
	jor g22221(.dina(n22478),.dinb(n22383),.dout(n22479),.clk(gclk));
	jor g22222(.dina(n22479),.dinb(w_asqrt26_13[2]),.dout(n22480),.clk(gclk));
	jnot g22223(.din(w_n22049_0[1]),.dout(n22481),.clk(gclk));
	jand g22224(.dina(n22481),.dinb(n22480),.dout(n22482),.clk(gclk));
	jor g22225(.dina(n22482),.dinb(n22382),.dout(n22483),.clk(gclk));
	jor g22226(.dina(n22483),.dinb(w_asqrt27_8[1]),.dout(n22484),.clk(gclk));
	jand g22227(.dina(w_n22056_0[1]),.dinb(n22484),.dout(n22485),.clk(gclk));
	jor g22228(.dina(n22485),.dinb(n22381),.dout(n22486),.clk(gclk));
	jor g22229(.dina(n22486),.dinb(w_asqrt28_14[0]),.dout(n22487),.clk(gclk));
	jand g22230(.dina(w_n22064_0[1]),.dinb(n22487),.dout(n22488),.clk(gclk));
	jor g22231(.dina(n22488),.dinb(n22380),.dout(n22489),.clk(gclk));
	jor g22232(.dina(n22489),.dinb(w_asqrt29_8[2]),.dout(n22490),.clk(gclk));
	jnot g22233(.din(w_n22072_0[1]),.dout(n22491),.clk(gclk));
	jand g22234(.dina(n22491),.dinb(n22490),.dout(n22492),.clk(gclk));
	jor g22235(.dina(n22492),.dinb(n22379),.dout(n22493),.clk(gclk));
	jor g22236(.dina(n22493),.dinb(w_asqrt30_14[1]),.dout(n22494),.clk(gclk));
	jand g22237(.dina(w_n22079_0[1]),.dinb(n22494),.dout(n22495),.clk(gclk));
	jor g22238(.dina(n22495),.dinb(n22378),.dout(n22496),.clk(gclk));
	jor g22239(.dina(n22496),.dinb(w_asqrt31_9[1]),.dout(n22497),.clk(gclk));
	jnot g22240(.din(w_n22087_0[1]),.dout(n22498),.clk(gclk));
	jand g22241(.dina(n22498),.dinb(n22497),.dout(n22499),.clk(gclk));
	jor g22242(.dina(n22499),.dinb(n22377),.dout(n22500),.clk(gclk));
	jor g22243(.dina(n22500),.dinb(w_asqrt32_14[1]),.dout(n22501),.clk(gclk));
	jand g22244(.dina(w_n22094_0[1]),.dinb(n22501),.dout(n22502),.clk(gclk));
	jor g22245(.dina(n22502),.dinb(n22376),.dout(n22503),.clk(gclk));
	jor g22246(.dina(n22503),.dinb(w_asqrt33_10[0]),.dout(n22504),.clk(gclk));
	jnot g22247(.din(w_n22102_0[1]),.dout(n22505),.clk(gclk));
	jand g22248(.dina(n22505),.dinb(n22504),.dout(n22506),.clk(gclk));
	jor g22249(.dina(n22506),.dinb(n22375),.dout(n22507),.clk(gclk));
	jor g22250(.dina(n22507),.dinb(w_asqrt34_14[2]),.dout(n22508),.clk(gclk));
	jnot g22251(.din(w_n22109_0[1]),.dout(n22509),.clk(gclk));
	jand g22252(.dina(n22509),.dinb(n22508),.dout(n22510),.clk(gclk));
	jor g22253(.dina(n22510),.dinb(n22374),.dout(n22511),.clk(gclk));
	jor g22254(.dina(n22511),.dinb(w_asqrt35_10[2]),.dout(n22512),.clk(gclk));
	jnot g22255(.din(w_n22116_0[1]),.dout(n22513),.clk(gclk));
	jand g22256(.dina(n22513),.dinb(n22512),.dout(n22514),.clk(gclk));
	jor g22257(.dina(n22514),.dinb(n22373),.dout(n22515),.clk(gclk));
	jor g22258(.dina(n22515),.dinb(w_asqrt36_14[2]),.dout(n22516),.clk(gclk));
	jand g22259(.dina(w_n22123_0[1]),.dinb(n22516),.dout(n22517),.clk(gclk));
	jor g22260(.dina(n22517),.dinb(n22372),.dout(n22518),.clk(gclk));
	jor g22261(.dina(n22518),.dinb(w_asqrt37_11[0]),.dout(n22519),.clk(gclk));
	jnot g22262(.din(w_n22131_0[1]),.dout(n22520),.clk(gclk));
	jand g22263(.dina(n22520),.dinb(n22519),.dout(n22521),.clk(gclk));
	jor g22264(.dina(n22521),.dinb(n22371),.dout(n22522),.clk(gclk));
	jor g22265(.dina(n22522),.dinb(w_asqrt38_15[0]),.dout(n22523),.clk(gclk));
	jand g22266(.dina(w_n22138_0[1]),.dinb(n22523),.dout(n22524),.clk(gclk));
	jor g22267(.dina(n22524),.dinb(n22370),.dout(n22525),.clk(gclk));
	jor g22268(.dina(n22525),.dinb(w_asqrt39_11[2]),.dout(n22526),.clk(gclk));
	jnot g22269(.din(w_n22146_0[1]),.dout(n22527),.clk(gclk));
	jand g22270(.dina(n22527),.dinb(n22526),.dout(n22528),.clk(gclk));
	jor g22271(.dina(n22528),.dinb(n22369),.dout(n22529),.clk(gclk));
	jor g22272(.dina(n22529),.dinb(w_asqrt40_15[0]),.dout(n22530),.clk(gclk));
	jand g22273(.dina(w_n22153_0[1]),.dinb(n22530),.dout(n22531),.clk(gclk));
	jor g22274(.dina(n22531),.dinb(n22368),.dout(n22532),.clk(gclk));
	jor g22275(.dina(n22532),.dinb(w_asqrt41_12[0]),.dout(n22533),.clk(gclk));
	jnot g22276(.din(w_n22161_0[1]),.dout(n22534),.clk(gclk));
	jand g22277(.dina(n22534),.dinb(n22533),.dout(n22535),.clk(gclk));
	jor g22278(.dina(n22535),.dinb(n22367),.dout(n22536),.clk(gclk));
	jor g22279(.dina(n22536),.dinb(w_asqrt42_15[1]),.dout(n22537),.clk(gclk));
	jand g22280(.dina(w_n22168_0[1]),.dinb(n22537),.dout(n22538),.clk(gclk));
	jor g22281(.dina(n22538),.dinb(n22366),.dout(n22539),.clk(gclk));
	jor g22282(.dina(n22539),.dinb(w_asqrt43_12[1]),.dout(n22540),.clk(gclk));
	jnot g22283(.din(w_n22176_0[1]),.dout(n22541),.clk(gclk));
	jand g22284(.dina(n22541),.dinb(n22540),.dout(n22542),.clk(gclk));
	jor g22285(.dina(n22542),.dinb(n22365),.dout(n22543),.clk(gclk));
	jor g22286(.dina(n22543),.dinb(w_asqrt44_15[1]),.dout(n22544),.clk(gclk));
	jnot g22287(.din(w_n22183_0[1]),.dout(n22545),.clk(gclk));
	jand g22288(.dina(n22545),.dinb(n22544),.dout(n22546),.clk(gclk));
	jor g22289(.dina(n22546),.dinb(n22364),.dout(n22547),.clk(gclk));
	jor g22290(.dina(n22547),.dinb(w_asqrt45_13[0]),.dout(n22548),.clk(gclk));
	jnot g22291(.din(w_n22190_0[1]),.dout(n22549),.clk(gclk));
	jand g22292(.dina(n22549),.dinb(n22548),.dout(n22550),.clk(gclk));
	jor g22293(.dina(n22550),.dinb(n22363),.dout(n22551),.clk(gclk));
	jor g22294(.dina(n22551),.dinb(w_asqrt46_15[1]),.dout(n22552),.clk(gclk));
	jand g22295(.dina(w_n22197_0[1]),.dinb(n22552),.dout(n22553),.clk(gclk));
	jor g22296(.dina(n22553),.dinb(n22362),.dout(n22554),.clk(gclk));
	jor g22297(.dina(n22554),.dinb(w_asqrt47_13[2]),.dout(n22555),.clk(gclk));
	jnot g22298(.din(w_n22205_0[1]),.dout(n22556),.clk(gclk));
	jand g22299(.dina(n22556),.dinb(n22555),.dout(n22557),.clk(gclk));
	jor g22300(.dina(n22557),.dinb(n22361),.dout(n22558),.clk(gclk));
	jor g22301(.dina(n22558),.dinb(w_asqrt48_15[2]),.dout(n22559),.clk(gclk));
	jnot g22302(.din(w_n22212_0[1]),.dout(n22560),.clk(gclk));
	jand g22303(.dina(n22560),.dinb(n22559),.dout(n22561),.clk(gclk));
	jor g22304(.dina(n22561),.dinb(n22360),.dout(n22562),.clk(gclk));
	jor g22305(.dina(n22562),.dinb(w_asqrt49_14[0]),.dout(n22563),.clk(gclk));
	jnot g22306(.din(w_n22219_0[1]),.dout(n22564),.clk(gclk));
	jand g22307(.dina(n22564),.dinb(n22563),.dout(n22565),.clk(gclk));
	jor g22308(.dina(n22565),.dinb(n22359),.dout(n22566),.clk(gclk));
	jor g22309(.dina(n22566),.dinb(w_asqrt50_16[0]),.dout(n22567),.clk(gclk));
	jnot g22310(.din(w_n22226_0[1]),.dout(n22568),.clk(gclk));
	jand g22311(.dina(n22568),.dinb(n22567),.dout(n22569),.clk(gclk));
	jor g22312(.dina(n22569),.dinb(n22358),.dout(n22570),.clk(gclk));
	jor g22313(.dina(n22570),.dinb(w_asqrt51_14[1]),.dout(n22571),.clk(gclk));
	jnot g22314(.din(w_n22233_0[1]),.dout(n22572),.clk(gclk));
	jand g22315(.dina(n22572),.dinb(n22571),.dout(n22573),.clk(gclk));
	jor g22316(.dina(n22573),.dinb(n22357),.dout(n22574),.clk(gclk));
	jor g22317(.dina(n22574),.dinb(w_asqrt52_16[0]),.dout(n22575),.clk(gclk));
	jand g22318(.dina(w_n22240_0[1]),.dinb(n22575),.dout(n22576),.clk(gclk));
	jor g22319(.dina(n22576),.dinb(n22356),.dout(n22577),.clk(gclk));
	jor g22320(.dina(n22577),.dinb(w_asqrt53_15[0]),.dout(n22578),.clk(gclk));
	jnot g22321(.din(w_n22248_0[1]),.dout(n22579),.clk(gclk));
	jand g22322(.dina(n22579),.dinb(n22578),.dout(n22580),.clk(gclk));
	jor g22323(.dina(n22580),.dinb(n22355),.dout(n22581),.clk(gclk));
	jor g22324(.dina(n22581),.dinb(w_asqrt54_16[0]),.dout(n22582),.clk(gclk));
	jand g22325(.dina(w_n22255_0[1]),.dinb(n22582),.dout(n22583),.clk(gclk));
	jor g22326(.dina(n22583),.dinb(n22354),.dout(n22584),.clk(gclk));
	jor g22327(.dina(n22584),.dinb(w_asqrt55_15[1]),.dout(n22585),.clk(gclk));
	jnot g22328(.din(w_n22263_0[1]),.dout(n22586),.clk(gclk));
	jand g22329(.dina(n22586),.dinb(n22585),.dout(n22587),.clk(gclk));
	jor g22330(.dina(n22587),.dinb(n22353),.dout(n22588),.clk(gclk));
	jor g22331(.dina(n22588),.dinb(w_asqrt56_16[1]),.dout(n22589),.clk(gclk));
	jnot g22332(.din(w_n22270_0[1]),.dout(n22590),.clk(gclk));
	jand g22333(.dina(n22590),.dinb(n22589),.dout(n22591),.clk(gclk));
	jor g22334(.dina(n22591),.dinb(n22352),.dout(n22592),.clk(gclk));
	jor g22335(.dina(n22592),.dinb(w_asqrt57_16[0]),.dout(n22593),.clk(gclk));
	jand g22336(.dina(w_n22277_0[1]),.dinb(n22593),.dout(n22594),.clk(gclk));
	jor g22337(.dina(n22594),.dinb(n22351),.dout(n22595),.clk(gclk));
	jor g22338(.dina(n22595),.dinb(w_asqrt58_16[2]),.dout(n22596),.clk(gclk));
	jand g22339(.dina(w_n22285_0[1]),.dinb(n22596),.dout(n22597),.clk(gclk));
	jor g22340(.dina(n22597),.dinb(n22350),.dout(n22598),.clk(gclk));
	jor g22341(.dina(n22598),.dinb(w_asqrt59_16[1]),.dout(n22599),.clk(gclk));
	jnot g22342(.din(w_n22293_0[1]),.dout(n22600),.clk(gclk));
	jand g22343(.dina(n22600),.dinb(n22599),.dout(n22601),.clk(gclk));
	jor g22344(.dina(n22601),.dinb(n22349),.dout(n22602),.clk(gclk));
	jor g22345(.dina(n22602),.dinb(w_asqrt60_16[2]),.dout(n22603),.clk(gclk));
	jnot g22346(.din(w_n22300_0[1]),.dout(n22604),.clk(gclk));
	jand g22347(.dina(n22604),.dinb(n22603),.dout(n22605),.clk(gclk));
	jor g22348(.dina(n22605),.dinb(n22348),.dout(n22606),.clk(gclk));
	jor g22349(.dina(n22606),.dinb(w_asqrt61_16[2]),.dout(n22607),.clk(gclk));
	jnot g22350(.din(w_n22307_0[1]),.dout(n22608),.clk(gclk));
	jand g22351(.dina(n22608),.dinb(n22607),.dout(n22609),.clk(gclk));
	jor g22352(.dina(n22609),.dinb(n22347),.dout(n22610),.clk(gclk));
	jor g22353(.dina(n22610),.dinb(w_asqrt62_16[2]),.dout(n22611),.clk(gclk));
	jand g22354(.dina(w_n22314_0[0]),.dinb(n22611),.dout(n22612),.clk(gclk));
	jor g22355(.dina(n22612),.dinb(n22346),.dout(n22613),.clk(gclk));
	jnot g22356(.din(w_n22320_0[2]),.dout(n22614),.clk(gclk));
	jand g22357(.dina(n22614),.dinb(n22613),.dout(n22615),.clk(gclk));
	jnot g22358(.din(w_n22325_0[0]),.dout(n22616),.clk(gclk));
	jand g22359(.dina(n22616),.dinb(w_n22615_0[1]),.dout(n22617),.clk(gclk));
	jor g22360(.dina(n22617),.dinb(w_asqrt63_20[2]),.dout(n22618),.clk(gclk));
	jand g22361(.dina(w_n22330_0[0]),.dinb(n22618),.dout(n22619),.clk(gclk));
	jand g22362(.dina(w_n22619_0[1]),.dinb(w_n22345_0[1]),.dout(n22620),.clk(gclk));
	jor g22363(.dina(w_n22620_4[2]),.dinb(n22344),.dout(n22621),.clk(gclk));
	jand g22364(.dina(w_n22621_0[1]),.dinb(n22343),.dout(n22622),.clk(gclk));
	jand g22365(.dina(w_n22622_0[1]),.dinb(n22341),.dout(n22623),.clk(gclk));
	jor g22366(.dina(n22623),.dinb(w_n22340_0[1]),.dout(n22624),.clk(gclk));
	jand g22367(.dina(w_n22624_0[2]),.dinb(w_asqrt6_12[0]),.dout(n22625),.clk(gclk));
	jor g22368(.dina(w_n22624_0[1]),.dinb(w_asqrt6_11[2]),.dout(n22626),.clk(gclk));
	jor g22369(.dina(w_asqrt4_30[2]),.dinb(w_n21887_14[1]),.dout(n22627),.clk(gclk));
	jand g22370(.dina(n22627),.dinb(w_n22621_0[0]),.dout(n22628),.clk(gclk));
	jxor g22371(.dina(n22628),.dinb(w_n20907_0[1]),.dout(n22629),.clk(gclk));
	jnot g22372(.din(w_n22629_0[1]),.dout(n22630),.clk(gclk));
	jand g22373(.dina(w_n22630_0[1]),.dinb(n22626),.dout(n22631),.clk(gclk));
	jor g22374(.dina(n22631),.dinb(w_n22625_0[1]),.dout(n22632),.clk(gclk));
	jand g22375(.dina(w_n22632_0[2]),.dinb(w_asqrt7_3[1]),.dout(n22633),.clk(gclk));
	jor g22376(.dina(w_n22632_0[1]),.dinb(w_asqrt7_3[0]),.dout(n22634),.clk(gclk));
	jxor g22377(.dina(w_n21894_0[0]),.dinb(w_n21184_5[1]),.dout(n22635),.clk(gclk));
	jand g22378(.dina(n22635),.dinb(w_asqrt4_30[1]),.dout(n22636),.clk(gclk));
	jxor g22379(.dina(n22636),.dinb(w_n22408_0[0]),.dout(n22637),.clk(gclk));
	jand g22380(.dina(w_n22637_0[1]),.dinb(n22634),.dout(n22638),.clk(gclk));
	jor g22381(.dina(n22638),.dinb(w_n22633_0[1]),.dout(n22639),.clk(gclk));
	jand g22382(.dina(w_n22639_0[2]),.dinb(w_asqrt8_12[0]),.dout(n22640),.clk(gclk));
	jor g22383(.dina(w_n22639_0[1]),.dinb(w_asqrt8_11[2]),.dout(n22641),.clk(gclk));
	jxor g22384(.dina(w_n21902_0[0]),.dinb(w_n20468_14[2]),.dout(n22642),.clk(gclk));
	jand g22385(.dina(n22642),.dinb(w_asqrt4_30[0]),.dout(n22643),.clk(gclk));
	jxor g22386(.dina(n22643),.dinb(w_n22412_0[0]),.dout(n22644),.clk(gclk));
	jand g22387(.dina(w_n22644_0[1]),.dinb(n22641),.dout(n22645),.clk(gclk));
	jor g22388(.dina(n22645),.dinb(w_n22640_0[1]),.dout(n22646),.clk(gclk));
	jand g22389(.dina(w_n22646_0[2]),.dinb(w_asqrt9_4[0]),.dout(n22647),.clk(gclk));
	jor g22390(.dina(w_n22646_0[1]),.dinb(w_asqrt9_3[2]),.dout(n22648),.clk(gclk));
	jxor g22391(.dina(w_n21911_0[0]),.dinb(w_n19791_6[1]),.dout(n22649),.clk(gclk));
	jand g22392(.dina(n22649),.dinb(w_asqrt4_29[2]),.dout(n22650),.clk(gclk));
	jxor g22393(.dina(n22650),.dinb(w_n21916_0[0]),.dout(n22651),.clk(gclk));
	jand g22394(.dina(w_n22651_0[1]),.dinb(n22648),.dout(n22652),.clk(gclk));
	jor g22395(.dina(n22652),.dinb(w_n22647_0[1]),.dout(n22653),.clk(gclk));
	jand g22396(.dina(w_n22653_0[2]),.dinb(w_asqrt10_12[0]),.dout(n22654),.clk(gclk));
	jor g22397(.dina(w_n22653_0[1]),.dinb(w_asqrt10_11[2]),.dout(n22655),.clk(gclk));
	jxor g22398(.dina(w_n21919_0[0]),.dinb(w_n19096_15[0]),.dout(n22656),.clk(gclk));
	jand g22399(.dina(n22656),.dinb(w_asqrt4_29[1]),.dout(n22657),.clk(gclk));
	jxor g22400(.dina(n22657),.dinb(w_n21924_0[0]),.dout(n22658),.clk(gclk));
	jnot g22401(.din(w_n22658_0[1]),.dout(n22659),.clk(gclk));
	jand g22402(.dina(w_n22659_0[1]),.dinb(n22655),.dout(n22660),.clk(gclk));
	jor g22403(.dina(n22660),.dinb(w_n22654_0[1]),.dout(n22661),.clk(gclk));
	jand g22404(.dina(w_n22661_0[2]),.dinb(w_asqrt11_4[0]),.dout(n22662),.clk(gclk));
	jor g22405(.dina(w_n22661_0[1]),.dinb(w_asqrt11_3[2]),.dout(n22663),.clk(gclk));
	jxor g22406(.dina(w_n21926_0[0]),.dinb(w_n18442_7[0]),.dout(n22664),.clk(gclk));
	jand g22407(.dina(n22664),.dinb(w_asqrt4_29[0]),.dout(n22665),.clk(gclk));
	jxor g22408(.dina(n22665),.dinb(w_n21931_0[0]),.dout(n22666),.clk(gclk));
	jand g22409(.dina(w_n22666_0[1]),.dinb(n22663),.dout(n22667),.clk(gclk));
	jor g22410(.dina(n22667),.dinb(w_n22662_0[1]),.dout(n22668),.clk(gclk));
	jand g22411(.dina(w_n22668_0[2]),.dinb(w_asqrt12_12[1]),.dout(n22669),.clk(gclk));
	jor g22412(.dina(w_n22668_0[1]),.dinb(w_asqrt12_12[0]),.dout(n22670),.clk(gclk));
	jxor g22413(.dina(w_n21934_0[0]),.dinb(w_n17769_15[2]),.dout(n22671),.clk(gclk));
	jand g22414(.dina(n22671),.dinb(w_asqrt4_28[2]),.dout(n22672),.clk(gclk));
	jxor g22415(.dina(n22672),.dinb(w_n21939_0[0]),.dout(n22673),.clk(gclk));
	jnot g22416(.din(w_n22673_0[1]),.dout(n22674),.clk(gclk));
	jand g22417(.dina(w_n22674_0[1]),.dinb(n22670),.dout(n22675),.clk(gclk));
	jor g22418(.dina(n22675),.dinb(w_n22669_0[1]),.dout(n22676),.clk(gclk));
	jand g22419(.dina(w_n22676_0[2]),.dinb(w_asqrt13_4[2]),.dout(n22677),.clk(gclk));
	jor g22420(.dina(w_n22676_0[1]),.dinb(w_asqrt13_4[1]),.dout(n22678),.clk(gclk));
	jxor g22421(.dina(w_n21941_0[0]),.dinb(w_n17134_8[0]),.dout(n22679),.clk(gclk));
	jand g22422(.dina(n22679),.dinb(w_asqrt4_28[1]),.dout(n22680),.clk(gclk));
	jxor g22423(.dina(n22680),.dinb(w_n21946_0[0]),.dout(n22681),.clk(gclk));
	jand g22424(.dina(w_n22681_0[1]),.dinb(n22678),.dout(n22682),.clk(gclk));
	jor g22425(.dina(n22682),.dinb(w_n22677_0[1]),.dout(n22683),.clk(gclk));
	jand g22426(.dina(w_n22683_0[2]),.dinb(w_asqrt14_12[2]),.dout(n22684),.clk(gclk));
	jor g22427(.dina(w_n22683_0[1]),.dinb(w_asqrt14_12[1]),.dout(n22685),.clk(gclk));
	jxor g22428(.dina(w_n21949_0[0]),.dinb(w_n16489_16[0]),.dout(n22686),.clk(gclk));
	jand g22429(.dina(n22686),.dinb(w_asqrt4_28[0]),.dout(n22687),.clk(gclk));
	jxor g22430(.dina(n22687),.dinb(w_n21954_0[0]),.dout(n22688),.clk(gclk));
	jnot g22431(.din(w_n22688_0[1]),.dout(n22689),.clk(gclk));
	jand g22432(.dina(w_n22689_0[1]),.dinb(n22685),.dout(n22690),.clk(gclk));
	jor g22433(.dina(n22690),.dinb(w_n22684_0[1]),.dout(n22691),.clk(gclk));
	jand g22434(.dina(w_n22691_0[2]),.dinb(w_asqrt15_5[1]),.dout(n22692),.clk(gclk));
	jor g22435(.dina(w_n22691_0[1]),.dinb(w_asqrt15_5[0]),.dout(n22693),.clk(gclk));
	jxor g22436(.dina(w_n21956_0[0]),.dinb(w_n15878_9[0]),.dout(n22694),.clk(gclk));
	jand g22437(.dina(n22694),.dinb(w_asqrt4_27[2]),.dout(n22695),.clk(gclk));
	jxor g22438(.dina(n22695),.dinb(w_n21961_0[0]),.dout(n22696),.clk(gclk));
	jnot g22439(.din(w_n22696_0[1]),.dout(n22697),.clk(gclk));
	jand g22440(.dina(w_n22697_0[1]),.dinb(n22693),.dout(n22698),.clk(gclk));
	jor g22441(.dina(n22698),.dinb(w_n22692_0[1]),.dout(n22699),.clk(gclk));
	jand g22442(.dina(w_n22699_0[2]),.dinb(w_asqrt16_12[2]),.dout(n22700),.clk(gclk));
	jor g22443(.dina(w_n22699_0[1]),.dinb(w_asqrt16_12[1]),.dout(n22701),.clk(gclk));
	jxor g22444(.dina(w_n21963_0[0]),.dinb(w_n15260_16[2]),.dout(n22702),.clk(gclk));
	jand g22445(.dina(n22702),.dinb(w_asqrt4_27[1]),.dout(n22703),.clk(gclk));
	jxor g22446(.dina(n22703),.dinb(w_n21968_0[0]),.dout(n22704),.clk(gclk));
	jnot g22447(.din(w_n22704_0[1]),.dout(n22705),.clk(gclk));
	jand g22448(.dina(w_n22705_0[1]),.dinb(n22701),.dout(n22706),.clk(gclk));
	jor g22449(.dina(n22706),.dinb(w_n22700_0[1]),.dout(n22707),.clk(gclk));
	jand g22450(.dina(w_n22707_0[2]),.dinb(w_asqrt17_5[2]),.dout(n22708),.clk(gclk));
	jor g22451(.dina(w_n22707_0[1]),.dinb(w_asqrt17_5[1]),.dout(n22709),.clk(gclk));
	jxor g22452(.dina(w_n21970_0[0]),.dinb(w_n14674_9[2]),.dout(n22710),.clk(gclk));
	jand g22453(.dina(n22710),.dinb(w_asqrt4_27[0]),.dout(n22711),.clk(gclk));
	jxor g22454(.dina(n22711),.dinb(w_n21975_0[0]),.dout(n22712),.clk(gclk));
	jand g22455(.dina(w_n22712_0[1]),.dinb(n22709),.dout(n22713),.clk(gclk));
	jor g22456(.dina(n22713),.dinb(w_n22708_0[1]),.dout(n22714),.clk(gclk));
	jand g22457(.dina(w_n22714_0[2]),.dinb(w_asqrt18_13[0]),.dout(n22715),.clk(gclk));
	jor g22458(.dina(w_n22714_0[1]),.dinb(w_asqrt18_12[2]),.dout(n22716),.clk(gclk));
	jxor g22459(.dina(w_n21978_0[0]),.dinb(w_n14078_17[0]),.dout(n22717),.clk(gclk));
	jand g22460(.dina(n22717),.dinb(w_asqrt4_26[2]),.dout(n22718),.clk(gclk));
	jxor g22461(.dina(n22718),.dinb(w_n21983_0[0]),.dout(n22719),.clk(gclk));
	jnot g22462(.din(w_n22719_0[1]),.dout(n22720),.clk(gclk));
	jand g22463(.dina(w_n22720_0[1]),.dinb(n22716),.dout(n22721),.clk(gclk));
	jor g22464(.dina(n22721),.dinb(w_n22715_0[1]),.dout(n22722),.clk(gclk));
	jand g22465(.dina(w_n22722_0[2]),.dinb(w_asqrt19_6[0]),.dout(n22723),.clk(gclk));
	jor g22466(.dina(w_n22722_0[1]),.dinb(w_asqrt19_5[2]),.dout(n22724),.clk(gclk));
	jxor g22467(.dina(w_n21985_0[0]),.dinb(w_n13515_10[2]),.dout(n22725),.clk(gclk));
	jand g22468(.dina(n22725),.dinb(w_asqrt4_26[1]),.dout(n22726),.clk(gclk));
	jxor g22469(.dina(n22726),.dinb(w_n21990_0[0]),.dout(n22727),.clk(gclk));
	jnot g22470(.din(w_n22727_0[1]),.dout(n22728),.clk(gclk));
	jand g22471(.dina(w_n22728_0[1]),.dinb(n22724),.dout(n22729),.clk(gclk));
	jor g22472(.dina(n22729),.dinb(w_n22723_0[1]),.dout(n22730),.clk(gclk));
	jand g22473(.dina(w_n22730_0[2]),.dinb(w_asqrt20_13[0]),.dout(n22731),.clk(gclk));
	jor g22474(.dina(w_n22730_0[1]),.dinb(w_asqrt20_12[2]),.dout(n22732),.clk(gclk));
	jxor g22475(.dina(w_n21992_0[0]),.dinb(w_n12947_17[2]),.dout(n22733),.clk(gclk));
	jand g22476(.dina(n22733),.dinb(w_asqrt4_26[0]),.dout(n22734),.clk(gclk));
	jxor g22477(.dina(n22734),.dinb(w_n21997_0[0]),.dout(n22735),.clk(gclk));
	jnot g22478(.din(w_n22735_0[1]),.dout(n22736),.clk(gclk));
	jand g22479(.dina(w_n22736_0[1]),.dinb(n22732),.dout(n22737),.clk(gclk));
	jor g22480(.dina(n22737),.dinb(w_n22731_0[1]),.dout(n22738),.clk(gclk));
	jand g22481(.dina(w_n22738_0[2]),.dinb(w_asqrt21_6[2]),.dout(n22739),.clk(gclk));
	jor g22482(.dina(w_n22738_0[1]),.dinb(w_asqrt21_6[1]),.dout(n22740),.clk(gclk));
	jxor g22483(.dina(w_n21999_0[0]),.dinb(w_n12410_11[1]),.dout(n22741),.clk(gclk));
	jand g22484(.dina(n22741),.dinb(w_asqrt4_25[2]),.dout(n22742),.clk(gclk));
	jxor g22485(.dina(n22742),.dinb(w_n22004_0[0]),.dout(n22743),.clk(gclk));
	jand g22486(.dina(w_n22743_0[1]),.dinb(n22740),.dout(n22744),.clk(gclk));
	jor g22487(.dina(n22744),.dinb(w_n22739_0[1]),.dout(n22745),.clk(gclk));
	jand g22488(.dina(w_n22745_0[2]),.dinb(w_asqrt22_13[1]),.dout(n22746),.clk(gclk));
	jor g22489(.dina(w_n22745_0[1]),.dinb(w_asqrt22_13[0]),.dout(n22747),.clk(gclk));
	jxor g22490(.dina(w_n22007_0[0]),.dinb(w_n11858_18[0]),.dout(n22748),.clk(gclk));
	jand g22491(.dina(n22748),.dinb(w_asqrt4_25[1]),.dout(n22749),.clk(gclk));
	jxor g22492(.dina(n22749),.dinb(w_n22012_0[0]),.dout(n22750),.clk(gclk));
	jnot g22493(.din(w_n22750_0[1]),.dout(n22751),.clk(gclk));
	jand g22494(.dina(w_n22751_0[1]),.dinb(n22747),.dout(n22752),.clk(gclk));
	jor g22495(.dina(n22752),.dinb(w_n22746_0[1]),.dout(n22753),.clk(gclk));
	jand g22496(.dina(w_n22753_0[2]),.dinb(w_asqrt23_7[1]),.dout(n22754),.clk(gclk));
	jor g22497(.dina(w_n22753_0[1]),.dinb(w_asqrt23_7[0]),.dout(n22755),.clk(gclk));
	jxor g22498(.dina(w_n22014_0[0]),.dinb(w_n11347_12[0]),.dout(n22756),.clk(gclk));
	jand g22499(.dina(n22756),.dinb(w_asqrt4_25[0]),.dout(n22757),.clk(gclk));
	jxor g22500(.dina(n22757),.dinb(w_n22019_0[0]),.dout(n22758),.clk(gclk));
	jand g22501(.dina(w_n22758_0[1]),.dinb(n22755),.dout(n22759),.clk(gclk));
	jor g22502(.dina(n22759),.dinb(w_n22754_0[1]),.dout(n22760),.clk(gclk));
	jand g22503(.dina(w_n22760_0[2]),.dinb(w_asqrt24_13[1]),.dout(n22761),.clk(gclk));
	jor g22504(.dina(w_n22760_0[1]),.dinb(w_asqrt24_13[0]),.dout(n22762),.clk(gclk));
	jxor g22505(.dina(w_n22022_0[0]),.dinb(w_n10824_18[2]),.dout(n22763),.clk(gclk));
	jand g22506(.dina(n22763),.dinb(w_asqrt4_24[2]),.dout(n22764),.clk(gclk));
	jxor g22507(.dina(n22764),.dinb(w_n22027_0[0]),.dout(n22765),.clk(gclk));
	jnot g22508(.din(w_n22765_0[1]),.dout(n22766),.clk(gclk));
	jand g22509(.dina(w_n22766_0[1]),.dinb(n22762),.dout(n22767),.clk(gclk));
	jor g22510(.dina(n22767),.dinb(w_n22761_0[1]),.dout(n22768),.clk(gclk));
	jand g22511(.dina(w_n22768_0[2]),.dinb(w_asqrt25_7[1]),.dout(n22769),.clk(gclk));
	jor g22512(.dina(w_n22768_0[1]),.dinb(w_asqrt25_7[0]),.dout(n22770),.clk(gclk));
	jxor g22513(.dina(w_n22029_0[0]),.dinb(w_n10328_13[0]),.dout(n22771),.clk(gclk));
	jand g22514(.dina(n22771),.dinb(w_asqrt4_24[1]),.dout(n22772),.clk(gclk));
	jxor g22515(.dina(n22772),.dinb(w_n22034_0[0]),.dout(n22773),.clk(gclk));
	jand g22516(.dina(w_n22773_0[1]),.dinb(n22770),.dout(n22774),.clk(gclk));
	jor g22517(.dina(n22774),.dinb(w_n22769_0[1]),.dout(n22775),.clk(gclk));
	jand g22518(.dina(w_n22775_0[2]),.dinb(w_asqrt26_13[1]),.dout(n22776),.clk(gclk));
	jor g22519(.dina(w_n22775_0[1]),.dinb(w_asqrt26_13[0]),.dout(n22777),.clk(gclk));
	jxor g22520(.dina(w_n22037_0[0]),.dinb(w_n9832_19[1]),.dout(n22778),.clk(gclk));
	jand g22521(.dina(n22778),.dinb(w_asqrt4_24[0]),.dout(n22779),.clk(gclk));
	jxor g22522(.dina(n22779),.dinb(w_n22042_0[0]),.dout(n22780),.clk(gclk));
	jnot g22523(.din(w_n22780_0[1]),.dout(n22781),.clk(gclk));
	jand g22524(.dina(w_n22781_0[1]),.dinb(n22777),.dout(n22782),.clk(gclk));
	jor g22525(.dina(n22782),.dinb(w_n22776_0[1]),.dout(n22783),.clk(gclk));
	jand g22526(.dina(w_n22783_0[2]),.dinb(w_asqrt27_8[0]),.dout(n22784),.clk(gclk));
	jor g22527(.dina(w_n22783_0[1]),.dinb(w_asqrt27_7[2]),.dout(n22785),.clk(gclk));
	jxor g22528(.dina(w_n22044_0[0]),.dinb(w_n9369_14[0]),.dout(n22786),.clk(gclk));
	jand g22529(.dina(n22786),.dinb(w_asqrt4_23[2]),.dout(n22787),.clk(gclk));
	jxor g22530(.dina(n22787),.dinb(w_n22049_0[0]),.dout(n22788),.clk(gclk));
	jnot g22531(.din(w_n22788_0[1]),.dout(n22789),.clk(gclk));
	jand g22532(.dina(w_n22789_0[1]),.dinb(n22785),.dout(n22790),.clk(gclk));
	jor g22533(.dina(n22790),.dinb(w_n22784_0[1]),.dout(n22791),.clk(gclk));
	jand g22534(.dina(w_n22791_0[2]),.dinb(w_asqrt28_13[2]),.dout(n22792),.clk(gclk));
	jor g22535(.dina(w_n22791_0[1]),.dinb(w_asqrt28_13[1]),.dout(n22793),.clk(gclk));
	jxor g22536(.dina(w_n22051_0[0]),.dinb(w_n8890_19[2]),.dout(n22794),.clk(gclk));
	jand g22537(.dina(n22794),.dinb(w_asqrt4_23[1]),.dout(n22795),.clk(gclk));
	jxor g22538(.dina(n22795),.dinb(w_n22056_0[0]),.dout(n22796),.clk(gclk));
	jand g22539(.dina(w_n22796_0[1]),.dinb(n22793),.dout(n22797),.clk(gclk));
	jor g22540(.dina(n22797),.dinb(w_n22792_0[1]),.dout(n22798),.clk(gclk));
	jand g22541(.dina(w_n22798_0[2]),.dinb(w_asqrt29_8[1]),.dout(n22799),.clk(gclk));
	jor g22542(.dina(w_n22798_0[1]),.dinb(w_asqrt29_8[0]),.dout(n22800),.clk(gclk));
	jxor g22543(.dina(w_n22059_0[0]),.dinb(w_n8449_14[2]),.dout(n22801),.clk(gclk));
	jand g22544(.dina(n22801),.dinb(w_asqrt4_23[0]),.dout(n22802),.clk(gclk));
	jxor g22545(.dina(n22802),.dinb(w_n22064_0[0]),.dout(n22803),.clk(gclk));
	jand g22546(.dina(w_n22803_0[1]),.dinb(n22800),.dout(n22804),.clk(gclk));
	jor g22547(.dina(n22804),.dinb(w_n22799_0[1]),.dout(n22805),.clk(gclk));
	jand g22548(.dina(w_n22805_0[2]),.dinb(w_asqrt30_14[0]),.dout(n22806),.clk(gclk));
	jor g22549(.dina(w_n22805_0[1]),.dinb(w_asqrt30_13[2]),.dout(n22807),.clk(gclk));
	jxor g22550(.dina(w_n22067_0[0]),.dinb(w_n8003_20[1]),.dout(n22808),.clk(gclk));
	jand g22551(.dina(n22808),.dinb(w_asqrt4_22[2]),.dout(n22809),.clk(gclk));
	jxor g22552(.dina(n22809),.dinb(w_n22072_0[0]),.dout(n22810),.clk(gclk));
	jnot g22553(.din(w_n22810_0[1]),.dout(n22811),.clk(gclk));
	jand g22554(.dina(w_n22811_0[1]),.dinb(n22807),.dout(n22812),.clk(gclk));
	jor g22555(.dina(n22812),.dinb(w_n22806_0[1]),.dout(n22813),.clk(gclk));
	jand g22556(.dina(w_n22813_0[2]),.dinb(w_asqrt31_9[0]),.dout(n22814),.clk(gclk));
	jor g22557(.dina(w_n22813_0[1]),.dinb(w_asqrt31_8[2]),.dout(n22815),.clk(gclk));
	jxor g22558(.dina(w_n22074_0[0]),.dinb(w_n7581_15[2]),.dout(n22816),.clk(gclk));
	jand g22559(.dina(n22816),.dinb(w_asqrt4_22[1]),.dout(n22817),.clk(gclk));
	jxor g22560(.dina(n22817),.dinb(w_n22079_0[0]),.dout(n22818),.clk(gclk));
	jand g22561(.dina(w_n22818_0[1]),.dinb(n22815),.dout(n22819),.clk(gclk));
	jor g22562(.dina(n22819),.dinb(w_n22814_0[1]),.dout(n22820),.clk(gclk));
	jand g22563(.dina(w_n22820_0[2]),.dinb(w_asqrt32_14[0]),.dout(n22821),.clk(gclk));
	jor g22564(.dina(w_n22820_0[1]),.dinb(w_asqrt32_13[2]),.dout(n22822),.clk(gclk));
	jxor g22565(.dina(w_n22082_0[0]),.dinb(w_n7154_20[2]),.dout(n22823),.clk(gclk));
	jand g22566(.dina(n22823),.dinb(w_asqrt4_22[0]),.dout(n22824),.clk(gclk));
	jxor g22567(.dina(n22824),.dinb(w_n22087_0[0]),.dout(n22825),.clk(gclk));
	jnot g22568(.din(w_n22825_0[1]),.dout(n22826),.clk(gclk));
	jand g22569(.dina(w_n22826_0[1]),.dinb(n22822),.dout(n22827),.clk(gclk));
	jor g22570(.dina(n22827),.dinb(w_n22821_0[1]),.dout(n22828),.clk(gclk));
	jand g22571(.dina(w_n22828_0[2]),.dinb(w_asqrt33_9[2]),.dout(n22829),.clk(gclk));
	jor g22572(.dina(w_n22828_0[1]),.dinb(w_asqrt33_9[1]),.dout(n22830),.clk(gclk));
	jxor g22573(.dina(w_n22089_0[0]),.dinb(w_n6758_16[1]),.dout(n22831),.clk(gclk));
	jand g22574(.dina(n22831),.dinb(w_asqrt4_21[2]),.dout(n22832),.clk(gclk));
	jxor g22575(.dina(n22832),.dinb(w_n22094_0[0]),.dout(n22833),.clk(gclk));
	jand g22576(.dina(w_n22833_0[1]),.dinb(n22830),.dout(n22834),.clk(gclk));
	jor g22577(.dina(n22834),.dinb(w_n22829_0[1]),.dout(n22835),.clk(gclk));
	jand g22578(.dina(w_n22835_0[2]),.dinb(w_asqrt34_14[1]),.dout(n22836),.clk(gclk));
	jor g22579(.dina(w_n22835_0[1]),.dinb(w_asqrt34_14[0]),.dout(n22837),.clk(gclk));
	jxor g22580(.dina(w_n22097_0[0]),.dinb(w_n6357_21[0]),.dout(n22838),.clk(gclk));
	jand g22581(.dina(n22838),.dinb(w_asqrt4_21[1]),.dout(n22839),.clk(gclk));
	jxor g22582(.dina(n22839),.dinb(w_n22102_0[0]),.dout(n22840),.clk(gclk));
	jnot g22583(.din(w_n22840_0[1]),.dout(n22841),.clk(gclk));
	jand g22584(.dina(w_n22841_0[1]),.dinb(n22837),.dout(n22842),.clk(gclk));
	jor g22585(.dina(n22842),.dinb(w_n22836_0[1]),.dout(n22843),.clk(gclk));
	jand g22586(.dina(w_n22843_0[2]),.dinb(w_asqrt35_10[1]),.dout(n22844),.clk(gclk));
	jor g22587(.dina(w_n22843_0[1]),.dinb(w_asqrt35_10[0]),.dout(n22845),.clk(gclk));
	jxor g22588(.dina(w_n22104_0[0]),.dinb(w_n5989_17[0]),.dout(n22846),.clk(gclk));
	jand g22589(.dina(n22846),.dinb(w_asqrt4_21[0]),.dout(n22847),.clk(gclk));
	jxor g22590(.dina(n22847),.dinb(w_n22109_0[0]),.dout(n22848),.clk(gclk));
	jnot g22591(.din(w_n22848_0[1]),.dout(n22849),.clk(gclk));
	jand g22592(.dina(w_n22849_0[1]),.dinb(n22845),.dout(n22850),.clk(gclk));
	jor g22593(.dina(n22850),.dinb(w_n22844_0[1]),.dout(n22851),.clk(gclk));
	jand g22594(.dina(w_n22851_0[2]),.dinb(w_asqrt36_14[1]),.dout(n22852),.clk(gclk));
	jor g22595(.dina(w_n22851_0[1]),.dinb(w_asqrt36_14[0]),.dout(n22853),.clk(gclk));
	jxor g22596(.dina(w_n22111_0[0]),.dinb(w_n5606_21[1]),.dout(n22854),.clk(gclk));
	jand g22597(.dina(n22854),.dinb(w_asqrt4_20[2]),.dout(n22855),.clk(gclk));
	jxor g22598(.dina(n22855),.dinb(w_n22116_0[0]),.dout(n22856),.clk(gclk));
	jnot g22599(.din(w_n22856_0[1]),.dout(n22857),.clk(gclk));
	jand g22600(.dina(w_n22857_0[1]),.dinb(n22853),.dout(n22858),.clk(gclk));
	jor g22601(.dina(n22858),.dinb(w_n22852_0[1]),.dout(n22859),.clk(gclk));
	jand g22602(.dina(w_n22859_0[2]),.dinb(w_asqrt37_10[2]),.dout(n22860),.clk(gclk));
	jor g22603(.dina(w_n22859_0[1]),.dinb(w_asqrt37_10[1]),.dout(n22861),.clk(gclk));
	jxor g22604(.dina(w_n22118_0[0]),.dinb(w_n5259_18[0]),.dout(n22862),.clk(gclk));
	jand g22605(.dina(n22862),.dinb(w_asqrt4_20[1]),.dout(n22863),.clk(gclk));
	jxor g22606(.dina(n22863),.dinb(w_n22123_0[0]),.dout(n22864),.clk(gclk));
	jand g22607(.dina(w_n22864_0[1]),.dinb(n22861),.dout(n22865),.clk(gclk));
	jor g22608(.dina(n22865),.dinb(w_n22860_0[1]),.dout(n22866),.clk(gclk));
	jand g22609(.dina(w_n22866_0[2]),.dinb(w_asqrt38_14[2]),.dout(n22867),.clk(gclk));
	jor g22610(.dina(w_n22866_0[1]),.dinb(w_asqrt38_14[1]),.dout(n22868),.clk(gclk));
	jxor g22611(.dina(w_n22126_0[0]),.dinb(w_n4902_22[0]),.dout(n22869),.clk(gclk));
	jand g22612(.dina(n22869),.dinb(w_asqrt4_20[0]),.dout(n22870),.clk(gclk));
	jxor g22613(.dina(n22870),.dinb(w_n22131_0[0]),.dout(n22871),.clk(gclk));
	jnot g22614(.din(w_n22871_0[1]),.dout(n22872),.clk(gclk));
	jand g22615(.dina(w_n22872_0[1]),.dinb(n22868),.dout(n22873),.clk(gclk));
	jor g22616(.dina(n22873),.dinb(w_n22867_0[1]),.dout(n22874),.clk(gclk));
	jand g22617(.dina(w_n22874_0[2]),.dinb(w_asqrt39_11[1]),.dout(n22875),.clk(gclk));
	jor g22618(.dina(w_n22874_0[1]),.dinb(w_asqrt39_11[0]),.dout(n22876),.clk(gclk));
	jxor g22619(.dina(w_n22133_0[0]),.dinb(w_n4582_19[0]),.dout(n22877),.clk(gclk));
	jand g22620(.dina(n22877),.dinb(w_asqrt4_19[2]),.dout(n22878),.clk(gclk));
	jxor g22621(.dina(n22878),.dinb(w_n22138_0[0]),.dout(n22879),.clk(gclk));
	jand g22622(.dina(w_n22879_0[1]),.dinb(n22876),.dout(n22880),.clk(gclk));
	jor g22623(.dina(n22880),.dinb(w_n22875_0[1]),.dout(n22881),.clk(gclk));
	jand g22624(.dina(w_n22881_0[2]),.dinb(w_asqrt40_14[2]),.dout(n22882),.clk(gclk));
	jor g22625(.dina(w_n22881_0[1]),.dinb(w_asqrt40_14[1]),.dout(n22883),.clk(gclk));
	jxor g22626(.dina(w_n22141_0[0]),.dinb(w_n4249_22[2]),.dout(n22884),.clk(gclk));
	jand g22627(.dina(n22884),.dinb(w_asqrt4_19[1]),.dout(n22885),.clk(gclk));
	jxor g22628(.dina(n22885),.dinb(w_n22146_0[0]),.dout(n22886),.clk(gclk));
	jnot g22629(.din(w_n22886_0[1]),.dout(n22887),.clk(gclk));
	jand g22630(.dina(w_n22887_0[1]),.dinb(n22883),.dout(n22888),.clk(gclk));
	jor g22631(.dina(n22888),.dinb(w_n22882_0[1]),.dout(n22889),.clk(gclk));
	jand g22632(.dina(w_n22889_0[2]),.dinb(w_asqrt41_11[2]),.dout(n22890),.clk(gclk));
	jor g22633(.dina(w_n22889_0[1]),.dinb(w_asqrt41_11[1]),.dout(n22891),.clk(gclk));
	jxor g22634(.dina(w_n22148_0[0]),.dinb(w_n3955_19[2]),.dout(n22892),.clk(gclk));
	jand g22635(.dina(n22892),.dinb(w_asqrt4_19[0]),.dout(n22893),.clk(gclk));
	jxor g22636(.dina(n22893),.dinb(w_n22153_0[0]),.dout(n22894),.clk(gclk));
	jand g22637(.dina(w_n22894_0[1]),.dinb(n22891),.dout(n22895),.clk(gclk));
	jor g22638(.dina(n22895),.dinb(w_n22890_0[1]),.dout(n22896),.clk(gclk));
	jand g22639(.dina(w_n22896_0[2]),.dinb(w_asqrt42_15[0]),.dout(n22897),.clk(gclk));
	jor g22640(.dina(w_n22896_0[1]),.dinb(w_asqrt42_14[2]),.dout(n22898),.clk(gclk));
	jxor g22641(.dina(w_n22156_0[0]),.dinb(w_n3642_23[0]),.dout(n22899),.clk(gclk));
	jand g22642(.dina(n22899),.dinb(w_asqrt4_18[2]),.dout(n22900),.clk(gclk));
	jxor g22643(.dina(n22900),.dinb(w_n22161_0[0]),.dout(n22901),.clk(gclk));
	jnot g22644(.din(w_n22901_0[1]),.dout(n22902),.clk(gclk));
	jand g22645(.dina(w_n22902_0[1]),.dinb(n22898),.dout(n22903),.clk(gclk));
	jor g22646(.dina(n22903),.dinb(w_n22897_0[1]),.dout(n22904),.clk(gclk));
	jand g22647(.dina(w_n22904_0[2]),.dinb(w_asqrt43_12[0]),.dout(n22905),.clk(gclk));
	jor g22648(.dina(w_n22904_0[1]),.dinb(w_asqrt43_11[2]),.dout(n22906),.clk(gclk));
	jxor g22649(.dina(w_n22163_0[0]),.dinb(w_n3368_20[1]),.dout(n22907),.clk(gclk));
	jand g22650(.dina(n22907),.dinb(w_asqrt4_18[1]),.dout(n22908),.clk(gclk));
	jxor g22651(.dina(n22908),.dinb(w_n22168_0[0]),.dout(n22909),.clk(gclk));
	jand g22652(.dina(w_n22909_0[1]),.dinb(n22906),.dout(n22910),.clk(gclk));
	jor g22653(.dina(n22910),.dinb(w_n22905_0[1]),.dout(n22911),.clk(gclk));
	jand g22654(.dina(w_n22911_0[2]),.dinb(w_asqrt44_15[0]),.dout(n22912),.clk(gclk));
	jor g22655(.dina(w_n22911_0[1]),.dinb(w_asqrt44_14[2]),.dout(n22913),.clk(gclk));
	jxor g22656(.dina(w_n22171_0[0]),.dinb(w_n3089_23[2]),.dout(n22914),.clk(gclk));
	jand g22657(.dina(n22914),.dinb(w_asqrt4_18[0]),.dout(n22915),.clk(gclk));
	jxor g22658(.dina(n22915),.dinb(w_n22176_0[0]),.dout(n22916),.clk(gclk));
	jnot g22659(.din(w_n22916_0[1]),.dout(n22917),.clk(gclk));
	jand g22660(.dina(w_n22917_0[1]),.dinb(n22913),.dout(n22918),.clk(gclk));
	jor g22661(.dina(n22918),.dinb(w_n22912_0[1]),.dout(n22919),.clk(gclk));
	jand g22662(.dina(w_n22919_0[2]),.dinb(w_asqrt45_12[2]),.dout(n22920),.clk(gclk));
	jor g22663(.dina(w_n22919_0[1]),.dinb(w_asqrt45_12[1]),.dout(n22921),.clk(gclk));
	jxor g22664(.dina(w_n22178_0[0]),.dinb(w_n2833_21[1]),.dout(n22922),.clk(gclk));
	jand g22665(.dina(n22922),.dinb(w_asqrt4_17[2]),.dout(n22923),.clk(gclk));
	jxor g22666(.dina(n22923),.dinb(w_n22183_0[0]),.dout(n22924),.clk(gclk));
	jnot g22667(.din(w_n22924_0[1]),.dout(n22925),.clk(gclk));
	jand g22668(.dina(w_n22925_0[1]),.dinb(n22921),.dout(n22926),.clk(gclk));
	jor g22669(.dina(n22926),.dinb(w_n22920_0[1]),.dout(n22927),.clk(gclk));
	jand g22670(.dina(w_n22927_0[2]),.dinb(w_asqrt46_15[0]),.dout(n22928),.clk(gclk));
	jor g22671(.dina(w_n22927_0[1]),.dinb(w_asqrt46_14[2]),.dout(n22929),.clk(gclk));
	jxor g22672(.dina(w_n22185_0[0]),.dinb(w_n2572_24[0]),.dout(n22930),.clk(gclk));
	jand g22673(.dina(n22930),.dinb(w_asqrt4_17[1]),.dout(n22931),.clk(gclk));
	jxor g22674(.dina(n22931),.dinb(w_n22190_0[0]),.dout(n22932),.clk(gclk));
	jnot g22675(.din(w_n22932_0[1]),.dout(n22933),.clk(gclk));
	jand g22676(.dina(w_n22933_0[1]),.dinb(n22929),.dout(n22934),.clk(gclk));
	jor g22677(.dina(n22934),.dinb(w_n22928_0[1]),.dout(n22935),.clk(gclk));
	jand g22678(.dina(w_n22935_0[2]),.dinb(w_asqrt47_13[1]),.dout(n22936),.clk(gclk));
	jor g22679(.dina(w_n22935_0[1]),.dinb(w_asqrt47_13[0]),.dout(n22937),.clk(gclk));
	jxor g22680(.dina(w_n22192_0[0]),.dinb(w_n2345_22[0]),.dout(n22938),.clk(gclk));
	jand g22681(.dina(n22938),.dinb(w_asqrt4_17[0]),.dout(n22939),.clk(gclk));
	jxor g22682(.dina(n22939),.dinb(w_n22197_0[0]),.dout(n22940),.clk(gclk));
	jand g22683(.dina(w_n22940_0[1]),.dinb(n22937),.dout(n22941),.clk(gclk));
	jor g22684(.dina(n22941),.dinb(w_n22936_0[1]),.dout(n22942),.clk(gclk));
	jand g22685(.dina(w_n22942_0[2]),.dinb(w_asqrt48_15[1]),.dout(n22943),.clk(gclk));
	jor g22686(.dina(w_n22942_0[1]),.dinb(w_asqrt48_15[0]),.dout(n22944),.clk(gclk));
	jxor g22687(.dina(w_n22200_0[0]),.dinb(w_n2108_24[2]),.dout(n22945),.clk(gclk));
	jand g22688(.dina(n22945),.dinb(w_asqrt4_16[2]),.dout(n22946),.clk(gclk));
	jxor g22689(.dina(n22946),.dinb(w_n22205_0[0]),.dout(n22947),.clk(gclk));
	jnot g22690(.din(w_n22947_0[1]),.dout(n22948),.clk(gclk));
	jand g22691(.dina(w_n22948_0[1]),.dinb(n22944),.dout(n22949),.clk(gclk));
	jor g22692(.dina(n22949),.dinb(w_n22943_0[1]),.dout(n22950),.clk(gclk));
	jand g22693(.dina(w_n22950_0[2]),.dinb(w_asqrt49_13[2]),.dout(n22951),.clk(gclk));
	jor g22694(.dina(w_n22950_0[1]),.dinb(w_asqrt49_13[1]),.dout(n22952),.clk(gclk));
	jxor g22695(.dina(w_n22207_0[0]),.dinb(w_n1912_23[0]),.dout(n22953),.clk(gclk));
	jand g22696(.dina(n22953),.dinb(w_asqrt4_16[1]),.dout(n22954),.clk(gclk));
	jxor g22697(.dina(n22954),.dinb(w_n22212_0[0]),.dout(n22955),.clk(gclk));
	jnot g22698(.din(w_n22955_0[1]),.dout(n22956),.clk(gclk));
	jand g22699(.dina(w_n22956_0[1]),.dinb(n22952),.dout(n22957),.clk(gclk));
	jor g22700(.dina(n22957),.dinb(w_n22951_0[1]),.dout(n22958),.clk(gclk));
	jand g22701(.dina(w_n22958_0[2]),.dinb(w_asqrt50_15[2]),.dout(n22959),.clk(gclk));
	jor g22702(.dina(w_n22958_0[1]),.dinb(w_asqrt50_15[1]),.dout(n22960),.clk(gclk));
	jxor g22703(.dina(w_n22214_0[0]),.dinb(w_n1699_25[1]),.dout(n22961),.clk(gclk));
	jand g22704(.dina(n22961),.dinb(w_asqrt4_16[0]),.dout(n22962),.clk(gclk));
	jxor g22705(.dina(n22962),.dinb(w_n22219_0[0]),.dout(n22963),.clk(gclk));
	jnot g22706(.din(w_n22963_0[1]),.dout(n22964),.clk(gclk));
	jand g22707(.dina(w_n22964_0[1]),.dinb(n22960),.dout(n22965),.clk(gclk));
	jor g22708(.dina(n22965),.dinb(w_n22959_0[1]),.dout(n22966),.clk(gclk));
	jand g22709(.dina(w_n22966_0[2]),.dinb(w_asqrt51_14[0]),.dout(n22967),.clk(gclk));
	jor g22710(.dina(w_n22966_0[1]),.dinb(w_asqrt51_13[2]),.dout(n22968),.clk(gclk));
	jxor g22711(.dina(w_n22221_0[0]),.dinb(w_n1516_23[2]),.dout(n22969),.clk(gclk));
	jand g22712(.dina(n22969),.dinb(w_asqrt4_15[2]),.dout(n22970),.clk(gclk));
	jxor g22713(.dina(n22970),.dinb(w_n22226_0[0]),.dout(n22971),.clk(gclk));
	jnot g22714(.din(w_n22971_0[1]),.dout(n22972),.clk(gclk));
	jand g22715(.dina(w_n22972_0[1]),.dinb(n22968),.dout(n22973),.clk(gclk));
	jor g22716(.dina(n22973),.dinb(w_n22967_0[1]),.dout(n22974),.clk(gclk));
	jand g22717(.dina(w_n22974_0[2]),.dinb(w_asqrt52_15[2]),.dout(n22975),.clk(gclk));
	jor g22718(.dina(w_n22974_0[1]),.dinb(w_asqrt52_15[1]),.dout(n22976),.clk(gclk));
	jxor g22719(.dina(w_n22228_0[0]),.dinb(w_n1332_25[1]),.dout(n22977),.clk(gclk));
	jand g22720(.dina(n22977),.dinb(w_asqrt4_15[1]),.dout(n22978),.clk(gclk));
	jxor g22721(.dina(n22978),.dinb(w_n22233_0[0]),.dout(n22979),.clk(gclk));
	jnot g22722(.din(w_n22979_0[1]),.dout(n22980),.clk(gclk));
	jand g22723(.dina(w_n22980_0[1]),.dinb(n22976),.dout(n22981),.clk(gclk));
	jor g22724(.dina(n22981),.dinb(w_n22975_0[1]),.dout(n22982),.clk(gclk));
	jand g22725(.dina(w_n22982_0[2]),.dinb(w_asqrt53_14[2]),.dout(n22983),.clk(gclk));
	jor g22726(.dina(w_n22982_0[1]),.dinb(w_asqrt53_14[1]),.dout(n22984),.clk(gclk));
	jxor g22727(.dina(w_n22235_0[0]),.dinb(w_n1173_24[1]),.dout(n22985),.clk(gclk));
	jand g22728(.dina(n22985),.dinb(w_asqrt4_15[0]),.dout(n22986),.clk(gclk));
	jxor g22729(.dina(n22986),.dinb(w_n22240_0[0]),.dout(n22987),.clk(gclk));
	jand g22730(.dina(w_n22987_0[1]),.dinb(n22984),.dout(n22988),.clk(gclk));
	jor g22731(.dina(n22988),.dinb(w_n22983_0[1]),.dout(n22989),.clk(gclk));
	jand g22732(.dina(w_n22989_0[2]),.dinb(w_asqrt54_15[2]),.dout(n22990),.clk(gclk));
	jor g22733(.dina(w_n22989_0[1]),.dinb(w_asqrt54_15[1]),.dout(n22991),.clk(gclk));
	jxor g22734(.dina(w_n22243_0[0]),.dinb(w_n1008_26[1]),.dout(n22992),.clk(gclk));
	jand g22735(.dina(n22992),.dinb(w_asqrt4_14[2]),.dout(n22993),.clk(gclk));
	jxor g22736(.dina(n22993),.dinb(w_n22248_0[0]),.dout(n22994),.clk(gclk));
	jnot g22737(.din(w_n22994_0[1]),.dout(n22995),.clk(gclk));
	jand g22738(.dina(w_n22995_0[1]),.dinb(n22991),.dout(n22996),.clk(gclk));
	jor g22739(.dina(n22996),.dinb(w_n22990_0[1]),.dout(n22997),.clk(gclk));
	jand g22740(.dina(w_n22997_0[2]),.dinb(w_asqrt55_15[0]),.dout(n22998),.clk(gclk));
	jor g22741(.dina(w_n22997_0[1]),.dinb(w_asqrt55_14[2]),.dout(n22999),.clk(gclk));
	jxor g22742(.dina(w_n22250_0[0]),.dinb(w_n884_25[1]),.dout(n23000),.clk(gclk));
	jand g22743(.dina(n23000),.dinb(w_asqrt4_14[1]),.dout(n23001),.clk(gclk));
	jxor g22744(.dina(n23001),.dinb(w_n22255_0[0]),.dout(n23002),.clk(gclk));
	jand g22745(.dina(w_n23002_0[1]),.dinb(n22999),.dout(n23003),.clk(gclk));
	jor g22746(.dina(n23003),.dinb(w_n22998_0[1]),.dout(n23004),.clk(gclk));
	jand g22747(.dina(w_n23004_0[2]),.dinb(w_asqrt56_16[0]),.dout(n23005),.clk(gclk));
	jor g22748(.dina(w_n23004_0[1]),.dinb(w_asqrt56_15[2]),.dout(n23006),.clk(gclk));
	jxor g22749(.dina(w_n22258_0[0]),.dinb(w_n743_26[1]),.dout(n23007),.clk(gclk));
	jand g22750(.dina(n23007),.dinb(w_asqrt4_14[0]),.dout(n23008),.clk(gclk));
	jxor g22751(.dina(n23008),.dinb(w_n22263_0[0]),.dout(n23009),.clk(gclk));
	jnot g22752(.din(w_n23009_0[1]),.dout(n23010),.clk(gclk));
	jand g22753(.dina(w_n23010_0[1]),.dinb(n23006),.dout(n23011),.clk(gclk));
	jor g22754(.dina(n23011),.dinb(w_n23005_0[1]),.dout(n23012),.clk(gclk));
	jand g22755(.dina(w_n23012_0[2]),.dinb(w_asqrt57_15[2]),.dout(n23013),.clk(gclk));
	jor g22756(.dina(w_n23012_0[1]),.dinb(w_asqrt57_15[1]),.dout(n23014),.clk(gclk));
	jxor g22757(.dina(w_n22265_0[0]),.dinb(w_n635_26[1]),.dout(n23015),.clk(gclk));
	jand g22758(.dina(n23015),.dinb(w_asqrt4_13[2]),.dout(n23016),.clk(gclk));
	jxor g22759(.dina(n23016),.dinb(w_n22270_0[0]),.dout(n23017),.clk(gclk));
	jnot g22760(.din(w_n23017_0[1]),.dout(n23018),.clk(gclk));
	jand g22761(.dina(w_n23018_0[1]),.dinb(n23014),.dout(n23019),.clk(gclk));
	jor g22762(.dina(n23019),.dinb(w_n23013_0[1]),.dout(n23020),.clk(gclk));
	jand g22763(.dina(w_n23020_0[2]),.dinb(w_asqrt58_16[1]),.dout(n23021),.clk(gclk));
	jor g22764(.dina(w_n23020_0[1]),.dinb(w_asqrt58_16[0]),.dout(n23022),.clk(gclk));
	jxor g22765(.dina(w_n22272_0[0]),.dinb(w_n515_27[1]),.dout(n23023),.clk(gclk));
	jand g22766(.dina(n23023),.dinb(w_asqrt4_13[1]),.dout(n23024),.clk(gclk));
	jxor g22767(.dina(n23024),.dinb(w_n22277_0[0]),.dout(n23025),.clk(gclk));
	jand g22768(.dina(w_n23025_0[1]),.dinb(n23022),.dout(n23026),.clk(gclk));
	jor g22769(.dina(n23026),.dinb(w_n23021_0[1]),.dout(n23027),.clk(gclk));
	jand g22770(.dina(w_n23027_0[2]),.dinb(w_asqrt59_16[0]),.dout(n23028),.clk(gclk));
	jor g22771(.dina(w_n23027_0[1]),.dinb(w_asqrt59_15[2]),.dout(n23029),.clk(gclk));
	jxor g22772(.dina(w_n22280_0[0]),.dinb(w_n443_27[1]),.dout(n23030),.clk(gclk));
	jand g22773(.dina(n23030),.dinb(w_asqrt4_13[0]),.dout(n23031),.clk(gclk));
	jxor g22774(.dina(n23031),.dinb(w_n22285_0[0]),.dout(n23032),.clk(gclk));
	jand g22775(.dina(w_n23032_0[1]),.dinb(n23029),.dout(n23033),.clk(gclk));
	jor g22776(.dina(n23033),.dinb(w_n23028_0[1]),.dout(n23034),.clk(gclk));
	jand g22777(.dina(w_n23034_0[2]),.dinb(w_asqrt60_16[1]),.dout(n23035),.clk(gclk));
	jor g22778(.dina(w_n23034_0[1]),.dinb(w_asqrt60_16[0]),.dout(n23036),.clk(gclk));
	jxor g22779(.dina(w_n22288_0[0]),.dinb(w_n352_27[2]),.dout(n23037),.clk(gclk));
	jand g22780(.dina(n23037),.dinb(w_asqrt4_12[2]),.dout(n23038),.clk(gclk));
	jxor g22781(.dina(n23038),.dinb(w_n22293_0[0]),.dout(n23039),.clk(gclk));
	jnot g22782(.din(w_n23039_0[1]),.dout(n23040),.clk(gclk));
	jand g22783(.dina(w_n23040_0[1]),.dinb(n23036),.dout(n23041),.clk(gclk));
	jor g22784(.dina(n23041),.dinb(w_n23035_0[1]),.dout(n23042),.clk(gclk));
	jand g22785(.dina(w_n23042_0[2]),.dinb(w_asqrt61_16[1]),.dout(n23043),.clk(gclk));
	jor g22786(.dina(w_n23042_0[1]),.dinb(w_asqrt61_16[0]),.dout(n23044),.clk(gclk));
	jxor g22787(.dina(w_n22295_0[0]),.dinb(w_n294_28[0]),.dout(n23045),.clk(gclk));
	jand g22788(.dina(n23045),.dinb(w_asqrt4_12[1]),.dout(n23046),.clk(gclk));
	jxor g22789(.dina(n23046),.dinb(w_n22300_0[0]),.dout(n23047),.clk(gclk));
	jnot g22790(.din(w_n23047_0[1]),.dout(n23048),.clk(gclk));
	jand g22791(.dina(w_n23048_0[1]),.dinb(n23044),.dout(n23049),.clk(gclk));
	jor g22792(.dina(n23049),.dinb(w_n23043_0[1]),.dout(n23050),.clk(gclk));
	jand g22793(.dina(w_n23050_0[2]),.dinb(w_asqrt62_16[1]),.dout(n23051),.clk(gclk));
	jor g22794(.dina(w_n23050_0[1]),.dinb(w_asqrt62_16[0]),.dout(n23052),.clk(gclk));
	jxor g22795(.dina(w_n22302_0[0]),.dinb(w_n239_28[0]),.dout(n23053),.clk(gclk));
	jand g22796(.dina(n23053),.dinb(w_asqrt4_12[0]),.dout(n23054),.clk(gclk));
	jxor g22797(.dina(n23054),.dinb(w_n22307_0[0]),.dout(n23055),.clk(gclk));
	jnot g22798(.din(w_n23055_0[2]),.dout(n23056),.clk(gclk));
	jand g22799(.dina(n23056),.dinb(n23052),.dout(n23057),.clk(gclk));
	jor g22800(.dina(n23057),.dinb(w_n23051_0[1]),.dout(n23058),.clk(gclk));
	jxor g22801(.dina(w_n22309_0[0]),.dinb(w_n221_28[1]),.dout(n23059),.clk(gclk));
	jand g22802(.dina(n23059),.dinb(w_asqrt4_11[2]),.dout(n23060),.clk(gclk));
	jxor g22803(.dina(n23060),.dinb(w_n22315_0[0]),.dout(n23061),.clk(gclk));
	jnot g22804(.din(w_n23061_0[1]),.dout(n23062),.clk(gclk));
	jor g22805(.dina(w_n23062_0[1]),.dinb(w_n23058_0[1]),.dout(n23063),.clk(gclk));
	jnot g22806(.din(w_n23063_1[1]),.dout(n23064),.clk(gclk));
	jand g22807(.dina(w_n22332_0[0]),.dinb(w_n22615_0[0]),.dout(n23065),.clk(gclk));
	jnot g22808(.din(w_n23051_0[0]),.dout(n23066),.clk(gclk));
	jnot g22809(.din(w_n23043_0[0]),.dout(n23067),.clk(gclk));
	jnot g22810(.din(w_n23035_0[0]),.dout(n23068),.clk(gclk));
	jnot g22811(.din(w_n23028_0[0]),.dout(n23069),.clk(gclk));
	jnot g22812(.din(w_n23021_0[0]),.dout(n23070),.clk(gclk));
	jnot g22813(.din(w_n23013_0[0]),.dout(n23071),.clk(gclk));
	jnot g22814(.din(w_n23005_0[0]),.dout(n23072),.clk(gclk));
	jnot g22815(.din(w_n22998_0[0]),.dout(n23073),.clk(gclk));
	jnot g22816(.din(w_n22990_0[0]),.dout(n23074),.clk(gclk));
	jnot g22817(.din(w_n22983_0[0]),.dout(n23075),.clk(gclk));
	jnot g22818(.din(w_n22975_0[0]),.dout(n23076),.clk(gclk));
	jnot g22819(.din(w_n22967_0[0]),.dout(n23077),.clk(gclk));
	jnot g22820(.din(w_n22959_0[0]),.dout(n23078),.clk(gclk));
	jnot g22821(.din(w_n22951_0[0]),.dout(n23079),.clk(gclk));
	jnot g22822(.din(w_n22943_0[0]),.dout(n23080),.clk(gclk));
	jnot g22823(.din(w_n22936_0[0]),.dout(n23081),.clk(gclk));
	jnot g22824(.din(w_n22928_0[0]),.dout(n23082),.clk(gclk));
	jnot g22825(.din(w_n22920_0[0]),.dout(n23083),.clk(gclk));
	jnot g22826(.din(w_n22912_0[0]),.dout(n23084),.clk(gclk));
	jnot g22827(.din(w_n22905_0[0]),.dout(n23085),.clk(gclk));
	jnot g22828(.din(w_n22897_0[0]),.dout(n23086),.clk(gclk));
	jnot g22829(.din(w_n22890_0[0]),.dout(n23087),.clk(gclk));
	jnot g22830(.din(w_n22882_0[0]),.dout(n23088),.clk(gclk));
	jnot g22831(.din(w_n22875_0[0]),.dout(n23089),.clk(gclk));
	jnot g22832(.din(w_n22867_0[0]),.dout(n23090),.clk(gclk));
	jnot g22833(.din(w_n22860_0[0]),.dout(n23091),.clk(gclk));
	jnot g22834(.din(w_n22852_0[0]),.dout(n23092),.clk(gclk));
	jnot g22835(.din(w_n22844_0[0]),.dout(n23093),.clk(gclk));
	jnot g22836(.din(w_n22836_0[0]),.dout(n23094),.clk(gclk));
	jnot g22837(.din(w_n22829_0[0]),.dout(n23095),.clk(gclk));
	jnot g22838(.din(w_n22821_0[0]),.dout(n23096),.clk(gclk));
	jnot g22839(.din(w_n22814_0[0]),.dout(n23097),.clk(gclk));
	jnot g22840(.din(w_n22806_0[0]),.dout(n23098),.clk(gclk));
	jnot g22841(.din(w_n22799_0[0]),.dout(n23099),.clk(gclk));
	jnot g22842(.din(w_n22792_0[0]),.dout(n23100),.clk(gclk));
	jnot g22843(.din(w_n22784_0[0]),.dout(n23101),.clk(gclk));
	jnot g22844(.din(w_n22776_0[0]),.dout(n23102),.clk(gclk));
	jnot g22845(.din(w_n22769_0[0]),.dout(n23103),.clk(gclk));
	jnot g22846(.din(w_n22761_0[0]),.dout(n23104),.clk(gclk));
	jnot g22847(.din(w_n22754_0[0]),.dout(n23105),.clk(gclk));
	jnot g22848(.din(w_n22746_0[0]),.dout(n23106),.clk(gclk));
	jnot g22849(.din(w_n22739_0[0]),.dout(n23107),.clk(gclk));
	jnot g22850(.din(w_n22731_0[0]),.dout(n23108),.clk(gclk));
	jnot g22851(.din(w_n22723_0[0]),.dout(n23109),.clk(gclk));
	jnot g22852(.din(w_n22715_0[0]),.dout(n23110),.clk(gclk));
	jnot g22853(.din(w_n22708_0[0]),.dout(n23111),.clk(gclk));
	jnot g22854(.din(w_n22700_0[0]),.dout(n23112),.clk(gclk));
	jnot g22855(.din(w_n22692_0[0]),.dout(n23113),.clk(gclk));
	jnot g22856(.din(w_n22684_0[0]),.dout(n23114),.clk(gclk));
	jnot g22857(.din(w_n22677_0[0]),.dout(n23115),.clk(gclk));
	jnot g22858(.din(w_n22669_0[0]),.dout(n23116),.clk(gclk));
	jnot g22859(.din(w_n22662_0[0]),.dout(n23117),.clk(gclk));
	jnot g22860(.din(w_n22654_0[0]),.dout(n23118),.clk(gclk));
	jnot g22861(.din(w_n22647_0[0]),.dout(n23119),.clk(gclk));
	jnot g22862(.din(w_n22640_0[0]),.dout(n23120),.clk(gclk));
	jnot g22863(.din(w_n22633_0[0]),.dout(n23121),.clk(gclk));
	jnot g22864(.din(w_n22625_0[0]),.dout(n23122),.clk(gclk));
	jnot g22865(.din(w_n22340_0[0]),.dout(n23123),.clk(gclk));
	jnot g22866(.din(w_n22337_0[0]),.dout(n23124),.clk(gclk));
	jor g22867(.dina(w_n22620_4[1]),.dinb(w_n21889_0[2]),.dout(n23125),.clk(gclk));
	jand g22868(.dina(n23125),.dinb(n23124),.dout(n23126),.clk(gclk));
	jand g22869(.dina(n23126),.dinb(w_n21887_14[0]),.dout(n23127),.clk(gclk));
	jor g22870(.dina(w_n22620_4[0]),.dinb(w_a8_0[0]),.dout(n23128),.clk(gclk));
	jand g22871(.dina(n23128),.dinb(w_a9_0[0]),.dout(n23129),.clk(gclk));
	jand g22872(.dina(w_asqrt4_11[1]),.dinb(w_n21891_0[0]),.dout(n23130),.clk(gclk));
	jor g22873(.dina(n23130),.dinb(n23129),.dout(n23131),.clk(gclk));
	jor g22874(.dina(n23131),.dinb(n23127),.dout(n23132),.clk(gclk));
	jand g22875(.dina(n23132),.dinb(n23123),.dout(n23133),.clk(gclk));
	jand g22876(.dina(n23133),.dinb(w_n21184_5[0]),.dout(n23134),.clk(gclk));
	jor g22877(.dina(w_n22629_0[0]),.dinb(n23134),.dout(n23135),.clk(gclk));
	jand g22878(.dina(n23135),.dinb(n23122),.dout(n23136),.clk(gclk));
	jand g22879(.dina(n23136),.dinb(w_n20468_14[1]),.dout(n23137),.clk(gclk));
	jnot g22880(.din(w_n22637_0[0]),.dout(n23138),.clk(gclk));
	jor g22881(.dina(w_n23138_0[1]),.dinb(n23137),.dout(n23139),.clk(gclk));
	jand g22882(.dina(n23139),.dinb(n23121),.dout(n23140),.clk(gclk));
	jand g22883(.dina(n23140),.dinb(w_n19791_6[0]),.dout(n23141),.clk(gclk));
	jnot g22884(.din(w_n22644_0[0]),.dout(n23142),.clk(gclk));
	jor g22885(.dina(w_n23142_0[1]),.dinb(n23141),.dout(n23143),.clk(gclk));
	jand g22886(.dina(n23143),.dinb(n23120),.dout(n23144),.clk(gclk));
	jand g22887(.dina(n23144),.dinb(w_n19096_14[2]),.dout(n23145),.clk(gclk));
	jnot g22888(.din(w_n22651_0[0]),.dout(n23146),.clk(gclk));
	jor g22889(.dina(w_n23146_0[1]),.dinb(n23145),.dout(n23147),.clk(gclk));
	jand g22890(.dina(n23147),.dinb(n23119),.dout(n23148),.clk(gclk));
	jand g22891(.dina(n23148),.dinb(w_n18442_6[2]),.dout(n23149),.clk(gclk));
	jor g22892(.dina(w_n22658_0[0]),.dinb(n23149),.dout(n23150),.clk(gclk));
	jand g22893(.dina(n23150),.dinb(n23118),.dout(n23151),.clk(gclk));
	jand g22894(.dina(n23151),.dinb(w_n17769_15[1]),.dout(n23152),.clk(gclk));
	jnot g22895(.din(w_n22666_0[0]),.dout(n23153),.clk(gclk));
	jor g22896(.dina(w_n23153_0[1]),.dinb(n23152),.dout(n23154),.clk(gclk));
	jand g22897(.dina(n23154),.dinb(n23117),.dout(n23155),.clk(gclk));
	jand g22898(.dina(n23155),.dinb(w_n17134_7[2]),.dout(n23156),.clk(gclk));
	jor g22899(.dina(w_n22673_0[0]),.dinb(n23156),.dout(n23157),.clk(gclk));
	jand g22900(.dina(n23157),.dinb(n23116),.dout(n23158),.clk(gclk));
	jand g22901(.dina(n23158),.dinb(w_n16489_15[2]),.dout(n23159),.clk(gclk));
	jnot g22902(.din(w_n22681_0[0]),.dout(n23160),.clk(gclk));
	jor g22903(.dina(w_n23160_0[1]),.dinb(n23159),.dout(n23161),.clk(gclk));
	jand g22904(.dina(n23161),.dinb(n23115),.dout(n23162),.clk(gclk));
	jand g22905(.dina(n23162),.dinb(w_n15878_8[2]),.dout(n23163),.clk(gclk));
	jor g22906(.dina(w_n22688_0[0]),.dinb(n23163),.dout(n23164),.clk(gclk));
	jand g22907(.dina(n23164),.dinb(n23114),.dout(n23165),.clk(gclk));
	jand g22908(.dina(n23165),.dinb(w_n15260_16[1]),.dout(n23166),.clk(gclk));
	jor g22909(.dina(w_n22696_0[0]),.dinb(n23166),.dout(n23167),.clk(gclk));
	jand g22910(.dina(n23167),.dinb(n23113),.dout(n23168),.clk(gclk));
	jand g22911(.dina(n23168),.dinb(w_n14674_9[1]),.dout(n23169),.clk(gclk));
	jor g22912(.dina(w_n22704_0[0]),.dinb(n23169),.dout(n23170),.clk(gclk));
	jand g22913(.dina(n23170),.dinb(n23112),.dout(n23171),.clk(gclk));
	jand g22914(.dina(n23171),.dinb(w_n14078_16[2]),.dout(n23172),.clk(gclk));
	jnot g22915(.din(w_n22712_0[0]),.dout(n23173),.clk(gclk));
	jor g22916(.dina(w_n23173_0[1]),.dinb(n23172),.dout(n23174),.clk(gclk));
	jand g22917(.dina(n23174),.dinb(n23111),.dout(n23175),.clk(gclk));
	jand g22918(.dina(n23175),.dinb(w_n13515_10[1]),.dout(n23176),.clk(gclk));
	jor g22919(.dina(w_n22719_0[0]),.dinb(n23176),.dout(n23177),.clk(gclk));
	jand g22920(.dina(n23177),.dinb(n23110),.dout(n23178),.clk(gclk));
	jand g22921(.dina(n23178),.dinb(w_n12947_17[1]),.dout(n23179),.clk(gclk));
	jor g22922(.dina(w_n22727_0[0]),.dinb(n23179),.dout(n23180),.clk(gclk));
	jand g22923(.dina(n23180),.dinb(n23109),.dout(n23181),.clk(gclk));
	jand g22924(.dina(n23181),.dinb(w_n12410_11[0]),.dout(n23182),.clk(gclk));
	jor g22925(.dina(w_n22735_0[0]),.dinb(n23182),.dout(n23183),.clk(gclk));
	jand g22926(.dina(n23183),.dinb(n23108),.dout(n23184),.clk(gclk));
	jand g22927(.dina(n23184),.dinb(w_n11858_17[2]),.dout(n23185),.clk(gclk));
	jnot g22928(.din(w_n22743_0[0]),.dout(n23186),.clk(gclk));
	jor g22929(.dina(w_n23186_0[1]),.dinb(n23185),.dout(n23187),.clk(gclk));
	jand g22930(.dina(n23187),.dinb(n23107),.dout(n23188),.clk(gclk));
	jand g22931(.dina(n23188),.dinb(w_n11347_11[2]),.dout(n23189),.clk(gclk));
	jor g22932(.dina(w_n22750_0[0]),.dinb(n23189),.dout(n23190),.clk(gclk));
	jand g22933(.dina(n23190),.dinb(n23106),.dout(n23191),.clk(gclk));
	jand g22934(.dina(n23191),.dinb(w_n10824_18[1]),.dout(n23192),.clk(gclk));
	jnot g22935(.din(w_n22758_0[0]),.dout(n23193),.clk(gclk));
	jor g22936(.dina(w_n23193_0[1]),.dinb(n23192),.dout(n23194),.clk(gclk));
	jand g22937(.dina(n23194),.dinb(n23105),.dout(n23195),.clk(gclk));
	jand g22938(.dina(n23195),.dinb(w_n10328_12[2]),.dout(n23196),.clk(gclk));
	jor g22939(.dina(w_n22765_0[0]),.dinb(n23196),.dout(n23197),.clk(gclk));
	jand g22940(.dina(n23197),.dinb(n23104),.dout(n23198),.clk(gclk));
	jand g22941(.dina(n23198),.dinb(w_n9832_19[0]),.dout(n23199),.clk(gclk));
	jnot g22942(.din(w_n22773_0[0]),.dout(n23200),.clk(gclk));
	jor g22943(.dina(w_n23200_0[1]),.dinb(n23199),.dout(n23201),.clk(gclk));
	jand g22944(.dina(n23201),.dinb(n23103),.dout(n23202),.clk(gclk));
	jand g22945(.dina(n23202),.dinb(w_n9369_13[2]),.dout(n23203),.clk(gclk));
	jor g22946(.dina(w_n22780_0[0]),.dinb(n23203),.dout(n23204),.clk(gclk));
	jand g22947(.dina(n23204),.dinb(n23102),.dout(n23205),.clk(gclk));
	jand g22948(.dina(n23205),.dinb(w_n8890_19[1]),.dout(n23206),.clk(gclk));
	jor g22949(.dina(w_n22788_0[0]),.dinb(n23206),.dout(n23207),.clk(gclk));
	jand g22950(.dina(n23207),.dinb(n23101),.dout(n23208),.clk(gclk));
	jand g22951(.dina(n23208),.dinb(w_n8449_14[1]),.dout(n23209),.clk(gclk));
	jnot g22952(.din(w_n22796_0[0]),.dout(n23210),.clk(gclk));
	jor g22953(.dina(w_n23210_0[1]),.dinb(n23209),.dout(n23211),.clk(gclk));
	jand g22954(.dina(n23211),.dinb(n23100),.dout(n23212),.clk(gclk));
	jand g22955(.dina(n23212),.dinb(w_n8003_20[0]),.dout(n23213),.clk(gclk));
	jnot g22956(.din(w_n22803_0[0]),.dout(n23214),.clk(gclk));
	jor g22957(.dina(w_n23214_0[1]),.dinb(n23213),.dout(n23215),.clk(gclk));
	jand g22958(.dina(n23215),.dinb(n23099),.dout(n23216),.clk(gclk));
	jand g22959(.dina(n23216),.dinb(w_n7581_15[1]),.dout(n23217),.clk(gclk));
	jor g22960(.dina(w_n22810_0[0]),.dinb(n23217),.dout(n23218),.clk(gclk));
	jand g22961(.dina(n23218),.dinb(n23098),.dout(n23219),.clk(gclk));
	jand g22962(.dina(n23219),.dinb(w_n7154_20[1]),.dout(n23220),.clk(gclk));
	jnot g22963(.din(w_n22818_0[0]),.dout(n23221),.clk(gclk));
	jor g22964(.dina(w_n23221_0[1]),.dinb(n23220),.dout(n23222),.clk(gclk));
	jand g22965(.dina(n23222),.dinb(n23097),.dout(n23223),.clk(gclk));
	jand g22966(.dina(n23223),.dinb(w_n6758_16[0]),.dout(n23224),.clk(gclk));
	jor g22967(.dina(w_n22825_0[0]),.dinb(n23224),.dout(n23225),.clk(gclk));
	jand g22968(.dina(n23225),.dinb(n23096),.dout(n23226),.clk(gclk));
	jand g22969(.dina(n23226),.dinb(w_n6357_20[2]),.dout(n23227),.clk(gclk));
	jnot g22970(.din(w_n22833_0[0]),.dout(n23228),.clk(gclk));
	jor g22971(.dina(w_n23228_0[1]),.dinb(n23227),.dout(n23229),.clk(gclk));
	jand g22972(.dina(n23229),.dinb(n23095),.dout(n23230),.clk(gclk));
	jand g22973(.dina(n23230),.dinb(w_n5989_16[2]),.dout(n23231),.clk(gclk));
	jor g22974(.dina(w_n22840_0[0]),.dinb(n23231),.dout(n23232),.clk(gclk));
	jand g22975(.dina(n23232),.dinb(n23094),.dout(n23233),.clk(gclk));
	jand g22976(.dina(n23233),.dinb(w_n5606_21[0]),.dout(n23234),.clk(gclk));
	jor g22977(.dina(w_n22848_0[0]),.dinb(n23234),.dout(n23235),.clk(gclk));
	jand g22978(.dina(n23235),.dinb(n23093),.dout(n23236),.clk(gclk));
	jand g22979(.dina(n23236),.dinb(w_n5259_17[2]),.dout(n23237),.clk(gclk));
	jor g22980(.dina(w_n22856_0[0]),.dinb(n23237),.dout(n23238),.clk(gclk));
	jand g22981(.dina(n23238),.dinb(n23092),.dout(n23239),.clk(gclk));
	jand g22982(.dina(n23239),.dinb(w_n4902_21[2]),.dout(n23240),.clk(gclk));
	jnot g22983(.din(w_n22864_0[0]),.dout(n23241),.clk(gclk));
	jor g22984(.dina(w_n23241_0[1]),.dinb(n23240),.dout(n23242),.clk(gclk));
	jand g22985(.dina(n23242),.dinb(n23091),.dout(n23243),.clk(gclk));
	jand g22986(.dina(n23243),.dinb(w_n4582_18[2]),.dout(n23244),.clk(gclk));
	jor g22987(.dina(w_n22871_0[0]),.dinb(n23244),.dout(n23245),.clk(gclk));
	jand g22988(.dina(n23245),.dinb(n23090),.dout(n23246),.clk(gclk));
	jand g22989(.dina(n23246),.dinb(w_n4249_22[1]),.dout(n23247),.clk(gclk));
	jnot g22990(.din(w_n22879_0[0]),.dout(n23248),.clk(gclk));
	jor g22991(.dina(w_n23248_0[1]),.dinb(n23247),.dout(n23249),.clk(gclk));
	jand g22992(.dina(n23249),.dinb(n23089),.dout(n23250),.clk(gclk));
	jand g22993(.dina(n23250),.dinb(w_n3955_19[1]),.dout(n23251),.clk(gclk));
	jor g22994(.dina(w_n22886_0[0]),.dinb(n23251),.dout(n23252),.clk(gclk));
	jand g22995(.dina(n23252),.dinb(n23088),.dout(n23253),.clk(gclk));
	jand g22996(.dina(n23253),.dinb(w_n3642_22[2]),.dout(n23254),.clk(gclk));
	jnot g22997(.din(w_n22894_0[0]),.dout(n23255),.clk(gclk));
	jor g22998(.dina(w_n23255_0[1]),.dinb(n23254),.dout(n23256),.clk(gclk));
	jand g22999(.dina(n23256),.dinb(n23087),.dout(n23257),.clk(gclk));
	jand g23000(.dina(n23257),.dinb(w_n3368_20[0]),.dout(n23258),.clk(gclk));
	jor g23001(.dina(w_n22901_0[0]),.dinb(n23258),.dout(n23259),.clk(gclk));
	jand g23002(.dina(n23259),.dinb(n23086),.dout(n23260),.clk(gclk));
	jand g23003(.dina(n23260),.dinb(w_n3089_23[1]),.dout(n23261),.clk(gclk));
	jnot g23004(.din(w_n22909_0[0]),.dout(n23262),.clk(gclk));
	jor g23005(.dina(w_n23262_0[1]),.dinb(n23261),.dout(n23263),.clk(gclk));
	jand g23006(.dina(n23263),.dinb(n23085),.dout(n23264),.clk(gclk));
	jand g23007(.dina(n23264),.dinb(w_n2833_21[0]),.dout(n23265),.clk(gclk));
	jor g23008(.dina(w_n22916_0[0]),.dinb(n23265),.dout(n23266),.clk(gclk));
	jand g23009(.dina(n23266),.dinb(n23084),.dout(n23267),.clk(gclk));
	jand g23010(.dina(n23267),.dinb(w_n2572_23[2]),.dout(n23268),.clk(gclk));
	jor g23011(.dina(w_n22924_0[0]),.dinb(n23268),.dout(n23269),.clk(gclk));
	jand g23012(.dina(n23269),.dinb(n23083),.dout(n23270),.clk(gclk));
	jand g23013(.dina(n23270),.dinb(w_n2345_21[2]),.dout(n23271),.clk(gclk));
	jor g23014(.dina(w_n22932_0[0]),.dinb(n23271),.dout(n23272),.clk(gclk));
	jand g23015(.dina(n23272),.dinb(n23082),.dout(n23273),.clk(gclk));
	jand g23016(.dina(n23273),.dinb(w_n2108_24[1]),.dout(n23274),.clk(gclk));
	jnot g23017(.din(w_n22940_0[0]),.dout(n23275),.clk(gclk));
	jor g23018(.dina(w_n23275_0[1]),.dinb(n23274),.dout(n23276),.clk(gclk));
	jand g23019(.dina(n23276),.dinb(n23081),.dout(n23277),.clk(gclk));
	jand g23020(.dina(n23277),.dinb(w_n1912_22[2]),.dout(n23278),.clk(gclk));
	jor g23021(.dina(w_n22947_0[0]),.dinb(n23278),.dout(n23279),.clk(gclk));
	jand g23022(.dina(n23279),.dinb(n23080),.dout(n23280),.clk(gclk));
	jand g23023(.dina(n23280),.dinb(w_n1699_25[0]),.dout(n23281),.clk(gclk));
	jor g23024(.dina(w_n22955_0[0]),.dinb(n23281),.dout(n23282),.clk(gclk));
	jand g23025(.dina(n23282),.dinb(n23079),.dout(n23283),.clk(gclk));
	jand g23026(.dina(n23283),.dinb(w_n1516_23[1]),.dout(n23284),.clk(gclk));
	jor g23027(.dina(w_n22963_0[0]),.dinb(n23284),.dout(n23285),.clk(gclk));
	jand g23028(.dina(n23285),.dinb(n23078),.dout(n23286),.clk(gclk));
	jand g23029(.dina(n23286),.dinb(w_n1332_25[0]),.dout(n23287),.clk(gclk));
	jor g23030(.dina(w_n22971_0[0]),.dinb(n23287),.dout(n23288),.clk(gclk));
	jand g23031(.dina(n23288),.dinb(n23077),.dout(n23289),.clk(gclk));
	jand g23032(.dina(n23289),.dinb(w_n1173_24[0]),.dout(n23290),.clk(gclk));
	jor g23033(.dina(w_n22979_0[0]),.dinb(n23290),.dout(n23291),.clk(gclk));
	jand g23034(.dina(n23291),.dinb(n23076),.dout(n23292),.clk(gclk));
	jand g23035(.dina(n23292),.dinb(w_n1008_26[0]),.dout(n23293),.clk(gclk));
	jnot g23036(.din(w_n22987_0[0]),.dout(n23294),.clk(gclk));
	jor g23037(.dina(w_n23294_0[1]),.dinb(n23293),.dout(n23295),.clk(gclk));
	jand g23038(.dina(n23295),.dinb(n23075),.dout(n23296),.clk(gclk));
	jand g23039(.dina(n23296),.dinb(w_n884_25[0]),.dout(n23297),.clk(gclk));
	jor g23040(.dina(w_n22994_0[0]),.dinb(n23297),.dout(n23298),.clk(gclk));
	jand g23041(.dina(n23298),.dinb(n23074),.dout(n23299),.clk(gclk));
	jand g23042(.dina(n23299),.dinb(w_n743_26[0]),.dout(n23300),.clk(gclk));
	jnot g23043(.din(w_n23002_0[0]),.dout(n23301),.clk(gclk));
	jor g23044(.dina(w_n23301_0[1]),.dinb(n23300),.dout(n23302),.clk(gclk));
	jand g23045(.dina(n23302),.dinb(n23073),.dout(n23303),.clk(gclk));
	jand g23046(.dina(n23303),.dinb(w_n635_26[0]),.dout(n23304),.clk(gclk));
	jor g23047(.dina(w_n23009_0[0]),.dinb(n23304),.dout(n23305),.clk(gclk));
	jand g23048(.dina(n23305),.dinb(n23072),.dout(n23306),.clk(gclk));
	jand g23049(.dina(n23306),.dinb(w_n515_27[0]),.dout(n23307),.clk(gclk));
	jor g23050(.dina(w_n23017_0[0]),.dinb(n23307),.dout(n23308),.clk(gclk));
	jand g23051(.dina(n23308),.dinb(n23071),.dout(n23309),.clk(gclk));
	jand g23052(.dina(n23309),.dinb(w_n443_27[0]),.dout(n23310),.clk(gclk));
	jnot g23053(.din(w_n23025_0[0]),.dout(n23311),.clk(gclk));
	jor g23054(.dina(w_n23311_0[1]),.dinb(n23310),.dout(n23312),.clk(gclk));
	jand g23055(.dina(n23312),.dinb(n23070),.dout(n23313),.clk(gclk));
	jand g23056(.dina(n23313),.dinb(w_n352_27[1]),.dout(n23314),.clk(gclk));
	jnot g23057(.din(w_n23032_0[0]),.dout(n23315),.clk(gclk));
	jor g23058(.dina(w_n23315_0[1]),.dinb(n23314),.dout(n23316),.clk(gclk));
	jand g23059(.dina(n23316),.dinb(n23069),.dout(n23317),.clk(gclk));
	jand g23060(.dina(n23317),.dinb(w_n294_27[2]),.dout(n23318),.clk(gclk));
	jor g23061(.dina(w_n23039_0[0]),.dinb(n23318),.dout(n23319),.clk(gclk));
	jand g23062(.dina(n23319),.dinb(n23068),.dout(n23320),.clk(gclk));
	jand g23063(.dina(n23320),.dinb(w_n239_27[2]),.dout(n23321),.clk(gclk));
	jor g23064(.dina(w_n23047_0[0]),.dinb(n23321),.dout(n23322),.clk(gclk));
	jand g23065(.dina(n23322),.dinb(n23067),.dout(n23323),.clk(gclk));
	jand g23066(.dina(n23323),.dinb(w_n221_28[0]),.dout(n23324),.clk(gclk));
	jor g23067(.dina(w_n23055_0[1]),.dinb(n23324),.dout(n23325),.clk(gclk));
	jand g23068(.dina(n23325),.dinb(n23066),.dout(n23326),.clk(gclk));
	jor g23069(.dina(w_n23061_0[0]),.dinb(w_n23326_0[1]),.dout(n23327),.clk(gclk));
	jor g23070(.dina(w_n23327_0[1]),.dinb(w_n22321_0[0]),.dout(n23328),.clk(gclk));
	jor g23071(.dina(n23328),.dinb(w_n23065_0[1]),.dout(n23329),.clk(gclk));
	jand g23072(.dina(n23329),.dinb(w_n218_11[2]),.dout(n23330),.clk(gclk));
	jand g23073(.dina(w_n22619_0[0]),.dinb(w_n22317_0[2]),.dout(n23331),.clk(gclk));
	jnot g23074(.din(n23331),.dout(n23332),.clk(gclk));
	jxor g23075(.dina(w_n22320_0[1]),.dinb(w_n22317_0[1]),.dout(n23333),.clk(gclk));
	jand g23076(.dina(n23333),.dinb(n23332),.dout(n23334),.clk(gclk));
	jand g23077(.dina(n23334),.dinb(w_asqrt63_20[1]),.dout(n23335),.clk(gclk));
	jor g23078(.dina(w_n23335_0[1]),.dinb(n23330),.dout(n23336),.clk(gclk));
	jor g23079(.dina(w_n23336_0[1]),.dinb(w_n23064_0[1]),.dout(asqrt_fa_4),.clk(gclk));
	jnot g23080(.din(w_n23065_0[0]),.dout(n23338),.clk(gclk));
	jand g23081(.dina(w_n23062_0[0]),.dinb(w_n23058_0[0]),.dout(n23339),.clk(gclk));
	jand g23082(.dina(w_n23339_0[1]),.dinb(w_n22345_0[0]),.dout(n23340),.clk(gclk));
	jand g23083(.dina(n23340),.dinb(n23338),.dout(n23341),.clk(gclk));
	jor g23084(.dina(n23341),.dinb(w_asqrt63_20[0]),.dout(n23342),.clk(gclk));
	jnot g23085(.din(w_n23335_0[0]),.dout(n23343),.clk(gclk));
	jand g23086(.dina(n23343),.dinb(n23342),.dout(n23344),.clk(gclk));
	jand g23087(.dina(w_n23344_0[1]),.dinb(w_n23063_1[0]),.dout(n23345),.clk(gclk));
	jxor g23088(.dina(w_n23050_0[0]),.dinb(w_n221_27[2]),.dout(n23346),.clk(gclk));
	jor g23089(.dina(n23346),.dinb(w_n23345_32[1]),.dout(n23347),.clk(gclk));
	jxor g23090(.dina(n23347),.dinb(w_n23055_0[0]),.dout(n23348),.clk(gclk));
	jnot g23091(.din(w_n23348_0[1]),.dout(n23349),.clk(gclk));
	jor g23092(.dina(w_n23345_32[0]),.dinb(w_n22334_1[1]),.dout(n23350),.clk(gclk));
	jnot g23093(.din(w_a4_1[1]),.dout(n23351),.clk(gclk));
	jnot g23094(.din(w_a5_0[1]),.dout(n23352),.clk(gclk));
	jand g23095(.dina(w_n23352_0[1]),.dinb(w_n23351_1[1]),.dout(n23353),.clk(gclk));
	jand g23096(.dina(w_n23353_0[2]),.dinb(w_n22334_1[0]),.dout(n23354),.clk(gclk));
	jnot g23097(.din(w_n23354_0[1]),.dout(n23355),.clk(gclk));
	jand g23098(.dina(n23355),.dinb(n23350),.dout(n23356),.clk(gclk));
	jor g23099(.dina(w_n23356_0[2]),.dinb(w_n22620_3[2]),.dout(n23357),.clk(gclk));
	jand g23100(.dina(w_n23356_0[1]),.dinb(w_n22620_3[1]),.dout(n23358),.clk(gclk));
	jor g23101(.dina(w_n23345_31[2]),.dinb(w_a6_0[1]),.dout(n23359),.clk(gclk));
	jand g23102(.dina(n23359),.dinb(w_a7_0[0]),.dout(n23360),.clk(gclk));
	jand g23103(.dina(w_asqrt3_2[1]),.dinb(w_n22336_0[1]),.dout(n23361),.clk(gclk));
	jor g23104(.dina(n23361),.dinb(n23360),.dout(n23362),.clk(gclk));
	jor g23105(.dina(n23362),.dinb(n23358),.dout(n23363),.clk(gclk));
	jand g23106(.dina(n23363),.dinb(w_n23357_0[1]),.dout(n23364),.clk(gclk));
	jor g23107(.dina(w_n23364_0[2]),.dinb(w_n21887_13[2]),.dout(n23365),.clk(gclk));
	jand g23108(.dina(w_n23364_0[1]),.dinb(w_n21887_13[1]),.dout(n23366),.clk(gclk));
	jnot g23109(.din(w_n22336_0[0]),.dout(n23367),.clk(gclk));
	jor g23110(.dina(w_n23345_31[1]),.dinb(n23367),.dout(n23368),.clk(gclk));
	jor g23111(.dina(w_asqrt3_2[0]),.dinb(w_n22620_3[0]),.dout(n23369),.clk(gclk));
	jand g23112(.dina(n23369),.dinb(w_n23368_0[1]),.dout(n23370),.clk(gclk));
	jxor g23113(.dina(n23370),.dinb(w_n21889_0[1]),.dout(n23371),.clk(gclk));
	jor g23114(.dina(w_n23371_0[1]),.dinb(n23366),.dout(n23372),.clk(gclk));
	jand g23115(.dina(n23372),.dinb(w_n23365_0[1]),.dout(n23373),.clk(gclk));
	jor g23116(.dina(w_n23373_0[2]),.dinb(w_n21184_4[2]),.dout(n23374),.clk(gclk));
	jand g23117(.dina(w_n23373_0[1]),.dinb(w_n21184_4[1]),.dout(n23375),.clk(gclk));
	jxor g23118(.dina(w_n22339_0[0]),.dinb(w_n21887_13[0]),.dout(n23376),.clk(gclk));
	jor g23119(.dina(n23376),.dinb(w_n23345_31[0]),.dout(n23377),.clk(gclk));
	jxor g23120(.dina(n23377),.dinb(w_n22622_0[0]),.dout(n23378),.clk(gclk));
	jor g23121(.dina(w_n23378_0[2]),.dinb(n23375),.dout(n23379),.clk(gclk));
	jand g23122(.dina(n23379),.dinb(w_n23374_0[1]),.dout(n23380),.clk(gclk));
	jor g23123(.dina(w_n23380_0[2]),.dinb(w_n20468_14[0]),.dout(n23381),.clk(gclk));
	jand g23124(.dina(w_n23380_0[1]),.dinb(w_n20468_13[2]),.dout(n23382),.clk(gclk));
	jxor g23125(.dina(w_n22624_0[0]),.dinb(w_n21184_4[0]),.dout(n23383),.clk(gclk));
	jor g23126(.dina(n23383),.dinb(w_n23345_30[2]),.dout(n23384),.clk(gclk));
	jxor g23127(.dina(n23384),.dinb(w_n22630_0[0]),.dout(n23385),.clk(gclk));
	jor g23128(.dina(w_n23385_0[2]),.dinb(n23382),.dout(n23386),.clk(gclk));
	jand g23129(.dina(n23386),.dinb(w_n23381_0[1]),.dout(n23387),.clk(gclk));
	jor g23130(.dina(w_n23387_0[2]),.dinb(w_n19791_5[2]),.dout(n23388),.clk(gclk));
	jand g23131(.dina(w_n23387_0[1]),.dinb(w_n19791_5[1]),.dout(n23389),.clk(gclk));
	jxor g23132(.dina(w_n22632_0[0]),.dinb(w_n20468_13[1]),.dout(n23390),.clk(gclk));
	jor g23133(.dina(n23390),.dinb(w_n23345_30[1]),.dout(n23391),.clk(gclk));
	jxor g23134(.dina(n23391),.dinb(w_n23138_0[0]),.dout(n23392),.clk(gclk));
	jnot g23135(.din(w_n23392_0[2]),.dout(n23393),.clk(gclk));
	jor g23136(.dina(n23393),.dinb(n23389),.dout(n23394),.clk(gclk));
	jand g23137(.dina(n23394),.dinb(w_n23388_0[1]),.dout(n23395),.clk(gclk));
	jor g23138(.dina(w_n23395_0[2]),.dinb(w_n19096_14[1]),.dout(n23396),.clk(gclk));
	jand g23139(.dina(w_n23395_0[1]),.dinb(w_n19096_14[0]),.dout(n23397),.clk(gclk));
	jxor g23140(.dina(w_n22639_0[0]),.dinb(w_n19791_5[0]),.dout(n23398),.clk(gclk));
	jor g23141(.dina(n23398),.dinb(w_n23345_30[0]),.dout(n23399),.clk(gclk));
	jxor g23142(.dina(n23399),.dinb(w_n23142_0[0]),.dout(n23400),.clk(gclk));
	jnot g23143(.din(w_n23400_0[2]),.dout(n23401),.clk(gclk));
	jor g23144(.dina(n23401),.dinb(n23397),.dout(n23402),.clk(gclk));
	jand g23145(.dina(n23402),.dinb(w_n23396_0[1]),.dout(n23403),.clk(gclk));
	jor g23146(.dina(w_n23403_0[2]),.dinb(w_n18442_6[1]),.dout(n23404),.clk(gclk));
	jand g23147(.dina(w_n23403_0[1]),.dinb(w_n18442_6[0]),.dout(n23405),.clk(gclk));
	jxor g23148(.dina(w_n22646_0[0]),.dinb(w_n19096_13[2]),.dout(n23406),.clk(gclk));
	jor g23149(.dina(n23406),.dinb(w_n23345_29[2]),.dout(n23407),.clk(gclk));
	jxor g23150(.dina(n23407),.dinb(w_n23146_0[0]),.dout(n23408),.clk(gclk));
	jnot g23151(.din(w_n23408_0[2]),.dout(n23409),.clk(gclk));
	jor g23152(.dina(n23409),.dinb(n23405),.dout(n23410),.clk(gclk));
	jand g23153(.dina(n23410),.dinb(w_n23404_0[1]),.dout(n23411),.clk(gclk));
	jor g23154(.dina(w_n23411_0[2]),.dinb(w_n17769_15[0]),.dout(n23412),.clk(gclk));
	jand g23155(.dina(w_n23411_0[1]),.dinb(w_n17769_14[2]),.dout(n23413),.clk(gclk));
	jxor g23156(.dina(w_n22653_0[0]),.dinb(w_n18442_5[2]),.dout(n23414),.clk(gclk));
	jor g23157(.dina(n23414),.dinb(w_n23345_29[1]),.dout(n23415),.clk(gclk));
	jxor g23158(.dina(n23415),.dinb(w_n22659_0[0]),.dout(n23416),.clk(gclk));
	jor g23159(.dina(w_n23416_0[2]),.dinb(n23413),.dout(n23417),.clk(gclk));
	jand g23160(.dina(n23417),.dinb(w_n23412_0[1]),.dout(n23418),.clk(gclk));
	jor g23161(.dina(w_n23418_0[2]),.dinb(w_n17134_7[1]),.dout(n23419),.clk(gclk));
	jand g23162(.dina(w_n23418_0[1]),.dinb(w_n17134_7[0]),.dout(n23420),.clk(gclk));
	jxor g23163(.dina(w_n22661_0[0]),.dinb(w_n17769_14[1]),.dout(n23421),.clk(gclk));
	jor g23164(.dina(n23421),.dinb(w_n23345_29[0]),.dout(n23422),.clk(gclk));
	jxor g23165(.dina(n23422),.dinb(w_n23153_0[0]),.dout(n23423),.clk(gclk));
	jnot g23166(.din(w_n23423_0[2]),.dout(n23424),.clk(gclk));
	jor g23167(.dina(n23424),.dinb(n23420),.dout(n23425),.clk(gclk));
	jand g23168(.dina(n23425),.dinb(w_n23419_0[1]),.dout(n23426),.clk(gclk));
	jor g23169(.dina(w_n23426_0[2]),.dinb(w_n16489_15[1]),.dout(n23427),.clk(gclk));
	jand g23170(.dina(w_n23426_0[1]),.dinb(w_n16489_15[0]),.dout(n23428),.clk(gclk));
	jxor g23171(.dina(w_n22668_0[0]),.dinb(w_n17134_6[2]),.dout(n23429),.clk(gclk));
	jor g23172(.dina(n23429),.dinb(w_n23345_28[2]),.dout(n23430),.clk(gclk));
	jxor g23173(.dina(n23430),.dinb(w_n22674_0[0]),.dout(n23431),.clk(gclk));
	jor g23174(.dina(w_n23431_0[2]),.dinb(n23428),.dout(n23432),.clk(gclk));
	jand g23175(.dina(n23432),.dinb(w_n23427_0[1]),.dout(n23433),.clk(gclk));
	jor g23176(.dina(w_n23433_0[2]),.dinb(w_n15878_8[1]),.dout(n23434),.clk(gclk));
	jand g23177(.dina(w_n23433_0[1]),.dinb(w_n15878_8[0]),.dout(n23435),.clk(gclk));
	jxor g23178(.dina(w_n22676_0[0]),.dinb(w_n16489_14[2]),.dout(n23436),.clk(gclk));
	jor g23179(.dina(n23436),.dinb(w_n23345_28[1]),.dout(n23437),.clk(gclk));
	jxor g23180(.dina(n23437),.dinb(w_n23160_0[0]),.dout(n23438),.clk(gclk));
	jnot g23181(.din(w_n23438_0[2]),.dout(n23439),.clk(gclk));
	jor g23182(.dina(n23439),.dinb(n23435),.dout(n23440),.clk(gclk));
	jand g23183(.dina(n23440),.dinb(w_n23434_0[1]),.dout(n23441),.clk(gclk));
	jor g23184(.dina(w_n23441_0[2]),.dinb(w_n15260_16[0]),.dout(n23442),.clk(gclk));
	jand g23185(.dina(w_n23441_0[1]),.dinb(w_n15260_15[2]),.dout(n23443),.clk(gclk));
	jxor g23186(.dina(w_n22683_0[0]),.dinb(w_n15878_7[2]),.dout(n23444),.clk(gclk));
	jor g23187(.dina(n23444),.dinb(w_n23345_28[0]),.dout(n23445),.clk(gclk));
	jxor g23188(.dina(n23445),.dinb(w_n22689_0[0]),.dout(n23446),.clk(gclk));
	jor g23189(.dina(w_n23446_0[2]),.dinb(n23443),.dout(n23447),.clk(gclk));
	jand g23190(.dina(n23447),.dinb(w_n23442_0[1]),.dout(n23448),.clk(gclk));
	jor g23191(.dina(w_n23448_0[2]),.dinb(w_n14674_9[0]),.dout(n23449),.clk(gclk));
	jand g23192(.dina(w_n23448_0[1]),.dinb(w_n14674_8[2]),.dout(n23450),.clk(gclk));
	jxor g23193(.dina(w_n22691_0[0]),.dinb(w_n15260_15[1]),.dout(n23451),.clk(gclk));
	jor g23194(.dina(n23451),.dinb(w_n23345_27[2]),.dout(n23452),.clk(gclk));
	jxor g23195(.dina(n23452),.dinb(w_n22697_0[0]),.dout(n23453),.clk(gclk));
	jor g23196(.dina(w_n23453_0[2]),.dinb(n23450),.dout(n23454),.clk(gclk));
	jand g23197(.dina(n23454),.dinb(w_n23449_0[1]),.dout(n23455),.clk(gclk));
	jor g23198(.dina(w_n23455_0[2]),.dinb(w_n14078_16[1]),.dout(n23456),.clk(gclk));
	jand g23199(.dina(w_n23455_0[1]),.dinb(w_n14078_16[0]),.dout(n23457),.clk(gclk));
	jxor g23200(.dina(w_n22699_0[0]),.dinb(w_n14674_8[1]),.dout(n23458),.clk(gclk));
	jor g23201(.dina(n23458),.dinb(w_n23345_27[1]),.dout(n23459),.clk(gclk));
	jxor g23202(.dina(n23459),.dinb(w_n22705_0[0]),.dout(n23460),.clk(gclk));
	jor g23203(.dina(w_n23460_0[2]),.dinb(n23457),.dout(n23461),.clk(gclk));
	jand g23204(.dina(n23461),.dinb(w_n23456_0[1]),.dout(n23462),.clk(gclk));
	jor g23205(.dina(w_n23462_0[2]),.dinb(w_n13515_10[0]),.dout(n23463),.clk(gclk));
	jand g23206(.dina(w_n23462_0[1]),.dinb(w_n13515_9[2]),.dout(n23464),.clk(gclk));
	jxor g23207(.dina(w_n22707_0[0]),.dinb(w_n14078_15[2]),.dout(n23465),.clk(gclk));
	jor g23208(.dina(n23465),.dinb(w_n23345_27[0]),.dout(n23466),.clk(gclk));
	jxor g23209(.dina(n23466),.dinb(w_n23173_0[0]),.dout(n23467),.clk(gclk));
	jnot g23210(.din(w_n23467_0[2]),.dout(n23468),.clk(gclk));
	jor g23211(.dina(n23468),.dinb(n23464),.dout(n23469),.clk(gclk));
	jand g23212(.dina(n23469),.dinb(w_n23463_0[1]),.dout(n23470),.clk(gclk));
	jor g23213(.dina(w_n23470_0[2]),.dinb(w_n12947_17[0]),.dout(n23471),.clk(gclk));
	jand g23214(.dina(w_n23470_0[1]),.dinb(w_n12947_16[2]),.dout(n23472),.clk(gclk));
	jxor g23215(.dina(w_n22714_0[0]),.dinb(w_n13515_9[1]),.dout(n23473),.clk(gclk));
	jor g23216(.dina(n23473),.dinb(w_n23345_26[2]),.dout(n23474),.clk(gclk));
	jxor g23217(.dina(n23474),.dinb(w_n22720_0[0]),.dout(n23475),.clk(gclk));
	jor g23218(.dina(w_n23475_0[2]),.dinb(n23472),.dout(n23476),.clk(gclk));
	jand g23219(.dina(n23476),.dinb(w_n23471_0[1]),.dout(n23477),.clk(gclk));
	jor g23220(.dina(w_n23477_0[2]),.dinb(w_n12410_10[2]),.dout(n23478),.clk(gclk));
	jand g23221(.dina(w_n23477_0[1]),.dinb(w_n12410_10[1]),.dout(n23479),.clk(gclk));
	jxor g23222(.dina(w_n22722_0[0]),.dinb(w_n12947_16[1]),.dout(n23480),.clk(gclk));
	jor g23223(.dina(n23480),.dinb(w_n23345_26[1]),.dout(n23481),.clk(gclk));
	jxor g23224(.dina(n23481),.dinb(w_n22728_0[0]),.dout(n23482),.clk(gclk));
	jor g23225(.dina(w_n23482_0[2]),.dinb(n23479),.dout(n23483),.clk(gclk));
	jand g23226(.dina(n23483),.dinb(w_n23478_0[1]),.dout(n23484),.clk(gclk));
	jor g23227(.dina(w_n23484_0[2]),.dinb(w_n11858_17[1]),.dout(n23485),.clk(gclk));
	jand g23228(.dina(w_n23484_0[1]),.dinb(w_n11858_17[0]),.dout(n23486),.clk(gclk));
	jxor g23229(.dina(w_n22730_0[0]),.dinb(w_n12410_10[0]),.dout(n23487),.clk(gclk));
	jor g23230(.dina(n23487),.dinb(w_n23345_26[0]),.dout(n23488),.clk(gclk));
	jxor g23231(.dina(n23488),.dinb(w_n22736_0[0]),.dout(n23489),.clk(gclk));
	jor g23232(.dina(w_n23489_0[2]),.dinb(n23486),.dout(n23490),.clk(gclk));
	jand g23233(.dina(n23490),.dinb(w_n23485_0[1]),.dout(n23491),.clk(gclk));
	jor g23234(.dina(w_n23491_0[2]),.dinb(w_n11347_11[1]),.dout(n23492),.clk(gclk));
	jand g23235(.dina(w_n23491_0[1]),.dinb(w_n11347_11[0]),.dout(n23493),.clk(gclk));
	jxor g23236(.dina(w_n22738_0[0]),.dinb(w_n11858_16[2]),.dout(n23494),.clk(gclk));
	jor g23237(.dina(n23494),.dinb(w_n23345_25[2]),.dout(n23495),.clk(gclk));
	jxor g23238(.dina(n23495),.dinb(w_n23186_0[0]),.dout(n23496),.clk(gclk));
	jnot g23239(.din(w_n23496_0[2]),.dout(n23497),.clk(gclk));
	jor g23240(.dina(n23497),.dinb(n23493),.dout(n23498),.clk(gclk));
	jand g23241(.dina(n23498),.dinb(w_n23492_0[1]),.dout(n23499),.clk(gclk));
	jor g23242(.dina(w_n23499_0[2]),.dinb(w_n10824_18[0]),.dout(n23500),.clk(gclk));
	jand g23243(.dina(w_n23499_0[1]),.dinb(w_n10824_17[2]),.dout(n23501),.clk(gclk));
	jxor g23244(.dina(w_n22745_0[0]),.dinb(w_n11347_10[2]),.dout(n23502),.clk(gclk));
	jor g23245(.dina(n23502),.dinb(w_n23345_25[1]),.dout(n23503),.clk(gclk));
	jxor g23246(.dina(n23503),.dinb(w_n22751_0[0]),.dout(n23504),.clk(gclk));
	jor g23247(.dina(w_n23504_0[2]),.dinb(n23501),.dout(n23505),.clk(gclk));
	jand g23248(.dina(n23505),.dinb(w_n23500_0[1]),.dout(n23506),.clk(gclk));
	jor g23249(.dina(w_n23506_0[2]),.dinb(w_n10328_12[1]),.dout(n23507),.clk(gclk));
	jand g23250(.dina(w_n23506_0[1]),.dinb(w_n10328_12[0]),.dout(n23508),.clk(gclk));
	jxor g23251(.dina(w_n22753_0[0]),.dinb(w_n10824_17[1]),.dout(n23509),.clk(gclk));
	jor g23252(.dina(n23509),.dinb(w_n23345_25[0]),.dout(n23510),.clk(gclk));
	jxor g23253(.dina(n23510),.dinb(w_n23193_0[0]),.dout(n23511),.clk(gclk));
	jnot g23254(.din(w_n23511_0[2]),.dout(n23512),.clk(gclk));
	jor g23255(.dina(n23512),.dinb(n23508),.dout(n23513),.clk(gclk));
	jand g23256(.dina(n23513),.dinb(w_n23507_0[1]),.dout(n23514),.clk(gclk));
	jor g23257(.dina(w_n23514_0[2]),.dinb(w_n9832_18[2]),.dout(n23515),.clk(gclk));
	jand g23258(.dina(w_n23514_0[1]),.dinb(w_n9832_18[1]),.dout(n23516),.clk(gclk));
	jxor g23259(.dina(w_n22760_0[0]),.dinb(w_n10328_11[2]),.dout(n23517),.clk(gclk));
	jor g23260(.dina(n23517),.dinb(w_n23345_24[2]),.dout(n23518),.clk(gclk));
	jxor g23261(.dina(n23518),.dinb(w_n22766_0[0]),.dout(n23519),.clk(gclk));
	jor g23262(.dina(w_n23519_0[2]),.dinb(n23516),.dout(n23520),.clk(gclk));
	jand g23263(.dina(n23520),.dinb(w_n23515_0[1]),.dout(n23521),.clk(gclk));
	jor g23264(.dina(w_n23521_0[2]),.dinb(w_n9369_13[1]),.dout(n23522),.clk(gclk));
	jand g23265(.dina(w_n23521_0[1]),.dinb(w_n9369_13[0]),.dout(n23523),.clk(gclk));
	jxor g23266(.dina(w_n22768_0[0]),.dinb(w_n9832_18[0]),.dout(n23524),.clk(gclk));
	jor g23267(.dina(n23524),.dinb(w_n23345_24[1]),.dout(n23525),.clk(gclk));
	jxor g23268(.dina(n23525),.dinb(w_n23200_0[0]),.dout(n23526),.clk(gclk));
	jnot g23269(.din(w_n23526_0[2]),.dout(n23527),.clk(gclk));
	jor g23270(.dina(n23527),.dinb(n23523),.dout(n23528),.clk(gclk));
	jand g23271(.dina(n23528),.dinb(w_n23522_0[1]),.dout(n23529),.clk(gclk));
	jor g23272(.dina(w_n23529_0[2]),.dinb(w_n8890_19[0]),.dout(n23530),.clk(gclk));
	jand g23273(.dina(w_n23529_0[1]),.dinb(w_n8890_18[2]),.dout(n23531),.clk(gclk));
	jxor g23274(.dina(w_n22775_0[0]),.dinb(w_n9369_12[2]),.dout(n23532),.clk(gclk));
	jor g23275(.dina(n23532),.dinb(w_n23345_24[0]),.dout(n23533),.clk(gclk));
	jxor g23276(.dina(n23533),.dinb(w_n22781_0[0]),.dout(n23534),.clk(gclk));
	jor g23277(.dina(w_n23534_0[2]),.dinb(n23531),.dout(n23535),.clk(gclk));
	jand g23278(.dina(n23535),.dinb(w_n23530_0[1]),.dout(n23536),.clk(gclk));
	jor g23279(.dina(w_n23536_0[2]),.dinb(w_n8449_14[0]),.dout(n23537),.clk(gclk));
	jand g23280(.dina(w_n23536_0[1]),.dinb(w_n8449_13[2]),.dout(n23538),.clk(gclk));
	jxor g23281(.dina(w_n22783_0[0]),.dinb(w_n8890_18[1]),.dout(n23539),.clk(gclk));
	jor g23282(.dina(n23539),.dinb(w_n23345_23[2]),.dout(n23540),.clk(gclk));
	jxor g23283(.dina(n23540),.dinb(w_n22789_0[0]),.dout(n23541),.clk(gclk));
	jor g23284(.dina(w_n23541_0[2]),.dinb(n23538),.dout(n23542),.clk(gclk));
	jand g23285(.dina(n23542),.dinb(w_n23537_0[1]),.dout(n23543),.clk(gclk));
	jor g23286(.dina(w_n23543_0[2]),.dinb(w_n8003_19[2]),.dout(n23544),.clk(gclk));
	jand g23287(.dina(w_n23543_0[1]),.dinb(w_n8003_19[1]),.dout(n23545),.clk(gclk));
	jxor g23288(.dina(w_n22791_0[0]),.dinb(w_n8449_13[1]),.dout(n23546),.clk(gclk));
	jor g23289(.dina(n23546),.dinb(w_n23345_23[1]),.dout(n23547),.clk(gclk));
	jxor g23290(.dina(n23547),.dinb(w_n23210_0[0]),.dout(n23548),.clk(gclk));
	jnot g23291(.din(w_n23548_0[2]),.dout(n23549),.clk(gclk));
	jor g23292(.dina(n23549),.dinb(n23545),.dout(n23550),.clk(gclk));
	jand g23293(.dina(n23550),.dinb(w_n23544_0[1]),.dout(n23551),.clk(gclk));
	jor g23294(.dina(w_n23551_0[2]),.dinb(w_n7581_15[0]),.dout(n23552),.clk(gclk));
	jand g23295(.dina(w_n23551_0[1]),.dinb(w_n7581_14[2]),.dout(n23553),.clk(gclk));
	jxor g23296(.dina(w_n22798_0[0]),.dinb(w_n8003_19[0]),.dout(n23554),.clk(gclk));
	jor g23297(.dina(n23554),.dinb(w_n23345_23[0]),.dout(n23555),.clk(gclk));
	jxor g23298(.dina(n23555),.dinb(w_n23214_0[0]),.dout(n23556),.clk(gclk));
	jnot g23299(.din(w_n23556_0[2]),.dout(n23557),.clk(gclk));
	jor g23300(.dina(n23557),.dinb(n23553),.dout(n23558),.clk(gclk));
	jand g23301(.dina(n23558),.dinb(w_n23552_0[1]),.dout(n23559),.clk(gclk));
	jor g23302(.dina(w_n23559_0[2]),.dinb(w_n7154_20[0]),.dout(n23560),.clk(gclk));
	jand g23303(.dina(w_n23559_0[1]),.dinb(w_n7154_19[2]),.dout(n23561),.clk(gclk));
	jxor g23304(.dina(w_n22805_0[0]),.dinb(w_n7581_14[1]),.dout(n23562),.clk(gclk));
	jor g23305(.dina(n23562),.dinb(w_n23345_22[2]),.dout(n23563),.clk(gclk));
	jxor g23306(.dina(n23563),.dinb(w_n22811_0[0]),.dout(n23564),.clk(gclk));
	jor g23307(.dina(w_n23564_0[2]),.dinb(n23561),.dout(n23565),.clk(gclk));
	jand g23308(.dina(n23565),.dinb(w_n23560_0[1]),.dout(n23566),.clk(gclk));
	jor g23309(.dina(w_n23566_0[2]),.dinb(w_n6758_15[2]),.dout(n23567),.clk(gclk));
	jand g23310(.dina(w_n23566_0[1]),.dinb(w_n6758_15[1]),.dout(n23568),.clk(gclk));
	jxor g23311(.dina(w_n22813_0[0]),.dinb(w_n7154_19[1]),.dout(n23569),.clk(gclk));
	jor g23312(.dina(n23569),.dinb(w_n23345_22[1]),.dout(n23570),.clk(gclk));
	jxor g23313(.dina(n23570),.dinb(w_n23221_0[0]),.dout(n23571),.clk(gclk));
	jnot g23314(.din(w_n23571_0[2]),.dout(n23572),.clk(gclk));
	jor g23315(.dina(n23572),.dinb(n23568),.dout(n23573),.clk(gclk));
	jand g23316(.dina(n23573),.dinb(w_n23567_0[1]),.dout(n23574),.clk(gclk));
	jor g23317(.dina(w_n23574_0[2]),.dinb(w_n6357_20[1]),.dout(n23575),.clk(gclk));
	jand g23318(.dina(w_n23574_0[1]),.dinb(w_n6357_20[0]),.dout(n23576),.clk(gclk));
	jxor g23319(.dina(w_n22820_0[0]),.dinb(w_n6758_15[0]),.dout(n23577),.clk(gclk));
	jor g23320(.dina(n23577),.dinb(w_n23345_22[0]),.dout(n23578),.clk(gclk));
	jxor g23321(.dina(n23578),.dinb(w_n22826_0[0]),.dout(n23579),.clk(gclk));
	jor g23322(.dina(w_n23579_0[2]),.dinb(n23576),.dout(n23580),.clk(gclk));
	jand g23323(.dina(n23580),.dinb(w_n23575_0[1]),.dout(n23581),.clk(gclk));
	jor g23324(.dina(w_n23581_0[2]),.dinb(w_n5989_16[1]),.dout(n23582),.clk(gclk));
	jand g23325(.dina(w_n23581_0[1]),.dinb(w_n5989_16[0]),.dout(n23583),.clk(gclk));
	jxor g23326(.dina(w_n22828_0[0]),.dinb(w_n6357_19[2]),.dout(n23584),.clk(gclk));
	jor g23327(.dina(n23584),.dinb(w_n23345_21[2]),.dout(n23585),.clk(gclk));
	jxor g23328(.dina(n23585),.dinb(w_n23228_0[0]),.dout(n23586),.clk(gclk));
	jnot g23329(.din(w_n23586_0[2]),.dout(n23587),.clk(gclk));
	jor g23330(.dina(n23587),.dinb(n23583),.dout(n23588),.clk(gclk));
	jand g23331(.dina(n23588),.dinb(w_n23582_0[1]),.dout(n23589),.clk(gclk));
	jor g23332(.dina(w_n23589_0[2]),.dinb(w_n5606_20[2]),.dout(n23590),.clk(gclk));
	jand g23333(.dina(w_n23589_0[1]),.dinb(w_n5606_20[1]),.dout(n23591),.clk(gclk));
	jxor g23334(.dina(w_n22835_0[0]),.dinb(w_n5989_15[2]),.dout(n23592),.clk(gclk));
	jor g23335(.dina(n23592),.dinb(w_n23345_21[1]),.dout(n23593),.clk(gclk));
	jxor g23336(.dina(n23593),.dinb(w_n22841_0[0]),.dout(n23594),.clk(gclk));
	jor g23337(.dina(w_n23594_0[2]),.dinb(n23591),.dout(n23595),.clk(gclk));
	jand g23338(.dina(n23595),.dinb(w_n23590_0[1]),.dout(n23596),.clk(gclk));
	jor g23339(.dina(w_n23596_0[2]),.dinb(w_n5259_17[1]),.dout(n23597),.clk(gclk));
	jand g23340(.dina(w_n23596_0[1]),.dinb(w_n5259_17[0]),.dout(n23598),.clk(gclk));
	jxor g23341(.dina(w_n22843_0[0]),.dinb(w_n5606_20[0]),.dout(n23599),.clk(gclk));
	jor g23342(.dina(n23599),.dinb(w_n23345_21[0]),.dout(n23600),.clk(gclk));
	jxor g23343(.dina(n23600),.dinb(w_n22849_0[0]),.dout(n23601),.clk(gclk));
	jor g23344(.dina(w_n23601_0[2]),.dinb(n23598),.dout(n23602),.clk(gclk));
	jand g23345(.dina(n23602),.dinb(w_n23597_0[1]),.dout(n23603),.clk(gclk));
	jor g23346(.dina(w_n23603_0[2]),.dinb(w_n4902_21[1]),.dout(n23604),.clk(gclk));
	jand g23347(.dina(w_n23603_0[1]),.dinb(w_n4902_21[0]),.dout(n23605),.clk(gclk));
	jxor g23348(.dina(w_n22851_0[0]),.dinb(w_n5259_16[2]),.dout(n23606),.clk(gclk));
	jor g23349(.dina(n23606),.dinb(w_n23345_20[2]),.dout(n23607),.clk(gclk));
	jxor g23350(.dina(n23607),.dinb(w_n22857_0[0]),.dout(n23608),.clk(gclk));
	jor g23351(.dina(w_n23608_0[2]),.dinb(n23605),.dout(n23609),.clk(gclk));
	jand g23352(.dina(n23609),.dinb(w_n23604_0[1]),.dout(n23610),.clk(gclk));
	jor g23353(.dina(w_n23610_0[2]),.dinb(w_n4582_18[1]),.dout(n23611),.clk(gclk));
	jand g23354(.dina(w_n23610_0[1]),.dinb(w_n4582_18[0]),.dout(n23612),.clk(gclk));
	jxor g23355(.dina(w_n22859_0[0]),.dinb(w_n4902_20[2]),.dout(n23613),.clk(gclk));
	jor g23356(.dina(n23613),.dinb(w_n23345_20[1]),.dout(n23614),.clk(gclk));
	jxor g23357(.dina(n23614),.dinb(w_n23241_0[0]),.dout(n23615),.clk(gclk));
	jnot g23358(.din(w_n23615_0[2]),.dout(n23616),.clk(gclk));
	jor g23359(.dina(n23616),.dinb(n23612),.dout(n23617),.clk(gclk));
	jand g23360(.dina(n23617),.dinb(w_n23611_0[1]),.dout(n23618),.clk(gclk));
	jor g23361(.dina(w_n23618_0[2]),.dinb(w_n4249_22[0]),.dout(n23619),.clk(gclk));
	jand g23362(.dina(w_n23618_0[1]),.dinb(w_n4249_21[2]),.dout(n23620),.clk(gclk));
	jxor g23363(.dina(w_n22866_0[0]),.dinb(w_n4582_17[2]),.dout(n23621),.clk(gclk));
	jor g23364(.dina(n23621),.dinb(w_n23345_20[0]),.dout(n23622),.clk(gclk));
	jxor g23365(.dina(n23622),.dinb(w_n22872_0[0]),.dout(n23623),.clk(gclk));
	jor g23366(.dina(w_n23623_0[2]),.dinb(n23620),.dout(n23624),.clk(gclk));
	jand g23367(.dina(n23624),.dinb(w_n23619_0[1]),.dout(n23625),.clk(gclk));
	jor g23368(.dina(w_n23625_0[2]),.dinb(w_n3955_19[0]),.dout(n23626),.clk(gclk));
	jand g23369(.dina(w_n23625_0[1]),.dinb(w_n3955_18[2]),.dout(n23627),.clk(gclk));
	jxor g23370(.dina(w_n22874_0[0]),.dinb(w_n4249_21[1]),.dout(n23628),.clk(gclk));
	jor g23371(.dina(n23628),.dinb(w_n23345_19[2]),.dout(n23629),.clk(gclk));
	jxor g23372(.dina(n23629),.dinb(w_n23248_0[0]),.dout(n23630),.clk(gclk));
	jnot g23373(.din(w_n23630_0[2]),.dout(n23631),.clk(gclk));
	jor g23374(.dina(n23631),.dinb(n23627),.dout(n23632),.clk(gclk));
	jand g23375(.dina(n23632),.dinb(w_n23626_0[1]),.dout(n23633),.clk(gclk));
	jor g23376(.dina(w_n23633_0[2]),.dinb(w_n3642_22[1]),.dout(n23634),.clk(gclk));
	jand g23377(.dina(w_n23633_0[1]),.dinb(w_n3642_22[0]),.dout(n23635),.clk(gclk));
	jxor g23378(.dina(w_n22881_0[0]),.dinb(w_n3955_18[1]),.dout(n23636),.clk(gclk));
	jor g23379(.dina(n23636),.dinb(w_n23345_19[1]),.dout(n23637),.clk(gclk));
	jxor g23380(.dina(n23637),.dinb(w_n22887_0[0]),.dout(n23638),.clk(gclk));
	jor g23381(.dina(w_n23638_0[2]),.dinb(n23635),.dout(n23639),.clk(gclk));
	jand g23382(.dina(n23639),.dinb(w_n23634_0[1]),.dout(n23640),.clk(gclk));
	jor g23383(.dina(w_n23640_0[2]),.dinb(w_n3368_19[2]),.dout(n23641),.clk(gclk));
	jand g23384(.dina(w_n23640_0[1]),.dinb(w_n3368_19[1]),.dout(n23642),.clk(gclk));
	jxor g23385(.dina(w_n22889_0[0]),.dinb(w_n3642_21[2]),.dout(n23643),.clk(gclk));
	jor g23386(.dina(n23643),.dinb(w_n23345_19[0]),.dout(n23644),.clk(gclk));
	jxor g23387(.dina(n23644),.dinb(w_n23255_0[0]),.dout(n23645),.clk(gclk));
	jnot g23388(.din(w_n23645_0[2]),.dout(n23646),.clk(gclk));
	jor g23389(.dina(n23646),.dinb(n23642),.dout(n23647),.clk(gclk));
	jand g23390(.dina(n23647),.dinb(w_n23641_0[1]),.dout(n23648),.clk(gclk));
	jor g23391(.dina(w_n23648_0[2]),.dinb(w_n3089_23[0]),.dout(n23649),.clk(gclk));
	jand g23392(.dina(w_n23648_0[1]),.dinb(w_n3089_22[2]),.dout(n23650),.clk(gclk));
	jxor g23393(.dina(w_n22896_0[0]),.dinb(w_n3368_19[0]),.dout(n23651),.clk(gclk));
	jor g23394(.dina(n23651),.dinb(w_n23345_18[2]),.dout(n23652),.clk(gclk));
	jxor g23395(.dina(n23652),.dinb(w_n22902_0[0]),.dout(n23653),.clk(gclk));
	jor g23396(.dina(w_n23653_0[2]),.dinb(n23650),.dout(n23654),.clk(gclk));
	jand g23397(.dina(n23654),.dinb(w_n23649_0[1]),.dout(n23655),.clk(gclk));
	jor g23398(.dina(w_n23655_0[2]),.dinb(w_n2833_20[2]),.dout(n23656),.clk(gclk));
	jand g23399(.dina(w_n23655_0[1]),.dinb(w_n2833_20[1]),.dout(n23657),.clk(gclk));
	jxor g23400(.dina(w_n22904_0[0]),.dinb(w_n3089_22[1]),.dout(n23658),.clk(gclk));
	jor g23401(.dina(n23658),.dinb(w_n23345_18[1]),.dout(n23659),.clk(gclk));
	jxor g23402(.dina(n23659),.dinb(w_n23262_0[0]),.dout(n23660),.clk(gclk));
	jnot g23403(.din(w_n23660_0[2]),.dout(n23661),.clk(gclk));
	jor g23404(.dina(n23661),.dinb(n23657),.dout(n23662),.clk(gclk));
	jand g23405(.dina(n23662),.dinb(w_n23656_0[1]),.dout(n23663),.clk(gclk));
	jor g23406(.dina(w_n23663_0[2]),.dinb(w_n2572_23[1]),.dout(n23664),.clk(gclk));
	jand g23407(.dina(w_n23663_0[1]),.dinb(w_n2572_23[0]),.dout(n23665),.clk(gclk));
	jxor g23408(.dina(w_n22911_0[0]),.dinb(w_n2833_20[0]),.dout(n23666),.clk(gclk));
	jor g23409(.dina(n23666),.dinb(w_n23345_18[0]),.dout(n23667),.clk(gclk));
	jxor g23410(.dina(n23667),.dinb(w_n22917_0[0]),.dout(n23668),.clk(gclk));
	jor g23411(.dina(w_n23668_0[2]),.dinb(n23665),.dout(n23669),.clk(gclk));
	jand g23412(.dina(n23669),.dinb(w_n23664_0[1]),.dout(n23670),.clk(gclk));
	jor g23413(.dina(w_n23670_0[2]),.dinb(w_n2345_21[1]),.dout(n23671),.clk(gclk));
	jand g23414(.dina(w_n23670_0[1]),.dinb(w_n2345_21[0]),.dout(n23672),.clk(gclk));
	jxor g23415(.dina(w_n22919_0[0]),.dinb(w_n2572_22[2]),.dout(n23673),.clk(gclk));
	jor g23416(.dina(n23673),.dinb(w_n23345_17[2]),.dout(n23674),.clk(gclk));
	jxor g23417(.dina(n23674),.dinb(w_n22925_0[0]),.dout(n23675),.clk(gclk));
	jor g23418(.dina(w_n23675_0[2]),.dinb(n23672),.dout(n23676),.clk(gclk));
	jand g23419(.dina(n23676),.dinb(w_n23671_0[1]),.dout(n23677),.clk(gclk));
	jor g23420(.dina(w_n23677_0[2]),.dinb(w_n2108_24[0]),.dout(n23678),.clk(gclk));
	jand g23421(.dina(w_n23677_0[1]),.dinb(w_n2108_23[2]),.dout(n23679),.clk(gclk));
	jxor g23422(.dina(w_n22927_0[0]),.dinb(w_n2345_20[2]),.dout(n23680),.clk(gclk));
	jor g23423(.dina(n23680),.dinb(w_n23345_17[1]),.dout(n23681),.clk(gclk));
	jxor g23424(.dina(n23681),.dinb(w_n22933_0[0]),.dout(n23682),.clk(gclk));
	jor g23425(.dina(w_n23682_0[2]),.dinb(n23679),.dout(n23683),.clk(gclk));
	jand g23426(.dina(n23683),.dinb(w_n23678_0[1]),.dout(n23684),.clk(gclk));
	jor g23427(.dina(w_n23684_0[2]),.dinb(w_n1912_22[1]),.dout(n23685),.clk(gclk));
	jand g23428(.dina(w_n23684_0[1]),.dinb(w_n1912_22[0]),.dout(n23686),.clk(gclk));
	jxor g23429(.dina(w_n22935_0[0]),.dinb(w_n2108_23[1]),.dout(n23687),.clk(gclk));
	jor g23430(.dina(n23687),.dinb(w_n23345_17[0]),.dout(n23688),.clk(gclk));
	jxor g23431(.dina(n23688),.dinb(w_n23275_0[0]),.dout(n23689),.clk(gclk));
	jnot g23432(.din(w_n23689_0[2]),.dout(n23690),.clk(gclk));
	jor g23433(.dina(n23690),.dinb(n23686),.dout(n23691),.clk(gclk));
	jand g23434(.dina(n23691),.dinb(w_n23685_0[1]),.dout(n23692),.clk(gclk));
	jor g23435(.dina(w_n23692_0[2]),.dinb(w_n1699_24[2]),.dout(n23693),.clk(gclk));
	jand g23436(.dina(w_n23692_0[1]),.dinb(w_n1699_24[1]),.dout(n23694),.clk(gclk));
	jxor g23437(.dina(w_n22942_0[0]),.dinb(w_n1912_21[2]),.dout(n23695),.clk(gclk));
	jor g23438(.dina(n23695),.dinb(w_n23345_16[2]),.dout(n23696),.clk(gclk));
	jxor g23439(.dina(n23696),.dinb(w_n22948_0[0]),.dout(n23697),.clk(gclk));
	jor g23440(.dina(w_n23697_0[2]),.dinb(n23694),.dout(n23698),.clk(gclk));
	jand g23441(.dina(n23698),.dinb(w_n23693_0[1]),.dout(n23699),.clk(gclk));
	jor g23442(.dina(w_n23699_0[2]),.dinb(w_n1516_23[0]),.dout(n23700),.clk(gclk));
	jand g23443(.dina(w_n23699_0[1]),.dinb(w_n1516_22[2]),.dout(n23701),.clk(gclk));
	jxor g23444(.dina(w_n22950_0[0]),.dinb(w_n1699_24[0]),.dout(n23702),.clk(gclk));
	jor g23445(.dina(n23702),.dinb(w_n23345_16[1]),.dout(n23703),.clk(gclk));
	jxor g23446(.dina(n23703),.dinb(w_n22956_0[0]),.dout(n23704),.clk(gclk));
	jor g23447(.dina(w_n23704_0[2]),.dinb(n23701),.dout(n23705),.clk(gclk));
	jand g23448(.dina(n23705),.dinb(w_n23700_0[1]),.dout(n23706),.clk(gclk));
	jor g23449(.dina(w_n23706_0[2]),.dinb(w_n1332_24[2]),.dout(n23707),.clk(gclk));
	jand g23450(.dina(w_n23706_0[1]),.dinb(w_n1332_24[1]),.dout(n23708),.clk(gclk));
	jxor g23451(.dina(w_n22958_0[0]),.dinb(w_n1516_22[1]),.dout(n23709),.clk(gclk));
	jor g23452(.dina(n23709),.dinb(w_n23345_16[0]),.dout(n23710),.clk(gclk));
	jxor g23453(.dina(n23710),.dinb(w_n22964_0[0]),.dout(n23711),.clk(gclk));
	jor g23454(.dina(w_n23711_0[2]),.dinb(n23708),.dout(n23712),.clk(gclk));
	jand g23455(.dina(n23712),.dinb(w_n23707_0[1]),.dout(n23713),.clk(gclk));
	jor g23456(.dina(w_n23713_0[2]),.dinb(w_n1173_23[2]),.dout(n23714),.clk(gclk));
	jand g23457(.dina(w_n23713_0[1]),.dinb(w_n1173_23[1]),.dout(n23715),.clk(gclk));
	jxor g23458(.dina(w_n22966_0[0]),.dinb(w_n1332_24[0]),.dout(n23716),.clk(gclk));
	jor g23459(.dina(n23716),.dinb(w_n23345_15[2]),.dout(n23717),.clk(gclk));
	jxor g23460(.dina(n23717),.dinb(w_n22972_0[0]),.dout(n23718),.clk(gclk));
	jor g23461(.dina(w_n23718_0[2]),.dinb(n23715),.dout(n23719),.clk(gclk));
	jand g23462(.dina(n23719),.dinb(w_n23714_0[1]),.dout(n23720),.clk(gclk));
	jor g23463(.dina(w_n23720_0[2]),.dinb(w_n1008_25[2]),.dout(n23721),.clk(gclk));
	jand g23464(.dina(w_n23720_0[1]),.dinb(w_n1008_25[1]),.dout(n23722),.clk(gclk));
	jxor g23465(.dina(w_n22974_0[0]),.dinb(w_n1173_23[0]),.dout(n23723),.clk(gclk));
	jor g23466(.dina(n23723),.dinb(w_n23345_15[1]),.dout(n23724),.clk(gclk));
	jxor g23467(.dina(n23724),.dinb(w_n22980_0[0]),.dout(n23725),.clk(gclk));
	jor g23468(.dina(w_n23725_0[2]),.dinb(n23722),.dout(n23726),.clk(gclk));
	jand g23469(.dina(n23726),.dinb(w_n23721_0[1]),.dout(n23727),.clk(gclk));
	jor g23470(.dina(w_n23727_0[2]),.dinb(w_n884_24[2]),.dout(n23728),.clk(gclk));
	jand g23471(.dina(w_n23727_0[1]),.dinb(w_n884_24[1]),.dout(n23729),.clk(gclk));
	jxor g23472(.dina(w_n22982_0[0]),.dinb(w_n1008_25[0]),.dout(n23730),.clk(gclk));
	jor g23473(.dina(n23730),.dinb(w_n23345_15[0]),.dout(n23731),.clk(gclk));
	jxor g23474(.dina(n23731),.dinb(w_n23294_0[0]),.dout(n23732),.clk(gclk));
	jnot g23475(.din(w_n23732_0[2]),.dout(n23733),.clk(gclk));
	jor g23476(.dina(n23733),.dinb(n23729),.dout(n23734),.clk(gclk));
	jand g23477(.dina(n23734),.dinb(w_n23728_0[1]),.dout(n23735),.clk(gclk));
	jor g23478(.dina(w_n23735_0[2]),.dinb(w_n743_25[2]),.dout(n23736),.clk(gclk));
	jand g23479(.dina(w_n23735_0[1]),.dinb(w_n743_25[1]),.dout(n23737),.clk(gclk));
	jxor g23480(.dina(w_n22989_0[0]),.dinb(w_n884_24[0]),.dout(n23738),.clk(gclk));
	jor g23481(.dina(n23738),.dinb(w_n23345_14[2]),.dout(n23739),.clk(gclk));
	jxor g23482(.dina(n23739),.dinb(w_n22995_0[0]),.dout(n23740),.clk(gclk));
	jor g23483(.dina(w_n23740_0[2]),.dinb(n23737),.dout(n23741),.clk(gclk));
	jand g23484(.dina(n23741),.dinb(w_n23736_0[1]),.dout(n23742),.clk(gclk));
	jor g23485(.dina(w_n23742_0[2]),.dinb(w_n635_25[2]),.dout(n23743),.clk(gclk));
	jand g23486(.dina(w_n23742_0[1]),.dinb(w_n635_25[1]),.dout(n23744),.clk(gclk));
	jxor g23487(.dina(w_n22997_0[0]),.dinb(w_n743_25[0]),.dout(n23745),.clk(gclk));
	jor g23488(.dina(n23745),.dinb(w_n23345_14[1]),.dout(n23746),.clk(gclk));
	jxor g23489(.dina(n23746),.dinb(w_n23301_0[0]),.dout(n23747),.clk(gclk));
	jnot g23490(.din(w_n23747_0[2]),.dout(n23748),.clk(gclk));
	jor g23491(.dina(n23748),.dinb(n23744),.dout(n23749),.clk(gclk));
	jand g23492(.dina(n23749),.dinb(w_n23743_0[1]),.dout(n23750),.clk(gclk));
	jor g23493(.dina(w_n23750_0[2]),.dinb(w_n515_26[2]),.dout(n23751),.clk(gclk));
	jand g23494(.dina(w_n23750_0[1]),.dinb(w_n515_26[1]),.dout(n23752),.clk(gclk));
	jxor g23495(.dina(w_n23004_0[0]),.dinb(w_n635_25[0]),.dout(n23753),.clk(gclk));
	jor g23496(.dina(n23753),.dinb(w_n23345_14[0]),.dout(n23754),.clk(gclk));
	jxor g23497(.dina(n23754),.dinb(w_n23010_0[0]),.dout(n23755),.clk(gclk));
	jor g23498(.dina(w_n23755_0[2]),.dinb(n23752),.dout(n23756),.clk(gclk));
	jand g23499(.dina(n23756),.dinb(w_n23751_0[1]),.dout(n23757),.clk(gclk));
	jor g23500(.dina(w_n23757_0[2]),.dinb(w_n443_26[2]),.dout(n23758),.clk(gclk));
	jand g23501(.dina(w_n23757_0[1]),.dinb(w_n443_26[1]),.dout(n23759),.clk(gclk));
	jxor g23502(.dina(w_n23012_0[0]),.dinb(w_n515_26[0]),.dout(n23760),.clk(gclk));
	jor g23503(.dina(n23760),.dinb(w_n23345_13[2]),.dout(n23761),.clk(gclk));
	jxor g23504(.dina(n23761),.dinb(w_n23018_0[0]),.dout(n23762),.clk(gclk));
	jor g23505(.dina(w_n23762_0[1]),.dinb(n23759),.dout(n23763),.clk(gclk));
	jand g23506(.dina(n23763),.dinb(w_n23758_0[1]),.dout(n23764),.clk(gclk));
	jor g23507(.dina(w_n23764_0[2]),.dinb(w_n352_27[0]),.dout(n23765),.clk(gclk));
	jand g23508(.dina(w_n23764_0[1]),.dinb(w_n352_26[2]),.dout(n23766),.clk(gclk));
	jxor g23509(.dina(w_n23020_0[0]),.dinb(w_n443_26[0]),.dout(n23767),.clk(gclk));
	jor g23510(.dina(n23767),.dinb(w_n23345_13[1]),.dout(n23768),.clk(gclk));
	jxor g23511(.dina(n23768),.dinb(w_n23311_0[0]),.dout(n23769),.clk(gclk));
	jnot g23512(.din(w_n23769_0[2]),.dout(n23770),.clk(gclk));
	jor g23513(.dina(n23770),.dinb(n23766),.dout(n23771),.clk(gclk));
	jand g23514(.dina(n23771),.dinb(w_n23765_0[1]),.dout(n23772),.clk(gclk));
	jor g23515(.dina(w_n23772_0[2]),.dinb(w_n294_27[1]),.dout(n23773),.clk(gclk));
	jand g23516(.dina(w_n23772_0[1]),.dinb(w_n294_27[0]),.dout(n23774),.clk(gclk));
	jxor g23517(.dina(w_n23027_0[0]),.dinb(w_n352_26[1]),.dout(n23775),.clk(gclk));
	jor g23518(.dina(n23775),.dinb(w_n23345_13[0]),.dout(n23776),.clk(gclk));
	jxor g23519(.dina(n23776),.dinb(w_n23315_0[0]),.dout(n23777),.clk(gclk));
	jnot g23520(.din(w_n23777_0[2]),.dout(n23778),.clk(gclk));
	jor g23521(.dina(n23778),.dinb(n23774),.dout(n23779),.clk(gclk));
	jand g23522(.dina(n23779),.dinb(w_n23773_0[1]),.dout(n23780),.clk(gclk));
	jor g23523(.dina(w_n23780_0[2]),.dinb(w_n239_27[1]),.dout(n23781),.clk(gclk));
	jand g23524(.dina(w_n23780_0[1]),.dinb(w_n239_27[0]),.dout(n23782),.clk(gclk));
	jxor g23525(.dina(w_n23034_0[0]),.dinb(w_n294_26[2]),.dout(n23783),.clk(gclk));
	jor g23526(.dina(n23783),.dinb(w_n23345_12[2]),.dout(n23784),.clk(gclk));
	jxor g23527(.dina(n23784),.dinb(w_n23040_0[0]),.dout(n23785),.clk(gclk));
	jor g23528(.dina(w_n23785_0[2]),.dinb(n23782),.dout(n23786),.clk(gclk));
	jand g23529(.dina(n23786),.dinb(w_n23781_0[1]),.dout(n23787),.clk(gclk));
	jor g23530(.dina(w_n23787_0[2]),.dinb(w_n221_27[1]),.dout(n23788),.clk(gclk));
	jand g23531(.dina(w_n23787_0[1]),.dinb(w_n221_27[0]),.dout(n23789),.clk(gclk));
	jxor g23532(.dina(w_n23042_0[0]),.dinb(w_n239_26[2]),.dout(n23790),.clk(gclk));
	jor g23533(.dina(n23790),.dinb(w_n23345_12[1]),.dout(n23791),.clk(gclk));
	jxor g23534(.dina(n23791),.dinb(w_n23048_0[0]),.dout(n23792),.clk(gclk));
	jor g23535(.dina(w_n23792_0[2]),.dinb(n23789),.dout(n23793),.clk(gclk));
	jand g23536(.dina(n23793),.dinb(w_n23788_0[1]),.dout(n23794),.clk(gclk));
	jand g23537(.dina(w_n23794_1[1]),.dinb(w_n23349_0[2]),.dout(n23795),.clk(gclk));
	jand g23538(.dina(w_n23336_0[0]),.dinb(w_n23339_0[0]),.dout(n23796),.clk(gclk));
	jor g23539(.dina(w_n23794_1[0]),.dinb(w_n23349_0[1]),.dout(n23797),.clk(gclk));
	jor g23540(.dina(n23797),.dinb(w_n23064_0[0]),.dout(n23798),.clk(gclk));
	jor g23541(.dina(n23798),.dinb(w_n23796_0[1]),.dout(n23799),.clk(gclk));
	jand g23542(.dina(n23799),.dinb(w_n218_11[1]),.dout(n23800),.clk(gclk));
	jand g23543(.dina(w_n23344_0[0]),.dinb(w_n23326_0[0]),.dout(n23801),.clk(gclk));
	jnot g23544(.din(n23801),.dout(n23802),.clk(gclk));
	jand g23545(.dina(w_n23063_0[2]),.dinb(w_asqrt63_19[2]),.dout(n23803),.clk(gclk));
	jand g23546(.dina(n23803),.dinb(w_n23327_0[0]),.dout(n23804),.clk(gclk));
	jand g23547(.dina(n23804),.dinb(n23802),.dout(n23805),.clk(gclk));
	jor g23548(.dina(w_n23805_0[1]),.dinb(n23800),.dout(n23806),.clk(gclk));
	jor g23549(.dina(w_n23806_0[1]),.dinb(w_n23795_0[2]),.dout(asqrt_fa_3),.clk(gclk));
	jand g23550(.dina(w_asqrt2_31[1]),.dinb(w_a4_1[0]),.dout(n23808),.clk(gclk));
	jor g23551(.dina(w_a3_0[1]),.dinb(w_a2_1[1]),.dout(n23809),.clk(gclk));
	jnot g23552(.din(n23809),.dout(n23810),.clk(gclk));
	jand g23553(.dina(w_n23810_0[1]),.dinb(w_n23351_1[0]),.dout(n23811),.clk(gclk));
	jor g23554(.dina(w_n23811_0[1]),.dinb(n23808),.dout(n23812),.clk(gclk));
	jand g23555(.dina(w_n23812_0[2]),.dinb(w_asqrt3_1[2]),.dout(n23813),.clk(gclk));
	jor g23556(.dina(w_n23812_0[1]),.dinb(w_asqrt3_1[1]),.dout(n23814),.clk(gclk));
	jand g23557(.dina(w_asqrt2_31[0]),.dinb(w_n23351_0[2]),.dout(n23815),.clk(gclk));
	jor g23558(.dina(n23815),.dinb(w_n23352_0[0]),.dout(n23816),.clk(gclk));
	jnot g23559(.din(w_n23353_0[1]),.dout(n23817),.clk(gclk));
	jnot g23560(.din(w_n23795_0[1]),.dout(n23818),.clk(gclk));
	jnot g23561(.din(w_n23796_0[0]),.dout(n23819),.clk(gclk));
	jnot g23562(.din(w_n23788_0[0]),.dout(n23820),.clk(gclk));
	jnot g23563(.din(w_n23781_0[0]),.dout(n23821),.clk(gclk));
	jnot g23564(.din(w_n23773_0[0]),.dout(n23822),.clk(gclk));
	jnot g23565(.din(w_n23765_0[0]),.dout(n23823),.clk(gclk));
	jnot g23566(.din(w_n23758_0[0]),.dout(n23824),.clk(gclk));
	jnot g23567(.din(w_n23751_0[0]),.dout(n23825),.clk(gclk));
	jnot g23568(.din(w_n23743_0[0]),.dout(n23826),.clk(gclk));
	jnot g23569(.din(w_n23736_0[0]),.dout(n23827),.clk(gclk));
	jnot g23570(.din(w_n23728_0[0]),.dout(n23828),.clk(gclk));
	jnot g23571(.din(w_n23721_0[0]),.dout(n23829),.clk(gclk));
	jnot g23572(.din(w_n23714_0[0]),.dout(n23830),.clk(gclk));
	jnot g23573(.din(w_n23707_0[0]),.dout(n23831),.clk(gclk));
	jnot g23574(.din(w_n23700_0[0]),.dout(n23832),.clk(gclk));
	jnot g23575(.din(w_n23693_0[0]),.dout(n23833),.clk(gclk));
	jnot g23576(.din(w_n23685_0[0]),.dout(n23834),.clk(gclk));
	jnot g23577(.din(w_n23678_0[0]),.dout(n23835),.clk(gclk));
	jnot g23578(.din(w_n23671_0[0]),.dout(n23836),.clk(gclk));
	jnot g23579(.din(w_n23664_0[0]),.dout(n23837),.clk(gclk));
	jnot g23580(.din(w_n23656_0[0]),.dout(n23838),.clk(gclk));
	jnot g23581(.din(w_n23649_0[0]),.dout(n23839),.clk(gclk));
	jnot g23582(.din(w_n23641_0[0]),.dout(n23840),.clk(gclk));
	jnot g23583(.din(w_n23634_0[0]),.dout(n23841),.clk(gclk));
	jnot g23584(.din(w_n23626_0[0]),.dout(n23842),.clk(gclk));
	jnot g23585(.din(w_n23619_0[0]),.dout(n23843),.clk(gclk));
	jnot g23586(.din(w_n23611_0[0]),.dout(n23844),.clk(gclk));
	jnot g23587(.din(w_n23604_0[0]),.dout(n23845),.clk(gclk));
	jnot g23588(.din(w_n23597_0[0]),.dout(n23846),.clk(gclk));
	jnot g23589(.din(w_n23590_0[0]),.dout(n23847),.clk(gclk));
	jnot g23590(.din(w_n23582_0[0]),.dout(n23848),.clk(gclk));
	jnot g23591(.din(w_n23575_0[0]),.dout(n23849),.clk(gclk));
	jnot g23592(.din(w_n23567_0[0]),.dout(n23850),.clk(gclk));
	jnot g23593(.din(w_n23560_0[0]),.dout(n23851),.clk(gclk));
	jnot g23594(.din(w_n23552_0[0]),.dout(n23852),.clk(gclk));
	jnot g23595(.din(w_n23544_0[0]),.dout(n23853),.clk(gclk));
	jnot g23596(.din(w_n23537_0[0]),.dout(n23854),.clk(gclk));
	jnot g23597(.din(w_n23530_0[0]),.dout(n23855),.clk(gclk));
	jnot g23598(.din(w_n23522_0[0]),.dout(n23856),.clk(gclk));
	jnot g23599(.din(w_n23515_0[0]),.dout(n23857),.clk(gclk));
	jnot g23600(.din(w_n23507_0[0]),.dout(n23858),.clk(gclk));
	jnot g23601(.din(w_n23500_0[0]),.dout(n23859),.clk(gclk));
	jnot g23602(.din(w_n23492_0[0]),.dout(n23860),.clk(gclk));
	jnot g23603(.din(w_n23485_0[0]),.dout(n23861),.clk(gclk));
	jnot g23604(.din(w_n23478_0[0]),.dout(n23862),.clk(gclk));
	jnot g23605(.din(w_n23471_0[0]),.dout(n23863),.clk(gclk));
	jnot g23606(.din(w_n23463_0[0]),.dout(n23864),.clk(gclk));
	jnot g23607(.din(w_n23456_0[0]),.dout(n23865),.clk(gclk));
	jnot g23608(.din(w_n23449_0[0]),.dout(n23866),.clk(gclk));
	jnot g23609(.din(w_n23442_0[0]),.dout(n23867),.clk(gclk));
	jnot g23610(.din(w_n23434_0[0]),.dout(n23868),.clk(gclk));
	jnot g23611(.din(w_n23427_0[0]),.dout(n23869),.clk(gclk));
	jnot g23612(.din(w_n23419_0[0]),.dout(n23870),.clk(gclk));
	jnot g23613(.din(w_n23412_0[0]),.dout(n23871),.clk(gclk));
	jnot g23614(.din(w_n23404_0[0]),.dout(n23872),.clk(gclk));
	jnot g23615(.din(w_n23396_0[0]),.dout(n23873),.clk(gclk));
	jnot g23616(.din(w_n23388_0[0]),.dout(n23874),.clk(gclk));
	jnot g23617(.din(w_n23381_0[0]),.dout(n23875),.clk(gclk));
	jnot g23618(.din(w_n23374_0[0]),.dout(n23876),.clk(gclk));
	jnot g23619(.din(w_n23365_0[0]),.dout(n23877),.clk(gclk));
	jnot g23620(.din(w_n23357_0[0]),.dout(n23878),.clk(gclk));
	jand g23621(.dina(w_asqrt3_1[0]),.dinb(w_a6_0[0]),.dout(n23879),.clk(gclk));
	jor g23622(.dina(w_n23354_0[0]),.dinb(n23879),.dout(n23880),.clk(gclk));
	jor g23623(.dina(n23880),.dinb(w_asqrt4_11[0]),.dout(n23881),.clk(gclk));
	jand g23624(.dina(w_asqrt3_0[2]),.dinb(w_n22334_0[2]),.dout(n23882),.clk(gclk));
	jor g23625(.dina(n23882),.dinb(w_n22335_0[0]),.dout(n23883),.clk(gclk));
	jand g23626(.dina(w_n23368_0[0]),.dinb(n23883),.dout(n23884),.clk(gclk));
	jand g23627(.dina(w_n23884_0[1]),.dinb(n23881),.dout(n23885),.clk(gclk));
	jor g23628(.dina(n23885),.dinb(n23878),.dout(n23886),.clk(gclk));
	jor g23629(.dina(n23886),.dinb(w_asqrt5_2[0]),.dout(n23887),.clk(gclk));
	jnot g23630(.din(w_n23371_0[0]),.dout(n23888),.clk(gclk));
	jand g23631(.dina(w_n23888_0[1]),.dinb(n23887),.dout(n23889),.clk(gclk));
	jor g23632(.dina(n23889),.dinb(n23877),.dout(n23890),.clk(gclk));
	jor g23633(.dina(n23890),.dinb(w_asqrt6_11[1]),.dout(n23891),.clk(gclk));
	jnot g23634(.din(w_n23378_0[1]),.dout(n23892),.clk(gclk));
	jand g23635(.dina(n23892),.dinb(n23891),.dout(n23893),.clk(gclk));
	jor g23636(.dina(n23893),.dinb(n23876),.dout(n23894),.clk(gclk));
	jor g23637(.dina(n23894),.dinb(w_asqrt7_2[2]),.dout(n23895),.clk(gclk));
	jnot g23638(.din(w_n23385_0[1]),.dout(n23896),.clk(gclk));
	jand g23639(.dina(n23896),.dinb(n23895),.dout(n23897),.clk(gclk));
	jor g23640(.dina(n23897),.dinb(n23875),.dout(n23898),.clk(gclk));
	jor g23641(.dina(n23898),.dinb(w_asqrt8_11[1]),.dout(n23899),.clk(gclk));
	jand g23642(.dina(w_n23392_0[1]),.dinb(n23899),.dout(n23900),.clk(gclk));
	jor g23643(.dina(n23900),.dinb(n23874),.dout(n23901),.clk(gclk));
	jor g23644(.dina(n23901),.dinb(w_asqrt9_3[1]),.dout(n23902),.clk(gclk));
	jand g23645(.dina(w_n23400_0[1]),.dinb(n23902),.dout(n23903),.clk(gclk));
	jor g23646(.dina(n23903),.dinb(n23873),.dout(n23904),.clk(gclk));
	jor g23647(.dina(n23904),.dinb(w_asqrt10_11[1]),.dout(n23905),.clk(gclk));
	jand g23648(.dina(w_n23408_0[1]),.dinb(n23905),.dout(n23906),.clk(gclk));
	jor g23649(.dina(n23906),.dinb(n23872),.dout(n23907),.clk(gclk));
	jor g23650(.dina(n23907),.dinb(w_asqrt11_3[1]),.dout(n23908),.clk(gclk));
	jnot g23651(.din(w_n23416_0[1]),.dout(n23909),.clk(gclk));
	jand g23652(.dina(n23909),.dinb(n23908),.dout(n23910),.clk(gclk));
	jor g23653(.dina(n23910),.dinb(n23871),.dout(n23911),.clk(gclk));
	jor g23654(.dina(n23911),.dinb(w_asqrt12_11[2]),.dout(n23912),.clk(gclk));
	jand g23655(.dina(w_n23423_0[1]),.dinb(n23912),.dout(n23913),.clk(gclk));
	jor g23656(.dina(n23913),.dinb(n23870),.dout(n23914),.clk(gclk));
	jor g23657(.dina(n23914),.dinb(w_asqrt13_4[0]),.dout(n23915),.clk(gclk));
	jnot g23658(.din(w_n23431_0[1]),.dout(n23916),.clk(gclk));
	jand g23659(.dina(n23916),.dinb(n23915),.dout(n23917),.clk(gclk));
	jor g23660(.dina(n23917),.dinb(n23869),.dout(n23918),.clk(gclk));
	jor g23661(.dina(n23918),.dinb(w_asqrt14_12[0]),.dout(n23919),.clk(gclk));
	jand g23662(.dina(w_n23438_0[1]),.dinb(n23919),.dout(n23920),.clk(gclk));
	jor g23663(.dina(n23920),.dinb(n23868),.dout(n23921),.clk(gclk));
	jor g23664(.dina(n23921),.dinb(w_asqrt15_4[2]),.dout(n23922),.clk(gclk));
	jnot g23665(.din(w_n23446_0[1]),.dout(n23923),.clk(gclk));
	jand g23666(.dina(n23923),.dinb(n23922),.dout(n23924),.clk(gclk));
	jor g23667(.dina(n23924),.dinb(n23867),.dout(n23925),.clk(gclk));
	jor g23668(.dina(n23925),.dinb(w_asqrt16_12[0]),.dout(n23926),.clk(gclk));
	jnot g23669(.din(w_n23453_0[1]),.dout(n23927),.clk(gclk));
	jand g23670(.dina(n23927),.dinb(n23926),.dout(n23928),.clk(gclk));
	jor g23671(.dina(n23928),.dinb(n23866),.dout(n23929),.clk(gclk));
	jor g23672(.dina(n23929),.dinb(w_asqrt17_5[0]),.dout(n23930),.clk(gclk));
	jnot g23673(.din(w_n23460_0[1]),.dout(n23931),.clk(gclk));
	jand g23674(.dina(n23931),.dinb(n23930),.dout(n23932),.clk(gclk));
	jor g23675(.dina(n23932),.dinb(n23865),.dout(n23933),.clk(gclk));
	jor g23676(.dina(n23933),.dinb(w_asqrt18_12[1]),.dout(n23934),.clk(gclk));
	jand g23677(.dina(w_n23467_0[1]),.dinb(n23934),.dout(n23935),.clk(gclk));
	jor g23678(.dina(n23935),.dinb(n23864),.dout(n23936),.clk(gclk));
	jor g23679(.dina(n23936),.dinb(w_asqrt19_5[1]),.dout(n23937),.clk(gclk));
	jnot g23680(.din(w_n23475_0[1]),.dout(n23938),.clk(gclk));
	jand g23681(.dina(n23938),.dinb(n23937),.dout(n23939),.clk(gclk));
	jor g23682(.dina(n23939),.dinb(n23863),.dout(n23940),.clk(gclk));
	jor g23683(.dina(n23940),.dinb(w_asqrt20_12[1]),.dout(n23941),.clk(gclk));
	jnot g23684(.din(w_n23482_0[1]),.dout(n23942),.clk(gclk));
	jand g23685(.dina(n23942),.dinb(n23941),.dout(n23943),.clk(gclk));
	jor g23686(.dina(n23943),.dinb(n23862),.dout(n23944),.clk(gclk));
	jor g23687(.dina(n23944),.dinb(w_asqrt21_6[0]),.dout(n23945),.clk(gclk));
	jnot g23688(.din(w_n23489_0[1]),.dout(n23946),.clk(gclk));
	jand g23689(.dina(n23946),.dinb(n23945),.dout(n23947),.clk(gclk));
	jor g23690(.dina(n23947),.dinb(n23861),.dout(n23948),.clk(gclk));
	jor g23691(.dina(n23948),.dinb(w_asqrt22_12[2]),.dout(n23949),.clk(gclk));
	jand g23692(.dina(w_n23496_0[1]),.dinb(n23949),.dout(n23950),.clk(gclk));
	jor g23693(.dina(n23950),.dinb(n23860),.dout(n23951),.clk(gclk));
	jor g23694(.dina(n23951),.dinb(w_asqrt23_6[2]),.dout(n23952),.clk(gclk));
	jnot g23695(.din(w_n23504_0[1]),.dout(n23953),.clk(gclk));
	jand g23696(.dina(n23953),.dinb(n23952),.dout(n23954),.clk(gclk));
	jor g23697(.dina(n23954),.dinb(n23859),.dout(n23955),.clk(gclk));
	jor g23698(.dina(n23955),.dinb(w_asqrt24_12[2]),.dout(n23956),.clk(gclk));
	jand g23699(.dina(w_n23511_0[1]),.dinb(n23956),.dout(n23957),.clk(gclk));
	jor g23700(.dina(n23957),.dinb(n23858),.dout(n23958),.clk(gclk));
	jor g23701(.dina(n23958),.dinb(w_asqrt25_6[2]),.dout(n23959),.clk(gclk));
	jnot g23702(.din(w_n23519_0[1]),.dout(n23960),.clk(gclk));
	jand g23703(.dina(n23960),.dinb(n23959),.dout(n23961),.clk(gclk));
	jor g23704(.dina(n23961),.dinb(n23857),.dout(n23962),.clk(gclk));
	jor g23705(.dina(n23962),.dinb(w_asqrt26_12[2]),.dout(n23963),.clk(gclk));
	jand g23706(.dina(w_n23526_0[1]),.dinb(n23963),.dout(n23964),.clk(gclk));
	jor g23707(.dina(n23964),.dinb(n23856),.dout(n23965),.clk(gclk));
	jor g23708(.dina(n23965),.dinb(w_asqrt27_7[1]),.dout(n23966),.clk(gclk));
	jnot g23709(.din(w_n23534_0[1]),.dout(n23967),.clk(gclk));
	jand g23710(.dina(n23967),.dinb(n23966),.dout(n23968),.clk(gclk));
	jor g23711(.dina(n23968),.dinb(n23855),.dout(n23969),.clk(gclk));
	jor g23712(.dina(n23969),.dinb(w_asqrt28_13[0]),.dout(n23970),.clk(gclk));
	jnot g23713(.din(w_n23541_0[1]),.dout(n23971),.clk(gclk));
	jand g23714(.dina(n23971),.dinb(n23970),.dout(n23972),.clk(gclk));
	jor g23715(.dina(n23972),.dinb(n23854),.dout(n23973),.clk(gclk));
	jor g23716(.dina(n23973),.dinb(w_asqrt29_7[2]),.dout(n23974),.clk(gclk));
	jand g23717(.dina(w_n23548_0[1]),.dinb(n23974),.dout(n23975),.clk(gclk));
	jor g23718(.dina(n23975),.dinb(n23853),.dout(n23976),.clk(gclk));
	jor g23719(.dina(n23976),.dinb(w_asqrt30_13[1]),.dout(n23977),.clk(gclk));
	jand g23720(.dina(w_n23556_0[1]),.dinb(n23977),.dout(n23978),.clk(gclk));
	jor g23721(.dina(n23978),.dinb(n23852),.dout(n23979),.clk(gclk));
	jor g23722(.dina(n23979),.dinb(w_asqrt31_8[1]),.dout(n23980),.clk(gclk));
	jnot g23723(.din(w_n23564_0[1]),.dout(n23981),.clk(gclk));
	jand g23724(.dina(n23981),.dinb(n23980),.dout(n23982),.clk(gclk));
	jor g23725(.dina(n23982),.dinb(n23851),.dout(n23983),.clk(gclk));
	jor g23726(.dina(n23983),.dinb(w_asqrt32_13[1]),.dout(n23984),.clk(gclk));
	jand g23727(.dina(w_n23571_0[1]),.dinb(n23984),.dout(n23985),.clk(gclk));
	jor g23728(.dina(n23985),.dinb(n23850),.dout(n23986),.clk(gclk));
	jor g23729(.dina(n23986),.dinb(w_asqrt33_9[0]),.dout(n23987),.clk(gclk));
	jnot g23730(.din(w_n23579_0[1]),.dout(n23988),.clk(gclk));
	jand g23731(.dina(n23988),.dinb(n23987),.dout(n23989),.clk(gclk));
	jor g23732(.dina(n23989),.dinb(n23849),.dout(n23990),.clk(gclk));
	jor g23733(.dina(n23990),.dinb(w_asqrt34_13[2]),.dout(n23991),.clk(gclk));
	jand g23734(.dina(w_n23586_0[1]),.dinb(n23991),.dout(n23992),.clk(gclk));
	jor g23735(.dina(n23992),.dinb(n23848),.dout(n23993),.clk(gclk));
	jor g23736(.dina(n23993),.dinb(w_asqrt35_9[2]),.dout(n23994),.clk(gclk));
	jnot g23737(.din(w_n23594_0[1]),.dout(n23995),.clk(gclk));
	jand g23738(.dina(n23995),.dinb(n23994),.dout(n23996),.clk(gclk));
	jor g23739(.dina(n23996),.dinb(n23847),.dout(n23997),.clk(gclk));
	jor g23740(.dina(n23997),.dinb(w_asqrt36_13[2]),.dout(n23998),.clk(gclk));
	jnot g23741(.din(w_n23601_0[1]),.dout(n23999),.clk(gclk));
	jand g23742(.dina(n23999),.dinb(n23998),.dout(n24000),.clk(gclk));
	jor g23743(.dina(n24000),.dinb(n23846),.dout(n24001),.clk(gclk));
	jor g23744(.dina(n24001),.dinb(w_asqrt37_10[0]),.dout(n24002),.clk(gclk));
	jnot g23745(.din(w_n23608_0[1]),.dout(n24003),.clk(gclk));
	jand g23746(.dina(n24003),.dinb(n24002),.dout(n24004),.clk(gclk));
	jor g23747(.dina(n24004),.dinb(n23845),.dout(n24005),.clk(gclk));
	jor g23748(.dina(n24005),.dinb(w_asqrt38_14[0]),.dout(n24006),.clk(gclk));
	jand g23749(.dina(w_n23615_0[1]),.dinb(n24006),.dout(n24007),.clk(gclk));
	jor g23750(.dina(n24007),.dinb(n23844),.dout(n24008),.clk(gclk));
	jor g23751(.dina(n24008),.dinb(w_asqrt39_10[2]),.dout(n24009),.clk(gclk));
	jnot g23752(.din(w_n23623_0[1]),.dout(n24010),.clk(gclk));
	jand g23753(.dina(n24010),.dinb(n24009),.dout(n24011),.clk(gclk));
	jor g23754(.dina(n24011),.dinb(n23843),.dout(n24012),.clk(gclk));
	jor g23755(.dina(n24012),.dinb(w_asqrt40_14[0]),.dout(n24013),.clk(gclk));
	jand g23756(.dina(w_n23630_0[1]),.dinb(n24013),.dout(n24014),.clk(gclk));
	jor g23757(.dina(n24014),.dinb(n23842),.dout(n24015),.clk(gclk));
	jor g23758(.dina(n24015),.dinb(w_asqrt41_11[0]),.dout(n24016),.clk(gclk));
	jnot g23759(.din(w_n23638_0[1]),.dout(n24017),.clk(gclk));
	jand g23760(.dina(n24017),.dinb(n24016),.dout(n24018),.clk(gclk));
	jor g23761(.dina(n24018),.dinb(n23841),.dout(n24019),.clk(gclk));
	jor g23762(.dina(n24019),.dinb(w_asqrt42_14[1]),.dout(n24020),.clk(gclk));
	jand g23763(.dina(w_n23645_0[1]),.dinb(n24020),.dout(n24021),.clk(gclk));
	jor g23764(.dina(n24021),.dinb(n23840),.dout(n24022),.clk(gclk));
	jor g23765(.dina(n24022),.dinb(w_asqrt43_11[1]),.dout(n24023),.clk(gclk));
	jnot g23766(.din(w_n23653_0[1]),.dout(n24024),.clk(gclk));
	jand g23767(.dina(n24024),.dinb(n24023),.dout(n24025),.clk(gclk));
	jor g23768(.dina(n24025),.dinb(n23839),.dout(n24026),.clk(gclk));
	jor g23769(.dina(n24026),.dinb(w_asqrt44_14[1]),.dout(n24027),.clk(gclk));
	jand g23770(.dina(w_n23660_0[1]),.dinb(n24027),.dout(n24028),.clk(gclk));
	jor g23771(.dina(n24028),.dinb(n23838),.dout(n24029),.clk(gclk));
	jor g23772(.dina(n24029),.dinb(w_asqrt45_12[0]),.dout(n24030),.clk(gclk));
	jnot g23773(.din(w_n23668_0[1]),.dout(n24031),.clk(gclk));
	jand g23774(.dina(n24031),.dinb(n24030),.dout(n24032),.clk(gclk));
	jor g23775(.dina(n24032),.dinb(n23837),.dout(n24033),.clk(gclk));
	jor g23776(.dina(n24033),.dinb(w_asqrt46_14[1]),.dout(n24034),.clk(gclk));
	jnot g23777(.din(w_n23675_0[1]),.dout(n24035),.clk(gclk));
	jand g23778(.dina(n24035),.dinb(n24034),.dout(n24036),.clk(gclk));
	jor g23779(.dina(n24036),.dinb(n23836),.dout(n24037),.clk(gclk));
	jor g23780(.dina(n24037),.dinb(w_asqrt47_12[2]),.dout(n24038),.clk(gclk));
	jnot g23781(.din(w_n23682_0[1]),.dout(n24039),.clk(gclk));
	jand g23782(.dina(n24039),.dinb(n24038),.dout(n24040),.clk(gclk));
	jor g23783(.dina(n24040),.dinb(n23835),.dout(n24041),.clk(gclk));
	jor g23784(.dina(n24041),.dinb(w_asqrt48_14[2]),.dout(n24042),.clk(gclk));
	jand g23785(.dina(w_n23689_0[1]),.dinb(n24042),.dout(n24043),.clk(gclk));
	jor g23786(.dina(n24043),.dinb(n23834),.dout(n24044),.clk(gclk));
	jor g23787(.dina(n24044),.dinb(w_asqrt49_13[0]),.dout(n24045),.clk(gclk));
	jnot g23788(.din(w_n23697_0[1]),.dout(n24046),.clk(gclk));
	jand g23789(.dina(n24046),.dinb(n24045),.dout(n24047),.clk(gclk));
	jor g23790(.dina(n24047),.dinb(n23833),.dout(n24048),.clk(gclk));
	jor g23791(.dina(n24048),.dinb(w_asqrt50_15[0]),.dout(n24049),.clk(gclk));
	jnot g23792(.din(w_n23704_0[1]),.dout(n24050),.clk(gclk));
	jand g23793(.dina(n24050),.dinb(n24049),.dout(n24051),.clk(gclk));
	jor g23794(.dina(n24051),.dinb(n23832),.dout(n24052),.clk(gclk));
	jor g23795(.dina(n24052),.dinb(w_asqrt51_13[1]),.dout(n24053),.clk(gclk));
	jnot g23796(.din(w_n23711_0[1]),.dout(n24054),.clk(gclk));
	jand g23797(.dina(n24054),.dinb(n24053),.dout(n24055),.clk(gclk));
	jor g23798(.dina(n24055),.dinb(n23831),.dout(n24056),.clk(gclk));
	jor g23799(.dina(n24056),.dinb(w_asqrt52_15[0]),.dout(n24057),.clk(gclk));
	jnot g23800(.din(w_n23718_0[1]),.dout(n24058),.clk(gclk));
	jand g23801(.dina(n24058),.dinb(n24057),.dout(n24059),.clk(gclk));
	jor g23802(.dina(n24059),.dinb(n23830),.dout(n24060),.clk(gclk));
	jor g23803(.dina(n24060),.dinb(w_asqrt53_14[0]),.dout(n24061),.clk(gclk));
	jnot g23804(.din(w_n23725_0[1]),.dout(n24062),.clk(gclk));
	jand g23805(.dina(n24062),.dinb(n24061),.dout(n24063),.clk(gclk));
	jor g23806(.dina(n24063),.dinb(n23829),.dout(n24064),.clk(gclk));
	jor g23807(.dina(n24064),.dinb(w_asqrt54_15[0]),.dout(n24065),.clk(gclk));
	jand g23808(.dina(w_n23732_0[1]),.dinb(n24065),.dout(n24066),.clk(gclk));
	jor g23809(.dina(n24066),.dinb(n23828),.dout(n24067),.clk(gclk));
	jor g23810(.dina(n24067),.dinb(w_asqrt55_14[1]),.dout(n24068),.clk(gclk));
	jnot g23811(.din(w_n23740_0[1]),.dout(n24069),.clk(gclk));
	jand g23812(.dina(n24069),.dinb(n24068),.dout(n24070),.clk(gclk));
	jor g23813(.dina(n24070),.dinb(n23827),.dout(n24071),.clk(gclk));
	jor g23814(.dina(n24071),.dinb(w_asqrt56_15[1]),.dout(n24072),.clk(gclk));
	jand g23815(.dina(w_n23747_0[1]),.dinb(n24072),.dout(n24073),.clk(gclk));
	jor g23816(.dina(n24073),.dinb(n23826),.dout(n24074),.clk(gclk));
	jor g23817(.dina(n24074),.dinb(w_asqrt57_15[0]),.dout(n24075),.clk(gclk));
	jnot g23818(.din(w_n23755_0[1]),.dout(n24076),.clk(gclk));
	jand g23819(.dina(n24076),.dinb(n24075),.dout(n24077),.clk(gclk));
	jor g23820(.dina(n24077),.dinb(n23825),.dout(n24078),.clk(gclk));
	jor g23821(.dina(n24078),.dinb(w_asqrt58_15[2]),.dout(n24079),.clk(gclk));
	jnot g23822(.din(w_n23762_0[0]),.dout(n24080),.clk(gclk));
	jand g23823(.dina(w_n24080_0[1]),.dinb(n24079),.dout(n24081),.clk(gclk));
	jor g23824(.dina(n24081),.dinb(n23824),.dout(n24082),.clk(gclk));
	jor g23825(.dina(n24082),.dinb(w_asqrt59_15[1]),.dout(n24083),.clk(gclk));
	jand g23826(.dina(w_n23769_0[1]),.dinb(n24083),.dout(n24084),.clk(gclk));
	jor g23827(.dina(n24084),.dinb(n23823),.dout(n24085),.clk(gclk));
	jor g23828(.dina(n24085),.dinb(w_asqrt60_15[2]),.dout(n24086),.clk(gclk));
	jand g23829(.dina(w_n23777_0[1]),.dinb(n24086),.dout(n24087),.clk(gclk));
	jor g23830(.dina(n24087),.dinb(n23822),.dout(n24088),.clk(gclk));
	jor g23831(.dina(n24088),.dinb(w_asqrt61_15[2]),.dout(n24089),.clk(gclk));
	jnot g23832(.din(w_n23785_0[1]),.dout(n24090),.clk(gclk));
	jand g23833(.dina(n24090),.dinb(n24089),.dout(n24091),.clk(gclk));
	jor g23834(.dina(n24091),.dinb(n23821),.dout(n24092),.clk(gclk));
	jor g23835(.dina(n24092),.dinb(w_asqrt62_15[2]),.dout(n24093),.clk(gclk));
	jnot g23836(.din(w_n23792_0[1]),.dout(n24094),.clk(gclk));
	jand g23837(.dina(n24094),.dinb(n24093),.dout(n24095),.clk(gclk));
	jor g23838(.dina(n24095),.dinb(n23820),.dout(n24096),.clk(gclk));
	jand g23839(.dina(n24096),.dinb(w_n23348_0[0]),.dout(n24097),.clk(gclk));
	jand g23840(.dina(w_n24097_0[1]),.dinb(w_n23063_0[1]),.dout(n24098),.clk(gclk));
	jand g23841(.dina(n24098),.dinb(n23819),.dout(n24099),.clk(gclk));
	jor g23842(.dina(n24099),.dinb(w_asqrt63_19[1]),.dout(n24100),.clk(gclk));
	jnot g23843(.din(w_n23805_0[0]),.dout(n24101),.clk(gclk));
	jand g23844(.dina(n24101),.dinb(n24100),.dout(n24102),.clk(gclk));
	jand g23845(.dina(w_n24102_0[1]),.dinb(w_n23818_0[1]),.dout(n24103),.clk(gclk));
	jor g23846(.dina(w_n24103_1[2]),.dinb(n23817),.dout(n24104),.clk(gclk));
	jand g23847(.dina(w_n24104_0[1]),.dinb(n23816),.dout(n24105),.clk(gclk));
	jand g23848(.dina(w_n24105_0[1]),.dinb(n23814),.dout(n24106),.clk(gclk));
	jor g23849(.dina(n24106),.dinb(w_n23813_0[1]),.dout(n24107),.clk(gclk));
	jand g23850(.dina(w_n24107_0[2]),.dinb(w_asqrt4_10[2]),.dout(n24108),.clk(gclk));
	jor g23851(.dina(w_n24107_0[1]),.dinb(w_asqrt4_10[1]),.dout(n24109),.clk(gclk));
	jor g23852(.dina(w_asqrt2_30[2]),.dinb(w_n23345_12[0]),.dout(n24110),.clk(gclk));
	jand g23853(.dina(n24110),.dinb(w_n24104_0[0]),.dout(n24111),.clk(gclk));
	jxor g23854(.dina(n24111),.dinb(w_n22334_0[1]),.dout(n24112),.clk(gclk));
	jnot g23855(.din(w_n24112_0[1]),.dout(n24113),.clk(gclk));
	jand g23856(.dina(w_n24113_0[1]),.dinb(n24109),.dout(n24114),.clk(gclk));
	jor g23857(.dina(n24114),.dinb(w_n24108_0[1]),.dout(n24115),.clk(gclk));
	jand g23858(.dina(w_n24115_0[2]),.dinb(w_asqrt5_1[2]),.dout(n24116),.clk(gclk));
	jor g23859(.dina(w_n24115_0[1]),.dinb(w_asqrt5_1[1]),.dout(n24117),.clk(gclk));
	jxor g23860(.dina(w_n23356_0[0]),.dinb(w_n22620_2[2]),.dout(n24118),.clk(gclk));
	jand g23861(.dina(n24118),.dinb(w_asqrt2_30[1]),.dout(n24119),.clk(gclk));
	jxor g23862(.dina(n24119),.dinb(w_n23884_0[0]),.dout(n24120),.clk(gclk));
	jand g23863(.dina(w_n24120_0[2]),.dinb(n24117),.dout(n24121),.clk(gclk));
	jor g23864(.dina(n24121),.dinb(w_n24116_0[1]),.dout(n24122),.clk(gclk));
	jand g23865(.dina(w_n24122_0[2]),.dinb(w_asqrt6_11[0]),.dout(n24123),.clk(gclk));
	jor g23866(.dina(w_n24122_0[1]),.dinb(w_asqrt6_10[2]),.dout(n24124),.clk(gclk));
	jxor g23867(.dina(w_n23364_0[0]),.dinb(w_n21887_12[2]),.dout(n24125),.clk(gclk));
	jand g23868(.dina(n24125),.dinb(w_asqrt2_30[0]),.dout(n24126),.clk(gclk));
	jxor g23869(.dina(n24126),.dinb(w_n23888_0[0]),.dout(n24127),.clk(gclk));
	jand g23870(.dina(w_n24127_0[2]),.dinb(n24124),.dout(n24128),.clk(gclk));
	jor g23871(.dina(n24128),.dinb(w_n24123_0[1]),.dout(n24129),.clk(gclk));
	jand g23872(.dina(w_n24129_0[2]),.dinb(w_asqrt7_2[1]),.dout(n24130),.clk(gclk));
	jor g23873(.dina(w_n24129_0[1]),.dinb(w_asqrt7_2[0]),.dout(n24131),.clk(gclk));
	jxor g23874(.dina(w_n23373_0[0]),.dinb(w_n21184_3[2]),.dout(n24132),.clk(gclk));
	jand g23875(.dina(n24132),.dinb(w_asqrt2_29[2]),.dout(n24133),.clk(gclk));
	jxor g23876(.dina(n24133),.dinb(w_n23378_0[0]),.dout(n24134),.clk(gclk));
	jnot g23877(.din(w_n24134_0[1]),.dout(n24135),.clk(gclk));
	jand g23878(.dina(w_n24135_0[1]),.dinb(n24131),.dout(n24136),.clk(gclk));
	jor g23879(.dina(n24136),.dinb(w_n24130_0[1]),.dout(n24137),.clk(gclk));
	jand g23880(.dina(w_n24137_0[2]),.dinb(w_asqrt8_11[0]),.dout(n24138),.clk(gclk));
	jor g23881(.dina(w_n24137_0[1]),.dinb(w_asqrt8_10[2]),.dout(n24139),.clk(gclk));
	jxor g23882(.dina(w_n23380_0[0]),.dinb(w_n20468_13[0]),.dout(n24140),.clk(gclk));
	jand g23883(.dina(n24140),.dinb(w_asqrt2_29[1]),.dout(n24141),.clk(gclk));
	jxor g23884(.dina(n24141),.dinb(w_n23385_0[0]),.dout(n24142),.clk(gclk));
	jnot g23885(.din(w_n24142_0[1]),.dout(n24143),.clk(gclk));
	jand g23886(.dina(w_n24143_0[1]),.dinb(n24139),.dout(n24144),.clk(gclk));
	jor g23887(.dina(n24144),.dinb(w_n24138_0[1]),.dout(n24145),.clk(gclk));
	jand g23888(.dina(w_n24145_0[2]),.dinb(w_asqrt9_3[0]),.dout(n24146),.clk(gclk));
	jor g23889(.dina(w_n24145_0[1]),.dinb(w_asqrt9_2[2]),.dout(n24147),.clk(gclk));
	jxor g23890(.dina(w_n23387_0[0]),.dinb(w_n19791_4[2]),.dout(n24148),.clk(gclk));
	jand g23891(.dina(n24148),.dinb(w_asqrt2_29[0]),.dout(n24149),.clk(gclk));
	jxor g23892(.dina(n24149),.dinb(w_n23392_0[0]),.dout(n24150),.clk(gclk));
	jand g23893(.dina(w_n24150_0[2]),.dinb(n24147),.dout(n24151),.clk(gclk));
	jor g23894(.dina(n24151),.dinb(w_n24146_0[1]),.dout(n24152),.clk(gclk));
	jand g23895(.dina(w_n24152_0[2]),.dinb(w_asqrt10_11[0]),.dout(n24153),.clk(gclk));
	jor g23896(.dina(w_n24152_0[1]),.dinb(w_asqrt10_10[2]),.dout(n24154),.clk(gclk));
	jxor g23897(.dina(w_n23395_0[0]),.dinb(w_n19096_13[1]),.dout(n24155),.clk(gclk));
	jand g23898(.dina(n24155),.dinb(w_asqrt2_28[2]),.dout(n24156),.clk(gclk));
	jxor g23899(.dina(n24156),.dinb(w_n23400_0[0]),.dout(n24157),.clk(gclk));
	jand g23900(.dina(w_n24157_0[2]),.dinb(n24154),.dout(n24158),.clk(gclk));
	jor g23901(.dina(n24158),.dinb(w_n24153_0[1]),.dout(n24159),.clk(gclk));
	jand g23902(.dina(w_n24159_0[2]),.dinb(w_asqrt11_3[0]),.dout(n24160),.clk(gclk));
	jor g23903(.dina(w_n24159_0[1]),.dinb(w_asqrt11_2[2]),.dout(n24161),.clk(gclk));
	jxor g23904(.dina(w_n23403_0[0]),.dinb(w_n18442_5[1]),.dout(n24162),.clk(gclk));
	jand g23905(.dina(n24162),.dinb(w_asqrt2_28[1]),.dout(n24163),.clk(gclk));
	jxor g23906(.dina(n24163),.dinb(w_n23408_0[0]),.dout(n24164),.clk(gclk));
	jand g23907(.dina(w_n24164_0[2]),.dinb(n24161),.dout(n24165),.clk(gclk));
	jor g23908(.dina(n24165),.dinb(w_n24160_0[1]),.dout(n24166),.clk(gclk));
	jand g23909(.dina(w_n24166_0[2]),.dinb(w_asqrt12_11[1]),.dout(n24167),.clk(gclk));
	jor g23910(.dina(w_n24166_0[1]),.dinb(w_asqrt12_11[0]),.dout(n24168),.clk(gclk));
	jxor g23911(.dina(w_n23411_0[0]),.dinb(w_n17769_14[0]),.dout(n24169),.clk(gclk));
	jand g23912(.dina(n24169),.dinb(w_asqrt2_28[0]),.dout(n24170),.clk(gclk));
	jxor g23913(.dina(n24170),.dinb(w_n23416_0[0]),.dout(n24171),.clk(gclk));
	jnot g23914(.din(w_n24171_0[1]),.dout(n24172),.clk(gclk));
	jand g23915(.dina(w_n24172_0[1]),.dinb(n24168),.dout(n24173),.clk(gclk));
	jor g23916(.dina(n24173),.dinb(w_n24167_0[1]),.dout(n24174),.clk(gclk));
	jand g23917(.dina(w_n24174_0[2]),.dinb(w_asqrt13_3[2]),.dout(n24175),.clk(gclk));
	jor g23918(.dina(w_n24174_0[1]),.dinb(w_asqrt13_3[1]),.dout(n24176),.clk(gclk));
	jxor g23919(.dina(w_n23418_0[0]),.dinb(w_n17134_6[1]),.dout(n24177),.clk(gclk));
	jand g23920(.dina(n24177),.dinb(w_asqrt2_27[2]),.dout(n24178),.clk(gclk));
	jxor g23921(.dina(n24178),.dinb(w_n23423_0[0]),.dout(n24179),.clk(gclk));
	jand g23922(.dina(w_n24179_0[2]),.dinb(n24176),.dout(n24180),.clk(gclk));
	jor g23923(.dina(n24180),.dinb(w_n24175_0[1]),.dout(n24181),.clk(gclk));
	jand g23924(.dina(w_n24181_0[2]),.dinb(w_asqrt14_11[2]),.dout(n24182),.clk(gclk));
	jor g23925(.dina(w_n24181_0[1]),.dinb(w_asqrt14_11[1]),.dout(n24183),.clk(gclk));
	jxor g23926(.dina(w_n23426_0[0]),.dinb(w_n16489_14[1]),.dout(n24184),.clk(gclk));
	jand g23927(.dina(n24184),.dinb(w_asqrt2_27[1]),.dout(n24185),.clk(gclk));
	jxor g23928(.dina(n24185),.dinb(w_n23431_0[0]),.dout(n24186),.clk(gclk));
	jnot g23929(.din(w_n24186_0[1]),.dout(n24187),.clk(gclk));
	jand g23930(.dina(w_n24187_0[1]),.dinb(n24183),.dout(n24188),.clk(gclk));
	jor g23931(.dina(n24188),.dinb(w_n24182_0[1]),.dout(n24189),.clk(gclk));
	jand g23932(.dina(w_n24189_0[2]),.dinb(w_asqrt15_4[1]),.dout(n24190),.clk(gclk));
	jor g23933(.dina(w_n24189_0[1]),.dinb(w_asqrt15_4[0]),.dout(n24191),.clk(gclk));
	jxor g23934(.dina(w_n23433_0[0]),.dinb(w_n15878_7[1]),.dout(n24192),.clk(gclk));
	jand g23935(.dina(n24192),.dinb(w_asqrt2_27[0]),.dout(n24193),.clk(gclk));
	jxor g23936(.dina(n24193),.dinb(w_n23438_0[0]),.dout(n24194),.clk(gclk));
	jand g23937(.dina(w_n24194_0[2]),.dinb(n24191),.dout(n24195),.clk(gclk));
	jor g23938(.dina(n24195),.dinb(w_n24190_0[1]),.dout(n24196),.clk(gclk));
	jand g23939(.dina(w_n24196_0[2]),.dinb(w_asqrt16_11[2]),.dout(n24197),.clk(gclk));
	jor g23940(.dina(w_n24196_0[1]),.dinb(w_asqrt16_11[1]),.dout(n24198),.clk(gclk));
	jxor g23941(.dina(w_n23441_0[0]),.dinb(w_n15260_15[0]),.dout(n24199),.clk(gclk));
	jand g23942(.dina(n24199),.dinb(w_asqrt2_26[2]),.dout(n24200),.clk(gclk));
	jxor g23943(.dina(n24200),.dinb(w_n23446_0[0]),.dout(n24201),.clk(gclk));
	jnot g23944(.din(w_n24201_0[1]),.dout(n24202),.clk(gclk));
	jand g23945(.dina(w_n24202_0[1]),.dinb(n24198),.dout(n24203),.clk(gclk));
	jor g23946(.dina(n24203),.dinb(w_n24197_0[1]),.dout(n24204),.clk(gclk));
	jand g23947(.dina(w_n24204_0[2]),.dinb(w_asqrt17_4[2]),.dout(n24205),.clk(gclk));
	jor g23948(.dina(w_n24204_0[1]),.dinb(w_asqrt17_4[1]),.dout(n24206),.clk(gclk));
	jxor g23949(.dina(w_n23448_0[0]),.dinb(w_n14674_8[0]),.dout(n24207),.clk(gclk));
	jand g23950(.dina(n24207),.dinb(w_asqrt2_26[1]),.dout(n24208),.clk(gclk));
	jxor g23951(.dina(n24208),.dinb(w_n23453_0[0]),.dout(n24209),.clk(gclk));
	jnot g23952(.din(w_n24209_0[1]),.dout(n24210),.clk(gclk));
	jand g23953(.dina(w_n24210_0[1]),.dinb(n24206),.dout(n24211),.clk(gclk));
	jor g23954(.dina(n24211),.dinb(w_n24205_0[1]),.dout(n24212),.clk(gclk));
	jand g23955(.dina(w_n24212_0[2]),.dinb(w_asqrt18_12[0]),.dout(n24213),.clk(gclk));
	jor g23956(.dina(w_n24212_0[1]),.dinb(w_asqrt18_11[2]),.dout(n24214),.clk(gclk));
	jxor g23957(.dina(w_n23455_0[0]),.dinb(w_n14078_15[1]),.dout(n24215),.clk(gclk));
	jand g23958(.dina(n24215),.dinb(w_asqrt2_26[0]),.dout(n24216),.clk(gclk));
	jxor g23959(.dina(n24216),.dinb(w_n23460_0[0]),.dout(n24217),.clk(gclk));
	jnot g23960(.din(w_n24217_0[1]),.dout(n24218),.clk(gclk));
	jand g23961(.dina(w_n24218_0[1]),.dinb(n24214),.dout(n24219),.clk(gclk));
	jor g23962(.dina(n24219),.dinb(w_n24213_0[1]),.dout(n24220),.clk(gclk));
	jand g23963(.dina(w_n24220_0[2]),.dinb(w_asqrt19_5[0]),.dout(n24221),.clk(gclk));
	jor g23964(.dina(w_n24220_0[1]),.dinb(w_asqrt19_4[2]),.dout(n24222),.clk(gclk));
	jxor g23965(.dina(w_n23462_0[0]),.dinb(w_n13515_9[0]),.dout(n24223),.clk(gclk));
	jand g23966(.dina(n24223),.dinb(w_asqrt2_25[2]),.dout(n24224),.clk(gclk));
	jxor g23967(.dina(n24224),.dinb(w_n23467_0[0]),.dout(n24225),.clk(gclk));
	jand g23968(.dina(w_n24225_0[2]),.dinb(n24222),.dout(n24226),.clk(gclk));
	jor g23969(.dina(n24226),.dinb(w_n24221_0[1]),.dout(n24227),.clk(gclk));
	jand g23970(.dina(w_n24227_0[2]),.dinb(w_asqrt20_12[0]),.dout(n24228),.clk(gclk));
	jor g23971(.dina(w_n24227_0[1]),.dinb(w_asqrt20_11[2]),.dout(n24229),.clk(gclk));
	jxor g23972(.dina(w_n23470_0[0]),.dinb(w_n12947_16[0]),.dout(n24230),.clk(gclk));
	jand g23973(.dina(n24230),.dinb(w_asqrt2_25[1]),.dout(n24231),.clk(gclk));
	jxor g23974(.dina(n24231),.dinb(w_n23475_0[0]),.dout(n24232),.clk(gclk));
	jnot g23975(.din(w_n24232_0[1]),.dout(n24233),.clk(gclk));
	jand g23976(.dina(w_n24233_0[1]),.dinb(n24229),.dout(n24234),.clk(gclk));
	jor g23977(.dina(n24234),.dinb(w_n24228_0[1]),.dout(n24235),.clk(gclk));
	jand g23978(.dina(w_n24235_0[2]),.dinb(w_asqrt21_5[2]),.dout(n24236),.clk(gclk));
	jor g23979(.dina(w_n24235_0[1]),.dinb(w_asqrt21_5[1]),.dout(n24237),.clk(gclk));
	jxor g23980(.dina(w_n23477_0[0]),.dinb(w_n12410_9[2]),.dout(n24238),.clk(gclk));
	jand g23981(.dina(n24238),.dinb(w_asqrt2_25[0]),.dout(n24239),.clk(gclk));
	jxor g23982(.dina(n24239),.dinb(w_n23482_0[0]),.dout(n24240),.clk(gclk));
	jnot g23983(.din(w_n24240_0[1]),.dout(n24241),.clk(gclk));
	jand g23984(.dina(w_n24241_0[1]),.dinb(n24237),.dout(n24242),.clk(gclk));
	jor g23985(.dina(n24242),.dinb(w_n24236_0[1]),.dout(n24243),.clk(gclk));
	jand g23986(.dina(w_n24243_0[2]),.dinb(w_asqrt22_12[1]),.dout(n24244),.clk(gclk));
	jor g23987(.dina(w_n24243_0[1]),.dinb(w_asqrt22_12[0]),.dout(n24245),.clk(gclk));
	jxor g23988(.dina(w_n23484_0[0]),.dinb(w_n11858_16[1]),.dout(n24246),.clk(gclk));
	jand g23989(.dina(n24246),.dinb(w_asqrt2_24[2]),.dout(n24247),.clk(gclk));
	jxor g23990(.dina(n24247),.dinb(w_n23489_0[0]),.dout(n24248),.clk(gclk));
	jnot g23991(.din(w_n24248_0[1]),.dout(n24249),.clk(gclk));
	jand g23992(.dina(w_n24249_0[1]),.dinb(n24245),.dout(n24250),.clk(gclk));
	jor g23993(.dina(n24250),.dinb(w_n24244_0[1]),.dout(n24251),.clk(gclk));
	jand g23994(.dina(w_n24251_0[2]),.dinb(w_asqrt23_6[1]),.dout(n24252),.clk(gclk));
	jor g23995(.dina(w_n24251_0[1]),.dinb(w_asqrt23_6[0]),.dout(n24253),.clk(gclk));
	jxor g23996(.dina(w_n23491_0[0]),.dinb(w_n11347_10[1]),.dout(n24254),.clk(gclk));
	jand g23997(.dina(n24254),.dinb(w_asqrt2_24[1]),.dout(n24255),.clk(gclk));
	jxor g23998(.dina(n24255),.dinb(w_n23496_0[0]),.dout(n24256),.clk(gclk));
	jand g23999(.dina(w_n24256_0[2]),.dinb(n24253),.dout(n24257),.clk(gclk));
	jor g24000(.dina(n24257),.dinb(w_n24252_0[1]),.dout(n24258),.clk(gclk));
	jand g24001(.dina(w_n24258_0[2]),.dinb(w_asqrt24_12[1]),.dout(n24259),.clk(gclk));
	jor g24002(.dina(w_n24258_0[1]),.dinb(w_asqrt24_12[0]),.dout(n24260),.clk(gclk));
	jxor g24003(.dina(w_n23499_0[0]),.dinb(w_n10824_17[0]),.dout(n24261),.clk(gclk));
	jand g24004(.dina(n24261),.dinb(w_asqrt2_24[0]),.dout(n24262),.clk(gclk));
	jxor g24005(.dina(n24262),.dinb(w_n23504_0[0]),.dout(n24263),.clk(gclk));
	jnot g24006(.din(w_n24263_0[1]),.dout(n24264),.clk(gclk));
	jand g24007(.dina(w_n24264_0[1]),.dinb(n24260),.dout(n24265),.clk(gclk));
	jor g24008(.dina(n24265),.dinb(w_n24259_0[1]),.dout(n24266),.clk(gclk));
	jand g24009(.dina(w_n24266_0[2]),.dinb(w_asqrt25_6[1]),.dout(n24267),.clk(gclk));
	jor g24010(.dina(w_n24266_0[1]),.dinb(w_asqrt25_6[0]),.dout(n24268),.clk(gclk));
	jxor g24011(.dina(w_n23506_0[0]),.dinb(w_n10328_11[1]),.dout(n24269),.clk(gclk));
	jand g24012(.dina(n24269),.dinb(w_asqrt2_23[2]),.dout(n24270),.clk(gclk));
	jxor g24013(.dina(n24270),.dinb(w_n23511_0[0]),.dout(n24271),.clk(gclk));
	jand g24014(.dina(w_n24271_0[2]),.dinb(n24268),.dout(n24272),.clk(gclk));
	jor g24015(.dina(n24272),.dinb(w_n24267_0[1]),.dout(n24273),.clk(gclk));
	jand g24016(.dina(w_n24273_0[2]),.dinb(w_asqrt26_12[1]),.dout(n24274),.clk(gclk));
	jor g24017(.dina(w_n24273_0[1]),.dinb(w_asqrt26_12[0]),.dout(n24275),.clk(gclk));
	jxor g24018(.dina(w_n23514_0[0]),.dinb(w_n9832_17[2]),.dout(n24276),.clk(gclk));
	jand g24019(.dina(n24276),.dinb(w_asqrt2_23[1]),.dout(n24277),.clk(gclk));
	jxor g24020(.dina(n24277),.dinb(w_n23519_0[0]),.dout(n24278),.clk(gclk));
	jnot g24021(.din(w_n24278_0[1]),.dout(n24279),.clk(gclk));
	jand g24022(.dina(w_n24279_0[1]),.dinb(n24275),.dout(n24280),.clk(gclk));
	jor g24023(.dina(n24280),.dinb(w_n24274_0[1]),.dout(n24281),.clk(gclk));
	jand g24024(.dina(w_n24281_0[2]),.dinb(w_asqrt27_7[0]),.dout(n24282),.clk(gclk));
	jor g24025(.dina(w_n24281_0[1]),.dinb(w_asqrt27_6[2]),.dout(n24283),.clk(gclk));
	jxor g24026(.dina(w_n23521_0[0]),.dinb(w_n9369_12[1]),.dout(n24284),.clk(gclk));
	jand g24027(.dina(n24284),.dinb(w_asqrt2_23[0]),.dout(n24285),.clk(gclk));
	jxor g24028(.dina(n24285),.dinb(w_n23526_0[0]),.dout(n24286),.clk(gclk));
	jand g24029(.dina(w_n24286_0[2]),.dinb(n24283),.dout(n24287),.clk(gclk));
	jor g24030(.dina(n24287),.dinb(w_n24282_0[1]),.dout(n24288),.clk(gclk));
	jand g24031(.dina(w_n24288_0[2]),.dinb(w_asqrt28_12[2]),.dout(n24289),.clk(gclk));
	jor g24032(.dina(w_n24288_0[1]),.dinb(w_asqrt28_12[1]),.dout(n24290),.clk(gclk));
	jxor g24033(.dina(w_n23529_0[0]),.dinb(w_n8890_18[0]),.dout(n24291),.clk(gclk));
	jand g24034(.dina(n24291),.dinb(w_asqrt2_22[2]),.dout(n24292),.clk(gclk));
	jxor g24035(.dina(n24292),.dinb(w_n23534_0[0]),.dout(n24293),.clk(gclk));
	jnot g24036(.din(w_n24293_0[1]),.dout(n24294),.clk(gclk));
	jand g24037(.dina(w_n24294_0[1]),.dinb(n24290),.dout(n24295),.clk(gclk));
	jor g24038(.dina(n24295),.dinb(w_n24289_0[1]),.dout(n24296),.clk(gclk));
	jand g24039(.dina(w_n24296_0[2]),.dinb(w_asqrt29_7[1]),.dout(n24297),.clk(gclk));
	jor g24040(.dina(w_n24296_0[1]),.dinb(w_asqrt29_7[0]),.dout(n24298),.clk(gclk));
	jxor g24041(.dina(w_n23536_0[0]),.dinb(w_n8449_13[0]),.dout(n24299),.clk(gclk));
	jand g24042(.dina(n24299),.dinb(w_asqrt2_22[1]),.dout(n24300),.clk(gclk));
	jxor g24043(.dina(n24300),.dinb(w_n23541_0[0]),.dout(n24301),.clk(gclk));
	jnot g24044(.din(w_n24301_0[1]),.dout(n24302),.clk(gclk));
	jand g24045(.dina(w_n24302_0[1]),.dinb(n24298),.dout(n24303),.clk(gclk));
	jor g24046(.dina(n24303),.dinb(w_n24297_0[1]),.dout(n24304),.clk(gclk));
	jand g24047(.dina(w_n24304_0[2]),.dinb(w_asqrt30_13[0]),.dout(n24305),.clk(gclk));
	jor g24048(.dina(w_n24304_0[1]),.dinb(w_asqrt30_12[2]),.dout(n24306),.clk(gclk));
	jxor g24049(.dina(w_n23543_0[0]),.dinb(w_n8003_18[2]),.dout(n24307),.clk(gclk));
	jand g24050(.dina(n24307),.dinb(w_asqrt2_22[0]),.dout(n24308),.clk(gclk));
	jxor g24051(.dina(n24308),.dinb(w_n23548_0[0]),.dout(n24309),.clk(gclk));
	jand g24052(.dina(w_n24309_0[2]),.dinb(n24306),.dout(n24310),.clk(gclk));
	jor g24053(.dina(n24310),.dinb(w_n24305_0[1]),.dout(n24311),.clk(gclk));
	jand g24054(.dina(w_n24311_0[2]),.dinb(w_asqrt31_8[0]),.dout(n24312),.clk(gclk));
	jor g24055(.dina(w_n24311_0[1]),.dinb(w_asqrt31_7[2]),.dout(n24313),.clk(gclk));
	jxor g24056(.dina(w_n23551_0[0]),.dinb(w_n7581_14[0]),.dout(n24314),.clk(gclk));
	jand g24057(.dina(n24314),.dinb(w_asqrt2_21[2]),.dout(n24315),.clk(gclk));
	jxor g24058(.dina(n24315),.dinb(w_n23556_0[0]),.dout(n24316),.clk(gclk));
	jand g24059(.dina(w_n24316_0[2]),.dinb(n24313),.dout(n24317),.clk(gclk));
	jor g24060(.dina(n24317),.dinb(w_n24312_0[1]),.dout(n24318),.clk(gclk));
	jand g24061(.dina(w_n24318_0[2]),.dinb(w_asqrt32_13[0]),.dout(n24319),.clk(gclk));
	jor g24062(.dina(w_n24318_0[1]),.dinb(w_asqrt32_12[2]),.dout(n24320),.clk(gclk));
	jxor g24063(.dina(w_n23559_0[0]),.dinb(w_n7154_19[0]),.dout(n24321),.clk(gclk));
	jand g24064(.dina(n24321),.dinb(w_asqrt2_21[1]),.dout(n24322),.clk(gclk));
	jxor g24065(.dina(n24322),.dinb(w_n23564_0[0]),.dout(n24323),.clk(gclk));
	jnot g24066(.din(w_n24323_0[1]),.dout(n24324),.clk(gclk));
	jand g24067(.dina(w_n24324_0[1]),.dinb(n24320),.dout(n24325),.clk(gclk));
	jor g24068(.dina(n24325),.dinb(w_n24319_0[1]),.dout(n24326),.clk(gclk));
	jand g24069(.dina(w_n24326_0[2]),.dinb(w_asqrt33_8[2]),.dout(n24327),.clk(gclk));
	jor g24070(.dina(w_n24326_0[1]),.dinb(w_asqrt33_8[1]),.dout(n24328),.clk(gclk));
	jxor g24071(.dina(w_n23566_0[0]),.dinb(w_n6758_14[2]),.dout(n24329),.clk(gclk));
	jand g24072(.dina(n24329),.dinb(w_asqrt2_21[0]),.dout(n24330),.clk(gclk));
	jxor g24073(.dina(n24330),.dinb(w_n23571_0[0]),.dout(n24331),.clk(gclk));
	jand g24074(.dina(w_n24331_0[2]),.dinb(n24328),.dout(n24332),.clk(gclk));
	jor g24075(.dina(n24332),.dinb(w_n24327_0[1]),.dout(n24333),.clk(gclk));
	jand g24076(.dina(w_n24333_0[2]),.dinb(w_asqrt34_13[1]),.dout(n24334),.clk(gclk));
	jor g24077(.dina(w_n24333_0[1]),.dinb(w_asqrt34_13[0]),.dout(n24335),.clk(gclk));
	jxor g24078(.dina(w_n23574_0[0]),.dinb(w_n6357_19[1]),.dout(n24336),.clk(gclk));
	jand g24079(.dina(n24336),.dinb(w_asqrt2_20[2]),.dout(n24337),.clk(gclk));
	jxor g24080(.dina(n24337),.dinb(w_n23579_0[0]),.dout(n24338),.clk(gclk));
	jnot g24081(.din(w_n24338_0[1]),.dout(n24339),.clk(gclk));
	jand g24082(.dina(w_n24339_0[1]),.dinb(n24335),.dout(n24340),.clk(gclk));
	jor g24083(.dina(n24340),.dinb(w_n24334_0[1]),.dout(n24341),.clk(gclk));
	jand g24084(.dina(w_n24341_0[2]),.dinb(w_asqrt35_9[1]),.dout(n24342),.clk(gclk));
	jor g24085(.dina(w_n24341_0[1]),.dinb(w_asqrt35_9[0]),.dout(n24343),.clk(gclk));
	jxor g24086(.dina(w_n23581_0[0]),.dinb(w_n5989_15[1]),.dout(n24344),.clk(gclk));
	jand g24087(.dina(n24344),.dinb(w_asqrt2_20[1]),.dout(n24345),.clk(gclk));
	jxor g24088(.dina(n24345),.dinb(w_n23586_0[0]),.dout(n24346),.clk(gclk));
	jand g24089(.dina(w_n24346_0[2]),.dinb(n24343),.dout(n24347),.clk(gclk));
	jor g24090(.dina(n24347),.dinb(w_n24342_0[1]),.dout(n24348),.clk(gclk));
	jand g24091(.dina(w_n24348_0[2]),.dinb(w_asqrt36_13[1]),.dout(n24349),.clk(gclk));
	jor g24092(.dina(w_n24348_0[1]),.dinb(w_asqrt36_13[0]),.dout(n24350),.clk(gclk));
	jxor g24093(.dina(w_n23589_0[0]),.dinb(w_n5606_19[2]),.dout(n24351),.clk(gclk));
	jand g24094(.dina(n24351),.dinb(w_asqrt2_20[0]),.dout(n24352),.clk(gclk));
	jxor g24095(.dina(n24352),.dinb(w_n23594_0[0]),.dout(n24353),.clk(gclk));
	jnot g24096(.din(w_n24353_0[1]),.dout(n24354),.clk(gclk));
	jand g24097(.dina(w_n24354_0[1]),.dinb(n24350),.dout(n24355),.clk(gclk));
	jor g24098(.dina(n24355),.dinb(w_n24349_0[1]),.dout(n24356),.clk(gclk));
	jand g24099(.dina(w_n24356_0[2]),.dinb(w_asqrt37_9[2]),.dout(n24357),.clk(gclk));
	jor g24100(.dina(w_n24356_0[1]),.dinb(w_asqrt37_9[1]),.dout(n24358),.clk(gclk));
	jxor g24101(.dina(w_n23596_0[0]),.dinb(w_n5259_16[1]),.dout(n24359),.clk(gclk));
	jand g24102(.dina(n24359),.dinb(w_asqrt2_19[2]),.dout(n24360),.clk(gclk));
	jxor g24103(.dina(n24360),.dinb(w_n23601_0[0]),.dout(n24361),.clk(gclk));
	jnot g24104(.din(w_n24361_0[1]),.dout(n24362),.clk(gclk));
	jand g24105(.dina(w_n24362_0[1]),.dinb(n24358),.dout(n24363),.clk(gclk));
	jor g24106(.dina(n24363),.dinb(w_n24357_0[1]),.dout(n24364),.clk(gclk));
	jand g24107(.dina(w_n24364_0[2]),.dinb(w_asqrt38_13[2]),.dout(n24365),.clk(gclk));
	jor g24108(.dina(w_n24364_0[1]),.dinb(w_asqrt38_13[1]),.dout(n24366),.clk(gclk));
	jxor g24109(.dina(w_n23603_0[0]),.dinb(w_n4902_20[1]),.dout(n24367),.clk(gclk));
	jand g24110(.dina(n24367),.dinb(w_asqrt2_19[1]),.dout(n24368),.clk(gclk));
	jxor g24111(.dina(n24368),.dinb(w_n23608_0[0]),.dout(n24369),.clk(gclk));
	jnot g24112(.din(w_n24369_0[1]),.dout(n24370),.clk(gclk));
	jand g24113(.dina(w_n24370_0[1]),.dinb(n24366),.dout(n24371),.clk(gclk));
	jor g24114(.dina(n24371),.dinb(w_n24365_0[1]),.dout(n24372),.clk(gclk));
	jand g24115(.dina(w_n24372_0[2]),.dinb(w_asqrt39_10[1]),.dout(n24373),.clk(gclk));
	jor g24116(.dina(w_n24372_0[1]),.dinb(w_asqrt39_10[0]),.dout(n24374),.clk(gclk));
	jxor g24117(.dina(w_n23610_0[0]),.dinb(w_n4582_17[1]),.dout(n24375),.clk(gclk));
	jand g24118(.dina(n24375),.dinb(w_asqrt2_19[0]),.dout(n24376),.clk(gclk));
	jxor g24119(.dina(n24376),.dinb(w_n23615_0[0]),.dout(n24377),.clk(gclk));
	jand g24120(.dina(w_n24377_0[2]),.dinb(n24374),.dout(n24378),.clk(gclk));
	jor g24121(.dina(n24378),.dinb(w_n24373_0[1]),.dout(n24379),.clk(gclk));
	jand g24122(.dina(w_n24379_0[2]),.dinb(w_asqrt40_13[2]),.dout(n24380),.clk(gclk));
	jor g24123(.dina(w_n24379_0[1]),.dinb(w_asqrt40_13[1]),.dout(n24381),.clk(gclk));
	jxor g24124(.dina(w_n23618_0[0]),.dinb(w_n4249_21[0]),.dout(n24382),.clk(gclk));
	jand g24125(.dina(n24382),.dinb(w_asqrt2_18[2]),.dout(n24383),.clk(gclk));
	jxor g24126(.dina(n24383),.dinb(w_n23623_0[0]),.dout(n24384),.clk(gclk));
	jnot g24127(.din(w_n24384_0[1]),.dout(n24385),.clk(gclk));
	jand g24128(.dina(w_n24385_0[1]),.dinb(n24381),.dout(n24386),.clk(gclk));
	jor g24129(.dina(n24386),.dinb(w_n24380_0[1]),.dout(n24387),.clk(gclk));
	jand g24130(.dina(w_n24387_0[2]),.dinb(w_asqrt41_10[2]),.dout(n24388),.clk(gclk));
	jor g24131(.dina(w_n24387_0[1]),.dinb(w_asqrt41_10[1]),.dout(n24389),.clk(gclk));
	jxor g24132(.dina(w_n23625_0[0]),.dinb(w_n3955_18[0]),.dout(n24390),.clk(gclk));
	jand g24133(.dina(n24390),.dinb(w_asqrt2_18[1]),.dout(n24391),.clk(gclk));
	jxor g24134(.dina(n24391),.dinb(w_n23630_0[0]),.dout(n24392),.clk(gclk));
	jand g24135(.dina(w_n24392_0[2]),.dinb(n24389),.dout(n24393),.clk(gclk));
	jor g24136(.dina(n24393),.dinb(w_n24388_0[1]),.dout(n24394),.clk(gclk));
	jand g24137(.dina(w_n24394_0[2]),.dinb(w_asqrt42_14[0]),.dout(n24395),.clk(gclk));
	jor g24138(.dina(w_n24394_0[1]),.dinb(w_asqrt42_13[2]),.dout(n24396),.clk(gclk));
	jxor g24139(.dina(w_n23633_0[0]),.dinb(w_n3642_21[1]),.dout(n24397),.clk(gclk));
	jand g24140(.dina(n24397),.dinb(w_asqrt2_18[0]),.dout(n24398),.clk(gclk));
	jxor g24141(.dina(n24398),.dinb(w_n23638_0[0]),.dout(n24399),.clk(gclk));
	jnot g24142(.din(w_n24399_0[1]),.dout(n24400),.clk(gclk));
	jand g24143(.dina(w_n24400_0[1]),.dinb(n24396),.dout(n24401),.clk(gclk));
	jor g24144(.dina(n24401),.dinb(w_n24395_0[1]),.dout(n24402),.clk(gclk));
	jand g24145(.dina(w_n24402_0[2]),.dinb(w_asqrt43_11[0]),.dout(n24403),.clk(gclk));
	jor g24146(.dina(w_n24402_0[1]),.dinb(w_asqrt43_10[2]),.dout(n24404),.clk(gclk));
	jxor g24147(.dina(w_n23640_0[0]),.dinb(w_n3368_18[2]),.dout(n24405),.clk(gclk));
	jand g24148(.dina(n24405),.dinb(w_asqrt2_17[2]),.dout(n24406),.clk(gclk));
	jxor g24149(.dina(n24406),.dinb(w_n23645_0[0]),.dout(n24407),.clk(gclk));
	jand g24150(.dina(w_n24407_0[2]),.dinb(n24404),.dout(n24408),.clk(gclk));
	jor g24151(.dina(n24408),.dinb(w_n24403_0[1]),.dout(n24409),.clk(gclk));
	jand g24152(.dina(w_n24409_0[2]),.dinb(w_asqrt44_14[0]),.dout(n24410),.clk(gclk));
	jor g24153(.dina(w_n24409_0[1]),.dinb(w_asqrt44_13[2]),.dout(n24411),.clk(gclk));
	jxor g24154(.dina(w_n23648_0[0]),.dinb(w_n3089_22[0]),.dout(n24412),.clk(gclk));
	jand g24155(.dina(n24412),.dinb(w_asqrt2_17[1]),.dout(n24413),.clk(gclk));
	jxor g24156(.dina(n24413),.dinb(w_n23653_0[0]),.dout(n24414),.clk(gclk));
	jnot g24157(.din(w_n24414_0[1]),.dout(n24415),.clk(gclk));
	jand g24158(.dina(w_n24415_0[1]),.dinb(n24411),.dout(n24416),.clk(gclk));
	jor g24159(.dina(n24416),.dinb(w_n24410_0[1]),.dout(n24417),.clk(gclk));
	jand g24160(.dina(w_n24417_0[2]),.dinb(w_asqrt45_11[2]),.dout(n24418),.clk(gclk));
	jor g24161(.dina(w_n24417_0[1]),.dinb(w_asqrt45_11[1]),.dout(n24419),.clk(gclk));
	jxor g24162(.dina(w_n23655_0[0]),.dinb(w_n2833_19[2]),.dout(n24420),.clk(gclk));
	jand g24163(.dina(n24420),.dinb(w_asqrt2_17[0]),.dout(n24421),.clk(gclk));
	jxor g24164(.dina(n24421),.dinb(w_n23660_0[0]),.dout(n24422),.clk(gclk));
	jand g24165(.dina(w_n24422_0[2]),.dinb(n24419),.dout(n24423),.clk(gclk));
	jor g24166(.dina(n24423),.dinb(w_n24418_0[1]),.dout(n24424),.clk(gclk));
	jand g24167(.dina(w_n24424_0[2]),.dinb(w_asqrt46_14[0]),.dout(n24425),.clk(gclk));
	jor g24168(.dina(w_n24424_0[1]),.dinb(w_asqrt46_13[2]),.dout(n24426),.clk(gclk));
	jxor g24169(.dina(w_n23663_0[0]),.dinb(w_n2572_22[1]),.dout(n24427),.clk(gclk));
	jand g24170(.dina(n24427),.dinb(w_asqrt2_16[2]),.dout(n24428),.clk(gclk));
	jxor g24171(.dina(n24428),.dinb(w_n23668_0[0]),.dout(n24429),.clk(gclk));
	jnot g24172(.din(w_n24429_0[1]),.dout(n24430),.clk(gclk));
	jand g24173(.dina(w_n24430_0[1]),.dinb(n24426),.dout(n24431),.clk(gclk));
	jor g24174(.dina(n24431),.dinb(w_n24425_0[1]),.dout(n24432),.clk(gclk));
	jand g24175(.dina(w_n24432_0[2]),.dinb(w_asqrt47_12[1]),.dout(n24433),.clk(gclk));
	jor g24176(.dina(w_n24432_0[1]),.dinb(w_asqrt47_12[0]),.dout(n24434),.clk(gclk));
	jxor g24177(.dina(w_n23670_0[0]),.dinb(w_n2345_20[1]),.dout(n24435),.clk(gclk));
	jand g24178(.dina(n24435),.dinb(w_asqrt2_16[1]),.dout(n24436),.clk(gclk));
	jxor g24179(.dina(n24436),.dinb(w_n23675_0[0]),.dout(n24437),.clk(gclk));
	jnot g24180(.din(w_n24437_0[1]),.dout(n24438),.clk(gclk));
	jand g24181(.dina(w_n24438_0[1]),.dinb(n24434),.dout(n24439),.clk(gclk));
	jor g24182(.dina(n24439),.dinb(w_n24433_0[1]),.dout(n24440),.clk(gclk));
	jand g24183(.dina(w_n24440_0[2]),.dinb(w_asqrt48_14[1]),.dout(n24441),.clk(gclk));
	jor g24184(.dina(w_n24440_0[1]),.dinb(w_asqrt48_14[0]),.dout(n24442),.clk(gclk));
	jxor g24185(.dina(w_n23677_0[0]),.dinb(w_n2108_23[0]),.dout(n24443),.clk(gclk));
	jand g24186(.dina(n24443),.dinb(w_asqrt2_16[0]),.dout(n24444),.clk(gclk));
	jxor g24187(.dina(n24444),.dinb(w_n23682_0[0]),.dout(n24445),.clk(gclk));
	jnot g24188(.din(w_n24445_0[1]),.dout(n24446),.clk(gclk));
	jand g24189(.dina(w_n24446_0[1]),.dinb(n24442),.dout(n24447),.clk(gclk));
	jor g24190(.dina(n24447),.dinb(w_n24441_0[1]),.dout(n24448),.clk(gclk));
	jand g24191(.dina(w_n24448_0[2]),.dinb(w_asqrt49_12[2]),.dout(n24449),.clk(gclk));
	jor g24192(.dina(w_n24448_0[1]),.dinb(w_asqrt49_12[1]),.dout(n24450),.clk(gclk));
	jxor g24193(.dina(w_n23684_0[0]),.dinb(w_n1912_21[1]),.dout(n24451),.clk(gclk));
	jand g24194(.dina(n24451),.dinb(w_asqrt2_15[2]),.dout(n24452),.clk(gclk));
	jxor g24195(.dina(n24452),.dinb(w_n23689_0[0]),.dout(n24453),.clk(gclk));
	jand g24196(.dina(w_n24453_0[2]),.dinb(n24450),.dout(n24454),.clk(gclk));
	jor g24197(.dina(n24454),.dinb(w_n24449_0[1]),.dout(n24455),.clk(gclk));
	jand g24198(.dina(w_n24455_0[2]),.dinb(w_asqrt50_14[2]),.dout(n24456),.clk(gclk));
	jor g24199(.dina(w_n24455_0[1]),.dinb(w_asqrt50_14[1]),.dout(n24457),.clk(gclk));
	jxor g24200(.dina(w_n23692_0[0]),.dinb(w_n1699_23[2]),.dout(n24458),.clk(gclk));
	jand g24201(.dina(n24458),.dinb(w_asqrt2_15[1]),.dout(n24459),.clk(gclk));
	jxor g24202(.dina(n24459),.dinb(w_n23697_0[0]),.dout(n24460),.clk(gclk));
	jnot g24203(.din(w_n24460_0[1]),.dout(n24461),.clk(gclk));
	jand g24204(.dina(w_n24461_0[1]),.dinb(n24457),.dout(n24462),.clk(gclk));
	jor g24205(.dina(n24462),.dinb(w_n24456_0[1]),.dout(n24463),.clk(gclk));
	jand g24206(.dina(w_n24463_0[2]),.dinb(w_asqrt51_13[0]),.dout(n24464),.clk(gclk));
	jor g24207(.dina(w_n24463_0[1]),.dinb(w_asqrt51_12[2]),.dout(n24465),.clk(gclk));
	jxor g24208(.dina(w_n23699_0[0]),.dinb(w_n1516_22[0]),.dout(n24466),.clk(gclk));
	jand g24209(.dina(n24466),.dinb(w_asqrt2_15[0]),.dout(n24467),.clk(gclk));
	jxor g24210(.dina(n24467),.dinb(w_n23704_0[0]),.dout(n24468),.clk(gclk));
	jnot g24211(.din(w_n24468_0[1]),.dout(n24469),.clk(gclk));
	jand g24212(.dina(w_n24469_0[1]),.dinb(n24465),.dout(n24470),.clk(gclk));
	jor g24213(.dina(n24470),.dinb(w_n24464_0[1]),.dout(n24471),.clk(gclk));
	jand g24214(.dina(w_n24471_0[2]),.dinb(w_asqrt52_14[2]),.dout(n24472),.clk(gclk));
	jor g24215(.dina(w_n24471_0[1]),.dinb(w_asqrt52_14[1]),.dout(n24473),.clk(gclk));
	jxor g24216(.dina(w_n23706_0[0]),.dinb(w_n1332_23[2]),.dout(n24474),.clk(gclk));
	jand g24217(.dina(n24474),.dinb(w_asqrt2_14[2]),.dout(n24475),.clk(gclk));
	jxor g24218(.dina(n24475),.dinb(w_n23711_0[0]),.dout(n24476),.clk(gclk));
	jnot g24219(.din(w_n24476_0[1]),.dout(n24477),.clk(gclk));
	jand g24220(.dina(w_n24477_0[1]),.dinb(n24473),.dout(n24478),.clk(gclk));
	jor g24221(.dina(n24478),.dinb(w_n24472_0[1]),.dout(n24479),.clk(gclk));
	jand g24222(.dina(w_n24479_0[2]),.dinb(w_asqrt53_13[2]),.dout(n24480),.clk(gclk));
	jor g24223(.dina(w_n24479_0[1]),.dinb(w_asqrt53_13[1]),.dout(n24481),.clk(gclk));
	jxor g24224(.dina(w_n23713_0[0]),.dinb(w_n1173_22[2]),.dout(n24482),.clk(gclk));
	jand g24225(.dina(n24482),.dinb(w_asqrt2_14[1]),.dout(n24483),.clk(gclk));
	jxor g24226(.dina(n24483),.dinb(w_n23718_0[0]),.dout(n24484),.clk(gclk));
	jnot g24227(.din(w_n24484_0[1]),.dout(n24485),.clk(gclk));
	jand g24228(.dina(w_n24485_0[1]),.dinb(n24481),.dout(n24486),.clk(gclk));
	jor g24229(.dina(n24486),.dinb(w_n24480_0[1]),.dout(n24487),.clk(gclk));
	jand g24230(.dina(w_n24487_0[2]),.dinb(w_asqrt54_14[2]),.dout(n24488),.clk(gclk));
	jor g24231(.dina(w_n24487_0[1]),.dinb(w_asqrt54_14[1]),.dout(n24489),.clk(gclk));
	jxor g24232(.dina(w_n23720_0[0]),.dinb(w_n1008_24[2]),.dout(n24490),.clk(gclk));
	jand g24233(.dina(n24490),.dinb(w_asqrt2_14[0]),.dout(n24491),.clk(gclk));
	jxor g24234(.dina(n24491),.dinb(w_n23725_0[0]),.dout(n24492),.clk(gclk));
	jnot g24235(.din(w_n24492_0[1]),.dout(n24493),.clk(gclk));
	jand g24236(.dina(w_n24493_0[1]),.dinb(n24489),.dout(n24494),.clk(gclk));
	jor g24237(.dina(n24494),.dinb(w_n24488_0[1]),.dout(n24495),.clk(gclk));
	jand g24238(.dina(w_n24495_0[2]),.dinb(w_asqrt55_14[0]),.dout(n24496),.clk(gclk));
	jor g24239(.dina(w_n24495_0[1]),.dinb(w_asqrt55_13[2]),.dout(n24497),.clk(gclk));
	jxor g24240(.dina(w_n23727_0[0]),.dinb(w_n884_23[2]),.dout(n24498),.clk(gclk));
	jand g24241(.dina(n24498),.dinb(w_asqrt2_13[2]),.dout(n24499),.clk(gclk));
	jxor g24242(.dina(n24499),.dinb(w_n23732_0[0]),.dout(n24500),.clk(gclk));
	jand g24243(.dina(w_n24500_0[2]),.dinb(n24497),.dout(n24501),.clk(gclk));
	jor g24244(.dina(n24501),.dinb(w_n24496_0[1]),.dout(n24502),.clk(gclk));
	jand g24245(.dina(w_n24502_0[2]),.dinb(w_asqrt56_15[0]),.dout(n24503),.clk(gclk));
	jor g24246(.dina(w_n24502_0[1]),.dinb(w_asqrt56_14[2]),.dout(n24504),.clk(gclk));
	jxor g24247(.dina(w_n23735_0[0]),.dinb(w_n743_24[2]),.dout(n24505),.clk(gclk));
	jand g24248(.dina(n24505),.dinb(w_asqrt2_13[1]),.dout(n24506),.clk(gclk));
	jxor g24249(.dina(n24506),.dinb(w_n23740_0[0]),.dout(n24507),.clk(gclk));
	jnot g24250(.din(w_n24507_0[1]),.dout(n24508),.clk(gclk));
	jand g24251(.dina(w_n24508_0[1]),.dinb(n24504),.dout(n24509),.clk(gclk));
	jor g24252(.dina(n24509),.dinb(w_n24503_0[1]),.dout(n24510),.clk(gclk));
	jand g24253(.dina(w_n24510_0[2]),.dinb(w_asqrt57_14[2]),.dout(n24511),.clk(gclk));
	jor g24254(.dina(w_n24510_0[1]),.dinb(w_asqrt57_14[1]),.dout(n24512),.clk(gclk));
	jxor g24255(.dina(w_n23742_0[0]),.dinb(w_n635_24[2]),.dout(n24513),.clk(gclk));
	jand g24256(.dina(n24513),.dinb(w_asqrt2_13[0]),.dout(n24514),.clk(gclk));
	jxor g24257(.dina(n24514),.dinb(w_n23747_0[0]),.dout(n24515),.clk(gclk));
	jand g24258(.dina(w_n24515_0[2]),.dinb(n24512),.dout(n24516),.clk(gclk));
	jor g24259(.dina(n24516),.dinb(w_n24511_0[1]),.dout(n24517),.clk(gclk));
	jand g24260(.dina(w_n24517_0[2]),.dinb(w_asqrt58_15[1]),.dout(n24518),.clk(gclk));
	jor g24261(.dina(w_n24517_0[1]),.dinb(w_asqrt58_15[0]),.dout(n24519),.clk(gclk));
	jxor g24262(.dina(w_n23750_0[0]),.dinb(w_n515_25[2]),.dout(n24520),.clk(gclk));
	jand g24263(.dina(n24520),.dinb(w_asqrt2_12[2]),.dout(n24521),.clk(gclk));
	jxor g24264(.dina(n24521),.dinb(w_n23755_0[0]),.dout(n24522),.clk(gclk));
	jnot g24265(.din(w_n24522_0[1]),.dout(n24523),.clk(gclk));
	jand g24266(.dina(w_n24523_0[1]),.dinb(n24519),.dout(n24524),.clk(gclk));
	jor g24267(.dina(n24524),.dinb(w_n24518_0[1]),.dout(n24525),.clk(gclk));
	jand g24268(.dina(w_n24525_0[2]),.dinb(w_asqrt59_15[0]),.dout(n24526),.clk(gclk));
	jor g24269(.dina(w_n24525_0[1]),.dinb(w_asqrt59_14[2]),.dout(n24527),.clk(gclk));
	jxor g24270(.dina(w_n23757_0[0]),.dinb(w_n443_25[2]),.dout(n24528),.clk(gclk));
	jand g24271(.dina(n24528),.dinb(w_asqrt2_12[1]),.dout(n24529),.clk(gclk));
	jxor g24272(.dina(n24529),.dinb(w_n24080_0[0]),.dout(n24530),.clk(gclk));
	jand g24273(.dina(w_n24530_0[2]),.dinb(n24527),.dout(n24531),.clk(gclk));
	jor g24274(.dina(n24531),.dinb(w_n24526_0[1]),.dout(n24532),.clk(gclk));
	jand g24275(.dina(w_n24532_0[2]),.dinb(w_asqrt60_15[1]),.dout(n24533),.clk(gclk));
	jor g24276(.dina(w_n24532_0[1]),.dinb(w_asqrt60_15[0]),.dout(n24534),.clk(gclk));
	jxor g24277(.dina(w_n23764_0[0]),.dinb(w_n352_26[0]),.dout(n24535),.clk(gclk));
	jand g24278(.dina(n24535),.dinb(w_asqrt2_12[0]),.dout(n24536),.clk(gclk));
	jxor g24279(.dina(n24536),.dinb(w_n23769_0[0]),.dout(n24537),.clk(gclk));
	jand g24280(.dina(w_n24537_0[2]),.dinb(n24534),.dout(n24538),.clk(gclk));
	jor g24281(.dina(n24538),.dinb(w_n24533_0[1]),.dout(n24539),.clk(gclk));
	jand g24282(.dina(w_n24539_0[2]),.dinb(w_asqrt61_15[1]),.dout(n24540),.clk(gclk));
	jor g24283(.dina(w_n24539_0[1]),.dinb(w_asqrt61_15[0]),.dout(n24541),.clk(gclk));
	jxor g24284(.dina(w_n23772_0[0]),.dinb(w_n294_26[1]),.dout(n24542),.clk(gclk));
	jand g24285(.dina(n24542),.dinb(w_asqrt2_11[2]),.dout(n24543),.clk(gclk));
	jxor g24286(.dina(n24543),.dinb(w_n23777_0[0]),.dout(n24544),.clk(gclk));
	jand g24287(.dina(w_n24544_0[2]),.dinb(n24541),.dout(n24545),.clk(gclk));
	jor g24288(.dina(n24545),.dinb(w_n24540_0[1]),.dout(n24546),.clk(gclk));
	jand g24289(.dina(w_n24546_0[2]),.dinb(w_asqrt62_15[1]),.dout(n24547),.clk(gclk));
	jor g24290(.dina(w_n24546_0[1]),.dinb(w_asqrt62_15[0]),.dout(n24548),.clk(gclk));
	jxor g24291(.dina(w_n23780_0[0]),.dinb(w_n239_26[1]),.dout(n24549),.clk(gclk));
	jand g24292(.dina(n24549),.dinb(w_asqrt2_11[1]),.dout(n24550),.clk(gclk));
	jxor g24293(.dina(n24550),.dinb(w_n23785_0[0]),.dout(n24551),.clk(gclk));
	jnot g24294(.din(w_n24551_0[1]),.dout(n24552),.clk(gclk));
	jand g24295(.dina(w_n24552_0[1]),.dinb(n24548),.dout(n24553),.clk(gclk));
	jor g24296(.dina(n24553),.dinb(w_n24547_0[1]),.dout(n24554),.clk(gclk));
	jand g24297(.dina(w_n23806_0[0]),.dinb(w_n24097_0[0]),.dout(n24555),.clk(gclk));
	jnot g24298(.din(w_n24547_0[0]),.dout(n24556),.clk(gclk));
	jnot g24299(.din(w_n24540_0[0]),.dout(n24557),.clk(gclk));
	jnot g24300(.din(w_n24533_0[0]),.dout(n24558),.clk(gclk));
	jnot g24301(.din(w_n24526_0[0]),.dout(n24559),.clk(gclk));
	jnot g24302(.din(w_n24518_0[0]),.dout(n24560),.clk(gclk));
	jnot g24303(.din(w_n24511_0[0]),.dout(n24561),.clk(gclk));
	jnot g24304(.din(w_n24503_0[0]),.dout(n24562),.clk(gclk));
	jnot g24305(.din(w_n24496_0[0]),.dout(n24563),.clk(gclk));
	jnot g24306(.din(w_n24488_0[0]),.dout(n24564),.clk(gclk));
	jnot g24307(.din(w_n24480_0[0]),.dout(n24565),.clk(gclk));
	jnot g24308(.din(w_n24472_0[0]),.dout(n24566),.clk(gclk));
	jnot g24309(.din(w_n24464_0[0]),.dout(n24567),.clk(gclk));
	jnot g24310(.din(w_n24456_0[0]),.dout(n24568),.clk(gclk));
	jnot g24311(.din(w_n24449_0[0]),.dout(n24569),.clk(gclk));
	jnot g24312(.din(w_n24441_0[0]),.dout(n24570),.clk(gclk));
	jnot g24313(.din(w_n24433_0[0]),.dout(n24571),.clk(gclk));
	jnot g24314(.din(w_n24425_0[0]),.dout(n24572),.clk(gclk));
	jnot g24315(.din(w_n24418_0[0]),.dout(n24573),.clk(gclk));
	jnot g24316(.din(w_n24410_0[0]),.dout(n24574),.clk(gclk));
	jnot g24317(.din(w_n24403_0[0]),.dout(n24575),.clk(gclk));
	jnot g24318(.din(w_n24395_0[0]),.dout(n24576),.clk(gclk));
	jnot g24319(.din(w_n24388_0[0]),.dout(n24577),.clk(gclk));
	jnot g24320(.din(w_n24380_0[0]),.dout(n24578),.clk(gclk));
	jnot g24321(.din(w_n24373_0[0]),.dout(n24579),.clk(gclk));
	jnot g24322(.din(w_n24365_0[0]),.dout(n24580),.clk(gclk));
	jnot g24323(.din(w_n24357_0[0]),.dout(n24581),.clk(gclk));
	jnot g24324(.din(w_n24349_0[0]),.dout(n24582),.clk(gclk));
	jnot g24325(.din(w_n24342_0[0]),.dout(n24583),.clk(gclk));
	jnot g24326(.din(w_n24334_0[0]),.dout(n24584),.clk(gclk));
	jnot g24327(.din(w_n24327_0[0]),.dout(n24585),.clk(gclk));
	jnot g24328(.din(w_n24319_0[0]),.dout(n24586),.clk(gclk));
	jnot g24329(.din(w_n24312_0[0]),.dout(n24587),.clk(gclk));
	jnot g24330(.din(w_n24305_0[0]),.dout(n24588),.clk(gclk));
	jnot g24331(.din(w_n24297_0[0]),.dout(n24589),.clk(gclk));
	jnot g24332(.din(w_n24289_0[0]),.dout(n24590),.clk(gclk));
	jnot g24333(.din(w_n24282_0[0]),.dout(n24591),.clk(gclk));
	jnot g24334(.din(w_n24274_0[0]),.dout(n24592),.clk(gclk));
	jnot g24335(.din(w_n24267_0[0]),.dout(n24593),.clk(gclk));
	jnot g24336(.din(w_n24259_0[0]),.dout(n24594),.clk(gclk));
	jnot g24337(.din(w_n24252_0[0]),.dout(n24595),.clk(gclk));
	jnot g24338(.din(w_n24244_0[0]),.dout(n24596),.clk(gclk));
	jnot g24339(.din(w_n24236_0[0]),.dout(n24597),.clk(gclk));
	jnot g24340(.din(w_n24228_0[0]),.dout(n24598),.clk(gclk));
	jnot g24341(.din(w_n24221_0[0]),.dout(n24599),.clk(gclk));
	jnot g24342(.din(w_n24213_0[0]),.dout(n24600),.clk(gclk));
	jnot g24343(.din(w_n24205_0[0]),.dout(n24601),.clk(gclk));
	jnot g24344(.din(w_n24197_0[0]),.dout(n24602),.clk(gclk));
	jnot g24345(.din(w_n24190_0[0]),.dout(n24603),.clk(gclk));
	jnot g24346(.din(w_n24182_0[0]),.dout(n24604),.clk(gclk));
	jnot g24347(.din(w_n24175_0[0]),.dout(n24605),.clk(gclk));
	jnot g24348(.din(w_n24167_0[0]),.dout(n24606),.clk(gclk));
	jnot g24349(.din(w_n24160_0[0]),.dout(n24607),.clk(gclk));
	jnot g24350(.din(w_n24153_0[0]),.dout(n24608),.clk(gclk));
	jnot g24351(.din(w_n24146_0[0]),.dout(n24609),.clk(gclk));
	jnot g24352(.din(w_n24138_0[0]),.dout(n24610),.clk(gclk));
	jnot g24353(.din(w_n24130_0[0]),.dout(n24611),.clk(gclk));
	jnot g24354(.din(w_n24123_0[0]),.dout(n24612),.clk(gclk));
	jnot g24355(.din(w_n24116_0[0]),.dout(n24613),.clk(gclk));
	jnot g24356(.din(w_n24108_0[0]),.dout(n24614),.clk(gclk));
	jnot g24357(.din(w_n23813_0[0]),.dout(n24615),.clk(gclk));
	jor g24358(.dina(w_n24103_1[1]),.dinb(w_n23351_0[1]),.dout(n24616),.clk(gclk));
	jnot g24359(.din(w_n23811_0[0]),.dout(n24617),.clk(gclk));
	jand g24360(.dina(n24617),.dinb(n24616),.dout(n24618),.clk(gclk));
	jand g24361(.dina(n24618),.dinb(w_n23345_11[2]),.dout(n24619),.clk(gclk));
	jor g24362(.dina(w_n24103_1[0]),.dinb(w_a4_0[2]),.dout(n24620),.clk(gclk));
	jand g24363(.dina(n24620),.dinb(w_a5_0[0]),.dout(n24621),.clk(gclk));
	jand g24364(.dina(w_asqrt2_11[0]),.dinb(w_n23353_0[0]),.dout(n24622),.clk(gclk));
	jor g24365(.dina(n24622),.dinb(n24621),.dout(n24623),.clk(gclk));
	jor g24366(.dina(n24623),.dinb(n24619),.dout(n24624),.clk(gclk));
	jand g24367(.dina(n24624),.dinb(n24615),.dout(n24625),.clk(gclk));
	jand g24368(.dina(n24625),.dinb(w_n22620_2[1]),.dout(n24626),.clk(gclk));
	jor g24369(.dina(w_n24112_0[0]),.dinb(n24626),.dout(n24627),.clk(gclk));
	jand g24370(.dina(n24627),.dinb(n24614),.dout(n24628),.clk(gclk));
	jand g24371(.dina(n24628),.dinb(w_n21887_12[1]),.dout(n24629),.clk(gclk));
	jnot g24372(.din(w_n24120_0[1]),.dout(n24630),.clk(gclk));
	jor g24373(.dina(n24630),.dinb(n24629),.dout(n24631),.clk(gclk));
	jand g24374(.dina(n24631),.dinb(n24613),.dout(n24632),.clk(gclk));
	jand g24375(.dina(n24632),.dinb(w_n21184_3[1]),.dout(n24633),.clk(gclk));
	jnot g24376(.din(w_n24127_0[1]),.dout(n24634),.clk(gclk));
	jor g24377(.dina(n24634),.dinb(n24633),.dout(n24635),.clk(gclk));
	jand g24378(.dina(n24635),.dinb(n24612),.dout(n24636),.clk(gclk));
	jand g24379(.dina(n24636),.dinb(w_n20468_12[2]),.dout(n24637),.clk(gclk));
	jor g24380(.dina(w_n24134_0[0]),.dinb(n24637),.dout(n24638),.clk(gclk));
	jand g24381(.dina(n24638),.dinb(n24611),.dout(n24639),.clk(gclk));
	jand g24382(.dina(n24639),.dinb(w_n19791_4[1]),.dout(n24640),.clk(gclk));
	jor g24383(.dina(w_n24142_0[0]),.dinb(n24640),.dout(n24641),.clk(gclk));
	jand g24384(.dina(n24641),.dinb(n24610),.dout(n24642),.clk(gclk));
	jand g24385(.dina(n24642),.dinb(w_n19096_13[0]),.dout(n24643),.clk(gclk));
	jnot g24386(.din(w_n24150_0[1]),.dout(n24644),.clk(gclk));
	jor g24387(.dina(n24644),.dinb(n24643),.dout(n24645),.clk(gclk));
	jand g24388(.dina(n24645),.dinb(n24609),.dout(n24646),.clk(gclk));
	jand g24389(.dina(n24646),.dinb(w_n18442_5[0]),.dout(n24647),.clk(gclk));
	jnot g24390(.din(w_n24157_0[1]),.dout(n24648),.clk(gclk));
	jor g24391(.dina(n24648),.dinb(n24647),.dout(n24649),.clk(gclk));
	jand g24392(.dina(n24649),.dinb(n24608),.dout(n24650),.clk(gclk));
	jand g24393(.dina(n24650),.dinb(w_n17769_13[2]),.dout(n24651),.clk(gclk));
	jnot g24394(.din(w_n24164_0[1]),.dout(n24652),.clk(gclk));
	jor g24395(.dina(n24652),.dinb(n24651),.dout(n24653),.clk(gclk));
	jand g24396(.dina(n24653),.dinb(n24607),.dout(n24654),.clk(gclk));
	jand g24397(.dina(n24654),.dinb(w_n17134_6[0]),.dout(n24655),.clk(gclk));
	jor g24398(.dina(w_n24171_0[0]),.dinb(n24655),.dout(n24656),.clk(gclk));
	jand g24399(.dina(n24656),.dinb(n24606),.dout(n24657),.clk(gclk));
	jand g24400(.dina(n24657),.dinb(w_n16489_14[0]),.dout(n24658),.clk(gclk));
	jnot g24401(.din(w_n24179_0[1]),.dout(n24659),.clk(gclk));
	jor g24402(.dina(n24659),.dinb(n24658),.dout(n24660),.clk(gclk));
	jand g24403(.dina(n24660),.dinb(n24605),.dout(n24661),.clk(gclk));
	jand g24404(.dina(n24661),.dinb(w_n15878_7[0]),.dout(n24662),.clk(gclk));
	jor g24405(.dina(w_n24186_0[0]),.dinb(n24662),.dout(n24663),.clk(gclk));
	jand g24406(.dina(n24663),.dinb(n24604),.dout(n24664),.clk(gclk));
	jand g24407(.dina(n24664),.dinb(w_n15260_14[2]),.dout(n24665),.clk(gclk));
	jnot g24408(.din(w_n24194_0[1]),.dout(n24666),.clk(gclk));
	jor g24409(.dina(n24666),.dinb(n24665),.dout(n24667),.clk(gclk));
	jand g24410(.dina(n24667),.dinb(n24603),.dout(n24668),.clk(gclk));
	jand g24411(.dina(n24668),.dinb(w_n14674_7[2]),.dout(n24669),.clk(gclk));
	jor g24412(.dina(w_n24201_0[0]),.dinb(n24669),.dout(n24670),.clk(gclk));
	jand g24413(.dina(n24670),.dinb(n24602),.dout(n24671),.clk(gclk));
	jand g24414(.dina(n24671),.dinb(w_n14078_15[0]),.dout(n24672),.clk(gclk));
	jor g24415(.dina(w_n24209_0[0]),.dinb(n24672),.dout(n24673),.clk(gclk));
	jand g24416(.dina(n24673),.dinb(n24601),.dout(n24674),.clk(gclk));
	jand g24417(.dina(n24674),.dinb(w_n13515_8[2]),.dout(n24675),.clk(gclk));
	jor g24418(.dina(w_n24217_0[0]),.dinb(n24675),.dout(n24676),.clk(gclk));
	jand g24419(.dina(n24676),.dinb(n24600),.dout(n24677),.clk(gclk));
	jand g24420(.dina(n24677),.dinb(w_n12947_15[2]),.dout(n24678),.clk(gclk));
	jnot g24421(.din(w_n24225_0[1]),.dout(n24679),.clk(gclk));
	jor g24422(.dina(n24679),.dinb(n24678),.dout(n24680),.clk(gclk));
	jand g24423(.dina(n24680),.dinb(n24599),.dout(n24681),.clk(gclk));
	jand g24424(.dina(n24681),.dinb(w_n12410_9[1]),.dout(n24682),.clk(gclk));
	jor g24425(.dina(w_n24232_0[0]),.dinb(n24682),.dout(n24683),.clk(gclk));
	jand g24426(.dina(n24683),.dinb(n24598),.dout(n24684),.clk(gclk));
	jand g24427(.dina(n24684),.dinb(w_n11858_16[0]),.dout(n24685),.clk(gclk));
	jor g24428(.dina(w_n24240_0[0]),.dinb(n24685),.dout(n24686),.clk(gclk));
	jand g24429(.dina(n24686),.dinb(n24597),.dout(n24687),.clk(gclk));
	jand g24430(.dina(n24687),.dinb(w_n11347_10[0]),.dout(n24688),.clk(gclk));
	jor g24431(.dina(w_n24248_0[0]),.dinb(n24688),.dout(n24689),.clk(gclk));
	jand g24432(.dina(n24689),.dinb(n24596),.dout(n24690),.clk(gclk));
	jand g24433(.dina(n24690),.dinb(w_n10824_16[2]),.dout(n24691),.clk(gclk));
	jnot g24434(.din(w_n24256_0[1]),.dout(n24692),.clk(gclk));
	jor g24435(.dina(n24692),.dinb(n24691),.dout(n24693),.clk(gclk));
	jand g24436(.dina(n24693),.dinb(n24595),.dout(n24694),.clk(gclk));
	jand g24437(.dina(n24694),.dinb(w_n10328_11[0]),.dout(n24695),.clk(gclk));
	jor g24438(.dina(w_n24263_0[0]),.dinb(n24695),.dout(n24696),.clk(gclk));
	jand g24439(.dina(n24696),.dinb(n24594),.dout(n24697),.clk(gclk));
	jand g24440(.dina(n24697),.dinb(w_n9832_17[1]),.dout(n24698),.clk(gclk));
	jnot g24441(.din(w_n24271_0[1]),.dout(n24699),.clk(gclk));
	jor g24442(.dina(n24699),.dinb(n24698),.dout(n24700),.clk(gclk));
	jand g24443(.dina(n24700),.dinb(n24593),.dout(n24701),.clk(gclk));
	jand g24444(.dina(n24701),.dinb(w_n9369_12[0]),.dout(n24702),.clk(gclk));
	jor g24445(.dina(w_n24278_0[0]),.dinb(n24702),.dout(n24703),.clk(gclk));
	jand g24446(.dina(n24703),.dinb(n24592),.dout(n24704),.clk(gclk));
	jand g24447(.dina(n24704),.dinb(w_n8890_17[2]),.dout(n24705),.clk(gclk));
	jnot g24448(.din(w_n24286_0[1]),.dout(n24706),.clk(gclk));
	jor g24449(.dina(n24706),.dinb(n24705),.dout(n24707),.clk(gclk));
	jand g24450(.dina(n24707),.dinb(n24591),.dout(n24708),.clk(gclk));
	jand g24451(.dina(n24708),.dinb(w_n8449_12[2]),.dout(n24709),.clk(gclk));
	jor g24452(.dina(w_n24293_0[0]),.dinb(n24709),.dout(n24710),.clk(gclk));
	jand g24453(.dina(n24710),.dinb(n24590),.dout(n24711),.clk(gclk));
	jand g24454(.dina(n24711),.dinb(w_n8003_18[1]),.dout(n24712),.clk(gclk));
	jor g24455(.dina(w_n24301_0[0]),.dinb(n24712),.dout(n24713),.clk(gclk));
	jand g24456(.dina(n24713),.dinb(n24589),.dout(n24714),.clk(gclk));
	jand g24457(.dina(n24714),.dinb(w_n7581_13[2]),.dout(n24715),.clk(gclk));
	jnot g24458(.din(w_n24309_0[1]),.dout(n24716),.clk(gclk));
	jor g24459(.dina(n24716),.dinb(n24715),.dout(n24717),.clk(gclk));
	jand g24460(.dina(n24717),.dinb(n24588),.dout(n24718),.clk(gclk));
	jand g24461(.dina(n24718),.dinb(w_n7154_18[2]),.dout(n24719),.clk(gclk));
	jnot g24462(.din(w_n24316_0[1]),.dout(n24720),.clk(gclk));
	jor g24463(.dina(n24720),.dinb(n24719),.dout(n24721),.clk(gclk));
	jand g24464(.dina(n24721),.dinb(n24587),.dout(n24722),.clk(gclk));
	jand g24465(.dina(n24722),.dinb(w_n6758_14[1]),.dout(n24723),.clk(gclk));
	jor g24466(.dina(w_n24323_0[0]),.dinb(n24723),.dout(n24724),.clk(gclk));
	jand g24467(.dina(n24724),.dinb(n24586),.dout(n24725),.clk(gclk));
	jand g24468(.dina(n24725),.dinb(w_n6357_19[0]),.dout(n24726),.clk(gclk));
	jnot g24469(.din(w_n24331_0[1]),.dout(n24727),.clk(gclk));
	jor g24470(.dina(n24727),.dinb(n24726),.dout(n24728),.clk(gclk));
	jand g24471(.dina(n24728),.dinb(n24585),.dout(n24729),.clk(gclk));
	jand g24472(.dina(n24729),.dinb(w_n5989_15[0]),.dout(n24730),.clk(gclk));
	jor g24473(.dina(w_n24338_0[0]),.dinb(n24730),.dout(n24731),.clk(gclk));
	jand g24474(.dina(n24731),.dinb(n24584),.dout(n24732),.clk(gclk));
	jand g24475(.dina(n24732),.dinb(w_n5606_19[1]),.dout(n24733),.clk(gclk));
	jnot g24476(.din(w_n24346_0[1]),.dout(n24734),.clk(gclk));
	jor g24477(.dina(n24734),.dinb(n24733),.dout(n24735),.clk(gclk));
	jand g24478(.dina(n24735),.dinb(n24583),.dout(n24736),.clk(gclk));
	jand g24479(.dina(n24736),.dinb(w_n5259_16[0]),.dout(n24737),.clk(gclk));
	jor g24480(.dina(w_n24353_0[0]),.dinb(n24737),.dout(n24738),.clk(gclk));
	jand g24481(.dina(n24738),.dinb(n24582),.dout(n24739),.clk(gclk));
	jand g24482(.dina(n24739),.dinb(w_n4902_20[0]),.dout(n24740),.clk(gclk));
	jor g24483(.dina(w_n24361_0[0]),.dinb(n24740),.dout(n24741),.clk(gclk));
	jand g24484(.dina(n24741),.dinb(n24581),.dout(n24742),.clk(gclk));
	jand g24485(.dina(n24742),.dinb(w_n4582_17[0]),.dout(n24743),.clk(gclk));
	jor g24486(.dina(w_n24369_0[0]),.dinb(n24743),.dout(n24744),.clk(gclk));
	jand g24487(.dina(n24744),.dinb(n24580),.dout(n24745),.clk(gclk));
	jand g24488(.dina(n24745),.dinb(w_n4249_20[2]),.dout(n24746),.clk(gclk));
	jnot g24489(.din(w_n24377_0[1]),.dout(n24747),.clk(gclk));
	jor g24490(.dina(n24747),.dinb(n24746),.dout(n24748),.clk(gclk));
	jand g24491(.dina(n24748),.dinb(n24579),.dout(n24749),.clk(gclk));
	jand g24492(.dina(n24749),.dinb(w_n3955_17[2]),.dout(n24750),.clk(gclk));
	jor g24493(.dina(w_n24384_0[0]),.dinb(n24750),.dout(n24751),.clk(gclk));
	jand g24494(.dina(n24751),.dinb(n24578),.dout(n24752),.clk(gclk));
	jand g24495(.dina(n24752),.dinb(w_n3642_21[0]),.dout(n24753),.clk(gclk));
	jnot g24496(.din(w_n24392_0[1]),.dout(n24754),.clk(gclk));
	jor g24497(.dina(n24754),.dinb(n24753),.dout(n24755),.clk(gclk));
	jand g24498(.dina(n24755),.dinb(n24577),.dout(n24756),.clk(gclk));
	jand g24499(.dina(n24756),.dinb(w_n3368_18[1]),.dout(n24757),.clk(gclk));
	jor g24500(.dina(w_n24399_0[0]),.dinb(n24757),.dout(n24758),.clk(gclk));
	jand g24501(.dina(n24758),.dinb(n24576),.dout(n24759),.clk(gclk));
	jand g24502(.dina(n24759),.dinb(w_n3089_21[2]),.dout(n24760),.clk(gclk));
	jnot g24503(.din(w_n24407_0[1]),.dout(n24761),.clk(gclk));
	jor g24504(.dina(n24761),.dinb(n24760),.dout(n24762),.clk(gclk));
	jand g24505(.dina(n24762),.dinb(n24575),.dout(n24763),.clk(gclk));
	jand g24506(.dina(n24763),.dinb(w_n2833_19[1]),.dout(n24764),.clk(gclk));
	jor g24507(.dina(w_n24414_0[0]),.dinb(n24764),.dout(n24765),.clk(gclk));
	jand g24508(.dina(n24765),.dinb(n24574),.dout(n24766),.clk(gclk));
	jand g24509(.dina(n24766),.dinb(w_n2572_22[0]),.dout(n24767),.clk(gclk));
	jnot g24510(.din(w_n24422_0[1]),.dout(n24768),.clk(gclk));
	jor g24511(.dina(n24768),.dinb(n24767),.dout(n24769),.clk(gclk));
	jand g24512(.dina(n24769),.dinb(n24573),.dout(n24770),.clk(gclk));
	jand g24513(.dina(n24770),.dinb(w_n2345_20[0]),.dout(n24771),.clk(gclk));
	jor g24514(.dina(w_n24429_0[0]),.dinb(n24771),.dout(n24772),.clk(gclk));
	jand g24515(.dina(n24772),.dinb(n24572),.dout(n24773),.clk(gclk));
	jand g24516(.dina(n24773),.dinb(w_n2108_22[2]),.dout(n24774),.clk(gclk));
	jor g24517(.dina(w_n24437_0[0]),.dinb(n24774),.dout(n24775),.clk(gclk));
	jand g24518(.dina(n24775),.dinb(n24571),.dout(n24776),.clk(gclk));
	jand g24519(.dina(n24776),.dinb(w_n1912_21[0]),.dout(n24777),.clk(gclk));
	jor g24520(.dina(w_n24445_0[0]),.dinb(n24777),.dout(n24778),.clk(gclk));
	jand g24521(.dina(n24778),.dinb(n24570),.dout(n24779),.clk(gclk));
	jand g24522(.dina(n24779),.dinb(w_n1699_23[1]),.dout(n24780),.clk(gclk));
	jnot g24523(.din(w_n24453_0[1]),.dout(n24781),.clk(gclk));
	jor g24524(.dina(n24781),.dinb(n24780),.dout(n24782),.clk(gclk));
	jand g24525(.dina(n24782),.dinb(n24569),.dout(n24783),.clk(gclk));
	jand g24526(.dina(n24783),.dinb(w_n1516_21[2]),.dout(n24784),.clk(gclk));
	jor g24527(.dina(w_n24460_0[0]),.dinb(n24784),.dout(n24785),.clk(gclk));
	jand g24528(.dina(n24785),.dinb(n24568),.dout(n24786),.clk(gclk));
	jand g24529(.dina(n24786),.dinb(w_n1332_23[1]),.dout(n24787),.clk(gclk));
	jor g24530(.dina(w_n24468_0[0]),.dinb(n24787),.dout(n24788),.clk(gclk));
	jand g24531(.dina(n24788),.dinb(n24567),.dout(n24789),.clk(gclk));
	jand g24532(.dina(n24789),.dinb(w_n1173_22[1]),.dout(n24790),.clk(gclk));
	jor g24533(.dina(w_n24476_0[0]),.dinb(n24790),.dout(n24791),.clk(gclk));
	jand g24534(.dina(n24791),.dinb(n24566),.dout(n24792),.clk(gclk));
	jand g24535(.dina(n24792),.dinb(w_n1008_24[1]),.dout(n24793),.clk(gclk));
	jor g24536(.dina(w_n24484_0[0]),.dinb(n24793),.dout(n24794),.clk(gclk));
	jand g24537(.dina(n24794),.dinb(n24565),.dout(n24795),.clk(gclk));
	jand g24538(.dina(n24795),.dinb(w_n884_23[1]),.dout(n24796),.clk(gclk));
	jor g24539(.dina(w_n24492_0[0]),.dinb(n24796),.dout(n24797),.clk(gclk));
	jand g24540(.dina(n24797),.dinb(n24564),.dout(n24798),.clk(gclk));
	jand g24541(.dina(n24798),.dinb(w_n743_24[1]),.dout(n24799),.clk(gclk));
	jnot g24542(.din(w_n24500_0[1]),.dout(n24800),.clk(gclk));
	jor g24543(.dina(n24800),.dinb(n24799),.dout(n24801),.clk(gclk));
	jand g24544(.dina(n24801),.dinb(n24563),.dout(n24802),.clk(gclk));
	jand g24545(.dina(n24802),.dinb(w_n635_24[1]),.dout(n24803),.clk(gclk));
	jor g24546(.dina(w_n24507_0[0]),.dinb(n24803),.dout(n24804),.clk(gclk));
	jand g24547(.dina(n24804),.dinb(n24562),.dout(n24805),.clk(gclk));
	jand g24548(.dina(n24805),.dinb(w_n515_25[1]),.dout(n24806),.clk(gclk));
	jnot g24549(.din(w_n24515_0[1]),.dout(n24807),.clk(gclk));
	jor g24550(.dina(n24807),.dinb(n24806),.dout(n24808),.clk(gclk));
	jand g24551(.dina(n24808),.dinb(n24561),.dout(n24809),.clk(gclk));
	jand g24552(.dina(n24809),.dinb(w_n443_25[1]),.dout(n24810),.clk(gclk));
	jor g24553(.dina(w_n24522_0[0]),.dinb(n24810),.dout(n24811),.clk(gclk));
	jand g24554(.dina(n24811),.dinb(n24560),.dout(n24812),.clk(gclk));
	jand g24555(.dina(n24812),.dinb(w_n352_25[2]),.dout(n24813),.clk(gclk));
	jnot g24556(.din(w_n24530_0[1]),.dout(n24814),.clk(gclk));
	jor g24557(.dina(n24814),.dinb(n24813),.dout(n24815),.clk(gclk));
	jand g24558(.dina(n24815),.dinb(n24559),.dout(n24816),.clk(gclk));
	jand g24559(.dina(n24816),.dinb(w_n294_26[0]),.dout(n24817),.clk(gclk));
	jnot g24560(.din(w_n24537_0[1]),.dout(n24818),.clk(gclk));
	jor g24561(.dina(n24818),.dinb(n24817),.dout(n24819),.clk(gclk));
	jand g24562(.dina(n24819),.dinb(n24558),.dout(n24820),.clk(gclk));
	jand g24563(.dina(n24820),.dinb(w_n239_26[0]),.dout(n24821),.clk(gclk));
	jnot g24564(.din(w_n24544_0[1]),.dout(n24822),.clk(gclk));
	jor g24565(.dina(n24822),.dinb(n24821),.dout(n24823),.clk(gclk));
	jand g24566(.dina(n24823),.dinb(n24557),.dout(n24824),.clk(gclk));
	jand g24567(.dina(n24824),.dinb(w_n221_26[2]),.dout(n24825),.clk(gclk));
	jor g24568(.dina(w_n24551_0[0]),.dinb(n24825),.dout(n24826),.clk(gclk));
	jand g24569(.dina(n24826),.dinb(n24556),.dout(n24827),.clk(gclk));
	jxor g24570(.dina(w_n23787_0[0]),.dinb(w_n221_26[1]),.dout(n24828),.clk(gclk));
	jand g24571(.dina(n24828),.dinb(w_asqrt2_10[2]),.dout(n24829),.clk(gclk));
	jxor g24572(.dina(n24829),.dinb(w_n23792_0[0]),.dout(n24830),.clk(gclk));
	jor g24573(.dina(w_n24830_0[1]),.dinb(n24827),.dout(n24831),.clk(gclk));
	jor g24574(.dina(w_n24831_0[1]),.dinb(w_n23795_0[0]),.dout(n24832),.clk(gclk));
	jor g24575(.dina(n24832),.dinb(w_n24555_0[1]),.dout(n24833),.clk(gclk));
	jnot g24576(.din(w_n24830_0[0]),.dout(n24834),.clk(gclk));
	jor g24577(.dina(w_n24834_0[1]),.dinb(w_n24554_0[2]),.dout(n24835),.clk(gclk));
	jand g24578(.dina(w_n24835_0[2]),.dinb(w_n218_11[0]),.dout(n24836),.clk(gclk));
	jnot g24579(.din(w_n24836_0[1]),.dout(n24837),.clk(gclk));
	jor g24580(.dina(n24837),.dinb(n24833),.dout(n24838),.clk(gclk));
	jand g24581(.dina(w_n24835_0[1]),.dinb(w_asqrt63_19[0]),.dout(n24839),.clk(gclk));
	jand g24582(.dina(w_n24102_0[0]),.dinb(w_n23794_0[2]),.dout(n24840),.clk(gclk));
	jnot g24583(.din(n24840),.dout(n24841),.clk(gclk));
	jxor g24584(.dina(w_n23794_0[1]),.dinb(w_n23349_0[0]),.dout(n24842),.clk(gclk));
	jand g24585(.dina(n24842),.dinb(n24841),.dout(n24843),.clk(gclk));
	jnot g24586(.din(n24843),.dout(n24844),.clk(gclk));
	jand g24587(.dina(n24844),.dinb(w_n24839_0[1]),.dout(n24845),.clk(gclk));
	jnot g24588(.din(w_n24845_0[1]),.dout(n24846),.clk(gclk));
	jand g24589(.dina(n24846),.dinb(n24838),.dout(asqrt_fa_2),.clk(gclk));
	jor g24590(.dina(w_asqrt1_1),.dinb(w_n24554_0[1]),.dout(n24848),.clk(gclk));
	jand g24591(.dina(w_n24839_0[0]),.dinb(w_n24831_0[0]),.dout(n24849),.clk(gclk));
	jand g24592(.dina(n24849),.dinb(n24848),.dout(n24850),.clk(gclk));
	jnot g24593(.din(w_n24555_0[0]),.dout(n24851),.clk(gclk));
	jand g24594(.dina(w_n24834_0[0]),.dinb(w_n24554_0[0]),.dout(n24852),.clk(gclk));
	jand g24595(.dina(w_n24852_0[1]),.dinb(w_n23818_0[0]),.dout(n24853),.clk(gclk));
	jand g24596(.dina(n24853),.dinb(n24851),.dout(n24854),.clk(gclk));
	jand g24597(.dina(w_n24836_0[0]),.dinb(n24854),.dout(n24855),.clk(gclk));
	jor g24598(.dina(w_n24845_0[0]),.dinb(n24855),.dout(n24856),.clk(gclk));
	jxor g24599(.dina(w_n24539_0[0]),.dinb(w_n239_25[2]),.dout(n24857),.clk(gclk));
	jor g24600(.dina(n24857),.dinb(w_n24856_30[2]),.dout(n24858),.clk(gclk));
	jxor g24601(.dina(n24858),.dinb(w_n24544_0[0]),.dout(n24859),.clk(gclk));
	jand g24602(.dina(w_n24859_0[1]),.dinb(w_n221_26[0]),.dout(n24860),.clk(gclk));
	jxor g24603(.dina(w_n24487_0[0]),.dinb(w_n884_23[0]),.dout(n24861),.clk(gclk));
	jor g24604(.dina(n24861),.dinb(w_n24856_30[1]),.dout(n24862),.clk(gclk));
	jxor g24605(.dina(n24862),.dinb(w_n24493_0[0]),.dout(n24863),.clk(gclk));
	jor g24606(.dina(w_n24863_0[1]),.dinb(w_n743_24[0]),.dout(n24864),.clk(gclk));
	jxor g24607(.dina(w_n24479_0[0]),.dinb(w_n1008_24[0]),.dout(n24865),.clk(gclk));
	jor g24608(.dina(n24865),.dinb(w_n24856_30[0]),.dout(n24866),.clk(gclk));
	jxor g24609(.dina(n24866),.dinb(w_n24485_0[0]),.dout(n24867),.clk(gclk));
	jand g24610(.dina(w_n24867_0[1]),.dinb(w_n884_22[2]),.dout(n24868),.clk(gclk));
	jand g24611(.dina(w_n24863_0[0]),.dinb(w_n743_23[2]),.dout(n24869),.clk(gclk));
	jor g24612(.dina(n24869),.dinb(n24868),.dout(n24870),.clk(gclk));
	jxor g24613(.dina(w_n24463_0[0]),.dinb(w_n1332_23[0]),.dout(n24871),.clk(gclk));
	jor g24614(.dina(n24871),.dinb(w_n24856_29[2]),.dout(n24872),.clk(gclk));
	jxor g24615(.dina(n24872),.dinb(w_n24469_0[0]),.dout(n24873),.clk(gclk));
	jand g24616(.dina(w_n24873_0[1]),.dinb(w_n1173_22[0]),.dout(n24874),.clk(gclk));
	jxor g24617(.dina(w_n24455_0[0]),.dinb(w_n1516_21[1]),.dout(n24875),.clk(gclk));
	jor g24618(.dina(n24875),.dinb(w_n24856_29[1]),.dout(n24876),.clk(gclk));
	jxor g24619(.dina(n24876),.dinb(w_n24461_0[0]),.dout(n24877),.clk(gclk));
	jand g24620(.dina(w_n24877_0[1]),.dinb(w_n1332_22[2]),.dout(n24878),.clk(gclk));
	jxor g24621(.dina(w_n24424_0[0]),.dinb(w_n2345_19[2]),.dout(n24879),.clk(gclk));
	jor g24622(.dina(n24879),.dinb(w_n24856_29[0]),.dout(n24880),.clk(gclk));
	jxor g24623(.dina(n24880),.dinb(w_n24430_0[0]),.dout(n24881),.clk(gclk));
	jor g24624(.dina(w_n24881_0[1]),.dinb(w_n2108_22[1]),.dout(n24882),.clk(gclk));
	jxor g24625(.dina(w_n24417_0[0]),.dinb(w_n2572_21[2]),.dout(n24883),.clk(gclk));
	jor g24626(.dina(n24883),.dinb(w_n24856_28[2]),.dout(n24884),.clk(gclk));
	jxor g24627(.dina(n24884),.dinb(w_n24422_0[0]),.dout(n24885),.clk(gclk));
	jand g24628(.dina(w_n24885_0[1]),.dinb(w_n2345_19[1]),.dout(n24886),.clk(gclk));
	jxor g24629(.dina(w_n24394_0[0]),.dinb(w_n3368_18[0]),.dout(n24887),.clk(gclk));
	jor g24630(.dina(n24887),.dinb(w_n24856_28[1]),.dout(n24888),.clk(gclk));
	jxor g24631(.dina(n24888),.dinb(w_n24400_0[0]),.dout(n24889),.clk(gclk));
	jand g24632(.dina(w_n24889_0[1]),.dinb(w_n3089_21[1]),.dout(n24890),.clk(gclk));
	jxor g24633(.dina(w_n24364_0[0]),.dinb(w_n4582_16[2]),.dout(n24891),.clk(gclk));
	jor g24634(.dina(n24891),.dinb(w_n24856_28[0]),.dout(n24892),.clk(gclk));
	jxor g24635(.dina(n24892),.dinb(w_n24370_0[0]),.dout(n24893),.clk(gclk));
	jor g24636(.dina(w_n24893_0[1]),.dinb(w_n4249_20[1]),.dout(n24894),.clk(gclk));
	jxor g24637(.dina(w_n24356_0[0]),.dinb(w_n4902_19[2]),.dout(n24895),.clk(gclk));
	jor g24638(.dina(n24895),.dinb(w_n24856_27[2]),.dout(n24896),.clk(gclk));
	jxor g24639(.dina(n24896),.dinb(w_n24362_0[0]),.dout(n24897),.clk(gclk));
	jand g24640(.dina(w_n24897_0[1]),.dinb(w_n4582_16[1]),.dout(n24898),.clk(gclk));
	jxor g24641(.dina(w_n24318_0[0]),.dinb(w_n6758_14[0]),.dout(n24899),.clk(gclk));
	jor g24642(.dina(n24899),.dinb(w_n24856_27[1]),.dout(n24900),.clk(gclk));
	jxor g24643(.dina(n24900),.dinb(w_n24324_0[0]),.dout(n24901),.clk(gclk));
	jor g24644(.dina(w_n24901_0[1]),.dinb(w_n6357_18[2]),.dout(n24902),.clk(gclk));
	jxor g24645(.dina(w_n24296_0[0]),.dinb(w_n8003_18[0]),.dout(n24903),.clk(gclk));
	jor g24646(.dina(n24903),.dinb(w_n24856_27[0]),.dout(n24904),.clk(gclk));
	jxor g24647(.dina(n24904),.dinb(w_n24302_0[0]),.dout(n24905),.clk(gclk));
	jand g24648(.dina(w_n24905_0[1]),.dinb(w_n7581_13[1]),.dout(n24906),.clk(gclk));
	jxor g24649(.dina(w_n24288_0[0]),.dinb(w_n8449_12[1]),.dout(n24907),.clk(gclk));
	jor g24650(.dina(n24907),.dinb(w_n24856_26[2]),.dout(n24908),.clk(gclk));
	jxor g24651(.dina(n24908),.dinb(w_n24294_0[0]),.dout(n24909),.clk(gclk));
	jand g24652(.dina(w_n24909_0[1]),.dinb(w_n8003_17[2]),.dout(n24910),.clk(gclk));
	jxor g24653(.dina(w_n24281_0[0]),.dinb(w_n8890_17[1]),.dout(n24911),.clk(gclk));
	jor g24654(.dina(n24911),.dinb(w_n24856_26[1]),.dout(n24912),.clk(gclk));
	jxor g24655(.dina(n24912),.dinb(w_n24286_0[0]),.dout(n24913),.clk(gclk));
	jor g24656(.dina(w_n24913_0[1]),.dinb(w_n8449_12[0]),.dout(n24914),.clk(gclk));
	jxor g24657(.dina(w_n24251_0[0]),.dinb(w_n10824_16[1]),.dout(n24915),.clk(gclk));
	jor g24658(.dina(n24915),.dinb(w_n24856_26[0]),.dout(n24916),.clk(gclk));
	jxor g24659(.dina(n24916),.dinb(w_n24256_0[0]),.dout(n24917),.clk(gclk));
	jand g24660(.dina(w_n24917_0[1]),.dinb(w_n10328_10[2]),.dout(n24918),.clk(gclk));
	jxor g24661(.dina(w_n24243_0[0]),.dinb(w_n11347_9[2]),.dout(n24919),.clk(gclk));
	jor g24662(.dina(n24919),.dinb(w_n24856_25[2]),.dout(n24920),.clk(gclk));
	jxor g24663(.dina(n24920),.dinb(w_n24249_0[0]),.dout(n24921),.clk(gclk));
	jand g24664(.dina(w_n24921_0[1]),.dinb(w_n10824_16[0]),.dout(n24922),.clk(gclk));
	jxor g24665(.dina(w_n24227_0[0]),.dinb(w_n12410_9[0]),.dout(n24923),.clk(gclk));
	jor g24666(.dina(n24923),.dinb(w_n24856_25[1]),.dout(n24924),.clk(gclk));
	jxor g24667(.dina(n24924),.dinb(w_n24233_0[0]),.dout(n24925),.clk(gclk));
	jor g24668(.dina(w_n24925_0[1]),.dinb(w_n11858_15[2]),.dout(n24926),.clk(gclk));
	jxor g24669(.dina(w_n24220_0[0]),.dinb(w_n12947_15[1]),.dout(n24927),.clk(gclk));
	jor g24670(.dina(n24927),.dinb(w_n24856_25[0]),.dout(n24928),.clk(gclk));
	jxor g24671(.dina(n24928),.dinb(w_n24225_0[0]),.dout(n24929),.clk(gclk));
	jand g24672(.dina(w_n24929_0[1]),.dinb(w_n12410_8[2]),.dout(n24930),.clk(gclk));
	jxor g24673(.dina(w_n24196_0[0]),.dinb(w_n14674_7[1]),.dout(n24931),.clk(gclk));
	jor g24674(.dina(n24931),.dinb(w_n24856_24[2]),.dout(n24932),.clk(gclk));
	jxor g24675(.dina(n24932),.dinb(w_n24202_0[0]),.dout(n24933),.clk(gclk));
	jor g24676(.dina(w_n24933_0[1]),.dinb(w_n14078_14[2]),.dout(n24934),.clk(gclk));
	jxor g24677(.dina(w_n24189_0[0]),.dinb(w_n15260_14[1]),.dout(n24935),.clk(gclk));
	jor g24678(.dina(n24935),.dinb(w_n24856_24[1]),.dout(n24936),.clk(gclk));
	jxor g24679(.dina(n24936),.dinb(w_n24194_0[0]),.dout(n24937),.clk(gclk));
	jor g24680(.dina(w_n24937_0[1]),.dinb(w_n14674_7[0]),.dout(n24938),.clk(gclk));
	jxor g24681(.dina(w_n24174_0[0]),.dinb(w_n16489_13[2]),.dout(n24939),.clk(gclk));
	jor g24682(.dina(n24939),.dinb(w_n24856_24[0]),.dout(n24940),.clk(gclk));
	jxor g24683(.dina(n24940),.dinb(w_n24179_0[0]),.dout(n24941),.clk(gclk));
	jor g24684(.dina(w_n24941_0[1]),.dinb(w_n15878_6[2]),.dout(n24942),.clk(gclk));
	jxor g24685(.dina(w_n24166_0[0]),.dinb(w_n17134_5[2]),.dout(n24943),.clk(gclk));
	jor g24686(.dina(n24943),.dinb(w_n24856_23[2]),.dout(n24944),.clk(gclk));
	jxor g24687(.dina(n24944),.dinb(w_n24172_0[0]),.dout(n24945),.clk(gclk));
	jor g24688(.dina(w_n24945_0[1]),.dinb(w_n16489_13[1]),.dout(n24946),.clk(gclk));
	jxor g24689(.dina(w_n24159_0[0]),.dinb(w_n17769_13[1]),.dout(n24947),.clk(gclk));
	jor g24690(.dina(n24947),.dinb(w_n24856_23[1]),.dout(n24948),.clk(gclk));
	jxor g24691(.dina(n24948),.dinb(w_n24164_0[0]),.dout(n24949),.clk(gclk));
	jand g24692(.dina(w_n24949_0[1]),.dinb(w_n17134_5[1]),.dout(n24950),.clk(gclk));
	jxor g24693(.dina(w_n24137_0[0]),.dinb(w_n19791_4[0]),.dout(n24951),.clk(gclk));
	jor g24694(.dina(n24951),.dinb(w_n24856_23[0]),.dout(n24952),.clk(gclk));
	jxor g24695(.dina(n24952),.dinb(w_n24143_0[0]),.dout(n24953),.clk(gclk));
	jor g24696(.dina(w_n24953_0[1]),.dinb(w_n19096_12[2]),.dout(n24954),.clk(gclk));
	jand g24697(.dina(w_n24953_0[0]),.dinb(w_n19096_12[1]),.dout(n24955),.clk(gclk));
	jxor g24698(.dina(w_n24129_0[0]),.dinb(w_n20468_12[1]),.dout(n24956),.clk(gclk));
	jor g24699(.dina(n24956),.dinb(w_n24856_22[2]),.dout(n24957),.clk(gclk));
	jxor g24700(.dina(n24957),.dinb(w_n24135_0[0]),.dout(n24958),.clk(gclk));
	jor g24701(.dina(w_n24958_0[1]),.dinb(w_n19791_3[2]),.dout(n24959),.clk(gclk));
	jxor g24702(.dina(w_n24122_0[0]),.dinb(w_n21184_3[0]),.dout(n24960),.clk(gclk));
	jor g24703(.dina(n24960),.dinb(w_n24856_22[1]),.dout(n24961),.clk(gclk));
	jxor g24704(.dina(n24961),.dinb(w_n24127_0[0]),.dout(n24962),.clk(gclk));
	jor g24705(.dina(w_n24962_0[1]),.dinb(w_n20468_12[0]),.dout(n24963),.clk(gclk));
	jxor g24706(.dina(w_n24115_0[0]),.dinb(w_n21887_12[0]),.dout(n24964),.clk(gclk));
	jor g24707(.dina(n24964),.dinb(w_n24856_22[0]),.dout(n24965),.clk(gclk));
	jxor g24708(.dina(n24965),.dinb(w_n24120_0[0]),.dout(n24966),.clk(gclk));
	jor g24709(.dina(w_n24966_0[1]),.dinb(w_n21184_2[2]),.dout(n24967),.clk(gclk));
	jand g24710(.dina(w_asqrt1_0[2]),.dinb(w_n23810_0[0]),.dout(n24968),.clk(gclk));
	jand g24711(.dina(w_n24856_21[2]),.dinb(w_asqrt2_10[1]),.dout(n24969),.clk(gclk));
	jor g24712(.dina(n24969),.dinb(w_n24968_0[1]),.dout(n24970),.clk(gclk));
	jxor g24713(.dina(n24970),.dinb(w_a4_0[1]),.dout(n24971),.clk(gclk));
	jor g24714(.dina(w_n24971_0[1]),.dinb(w_n23345_11[1]),.dout(n24972),.clk(gclk));
	jnot g24715(.din(w_a2_1[0]),.dout(n24973),.clk(gclk));
	jor g24716(.dina(a[1]),.dinb(a[0]),.dout(n24974),.clk(gclk));
	jand g24717(.dina(n24974),.dinb(n24973),.dout(n24975),.clk(gclk));
	jand g24718(.dina(w_n24856_21[1]),.dinb(w_a2_0[2]),.dout(n24976),.clk(gclk));
	jor g24719(.dina(n24976),.dinb(n24975),.dout(n24977),.clk(gclk));
	jor g24720(.dina(w_n24977_0[1]),.dinb(w_n24103_0[2]),.dout(n24978),.clk(gclk));
	jand g24721(.dina(w_n24977_0[0]),.dinb(w_n24103_0[1]),.dout(n24979),.clk(gclk));
	jor g24722(.dina(w_n24856_21[0]),.dinb(w_a2_0[1]),.dout(n24980),.clk(gclk));
	jand g24723(.dina(n24980),.dinb(w_a3_0[0]),.dout(n24981),.clk(gclk));
	jor g24724(.dina(n24981),.dinb(w_n24968_0[0]),.dout(n24982),.clk(gclk));
	jor g24725(.dina(n24982),.dinb(n24979),.dout(n24983),.clk(gclk));
	jand g24726(.dina(n24983),.dinb(n24978),.dout(n24984),.clk(gclk));
	jand g24727(.dina(n24984),.dinb(n24972),.dout(n24985),.clk(gclk));
	jxor g24728(.dina(w_n23812_0[0]),.dinb(w_n23345_11[0]),.dout(n24986),.clk(gclk));
	jor g24729(.dina(n24986),.dinb(w_n24856_20[2]),.dout(n24987),.clk(gclk));
	jxor g24730(.dina(n24987),.dinb(w_n24105_0[0]),.dout(n24988),.clk(gclk));
	jand g24731(.dina(w_n24988_0[1]),.dinb(w_n22620_2[0]),.dout(n24989),.clk(gclk));
	jand g24732(.dina(w_n24971_0[0]),.dinb(w_n23345_10[2]),.dout(n24990),.clk(gclk));
	jor g24733(.dina(n24990),.dinb(n24989),.dout(n24991),.clk(gclk));
	jor g24734(.dina(n24991),.dinb(n24985),.dout(n24992),.clk(gclk));
	jxor g24735(.dina(w_n24107_0[0]),.dinb(w_n22620_1[2]),.dout(n24993),.clk(gclk));
	jor g24736(.dina(n24993),.dinb(w_n24856_20[1]),.dout(n24994),.clk(gclk));
	jxor g24737(.dina(n24994),.dinb(w_n24113_0[0]),.dout(n24995),.clk(gclk));
	jor g24738(.dina(w_n24995_0[1]),.dinb(w_n21887_11[2]),.dout(n24996),.clk(gclk));
	jor g24739(.dina(w_n24988_0[0]),.dinb(w_n22620_1[1]),.dout(n24997),.clk(gclk));
	jand g24740(.dina(n24997),.dinb(n24996),.dout(n24998),.clk(gclk));
	jand g24741(.dina(n24998),.dinb(n24992),.dout(n24999),.clk(gclk));
	jand g24742(.dina(w_n24966_0[0]),.dinb(w_n21184_2[1]),.dout(n25000),.clk(gclk));
	jand g24743(.dina(w_n24995_0[0]),.dinb(w_n21887_11[1]),.dout(n25001),.clk(gclk));
	jor g24744(.dina(n25001),.dinb(n25000),.dout(n25002),.clk(gclk));
	jor g24745(.dina(n25002),.dinb(n24999),.dout(n25003),.clk(gclk));
	jand g24746(.dina(n25003),.dinb(n24967),.dout(n25004),.clk(gclk));
	jand g24747(.dina(n25004),.dinb(n24963),.dout(n25005),.clk(gclk));
	jand g24748(.dina(w_n24962_0[0]),.dinb(w_n20468_11[2]),.dout(n25006),.clk(gclk));
	jand g24749(.dina(w_n24958_0[0]),.dinb(w_n19791_3[1]),.dout(n25007),.clk(gclk));
	jor g24750(.dina(n25007),.dinb(n25006),.dout(n25008),.clk(gclk));
	jor g24751(.dina(n25008),.dinb(n25005),.dout(n25009),.clk(gclk));
	jand g24752(.dina(n25009),.dinb(n24959),.dout(n25010),.clk(gclk));
	jor g24753(.dina(n25010),.dinb(n24955),.dout(n25011),.clk(gclk));
	jxor g24754(.dina(w_n24145_0[0]),.dinb(w_n19096_12[0]),.dout(n25012),.clk(gclk));
	jor g24755(.dina(n25012),.dinb(w_n24856_20[0]),.dout(n25013),.clk(gclk));
	jxor g24756(.dina(n25013),.dinb(w_n24150_0[0]),.dout(n25014),.clk(gclk));
	jor g24757(.dina(w_n25014_0[1]),.dinb(w_n18442_4[2]),.dout(n25015),.clk(gclk));
	jand g24758(.dina(n25015),.dinb(n25011),.dout(n25016),.clk(gclk));
	jand g24759(.dina(n25016),.dinb(n24954),.dout(n25017),.clk(gclk));
	jand g24760(.dina(w_n25014_0[0]),.dinb(w_n18442_4[1]),.dout(n25018),.clk(gclk));
	jxor g24761(.dina(w_n24152_0[0]),.dinb(w_n18442_4[0]),.dout(n25019),.clk(gclk));
	jor g24762(.dina(n25019),.dinb(w_n24856_19[2]),.dout(n25020),.clk(gclk));
	jxor g24763(.dina(n25020),.dinb(w_n24157_0[0]),.dout(n25021),.clk(gclk));
	jand g24764(.dina(w_n25021_0[1]),.dinb(w_n17769_13[0]),.dout(n25022),.clk(gclk));
	jor g24765(.dina(n25022),.dinb(n25018),.dout(n25023),.clk(gclk));
	jor g24766(.dina(n25023),.dinb(n25017),.dout(n25024),.clk(gclk));
	jor g24767(.dina(w_n25021_0[0]),.dinb(w_n17769_12[2]),.dout(n25025),.clk(gclk));
	jor g24768(.dina(w_n24949_0[0]),.dinb(w_n17134_5[0]),.dout(n25026),.clk(gclk));
	jand g24769(.dina(n25026),.dinb(n25025),.dout(n25027),.clk(gclk));
	jand g24770(.dina(n25027),.dinb(n25024),.dout(n25028),.clk(gclk));
	jor g24771(.dina(n25028),.dinb(n24950),.dout(n25029),.clk(gclk));
	jand g24772(.dina(n25029),.dinb(n24946),.dout(n25030),.clk(gclk));
	jand g24773(.dina(w_n24945_0[0]),.dinb(w_n16489_13[0]),.dout(n25031),.clk(gclk));
	jand g24774(.dina(w_n24941_0[0]),.dinb(w_n15878_6[1]),.dout(n25032),.clk(gclk));
	jor g24775(.dina(n25032),.dinb(n25031),.dout(n25033),.clk(gclk));
	jor g24776(.dina(n25033),.dinb(n25030),.dout(n25034),.clk(gclk));
	jxor g24777(.dina(w_n24181_0[0]),.dinb(w_n15878_6[0]),.dout(n25035),.clk(gclk));
	jor g24778(.dina(n25035),.dinb(w_n24856_19[1]),.dout(n25036),.clk(gclk));
	jxor g24779(.dina(n25036),.dinb(w_n24187_0[0]),.dout(n25037),.clk(gclk));
	jor g24780(.dina(w_n25037_0[1]),.dinb(w_n15260_14[0]),.dout(n25038),.clk(gclk));
	jand g24781(.dina(n25038),.dinb(n25034),.dout(n25039),.clk(gclk));
	jand g24782(.dina(n25039),.dinb(n24942),.dout(n25040),.clk(gclk));
	jand g24783(.dina(w_n25037_0[0]),.dinb(w_n15260_13[2]),.dout(n25041),.clk(gclk));
	jand g24784(.dina(w_n24937_0[0]),.dinb(w_n14674_6[2]),.dout(n25042),.clk(gclk));
	jor g24785(.dina(n25042),.dinb(n25041),.dout(n25043),.clk(gclk));
	jor g24786(.dina(n25043),.dinb(n25040),.dout(n25044),.clk(gclk));
	jand g24787(.dina(n25044),.dinb(n24938),.dout(n25045),.clk(gclk));
	jand g24788(.dina(w_n24933_0[0]),.dinb(w_n14078_14[1]),.dout(n25046),.clk(gclk));
	jor g24789(.dina(n25046),.dinb(n25045),.dout(n25047),.clk(gclk));
	jxor g24790(.dina(w_n24204_0[0]),.dinb(w_n14078_14[0]),.dout(n25048),.clk(gclk));
	jor g24791(.dina(n25048),.dinb(w_n24856_19[0]),.dout(n25049),.clk(gclk));
	jxor g24792(.dina(n25049),.dinb(w_n24210_0[0]),.dout(n25050),.clk(gclk));
	jor g24793(.dina(w_n25050_0[1]),.dinb(w_n13515_8[1]),.dout(n25051),.clk(gclk));
	jand g24794(.dina(n25051),.dinb(n25047),.dout(n25052),.clk(gclk));
	jand g24795(.dina(n25052),.dinb(n24934),.dout(n25053),.clk(gclk));
	jand g24796(.dina(w_n25050_0[0]),.dinb(w_n13515_8[0]),.dout(n25054),.clk(gclk));
	jxor g24797(.dina(w_n24212_0[0]),.dinb(w_n13515_7[2]),.dout(n25055),.clk(gclk));
	jor g24798(.dina(n25055),.dinb(w_n24856_18[2]),.dout(n25056),.clk(gclk));
	jxor g24799(.dina(n25056),.dinb(w_n24218_0[0]),.dout(n25057),.clk(gclk));
	jand g24800(.dina(w_n25057_0[1]),.dinb(w_n12947_15[0]),.dout(n25058),.clk(gclk));
	jor g24801(.dina(n25058),.dinb(n25054),.dout(n25059),.clk(gclk));
	jor g24802(.dina(n25059),.dinb(n25053),.dout(n25060),.clk(gclk));
	jor g24803(.dina(w_n24929_0[0]),.dinb(w_n12410_8[1]),.dout(n25061),.clk(gclk));
	jor g24804(.dina(w_n25057_0[0]),.dinb(w_n12947_14[2]),.dout(n25062),.clk(gclk));
	jand g24805(.dina(n25062),.dinb(n25061),.dout(n25063),.clk(gclk));
	jand g24806(.dina(n25063),.dinb(n25060),.dout(n25064),.clk(gclk));
	jor g24807(.dina(n25064),.dinb(n24930),.dout(n25065),.clk(gclk));
	jand g24808(.dina(n25065),.dinb(n24926),.dout(n25066),.clk(gclk));
	jand g24809(.dina(w_n24925_0[0]),.dinb(w_n11858_15[1]),.dout(n25067),.clk(gclk));
	jxor g24810(.dina(w_n24235_0[0]),.dinb(w_n11858_15[0]),.dout(n25068),.clk(gclk));
	jor g24811(.dina(n25068),.dinb(w_n24856_18[1]),.dout(n25069),.clk(gclk));
	jxor g24812(.dina(n25069),.dinb(w_n24241_0[0]),.dout(n25070),.clk(gclk));
	jand g24813(.dina(w_n25070_0[1]),.dinb(w_n11347_9[1]),.dout(n25071),.clk(gclk));
	jor g24814(.dina(n25071),.dinb(n25067),.dout(n25072),.clk(gclk));
	jor g24815(.dina(n25072),.dinb(n25066),.dout(n25073),.clk(gclk));
	jor g24816(.dina(w_n25070_0[0]),.dinb(w_n11347_9[0]),.dout(n25074),.clk(gclk));
	jor g24817(.dina(w_n24921_0[0]),.dinb(w_n10824_15[2]),.dout(n25075),.clk(gclk));
	jand g24818(.dina(n25075),.dinb(n25074),.dout(n25076),.clk(gclk));
	jand g24819(.dina(n25076),.dinb(n25073),.dout(n25077),.clk(gclk));
	jor g24820(.dina(n25077),.dinb(n24922),.dout(n25078),.clk(gclk));
	jor g24821(.dina(w_n24917_0[0]),.dinb(w_n10328_10[1]),.dout(n25079),.clk(gclk));
	jand g24822(.dina(n25079),.dinb(n25078),.dout(n25080),.clk(gclk));
	jxor g24823(.dina(w_n24258_0[0]),.dinb(w_n10328_10[0]),.dout(n25081),.clk(gclk));
	jor g24824(.dina(n25081),.dinb(w_n24856_18[0]),.dout(n25082),.clk(gclk));
	jxor g24825(.dina(n25082),.dinb(w_n24264_0[0]),.dout(n25083),.clk(gclk));
	jand g24826(.dina(w_n25083_0[1]),.dinb(w_n9832_17[0]),.dout(n25084),.clk(gclk));
	jor g24827(.dina(n25084),.dinb(n25080),.dout(n25085),.clk(gclk));
	jor g24828(.dina(n25085),.dinb(n24918),.dout(n25086),.clk(gclk));
	jor g24829(.dina(w_n25083_0[0]),.dinb(w_n9832_16[2]),.dout(n25087),.clk(gclk));
	jxor g24830(.dina(w_n24266_0[0]),.dinb(w_n9832_16[1]),.dout(n25088),.clk(gclk));
	jor g24831(.dina(n25088),.dinb(w_n24856_17[2]),.dout(n25089),.clk(gclk));
	jxor g24832(.dina(n25089),.dinb(w_n24271_0[0]),.dout(n25090),.clk(gclk));
	jor g24833(.dina(w_n25090_0[1]),.dinb(w_n9369_11[2]),.dout(n25091),.clk(gclk));
	jand g24834(.dina(n25091),.dinb(n25087),.dout(n25092),.clk(gclk));
	jand g24835(.dina(n25092),.dinb(n25086),.dout(n25093),.clk(gclk));
	jand g24836(.dina(w_n25090_0[0]),.dinb(w_n9369_11[1]),.dout(n25094),.clk(gclk));
	jxor g24837(.dina(w_n24273_0[0]),.dinb(w_n9369_11[0]),.dout(n25095),.clk(gclk));
	jor g24838(.dina(n25095),.dinb(w_n24856_17[1]),.dout(n25096),.clk(gclk));
	jxor g24839(.dina(n25096),.dinb(w_n24279_0[0]),.dout(n25097),.clk(gclk));
	jand g24840(.dina(w_n25097_0[1]),.dinb(w_n8890_17[0]),.dout(n25098),.clk(gclk));
	jor g24841(.dina(n25098),.dinb(n25094),.dout(n25099),.clk(gclk));
	jor g24842(.dina(n25099),.dinb(n25093),.dout(n25100),.clk(gclk));
	jor g24843(.dina(w_n25097_0[0]),.dinb(w_n8890_16[2]),.dout(n25101),.clk(gclk));
	jand g24844(.dina(n25101),.dinb(n25100),.dout(n25102),.clk(gclk));
	jand g24845(.dina(w_n24913_0[0]),.dinb(w_n8449_11[2]),.dout(n25103),.clk(gclk));
	jor g24846(.dina(n25103),.dinb(n25102),.dout(n25104),.clk(gclk));
	jor g24847(.dina(w_n24909_0[0]),.dinb(w_n8003_17[1]),.dout(n25105),.clk(gclk));
	jand g24848(.dina(n25105),.dinb(n25104),.dout(n25106),.clk(gclk));
	jand g24849(.dina(n25106),.dinb(n24914),.dout(n25107),.clk(gclk));
	jor g24850(.dina(n25107),.dinb(n24910),.dout(n25108),.clk(gclk));
	jor g24851(.dina(w_n24905_0[0]),.dinb(w_n7581_13[0]),.dout(n25109),.clk(gclk));
	jand g24852(.dina(n25109),.dinb(n25108),.dout(n25110),.clk(gclk));
	jxor g24853(.dina(w_n24304_0[0]),.dinb(w_n7581_12[2]),.dout(n25111),.clk(gclk));
	jor g24854(.dina(n25111),.dinb(w_n24856_17[0]),.dout(n25112),.clk(gclk));
	jxor g24855(.dina(n25112),.dinb(w_n24309_0[0]),.dout(n25113),.clk(gclk));
	jand g24856(.dina(w_n25113_0[1]),.dinb(w_n7154_18[1]),.dout(n25114),.clk(gclk));
	jor g24857(.dina(n25114),.dinb(n25110),.dout(n25115),.clk(gclk));
	jor g24858(.dina(n25115),.dinb(n24906),.dout(n25116),.clk(gclk));
	jxor g24859(.dina(w_n24311_0[0]),.dinb(w_n7154_18[0]),.dout(n25117),.clk(gclk));
	jor g24860(.dina(n25117),.dinb(w_n24856_16[2]),.dout(n25118),.clk(gclk));
	jxor g24861(.dina(n25118),.dinb(w_n24316_0[0]),.dout(n25119),.clk(gclk));
	jor g24862(.dina(w_n25119_0[1]),.dinb(w_n6758_13[2]),.dout(n25120),.clk(gclk));
	jor g24863(.dina(w_n25113_0[0]),.dinb(w_n7154_17[2]),.dout(n25121),.clk(gclk));
	jand g24864(.dina(n25121),.dinb(n25120),.dout(n25122),.clk(gclk));
	jand g24865(.dina(n25122),.dinb(n25116),.dout(n25123),.clk(gclk));
	jand g24866(.dina(w_n25119_0[0]),.dinb(w_n6758_13[1]),.dout(n25124),.clk(gclk));
	jand g24867(.dina(w_n24901_0[0]),.dinb(w_n6357_18[1]),.dout(n25125),.clk(gclk));
	jor g24868(.dina(n25125),.dinb(n25124),.dout(n25126),.clk(gclk));
	jor g24869(.dina(n25126),.dinb(n25123),.dout(n25127),.clk(gclk));
	jxor g24870(.dina(w_n24326_0[0]),.dinb(w_n6357_18[0]),.dout(n25128),.clk(gclk));
	jor g24871(.dina(n25128),.dinb(w_n24856_16[1]),.dout(n25129),.clk(gclk));
	jxor g24872(.dina(n25129),.dinb(w_n24331_0[0]),.dout(n25130),.clk(gclk));
	jor g24873(.dina(w_n25130_0[1]),.dinb(w_n5989_14[2]),.dout(n25131),.clk(gclk));
	jand g24874(.dina(n25131),.dinb(n25127),.dout(n25132),.clk(gclk));
	jand g24875(.dina(n25132),.dinb(n24902),.dout(n25133),.clk(gclk));
	jand g24876(.dina(w_n25130_0[0]),.dinb(w_n5989_14[1]),.dout(n25134),.clk(gclk));
	jxor g24877(.dina(w_n24333_0[0]),.dinb(w_n5989_14[0]),.dout(n25135),.clk(gclk));
	jor g24878(.dina(n25135),.dinb(w_n24856_16[0]),.dout(n25136),.clk(gclk));
	jxor g24879(.dina(n25136),.dinb(w_n24339_0[0]),.dout(n25137),.clk(gclk));
	jand g24880(.dina(w_n25137_0[1]),.dinb(w_n5606_19[0]),.dout(n25138),.clk(gclk));
	jor g24881(.dina(n25138),.dinb(n25134),.dout(n25139),.clk(gclk));
	jor g24882(.dina(n25139),.dinb(n25133),.dout(n25140),.clk(gclk));
	jxor g24883(.dina(w_n24341_0[0]),.dinb(w_n5606_18[2]),.dout(n25141),.clk(gclk));
	jor g24884(.dina(n25141),.dinb(w_n24856_15[2]),.dout(n25142),.clk(gclk));
	jxor g24885(.dina(n25142),.dinb(w_n24346_0[0]),.dout(n25143),.clk(gclk));
	jor g24886(.dina(w_n25143_0[1]),.dinb(w_n5259_15[2]),.dout(n25144),.clk(gclk));
	jor g24887(.dina(w_n25137_0[0]),.dinb(w_n5606_18[1]),.dout(n25145),.clk(gclk));
	jand g24888(.dina(n25145),.dinb(n25144),.dout(n25146),.clk(gclk));
	jand g24889(.dina(n25146),.dinb(n25140),.dout(n25147),.clk(gclk));
	jand g24890(.dina(w_n25143_0[0]),.dinb(w_n5259_15[1]),.dout(n25148),.clk(gclk));
	jxor g24891(.dina(w_n24348_0[0]),.dinb(w_n5259_15[0]),.dout(n25149),.clk(gclk));
	jor g24892(.dina(n25149),.dinb(w_n24856_15[1]),.dout(n25150),.clk(gclk));
	jxor g24893(.dina(n25150),.dinb(w_n24354_0[0]),.dout(n25151),.clk(gclk));
	jand g24894(.dina(w_n25151_0[1]),.dinb(w_n4902_19[1]),.dout(n25152),.clk(gclk));
	jor g24895(.dina(n25152),.dinb(n25148),.dout(n25153),.clk(gclk));
	jor g24896(.dina(n25153),.dinb(n25147),.dout(n25154),.clk(gclk));
	jor g24897(.dina(w_n25151_0[0]),.dinb(w_n4902_19[0]),.dout(n25155),.clk(gclk));
	jor g24898(.dina(w_n24897_0[0]),.dinb(w_n4582_16[0]),.dout(n25156),.clk(gclk));
	jand g24899(.dina(n25156),.dinb(n25155),.dout(n25157),.clk(gclk));
	jand g24900(.dina(n25157),.dinb(n25154),.dout(n25158),.clk(gclk));
	jor g24901(.dina(n25158),.dinb(n24898),.dout(n25159),.clk(gclk));
	jand g24902(.dina(n25159),.dinb(n24894),.dout(n25160),.clk(gclk));
	jand g24903(.dina(w_n24893_0[0]),.dinb(w_n4249_20[0]),.dout(n25161),.clk(gclk));
	jxor g24904(.dina(w_n24372_0[0]),.dinb(w_n4249_19[2]),.dout(n25162),.clk(gclk));
	jor g24905(.dina(n25162),.dinb(w_n24856_15[0]),.dout(n25163),.clk(gclk));
	jxor g24906(.dina(n25163),.dinb(w_n24377_0[0]),.dout(n25164),.clk(gclk));
	jand g24907(.dina(w_n25164_0[1]),.dinb(w_n3955_17[1]),.dout(n25165),.clk(gclk));
	jor g24908(.dina(n25165),.dinb(n25161),.dout(n25166),.clk(gclk));
	jor g24909(.dina(n25166),.dinb(n25160),.dout(n25167),.clk(gclk));
	jor g24910(.dina(w_n25164_0[0]),.dinb(w_n3955_17[0]),.dout(n25168),.clk(gclk));
	jxor g24911(.dina(w_n24379_0[0]),.dinb(w_n3955_16[2]),.dout(n25169),.clk(gclk));
	jor g24912(.dina(n25169),.dinb(w_n24856_14[2]),.dout(n25170),.clk(gclk));
	jxor g24913(.dina(n25170),.dinb(w_n24385_0[0]),.dout(n25171),.clk(gclk));
	jor g24914(.dina(w_n25171_0[1]),.dinb(w_n3642_20[2]),.dout(n25172),.clk(gclk));
	jand g24915(.dina(n25172),.dinb(n25168),.dout(n25173),.clk(gclk));
	jand g24916(.dina(n25173),.dinb(n25167),.dout(n25174),.clk(gclk));
	jand g24917(.dina(w_n25171_0[0]),.dinb(w_n3642_20[1]),.dout(n25175),.clk(gclk));
	jxor g24918(.dina(w_n24387_0[0]),.dinb(w_n3642_20[0]),.dout(n25176),.clk(gclk));
	jor g24919(.dina(n25176),.dinb(w_n24856_14[1]),.dout(n25177),.clk(gclk));
	jxor g24920(.dina(n25177),.dinb(w_n24392_0[0]),.dout(n25178),.clk(gclk));
	jand g24921(.dina(w_n25178_0[1]),.dinb(w_n3368_17[2]),.dout(n25179),.clk(gclk));
	jor g24922(.dina(n25179),.dinb(n25175),.dout(n25180),.clk(gclk));
	jor g24923(.dina(n25180),.dinb(n25174),.dout(n25181),.clk(gclk));
	jor g24924(.dina(w_n25178_0[0]),.dinb(w_n3368_17[1]),.dout(n25182),.clk(gclk));
	jor g24925(.dina(w_n24889_0[0]),.dinb(w_n3089_21[0]),.dout(n25183),.clk(gclk));
	jand g24926(.dina(n25183),.dinb(n25182),.dout(n25184),.clk(gclk));
	jand g24927(.dina(n25184),.dinb(n25181),.dout(n25185),.clk(gclk));
	jor g24928(.dina(n25185),.dinb(n24890),.dout(n25186),.clk(gclk));
	jxor g24929(.dina(w_n24402_0[0]),.dinb(w_n3089_20[2]),.dout(n25187),.clk(gclk));
	jor g24930(.dina(n25187),.dinb(w_n24856_14[0]),.dout(n25188),.clk(gclk));
	jxor g24931(.dina(n25188),.dinb(w_n24407_0[0]),.dout(n25189),.clk(gclk));
	jor g24932(.dina(w_n25189_0[1]),.dinb(w_n2833_19[0]),.dout(n25190),.clk(gclk));
	jand g24933(.dina(n25190),.dinb(n25186),.dout(n25191),.clk(gclk));
	jand g24934(.dina(w_n25189_0[0]),.dinb(w_n2833_18[2]),.dout(n25192),.clk(gclk));
	jxor g24935(.dina(w_n24409_0[0]),.dinb(w_n2833_18[1]),.dout(n25193),.clk(gclk));
	jor g24936(.dina(n25193),.dinb(w_n24856_13[2]),.dout(n25194),.clk(gclk));
	jxor g24937(.dina(n25194),.dinb(w_n24415_0[0]),.dout(n25195),.clk(gclk));
	jand g24938(.dina(w_n25195_0[1]),.dinb(w_n2572_21[1]),.dout(n25196),.clk(gclk));
	jor g24939(.dina(n25196),.dinb(n25192),.dout(n25197),.clk(gclk));
	jor g24940(.dina(n25197),.dinb(n25191),.dout(n25198),.clk(gclk));
	jor g24941(.dina(w_n25195_0[0]),.dinb(w_n2572_21[0]),.dout(n25199),.clk(gclk));
	jor g24942(.dina(w_n24885_0[0]),.dinb(w_n2345_19[0]),.dout(n25200),.clk(gclk));
	jand g24943(.dina(n25200),.dinb(n25199),.dout(n25201),.clk(gclk));
	jand g24944(.dina(n25201),.dinb(n25198),.dout(n25202),.clk(gclk));
	jor g24945(.dina(n25202),.dinb(n24886),.dout(n25203),.clk(gclk));
	jand g24946(.dina(n25203),.dinb(n24882),.dout(n25204),.clk(gclk));
	jand g24947(.dina(w_n24881_0[0]),.dinb(w_n2108_22[0]),.dout(n25205),.clk(gclk));
	jxor g24948(.dina(w_n24432_0[0]),.dinb(w_n2108_21[2]),.dout(n25206),.clk(gclk));
	jor g24949(.dina(n25206),.dinb(w_n24856_13[1]),.dout(n25207),.clk(gclk));
	jxor g24950(.dina(n25207),.dinb(w_n24438_0[0]),.dout(n25208),.clk(gclk));
	jand g24951(.dina(w_n25208_0[1]),.dinb(w_n1912_20[2]),.dout(n25209),.clk(gclk));
	jor g24952(.dina(n25209),.dinb(n25205),.dout(n25210),.clk(gclk));
	jor g24953(.dina(n25210),.dinb(n25204),.dout(n25211),.clk(gclk));
	jor g24954(.dina(w_n25208_0[0]),.dinb(w_n1912_20[1]),.dout(n25212),.clk(gclk));
	jxor g24955(.dina(w_n24440_0[0]),.dinb(w_n1912_20[0]),.dout(n25213),.clk(gclk));
	jor g24956(.dina(n25213),.dinb(w_n24856_13[0]),.dout(n25214),.clk(gclk));
	jxor g24957(.dina(n25214),.dinb(w_n24446_0[0]),.dout(n25215),.clk(gclk));
	jor g24958(.dina(w_n25215_0[1]),.dinb(w_n1699_23[0]),.dout(n25216),.clk(gclk));
	jand g24959(.dina(n25216),.dinb(n25212),.dout(n25217),.clk(gclk));
	jand g24960(.dina(n25217),.dinb(n25211),.dout(n25218),.clk(gclk));
	jand g24961(.dina(w_n25215_0[0]),.dinb(w_n1699_22[2]),.dout(n25219),.clk(gclk));
	jxor g24962(.dina(w_n24448_0[0]),.dinb(w_n1699_22[1]),.dout(n25220),.clk(gclk));
	jor g24963(.dina(n25220),.dinb(w_n24856_12[2]),.dout(n25221),.clk(gclk));
	jxor g24964(.dina(n25221),.dinb(w_n24453_0[0]),.dout(n25222),.clk(gclk));
	jand g24965(.dina(w_n25222_0[1]),.dinb(w_n1516_21[0]),.dout(n25223),.clk(gclk));
	jor g24966(.dina(n25223),.dinb(n25219),.dout(n25224),.clk(gclk));
	jor g24967(.dina(n25224),.dinb(n25218),.dout(n25225),.clk(gclk));
	jor g24968(.dina(w_n25222_0[0]),.dinb(w_n1516_20[2]),.dout(n25226),.clk(gclk));
	jor g24969(.dina(w_n24877_0[0]),.dinb(w_n1332_22[1]),.dout(n25227),.clk(gclk));
	jand g24970(.dina(n25227),.dinb(n25226),.dout(n25228),.clk(gclk));
	jand g24971(.dina(n25228),.dinb(n25225),.dout(n25229),.clk(gclk));
	jor g24972(.dina(n25229),.dinb(n24878),.dout(n25230),.clk(gclk));
	jor g24973(.dina(w_n24873_0[0]),.dinb(w_n1173_21[2]),.dout(n25231),.clk(gclk));
	jand g24974(.dina(n25231),.dinb(n25230),.dout(n25232),.clk(gclk));
	jxor g24975(.dina(w_n24471_0[0]),.dinb(w_n1173_21[1]),.dout(n25233),.clk(gclk));
	jor g24976(.dina(n25233),.dinb(w_n24856_12[1]),.dout(n25234),.clk(gclk));
	jxor g24977(.dina(n25234),.dinb(w_n24477_0[0]),.dout(n25235),.clk(gclk));
	jand g24978(.dina(w_n25235_0[1]),.dinb(w_n1008_23[2]),.dout(n25236),.clk(gclk));
	jor g24979(.dina(n25236),.dinb(n25232),.dout(n25237),.clk(gclk));
	jor g24980(.dina(n25237),.dinb(n24874),.dout(n25238),.clk(gclk));
	jor g24981(.dina(w_n25235_0[0]),.dinb(w_n1008_23[1]),.dout(n25239),.clk(gclk));
	jor g24982(.dina(w_n24867_0[0]),.dinb(w_n884_22[1]),.dout(n25240),.clk(gclk));
	jand g24983(.dina(n25240),.dinb(n25239),.dout(n25241),.clk(gclk));
	jand g24984(.dina(n25241),.dinb(n25238),.dout(n25242),.clk(gclk));
	jor g24985(.dina(n25242),.dinb(n24870),.dout(n25243),.clk(gclk));
	jxor g24986(.dina(w_n24495_0[0]),.dinb(w_n743_23[1]),.dout(n25244),.clk(gclk));
	jor g24987(.dina(n25244),.dinb(w_n24856_12[0]),.dout(n25245),.clk(gclk));
	jxor g24988(.dina(n25245),.dinb(w_n24500_0[0]),.dout(n25246),.clk(gclk));
	jor g24989(.dina(w_n25246_0[1]),.dinb(w_n635_24[0]),.dout(n25247),.clk(gclk));
	jand g24990(.dina(n25247),.dinb(n25243),.dout(n25248),.clk(gclk));
	jand g24991(.dina(n25248),.dinb(n24864),.dout(n25249),.clk(gclk));
	jand g24992(.dina(w_n25246_0[0]),.dinb(w_n635_23[2]),.dout(n25250),.clk(gclk));
	jxor g24993(.dina(w_n24502_0[0]),.dinb(w_n635_23[1]),.dout(n25251),.clk(gclk));
	jor g24994(.dina(n25251),.dinb(w_n24856_11[2]),.dout(n25252),.clk(gclk));
	jxor g24995(.dina(n25252),.dinb(w_n24508_0[0]),.dout(n25253),.clk(gclk));
	jand g24996(.dina(w_n25253_0[1]),.dinb(w_n515_25[0]),.dout(n25254),.clk(gclk));
	jor g24997(.dina(n25254),.dinb(n25250),.dout(n25255),.clk(gclk));
	jor g24998(.dina(n25255),.dinb(n25249),.dout(n25256),.clk(gclk));
	jor g24999(.dina(w_n25253_0[0]),.dinb(w_n515_24[2]),.dout(n25257),.clk(gclk));
	jxor g25000(.dina(w_n24510_0[0]),.dinb(w_n515_24[1]),.dout(n25258),.clk(gclk));
	jor g25001(.dina(n25258),.dinb(w_n24856_11[1]),.dout(n25259),.clk(gclk));
	jxor g25002(.dina(n25259),.dinb(w_n24515_0[0]),.dout(n25260),.clk(gclk));
	jor g25003(.dina(w_n25260_0[1]),.dinb(w_n443_25[0]),.dout(n25261),.clk(gclk));
	jand g25004(.dina(n25261),.dinb(n25257),.dout(n25262),.clk(gclk));
	jand g25005(.dina(n25262),.dinb(n25256),.dout(n25263),.clk(gclk));
	jand g25006(.dina(w_n25260_0[0]),.dinb(w_n443_24[2]),.dout(n25264),.clk(gclk));
	jxor g25007(.dina(w_n24517_0[0]),.dinb(w_n443_24[1]),.dout(n25265),.clk(gclk));
	jor g25008(.dina(n25265),.dinb(w_n24856_11[0]),.dout(n25266),.clk(gclk));
	jxor g25009(.dina(n25266),.dinb(w_n24523_0[0]),.dout(n25267),.clk(gclk));
	jand g25010(.dina(w_n25267_0[1]),.dinb(w_n352_25[1]),.dout(n25268),.clk(gclk));
	jor g25011(.dina(n25268),.dinb(n25264),.dout(n25269),.clk(gclk));
	jor g25012(.dina(n25269),.dinb(n25263),.dout(n25270),.clk(gclk));
	jxor g25013(.dina(w_n24525_0[0]),.dinb(w_n352_25[0]),.dout(n25271),.clk(gclk));
	jor g25014(.dina(n25271),.dinb(w_n24856_10[2]),.dout(n25272),.clk(gclk));
	jxor g25015(.dina(n25272),.dinb(w_n24530_0[0]),.dout(n25273),.clk(gclk));
	jor g25016(.dina(w_n25273_0[1]),.dinb(w_n294_25[2]),.dout(n25274),.clk(gclk));
	jor g25017(.dina(w_n25267_0[0]),.dinb(w_n352_24[2]),.dout(n25275),.clk(gclk));
	jand g25018(.dina(n25275),.dinb(n25274),.dout(n25276),.clk(gclk));
	jand g25019(.dina(n25276),.dinb(n25270),.dout(n25277),.clk(gclk));
	jand g25020(.dina(w_n25273_0[0]),.dinb(w_n294_25[1]),.dout(n25278),.clk(gclk));
	jxor g25021(.dina(w_n24532_0[0]),.dinb(w_n294_25[0]),.dout(n25279),.clk(gclk));
	jor g25022(.dina(n25279),.dinb(w_n24856_10[1]),.dout(n25280),.clk(gclk));
	jxor g25023(.dina(n25280),.dinb(w_n24537_0[0]),.dout(n25281),.clk(gclk));
	jand g25024(.dina(w_n25281_0[1]),.dinb(w_n239_25[1]),.dout(n25282),.clk(gclk));
	jor g25025(.dina(n25282),.dinb(n25278),.dout(n25283),.clk(gclk));
	jor g25026(.dina(n25283),.dinb(n25277),.dout(n25284),.clk(gclk));
	jor g25027(.dina(w_n25281_0[0]),.dinb(w_n239_25[0]),.dout(n25285),.clk(gclk));
	jor g25028(.dina(w_n24859_0[0]),.dinb(w_n221_25[2]),.dout(n25286),.clk(gclk));
	jand g25029(.dina(n25286),.dinb(n25285),.dout(n25287),.clk(gclk));
	jand g25030(.dina(n25287),.dinb(n25284),.dout(n25288),.clk(gclk));
	jor g25031(.dina(n25288),.dinb(n24860),.dout(n25289),.clk(gclk));
	jxor g25032(.dina(w_n24546_0[0]),.dinb(w_n221_25[1]),.dout(n25290),.clk(gclk));
	jor g25033(.dina(n25290),.dinb(w_n24856_10[0]),.dout(n25291),.clk(gclk));
	jxor g25034(.dina(n25291),.dinb(w_n24552_0[0]),.dout(n25292),.clk(gclk));
	jor g25035(.dina(w_n25292_0[1]),.dinb(w_n218_10[2]),.dout(n25293),.clk(gclk));
	jand g25036(.dina(n25293),.dinb(n25289),.dout(n25294),.clk(gclk));
	jand g25037(.dina(w_asqrt1_0[1]),.dinb(w_n24852_0[0]),.dout(n25295),.clk(gclk));
	jnot g25038(.din(w_n24835_0[0]),.dout(n25296),.clk(gclk));
	jor g25039(.dina(w_n25292_0[0]),.dinb(n25296),.dout(n25297),.clk(gclk));
	jor g25040(.dina(n25297),.dinb(n25295),.dout(n25298),.clk(gclk));
	jand g25041(.dina(n25298),.dinb(w_n218_10[1]),.dout(n25299),.clk(gclk));
	jor g25042(.dina(n25299),.dinb(n25294),.dout(n25300),.clk(gclk));
	jor g25043(.dina(n25300),.dinb(n24850),.dout(asqrt_fa_1),.clk(gclk));
	jspl3 jspl3_w_a2_0(.douta(w_a2_0[0]),.doutb(w_a2_0[1]),.doutc(w_a2_0[2]),.din(a[2]));
	jspl jspl_w_a2_1(.douta(w_a2_1[0]),.doutb(w_a2_1[1]),.din(w_a2_0[0]));
	jspl jspl_w_a3_0(.douta(w_a3_0[0]),.doutb(w_a3_0[1]),.din(a[3]));
	jspl3 jspl3_w_a4_0(.douta(w_a4_0[0]),.doutb(w_a4_0[1]),.doutc(w_a4_0[2]),.din(a[4]));
	jspl jspl_w_a4_1(.douta(w_a4_1[0]),.doutb(w_a4_1[1]),.din(w_a4_0[0]));
	jspl jspl_w_a5_0(.douta(w_a5_0[0]),.doutb(w_a5_0[1]),.din(a[5]));
	jspl3 jspl3_w_a6_0(.douta(w_a6_0[0]),.doutb(w_a6_0[1]),.doutc(w_a6_0[2]),.din(a[6]));
	jspl jspl_w_a7_0(.douta(w_a7_0[0]),.doutb(w_a7_0[1]),.din(a[7]));
	jspl3 jspl3_w_a8_0(.douta(w_a8_0[0]),.doutb(w_a8_0[1]),.doutc(w_a8_0[2]),.din(a[8]));
	jspl jspl_w_a9_0(.douta(w_a9_0[0]),.doutb(w_a9_0[1]),.din(a[9]));
	jspl3 jspl3_w_a10_0(.douta(w_a10_0[0]),.doutb(w_a10_0[1]),.doutc(w_a10_0[2]),.din(a[10]));
	jspl jspl_w_a11_0(.douta(w_a11_0[0]),.doutb(w_a11_0[1]),.din(a[11]));
	jspl3 jspl3_w_a12_0(.douta(w_a12_0[0]),.doutb(w_a12_0[1]),.doutc(w_a12_0[2]),.din(a[12]));
	jspl jspl_w_a13_0(.douta(w_a13_0[0]),.doutb(w_a13_0[1]),.din(a[13]));
	jspl3 jspl3_w_a14_0(.douta(w_a14_0[0]),.doutb(w_a14_0[1]),.doutc(w_a14_0[2]),.din(a[14]));
	jspl jspl_w_a14_1(.douta(w_a14_1[0]),.doutb(w_a14_1[1]),.din(w_a14_0[0]));
	jspl jspl_w_a15_0(.douta(w_a15_0[0]),.doutb(w_a15_0[1]),.din(a[15]));
	jspl3 jspl3_w_a16_0(.douta(w_a16_0[0]),.doutb(w_a16_0[1]),.doutc(w_a16_0[2]),.din(a[16]));
	jspl jspl_w_a17_0(.douta(w_a17_0[0]),.doutb(w_a17_0[1]),.din(a[17]));
	jspl3 jspl3_w_a18_0(.douta(w_a18_0[0]),.doutb(w_a18_0[1]),.doutc(w_a18_0[2]),.din(a[18]));
	jspl jspl_w_a18_1(.douta(w_a18_1[0]),.doutb(w_a18_1[1]),.din(w_a18_0[0]));
	jspl jspl_w_a19_0(.douta(w_a19_0[0]),.doutb(w_a19_0[1]),.din(a[19]));
	jspl3 jspl3_w_a20_0(.douta(w_a20_0[0]),.doutb(w_a20_0[1]),.doutc(w_a20_0[2]),.din(a[20]));
	jspl jspl_w_a21_0(.douta(w_a21_0[0]),.doutb(w_a21_0[1]),.din(a[21]));
	jspl3 jspl3_w_a22_0(.douta(w_a22_0[0]),.doutb(w_a22_0[1]),.doutc(w_a22_0[2]),.din(a[22]));
	jspl jspl_w_a22_1(.douta(w_a22_1[0]),.doutb(w_a22_1[1]),.din(w_a22_0[0]));
	jspl jspl_w_a23_0(.douta(w_a23_0[0]),.doutb(w_a23_0[1]),.din(a[23]));
	jspl3 jspl3_w_a24_0(.douta(w_a24_0[0]),.doutb(w_a24_0[1]),.doutc(w_a24_0[2]),.din(a[24]));
	jspl jspl_w_a25_0(.douta(w_a25_0[0]),.doutb(w_a25_0[1]),.din(a[25]));
	jspl3 jspl3_w_a26_0(.douta(w_a26_0[0]),.doutb(w_a26_0[1]),.doutc(w_a26_0[2]),.din(a[26]));
	jspl jspl_w_a26_1(.douta(w_a26_1[0]),.doutb(w_a26_1[1]),.din(w_a26_0[0]));
	jspl jspl_w_a27_0(.douta(w_a27_0[0]),.doutb(w_a27_0[1]),.din(a[27]));
	jspl3 jspl3_w_a28_0(.douta(w_a28_0[0]),.doutb(w_a28_0[1]),.doutc(w_a28_0[2]),.din(a[28]));
	jspl jspl_w_a29_0(.douta(w_a29_0[0]),.doutb(w_a29_0[1]),.din(a[29]));
	jspl3 jspl3_w_a30_0(.douta(w_a30_0[0]),.doutb(w_a30_0[1]),.doutc(w_a30_0[2]),.din(a[30]));
	jspl jspl_w_a30_1(.douta(w_a30_1[0]),.doutb(w_a30_1[1]),.din(w_a30_0[0]));
	jspl jspl_w_a31_0(.douta(w_a31_0[0]),.doutb(w_a31_0[1]),.din(a[31]));
	jspl3 jspl3_w_a32_0(.douta(w_a32_0[0]),.doutb(w_a32_0[1]),.doutc(w_a32_0[2]),.din(a[32]));
	jspl jspl_w_a33_0(.douta(w_a33_0[0]),.doutb(w_a33_0[1]),.din(a[33]));
	jspl3 jspl3_w_a34_0(.douta(w_a34_0[0]),.doutb(w_a34_0[1]),.doutc(w_a34_0[2]),.din(a[34]));
	jspl jspl_w_a34_1(.douta(w_a34_1[0]),.doutb(w_a34_1[1]),.din(w_a34_0[0]));
	jspl jspl_w_a35_0(.douta(w_a35_0[0]),.doutb(w_a35_0[1]),.din(a[35]));
	jspl3 jspl3_w_a36_0(.douta(w_a36_0[0]),.doutb(w_a36_0[1]),.doutc(w_a36_0[2]),.din(a[36]));
	jspl jspl_w_a37_0(.douta(w_a37_0[0]),.doutb(w_a37_0[1]),.din(a[37]));
	jspl3 jspl3_w_a38_0(.douta(w_a38_0[0]),.doutb(w_a38_0[1]),.doutc(w_a38_0[2]),.din(a[38]));
	jspl jspl_w_a39_0(.douta(w_a39_0[0]),.doutb(w_a39_0[1]),.din(a[39]));
	jspl3 jspl3_w_a40_0(.douta(w_a40_0[0]),.doutb(w_a40_0[1]),.doutc(w_a40_0[2]),.din(a[40]));
	jspl jspl_w_a41_0(.douta(w_a41_0[0]),.doutb(w_a41_0[1]),.din(a[41]));
	jspl3 jspl3_w_a42_0(.douta(w_a42_0[0]),.doutb(w_a42_0[1]),.doutc(w_a42_0[2]),.din(a[42]));
	jspl jspl_w_a42_1(.douta(w_a42_1[0]),.doutb(w_a42_1[1]),.din(w_a42_0[0]));
	jspl jspl_w_a43_0(.douta(w_a43_0[0]),.doutb(w_a43_0[1]),.din(a[43]));
	jspl3 jspl3_w_a44_0(.douta(w_a44_0[0]),.doutb(w_a44_0[1]),.doutc(w_a44_0[2]),.din(a[44]));
	jspl jspl_w_a45_0(.douta(w_a45_0[0]),.doutb(w_a45_0[1]),.din(a[45]));
	jspl3 jspl3_w_a46_0(.douta(w_a46_0[0]),.doutb(w_a46_0[1]),.doutc(w_a46_0[2]),.din(a[46]));
	jspl jspl_w_a46_1(.douta(w_a46_1[0]),.doutb(w_a46_1[1]),.din(w_a46_0[0]));
	jspl jspl_w_a47_0(.douta(w_a47_0[0]),.doutb(w_a47_0[1]),.din(a[47]));
	jspl3 jspl3_w_a48_0(.douta(w_a48_0[0]),.doutb(w_a48_0[1]),.doutc(w_a48_0[2]),.din(a[48]));
	jspl jspl_w_a49_0(.douta(w_a49_0[0]),.doutb(w_a49_0[1]),.din(a[49]));
	jspl3 jspl3_w_a50_0(.douta(w_a50_0[0]),.doutb(w_a50_0[1]),.doutc(w_a50_0[2]),.din(a[50]));
	jspl jspl_w_a51_0(.douta(w_a51_0[0]),.doutb(w_a51_0[1]),.din(a[51]));
	jspl3 jspl3_w_a52_0(.douta(w_a52_0[0]),.doutb(w_a52_0[1]),.doutc(w_a52_0[2]),.din(a[52]));
	jspl jspl_w_a53_0(.douta(w_a53_0[0]),.doutb(w_a53_0[1]),.din(a[53]));
	jspl3 jspl3_w_a54_0(.douta(w_a54_0[0]),.doutb(w_a54_0[1]),.doutc(w_a54_0[2]),.din(a[54]));
	jspl jspl_w_a54_1(.douta(w_a54_1[0]),.doutb(w_a54_1[1]),.din(w_a54_0[0]));
	jspl jspl_w_a55_0(.douta(w_a55_0[0]),.doutb(w_a55_0[1]),.din(a[55]));
	jspl3 jspl3_w_a56_0(.douta(w_a56_0[0]),.doutb(w_a56_0[1]),.doutc(w_a56_0[2]),.din(a[56]));
	jspl jspl_w_a57_0(.douta(w_a57_0[0]),.doutb(w_a57_0[1]),.din(a[57]));
	jspl3 jspl3_w_a58_0(.douta(w_a58_0[0]),.doutb(w_a58_0[1]),.doutc(w_a58_0[2]),.din(a[58]));
	jspl jspl_w_a59_0(.douta(w_a59_0[0]),.doutb(w_a59_0[1]),.din(a[59]));
	jspl3 jspl3_w_a60_0(.douta(w_a60_0[0]),.doutb(w_a60_0[1]),.doutc(w_a60_0[2]),.din(a[60]));
	jspl jspl_w_a61_0(.douta(w_a61_0[0]),.doutb(w_a61_0[1]),.din(a[61]));
	jspl3 jspl3_w_a62_0(.douta(w_a62_0[0]),.doutb(w_a62_0[1]),.doutc(w_a62_0[2]),.din(a[62]));
	jspl jspl_w_a63_0(.douta(w_a63_0[0]),.doutb(w_a63_0[1]),.din(a[63]));
	jspl3 jspl3_w_a64_0(.douta(w_a64_0[0]),.doutb(w_a64_0[1]),.doutc(w_a64_0[2]),.din(a[64]));
	jspl jspl_w_a65_0(.douta(w_a65_0[0]),.doutb(w_a65_0[1]),.din(a[65]));
	jspl3 jspl3_w_a66_0(.douta(w_a66_0[0]),.doutb(w_a66_0[1]),.doutc(w_a66_0[2]),.din(a[66]));
	jspl jspl_w_a66_1(.douta(w_a66_1[0]),.doutb(w_a66_1[1]),.din(w_a66_0[0]));
	jspl jspl_w_a67_0(.douta(w_a67_0[0]),.doutb(w_a67_0[1]),.din(a[67]));
	jspl3 jspl3_w_a68_0(.douta(w_a68_0[0]),.doutb(w_a68_0[1]),.doutc(w_a68_0[2]),.din(a[68]));
	jspl jspl_w_a69_0(.douta(w_a69_0[0]),.doutb(w_a69_0[1]),.din(a[69]));
	jspl3 jspl3_w_a70_0(.douta(w_a70_0[0]),.doutb(w_a70_0[1]),.doutc(w_a70_0[2]),.din(a[70]));
	jspl jspl_w_a70_1(.douta(w_a70_1[0]),.doutb(w_a70_1[1]),.din(w_a70_0[0]));
	jspl jspl_w_a71_0(.douta(w_a71_0[0]),.doutb(w_a71_0[1]),.din(a[71]));
	jspl3 jspl3_w_a72_0(.douta(w_a72_0[0]),.doutb(w_a72_0[1]),.doutc(w_a72_0[2]),.din(a[72]));
	jspl jspl_w_a73_0(.douta(w_a73_0[0]),.doutb(w_a73_0[1]),.din(a[73]));
	jspl3 jspl3_w_a74_0(.douta(w_a74_0[0]),.doutb(w_a74_0[1]),.doutc(w_a74_0[2]),.din(a[74]));
	jspl jspl_w_a74_1(.douta(w_a74_1[0]),.doutb(w_a74_1[1]),.din(w_a74_0[0]));
	jspl jspl_w_a75_0(.douta(w_a75_0[0]),.doutb(w_a75_0[1]),.din(a[75]));
	jspl3 jspl3_w_a76_0(.douta(w_a76_0[0]),.doutb(w_a76_0[1]),.doutc(w_a76_0[2]),.din(a[76]));
	jspl jspl_w_a77_0(.douta(w_a77_0[0]),.doutb(w_a77_0[1]),.din(a[77]));
	jspl3 jspl3_w_a78_0(.douta(w_a78_0[0]),.doutb(w_a78_0[1]),.doutc(w_a78_0[2]),.din(a[78]));
	jspl jspl_w_a78_1(.douta(w_a78_1[0]),.doutb(w_a78_1[1]),.din(w_a78_0[0]));
	jspl jspl_w_a79_0(.douta(w_a79_0[0]),.doutb(w_a79_0[1]),.din(a[79]));
	jspl3 jspl3_w_a80_0(.douta(w_a80_0[0]),.doutb(w_a80_0[1]),.doutc(w_a80_0[2]),.din(a[80]));
	jspl jspl_w_a81_0(.douta(w_a81_0[0]),.doutb(w_a81_0[1]),.din(a[81]));
	jspl3 jspl3_w_a82_0(.douta(w_a82_0[0]),.doutb(w_a82_0[1]),.doutc(w_a82_0[2]),.din(a[82]));
	jspl jspl_w_a82_1(.douta(w_a82_1[0]),.doutb(w_a82_1[1]),.din(w_a82_0[0]));
	jspl jspl_w_a83_0(.douta(w_a83_0[0]),.doutb(w_a83_0[1]),.din(a[83]));
	jspl3 jspl3_w_a84_0(.douta(w_a84_0[0]),.doutb(w_a84_0[1]),.doutc(w_a84_0[2]),.din(a[84]));
	jspl jspl_w_a85_0(.douta(w_a85_0[0]),.doutb(w_a85_0[1]),.din(a[85]));
	jspl3 jspl3_w_a86_0(.douta(w_a86_0[0]),.doutb(w_a86_0[1]),.doutc(w_a86_0[2]),.din(a[86]));
	jspl jspl_w_a86_1(.douta(w_a86_1[0]),.doutb(w_a86_1[1]),.din(w_a86_0[0]));
	jspl jspl_w_a87_0(.douta(w_a87_0[0]),.doutb(w_a87_0[1]),.din(a[87]));
	jspl3 jspl3_w_a88_0(.douta(w_a88_0[0]),.doutb(w_a88_0[1]),.doutc(w_a88_0[2]),.din(a[88]));
	jspl jspl_w_a89_0(.douta(w_a89_0[0]),.doutb(w_a89_0[1]),.din(a[89]));
	jspl3 jspl3_w_a90_0(.douta(w_a90_0[0]),.doutb(w_a90_0[1]),.doutc(w_a90_0[2]),.din(a[90]));
	jspl jspl_w_a90_1(.douta(w_a90_1[0]),.doutb(w_a90_1[1]),.din(w_a90_0[0]));
	jspl jspl_w_a91_0(.douta(w_a91_0[0]),.doutb(w_a91_0[1]),.din(a[91]));
	jspl3 jspl3_w_a92_0(.douta(w_a92_0[0]),.doutb(w_a92_0[1]),.doutc(w_a92_0[2]),.din(a[92]));
	jspl jspl_w_a93_0(.douta(w_a93_0[0]),.doutb(w_a93_0[1]),.din(a[93]));
	jspl3 jspl3_w_a94_0(.douta(w_a94_0[0]),.doutb(w_a94_0[1]),.doutc(w_a94_0[2]),.din(a[94]));
	jspl jspl_w_a94_1(.douta(w_a94_1[0]),.doutb(w_a94_1[1]),.din(w_a94_0[0]));
	jspl jspl_w_a95_0(.douta(w_a95_0[0]),.doutb(w_a95_0[1]),.din(a[95]));
	jspl3 jspl3_w_a96_0(.douta(w_a96_0[0]),.doutb(w_a96_0[1]),.doutc(w_a96_0[2]),.din(a[96]));
	jspl jspl_w_a97_0(.douta(w_a97_0[0]),.doutb(w_a97_0[1]),.din(a[97]));
	jspl3 jspl3_w_a98_0(.douta(w_a98_0[0]),.doutb(w_a98_0[1]),.doutc(w_a98_0[2]),.din(a[98]));
	jspl jspl_w_a98_1(.douta(w_a98_1[0]),.doutb(w_a98_1[1]),.din(w_a98_0[0]));
	jspl jspl_w_a99_0(.douta(w_a99_0[0]),.doutb(w_a99_0[1]),.din(a[99]));
	jspl3 jspl3_w_a100_0(.douta(w_a100_0[0]),.doutb(w_a100_0[1]),.doutc(w_a100_0[2]),.din(a[100]));
	jspl jspl_w_a101_0(.douta(w_a101_0[0]),.doutb(w_a101_0[1]),.din(a[101]));
	jspl3 jspl3_w_a102_0(.douta(w_a102_0[0]),.doutb(w_a102_0[1]),.doutc(w_a102_0[2]),.din(a[102]));
	jspl jspl_w_a102_1(.douta(w_a102_1[0]),.doutb(w_a102_1[1]),.din(w_a102_0[0]));
	jspl jspl_w_a103_0(.douta(w_a103_0[0]),.doutb(w_a103_0[1]),.din(a[103]));
	jspl3 jspl3_w_a104_0(.douta(w_a104_0[0]),.doutb(w_a104_0[1]),.doutc(w_a104_0[2]),.din(a[104]));
	jspl jspl_w_a105_0(.douta(w_a105_0[0]),.doutb(w_a105_0[1]),.din(a[105]));
	jspl3 jspl3_w_a106_0(.douta(w_a106_0[0]),.doutb(w_a106_0[1]),.doutc(w_a106_0[2]),.din(a[106]));
	jspl jspl_w_a106_1(.douta(w_a106_1[0]),.doutb(w_a106_1[1]),.din(w_a106_0[0]));
	jspl jspl_w_a107_0(.douta(w_a107_0[0]),.doutb(w_a107_0[1]),.din(a[107]));
	jspl3 jspl3_w_a108_0(.douta(w_a108_0[0]),.doutb(w_a108_0[1]),.doutc(w_a108_0[2]),.din(a[108]));
	jspl jspl_w_a109_0(.douta(w_a109_0[0]),.doutb(w_a109_0[1]),.din(a[109]));
	jspl3 jspl3_w_a110_0(.douta(w_a110_0[0]),.doutb(w_a110_0[1]),.doutc(w_a110_0[2]),.din(a[110]));
	jspl jspl_w_a110_1(.douta(w_a110_1[0]),.doutb(w_a110_1[1]),.din(w_a110_0[0]));
	jspl jspl_w_a111_0(.douta(w_a111_0[0]),.doutb(w_a111_0[1]),.din(a[111]));
	jspl3 jspl3_w_a112_0(.douta(w_a112_0[0]),.doutb(w_a112_0[1]),.doutc(w_a112_0[2]),.din(a[112]));
	jspl jspl_w_a113_0(.douta(w_a113_0[0]),.doutb(w_a113_0[1]),.din(a[113]));
	jspl3 jspl3_w_a114_0(.douta(w_a114_0[0]),.doutb(w_a114_0[1]),.doutc(w_a114_0[2]),.din(a[114]));
	jspl jspl_w_a114_1(.douta(w_a114_1[0]),.doutb(w_a114_1[1]),.din(w_a114_0[0]));
	jspl jspl_w_a115_0(.douta(w_a115_0[0]),.doutb(w_a115_0[1]),.din(a[115]));
	jspl3 jspl3_w_a116_0(.douta(w_a116_0[0]),.doutb(w_a116_0[1]),.doutc(w_a116_0[2]),.din(a[116]));
	jspl jspl_w_a117_0(.douta(w_a117_0[0]),.doutb(w_a117_0[1]),.din(a[117]));
	jspl3 jspl3_w_a118_0(.douta(w_a118_0[0]),.doutb(w_a118_0[1]),.doutc(w_a118_0[2]),.din(a[118]));
	jspl jspl_w_a118_1(.douta(w_a118_1[0]),.doutb(w_a118_1[1]),.din(w_a118_0[0]));
	jspl jspl_w_a119_0(.douta(w_a119_0[0]),.doutb(w_a119_0[1]),.din(a[119]));
	jspl3 jspl3_w_a120_0(.douta(w_a120_0[0]),.doutb(w_a120_0[1]),.doutc(w_a120_0[2]),.din(a[120]));
	jspl jspl_w_a121_0(.douta(w_a121_0[0]),.doutb(w_a121_0[1]),.din(a[121]));
	jspl3 jspl3_w_a122_0(.douta(w_a122_0[0]),.doutb(w_a122_0[1]),.doutc(w_a122_0[2]),.din(a[122]));
	jspl jspl_w_a123_0(.douta(w_a123_0[0]),.doutb(w_a123_0[1]),.din(a[123]));
	jspl3 jspl3_w_a124_0(.douta(w_a124_0[0]),.doutb(w_a124_0[1]),.doutc(w_a124_0[2]),.din(a[124]));
	jspl jspl_w_a124_1(.douta(w_a124_1[0]),.doutb(w_a124_1[1]),.din(w_a124_0[0]));
	jspl3 jspl3_w_a125_0(.douta(w_a125_0[0]),.doutb(w_a125_0[1]),.doutc(w_a125_0[2]),.din(a[125]));
	jspl3 jspl3_w_a126_0(.douta(w_a126_0[0]),.doutb(w_a126_0[1]),.doutc(w_a126_0[2]),.din(a[126]));
	jspl jspl_w_a126_1(.douta(w_a126_1[0]),.doutb(w_a126_1[1]),.din(w_a126_0[0]));
	jspl jspl_w_a127_0(.douta(w_a127_0[0]),.doutb(w_a127_0[1]),.din(a[127]));
	jspl3 jspl3_w_asqrt1_0(.douta(w_asqrt1_0[0]),.doutb(w_asqrt1_0[1]),.doutc(w_asqrt1_0[2]),.din(asqrt_fa_1));
	jspl jspl_w_asqrt1_1(.douta(w_asqrt1_1),.doutb(asqrt[0]),.din(w_asqrt1_0[0]));
	jspl3 jspl3_w_asqrt2_0(.douta(w_asqrt2_0[0]),.doutb(w_asqrt2_0[1]),.doutc(w_asqrt2_0[2]),.din(asqrt_fa_2));
	jspl3 jspl3_w_asqrt2_1(.douta(w_asqrt2_1[0]),.doutb(w_asqrt2_1[1]),.doutc(w_asqrt2_1[2]),.din(w_asqrt2_0[0]));
	jspl3 jspl3_w_asqrt2_2(.douta(w_asqrt2_2[0]),.doutb(w_asqrt2_2[1]),.doutc(w_asqrt2_2[2]),.din(w_asqrt2_0[1]));
	jspl3 jspl3_w_asqrt2_3(.douta(w_asqrt2_3[0]),.doutb(w_asqrt2_3[1]),.doutc(w_asqrt2_3[2]),.din(w_asqrt2_0[2]));
	jspl3 jspl3_w_asqrt2_4(.douta(w_asqrt2_4[0]),.doutb(w_asqrt2_4[1]),.doutc(w_asqrt2_4[2]),.din(w_asqrt2_1[0]));
	jspl3 jspl3_w_asqrt2_5(.douta(w_asqrt2_5[0]),.doutb(w_asqrt2_5[1]),.doutc(w_asqrt2_5[2]),.din(w_asqrt2_1[1]));
	jspl3 jspl3_w_asqrt2_6(.douta(w_asqrt2_6[0]),.doutb(w_asqrt2_6[1]),.doutc(w_asqrt2_6[2]),.din(w_asqrt2_1[2]));
	jspl3 jspl3_w_asqrt2_7(.douta(w_asqrt2_7[0]),.doutb(w_asqrt2_7[1]),.doutc(w_asqrt2_7[2]),.din(w_asqrt2_2[0]));
	jspl3 jspl3_w_asqrt2_8(.douta(w_asqrt2_8[0]),.doutb(w_asqrt2_8[1]),.doutc(w_asqrt2_8[2]),.din(w_asqrt2_2[1]));
	jspl3 jspl3_w_asqrt2_9(.douta(w_asqrt2_9[0]),.doutb(w_asqrt2_9[1]),.doutc(w_asqrt2_9[2]),.din(w_asqrt2_2[2]));
	jspl3 jspl3_w_asqrt2_10(.douta(w_asqrt2_10[0]),.doutb(w_asqrt2_10[1]),.doutc(w_asqrt2_10[2]),.din(w_asqrt2_3[0]));
	jspl3 jspl3_w_asqrt2_11(.douta(w_asqrt2_11[0]),.doutb(w_asqrt2_11[1]),.doutc(w_asqrt2_11[2]),.din(w_asqrt2_3[1]));
	jspl3 jspl3_w_asqrt2_12(.douta(w_asqrt2_12[0]),.doutb(w_asqrt2_12[1]),.doutc(w_asqrt2_12[2]),.din(w_asqrt2_3[2]));
	jspl3 jspl3_w_asqrt2_13(.douta(w_asqrt2_13[0]),.doutb(w_asqrt2_13[1]),.doutc(w_asqrt2_13[2]),.din(w_asqrt2_4[0]));
	jspl3 jspl3_w_asqrt2_14(.douta(w_asqrt2_14[0]),.doutb(w_asqrt2_14[1]),.doutc(w_asqrt2_14[2]),.din(w_asqrt2_4[1]));
	jspl3 jspl3_w_asqrt2_15(.douta(w_asqrt2_15[0]),.doutb(w_asqrt2_15[1]),.doutc(w_asqrt2_15[2]),.din(w_asqrt2_4[2]));
	jspl3 jspl3_w_asqrt2_16(.douta(w_asqrt2_16[0]),.doutb(w_asqrt2_16[1]),.doutc(w_asqrt2_16[2]),.din(w_asqrt2_5[0]));
	jspl3 jspl3_w_asqrt2_17(.douta(w_asqrt2_17[0]),.doutb(w_asqrt2_17[1]),.doutc(w_asqrt2_17[2]),.din(w_asqrt2_5[1]));
	jspl3 jspl3_w_asqrt2_18(.douta(w_asqrt2_18[0]),.doutb(w_asqrt2_18[1]),.doutc(w_asqrt2_18[2]),.din(w_asqrt2_5[2]));
	jspl3 jspl3_w_asqrt2_19(.douta(w_asqrt2_19[0]),.doutb(w_asqrt2_19[1]),.doutc(w_asqrt2_19[2]),.din(w_asqrt2_6[0]));
	jspl3 jspl3_w_asqrt2_20(.douta(w_asqrt2_20[0]),.doutb(w_asqrt2_20[1]),.doutc(w_asqrt2_20[2]),.din(w_asqrt2_6[1]));
	jspl3 jspl3_w_asqrt2_21(.douta(w_asqrt2_21[0]),.doutb(w_asqrt2_21[1]),.doutc(w_asqrt2_21[2]),.din(w_asqrt2_6[2]));
	jspl3 jspl3_w_asqrt2_22(.douta(w_asqrt2_22[0]),.doutb(w_asqrt2_22[1]),.doutc(w_asqrt2_22[2]),.din(w_asqrt2_7[0]));
	jspl3 jspl3_w_asqrt2_23(.douta(w_asqrt2_23[0]),.doutb(w_asqrt2_23[1]),.doutc(w_asqrt2_23[2]),.din(w_asqrt2_7[1]));
	jspl3 jspl3_w_asqrt2_24(.douta(w_asqrt2_24[0]),.doutb(w_asqrt2_24[1]),.doutc(w_asqrt2_24[2]),.din(w_asqrt2_7[2]));
	jspl3 jspl3_w_asqrt2_25(.douta(w_asqrt2_25[0]),.doutb(w_asqrt2_25[1]),.doutc(w_asqrt2_25[2]),.din(w_asqrt2_8[0]));
	jspl3 jspl3_w_asqrt2_26(.douta(w_asqrt2_26[0]),.doutb(w_asqrt2_26[1]),.doutc(w_asqrt2_26[2]),.din(w_asqrt2_8[1]));
	jspl3 jspl3_w_asqrt2_27(.douta(w_asqrt2_27[0]),.doutb(w_asqrt2_27[1]),.doutc(w_asqrt2_27[2]),.din(w_asqrt2_8[2]));
	jspl3 jspl3_w_asqrt2_28(.douta(w_asqrt2_28[0]),.doutb(w_asqrt2_28[1]),.doutc(w_asqrt2_28[2]),.din(w_asqrt2_9[0]));
	jspl3 jspl3_w_asqrt2_29(.douta(w_asqrt2_29[0]),.doutb(w_asqrt2_29[1]),.doutc(w_asqrt2_29[2]),.din(w_asqrt2_9[1]));
	jspl3 jspl3_w_asqrt2_30(.douta(w_asqrt2_30[0]),.doutb(w_asqrt2_30[1]),.doutc(w_asqrt2_30[2]),.din(w_asqrt2_9[2]));
	jspl3 jspl3_w_asqrt2_31(.douta(w_asqrt2_31[0]),.doutb(w_asqrt2_31[1]),.doutc(asqrt[1]),.din(w_asqrt2_10[0]));
	jspl3 jspl3_w_asqrt3_0(.douta(w_asqrt3_0[0]),.doutb(w_asqrt3_0[1]),.doutc(w_asqrt3_0[2]),.din(asqrt_fa_3));
	jspl3 jspl3_w_asqrt3_1(.douta(w_asqrt3_1[0]),.doutb(w_asqrt3_1[1]),.doutc(w_asqrt3_1[2]),.din(w_asqrt3_0[0]));
	jspl3 jspl3_w_asqrt3_2(.douta(w_asqrt3_2[0]),.doutb(w_asqrt3_2[1]),.doutc(asqrt[2]),.din(w_asqrt3_0[1]));
	jspl3 jspl3_w_asqrt4_0(.douta(w_asqrt4_0[0]),.doutb(w_asqrt4_0[1]),.doutc(w_asqrt4_0[2]),.din(asqrt_fa_4));
	jspl3 jspl3_w_asqrt4_1(.douta(w_asqrt4_1[0]),.doutb(w_asqrt4_1[1]),.doutc(w_asqrt4_1[2]),.din(w_asqrt4_0[0]));
	jspl3 jspl3_w_asqrt4_2(.douta(w_asqrt4_2[0]),.doutb(w_asqrt4_2[1]),.doutc(w_asqrt4_2[2]),.din(w_asqrt4_0[1]));
	jspl3 jspl3_w_asqrt4_3(.douta(w_asqrt4_3[0]),.doutb(w_asqrt4_3[1]),.doutc(w_asqrt4_3[2]),.din(w_asqrt4_0[2]));
	jspl3 jspl3_w_asqrt4_4(.douta(w_asqrt4_4[0]),.doutb(w_asqrt4_4[1]),.doutc(w_asqrt4_4[2]),.din(w_asqrt4_1[0]));
	jspl3 jspl3_w_asqrt4_5(.douta(w_asqrt4_5[0]),.doutb(w_asqrt4_5[1]),.doutc(w_asqrt4_5[2]),.din(w_asqrt4_1[1]));
	jspl3 jspl3_w_asqrt4_6(.douta(w_asqrt4_6[0]),.doutb(w_asqrt4_6[1]),.doutc(w_asqrt4_6[2]),.din(w_asqrt4_1[2]));
	jspl3 jspl3_w_asqrt4_7(.douta(w_asqrt4_7[0]),.doutb(w_asqrt4_7[1]),.doutc(w_asqrt4_7[2]),.din(w_asqrt4_2[0]));
	jspl3 jspl3_w_asqrt4_8(.douta(w_asqrt4_8[0]),.doutb(w_asqrt4_8[1]),.doutc(w_asqrt4_8[2]),.din(w_asqrt4_2[1]));
	jspl3 jspl3_w_asqrt4_9(.douta(w_asqrt4_9[0]),.doutb(w_asqrt4_9[1]),.doutc(w_asqrt4_9[2]),.din(w_asqrt4_2[2]));
	jspl3 jspl3_w_asqrt4_10(.douta(w_asqrt4_10[0]),.doutb(w_asqrt4_10[1]),.doutc(w_asqrt4_10[2]),.din(w_asqrt4_3[0]));
	jspl3 jspl3_w_asqrt4_11(.douta(w_asqrt4_11[0]),.doutb(w_asqrt4_11[1]),.doutc(w_asqrt4_11[2]),.din(w_asqrt4_3[1]));
	jspl3 jspl3_w_asqrt4_12(.douta(w_asqrt4_12[0]),.doutb(w_asqrt4_12[1]),.doutc(w_asqrt4_12[2]),.din(w_asqrt4_3[2]));
	jspl3 jspl3_w_asqrt4_13(.douta(w_asqrt4_13[0]),.doutb(w_asqrt4_13[1]),.doutc(w_asqrt4_13[2]),.din(w_asqrt4_4[0]));
	jspl3 jspl3_w_asqrt4_14(.douta(w_asqrt4_14[0]),.doutb(w_asqrt4_14[1]),.doutc(w_asqrt4_14[2]),.din(w_asqrt4_4[1]));
	jspl3 jspl3_w_asqrt4_15(.douta(w_asqrt4_15[0]),.doutb(w_asqrt4_15[1]),.doutc(w_asqrt4_15[2]),.din(w_asqrt4_4[2]));
	jspl3 jspl3_w_asqrt4_16(.douta(w_asqrt4_16[0]),.doutb(w_asqrt4_16[1]),.doutc(w_asqrt4_16[2]),.din(w_asqrt4_5[0]));
	jspl3 jspl3_w_asqrt4_17(.douta(w_asqrt4_17[0]),.doutb(w_asqrt4_17[1]),.doutc(w_asqrt4_17[2]),.din(w_asqrt4_5[1]));
	jspl3 jspl3_w_asqrt4_18(.douta(w_asqrt4_18[0]),.doutb(w_asqrt4_18[1]),.doutc(w_asqrt4_18[2]),.din(w_asqrt4_5[2]));
	jspl3 jspl3_w_asqrt4_19(.douta(w_asqrt4_19[0]),.doutb(w_asqrt4_19[1]),.doutc(w_asqrt4_19[2]),.din(w_asqrt4_6[0]));
	jspl3 jspl3_w_asqrt4_20(.douta(w_asqrt4_20[0]),.doutb(w_asqrt4_20[1]),.doutc(w_asqrt4_20[2]),.din(w_asqrt4_6[1]));
	jspl3 jspl3_w_asqrt4_21(.douta(w_asqrt4_21[0]),.doutb(w_asqrt4_21[1]),.doutc(w_asqrt4_21[2]),.din(w_asqrt4_6[2]));
	jspl3 jspl3_w_asqrt4_22(.douta(w_asqrt4_22[0]),.doutb(w_asqrt4_22[1]),.doutc(w_asqrt4_22[2]),.din(w_asqrt4_7[0]));
	jspl3 jspl3_w_asqrt4_23(.douta(w_asqrt4_23[0]),.doutb(w_asqrt4_23[1]),.doutc(w_asqrt4_23[2]),.din(w_asqrt4_7[1]));
	jspl3 jspl3_w_asqrt4_24(.douta(w_asqrt4_24[0]),.doutb(w_asqrt4_24[1]),.doutc(w_asqrt4_24[2]),.din(w_asqrt4_7[2]));
	jspl3 jspl3_w_asqrt4_25(.douta(w_asqrt4_25[0]),.doutb(w_asqrt4_25[1]),.doutc(w_asqrt4_25[2]),.din(w_asqrt4_8[0]));
	jspl3 jspl3_w_asqrt4_26(.douta(w_asqrt4_26[0]),.doutb(w_asqrt4_26[1]),.doutc(w_asqrt4_26[2]),.din(w_asqrt4_8[1]));
	jspl3 jspl3_w_asqrt4_27(.douta(w_asqrt4_27[0]),.doutb(w_asqrt4_27[1]),.doutc(w_asqrt4_27[2]),.din(w_asqrt4_8[2]));
	jspl3 jspl3_w_asqrt4_28(.douta(w_asqrt4_28[0]),.doutb(w_asqrt4_28[1]),.doutc(w_asqrt4_28[2]),.din(w_asqrt4_9[0]));
	jspl3 jspl3_w_asqrt4_29(.douta(w_asqrt4_29[0]),.doutb(w_asqrt4_29[1]),.doutc(w_asqrt4_29[2]),.din(w_asqrt4_9[1]));
	jspl3 jspl3_w_asqrt4_30(.douta(w_asqrt4_30[0]),.doutb(w_asqrt4_30[1]),.doutc(w_asqrt4_30[2]),.din(w_asqrt4_9[2]));
	jspl3 jspl3_w_asqrt4_31(.douta(w_asqrt4_31[0]),.doutb(w_asqrt4_31[1]),.doutc(asqrt[3]),.din(w_asqrt4_10[0]));
	jspl3 jspl3_w_asqrt5_0(.douta(w_asqrt5_0[0]),.doutb(w_asqrt5_0[1]),.doutc(w_asqrt5_0[2]),.din(asqrt_fa_5));
	jspl3 jspl3_w_asqrt5_1(.douta(w_asqrt5_1[0]),.doutb(w_asqrt5_1[1]),.doutc(w_asqrt5_1[2]),.din(w_asqrt5_0[0]));
	jspl3 jspl3_w_asqrt5_2(.douta(w_asqrt5_2[0]),.doutb(w_asqrt5_2[1]),.doutc(w_asqrt5_2[2]),.din(w_asqrt5_0[1]));
	jspl3 jspl3_w_asqrt5_3(.douta(w_asqrt5_3[0]),.doutb(w_asqrt5_3[1]),.doutc(w_asqrt5_3[2]),.din(w_asqrt5_0[2]));
	jspl3 jspl3_w_asqrt5_4(.douta(w_asqrt5_4[0]),.doutb(w_asqrt5_4[1]),.doutc(asqrt[4]),.din(w_asqrt5_1[0]));
	jspl3 jspl3_w_asqrt6_0(.douta(w_asqrt6_0[0]),.doutb(w_asqrt6_0[1]),.doutc(w_asqrt6_0[2]),.din(asqrt_fa_6));
	jspl3 jspl3_w_asqrt6_1(.douta(w_asqrt6_1[0]),.doutb(w_asqrt6_1[1]),.doutc(w_asqrt6_1[2]),.din(w_asqrt6_0[0]));
	jspl3 jspl3_w_asqrt6_2(.douta(w_asqrt6_2[0]),.doutb(w_asqrt6_2[1]),.doutc(w_asqrt6_2[2]),.din(w_asqrt6_0[1]));
	jspl3 jspl3_w_asqrt6_3(.douta(w_asqrt6_3[0]),.doutb(w_asqrt6_3[1]),.doutc(w_asqrt6_3[2]),.din(w_asqrt6_0[2]));
	jspl3 jspl3_w_asqrt6_4(.douta(w_asqrt6_4[0]),.doutb(w_asqrt6_4[1]),.doutc(w_asqrt6_4[2]),.din(w_asqrt6_1[0]));
	jspl3 jspl3_w_asqrt6_5(.douta(w_asqrt6_5[0]),.doutb(w_asqrt6_5[1]),.doutc(w_asqrt6_5[2]),.din(w_asqrt6_1[1]));
	jspl3 jspl3_w_asqrt6_6(.douta(w_asqrt6_6[0]),.doutb(w_asqrt6_6[1]),.doutc(w_asqrt6_6[2]),.din(w_asqrt6_1[2]));
	jspl3 jspl3_w_asqrt6_7(.douta(w_asqrt6_7[0]),.doutb(w_asqrt6_7[1]),.doutc(w_asqrt6_7[2]),.din(w_asqrt6_2[0]));
	jspl3 jspl3_w_asqrt6_8(.douta(w_asqrt6_8[0]),.doutb(w_asqrt6_8[1]),.doutc(w_asqrt6_8[2]),.din(w_asqrt6_2[1]));
	jspl3 jspl3_w_asqrt6_9(.douta(w_asqrt6_9[0]),.doutb(w_asqrt6_9[1]),.doutc(w_asqrt6_9[2]),.din(w_asqrt6_2[2]));
	jspl3 jspl3_w_asqrt6_10(.douta(w_asqrt6_10[0]),.doutb(w_asqrt6_10[1]),.doutc(w_asqrt6_10[2]),.din(w_asqrt6_3[0]));
	jspl3 jspl3_w_asqrt6_11(.douta(w_asqrt6_11[0]),.doutb(w_asqrt6_11[1]),.doutc(w_asqrt6_11[2]),.din(w_asqrt6_3[1]));
	jspl3 jspl3_w_asqrt6_12(.douta(w_asqrt6_12[0]),.doutb(w_asqrt6_12[1]),.doutc(w_asqrt6_12[2]),.din(w_asqrt6_3[2]));
	jspl3 jspl3_w_asqrt6_13(.douta(w_asqrt6_13[0]),.doutb(w_asqrt6_13[1]),.doutc(w_asqrt6_13[2]),.din(w_asqrt6_4[0]));
	jspl3 jspl3_w_asqrt6_14(.douta(w_asqrt6_14[0]),.doutb(w_asqrt6_14[1]),.doutc(w_asqrt6_14[2]),.din(w_asqrt6_4[1]));
	jspl3 jspl3_w_asqrt6_15(.douta(w_asqrt6_15[0]),.doutb(w_asqrt6_15[1]),.doutc(w_asqrt6_15[2]),.din(w_asqrt6_4[2]));
	jspl3 jspl3_w_asqrt6_16(.douta(w_asqrt6_16[0]),.doutb(w_asqrt6_16[1]),.doutc(w_asqrt6_16[2]),.din(w_asqrt6_5[0]));
	jspl3 jspl3_w_asqrt6_17(.douta(w_asqrt6_17[0]),.doutb(w_asqrt6_17[1]),.doutc(w_asqrt6_17[2]),.din(w_asqrt6_5[1]));
	jspl3 jspl3_w_asqrt6_18(.douta(w_asqrt6_18[0]),.doutb(w_asqrt6_18[1]),.doutc(w_asqrt6_18[2]),.din(w_asqrt6_5[2]));
	jspl3 jspl3_w_asqrt6_19(.douta(w_asqrt6_19[0]),.doutb(w_asqrt6_19[1]),.doutc(w_asqrt6_19[2]),.din(w_asqrt6_6[0]));
	jspl3 jspl3_w_asqrt6_20(.douta(w_asqrt6_20[0]),.doutb(w_asqrt6_20[1]),.doutc(w_asqrt6_20[2]),.din(w_asqrt6_6[1]));
	jspl3 jspl3_w_asqrt6_21(.douta(w_asqrt6_21[0]),.doutb(w_asqrt6_21[1]),.doutc(w_asqrt6_21[2]),.din(w_asqrt6_6[2]));
	jspl3 jspl3_w_asqrt6_22(.douta(w_asqrt6_22[0]),.doutb(w_asqrt6_22[1]),.doutc(w_asqrt6_22[2]),.din(w_asqrt6_7[0]));
	jspl3 jspl3_w_asqrt6_23(.douta(w_asqrt6_23[0]),.doutb(w_asqrt6_23[1]),.doutc(w_asqrt6_23[2]),.din(w_asqrt6_7[1]));
	jspl3 jspl3_w_asqrt6_24(.douta(w_asqrt6_24[0]),.doutb(w_asqrt6_24[1]),.doutc(w_asqrt6_24[2]),.din(w_asqrt6_7[2]));
	jspl3 jspl3_w_asqrt6_25(.douta(w_asqrt6_25[0]),.doutb(w_asqrt6_25[1]),.doutc(w_asqrt6_25[2]),.din(w_asqrt6_8[0]));
	jspl3 jspl3_w_asqrt6_26(.douta(w_asqrt6_26[0]),.doutb(w_asqrt6_26[1]),.doutc(w_asqrt6_26[2]),.din(w_asqrt6_8[1]));
	jspl3 jspl3_w_asqrt6_27(.douta(w_asqrt6_27[0]),.doutb(w_asqrt6_27[1]),.doutc(w_asqrt6_27[2]),.din(w_asqrt6_8[2]));
	jspl3 jspl3_w_asqrt6_28(.douta(w_asqrt6_28[0]),.doutb(w_asqrt6_28[1]),.doutc(w_asqrt6_28[2]),.din(w_asqrt6_9[0]));
	jspl3 jspl3_w_asqrt6_29(.douta(w_asqrt6_29[0]),.doutb(w_asqrt6_29[1]),.doutc(w_asqrt6_29[2]),.din(w_asqrt6_9[1]));
	jspl3 jspl3_w_asqrt6_30(.douta(w_asqrt6_30[0]),.doutb(w_asqrt6_30[1]),.doutc(w_asqrt6_30[2]),.din(w_asqrt6_9[2]));
	jspl3 jspl3_w_asqrt6_31(.douta(w_asqrt6_31[0]),.doutb(w_asqrt6_31[1]),.doutc(w_asqrt6_31[2]),.din(w_asqrt6_10[0]));
	jspl jspl_w_asqrt6_32(.douta(w_asqrt6_32),.doutb(asqrt[5]),.din(w_asqrt6_10[1]));
	jspl3 jspl3_w_asqrt7_0(.douta(w_asqrt7_0[0]),.doutb(w_asqrt7_0[1]),.doutc(w_asqrt7_0[2]),.din(asqrt_fa_7));
	jspl3 jspl3_w_asqrt7_1(.douta(w_asqrt7_1[0]),.doutb(w_asqrt7_1[1]),.doutc(w_asqrt7_1[2]),.din(w_asqrt7_0[0]));
	jspl3 jspl3_w_asqrt7_2(.douta(w_asqrt7_2[0]),.doutb(w_asqrt7_2[1]),.doutc(w_asqrt7_2[2]),.din(w_asqrt7_0[1]));
	jspl3 jspl3_w_asqrt7_3(.douta(w_asqrt7_3[0]),.doutb(w_asqrt7_3[1]),.doutc(w_asqrt7_3[2]),.din(w_asqrt7_0[2]));
	jspl3 jspl3_w_asqrt7_4(.douta(w_asqrt7_4[0]),.doutb(w_asqrt7_4[1]),.doutc(w_asqrt7_4[2]),.din(w_asqrt7_1[0]));
	jspl3 jspl3_w_asqrt7_5(.douta(w_asqrt7_5[0]),.doutb(w_asqrt7_5[1]),.doutc(w_asqrt7_5[2]),.din(w_asqrt7_1[1]));
	jspl jspl_w_asqrt7_6(.douta(w_asqrt7_6),.doutb(asqrt[6]),.din(w_asqrt7_1[2]));
	jspl3 jspl3_w_asqrt8_0(.douta(w_asqrt8_0[0]),.doutb(w_asqrt8_0[1]),.doutc(w_asqrt8_0[2]),.din(asqrt_fa_8));
	jspl3 jspl3_w_asqrt8_1(.douta(w_asqrt8_1[0]),.doutb(w_asqrt8_1[1]),.doutc(w_asqrt8_1[2]),.din(w_asqrt8_0[0]));
	jspl3 jspl3_w_asqrt8_2(.douta(w_asqrt8_2[0]),.doutb(w_asqrt8_2[1]),.doutc(w_asqrt8_2[2]),.din(w_asqrt8_0[1]));
	jspl3 jspl3_w_asqrt8_3(.douta(w_asqrt8_3[0]),.doutb(w_asqrt8_3[1]),.doutc(w_asqrt8_3[2]),.din(w_asqrt8_0[2]));
	jspl3 jspl3_w_asqrt8_4(.douta(w_asqrt8_4[0]),.doutb(w_asqrt8_4[1]),.doutc(w_asqrt8_4[2]),.din(w_asqrt8_1[0]));
	jspl3 jspl3_w_asqrt8_5(.douta(w_asqrt8_5[0]),.doutb(w_asqrt8_5[1]),.doutc(w_asqrt8_5[2]),.din(w_asqrt8_1[1]));
	jspl3 jspl3_w_asqrt8_6(.douta(w_asqrt8_6[0]),.doutb(w_asqrt8_6[1]),.doutc(w_asqrt8_6[2]),.din(w_asqrt8_1[2]));
	jspl3 jspl3_w_asqrt8_7(.douta(w_asqrt8_7[0]),.doutb(w_asqrt8_7[1]),.doutc(w_asqrt8_7[2]),.din(w_asqrt8_2[0]));
	jspl3 jspl3_w_asqrt8_8(.douta(w_asqrt8_8[0]),.doutb(w_asqrt8_8[1]),.doutc(w_asqrt8_8[2]),.din(w_asqrt8_2[1]));
	jspl3 jspl3_w_asqrt8_9(.douta(w_asqrt8_9[0]),.doutb(w_asqrt8_9[1]),.doutc(w_asqrt8_9[2]),.din(w_asqrt8_2[2]));
	jspl3 jspl3_w_asqrt8_10(.douta(w_asqrt8_10[0]),.doutb(w_asqrt8_10[1]),.doutc(w_asqrt8_10[2]),.din(w_asqrt8_3[0]));
	jspl3 jspl3_w_asqrt8_11(.douta(w_asqrt8_11[0]),.doutb(w_asqrt8_11[1]),.doutc(w_asqrt8_11[2]),.din(w_asqrt8_3[1]));
	jspl3 jspl3_w_asqrt8_12(.douta(w_asqrt8_12[0]),.doutb(w_asqrt8_12[1]),.doutc(w_asqrt8_12[2]),.din(w_asqrt8_3[2]));
	jspl3 jspl3_w_asqrt8_13(.douta(w_asqrt8_13[0]),.doutb(w_asqrt8_13[1]),.doutc(w_asqrt8_13[2]),.din(w_asqrt8_4[0]));
	jspl3 jspl3_w_asqrt8_14(.douta(w_asqrt8_14[0]),.doutb(w_asqrt8_14[1]),.doutc(w_asqrt8_14[2]),.din(w_asqrt8_4[1]));
	jspl3 jspl3_w_asqrt8_15(.douta(w_asqrt8_15[0]),.doutb(w_asqrt8_15[1]),.doutc(w_asqrt8_15[2]),.din(w_asqrt8_4[2]));
	jspl3 jspl3_w_asqrt8_16(.douta(w_asqrt8_16[0]),.doutb(w_asqrt8_16[1]),.doutc(w_asqrt8_16[2]),.din(w_asqrt8_5[0]));
	jspl3 jspl3_w_asqrt8_17(.douta(w_asqrt8_17[0]),.doutb(w_asqrt8_17[1]),.doutc(w_asqrt8_17[2]),.din(w_asqrt8_5[1]));
	jspl3 jspl3_w_asqrt8_18(.douta(w_asqrt8_18[0]),.doutb(w_asqrt8_18[1]),.doutc(w_asqrt8_18[2]),.din(w_asqrt8_5[2]));
	jspl3 jspl3_w_asqrt8_19(.douta(w_asqrt8_19[0]),.doutb(w_asqrt8_19[1]),.doutc(w_asqrt8_19[2]),.din(w_asqrt8_6[0]));
	jspl3 jspl3_w_asqrt8_20(.douta(w_asqrt8_20[0]),.doutb(w_asqrt8_20[1]),.doutc(w_asqrt8_20[2]),.din(w_asqrt8_6[1]));
	jspl3 jspl3_w_asqrt8_21(.douta(w_asqrt8_21[0]),.doutb(w_asqrt8_21[1]),.doutc(w_asqrt8_21[2]),.din(w_asqrt8_6[2]));
	jspl3 jspl3_w_asqrt8_22(.douta(w_asqrt8_22[0]),.doutb(w_asqrt8_22[1]),.doutc(w_asqrt8_22[2]),.din(w_asqrt8_7[0]));
	jspl3 jspl3_w_asqrt8_23(.douta(w_asqrt8_23[0]),.doutb(w_asqrt8_23[1]),.doutc(w_asqrt8_23[2]),.din(w_asqrt8_7[1]));
	jspl3 jspl3_w_asqrt8_24(.douta(w_asqrt8_24[0]),.doutb(w_asqrt8_24[1]),.doutc(w_asqrt8_24[2]),.din(w_asqrt8_7[2]));
	jspl3 jspl3_w_asqrt8_25(.douta(w_asqrt8_25[0]),.doutb(w_asqrt8_25[1]),.doutc(w_asqrt8_25[2]),.din(w_asqrt8_8[0]));
	jspl3 jspl3_w_asqrt8_26(.douta(w_asqrt8_26[0]),.doutb(w_asqrt8_26[1]),.doutc(w_asqrt8_26[2]),.din(w_asqrt8_8[1]));
	jspl3 jspl3_w_asqrt8_27(.douta(w_asqrt8_27[0]),.doutb(w_asqrt8_27[1]),.doutc(w_asqrt8_27[2]),.din(w_asqrt8_8[2]));
	jspl3 jspl3_w_asqrt8_28(.douta(w_asqrt8_28[0]),.doutb(w_asqrt8_28[1]),.doutc(w_asqrt8_28[2]),.din(w_asqrt8_9[0]));
	jspl3 jspl3_w_asqrt8_29(.douta(w_asqrt8_29[0]),.doutb(w_asqrt8_29[1]),.doutc(w_asqrt8_29[2]),.din(w_asqrt8_9[1]));
	jspl3 jspl3_w_asqrt8_30(.douta(w_asqrt8_30[0]),.doutb(w_asqrt8_30[1]),.doutc(w_asqrt8_30[2]),.din(w_asqrt8_9[2]));
	jspl3 jspl3_w_asqrt8_31(.douta(w_asqrt8_31[0]),.doutb(w_asqrt8_31[1]),.doutc(w_asqrt8_31[2]),.din(w_asqrt8_10[0]));
	jspl3 jspl3_w_asqrt8_32(.douta(w_asqrt8_32[0]),.doutb(w_asqrt8_32[1]),.doutc(asqrt[7]),.din(w_asqrt8_10[1]));
	jspl3 jspl3_w_asqrt9_0(.douta(w_asqrt9_0[0]),.doutb(w_asqrt9_0[1]),.doutc(w_asqrt9_0[2]),.din(asqrt_fa_9));
	jspl3 jspl3_w_asqrt9_1(.douta(w_asqrt9_1[0]),.doutb(w_asqrt9_1[1]),.doutc(w_asqrt9_1[2]),.din(w_asqrt9_0[0]));
	jspl3 jspl3_w_asqrt9_2(.douta(w_asqrt9_2[0]),.doutb(w_asqrt9_2[1]),.doutc(w_asqrt9_2[2]),.din(w_asqrt9_0[1]));
	jspl3 jspl3_w_asqrt9_3(.douta(w_asqrt9_3[0]),.doutb(w_asqrt9_3[1]),.doutc(w_asqrt9_3[2]),.din(w_asqrt9_0[2]));
	jspl3 jspl3_w_asqrt9_4(.douta(w_asqrt9_4[0]),.doutb(w_asqrt9_4[1]),.doutc(w_asqrt9_4[2]),.din(w_asqrt9_1[0]));
	jspl3 jspl3_w_asqrt9_5(.douta(w_asqrt9_5[0]),.doutb(w_asqrt9_5[1]),.doutc(w_asqrt9_5[2]),.din(w_asqrt9_1[1]));
	jspl3 jspl3_w_asqrt9_6(.douta(w_asqrt9_6[0]),.doutb(w_asqrt9_6[1]),.doutc(w_asqrt9_6[2]),.din(w_asqrt9_1[2]));
	jspl3 jspl3_w_asqrt9_7(.douta(w_asqrt9_7[0]),.doutb(w_asqrt9_7[1]),.doutc(w_asqrt9_7[2]),.din(w_asqrt9_2[0]));
	jspl jspl_w_asqrt9_8(.douta(w_asqrt9_8),.doutb(asqrt[8]),.din(w_asqrt9_2[1]));
	jspl3 jspl3_w_asqrt10_0(.douta(w_asqrt10_0[0]),.doutb(w_asqrt10_0[1]),.doutc(w_asqrt10_0[2]),.din(asqrt_fa_10));
	jspl3 jspl3_w_asqrt10_1(.douta(w_asqrt10_1[0]),.doutb(w_asqrt10_1[1]),.doutc(w_asqrt10_1[2]),.din(w_asqrt10_0[0]));
	jspl3 jspl3_w_asqrt10_2(.douta(w_asqrt10_2[0]),.doutb(w_asqrt10_2[1]),.doutc(w_asqrt10_2[2]),.din(w_asqrt10_0[1]));
	jspl3 jspl3_w_asqrt10_3(.douta(w_asqrt10_3[0]),.doutb(w_asqrt10_3[1]),.doutc(w_asqrt10_3[2]),.din(w_asqrt10_0[2]));
	jspl3 jspl3_w_asqrt10_4(.douta(w_asqrt10_4[0]),.doutb(w_asqrt10_4[1]),.doutc(w_asqrt10_4[2]),.din(w_asqrt10_1[0]));
	jspl3 jspl3_w_asqrt10_5(.douta(w_asqrt10_5[0]),.doutb(w_asqrt10_5[1]),.doutc(w_asqrt10_5[2]),.din(w_asqrt10_1[1]));
	jspl3 jspl3_w_asqrt10_6(.douta(w_asqrt10_6[0]),.doutb(w_asqrt10_6[1]),.doutc(w_asqrt10_6[2]),.din(w_asqrt10_1[2]));
	jspl3 jspl3_w_asqrt10_7(.douta(w_asqrt10_7[0]),.doutb(w_asqrt10_7[1]),.doutc(w_asqrt10_7[2]),.din(w_asqrt10_2[0]));
	jspl3 jspl3_w_asqrt10_8(.douta(w_asqrt10_8[0]),.doutb(w_asqrt10_8[1]),.doutc(w_asqrt10_8[2]),.din(w_asqrt10_2[1]));
	jspl3 jspl3_w_asqrt10_9(.douta(w_asqrt10_9[0]),.doutb(w_asqrt10_9[1]),.doutc(w_asqrt10_9[2]),.din(w_asqrt10_2[2]));
	jspl3 jspl3_w_asqrt10_10(.douta(w_asqrt10_10[0]),.doutb(w_asqrt10_10[1]),.doutc(w_asqrt10_10[2]),.din(w_asqrt10_3[0]));
	jspl3 jspl3_w_asqrt10_11(.douta(w_asqrt10_11[0]),.doutb(w_asqrt10_11[1]),.doutc(w_asqrt10_11[2]),.din(w_asqrt10_3[1]));
	jspl3 jspl3_w_asqrt10_12(.douta(w_asqrt10_12[0]),.doutb(w_asqrt10_12[1]),.doutc(w_asqrt10_12[2]),.din(w_asqrt10_3[2]));
	jspl3 jspl3_w_asqrt10_13(.douta(w_asqrt10_13[0]),.doutb(w_asqrt10_13[1]),.doutc(w_asqrt10_13[2]),.din(w_asqrt10_4[0]));
	jspl3 jspl3_w_asqrt10_14(.douta(w_asqrt10_14[0]),.doutb(w_asqrt10_14[1]),.doutc(w_asqrt10_14[2]),.din(w_asqrt10_4[1]));
	jspl3 jspl3_w_asqrt10_15(.douta(w_asqrt10_15[0]),.doutb(w_asqrt10_15[1]),.doutc(w_asqrt10_15[2]),.din(w_asqrt10_4[2]));
	jspl3 jspl3_w_asqrt10_16(.douta(w_asqrt10_16[0]),.doutb(w_asqrt10_16[1]),.doutc(w_asqrt10_16[2]),.din(w_asqrt10_5[0]));
	jspl3 jspl3_w_asqrt10_17(.douta(w_asqrt10_17[0]),.doutb(w_asqrt10_17[1]),.doutc(w_asqrt10_17[2]),.din(w_asqrt10_5[1]));
	jspl3 jspl3_w_asqrt10_18(.douta(w_asqrt10_18[0]),.doutb(w_asqrt10_18[1]),.doutc(w_asqrt10_18[2]),.din(w_asqrt10_5[2]));
	jspl3 jspl3_w_asqrt10_19(.douta(w_asqrt10_19[0]),.doutb(w_asqrt10_19[1]),.doutc(w_asqrt10_19[2]),.din(w_asqrt10_6[0]));
	jspl3 jspl3_w_asqrt10_20(.douta(w_asqrt10_20[0]),.doutb(w_asqrt10_20[1]),.doutc(w_asqrt10_20[2]),.din(w_asqrt10_6[1]));
	jspl3 jspl3_w_asqrt10_21(.douta(w_asqrt10_21[0]),.doutb(w_asqrt10_21[1]),.doutc(w_asqrt10_21[2]),.din(w_asqrt10_6[2]));
	jspl3 jspl3_w_asqrt10_22(.douta(w_asqrt10_22[0]),.doutb(w_asqrt10_22[1]),.doutc(w_asqrt10_22[2]),.din(w_asqrt10_7[0]));
	jspl3 jspl3_w_asqrt10_23(.douta(w_asqrt10_23[0]),.doutb(w_asqrt10_23[1]),.doutc(w_asqrt10_23[2]),.din(w_asqrt10_7[1]));
	jspl3 jspl3_w_asqrt10_24(.douta(w_asqrt10_24[0]),.doutb(w_asqrt10_24[1]),.doutc(w_asqrt10_24[2]),.din(w_asqrt10_7[2]));
	jspl3 jspl3_w_asqrt10_25(.douta(w_asqrt10_25[0]),.doutb(w_asqrt10_25[1]),.doutc(w_asqrt10_25[2]),.din(w_asqrt10_8[0]));
	jspl3 jspl3_w_asqrt10_26(.douta(w_asqrt10_26[0]),.doutb(w_asqrt10_26[1]),.doutc(w_asqrt10_26[2]),.din(w_asqrt10_8[1]));
	jspl3 jspl3_w_asqrt10_27(.douta(w_asqrt10_27[0]),.doutb(w_asqrt10_27[1]),.doutc(w_asqrt10_27[2]),.din(w_asqrt10_8[2]));
	jspl3 jspl3_w_asqrt10_28(.douta(w_asqrt10_28[0]),.doutb(w_asqrt10_28[1]),.doutc(w_asqrt10_28[2]),.din(w_asqrt10_9[0]));
	jspl3 jspl3_w_asqrt10_29(.douta(w_asqrt10_29[0]),.doutb(w_asqrt10_29[1]),.doutc(w_asqrt10_29[2]),.din(w_asqrt10_9[1]));
	jspl3 jspl3_w_asqrt10_30(.douta(w_asqrt10_30[0]),.doutb(w_asqrt10_30[1]),.doutc(w_asqrt10_30[2]),.din(w_asqrt10_9[2]));
	jspl3 jspl3_w_asqrt10_31(.douta(w_asqrt10_31[0]),.doutb(w_asqrt10_31[1]),.doutc(w_asqrt10_31[2]),.din(w_asqrt10_10[0]));
	jspl3 jspl3_w_asqrt10_32(.douta(w_asqrt10_32[0]),.doutb(w_asqrt10_32[1]),.doutc(asqrt[9]),.din(w_asqrt10_10[1]));
	jspl3 jspl3_w_asqrt11_0(.douta(w_asqrt11_0[0]),.doutb(w_asqrt11_0[1]),.doutc(w_asqrt11_0[2]),.din(asqrt_fa_11));
	jspl3 jspl3_w_asqrt11_1(.douta(w_asqrt11_1[0]),.doutb(w_asqrt11_1[1]),.doutc(w_asqrt11_1[2]),.din(w_asqrt11_0[0]));
	jspl3 jspl3_w_asqrt11_2(.douta(w_asqrt11_2[0]),.doutb(w_asqrt11_2[1]),.doutc(w_asqrt11_2[2]),.din(w_asqrt11_0[1]));
	jspl3 jspl3_w_asqrt11_3(.douta(w_asqrt11_3[0]),.doutb(w_asqrt11_3[1]),.doutc(w_asqrt11_3[2]),.din(w_asqrt11_0[2]));
	jspl3 jspl3_w_asqrt11_4(.douta(w_asqrt11_4[0]),.doutb(w_asqrt11_4[1]),.doutc(w_asqrt11_4[2]),.din(w_asqrt11_1[0]));
	jspl3 jspl3_w_asqrt11_5(.douta(w_asqrt11_5[0]),.doutb(w_asqrt11_5[1]),.doutc(w_asqrt11_5[2]),.din(w_asqrt11_1[1]));
	jspl3 jspl3_w_asqrt11_6(.douta(w_asqrt11_6[0]),.doutb(w_asqrt11_6[1]),.doutc(w_asqrt11_6[2]),.din(w_asqrt11_1[2]));
	jspl3 jspl3_w_asqrt11_7(.douta(w_asqrt11_7[0]),.doutb(w_asqrt11_7[1]),.doutc(w_asqrt11_7[2]),.din(w_asqrt11_2[0]));
	jspl3 jspl3_w_asqrt11_8(.douta(w_asqrt11_8[0]),.doutb(w_asqrt11_8[1]),.doutc(asqrt[10]),.din(w_asqrt11_2[1]));
	jspl3 jspl3_w_asqrt12_0(.douta(w_asqrt12_0[0]),.doutb(w_asqrt12_0[1]),.doutc(w_asqrt12_0[2]),.din(asqrt_fa_12));
	jspl3 jspl3_w_asqrt12_1(.douta(w_asqrt12_1[0]),.doutb(w_asqrt12_1[1]),.doutc(w_asqrt12_1[2]),.din(w_asqrt12_0[0]));
	jspl3 jspl3_w_asqrt12_2(.douta(w_asqrt12_2[0]),.doutb(w_asqrt12_2[1]),.doutc(w_asqrt12_2[2]),.din(w_asqrt12_0[1]));
	jspl3 jspl3_w_asqrt12_3(.douta(w_asqrt12_3[0]),.doutb(w_asqrt12_3[1]),.doutc(w_asqrt12_3[2]),.din(w_asqrt12_0[2]));
	jspl3 jspl3_w_asqrt12_4(.douta(w_asqrt12_4[0]),.doutb(w_asqrt12_4[1]),.doutc(w_asqrt12_4[2]),.din(w_asqrt12_1[0]));
	jspl3 jspl3_w_asqrt12_5(.douta(w_asqrt12_5[0]),.doutb(w_asqrt12_5[1]),.doutc(w_asqrt12_5[2]),.din(w_asqrt12_1[1]));
	jspl3 jspl3_w_asqrt12_6(.douta(w_asqrt12_6[0]),.doutb(w_asqrt12_6[1]),.doutc(w_asqrt12_6[2]),.din(w_asqrt12_1[2]));
	jspl3 jspl3_w_asqrt12_7(.douta(w_asqrt12_7[0]),.doutb(w_asqrt12_7[1]),.doutc(w_asqrt12_7[2]),.din(w_asqrt12_2[0]));
	jspl3 jspl3_w_asqrt12_8(.douta(w_asqrt12_8[0]),.doutb(w_asqrt12_8[1]),.doutc(w_asqrt12_8[2]),.din(w_asqrt12_2[1]));
	jspl3 jspl3_w_asqrt12_9(.douta(w_asqrt12_9[0]),.doutb(w_asqrt12_9[1]),.doutc(w_asqrt12_9[2]),.din(w_asqrt12_2[2]));
	jspl3 jspl3_w_asqrt12_10(.douta(w_asqrt12_10[0]),.doutb(w_asqrt12_10[1]),.doutc(w_asqrt12_10[2]),.din(w_asqrt12_3[0]));
	jspl3 jspl3_w_asqrt12_11(.douta(w_asqrt12_11[0]),.doutb(w_asqrt12_11[1]),.doutc(w_asqrt12_11[2]),.din(w_asqrt12_3[1]));
	jspl3 jspl3_w_asqrt12_12(.douta(w_asqrt12_12[0]),.doutb(w_asqrt12_12[1]),.doutc(w_asqrt12_12[2]),.din(w_asqrt12_3[2]));
	jspl3 jspl3_w_asqrt12_13(.douta(w_asqrt12_13[0]),.doutb(w_asqrt12_13[1]),.doutc(w_asqrt12_13[2]),.din(w_asqrt12_4[0]));
	jspl3 jspl3_w_asqrt12_14(.douta(w_asqrt12_14[0]),.doutb(w_asqrt12_14[1]),.doutc(w_asqrt12_14[2]),.din(w_asqrt12_4[1]));
	jspl3 jspl3_w_asqrt12_15(.douta(w_asqrt12_15[0]),.doutb(w_asqrt12_15[1]),.doutc(w_asqrt12_15[2]),.din(w_asqrt12_4[2]));
	jspl3 jspl3_w_asqrt12_16(.douta(w_asqrt12_16[0]),.doutb(w_asqrt12_16[1]),.doutc(w_asqrt12_16[2]),.din(w_asqrt12_5[0]));
	jspl3 jspl3_w_asqrt12_17(.douta(w_asqrt12_17[0]),.doutb(w_asqrt12_17[1]),.doutc(w_asqrt12_17[2]),.din(w_asqrt12_5[1]));
	jspl3 jspl3_w_asqrt12_18(.douta(w_asqrt12_18[0]),.doutb(w_asqrt12_18[1]),.doutc(w_asqrt12_18[2]),.din(w_asqrt12_5[2]));
	jspl3 jspl3_w_asqrt12_19(.douta(w_asqrt12_19[0]),.doutb(w_asqrt12_19[1]),.doutc(w_asqrt12_19[2]),.din(w_asqrt12_6[0]));
	jspl3 jspl3_w_asqrt12_20(.douta(w_asqrt12_20[0]),.doutb(w_asqrt12_20[1]),.doutc(w_asqrt12_20[2]),.din(w_asqrt12_6[1]));
	jspl3 jspl3_w_asqrt12_21(.douta(w_asqrt12_21[0]),.doutb(w_asqrt12_21[1]),.doutc(w_asqrt12_21[2]),.din(w_asqrt12_6[2]));
	jspl3 jspl3_w_asqrt12_22(.douta(w_asqrt12_22[0]),.doutb(w_asqrt12_22[1]),.doutc(w_asqrt12_22[2]),.din(w_asqrt12_7[0]));
	jspl3 jspl3_w_asqrt12_23(.douta(w_asqrt12_23[0]),.doutb(w_asqrt12_23[1]),.doutc(w_asqrt12_23[2]),.din(w_asqrt12_7[1]));
	jspl3 jspl3_w_asqrt12_24(.douta(w_asqrt12_24[0]),.doutb(w_asqrt12_24[1]),.doutc(w_asqrt12_24[2]),.din(w_asqrt12_7[2]));
	jspl3 jspl3_w_asqrt12_25(.douta(w_asqrt12_25[0]),.doutb(w_asqrt12_25[1]),.doutc(w_asqrt12_25[2]),.din(w_asqrt12_8[0]));
	jspl3 jspl3_w_asqrt12_26(.douta(w_asqrt12_26[0]),.doutb(w_asqrt12_26[1]),.doutc(w_asqrt12_26[2]),.din(w_asqrt12_8[1]));
	jspl3 jspl3_w_asqrt12_27(.douta(w_asqrt12_27[0]),.doutb(w_asqrt12_27[1]),.doutc(w_asqrt12_27[2]),.din(w_asqrt12_8[2]));
	jspl3 jspl3_w_asqrt12_28(.douta(w_asqrt12_28[0]),.doutb(w_asqrt12_28[1]),.doutc(w_asqrt12_28[2]),.din(w_asqrt12_9[0]));
	jspl3 jspl3_w_asqrt12_29(.douta(w_asqrt12_29[0]),.doutb(w_asqrt12_29[1]),.doutc(w_asqrt12_29[2]),.din(w_asqrt12_9[1]));
	jspl3 jspl3_w_asqrt12_30(.douta(w_asqrt12_30[0]),.doutb(w_asqrt12_30[1]),.doutc(w_asqrt12_30[2]),.din(w_asqrt12_9[2]));
	jspl3 jspl3_w_asqrt12_31(.douta(w_asqrt12_31[0]),.doutb(w_asqrt12_31[1]),.doutc(w_asqrt12_31[2]),.din(w_asqrt12_10[0]));
	jspl3 jspl3_w_asqrt12_32(.douta(w_asqrt12_32[0]),.doutb(w_asqrt12_32[1]),.doutc(w_asqrt12_32[2]),.din(w_asqrt12_10[1]));
	jspl jspl_w_asqrt12_33(.douta(w_asqrt12_33),.doutb(asqrt[11]),.din(w_asqrt12_10[2]));
	jspl3 jspl3_w_asqrt13_0(.douta(w_asqrt13_0[0]),.doutb(w_asqrt13_0[1]),.doutc(w_asqrt13_0[2]),.din(asqrt_fa_13));
	jspl3 jspl3_w_asqrt13_1(.douta(w_asqrt13_1[0]),.doutb(w_asqrt13_1[1]),.doutc(w_asqrt13_1[2]),.din(w_asqrt13_0[0]));
	jspl3 jspl3_w_asqrt13_2(.douta(w_asqrt13_2[0]),.doutb(w_asqrt13_2[1]),.doutc(w_asqrt13_2[2]),.din(w_asqrt13_0[1]));
	jspl3 jspl3_w_asqrt13_3(.douta(w_asqrt13_3[0]),.doutb(w_asqrt13_3[1]),.doutc(w_asqrt13_3[2]),.din(w_asqrt13_0[2]));
	jspl3 jspl3_w_asqrt13_4(.douta(w_asqrt13_4[0]),.doutb(w_asqrt13_4[1]),.doutc(w_asqrt13_4[2]),.din(w_asqrt13_1[0]));
	jspl3 jspl3_w_asqrt13_5(.douta(w_asqrt13_5[0]),.doutb(w_asqrt13_5[1]),.doutc(w_asqrt13_5[2]),.din(w_asqrt13_1[1]));
	jspl3 jspl3_w_asqrt13_6(.douta(w_asqrt13_6[0]),.doutb(w_asqrt13_6[1]),.doutc(w_asqrt13_6[2]),.din(w_asqrt13_1[2]));
	jspl3 jspl3_w_asqrt13_7(.douta(w_asqrt13_7[0]),.doutb(w_asqrt13_7[1]),.doutc(w_asqrt13_7[2]),.din(w_asqrt13_2[0]));
	jspl3 jspl3_w_asqrt13_8(.douta(w_asqrt13_8[0]),.doutb(w_asqrt13_8[1]),.doutc(w_asqrt13_8[2]),.din(w_asqrt13_2[1]));
	jspl3 jspl3_w_asqrt13_9(.douta(w_asqrt13_9[0]),.doutb(w_asqrt13_9[1]),.doutc(w_asqrt13_9[2]),.din(w_asqrt13_2[2]));
	jspl3 jspl3_w_asqrt13_10(.douta(w_asqrt13_10[0]),.doutb(w_asqrt13_10[1]),.doutc(asqrt[12]),.din(w_asqrt13_3[0]));
	jspl3 jspl3_w_asqrt14_0(.douta(w_asqrt14_0[0]),.doutb(w_asqrt14_0[1]),.doutc(w_asqrt14_0[2]),.din(asqrt_fa_14));
	jspl3 jspl3_w_asqrt14_1(.douta(w_asqrt14_1[0]),.doutb(w_asqrt14_1[1]),.doutc(w_asqrt14_1[2]),.din(w_asqrt14_0[0]));
	jspl3 jspl3_w_asqrt14_2(.douta(w_asqrt14_2[0]),.doutb(w_asqrt14_2[1]),.doutc(w_asqrt14_2[2]),.din(w_asqrt14_0[1]));
	jspl3 jspl3_w_asqrt14_3(.douta(w_asqrt14_3[0]),.doutb(w_asqrt14_3[1]),.doutc(w_asqrt14_3[2]),.din(w_asqrt14_0[2]));
	jspl3 jspl3_w_asqrt14_4(.douta(w_asqrt14_4[0]),.doutb(w_asqrt14_4[1]),.doutc(w_asqrt14_4[2]),.din(w_asqrt14_1[0]));
	jspl3 jspl3_w_asqrt14_5(.douta(w_asqrt14_5[0]),.doutb(w_asqrt14_5[1]),.doutc(w_asqrt14_5[2]),.din(w_asqrt14_1[1]));
	jspl3 jspl3_w_asqrt14_6(.douta(w_asqrt14_6[0]),.doutb(w_asqrt14_6[1]),.doutc(w_asqrt14_6[2]),.din(w_asqrt14_1[2]));
	jspl3 jspl3_w_asqrt14_7(.douta(w_asqrt14_7[0]),.doutb(w_asqrt14_7[1]),.doutc(w_asqrt14_7[2]),.din(w_asqrt14_2[0]));
	jspl3 jspl3_w_asqrt14_8(.douta(w_asqrt14_8[0]),.doutb(w_asqrt14_8[1]),.doutc(w_asqrt14_8[2]),.din(w_asqrt14_2[1]));
	jspl3 jspl3_w_asqrt14_9(.douta(w_asqrt14_9[0]),.doutb(w_asqrt14_9[1]),.doutc(w_asqrt14_9[2]),.din(w_asqrt14_2[2]));
	jspl3 jspl3_w_asqrt14_10(.douta(w_asqrt14_10[0]),.doutb(w_asqrt14_10[1]),.doutc(w_asqrt14_10[2]),.din(w_asqrt14_3[0]));
	jspl3 jspl3_w_asqrt14_11(.douta(w_asqrt14_11[0]),.doutb(w_asqrt14_11[1]),.doutc(w_asqrt14_11[2]),.din(w_asqrt14_3[1]));
	jspl3 jspl3_w_asqrt14_12(.douta(w_asqrt14_12[0]),.doutb(w_asqrt14_12[1]),.doutc(w_asqrt14_12[2]),.din(w_asqrt14_3[2]));
	jspl3 jspl3_w_asqrt14_13(.douta(w_asqrt14_13[0]),.doutb(w_asqrt14_13[1]),.doutc(w_asqrt14_13[2]),.din(w_asqrt14_4[0]));
	jspl3 jspl3_w_asqrt14_14(.douta(w_asqrt14_14[0]),.doutb(w_asqrt14_14[1]),.doutc(w_asqrt14_14[2]),.din(w_asqrt14_4[1]));
	jspl3 jspl3_w_asqrt14_15(.douta(w_asqrt14_15[0]),.doutb(w_asqrt14_15[1]),.doutc(w_asqrt14_15[2]),.din(w_asqrt14_4[2]));
	jspl3 jspl3_w_asqrt14_16(.douta(w_asqrt14_16[0]),.doutb(w_asqrt14_16[1]),.doutc(w_asqrt14_16[2]),.din(w_asqrt14_5[0]));
	jspl3 jspl3_w_asqrt14_17(.douta(w_asqrt14_17[0]),.doutb(w_asqrt14_17[1]),.doutc(w_asqrt14_17[2]),.din(w_asqrt14_5[1]));
	jspl3 jspl3_w_asqrt14_18(.douta(w_asqrt14_18[0]),.doutb(w_asqrt14_18[1]),.doutc(w_asqrt14_18[2]),.din(w_asqrt14_5[2]));
	jspl3 jspl3_w_asqrt14_19(.douta(w_asqrt14_19[0]),.doutb(w_asqrt14_19[1]),.doutc(w_asqrt14_19[2]),.din(w_asqrt14_6[0]));
	jspl3 jspl3_w_asqrt14_20(.douta(w_asqrt14_20[0]),.doutb(w_asqrt14_20[1]),.doutc(w_asqrt14_20[2]),.din(w_asqrt14_6[1]));
	jspl3 jspl3_w_asqrt14_21(.douta(w_asqrt14_21[0]),.doutb(w_asqrt14_21[1]),.doutc(w_asqrt14_21[2]),.din(w_asqrt14_6[2]));
	jspl3 jspl3_w_asqrt14_22(.douta(w_asqrt14_22[0]),.doutb(w_asqrt14_22[1]),.doutc(w_asqrt14_22[2]),.din(w_asqrt14_7[0]));
	jspl3 jspl3_w_asqrt14_23(.douta(w_asqrt14_23[0]),.doutb(w_asqrt14_23[1]),.doutc(w_asqrt14_23[2]),.din(w_asqrt14_7[1]));
	jspl3 jspl3_w_asqrt14_24(.douta(w_asqrt14_24[0]),.doutb(w_asqrt14_24[1]),.doutc(w_asqrt14_24[2]),.din(w_asqrt14_7[2]));
	jspl3 jspl3_w_asqrt14_25(.douta(w_asqrt14_25[0]),.doutb(w_asqrt14_25[1]),.doutc(w_asqrt14_25[2]),.din(w_asqrt14_8[0]));
	jspl3 jspl3_w_asqrt14_26(.douta(w_asqrt14_26[0]),.doutb(w_asqrt14_26[1]),.doutc(w_asqrt14_26[2]),.din(w_asqrt14_8[1]));
	jspl3 jspl3_w_asqrt14_27(.douta(w_asqrt14_27[0]),.doutb(w_asqrt14_27[1]),.doutc(w_asqrt14_27[2]),.din(w_asqrt14_8[2]));
	jspl3 jspl3_w_asqrt14_28(.douta(w_asqrt14_28[0]),.doutb(w_asqrt14_28[1]),.doutc(w_asqrt14_28[2]),.din(w_asqrt14_9[0]));
	jspl3 jspl3_w_asqrt14_29(.douta(w_asqrt14_29[0]),.doutb(w_asqrt14_29[1]),.doutc(w_asqrt14_29[2]),.din(w_asqrt14_9[1]));
	jspl3 jspl3_w_asqrt14_30(.douta(w_asqrt14_30[0]),.doutb(w_asqrt14_30[1]),.doutc(w_asqrt14_30[2]),.din(w_asqrt14_9[2]));
	jspl3 jspl3_w_asqrt14_31(.douta(w_asqrt14_31[0]),.doutb(w_asqrt14_31[1]),.doutc(w_asqrt14_31[2]),.din(w_asqrt14_10[0]));
	jspl3 jspl3_w_asqrt14_32(.douta(w_asqrt14_32[0]),.doutb(w_asqrt14_32[1]),.doutc(w_asqrt14_32[2]),.din(w_asqrt14_10[1]));
	jspl3 jspl3_w_asqrt14_33(.douta(w_asqrt14_33[0]),.doutb(w_asqrt14_33[1]),.doutc(w_asqrt14_33[2]),.din(w_asqrt14_10[2]));
	jspl jspl_w_asqrt14_34(.douta(w_asqrt14_34),.doutb(asqrt[13]),.din(w_asqrt14_11[0]));
	jspl3 jspl3_w_asqrt15_0(.douta(w_asqrt15_0[0]),.doutb(w_asqrt15_0[1]),.doutc(w_asqrt15_0[2]),.din(asqrt_fa_15));
	jspl3 jspl3_w_asqrt15_1(.douta(w_asqrt15_1[0]),.doutb(w_asqrt15_1[1]),.doutc(w_asqrt15_1[2]),.din(w_asqrt15_0[0]));
	jspl3 jspl3_w_asqrt15_2(.douta(w_asqrt15_2[0]),.doutb(w_asqrt15_2[1]),.doutc(w_asqrt15_2[2]),.din(w_asqrt15_0[1]));
	jspl3 jspl3_w_asqrt15_3(.douta(w_asqrt15_3[0]),.doutb(w_asqrt15_3[1]),.doutc(w_asqrt15_3[2]),.din(w_asqrt15_0[2]));
	jspl3 jspl3_w_asqrt15_4(.douta(w_asqrt15_4[0]),.doutb(w_asqrt15_4[1]),.doutc(w_asqrt15_4[2]),.din(w_asqrt15_1[0]));
	jspl3 jspl3_w_asqrt15_5(.douta(w_asqrt15_5[0]),.doutb(w_asqrt15_5[1]),.doutc(w_asqrt15_5[2]),.din(w_asqrt15_1[1]));
	jspl3 jspl3_w_asqrt15_6(.douta(w_asqrt15_6[0]),.doutb(w_asqrt15_6[1]),.doutc(w_asqrt15_6[2]),.din(w_asqrt15_1[2]));
	jspl3 jspl3_w_asqrt15_7(.douta(w_asqrt15_7[0]),.doutb(w_asqrt15_7[1]),.doutc(w_asqrt15_7[2]),.din(w_asqrt15_2[0]));
	jspl3 jspl3_w_asqrt15_8(.douta(w_asqrt15_8[0]),.doutb(w_asqrt15_8[1]),.doutc(w_asqrt15_8[2]),.din(w_asqrt15_2[1]));
	jspl3 jspl3_w_asqrt15_9(.douta(w_asqrt15_9[0]),.doutb(w_asqrt15_9[1]),.doutc(w_asqrt15_9[2]),.din(w_asqrt15_2[2]));
	jspl3 jspl3_w_asqrt15_10(.douta(w_asqrt15_10[0]),.doutb(w_asqrt15_10[1]),.doutc(w_asqrt15_10[2]),.din(w_asqrt15_3[0]));
	jspl3 jspl3_w_asqrt15_11(.douta(w_asqrt15_11[0]),.doutb(w_asqrt15_11[1]),.doutc(w_asqrt15_11[2]),.din(w_asqrt15_3[1]));
	jspl jspl_w_asqrt15_12(.douta(w_asqrt15_12),.doutb(asqrt[14]),.din(w_asqrt15_3[2]));
	jspl3 jspl3_w_asqrt16_0(.douta(w_asqrt16_0[0]),.doutb(w_asqrt16_0[1]),.doutc(w_asqrt16_0[2]),.din(asqrt_fa_16));
	jspl3 jspl3_w_asqrt16_1(.douta(w_asqrt16_1[0]),.doutb(w_asqrt16_1[1]),.doutc(w_asqrt16_1[2]),.din(w_asqrt16_0[0]));
	jspl3 jspl3_w_asqrt16_2(.douta(w_asqrt16_2[0]),.doutb(w_asqrt16_2[1]),.doutc(w_asqrt16_2[2]),.din(w_asqrt16_0[1]));
	jspl3 jspl3_w_asqrt16_3(.douta(w_asqrt16_3[0]),.doutb(w_asqrt16_3[1]),.doutc(w_asqrt16_3[2]),.din(w_asqrt16_0[2]));
	jspl3 jspl3_w_asqrt16_4(.douta(w_asqrt16_4[0]),.doutb(w_asqrt16_4[1]),.doutc(w_asqrt16_4[2]),.din(w_asqrt16_1[0]));
	jspl3 jspl3_w_asqrt16_5(.douta(w_asqrt16_5[0]),.doutb(w_asqrt16_5[1]),.doutc(w_asqrt16_5[2]),.din(w_asqrt16_1[1]));
	jspl3 jspl3_w_asqrt16_6(.douta(w_asqrt16_6[0]),.doutb(w_asqrt16_6[1]),.doutc(w_asqrt16_6[2]),.din(w_asqrt16_1[2]));
	jspl3 jspl3_w_asqrt16_7(.douta(w_asqrt16_7[0]),.doutb(w_asqrt16_7[1]),.doutc(w_asqrt16_7[2]),.din(w_asqrt16_2[0]));
	jspl3 jspl3_w_asqrt16_8(.douta(w_asqrt16_8[0]),.doutb(w_asqrt16_8[1]),.doutc(w_asqrt16_8[2]),.din(w_asqrt16_2[1]));
	jspl3 jspl3_w_asqrt16_9(.douta(w_asqrt16_9[0]),.doutb(w_asqrt16_9[1]),.doutc(w_asqrt16_9[2]),.din(w_asqrt16_2[2]));
	jspl3 jspl3_w_asqrt16_10(.douta(w_asqrt16_10[0]),.doutb(w_asqrt16_10[1]),.doutc(w_asqrt16_10[2]),.din(w_asqrt16_3[0]));
	jspl3 jspl3_w_asqrt16_11(.douta(w_asqrt16_11[0]),.doutb(w_asqrt16_11[1]),.doutc(w_asqrt16_11[2]),.din(w_asqrt16_3[1]));
	jspl3 jspl3_w_asqrt16_12(.douta(w_asqrt16_12[0]),.doutb(w_asqrt16_12[1]),.doutc(w_asqrt16_12[2]),.din(w_asqrt16_3[2]));
	jspl3 jspl3_w_asqrt16_13(.douta(w_asqrt16_13[0]),.doutb(w_asqrt16_13[1]),.doutc(w_asqrt16_13[2]),.din(w_asqrt16_4[0]));
	jspl3 jspl3_w_asqrt16_14(.douta(w_asqrt16_14[0]),.doutb(w_asqrt16_14[1]),.doutc(w_asqrt16_14[2]),.din(w_asqrt16_4[1]));
	jspl3 jspl3_w_asqrt16_15(.douta(w_asqrt16_15[0]),.doutb(w_asqrt16_15[1]),.doutc(w_asqrt16_15[2]),.din(w_asqrt16_4[2]));
	jspl3 jspl3_w_asqrt16_16(.douta(w_asqrt16_16[0]),.doutb(w_asqrt16_16[1]),.doutc(w_asqrt16_16[2]),.din(w_asqrt16_5[0]));
	jspl3 jspl3_w_asqrt16_17(.douta(w_asqrt16_17[0]),.doutb(w_asqrt16_17[1]),.doutc(w_asqrt16_17[2]),.din(w_asqrt16_5[1]));
	jspl3 jspl3_w_asqrt16_18(.douta(w_asqrt16_18[0]),.doutb(w_asqrt16_18[1]),.doutc(w_asqrt16_18[2]),.din(w_asqrt16_5[2]));
	jspl3 jspl3_w_asqrt16_19(.douta(w_asqrt16_19[0]),.doutb(w_asqrt16_19[1]),.doutc(w_asqrt16_19[2]),.din(w_asqrt16_6[0]));
	jspl3 jspl3_w_asqrt16_20(.douta(w_asqrt16_20[0]),.doutb(w_asqrt16_20[1]),.doutc(w_asqrt16_20[2]),.din(w_asqrt16_6[1]));
	jspl3 jspl3_w_asqrt16_21(.douta(w_asqrt16_21[0]),.doutb(w_asqrt16_21[1]),.doutc(w_asqrt16_21[2]),.din(w_asqrt16_6[2]));
	jspl3 jspl3_w_asqrt16_22(.douta(w_asqrt16_22[0]),.doutb(w_asqrt16_22[1]),.doutc(w_asqrt16_22[2]),.din(w_asqrt16_7[0]));
	jspl3 jspl3_w_asqrt16_23(.douta(w_asqrt16_23[0]),.doutb(w_asqrt16_23[1]),.doutc(w_asqrt16_23[2]),.din(w_asqrt16_7[1]));
	jspl3 jspl3_w_asqrt16_24(.douta(w_asqrt16_24[0]),.doutb(w_asqrt16_24[1]),.doutc(w_asqrt16_24[2]),.din(w_asqrt16_7[2]));
	jspl3 jspl3_w_asqrt16_25(.douta(w_asqrt16_25[0]),.doutb(w_asqrt16_25[1]),.doutc(w_asqrt16_25[2]),.din(w_asqrt16_8[0]));
	jspl3 jspl3_w_asqrt16_26(.douta(w_asqrt16_26[0]),.doutb(w_asqrt16_26[1]),.doutc(w_asqrt16_26[2]),.din(w_asqrt16_8[1]));
	jspl3 jspl3_w_asqrt16_27(.douta(w_asqrt16_27[0]),.doutb(w_asqrt16_27[1]),.doutc(w_asqrt16_27[2]),.din(w_asqrt16_8[2]));
	jspl3 jspl3_w_asqrt16_28(.douta(w_asqrt16_28[0]),.doutb(w_asqrt16_28[1]),.doutc(w_asqrt16_28[2]),.din(w_asqrt16_9[0]));
	jspl3 jspl3_w_asqrt16_29(.douta(w_asqrt16_29[0]),.doutb(w_asqrt16_29[1]),.doutc(w_asqrt16_29[2]),.din(w_asqrt16_9[1]));
	jspl3 jspl3_w_asqrt16_30(.douta(w_asqrt16_30[0]),.doutb(w_asqrt16_30[1]),.doutc(w_asqrt16_30[2]),.din(w_asqrt16_9[2]));
	jspl3 jspl3_w_asqrt16_31(.douta(w_asqrt16_31[0]),.doutb(w_asqrt16_31[1]),.doutc(w_asqrt16_31[2]),.din(w_asqrt16_10[0]));
	jspl3 jspl3_w_asqrt16_32(.douta(w_asqrt16_32[0]),.doutb(w_asqrt16_32[1]),.doutc(w_asqrt16_32[2]),.din(w_asqrt16_10[1]));
	jspl3 jspl3_w_asqrt16_33(.douta(w_asqrt16_33[0]),.doutb(w_asqrt16_33[1]),.doutc(w_asqrt16_33[2]),.din(w_asqrt16_10[2]));
	jspl3 jspl3_w_asqrt16_34(.douta(w_asqrt16_34[0]),.doutb(w_asqrt16_34[1]),.doutc(asqrt[15]),.din(w_asqrt16_11[0]));
	jspl3 jspl3_w_asqrt17_0(.douta(w_asqrt17_0[0]),.doutb(w_asqrt17_0[1]),.doutc(w_asqrt17_0[2]),.din(asqrt_fa_17));
	jspl3 jspl3_w_asqrt17_1(.douta(w_asqrt17_1[0]),.doutb(w_asqrt17_1[1]),.doutc(w_asqrt17_1[2]),.din(w_asqrt17_0[0]));
	jspl3 jspl3_w_asqrt17_2(.douta(w_asqrt17_2[0]),.doutb(w_asqrt17_2[1]),.doutc(w_asqrt17_2[2]),.din(w_asqrt17_0[1]));
	jspl3 jspl3_w_asqrt17_3(.douta(w_asqrt17_3[0]),.doutb(w_asqrt17_3[1]),.doutc(w_asqrt17_3[2]),.din(w_asqrt17_0[2]));
	jspl3 jspl3_w_asqrt17_4(.douta(w_asqrt17_4[0]),.doutb(w_asqrt17_4[1]),.doutc(w_asqrt17_4[2]),.din(w_asqrt17_1[0]));
	jspl3 jspl3_w_asqrt17_5(.douta(w_asqrt17_5[0]),.doutb(w_asqrt17_5[1]),.doutc(w_asqrt17_5[2]),.din(w_asqrt17_1[1]));
	jspl3 jspl3_w_asqrt17_6(.douta(w_asqrt17_6[0]),.doutb(w_asqrt17_6[1]),.doutc(w_asqrt17_6[2]),.din(w_asqrt17_1[2]));
	jspl3 jspl3_w_asqrt17_7(.douta(w_asqrt17_7[0]),.doutb(w_asqrt17_7[1]),.doutc(w_asqrt17_7[2]),.din(w_asqrt17_2[0]));
	jspl3 jspl3_w_asqrt17_8(.douta(w_asqrt17_8[0]),.doutb(w_asqrt17_8[1]),.doutc(w_asqrt17_8[2]),.din(w_asqrt17_2[1]));
	jspl3 jspl3_w_asqrt17_9(.douta(w_asqrt17_9[0]),.doutb(w_asqrt17_9[1]),.doutc(w_asqrt17_9[2]),.din(w_asqrt17_2[2]));
	jspl3 jspl3_w_asqrt17_10(.douta(w_asqrt17_10[0]),.doutb(w_asqrt17_10[1]),.doutc(w_asqrt17_10[2]),.din(w_asqrt17_3[0]));
	jspl3 jspl3_w_asqrt17_11(.douta(w_asqrt17_11[0]),.doutb(w_asqrt17_11[1]),.doutc(w_asqrt17_11[2]),.din(w_asqrt17_3[1]));
	jspl3 jspl3_w_asqrt17_12(.douta(w_asqrt17_12[0]),.doutb(w_asqrt17_12[1]),.doutc(w_asqrt17_12[2]),.din(w_asqrt17_3[2]));
	jspl3 jspl3_w_asqrt17_13(.douta(w_asqrt17_13[0]),.doutb(w_asqrt17_13[1]),.doutc(asqrt[16]),.din(w_asqrt17_4[0]));
	jspl3 jspl3_w_asqrt18_0(.douta(w_asqrt18_0[0]),.doutb(w_asqrt18_0[1]),.doutc(w_asqrt18_0[2]),.din(asqrt_fa_18));
	jspl3 jspl3_w_asqrt18_1(.douta(w_asqrt18_1[0]),.doutb(w_asqrt18_1[1]),.doutc(w_asqrt18_1[2]),.din(w_asqrt18_0[0]));
	jspl3 jspl3_w_asqrt18_2(.douta(w_asqrt18_2[0]),.doutb(w_asqrt18_2[1]),.doutc(w_asqrt18_2[2]),.din(w_asqrt18_0[1]));
	jspl3 jspl3_w_asqrt18_3(.douta(w_asqrt18_3[0]),.doutb(w_asqrt18_3[1]),.doutc(w_asqrt18_3[2]),.din(w_asqrt18_0[2]));
	jspl3 jspl3_w_asqrt18_4(.douta(w_asqrt18_4[0]),.doutb(w_asqrt18_4[1]),.doutc(w_asqrt18_4[2]),.din(w_asqrt18_1[0]));
	jspl3 jspl3_w_asqrt18_5(.douta(w_asqrt18_5[0]),.doutb(w_asqrt18_5[1]),.doutc(w_asqrt18_5[2]),.din(w_asqrt18_1[1]));
	jspl3 jspl3_w_asqrt18_6(.douta(w_asqrt18_6[0]),.doutb(w_asqrt18_6[1]),.doutc(w_asqrt18_6[2]),.din(w_asqrt18_1[2]));
	jspl3 jspl3_w_asqrt18_7(.douta(w_asqrt18_7[0]),.doutb(w_asqrt18_7[1]),.doutc(w_asqrt18_7[2]),.din(w_asqrt18_2[0]));
	jspl3 jspl3_w_asqrt18_8(.douta(w_asqrt18_8[0]),.doutb(w_asqrt18_8[1]),.doutc(w_asqrt18_8[2]),.din(w_asqrt18_2[1]));
	jspl3 jspl3_w_asqrt18_9(.douta(w_asqrt18_9[0]),.doutb(w_asqrt18_9[1]),.doutc(w_asqrt18_9[2]),.din(w_asqrt18_2[2]));
	jspl3 jspl3_w_asqrt18_10(.douta(w_asqrt18_10[0]),.doutb(w_asqrt18_10[1]),.doutc(w_asqrt18_10[2]),.din(w_asqrt18_3[0]));
	jspl3 jspl3_w_asqrt18_11(.douta(w_asqrt18_11[0]),.doutb(w_asqrt18_11[1]),.doutc(w_asqrt18_11[2]),.din(w_asqrt18_3[1]));
	jspl3 jspl3_w_asqrt18_12(.douta(w_asqrt18_12[0]),.doutb(w_asqrt18_12[1]),.doutc(w_asqrt18_12[2]),.din(w_asqrt18_3[2]));
	jspl3 jspl3_w_asqrt18_13(.douta(w_asqrt18_13[0]),.doutb(w_asqrt18_13[1]),.doutc(w_asqrt18_13[2]),.din(w_asqrt18_4[0]));
	jspl3 jspl3_w_asqrt18_14(.douta(w_asqrt18_14[0]),.doutb(w_asqrt18_14[1]),.doutc(w_asqrt18_14[2]),.din(w_asqrt18_4[1]));
	jspl3 jspl3_w_asqrt18_15(.douta(w_asqrt18_15[0]),.doutb(w_asqrt18_15[1]),.doutc(w_asqrt18_15[2]),.din(w_asqrt18_4[2]));
	jspl3 jspl3_w_asqrt18_16(.douta(w_asqrt18_16[0]),.doutb(w_asqrt18_16[1]),.doutc(w_asqrt18_16[2]),.din(w_asqrt18_5[0]));
	jspl3 jspl3_w_asqrt18_17(.douta(w_asqrt18_17[0]),.doutb(w_asqrt18_17[1]),.doutc(w_asqrt18_17[2]),.din(w_asqrt18_5[1]));
	jspl3 jspl3_w_asqrt18_18(.douta(w_asqrt18_18[0]),.doutb(w_asqrt18_18[1]),.doutc(w_asqrt18_18[2]),.din(w_asqrt18_5[2]));
	jspl3 jspl3_w_asqrt18_19(.douta(w_asqrt18_19[0]),.doutb(w_asqrt18_19[1]),.doutc(w_asqrt18_19[2]),.din(w_asqrt18_6[0]));
	jspl3 jspl3_w_asqrt18_20(.douta(w_asqrt18_20[0]),.doutb(w_asqrt18_20[1]),.doutc(w_asqrt18_20[2]),.din(w_asqrt18_6[1]));
	jspl3 jspl3_w_asqrt18_21(.douta(w_asqrt18_21[0]),.doutb(w_asqrt18_21[1]),.doutc(w_asqrt18_21[2]),.din(w_asqrt18_6[2]));
	jspl3 jspl3_w_asqrt18_22(.douta(w_asqrt18_22[0]),.doutb(w_asqrt18_22[1]),.doutc(w_asqrt18_22[2]),.din(w_asqrt18_7[0]));
	jspl3 jspl3_w_asqrt18_23(.douta(w_asqrt18_23[0]),.doutb(w_asqrt18_23[1]),.doutc(w_asqrt18_23[2]),.din(w_asqrt18_7[1]));
	jspl3 jspl3_w_asqrt18_24(.douta(w_asqrt18_24[0]),.doutb(w_asqrt18_24[1]),.doutc(w_asqrt18_24[2]),.din(w_asqrt18_7[2]));
	jspl3 jspl3_w_asqrt18_25(.douta(w_asqrt18_25[0]),.doutb(w_asqrt18_25[1]),.doutc(w_asqrt18_25[2]),.din(w_asqrt18_8[0]));
	jspl3 jspl3_w_asqrt18_26(.douta(w_asqrt18_26[0]),.doutb(w_asqrt18_26[1]),.doutc(w_asqrt18_26[2]),.din(w_asqrt18_8[1]));
	jspl3 jspl3_w_asqrt18_27(.douta(w_asqrt18_27[0]),.doutb(w_asqrt18_27[1]),.doutc(w_asqrt18_27[2]),.din(w_asqrt18_8[2]));
	jspl3 jspl3_w_asqrt18_28(.douta(w_asqrt18_28[0]),.doutb(w_asqrt18_28[1]),.doutc(w_asqrt18_28[2]),.din(w_asqrt18_9[0]));
	jspl3 jspl3_w_asqrt18_29(.douta(w_asqrt18_29[0]),.doutb(w_asqrt18_29[1]),.doutc(w_asqrt18_29[2]),.din(w_asqrt18_9[1]));
	jspl3 jspl3_w_asqrt18_30(.douta(w_asqrt18_30[0]),.doutb(w_asqrt18_30[1]),.doutc(w_asqrt18_30[2]),.din(w_asqrt18_9[2]));
	jspl3 jspl3_w_asqrt18_31(.douta(w_asqrt18_31[0]),.doutb(w_asqrt18_31[1]),.doutc(w_asqrt18_31[2]),.din(w_asqrt18_10[0]));
	jspl3 jspl3_w_asqrt18_32(.douta(w_asqrt18_32[0]),.doutb(w_asqrt18_32[1]),.doutc(w_asqrt18_32[2]),.din(w_asqrt18_10[1]));
	jspl3 jspl3_w_asqrt18_33(.douta(w_asqrt18_33[0]),.doutb(w_asqrt18_33[1]),.doutc(w_asqrt18_33[2]),.din(w_asqrt18_10[2]));
	jspl3 jspl3_w_asqrt18_34(.douta(w_asqrt18_34[0]),.doutb(w_asqrt18_34[1]),.doutc(w_asqrt18_34[2]),.din(w_asqrt18_11[0]));
	jspl jspl_w_asqrt18_35(.douta(w_asqrt18_35),.doutb(asqrt[17]),.din(w_asqrt18_11[1]));
	jspl3 jspl3_w_asqrt19_0(.douta(w_asqrt19_0[0]),.doutb(w_asqrt19_0[1]),.doutc(w_asqrt19_0[2]),.din(asqrt_fa_19));
	jspl3 jspl3_w_asqrt19_1(.douta(w_asqrt19_1[0]),.doutb(w_asqrt19_1[1]),.doutc(w_asqrt19_1[2]),.din(w_asqrt19_0[0]));
	jspl3 jspl3_w_asqrt19_2(.douta(w_asqrt19_2[0]),.doutb(w_asqrt19_2[1]),.doutc(w_asqrt19_2[2]),.din(w_asqrt19_0[1]));
	jspl3 jspl3_w_asqrt19_3(.douta(w_asqrt19_3[0]),.doutb(w_asqrt19_3[1]),.doutc(w_asqrt19_3[2]),.din(w_asqrt19_0[2]));
	jspl3 jspl3_w_asqrt19_4(.douta(w_asqrt19_4[0]),.doutb(w_asqrt19_4[1]),.doutc(w_asqrt19_4[2]),.din(w_asqrt19_1[0]));
	jspl3 jspl3_w_asqrt19_5(.douta(w_asqrt19_5[0]),.doutb(w_asqrt19_5[1]),.doutc(w_asqrt19_5[2]),.din(w_asqrt19_1[1]));
	jspl3 jspl3_w_asqrt19_6(.douta(w_asqrt19_6[0]),.doutb(w_asqrt19_6[1]),.doutc(w_asqrt19_6[2]),.din(w_asqrt19_1[2]));
	jspl3 jspl3_w_asqrt19_7(.douta(w_asqrt19_7[0]),.doutb(w_asqrt19_7[1]),.doutc(w_asqrt19_7[2]),.din(w_asqrt19_2[0]));
	jspl3 jspl3_w_asqrt19_8(.douta(w_asqrt19_8[0]),.doutb(w_asqrt19_8[1]),.doutc(w_asqrt19_8[2]),.din(w_asqrt19_2[1]));
	jspl3 jspl3_w_asqrt19_9(.douta(w_asqrt19_9[0]),.doutb(w_asqrt19_9[1]),.doutc(w_asqrt19_9[2]),.din(w_asqrt19_2[2]));
	jspl3 jspl3_w_asqrt19_10(.douta(w_asqrt19_10[0]),.doutb(w_asqrt19_10[1]),.doutc(w_asqrt19_10[2]),.din(w_asqrt19_3[0]));
	jspl3 jspl3_w_asqrt19_11(.douta(w_asqrt19_11[0]),.doutb(w_asqrt19_11[1]),.doutc(w_asqrt19_11[2]),.din(w_asqrt19_3[1]));
	jspl3 jspl3_w_asqrt19_12(.douta(w_asqrt19_12[0]),.doutb(w_asqrt19_12[1]),.doutc(w_asqrt19_12[2]),.din(w_asqrt19_3[2]));
	jspl3 jspl3_w_asqrt19_13(.douta(w_asqrt19_13[0]),.doutb(w_asqrt19_13[1]),.doutc(w_asqrt19_13[2]),.din(w_asqrt19_4[0]));
	jspl jspl_w_asqrt19_14(.douta(w_asqrt19_14),.doutb(asqrt[18]),.din(w_asqrt19_4[1]));
	jspl3 jspl3_w_asqrt20_0(.douta(w_asqrt20_0[0]),.doutb(w_asqrt20_0[1]),.doutc(w_asqrt20_0[2]),.din(asqrt_fa_20));
	jspl3 jspl3_w_asqrt20_1(.douta(w_asqrt20_1[0]),.doutb(w_asqrt20_1[1]),.doutc(w_asqrt20_1[2]),.din(w_asqrt20_0[0]));
	jspl3 jspl3_w_asqrt20_2(.douta(w_asqrt20_2[0]),.doutb(w_asqrt20_2[1]),.doutc(w_asqrt20_2[2]),.din(w_asqrt20_0[1]));
	jspl3 jspl3_w_asqrt20_3(.douta(w_asqrt20_3[0]),.doutb(w_asqrt20_3[1]),.doutc(w_asqrt20_3[2]),.din(w_asqrt20_0[2]));
	jspl3 jspl3_w_asqrt20_4(.douta(w_asqrt20_4[0]),.doutb(w_asqrt20_4[1]),.doutc(w_asqrt20_4[2]),.din(w_asqrt20_1[0]));
	jspl3 jspl3_w_asqrt20_5(.douta(w_asqrt20_5[0]),.doutb(w_asqrt20_5[1]),.doutc(w_asqrt20_5[2]),.din(w_asqrt20_1[1]));
	jspl3 jspl3_w_asqrt20_6(.douta(w_asqrt20_6[0]),.doutb(w_asqrt20_6[1]),.doutc(w_asqrt20_6[2]),.din(w_asqrt20_1[2]));
	jspl3 jspl3_w_asqrt20_7(.douta(w_asqrt20_7[0]),.doutb(w_asqrt20_7[1]),.doutc(w_asqrt20_7[2]),.din(w_asqrt20_2[0]));
	jspl3 jspl3_w_asqrt20_8(.douta(w_asqrt20_8[0]),.doutb(w_asqrt20_8[1]),.doutc(w_asqrt20_8[2]),.din(w_asqrt20_2[1]));
	jspl3 jspl3_w_asqrt20_9(.douta(w_asqrt20_9[0]),.doutb(w_asqrt20_9[1]),.doutc(w_asqrt20_9[2]),.din(w_asqrt20_2[2]));
	jspl3 jspl3_w_asqrt20_10(.douta(w_asqrt20_10[0]),.doutb(w_asqrt20_10[1]),.doutc(w_asqrt20_10[2]),.din(w_asqrt20_3[0]));
	jspl3 jspl3_w_asqrt20_11(.douta(w_asqrt20_11[0]),.doutb(w_asqrt20_11[1]),.doutc(w_asqrt20_11[2]),.din(w_asqrt20_3[1]));
	jspl3 jspl3_w_asqrt20_12(.douta(w_asqrt20_12[0]),.doutb(w_asqrt20_12[1]),.doutc(w_asqrt20_12[2]),.din(w_asqrt20_3[2]));
	jspl3 jspl3_w_asqrt20_13(.douta(w_asqrt20_13[0]),.doutb(w_asqrt20_13[1]),.doutc(w_asqrt20_13[2]),.din(w_asqrt20_4[0]));
	jspl3 jspl3_w_asqrt20_14(.douta(w_asqrt20_14[0]),.doutb(w_asqrt20_14[1]),.doutc(w_asqrt20_14[2]),.din(w_asqrt20_4[1]));
	jspl3 jspl3_w_asqrt20_15(.douta(w_asqrt20_15[0]),.doutb(w_asqrt20_15[1]),.doutc(w_asqrt20_15[2]),.din(w_asqrt20_4[2]));
	jspl3 jspl3_w_asqrt20_16(.douta(w_asqrt20_16[0]),.doutb(w_asqrt20_16[1]),.doutc(w_asqrt20_16[2]),.din(w_asqrt20_5[0]));
	jspl3 jspl3_w_asqrt20_17(.douta(w_asqrt20_17[0]),.doutb(w_asqrt20_17[1]),.doutc(w_asqrt20_17[2]),.din(w_asqrt20_5[1]));
	jspl3 jspl3_w_asqrt20_18(.douta(w_asqrt20_18[0]),.doutb(w_asqrt20_18[1]),.doutc(w_asqrt20_18[2]),.din(w_asqrt20_5[2]));
	jspl3 jspl3_w_asqrt20_19(.douta(w_asqrt20_19[0]),.doutb(w_asqrt20_19[1]),.doutc(w_asqrt20_19[2]),.din(w_asqrt20_6[0]));
	jspl3 jspl3_w_asqrt20_20(.douta(w_asqrt20_20[0]),.doutb(w_asqrt20_20[1]),.doutc(w_asqrt20_20[2]),.din(w_asqrt20_6[1]));
	jspl3 jspl3_w_asqrt20_21(.douta(w_asqrt20_21[0]),.doutb(w_asqrt20_21[1]),.doutc(w_asqrt20_21[2]),.din(w_asqrt20_6[2]));
	jspl3 jspl3_w_asqrt20_22(.douta(w_asqrt20_22[0]),.doutb(w_asqrt20_22[1]),.doutc(w_asqrt20_22[2]),.din(w_asqrt20_7[0]));
	jspl3 jspl3_w_asqrt20_23(.douta(w_asqrt20_23[0]),.doutb(w_asqrt20_23[1]),.doutc(w_asqrt20_23[2]),.din(w_asqrt20_7[1]));
	jspl3 jspl3_w_asqrt20_24(.douta(w_asqrt20_24[0]),.doutb(w_asqrt20_24[1]),.doutc(w_asqrt20_24[2]),.din(w_asqrt20_7[2]));
	jspl3 jspl3_w_asqrt20_25(.douta(w_asqrt20_25[0]),.doutb(w_asqrt20_25[1]),.doutc(w_asqrt20_25[2]),.din(w_asqrt20_8[0]));
	jspl3 jspl3_w_asqrt20_26(.douta(w_asqrt20_26[0]),.doutb(w_asqrt20_26[1]),.doutc(w_asqrt20_26[2]),.din(w_asqrt20_8[1]));
	jspl3 jspl3_w_asqrt20_27(.douta(w_asqrt20_27[0]),.doutb(w_asqrt20_27[1]),.doutc(w_asqrt20_27[2]),.din(w_asqrt20_8[2]));
	jspl3 jspl3_w_asqrt20_28(.douta(w_asqrt20_28[0]),.doutb(w_asqrt20_28[1]),.doutc(w_asqrt20_28[2]),.din(w_asqrt20_9[0]));
	jspl3 jspl3_w_asqrt20_29(.douta(w_asqrt20_29[0]),.doutb(w_asqrt20_29[1]),.doutc(w_asqrt20_29[2]),.din(w_asqrt20_9[1]));
	jspl3 jspl3_w_asqrt20_30(.douta(w_asqrt20_30[0]),.doutb(w_asqrt20_30[1]),.doutc(w_asqrt20_30[2]),.din(w_asqrt20_9[2]));
	jspl3 jspl3_w_asqrt20_31(.douta(w_asqrt20_31[0]),.doutb(w_asqrt20_31[1]),.doutc(w_asqrt20_31[2]),.din(w_asqrt20_10[0]));
	jspl3 jspl3_w_asqrt20_32(.douta(w_asqrt20_32[0]),.doutb(w_asqrt20_32[1]),.doutc(w_asqrt20_32[2]),.din(w_asqrt20_10[1]));
	jspl3 jspl3_w_asqrt20_33(.douta(w_asqrt20_33[0]),.doutb(w_asqrt20_33[1]),.doutc(w_asqrt20_33[2]),.din(w_asqrt20_10[2]));
	jspl3 jspl3_w_asqrt20_34(.douta(w_asqrt20_34[0]),.doutb(w_asqrt20_34[1]),.doutc(w_asqrt20_34[2]),.din(w_asqrt20_11[0]));
	jspl jspl_w_asqrt20_35(.douta(w_asqrt20_35),.doutb(asqrt[19]),.din(w_asqrt20_11[1]));
	jspl3 jspl3_w_asqrt21_0(.douta(w_asqrt21_0[0]),.doutb(w_asqrt21_0[1]),.doutc(w_asqrt21_0[2]),.din(asqrt_fa_21));
	jspl3 jspl3_w_asqrt21_1(.douta(w_asqrt21_1[0]),.doutb(w_asqrt21_1[1]),.doutc(w_asqrt21_1[2]),.din(w_asqrt21_0[0]));
	jspl3 jspl3_w_asqrt21_2(.douta(w_asqrt21_2[0]),.doutb(w_asqrt21_2[1]),.doutc(w_asqrt21_2[2]),.din(w_asqrt21_0[1]));
	jspl3 jspl3_w_asqrt21_3(.douta(w_asqrt21_3[0]),.doutb(w_asqrt21_3[1]),.doutc(w_asqrt21_3[2]),.din(w_asqrt21_0[2]));
	jspl3 jspl3_w_asqrt21_4(.douta(w_asqrt21_4[0]),.doutb(w_asqrt21_4[1]),.doutc(w_asqrt21_4[2]),.din(w_asqrt21_1[0]));
	jspl3 jspl3_w_asqrt21_5(.douta(w_asqrt21_5[0]),.doutb(w_asqrt21_5[1]),.doutc(w_asqrt21_5[2]),.din(w_asqrt21_1[1]));
	jspl3 jspl3_w_asqrt21_6(.douta(w_asqrt21_6[0]),.doutb(w_asqrt21_6[1]),.doutc(w_asqrt21_6[2]),.din(w_asqrt21_1[2]));
	jspl3 jspl3_w_asqrt21_7(.douta(w_asqrt21_7[0]),.doutb(w_asqrt21_7[1]),.doutc(w_asqrt21_7[2]),.din(w_asqrt21_2[0]));
	jspl3 jspl3_w_asqrt21_8(.douta(w_asqrt21_8[0]),.doutb(w_asqrt21_8[1]),.doutc(w_asqrt21_8[2]),.din(w_asqrt21_2[1]));
	jspl3 jspl3_w_asqrt21_9(.douta(w_asqrt21_9[0]),.doutb(w_asqrt21_9[1]),.doutc(w_asqrt21_9[2]),.din(w_asqrt21_2[2]));
	jspl3 jspl3_w_asqrt21_10(.douta(w_asqrt21_10[0]),.doutb(w_asqrt21_10[1]),.doutc(w_asqrt21_10[2]),.din(w_asqrt21_3[0]));
	jspl3 jspl3_w_asqrt21_11(.douta(w_asqrt21_11[0]),.doutb(w_asqrt21_11[1]),.doutc(w_asqrt21_11[2]),.din(w_asqrt21_3[1]));
	jspl3 jspl3_w_asqrt21_12(.douta(w_asqrt21_12[0]),.doutb(w_asqrt21_12[1]),.doutc(w_asqrt21_12[2]),.din(w_asqrt21_3[2]));
	jspl3 jspl3_w_asqrt21_13(.douta(w_asqrt21_13[0]),.doutb(w_asqrt21_13[1]),.doutc(w_asqrt21_13[2]),.din(w_asqrt21_4[0]));
	jspl3 jspl3_w_asqrt21_14(.douta(w_asqrt21_14[0]),.doutb(w_asqrt21_14[1]),.doutc(w_asqrt21_14[2]),.din(w_asqrt21_4[1]));
	jspl3 jspl3_w_asqrt21_15(.douta(w_asqrt21_15[0]),.doutb(w_asqrt21_15[1]),.doutc(w_asqrt21_15[2]),.din(w_asqrt21_4[2]));
	jspl jspl_w_asqrt21_16(.douta(w_asqrt21_16),.doutb(asqrt[20]),.din(w_asqrt21_5[0]));
	jspl3 jspl3_w_asqrt22_0(.douta(w_asqrt22_0[0]),.doutb(w_asqrt22_0[1]),.doutc(w_asqrt22_0[2]),.din(asqrt_fa_22));
	jspl3 jspl3_w_asqrt22_1(.douta(w_asqrt22_1[0]),.doutb(w_asqrt22_1[1]),.doutc(w_asqrt22_1[2]),.din(w_asqrt22_0[0]));
	jspl3 jspl3_w_asqrt22_2(.douta(w_asqrt22_2[0]),.doutb(w_asqrt22_2[1]),.doutc(w_asqrt22_2[2]),.din(w_asqrt22_0[1]));
	jspl3 jspl3_w_asqrt22_3(.douta(w_asqrt22_3[0]),.doutb(w_asqrt22_3[1]),.doutc(w_asqrt22_3[2]),.din(w_asqrt22_0[2]));
	jspl3 jspl3_w_asqrt22_4(.douta(w_asqrt22_4[0]),.doutb(w_asqrt22_4[1]),.doutc(w_asqrt22_4[2]),.din(w_asqrt22_1[0]));
	jspl3 jspl3_w_asqrt22_5(.douta(w_asqrt22_5[0]),.doutb(w_asqrt22_5[1]),.doutc(w_asqrt22_5[2]),.din(w_asqrt22_1[1]));
	jspl3 jspl3_w_asqrt22_6(.douta(w_asqrt22_6[0]),.doutb(w_asqrt22_6[1]),.doutc(w_asqrt22_6[2]),.din(w_asqrt22_1[2]));
	jspl3 jspl3_w_asqrt22_7(.douta(w_asqrt22_7[0]),.doutb(w_asqrt22_7[1]),.doutc(w_asqrt22_7[2]),.din(w_asqrt22_2[0]));
	jspl3 jspl3_w_asqrt22_8(.douta(w_asqrt22_8[0]),.doutb(w_asqrt22_8[1]),.doutc(w_asqrt22_8[2]),.din(w_asqrt22_2[1]));
	jspl3 jspl3_w_asqrt22_9(.douta(w_asqrt22_9[0]),.doutb(w_asqrt22_9[1]),.doutc(w_asqrt22_9[2]),.din(w_asqrt22_2[2]));
	jspl3 jspl3_w_asqrt22_10(.douta(w_asqrt22_10[0]),.doutb(w_asqrt22_10[1]),.doutc(w_asqrt22_10[2]),.din(w_asqrt22_3[0]));
	jspl3 jspl3_w_asqrt22_11(.douta(w_asqrt22_11[0]),.doutb(w_asqrt22_11[1]),.doutc(w_asqrt22_11[2]),.din(w_asqrt22_3[1]));
	jspl3 jspl3_w_asqrt22_12(.douta(w_asqrt22_12[0]),.doutb(w_asqrt22_12[1]),.doutc(w_asqrt22_12[2]),.din(w_asqrt22_3[2]));
	jspl3 jspl3_w_asqrt22_13(.douta(w_asqrt22_13[0]),.doutb(w_asqrt22_13[1]),.doutc(w_asqrt22_13[2]),.din(w_asqrt22_4[0]));
	jspl3 jspl3_w_asqrt22_14(.douta(w_asqrt22_14[0]),.doutb(w_asqrt22_14[1]),.doutc(w_asqrt22_14[2]),.din(w_asqrt22_4[1]));
	jspl3 jspl3_w_asqrt22_15(.douta(w_asqrt22_15[0]),.doutb(w_asqrt22_15[1]),.doutc(w_asqrt22_15[2]),.din(w_asqrt22_4[2]));
	jspl3 jspl3_w_asqrt22_16(.douta(w_asqrt22_16[0]),.doutb(w_asqrt22_16[1]),.doutc(w_asqrt22_16[2]),.din(w_asqrt22_5[0]));
	jspl3 jspl3_w_asqrt22_17(.douta(w_asqrt22_17[0]),.doutb(w_asqrt22_17[1]),.doutc(w_asqrt22_17[2]),.din(w_asqrt22_5[1]));
	jspl3 jspl3_w_asqrt22_18(.douta(w_asqrt22_18[0]),.doutb(w_asqrt22_18[1]),.doutc(w_asqrt22_18[2]),.din(w_asqrt22_5[2]));
	jspl3 jspl3_w_asqrt22_19(.douta(w_asqrt22_19[0]),.doutb(w_asqrt22_19[1]),.doutc(w_asqrt22_19[2]),.din(w_asqrt22_6[0]));
	jspl3 jspl3_w_asqrt22_20(.douta(w_asqrt22_20[0]),.doutb(w_asqrt22_20[1]),.doutc(w_asqrt22_20[2]),.din(w_asqrt22_6[1]));
	jspl3 jspl3_w_asqrt22_21(.douta(w_asqrt22_21[0]),.doutb(w_asqrt22_21[1]),.doutc(w_asqrt22_21[2]),.din(w_asqrt22_6[2]));
	jspl3 jspl3_w_asqrt22_22(.douta(w_asqrt22_22[0]),.doutb(w_asqrt22_22[1]),.doutc(w_asqrt22_22[2]),.din(w_asqrt22_7[0]));
	jspl3 jspl3_w_asqrt22_23(.douta(w_asqrt22_23[0]),.doutb(w_asqrt22_23[1]),.doutc(w_asqrt22_23[2]),.din(w_asqrt22_7[1]));
	jspl3 jspl3_w_asqrt22_24(.douta(w_asqrt22_24[0]),.doutb(w_asqrt22_24[1]),.doutc(w_asqrt22_24[2]),.din(w_asqrt22_7[2]));
	jspl3 jspl3_w_asqrt22_25(.douta(w_asqrt22_25[0]),.doutb(w_asqrt22_25[1]),.doutc(w_asqrt22_25[2]),.din(w_asqrt22_8[0]));
	jspl3 jspl3_w_asqrt22_26(.douta(w_asqrt22_26[0]),.doutb(w_asqrt22_26[1]),.doutc(w_asqrt22_26[2]),.din(w_asqrt22_8[1]));
	jspl3 jspl3_w_asqrt22_27(.douta(w_asqrt22_27[0]),.doutb(w_asqrt22_27[1]),.doutc(w_asqrt22_27[2]),.din(w_asqrt22_8[2]));
	jspl3 jspl3_w_asqrt22_28(.douta(w_asqrt22_28[0]),.doutb(w_asqrt22_28[1]),.doutc(w_asqrt22_28[2]),.din(w_asqrt22_9[0]));
	jspl3 jspl3_w_asqrt22_29(.douta(w_asqrt22_29[0]),.doutb(w_asqrt22_29[1]),.doutc(w_asqrt22_29[2]),.din(w_asqrt22_9[1]));
	jspl3 jspl3_w_asqrt22_30(.douta(w_asqrt22_30[0]),.doutb(w_asqrt22_30[1]),.doutc(w_asqrt22_30[2]),.din(w_asqrt22_9[2]));
	jspl3 jspl3_w_asqrt22_31(.douta(w_asqrt22_31[0]),.doutb(w_asqrt22_31[1]),.doutc(w_asqrt22_31[2]),.din(w_asqrt22_10[0]));
	jspl3 jspl3_w_asqrt22_32(.douta(w_asqrt22_32[0]),.doutb(w_asqrt22_32[1]),.doutc(w_asqrt22_32[2]),.din(w_asqrt22_10[1]));
	jspl3 jspl3_w_asqrt22_33(.douta(w_asqrt22_33[0]),.doutb(w_asqrt22_33[1]),.doutc(w_asqrt22_33[2]),.din(w_asqrt22_10[2]));
	jspl3 jspl3_w_asqrt22_34(.douta(w_asqrt22_34[0]),.doutb(w_asqrt22_34[1]),.doutc(w_asqrt22_34[2]),.din(w_asqrt22_11[0]));
	jspl3 jspl3_w_asqrt22_35(.douta(w_asqrt22_35[0]),.doutb(w_asqrt22_35[1]),.doutc(w_asqrt22_35[2]),.din(w_asqrt22_11[1]));
	jspl jspl_w_asqrt22_36(.douta(w_asqrt22_36),.doutb(asqrt[21]),.din(w_asqrt22_11[2]));
	jspl3 jspl3_w_asqrt23_0(.douta(w_asqrt23_0[0]),.doutb(w_asqrt23_0[1]),.doutc(w_asqrt23_0[2]),.din(asqrt_fa_23));
	jspl3 jspl3_w_asqrt23_1(.douta(w_asqrt23_1[0]),.doutb(w_asqrt23_1[1]),.doutc(w_asqrt23_1[2]),.din(w_asqrt23_0[0]));
	jspl3 jspl3_w_asqrt23_2(.douta(w_asqrt23_2[0]),.doutb(w_asqrt23_2[1]),.doutc(w_asqrt23_2[2]),.din(w_asqrt23_0[1]));
	jspl3 jspl3_w_asqrt23_3(.douta(w_asqrt23_3[0]),.doutb(w_asqrt23_3[1]),.doutc(w_asqrt23_3[2]),.din(w_asqrt23_0[2]));
	jspl3 jspl3_w_asqrt23_4(.douta(w_asqrt23_4[0]),.doutb(w_asqrt23_4[1]),.doutc(w_asqrt23_4[2]),.din(w_asqrt23_1[0]));
	jspl3 jspl3_w_asqrt23_5(.douta(w_asqrt23_5[0]),.doutb(w_asqrt23_5[1]),.doutc(w_asqrt23_5[2]),.din(w_asqrt23_1[1]));
	jspl3 jspl3_w_asqrt23_6(.douta(w_asqrt23_6[0]),.doutb(w_asqrt23_6[1]),.doutc(w_asqrt23_6[2]),.din(w_asqrt23_1[2]));
	jspl3 jspl3_w_asqrt23_7(.douta(w_asqrt23_7[0]),.doutb(w_asqrt23_7[1]),.doutc(w_asqrt23_7[2]),.din(w_asqrt23_2[0]));
	jspl3 jspl3_w_asqrt23_8(.douta(w_asqrt23_8[0]),.doutb(w_asqrt23_8[1]),.doutc(w_asqrt23_8[2]),.din(w_asqrt23_2[1]));
	jspl3 jspl3_w_asqrt23_9(.douta(w_asqrt23_9[0]),.doutb(w_asqrt23_9[1]),.doutc(w_asqrt23_9[2]),.din(w_asqrt23_2[2]));
	jspl3 jspl3_w_asqrt23_10(.douta(w_asqrt23_10[0]),.doutb(w_asqrt23_10[1]),.doutc(w_asqrt23_10[2]),.din(w_asqrt23_3[0]));
	jspl3 jspl3_w_asqrt23_11(.douta(w_asqrt23_11[0]),.doutb(w_asqrt23_11[1]),.doutc(w_asqrt23_11[2]),.din(w_asqrt23_3[1]));
	jspl3 jspl3_w_asqrt23_12(.douta(w_asqrt23_12[0]),.doutb(w_asqrt23_12[1]),.doutc(w_asqrt23_12[2]),.din(w_asqrt23_3[2]));
	jspl3 jspl3_w_asqrt23_13(.douta(w_asqrt23_13[0]),.doutb(w_asqrt23_13[1]),.doutc(w_asqrt23_13[2]),.din(w_asqrt23_4[0]));
	jspl3 jspl3_w_asqrt23_14(.douta(w_asqrt23_14[0]),.doutb(w_asqrt23_14[1]),.doutc(w_asqrt23_14[2]),.din(w_asqrt23_4[1]));
	jspl3 jspl3_w_asqrt23_15(.douta(w_asqrt23_15[0]),.doutb(w_asqrt23_15[1]),.doutc(w_asqrt23_15[2]),.din(w_asqrt23_4[2]));
	jspl3 jspl3_w_asqrt23_16(.douta(w_asqrt23_16[0]),.doutb(w_asqrt23_16[1]),.doutc(w_asqrt23_16[2]),.din(w_asqrt23_5[0]));
	jspl3 jspl3_w_asqrt23_17(.douta(w_asqrt23_17[0]),.doutb(w_asqrt23_17[1]),.doutc(w_asqrt23_17[2]),.din(w_asqrt23_5[1]));
	jspl jspl_w_asqrt23_18(.douta(w_asqrt23_18),.doutb(asqrt[22]),.din(w_asqrt23_5[2]));
	jspl3 jspl3_w_asqrt24_0(.douta(w_asqrt24_0[0]),.doutb(w_asqrt24_0[1]),.doutc(w_asqrt24_0[2]),.din(asqrt_fa_24));
	jspl3 jspl3_w_asqrt24_1(.douta(w_asqrt24_1[0]),.doutb(w_asqrt24_1[1]),.doutc(w_asqrt24_1[2]),.din(w_asqrt24_0[0]));
	jspl3 jspl3_w_asqrt24_2(.douta(w_asqrt24_2[0]),.doutb(w_asqrt24_2[1]),.doutc(w_asqrt24_2[2]),.din(w_asqrt24_0[1]));
	jspl3 jspl3_w_asqrt24_3(.douta(w_asqrt24_3[0]),.doutb(w_asqrt24_3[1]),.doutc(w_asqrt24_3[2]),.din(w_asqrt24_0[2]));
	jspl3 jspl3_w_asqrt24_4(.douta(w_asqrt24_4[0]),.doutb(w_asqrt24_4[1]),.doutc(w_asqrt24_4[2]),.din(w_asqrt24_1[0]));
	jspl3 jspl3_w_asqrt24_5(.douta(w_asqrt24_5[0]),.doutb(w_asqrt24_5[1]),.doutc(w_asqrt24_5[2]),.din(w_asqrt24_1[1]));
	jspl3 jspl3_w_asqrt24_6(.douta(w_asqrt24_6[0]),.doutb(w_asqrt24_6[1]),.doutc(w_asqrt24_6[2]),.din(w_asqrt24_1[2]));
	jspl3 jspl3_w_asqrt24_7(.douta(w_asqrt24_7[0]),.doutb(w_asqrt24_7[1]),.doutc(w_asqrt24_7[2]),.din(w_asqrt24_2[0]));
	jspl3 jspl3_w_asqrt24_8(.douta(w_asqrt24_8[0]),.doutb(w_asqrt24_8[1]),.doutc(w_asqrt24_8[2]),.din(w_asqrt24_2[1]));
	jspl3 jspl3_w_asqrt24_9(.douta(w_asqrt24_9[0]),.doutb(w_asqrt24_9[1]),.doutc(w_asqrt24_9[2]),.din(w_asqrt24_2[2]));
	jspl3 jspl3_w_asqrt24_10(.douta(w_asqrt24_10[0]),.doutb(w_asqrt24_10[1]),.doutc(w_asqrt24_10[2]),.din(w_asqrt24_3[0]));
	jspl3 jspl3_w_asqrt24_11(.douta(w_asqrt24_11[0]),.doutb(w_asqrt24_11[1]),.doutc(w_asqrt24_11[2]),.din(w_asqrt24_3[1]));
	jspl3 jspl3_w_asqrt24_12(.douta(w_asqrt24_12[0]),.doutb(w_asqrt24_12[1]),.doutc(w_asqrt24_12[2]),.din(w_asqrt24_3[2]));
	jspl3 jspl3_w_asqrt24_13(.douta(w_asqrt24_13[0]),.doutb(w_asqrt24_13[1]),.doutc(w_asqrt24_13[2]),.din(w_asqrt24_4[0]));
	jspl3 jspl3_w_asqrt24_14(.douta(w_asqrt24_14[0]),.doutb(w_asqrt24_14[1]),.doutc(w_asqrt24_14[2]),.din(w_asqrt24_4[1]));
	jspl3 jspl3_w_asqrt24_15(.douta(w_asqrt24_15[0]),.doutb(w_asqrt24_15[1]),.doutc(w_asqrt24_15[2]),.din(w_asqrt24_4[2]));
	jspl3 jspl3_w_asqrt24_16(.douta(w_asqrt24_16[0]),.doutb(w_asqrt24_16[1]),.doutc(w_asqrt24_16[2]),.din(w_asqrt24_5[0]));
	jspl3 jspl3_w_asqrt24_17(.douta(w_asqrt24_17[0]),.doutb(w_asqrt24_17[1]),.doutc(w_asqrt24_17[2]),.din(w_asqrt24_5[1]));
	jspl3 jspl3_w_asqrt24_18(.douta(w_asqrt24_18[0]),.doutb(w_asqrt24_18[1]),.doutc(w_asqrt24_18[2]),.din(w_asqrt24_5[2]));
	jspl3 jspl3_w_asqrt24_19(.douta(w_asqrt24_19[0]),.doutb(w_asqrt24_19[1]),.doutc(w_asqrt24_19[2]),.din(w_asqrt24_6[0]));
	jspl3 jspl3_w_asqrt24_20(.douta(w_asqrt24_20[0]),.doutb(w_asqrt24_20[1]),.doutc(w_asqrt24_20[2]),.din(w_asqrt24_6[1]));
	jspl3 jspl3_w_asqrt24_21(.douta(w_asqrt24_21[0]),.doutb(w_asqrt24_21[1]),.doutc(w_asqrt24_21[2]),.din(w_asqrt24_6[2]));
	jspl3 jspl3_w_asqrt24_22(.douta(w_asqrt24_22[0]),.doutb(w_asqrt24_22[1]),.doutc(w_asqrt24_22[2]),.din(w_asqrt24_7[0]));
	jspl3 jspl3_w_asqrt24_23(.douta(w_asqrt24_23[0]),.doutb(w_asqrt24_23[1]),.doutc(w_asqrt24_23[2]),.din(w_asqrt24_7[1]));
	jspl3 jspl3_w_asqrt24_24(.douta(w_asqrt24_24[0]),.doutb(w_asqrt24_24[1]),.doutc(w_asqrt24_24[2]),.din(w_asqrt24_7[2]));
	jspl3 jspl3_w_asqrt24_25(.douta(w_asqrt24_25[0]),.doutb(w_asqrt24_25[1]),.doutc(w_asqrt24_25[2]),.din(w_asqrt24_8[0]));
	jspl3 jspl3_w_asqrt24_26(.douta(w_asqrt24_26[0]),.doutb(w_asqrt24_26[1]),.doutc(w_asqrt24_26[2]),.din(w_asqrt24_8[1]));
	jspl3 jspl3_w_asqrt24_27(.douta(w_asqrt24_27[0]),.doutb(w_asqrt24_27[1]),.doutc(w_asqrt24_27[2]),.din(w_asqrt24_8[2]));
	jspl3 jspl3_w_asqrt24_28(.douta(w_asqrt24_28[0]),.doutb(w_asqrt24_28[1]),.doutc(w_asqrt24_28[2]),.din(w_asqrt24_9[0]));
	jspl3 jspl3_w_asqrt24_29(.douta(w_asqrt24_29[0]),.doutb(w_asqrt24_29[1]),.doutc(w_asqrt24_29[2]),.din(w_asqrt24_9[1]));
	jspl3 jspl3_w_asqrt24_30(.douta(w_asqrt24_30[0]),.doutb(w_asqrt24_30[1]),.doutc(w_asqrt24_30[2]),.din(w_asqrt24_9[2]));
	jspl3 jspl3_w_asqrt24_31(.douta(w_asqrt24_31[0]),.doutb(w_asqrt24_31[1]),.doutc(w_asqrt24_31[2]),.din(w_asqrt24_10[0]));
	jspl3 jspl3_w_asqrt24_32(.douta(w_asqrt24_32[0]),.doutb(w_asqrt24_32[1]),.doutc(w_asqrt24_32[2]),.din(w_asqrt24_10[1]));
	jspl3 jspl3_w_asqrt24_33(.douta(w_asqrt24_33[0]),.doutb(w_asqrt24_33[1]),.doutc(w_asqrt24_33[2]),.din(w_asqrt24_10[2]));
	jspl3 jspl3_w_asqrt24_34(.douta(w_asqrt24_34[0]),.doutb(w_asqrt24_34[1]),.doutc(w_asqrt24_34[2]),.din(w_asqrt24_11[0]));
	jspl3 jspl3_w_asqrt24_35(.douta(w_asqrt24_35[0]),.doutb(w_asqrt24_35[1]),.doutc(w_asqrt24_35[2]),.din(w_asqrt24_11[1]));
	jspl3 jspl3_w_asqrt24_36(.douta(w_asqrt24_36[0]),.doutb(w_asqrt24_36[1]),.doutc(asqrt[23]),.din(w_asqrt24_11[2]));
	jspl3 jspl3_w_asqrt25_0(.douta(w_asqrt25_0[0]),.doutb(w_asqrt25_0[1]),.doutc(w_asqrt25_0[2]),.din(asqrt_fa_25));
	jspl3 jspl3_w_asqrt25_1(.douta(w_asqrt25_1[0]),.doutb(w_asqrt25_1[1]),.doutc(w_asqrt25_1[2]),.din(w_asqrt25_0[0]));
	jspl3 jspl3_w_asqrt25_2(.douta(w_asqrt25_2[0]),.doutb(w_asqrt25_2[1]),.doutc(w_asqrt25_2[2]),.din(w_asqrt25_0[1]));
	jspl3 jspl3_w_asqrt25_3(.douta(w_asqrt25_3[0]),.doutb(w_asqrt25_3[1]),.doutc(w_asqrt25_3[2]),.din(w_asqrt25_0[2]));
	jspl3 jspl3_w_asqrt25_4(.douta(w_asqrt25_4[0]),.doutb(w_asqrt25_4[1]),.doutc(w_asqrt25_4[2]),.din(w_asqrt25_1[0]));
	jspl3 jspl3_w_asqrt25_5(.douta(w_asqrt25_5[0]),.doutb(w_asqrt25_5[1]),.doutc(w_asqrt25_5[2]),.din(w_asqrt25_1[1]));
	jspl3 jspl3_w_asqrt25_6(.douta(w_asqrt25_6[0]),.doutb(w_asqrt25_6[1]),.doutc(w_asqrt25_6[2]),.din(w_asqrt25_1[2]));
	jspl3 jspl3_w_asqrt25_7(.douta(w_asqrt25_7[0]),.doutb(w_asqrt25_7[1]),.doutc(w_asqrt25_7[2]),.din(w_asqrt25_2[0]));
	jspl3 jspl3_w_asqrt25_8(.douta(w_asqrt25_8[0]),.doutb(w_asqrt25_8[1]),.doutc(w_asqrt25_8[2]),.din(w_asqrt25_2[1]));
	jspl3 jspl3_w_asqrt25_9(.douta(w_asqrt25_9[0]),.doutb(w_asqrt25_9[1]),.doutc(w_asqrt25_9[2]),.din(w_asqrt25_2[2]));
	jspl3 jspl3_w_asqrt25_10(.douta(w_asqrt25_10[0]),.doutb(w_asqrt25_10[1]),.doutc(w_asqrt25_10[2]),.din(w_asqrt25_3[0]));
	jspl3 jspl3_w_asqrt25_11(.douta(w_asqrt25_11[0]),.doutb(w_asqrt25_11[1]),.doutc(w_asqrt25_11[2]),.din(w_asqrt25_3[1]));
	jspl3 jspl3_w_asqrt25_12(.douta(w_asqrt25_12[0]),.doutb(w_asqrt25_12[1]),.doutc(w_asqrt25_12[2]),.din(w_asqrt25_3[2]));
	jspl3 jspl3_w_asqrt25_13(.douta(w_asqrt25_13[0]),.doutb(w_asqrt25_13[1]),.doutc(w_asqrt25_13[2]),.din(w_asqrt25_4[0]));
	jspl3 jspl3_w_asqrt25_14(.douta(w_asqrt25_14[0]),.doutb(w_asqrt25_14[1]),.doutc(w_asqrt25_14[2]),.din(w_asqrt25_4[1]));
	jspl3 jspl3_w_asqrt25_15(.douta(w_asqrt25_15[0]),.doutb(w_asqrt25_15[1]),.doutc(w_asqrt25_15[2]),.din(w_asqrt25_4[2]));
	jspl3 jspl3_w_asqrt25_16(.douta(w_asqrt25_16[0]),.doutb(w_asqrt25_16[1]),.doutc(w_asqrt25_16[2]),.din(w_asqrt25_5[0]));
	jspl3 jspl3_w_asqrt25_17(.douta(w_asqrt25_17[0]),.doutb(w_asqrt25_17[1]),.doutc(w_asqrt25_17[2]),.din(w_asqrt25_5[1]));
	jspl3 jspl3_w_asqrt25_18(.douta(w_asqrt25_18[0]),.doutb(w_asqrt25_18[1]),.doutc(asqrt[24]),.din(w_asqrt25_5[2]));
	jspl3 jspl3_w_asqrt26_0(.douta(w_asqrt26_0[0]),.doutb(w_asqrt26_0[1]),.doutc(w_asqrt26_0[2]),.din(asqrt_fa_26));
	jspl3 jspl3_w_asqrt26_1(.douta(w_asqrt26_1[0]),.doutb(w_asqrt26_1[1]),.doutc(w_asqrt26_1[2]),.din(w_asqrt26_0[0]));
	jspl3 jspl3_w_asqrt26_2(.douta(w_asqrt26_2[0]),.doutb(w_asqrt26_2[1]),.doutc(w_asqrt26_2[2]),.din(w_asqrt26_0[1]));
	jspl3 jspl3_w_asqrt26_3(.douta(w_asqrt26_3[0]),.doutb(w_asqrt26_3[1]),.doutc(w_asqrt26_3[2]),.din(w_asqrt26_0[2]));
	jspl3 jspl3_w_asqrt26_4(.douta(w_asqrt26_4[0]),.doutb(w_asqrt26_4[1]),.doutc(w_asqrt26_4[2]),.din(w_asqrt26_1[0]));
	jspl3 jspl3_w_asqrt26_5(.douta(w_asqrt26_5[0]),.doutb(w_asqrt26_5[1]),.doutc(w_asqrt26_5[2]),.din(w_asqrt26_1[1]));
	jspl3 jspl3_w_asqrt26_6(.douta(w_asqrt26_6[0]),.doutb(w_asqrt26_6[1]),.doutc(w_asqrt26_6[2]),.din(w_asqrt26_1[2]));
	jspl3 jspl3_w_asqrt26_7(.douta(w_asqrt26_7[0]),.doutb(w_asqrt26_7[1]),.doutc(w_asqrt26_7[2]),.din(w_asqrt26_2[0]));
	jspl3 jspl3_w_asqrt26_8(.douta(w_asqrt26_8[0]),.doutb(w_asqrt26_8[1]),.doutc(w_asqrt26_8[2]),.din(w_asqrt26_2[1]));
	jspl3 jspl3_w_asqrt26_9(.douta(w_asqrt26_9[0]),.doutb(w_asqrt26_9[1]),.doutc(w_asqrt26_9[2]),.din(w_asqrt26_2[2]));
	jspl3 jspl3_w_asqrt26_10(.douta(w_asqrt26_10[0]),.doutb(w_asqrt26_10[1]),.doutc(w_asqrt26_10[2]),.din(w_asqrt26_3[0]));
	jspl3 jspl3_w_asqrt26_11(.douta(w_asqrt26_11[0]),.doutb(w_asqrt26_11[1]),.doutc(w_asqrt26_11[2]),.din(w_asqrt26_3[1]));
	jspl3 jspl3_w_asqrt26_12(.douta(w_asqrt26_12[0]),.doutb(w_asqrt26_12[1]),.doutc(w_asqrt26_12[2]),.din(w_asqrt26_3[2]));
	jspl3 jspl3_w_asqrt26_13(.douta(w_asqrt26_13[0]),.doutb(w_asqrt26_13[1]),.doutc(w_asqrt26_13[2]),.din(w_asqrt26_4[0]));
	jspl3 jspl3_w_asqrt26_14(.douta(w_asqrt26_14[0]),.doutb(w_asqrt26_14[1]),.doutc(w_asqrt26_14[2]),.din(w_asqrt26_4[1]));
	jspl3 jspl3_w_asqrt26_15(.douta(w_asqrt26_15[0]),.doutb(w_asqrt26_15[1]),.doutc(w_asqrt26_15[2]),.din(w_asqrt26_4[2]));
	jspl3 jspl3_w_asqrt26_16(.douta(w_asqrt26_16[0]),.doutb(w_asqrt26_16[1]),.doutc(w_asqrt26_16[2]),.din(w_asqrt26_5[0]));
	jspl3 jspl3_w_asqrt26_17(.douta(w_asqrt26_17[0]),.doutb(w_asqrt26_17[1]),.doutc(w_asqrt26_17[2]),.din(w_asqrt26_5[1]));
	jspl3 jspl3_w_asqrt26_18(.douta(w_asqrt26_18[0]),.doutb(w_asqrt26_18[1]),.doutc(w_asqrt26_18[2]),.din(w_asqrt26_5[2]));
	jspl3 jspl3_w_asqrt26_19(.douta(w_asqrt26_19[0]),.doutb(w_asqrt26_19[1]),.doutc(w_asqrt26_19[2]),.din(w_asqrt26_6[0]));
	jspl3 jspl3_w_asqrt26_20(.douta(w_asqrt26_20[0]),.doutb(w_asqrt26_20[1]),.doutc(w_asqrt26_20[2]),.din(w_asqrt26_6[1]));
	jspl3 jspl3_w_asqrt26_21(.douta(w_asqrt26_21[0]),.doutb(w_asqrt26_21[1]),.doutc(w_asqrt26_21[2]),.din(w_asqrt26_6[2]));
	jspl3 jspl3_w_asqrt26_22(.douta(w_asqrt26_22[0]),.doutb(w_asqrt26_22[1]),.doutc(w_asqrt26_22[2]),.din(w_asqrt26_7[0]));
	jspl3 jspl3_w_asqrt26_23(.douta(w_asqrt26_23[0]),.doutb(w_asqrt26_23[1]),.doutc(w_asqrt26_23[2]),.din(w_asqrt26_7[1]));
	jspl3 jspl3_w_asqrt26_24(.douta(w_asqrt26_24[0]),.doutb(w_asqrt26_24[1]),.doutc(w_asqrt26_24[2]),.din(w_asqrt26_7[2]));
	jspl3 jspl3_w_asqrt26_25(.douta(w_asqrt26_25[0]),.doutb(w_asqrt26_25[1]),.doutc(w_asqrt26_25[2]),.din(w_asqrt26_8[0]));
	jspl3 jspl3_w_asqrt26_26(.douta(w_asqrt26_26[0]),.doutb(w_asqrt26_26[1]),.doutc(w_asqrt26_26[2]),.din(w_asqrt26_8[1]));
	jspl3 jspl3_w_asqrt26_27(.douta(w_asqrt26_27[0]),.doutb(w_asqrt26_27[1]),.doutc(w_asqrt26_27[2]),.din(w_asqrt26_8[2]));
	jspl3 jspl3_w_asqrt26_28(.douta(w_asqrt26_28[0]),.doutb(w_asqrt26_28[1]),.doutc(w_asqrt26_28[2]),.din(w_asqrt26_9[0]));
	jspl3 jspl3_w_asqrt26_29(.douta(w_asqrt26_29[0]),.doutb(w_asqrt26_29[1]),.doutc(w_asqrt26_29[2]),.din(w_asqrt26_9[1]));
	jspl3 jspl3_w_asqrt26_30(.douta(w_asqrt26_30[0]),.doutb(w_asqrt26_30[1]),.doutc(w_asqrt26_30[2]),.din(w_asqrt26_9[2]));
	jspl3 jspl3_w_asqrt26_31(.douta(w_asqrt26_31[0]),.doutb(w_asqrt26_31[1]),.doutc(w_asqrt26_31[2]),.din(w_asqrt26_10[0]));
	jspl3 jspl3_w_asqrt26_32(.douta(w_asqrt26_32[0]),.doutb(w_asqrt26_32[1]),.doutc(w_asqrt26_32[2]),.din(w_asqrt26_10[1]));
	jspl3 jspl3_w_asqrt26_33(.douta(w_asqrt26_33[0]),.doutb(w_asqrt26_33[1]),.doutc(w_asqrt26_33[2]),.din(w_asqrt26_10[2]));
	jspl3 jspl3_w_asqrt26_34(.douta(w_asqrt26_34[0]),.doutb(w_asqrt26_34[1]),.doutc(w_asqrt26_34[2]),.din(w_asqrt26_11[0]));
	jspl3 jspl3_w_asqrt26_35(.douta(w_asqrt26_35[0]),.doutb(w_asqrt26_35[1]),.doutc(w_asqrt26_35[2]),.din(w_asqrt26_11[1]));
	jspl3 jspl3_w_asqrt26_36(.douta(w_asqrt26_36[0]),.doutb(w_asqrt26_36[1]),.doutc(asqrt[25]),.din(w_asqrt26_11[2]));
	jspl3 jspl3_w_asqrt27_0(.douta(w_asqrt27_0[0]),.doutb(w_asqrt27_0[1]),.doutc(w_asqrt27_0[2]),.din(asqrt_fa_27));
	jspl3 jspl3_w_asqrt27_1(.douta(w_asqrt27_1[0]),.doutb(w_asqrt27_1[1]),.doutc(w_asqrt27_1[2]),.din(w_asqrt27_0[0]));
	jspl3 jspl3_w_asqrt27_2(.douta(w_asqrt27_2[0]),.doutb(w_asqrt27_2[1]),.doutc(w_asqrt27_2[2]),.din(w_asqrt27_0[1]));
	jspl3 jspl3_w_asqrt27_3(.douta(w_asqrt27_3[0]),.doutb(w_asqrt27_3[1]),.doutc(w_asqrt27_3[2]),.din(w_asqrt27_0[2]));
	jspl3 jspl3_w_asqrt27_4(.douta(w_asqrt27_4[0]),.doutb(w_asqrt27_4[1]),.doutc(w_asqrt27_4[2]),.din(w_asqrt27_1[0]));
	jspl3 jspl3_w_asqrt27_5(.douta(w_asqrt27_5[0]),.doutb(w_asqrt27_5[1]),.doutc(w_asqrt27_5[2]),.din(w_asqrt27_1[1]));
	jspl3 jspl3_w_asqrt27_6(.douta(w_asqrt27_6[0]),.doutb(w_asqrt27_6[1]),.doutc(w_asqrt27_6[2]),.din(w_asqrt27_1[2]));
	jspl3 jspl3_w_asqrt27_7(.douta(w_asqrt27_7[0]),.doutb(w_asqrt27_7[1]),.doutc(w_asqrt27_7[2]),.din(w_asqrt27_2[0]));
	jspl3 jspl3_w_asqrt27_8(.douta(w_asqrt27_8[0]),.doutb(w_asqrt27_8[1]),.doutc(w_asqrt27_8[2]),.din(w_asqrt27_2[1]));
	jspl3 jspl3_w_asqrt27_9(.douta(w_asqrt27_9[0]),.doutb(w_asqrt27_9[1]),.doutc(w_asqrt27_9[2]),.din(w_asqrt27_2[2]));
	jspl3 jspl3_w_asqrt27_10(.douta(w_asqrt27_10[0]),.doutb(w_asqrt27_10[1]),.doutc(w_asqrt27_10[2]),.din(w_asqrt27_3[0]));
	jspl3 jspl3_w_asqrt27_11(.douta(w_asqrt27_11[0]),.doutb(w_asqrt27_11[1]),.doutc(w_asqrt27_11[2]),.din(w_asqrt27_3[1]));
	jspl3 jspl3_w_asqrt27_12(.douta(w_asqrt27_12[0]),.doutb(w_asqrt27_12[1]),.doutc(w_asqrt27_12[2]),.din(w_asqrt27_3[2]));
	jspl3 jspl3_w_asqrt27_13(.douta(w_asqrt27_13[0]),.doutb(w_asqrt27_13[1]),.doutc(w_asqrt27_13[2]),.din(w_asqrt27_4[0]));
	jspl3 jspl3_w_asqrt27_14(.douta(w_asqrt27_14[0]),.doutb(w_asqrt27_14[1]),.doutc(w_asqrt27_14[2]),.din(w_asqrt27_4[1]));
	jspl3 jspl3_w_asqrt27_15(.douta(w_asqrt27_15[0]),.doutb(w_asqrt27_15[1]),.doutc(w_asqrt27_15[2]),.din(w_asqrt27_4[2]));
	jspl3 jspl3_w_asqrt27_16(.douta(w_asqrt27_16[0]),.doutb(w_asqrt27_16[1]),.doutc(w_asqrt27_16[2]),.din(w_asqrt27_5[0]));
	jspl3 jspl3_w_asqrt27_17(.douta(w_asqrt27_17[0]),.doutb(w_asqrt27_17[1]),.doutc(w_asqrt27_17[2]),.din(w_asqrt27_5[1]));
	jspl3 jspl3_w_asqrt27_18(.douta(w_asqrt27_18[0]),.doutb(w_asqrt27_18[1]),.doutc(w_asqrt27_18[2]),.din(w_asqrt27_5[2]));
	jspl3 jspl3_w_asqrt27_19(.douta(w_asqrt27_19[0]),.doutb(w_asqrt27_19[1]),.doutc(w_asqrt27_19[2]),.din(w_asqrt27_6[0]));
	jspl3 jspl3_w_asqrt27_20(.douta(w_asqrt27_20[0]),.doutb(w_asqrt27_20[1]),.doutc(asqrt[26]),.din(w_asqrt27_6[1]));
	jspl3 jspl3_w_asqrt28_0(.douta(w_asqrt28_0[0]),.doutb(w_asqrt28_0[1]),.doutc(w_asqrt28_0[2]),.din(asqrt_fa_28));
	jspl3 jspl3_w_asqrt28_1(.douta(w_asqrt28_1[0]),.doutb(w_asqrt28_1[1]),.doutc(w_asqrt28_1[2]),.din(w_asqrt28_0[0]));
	jspl3 jspl3_w_asqrt28_2(.douta(w_asqrt28_2[0]),.doutb(w_asqrt28_2[1]),.doutc(w_asqrt28_2[2]),.din(w_asqrt28_0[1]));
	jspl3 jspl3_w_asqrt28_3(.douta(w_asqrt28_3[0]),.doutb(w_asqrt28_3[1]),.doutc(w_asqrt28_3[2]),.din(w_asqrt28_0[2]));
	jspl3 jspl3_w_asqrt28_4(.douta(w_asqrt28_4[0]),.doutb(w_asqrt28_4[1]),.doutc(w_asqrt28_4[2]),.din(w_asqrt28_1[0]));
	jspl3 jspl3_w_asqrt28_5(.douta(w_asqrt28_5[0]),.doutb(w_asqrt28_5[1]),.doutc(w_asqrt28_5[2]),.din(w_asqrt28_1[1]));
	jspl3 jspl3_w_asqrt28_6(.douta(w_asqrt28_6[0]),.doutb(w_asqrt28_6[1]),.doutc(w_asqrt28_6[2]),.din(w_asqrt28_1[2]));
	jspl3 jspl3_w_asqrt28_7(.douta(w_asqrt28_7[0]),.doutb(w_asqrt28_7[1]),.doutc(w_asqrt28_7[2]),.din(w_asqrt28_2[0]));
	jspl3 jspl3_w_asqrt28_8(.douta(w_asqrt28_8[0]),.doutb(w_asqrt28_8[1]),.doutc(w_asqrt28_8[2]),.din(w_asqrt28_2[1]));
	jspl3 jspl3_w_asqrt28_9(.douta(w_asqrt28_9[0]),.doutb(w_asqrt28_9[1]),.doutc(w_asqrt28_9[2]),.din(w_asqrt28_2[2]));
	jspl3 jspl3_w_asqrt28_10(.douta(w_asqrt28_10[0]),.doutb(w_asqrt28_10[1]),.doutc(w_asqrt28_10[2]),.din(w_asqrt28_3[0]));
	jspl3 jspl3_w_asqrt28_11(.douta(w_asqrt28_11[0]),.doutb(w_asqrt28_11[1]),.doutc(w_asqrt28_11[2]),.din(w_asqrt28_3[1]));
	jspl3 jspl3_w_asqrt28_12(.douta(w_asqrt28_12[0]),.doutb(w_asqrt28_12[1]),.doutc(w_asqrt28_12[2]),.din(w_asqrt28_3[2]));
	jspl3 jspl3_w_asqrt28_13(.douta(w_asqrt28_13[0]),.doutb(w_asqrt28_13[1]),.doutc(w_asqrt28_13[2]),.din(w_asqrt28_4[0]));
	jspl3 jspl3_w_asqrt28_14(.douta(w_asqrt28_14[0]),.doutb(w_asqrt28_14[1]),.doutc(w_asqrt28_14[2]),.din(w_asqrt28_4[1]));
	jspl3 jspl3_w_asqrt28_15(.douta(w_asqrt28_15[0]),.doutb(w_asqrt28_15[1]),.doutc(w_asqrt28_15[2]),.din(w_asqrt28_4[2]));
	jspl3 jspl3_w_asqrt28_16(.douta(w_asqrt28_16[0]),.doutb(w_asqrt28_16[1]),.doutc(w_asqrt28_16[2]),.din(w_asqrt28_5[0]));
	jspl3 jspl3_w_asqrt28_17(.douta(w_asqrt28_17[0]),.doutb(w_asqrt28_17[1]),.doutc(w_asqrt28_17[2]),.din(w_asqrt28_5[1]));
	jspl3 jspl3_w_asqrt28_18(.douta(w_asqrt28_18[0]),.doutb(w_asqrt28_18[1]),.doutc(w_asqrt28_18[2]),.din(w_asqrt28_5[2]));
	jspl3 jspl3_w_asqrt28_19(.douta(w_asqrt28_19[0]),.doutb(w_asqrt28_19[1]),.doutc(w_asqrt28_19[2]),.din(w_asqrt28_6[0]));
	jspl3 jspl3_w_asqrt28_20(.douta(w_asqrt28_20[0]),.doutb(w_asqrt28_20[1]),.doutc(w_asqrt28_20[2]),.din(w_asqrt28_6[1]));
	jspl3 jspl3_w_asqrt28_21(.douta(w_asqrt28_21[0]),.doutb(w_asqrt28_21[1]),.doutc(w_asqrt28_21[2]),.din(w_asqrt28_6[2]));
	jspl3 jspl3_w_asqrt28_22(.douta(w_asqrt28_22[0]),.doutb(w_asqrt28_22[1]),.doutc(w_asqrt28_22[2]),.din(w_asqrt28_7[0]));
	jspl3 jspl3_w_asqrt28_23(.douta(w_asqrt28_23[0]),.doutb(w_asqrt28_23[1]),.doutc(w_asqrt28_23[2]),.din(w_asqrt28_7[1]));
	jspl3 jspl3_w_asqrt28_24(.douta(w_asqrt28_24[0]),.doutb(w_asqrt28_24[1]),.doutc(w_asqrt28_24[2]),.din(w_asqrt28_7[2]));
	jspl3 jspl3_w_asqrt28_25(.douta(w_asqrt28_25[0]),.doutb(w_asqrt28_25[1]),.doutc(w_asqrt28_25[2]),.din(w_asqrt28_8[0]));
	jspl3 jspl3_w_asqrt28_26(.douta(w_asqrt28_26[0]),.doutb(w_asqrt28_26[1]),.doutc(w_asqrt28_26[2]),.din(w_asqrt28_8[1]));
	jspl3 jspl3_w_asqrt28_27(.douta(w_asqrt28_27[0]),.doutb(w_asqrt28_27[1]),.doutc(w_asqrt28_27[2]),.din(w_asqrt28_8[2]));
	jspl3 jspl3_w_asqrt28_28(.douta(w_asqrt28_28[0]),.doutb(w_asqrt28_28[1]),.doutc(w_asqrt28_28[2]),.din(w_asqrt28_9[0]));
	jspl3 jspl3_w_asqrt28_29(.douta(w_asqrt28_29[0]),.doutb(w_asqrt28_29[1]),.doutc(w_asqrt28_29[2]),.din(w_asqrt28_9[1]));
	jspl3 jspl3_w_asqrt28_30(.douta(w_asqrt28_30[0]),.doutb(w_asqrt28_30[1]),.doutc(w_asqrt28_30[2]),.din(w_asqrt28_9[2]));
	jspl3 jspl3_w_asqrt28_31(.douta(w_asqrt28_31[0]),.doutb(w_asqrt28_31[1]),.doutc(w_asqrt28_31[2]),.din(w_asqrt28_10[0]));
	jspl3 jspl3_w_asqrt28_32(.douta(w_asqrt28_32[0]),.doutb(w_asqrt28_32[1]),.doutc(w_asqrt28_32[2]),.din(w_asqrt28_10[1]));
	jspl3 jspl3_w_asqrt28_33(.douta(w_asqrt28_33[0]),.doutb(w_asqrt28_33[1]),.doutc(w_asqrt28_33[2]),.din(w_asqrt28_10[2]));
	jspl3 jspl3_w_asqrt28_34(.douta(w_asqrt28_34[0]),.doutb(w_asqrt28_34[1]),.doutc(w_asqrt28_34[2]),.din(w_asqrt28_11[0]));
	jspl3 jspl3_w_asqrt28_35(.douta(w_asqrt28_35[0]),.doutb(w_asqrt28_35[1]),.doutc(w_asqrt28_35[2]),.din(w_asqrt28_11[1]));
	jspl3 jspl3_w_asqrt28_36(.douta(w_asqrt28_36[0]),.doutb(w_asqrt28_36[1]),.doutc(w_asqrt28_36[2]),.din(w_asqrt28_11[2]));
	jspl3 jspl3_w_asqrt28_37(.douta(w_asqrt28_37[0]),.doutb(w_asqrt28_37[1]),.doutc(asqrt[27]),.din(w_asqrt28_12[0]));
	jspl3 jspl3_w_asqrt29_0(.douta(w_asqrt29_0[0]),.doutb(w_asqrt29_0[1]),.doutc(w_asqrt29_0[2]),.din(asqrt_fa_29));
	jspl3 jspl3_w_asqrt29_1(.douta(w_asqrt29_1[0]),.doutb(w_asqrt29_1[1]),.doutc(w_asqrt29_1[2]),.din(w_asqrt29_0[0]));
	jspl3 jspl3_w_asqrt29_2(.douta(w_asqrt29_2[0]),.doutb(w_asqrt29_2[1]),.doutc(w_asqrt29_2[2]),.din(w_asqrt29_0[1]));
	jspl3 jspl3_w_asqrt29_3(.douta(w_asqrt29_3[0]),.doutb(w_asqrt29_3[1]),.doutc(w_asqrt29_3[2]),.din(w_asqrt29_0[2]));
	jspl3 jspl3_w_asqrt29_4(.douta(w_asqrt29_4[0]),.doutb(w_asqrt29_4[1]),.doutc(w_asqrt29_4[2]),.din(w_asqrt29_1[0]));
	jspl3 jspl3_w_asqrt29_5(.douta(w_asqrt29_5[0]),.doutb(w_asqrt29_5[1]),.doutc(w_asqrt29_5[2]),.din(w_asqrt29_1[1]));
	jspl3 jspl3_w_asqrt29_6(.douta(w_asqrt29_6[0]),.doutb(w_asqrt29_6[1]),.doutc(w_asqrt29_6[2]),.din(w_asqrt29_1[2]));
	jspl3 jspl3_w_asqrt29_7(.douta(w_asqrt29_7[0]),.doutb(w_asqrt29_7[1]),.doutc(w_asqrt29_7[2]),.din(w_asqrt29_2[0]));
	jspl3 jspl3_w_asqrt29_8(.douta(w_asqrt29_8[0]),.doutb(w_asqrt29_8[1]),.doutc(w_asqrt29_8[2]),.din(w_asqrt29_2[1]));
	jspl3 jspl3_w_asqrt29_9(.douta(w_asqrt29_9[0]),.doutb(w_asqrt29_9[1]),.doutc(w_asqrt29_9[2]),.din(w_asqrt29_2[2]));
	jspl3 jspl3_w_asqrt29_10(.douta(w_asqrt29_10[0]),.doutb(w_asqrt29_10[1]),.doutc(w_asqrt29_10[2]),.din(w_asqrt29_3[0]));
	jspl3 jspl3_w_asqrt29_11(.douta(w_asqrt29_11[0]),.doutb(w_asqrt29_11[1]),.doutc(w_asqrt29_11[2]),.din(w_asqrt29_3[1]));
	jspl3 jspl3_w_asqrt29_12(.douta(w_asqrt29_12[0]),.doutb(w_asqrt29_12[1]),.doutc(w_asqrt29_12[2]),.din(w_asqrt29_3[2]));
	jspl3 jspl3_w_asqrt29_13(.douta(w_asqrt29_13[0]),.doutb(w_asqrt29_13[1]),.doutc(w_asqrt29_13[2]),.din(w_asqrt29_4[0]));
	jspl3 jspl3_w_asqrt29_14(.douta(w_asqrt29_14[0]),.doutb(w_asqrt29_14[1]),.doutc(w_asqrt29_14[2]),.din(w_asqrt29_4[1]));
	jspl3 jspl3_w_asqrt29_15(.douta(w_asqrt29_15[0]),.doutb(w_asqrt29_15[1]),.doutc(w_asqrt29_15[2]),.din(w_asqrt29_4[2]));
	jspl3 jspl3_w_asqrt29_16(.douta(w_asqrt29_16[0]),.doutb(w_asqrt29_16[1]),.doutc(w_asqrt29_16[2]),.din(w_asqrt29_5[0]));
	jspl3 jspl3_w_asqrt29_17(.douta(w_asqrt29_17[0]),.doutb(w_asqrt29_17[1]),.doutc(w_asqrt29_17[2]),.din(w_asqrt29_5[1]));
	jspl3 jspl3_w_asqrt29_18(.douta(w_asqrt29_18[0]),.doutb(w_asqrt29_18[1]),.doutc(w_asqrt29_18[2]),.din(w_asqrt29_5[2]));
	jspl3 jspl3_w_asqrt29_19(.douta(w_asqrt29_19[0]),.doutb(w_asqrt29_19[1]),.doutc(w_asqrt29_19[2]),.din(w_asqrt29_6[0]));
	jspl3 jspl3_w_asqrt29_20(.douta(w_asqrt29_20[0]),.doutb(w_asqrt29_20[1]),.doutc(w_asqrt29_20[2]),.din(w_asqrt29_6[1]));
	jspl3 jspl3_w_asqrt29_21(.douta(w_asqrt29_21[0]),.doutb(w_asqrt29_21[1]),.doutc(asqrt[28]),.din(w_asqrt29_6[2]));
	jspl3 jspl3_w_asqrt30_0(.douta(w_asqrt30_0[0]),.doutb(w_asqrt30_0[1]),.doutc(w_asqrt30_0[2]),.din(asqrt_fa_30));
	jspl3 jspl3_w_asqrt30_1(.douta(w_asqrt30_1[0]),.doutb(w_asqrt30_1[1]),.doutc(w_asqrt30_1[2]),.din(w_asqrt30_0[0]));
	jspl3 jspl3_w_asqrt30_2(.douta(w_asqrt30_2[0]),.doutb(w_asqrt30_2[1]),.doutc(w_asqrt30_2[2]),.din(w_asqrt30_0[1]));
	jspl3 jspl3_w_asqrt30_3(.douta(w_asqrt30_3[0]),.doutb(w_asqrt30_3[1]),.doutc(w_asqrt30_3[2]),.din(w_asqrt30_0[2]));
	jspl3 jspl3_w_asqrt30_4(.douta(w_asqrt30_4[0]),.doutb(w_asqrt30_4[1]),.doutc(w_asqrt30_4[2]),.din(w_asqrt30_1[0]));
	jspl3 jspl3_w_asqrt30_5(.douta(w_asqrt30_5[0]),.doutb(w_asqrt30_5[1]),.doutc(w_asqrt30_5[2]),.din(w_asqrt30_1[1]));
	jspl3 jspl3_w_asqrt30_6(.douta(w_asqrt30_6[0]),.doutb(w_asqrt30_6[1]),.doutc(w_asqrt30_6[2]),.din(w_asqrt30_1[2]));
	jspl3 jspl3_w_asqrt30_7(.douta(w_asqrt30_7[0]),.doutb(w_asqrt30_7[1]),.doutc(w_asqrt30_7[2]),.din(w_asqrt30_2[0]));
	jspl3 jspl3_w_asqrt30_8(.douta(w_asqrt30_8[0]),.doutb(w_asqrt30_8[1]),.doutc(w_asqrt30_8[2]),.din(w_asqrt30_2[1]));
	jspl3 jspl3_w_asqrt30_9(.douta(w_asqrt30_9[0]),.doutb(w_asqrt30_9[1]),.doutc(w_asqrt30_9[2]),.din(w_asqrt30_2[2]));
	jspl3 jspl3_w_asqrt30_10(.douta(w_asqrt30_10[0]),.doutb(w_asqrt30_10[1]),.doutc(w_asqrt30_10[2]),.din(w_asqrt30_3[0]));
	jspl3 jspl3_w_asqrt30_11(.douta(w_asqrt30_11[0]),.doutb(w_asqrt30_11[1]),.doutc(w_asqrt30_11[2]),.din(w_asqrt30_3[1]));
	jspl3 jspl3_w_asqrt30_12(.douta(w_asqrt30_12[0]),.doutb(w_asqrt30_12[1]),.doutc(w_asqrt30_12[2]),.din(w_asqrt30_3[2]));
	jspl3 jspl3_w_asqrt30_13(.douta(w_asqrt30_13[0]),.doutb(w_asqrt30_13[1]),.doutc(w_asqrt30_13[2]),.din(w_asqrt30_4[0]));
	jspl3 jspl3_w_asqrt30_14(.douta(w_asqrt30_14[0]),.doutb(w_asqrt30_14[1]),.doutc(w_asqrt30_14[2]),.din(w_asqrt30_4[1]));
	jspl3 jspl3_w_asqrt30_15(.douta(w_asqrt30_15[0]),.doutb(w_asqrt30_15[1]),.doutc(w_asqrt30_15[2]),.din(w_asqrt30_4[2]));
	jspl3 jspl3_w_asqrt30_16(.douta(w_asqrt30_16[0]),.doutb(w_asqrt30_16[1]),.doutc(w_asqrt30_16[2]),.din(w_asqrt30_5[0]));
	jspl3 jspl3_w_asqrt30_17(.douta(w_asqrt30_17[0]),.doutb(w_asqrt30_17[1]),.doutc(w_asqrt30_17[2]),.din(w_asqrt30_5[1]));
	jspl3 jspl3_w_asqrt30_18(.douta(w_asqrt30_18[0]),.doutb(w_asqrt30_18[1]),.doutc(w_asqrt30_18[2]),.din(w_asqrt30_5[2]));
	jspl3 jspl3_w_asqrt30_19(.douta(w_asqrt30_19[0]),.doutb(w_asqrt30_19[1]),.doutc(w_asqrt30_19[2]),.din(w_asqrt30_6[0]));
	jspl3 jspl3_w_asqrt30_20(.douta(w_asqrt30_20[0]),.doutb(w_asqrt30_20[1]),.doutc(w_asqrt30_20[2]),.din(w_asqrt30_6[1]));
	jspl3 jspl3_w_asqrt30_21(.douta(w_asqrt30_21[0]),.doutb(w_asqrt30_21[1]),.doutc(w_asqrt30_21[2]),.din(w_asqrt30_6[2]));
	jspl3 jspl3_w_asqrt30_22(.douta(w_asqrt30_22[0]),.doutb(w_asqrt30_22[1]),.doutc(w_asqrt30_22[2]),.din(w_asqrt30_7[0]));
	jspl3 jspl3_w_asqrt30_23(.douta(w_asqrt30_23[0]),.doutb(w_asqrt30_23[1]),.doutc(w_asqrt30_23[2]),.din(w_asqrt30_7[1]));
	jspl3 jspl3_w_asqrt30_24(.douta(w_asqrt30_24[0]),.doutb(w_asqrt30_24[1]),.doutc(w_asqrt30_24[2]),.din(w_asqrt30_7[2]));
	jspl3 jspl3_w_asqrt30_25(.douta(w_asqrt30_25[0]),.doutb(w_asqrt30_25[1]),.doutc(w_asqrt30_25[2]),.din(w_asqrt30_8[0]));
	jspl3 jspl3_w_asqrt30_26(.douta(w_asqrt30_26[0]),.doutb(w_asqrt30_26[1]),.doutc(w_asqrt30_26[2]),.din(w_asqrt30_8[1]));
	jspl3 jspl3_w_asqrt30_27(.douta(w_asqrt30_27[0]),.doutb(w_asqrt30_27[1]),.doutc(w_asqrt30_27[2]),.din(w_asqrt30_8[2]));
	jspl3 jspl3_w_asqrt30_28(.douta(w_asqrt30_28[0]),.doutb(w_asqrt30_28[1]),.doutc(w_asqrt30_28[2]),.din(w_asqrt30_9[0]));
	jspl3 jspl3_w_asqrt30_29(.douta(w_asqrt30_29[0]),.doutb(w_asqrt30_29[1]),.doutc(w_asqrt30_29[2]),.din(w_asqrt30_9[1]));
	jspl3 jspl3_w_asqrt30_30(.douta(w_asqrt30_30[0]),.doutb(w_asqrt30_30[1]),.doutc(w_asqrt30_30[2]),.din(w_asqrt30_9[2]));
	jspl3 jspl3_w_asqrt30_31(.douta(w_asqrt30_31[0]),.doutb(w_asqrt30_31[1]),.doutc(w_asqrt30_31[2]),.din(w_asqrt30_10[0]));
	jspl3 jspl3_w_asqrt30_32(.douta(w_asqrt30_32[0]),.doutb(w_asqrt30_32[1]),.doutc(w_asqrt30_32[2]),.din(w_asqrt30_10[1]));
	jspl3 jspl3_w_asqrt30_33(.douta(w_asqrt30_33[0]),.doutb(w_asqrt30_33[1]),.doutc(w_asqrt30_33[2]),.din(w_asqrt30_10[2]));
	jspl3 jspl3_w_asqrt30_34(.douta(w_asqrt30_34[0]),.doutb(w_asqrt30_34[1]),.doutc(w_asqrt30_34[2]),.din(w_asqrt30_11[0]));
	jspl3 jspl3_w_asqrt30_35(.douta(w_asqrt30_35[0]),.doutb(w_asqrt30_35[1]),.doutc(w_asqrt30_35[2]),.din(w_asqrt30_11[1]));
	jspl3 jspl3_w_asqrt30_36(.douta(w_asqrt30_36[0]),.doutb(w_asqrt30_36[1]),.doutc(w_asqrt30_36[2]),.din(w_asqrt30_11[2]));
	jspl3 jspl3_w_asqrt30_37(.douta(w_asqrt30_37[0]),.doutb(w_asqrt30_37[1]),.doutc(w_asqrt30_37[2]),.din(w_asqrt30_12[0]));
	jspl jspl_w_asqrt30_38(.douta(w_asqrt30_38),.doutb(asqrt[29]),.din(w_asqrt30_12[1]));
	jspl3 jspl3_w_asqrt31_0(.douta(w_asqrt31_0[0]),.doutb(w_asqrt31_0[1]),.doutc(w_asqrt31_0[2]),.din(asqrt_fa_31));
	jspl3 jspl3_w_asqrt31_1(.douta(w_asqrt31_1[0]),.doutb(w_asqrt31_1[1]),.doutc(w_asqrt31_1[2]),.din(w_asqrt31_0[0]));
	jspl3 jspl3_w_asqrt31_2(.douta(w_asqrt31_2[0]),.doutb(w_asqrt31_2[1]),.doutc(w_asqrt31_2[2]),.din(w_asqrt31_0[1]));
	jspl3 jspl3_w_asqrt31_3(.douta(w_asqrt31_3[0]),.doutb(w_asqrt31_3[1]),.doutc(w_asqrt31_3[2]),.din(w_asqrt31_0[2]));
	jspl3 jspl3_w_asqrt31_4(.douta(w_asqrt31_4[0]),.doutb(w_asqrt31_4[1]),.doutc(w_asqrt31_4[2]),.din(w_asqrt31_1[0]));
	jspl3 jspl3_w_asqrt31_5(.douta(w_asqrt31_5[0]),.doutb(w_asqrt31_5[1]),.doutc(w_asqrt31_5[2]),.din(w_asqrt31_1[1]));
	jspl3 jspl3_w_asqrt31_6(.douta(w_asqrt31_6[0]),.doutb(w_asqrt31_6[1]),.doutc(w_asqrt31_6[2]),.din(w_asqrt31_1[2]));
	jspl3 jspl3_w_asqrt31_7(.douta(w_asqrt31_7[0]),.doutb(w_asqrt31_7[1]),.doutc(w_asqrt31_7[2]),.din(w_asqrt31_2[0]));
	jspl3 jspl3_w_asqrt31_8(.douta(w_asqrt31_8[0]),.doutb(w_asqrt31_8[1]),.doutc(w_asqrt31_8[2]),.din(w_asqrt31_2[1]));
	jspl3 jspl3_w_asqrt31_9(.douta(w_asqrt31_9[0]),.doutb(w_asqrt31_9[1]),.doutc(w_asqrt31_9[2]),.din(w_asqrt31_2[2]));
	jspl3 jspl3_w_asqrt31_10(.douta(w_asqrt31_10[0]),.doutb(w_asqrt31_10[1]),.doutc(w_asqrt31_10[2]),.din(w_asqrt31_3[0]));
	jspl3 jspl3_w_asqrt31_11(.douta(w_asqrt31_11[0]),.doutb(w_asqrt31_11[1]),.doutc(w_asqrt31_11[2]),.din(w_asqrt31_3[1]));
	jspl3 jspl3_w_asqrt31_12(.douta(w_asqrt31_12[0]),.doutb(w_asqrt31_12[1]),.doutc(w_asqrt31_12[2]),.din(w_asqrt31_3[2]));
	jspl3 jspl3_w_asqrt31_13(.douta(w_asqrt31_13[0]),.doutb(w_asqrt31_13[1]),.doutc(w_asqrt31_13[2]),.din(w_asqrt31_4[0]));
	jspl3 jspl3_w_asqrt31_14(.douta(w_asqrt31_14[0]),.doutb(w_asqrt31_14[1]),.doutc(w_asqrt31_14[2]),.din(w_asqrt31_4[1]));
	jspl3 jspl3_w_asqrt31_15(.douta(w_asqrt31_15[0]),.doutb(w_asqrt31_15[1]),.doutc(w_asqrt31_15[2]),.din(w_asqrt31_4[2]));
	jspl3 jspl3_w_asqrt31_16(.douta(w_asqrt31_16[0]),.doutb(w_asqrt31_16[1]),.doutc(w_asqrt31_16[2]),.din(w_asqrt31_5[0]));
	jspl3 jspl3_w_asqrt31_17(.douta(w_asqrt31_17[0]),.doutb(w_asqrt31_17[1]),.doutc(w_asqrt31_17[2]),.din(w_asqrt31_5[1]));
	jspl3 jspl3_w_asqrt31_18(.douta(w_asqrt31_18[0]),.doutb(w_asqrt31_18[1]),.doutc(w_asqrt31_18[2]),.din(w_asqrt31_5[2]));
	jspl3 jspl3_w_asqrt31_19(.douta(w_asqrt31_19[0]),.doutb(w_asqrt31_19[1]),.doutc(w_asqrt31_19[2]),.din(w_asqrt31_6[0]));
	jspl3 jspl3_w_asqrt31_20(.douta(w_asqrt31_20[0]),.doutb(w_asqrt31_20[1]),.doutc(w_asqrt31_20[2]),.din(w_asqrt31_6[1]));
	jspl3 jspl3_w_asqrt31_21(.douta(w_asqrt31_21[0]),.doutb(w_asqrt31_21[1]),.doutc(w_asqrt31_21[2]),.din(w_asqrt31_6[2]));
	jspl3 jspl3_w_asqrt31_22(.douta(w_asqrt31_22[0]),.doutb(w_asqrt31_22[1]),.doutc(w_asqrt31_22[2]),.din(w_asqrt31_7[0]));
	jspl jspl_w_asqrt31_23(.douta(w_asqrt31_23),.doutb(asqrt[30]),.din(w_asqrt31_7[1]));
	jspl3 jspl3_w_asqrt32_0(.douta(w_asqrt32_0[0]),.doutb(w_asqrt32_0[1]),.doutc(w_asqrt32_0[2]),.din(asqrt_fa_32));
	jspl3 jspl3_w_asqrt32_1(.douta(w_asqrt32_1[0]),.doutb(w_asqrt32_1[1]),.doutc(w_asqrt32_1[2]),.din(w_asqrt32_0[0]));
	jspl3 jspl3_w_asqrt32_2(.douta(w_asqrt32_2[0]),.doutb(w_asqrt32_2[1]),.doutc(w_asqrt32_2[2]),.din(w_asqrt32_0[1]));
	jspl3 jspl3_w_asqrt32_3(.douta(w_asqrt32_3[0]),.doutb(w_asqrt32_3[1]),.doutc(w_asqrt32_3[2]),.din(w_asqrt32_0[2]));
	jspl3 jspl3_w_asqrt32_4(.douta(w_asqrt32_4[0]),.doutb(w_asqrt32_4[1]),.doutc(w_asqrt32_4[2]),.din(w_asqrt32_1[0]));
	jspl3 jspl3_w_asqrt32_5(.douta(w_asqrt32_5[0]),.doutb(w_asqrt32_5[1]),.doutc(w_asqrt32_5[2]),.din(w_asqrt32_1[1]));
	jspl3 jspl3_w_asqrt32_6(.douta(w_asqrt32_6[0]),.doutb(w_asqrt32_6[1]),.doutc(w_asqrt32_6[2]),.din(w_asqrt32_1[2]));
	jspl3 jspl3_w_asqrt32_7(.douta(w_asqrt32_7[0]),.doutb(w_asqrt32_7[1]),.doutc(w_asqrt32_7[2]),.din(w_asqrt32_2[0]));
	jspl3 jspl3_w_asqrt32_8(.douta(w_asqrt32_8[0]),.doutb(w_asqrt32_8[1]),.doutc(w_asqrt32_8[2]),.din(w_asqrt32_2[1]));
	jspl3 jspl3_w_asqrt32_9(.douta(w_asqrt32_9[0]),.doutb(w_asqrt32_9[1]),.doutc(w_asqrt32_9[2]),.din(w_asqrt32_2[2]));
	jspl3 jspl3_w_asqrt32_10(.douta(w_asqrt32_10[0]),.doutb(w_asqrt32_10[1]),.doutc(w_asqrt32_10[2]),.din(w_asqrt32_3[0]));
	jspl3 jspl3_w_asqrt32_11(.douta(w_asqrt32_11[0]),.doutb(w_asqrt32_11[1]),.doutc(w_asqrt32_11[2]),.din(w_asqrt32_3[1]));
	jspl3 jspl3_w_asqrt32_12(.douta(w_asqrt32_12[0]),.doutb(w_asqrt32_12[1]),.doutc(w_asqrt32_12[2]),.din(w_asqrt32_3[2]));
	jspl3 jspl3_w_asqrt32_13(.douta(w_asqrt32_13[0]),.doutb(w_asqrt32_13[1]),.doutc(w_asqrt32_13[2]),.din(w_asqrt32_4[0]));
	jspl3 jspl3_w_asqrt32_14(.douta(w_asqrt32_14[0]),.doutb(w_asqrt32_14[1]),.doutc(w_asqrt32_14[2]),.din(w_asqrt32_4[1]));
	jspl3 jspl3_w_asqrt32_15(.douta(w_asqrt32_15[0]),.doutb(w_asqrt32_15[1]),.doutc(w_asqrt32_15[2]),.din(w_asqrt32_4[2]));
	jspl3 jspl3_w_asqrt32_16(.douta(w_asqrt32_16[0]),.doutb(w_asqrt32_16[1]),.doutc(w_asqrt32_16[2]),.din(w_asqrt32_5[0]));
	jspl3 jspl3_w_asqrt32_17(.douta(w_asqrt32_17[0]),.doutb(w_asqrt32_17[1]),.doutc(w_asqrt32_17[2]),.din(w_asqrt32_5[1]));
	jspl3 jspl3_w_asqrt32_18(.douta(w_asqrt32_18[0]),.doutb(w_asqrt32_18[1]),.doutc(w_asqrt32_18[2]),.din(w_asqrt32_5[2]));
	jspl3 jspl3_w_asqrt32_19(.douta(w_asqrt32_19[0]),.doutb(w_asqrt32_19[1]),.doutc(w_asqrt32_19[2]),.din(w_asqrt32_6[0]));
	jspl3 jspl3_w_asqrt32_20(.douta(w_asqrt32_20[0]),.doutb(w_asqrt32_20[1]),.doutc(w_asqrt32_20[2]),.din(w_asqrt32_6[1]));
	jspl3 jspl3_w_asqrt32_21(.douta(w_asqrt32_21[0]),.doutb(w_asqrt32_21[1]),.doutc(w_asqrt32_21[2]),.din(w_asqrt32_6[2]));
	jspl3 jspl3_w_asqrt32_22(.douta(w_asqrt32_22[0]),.doutb(w_asqrt32_22[1]),.doutc(w_asqrt32_22[2]),.din(w_asqrt32_7[0]));
	jspl3 jspl3_w_asqrt32_23(.douta(w_asqrt32_23[0]),.doutb(w_asqrt32_23[1]),.doutc(w_asqrt32_23[2]),.din(w_asqrt32_7[1]));
	jspl3 jspl3_w_asqrt32_24(.douta(w_asqrt32_24[0]),.doutb(w_asqrt32_24[1]),.doutc(w_asqrt32_24[2]),.din(w_asqrt32_7[2]));
	jspl3 jspl3_w_asqrt32_25(.douta(w_asqrt32_25[0]),.doutb(w_asqrt32_25[1]),.doutc(w_asqrt32_25[2]),.din(w_asqrt32_8[0]));
	jspl3 jspl3_w_asqrt32_26(.douta(w_asqrt32_26[0]),.doutb(w_asqrt32_26[1]),.doutc(w_asqrt32_26[2]),.din(w_asqrt32_8[1]));
	jspl3 jspl3_w_asqrt32_27(.douta(w_asqrt32_27[0]),.doutb(w_asqrt32_27[1]),.doutc(w_asqrt32_27[2]),.din(w_asqrt32_8[2]));
	jspl3 jspl3_w_asqrt32_28(.douta(w_asqrt32_28[0]),.doutb(w_asqrt32_28[1]),.doutc(w_asqrt32_28[2]),.din(w_asqrt32_9[0]));
	jspl3 jspl3_w_asqrt32_29(.douta(w_asqrt32_29[0]),.doutb(w_asqrt32_29[1]),.doutc(w_asqrt32_29[2]),.din(w_asqrt32_9[1]));
	jspl3 jspl3_w_asqrt32_30(.douta(w_asqrt32_30[0]),.doutb(w_asqrt32_30[1]),.doutc(w_asqrt32_30[2]),.din(w_asqrt32_9[2]));
	jspl3 jspl3_w_asqrt32_31(.douta(w_asqrt32_31[0]),.doutb(w_asqrt32_31[1]),.doutc(w_asqrt32_31[2]),.din(w_asqrt32_10[0]));
	jspl3 jspl3_w_asqrt32_32(.douta(w_asqrt32_32[0]),.doutb(w_asqrt32_32[1]),.doutc(w_asqrt32_32[2]),.din(w_asqrt32_10[1]));
	jspl3 jspl3_w_asqrt32_33(.douta(w_asqrt32_33[0]),.doutb(w_asqrt32_33[1]),.doutc(w_asqrt32_33[2]),.din(w_asqrt32_10[2]));
	jspl3 jspl3_w_asqrt32_34(.douta(w_asqrt32_34[0]),.doutb(w_asqrt32_34[1]),.doutc(w_asqrt32_34[2]),.din(w_asqrt32_11[0]));
	jspl3 jspl3_w_asqrt32_35(.douta(w_asqrt32_35[0]),.doutb(w_asqrt32_35[1]),.doutc(w_asqrt32_35[2]),.din(w_asqrt32_11[1]));
	jspl3 jspl3_w_asqrt32_36(.douta(w_asqrt32_36[0]),.doutb(w_asqrt32_36[1]),.doutc(w_asqrt32_36[2]),.din(w_asqrt32_11[2]));
	jspl3 jspl3_w_asqrt32_37(.douta(w_asqrt32_37[0]),.doutb(w_asqrt32_37[1]),.doutc(w_asqrt32_37[2]),.din(w_asqrt32_12[0]));
	jspl3 jspl3_w_asqrt32_38(.douta(w_asqrt32_38[0]),.doutb(w_asqrt32_38[1]),.doutc(asqrt[31]),.din(w_asqrt32_12[1]));
	jspl3 jspl3_w_asqrt33_0(.douta(w_asqrt33_0[0]),.doutb(w_asqrt33_0[1]),.doutc(w_asqrt33_0[2]),.din(asqrt_fa_33));
	jspl3 jspl3_w_asqrt33_1(.douta(w_asqrt33_1[0]),.doutb(w_asqrt33_1[1]),.doutc(w_asqrt33_1[2]),.din(w_asqrt33_0[0]));
	jspl3 jspl3_w_asqrt33_2(.douta(w_asqrt33_2[0]),.doutb(w_asqrt33_2[1]),.doutc(w_asqrt33_2[2]),.din(w_asqrt33_0[1]));
	jspl3 jspl3_w_asqrt33_3(.douta(w_asqrt33_3[0]),.doutb(w_asqrt33_3[1]),.doutc(w_asqrt33_3[2]),.din(w_asqrt33_0[2]));
	jspl3 jspl3_w_asqrt33_4(.douta(w_asqrt33_4[0]),.doutb(w_asqrt33_4[1]),.doutc(w_asqrt33_4[2]),.din(w_asqrt33_1[0]));
	jspl3 jspl3_w_asqrt33_5(.douta(w_asqrt33_5[0]),.doutb(w_asqrt33_5[1]),.doutc(w_asqrt33_5[2]),.din(w_asqrt33_1[1]));
	jspl3 jspl3_w_asqrt33_6(.douta(w_asqrt33_6[0]),.doutb(w_asqrt33_6[1]),.doutc(w_asqrt33_6[2]),.din(w_asqrt33_1[2]));
	jspl3 jspl3_w_asqrt33_7(.douta(w_asqrt33_7[0]),.doutb(w_asqrt33_7[1]),.doutc(w_asqrt33_7[2]),.din(w_asqrt33_2[0]));
	jspl3 jspl3_w_asqrt33_8(.douta(w_asqrt33_8[0]),.doutb(w_asqrt33_8[1]),.doutc(w_asqrt33_8[2]),.din(w_asqrt33_2[1]));
	jspl3 jspl3_w_asqrt33_9(.douta(w_asqrt33_9[0]),.doutb(w_asqrt33_9[1]),.doutc(w_asqrt33_9[2]),.din(w_asqrt33_2[2]));
	jspl3 jspl3_w_asqrt33_10(.douta(w_asqrt33_10[0]),.doutb(w_asqrt33_10[1]),.doutc(w_asqrt33_10[2]),.din(w_asqrt33_3[0]));
	jspl3 jspl3_w_asqrt33_11(.douta(w_asqrt33_11[0]),.doutb(w_asqrt33_11[1]),.doutc(w_asqrt33_11[2]),.din(w_asqrt33_3[1]));
	jspl3 jspl3_w_asqrt33_12(.douta(w_asqrt33_12[0]),.doutb(w_asqrt33_12[1]),.doutc(w_asqrt33_12[2]),.din(w_asqrt33_3[2]));
	jspl3 jspl3_w_asqrt33_13(.douta(w_asqrt33_13[0]),.doutb(w_asqrt33_13[1]),.doutc(w_asqrt33_13[2]),.din(w_asqrt33_4[0]));
	jspl3 jspl3_w_asqrt33_14(.douta(w_asqrt33_14[0]),.doutb(w_asqrt33_14[1]),.doutc(w_asqrt33_14[2]),.din(w_asqrt33_4[1]));
	jspl3 jspl3_w_asqrt33_15(.douta(w_asqrt33_15[0]),.doutb(w_asqrt33_15[1]),.doutc(w_asqrt33_15[2]),.din(w_asqrt33_4[2]));
	jspl3 jspl3_w_asqrt33_16(.douta(w_asqrt33_16[0]),.doutb(w_asqrt33_16[1]),.doutc(w_asqrt33_16[2]),.din(w_asqrt33_5[0]));
	jspl3 jspl3_w_asqrt33_17(.douta(w_asqrt33_17[0]),.doutb(w_asqrt33_17[1]),.doutc(w_asqrt33_17[2]),.din(w_asqrt33_5[1]));
	jspl3 jspl3_w_asqrt33_18(.douta(w_asqrt33_18[0]),.doutb(w_asqrt33_18[1]),.doutc(w_asqrt33_18[2]),.din(w_asqrt33_5[2]));
	jspl3 jspl3_w_asqrt33_19(.douta(w_asqrt33_19[0]),.doutb(w_asqrt33_19[1]),.doutc(w_asqrt33_19[2]),.din(w_asqrt33_6[0]));
	jspl3 jspl3_w_asqrt33_20(.douta(w_asqrt33_20[0]),.doutb(w_asqrt33_20[1]),.doutc(w_asqrt33_20[2]),.din(w_asqrt33_6[1]));
	jspl3 jspl3_w_asqrt33_21(.douta(w_asqrt33_21[0]),.doutb(w_asqrt33_21[1]),.doutc(w_asqrt33_21[2]),.din(w_asqrt33_6[2]));
	jspl3 jspl3_w_asqrt33_22(.douta(w_asqrt33_22[0]),.doutb(w_asqrt33_22[1]),.doutc(w_asqrt33_22[2]),.din(w_asqrt33_7[0]));
	jspl3 jspl3_w_asqrt33_23(.douta(w_asqrt33_23[0]),.doutb(w_asqrt33_23[1]),.doutc(w_asqrt33_23[2]),.din(w_asqrt33_7[1]));
	jspl3 jspl3_w_asqrt33_24(.douta(w_asqrt33_24[0]),.doutb(w_asqrt33_24[1]),.doutc(w_asqrt33_24[2]),.din(w_asqrt33_7[2]));
	jspl jspl_w_asqrt33_25(.douta(w_asqrt33_25),.doutb(asqrt[32]),.din(w_asqrt33_8[0]));
	jspl3 jspl3_w_asqrt34_0(.douta(w_asqrt34_0[0]),.doutb(w_asqrt34_0[1]),.doutc(w_asqrt34_0[2]),.din(asqrt_fa_34));
	jspl3 jspl3_w_asqrt34_1(.douta(w_asqrt34_1[0]),.doutb(w_asqrt34_1[1]),.doutc(w_asqrt34_1[2]),.din(w_asqrt34_0[0]));
	jspl3 jspl3_w_asqrt34_2(.douta(w_asqrt34_2[0]),.doutb(w_asqrt34_2[1]),.doutc(w_asqrt34_2[2]),.din(w_asqrt34_0[1]));
	jspl3 jspl3_w_asqrt34_3(.douta(w_asqrt34_3[0]),.doutb(w_asqrt34_3[1]),.doutc(w_asqrt34_3[2]),.din(w_asqrt34_0[2]));
	jspl3 jspl3_w_asqrt34_4(.douta(w_asqrt34_4[0]),.doutb(w_asqrt34_4[1]),.doutc(w_asqrt34_4[2]),.din(w_asqrt34_1[0]));
	jspl3 jspl3_w_asqrt34_5(.douta(w_asqrt34_5[0]),.doutb(w_asqrt34_5[1]),.doutc(w_asqrt34_5[2]),.din(w_asqrt34_1[1]));
	jspl3 jspl3_w_asqrt34_6(.douta(w_asqrt34_6[0]),.doutb(w_asqrt34_6[1]),.doutc(w_asqrt34_6[2]),.din(w_asqrt34_1[2]));
	jspl3 jspl3_w_asqrt34_7(.douta(w_asqrt34_7[0]),.doutb(w_asqrt34_7[1]),.doutc(w_asqrt34_7[2]),.din(w_asqrt34_2[0]));
	jspl3 jspl3_w_asqrt34_8(.douta(w_asqrt34_8[0]),.doutb(w_asqrt34_8[1]),.doutc(w_asqrt34_8[2]),.din(w_asqrt34_2[1]));
	jspl3 jspl3_w_asqrt34_9(.douta(w_asqrt34_9[0]),.doutb(w_asqrt34_9[1]),.doutc(w_asqrt34_9[2]),.din(w_asqrt34_2[2]));
	jspl3 jspl3_w_asqrt34_10(.douta(w_asqrt34_10[0]),.doutb(w_asqrt34_10[1]),.doutc(w_asqrt34_10[2]),.din(w_asqrt34_3[0]));
	jspl3 jspl3_w_asqrt34_11(.douta(w_asqrt34_11[0]),.doutb(w_asqrt34_11[1]),.doutc(w_asqrt34_11[2]),.din(w_asqrt34_3[1]));
	jspl3 jspl3_w_asqrt34_12(.douta(w_asqrt34_12[0]),.doutb(w_asqrt34_12[1]),.doutc(w_asqrt34_12[2]),.din(w_asqrt34_3[2]));
	jspl3 jspl3_w_asqrt34_13(.douta(w_asqrt34_13[0]),.doutb(w_asqrt34_13[1]),.doutc(w_asqrt34_13[2]),.din(w_asqrt34_4[0]));
	jspl3 jspl3_w_asqrt34_14(.douta(w_asqrt34_14[0]),.doutb(w_asqrt34_14[1]),.doutc(w_asqrt34_14[2]),.din(w_asqrt34_4[1]));
	jspl3 jspl3_w_asqrt34_15(.douta(w_asqrt34_15[0]),.doutb(w_asqrt34_15[1]),.doutc(w_asqrt34_15[2]),.din(w_asqrt34_4[2]));
	jspl3 jspl3_w_asqrt34_16(.douta(w_asqrt34_16[0]),.doutb(w_asqrt34_16[1]),.doutc(w_asqrt34_16[2]),.din(w_asqrt34_5[0]));
	jspl3 jspl3_w_asqrt34_17(.douta(w_asqrt34_17[0]),.doutb(w_asqrt34_17[1]),.doutc(w_asqrt34_17[2]),.din(w_asqrt34_5[1]));
	jspl3 jspl3_w_asqrt34_18(.douta(w_asqrt34_18[0]),.doutb(w_asqrt34_18[1]),.doutc(w_asqrt34_18[2]),.din(w_asqrt34_5[2]));
	jspl3 jspl3_w_asqrt34_19(.douta(w_asqrt34_19[0]),.doutb(w_asqrt34_19[1]),.doutc(w_asqrt34_19[2]),.din(w_asqrt34_6[0]));
	jspl3 jspl3_w_asqrt34_20(.douta(w_asqrt34_20[0]),.doutb(w_asqrt34_20[1]),.doutc(w_asqrt34_20[2]),.din(w_asqrt34_6[1]));
	jspl3 jspl3_w_asqrt34_21(.douta(w_asqrt34_21[0]),.doutb(w_asqrt34_21[1]),.doutc(w_asqrt34_21[2]),.din(w_asqrt34_6[2]));
	jspl3 jspl3_w_asqrt34_22(.douta(w_asqrt34_22[0]),.doutb(w_asqrt34_22[1]),.doutc(w_asqrt34_22[2]),.din(w_asqrt34_7[0]));
	jspl3 jspl3_w_asqrt34_23(.douta(w_asqrt34_23[0]),.doutb(w_asqrt34_23[1]),.doutc(w_asqrt34_23[2]),.din(w_asqrt34_7[1]));
	jspl3 jspl3_w_asqrt34_24(.douta(w_asqrt34_24[0]),.doutb(w_asqrt34_24[1]),.doutc(w_asqrt34_24[2]),.din(w_asqrt34_7[2]));
	jspl3 jspl3_w_asqrt34_25(.douta(w_asqrt34_25[0]),.doutb(w_asqrt34_25[1]),.doutc(w_asqrt34_25[2]),.din(w_asqrt34_8[0]));
	jspl3 jspl3_w_asqrt34_26(.douta(w_asqrt34_26[0]),.doutb(w_asqrt34_26[1]),.doutc(w_asqrt34_26[2]),.din(w_asqrt34_8[1]));
	jspl3 jspl3_w_asqrt34_27(.douta(w_asqrt34_27[0]),.doutb(w_asqrt34_27[1]),.doutc(w_asqrt34_27[2]),.din(w_asqrt34_8[2]));
	jspl3 jspl3_w_asqrt34_28(.douta(w_asqrt34_28[0]),.doutb(w_asqrt34_28[1]),.doutc(w_asqrt34_28[2]),.din(w_asqrt34_9[0]));
	jspl3 jspl3_w_asqrt34_29(.douta(w_asqrt34_29[0]),.doutb(w_asqrt34_29[1]),.doutc(w_asqrt34_29[2]),.din(w_asqrt34_9[1]));
	jspl3 jspl3_w_asqrt34_30(.douta(w_asqrt34_30[0]),.doutb(w_asqrt34_30[1]),.doutc(w_asqrt34_30[2]),.din(w_asqrt34_9[2]));
	jspl3 jspl3_w_asqrt34_31(.douta(w_asqrt34_31[0]),.doutb(w_asqrt34_31[1]),.doutc(w_asqrt34_31[2]),.din(w_asqrt34_10[0]));
	jspl3 jspl3_w_asqrt34_32(.douta(w_asqrt34_32[0]),.doutb(w_asqrt34_32[1]),.doutc(w_asqrt34_32[2]),.din(w_asqrt34_10[1]));
	jspl3 jspl3_w_asqrt34_33(.douta(w_asqrt34_33[0]),.doutb(w_asqrt34_33[1]),.doutc(w_asqrt34_33[2]),.din(w_asqrt34_10[2]));
	jspl3 jspl3_w_asqrt34_34(.douta(w_asqrt34_34[0]),.doutb(w_asqrt34_34[1]),.doutc(w_asqrt34_34[2]),.din(w_asqrt34_11[0]));
	jspl3 jspl3_w_asqrt34_35(.douta(w_asqrt34_35[0]),.doutb(w_asqrt34_35[1]),.doutc(w_asqrt34_35[2]),.din(w_asqrt34_11[1]));
	jspl3 jspl3_w_asqrt34_36(.douta(w_asqrt34_36[0]),.doutb(w_asqrt34_36[1]),.doutc(w_asqrt34_36[2]),.din(w_asqrt34_11[2]));
	jspl3 jspl3_w_asqrt34_37(.douta(w_asqrt34_37[0]),.doutb(w_asqrt34_37[1]),.doutc(w_asqrt34_37[2]),.din(w_asqrt34_12[0]));
	jspl3 jspl3_w_asqrt34_38(.douta(w_asqrt34_38[0]),.doutb(w_asqrt34_38[1]),.doutc(w_asqrt34_38[2]),.din(w_asqrt34_12[1]));
	jspl jspl_w_asqrt34_39(.douta(w_asqrt34_39),.doutb(asqrt[33]),.din(w_asqrt34_12[2]));
	jspl3 jspl3_w_asqrt35_0(.douta(w_asqrt35_0[0]),.doutb(w_asqrt35_0[1]),.doutc(w_asqrt35_0[2]),.din(asqrt_fa_35));
	jspl3 jspl3_w_asqrt35_1(.douta(w_asqrt35_1[0]),.doutb(w_asqrt35_1[1]),.doutc(w_asqrt35_1[2]),.din(w_asqrt35_0[0]));
	jspl3 jspl3_w_asqrt35_2(.douta(w_asqrt35_2[0]),.doutb(w_asqrt35_2[1]),.doutc(w_asqrt35_2[2]),.din(w_asqrt35_0[1]));
	jspl3 jspl3_w_asqrt35_3(.douta(w_asqrt35_3[0]),.doutb(w_asqrt35_3[1]),.doutc(w_asqrt35_3[2]),.din(w_asqrt35_0[2]));
	jspl3 jspl3_w_asqrt35_4(.douta(w_asqrt35_4[0]),.doutb(w_asqrt35_4[1]),.doutc(w_asqrt35_4[2]),.din(w_asqrt35_1[0]));
	jspl3 jspl3_w_asqrt35_5(.douta(w_asqrt35_5[0]),.doutb(w_asqrt35_5[1]),.doutc(w_asqrt35_5[2]),.din(w_asqrt35_1[1]));
	jspl3 jspl3_w_asqrt35_6(.douta(w_asqrt35_6[0]),.doutb(w_asqrt35_6[1]),.doutc(w_asqrt35_6[2]),.din(w_asqrt35_1[2]));
	jspl3 jspl3_w_asqrt35_7(.douta(w_asqrt35_7[0]),.doutb(w_asqrt35_7[1]),.doutc(w_asqrt35_7[2]),.din(w_asqrt35_2[0]));
	jspl3 jspl3_w_asqrt35_8(.douta(w_asqrt35_8[0]),.doutb(w_asqrt35_8[1]),.doutc(w_asqrt35_8[2]),.din(w_asqrt35_2[1]));
	jspl3 jspl3_w_asqrt35_9(.douta(w_asqrt35_9[0]),.doutb(w_asqrt35_9[1]),.doutc(w_asqrt35_9[2]),.din(w_asqrt35_2[2]));
	jspl3 jspl3_w_asqrt35_10(.douta(w_asqrt35_10[0]),.doutb(w_asqrt35_10[1]),.doutc(w_asqrt35_10[2]),.din(w_asqrt35_3[0]));
	jspl3 jspl3_w_asqrt35_11(.douta(w_asqrt35_11[0]),.doutb(w_asqrt35_11[1]),.doutc(w_asqrt35_11[2]),.din(w_asqrt35_3[1]));
	jspl3 jspl3_w_asqrt35_12(.douta(w_asqrt35_12[0]),.doutb(w_asqrt35_12[1]),.doutc(w_asqrt35_12[2]),.din(w_asqrt35_3[2]));
	jspl3 jspl3_w_asqrt35_13(.douta(w_asqrt35_13[0]),.doutb(w_asqrt35_13[1]),.doutc(w_asqrt35_13[2]),.din(w_asqrt35_4[0]));
	jspl3 jspl3_w_asqrt35_14(.douta(w_asqrt35_14[0]),.doutb(w_asqrt35_14[1]),.doutc(w_asqrt35_14[2]),.din(w_asqrt35_4[1]));
	jspl3 jspl3_w_asqrt35_15(.douta(w_asqrt35_15[0]),.doutb(w_asqrt35_15[1]),.doutc(w_asqrt35_15[2]),.din(w_asqrt35_4[2]));
	jspl3 jspl3_w_asqrt35_16(.douta(w_asqrt35_16[0]),.doutb(w_asqrt35_16[1]),.doutc(w_asqrt35_16[2]),.din(w_asqrt35_5[0]));
	jspl3 jspl3_w_asqrt35_17(.douta(w_asqrt35_17[0]),.doutb(w_asqrt35_17[1]),.doutc(w_asqrt35_17[2]),.din(w_asqrt35_5[1]));
	jspl3 jspl3_w_asqrt35_18(.douta(w_asqrt35_18[0]),.doutb(w_asqrt35_18[1]),.doutc(w_asqrt35_18[2]),.din(w_asqrt35_5[2]));
	jspl3 jspl3_w_asqrt35_19(.douta(w_asqrt35_19[0]),.doutb(w_asqrt35_19[1]),.doutc(w_asqrt35_19[2]),.din(w_asqrt35_6[0]));
	jspl3 jspl3_w_asqrt35_20(.douta(w_asqrt35_20[0]),.doutb(w_asqrt35_20[1]),.doutc(w_asqrt35_20[2]),.din(w_asqrt35_6[1]));
	jspl3 jspl3_w_asqrt35_21(.douta(w_asqrt35_21[0]),.doutb(w_asqrt35_21[1]),.doutc(w_asqrt35_21[2]),.din(w_asqrt35_6[2]));
	jspl3 jspl3_w_asqrt35_22(.douta(w_asqrt35_22[0]),.doutb(w_asqrt35_22[1]),.doutc(w_asqrt35_22[2]),.din(w_asqrt35_7[0]));
	jspl3 jspl3_w_asqrt35_23(.douta(w_asqrt35_23[0]),.doutb(w_asqrt35_23[1]),.doutc(w_asqrt35_23[2]),.din(w_asqrt35_7[1]));
	jspl3 jspl3_w_asqrt35_24(.douta(w_asqrt35_24[0]),.doutb(w_asqrt35_24[1]),.doutc(w_asqrt35_24[2]),.din(w_asqrt35_7[2]));
	jspl3 jspl3_w_asqrt35_25(.douta(w_asqrt35_25[0]),.doutb(w_asqrt35_25[1]),.doutc(w_asqrt35_25[2]),.din(w_asqrt35_8[0]));
	jspl3 jspl3_w_asqrt35_26(.douta(w_asqrt35_26[0]),.doutb(w_asqrt35_26[1]),.doutc(w_asqrt35_26[2]),.din(w_asqrt35_8[1]));
	jspl jspl_w_asqrt35_27(.douta(w_asqrt35_27),.doutb(asqrt[34]),.din(w_asqrt35_8[2]));
	jspl3 jspl3_w_asqrt36_0(.douta(w_asqrt36_0[0]),.doutb(w_asqrt36_0[1]),.doutc(w_asqrt36_0[2]),.din(asqrt_fa_36));
	jspl3 jspl3_w_asqrt36_1(.douta(w_asqrt36_1[0]),.doutb(w_asqrt36_1[1]),.doutc(w_asqrt36_1[2]),.din(w_asqrt36_0[0]));
	jspl3 jspl3_w_asqrt36_2(.douta(w_asqrt36_2[0]),.doutb(w_asqrt36_2[1]),.doutc(w_asqrt36_2[2]),.din(w_asqrt36_0[1]));
	jspl3 jspl3_w_asqrt36_3(.douta(w_asqrt36_3[0]),.doutb(w_asqrt36_3[1]),.doutc(w_asqrt36_3[2]),.din(w_asqrt36_0[2]));
	jspl3 jspl3_w_asqrt36_4(.douta(w_asqrt36_4[0]),.doutb(w_asqrt36_4[1]),.doutc(w_asqrt36_4[2]),.din(w_asqrt36_1[0]));
	jspl3 jspl3_w_asqrt36_5(.douta(w_asqrt36_5[0]),.doutb(w_asqrt36_5[1]),.doutc(w_asqrt36_5[2]),.din(w_asqrt36_1[1]));
	jspl3 jspl3_w_asqrt36_6(.douta(w_asqrt36_6[0]),.doutb(w_asqrt36_6[1]),.doutc(w_asqrt36_6[2]),.din(w_asqrt36_1[2]));
	jspl3 jspl3_w_asqrt36_7(.douta(w_asqrt36_7[0]),.doutb(w_asqrt36_7[1]),.doutc(w_asqrt36_7[2]),.din(w_asqrt36_2[0]));
	jspl3 jspl3_w_asqrt36_8(.douta(w_asqrt36_8[0]),.doutb(w_asqrt36_8[1]),.doutc(w_asqrt36_8[2]),.din(w_asqrt36_2[1]));
	jspl3 jspl3_w_asqrt36_9(.douta(w_asqrt36_9[0]),.doutb(w_asqrt36_9[1]),.doutc(w_asqrt36_9[2]),.din(w_asqrt36_2[2]));
	jspl3 jspl3_w_asqrt36_10(.douta(w_asqrt36_10[0]),.doutb(w_asqrt36_10[1]),.doutc(w_asqrt36_10[2]),.din(w_asqrt36_3[0]));
	jspl3 jspl3_w_asqrt36_11(.douta(w_asqrt36_11[0]),.doutb(w_asqrt36_11[1]),.doutc(w_asqrt36_11[2]),.din(w_asqrt36_3[1]));
	jspl3 jspl3_w_asqrt36_12(.douta(w_asqrt36_12[0]),.doutb(w_asqrt36_12[1]),.doutc(w_asqrt36_12[2]),.din(w_asqrt36_3[2]));
	jspl3 jspl3_w_asqrt36_13(.douta(w_asqrt36_13[0]),.doutb(w_asqrt36_13[1]),.doutc(w_asqrt36_13[2]),.din(w_asqrt36_4[0]));
	jspl3 jspl3_w_asqrt36_14(.douta(w_asqrt36_14[0]),.doutb(w_asqrt36_14[1]),.doutc(w_asqrt36_14[2]),.din(w_asqrt36_4[1]));
	jspl3 jspl3_w_asqrt36_15(.douta(w_asqrt36_15[0]),.doutb(w_asqrt36_15[1]),.doutc(w_asqrt36_15[2]),.din(w_asqrt36_4[2]));
	jspl3 jspl3_w_asqrt36_16(.douta(w_asqrt36_16[0]),.doutb(w_asqrt36_16[1]),.doutc(w_asqrt36_16[2]),.din(w_asqrt36_5[0]));
	jspl3 jspl3_w_asqrt36_17(.douta(w_asqrt36_17[0]),.doutb(w_asqrt36_17[1]),.doutc(w_asqrt36_17[2]),.din(w_asqrt36_5[1]));
	jspl3 jspl3_w_asqrt36_18(.douta(w_asqrt36_18[0]),.doutb(w_asqrt36_18[1]),.doutc(w_asqrt36_18[2]),.din(w_asqrt36_5[2]));
	jspl3 jspl3_w_asqrt36_19(.douta(w_asqrt36_19[0]),.doutb(w_asqrt36_19[1]),.doutc(w_asqrt36_19[2]),.din(w_asqrt36_6[0]));
	jspl3 jspl3_w_asqrt36_20(.douta(w_asqrt36_20[0]),.doutb(w_asqrt36_20[1]),.doutc(w_asqrt36_20[2]),.din(w_asqrt36_6[1]));
	jspl3 jspl3_w_asqrt36_21(.douta(w_asqrt36_21[0]),.doutb(w_asqrt36_21[1]),.doutc(w_asqrt36_21[2]),.din(w_asqrt36_6[2]));
	jspl3 jspl3_w_asqrt36_22(.douta(w_asqrt36_22[0]),.doutb(w_asqrt36_22[1]),.doutc(w_asqrt36_22[2]),.din(w_asqrt36_7[0]));
	jspl3 jspl3_w_asqrt36_23(.douta(w_asqrt36_23[0]),.doutb(w_asqrt36_23[1]),.doutc(w_asqrt36_23[2]),.din(w_asqrt36_7[1]));
	jspl3 jspl3_w_asqrt36_24(.douta(w_asqrt36_24[0]),.doutb(w_asqrt36_24[1]),.doutc(w_asqrt36_24[2]),.din(w_asqrt36_7[2]));
	jspl3 jspl3_w_asqrt36_25(.douta(w_asqrt36_25[0]),.doutb(w_asqrt36_25[1]),.doutc(w_asqrt36_25[2]),.din(w_asqrt36_8[0]));
	jspl3 jspl3_w_asqrt36_26(.douta(w_asqrt36_26[0]),.doutb(w_asqrt36_26[1]),.doutc(w_asqrt36_26[2]),.din(w_asqrt36_8[1]));
	jspl3 jspl3_w_asqrt36_27(.douta(w_asqrt36_27[0]),.doutb(w_asqrt36_27[1]),.doutc(w_asqrt36_27[2]),.din(w_asqrt36_8[2]));
	jspl3 jspl3_w_asqrt36_28(.douta(w_asqrt36_28[0]),.doutb(w_asqrt36_28[1]),.doutc(w_asqrt36_28[2]),.din(w_asqrt36_9[0]));
	jspl3 jspl3_w_asqrt36_29(.douta(w_asqrt36_29[0]),.doutb(w_asqrt36_29[1]),.doutc(w_asqrt36_29[2]),.din(w_asqrt36_9[1]));
	jspl3 jspl3_w_asqrt36_30(.douta(w_asqrt36_30[0]),.doutb(w_asqrt36_30[1]),.doutc(w_asqrt36_30[2]),.din(w_asqrt36_9[2]));
	jspl3 jspl3_w_asqrt36_31(.douta(w_asqrt36_31[0]),.doutb(w_asqrt36_31[1]),.doutc(w_asqrt36_31[2]),.din(w_asqrt36_10[0]));
	jspl3 jspl3_w_asqrt36_32(.douta(w_asqrt36_32[0]),.doutb(w_asqrt36_32[1]),.doutc(w_asqrt36_32[2]),.din(w_asqrt36_10[1]));
	jspl3 jspl3_w_asqrt36_33(.douta(w_asqrt36_33[0]),.doutb(w_asqrt36_33[1]),.doutc(w_asqrt36_33[2]),.din(w_asqrt36_10[2]));
	jspl3 jspl3_w_asqrt36_34(.douta(w_asqrt36_34[0]),.doutb(w_asqrt36_34[1]),.doutc(w_asqrt36_34[2]),.din(w_asqrt36_11[0]));
	jspl3 jspl3_w_asqrt36_35(.douta(w_asqrt36_35[0]),.doutb(w_asqrt36_35[1]),.doutc(w_asqrt36_35[2]),.din(w_asqrt36_11[1]));
	jspl3 jspl3_w_asqrt36_36(.douta(w_asqrt36_36[0]),.doutb(w_asqrt36_36[1]),.doutc(w_asqrt36_36[2]),.din(w_asqrt36_11[2]));
	jspl3 jspl3_w_asqrt36_37(.douta(w_asqrt36_37[0]),.doutb(w_asqrt36_37[1]),.doutc(w_asqrt36_37[2]),.din(w_asqrt36_12[0]));
	jspl3 jspl3_w_asqrt36_38(.douta(w_asqrt36_38[0]),.doutb(w_asqrt36_38[1]),.doutc(w_asqrt36_38[2]),.din(w_asqrt36_12[1]));
	jspl jspl_w_asqrt36_39(.douta(w_asqrt36_39),.doutb(asqrt[35]),.din(w_asqrt36_12[2]));
	jspl3 jspl3_w_asqrt37_0(.douta(w_asqrt37_0[0]),.doutb(w_asqrt37_0[1]),.doutc(w_asqrt37_0[2]),.din(asqrt_fa_37));
	jspl3 jspl3_w_asqrt37_1(.douta(w_asqrt37_1[0]),.doutb(w_asqrt37_1[1]),.doutc(w_asqrt37_1[2]),.din(w_asqrt37_0[0]));
	jspl3 jspl3_w_asqrt37_2(.douta(w_asqrt37_2[0]),.doutb(w_asqrt37_2[1]),.doutc(w_asqrt37_2[2]),.din(w_asqrt37_0[1]));
	jspl3 jspl3_w_asqrt37_3(.douta(w_asqrt37_3[0]),.doutb(w_asqrt37_3[1]),.doutc(w_asqrt37_3[2]),.din(w_asqrt37_0[2]));
	jspl3 jspl3_w_asqrt37_4(.douta(w_asqrt37_4[0]),.doutb(w_asqrt37_4[1]),.doutc(w_asqrt37_4[2]),.din(w_asqrt37_1[0]));
	jspl3 jspl3_w_asqrt37_5(.douta(w_asqrt37_5[0]),.doutb(w_asqrt37_5[1]),.doutc(w_asqrt37_5[2]),.din(w_asqrt37_1[1]));
	jspl3 jspl3_w_asqrt37_6(.douta(w_asqrt37_6[0]),.doutb(w_asqrt37_6[1]),.doutc(w_asqrt37_6[2]),.din(w_asqrt37_1[2]));
	jspl3 jspl3_w_asqrt37_7(.douta(w_asqrt37_7[0]),.doutb(w_asqrt37_7[1]),.doutc(w_asqrt37_7[2]),.din(w_asqrt37_2[0]));
	jspl3 jspl3_w_asqrt37_8(.douta(w_asqrt37_8[0]),.doutb(w_asqrt37_8[1]),.doutc(w_asqrt37_8[2]),.din(w_asqrt37_2[1]));
	jspl3 jspl3_w_asqrt37_9(.douta(w_asqrt37_9[0]),.doutb(w_asqrt37_9[1]),.doutc(w_asqrt37_9[2]),.din(w_asqrt37_2[2]));
	jspl3 jspl3_w_asqrt37_10(.douta(w_asqrt37_10[0]),.doutb(w_asqrt37_10[1]),.doutc(w_asqrt37_10[2]),.din(w_asqrt37_3[0]));
	jspl3 jspl3_w_asqrt37_11(.douta(w_asqrt37_11[0]),.doutb(w_asqrt37_11[1]),.doutc(w_asqrt37_11[2]),.din(w_asqrt37_3[1]));
	jspl3 jspl3_w_asqrt37_12(.douta(w_asqrt37_12[0]),.doutb(w_asqrt37_12[1]),.doutc(w_asqrt37_12[2]),.din(w_asqrt37_3[2]));
	jspl3 jspl3_w_asqrt37_13(.douta(w_asqrt37_13[0]),.doutb(w_asqrt37_13[1]),.doutc(w_asqrt37_13[2]),.din(w_asqrt37_4[0]));
	jspl3 jspl3_w_asqrt37_14(.douta(w_asqrt37_14[0]),.doutb(w_asqrt37_14[1]),.doutc(w_asqrt37_14[2]),.din(w_asqrt37_4[1]));
	jspl3 jspl3_w_asqrt37_15(.douta(w_asqrt37_15[0]),.doutb(w_asqrt37_15[1]),.doutc(w_asqrt37_15[2]),.din(w_asqrt37_4[2]));
	jspl3 jspl3_w_asqrt37_16(.douta(w_asqrt37_16[0]),.doutb(w_asqrt37_16[1]),.doutc(w_asqrt37_16[2]),.din(w_asqrt37_5[0]));
	jspl3 jspl3_w_asqrt37_17(.douta(w_asqrt37_17[0]),.doutb(w_asqrt37_17[1]),.doutc(w_asqrt37_17[2]),.din(w_asqrt37_5[1]));
	jspl3 jspl3_w_asqrt37_18(.douta(w_asqrt37_18[0]),.doutb(w_asqrt37_18[1]),.doutc(w_asqrt37_18[2]),.din(w_asqrt37_5[2]));
	jspl3 jspl3_w_asqrt37_19(.douta(w_asqrt37_19[0]),.doutb(w_asqrt37_19[1]),.doutc(w_asqrt37_19[2]),.din(w_asqrt37_6[0]));
	jspl3 jspl3_w_asqrt37_20(.douta(w_asqrt37_20[0]),.doutb(w_asqrt37_20[1]),.doutc(w_asqrt37_20[2]),.din(w_asqrt37_6[1]));
	jspl3 jspl3_w_asqrt37_21(.douta(w_asqrt37_21[0]),.doutb(w_asqrt37_21[1]),.doutc(w_asqrt37_21[2]),.din(w_asqrt37_6[2]));
	jspl3 jspl3_w_asqrt37_22(.douta(w_asqrt37_22[0]),.doutb(w_asqrt37_22[1]),.doutc(w_asqrt37_22[2]),.din(w_asqrt37_7[0]));
	jspl3 jspl3_w_asqrt37_23(.douta(w_asqrt37_23[0]),.doutb(w_asqrt37_23[1]),.doutc(w_asqrt37_23[2]),.din(w_asqrt37_7[1]));
	jspl3 jspl3_w_asqrt37_24(.douta(w_asqrt37_24[0]),.doutb(w_asqrt37_24[1]),.doutc(w_asqrt37_24[2]),.din(w_asqrt37_7[2]));
	jspl3 jspl3_w_asqrt37_25(.douta(w_asqrt37_25[0]),.doutb(w_asqrt37_25[1]),.doutc(w_asqrt37_25[2]),.din(w_asqrt37_8[0]));
	jspl3 jspl3_w_asqrt37_26(.douta(w_asqrt37_26[0]),.doutb(w_asqrt37_26[1]),.doutc(w_asqrt37_26[2]),.din(w_asqrt37_8[1]));
	jspl3 jspl3_w_asqrt37_27(.douta(w_asqrt37_27[0]),.doutb(w_asqrt37_27[1]),.doutc(w_asqrt37_27[2]),.din(w_asqrt37_8[2]));
	jspl jspl_w_asqrt37_28(.douta(w_asqrt37_28),.doutb(asqrt[36]),.din(w_asqrt37_9[0]));
	jspl3 jspl3_w_asqrt38_0(.douta(w_asqrt38_0[0]),.doutb(w_asqrt38_0[1]),.doutc(w_asqrt38_0[2]),.din(asqrt_fa_38));
	jspl3 jspl3_w_asqrt38_1(.douta(w_asqrt38_1[0]),.doutb(w_asqrt38_1[1]),.doutc(w_asqrt38_1[2]),.din(w_asqrt38_0[0]));
	jspl3 jspl3_w_asqrt38_2(.douta(w_asqrt38_2[0]),.doutb(w_asqrt38_2[1]),.doutc(w_asqrt38_2[2]),.din(w_asqrt38_0[1]));
	jspl3 jspl3_w_asqrt38_3(.douta(w_asqrt38_3[0]),.doutb(w_asqrt38_3[1]),.doutc(w_asqrt38_3[2]),.din(w_asqrt38_0[2]));
	jspl3 jspl3_w_asqrt38_4(.douta(w_asqrt38_4[0]),.doutb(w_asqrt38_4[1]),.doutc(w_asqrt38_4[2]),.din(w_asqrt38_1[0]));
	jspl3 jspl3_w_asqrt38_5(.douta(w_asqrt38_5[0]),.doutb(w_asqrt38_5[1]),.doutc(w_asqrt38_5[2]),.din(w_asqrt38_1[1]));
	jspl3 jspl3_w_asqrt38_6(.douta(w_asqrt38_6[0]),.doutb(w_asqrt38_6[1]),.doutc(w_asqrt38_6[2]),.din(w_asqrt38_1[2]));
	jspl3 jspl3_w_asqrt38_7(.douta(w_asqrt38_7[0]),.doutb(w_asqrt38_7[1]),.doutc(w_asqrt38_7[2]),.din(w_asqrt38_2[0]));
	jspl3 jspl3_w_asqrt38_8(.douta(w_asqrt38_8[0]),.doutb(w_asqrt38_8[1]),.doutc(w_asqrt38_8[2]),.din(w_asqrt38_2[1]));
	jspl3 jspl3_w_asqrt38_9(.douta(w_asqrt38_9[0]),.doutb(w_asqrt38_9[1]),.doutc(w_asqrt38_9[2]),.din(w_asqrt38_2[2]));
	jspl3 jspl3_w_asqrt38_10(.douta(w_asqrt38_10[0]),.doutb(w_asqrt38_10[1]),.doutc(w_asqrt38_10[2]),.din(w_asqrt38_3[0]));
	jspl3 jspl3_w_asqrt38_11(.douta(w_asqrt38_11[0]),.doutb(w_asqrt38_11[1]),.doutc(w_asqrt38_11[2]),.din(w_asqrt38_3[1]));
	jspl3 jspl3_w_asqrt38_12(.douta(w_asqrt38_12[0]),.doutb(w_asqrt38_12[1]),.doutc(w_asqrt38_12[2]),.din(w_asqrt38_3[2]));
	jspl3 jspl3_w_asqrt38_13(.douta(w_asqrt38_13[0]),.doutb(w_asqrt38_13[1]),.doutc(w_asqrt38_13[2]),.din(w_asqrt38_4[0]));
	jspl3 jspl3_w_asqrt38_14(.douta(w_asqrt38_14[0]),.doutb(w_asqrt38_14[1]),.doutc(w_asqrt38_14[2]),.din(w_asqrt38_4[1]));
	jspl3 jspl3_w_asqrt38_15(.douta(w_asqrt38_15[0]),.doutb(w_asqrt38_15[1]),.doutc(w_asqrt38_15[2]),.din(w_asqrt38_4[2]));
	jspl3 jspl3_w_asqrt38_16(.douta(w_asqrt38_16[0]),.doutb(w_asqrt38_16[1]),.doutc(w_asqrt38_16[2]),.din(w_asqrt38_5[0]));
	jspl3 jspl3_w_asqrt38_17(.douta(w_asqrt38_17[0]),.doutb(w_asqrt38_17[1]),.doutc(w_asqrt38_17[2]),.din(w_asqrt38_5[1]));
	jspl3 jspl3_w_asqrt38_18(.douta(w_asqrt38_18[0]),.doutb(w_asqrt38_18[1]),.doutc(w_asqrt38_18[2]),.din(w_asqrt38_5[2]));
	jspl3 jspl3_w_asqrt38_19(.douta(w_asqrt38_19[0]),.doutb(w_asqrt38_19[1]),.doutc(w_asqrt38_19[2]),.din(w_asqrt38_6[0]));
	jspl3 jspl3_w_asqrt38_20(.douta(w_asqrt38_20[0]),.doutb(w_asqrt38_20[1]),.doutc(w_asqrt38_20[2]),.din(w_asqrt38_6[1]));
	jspl3 jspl3_w_asqrt38_21(.douta(w_asqrt38_21[0]),.doutb(w_asqrt38_21[1]),.doutc(w_asqrt38_21[2]),.din(w_asqrt38_6[2]));
	jspl3 jspl3_w_asqrt38_22(.douta(w_asqrt38_22[0]),.doutb(w_asqrt38_22[1]),.doutc(w_asqrt38_22[2]),.din(w_asqrt38_7[0]));
	jspl3 jspl3_w_asqrt38_23(.douta(w_asqrt38_23[0]),.doutb(w_asqrt38_23[1]),.doutc(w_asqrt38_23[2]),.din(w_asqrt38_7[1]));
	jspl3 jspl3_w_asqrt38_24(.douta(w_asqrt38_24[0]),.doutb(w_asqrt38_24[1]),.doutc(w_asqrt38_24[2]),.din(w_asqrt38_7[2]));
	jspl3 jspl3_w_asqrt38_25(.douta(w_asqrt38_25[0]),.doutb(w_asqrt38_25[1]),.doutc(w_asqrt38_25[2]),.din(w_asqrt38_8[0]));
	jspl3 jspl3_w_asqrt38_26(.douta(w_asqrt38_26[0]),.doutb(w_asqrt38_26[1]),.doutc(w_asqrt38_26[2]),.din(w_asqrt38_8[1]));
	jspl3 jspl3_w_asqrt38_27(.douta(w_asqrt38_27[0]),.doutb(w_asqrt38_27[1]),.doutc(w_asqrt38_27[2]),.din(w_asqrt38_8[2]));
	jspl3 jspl3_w_asqrt38_28(.douta(w_asqrt38_28[0]),.doutb(w_asqrt38_28[1]),.doutc(w_asqrt38_28[2]),.din(w_asqrt38_9[0]));
	jspl3 jspl3_w_asqrt38_29(.douta(w_asqrt38_29[0]),.doutb(w_asqrt38_29[1]),.doutc(w_asqrt38_29[2]),.din(w_asqrt38_9[1]));
	jspl3 jspl3_w_asqrt38_30(.douta(w_asqrt38_30[0]),.doutb(w_asqrt38_30[1]),.doutc(w_asqrt38_30[2]),.din(w_asqrt38_9[2]));
	jspl3 jspl3_w_asqrt38_31(.douta(w_asqrt38_31[0]),.doutb(w_asqrt38_31[1]),.doutc(w_asqrt38_31[2]),.din(w_asqrt38_10[0]));
	jspl3 jspl3_w_asqrt38_32(.douta(w_asqrt38_32[0]),.doutb(w_asqrt38_32[1]),.doutc(w_asqrt38_32[2]),.din(w_asqrt38_10[1]));
	jspl3 jspl3_w_asqrt38_33(.douta(w_asqrt38_33[0]),.doutb(w_asqrt38_33[1]),.doutc(w_asqrt38_33[2]),.din(w_asqrt38_10[2]));
	jspl3 jspl3_w_asqrt38_34(.douta(w_asqrt38_34[0]),.doutb(w_asqrt38_34[1]),.doutc(w_asqrt38_34[2]),.din(w_asqrt38_11[0]));
	jspl3 jspl3_w_asqrt38_35(.douta(w_asqrt38_35[0]),.doutb(w_asqrt38_35[1]),.doutc(w_asqrt38_35[2]),.din(w_asqrt38_11[1]));
	jspl3 jspl3_w_asqrt38_36(.douta(w_asqrt38_36[0]),.doutb(w_asqrt38_36[1]),.doutc(w_asqrt38_36[2]),.din(w_asqrt38_11[2]));
	jspl3 jspl3_w_asqrt38_37(.douta(w_asqrt38_37[0]),.doutb(w_asqrt38_37[1]),.doutc(w_asqrt38_37[2]),.din(w_asqrt38_12[0]));
	jspl3 jspl3_w_asqrt38_38(.douta(w_asqrt38_38[0]),.doutb(w_asqrt38_38[1]),.doutc(w_asqrt38_38[2]),.din(w_asqrt38_12[1]));
	jspl3 jspl3_w_asqrt38_39(.douta(w_asqrt38_39[0]),.doutb(w_asqrt38_39[1]),.doutc(w_asqrt38_39[2]),.din(w_asqrt38_12[2]));
	jspl jspl_w_asqrt38_40(.douta(w_asqrt38_40),.doutb(asqrt[37]),.din(w_asqrt38_13[0]));
	jspl3 jspl3_w_asqrt39_0(.douta(w_asqrt39_0[0]),.doutb(w_asqrt39_0[1]),.doutc(w_asqrt39_0[2]),.din(asqrt_fa_39));
	jspl3 jspl3_w_asqrt39_1(.douta(w_asqrt39_1[0]),.doutb(w_asqrt39_1[1]),.doutc(w_asqrt39_1[2]),.din(w_asqrt39_0[0]));
	jspl3 jspl3_w_asqrt39_2(.douta(w_asqrt39_2[0]),.doutb(w_asqrt39_2[1]),.doutc(w_asqrt39_2[2]),.din(w_asqrt39_0[1]));
	jspl3 jspl3_w_asqrt39_3(.douta(w_asqrt39_3[0]),.doutb(w_asqrt39_3[1]),.doutc(w_asqrt39_3[2]),.din(w_asqrt39_0[2]));
	jspl3 jspl3_w_asqrt39_4(.douta(w_asqrt39_4[0]),.doutb(w_asqrt39_4[1]),.doutc(w_asqrt39_4[2]),.din(w_asqrt39_1[0]));
	jspl3 jspl3_w_asqrt39_5(.douta(w_asqrt39_5[0]),.doutb(w_asqrt39_5[1]),.doutc(w_asqrt39_5[2]),.din(w_asqrt39_1[1]));
	jspl3 jspl3_w_asqrt39_6(.douta(w_asqrt39_6[0]),.doutb(w_asqrt39_6[1]),.doutc(w_asqrt39_6[2]),.din(w_asqrt39_1[2]));
	jspl3 jspl3_w_asqrt39_7(.douta(w_asqrt39_7[0]),.doutb(w_asqrt39_7[1]),.doutc(w_asqrt39_7[2]),.din(w_asqrt39_2[0]));
	jspl3 jspl3_w_asqrt39_8(.douta(w_asqrt39_8[0]),.doutb(w_asqrt39_8[1]),.doutc(w_asqrt39_8[2]),.din(w_asqrt39_2[1]));
	jspl3 jspl3_w_asqrt39_9(.douta(w_asqrt39_9[0]),.doutb(w_asqrt39_9[1]),.doutc(w_asqrt39_9[2]),.din(w_asqrt39_2[2]));
	jspl3 jspl3_w_asqrt39_10(.douta(w_asqrt39_10[0]),.doutb(w_asqrt39_10[1]),.doutc(w_asqrt39_10[2]),.din(w_asqrt39_3[0]));
	jspl3 jspl3_w_asqrt39_11(.douta(w_asqrt39_11[0]),.doutb(w_asqrt39_11[1]),.doutc(w_asqrt39_11[2]),.din(w_asqrt39_3[1]));
	jspl3 jspl3_w_asqrt39_12(.douta(w_asqrt39_12[0]),.doutb(w_asqrt39_12[1]),.doutc(w_asqrt39_12[2]),.din(w_asqrt39_3[2]));
	jspl3 jspl3_w_asqrt39_13(.douta(w_asqrt39_13[0]),.doutb(w_asqrt39_13[1]),.doutc(w_asqrt39_13[2]),.din(w_asqrt39_4[0]));
	jspl3 jspl3_w_asqrt39_14(.douta(w_asqrt39_14[0]),.doutb(w_asqrt39_14[1]),.doutc(w_asqrt39_14[2]),.din(w_asqrt39_4[1]));
	jspl3 jspl3_w_asqrt39_15(.douta(w_asqrt39_15[0]),.doutb(w_asqrt39_15[1]),.doutc(w_asqrt39_15[2]),.din(w_asqrt39_4[2]));
	jspl3 jspl3_w_asqrt39_16(.douta(w_asqrt39_16[0]),.doutb(w_asqrt39_16[1]),.doutc(w_asqrt39_16[2]),.din(w_asqrt39_5[0]));
	jspl3 jspl3_w_asqrt39_17(.douta(w_asqrt39_17[0]),.doutb(w_asqrt39_17[1]),.doutc(w_asqrt39_17[2]),.din(w_asqrt39_5[1]));
	jspl3 jspl3_w_asqrt39_18(.douta(w_asqrt39_18[0]),.doutb(w_asqrt39_18[1]),.doutc(w_asqrt39_18[2]),.din(w_asqrt39_5[2]));
	jspl3 jspl3_w_asqrt39_19(.douta(w_asqrt39_19[0]),.doutb(w_asqrt39_19[1]),.doutc(w_asqrt39_19[2]),.din(w_asqrt39_6[0]));
	jspl3 jspl3_w_asqrt39_20(.douta(w_asqrt39_20[0]),.doutb(w_asqrt39_20[1]),.doutc(w_asqrt39_20[2]),.din(w_asqrt39_6[1]));
	jspl3 jspl3_w_asqrt39_21(.douta(w_asqrt39_21[0]),.doutb(w_asqrt39_21[1]),.doutc(w_asqrt39_21[2]),.din(w_asqrt39_6[2]));
	jspl3 jspl3_w_asqrt39_22(.douta(w_asqrt39_22[0]),.doutb(w_asqrt39_22[1]),.doutc(w_asqrt39_22[2]),.din(w_asqrt39_7[0]));
	jspl3 jspl3_w_asqrt39_23(.douta(w_asqrt39_23[0]),.doutb(w_asqrt39_23[1]),.doutc(w_asqrt39_23[2]),.din(w_asqrt39_7[1]));
	jspl3 jspl3_w_asqrt39_24(.douta(w_asqrt39_24[0]),.doutb(w_asqrt39_24[1]),.doutc(w_asqrt39_24[2]),.din(w_asqrt39_7[2]));
	jspl3 jspl3_w_asqrt39_25(.douta(w_asqrt39_25[0]),.doutb(w_asqrt39_25[1]),.doutc(w_asqrt39_25[2]),.din(w_asqrt39_8[0]));
	jspl3 jspl3_w_asqrt39_26(.douta(w_asqrt39_26[0]),.doutb(w_asqrt39_26[1]),.doutc(w_asqrt39_26[2]),.din(w_asqrt39_8[1]));
	jspl3 jspl3_w_asqrt39_27(.douta(w_asqrt39_27[0]),.doutb(w_asqrt39_27[1]),.doutc(w_asqrt39_27[2]),.din(w_asqrt39_8[2]));
	jspl3 jspl3_w_asqrt39_28(.douta(w_asqrt39_28[0]),.doutb(w_asqrt39_28[1]),.doutc(w_asqrt39_28[2]),.din(w_asqrt39_9[0]));
	jspl3 jspl3_w_asqrt39_29(.douta(w_asqrt39_29[0]),.doutb(w_asqrt39_29[1]),.doutc(w_asqrt39_29[2]),.din(w_asqrt39_9[1]));
	jspl jspl_w_asqrt39_30(.douta(w_asqrt39_30),.doutb(asqrt[38]),.din(w_asqrt39_9[2]));
	jspl3 jspl3_w_asqrt40_0(.douta(w_asqrt40_0[0]),.doutb(w_asqrt40_0[1]),.doutc(w_asqrt40_0[2]),.din(asqrt_fa_40));
	jspl3 jspl3_w_asqrt40_1(.douta(w_asqrt40_1[0]),.doutb(w_asqrt40_1[1]),.doutc(w_asqrt40_1[2]),.din(w_asqrt40_0[0]));
	jspl3 jspl3_w_asqrt40_2(.douta(w_asqrt40_2[0]),.doutb(w_asqrt40_2[1]),.doutc(w_asqrt40_2[2]),.din(w_asqrt40_0[1]));
	jspl3 jspl3_w_asqrt40_3(.douta(w_asqrt40_3[0]),.doutb(w_asqrt40_3[1]),.doutc(w_asqrt40_3[2]),.din(w_asqrt40_0[2]));
	jspl3 jspl3_w_asqrt40_4(.douta(w_asqrt40_4[0]),.doutb(w_asqrt40_4[1]),.doutc(w_asqrt40_4[2]),.din(w_asqrt40_1[0]));
	jspl3 jspl3_w_asqrt40_5(.douta(w_asqrt40_5[0]),.doutb(w_asqrt40_5[1]),.doutc(w_asqrt40_5[2]),.din(w_asqrt40_1[1]));
	jspl3 jspl3_w_asqrt40_6(.douta(w_asqrt40_6[0]),.doutb(w_asqrt40_6[1]),.doutc(w_asqrt40_6[2]),.din(w_asqrt40_1[2]));
	jspl3 jspl3_w_asqrt40_7(.douta(w_asqrt40_7[0]),.doutb(w_asqrt40_7[1]),.doutc(w_asqrt40_7[2]),.din(w_asqrt40_2[0]));
	jspl3 jspl3_w_asqrt40_8(.douta(w_asqrt40_8[0]),.doutb(w_asqrt40_8[1]),.doutc(w_asqrt40_8[2]),.din(w_asqrt40_2[1]));
	jspl3 jspl3_w_asqrt40_9(.douta(w_asqrt40_9[0]),.doutb(w_asqrt40_9[1]),.doutc(w_asqrt40_9[2]),.din(w_asqrt40_2[2]));
	jspl3 jspl3_w_asqrt40_10(.douta(w_asqrt40_10[0]),.doutb(w_asqrt40_10[1]),.doutc(w_asqrt40_10[2]),.din(w_asqrt40_3[0]));
	jspl3 jspl3_w_asqrt40_11(.douta(w_asqrt40_11[0]),.doutb(w_asqrt40_11[1]),.doutc(w_asqrt40_11[2]),.din(w_asqrt40_3[1]));
	jspl3 jspl3_w_asqrt40_12(.douta(w_asqrt40_12[0]),.doutb(w_asqrt40_12[1]),.doutc(w_asqrt40_12[2]),.din(w_asqrt40_3[2]));
	jspl3 jspl3_w_asqrt40_13(.douta(w_asqrt40_13[0]),.doutb(w_asqrt40_13[1]),.doutc(w_asqrt40_13[2]),.din(w_asqrt40_4[0]));
	jspl3 jspl3_w_asqrt40_14(.douta(w_asqrt40_14[0]),.doutb(w_asqrt40_14[1]),.doutc(w_asqrt40_14[2]),.din(w_asqrt40_4[1]));
	jspl3 jspl3_w_asqrt40_15(.douta(w_asqrt40_15[0]),.doutb(w_asqrt40_15[1]),.doutc(w_asqrt40_15[2]),.din(w_asqrt40_4[2]));
	jspl3 jspl3_w_asqrt40_16(.douta(w_asqrt40_16[0]),.doutb(w_asqrt40_16[1]),.doutc(w_asqrt40_16[2]),.din(w_asqrt40_5[0]));
	jspl3 jspl3_w_asqrt40_17(.douta(w_asqrt40_17[0]),.doutb(w_asqrt40_17[1]),.doutc(w_asqrt40_17[2]),.din(w_asqrt40_5[1]));
	jspl3 jspl3_w_asqrt40_18(.douta(w_asqrt40_18[0]),.doutb(w_asqrt40_18[1]),.doutc(w_asqrt40_18[2]),.din(w_asqrt40_5[2]));
	jspl3 jspl3_w_asqrt40_19(.douta(w_asqrt40_19[0]),.doutb(w_asqrt40_19[1]),.doutc(w_asqrt40_19[2]),.din(w_asqrt40_6[0]));
	jspl3 jspl3_w_asqrt40_20(.douta(w_asqrt40_20[0]),.doutb(w_asqrt40_20[1]),.doutc(w_asqrt40_20[2]),.din(w_asqrt40_6[1]));
	jspl3 jspl3_w_asqrt40_21(.douta(w_asqrt40_21[0]),.doutb(w_asqrt40_21[1]),.doutc(w_asqrt40_21[2]),.din(w_asqrt40_6[2]));
	jspl3 jspl3_w_asqrt40_22(.douta(w_asqrt40_22[0]),.doutb(w_asqrt40_22[1]),.doutc(w_asqrt40_22[2]),.din(w_asqrt40_7[0]));
	jspl3 jspl3_w_asqrt40_23(.douta(w_asqrt40_23[0]),.doutb(w_asqrt40_23[1]),.doutc(w_asqrt40_23[2]),.din(w_asqrt40_7[1]));
	jspl3 jspl3_w_asqrt40_24(.douta(w_asqrt40_24[0]),.doutb(w_asqrt40_24[1]),.doutc(w_asqrt40_24[2]),.din(w_asqrt40_7[2]));
	jspl3 jspl3_w_asqrt40_25(.douta(w_asqrt40_25[0]),.doutb(w_asqrt40_25[1]),.doutc(w_asqrt40_25[2]),.din(w_asqrt40_8[0]));
	jspl3 jspl3_w_asqrt40_26(.douta(w_asqrt40_26[0]),.doutb(w_asqrt40_26[1]),.doutc(w_asqrt40_26[2]),.din(w_asqrt40_8[1]));
	jspl3 jspl3_w_asqrt40_27(.douta(w_asqrt40_27[0]),.doutb(w_asqrt40_27[1]),.doutc(w_asqrt40_27[2]),.din(w_asqrt40_8[2]));
	jspl3 jspl3_w_asqrt40_28(.douta(w_asqrt40_28[0]),.doutb(w_asqrt40_28[1]),.doutc(w_asqrt40_28[2]),.din(w_asqrt40_9[0]));
	jspl3 jspl3_w_asqrt40_29(.douta(w_asqrt40_29[0]),.doutb(w_asqrt40_29[1]),.doutc(w_asqrt40_29[2]),.din(w_asqrt40_9[1]));
	jspl3 jspl3_w_asqrt40_30(.douta(w_asqrt40_30[0]),.doutb(w_asqrt40_30[1]),.doutc(w_asqrt40_30[2]),.din(w_asqrt40_9[2]));
	jspl3 jspl3_w_asqrt40_31(.douta(w_asqrt40_31[0]),.doutb(w_asqrt40_31[1]),.doutc(w_asqrt40_31[2]),.din(w_asqrt40_10[0]));
	jspl3 jspl3_w_asqrt40_32(.douta(w_asqrt40_32[0]),.doutb(w_asqrt40_32[1]),.doutc(w_asqrt40_32[2]),.din(w_asqrt40_10[1]));
	jspl3 jspl3_w_asqrt40_33(.douta(w_asqrt40_33[0]),.doutb(w_asqrt40_33[1]),.doutc(w_asqrt40_33[2]),.din(w_asqrt40_10[2]));
	jspl3 jspl3_w_asqrt40_34(.douta(w_asqrt40_34[0]),.doutb(w_asqrt40_34[1]),.doutc(w_asqrt40_34[2]),.din(w_asqrt40_11[0]));
	jspl3 jspl3_w_asqrt40_35(.douta(w_asqrt40_35[0]),.doutb(w_asqrt40_35[1]),.doutc(w_asqrt40_35[2]),.din(w_asqrt40_11[1]));
	jspl3 jspl3_w_asqrt40_36(.douta(w_asqrt40_36[0]),.doutb(w_asqrt40_36[1]),.doutc(w_asqrt40_36[2]),.din(w_asqrt40_11[2]));
	jspl3 jspl3_w_asqrt40_37(.douta(w_asqrt40_37[0]),.doutb(w_asqrt40_37[1]),.doutc(w_asqrt40_37[2]),.din(w_asqrt40_12[0]));
	jspl3 jspl3_w_asqrt40_38(.douta(w_asqrt40_38[0]),.doutb(w_asqrt40_38[1]),.doutc(w_asqrt40_38[2]),.din(w_asqrt40_12[1]));
	jspl3 jspl3_w_asqrt40_39(.douta(w_asqrt40_39[0]),.doutb(w_asqrt40_39[1]),.doutc(w_asqrt40_39[2]),.din(w_asqrt40_12[2]));
	jspl3 jspl3_w_asqrt40_40(.douta(w_asqrt40_40[0]),.doutb(w_asqrt40_40[1]),.doutc(asqrt[39]),.din(w_asqrt40_13[0]));
	jspl3 jspl3_w_asqrt41_0(.douta(w_asqrt41_0[0]),.doutb(w_asqrt41_0[1]),.doutc(w_asqrt41_0[2]),.din(asqrt_fa_41));
	jspl3 jspl3_w_asqrt41_1(.douta(w_asqrt41_1[0]),.doutb(w_asqrt41_1[1]),.doutc(w_asqrt41_1[2]),.din(w_asqrt41_0[0]));
	jspl3 jspl3_w_asqrt41_2(.douta(w_asqrt41_2[0]),.doutb(w_asqrt41_2[1]),.doutc(w_asqrt41_2[2]),.din(w_asqrt41_0[1]));
	jspl3 jspl3_w_asqrt41_3(.douta(w_asqrt41_3[0]),.doutb(w_asqrt41_3[1]),.doutc(w_asqrt41_3[2]),.din(w_asqrt41_0[2]));
	jspl3 jspl3_w_asqrt41_4(.douta(w_asqrt41_4[0]),.doutb(w_asqrt41_4[1]),.doutc(w_asqrt41_4[2]),.din(w_asqrt41_1[0]));
	jspl3 jspl3_w_asqrt41_5(.douta(w_asqrt41_5[0]),.doutb(w_asqrt41_5[1]),.doutc(w_asqrt41_5[2]),.din(w_asqrt41_1[1]));
	jspl3 jspl3_w_asqrt41_6(.douta(w_asqrt41_6[0]),.doutb(w_asqrt41_6[1]),.doutc(w_asqrt41_6[2]),.din(w_asqrt41_1[2]));
	jspl3 jspl3_w_asqrt41_7(.douta(w_asqrt41_7[0]),.doutb(w_asqrt41_7[1]),.doutc(w_asqrt41_7[2]),.din(w_asqrt41_2[0]));
	jspl3 jspl3_w_asqrt41_8(.douta(w_asqrt41_8[0]),.doutb(w_asqrt41_8[1]),.doutc(w_asqrt41_8[2]),.din(w_asqrt41_2[1]));
	jspl3 jspl3_w_asqrt41_9(.douta(w_asqrt41_9[0]),.doutb(w_asqrt41_9[1]),.doutc(w_asqrt41_9[2]),.din(w_asqrt41_2[2]));
	jspl3 jspl3_w_asqrt41_10(.douta(w_asqrt41_10[0]),.doutb(w_asqrt41_10[1]),.doutc(w_asqrt41_10[2]),.din(w_asqrt41_3[0]));
	jspl3 jspl3_w_asqrt41_11(.douta(w_asqrt41_11[0]),.doutb(w_asqrt41_11[1]),.doutc(w_asqrt41_11[2]),.din(w_asqrt41_3[1]));
	jspl3 jspl3_w_asqrt41_12(.douta(w_asqrt41_12[0]),.doutb(w_asqrt41_12[1]),.doutc(w_asqrt41_12[2]),.din(w_asqrt41_3[2]));
	jspl3 jspl3_w_asqrt41_13(.douta(w_asqrt41_13[0]),.doutb(w_asqrt41_13[1]),.doutc(w_asqrt41_13[2]),.din(w_asqrt41_4[0]));
	jspl3 jspl3_w_asqrt41_14(.douta(w_asqrt41_14[0]),.doutb(w_asqrt41_14[1]),.doutc(w_asqrt41_14[2]),.din(w_asqrt41_4[1]));
	jspl3 jspl3_w_asqrt41_15(.douta(w_asqrt41_15[0]),.doutb(w_asqrt41_15[1]),.doutc(w_asqrt41_15[2]),.din(w_asqrt41_4[2]));
	jspl3 jspl3_w_asqrt41_16(.douta(w_asqrt41_16[0]),.doutb(w_asqrt41_16[1]),.doutc(w_asqrt41_16[2]),.din(w_asqrt41_5[0]));
	jspl3 jspl3_w_asqrt41_17(.douta(w_asqrt41_17[0]),.doutb(w_asqrt41_17[1]),.doutc(w_asqrt41_17[2]),.din(w_asqrt41_5[1]));
	jspl3 jspl3_w_asqrt41_18(.douta(w_asqrt41_18[0]),.doutb(w_asqrt41_18[1]),.doutc(w_asqrt41_18[2]),.din(w_asqrt41_5[2]));
	jspl3 jspl3_w_asqrt41_19(.douta(w_asqrt41_19[0]),.doutb(w_asqrt41_19[1]),.doutc(w_asqrt41_19[2]),.din(w_asqrt41_6[0]));
	jspl3 jspl3_w_asqrt41_20(.douta(w_asqrt41_20[0]),.doutb(w_asqrt41_20[1]),.doutc(w_asqrt41_20[2]),.din(w_asqrt41_6[1]));
	jspl3 jspl3_w_asqrt41_21(.douta(w_asqrt41_21[0]),.doutb(w_asqrt41_21[1]),.doutc(w_asqrt41_21[2]),.din(w_asqrt41_6[2]));
	jspl3 jspl3_w_asqrt41_22(.douta(w_asqrt41_22[0]),.doutb(w_asqrt41_22[1]),.doutc(w_asqrt41_22[2]),.din(w_asqrt41_7[0]));
	jspl3 jspl3_w_asqrt41_23(.douta(w_asqrt41_23[0]),.doutb(w_asqrt41_23[1]),.doutc(w_asqrt41_23[2]),.din(w_asqrt41_7[1]));
	jspl3 jspl3_w_asqrt41_24(.douta(w_asqrt41_24[0]),.doutb(w_asqrt41_24[1]),.doutc(w_asqrt41_24[2]),.din(w_asqrt41_7[2]));
	jspl3 jspl3_w_asqrt41_25(.douta(w_asqrt41_25[0]),.doutb(w_asqrt41_25[1]),.doutc(w_asqrt41_25[2]),.din(w_asqrt41_8[0]));
	jspl3 jspl3_w_asqrt41_26(.douta(w_asqrt41_26[0]),.doutb(w_asqrt41_26[1]),.doutc(w_asqrt41_26[2]),.din(w_asqrt41_8[1]));
	jspl3 jspl3_w_asqrt41_27(.douta(w_asqrt41_27[0]),.doutb(w_asqrt41_27[1]),.doutc(w_asqrt41_27[2]),.din(w_asqrt41_8[2]));
	jspl3 jspl3_w_asqrt41_28(.douta(w_asqrt41_28[0]),.doutb(w_asqrt41_28[1]),.doutc(w_asqrt41_28[2]),.din(w_asqrt41_9[0]));
	jspl3 jspl3_w_asqrt41_29(.douta(w_asqrt41_29[0]),.doutb(w_asqrt41_29[1]),.doutc(w_asqrt41_29[2]),.din(w_asqrt41_9[1]));
	jspl3 jspl3_w_asqrt41_30(.douta(w_asqrt41_30[0]),.doutb(w_asqrt41_30[1]),.doutc(w_asqrt41_30[2]),.din(w_asqrt41_9[2]));
	jspl jspl_w_asqrt41_31(.douta(w_asqrt41_31),.doutb(asqrt[40]),.din(w_asqrt41_10[0]));
	jspl3 jspl3_w_asqrt42_0(.douta(w_asqrt42_0[0]),.doutb(w_asqrt42_0[1]),.doutc(w_asqrt42_0[2]),.din(asqrt_fa_42));
	jspl3 jspl3_w_asqrt42_1(.douta(w_asqrt42_1[0]),.doutb(w_asqrt42_1[1]),.doutc(w_asqrt42_1[2]),.din(w_asqrt42_0[0]));
	jspl3 jspl3_w_asqrt42_2(.douta(w_asqrt42_2[0]),.doutb(w_asqrt42_2[1]),.doutc(w_asqrt42_2[2]),.din(w_asqrt42_0[1]));
	jspl3 jspl3_w_asqrt42_3(.douta(w_asqrt42_3[0]),.doutb(w_asqrt42_3[1]),.doutc(w_asqrt42_3[2]),.din(w_asqrt42_0[2]));
	jspl3 jspl3_w_asqrt42_4(.douta(w_asqrt42_4[0]),.doutb(w_asqrt42_4[1]),.doutc(w_asqrt42_4[2]),.din(w_asqrt42_1[0]));
	jspl3 jspl3_w_asqrt42_5(.douta(w_asqrt42_5[0]),.doutb(w_asqrt42_5[1]),.doutc(w_asqrt42_5[2]),.din(w_asqrt42_1[1]));
	jspl3 jspl3_w_asqrt42_6(.douta(w_asqrt42_6[0]),.doutb(w_asqrt42_6[1]),.doutc(w_asqrt42_6[2]),.din(w_asqrt42_1[2]));
	jspl3 jspl3_w_asqrt42_7(.douta(w_asqrt42_7[0]),.doutb(w_asqrt42_7[1]),.doutc(w_asqrt42_7[2]),.din(w_asqrt42_2[0]));
	jspl3 jspl3_w_asqrt42_8(.douta(w_asqrt42_8[0]),.doutb(w_asqrt42_8[1]),.doutc(w_asqrt42_8[2]),.din(w_asqrt42_2[1]));
	jspl3 jspl3_w_asqrt42_9(.douta(w_asqrt42_9[0]),.doutb(w_asqrt42_9[1]),.doutc(w_asqrt42_9[2]),.din(w_asqrt42_2[2]));
	jspl3 jspl3_w_asqrt42_10(.douta(w_asqrt42_10[0]),.doutb(w_asqrt42_10[1]),.doutc(w_asqrt42_10[2]),.din(w_asqrt42_3[0]));
	jspl3 jspl3_w_asqrt42_11(.douta(w_asqrt42_11[0]),.doutb(w_asqrt42_11[1]),.doutc(w_asqrt42_11[2]),.din(w_asqrt42_3[1]));
	jspl3 jspl3_w_asqrt42_12(.douta(w_asqrt42_12[0]),.doutb(w_asqrt42_12[1]),.doutc(w_asqrt42_12[2]),.din(w_asqrt42_3[2]));
	jspl3 jspl3_w_asqrt42_13(.douta(w_asqrt42_13[0]),.doutb(w_asqrt42_13[1]),.doutc(w_asqrt42_13[2]),.din(w_asqrt42_4[0]));
	jspl3 jspl3_w_asqrt42_14(.douta(w_asqrt42_14[0]),.doutb(w_asqrt42_14[1]),.doutc(w_asqrt42_14[2]),.din(w_asqrt42_4[1]));
	jspl3 jspl3_w_asqrt42_15(.douta(w_asqrt42_15[0]),.doutb(w_asqrt42_15[1]),.doutc(w_asqrt42_15[2]),.din(w_asqrt42_4[2]));
	jspl3 jspl3_w_asqrt42_16(.douta(w_asqrt42_16[0]),.doutb(w_asqrt42_16[1]),.doutc(w_asqrt42_16[2]),.din(w_asqrt42_5[0]));
	jspl3 jspl3_w_asqrt42_17(.douta(w_asqrt42_17[0]),.doutb(w_asqrt42_17[1]),.doutc(w_asqrt42_17[2]),.din(w_asqrt42_5[1]));
	jspl3 jspl3_w_asqrt42_18(.douta(w_asqrt42_18[0]),.doutb(w_asqrt42_18[1]),.doutc(w_asqrt42_18[2]),.din(w_asqrt42_5[2]));
	jspl3 jspl3_w_asqrt42_19(.douta(w_asqrt42_19[0]),.doutb(w_asqrt42_19[1]),.doutc(w_asqrt42_19[2]),.din(w_asqrt42_6[0]));
	jspl3 jspl3_w_asqrt42_20(.douta(w_asqrt42_20[0]),.doutb(w_asqrt42_20[1]),.doutc(w_asqrt42_20[2]),.din(w_asqrt42_6[1]));
	jspl3 jspl3_w_asqrt42_21(.douta(w_asqrt42_21[0]),.doutb(w_asqrt42_21[1]),.doutc(w_asqrt42_21[2]),.din(w_asqrt42_6[2]));
	jspl3 jspl3_w_asqrt42_22(.douta(w_asqrt42_22[0]),.doutb(w_asqrt42_22[1]),.doutc(w_asqrt42_22[2]),.din(w_asqrt42_7[0]));
	jspl3 jspl3_w_asqrt42_23(.douta(w_asqrt42_23[0]),.doutb(w_asqrt42_23[1]),.doutc(w_asqrt42_23[2]),.din(w_asqrt42_7[1]));
	jspl3 jspl3_w_asqrt42_24(.douta(w_asqrt42_24[0]),.doutb(w_asqrt42_24[1]),.doutc(w_asqrt42_24[2]),.din(w_asqrt42_7[2]));
	jspl3 jspl3_w_asqrt42_25(.douta(w_asqrt42_25[0]),.doutb(w_asqrt42_25[1]),.doutc(w_asqrt42_25[2]),.din(w_asqrt42_8[0]));
	jspl3 jspl3_w_asqrt42_26(.douta(w_asqrt42_26[0]),.doutb(w_asqrt42_26[1]),.doutc(w_asqrt42_26[2]),.din(w_asqrt42_8[1]));
	jspl3 jspl3_w_asqrt42_27(.douta(w_asqrt42_27[0]),.doutb(w_asqrt42_27[1]),.doutc(w_asqrt42_27[2]),.din(w_asqrt42_8[2]));
	jspl3 jspl3_w_asqrt42_28(.douta(w_asqrt42_28[0]),.doutb(w_asqrt42_28[1]),.doutc(w_asqrt42_28[2]),.din(w_asqrt42_9[0]));
	jspl3 jspl3_w_asqrt42_29(.douta(w_asqrt42_29[0]),.doutb(w_asqrt42_29[1]),.doutc(w_asqrt42_29[2]),.din(w_asqrt42_9[1]));
	jspl3 jspl3_w_asqrt42_30(.douta(w_asqrt42_30[0]),.doutb(w_asqrt42_30[1]),.doutc(w_asqrt42_30[2]),.din(w_asqrt42_9[2]));
	jspl3 jspl3_w_asqrt42_31(.douta(w_asqrt42_31[0]),.doutb(w_asqrt42_31[1]),.doutc(w_asqrt42_31[2]),.din(w_asqrt42_10[0]));
	jspl3 jspl3_w_asqrt42_32(.douta(w_asqrt42_32[0]),.doutb(w_asqrt42_32[1]),.doutc(w_asqrt42_32[2]),.din(w_asqrt42_10[1]));
	jspl3 jspl3_w_asqrt42_33(.douta(w_asqrt42_33[0]),.doutb(w_asqrt42_33[1]),.doutc(w_asqrt42_33[2]),.din(w_asqrt42_10[2]));
	jspl3 jspl3_w_asqrt42_34(.douta(w_asqrt42_34[0]),.doutb(w_asqrt42_34[1]),.doutc(w_asqrt42_34[2]),.din(w_asqrt42_11[0]));
	jspl3 jspl3_w_asqrt42_35(.douta(w_asqrt42_35[0]),.doutb(w_asqrt42_35[1]),.doutc(w_asqrt42_35[2]),.din(w_asqrt42_11[1]));
	jspl3 jspl3_w_asqrt42_36(.douta(w_asqrt42_36[0]),.doutb(w_asqrt42_36[1]),.doutc(w_asqrt42_36[2]),.din(w_asqrt42_11[2]));
	jspl3 jspl3_w_asqrt42_37(.douta(w_asqrt42_37[0]),.doutb(w_asqrt42_37[1]),.doutc(w_asqrt42_37[2]),.din(w_asqrt42_12[0]));
	jspl3 jspl3_w_asqrt42_38(.douta(w_asqrt42_38[0]),.doutb(w_asqrt42_38[1]),.doutc(w_asqrt42_38[2]),.din(w_asqrt42_12[1]));
	jspl3 jspl3_w_asqrt42_39(.douta(w_asqrt42_39[0]),.doutb(w_asqrt42_39[1]),.doutc(w_asqrt42_39[2]),.din(w_asqrt42_12[2]));
	jspl3 jspl3_w_asqrt42_40(.douta(w_asqrt42_40[0]),.doutb(w_asqrt42_40[1]),.doutc(w_asqrt42_40[2]),.din(w_asqrt42_13[0]));
	jspl jspl_w_asqrt42_41(.douta(w_asqrt42_41),.doutb(asqrt[41]),.din(w_asqrt42_13[1]));
	jspl3 jspl3_w_asqrt43_0(.douta(w_asqrt43_0[0]),.doutb(w_asqrt43_0[1]),.doutc(w_asqrt43_0[2]),.din(asqrt_fa_43));
	jspl3 jspl3_w_asqrt43_1(.douta(w_asqrt43_1[0]),.doutb(w_asqrt43_1[1]),.doutc(w_asqrt43_1[2]),.din(w_asqrt43_0[0]));
	jspl3 jspl3_w_asqrt43_2(.douta(w_asqrt43_2[0]),.doutb(w_asqrt43_2[1]),.doutc(w_asqrt43_2[2]),.din(w_asqrt43_0[1]));
	jspl3 jspl3_w_asqrt43_3(.douta(w_asqrt43_3[0]),.doutb(w_asqrt43_3[1]),.doutc(w_asqrt43_3[2]),.din(w_asqrt43_0[2]));
	jspl3 jspl3_w_asqrt43_4(.douta(w_asqrt43_4[0]),.doutb(w_asqrt43_4[1]),.doutc(w_asqrt43_4[2]),.din(w_asqrt43_1[0]));
	jspl3 jspl3_w_asqrt43_5(.douta(w_asqrt43_5[0]),.doutb(w_asqrt43_5[1]),.doutc(w_asqrt43_5[2]),.din(w_asqrt43_1[1]));
	jspl3 jspl3_w_asqrt43_6(.douta(w_asqrt43_6[0]),.doutb(w_asqrt43_6[1]),.doutc(w_asqrt43_6[2]),.din(w_asqrt43_1[2]));
	jspl3 jspl3_w_asqrt43_7(.douta(w_asqrt43_7[0]),.doutb(w_asqrt43_7[1]),.doutc(w_asqrt43_7[2]),.din(w_asqrt43_2[0]));
	jspl3 jspl3_w_asqrt43_8(.douta(w_asqrt43_8[0]),.doutb(w_asqrt43_8[1]),.doutc(w_asqrt43_8[2]),.din(w_asqrt43_2[1]));
	jspl3 jspl3_w_asqrt43_9(.douta(w_asqrt43_9[0]),.doutb(w_asqrt43_9[1]),.doutc(w_asqrt43_9[2]),.din(w_asqrt43_2[2]));
	jspl3 jspl3_w_asqrt43_10(.douta(w_asqrt43_10[0]),.doutb(w_asqrt43_10[1]),.doutc(w_asqrt43_10[2]),.din(w_asqrt43_3[0]));
	jspl3 jspl3_w_asqrt43_11(.douta(w_asqrt43_11[0]),.doutb(w_asqrt43_11[1]),.doutc(w_asqrt43_11[2]),.din(w_asqrt43_3[1]));
	jspl3 jspl3_w_asqrt43_12(.douta(w_asqrt43_12[0]),.doutb(w_asqrt43_12[1]),.doutc(w_asqrt43_12[2]),.din(w_asqrt43_3[2]));
	jspl3 jspl3_w_asqrt43_13(.douta(w_asqrt43_13[0]),.doutb(w_asqrt43_13[1]),.doutc(w_asqrt43_13[2]),.din(w_asqrt43_4[0]));
	jspl3 jspl3_w_asqrt43_14(.douta(w_asqrt43_14[0]),.doutb(w_asqrt43_14[1]),.doutc(w_asqrt43_14[2]),.din(w_asqrt43_4[1]));
	jspl3 jspl3_w_asqrt43_15(.douta(w_asqrt43_15[0]),.doutb(w_asqrt43_15[1]),.doutc(w_asqrt43_15[2]),.din(w_asqrt43_4[2]));
	jspl3 jspl3_w_asqrt43_16(.douta(w_asqrt43_16[0]),.doutb(w_asqrt43_16[1]),.doutc(w_asqrt43_16[2]),.din(w_asqrt43_5[0]));
	jspl3 jspl3_w_asqrt43_17(.douta(w_asqrt43_17[0]),.doutb(w_asqrt43_17[1]),.doutc(w_asqrt43_17[2]),.din(w_asqrt43_5[1]));
	jspl3 jspl3_w_asqrt43_18(.douta(w_asqrt43_18[0]),.doutb(w_asqrt43_18[1]),.doutc(w_asqrt43_18[2]),.din(w_asqrt43_5[2]));
	jspl3 jspl3_w_asqrt43_19(.douta(w_asqrt43_19[0]),.doutb(w_asqrt43_19[1]),.doutc(w_asqrt43_19[2]),.din(w_asqrt43_6[0]));
	jspl3 jspl3_w_asqrt43_20(.douta(w_asqrt43_20[0]),.doutb(w_asqrt43_20[1]),.doutc(w_asqrt43_20[2]),.din(w_asqrt43_6[1]));
	jspl3 jspl3_w_asqrt43_21(.douta(w_asqrt43_21[0]),.doutb(w_asqrt43_21[1]),.doutc(w_asqrt43_21[2]),.din(w_asqrt43_6[2]));
	jspl3 jspl3_w_asqrt43_22(.douta(w_asqrt43_22[0]),.doutb(w_asqrt43_22[1]),.doutc(w_asqrt43_22[2]),.din(w_asqrt43_7[0]));
	jspl3 jspl3_w_asqrt43_23(.douta(w_asqrt43_23[0]),.doutb(w_asqrt43_23[1]),.doutc(w_asqrt43_23[2]),.din(w_asqrt43_7[1]));
	jspl3 jspl3_w_asqrt43_24(.douta(w_asqrt43_24[0]),.doutb(w_asqrt43_24[1]),.doutc(w_asqrt43_24[2]),.din(w_asqrt43_7[2]));
	jspl3 jspl3_w_asqrt43_25(.douta(w_asqrt43_25[0]),.doutb(w_asqrt43_25[1]),.doutc(w_asqrt43_25[2]),.din(w_asqrt43_8[0]));
	jspl3 jspl3_w_asqrt43_26(.douta(w_asqrt43_26[0]),.doutb(w_asqrt43_26[1]),.doutc(w_asqrt43_26[2]),.din(w_asqrt43_8[1]));
	jspl3 jspl3_w_asqrt43_27(.douta(w_asqrt43_27[0]),.doutb(w_asqrt43_27[1]),.doutc(w_asqrt43_27[2]),.din(w_asqrt43_8[2]));
	jspl3 jspl3_w_asqrt43_28(.douta(w_asqrt43_28[0]),.doutb(w_asqrt43_28[1]),.doutc(w_asqrt43_28[2]),.din(w_asqrt43_9[0]));
	jspl3 jspl3_w_asqrt43_29(.douta(w_asqrt43_29[0]),.doutb(w_asqrt43_29[1]),.doutc(w_asqrt43_29[2]),.din(w_asqrt43_9[1]));
	jspl3 jspl3_w_asqrt43_30(.douta(w_asqrt43_30[0]),.doutb(w_asqrt43_30[1]),.doutc(w_asqrt43_30[2]),.din(w_asqrt43_9[2]));
	jspl3 jspl3_w_asqrt43_31(.douta(w_asqrt43_31[0]),.doutb(w_asqrt43_31[1]),.doutc(w_asqrt43_31[2]),.din(w_asqrt43_10[0]));
	jspl3 jspl3_w_asqrt43_32(.douta(w_asqrt43_32[0]),.doutb(w_asqrt43_32[1]),.doutc(asqrt[42]),.din(w_asqrt43_10[1]));
	jspl3 jspl3_w_asqrt44_0(.douta(w_asqrt44_0[0]),.doutb(w_asqrt44_0[1]),.doutc(w_asqrt44_0[2]),.din(asqrt_fa_44));
	jspl3 jspl3_w_asqrt44_1(.douta(w_asqrt44_1[0]),.doutb(w_asqrt44_1[1]),.doutc(w_asqrt44_1[2]),.din(w_asqrt44_0[0]));
	jspl3 jspl3_w_asqrt44_2(.douta(w_asqrt44_2[0]),.doutb(w_asqrt44_2[1]),.doutc(w_asqrt44_2[2]),.din(w_asqrt44_0[1]));
	jspl3 jspl3_w_asqrt44_3(.douta(w_asqrt44_3[0]),.doutb(w_asqrt44_3[1]),.doutc(w_asqrt44_3[2]),.din(w_asqrt44_0[2]));
	jspl3 jspl3_w_asqrt44_4(.douta(w_asqrt44_4[0]),.doutb(w_asqrt44_4[1]),.doutc(w_asqrt44_4[2]),.din(w_asqrt44_1[0]));
	jspl3 jspl3_w_asqrt44_5(.douta(w_asqrt44_5[0]),.doutb(w_asqrt44_5[1]),.doutc(w_asqrt44_5[2]),.din(w_asqrt44_1[1]));
	jspl3 jspl3_w_asqrt44_6(.douta(w_asqrt44_6[0]),.doutb(w_asqrt44_6[1]),.doutc(w_asqrt44_6[2]),.din(w_asqrt44_1[2]));
	jspl3 jspl3_w_asqrt44_7(.douta(w_asqrt44_7[0]),.doutb(w_asqrt44_7[1]),.doutc(w_asqrt44_7[2]),.din(w_asqrt44_2[0]));
	jspl3 jspl3_w_asqrt44_8(.douta(w_asqrt44_8[0]),.doutb(w_asqrt44_8[1]),.doutc(w_asqrt44_8[2]),.din(w_asqrt44_2[1]));
	jspl3 jspl3_w_asqrt44_9(.douta(w_asqrt44_9[0]),.doutb(w_asqrt44_9[1]),.doutc(w_asqrt44_9[2]),.din(w_asqrt44_2[2]));
	jspl3 jspl3_w_asqrt44_10(.douta(w_asqrt44_10[0]),.doutb(w_asqrt44_10[1]),.doutc(w_asqrt44_10[2]),.din(w_asqrt44_3[0]));
	jspl3 jspl3_w_asqrt44_11(.douta(w_asqrt44_11[0]),.doutb(w_asqrt44_11[1]),.doutc(w_asqrt44_11[2]),.din(w_asqrt44_3[1]));
	jspl3 jspl3_w_asqrt44_12(.douta(w_asqrt44_12[0]),.doutb(w_asqrt44_12[1]),.doutc(w_asqrt44_12[2]),.din(w_asqrt44_3[2]));
	jspl3 jspl3_w_asqrt44_13(.douta(w_asqrt44_13[0]),.doutb(w_asqrt44_13[1]),.doutc(w_asqrt44_13[2]),.din(w_asqrt44_4[0]));
	jspl3 jspl3_w_asqrt44_14(.douta(w_asqrt44_14[0]),.doutb(w_asqrt44_14[1]),.doutc(w_asqrt44_14[2]),.din(w_asqrt44_4[1]));
	jspl3 jspl3_w_asqrt44_15(.douta(w_asqrt44_15[0]),.doutb(w_asqrt44_15[1]),.doutc(w_asqrt44_15[2]),.din(w_asqrt44_4[2]));
	jspl3 jspl3_w_asqrt44_16(.douta(w_asqrt44_16[0]),.doutb(w_asqrt44_16[1]),.doutc(w_asqrt44_16[2]),.din(w_asqrt44_5[0]));
	jspl3 jspl3_w_asqrt44_17(.douta(w_asqrt44_17[0]),.doutb(w_asqrt44_17[1]),.doutc(w_asqrt44_17[2]),.din(w_asqrt44_5[1]));
	jspl3 jspl3_w_asqrt44_18(.douta(w_asqrt44_18[0]),.doutb(w_asqrt44_18[1]),.doutc(w_asqrt44_18[2]),.din(w_asqrt44_5[2]));
	jspl3 jspl3_w_asqrt44_19(.douta(w_asqrt44_19[0]),.doutb(w_asqrt44_19[1]),.doutc(w_asqrt44_19[2]),.din(w_asqrt44_6[0]));
	jspl3 jspl3_w_asqrt44_20(.douta(w_asqrt44_20[0]),.doutb(w_asqrt44_20[1]),.doutc(w_asqrt44_20[2]),.din(w_asqrt44_6[1]));
	jspl3 jspl3_w_asqrt44_21(.douta(w_asqrt44_21[0]),.doutb(w_asqrt44_21[1]),.doutc(w_asqrt44_21[2]),.din(w_asqrt44_6[2]));
	jspl3 jspl3_w_asqrt44_22(.douta(w_asqrt44_22[0]),.doutb(w_asqrt44_22[1]),.doutc(w_asqrt44_22[2]),.din(w_asqrt44_7[0]));
	jspl3 jspl3_w_asqrt44_23(.douta(w_asqrt44_23[0]),.doutb(w_asqrt44_23[1]),.doutc(w_asqrt44_23[2]),.din(w_asqrt44_7[1]));
	jspl3 jspl3_w_asqrt44_24(.douta(w_asqrt44_24[0]),.doutb(w_asqrt44_24[1]),.doutc(w_asqrt44_24[2]),.din(w_asqrt44_7[2]));
	jspl3 jspl3_w_asqrt44_25(.douta(w_asqrt44_25[0]),.doutb(w_asqrt44_25[1]),.doutc(w_asqrt44_25[2]),.din(w_asqrt44_8[0]));
	jspl3 jspl3_w_asqrt44_26(.douta(w_asqrt44_26[0]),.doutb(w_asqrt44_26[1]),.doutc(w_asqrt44_26[2]),.din(w_asqrt44_8[1]));
	jspl3 jspl3_w_asqrt44_27(.douta(w_asqrt44_27[0]),.doutb(w_asqrt44_27[1]),.doutc(w_asqrt44_27[2]),.din(w_asqrt44_8[2]));
	jspl3 jspl3_w_asqrt44_28(.douta(w_asqrt44_28[0]),.doutb(w_asqrt44_28[1]),.doutc(w_asqrt44_28[2]),.din(w_asqrt44_9[0]));
	jspl3 jspl3_w_asqrt44_29(.douta(w_asqrt44_29[0]),.doutb(w_asqrt44_29[1]),.doutc(w_asqrt44_29[2]),.din(w_asqrt44_9[1]));
	jspl3 jspl3_w_asqrt44_30(.douta(w_asqrt44_30[0]),.doutb(w_asqrt44_30[1]),.doutc(w_asqrt44_30[2]),.din(w_asqrt44_9[2]));
	jspl3 jspl3_w_asqrt44_31(.douta(w_asqrt44_31[0]),.doutb(w_asqrt44_31[1]),.doutc(w_asqrt44_31[2]),.din(w_asqrt44_10[0]));
	jspl3 jspl3_w_asqrt44_32(.douta(w_asqrt44_32[0]),.doutb(w_asqrt44_32[1]),.doutc(w_asqrt44_32[2]),.din(w_asqrt44_10[1]));
	jspl3 jspl3_w_asqrt44_33(.douta(w_asqrt44_33[0]),.doutb(w_asqrt44_33[1]),.doutc(w_asqrt44_33[2]),.din(w_asqrt44_10[2]));
	jspl3 jspl3_w_asqrt44_34(.douta(w_asqrt44_34[0]),.doutb(w_asqrt44_34[1]),.doutc(w_asqrt44_34[2]),.din(w_asqrt44_11[0]));
	jspl3 jspl3_w_asqrt44_35(.douta(w_asqrt44_35[0]),.doutb(w_asqrt44_35[1]),.doutc(w_asqrt44_35[2]),.din(w_asqrt44_11[1]));
	jspl3 jspl3_w_asqrt44_36(.douta(w_asqrt44_36[0]),.doutb(w_asqrt44_36[1]),.doutc(w_asqrt44_36[2]),.din(w_asqrt44_11[2]));
	jspl3 jspl3_w_asqrt44_37(.douta(w_asqrt44_37[0]),.doutb(w_asqrt44_37[1]),.doutc(w_asqrt44_37[2]),.din(w_asqrt44_12[0]));
	jspl3 jspl3_w_asqrt44_38(.douta(w_asqrt44_38[0]),.doutb(w_asqrt44_38[1]),.doutc(w_asqrt44_38[2]),.din(w_asqrt44_12[1]));
	jspl3 jspl3_w_asqrt44_39(.douta(w_asqrt44_39[0]),.doutb(w_asqrt44_39[1]),.doutc(w_asqrt44_39[2]),.din(w_asqrt44_12[2]));
	jspl3 jspl3_w_asqrt44_40(.douta(w_asqrt44_40[0]),.doutb(w_asqrt44_40[1]),.doutc(w_asqrt44_40[2]),.din(w_asqrt44_13[0]));
	jspl jspl_w_asqrt44_41(.douta(w_asqrt44_41),.doutb(asqrt[43]),.din(w_asqrt44_13[1]));
	jspl3 jspl3_w_asqrt45_0(.douta(w_asqrt45_0[0]),.doutb(w_asqrt45_0[1]),.doutc(w_asqrt45_0[2]),.din(asqrt_fa_45));
	jspl3 jspl3_w_asqrt45_1(.douta(w_asqrt45_1[0]),.doutb(w_asqrt45_1[1]),.doutc(w_asqrt45_1[2]),.din(w_asqrt45_0[0]));
	jspl3 jspl3_w_asqrt45_2(.douta(w_asqrt45_2[0]),.doutb(w_asqrt45_2[1]),.doutc(w_asqrt45_2[2]),.din(w_asqrt45_0[1]));
	jspl3 jspl3_w_asqrt45_3(.douta(w_asqrt45_3[0]),.doutb(w_asqrt45_3[1]),.doutc(w_asqrt45_3[2]),.din(w_asqrt45_0[2]));
	jspl3 jspl3_w_asqrt45_4(.douta(w_asqrt45_4[0]),.doutb(w_asqrt45_4[1]),.doutc(w_asqrt45_4[2]),.din(w_asqrt45_1[0]));
	jspl3 jspl3_w_asqrt45_5(.douta(w_asqrt45_5[0]),.doutb(w_asqrt45_5[1]),.doutc(w_asqrt45_5[2]),.din(w_asqrt45_1[1]));
	jspl3 jspl3_w_asqrt45_6(.douta(w_asqrt45_6[0]),.doutb(w_asqrt45_6[1]),.doutc(w_asqrt45_6[2]),.din(w_asqrt45_1[2]));
	jspl3 jspl3_w_asqrt45_7(.douta(w_asqrt45_7[0]),.doutb(w_asqrt45_7[1]),.doutc(w_asqrt45_7[2]),.din(w_asqrt45_2[0]));
	jspl3 jspl3_w_asqrt45_8(.douta(w_asqrt45_8[0]),.doutb(w_asqrt45_8[1]),.doutc(w_asqrt45_8[2]),.din(w_asqrt45_2[1]));
	jspl3 jspl3_w_asqrt45_9(.douta(w_asqrt45_9[0]),.doutb(w_asqrt45_9[1]),.doutc(w_asqrt45_9[2]),.din(w_asqrt45_2[2]));
	jspl3 jspl3_w_asqrt45_10(.douta(w_asqrt45_10[0]),.doutb(w_asqrt45_10[1]),.doutc(w_asqrt45_10[2]),.din(w_asqrt45_3[0]));
	jspl3 jspl3_w_asqrt45_11(.douta(w_asqrt45_11[0]),.doutb(w_asqrt45_11[1]),.doutc(w_asqrt45_11[2]),.din(w_asqrt45_3[1]));
	jspl3 jspl3_w_asqrt45_12(.douta(w_asqrt45_12[0]),.doutb(w_asqrt45_12[1]),.doutc(w_asqrt45_12[2]),.din(w_asqrt45_3[2]));
	jspl3 jspl3_w_asqrt45_13(.douta(w_asqrt45_13[0]),.doutb(w_asqrt45_13[1]),.doutc(w_asqrt45_13[2]),.din(w_asqrt45_4[0]));
	jspl3 jspl3_w_asqrt45_14(.douta(w_asqrt45_14[0]),.doutb(w_asqrt45_14[1]),.doutc(w_asqrt45_14[2]),.din(w_asqrt45_4[1]));
	jspl3 jspl3_w_asqrt45_15(.douta(w_asqrt45_15[0]),.doutb(w_asqrt45_15[1]),.doutc(w_asqrt45_15[2]),.din(w_asqrt45_4[2]));
	jspl3 jspl3_w_asqrt45_16(.douta(w_asqrt45_16[0]),.doutb(w_asqrt45_16[1]),.doutc(w_asqrt45_16[2]),.din(w_asqrt45_5[0]));
	jspl3 jspl3_w_asqrt45_17(.douta(w_asqrt45_17[0]),.doutb(w_asqrt45_17[1]),.doutc(w_asqrt45_17[2]),.din(w_asqrt45_5[1]));
	jspl3 jspl3_w_asqrt45_18(.douta(w_asqrt45_18[0]),.doutb(w_asqrt45_18[1]),.doutc(w_asqrt45_18[2]),.din(w_asqrt45_5[2]));
	jspl3 jspl3_w_asqrt45_19(.douta(w_asqrt45_19[0]),.doutb(w_asqrt45_19[1]),.doutc(w_asqrt45_19[2]),.din(w_asqrt45_6[0]));
	jspl3 jspl3_w_asqrt45_20(.douta(w_asqrt45_20[0]),.doutb(w_asqrt45_20[1]),.doutc(w_asqrt45_20[2]),.din(w_asqrt45_6[1]));
	jspl3 jspl3_w_asqrt45_21(.douta(w_asqrt45_21[0]),.doutb(w_asqrt45_21[1]),.doutc(w_asqrt45_21[2]),.din(w_asqrt45_6[2]));
	jspl3 jspl3_w_asqrt45_22(.douta(w_asqrt45_22[0]),.doutb(w_asqrt45_22[1]),.doutc(w_asqrt45_22[2]),.din(w_asqrt45_7[0]));
	jspl3 jspl3_w_asqrt45_23(.douta(w_asqrt45_23[0]),.doutb(w_asqrt45_23[1]),.doutc(w_asqrt45_23[2]),.din(w_asqrt45_7[1]));
	jspl3 jspl3_w_asqrt45_24(.douta(w_asqrt45_24[0]),.doutb(w_asqrt45_24[1]),.doutc(w_asqrt45_24[2]),.din(w_asqrt45_7[2]));
	jspl3 jspl3_w_asqrt45_25(.douta(w_asqrt45_25[0]),.doutb(w_asqrt45_25[1]),.doutc(w_asqrt45_25[2]),.din(w_asqrt45_8[0]));
	jspl3 jspl3_w_asqrt45_26(.douta(w_asqrt45_26[0]),.doutb(w_asqrt45_26[1]),.doutc(w_asqrt45_26[2]),.din(w_asqrt45_8[1]));
	jspl3 jspl3_w_asqrt45_27(.douta(w_asqrt45_27[0]),.doutb(w_asqrt45_27[1]),.doutc(w_asqrt45_27[2]),.din(w_asqrt45_8[2]));
	jspl3 jspl3_w_asqrt45_28(.douta(w_asqrt45_28[0]),.doutb(w_asqrt45_28[1]),.doutc(w_asqrt45_28[2]),.din(w_asqrt45_9[0]));
	jspl3 jspl3_w_asqrt45_29(.douta(w_asqrt45_29[0]),.doutb(w_asqrt45_29[1]),.doutc(w_asqrt45_29[2]),.din(w_asqrt45_9[1]));
	jspl3 jspl3_w_asqrt45_30(.douta(w_asqrt45_30[0]),.doutb(w_asqrt45_30[1]),.doutc(w_asqrt45_30[2]),.din(w_asqrt45_9[2]));
	jspl3 jspl3_w_asqrt45_31(.douta(w_asqrt45_31[0]),.doutb(w_asqrt45_31[1]),.doutc(w_asqrt45_31[2]),.din(w_asqrt45_10[0]));
	jspl3 jspl3_w_asqrt45_32(.douta(w_asqrt45_32[0]),.doutb(w_asqrt45_32[1]),.doutc(w_asqrt45_32[2]),.din(w_asqrt45_10[1]));
	jspl3 jspl3_w_asqrt45_33(.douta(w_asqrt45_33[0]),.doutb(w_asqrt45_33[1]),.doutc(w_asqrt45_33[2]),.din(w_asqrt45_10[2]));
	jspl jspl_w_asqrt45_34(.douta(w_asqrt45_34),.doutb(asqrt[44]),.din(w_asqrt45_11[0]));
	jspl3 jspl3_w_asqrt46_0(.douta(w_asqrt46_0[0]),.doutb(w_asqrt46_0[1]),.doutc(w_asqrt46_0[2]),.din(asqrt_fa_46));
	jspl3 jspl3_w_asqrt46_1(.douta(w_asqrt46_1[0]),.doutb(w_asqrt46_1[1]),.doutc(w_asqrt46_1[2]),.din(w_asqrt46_0[0]));
	jspl3 jspl3_w_asqrt46_2(.douta(w_asqrt46_2[0]),.doutb(w_asqrt46_2[1]),.doutc(w_asqrt46_2[2]),.din(w_asqrt46_0[1]));
	jspl3 jspl3_w_asqrt46_3(.douta(w_asqrt46_3[0]),.doutb(w_asqrt46_3[1]),.doutc(w_asqrt46_3[2]),.din(w_asqrt46_0[2]));
	jspl3 jspl3_w_asqrt46_4(.douta(w_asqrt46_4[0]),.doutb(w_asqrt46_4[1]),.doutc(w_asqrt46_4[2]),.din(w_asqrt46_1[0]));
	jspl3 jspl3_w_asqrt46_5(.douta(w_asqrt46_5[0]),.doutb(w_asqrt46_5[1]),.doutc(w_asqrt46_5[2]),.din(w_asqrt46_1[1]));
	jspl3 jspl3_w_asqrt46_6(.douta(w_asqrt46_6[0]),.doutb(w_asqrt46_6[1]),.doutc(w_asqrt46_6[2]),.din(w_asqrt46_1[2]));
	jspl3 jspl3_w_asqrt46_7(.douta(w_asqrt46_7[0]),.doutb(w_asqrt46_7[1]),.doutc(w_asqrt46_7[2]),.din(w_asqrt46_2[0]));
	jspl3 jspl3_w_asqrt46_8(.douta(w_asqrt46_8[0]),.doutb(w_asqrt46_8[1]),.doutc(w_asqrt46_8[2]),.din(w_asqrt46_2[1]));
	jspl3 jspl3_w_asqrt46_9(.douta(w_asqrt46_9[0]),.doutb(w_asqrt46_9[1]),.doutc(w_asqrt46_9[2]),.din(w_asqrt46_2[2]));
	jspl3 jspl3_w_asqrt46_10(.douta(w_asqrt46_10[0]),.doutb(w_asqrt46_10[1]),.doutc(w_asqrt46_10[2]),.din(w_asqrt46_3[0]));
	jspl3 jspl3_w_asqrt46_11(.douta(w_asqrt46_11[0]),.doutb(w_asqrt46_11[1]),.doutc(w_asqrt46_11[2]),.din(w_asqrt46_3[1]));
	jspl3 jspl3_w_asqrt46_12(.douta(w_asqrt46_12[0]),.doutb(w_asqrt46_12[1]),.doutc(w_asqrt46_12[2]),.din(w_asqrt46_3[2]));
	jspl3 jspl3_w_asqrt46_13(.douta(w_asqrt46_13[0]),.doutb(w_asqrt46_13[1]),.doutc(w_asqrt46_13[2]),.din(w_asqrt46_4[0]));
	jspl3 jspl3_w_asqrt46_14(.douta(w_asqrt46_14[0]),.doutb(w_asqrt46_14[1]),.doutc(w_asqrt46_14[2]),.din(w_asqrt46_4[1]));
	jspl3 jspl3_w_asqrt46_15(.douta(w_asqrt46_15[0]),.doutb(w_asqrt46_15[1]),.doutc(w_asqrt46_15[2]),.din(w_asqrt46_4[2]));
	jspl3 jspl3_w_asqrt46_16(.douta(w_asqrt46_16[0]),.doutb(w_asqrt46_16[1]),.doutc(w_asqrt46_16[2]),.din(w_asqrt46_5[0]));
	jspl3 jspl3_w_asqrt46_17(.douta(w_asqrt46_17[0]),.doutb(w_asqrt46_17[1]),.doutc(w_asqrt46_17[2]),.din(w_asqrt46_5[1]));
	jspl3 jspl3_w_asqrt46_18(.douta(w_asqrt46_18[0]),.doutb(w_asqrt46_18[1]),.doutc(w_asqrt46_18[2]),.din(w_asqrt46_5[2]));
	jspl3 jspl3_w_asqrt46_19(.douta(w_asqrt46_19[0]),.doutb(w_asqrt46_19[1]),.doutc(w_asqrt46_19[2]),.din(w_asqrt46_6[0]));
	jspl3 jspl3_w_asqrt46_20(.douta(w_asqrt46_20[0]),.doutb(w_asqrt46_20[1]),.doutc(w_asqrt46_20[2]),.din(w_asqrt46_6[1]));
	jspl3 jspl3_w_asqrt46_21(.douta(w_asqrt46_21[0]),.doutb(w_asqrt46_21[1]),.doutc(w_asqrt46_21[2]),.din(w_asqrt46_6[2]));
	jspl3 jspl3_w_asqrt46_22(.douta(w_asqrt46_22[0]),.doutb(w_asqrt46_22[1]),.doutc(w_asqrt46_22[2]),.din(w_asqrt46_7[0]));
	jspl3 jspl3_w_asqrt46_23(.douta(w_asqrt46_23[0]),.doutb(w_asqrt46_23[1]),.doutc(w_asqrt46_23[2]),.din(w_asqrt46_7[1]));
	jspl3 jspl3_w_asqrt46_24(.douta(w_asqrt46_24[0]),.doutb(w_asqrt46_24[1]),.doutc(w_asqrt46_24[2]),.din(w_asqrt46_7[2]));
	jspl3 jspl3_w_asqrt46_25(.douta(w_asqrt46_25[0]),.doutb(w_asqrt46_25[1]),.doutc(w_asqrt46_25[2]),.din(w_asqrt46_8[0]));
	jspl3 jspl3_w_asqrt46_26(.douta(w_asqrt46_26[0]),.doutb(w_asqrt46_26[1]),.doutc(w_asqrt46_26[2]),.din(w_asqrt46_8[1]));
	jspl3 jspl3_w_asqrt46_27(.douta(w_asqrt46_27[0]),.doutb(w_asqrt46_27[1]),.doutc(w_asqrt46_27[2]),.din(w_asqrt46_8[2]));
	jspl3 jspl3_w_asqrt46_28(.douta(w_asqrt46_28[0]),.doutb(w_asqrt46_28[1]),.doutc(w_asqrt46_28[2]),.din(w_asqrt46_9[0]));
	jspl3 jspl3_w_asqrt46_29(.douta(w_asqrt46_29[0]),.doutb(w_asqrt46_29[1]),.doutc(w_asqrt46_29[2]),.din(w_asqrt46_9[1]));
	jspl3 jspl3_w_asqrt46_30(.douta(w_asqrt46_30[0]),.doutb(w_asqrt46_30[1]),.doutc(w_asqrt46_30[2]),.din(w_asqrt46_9[2]));
	jspl3 jspl3_w_asqrt46_31(.douta(w_asqrt46_31[0]),.doutb(w_asqrt46_31[1]),.doutc(w_asqrt46_31[2]),.din(w_asqrt46_10[0]));
	jspl3 jspl3_w_asqrt46_32(.douta(w_asqrt46_32[0]),.doutb(w_asqrt46_32[1]),.doutc(w_asqrt46_32[2]),.din(w_asqrt46_10[1]));
	jspl3 jspl3_w_asqrt46_33(.douta(w_asqrt46_33[0]),.doutb(w_asqrt46_33[1]),.doutc(w_asqrt46_33[2]),.din(w_asqrt46_10[2]));
	jspl3 jspl3_w_asqrt46_34(.douta(w_asqrt46_34[0]),.doutb(w_asqrt46_34[1]),.doutc(w_asqrt46_34[2]),.din(w_asqrt46_11[0]));
	jspl3 jspl3_w_asqrt46_35(.douta(w_asqrt46_35[0]),.doutb(w_asqrt46_35[1]),.doutc(w_asqrt46_35[2]),.din(w_asqrt46_11[1]));
	jspl3 jspl3_w_asqrt46_36(.douta(w_asqrt46_36[0]),.doutb(w_asqrt46_36[1]),.doutc(w_asqrt46_36[2]),.din(w_asqrt46_11[2]));
	jspl3 jspl3_w_asqrt46_37(.douta(w_asqrt46_37[0]),.doutb(w_asqrt46_37[1]),.doutc(w_asqrt46_37[2]),.din(w_asqrt46_12[0]));
	jspl3 jspl3_w_asqrt46_38(.douta(w_asqrt46_38[0]),.doutb(w_asqrt46_38[1]),.doutc(w_asqrt46_38[2]),.din(w_asqrt46_12[1]));
	jspl3 jspl3_w_asqrt46_39(.douta(w_asqrt46_39[0]),.doutb(w_asqrt46_39[1]),.doutc(w_asqrt46_39[2]),.din(w_asqrt46_12[2]));
	jspl3 jspl3_w_asqrt46_40(.douta(w_asqrt46_40[0]),.doutb(w_asqrt46_40[1]),.doutc(w_asqrt46_40[2]),.din(w_asqrt46_13[0]));
	jspl3 jspl3_w_asqrt46_41(.douta(w_asqrt46_41[0]),.doutb(w_asqrt46_41[1]),.doutc(asqrt[45]),.din(w_asqrt46_13[1]));
	jspl3 jspl3_w_asqrt47_0(.douta(w_asqrt47_0[0]),.doutb(w_asqrt47_0[1]),.doutc(w_asqrt47_0[2]),.din(asqrt_fa_47));
	jspl3 jspl3_w_asqrt47_1(.douta(w_asqrt47_1[0]),.doutb(w_asqrt47_1[1]),.doutc(w_asqrt47_1[2]),.din(w_asqrt47_0[0]));
	jspl3 jspl3_w_asqrt47_2(.douta(w_asqrt47_2[0]),.doutb(w_asqrt47_2[1]),.doutc(w_asqrt47_2[2]),.din(w_asqrt47_0[1]));
	jspl3 jspl3_w_asqrt47_3(.douta(w_asqrt47_3[0]),.doutb(w_asqrt47_3[1]),.doutc(w_asqrt47_3[2]),.din(w_asqrt47_0[2]));
	jspl3 jspl3_w_asqrt47_4(.douta(w_asqrt47_4[0]),.doutb(w_asqrt47_4[1]),.doutc(w_asqrt47_4[2]),.din(w_asqrt47_1[0]));
	jspl3 jspl3_w_asqrt47_5(.douta(w_asqrt47_5[0]),.doutb(w_asqrt47_5[1]),.doutc(w_asqrt47_5[2]),.din(w_asqrt47_1[1]));
	jspl3 jspl3_w_asqrt47_6(.douta(w_asqrt47_6[0]),.doutb(w_asqrt47_6[1]),.doutc(w_asqrt47_6[2]),.din(w_asqrt47_1[2]));
	jspl3 jspl3_w_asqrt47_7(.douta(w_asqrt47_7[0]),.doutb(w_asqrt47_7[1]),.doutc(w_asqrt47_7[2]),.din(w_asqrt47_2[0]));
	jspl3 jspl3_w_asqrt47_8(.douta(w_asqrt47_8[0]),.doutb(w_asqrt47_8[1]),.doutc(w_asqrt47_8[2]),.din(w_asqrt47_2[1]));
	jspl3 jspl3_w_asqrt47_9(.douta(w_asqrt47_9[0]),.doutb(w_asqrt47_9[1]),.doutc(w_asqrt47_9[2]),.din(w_asqrt47_2[2]));
	jspl3 jspl3_w_asqrt47_10(.douta(w_asqrt47_10[0]),.doutb(w_asqrt47_10[1]),.doutc(w_asqrt47_10[2]),.din(w_asqrt47_3[0]));
	jspl3 jspl3_w_asqrt47_11(.douta(w_asqrt47_11[0]),.doutb(w_asqrt47_11[1]),.doutc(w_asqrt47_11[2]),.din(w_asqrt47_3[1]));
	jspl3 jspl3_w_asqrt47_12(.douta(w_asqrt47_12[0]),.doutb(w_asqrt47_12[1]),.doutc(w_asqrt47_12[2]),.din(w_asqrt47_3[2]));
	jspl3 jspl3_w_asqrt47_13(.douta(w_asqrt47_13[0]),.doutb(w_asqrt47_13[1]),.doutc(w_asqrt47_13[2]),.din(w_asqrt47_4[0]));
	jspl3 jspl3_w_asqrt47_14(.douta(w_asqrt47_14[0]),.doutb(w_asqrt47_14[1]),.doutc(w_asqrt47_14[2]),.din(w_asqrt47_4[1]));
	jspl3 jspl3_w_asqrt47_15(.douta(w_asqrt47_15[0]),.doutb(w_asqrt47_15[1]),.doutc(w_asqrt47_15[2]),.din(w_asqrt47_4[2]));
	jspl3 jspl3_w_asqrt47_16(.douta(w_asqrt47_16[0]),.doutb(w_asqrt47_16[1]),.doutc(w_asqrt47_16[2]),.din(w_asqrt47_5[0]));
	jspl3 jspl3_w_asqrt47_17(.douta(w_asqrt47_17[0]),.doutb(w_asqrt47_17[1]),.doutc(w_asqrt47_17[2]),.din(w_asqrt47_5[1]));
	jspl3 jspl3_w_asqrt47_18(.douta(w_asqrt47_18[0]),.doutb(w_asqrt47_18[1]),.doutc(w_asqrt47_18[2]),.din(w_asqrt47_5[2]));
	jspl3 jspl3_w_asqrt47_19(.douta(w_asqrt47_19[0]),.doutb(w_asqrt47_19[1]),.doutc(w_asqrt47_19[2]),.din(w_asqrt47_6[0]));
	jspl3 jspl3_w_asqrt47_20(.douta(w_asqrt47_20[0]),.doutb(w_asqrt47_20[1]),.doutc(w_asqrt47_20[2]),.din(w_asqrt47_6[1]));
	jspl3 jspl3_w_asqrt47_21(.douta(w_asqrt47_21[0]),.doutb(w_asqrt47_21[1]),.doutc(w_asqrt47_21[2]),.din(w_asqrt47_6[2]));
	jspl3 jspl3_w_asqrt47_22(.douta(w_asqrt47_22[0]),.doutb(w_asqrt47_22[1]),.doutc(w_asqrt47_22[2]),.din(w_asqrt47_7[0]));
	jspl3 jspl3_w_asqrt47_23(.douta(w_asqrt47_23[0]),.doutb(w_asqrt47_23[1]),.doutc(w_asqrt47_23[2]),.din(w_asqrt47_7[1]));
	jspl3 jspl3_w_asqrt47_24(.douta(w_asqrt47_24[0]),.doutb(w_asqrt47_24[1]),.doutc(w_asqrt47_24[2]),.din(w_asqrt47_7[2]));
	jspl3 jspl3_w_asqrt47_25(.douta(w_asqrt47_25[0]),.doutb(w_asqrt47_25[1]),.doutc(w_asqrt47_25[2]),.din(w_asqrt47_8[0]));
	jspl3 jspl3_w_asqrt47_26(.douta(w_asqrt47_26[0]),.doutb(w_asqrt47_26[1]),.doutc(w_asqrt47_26[2]),.din(w_asqrt47_8[1]));
	jspl3 jspl3_w_asqrt47_27(.douta(w_asqrt47_27[0]),.doutb(w_asqrt47_27[1]),.doutc(w_asqrt47_27[2]),.din(w_asqrt47_8[2]));
	jspl3 jspl3_w_asqrt47_28(.douta(w_asqrt47_28[0]),.doutb(w_asqrt47_28[1]),.doutc(w_asqrt47_28[2]),.din(w_asqrt47_9[0]));
	jspl3 jspl3_w_asqrt47_29(.douta(w_asqrt47_29[0]),.doutb(w_asqrt47_29[1]),.doutc(w_asqrt47_29[2]),.din(w_asqrt47_9[1]));
	jspl3 jspl3_w_asqrt47_30(.douta(w_asqrt47_30[0]),.doutb(w_asqrt47_30[1]),.doutc(w_asqrt47_30[2]),.din(w_asqrt47_9[2]));
	jspl3 jspl3_w_asqrt47_31(.douta(w_asqrt47_31[0]),.doutb(w_asqrt47_31[1]),.doutc(w_asqrt47_31[2]),.din(w_asqrt47_10[0]));
	jspl3 jspl3_w_asqrt47_32(.douta(w_asqrt47_32[0]),.doutb(w_asqrt47_32[1]),.doutc(w_asqrt47_32[2]),.din(w_asqrt47_10[1]));
	jspl3 jspl3_w_asqrt47_33(.douta(w_asqrt47_33[0]),.doutb(w_asqrt47_33[1]),.doutc(w_asqrt47_33[2]),.din(w_asqrt47_10[2]));
	jspl3 jspl3_w_asqrt47_34(.douta(w_asqrt47_34[0]),.doutb(w_asqrt47_34[1]),.doutc(w_asqrt47_34[2]),.din(w_asqrt47_11[0]));
	jspl3 jspl3_w_asqrt47_35(.douta(w_asqrt47_35[0]),.doutb(w_asqrt47_35[1]),.doutc(w_asqrt47_35[2]),.din(w_asqrt47_11[1]));
	jspl jspl_w_asqrt47_36(.douta(w_asqrt47_36),.doutb(asqrt[46]),.din(w_asqrt47_11[2]));
	jspl3 jspl3_w_asqrt48_0(.douta(w_asqrt48_0[0]),.doutb(w_asqrt48_0[1]),.doutc(w_asqrt48_0[2]),.din(asqrt_fa_48));
	jspl3 jspl3_w_asqrt48_1(.douta(w_asqrt48_1[0]),.doutb(w_asqrt48_1[1]),.doutc(w_asqrt48_1[2]),.din(w_asqrt48_0[0]));
	jspl3 jspl3_w_asqrt48_2(.douta(w_asqrt48_2[0]),.doutb(w_asqrt48_2[1]),.doutc(w_asqrt48_2[2]),.din(w_asqrt48_0[1]));
	jspl3 jspl3_w_asqrt48_3(.douta(w_asqrt48_3[0]),.doutb(w_asqrt48_3[1]),.doutc(w_asqrt48_3[2]),.din(w_asqrt48_0[2]));
	jspl3 jspl3_w_asqrt48_4(.douta(w_asqrt48_4[0]),.doutb(w_asqrt48_4[1]),.doutc(w_asqrt48_4[2]),.din(w_asqrt48_1[0]));
	jspl3 jspl3_w_asqrt48_5(.douta(w_asqrt48_5[0]),.doutb(w_asqrt48_5[1]),.doutc(w_asqrt48_5[2]),.din(w_asqrt48_1[1]));
	jspl3 jspl3_w_asqrt48_6(.douta(w_asqrt48_6[0]),.doutb(w_asqrt48_6[1]),.doutc(w_asqrt48_6[2]),.din(w_asqrt48_1[2]));
	jspl3 jspl3_w_asqrt48_7(.douta(w_asqrt48_7[0]),.doutb(w_asqrt48_7[1]),.doutc(w_asqrt48_7[2]),.din(w_asqrt48_2[0]));
	jspl3 jspl3_w_asqrt48_8(.douta(w_asqrt48_8[0]),.doutb(w_asqrt48_8[1]),.doutc(w_asqrt48_8[2]),.din(w_asqrt48_2[1]));
	jspl3 jspl3_w_asqrt48_9(.douta(w_asqrt48_9[0]),.doutb(w_asqrt48_9[1]),.doutc(w_asqrt48_9[2]),.din(w_asqrt48_2[2]));
	jspl3 jspl3_w_asqrt48_10(.douta(w_asqrt48_10[0]),.doutb(w_asqrt48_10[1]),.doutc(w_asqrt48_10[2]),.din(w_asqrt48_3[0]));
	jspl3 jspl3_w_asqrt48_11(.douta(w_asqrt48_11[0]),.doutb(w_asqrt48_11[1]),.doutc(w_asqrt48_11[2]),.din(w_asqrt48_3[1]));
	jspl3 jspl3_w_asqrt48_12(.douta(w_asqrt48_12[0]),.doutb(w_asqrt48_12[1]),.doutc(w_asqrt48_12[2]),.din(w_asqrt48_3[2]));
	jspl3 jspl3_w_asqrt48_13(.douta(w_asqrt48_13[0]),.doutb(w_asqrt48_13[1]),.doutc(w_asqrt48_13[2]),.din(w_asqrt48_4[0]));
	jspl3 jspl3_w_asqrt48_14(.douta(w_asqrt48_14[0]),.doutb(w_asqrt48_14[1]),.doutc(w_asqrt48_14[2]),.din(w_asqrt48_4[1]));
	jspl3 jspl3_w_asqrt48_15(.douta(w_asqrt48_15[0]),.doutb(w_asqrt48_15[1]),.doutc(w_asqrt48_15[2]),.din(w_asqrt48_4[2]));
	jspl3 jspl3_w_asqrt48_16(.douta(w_asqrt48_16[0]),.doutb(w_asqrt48_16[1]),.doutc(w_asqrt48_16[2]),.din(w_asqrt48_5[0]));
	jspl3 jspl3_w_asqrt48_17(.douta(w_asqrt48_17[0]),.doutb(w_asqrt48_17[1]),.doutc(w_asqrt48_17[2]),.din(w_asqrt48_5[1]));
	jspl3 jspl3_w_asqrt48_18(.douta(w_asqrt48_18[0]),.doutb(w_asqrt48_18[1]),.doutc(w_asqrt48_18[2]),.din(w_asqrt48_5[2]));
	jspl3 jspl3_w_asqrt48_19(.douta(w_asqrt48_19[0]),.doutb(w_asqrt48_19[1]),.doutc(w_asqrt48_19[2]),.din(w_asqrt48_6[0]));
	jspl3 jspl3_w_asqrt48_20(.douta(w_asqrt48_20[0]),.doutb(w_asqrt48_20[1]),.doutc(w_asqrt48_20[2]),.din(w_asqrt48_6[1]));
	jspl3 jspl3_w_asqrt48_21(.douta(w_asqrt48_21[0]),.doutb(w_asqrt48_21[1]),.doutc(w_asqrt48_21[2]),.din(w_asqrt48_6[2]));
	jspl3 jspl3_w_asqrt48_22(.douta(w_asqrt48_22[0]),.doutb(w_asqrt48_22[1]),.doutc(w_asqrt48_22[2]),.din(w_asqrt48_7[0]));
	jspl3 jspl3_w_asqrt48_23(.douta(w_asqrt48_23[0]),.doutb(w_asqrt48_23[1]),.doutc(w_asqrt48_23[2]),.din(w_asqrt48_7[1]));
	jspl3 jspl3_w_asqrt48_24(.douta(w_asqrt48_24[0]),.doutb(w_asqrt48_24[1]),.doutc(w_asqrt48_24[2]),.din(w_asqrt48_7[2]));
	jspl3 jspl3_w_asqrt48_25(.douta(w_asqrt48_25[0]),.doutb(w_asqrt48_25[1]),.doutc(w_asqrt48_25[2]),.din(w_asqrt48_8[0]));
	jspl3 jspl3_w_asqrt48_26(.douta(w_asqrt48_26[0]),.doutb(w_asqrt48_26[1]),.doutc(w_asqrt48_26[2]),.din(w_asqrt48_8[1]));
	jspl3 jspl3_w_asqrt48_27(.douta(w_asqrt48_27[0]),.doutb(w_asqrt48_27[1]),.doutc(w_asqrt48_27[2]),.din(w_asqrt48_8[2]));
	jspl3 jspl3_w_asqrt48_28(.douta(w_asqrt48_28[0]),.doutb(w_asqrt48_28[1]),.doutc(w_asqrt48_28[2]),.din(w_asqrt48_9[0]));
	jspl3 jspl3_w_asqrt48_29(.douta(w_asqrt48_29[0]),.doutb(w_asqrt48_29[1]),.doutc(w_asqrt48_29[2]),.din(w_asqrt48_9[1]));
	jspl3 jspl3_w_asqrt48_30(.douta(w_asqrt48_30[0]),.doutb(w_asqrt48_30[1]),.doutc(w_asqrt48_30[2]),.din(w_asqrt48_9[2]));
	jspl3 jspl3_w_asqrt48_31(.douta(w_asqrt48_31[0]),.doutb(w_asqrt48_31[1]),.doutc(w_asqrt48_31[2]),.din(w_asqrt48_10[0]));
	jspl3 jspl3_w_asqrt48_32(.douta(w_asqrt48_32[0]),.doutb(w_asqrt48_32[1]),.doutc(w_asqrt48_32[2]),.din(w_asqrt48_10[1]));
	jspl3 jspl3_w_asqrt48_33(.douta(w_asqrt48_33[0]),.doutb(w_asqrt48_33[1]),.doutc(w_asqrt48_33[2]),.din(w_asqrt48_10[2]));
	jspl3 jspl3_w_asqrt48_34(.douta(w_asqrt48_34[0]),.doutb(w_asqrt48_34[1]),.doutc(w_asqrt48_34[2]),.din(w_asqrt48_11[0]));
	jspl3 jspl3_w_asqrt48_35(.douta(w_asqrt48_35[0]),.doutb(w_asqrt48_35[1]),.doutc(w_asqrt48_35[2]),.din(w_asqrt48_11[1]));
	jspl3 jspl3_w_asqrt48_36(.douta(w_asqrt48_36[0]),.doutb(w_asqrt48_36[1]),.doutc(w_asqrt48_36[2]),.din(w_asqrt48_11[2]));
	jspl3 jspl3_w_asqrt48_37(.douta(w_asqrt48_37[0]),.doutb(w_asqrt48_37[1]),.doutc(w_asqrt48_37[2]),.din(w_asqrt48_12[0]));
	jspl3 jspl3_w_asqrt48_38(.douta(w_asqrt48_38[0]),.doutb(w_asqrt48_38[1]),.doutc(w_asqrt48_38[2]),.din(w_asqrt48_12[1]));
	jspl3 jspl3_w_asqrt48_39(.douta(w_asqrt48_39[0]),.doutb(w_asqrt48_39[1]),.doutc(w_asqrt48_39[2]),.din(w_asqrt48_12[2]));
	jspl3 jspl3_w_asqrt48_40(.douta(w_asqrt48_40[0]),.doutb(w_asqrt48_40[1]),.doutc(w_asqrt48_40[2]),.din(w_asqrt48_13[0]));
	jspl3 jspl3_w_asqrt48_41(.douta(w_asqrt48_41[0]),.doutb(w_asqrt48_41[1]),.doutc(w_asqrt48_41[2]),.din(w_asqrt48_13[1]));
	jspl jspl_w_asqrt48_42(.douta(w_asqrt48_42),.doutb(asqrt[47]),.din(w_asqrt48_13[2]));
	jspl3 jspl3_w_asqrt49_0(.douta(w_asqrt49_0[0]),.doutb(w_asqrt49_0[1]),.doutc(w_asqrt49_0[2]),.din(asqrt_fa_49));
	jspl3 jspl3_w_asqrt49_1(.douta(w_asqrt49_1[0]),.doutb(w_asqrt49_1[1]),.doutc(w_asqrt49_1[2]),.din(w_asqrt49_0[0]));
	jspl3 jspl3_w_asqrt49_2(.douta(w_asqrt49_2[0]),.doutb(w_asqrt49_2[1]),.doutc(w_asqrt49_2[2]),.din(w_asqrt49_0[1]));
	jspl3 jspl3_w_asqrt49_3(.douta(w_asqrt49_3[0]),.doutb(w_asqrt49_3[1]),.doutc(w_asqrt49_3[2]),.din(w_asqrt49_0[2]));
	jspl3 jspl3_w_asqrt49_4(.douta(w_asqrt49_4[0]),.doutb(w_asqrt49_4[1]),.doutc(w_asqrt49_4[2]),.din(w_asqrt49_1[0]));
	jspl3 jspl3_w_asqrt49_5(.douta(w_asqrt49_5[0]),.doutb(w_asqrt49_5[1]),.doutc(w_asqrt49_5[2]),.din(w_asqrt49_1[1]));
	jspl3 jspl3_w_asqrt49_6(.douta(w_asqrt49_6[0]),.doutb(w_asqrt49_6[1]),.doutc(w_asqrt49_6[2]),.din(w_asqrt49_1[2]));
	jspl3 jspl3_w_asqrt49_7(.douta(w_asqrt49_7[0]),.doutb(w_asqrt49_7[1]),.doutc(w_asqrt49_7[2]),.din(w_asqrt49_2[0]));
	jspl3 jspl3_w_asqrt49_8(.douta(w_asqrt49_8[0]),.doutb(w_asqrt49_8[1]),.doutc(w_asqrt49_8[2]),.din(w_asqrt49_2[1]));
	jspl3 jspl3_w_asqrt49_9(.douta(w_asqrt49_9[0]),.doutb(w_asqrt49_9[1]),.doutc(w_asqrt49_9[2]),.din(w_asqrt49_2[2]));
	jspl3 jspl3_w_asqrt49_10(.douta(w_asqrt49_10[0]),.doutb(w_asqrt49_10[1]),.doutc(w_asqrt49_10[2]),.din(w_asqrt49_3[0]));
	jspl3 jspl3_w_asqrt49_11(.douta(w_asqrt49_11[0]),.doutb(w_asqrt49_11[1]),.doutc(w_asqrt49_11[2]),.din(w_asqrt49_3[1]));
	jspl3 jspl3_w_asqrt49_12(.douta(w_asqrt49_12[0]),.doutb(w_asqrt49_12[1]),.doutc(w_asqrt49_12[2]),.din(w_asqrt49_3[2]));
	jspl3 jspl3_w_asqrt49_13(.douta(w_asqrt49_13[0]),.doutb(w_asqrt49_13[1]),.doutc(w_asqrt49_13[2]),.din(w_asqrt49_4[0]));
	jspl3 jspl3_w_asqrt49_14(.douta(w_asqrt49_14[0]),.doutb(w_asqrt49_14[1]),.doutc(w_asqrt49_14[2]),.din(w_asqrt49_4[1]));
	jspl3 jspl3_w_asqrt49_15(.douta(w_asqrt49_15[0]),.doutb(w_asqrt49_15[1]),.doutc(w_asqrt49_15[2]),.din(w_asqrt49_4[2]));
	jspl3 jspl3_w_asqrt49_16(.douta(w_asqrt49_16[0]),.doutb(w_asqrt49_16[1]),.doutc(w_asqrt49_16[2]),.din(w_asqrt49_5[0]));
	jspl3 jspl3_w_asqrt49_17(.douta(w_asqrt49_17[0]),.doutb(w_asqrt49_17[1]),.doutc(w_asqrt49_17[2]),.din(w_asqrt49_5[1]));
	jspl3 jspl3_w_asqrt49_18(.douta(w_asqrt49_18[0]),.doutb(w_asqrt49_18[1]),.doutc(w_asqrt49_18[2]),.din(w_asqrt49_5[2]));
	jspl3 jspl3_w_asqrt49_19(.douta(w_asqrt49_19[0]),.doutb(w_asqrt49_19[1]),.doutc(w_asqrt49_19[2]),.din(w_asqrt49_6[0]));
	jspl3 jspl3_w_asqrt49_20(.douta(w_asqrt49_20[0]),.doutb(w_asqrt49_20[1]),.doutc(w_asqrt49_20[2]),.din(w_asqrt49_6[1]));
	jspl3 jspl3_w_asqrt49_21(.douta(w_asqrt49_21[0]),.doutb(w_asqrt49_21[1]),.doutc(w_asqrt49_21[2]),.din(w_asqrt49_6[2]));
	jspl3 jspl3_w_asqrt49_22(.douta(w_asqrt49_22[0]),.doutb(w_asqrt49_22[1]),.doutc(w_asqrt49_22[2]),.din(w_asqrt49_7[0]));
	jspl3 jspl3_w_asqrt49_23(.douta(w_asqrt49_23[0]),.doutb(w_asqrt49_23[1]),.doutc(w_asqrt49_23[2]),.din(w_asqrt49_7[1]));
	jspl3 jspl3_w_asqrt49_24(.douta(w_asqrt49_24[0]),.doutb(w_asqrt49_24[1]),.doutc(w_asqrt49_24[2]),.din(w_asqrt49_7[2]));
	jspl3 jspl3_w_asqrt49_25(.douta(w_asqrt49_25[0]),.doutb(w_asqrt49_25[1]),.doutc(w_asqrt49_25[2]),.din(w_asqrt49_8[0]));
	jspl3 jspl3_w_asqrt49_26(.douta(w_asqrt49_26[0]),.doutb(w_asqrt49_26[1]),.doutc(w_asqrt49_26[2]),.din(w_asqrt49_8[1]));
	jspl3 jspl3_w_asqrt49_27(.douta(w_asqrt49_27[0]),.doutb(w_asqrt49_27[1]),.doutc(w_asqrt49_27[2]),.din(w_asqrt49_8[2]));
	jspl3 jspl3_w_asqrt49_28(.douta(w_asqrt49_28[0]),.doutb(w_asqrt49_28[1]),.doutc(w_asqrt49_28[2]),.din(w_asqrt49_9[0]));
	jspl3 jspl3_w_asqrt49_29(.douta(w_asqrt49_29[0]),.doutb(w_asqrt49_29[1]),.doutc(w_asqrt49_29[2]),.din(w_asqrt49_9[1]));
	jspl3 jspl3_w_asqrt49_30(.douta(w_asqrt49_30[0]),.doutb(w_asqrt49_30[1]),.doutc(w_asqrt49_30[2]),.din(w_asqrt49_9[2]));
	jspl3 jspl3_w_asqrt49_31(.douta(w_asqrt49_31[0]),.doutb(w_asqrt49_31[1]),.doutc(w_asqrt49_31[2]),.din(w_asqrt49_10[0]));
	jspl3 jspl3_w_asqrt49_32(.douta(w_asqrt49_32[0]),.doutb(w_asqrt49_32[1]),.doutc(w_asqrt49_32[2]),.din(w_asqrt49_10[1]));
	jspl3 jspl3_w_asqrt49_33(.douta(w_asqrt49_33[0]),.doutb(w_asqrt49_33[1]),.doutc(w_asqrt49_33[2]),.din(w_asqrt49_10[2]));
	jspl3 jspl3_w_asqrt49_34(.douta(w_asqrt49_34[0]),.doutb(w_asqrt49_34[1]),.doutc(w_asqrt49_34[2]),.din(w_asqrt49_11[0]));
	jspl3 jspl3_w_asqrt49_35(.douta(w_asqrt49_35[0]),.doutb(w_asqrt49_35[1]),.doutc(w_asqrt49_35[2]),.din(w_asqrt49_11[1]));
	jspl3 jspl3_w_asqrt49_36(.douta(w_asqrt49_36[0]),.doutb(w_asqrt49_36[1]),.doutc(w_asqrt49_36[2]),.din(w_asqrt49_11[2]));
	jspl3 jspl3_w_asqrt49_37(.douta(w_asqrt49_37[0]),.doutb(w_asqrt49_37[1]),.doutc(asqrt[48]),.din(w_asqrt49_12[0]));
	jspl3 jspl3_w_asqrt50_0(.douta(w_asqrt50_0[0]),.doutb(w_asqrt50_0[1]),.doutc(w_asqrt50_0[2]),.din(asqrt_fa_50));
	jspl3 jspl3_w_asqrt50_1(.douta(w_asqrt50_1[0]),.doutb(w_asqrt50_1[1]),.doutc(w_asqrt50_1[2]),.din(w_asqrt50_0[0]));
	jspl3 jspl3_w_asqrt50_2(.douta(w_asqrt50_2[0]),.doutb(w_asqrt50_2[1]),.doutc(w_asqrt50_2[2]),.din(w_asqrt50_0[1]));
	jspl3 jspl3_w_asqrt50_3(.douta(w_asqrt50_3[0]),.doutb(w_asqrt50_3[1]),.doutc(w_asqrt50_3[2]),.din(w_asqrt50_0[2]));
	jspl3 jspl3_w_asqrt50_4(.douta(w_asqrt50_4[0]),.doutb(w_asqrt50_4[1]),.doutc(w_asqrt50_4[2]),.din(w_asqrt50_1[0]));
	jspl3 jspl3_w_asqrt50_5(.douta(w_asqrt50_5[0]),.doutb(w_asqrt50_5[1]),.doutc(w_asqrt50_5[2]),.din(w_asqrt50_1[1]));
	jspl3 jspl3_w_asqrt50_6(.douta(w_asqrt50_6[0]),.doutb(w_asqrt50_6[1]),.doutc(w_asqrt50_6[2]),.din(w_asqrt50_1[2]));
	jspl3 jspl3_w_asqrt50_7(.douta(w_asqrt50_7[0]),.doutb(w_asqrt50_7[1]),.doutc(w_asqrt50_7[2]),.din(w_asqrt50_2[0]));
	jspl3 jspl3_w_asqrt50_8(.douta(w_asqrt50_8[0]),.doutb(w_asqrt50_8[1]),.doutc(w_asqrt50_8[2]),.din(w_asqrt50_2[1]));
	jspl3 jspl3_w_asqrt50_9(.douta(w_asqrt50_9[0]),.doutb(w_asqrt50_9[1]),.doutc(w_asqrt50_9[2]),.din(w_asqrt50_2[2]));
	jspl3 jspl3_w_asqrt50_10(.douta(w_asqrt50_10[0]),.doutb(w_asqrt50_10[1]),.doutc(w_asqrt50_10[2]),.din(w_asqrt50_3[0]));
	jspl3 jspl3_w_asqrt50_11(.douta(w_asqrt50_11[0]),.doutb(w_asqrt50_11[1]),.doutc(w_asqrt50_11[2]),.din(w_asqrt50_3[1]));
	jspl3 jspl3_w_asqrt50_12(.douta(w_asqrt50_12[0]),.doutb(w_asqrt50_12[1]),.doutc(w_asqrt50_12[2]),.din(w_asqrt50_3[2]));
	jspl3 jspl3_w_asqrt50_13(.douta(w_asqrt50_13[0]),.doutb(w_asqrt50_13[1]),.doutc(w_asqrt50_13[2]),.din(w_asqrt50_4[0]));
	jspl3 jspl3_w_asqrt50_14(.douta(w_asqrt50_14[0]),.doutb(w_asqrt50_14[1]),.doutc(w_asqrt50_14[2]),.din(w_asqrt50_4[1]));
	jspl3 jspl3_w_asqrt50_15(.douta(w_asqrt50_15[0]),.doutb(w_asqrt50_15[1]),.doutc(w_asqrt50_15[2]),.din(w_asqrt50_4[2]));
	jspl3 jspl3_w_asqrt50_16(.douta(w_asqrt50_16[0]),.doutb(w_asqrt50_16[1]),.doutc(w_asqrt50_16[2]),.din(w_asqrt50_5[0]));
	jspl3 jspl3_w_asqrt50_17(.douta(w_asqrt50_17[0]),.doutb(w_asqrt50_17[1]),.doutc(w_asqrt50_17[2]),.din(w_asqrt50_5[1]));
	jspl3 jspl3_w_asqrt50_18(.douta(w_asqrt50_18[0]),.doutb(w_asqrt50_18[1]),.doutc(w_asqrt50_18[2]),.din(w_asqrt50_5[2]));
	jspl3 jspl3_w_asqrt50_19(.douta(w_asqrt50_19[0]),.doutb(w_asqrt50_19[1]),.doutc(w_asqrt50_19[2]),.din(w_asqrt50_6[0]));
	jspl3 jspl3_w_asqrt50_20(.douta(w_asqrt50_20[0]),.doutb(w_asqrt50_20[1]),.doutc(w_asqrt50_20[2]),.din(w_asqrt50_6[1]));
	jspl3 jspl3_w_asqrt50_21(.douta(w_asqrt50_21[0]),.doutb(w_asqrt50_21[1]),.doutc(w_asqrt50_21[2]),.din(w_asqrt50_6[2]));
	jspl3 jspl3_w_asqrt50_22(.douta(w_asqrt50_22[0]),.doutb(w_asqrt50_22[1]),.doutc(w_asqrt50_22[2]),.din(w_asqrt50_7[0]));
	jspl3 jspl3_w_asqrt50_23(.douta(w_asqrt50_23[0]),.doutb(w_asqrt50_23[1]),.doutc(w_asqrt50_23[2]),.din(w_asqrt50_7[1]));
	jspl3 jspl3_w_asqrt50_24(.douta(w_asqrt50_24[0]),.doutb(w_asqrt50_24[1]),.doutc(w_asqrt50_24[2]),.din(w_asqrt50_7[2]));
	jspl3 jspl3_w_asqrt50_25(.douta(w_asqrt50_25[0]),.doutb(w_asqrt50_25[1]),.doutc(w_asqrt50_25[2]),.din(w_asqrt50_8[0]));
	jspl3 jspl3_w_asqrt50_26(.douta(w_asqrt50_26[0]),.doutb(w_asqrt50_26[1]),.doutc(w_asqrt50_26[2]),.din(w_asqrt50_8[1]));
	jspl3 jspl3_w_asqrt50_27(.douta(w_asqrt50_27[0]),.doutb(w_asqrt50_27[1]),.doutc(w_asqrt50_27[2]),.din(w_asqrt50_8[2]));
	jspl3 jspl3_w_asqrt50_28(.douta(w_asqrt50_28[0]),.doutb(w_asqrt50_28[1]),.doutc(w_asqrt50_28[2]),.din(w_asqrt50_9[0]));
	jspl3 jspl3_w_asqrt50_29(.douta(w_asqrt50_29[0]),.doutb(w_asqrt50_29[1]),.doutc(w_asqrt50_29[2]),.din(w_asqrt50_9[1]));
	jspl3 jspl3_w_asqrt50_30(.douta(w_asqrt50_30[0]),.doutb(w_asqrt50_30[1]),.doutc(w_asqrt50_30[2]),.din(w_asqrt50_9[2]));
	jspl3 jspl3_w_asqrt50_31(.douta(w_asqrt50_31[0]),.doutb(w_asqrt50_31[1]),.doutc(w_asqrt50_31[2]),.din(w_asqrt50_10[0]));
	jspl3 jspl3_w_asqrt50_32(.douta(w_asqrt50_32[0]),.doutb(w_asqrt50_32[1]),.doutc(w_asqrt50_32[2]),.din(w_asqrt50_10[1]));
	jspl3 jspl3_w_asqrt50_33(.douta(w_asqrt50_33[0]),.doutb(w_asqrt50_33[1]),.doutc(w_asqrt50_33[2]),.din(w_asqrt50_10[2]));
	jspl3 jspl3_w_asqrt50_34(.douta(w_asqrt50_34[0]),.doutb(w_asqrt50_34[1]),.doutc(w_asqrt50_34[2]),.din(w_asqrt50_11[0]));
	jspl3 jspl3_w_asqrt50_35(.douta(w_asqrt50_35[0]),.doutb(w_asqrt50_35[1]),.doutc(w_asqrt50_35[2]),.din(w_asqrt50_11[1]));
	jspl3 jspl3_w_asqrt50_36(.douta(w_asqrt50_36[0]),.doutb(w_asqrt50_36[1]),.doutc(w_asqrt50_36[2]),.din(w_asqrt50_11[2]));
	jspl3 jspl3_w_asqrt50_37(.douta(w_asqrt50_37[0]),.doutb(w_asqrt50_37[1]),.doutc(w_asqrt50_37[2]),.din(w_asqrt50_12[0]));
	jspl3 jspl3_w_asqrt50_38(.douta(w_asqrt50_38[0]),.doutb(w_asqrt50_38[1]),.doutc(w_asqrt50_38[2]),.din(w_asqrt50_12[1]));
	jspl3 jspl3_w_asqrt50_39(.douta(w_asqrt50_39[0]),.doutb(w_asqrt50_39[1]),.doutc(w_asqrt50_39[2]),.din(w_asqrt50_12[2]));
	jspl3 jspl3_w_asqrt50_40(.douta(w_asqrt50_40[0]),.doutb(w_asqrt50_40[1]),.doutc(w_asqrt50_40[2]),.din(w_asqrt50_13[0]));
	jspl3 jspl3_w_asqrt50_41(.douta(w_asqrt50_41[0]),.doutb(w_asqrt50_41[1]),.doutc(w_asqrt50_41[2]),.din(w_asqrt50_13[1]));
	jspl3 jspl3_w_asqrt50_42(.douta(w_asqrt50_42[0]),.doutb(w_asqrt50_42[1]),.doutc(w_asqrt50_42[2]),.din(w_asqrt50_13[2]));
	jspl jspl_w_asqrt50_43(.douta(w_asqrt50_43),.doutb(asqrt[49]),.din(w_asqrt50_14[0]));
	jspl3 jspl3_w_asqrt51_0(.douta(w_asqrt51_0[0]),.doutb(w_asqrt51_0[1]),.doutc(w_asqrt51_0[2]),.din(asqrt_fa_51));
	jspl3 jspl3_w_asqrt51_1(.douta(w_asqrt51_1[0]),.doutb(w_asqrt51_1[1]),.doutc(w_asqrt51_1[2]),.din(w_asqrt51_0[0]));
	jspl3 jspl3_w_asqrt51_2(.douta(w_asqrt51_2[0]),.doutb(w_asqrt51_2[1]),.doutc(w_asqrt51_2[2]),.din(w_asqrt51_0[1]));
	jspl3 jspl3_w_asqrt51_3(.douta(w_asqrt51_3[0]),.doutb(w_asqrt51_3[1]),.doutc(w_asqrt51_3[2]),.din(w_asqrt51_0[2]));
	jspl3 jspl3_w_asqrt51_4(.douta(w_asqrt51_4[0]),.doutb(w_asqrt51_4[1]),.doutc(w_asqrt51_4[2]),.din(w_asqrt51_1[0]));
	jspl3 jspl3_w_asqrt51_5(.douta(w_asqrt51_5[0]),.doutb(w_asqrt51_5[1]),.doutc(w_asqrt51_5[2]),.din(w_asqrt51_1[1]));
	jspl3 jspl3_w_asqrt51_6(.douta(w_asqrt51_6[0]),.doutb(w_asqrt51_6[1]),.doutc(w_asqrt51_6[2]),.din(w_asqrt51_1[2]));
	jspl3 jspl3_w_asqrt51_7(.douta(w_asqrt51_7[0]),.doutb(w_asqrt51_7[1]),.doutc(w_asqrt51_7[2]),.din(w_asqrt51_2[0]));
	jspl3 jspl3_w_asqrt51_8(.douta(w_asqrt51_8[0]),.doutb(w_asqrt51_8[1]),.doutc(w_asqrt51_8[2]),.din(w_asqrt51_2[1]));
	jspl3 jspl3_w_asqrt51_9(.douta(w_asqrt51_9[0]),.doutb(w_asqrt51_9[1]),.doutc(w_asqrt51_9[2]),.din(w_asqrt51_2[2]));
	jspl3 jspl3_w_asqrt51_10(.douta(w_asqrt51_10[0]),.doutb(w_asqrt51_10[1]),.doutc(w_asqrt51_10[2]),.din(w_asqrt51_3[0]));
	jspl3 jspl3_w_asqrt51_11(.douta(w_asqrt51_11[0]),.doutb(w_asqrt51_11[1]),.doutc(w_asqrt51_11[2]),.din(w_asqrt51_3[1]));
	jspl3 jspl3_w_asqrt51_12(.douta(w_asqrt51_12[0]),.doutb(w_asqrt51_12[1]),.doutc(w_asqrt51_12[2]),.din(w_asqrt51_3[2]));
	jspl3 jspl3_w_asqrt51_13(.douta(w_asqrt51_13[0]),.doutb(w_asqrt51_13[1]),.doutc(w_asqrt51_13[2]),.din(w_asqrt51_4[0]));
	jspl3 jspl3_w_asqrt51_14(.douta(w_asqrt51_14[0]),.doutb(w_asqrt51_14[1]),.doutc(w_asqrt51_14[2]),.din(w_asqrt51_4[1]));
	jspl3 jspl3_w_asqrt51_15(.douta(w_asqrt51_15[0]),.doutb(w_asqrt51_15[1]),.doutc(w_asqrt51_15[2]),.din(w_asqrt51_4[2]));
	jspl3 jspl3_w_asqrt51_16(.douta(w_asqrt51_16[0]),.doutb(w_asqrt51_16[1]),.doutc(w_asqrt51_16[2]),.din(w_asqrt51_5[0]));
	jspl3 jspl3_w_asqrt51_17(.douta(w_asqrt51_17[0]),.doutb(w_asqrt51_17[1]),.doutc(w_asqrt51_17[2]),.din(w_asqrt51_5[1]));
	jspl3 jspl3_w_asqrt51_18(.douta(w_asqrt51_18[0]),.doutb(w_asqrt51_18[1]),.doutc(w_asqrt51_18[2]),.din(w_asqrt51_5[2]));
	jspl3 jspl3_w_asqrt51_19(.douta(w_asqrt51_19[0]),.doutb(w_asqrt51_19[1]),.doutc(w_asqrt51_19[2]),.din(w_asqrt51_6[0]));
	jspl3 jspl3_w_asqrt51_20(.douta(w_asqrt51_20[0]),.doutb(w_asqrt51_20[1]),.doutc(w_asqrt51_20[2]),.din(w_asqrt51_6[1]));
	jspl3 jspl3_w_asqrt51_21(.douta(w_asqrt51_21[0]),.doutb(w_asqrt51_21[1]),.doutc(w_asqrt51_21[2]),.din(w_asqrt51_6[2]));
	jspl3 jspl3_w_asqrt51_22(.douta(w_asqrt51_22[0]),.doutb(w_asqrt51_22[1]),.doutc(w_asqrt51_22[2]),.din(w_asqrt51_7[0]));
	jspl3 jspl3_w_asqrt51_23(.douta(w_asqrt51_23[0]),.doutb(w_asqrt51_23[1]),.doutc(w_asqrt51_23[2]),.din(w_asqrt51_7[1]));
	jspl3 jspl3_w_asqrt51_24(.douta(w_asqrt51_24[0]),.doutb(w_asqrt51_24[1]),.doutc(w_asqrt51_24[2]),.din(w_asqrt51_7[2]));
	jspl3 jspl3_w_asqrt51_25(.douta(w_asqrt51_25[0]),.doutb(w_asqrt51_25[1]),.doutc(w_asqrt51_25[2]),.din(w_asqrt51_8[0]));
	jspl3 jspl3_w_asqrt51_26(.douta(w_asqrt51_26[0]),.doutb(w_asqrt51_26[1]),.doutc(w_asqrt51_26[2]),.din(w_asqrt51_8[1]));
	jspl3 jspl3_w_asqrt51_27(.douta(w_asqrt51_27[0]),.doutb(w_asqrt51_27[1]),.doutc(w_asqrt51_27[2]),.din(w_asqrt51_8[2]));
	jspl3 jspl3_w_asqrt51_28(.douta(w_asqrt51_28[0]),.doutb(w_asqrt51_28[1]),.doutc(w_asqrt51_28[2]),.din(w_asqrt51_9[0]));
	jspl3 jspl3_w_asqrt51_29(.douta(w_asqrt51_29[0]),.doutb(w_asqrt51_29[1]),.doutc(w_asqrt51_29[2]),.din(w_asqrt51_9[1]));
	jspl3 jspl3_w_asqrt51_30(.douta(w_asqrt51_30[0]),.doutb(w_asqrt51_30[1]),.doutc(w_asqrt51_30[2]),.din(w_asqrt51_9[2]));
	jspl3 jspl3_w_asqrt51_31(.douta(w_asqrt51_31[0]),.doutb(w_asqrt51_31[1]),.doutc(w_asqrt51_31[2]),.din(w_asqrt51_10[0]));
	jspl3 jspl3_w_asqrt51_32(.douta(w_asqrt51_32[0]),.doutb(w_asqrt51_32[1]),.doutc(w_asqrt51_32[2]),.din(w_asqrt51_10[1]));
	jspl3 jspl3_w_asqrt51_33(.douta(w_asqrt51_33[0]),.doutb(w_asqrt51_33[1]),.doutc(w_asqrt51_33[2]),.din(w_asqrt51_10[2]));
	jspl3 jspl3_w_asqrt51_34(.douta(w_asqrt51_34[0]),.doutb(w_asqrt51_34[1]),.doutc(w_asqrt51_34[2]),.din(w_asqrt51_11[0]));
	jspl3 jspl3_w_asqrt51_35(.douta(w_asqrt51_35[0]),.doutb(w_asqrt51_35[1]),.doutc(w_asqrt51_35[2]),.din(w_asqrt51_11[1]));
	jspl3 jspl3_w_asqrt51_36(.douta(w_asqrt51_36[0]),.doutb(w_asqrt51_36[1]),.doutc(w_asqrt51_36[2]),.din(w_asqrt51_11[2]));
	jspl3 jspl3_w_asqrt51_37(.douta(w_asqrt51_37[0]),.doutb(w_asqrt51_37[1]),.doutc(w_asqrt51_37[2]),.din(w_asqrt51_12[0]));
	jspl3 jspl3_w_asqrt51_38(.douta(w_asqrt51_38[0]),.doutb(w_asqrt51_38[1]),.doutc(asqrt[50]),.din(w_asqrt51_12[1]));
	jspl3 jspl3_w_asqrt52_0(.douta(w_asqrt52_0[0]),.doutb(w_asqrt52_0[1]),.doutc(w_asqrt52_0[2]),.din(asqrt_fa_52));
	jspl3 jspl3_w_asqrt52_1(.douta(w_asqrt52_1[0]),.doutb(w_asqrt52_1[1]),.doutc(w_asqrt52_1[2]),.din(w_asqrt52_0[0]));
	jspl3 jspl3_w_asqrt52_2(.douta(w_asqrt52_2[0]),.doutb(w_asqrt52_2[1]),.doutc(w_asqrt52_2[2]),.din(w_asqrt52_0[1]));
	jspl3 jspl3_w_asqrt52_3(.douta(w_asqrt52_3[0]),.doutb(w_asqrt52_3[1]),.doutc(w_asqrt52_3[2]),.din(w_asqrt52_0[2]));
	jspl3 jspl3_w_asqrt52_4(.douta(w_asqrt52_4[0]),.doutb(w_asqrt52_4[1]),.doutc(w_asqrt52_4[2]),.din(w_asqrt52_1[0]));
	jspl3 jspl3_w_asqrt52_5(.douta(w_asqrt52_5[0]),.doutb(w_asqrt52_5[1]),.doutc(w_asqrt52_5[2]),.din(w_asqrt52_1[1]));
	jspl3 jspl3_w_asqrt52_6(.douta(w_asqrt52_6[0]),.doutb(w_asqrt52_6[1]),.doutc(w_asqrt52_6[2]),.din(w_asqrt52_1[2]));
	jspl3 jspl3_w_asqrt52_7(.douta(w_asqrt52_7[0]),.doutb(w_asqrt52_7[1]),.doutc(w_asqrt52_7[2]),.din(w_asqrt52_2[0]));
	jspl3 jspl3_w_asqrt52_8(.douta(w_asqrt52_8[0]),.doutb(w_asqrt52_8[1]),.doutc(w_asqrt52_8[2]),.din(w_asqrt52_2[1]));
	jspl3 jspl3_w_asqrt52_9(.douta(w_asqrt52_9[0]),.doutb(w_asqrt52_9[1]),.doutc(w_asqrt52_9[2]),.din(w_asqrt52_2[2]));
	jspl3 jspl3_w_asqrt52_10(.douta(w_asqrt52_10[0]),.doutb(w_asqrt52_10[1]),.doutc(w_asqrt52_10[2]),.din(w_asqrt52_3[0]));
	jspl3 jspl3_w_asqrt52_11(.douta(w_asqrt52_11[0]),.doutb(w_asqrt52_11[1]),.doutc(w_asqrt52_11[2]),.din(w_asqrt52_3[1]));
	jspl3 jspl3_w_asqrt52_12(.douta(w_asqrt52_12[0]),.doutb(w_asqrt52_12[1]),.doutc(w_asqrt52_12[2]),.din(w_asqrt52_3[2]));
	jspl3 jspl3_w_asqrt52_13(.douta(w_asqrt52_13[0]),.doutb(w_asqrt52_13[1]),.doutc(w_asqrt52_13[2]),.din(w_asqrt52_4[0]));
	jspl3 jspl3_w_asqrt52_14(.douta(w_asqrt52_14[0]),.doutb(w_asqrt52_14[1]),.doutc(w_asqrt52_14[2]),.din(w_asqrt52_4[1]));
	jspl3 jspl3_w_asqrt52_15(.douta(w_asqrt52_15[0]),.doutb(w_asqrt52_15[1]),.doutc(w_asqrt52_15[2]),.din(w_asqrt52_4[2]));
	jspl3 jspl3_w_asqrt52_16(.douta(w_asqrt52_16[0]),.doutb(w_asqrt52_16[1]),.doutc(w_asqrt52_16[2]),.din(w_asqrt52_5[0]));
	jspl3 jspl3_w_asqrt52_17(.douta(w_asqrt52_17[0]),.doutb(w_asqrt52_17[1]),.doutc(w_asqrt52_17[2]),.din(w_asqrt52_5[1]));
	jspl3 jspl3_w_asqrt52_18(.douta(w_asqrt52_18[0]),.doutb(w_asqrt52_18[1]),.doutc(w_asqrt52_18[2]),.din(w_asqrt52_5[2]));
	jspl3 jspl3_w_asqrt52_19(.douta(w_asqrt52_19[0]),.doutb(w_asqrt52_19[1]),.doutc(w_asqrt52_19[2]),.din(w_asqrt52_6[0]));
	jspl3 jspl3_w_asqrt52_20(.douta(w_asqrt52_20[0]),.doutb(w_asqrt52_20[1]),.doutc(w_asqrt52_20[2]),.din(w_asqrt52_6[1]));
	jspl3 jspl3_w_asqrt52_21(.douta(w_asqrt52_21[0]),.doutb(w_asqrt52_21[1]),.doutc(w_asqrt52_21[2]),.din(w_asqrt52_6[2]));
	jspl3 jspl3_w_asqrt52_22(.douta(w_asqrt52_22[0]),.doutb(w_asqrt52_22[1]),.doutc(w_asqrt52_22[2]),.din(w_asqrt52_7[0]));
	jspl3 jspl3_w_asqrt52_23(.douta(w_asqrt52_23[0]),.doutb(w_asqrt52_23[1]),.doutc(w_asqrt52_23[2]),.din(w_asqrt52_7[1]));
	jspl3 jspl3_w_asqrt52_24(.douta(w_asqrt52_24[0]),.doutb(w_asqrt52_24[1]),.doutc(w_asqrt52_24[2]),.din(w_asqrt52_7[2]));
	jspl3 jspl3_w_asqrt52_25(.douta(w_asqrt52_25[0]),.doutb(w_asqrt52_25[1]),.doutc(w_asqrt52_25[2]),.din(w_asqrt52_8[0]));
	jspl3 jspl3_w_asqrt52_26(.douta(w_asqrt52_26[0]),.doutb(w_asqrt52_26[1]),.doutc(w_asqrt52_26[2]),.din(w_asqrt52_8[1]));
	jspl3 jspl3_w_asqrt52_27(.douta(w_asqrt52_27[0]),.doutb(w_asqrt52_27[1]),.doutc(w_asqrt52_27[2]),.din(w_asqrt52_8[2]));
	jspl3 jspl3_w_asqrt52_28(.douta(w_asqrt52_28[0]),.doutb(w_asqrt52_28[1]),.doutc(w_asqrt52_28[2]),.din(w_asqrt52_9[0]));
	jspl3 jspl3_w_asqrt52_29(.douta(w_asqrt52_29[0]),.doutb(w_asqrt52_29[1]),.doutc(w_asqrt52_29[2]),.din(w_asqrt52_9[1]));
	jspl3 jspl3_w_asqrt52_30(.douta(w_asqrt52_30[0]),.doutb(w_asqrt52_30[1]),.doutc(w_asqrt52_30[2]),.din(w_asqrt52_9[2]));
	jspl3 jspl3_w_asqrt52_31(.douta(w_asqrt52_31[0]),.doutb(w_asqrt52_31[1]),.doutc(w_asqrt52_31[2]),.din(w_asqrt52_10[0]));
	jspl3 jspl3_w_asqrt52_32(.douta(w_asqrt52_32[0]),.doutb(w_asqrt52_32[1]),.doutc(w_asqrt52_32[2]),.din(w_asqrt52_10[1]));
	jspl3 jspl3_w_asqrt52_33(.douta(w_asqrt52_33[0]),.doutb(w_asqrt52_33[1]),.doutc(w_asqrt52_33[2]),.din(w_asqrt52_10[2]));
	jspl3 jspl3_w_asqrt52_34(.douta(w_asqrt52_34[0]),.doutb(w_asqrt52_34[1]),.doutc(w_asqrt52_34[2]),.din(w_asqrt52_11[0]));
	jspl3 jspl3_w_asqrt52_35(.douta(w_asqrt52_35[0]),.doutb(w_asqrt52_35[1]),.doutc(w_asqrt52_35[2]),.din(w_asqrt52_11[1]));
	jspl3 jspl3_w_asqrt52_36(.douta(w_asqrt52_36[0]),.doutb(w_asqrt52_36[1]),.doutc(w_asqrt52_36[2]),.din(w_asqrt52_11[2]));
	jspl3 jspl3_w_asqrt52_37(.douta(w_asqrt52_37[0]),.doutb(w_asqrt52_37[1]),.doutc(w_asqrt52_37[2]),.din(w_asqrt52_12[0]));
	jspl3 jspl3_w_asqrt52_38(.douta(w_asqrt52_38[0]),.doutb(w_asqrt52_38[1]),.doutc(w_asqrt52_38[2]),.din(w_asqrt52_12[1]));
	jspl3 jspl3_w_asqrt52_39(.douta(w_asqrt52_39[0]),.doutb(w_asqrt52_39[1]),.doutc(w_asqrt52_39[2]),.din(w_asqrt52_12[2]));
	jspl3 jspl3_w_asqrt52_40(.douta(w_asqrt52_40[0]),.doutb(w_asqrt52_40[1]),.doutc(w_asqrt52_40[2]),.din(w_asqrt52_13[0]));
	jspl3 jspl3_w_asqrt52_41(.douta(w_asqrt52_41[0]),.doutb(w_asqrt52_41[1]),.doutc(w_asqrt52_41[2]),.din(w_asqrt52_13[1]));
	jspl3 jspl3_w_asqrt52_42(.douta(w_asqrt52_42[0]),.doutb(w_asqrt52_42[1]),.doutc(w_asqrt52_42[2]),.din(w_asqrt52_13[2]));
	jspl3 jspl3_w_asqrt52_43(.douta(w_asqrt52_43[0]),.doutb(w_asqrt52_43[1]),.doutc(asqrt[51]),.din(w_asqrt52_14[0]));
	jspl3 jspl3_w_asqrt53_0(.douta(w_asqrt53_0[0]),.doutb(w_asqrt53_0[1]),.doutc(w_asqrt53_0[2]),.din(asqrt_fa_53));
	jspl3 jspl3_w_asqrt53_1(.douta(w_asqrt53_1[0]),.doutb(w_asqrt53_1[1]),.doutc(w_asqrt53_1[2]),.din(w_asqrt53_0[0]));
	jspl3 jspl3_w_asqrt53_2(.douta(w_asqrt53_2[0]),.doutb(w_asqrt53_2[1]),.doutc(w_asqrt53_2[2]),.din(w_asqrt53_0[1]));
	jspl3 jspl3_w_asqrt53_3(.douta(w_asqrt53_3[0]),.doutb(w_asqrt53_3[1]),.doutc(w_asqrt53_3[2]),.din(w_asqrt53_0[2]));
	jspl3 jspl3_w_asqrt53_4(.douta(w_asqrt53_4[0]),.doutb(w_asqrt53_4[1]),.doutc(w_asqrt53_4[2]),.din(w_asqrt53_1[0]));
	jspl3 jspl3_w_asqrt53_5(.douta(w_asqrt53_5[0]),.doutb(w_asqrt53_5[1]),.doutc(w_asqrt53_5[2]),.din(w_asqrt53_1[1]));
	jspl3 jspl3_w_asqrt53_6(.douta(w_asqrt53_6[0]),.doutb(w_asqrt53_6[1]),.doutc(w_asqrt53_6[2]),.din(w_asqrt53_1[2]));
	jspl3 jspl3_w_asqrt53_7(.douta(w_asqrt53_7[0]),.doutb(w_asqrt53_7[1]),.doutc(w_asqrt53_7[2]),.din(w_asqrt53_2[0]));
	jspl3 jspl3_w_asqrt53_8(.douta(w_asqrt53_8[0]),.doutb(w_asqrt53_8[1]),.doutc(w_asqrt53_8[2]),.din(w_asqrt53_2[1]));
	jspl3 jspl3_w_asqrt53_9(.douta(w_asqrt53_9[0]),.doutb(w_asqrt53_9[1]),.doutc(w_asqrt53_9[2]),.din(w_asqrt53_2[2]));
	jspl3 jspl3_w_asqrt53_10(.douta(w_asqrt53_10[0]),.doutb(w_asqrt53_10[1]),.doutc(w_asqrt53_10[2]),.din(w_asqrt53_3[0]));
	jspl3 jspl3_w_asqrt53_11(.douta(w_asqrt53_11[0]),.doutb(w_asqrt53_11[1]),.doutc(w_asqrt53_11[2]),.din(w_asqrt53_3[1]));
	jspl3 jspl3_w_asqrt53_12(.douta(w_asqrt53_12[0]),.doutb(w_asqrt53_12[1]),.doutc(w_asqrt53_12[2]),.din(w_asqrt53_3[2]));
	jspl3 jspl3_w_asqrt53_13(.douta(w_asqrt53_13[0]),.doutb(w_asqrt53_13[1]),.doutc(w_asqrt53_13[2]),.din(w_asqrt53_4[0]));
	jspl3 jspl3_w_asqrt53_14(.douta(w_asqrt53_14[0]),.doutb(w_asqrt53_14[1]),.doutc(w_asqrt53_14[2]),.din(w_asqrt53_4[1]));
	jspl3 jspl3_w_asqrt53_15(.douta(w_asqrt53_15[0]),.doutb(w_asqrt53_15[1]),.doutc(w_asqrt53_15[2]),.din(w_asqrt53_4[2]));
	jspl3 jspl3_w_asqrt53_16(.douta(w_asqrt53_16[0]),.doutb(w_asqrt53_16[1]),.doutc(w_asqrt53_16[2]),.din(w_asqrt53_5[0]));
	jspl3 jspl3_w_asqrt53_17(.douta(w_asqrt53_17[0]),.doutb(w_asqrt53_17[1]),.doutc(w_asqrt53_17[2]),.din(w_asqrt53_5[1]));
	jspl3 jspl3_w_asqrt53_18(.douta(w_asqrt53_18[0]),.doutb(w_asqrt53_18[1]),.doutc(w_asqrt53_18[2]),.din(w_asqrt53_5[2]));
	jspl3 jspl3_w_asqrt53_19(.douta(w_asqrt53_19[0]),.doutb(w_asqrt53_19[1]),.doutc(w_asqrt53_19[2]),.din(w_asqrt53_6[0]));
	jspl3 jspl3_w_asqrt53_20(.douta(w_asqrt53_20[0]),.doutb(w_asqrt53_20[1]),.doutc(w_asqrt53_20[2]),.din(w_asqrt53_6[1]));
	jspl3 jspl3_w_asqrt53_21(.douta(w_asqrt53_21[0]),.doutb(w_asqrt53_21[1]),.doutc(w_asqrt53_21[2]),.din(w_asqrt53_6[2]));
	jspl3 jspl3_w_asqrt53_22(.douta(w_asqrt53_22[0]),.doutb(w_asqrt53_22[1]),.doutc(w_asqrt53_22[2]),.din(w_asqrt53_7[0]));
	jspl3 jspl3_w_asqrt53_23(.douta(w_asqrt53_23[0]),.doutb(w_asqrt53_23[1]),.doutc(w_asqrt53_23[2]),.din(w_asqrt53_7[1]));
	jspl3 jspl3_w_asqrt53_24(.douta(w_asqrt53_24[0]),.doutb(w_asqrt53_24[1]),.doutc(w_asqrt53_24[2]),.din(w_asqrt53_7[2]));
	jspl3 jspl3_w_asqrt53_25(.douta(w_asqrt53_25[0]),.doutb(w_asqrt53_25[1]),.doutc(w_asqrt53_25[2]),.din(w_asqrt53_8[0]));
	jspl3 jspl3_w_asqrt53_26(.douta(w_asqrt53_26[0]),.doutb(w_asqrt53_26[1]),.doutc(w_asqrt53_26[2]),.din(w_asqrt53_8[1]));
	jspl3 jspl3_w_asqrt53_27(.douta(w_asqrt53_27[0]),.doutb(w_asqrt53_27[1]),.doutc(w_asqrt53_27[2]),.din(w_asqrt53_8[2]));
	jspl3 jspl3_w_asqrt53_28(.douta(w_asqrt53_28[0]),.doutb(w_asqrt53_28[1]),.doutc(w_asqrt53_28[2]),.din(w_asqrt53_9[0]));
	jspl3 jspl3_w_asqrt53_29(.douta(w_asqrt53_29[0]),.doutb(w_asqrt53_29[1]),.doutc(w_asqrt53_29[2]),.din(w_asqrt53_9[1]));
	jspl3 jspl3_w_asqrt53_30(.douta(w_asqrt53_30[0]),.doutb(w_asqrt53_30[1]),.doutc(w_asqrt53_30[2]),.din(w_asqrt53_9[2]));
	jspl3 jspl3_w_asqrt53_31(.douta(w_asqrt53_31[0]),.doutb(w_asqrt53_31[1]),.doutc(w_asqrt53_31[2]),.din(w_asqrt53_10[0]));
	jspl3 jspl3_w_asqrt53_32(.douta(w_asqrt53_32[0]),.doutb(w_asqrt53_32[1]),.doutc(w_asqrt53_32[2]),.din(w_asqrt53_10[1]));
	jspl3 jspl3_w_asqrt53_33(.douta(w_asqrt53_33[0]),.doutb(w_asqrt53_33[1]),.doutc(w_asqrt53_33[2]),.din(w_asqrt53_10[2]));
	jspl3 jspl3_w_asqrt53_34(.douta(w_asqrt53_34[0]),.doutb(w_asqrt53_34[1]),.doutc(w_asqrt53_34[2]),.din(w_asqrt53_11[0]));
	jspl3 jspl3_w_asqrt53_35(.douta(w_asqrt53_35[0]),.doutb(w_asqrt53_35[1]),.doutc(w_asqrt53_35[2]),.din(w_asqrt53_11[1]));
	jspl3 jspl3_w_asqrt53_36(.douta(w_asqrt53_36[0]),.doutb(w_asqrt53_36[1]),.doutc(w_asqrt53_36[2]),.din(w_asqrt53_11[2]));
	jspl3 jspl3_w_asqrt53_37(.douta(w_asqrt53_37[0]),.doutb(w_asqrt53_37[1]),.doutc(w_asqrt53_37[2]),.din(w_asqrt53_12[0]));
	jspl3 jspl3_w_asqrt53_38(.douta(w_asqrt53_38[0]),.doutb(w_asqrt53_38[1]),.doutc(w_asqrt53_38[2]),.din(w_asqrt53_12[1]));
	jspl3 jspl3_w_asqrt53_39(.douta(w_asqrt53_39[0]),.doutb(w_asqrt53_39[1]),.doutc(w_asqrt53_39[2]),.din(w_asqrt53_12[2]));
	jspl3 jspl3_w_asqrt53_40(.douta(w_asqrt53_40[0]),.doutb(w_asqrt53_40[1]),.doutc(asqrt[52]),.din(w_asqrt53_13[0]));
	jspl3 jspl3_w_asqrt54_0(.douta(w_asqrt54_0[0]),.doutb(w_asqrt54_0[1]),.doutc(w_asqrt54_0[2]),.din(asqrt_fa_54));
	jspl3 jspl3_w_asqrt54_1(.douta(w_asqrt54_1[0]),.doutb(w_asqrt54_1[1]),.doutc(w_asqrt54_1[2]),.din(w_asqrt54_0[0]));
	jspl3 jspl3_w_asqrt54_2(.douta(w_asqrt54_2[0]),.doutb(w_asqrt54_2[1]),.doutc(w_asqrt54_2[2]),.din(w_asqrt54_0[1]));
	jspl3 jspl3_w_asqrt54_3(.douta(w_asqrt54_3[0]),.doutb(w_asqrt54_3[1]),.doutc(w_asqrt54_3[2]),.din(w_asqrt54_0[2]));
	jspl3 jspl3_w_asqrt54_4(.douta(w_asqrt54_4[0]),.doutb(w_asqrt54_4[1]),.doutc(w_asqrt54_4[2]),.din(w_asqrt54_1[0]));
	jspl3 jspl3_w_asqrt54_5(.douta(w_asqrt54_5[0]),.doutb(w_asqrt54_5[1]),.doutc(w_asqrt54_5[2]),.din(w_asqrt54_1[1]));
	jspl3 jspl3_w_asqrt54_6(.douta(w_asqrt54_6[0]),.doutb(w_asqrt54_6[1]),.doutc(w_asqrt54_6[2]),.din(w_asqrt54_1[2]));
	jspl3 jspl3_w_asqrt54_7(.douta(w_asqrt54_7[0]),.doutb(w_asqrt54_7[1]),.doutc(w_asqrt54_7[2]),.din(w_asqrt54_2[0]));
	jspl3 jspl3_w_asqrt54_8(.douta(w_asqrt54_8[0]),.doutb(w_asqrt54_8[1]),.doutc(w_asqrt54_8[2]),.din(w_asqrt54_2[1]));
	jspl3 jspl3_w_asqrt54_9(.douta(w_asqrt54_9[0]),.doutb(w_asqrt54_9[1]),.doutc(w_asqrt54_9[2]),.din(w_asqrt54_2[2]));
	jspl3 jspl3_w_asqrt54_10(.douta(w_asqrt54_10[0]),.doutb(w_asqrt54_10[1]),.doutc(w_asqrt54_10[2]),.din(w_asqrt54_3[0]));
	jspl3 jspl3_w_asqrt54_11(.douta(w_asqrt54_11[0]),.doutb(w_asqrt54_11[1]),.doutc(w_asqrt54_11[2]),.din(w_asqrt54_3[1]));
	jspl3 jspl3_w_asqrt54_12(.douta(w_asqrt54_12[0]),.doutb(w_asqrt54_12[1]),.doutc(w_asqrt54_12[2]),.din(w_asqrt54_3[2]));
	jspl3 jspl3_w_asqrt54_13(.douta(w_asqrt54_13[0]),.doutb(w_asqrt54_13[1]),.doutc(w_asqrt54_13[2]),.din(w_asqrt54_4[0]));
	jspl3 jspl3_w_asqrt54_14(.douta(w_asqrt54_14[0]),.doutb(w_asqrt54_14[1]),.doutc(w_asqrt54_14[2]),.din(w_asqrt54_4[1]));
	jspl3 jspl3_w_asqrt54_15(.douta(w_asqrt54_15[0]),.doutb(w_asqrt54_15[1]),.doutc(w_asqrt54_15[2]),.din(w_asqrt54_4[2]));
	jspl3 jspl3_w_asqrt54_16(.douta(w_asqrt54_16[0]),.doutb(w_asqrt54_16[1]),.doutc(w_asqrt54_16[2]),.din(w_asqrt54_5[0]));
	jspl3 jspl3_w_asqrt54_17(.douta(w_asqrt54_17[0]),.doutb(w_asqrt54_17[1]),.doutc(w_asqrt54_17[2]),.din(w_asqrt54_5[1]));
	jspl3 jspl3_w_asqrt54_18(.douta(w_asqrt54_18[0]),.doutb(w_asqrt54_18[1]),.doutc(w_asqrt54_18[2]),.din(w_asqrt54_5[2]));
	jspl3 jspl3_w_asqrt54_19(.douta(w_asqrt54_19[0]),.doutb(w_asqrt54_19[1]),.doutc(w_asqrt54_19[2]),.din(w_asqrt54_6[0]));
	jspl3 jspl3_w_asqrt54_20(.douta(w_asqrt54_20[0]),.doutb(w_asqrt54_20[1]),.doutc(w_asqrt54_20[2]),.din(w_asqrt54_6[1]));
	jspl3 jspl3_w_asqrt54_21(.douta(w_asqrt54_21[0]),.doutb(w_asqrt54_21[1]),.doutc(w_asqrt54_21[2]),.din(w_asqrt54_6[2]));
	jspl3 jspl3_w_asqrt54_22(.douta(w_asqrt54_22[0]),.doutb(w_asqrt54_22[1]),.doutc(w_asqrt54_22[2]),.din(w_asqrt54_7[0]));
	jspl3 jspl3_w_asqrt54_23(.douta(w_asqrt54_23[0]),.doutb(w_asqrt54_23[1]),.doutc(w_asqrt54_23[2]),.din(w_asqrt54_7[1]));
	jspl3 jspl3_w_asqrt54_24(.douta(w_asqrt54_24[0]),.doutb(w_asqrt54_24[1]),.doutc(w_asqrt54_24[2]),.din(w_asqrt54_7[2]));
	jspl3 jspl3_w_asqrt54_25(.douta(w_asqrt54_25[0]),.doutb(w_asqrt54_25[1]),.doutc(w_asqrt54_25[2]),.din(w_asqrt54_8[0]));
	jspl3 jspl3_w_asqrt54_26(.douta(w_asqrt54_26[0]),.doutb(w_asqrt54_26[1]),.doutc(w_asqrt54_26[2]),.din(w_asqrt54_8[1]));
	jspl3 jspl3_w_asqrt54_27(.douta(w_asqrt54_27[0]),.doutb(w_asqrt54_27[1]),.doutc(w_asqrt54_27[2]),.din(w_asqrt54_8[2]));
	jspl3 jspl3_w_asqrt54_28(.douta(w_asqrt54_28[0]),.doutb(w_asqrt54_28[1]),.doutc(w_asqrt54_28[2]),.din(w_asqrt54_9[0]));
	jspl3 jspl3_w_asqrt54_29(.douta(w_asqrt54_29[0]),.doutb(w_asqrt54_29[1]),.doutc(w_asqrt54_29[2]),.din(w_asqrt54_9[1]));
	jspl3 jspl3_w_asqrt54_30(.douta(w_asqrt54_30[0]),.doutb(w_asqrt54_30[1]),.doutc(w_asqrt54_30[2]),.din(w_asqrt54_9[2]));
	jspl3 jspl3_w_asqrt54_31(.douta(w_asqrt54_31[0]),.doutb(w_asqrt54_31[1]),.doutc(w_asqrt54_31[2]),.din(w_asqrt54_10[0]));
	jspl3 jspl3_w_asqrt54_32(.douta(w_asqrt54_32[0]),.doutb(w_asqrt54_32[1]),.doutc(w_asqrt54_32[2]),.din(w_asqrt54_10[1]));
	jspl3 jspl3_w_asqrt54_33(.douta(w_asqrt54_33[0]),.doutb(w_asqrt54_33[1]),.doutc(w_asqrt54_33[2]),.din(w_asqrt54_10[2]));
	jspl3 jspl3_w_asqrt54_34(.douta(w_asqrt54_34[0]),.doutb(w_asqrt54_34[1]),.doutc(w_asqrt54_34[2]),.din(w_asqrt54_11[0]));
	jspl3 jspl3_w_asqrt54_35(.douta(w_asqrt54_35[0]),.doutb(w_asqrt54_35[1]),.doutc(w_asqrt54_35[2]),.din(w_asqrt54_11[1]));
	jspl3 jspl3_w_asqrt54_36(.douta(w_asqrt54_36[0]),.doutb(w_asqrt54_36[1]),.doutc(w_asqrt54_36[2]),.din(w_asqrt54_11[2]));
	jspl3 jspl3_w_asqrt54_37(.douta(w_asqrt54_37[0]),.doutb(w_asqrt54_37[1]),.doutc(w_asqrt54_37[2]),.din(w_asqrt54_12[0]));
	jspl3 jspl3_w_asqrt54_38(.douta(w_asqrt54_38[0]),.doutb(w_asqrt54_38[1]),.doutc(w_asqrt54_38[2]),.din(w_asqrt54_12[1]));
	jspl3 jspl3_w_asqrt54_39(.douta(w_asqrt54_39[0]),.doutb(w_asqrt54_39[1]),.doutc(w_asqrt54_39[2]),.din(w_asqrt54_12[2]));
	jspl3 jspl3_w_asqrt54_40(.douta(w_asqrt54_40[0]),.doutb(w_asqrt54_40[1]),.doutc(w_asqrt54_40[2]),.din(w_asqrt54_13[0]));
	jspl3 jspl3_w_asqrt54_41(.douta(w_asqrt54_41[0]),.doutb(w_asqrt54_41[1]),.doutc(w_asqrt54_41[2]),.din(w_asqrt54_13[1]));
	jspl3 jspl3_w_asqrt54_42(.douta(w_asqrt54_42[0]),.doutb(w_asqrt54_42[1]),.doutc(w_asqrt54_42[2]),.din(w_asqrt54_13[2]));
	jspl3 jspl3_w_asqrt54_43(.douta(w_asqrt54_43[0]),.doutb(w_asqrt54_43[1]),.doutc(asqrt[53]),.din(w_asqrt54_14[0]));
	jspl3 jspl3_w_asqrt55_0(.douta(w_asqrt55_0[0]),.doutb(w_asqrt55_0[1]),.doutc(w_asqrt55_0[2]),.din(asqrt_fa_55));
	jspl3 jspl3_w_asqrt55_1(.douta(w_asqrt55_1[0]),.doutb(w_asqrt55_1[1]),.doutc(w_asqrt55_1[2]),.din(w_asqrt55_0[0]));
	jspl3 jspl3_w_asqrt55_2(.douta(w_asqrt55_2[0]),.doutb(w_asqrt55_2[1]),.doutc(w_asqrt55_2[2]),.din(w_asqrt55_0[1]));
	jspl3 jspl3_w_asqrt55_3(.douta(w_asqrt55_3[0]),.doutb(w_asqrt55_3[1]),.doutc(w_asqrt55_3[2]),.din(w_asqrt55_0[2]));
	jspl3 jspl3_w_asqrt55_4(.douta(w_asqrt55_4[0]),.doutb(w_asqrt55_4[1]),.doutc(w_asqrt55_4[2]),.din(w_asqrt55_1[0]));
	jspl3 jspl3_w_asqrt55_5(.douta(w_asqrt55_5[0]),.doutb(w_asqrt55_5[1]),.doutc(w_asqrt55_5[2]),.din(w_asqrt55_1[1]));
	jspl3 jspl3_w_asqrt55_6(.douta(w_asqrt55_6[0]),.doutb(w_asqrt55_6[1]),.doutc(w_asqrt55_6[2]),.din(w_asqrt55_1[2]));
	jspl3 jspl3_w_asqrt55_7(.douta(w_asqrt55_7[0]),.doutb(w_asqrt55_7[1]),.doutc(w_asqrt55_7[2]),.din(w_asqrt55_2[0]));
	jspl3 jspl3_w_asqrt55_8(.douta(w_asqrt55_8[0]),.doutb(w_asqrt55_8[1]),.doutc(w_asqrt55_8[2]),.din(w_asqrt55_2[1]));
	jspl3 jspl3_w_asqrt55_9(.douta(w_asqrt55_9[0]),.doutb(w_asqrt55_9[1]),.doutc(w_asqrt55_9[2]),.din(w_asqrt55_2[2]));
	jspl3 jspl3_w_asqrt55_10(.douta(w_asqrt55_10[0]),.doutb(w_asqrt55_10[1]),.doutc(w_asqrt55_10[2]),.din(w_asqrt55_3[0]));
	jspl3 jspl3_w_asqrt55_11(.douta(w_asqrt55_11[0]),.doutb(w_asqrt55_11[1]),.doutc(w_asqrt55_11[2]),.din(w_asqrt55_3[1]));
	jspl3 jspl3_w_asqrt55_12(.douta(w_asqrt55_12[0]),.doutb(w_asqrt55_12[1]),.doutc(w_asqrt55_12[2]),.din(w_asqrt55_3[2]));
	jspl3 jspl3_w_asqrt55_13(.douta(w_asqrt55_13[0]),.doutb(w_asqrt55_13[1]),.doutc(w_asqrt55_13[2]),.din(w_asqrt55_4[0]));
	jspl3 jspl3_w_asqrt55_14(.douta(w_asqrt55_14[0]),.doutb(w_asqrt55_14[1]),.doutc(w_asqrt55_14[2]),.din(w_asqrt55_4[1]));
	jspl3 jspl3_w_asqrt55_15(.douta(w_asqrt55_15[0]),.doutb(w_asqrt55_15[1]),.doutc(w_asqrt55_15[2]),.din(w_asqrt55_4[2]));
	jspl3 jspl3_w_asqrt55_16(.douta(w_asqrt55_16[0]),.doutb(w_asqrt55_16[1]),.doutc(w_asqrt55_16[2]),.din(w_asqrt55_5[0]));
	jspl3 jspl3_w_asqrt55_17(.douta(w_asqrt55_17[0]),.doutb(w_asqrt55_17[1]),.doutc(w_asqrt55_17[2]),.din(w_asqrt55_5[1]));
	jspl3 jspl3_w_asqrt55_18(.douta(w_asqrt55_18[0]),.doutb(w_asqrt55_18[1]),.doutc(w_asqrt55_18[2]),.din(w_asqrt55_5[2]));
	jspl3 jspl3_w_asqrt55_19(.douta(w_asqrt55_19[0]),.doutb(w_asqrt55_19[1]),.doutc(w_asqrt55_19[2]),.din(w_asqrt55_6[0]));
	jspl3 jspl3_w_asqrt55_20(.douta(w_asqrt55_20[0]),.doutb(w_asqrt55_20[1]),.doutc(w_asqrt55_20[2]),.din(w_asqrt55_6[1]));
	jspl3 jspl3_w_asqrt55_21(.douta(w_asqrt55_21[0]),.doutb(w_asqrt55_21[1]),.doutc(w_asqrt55_21[2]),.din(w_asqrt55_6[2]));
	jspl3 jspl3_w_asqrt55_22(.douta(w_asqrt55_22[0]),.doutb(w_asqrt55_22[1]),.doutc(w_asqrt55_22[2]),.din(w_asqrt55_7[0]));
	jspl3 jspl3_w_asqrt55_23(.douta(w_asqrt55_23[0]),.doutb(w_asqrt55_23[1]),.doutc(w_asqrt55_23[2]),.din(w_asqrt55_7[1]));
	jspl3 jspl3_w_asqrt55_24(.douta(w_asqrt55_24[0]),.doutb(w_asqrt55_24[1]),.doutc(w_asqrt55_24[2]),.din(w_asqrt55_7[2]));
	jspl3 jspl3_w_asqrt55_25(.douta(w_asqrt55_25[0]),.doutb(w_asqrt55_25[1]),.doutc(w_asqrt55_25[2]),.din(w_asqrt55_8[0]));
	jspl3 jspl3_w_asqrt55_26(.douta(w_asqrt55_26[0]),.doutb(w_asqrt55_26[1]),.doutc(w_asqrt55_26[2]),.din(w_asqrt55_8[1]));
	jspl3 jspl3_w_asqrt55_27(.douta(w_asqrt55_27[0]),.doutb(w_asqrt55_27[1]),.doutc(w_asqrt55_27[2]),.din(w_asqrt55_8[2]));
	jspl3 jspl3_w_asqrt55_28(.douta(w_asqrt55_28[0]),.doutb(w_asqrt55_28[1]),.doutc(w_asqrt55_28[2]),.din(w_asqrt55_9[0]));
	jspl3 jspl3_w_asqrt55_29(.douta(w_asqrt55_29[0]),.doutb(w_asqrt55_29[1]),.doutc(w_asqrt55_29[2]),.din(w_asqrt55_9[1]));
	jspl3 jspl3_w_asqrt55_30(.douta(w_asqrt55_30[0]),.doutb(w_asqrt55_30[1]),.doutc(w_asqrt55_30[2]),.din(w_asqrt55_9[2]));
	jspl3 jspl3_w_asqrt55_31(.douta(w_asqrt55_31[0]),.doutb(w_asqrt55_31[1]),.doutc(w_asqrt55_31[2]),.din(w_asqrt55_10[0]));
	jspl3 jspl3_w_asqrt55_32(.douta(w_asqrt55_32[0]),.doutb(w_asqrt55_32[1]),.doutc(w_asqrt55_32[2]),.din(w_asqrt55_10[1]));
	jspl3 jspl3_w_asqrt55_33(.douta(w_asqrt55_33[0]),.doutb(w_asqrt55_33[1]),.doutc(w_asqrt55_33[2]),.din(w_asqrt55_10[2]));
	jspl3 jspl3_w_asqrt55_34(.douta(w_asqrt55_34[0]),.doutb(w_asqrt55_34[1]),.doutc(w_asqrt55_34[2]),.din(w_asqrt55_11[0]));
	jspl3 jspl3_w_asqrt55_35(.douta(w_asqrt55_35[0]),.doutb(w_asqrt55_35[1]),.doutc(w_asqrt55_35[2]),.din(w_asqrt55_11[1]));
	jspl3 jspl3_w_asqrt55_36(.douta(w_asqrt55_36[0]),.doutb(w_asqrt55_36[1]),.doutc(w_asqrt55_36[2]),.din(w_asqrt55_11[2]));
	jspl3 jspl3_w_asqrt55_37(.douta(w_asqrt55_37[0]),.doutb(w_asqrt55_37[1]),.doutc(w_asqrt55_37[2]),.din(w_asqrt55_12[0]));
	jspl3 jspl3_w_asqrt55_38(.douta(w_asqrt55_38[0]),.doutb(w_asqrt55_38[1]),.doutc(w_asqrt55_38[2]),.din(w_asqrt55_12[1]));
	jspl3 jspl3_w_asqrt55_39(.douta(w_asqrt55_39[0]),.doutb(w_asqrt55_39[1]),.doutc(w_asqrt55_39[2]),.din(w_asqrt55_12[2]));
	jspl3 jspl3_w_asqrt55_40(.douta(w_asqrt55_40[0]),.doutb(w_asqrt55_40[1]),.doutc(w_asqrt55_40[2]),.din(w_asqrt55_13[0]));
	jspl3 jspl3_w_asqrt55_41(.douta(w_asqrt55_41[0]),.doutb(w_asqrt55_41[1]),.doutc(asqrt[54]),.din(w_asqrt55_13[1]));
	jspl3 jspl3_w_asqrt56_0(.douta(w_asqrt56_0[0]),.doutb(w_asqrt56_0[1]),.doutc(w_asqrt56_0[2]),.din(asqrt_fa_56));
	jspl3 jspl3_w_asqrt56_1(.douta(w_asqrt56_1[0]),.doutb(w_asqrt56_1[1]),.doutc(w_asqrt56_1[2]),.din(w_asqrt56_0[0]));
	jspl3 jspl3_w_asqrt56_2(.douta(w_asqrt56_2[0]),.doutb(w_asqrt56_2[1]),.doutc(w_asqrt56_2[2]),.din(w_asqrt56_0[1]));
	jspl3 jspl3_w_asqrt56_3(.douta(w_asqrt56_3[0]),.doutb(w_asqrt56_3[1]),.doutc(w_asqrt56_3[2]),.din(w_asqrt56_0[2]));
	jspl3 jspl3_w_asqrt56_4(.douta(w_asqrt56_4[0]),.doutb(w_asqrt56_4[1]),.doutc(w_asqrt56_4[2]),.din(w_asqrt56_1[0]));
	jspl3 jspl3_w_asqrt56_5(.douta(w_asqrt56_5[0]),.doutb(w_asqrt56_5[1]),.doutc(w_asqrt56_5[2]),.din(w_asqrt56_1[1]));
	jspl3 jspl3_w_asqrt56_6(.douta(w_asqrt56_6[0]),.doutb(w_asqrt56_6[1]),.doutc(w_asqrt56_6[2]),.din(w_asqrt56_1[2]));
	jspl3 jspl3_w_asqrt56_7(.douta(w_asqrt56_7[0]),.doutb(w_asqrt56_7[1]),.doutc(w_asqrt56_7[2]),.din(w_asqrt56_2[0]));
	jspl3 jspl3_w_asqrt56_8(.douta(w_asqrt56_8[0]),.doutb(w_asqrt56_8[1]),.doutc(w_asqrt56_8[2]),.din(w_asqrt56_2[1]));
	jspl3 jspl3_w_asqrt56_9(.douta(w_asqrt56_9[0]),.doutb(w_asqrt56_9[1]),.doutc(w_asqrt56_9[2]),.din(w_asqrt56_2[2]));
	jspl3 jspl3_w_asqrt56_10(.douta(w_asqrt56_10[0]),.doutb(w_asqrt56_10[1]),.doutc(w_asqrt56_10[2]),.din(w_asqrt56_3[0]));
	jspl3 jspl3_w_asqrt56_11(.douta(w_asqrt56_11[0]),.doutb(w_asqrt56_11[1]),.doutc(w_asqrt56_11[2]),.din(w_asqrt56_3[1]));
	jspl3 jspl3_w_asqrt56_12(.douta(w_asqrt56_12[0]),.doutb(w_asqrt56_12[1]),.doutc(w_asqrt56_12[2]),.din(w_asqrt56_3[2]));
	jspl3 jspl3_w_asqrt56_13(.douta(w_asqrt56_13[0]),.doutb(w_asqrt56_13[1]),.doutc(w_asqrt56_13[2]),.din(w_asqrt56_4[0]));
	jspl3 jspl3_w_asqrt56_14(.douta(w_asqrt56_14[0]),.doutb(w_asqrt56_14[1]),.doutc(w_asqrt56_14[2]),.din(w_asqrt56_4[1]));
	jspl3 jspl3_w_asqrt56_15(.douta(w_asqrt56_15[0]),.doutb(w_asqrt56_15[1]),.doutc(w_asqrt56_15[2]),.din(w_asqrt56_4[2]));
	jspl3 jspl3_w_asqrt56_16(.douta(w_asqrt56_16[0]),.doutb(w_asqrt56_16[1]),.doutc(w_asqrt56_16[2]),.din(w_asqrt56_5[0]));
	jspl3 jspl3_w_asqrt56_17(.douta(w_asqrt56_17[0]),.doutb(w_asqrt56_17[1]),.doutc(w_asqrt56_17[2]),.din(w_asqrt56_5[1]));
	jspl3 jspl3_w_asqrt56_18(.douta(w_asqrt56_18[0]),.doutb(w_asqrt56_18[1]),.doutc(w_asqrt56_18[2]),.din(w_asqrt56_5[2]));
	jspl3 jspl3_w_asqrt56_19(.douta(w_asqrt56_19[0]),.doutb(w_asqrt56_19[1]),.doutc(w_asqrt56_19[2]),.din(w_asqrt56_6[0]));
	jspl3 jspl3_w_asqrt56_20(.douta(w_asqrt56_20[0]),.doutb(w_asqrt56_20[1]),.doutc(w_asqrt56_20[2]),.din(w_asqrt56_6[1]));
	jspl3 jspl3_w_asqrt56_21(.douta(w_asqrt56_21[0]),.doutb(w_asqrt56_21[1]),.doutc(w_asqrt56_21[2]),.din(w_asqrt56_6[2]));
	jspl3 jspl3_w_asqrt56_22(.douta(w_asqrt56_22[0]),.doutb(w_asqrt56_22[1]),.doutc(w_asqrt56_22[2]),.din(w_asqrt56_7[0]));
	jspl3 jspl3_w_asqrt56_23(.douta(w_asqrt56_23[0]),.doutb(w_asqrt56_23[1]),.doutc(w_asqrt56_23[2]),.din(w_asqrt56_7[1]));
	jspl3 jspl3_w_asqrt56_24(.douta(w_asqrt56_24[0]),.doutb(w_asqrt56_24[1]),.doutc(w_asqrt56_24[2]),.din(w_asqrt56_7[2]));
	jspl3 jspl3_w_asqrt56_25(.douta(w_asqrt56_25[0]),.doutb(w_asqrt56_25[1]),.doutc(w_asqrt56_25[2]),.din(w_asqrt56_8[0]));
	jspl3 jspl3_w_asqrt56_26(.douta(w_asqrt56_26[0]),.doutb(w_asqrt56_26[1]),.doutc(w_asqrt56_26[2]),.din(w_asqrt56_8[1]));
	jspl3 jspl3_w_asqrt56_27(.douta(w_asqrt56_27[0]),.doutb(w_asqrt56_27[1]),.doutc(w_asqrt56_27[2]),.din(w_asqrt56_8[2]));
	jspl3 jspl3_w_asqrt56_28(.douta(w_asqrt56_28[0]),.doutb(w_asqrt56_28[1]),.doutc(w_asqrt56_28[2]),.din(w_asqrt56_9[0]));
	jspl3 jspl3_w_asqrt56_29(.douta(w_asqrt56_29[0]),.doutb(w_asqrt56_29[1]),.doutc(w_asqrt56_29[2]),.din(w_asqrt56_9[1]));
	jspl3 jspl3_w_asqrt56_30(.douta(w_asqrt56_30[0]),.doutb(w_asqrt56_30[1]),.doutc(w_asqrt56_30[2]),.din(w_asqrt56_9[2]));
	jspl3 jspl3_w_asqrt56_31(.douta(w_asqrt56_31[0]),.doutb(w_asqrt56_31[1]),.doutc(w_asqrt56_31[2]),.din(w_asqrt56_10[0]));
	jspl3 jspl3_w_asqrt56_32(.douta(w_asqrt56_32[0]),.doutb(w_asqrt56_32[1]),.doutc(w_asqrt56_32[2]),.din(w_asqrt56_10[1]));
	jspl3 jspl3_w_asqrt56_33(.douta(w_asqrt56_33[0]),.doutb(w_asqrt56_33[1]),.doutc(w_asqrt56_33[2]),.din(w_asqrt56_10[2]));
	jspl3 jspl3_w_asqrt56_34(.douta(w_asqrt56_34[0]),.doutb(w_asqrt56_34[1]),.doutc(w_asqrt56_34[2]),.din(w_asqrt56_11[0]));
	jspl3 jspl3_w_asqrt56_35(.douta(w_asqrt56_35[0]),.doutb(w_asqrt56_35[1]),.doutc(w_asqrt56_35[2]),.din(w_asqrt56_11[1]));
	jspl3 jspl3_w_asqrt56_36(.douta(w_asqrt56_36[0]),.doutb(w_asqrt56_36[1]),.doutc(w_asqrt56_36[2]),.din(w_asqrt56_11[2]));
	jspl3 jspl3_w_asqrt56_37(.douta(w_asqrt56_37[0]),.doutb(w_asqrt56_37[1]),.doutc(w_asqrt56_37[2]),.din(w_asqrt56_12[0]));
	jspl3 jspl3_w_asqrt56_38(.douta(w_asqrt56_38[0]),.doutb(w_asqrt56_38[1]),.doutc(w_asqrt56_38[2]),.din(w_asqrt56_12[1]));
	jspl3 jspl3_w_asqrt56_39(.douta(w_asqrt56_39[0]),.doutb(w_asqrt56_39[1]),.doutc(w_asqrt56_39[2]),.din(w_asqrt56_12[2]));
	jspl3 jspl3_w_asqrt56_40(.douta(w_asqrt56_40[0]),.doutb(w_asqrt56_40[1]),.doutc(w_asqrt56_40[2]),.din(w_asqrt56_13[0]));
	jspl3 jspl3_w_asqrt56_41(.douta(w_asqrt56_41[0]),.doutb(w_asqrt56_41[1]),.doutc(w_asqrt56_41[2]),.din(w_asqrt56_13[1]));
	jspl3 jspl3_w_asqrt56_42(.douta(w_asqrt56_42[0]),.doutb(w_asqrt56_42[1]),.doutc(w_asqrt56_42[2]),.din(w_asqrt56_13[2]));
	jspl3 jspl3_w_asqrt56_43(.douta(w_asqrt56_43[0]),.doutb(w_asqrt56_43[1]),.doutc(w_asqrt56_43[2]),.din(w_asqrt56_14[0]));
	jspl3 jspl3_w_asqrt56_44(.douta(w_asqrt56_44[0]),.doutb(w_asqrt56_44[1]),.doutc(asqrt[55]),.din(w_asqrt56_14[1]));
	jspl3 jspl3_w_asqrt57_0(.douta(w_asqrt57_0[0]),.doutb(w_asqrt57_0[1]),.doutc(w_asqrt57_0[2]),.din(asqrt_fa_57));
	jspl3 jspl3_w_asqrt57_1(.douta(w_asqrt57_1[0]),.doutb(w_asqrt57_1[1]),.doutc(w_asqrt57_1[2]),.din(w_asqrt57_0[0]));
	jspl3 jspl3_w_asqrt57_2(.douta(w_asqrt57_2[0]),.doutb(w_asqrt57_2[1]),.doutc(w_asqrt57_2[2]),.din(w_asqrt57_0[1]));
	jspl3 jspl3_w_asqrt57_3(.douta(w_asqrt57_3[0]),.doutb(w_asqrt57_3[1]),.doutc(w_asqrt57_3[2]),.din(w_asqrt57_0[2]));
	jspl3 jspl3_w_asqrt57_4(.douta(w_asqrt57_4[0]),.doutb(w_asqrt57_4[1]),.doutc(w_asqrt57_4[2]),.din(w_asqrt57_1[0]));
	jspl3 jspl3_w_asqrt57_5(.douta(w_asqrt57_5[0]),.doutb(w_asqrt57_5[1]),.doutc(w_asqrt57_5[2]),.din(w_asqrt57_1[1]));
	jspl3 jspl3_w_asqrt57_6(.douta(w_asqrt57_6[0]),.doutb(w_asqrt57_6[1]),.doutc(w_asqrt57_6[2]),.din(w_asqrt57_1[2]));
	jspl3 jspl3_w_asqrt57_7(.douta(w_asqrt57_7[0]),.doutb(w_asqrt57_7[1]),.doutc(w_asqrt57_7[2]),.din(w_asqrt57_2[0]));
	jspl3 jspl3_w_asqrt57_8(.douta(w_asqrt57_8[0]),.doutb(w_asqrt57_8[1]),.doutc(w_asqrt57_8[2]),.din(w_asqrt57_2[1]));
	jspl3 jspl3_w_asqrt57_9(.douta(w_asqrt57_9[0]),.doutb(w_asqrt57_9[1]),.doutc(w_asqrt57_9[2]),.din(w_asqrt57_2[2]));
	jspl3 jspl3_w_asqrt57_10(.douta(w_asqrt57_10[0]),.doutb(w_asqrt57_10[1]),.doutc(w_asqrt57_10[2]),.din(w_asqrt57_3[0]));
	jspl3 jspl3_w_asqrt57_11(.douta(w_asqrt57_11[0]),.doutb(w_asqrt57_11[1]),.doutc(w_asqrt57_11[2]),.din(w_asqrt57_3[1]));
	jspl3 jspl3_w_asqrt57_12(.douta(w_asqrt57_12[0]),.doutb(w_asqrt57_12[1]),.doutc(w_asqrt57_12[2]),.din(w_asqrt57_3[2]));
	jspl3 jspl3_w_asqrt57_13(.douta(w_asqrt57_13[0]),.doutb(w_asqrt57_13[1]),.doutc(w_asqrt57_13[2]),.din(w_asqrt57_4[0]));
	jspl3 jspl3_w_asqrt57_14(.douta(w_asqrt57_14[0]),.doutb(w_asqrt57_14[1]),.doutc(w_asqrt57_14[2]),.din(w_asqrt57_4[1]));
	jspl3 jspl3_w_asqrt57_15(.douta(w_asqrt57_15[0]),.doutb(w_asqrt57_15[1]),.doutc(w_asqrt57_15[2]),.din(w_asqrt57_4[2]));
	jspl3 jspl3_w_asqrt57_16(.douta(w_asqrt57_16[0]),.doutb(w_asqrt57_16[1]),.doutc(w_asqrt57_16[2]),.din(w_asqrt57_5[0]));
	jspl3 jspl3_w_asqrt57_17(.douta(w_asqrt57_17[0]),.doutb(w_asqrt57_17[1]),.doutc(w_asqrt57_17[2]),.din(w_asqrt57_5[1]));
	jspl3 jspl3_w_asqrt57_18(.douta(w_asqrt57_18[0]),.doutb(w_asqrt57_18[1]),.doutc(w_asqrt57_18[2]),.din(w_asqrt57_5[2]));
	jspl3 jspl3_w_asqrt57_19(.douta(w_asqrt57_19[0]),.doutb(w_asqrt57_19[1]),.doutc(w_asqrt57_19[2]),.din(w_asqrt57_6[0]));
	jspl3 jspl3_w_asqrt57_20(.douta(w_asqrt57_20[0]),.doutb(w_asqrt57_20[1]),.doutc(w_asqrt57_20[2]),.din(w_asqrt57_6[1]));
	jspl3 jspl3_w_asqrt57_21(.douta(w_asqrt57_21[0]),.doutb(w_asqrt57_21[1]),.doutc(w_asqrt57_21[2]),.din(w_asqrt57_6[2]));
	jspl3 jspl3_w_asqrt57_22(.douta(w_asqrt57_22[0]),.doutb(w_asqrt57_22[1]),.doutc(w_asqrt57_22[2]),.din(w_asqrt57_7[0]));
	jspl3 jspl3_w_asqrt57_23(.douta(w_asqrt57_23[0]),.doutb(w_asqrt57_23[1]),.doutc(w_asqrt57_23[2]),.din(w_asqrt57_7[1]));
	jspl3 jspl3_w_asqrt57_24(.douta(w_asqrt57_24[0]),.doutb(w_asqrt57_24[1]),.doutc(w_asqrt57_24[2]),.din(w_asqrt57_7[2]));
	jspl3 jspl3_w_asqrt57_25(.douta(w_asqrt57_25[0]),.doutb(w_asqrt57_25[1]),.doutc(w_asqrt57_25[2]),.din(w_asqrt57_8[0]));
	jspl3 jspl3_w_asqrt57_26(.douta(w_asqrt57_26[0]),.doutb(w_asqrt57_26[1]),.doutc(w_asqrt57_26[2]),.din(w_asqrt57_8[1]));
	jspl3 jspl3_w_asqrt57_27(.douta(w_asqrt57_27[0]),.doutb(w_asqrt57_27[1]),.doutc(w_asqrt57_27[2]),.din(w_asqrt57_8[2]));
	jspl3 jspl3_w_asqrt57_28(.douta(w_asqrt57_28[0]),.doutb(w_asqrt57_28[1]),.doutc(w_asqrt57_28[2]),.din(w_asqrt57_9[0]));
	jspl3 jspl3_w_asqrt57_29(.douta(w_asqrt57_29[0]),.doutb(w_asqrt57_29[1]),.doutc(w_asqrt57_29[2]),.din(w_asqrt57_9[1]));
	jspl3 jspl3_w_asqrt57_30(.douta(w_asqrt57_30[0]),.doutb(w_asqrt57_30[1]),.doutc(w_asqrt57_30[2]),.din(w_asqrt57_9[2]));
	jspl3 jspl3_w_asqrt57_31(.douta(w_asqrt57_31[0]),.doutb(w_asqrt57_31[1]),.doutc(w_asqrt57_31[2]),.din(w_asqrt57_10[0]));
	jspl3 jspl3_w_asqrt57_32(.douta(w_asqrt57_32[0]),.doutb(w_asqrt57_32[1]),.doutc(w_asqrt57_32[2]),.din(w_asqrt57_10[1]));
	jspl3 jspl3_w_asqrt57_33(.douta(w_asqrt57_33[0]),.doutb(w_asqrt57_33[1]),.doutc(w_asqrt57_33[2]),.din(w_asqrt57_10[2]));
	jspl3 jspl3_w_asqrt57_34(.douta(w_asqrt57_34[0]),.doutb(w_asqrt57_34[1]),.doutc(w_asqrt57_34[2]),.din(w_asqrt57_11[0]));
	jspl3 jspl3_w_asqrt57_35(.douta(w_asqrt57_35[0]),.doutb(w_asqrt57_35[1]),.doutc(w_asqrt57_35[2]),.din(w_asqrt57_11[1]));
	jspl3 jspl3_w_asqrt57_36(.douta(w_asqrt57_36[0]),.doutb(w_asqrt57_36[1]),.doutc(w_asqrt57_36[2]),.din(w_asqrt57_11[2]));
	jspl3 jspl3_w_asqrt57_37(.douta(w_asqrt57_37[0]),.doutb(w_asqrt57_37[1]),.doutc(w_asqrt57_37[2]),.din(w_asqrt57_12[0]));
	jspl3 jspl3_w_asqrt57_38(.douta(w_asqrt57_38[0]),.doutb(w_asqrt57_38[1]),.doutc(w_asqrt57_38[2]),.din(w_asqrt57_12[1]));
	jspl3 jspl3_w_asqrt57_39(.douta(w_asqrt57_39[0]),.doutb(w_asqrt57_39[1]),.doutc(w_asqrt57_39[2]),.din(w_asqrt57_12[2]));
	jspl3 jspl3_w_asqrt57_40(.douta(w_asqrt57_40[0]),.doutb(w_asqrt57_40[1]),.doutc(w_asqrt57_40[2]),.din(w_asqrt57_13[0]));
	jspl3 jspl3_w_asqrt57_41(.douta(w_asqrt57_41[0]),.doutb(w_asqrt57_41[1]),.doutc(w_asqrt57_41[2]),.din(w_asqrt57_13[1]));
	jspl3 jspl3_w_asqrt57_42(.douta(w_asqrt57_42[0]),.doutb(w_asqrt57_42[1]),.doutc(w_asqrt57_42[2]),.din(w_asqrt57_13[2]));
	jspl3 jspl3_w_asqrt57_43(.douta(w_asqrt57_43[0]),.doutb(w_asqrt57_43[1]),.doutc(asqrt[56]),.din(w_asqrt57_14[0]));
	jspl3 jspl3_w_asqrt58_0(.douta(w_asqrt58_0[0]),.doutb(w_asqrt58_0[1]),.doutc(w_asqrt58_0[2]),.din(asqrt_fa_58));
	jspl3 jspl3_w_asqrt58_1(.douta(w_asqrt58_1[0]),.doutb(w_asqrt58_1[1]),.doutc(w_asqrt58_1[2]),.din(w_asqrt58_0[0]));
	jspl3 jspl3_w_asqrt58_2(.douta(w_asqrt58_2[0]),.doutb(w_asqrt58_2[1]),.doutc(w_asqrt58_2[2]),.din(w_asqrt58_0[1]));
	jspl3 jspl3_w_asqrt58_3(.douta(w_asqrt58_3[0]),.doutb(w_asqrt58_3[1]),.doutc(w_asqrt58_3[2]),.din(w_asqrt58_0[2]));
	jspl3 jspl3_w_asqrt58_4(.douta(w_asqrt58_4[0]),.doutb(w_asqrt58_4[1]),.doutc(w_asqrt58_4[2]),.din(w_asqrt58_1[0]));
	jspl3 jspl3_w_asqrt58_5(.douta(w_asqrt58_5[0]),.doutb(w_asqrt58_5[1]),.doutc(w_asqrt58_5[2]),.din(w_asqrt58_1[1]));
	jspl3 jspl3_w_asqrt58_6(.douta(w_asqrt58_6[0]),.doutb(w_asqrt58_6[1]),.doutc(w_asqrt58_6[2]),.din(w_asqrt58_1[2]));
	jspl3 jspl3_w_asqrt58_7(.douta(w_asqrt58_7[0]),.doutb(w_asqrt58_7[1]),.doutc(w_asqrt58_7[2]),.din(w_asqrt58_2[0]));
	jspl3 jspl3_w_asqrt58_8(.douta(w_asqrt58_8[0]),.doutb(w_asqrt58_8[1]),.doutc(w_asqrt58_8[2]),.din(w_asqrt58_2[1]));
	jspl3 jspl3_w_asqrt58_9(.douta(w_asqrt58_9[0]),.doutb(w_asqrt58_9[1]),.doutc(w_asqrt58_9[2]),.din(w_asqrt58_2[2]));
	jspl3 jspl3_w_asqrt58_10(.douta(w_asqrt58_10[0]),.doutb(w_asqrt58_10[1]),.doutc(w_asqrt58_10[2]),.din(w_asqrt58_3[0]));
	jspl3 jspl3_w_asqrt58_11(.douta(w_asqrt58_11[0]),.doutb(w_asqrt58_11[1]),.doutc(w_asqrt58_11[2]),.din(w_asqrt58_3[1]));
	jspl3 jspl3_w_asqrt58_12(.douta(w_asqrt58_12[0]),.doutb(w_asqrt58_12[1]),.doutc(w_asqrt58_12[2]),.din(w_asqrt58_3[2]));
	jspl3 jspl3_w_asqrt58_13(.douta(w_asqrt58_13[0]),.doutb(w_asqrt58_13[1]),.doutc(w_asqrt58_13[2]),.din(w_asqrt58_4[0]));
	jspl3 jspl3_w_asqrt58_14(.douta(w_asqrt58_14[0]),.doutb(w_asqrt58_14[1]),.doutc(w_asqrt58_14[2]),.din(w_asqrt58_4[1]));
	jspl3 jspl3_w_asqrt58_15(.douta(w_asqrt58_15[0]),.doutb(w_asqrt58_15[1]),.doutc(w_asqrt58_15[2]),.din(w_asqrt58_4[2]));
	jspl3 jspl3_w_asqrt58_16(.douta(w_asqrt58_16[0]),.doutb(w_asqrt58_16[1]),.doutc(w_asqrt58_16[2]),.din(w_asqrt58_5[0]));
	jspl3 jspl3_w_asqrt58_17(.douta(w_asqrt58_17[0]),.doutb(w_asqrt58_17[1]),.doutc(w_asqrt58_17[2]),.din(w_asqrt58_5[1]));
	jspl3 jspl3_w_asqrt58_18(.douta(w_asqrt58_18[0]),.doutb(w_asqrt58_18[1]),.doutc(w_asqrt58_18[2]),.din(w_asqrt58_5[2]));
	jspl3 jspl3_w_asqrt58_19(.douta(w_asqrt58_19[0]),.doutb(w_asqrt58_19[1]),.doutc(w_asqrt58_19[2]),.din(w_asqrt58_6[0]));
	jspl3 jspl3_w_asqrt58_20(.douta(w_asqrt58_20[0]),.doutb(w_asqrt58_20[1]),.doutc(w_asqrt58_20[2]),.din(w_asqrt58_6[1]));
	jspl3 jspl3_w_asqrt58_21(.douta(w_asqrt58_21[0]),.doutb(w_asqrt58_21[1]),.doutc(w_asqrt58_21[2]),.din(w_asqrt58_6[2]));
	jspl3 jspl3_w_asqrt58_22(.douta(w_asqrt58_22[0]),.doutb(w_asqrt58_22[1]),.doutc(w_asqrt58_22[2]),.din(w_asqrt58_7[0]));
	jspl3 jspl3_w_asqrt58_23(.douta(w_asqrt58_23[0]),.doutb(w_asqrt58_23[1]),.doutc(w_asqrt58_23[2]),.din(w_asqrt58_7[1]));
	jspl3 jspl3_w_asqrt58_24(.douta(w_asqrt58_24[0]),.doutb(w_asqrt58_24[1]),.doutc(w_asqrt58_24[2]),.din(w_asqrt58_7[2]));
	jspl3 jspl3_w_asqrt58_25(.douta(w_asqrt58_25[0]),.doutb(w_asqrt58_25[1]),.doutc(w_asqrt58_25[2]),.din(w_asqrt58_8[0]));
	jspl3 jspl3_w_asqrt58_26(.douta(w_asqrt58_26[0]),.doutb(w_asqrt58_26[1]),.doutc(w_asqrt58_26[2]),.din(w_asqrt58_8[1]));
	jspl3 jspl3_w_asqrt58_27(.douta(w_asqrt58_27[0]),.doutb(w_asqrt58_27[1]),.doutc(w_asqrt58_27[2]),.din(w_asqrt58_8[2]));
	jspl3 jspl3_w_asqrt58_28(.douta(w_asqrt58_28[0]),.doutb(w_asqrt58_28[1]),.doutc(w_asqrt58_28[2]),.din(w_asqrt58_9[0]));
	jspl3 jspl3_w_asqrt58_29(.douta(w_asqrt58_29[0]),.doutb(w_asqrt58_29[1]),.doutc(w_asqrt58_29[2]),.din(w_asqrt58_9[1]));
	jspl3 jspl3_w_asqrt58_30(.douta(w_asqrt58_30[0]),.doutb(w_asqrt58_30[1]),.doutc(w_asqrt58_30[2]),.din(w_asqrt58_9[2]));
	jspl3 jspl3_w_asqrt58_31(.douta(w_asqrt58_31[0]),.doutb(w_asqrt58_31[1]),.doutc(w_asqrt58_31[2]),.din(w_asqrt58_10[0]));
	jspl3 jspl3_w_asqrt58_32(.douta(w_asqrt58_32[0]),.doutb(w_asqrt58_32[1]),.doutc(w_asqrt58_32[2]),.din(w_asqrt58_10[1]));
	jspl3 jspl3_w_asqrt58_33(.douta(w_asqrt58_33[0]),.doutb(w_asqrt58_33[1]),.doutc(w_asqrt58_33[2]),.din(w_asqrt58_10[2]));
	jspl3 jspl3_w_asqrt58_34(.douta(w_asqrt58_34[0]),.doutb(w_asqrt58_34[1]),.doutc(w_asqrt58_34[2]),.din(w_asqrt58_11[0]));
	jspl3 jspl3_w_asqrt58_35(.douta(w_asqrt58_35[0]),.doutb(w_asqrt58_35[1]),.doutc(w_asqrt58_35[2]),.din(w_asqrt58_11[1]));
	jspl3 jspl3_w_asqrt58_36(.douta(w_asqrt58_36[0]),.doutb(w_asqrt58_36[1]),.doutc(w_asqrt58_36[2]),.din(w_asqrt58_11[2]));
	jspl3 jspl3_w_asqrt58_37(.douta(w_asqrt58_37[0]),.doutb(w_asqrt58_37[1]),.doutc(w_asqrt58_37[2]),.din(w_asqrt58_12[0]));
	jspl3 jspl3_w_asqrt58_38(.douta(w_asqrt58_38[0]),.doutb(w_asqrt58_38[1]),.doutc(w_asqrt58_38[2]),.din(w_asqrt58_12[1]));
	jspl3 jspl3_w_asqrt58_39(.douta(w_asqrt58_39[0]),.doutb(w_asqrt58_39[1]),.doutc(w_asqrt58_39[2]),.din(w_asqrt58_12[2]));
	jspl3 jspl3_w_asqrt58_40(.douta(w_asqrt58_40[0]),.doutb(w_asqrt58_40[1]),.doutc(w_asqrt58_40[2]),.din(w_asqrt58_13[0]));
	jspl3 jspl3_w_asqrt58_41(.douta(w_asqrt58_41[0]),.doutb(w_asqrt58_41[1]),.doutc(w_asqrt58_41[2]),.din(w_asqrt58_13[1]));
	jspl3 jspl3_w_asqrt58_42(.douta(w_asqrt58_42[0]),.doutb(w_asqrt58_42[1]),.doutc(w_asqrt58_42[2]),.din(w_asqrt58_13[2]));
	jspl3 jspl3_w_asqrt58_43(.douta(w_asqrt58_43[0]),.doutb(w_asqrt58_43[1]),.doutc(w_asqrt58_43[2]),.din(w_asqrt58_14[0]));
	jspl3 jspl3_w_asqrt58_44(.douta(w_asqrt58_44[0]),.doutb(w_asqrt58_44[1]),.doutc(w_asqrt58_44[2]),.din(w_asqrt58_14[1]));
	jspl jspl_w_asqrt58_45(.douta(w_asqrt58_45),.doutb(asqrt[57]),.din(w_asqrt58_14[2]));
	jspl3 jspl3_w_asqrt59_0(.douta(w_asqrt59_0[0]),.doutb(w_asqrt59_0[1]),.doutc(w_asqrt59_0[2]),.din(asqrt_fa_59));
	jspl3 jspl3_w_asqrt59_1(.douta(w_asqrt59_1[0]),.doutb(w_asqrt59_1[1]),.doutc(w_asqrt59_1[2]),.din(w_asqrt59_0[0]));
	jspl3 jspl3_w_asqrt59_2(.douta(w_asqrt59_2[0]),.doutb(w_asqrt59_2[1]),.doutc(w_asqrt59_2[2]),.din(w_asqrt59_0[1]));
	jspl3 jspl3_w_asqrt59_3(.douta(w_asqrt59_3[0]),.doutb(w_asqrt59_3[1]),.doutc(w_asqrt59_3[2]),.din(w_asqrt59_0[2]));
	jspl3 jspl3_w_asqrt59_4(.douta(w_asqrt59_4[0]),.doutb(w_asqrt59_4[1]),.doutc(w_asqrt59_4[2]),.din(w_asqrt59_1[0]));
	jspl3 jspl3_w_asqrt59_5(.douta(w_asqrt59_5[0]),.doutb(w_asqrt59_5[1]),.doutc(w_asqrt59_5[2]),.din(w_asqrt59_1[1]));
	jspl3 jspl3_w_asqrt59_6(.douta(w_asqrt59_6[0]),.doutb(w_asqrt59_6[1]),.doutc(w_asqrt59_6[2]),.din(w_asqrt59_1[2]));
	jspl3 jspl3_w_asqrt59_7(.douta(w_asqrt59_7[0]),.doutb(w_asqrt59_7[1]),.doutc(w_asqrt59_7[2]),.din(w_asqrt59_2[0]));
	jspl3 jspl3_w_asqrt59_8(.douta(w_asqrt59_8[0]),.doutb(w_asqrt59_8[1]),.doutc(w_asqrt59_8[2]),.din(w_asqrt59_2[1]));
	jspl3 jspl3_w_asqrt59_9(.douta(w_asqrt59_9[0]),.doutb(w_asqrt59_9[1]),.doutc(w_asqrt59_9[2]),.din(w_asqrt59_2[2]));
	jspl3 jspl3_w_asqrt59_10(.douta(w_asqrt59_10[0]),.doutb(w_asqrt59_10[1]),.doutc(w_asqrt59_10[2]),.din(w_asqrt59_3[0]));
	jspl3 jspl3_w_asqrt59_11(.douta(w_asqrt59_11[0]),.doutb(w_asqrt59_11[1]),.doutc(w_asqrt59_11[2]),.din(w_asqrt59_3[1]));
	jspl3 jspl3_w_asqrt59_12(.douta(w_asqrt59_12[0]),.doutb(w_asqrt59_12[1]),.doutc(w_asqrt59_12[2]),.din(w_asqrt59_3[2]));
	jspl3 jspl3_w_asqrt59_13(.douta(w_asqrt59_13[0]),.doutb(w_asqrt59_13[1]),.doutc(w_asqrt59_13[2]),.din(w_asqrt59_4[0]));
	jspl3 jspl3_w_asqrt59_14(.douta(w_asqrt59_14[0]),.doutb(w_asqrt59_14[1]),.doutc(w_asqrt59_14[2]),.din(w_asqrt59_4[1]));
	jspl3 jspl3_w_asqrt59_15(.douta(w_asqrt59_15[0]),.doutb(w_asqrt59_15[1]),.doutc(w_asqrt59_15[2]),.din(w_asqrt59_4[2]));
	jspl3 jspl3_w_asqrt59_16(.douta(w_asqrt59_16[0]),.doutb(w_asqrt59_16[1]),.doutc(w_asqrt59_16[2]),.din(w_asqrt59_5[0]));
	jspl3 jspl3_w_asqrt59_17(.douta(w_asqrt59_17[0]),.doutb(w_asqrt59_17[1]),.doutc(w_asqrt59_17[2]),.din(w_asqrt59_5[1]));
	jspl3 jspl3_w_asqrt59_18(.douta(w_asqrt59_18[0]),.doutb(w_asqrt59_18[1]),.doutc(w_asqrt59_18[2]),.din(w_asqrt59_5[2]));
	jspl3 jspl3_w_asqrt59_19(.douta(w_asqrt59_19[0]),.doutb(w_asqrt59_19[1]),.doutc(w_asqrt59_19[2]),.din(w_asqrt59_6[0]));
	jspl3 jspl3_w_asqrt59_20(.douta(w_asqrt59_20[0]),.doutb(w_asqrt59_20[1]),.doutc(w_asqrt59_20[2]),.din(w_asqrt59_6[1]));
	jspl3 jspl3_w_asqrt59_21(.douta(w_asqrt59_21[0]),.doutb(w_asqrt59_21[1]),.doutc(w_asqrt59_21[2]),.din(w_asqrt59_6[2]));
	jspl3 jspl3_w_asqrt59_22(.douta(w_asqrt59_22[0]),.doutb(w_asqrt59_22[1]),.doutc(w_asqrt59_22[2]),.din(w_asqrt59_7[0]));
	jspl3 jspl3_w_asqrt59_23(.douta(w_asqrt59_23[0]),.doutb(w_asqrt59_23[1]),.doutc(w_asqrt59_23[2]),.din(w_asqrt59_7[1]));
	jspl3 jspl3_w_asqrt59_24(.douta(w_asqrt59_24[0]),.doutb(w_asqrt59_24[1]),.doutc(w_asqrt59_24[2]),.din(w_asqrt59_7[2]));
	jspl3 jspl3_w_asqrt59_25(.douta(w_asqrt59_25[0]),.doutb(w_asqrt59_25[1]),.doutc(w_asqrt59_25[2]),.din(w_asqrt59_8[0]));
	jspl3 jspl3_w_asqrt59_26(.douta(w_asqrt59_26[0]),.doutb(w_asqrt59_26[1]),.doutc(w_asqrt59_26[2]),.din(w_asqrt59_8[1]));
	jspl3 jspl3_w_asqrt59_27(.douta(w_asqrt59_27[0]),.doutb(w_asqrt59_27[1]),.doutc(w_asqrt59_27[2]),.din(w_asqrt59_8[2]));
	jspl3 jspl3_w_asqrt59_28(.douta(w_asqrt59_28[0]),.doutb(w_asqrt59_28[1]),.doutc(w_asqrt59_28[2]),.din(w_asqrt59_9[0]));
	jspl3 jspl3_w_asqrt59_29(.douta(w_asqrt59_29[0]),.doutb(w_asqrt59_29[1]),.doutc(w_asqrt59_29[2]),.din(w_asqrt59_9[1]));
	jspl3 jspl3_w_asqrt59_30(.douta(w_asqrt59_30[0]),.doutb(w_asqrt59_30[1]),.doutc(w_asqrt59_30[2]),.din(w_asqrt59_9[2]));
	jspl3 jspl3_w_asqrt59_31(.douta(w_asqrt59_31[0]),.doutb(w_asqrt59_31[1]),.doutc(w_asqrt59_31[2]),.din(w_asqrt59_10[0]));
	jspl3 jspl3_w_asqrt59_32(.douta(w_asqrt59_32[0]),.doutb(w_asqrt59_32[1]),.doutc(w_asqrt59_32[2]),.din(w_asqrt59_10[1]));
	jspl3 jspl3_w_asqrt59_33(.douta(w_asqrt59_33[0]),.doutb(w_asqrt59_33[1]),.doutc(w_asqrt59_33[2]),.din(w_asqrt59_10[2]));
	jspl3 jspl3_w_asqrt59_34(.douta(w_asqrt59_34[0]),.doutb(w_asqrt59_34[1]),.doutc(w_asqrt59_34[2]),.din(w_asqrt59_11[0]));
	jspl3 jspl3_w_asqrt59_35(.douta(w_asqrt59_35[0]),.doutb(w_asqrt59_35[1]),.doutc(w_asqrt59_35[2]),.din(w_asqrt59_11[1]));
	jspl3 jspl3_w_asqrt59_36(.douta(w_asqrt59_36[0]),.doutb(w_asqrt59_36[1]),.doutc(w_asqrt59_36[2]),.din(w_asqrt59_11[2]));
	jspl3 jspl3_w_asqrt59_37(.douta(w_asqrt59_37[0]),.doutb(w_asqrt59_37[1]),.doutc(w_asqrt59_37[2]),.din(w_asqrt59_12[0]));
	jspl3 jspl3_w_asqrt59_38(.douta(w_asqrt59_38[0]),.doutb(w_asqrt59_38[1]),.doutc(w_asqrt59_38[2]),.din(w_asqrt59_12[1]));
	jspl3 jspl3_w_asqrt59_39(.douta(w_asqrt59_39[0]),.doutb(w_asqrt59_39[1]),.doutc(w_asqrt59_39[2]),.din(w_asqrt59_12[2]));
	jspl3 jspl3_w_asqrt59_40(.douta(w_asqrt59_40[0]),.doutb(w_asqrt59_40[1]),.doutc(w_asqrt59_40[2]),.din(w_asqrt59_13[0]));
	jspl3 jspl3_w_asqrt59_41(.douta(w_asqrt59_41[0]),.doutb(w_asqrt59_41[1]),.doutc(w_asqrt59_41[2]),.din(w_asqrt59_13[1]));
	jspl3 jspl3_w_asqrt59_42(.douta(w_asqrt59_42[0]),.doutb(w_asqrt59_42[1]),.doutc(w_asqrt59_42[2]),.din(w_asqrt59_13[2]));
	jspl3 jspl3_w_asqrt59_43(.douta(w_asqrt59_43[0]),.doutb(w_asqrt59_43[1]),.doutc(w_asqrt59_43[2]),.din(w_asqrt59_14[0]));
	jspl3 jspl3_w_asqrt59_44(.douta(w_asqrt59_44[0]),.doutb(w_asqrt59_44[1]),.doutc(asqrt[58]),.din(w_asqrt59_14[1]));
	jspl3 jspl3_w_asqrt60_0(.douta(w_asqrt60_0[0]),.doutb(w_asqrt60_0[1]),.doutc(w_asqrt60_0[2]),.din(asqrt_fa_60));
	jspl3 jspl3_w_asqrt60_1(.douta(w_asqrt60_1[0]),.doutb(w_asqrt60_1[1]),.doutc(w_asqrt60_1[2]),.din(w_asqrt60_0[0]));
	jspl3 jspl3_w_asqrt60_2(.douta(w_asqrt60_2[0]),.doutb(w_asqrt60_2[1]),.doutc(w_asqrt60_2[2]),.din(w_asqrt60_0[1]));
	jspl3 jspl3_w_asqrt60_3(.douta(w_asqrt60_3[0]),.doutb(w_asqrt60_3[1]),.doutc(w_asqrt60_3[2]),.din(w_asqrt60_0[2]));
	jspl3 jspl3_w_asqrt60_4(.douta(w_asqrt60_4[0]),.doutb(w_asqrt60_4[1]),.doutc(w_asqrt60_4[2]),.din(w_asqrt60_1[0]));
	jspl3 jspl3_w_asqrt60_5(.douta(w_asqrt60_5[0]),.doutb(w_asqrt60_5[1]),.doutc(w_asqrt60_5[2]),.din(w_asqrt60_1[1]));
	jspl3 jspl3_w_asqrt60_6(.douta(w_asqrt60_6[0]),.doutb(w_asqrt60_6[1]),.doutc(w_asqrt60_6[2]),.din(w_asqrt60_1[2]));
	jspl3 jspl3_w_asqrt60_7(.douta(w_asqrt60_7[0]),.doutb(w_asqrt60_7[1]),.doutc(w_asqrt60_7[2]),.din(w_asqrt60_2[0]));
	jspl3 jspl3_w_asqrt60_8(.douta(w_asqrt60_8[0]),.doutb(w_asqrt60_8[1]),.doutc(w_asqrt60_8[2]),.din(w_asqrt60_2[1]));
	jspl3 jspl3_w_asqrt60_9(.douta(w_asqrt60_9[0]),.doutb(w_asqrt60_9[1]),.doutc(w_asqrt60_9[2]),.din(w_asqrt60_2[2]));
	jspl3 jspl3_w_asqrt60_10(.douta(w_asqrt60_10[0]),.doutb(w_asqrt60_10[1]),.doutc(w_asqrt60_10[2]),.din(w_asqrt60_3[0]));
	jspl3 jspl3_w_asqrt60_11(.douta(w_asqrt60_11[0]),.doutb(w_asqrt60_11[1]),.doutc(w_asqrt60_11[2]),.din(w_asqrt60_3[1]));
	jspl3 jspl3_w_asqrt60_12(.douta(w_asqrt60_12[0]),.doutb(w_asqrt60_12[1]),.doutc(w_asqrt60_12[2]),.din(w_asqrt60_3[2]));
	jspl3 jspl3_w_asqrt60_13(.douta(w_asqrt60_13[0]),.doutb(w_asqrt60_13[1]),.doutc(w_asqrt60_13[2]),.din(w_asqrt60_4[0]));
	jspl3 jspl3_w_asqrt60_14(.douta(w_asqrt60_14[0]),.doutb(w_asqrt60_14[1]),.doutc(w_asqrt60_14[2]),.din(w_asqrt60_4[1]));
	jspl3 jspl3_w_asqrt60_15(.douta(w_asqrt60_15[0]),.doutb(w_asqrt60_15[1]),.doutc(w_asqrt60_15[2]),.din(w_asqrt60_4[2]));
	jspl3 jspl3_w_asqrt60_16(.douta(w_asqrt60_16[0]),.doutb(w_asqrt60_16[1]),.doutc(w_asqrt60_16[2]),.din(w_asqrt60_5[0]));
	jspl3 jspl3_w_asqrt60_17(.douta(w_asqrt60_17[0]),.doutb(w_asqrt60_17[1]),.doutc(w_asqrt60_17[2]),.din(w_asqrt60_5[1]));
	jspl3 jspl3_w_asqrt60_18(.douta(w_asqrt60_18[0]),.doutb(w_asqrt60_18[1]),.doutc(w_asqrt60_18[2]),.din(w_asqrt60_5[2]));
	jspl3 jspl3_w_asqrt60_19(.douta(w_asqrt60_19[0]),.doutb(w_asqrt60_19[1]),.doutc(w_asqrt60_19[2]),.din(w_asqrt60_6[0]));
	jspl3 jspl3_w_asqrt60_20(.douta(w_asqrt60_20[0]),.doutb(w_asqrt60_20[1]),.doutc(w_asqrt60_20[2]),.din(w_asqrt60_6[1]));
	jspl3 jspl3_w_asqrt60_21(.douta(w_asqrt60_21[0]),.doutb(w_asqrt60_21[1]),.doutc(w_asqrt60_21[2]),.din(w_asqrt60_6[2]));
	jspl3 jspl3_w_asqrt60_22(.douta(w_asqrt60_22[0]),.doutb(w_asqrt60_22[1]),.doutc(w_asqrt60_22[2]),.din(w_asqrt60_7[0]));
	jspl3 jspl3_w_asqrt60_23(.douta(w_asqrt60_23[0]),.doutb(w_asqrt60_23[1]),.doutc(w_asqrt60_23[2]),.din(w_asqrt60_7[1]));
	jspl3 jspl3_w_asqrt60_24(.douta(w_asqrt60_24[0]),.doutb(w_asqrt60_24[1]),.doutc(w_asqrt60_24[2]),.din(w_asqrt60_7[2]));
	jspl3 jspl3_w_asqrt60_25(.douta(w_asqrt60_25[0]),.doutb(w_asqrt60_25[1]),.doutc(w_asqrt60_25[2]),.din(w_asqrt60_8[0]));
	jspl3 jspl3_w_asqrt60_26(.douta(w_asqrt60_26[0]),.doutb(w_asqrt60_26[1]),.doutc(w_asqrt60_26[2]),.din(w_asqrt60_8[1]));
	jspl3 jspl3_w_asqrt60_27(.douta(w_asqrt60_27[0]),.doutb(w_asqrt60_27[1]),.doutc(w_asqrt60_27[2]),.din(w_asqrt60_8[2]));
	jspl3 jspl3_w_asqrt60_28(.douta(w_asqrt60_28[0]),.doutb(w_asqrt60_28[1]),.doutc(w_asqrt60_28[2]),.din(w_asqrt60_9[0]));
	jspl3 jspl3_w_asqrt60_29(.douta(w_asqrt60_29[0]),.doutb(w_asqrt60_29[1]),.doutc(w_asqrt60_29[2]),.din(w_asqrt60_9[1]));
	jspl3 jspl3_w_asqrt60_30(.douta(w_asqrt60_30[0]),.doutb(w_asqrt60_30[1]),.doutc(w_asqrt60_30[2]),.din(w_asqrt60_9[2]));
	jspl3 jspl3_w_asqrt60_31(.douta(w_asqrt60_31[0]),.doutb(w_asqrt60_31[1]),.doutc(w_asqrt60_31[2]),.din(w_asqrt60_10[0]));
	jspl3 jspl3_w_asqrt60_32(.douta(w_asqrt60_32[0]),.doutb(w_asqrt60_32[1]),.doutc(w_asqrt60_32[2]),.din(w_asqrt60_10[1]));
	jspl3 jspl3_w_asqrt60_33(.douta(w_asqrt60_33[0]),.doutb(w_asqrt60_33[1]),.doutc(w_asqrt60_33[2]),.din(w_asqrt60_10[2]));
	jspl3 jspl3_w_asqrt60_34(.douta(w_asqrt60_34[0]),.doutb(w_asqrt60_34[1]),.doutc(w_asqrt60_34[2]),.din(w_asqrt60_11[0]));
	jspl3 jspl3_w_asqrt60_35(.douta(w_asqrt60_35[0]),.doutb(w_asqrt60_35[1]),.doutc(w_asqrt60_35[2]),.din(w_asqrt60_11[1]));
	jspl3 jspl3_w_asqrt60_36(.douta(w_asqrt60_36[0]),.doutb(w_asqrt60_36[1]),.doutc(w_asqrt60_36[2]),.din(w_asqrt60_11[2]));
	jspl3 jspl3_w_asqrt60_37(.douta(w_asqrt60_37[0]),.doutb(w_asqrt60_37[1]),.doutc(w_asqrt60_37[2]),.din(w_asqrt60_12[0]));
	jspl3 jspl3_w_asqrt60_38(.douta(w_asqrt60_38[0]),.doutb(w_asqrt60_38[1]),.doutc(w_asqrt60_38[2]),.din(w_asqrt60_12[1]));
	jspl3 jspl3_w_asqrt60_39(.douta(w_asqrt60_39[0]),.doutb(w_asqrt60_39[1]),.doutc(w_asqrt60_39[2]),.din(w_asqrt60_12[2]));
	jspl3 jspl3_w_asqrt60_40(.douta(w_asqrt60_40[0]),.doutb(w_asqrt60_40[1]),.doutc(w_asqrt60_40[2]),.din(w_asqrt60_13[0]));
	jspl3 jspl3_w_asqrt60_41(.douta(w_asqrt60_41[0]),.doutb(w_asqrt60_41[1]),.doutc(w_asqrt60_41[2]),.din(w_asqrt60_13[1]));
	jspl3 jspl3_w_asqrt60_42(.douta(w_asqrt60_42[0]),.doutb(w_asqrt60_42[1]),.doutc(w_asqrt60_42[2]),.din(w_asqrt60_13[2]));
	jspl3 jspl3_w_asqrt60_43(.douta(w_asqrt60_43[0]),.doutb(w_asqrt60_43[1]),.doutc(w_asqrt60_43[2]),.din(w_asqrt60_14[0]));
	jspl3 jspl3_w_asqrt60_44(.douta(w_asqrt60_44[0]),.doutb(w_asqrt60_44[1]),.doutc(w_asqrt60_44[2]),.din(w_asqrt60_14[1]));
	jspl3 jspl3_w_asqrt60_45(.douta(w_asqrt60_45[0]),.doutb(w_asqrt60_45[1]),.doutc(asqrt[59]),.din(w_asqrt60_14[2]));
	jspl3 jspl3_w_asqrt61_0(.douta(w_asqrt61_0[0]),.doutb(w_asqrt61_0[1]),.doutc(w_asqrt61_0[2]),.din(asqrt_fa_61));
	jspl3 jspl3_w_asqrt61_1(.douta(w_asqrt61_1[0]),.doutb(w_asqrt61_1[1]),.doutc(w_asqrt61_1[2]),.din(w_asqrt61_0[0]));
	jspl3 jspl3_w_asqrt61_2(.douta(w_asqrt61_2[0]),.doutb(w_asqrt61_2[1]),.doutc(w_asqrt61_2[2]),.din(w_asqrt61_0[1]));
	jspl3 jspl3_w_asqrt61_3(.douta(w_asqrt61_3[0]),.doutb(w_asqrt61_3[1]),.doutc(w_asqrt61_3[2]),.din(w_asqrt61_0[2]));
	jspl3 jspl3_w_asqrt61_4(.douta(w_asqrt61_4[0]),.doutb(w_asqrt61_4[1]),.doutc(w_asqrt61_4[2]),.din(w_asqrt61_1[0]));
	jspl3 jspl3_w_asqrt61_5(.douta(w_asqrt61_5[0]),.doutb(w_asqrt61_5[1]),.doutc(w_asqrt61_5[2]),.din(w_asqrt61_1[1]));
	jspl3 jspl3_w_asqrt61_6(.douta(w_asqrt61_6[0]),.doutb(w_asqrt61_6[1]),.doutc(w_asqrt61_6[2]),.din(w_asqrt61_1[2]));
	jspl3 jspl3_w_asqrt61_7(.douta(w_asqrt61_7[0]),.doutb(w_asqrt61_7[1]),.doutc(w_asqrt61_7[2]),.din(w_asqrt61_2[0]));
	jspl3 jspl3_w_asqrt61_8(.douta(w_asqrt61_8[0]),.doutb(w_asqrt61_8[1]),.doutc(w_asqrt61_8[2]),.din(w_asqrt61_2[1]));
	jspl3 jspl3_w_asqrt61_9(.douta(w_asqrt61_9[0]),.doutb(w_asqrt61_9[1]),.doutc(w_asqrt61_9[2]),.din(w_asqrt61_2[2]));
	jspl3 jspl3_w_asqrt61_10(.douta(w_asqrt61_10[0]),.doutb(w_asqrt61_10[1]),.doutc(w_asqrt61_10[2]),.din(w_asqrt61_3[0]));
	jspl3 jspl3_w_asqrt61_11(.douta(w_asqrt61_11[0]),.doutb(w_asqrt61_11[1]),.doutc(w_asqrt61_11[2]),.din(w_asqrt61_3[1]));
	jspl3 jspl3_w_asqrt61_12(.douta(w_asqrt61_12[0]),.doutb(w_asqrt61_12[1]),.doutc(w_asqrt61_12[2]),.din(w_asqrt61_3[2]));
	jspl3 jspl3_w_asqrt61_13(.douta(w_asqrt61_13[0]),.doutb(w_asqrt61_13[1]),.doutc(w_asqrt61_13[2]),.din(w_asqrt61_4[0]));
	jspl3 jspl3_w_asqrt61_14(.douta(w_asqrt61_14[0]),.doutb(w_asqrt61_14[1]),.doutc(w_asqrt61_14[2]),.din(w_asqrt61_4[1]));
	jspl3 jspl3_w_asqrt61_15(.douta(w_asqrt61_15[0]),.doutb(w_asqrt61_15[1]),.doutc(w_asqrt61_15[2]),.din(w_asqrt61_4[2]));
	jspl3 jspl3_w_asqrt61_16(.douta(w_asqrt61_16[0]),.doutb(w_asqrt61_16[1]),.doutc(w_asqrt61_16[2]),.din(w_asqrt61_5[0]));
	jspl3 jspl3_w_asqrt61_17(.douta(w_asqrt61_17[0]),.doutb(w_asqrt61_17[1]),.doutc(w_asqrt61_17[2]),.din(w_asqrt61_5[1]));
	jspl3 jspl3_w_asqrt61_18(.douta(w_asqrt61_18[0]),.doutb(w_asqrt61_18[1]),.doutc(w_asqrt61_18[2]),.din(w_asqrt61_5[2]));
	jspl3 jspl3_w_asqrt61_19(.douta(w_asqrt61_19[0]),.doutb(w_asqrt61_19[1]),.doutc(w_asqrt61_19[2]),.din(w_asqrt61_6[0]));
	jspl3 jspl3_w_asqrt61_20(.douta(w_asqrt61_20[0]),.doutb(w_asqrt61_20[1]),.doutc(w_asqrt61_20[2]),.din(w_asqrt61_6[1]));
	jspl3 jspl3_w_asqrt61_21(.douta(w_asqrt61_21[0]),.doutb(w_asqrt61_21[1]),.doutc(w_asqrt61_21[2]),.din(w_asqrt61_6[2]));
	jspl3 jspl3_w_asqrt61_22(.douta(w_asqrt61_22[0]),.doutb(w_asqrt61_22[1]),.doutc(w_asqrt61_22[2]),.din(w_asqrt61_7[0]));
	jspl3 jspl3_w_asqrt61_23(.douta(w_asqrt61_23[0]),.doutb(w_asqrt61_23[1]),.doutc(w_asqrt61_23[2]),.din(w_asqrt61_7[1]));
	jspl3 jspl3_w_asqrt61_24(.douta(w_asqrt61_24[0]),.doutb(w_asqrt61_24[1]),.doutc(w_asqrt61_24[2]),.din(w_asqrt61_7[2]));
	jspl3 jspl3_w_asqrt61_25(.douta(w_asqrt61_25[0]),.doutb(w_asqrt61_25[1]),.doutc(w_asqrt61_25[2]),.din(w_asqrt61_8[0]));
	jspl3 jspl3_w_asqrt61_26(.douta(w_asqrt61_26[0]),.doutb(w_asqrt61_26[1]),.doutc(w_asqrt61_26[2]),.din(w_asqrt61_8[1]));
	jspl3 jspl3_w_asqrt61_27(.douta(w_asqrt61_27[0]),.doutb(w_asqrt61_27[1]),.doutc(w_asqrt61_27[2]),.din(w_asqrt61_8[2]));
	jspl3 jspl3_w_asqrt61_28(.douta(w_asqrt61_28[0]),.doutb(w_asqrt61_28[1]),.doutc(w_asqrt61_28[2]),.din(w_asqrt61_9[0]));
	jspl3 jspl3_w_asqrt61_29(.douta(w_asqrt61_29[0]),.doutb(w_asqrt61_29[1]),.doutc(w_asqrt61_29[2]),.din(w_asqrt61_9[1]));
	jspl3 jspl3_w_asqrt61_30(.douta(w_asqrt61_30[0]),.doutb(w_asqrt61_30[1]),.doutc(w_asqrt61_30[2]),.din(w_asqrt61_9[2]));
	jspl3 jspl3_w_asqrt61_31(.douta(w_asqrt61_31[0]),.doutb(w_asqrt61_31[1]),.doutc(w_asqrt61_31[2]),.din(w_asqrt61_10[0]));
	jspl3 jspl3_w_asqrt61_32(.douta(w_asqrt61_32[0]),.doutb(w_asqrt61_32[1]),.doutc(w_asqrt61_32[2]),.din(w_asqrt61_10[1]));
	jspl3 jspl3_w_asqrt61_33(.douta(w_asqrt61_33[0]),.doutb(w_asqrt61_33[1]),.doutc(w_asqrt61_33[2]),.din(w_asqrt61_10[2]));
	jspl3 jspl3_w_asqrt61_34(.douta(w_asqrt61_34[0]),.doutb(w_asqrt61_34[1]),.doutc(w_asqrt61_34[2]),.din(w_asqrt61_11[0]));
	jspl3 jspl3_w_asqrt61_35(.douta(w_asqrt61_35[0]),.doutb(w_asqrt61_35[1]),.doutc(w_asqrt61_35[2]),.din(w_asqrt61_11[1]));
	jspl3 jspl3_w_asqrt61_36(.douta(w_asqrt61_36[0]),.doutb(w_asqrt61_36[1]),.doutc(w_asqrt61_36[2]),.din(w_asqrt61_11[2]));
	jspl3 jspl3_w_asqrt61_37(.douta(w_asqrt61_37[0]),.doutb(w_asqrt61_37[1]),.doutc(w_asqrt61_37[2]),.din(w_asqrt61_12[0]));
	jspl3 jspl3_w_asqrt61_38(.douta(w_asqrt61_38[0]),.doutb(w_asqrt61_38[1]),.doutc(w_asqrt61_38[2]),.din(w_asqrt61_12[1]));
	jspl3 jspl3_w_asqrt61_39(.douta(w_asqrt61_39[0]),.doutb(w_asqrt61_39[1]),.doutc(w_asqrt61_39[2]),.din(w_asqrt61_12[2]));
	jspl3 jspl3_w_asqrt61_40(.douta(w_asqrt61_40[0]),.doutb(w_asqrt61_40[1]),.doutc(w_asqrt61_40[2]),.din(w_asqrt61_13[0]));
	jspl3 jspl3_w_asqrt61_41(.douta(w_asqrt61_41[0]),.doutb(w_asqrt61_41[1]),.doutc(w_asqrt61_41[2]),.din(w_asqrt61_13[1]));
	jspl3 jspl3_w_asqrt61_42(.douta(w_asqrt61_42[0]),.doutb(w_asqrt61_42[1]),.doutc(w_asqrt61_42[2]),.din(w_asqrt61_13[2]));
	jspl3 jspl3_w_asqrt61_43(.douta(w_asqrt61_43[0]),.doutb(w_asqrt61_43[1]),.doutc(w_asqrt61_43[2]),.din(w_asqrt61_14[0]));
	jspl3 jspl3_w_asqrt61_44(.douta(w_asqrt61_44[0]),.doutb(w_asqrt61_44[1]),.doutc(w_asqrt61_44[2]),.din(w_asqrt61_14[1]));
	jspl jspl_w_asqrt61_45(.douta(w_asqrt61_45),.doutb(asqrt[60]),.din(w_asqrt61_14[2]));
	jspl3 jspl3_w_asqrt62_0(.douta(w_asqrt62_0[0]),.doutb(w_asqrt62_0[1]),.doutc(w_asqrt62_0[2]),.din(asqrt_fa_62));
	jspl3 jspl3_w_asqrt62_1(.douta(w_asqrt62_1[0]),.doutb(w_asqrt62_1[1]),.doutc(w_asqrt62_1[2]),.din(w_asqrt62_0[0]));
	jspl3 jspl3_w_asqrt62_2(.douta(w_asqrt62_2[0]),.doutb(w_asqrt62_2[1]),.doutc(w_asqrt62_2[2]),.din(w_asqrt62_0[1]));
	jspl3 jspl3_w_asqrt62_3(.douta(w_asqrt62_3[0]),.doutb(w_asqrt62_3[1]),.doutc(w_asqrt62_3[2]),.din(w_asqrt62_0[2]));
	jspl3 jspl3_w_asqrt62_4(.douta(w_asqrt62_4[0]),.doutb(w_asqrt62_4[1]),.doutc(w_asqrt62_4[2]),.din(w_asqrt62_1[0]));
	jspl3 jspl3_w_asqrt62_5(.douta(w_asqrt62_5[0]),.doutb(w_asqrt62_5[1]),.doutc(w_asqrt62_5[2]),.din(w_asqrt62_1[1]));
	jspl3 jspl3_w_asqrt62_6(.douta(w_asqrt62_6[0]),.doutb(w_asqrt62_6[1]),.doutc(w_asqrt62_6[2]),.din(w_asqrt62_1[2]));
	jspl3 jspl3_w_asqrt62_7(.douta(w_asqrt62_7[0]),.doutb(w_asqrt62_7[1]),.doutc(w_asqrt62_7[2]),.din(w_asqrt62_2[0]));
	jspl3 jspl3_w_asqrt62_8(.douta(w_asqrt62_8[0]),.doutb(w_asqrt62_8[1]),.doutc(w_asqrt62_8[2]),.din(w_asqrt62_2[1]));
	jspl3 jspl3_w_asqrt62_9(.douta(w_asqrt62_9[0]),.doutb(w_asqrt62_9[1]),.doutc(w_asqrt62_9[2]),.din(w_asqrt62_2[2]));
	jspl3 jspl3_w_asqrt62_10(.douta(w_asqrt62_10[0]),.doutb(w_asqrt62_10[1]),.doutc(w_asqrt62_10[2]),.din(w_asqrt62_3[0]));
	jspl3 jspl3_w_asqrt62_11(.douta(w_asqrt62_11[0]),.doutb(w_asqrt62_11[1]),.doutc(w_asqrt62_11[2]),.din(w_asqrt62_3[1]));
	jspl3 jspl3_w_asqrt62_12(.douta(w_asqrt62_12[0]),.doutb(w_asqrt62_12[1]),.doutc(w_asqrt62_12[2]),.din(w_asqrt62_3[2]));
	jspl3 jspl3_w_asqrt62_13(.douta(w_asqrt62_13[0]),.doutb(w_asqrt62_13[1]),.doutc(w_asqrt62_13[2]),.din(w_asqrt62_4[0]));
	jspl3 jspl3_w_asqrt62_14(.douta(w_asqrt62_14[0]),.doutb(w_asqrt62_14[1]),.doutc(w_asqrt62_14[2]),.din(w_asqrt62_4[1]));
	jspl3 jspl3_w_asqrt62_15(.douta(w_asqrt62_15[0]),.doutb(w_asqrt62_15[1]),.doutc(w_asqrt62_15[2]),.din(w_asqrt62_4[2]));
	jspl3 jspl3_w_asqrt62_16(.douta(w_asqrt62_16[0]),.doutb(w_asqrt62_16[1]),.doutc(w_asqrt62_16[2]),.din(w_asqrt62_5[0]));
	jspl3 jspl3_w_asqrt62_17(.douta(w_asqrt62_17[0]),.doutb(w_asqrt62_17[1]),.doutc(w_asqrt62_17[2]),.din(w_asqrt62_5[1]));
	jspl3 jspl3_w_asqrt62_18(.douta(w_asqrt62_18[0]),.doutb(w_asqrt62_18[1]),.doutc(w_asqrt62_18[2]),.din(w_asqrt62_5[2]));
	jspl3 jspl3_w_asqrt62_19(.douta(w_asqrt62_19[0]),.doutb(w_asqrt62_19[1]),.doutc(w_asqrt62_19[2]),.din(w_asqrt62_6[0]));
	jspl3 jspl3_w_asqrt62_20(.douta(w_asqrt62_20[0]),.doutb(w_asqrt62_20[1]),.doutc(w_asqrt62_20[2]),.din(w_asqrt62_6[1]));
	jspl3 jspl3_w_asqrt62_21(.douta(w_asqrt62_21[0]),.doutb(w_asqrt62_21[1]),.doutc(w_asqrt62_21[2]),.din(w_asqrt62_6[2]));
	jspl3 jspl3_w_asqrt62_22(.douta(w_asqrt62_22[0]),.doutb(w_asqrt62_22[1]),.doutc(w_asqrt62_22[2]),.din(w_asqrt62_7[0]));
	jspl3 jspl3_w_asqrt62_23(.douta(w_asqrt62_23[0]),.doutb(w_asqrt62_23[1]),.doutc(w_asqrt62_23[2]),.din(w_asqrt62_7[1]));
	jspl3 jspl3_w_asqrt62_24(.douta(w_asqrt62_24[0]),.doutb(w_asqrt62_24[1]),.doutc(w_asqrt62_24[2]),.din(w_asqrt62_7[2]));
	jspl3 jspl3_w_asqrt62_25(.douta(w_asqrt62_25[0]),.doutb(w_asqrt62_25[1]),.doutc(w_asqrt62_25[2]),.din(w_asqrt62_8[0]));
	jspl3 jspl3_w_asqrt62_26(.douta(w_asqrt62_26[0]),.doutb(w_asqrt62_26[1]),.doutc(w_asqrt62_26[2]),.din(w_asqrt62_8[1]));
	jspl3 jspl3_w_asqrt62_27(.douta(w_asqrt62_27[0]),.doutb(w_asqrt62_27[1]),.doutc(w_asqrt62_27[2]),.din(w_asqrt62_8[2]));
	jspl3 jspl3_w_asqrt62_28(.douta(w_asqrt62_28[0]),.doutb(w_asqrt62_28[1]),.doutc(w_asqrt62_28[2]),.din(w_asqrt62_9[0]));
	jspl3 jspl3_w_asqrt62_29(.douta(w_asqrt62_29[0]),.doutb(w_asqrt62_29[1]),.doutc(w_asqrt62_29[2]),.din(w_asqrt62_9[1]));
	jspl3 jspl3_w_asqrt62_30(.douta(w_asqrt62_30[0]),.doutb(w_asqrt62_30[1]),.doutc(w_asqrt62_30[2]),.din(w_asqrt62_9[2]));
	jspl3 jspl3_w_asqrt62_31(.douta(w_asqrt62_31[0]),.doutb(w_asqrt62_31[1]),.doutc(w_asqrt62_31[2]),.din(w_asqrt62_10[0]));
	jspl3 jspl3_w_asqrt62_32(.douta(w_asqrt62_32[0]),.doutb(w_asqrt62_32[1]),.doutc(w_asqrt62_32[2]),.din(w_asqrt62_10[1]));
	jspl3 jspl3_w_asqrt62_33(.douta(w_asqrt62_33[0]),.doutb(w_asqrt62_33[1]),.doutc(w_asqrt62_33[2]),.din(w_asqrt62_10[2]));
	jspl3 jspl3_w_asqrt62_34(.douta(w_asqrt62_34[0]),.doutb(w_asqrt62_34[1]),.doutc(w_asqrt62_34[2]),.din(w_asqrt62_11[0]));
	jspl3 jspl3_w_asqrt62_35(.douta(w_asqrt62_35[0]),.doutb(w_asqrt62_35[1]),.doutc(w_asqrt62_35[2]),.din(w_asqrt62_11[1]));
	jspl3 jspl3_w_asqrt62_36(.douta(w_asqrt62_36[0]),.doutb(w_asqrt62_36[1]),.doutc(w_asqrt62_36[2]),.din(w_asqrt62_11[2]));
	jspl3 jspl3_w_asqrt62_37(.douta(w_asqrt62_37[0]),.doutb(w_asqrt62_37[1]),.doutc(w_asqrt62_37[2]),.din(w_asqrt62_12[0]));
	jspl3 jspl3_w_asqrt62_38(.douta(w_asqrt62_38[0]),.doutb(w_asqrt62_38[1]),.doutc(w_asqrt62_38[2]),.din(w_asqrt62_12[1]));
	jspl3 jspl3_w_asqrt62_39(.douta(w_asqrt62_39[0]),.doutb(w_asqrt62_39[1]),.doutc(w_asqrt62_39[2]),.din(w_asqrt62_12[2]));
	jspl3 jspl3_w_asqrt62_40(.douta(w_asqrt62_40[0]),.doutb(w_asqrt62_40[1]),.doutc(w_asqrt62_40[2]),.din(w_asqrt62_13[0]));
	jspl3 jspl3_w_asqrt62_41(.douta(w_asqrt62_41[0]),.doutb(w_asqrt62_41[1]),.doutc(w_asqrt62_41[2]),.din(w_asqrt62_13[1]));
	jspl3 jspl3_w_asqrt62_42(.douta(w_asqrt62_42[0]),.doutb(w_asqrt62_42[1]),.doutc(w_asqrt62_42[2]),.din(w_asqrt62_13[2]));
	jspl3 jspl3_w_asqrt62_43(.douta(w_asqrt62_43[0]),.doutb(w_asqrt62_43[1]),.doutc(w_asqrt62_43[2]),.din(w_asqrt62_14[0]));
	jspl3 jspl3_w_asqrt62_44(.douta(w_asqrt62_44[0]),.doutb(w_asqrt62_44[1]),.doutc(w_asqrt62_44[2]),.din(w_asqrt62_14[1]));
	jspl3 jspl3_w_asqrt62_45(.douta(w_asqrt62_45[0]),.doutb(w_asqrt62_45[1]),.doutc(asqrt[61]),.din(w_asqrt62_14[2]));
	jspl3 jspl3_w_asqrt63_0(.douta(w_asqrt63_0[0]),.doutb(w_asqrt63_0[1]),.doutc(w_asqrt63_0[2]),.din(asqrt_fa_63));
	jspl3 jspl3_w_asqrt63_1(.douta(w_asqrt63_1[0]),.doutb(w_asqrt63_1[1]),.doutc(w_asqrt63_1[2]),.din(w_asqrt63_0[0]));
	jspl3 jspl3_w_asqrt63_2(.douta(w_asqrt63_2[0]),.doutb(w_asqrt63_2[1]),.doutc(w_asqrt63_2[2]),.din(w_asqrt63_0[1]));
	jspl3 jspl3_w_asqrt63_3(.douta(w_asqrt63_3[0]),.doutb(w_asqrt63_3[1]),.doutc(w_asqrt63_3[2]),.din(w_asqrt63_0[2]));
	jspl3 jspl3_w_asqrt63_4(.douta(w_asqrt63_4[0]),.doutb(w_asqrt63_4[1]),.doutc(w_asqrt63_4[2]),.din(w_asqrt63_1[0]));
	jspl3 jspl3_w_asqrt63_5(.douta(w_asqrt63_5[0]),.doutb(w_asqrt63_5[1]),.doutc(w_asqrt63_5[2]),.din(w_asqrt63_1[1]));
	jspl3 jspl3_w_asqrt63_6(.douta(w_asqrt63_6[0]),.doutb(w_asqrt63_6[1]),.doutc(w_asqrt63_6[2]),.din(w_asqrt63_1[2]));
	jspl3 jspl3_w_asqrt63_7(.douta(w_asqrt63_7[0]),.doutb(w_asqrt63_7[1]),.doutc(w_asqrt63_7[2]),.din(w_asqrt63_2[0]));
	jspl3 jspl3_w_asqrt63_8(.douta(w_asqrt63_8[0]),.doutb(w_asqrt63_8[1]),.doutc(w_asqrt63_8[2]),.din(w_asqrt63_2[1]));
	jspl3 jspl3_w_asqrt63_9(.douta(w_asqrt63_9[0]),.doutb(w_asqrt63_9[1]),.doutc(w_asqrt63_9[2]),.din(w_asqrt63_2[2]));
	jspl3 jspl3_w_asqrt63_10(.douta(w_asqrt63_10[0]),.doutb(w_asqrt63_10[1]),.doutc(w_asqrt63_10[2]),.din(w_asqrt63_3[0]));
	jspl3 jspl3_w_asqrt63_11(.douta(w_asqrt63_11[0]),.doutb(w_asqrt63_11[1]),.doutc(w_asqrt63_11[2]),.din(w_asqrt63_3[1]));
	jspl3 jspl3_w_asqrt63_12(.douta(w_asqrt63_12[0]),.doutb(w_asqrt63_12[1]),.doutc(w_asqrt63_12[2]),.din(w_asqrt63_3[2]));
	jspl3 jspl3_w_asqrt63_13(.douta(w_asqrt63_13[0]),.doutb(w_asqrt63_13[1]),.doutc(w_asqrt63_13[2]),.din(w_asqrt63_4[0]));
	jspl3 jspl3_w_asqrt63_14(.douta(w_asqrt63_14[0]),.doutb(w_asqrt63_14[1]),.doutc(w_asqrt63_14[2]),.din(w_asqrt63_4[1]));
	jspl3 jspl3_w_asqrt63_15(.douta(w_asqrt63_15[0]),.doutb(w_asqrt63_15[1]),.doutc(w_asqrt63_15[2]),.din(w_asqrt63_4[2]));
	jspl3 jspl3_w_asqrt63_16(.douta(w_asqrt63_16[0]),.doutb(w_asqrt63_16[1]),.doutc(w_asqrt63_16[2]),.din(w_asqrt63_5[0]));
	jspl3 jspl3_w_asqrt63_17(.douta(w_asqrt63_17[0]),.doutb(w_asqrt63_17[1]),.doutc(w_asqrt63_17[2]),.din(w_asqrt63_5[1]));
	jspl3 jspl3_w_asqrt63_18(.douta(w_asqrt63_18[0]),.doutb(w_asqrt63_18[1]),.doutc(w_asqrt63_18[2]),.din(w_asqrt63_5[2]));
	jspl3 jspl3_w_asqrt63_19(.douta(w_asqrt63_19[0]),.doutb(w_asqrt63_19[1]),.doutc(w_asqrt63_19[2]),.din(w_asqrt63_6[0]));
	jspl3 jspl3_w_asqrt63_20(.douta(w_asqrt63_20[0]),.doutb(w_asqrt63_20[1]),.doutc(w_asqrt63_20[2]),.din(w_asqrt63_6[1]));
	jspl3 jspl3_w_asqrt63_21(.douta(w_asqrt63_21[0]),.doutb(w_asqrt63_21[1]),.doutc(w_asqrt63_21[2]),.din(w_asqrt63_6[2]));
	jspl3 jspl3_w_asqrt63_22(.douta(w_asqrt63_22[0]),.doutb(w_asqrt63_22[1]),.doutc(w_asqrt63_22[2]),.din(w_asqrt63_7[0]));
	jspl3 jspl3_w_asqrt63_23(.douta(w_asqrt63_23[0]),.doutb(w_asqrt63_23[1]),.doutc(w_asqrt63_23[2]),.din(w_asqrt63_7[1]));
	jspl3 jspl3_w_asqrt63_24(.douta(w_asqrt63_24[0]),.doutb(w_asqrt63_24[1]),.doutc(w_asqrt63_24[2]),.din(w_asqrt63_7[2]));
	jspl3 jspl3_w_asqrt63_25(.douta(w_asqrt63_25[0]),.doutb(w_asqrt63_25[1]),.doutc(w_asqrt63_25[2]),.din(w_asqrt63_8[0]));
	jspl3 jspl3_w_asqrt63_26(.douta(w_asqrt63_26[0]),.doutb(w_asqrt63_26[1]),.doutc(w_asqrt63_26[2]),.din(w_asqrt63_8[1]));
	jspl3 jspl3_w_asqrt63_27(.douta(w_asqrt63_27[0]),.doutb(w_asqrt63_27[1]),.doutc(w_asqrt63_27[2]),.din(w_asqrt63_8[2]));
	jspl3 jspl3_w_asqrt63_28(.douta(w_asqrt63_28[0]),.doutb(w_asqrt63_28[1]),.doutc(w_asqrt63_28[2]),.din(w_asqrt63_9[0]));
	jspl3 jspl3_w_asqrt63_29(.douta(w_asqrt63_29[0]),.doutb(w_asqrt63_29[1]),.doutc(w_asqrt63_29[2]),.din(w_asqrt63_9[1]));
	jspl3 jspl3_w_asqrt63_30(.douta(w_asqrt63_30[0]),.doutb(w_asqrt63_30[1]),.doutc(w_asqrt63_30[2]),.din(w_asqrt63_9[2]));
	jspl3 jspl3_w_asqrt63_31(.douta(w_asqrt63_31[0]),.doutb(w_asqrt63_31[1]),.doutc(w_asqrt63_31[2]),.din(w_asqrt63_10[0]));
	jspl3 jspl3_w_asqrt63_32(.douta(w_asqrt63_32[0]),.doutb(w_asqrt63_32[1]),.doutc(w_asqrt63_32[2]),.din(w_asqrt63_10[1]));
	jspl3 jspl3_w_asqrt63_33(.douta(w_asqrt63_33[0]),.doutb(w_asqrt63_33[1]),.doutc(w_asqrt63_33[2]),.din(w_asqrt63_10[2]));
	jspl3 jspl3_w_asqrt63_34(.douta(w_asqrt63_34[0]),.doutb(w_asqrt63_34[1]),.doutc(w_asqrt63_34[2]),.din(w_asqrt63_11[0]));
	jspl3 jspl3_w_asqrt63_35(.douta(w_asqrt63_35[0]),.doutb(w_asqrt63_35[1]),.doutc(w_asqrt63_35[2]),.din(w_asqrt63_11[1]));
	jspl3 jspl3_w_asqrt63_36(.douta(w_asqrt63_36[0]),.doutb(w_asqrt63_36[1]),.doutc(w_asqrt63_36[2]),.din(w_asqrt63_11[2]));
	jspl3 jspl3_w_asqrt63_37(.douta(w_asqrt63_37[0]),.doutb(w_asqrt63_37[1]),.doutc(w_asqrt63_37[2]),.din(w_asqrt63_12[0]));
	jspl3 jspl3_w_asqrt63_38(.douta(w_asqrt63_38[0]),.doutb(w_asqrt63_38[1]),.doutc(w_asqrt63_38[2]),.din(w_asqrt63_12[1]));
	jspl3 jspl3_w_asqrt63_39(.douta(w_asqrt63_39[0]),.doutb(w_asqrt63_39[1]),.doutc(w_asqrt63_39[2]),.din(w_asqrt63_12[2]));
	jspl3 jspl3_w_asqrt63_40(.douta(w_asqrt63_40[0]),.doutb(w_asqrt63_40[1]),.doutc(w_asqrt63_40[2]),.din(w_asqrt63_13[0]));
	jspl3 jspl3_w_asqrt63_41(.douta(w_asqrt63_41[0]),.doutb(w_asqrt63_41[1]),.doutc(w_asqrt63_41[2]),.din(w_asqrt63_13[1]));
	jspl3 jspl3_w_asqrt63_42(.douta(w_asqrt63_42[0]),.doutb(w_asqrt63_42[1]),.doutc(w_asqrt63_42[2]),.din(w_asqrt63_13[2]));
	jspl3 jspl3_w_asqrt63_43(.douta(w_asqrt63_43[0]),.doutb(w_asqrt63_43[1]),.doutc(w_asqrt63_43[2]),.din(w_asqrt63_14[0]));
	jspl3 jspl3_w_asqrt63_44(.douta(w_asqrt63_44[0]),.doutb(w_asqrt63_44[1]),.doutc(w_asqrt63_44[2]),.din(w_asqrt63_14[1]));
	jspl3 jspl3_w_asqrt63_45(.douta(w_asqrt63_45[0]),.doutb(w_asqrt63_45[1]),.doutc(w_asqrt63_45[2]),.din(w_asqrt63_14[2]));
	jspl3 jspl3_w_asqrt63_46(.douta(w_asqrt63_46[0]),.doutb(w_asqrt63_46[1]),.doutc(w_asqrt63_46[2]),.din(w_asqrt63_15[0]));
	jspl3 jspl3_w_asqrt63_47(.douta(w_asqrt63_47[0]),.doutb(w_asqrt63_47[1]),.doutc(w_asqrt63_47[2]),.din(w_asqrt63_15[1]));
	jspl3 jspl3_w_asqrt63_48(.douta(w_asqrt63_48[0]),.doutb(w_asqrt63_48[1]),.doutc(w_asqrt63_48[2]),.din(w_asqrt63_15[2]));
	jspl3 jspl3_w_asqrt63_49(.douta(w_asqrt63_49[0]),.doutb(w_asqrt63_49[1]),.doutc(w_asqrt63_49[2]),.din(w_asqrt63_16[0]));
	jspl3 jspl3_w_asqrt63_50(.douta(w_asqrt63_50[0]),.doutb(w_asqrt63_50[1]),.doutc(w_asqrt63_50[2]),.din(w_asqrt63_16[1]));
	jspl3 jspl3_w_asqrt63_51(.douta(w_asqrt63_51[0]),.doutb(w_asqrt63_51[1]),.doutc(w_asqrt63_51[2]),.din(w_asqrt63_16[2]));
	jspl3 jspl3_w_asqrt63_52(.douta(w_asqrt63_52[0]),.doutb(w_asqrt63_52[1]),.doutc(w_asqrt63_52[2]),.din(w_asqrt63_17[0]));
	jspl3 jspl3_w_asqrt63_53(.douta(w_asqrt63_53[0]),.doutb(w_asqrt63_53[1]),.doutc(w_asqrt63_53[2]),.din(w_asqrt63_17[1]));
	jspl3 jspl3_w_asqrt63_54(.douta(w_asqrt63_54[0]),.doutb(w_asqrt63_54[1]),.doutc(w_asqrt63_54[2]),.din(w_asqrt63_17[2]));
	jspl3 jspl3_w_asqrt63_55(.douta(w_asqrt63_55[0]),.doutb(w_asqrt63_55[1]),.doutc(w_asqrt63_55[2]),.din(w_asqrt63_18[0]));
	jspl3 jspl3_w_asqrt63_56(.douta(w_asqrt63_56[0]),.doutb(w_asqrt63_56[1]),.doutc(w_asqrt63_56[2]),.din(w_asqrt63_18[1]));
	jspl jspl_w_asqrt63_57(.douta(w_asqrt63_57),.doutb(asqrt[62]),.din(w_asqrt63_18[2]));
	jspl3 jspl3_w_n192_0(.douta(w_n192_0[0]),.doutb(w_n192_0[1]),.doutc(w_n192_0[2]),.din(n192));
	jspl jspl_w_n193_0(.douta(w_n193_0[0]),.doutb(w_n193_0[1]),.din(n193));
	jspl jspl_w_n195_0(.douta(w_n195_0[0]),.doutb(w_n195_0[1]),.din(n195));
	jspl jspl_w_n197_0(.douta(w_n197_0[0]),.doutb(w_n197_0[1]),.din(n197));
	jspl3 jspl3_w_n198_0(.douta(w_n198_0[0]),.doutb(w_n198_0[1]),.doutc(w_n198_0[2]),.din(n198));
	jspl jspl_w_n198_1(.douta(w_n198_1[0]),.doutb(w_n198_1[1]),.din(w_n198_0[0]));
	jspl jspl_w_n199_0(.douta(w_n199_0[0]),.doutb(w_n199_0[1]),.din(n199));
	jspl3 jspl3_w_n200_0(.douta(w_n200_0[0]),.doutb(w_n200_0[1]),.doutc(w_n200_0[2]),.din(n200));
	jspl jspl_w_n203_0(.douta(w_n203_0[0]),.doutb(w_n203_0[1]),.din(n203));
	jspl3 jspl3_w_n204_0(.douta(w_n204_0[0]),.doutb(w_n204_0[1]),.doutc(w_n204_0[2]),.din(n204));
	jspl jspl_w_n207_0(.douta(w_n207_0[0]),.doutb(w_n207_0[1]),.din(n207));
	jspl jspl_w_n209_0(.douta(w_n209_0[0]),.doutb(w_n209_0[1]),.din(n209));
	jspl3 jspl3_w_n211_0(.douta(w_n211_0[0]),.doutb(w_n211_0[1]),.doutc(w_n211_0[2]),.din(n211));
	jspl jspl_w_n211_1(.douta(w_n211_1[0]),.doutb(w_n211_1[1]),.din(w_n211_0[0]));
	jspl jspl_w_n212_0(.douta(w_n212_0[0]),.doutb(w_n212_0[1]),.din(n212));
	jspl3 jspl3_w_n215_0(.douta(w_n215_0[0]),.doutb(w_n215_0[1]),.doutc(w_n215_0[2]),.din(n215));
	jspl3 jspl3_w_n216_0(.douta(w_n216_0[0]),.doutb(w_n216_0[1]),.doutc(w_n216_0[2]),.din(n216));
	jspl jspl_w_n216_1(.douta(w_n216_1[0]),.doutb(w_n216_1[1]),.din(w_n216_0[0]));
	jspl jspl_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.din(n217));
	jspl3 jspl3_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.doutc(w_n218_0[2]),.din(n218));
	jspl3 jspl3_w_n218_1(.douta(w_n218_1[0]),.doutb(w_n218_1[1]),.doutc(w_n218_1[2]),.din(w_n218_0[0]));
	jspl3 jspl3_w_n218_2(.douta(w_n218_2[0]),.doutb(w_n218_2[1]),.doutc(w_n218_2[2]),.din(w_n218_0[1]));
	jspl3 jspl3_w_n218_3(.douta(w_n218_3[0]),.doutb(w_n218_3[1]),.doutc(w_n218_3[2]),.din(w_n218_0[2]));
	jspl3 jspl3_w_n218_4(.douta(w_n218_4[0]),.doutb(w_n218_4[1]),.doutc(w_n218_4[2]),.din(w_n218_1[0]));
	jspl3 jspl3_w_n218_5(.douta(w_n218_5[0]),.doutb(w_n218_5[1]),.doutc(w_n218_5[2]),.din(w_n218_1[1]));
	jspl3 jspl3_w_n218_6(.douta(w_n218_6[0]),.doutb(w_n218_6[1]),.doutc(w_n218_6[2]),.din(w_n218_1[2]));
	jspl3 jspl3_w_n218_7(.douta(w_n218_7[0]),.doutb(w_n218_7[1]),.doutc(w_n218_7[2]),.din(w_n218_2[0]));
	jspl3 jspl3_w_n218_8(.douta(w_n218_8[0]),.doutb(w_n218_8[1]),.doutc(w_n218_8[2]),.din(w_n218_2[1]));
	jspl3 jspl3_w_n218_9(.douta(w_n218_9[0]),.doutb(w_n218_9[1]),.doutc(w_n218_9[2]),.din(w_n218_2[2]));
	jspl3 jspl3_w_n218_10(.douta(w_n218_10[0]),.doutb(w_n218_10[1]),.doutc(w_n218_10[2]),.din(w_n218_3[0]));
	jspl3 jspl3_w_n218_11(.douta(w_n218_11[0]),.doutb(w_n218_11[1]),.doutc(w_n218_11[2]),.din(w_n218_3[1]));
	jspl3 jspl3_w_n218_12(.douta(w_n218_12[0]),.doutb(w_n218_12[1]),.doutc(w_n218_12[2]),.din(w_n218_3[2]));
	jspl3 jspl3_w_n218_13(.douta(w_n218_13[0]),.doutb(w_n218_13[1]),.doutc(w_n218_13[2]),.din(w_n218_4[0]));
	jspl3 jspl3_w_n218_14(.douta(w_n218_14[0]),.doutb(w_n218_14[1]),.doutc(w_n218_14[2]),.din(w_n218_4[1]));
	jspl3 jspl3_w_n218_15(.douta(w_n218_15[0]),.doutb(w_n218_15[1]),.doutc(w_n218_15[2]),.din(w_n218_4[2]));
	jspl3 jspl3_w_n218_16(.douta(w_n218_16[0]),.doutb(w_n218_16[1]),.doutc(w_n218_16[2]),.din(w_n218_5[0]));
	jspl3 jspl3_w_n218_17(.douta(w_n218_17[0]),.doutb(w_n218_17[1]),.doutc(w_n218_17[2]),.din(w_n218_5[1]));
	jspl3 jspl3_w_n218_18(.douta(w_n218_18[0]),.doutb(w_n218_18[1]),.doutc(w_n218_18[2]),.din(w_n218_5[2]));
	jspl3 jspl3_w_n218_19(.douta(w_n218_19[0]),.doutb(w_n218_19[1]),.doutc(w_n218_19[2]),.din(w_n218_6[0]));
	jspl3 jspl3_w_n218_20(.douta(w_n218_20[0]),.doutb(w_n218_20[1]),.doutc(w_n218_20[2]),.din(w_n218_6[1]));
	jspl3 jspl3_w_n218_21(.douta(w_n218_21[0]),.doutb(w_n218_21[1]),.doutc(w_n218_21[2]),.din(w_n218_6[2]));
	jspl3 jspl3_w_n218_22(.douta(w_n218_22[0]),.doutb(w_n218_22[1]),.doutc(w_n218_22[2]),.din(w_n218_7[0]));
	jspl3 jspl3_w_n218_23(.douta(w_n218_23[0]),.doutb(w_n218_23[1]),.doutc(w_n218_23[2]),.din(w_n218_7[1]));
	jspl3 jspl3_w_n218_24(.douta(w_n218_24[0]),.doutb(w_n218_24[1]),.doutc(w_n218_24[2]),.din(w_n218_7[2]));
	jspl3 jspl3_w_n218_25(.douta(w_n218_25[0]),.doutb(w_n218_25[1]),.doutc(w_n218_25[2]),.din(w_n218_8[0]));
	jspl3 jspl3_w_n218_26(.douta(w_n218_26[0]),.doutb(w_n218_26[1]),.doutc(w_n218_26[2]),.din(w_n218_8[1]));
	jspl3 jspl3_w_n218_27(.douta(w_n218_27[0]),.doutb(w_n218_27[1]),.doutc(w_n218_27[2]),.din(w_n218_8[2]));
	jspl3 jspl3_w_n218_28(.douta(w_n218_28[0]),.doutb(w_n218_28[1]),.doutc(w_n218_28[2]),.din(w_n218_9[0]));
	jspl3 jspl3_w_n218_29(.douta(w_n218_29[0]),.doutb(w_n218_29[1]),.doutc(w_n218_29[2]),.din(w_n218_9[1]));
	jspl3 jspl3_w_n218_30(.douta(w_n218_30[0]),.doutb(w_n218_30[1]),.doutc(w_n218_30[2]),.din(w_n218_9[2]));
	jspl jspl_w_n218_31(.douta(w_n218_31[0]),.doutb(w_n218_31[1]),.din(w_n218_10[0]));
	jspl3 jspl3_w_n221_0(.douta(w_n221_0[0]),.doutb(w_n221_0[1]),.doutc(w_n221_0[2]),.din(n221));
	jspl3 jspl3_w_n221_1(.douta(w_n221_1[0]),.doutb(w_n221_1[1]),.doutc(w_n221_1[2]),.din(w_n221_0[0]));
	jspl3 jspl3_w_n221_2(.douta(w_n221_2[0]),.doutb(w_n221_2[1]),.doutc(w_n221_2[2]),.din(w_n221_0[1]));
	jspl3 jspl3_w_n221_3(.douta(w_n221_3[0]),.doutb(w_n221_3[1]),.doutc(w_n221_3[2]),.din(w_n221_0[2]));
	jspl3 jspl3_w_n221_4(.douta(w_n221_4[0]),.doutb(w_n221_4[1]),.doutc(w_n221_4[2]),.din(w_n221_1[0]));
	jspl3 jspl3_w_n221_5(.douta(w_n221_5[0]),.doutb(w_n221_5[1]),.doutc(w_n221_5[2]),.din(w_n221_1[1]));
	jspl3 jspl3_w_n221_6(.douta(w_n221_6[0]),.doutb(w_n221_6[1]),.doutc(w_n221_6[2]),.din(w_n221_1[2]));
	jspl3 jspl3_w_n221_7(.douta(w_n221_7[0]),.doutb(w_n221_7[1]),.doutc(w_n221_7[2]),.din(w_n221_2[0]));
	jspl3 jspl3_w_n221_8(.douta(w_n221_8[0]),.doutb(w_n221_8[1]),.doutc(w_n221_8[2]),.din(w_n221_2[1]));
	jspl3 jspl3_w_n221_9(.douta(w_n221_9[0]),.doutb(w_n221_9[1]),.doutc(w_n221_9[2]),.din(w_n221_2[2]));
	jspl3 jspl3_w_n221_10(.douta(w_n221_10[0]),.doutb(w_n221_10[1]),.doutc(w_n221_10[2]),.din(w_n221_3[0]));
	jspl3 jspl3_w_n221_11(.douta(w_n221_11[0]),.doutb(w_n221_11[1]),.doutc(w_n221_11[2]),.din(w_n221_3[1]));
	jspl3 jspl3_w_n221_12(.douta(w_n221_12[0]),.doutb(w_n221_12[1]),.doutc(w_n221_12[2]),.din(w_n221_3[2]));
	jspl3 jspl3_w_n221_13(.douta(w_n221_13[0]),.doutb(w_n221_13[1]),.doutc(w_n221_13[2]),.din(w_n221_4[0]));
	jspl3 jspl3_w_n221_14(.douta(w_n221_14[0]),.doutb(w_n221_14[1]),.doutc(w_n221_14[2]),.din(w_n221_4[1]));
	jspl3 jspl3_w_n221_15(.douta(w_n221_15[0]),.doutb(w_n221_15[1]),.doutc(w_n221_15[2]),.din(w_n221_4[2]));
	jspl3 jspl3_w_n221_16(.douta(w_n221_16[0]),.doutb(w_n221_16[1]),.doutc(w_n221_16[2]),.din(w_n221_5[0]));
	jspl3 jspl3_w_n221_17(.douta(w_n221_17[0]),.doutb(w_n221_17[1]),.doutc(w_n221_17[2]),.din(w_n221_5[1]));
	jspl3 jspl3_w_n221_18(.douta(w_n221_18[0]),.doutb(w_n221_18[1]),.doutc(w_n221_18[2]),.din(w_n221_5[2]));
	jspl3 jspl3_w_n221_19(.douta(w_n221_19[0]),.doutb(w_n221_19[1]),.doutc(w_n221_19[2]),.din(w_n221_6[0]));
	jspl3 jspl3_w_n221_20(.douta(w_n221_20[0]),.doutb(w_n221_20[1]),.doutc(w_n221_20[2]),.din(w_n221_6[1]));
	jspl3 jspl3_w_n221_21(.douta(w_n221_21[0]),.doutb(w_n221_21[1]),.doutc(w_n221_21[2]),.din(w_n221_6[2]));
	jspl3 jspl3_w_n221_22(.douta(w_n221_22[0]),.doutb(w_n221_22[1]),.doutc(w_n221_22[2]),.din(w_n221_7[0]));
	jspl3 jspl3_w_n221_23(.douta(w_n221_23[0]),.doutb(w_n221_23[1]),.doutc(w_n221_23[2]),.din(w_n221_7[1]));
	jspl3 jspl3_w_n221_24(.douta(w_n221_24[0]),.doutb(w_n221_24[1]),.doutc(w_n221_24[2]),.din(w_n221_7[2]));
	jspl3 jspl3_w_n221_25(.douta(w_n221_25[0]),.doutb(w_n221_25[1]),.doutc(w_n221_25[2]),.din(w_n221_8[0]));
	jspl3 jspl3_w_n221_26(.douta(w_n221_26[0]),.doutb(w_n221_26[1]),.doutc(w_n221_26[2]),.din(w_n221_8[1]));
	jspl3 jspl3_w_n221_27(.douta(w_n221_27[0]),.doutb(w_n221_27[1]),.doutc(w_n221_27[2]),.din(w_n221_8[2]));
	jspl3 jspl3_w_n221_28(.douta(w_n221_28[0]),.doutb(w_n221_28[1]),.doutc(w_n221_28[2]),.din(w_n221_9[0]));
	jspl3 jspl3_w_n221_29(.douta(w_n221_29[0]),.doutb(w_n221_29[1]),.doutc(w_n221_29[2]),.din(w_n221_9[1]));
	jspl3 jspl3_w_n221_30(.douta(w_n221_30[0]),.doutb(w_n221_30[1]),.doutc(w_n221_30[2]),.din(w_n221_9[2]));
	jspl3 jspl3_w_n221_31(.douta(w_n221_31[0]),.doutb(w_n221_31[1]),.doutc(w_n221_31[2]),.din(w_n221_10[0]));
	jspl3 jspl3_w_n221_32(.douta(w_n221_32[0]),.doutb(w_n221_32[1]),.doutc(w_n221_32[2]),.din(w_n221_10[1]));
	jspl3 jspl3_w_n221_33(.douta(w_n221_33[0]),.doutb(w_n221_33[1]),.doutc(w_n221_33[2]),.din(w_n221_10[2]));
	jspl3 jspl3_w_n221_34(.douta(w_n221_34[0]),.doutb(w_n221_34[1]),.doutc(w_n221_34[2]),.din(w_n221_11[0]));
	jspl3 jspl3_w_n221_35(.douta(w_n221_35[0]),.doutb(w_n221_35[1]),.doutc(w_n221_35[2]),.din(w_n221_11[1]));
	jspl3 jspl3_w_n221_36(.douta(w_n221_36[0]),.doutb(w_n221_36[1]),.doutc(w_n221_36[2]),.din(w_n221_11[2]));
	jspl3 jspl3_w_n221_37(.douta(w_n221_37[0]),.doutb(w_n221_37[1]),.doutc(w_n221_37[2]),.din(w_n221_12[0]));
	jspl3 jspl3_w_n221_38(.douta(w_n221_38[0]),.doutb(w_n221_38[1]),.doutc(w_n221_38[2]),.din(w_n221_12[1]));
	jspl3 jspl3_w_n221_39(.douta(w_n221_39[0]),.doutb(w_n221_39[1]),.doutc(w_n221_39[2]),.din(w_n221_12[2]));
	jspl3 jspl3_w_n221_40(.douta(w_n221_40[0]),.doutb(w_n221_40[1]),.doutc(w_n221_40[2]),.din(w_n221_13[0]));
	jspl3 jspl3_w_n221_41(.douta(w_n221_41[0]),.doutb(w_n221_41[1]),.doutc(w_n221_41[2]),.din(w_n221_13[1]));
	jspl3 jspl3_w_n221_42(.douta(w_n221_42[0]),.doutb(w_n221_42[1]),.doutc(w_n221_42[2]),.din(w_n221_13[2]));
	jspl3 jspl3_w_n221_43(.douta(w_n221_43[0]),.doutb(w_n221_43[1]),.doutc(w_n221_43[2]),.din(w_n221_14[0]));
	jspl3 jspl3_w_n221_44(.douta(w_n221_44[0]),.doutb(w_n221_44[1]),.doutc(w_n221_44[2]),.din(w_n221_14[1]));
	jspl3 jspl3_w_n221_45(.douta(w_n221_45[0]),.doutb(w_n221_45[1]),.doutc(w_n221_45[2]),.din(w_n221_14[2]));
	jspl3 jspl3_w_n221_46(.douta(w_n221_46[0]),.doutb(w_n221_46[1]),.doutc(w_n221_46[2]),.din(w_n221_15[0]));
	jspl3 jspl3_w_n221_47(.douta(w_n221_47[0]),.doutb(w_n221_47[1]),.doutc(w_n221_47[2]),.din(w_n221_15[1]));
	jspl3 jspl3_w_n221_48(.douta(w_n221_48[0]),.doutb(w_n221_48[1]),.doutc(w_n221_48[2]),.din(w_n221_15[2]));
	jspl3 jspl3_w_n221_49(.douta(w_n221_49[0]),.doutb(w_n221_49[1]),.doutc(w_n221_49[2]),.din(w_n221_16[0]));
	jspl3 jspl3_w_n221_50(.douta(w_n221_50[0]),.doutb(w_n221_50[1]),.doutc(w_n221_50[2]),.din(w_n221_16[1]));
	jspl3 jspl3_w_n221_51(.douta(w_n221_51[0]),.doutb(w_n221_51[1]),.doutc(w_n221_51[2]),.din(w_n221_16[2]));
	jspl3 jspl3_w_n221_52(.douta(w_n221_52[0]),.doutb(w_n221_52[1]),.doutc(w_n221_52[2]),.din(w_n221_17[0]));
	jspl3 jspl3_w_n221_53(.douta(w_n221_53[0]),.doutb(w_n221_53[1]),.doutc(w_n221_53[2]),.din(w_n221_17[1]));
	jspl3 jspl3_w_n221_54(.douta(w_n221_54[0]),.doutb(w_n221_54[1]),.doutc(w_n221_54[2]),.din(w_n221_17[2]));
	jspl3 jspl3_w_n221_55(.douta(w_n221_55[0]),.doutb(w_n221_55[1]),.doutc(w_n221_55[2]),.din(w_n221_18[0]));
	jspl3 jspl3_w_n221_56(.douta(w_n221_56[0]),.doutb(w_n221_56[1]),.doutc(w_n221_56[2]),.din(w_n221_18[1]));
	jspl3 jspl3_w_n221_57(.douta(w_n221_57[0]),.doutb(w_n221_57[1]),.doutc(w_n221_57[2]),.din(w_n221_18[2]));
	jspl3 jspl3_w_n221_58(.douta(w_n221_58[0]),.doutb(w_n221_58[1]),.doutc(w_n221_58[2]),.din(w_n221_19[0]));
	jspl3 jspl3_w_n221_59(.douta(w_n221_59[0]),.doutb(w_n221_59[1]),.doutc(w_n221_59[2]),.din(w_n221_19[1]));
	jspl3 jspl3_w_n221_60(.douta(w_n221_60[0]),.doutb(w_n221_60[1]),.doutc(w_n221_60[2]),.din(w_n221_19[2]));
	jspl3 jspl3_w_n221_61(.douta(w_n221_61[0]),.doutb(w_n221_61[1]),.doutc(w_n221_61[2]),.din(w_n221_20[0]));
	jspl3 jspl3_w_n221_62(.douta(w_n221_62[0]),.doutb(w_n221_62[1]),.doutc(w_n221_62[2]),.din(w_n221_20[1]));
	jspl3 jspl3_w_n221_63(.douta(w_n221_63[0]),.doutb(w_n221_63[1]),.doutc(w_n221_63[2]),.din(w_n221_20[2]));
	jspl3 jspl3_w_n221_64(.douta(w_n221_64[0]),.doutb(w_n221_64[1]),.doutc(w_n221_64[2]),.din(w_n221_21[0]));
	jspl3 jspl3_w_n221_65(.douta(w_n221_65[0]),.doutb(w_n221_65[1]),.doutc(w_n221_65[2]),.din(w_n221_21[1]));
	jspl3 jspl3_w_n221_66(.douta(w_n221_66[0]),.doutb(w_n221_66[1]),.doutc(w_n221_66[2]),.din(w_n221_21[2]));
	jspl3 jspl3_w_n221_67(.douta(w_n221_67[0]),.doutb(w_n221_67[1]),.doutc(w_n221_67[2]),.din(w_n221_22[0]));
	jspl3 jspl3_w_n221_68(.douta(w_n221_68[0]),.doutb(w_n221_68[1]),.doutc(w_n221_68[2]),.din(w_n221_22[1]));
	jspl3 jspl3_w_n221_69(.douta(w_n221_69[0]),.doutb(w_n221_69[1]),.doutc(w_n221_69[2]),.din(w_n221_22[2]));
	jspl3 jspl3_w_n221_70(.douta(w_n221_70[0]),.doutb(w_n221_70[1]),.doutc(w_n221_70[2]),.din(w_n221_23[0]));
	jspl3 jspl3_w_n221_71(.douta(w_n221_71[0]),.doutb(w_n221_71[1]),.doutc(w_n221_71[2]),.din(w_n221_23[1]));
	jspl3 jspl3_w_n221_72(.douta(w_n221_72[0]),.doutb(w_n221_72[1]),.doutc(w_n221_72[2]),.din(w_n221_23[2]));
	jspl3 jspl3_w_n221_73(.douta(w_n221_73[0]),.doutb(w_n221_73[1]),.doutc(w_n221_73[2]),.din(w_n221_24[0]));
	jspl3 jspl3_w_n221_74(.douta(w_n221_74[0]),.doutb(w_n221_74[1]),.doutc(w_n221_74[2]),.din(w_n221_24[1]));
	jspl3 jspl3_w_n221_75(.douta(w_n221_75[0]),.doutb(w_n221_75[1]),.doutc(w_n221_75[2]),.din(w_n221_24[2]));
	jspl jspl_w_n221_76(.douta(w_n221_76[0]),.doutb(w_n221_76[1]),.din(w_n221_25[0]));
	jspl jspl_w_n224_0(.douta(w_n224_0[0]),.doutb(w_n224_0[1]),.din(n224));
	jspl jspl_w_n225_0(.douta(w_n225_0[0]),.doutb(w_n225_0[1]),.din(n225));
	jspl jspl_w_n234_0(.douta(w_n234_0[0]),.doutb(w_n234_0[1]),.din(n234));
	jspl jspl_w_n235_0(.douta(w_n235_0[0]),.doutb(w_n235_0[1]),.din(n235));
	jspl jspl_w_n236_0(.douta(w_n236_0[0]),.doutb(w_n236_0[1]),.din(n236));
	jspl3 jspl3_w_n239_0(.douta(w_n239_0[0]),.doutb(w_n239_0[1]),.doutc(w_n239_0[2]),.din(n239));
	jspl3 jspl3_w_n239_1(.douta(w_n239_1[0]),.doutb(w_n239_1[1]),.doutc(w_n239_1[2]),.din(w_n239_0[0]));
	jspl3 jspl3_w_n239_2(.douta(w_n239_2[0]),.doutb(w_n239_2[1]),.doutc(w_n239_2[2]),.din(w_n239_0[1]));
	jspl3 jspl3_w_n239_3(.douta(w_n239_3[0]),.doutb(w_n239_3[1]),.doutc(w_n239_3[2]),.din(w_n239_0[2]));
	jspl3 jspl3_w_n239_4(.douta(w_n239_4[0]),.doutb(w_n239_4[1]),.doutc(w_n239_4[2]),.din(w_n239_1[0]));
	jspl3 jspl3_w_n239_5(.douta(w_n239_5[0]),.doutb(w_n239_5[1]),.doutc(w_n239_5[2]),.din(w_n239_1[1]));
	jspl3 jspl3_w_n239_6(.douta(w_n239_6[0]),.doutb(w_n239_6[1]),.doutc(w_n239_6[2]),.din(w_n239_1[2]));
	jspl3 jspl3_w_n239_7(.douta(w_n239_7[0]),.doutb(w_n239_7[1]),.doutc(w_n239_7[2]),.din(w_n239_2[0]));
	jspl3 jspl3_w_n239_8(.douta(w_n239_8[0]),.doutb(w_n239_8[1]),.doutc(w_n239_8[2]),.din(w_n239_2[1]));
	jspl3 jspl3_w_n239_9(.douta(w_n239_9[0]),.doutb(w_n239_9[1]),.doutc(w_n239_9[2]),.din(w_n239_2[2]));
	jspl3 jspl3_w_n239_10(.douta(w_n239_10[0]),.doutb(w_n239_10[1]),.doutc(w_n239_10[2]),.din(w_n239_3[0]));
	jspl3 jspl3_w_n239_11(.douta(w_n239_11[0]),.doutb(w_n239_11[1]),.doutc(w_n239_11[2]),.din(w_n239_3[1]));
	jspl3 jspl3_w_n239_12(.douta(w_n239_12[0]),.doutb(w_n239_12[1]),.doutc(w_n239_12[2]),.din(w_n239_3[2]));
	jspl3 jspl3_w_n239_13(.douta(w_n239_13[0]),.doutb(w_n239_13[1]),.doutc(w_n239_13[2]),.din(w_n239_4[0]));
	jspl3 jspl3_w_n239_14(.douta(w_n239_14[0]),.doutb(w_n239_14[1]),.doutc(w_n239_14[2]),.din(w_n239_4[1]));
	jspl3 jspl3_w_n239_15(.douta(w_n239_15[0]),.doutb(w_n239_15[1]),.doutc(w_n239_15[2]),.din(w_n239_4[2]));
	jspl3 jspl3_w_n239_16(.douta(w_n239_16[0]),.doutb(w_n239_16[1]),.doutc(w_n239_16[2]),.din(w_n239_5[0]));
	jspl3 jspl3_w_n239_17(.douta(w_n239_17[0]),.doutb(w_n239_17[1]),.doutc(w_n239_17[2]),.din(w_n239_5[1]));
	jspl3 jspl3_w_n239_18(.douta(w_n239_18[0]),.doutb(w_n239_18[1]),.doutc(w_n239_18[2]),.din(w_n239_5[2]));
	jspl3 jspl3_w_n239_19(.douta(w_n239_19[0]),.doutb(w_n239_19[1]),.doutc(w_n239_19[2]),.din(w_n239_6[0]));
	jspl3 jspl3_w_n239_20(.douta(w_n239_20[0]),.doutb(w_n239_20[1]),.doutc(w_n239_20[2]),.din(w_n239_6[1]));
	jspl3 jspl3_w_n239_21(.douta(w_n239_21[0]),.doutb(w_n239_21[1]),.doutc(w_n239_21[2]),.din(w_n239_6[2]));
	jspl3 jspl3_w_n239_22(.douta(w_n239_22[0]),.doutb(w_n239_22[1]),.doutc(w_n239_22[2]),.din(w_n239_7[0]));
	jspl3 jspl3_w_n239_23(.douta(w_n239_23[0]),.doutb(w_n239_23[1]),.doutc(w_n239_23[2]),.din(w_n239_7[1]));
	jspl3 jspl3_w_n239_24(.douta(w_n239_24[0]),.doutb(w_n239_24[1]),.doutc(w_n239_24[2]),.din(w_n239_7[2]));
	jspl3 jspl3_w_n239_25(.douta(w_n239_25[0]),.doutb(w_n239_25[1]),.doutc(w_n239_25[2]),.din(w_n239_8[0]));
	jspl3 jspl3_w_n239_26(.douta(w_n239_26[0]),.doutb(w_n239_26[1]),.doutc(w_n239_26[2]),.din(w_n239_8[1]));
	jspl3 jspl3_w_n239_27(.douta(w_n239_27[0]),.doutb(w_n239_27[1]),.doutc(w_n239_27[2]),.din(w_n239_8[2]));
	jspl3 jspl3_w_n239_28(.douta(w_n239_28[0]),.doutb(w_n239_28[1]),.doutc(w_n239_28[2]),.din(w_n239_9[0]));
	jspl3 jspl3_w_n239_29(.douta(w_n239_29[0]),.doutb(w_n239_29[1]),.doutc(w_n239_29[2]),.din(w_n239_9[1]));
	jspl3 jspl3_w_n239_30(.douta(w_n239_30[0]),.doutb(w_n239_30[1]),.doutc(w_n239_30[2]),.din(w_n239_9[2]));
	jspl3 jspl3_w_n239_31(.douta(w_n239_31[0]),.doutb(w_n239_31[1]),.doutc(w_n239_31[2]),.din(w_n239_10[0]));
	jspl3 jspl3_w_n239_32(.douta(w_n239_32[0]),.doutb(w_n239_32[1]),.doutc(w_n239_32[2]),.din(w_n239_10[1]));
	jspl3 jspl3_w_n239_33(.douta(w_n239_33[0]),.doutb(w_n239_33[1]),.doutc(w_n239_33[2]),.din(w_n239_10[2]));
	jspl3 jspl3_w_n239_34(.douta(w_n239_34[0]),.doutb(w_n239_34[1]),.doutc(w_n239_34[2]),.din(w_n239_11[0]));
	jspl3 jspl3_w_n239_35(.douta(w_n239_35[0]),.doutb(w_n239_35[1]),.doutc(w_n239_35[2]),.din(w_n239_11[1]));
	jspl3 jspl3_w_n239_36(.douta(w_n239_36[0]),.doutb(w_n239_36[1]),.doutc(w_n239_36[2]),.din(w_n239_11[2]));
	jspl3 jspl3_w_n239_37(.douta(w_n239_37[0]),.doutb(w_n239_37[1]),.doutc(w_n239_37[2]),.din(w_n239_12[0]));
	jspl3 jspl3_w_n239_38(.douta(w_n239_38[0]),.doutb(w_n239_38[1]),.doutc(w_n239_38[2]),.din(w_n239_12[1]));
	jspl3 jspl3_w_n239_39(.douta(w_n239_39[0]),.doutb(w_n239_39[1]),.doutc(w_n239_39[2]),.din(w_n239_12[2]));
	jspl3 jspl3_w_n239_40(.douta(w_n239_40[0]),.doutb(w_n239_40[1]),.doutc(w_n239_40[2]),.din(w_n239_13[0]));
	jspl3 jspl3_w_n239_41(.douta(w_n239_41[0]),.doutb(w_n239_41[1]),.doutc(w_n239_41[2]),.din(w_n239_13[1]));
	jspl3 jspl3_w_n239_42(.douta(w_n239_42[0]),.doutb(w_n239_42[1]),.doutc(w_n239_42[2]),.din(w_n239_13[2]));
	jspl3 jspl3_w_n239_43(.douta(w_n239_43[0]),.doutb(w_n239_43[1]),.doutc(w_n239_43[2]),.din(w_n239_14[0]));
	jspl3 jspl3_w_n239_44(.douta(w_n239_44[0]),.doutb(w_n239_44[1]),.doutc(w_n239_44[2]),.din(w_n239_14[1]));
	jspl3 jspl3_w_n239_45(.douta(w_n239_45[0]),.doutb(w_n239_45[1]),.doutc(w_n239_45[2]),.din(w_n239_14[2]));
	jspl3 jspl3_w_n239_46(.douta(w_n239_46[0]),.doutb(w_n239_46[1]),.doutc(w_n239_46[2]),.din(w_n239_15[0]));
	jspl3 jspl3_w_n239_47(.douta(w_n239_47[0]),.doutb(w_n239_47[1]),.doutc(w_n239_47[2]),.din(w_n239_15[1]));
	jspl3 jspl3_w_n239_48(.douta(w_n239_48[0]),.doutb(w_n239_48[1]),.doutc(w_n239_48[2]),.din(w_n239_15[2]));
	jspl3 jspl3_w_n239_49(.douta(w_n239_49[0]),.doutb(w_n239_49[1]),.doutc(w_n239_49[2]),.din(w_n239_16[0]));
	jspl3 jspl3_w_n239_50(.douta(w_n239_50[0]),.doutb(w_n239_50[1]),.doutc(w_n239_50[2]),.din(w_n239_16[1]));
	jspl3 jspl3_w_n239_51(.douta(w_n239_51[0]),.doutb(w_n239_51[1]),.doutc(w_n239_51[2]),.din(w_n239_16[2]));
	jspl3 jspl3_w_n239_52(.douta(w_n239_52[0]),.doutb(w_n239_52[1]),.doutc(w_n239_52[2]),.din(w_n239_17[0]));
	jspl3 jspl3_w_n239_53(.douta(w_n239_53[0]),.doutb(w_n239_53[1]),.doutc(w_n239_53[2]),.din(w_n239_17[1]));
	jspl3 jspl3_w_n239_54(.douta(w_n239_54[0]),.doutb(w_n239_54[1]),.doutc(w_n239_54[2]),.din(w_n239_17[2]));
	jspl3 jspl3_w_n239_55(.douta(w_n239_55[0]),.doutb(w_n239_55[1]),.doutc(w_n239_55[2]),.din(w_n239_18[0]));
	jspl3 jspl3_w_n239_56(.douta(w_n239_56[0]),.doutb(w_n239_56[1]),.doutc(w_n239_56[2]),.din(w_n239_18[1]));
	jspl3 jspl3_w_n239_57(.douta(w_n239_57[0]),.doutb(w_n239_57[1]),.doutc(w_n239_57[2]),.din(w_n239_18[2]));
	jspl3 jspl3_w_n239_58(.douta(w_n239_58[0]),.doutb(w_n239_58[1]),.doutc(w_n239_58[2]),.din(w_n239_19[0]));
	jspl3 jspl3_w_n239_59(.douta(w_n239_59[0]),.doutb(w_n239_59[1]),.doutc(w_n239_59[2]),.din(w_n239_19[1]));
	jspl3 jspl3_w_n239_60(.douta(w_n239_60[0]),.doutb(w_n239_60[1]),.doutc(w_n239_60[2]),.din(w_n239_19[2]));
	jspl3 jspl3_w_n239_61(.douta(w_n239_61[0]),.doutb(w_n239_61[1]),.doutc(w_n239_61[2]),.din(w_n239_20[0]));
	jspl3 jspl3_w_n239_62(.douta(w_n239_62[0]),.doutb(w_n239_62[1]),.doutc(w_n239_62[2]),.din(w_n239_20[1]));
	jspl3 jspl3_w_n239_63(.douta(w_n239_63[0]),.doutb(w_n239_63[1]),.doutc(w_n239_63[2]),.din(w_n239_20[2]));
	jspl3 jspl3_w_n239_64(.douta(w_n239_64[0]),.doutb(w_n239_64[1]),.doutc(w_n239_64[2]),.din(w_n239_21[0]));
	jspl3 jspl3_w_n239_65(.douta(w_n239_65[0]),.doutb(w_n239_65[1]),.doutc(w_n239_65[2]),.din(w_n239_21[1]));
	jspl3 jspl3_w_n239_66(.douta(w_n239_66[0]),.doutb(w_n239_66[1]),.doutc(w_n239_66[2]),.din(w_n239_21[2]));
	jspl3 jspl3_w_n239_67(.douta(w_n239_67[0]),.doutb(w_n239_67[1]),.doutc(w_n239_67[2]),.din(w_n239_22[0]));
	jspl3 jspl3_w_n239_68(.douta(w_n239_68[0]),.doutb(w_n239_68[1]),.doutc(w_n239_68[2]),.din(w_n239_22[1]));
	jspl3 jspl3_w_n239_69(.douta(w_n239_69[0]),.doutb(w_n239_69[1]),.doutc(w_n239_69[2]),.din(w_n239_22[2]));
	jspl3 jspl3_w_n239_70(.douta(w_n239_70[0]),.doutb(w_n239_70[1]),.doutc(w_n239_70[2]),.din(w_n239_23[0]));
	jspl3 jspl3_w_n239_71(.douta(w_n239_71[0]),.doutb(w_n239_71[1]),.doutc(w_n239_71[2]),.din(w_n239_23[1]));
	jspl3 jspl3_w_n239_72(.douta(w_n239_72[0]),.doutb(w_n239_72[1]),.doutc(w_n239_72[2]),.din(w_n239_23[2]));
	jspl3 jspl3_w_n239_73(.douta(w_n239_73[0]),.doutb(w_n239_73[1]),.doutc(w_n239_73[2]),.din(w_n239_24[0]));
	jspl3 jspl3_w_n239_74(.douta(w_n239_74[0]),.doutb(w_n239_74[1]),.doutc(w_n239_74[2]),.din(w_n239_24[1]));
	jspl jspl_w_n239_75(.douta(w_n239_75[0]),.doutb(w_n239_75[1]),.din(w_n239_24[2]));
	jspl3 jspl3_w_n241_0(.douta(w_n241_0[0]),.doutb(w_n241_0[1]),.doutc(w_n241_0[2]),.din(n241));
	jspl3 jspl3_w_n241_1(.douta(w_n241_1[0]),.doutb(w_n241_1[1]),.doutc(w_n241_1[2]),.din(w_n241_0[0]));
	jspl jspl_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.din(n242));
	jspl3 jspl3_w_n243_0(.douta(w_n243_0[0]),.doutb(w_n243_0[1]),.doutc(w_n243_0[2]),.din(n243));
	jspl jspl_w_n244_0(.douta(w_n244_0[0]),.doutb(w_n244_0[1]),.din(n244));
	jspl3 jspl3_w_n246_0(.douta(w_n246_0[0]),.doutb(w_n246_0[1]),.doutc(w_n246_0[2]),.din(n246));
	jspl jspl_w_n247_0(.douta(w_n247_0[0]),.doutb(w_n247_0[1]),.din(n247));
	jspl jspl_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.din(n249));
	jspl jspl_w_n250_0(.douta(w_n250_0[0]),.doutb(w_n250_0[1]),.din(n250));
	jspl3 jspl3_w_n252_0(.douta(w_n252_0[0]),.doutb(w_n252_0[1]),.doutc(w_n252_0[2]),.din(n252));
	jspl3 jspl3_w_n256_0(.douta(w_n256_0[0]),.doutb(w_n256_0[1]),.doutc(w_n256_0[2]),.din(n256));
	jspl jspl_w_n256_1(.douta(w_n256_1[0]),.doutb(w_n256_1[1]),.din(w_n256_0[0]));
	jspl jspl_w_n260_0(.douta(w_n260_0[0]),.doutb(w_n260_0[1]),.din(n260));
	jspl jspl_w_n261_0(.douta(w_n261_0[0]),.doutb(w_n261_0[1]),.din(n261));
	jspl jspl_w_n264_0(.douta(w_n264_0[0]),.doutb(w_n264_0[1]),.din(n264));
	jspl3 jspl3_w_n267_0(.douta(w_n267_0[0]),.doutb(w_n267_0[1]),.doutc(w_n267_0[2]),.din(n267));
	jspl jspl_w_n267_1(.douta(w_n267_1[0]),.doutb(w_n267_1[1]),.din(w_n267_0[0]));
	jspl3 jspl3_w_n268_0(.douta(w_n268_0[0]),.doutb(w_n268_0[1]),.doutc(w_n268_0[2]),.din(n268));
	jspl jspl_w_n268_1(.douta(w_n268_1[0]),.doutb(w_n268_1[1]),.din(w_n268_0[0]));
	jspl jspl_w_n269_0(.douta(w_n269_0[0]),.doutb(w_n269_0[1]),.din(n269));
	jspl3 jspl3_w_n270_0(.douta(w_n270_0[0]),.doutb(w_n270_0[1]),.doutc(w_n270_0[2]),.din(n270));
	jspl jspl_w_n271_0(.douta(w_n271_0[0]),.doutb(w_n271_0[1]),.din(n271));
	jspl3 jspl3_w_n273_0(.douta(w_n273_0[0]),.doutb(w_n273_0[1]),.doutc(w_n273_0[2]),.din(n273));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_n274_0[1]),.din(n274));
	jspl jspl_w_n287_0(.douta(w_n287_0[0]),.doutb(w_n287_0[1]),.din(n287));
	jspl3 jspl3_w_n294_0(.douta(w_n294_0[0]),.doutb(w_n294_0[1]),.doutc(w_n294_0[2]),.din(n294));
	jspl3 jspl3_w_n294_1(.douta(w_n294_1[0]),.doutb(w_n294_1[1]),.doutc(w_n294_1[2]),.din(w_n294_0[0]));
	jspl3 jspl3_w_n294_2(.douta(w_n294_2[0]),.doutb(w_n294_2[1]),.doutc(w_n294_2[2]),.din(w_n294_0[1]));
	jspl3 jspl3_w_n294_3(.douta(w_n294_3[0]),.doutb(w_n294_3[1]),.doutc(w_n294_3[2]),.din(w_n294_0[2]));
	jspl3 jspl3_w_n294_4(.douta(w_n294_4[0]),.doutb(w_n294_4[1]),.doutc(w_n294_4[2]),.din(w_n294_1[0]));
	jspl3 jspl3_w_n294_5(.douta(w_n294_5[0]),.doutb(w_n294_5[1]),.doutc(w_n294_5[2]),.din(w_n294_1[1]));
	jspl3 jspl3_w_n294_6(.douta(w_n294_6[0]),.doutb(w_n294_6[1]),.doutc(w_n294_6[2]),.din(w_n294_1[2]));
	jspl3 jspl3_w_n294_7(.douta(w_n294_7[0]),.doutb(w_n294_7[1]),.doutc(w_n294_7[2]),.din(w_n294_2[0]));
	jspl3 jspl3_w_n294_8(.douta(w_n294_8[0]),.doutb(w_n294_8[1]),.doutc(w_n294_8[2]),.din(w_n294_2[1]));
	jspl3 jspl3_w_n294_9(.douta(w_n294_9[0]),.doutb(w_n294_9[1]),.doutc(w_n294_9[2]),.din(w_n294_2[2]));
	jspl3 jspl3_w_n294_10(.douta(w_n294_10[0]),.doutb(w_n294_10[1]),.doutc(w_n294_10[2]),.din(w_n294_3[0]));
	jspl3 jspl3_w_n294_11(.douta(w_n294_11[0]),.doutb(w_n294_11[1]),.doutc(w_n294_11[2]),.din(w_n294_3[1]));
	jspl3 jspl3_w_n294_12(.douta(w_n294_12[0]),.doutb(w_n294_12[1]),.doutc(w_n294_12[2]),.din(w_n294_3[2]));
	jspl3 jspl3_w_n294_13(.douta(w_n294_13[0]),.doutb(w_n294_13[1]),.doutc(w_n294_13[2]),.din(w_n294_4[0]));
	jspl3 jspl3_w_n294_14(.douta(w_n294_14[0]),.doutb(w_n294_14[1]),.doutc(w_n294_14[2]),.din(w_n294_4[1]));
	jspl3 jspl3_w_n294_15(.douta(w_n294_15[0]),.doutb(w_n294_15[1]),.doutc(w_n294_15[2]),.din(w_n294_4[2]));
	jspl3 jspl3_w_n294_16(.douta(w_n294_16[0]),.doutb(w_n294_16[1]),.doutc(w_n294_16[2]),.din(w_n294_5[0]));
	jspl3 jspl3_w_n294_17(.douta(w_n294_17[0]),.doutb(w_n294_17[1]),.doutc(w_n294_17[2]),.din(w_n294_5[1]));
	jspl3 jspl3_w_n294_18(.douta(w_n294_18[0]),.doutb(w_n294_18[1]),.doutc(w_n294_18[2]),.din(w_n294_5[2]));
	jspl3 jspl3_w_n294_19(.douta(w_n294_19[0]),.doutb(w_n294_19[1]),.doutc(w_n294_19[2]),.din(w_n294_6[0]));
	jspl3 jspl3_w_n294_20(.douta(w_n294_20[0]),.doutb(w_n294_20[1]),.doutc(w_n294_20[2]),.din(w_n294_6[1]));
	jspl3 jspl3_w_n294_21(.douta(w_n294_21[0]),.doutb(w_n294_21[1]),.doutc(w_n294_21[2]),.din(w_n294_6[2]));
	jspl3 jspl3_w_n294_22(.douta(w_n294_22[0]),.doutb(w_n294_22[1]),.doutc(w_n294_22[2]),.din(w_n294_7[0]));
	jspl3 jspl3_w_n294_23(.douta(w_n294_23[0]),.doutb(w_n294_23[1]),.doutc(w_n294_23[2]),.din(w_n294_7[1]));
	jspl3 jspl3_w_n294_24(.douta(w_n294_24[0]),.doutb(w_n294_24[1]),.doutc(w_n294_24[2]),.din(w_n294_7[2]));
	jspl3 jspl3_w_n294_25(.douta(w_n294_25[0]),.doutb(w_n294_25[1]),.doutc(w_n294_25[2]),.din(w_n294_8[0]));
	jspl3 jspl3_w_n294_26(.douta(w_n294_26[0]),.doutb(w_n294_26[1]),.doutc(w_n294_26[2]),.din(w_n294_8[1]));
	jspl3 jspl3_w_n294_27(.douta(w_n294_27[0]),.doutb(w_n294_27[1]),.doutc(w_n294_27[2]),.din(w_n294_8[2]));
	jspl3 jspl3_w_n294_28(.douta(w_n294_28[0]),.doutb(w_n294_28[1]),.doutc(w_n294_28[2]),.din(w_n294_9[0]));
	jspl3 jspl3_w_n294_29(.douta(w_n294_29[0]),.doutb(w_n294_29[1]),.doutc(w_n294_29[2]),.din(w_n294_9[1]));
	jspl3 jspl3_w_n294_30(.douta(w_n294_30[0]),.doutb(w_n294_30[1]),.doutc(w_n294_30[2]),.din(w_n294_9[2]));
	jspl3 jspl3_w_n294_31(.douta(w_n294_31[0]),.doutb(w_n294_31[1]),.doutc(w_n294_31[2]),.din(w_n294_10[0]));
	jspl3 jspl3_w_n294_32(.douta(w_n294_32[0]),.doutb(w_n294_32[1]),.doutc(w_n294_32[2]),.din(w_n294_10[1]));
	jspl3 jspl3_w_n294_33(.douta(w_n294_33[0]),.doutb(w_n294_33[1]),.doutc(w_n294_33[2]),.din(w_n294_10[2]));
	jspl3 jspl3_w_n294_34(.douta(w_n294_34[0]),.doutb(w_n294_34[1]),.doutc(w_n294_34[2]),.din(w_n294_11[0]));
	jspl3 jspl3_w_n294_35(.douta(w_n294_35[0]),.doutb(w_n294_35[1]),.doutc(w_n294_35[2]),.din(w_n294_11[1]));
	jspl3 jspl3_w_n294_36(.douta(w_n294_36[0]),.doutb(w_n294_36[1]),.doutc(w_n294_36[2]),.din(w_n294_11[2]));
	jspl3 jspl3_w_n294_37(.douta(w_n294_37[0]),.doutb(w_n294_37[1]),.doutc(w_n294_37[2]),.din(w_n294_12[0]));
	jspl3 jspl3_w_n294_38(.douta(w_n294_38[0]),.doutb(w_n294_38[1]),.doutc(w_n294_38[2]),.din(w_n294_12[1]));
	jspl3 jspl3_w_n294_39(.douta(w_n294_39[0]),.doutb(w_n294_39[1]),.doutc(w_n294_39[2]),.din(w_n294_12[2]));
	jspl3 jspl3_w_n294_40(.douta(w_n294_40[0]),.doutb(w_n294_40[1]),.doutc(w_n294_40[2]),.din(w_n294_13[0]));
	jspl3 jspl3_w_n294_41(.douta(w_n294_41[0]),.doutb(w_n294_41[1]),.doutc(w_n294_41[2]),.din(w_n294_13[1]));
	jspl3 jspl3_w_n294_42(.douta(w_n294_42[0]),.doutb(w_n294_42[1]),.doutc(w_n294_42[2]),.din(w_n294_13[2]));
	jspl3 jspl3_w_n294_43(.douta(w_n294_43[0]),.doutb(w_n294_43[1]),.doutc(w_n294_43[2]),.din(w_n294_14[0]));
	jspl3 jspl3_w_n294_44(.douta(w_n294_44[0]),.doutb(w_n294_44[1]),.doutc(w_n294_44[2]),.din(w_n294_14[1]));
	jspl3 jspl3_w_n294_45(.douta(w_n294_45[0]),.doutb(w_n294_45[1]),.doutc(w_n294_45[2]),.din(w_n294_14[2]));
	jspl3 jspl3_w_n294_46(.douta(w_n294_46[0]),.doutb(w_n294_46[1]),.doutc(w_n294_46[2]),.din(w_n294_15[0]));
	jspl3 jspl3_w_n294_47(.douta(w_n294_47[0]),.doutb(w_n294_47[1]),.doutc(w_n294_47[2]),.din(w_n294_15[1]));
	jspl3 jspl3_w_n294_48(.douta(w_n294_48[0]),.doutb(w_n294_48[1]),.doutc(w_n294_48[2]),.din(w_n294_15[2]));
	jspl3 jspl3_w_n294_49(.douta(w_n294_49[0]),.doutb(w_n294_49[1]),.doutc(w_n294_49[2]),.din(w_n294_16[0]));
	jspl3 jspl3_w_n294_50(.douta(w_n294_50[0]),.doutb(w_n294_50[1]),.doutc(w_n294_50[2]),.din(w_n294_16[1]));
	jspl3 jspl3_w_n294_51(.douta(w_n294_51[0]),.doutb(w_n294_51[1]),.doutc(w_n294_51[2]),.din(w_n294_16[2]));
	jspl3 jspl3_w_n294_52(.douta(w_n294_52[0]),.doutb(w_n294_52[1]),.doutc(w_n294_52[2]),.din(w_n294_17[0]));
	jspl3 jspl3_w_n294_53(.douta(w_n294_53[0]),.doutb(w_n294_53[1]),.doutc(w_n294_53[2]),.din(w_n294_17[1]));
	jspl3 jspl3_w_n294_54(.douta(w_n294_54[0]),.doutb(w_n294_54[1]),.doutc(w_n294_54[2]),.din(w_n294_17[2]));
	jspl3 jspl3_w_n294_55(.douta(w_n294_55[0]),.doutb(w_n294_55[1]),.doutc(w_n294_55[2]),.din(w_n294_18[0]));
	jspl3 jspl3_w_n294_56(.douta(w_n294_56[0]),.doutb(w_n294_56[1]),.doutc(w_n294_56[2]),.din(w_n294_18[1]));
	jspl3 jspl3_w_n294_57(.douta(w_n294_57[0]),.doutb(w_n294_57[1]),.doutc(w_n294_57[2]),.din(w_n294_18[2]));
	jspl3 jspl3_w_n294_58(.douta(w_n294_58[0]),.doutb(w_n294_58[1]),.doutc(w_n294_58[2]),.din(w_n294_19[0]));
	jspl3 jspl3_w_n294_59(.douta(w_n294_59[0]),.doutb(w_n294_59[1]),.doutc(w_n294_59[2]),.din(w_n294_19[1]));
	jspl3 jspl3_w_n294_60(.douta(w_n294_60[0]),.doutb(w_n294_60[1]),.doutc(w_n294_60[2]),.din(w_n294_19[2]));
	jspl3 jspl3_w_n294_61(.douta(w_n294_61[0]),.doutb(w_n294_61[1]),.doutc(w_n294_61[2]),.din(w_n294_20[0]));
	jspl3 jspl3_w_n294_62(.douta(w_n294_62[0]),.doutb(w_n294_62[1]),.doutc(w_n294_62[2]),.din(w_n294_20[1]));
	jspl3 jspl3_w_n294_63(.douta(w_n294_63[0]),.doutb(w_n294_63[1]),.doutc(w_n294_63[2]),.din(w_n294_20[2]));
	jspl3 jspl3_w_n294_64(.douta(w_n294_64[0]),.doutb(w_n294_64[1]),.doutc(w_n294_64[2]),.din(w_n294_21[0]));
	jspl3 jspl3_w_n294_65(.douta(w_n294_65[0]),.doutb(w_n294_65[1]),.doutc(w_n294_65[2]),.din(w_n294_21[1]));
	jspl3 jspl3_w_n294_66(.douta(w_n294_66[0]),.doutb(w_n294_66[1]),.doutc(w_n294_66[2]),.din(w_n294_21[2]));
	jspl3 jspl3_w_n294_67(.douta(w_n294_67[0]),.doutb(w_n294_67[1]),.doutc(w_n294_67[2]),.din(w_n294_22[0]));
	jspl3 jspl3_w_n294_68(.douta(w_n294_68[0]),.doutb(w_n294_68[1]),.doutc(w_n294_68[2]),.din(w_n294_22[1]));
	jspl3 jspl3_w_n294_69(.douta(w_n294_69[0]),.doutb(w_n294_69[1]),.doutc(w_n294_69[2]),.din(w_n294_22[2]));
	jspl3 jspl3_w_n294_70(.douta(w_n294_70[0]),.doutb(w_n294_70[1]),.doutc(w_n294_70[2]),.din(w_n294_23[0]));
	jspl3 jspl3_w_n294_71(.douta(w_n294_71[0]),.doutb(w_n294_71[1]),.doutc(w_n294_71[2]),.din(w_n294_23[1]));
	jspl3 jspl3_w_n294_72(.douta(w_n294_72[0]),.doutb(w_n294_72[1]),.doutc(w_n294_72[2]),.din(w_n294_23[2]));
	jspl3 jspl3_w_n294_73(.douta(w_n294_73[0]),.doutb(w_n294_73[1]),.doutc(w_n294_73[2]),.din(w_n294_24[0]));
	jspl3 jspl3_w_n294_74(.douta(w_n294_74[0]),.doutb(w_n294_74[1]),.doutc(w_n294_74[2]),.din(w_n294_24[1]));
	jspl jspl_w_n294_75(.douta(w_n294_75[0]),.doutb(w_n294_75[1]),.din(w_n294_24[2]));
	jspl jspl_w_n295_0(.douta(w_n295_0[0]),.doutb(w_n295_0[1]),.din(n295));
	jspl3 jspl3_w_n298_0(.douta(w_n298_0[0]),.doutb(w_n298_0[1]),.doutc(w_n298_0[2]),.din(n298));
	jspl jspl_w_n299_0(.douta(w_n299_0[0]),.doutb(w_n299_0[1]),.din(n299));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.din(n303));
	jspl jspl_w_n304_0(.douta(w_n304_0[0]),.doutb(w_n304_0[1]),.din(n304));
	jspl jspl_w_n306_0(.douta(w_n306_0[0]),.doutb(w_n306_0[1]),.din(n306));
	jspl jspl_w_n307_0(.douta(w_n307_0[0]),.doutb(w_n307_0[1]),.din(n307));
	jspl jspl_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.din(n308));
	jspl jspl_w_n321_0(.douta(w_n321_0[0]),.doutb(w_n321_0[1]),.din(n321));
	jspl jspl_w_n329_0(.douta(w_n329_0[0]),.doutb(w_n329_0[1]),.din(n329));
	jspl jspl_w_n330_0(.douta(w_n330_0[0]),.doutb(w_n330_0[1]),.din(n330));
	jspl3 jspl3_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.doutc(w_n333_0[2]),.din(n333));
	jspl jspl_w_n335_0(.douta(w_n335_0[0]),.doutb(w_n335_0[1]),.din(n335));
	jspl jspl_w_n337_0(.douta(w_n337_0[0]),.doutb(w_n337_0[1]),.din(n337));
	jspl jspl_w_n338_0(.douta(w_n338_0[0]),.doutb(w_n338_0[1]),.din(n338));
	jspl jspl_w_n342_0(.douta(w_n342_0[0]),.doutb(w_n342_0[1]),.din(n342));
	jspl jspl_w_n343_0(.douta(w_n343_0[0]),.doutb(w_n343_0[1]),.din(n343));
	jspl jspl_w_n345_0(.douta(w_n345_0[0]),.doutb(w_n345_0[1]),.din(n345));
	jspl jspl_w_n349_0(.douta(w_n349_0[0]),.doutb(w_n349_0[1]),.din(n349));
	jspl3 jspl3_w_n352_0(.douta(w_n352_0[0]),.doutb(w_n352_0[1]),.doutc(w_n352_0[2]),.din(n352));
	jspl3 jspl3_w_n352_1(.douta(w_n352_1[0]),.doutb(w_n352_1[1]),.doutc(w_n352_1[2]),.din(w_n352_0[0]));
	jspl3 jspl3_w_n352_2(.douta(w_n352_2[0]),.doutb(w_n352_2[1]),.doutc(w_n352_2[2]),.din(w_n352_0[1]));
	jspl3 jspl3_w_n352_3(.douta(w_n352_3[0]),.doutb(w_n352_3[1]),.doutc(w_n352_3[2]),.din(w_n352_0[2]));
	jspl3 jspl3_w_n352_4(.douta(w_n352_4[0]),.doutb(w_n352_4[1]),.doutc(w_n352_4[2]),.din(w_n352_1[0]));
	jspl3 jspl3_w_n352_5(.douta(w_n352_5[0]),.doutb(w_n352_5[1]),.doutc(w_n352_5[2]),.din(w_n352_1[1]));
	jspl3 jspl3_w_n352_6(.douta(w_n352_6[0]),.doutb(w_n352_6[1]),.doutc(w_n352_6[2]),.din(w_n352_1[2]));
	jspl3 jspl3_w_n352_7(.douta(w_n352_7[0]),.doutb(w_n352_7[1]),.doutc(w_n352_7[2]),.din(w_n352_2[0]));
	jspl3 jspl3_w_n352_8(.douta(w_n352_8[0]),.doutb(w_n352_8[1]),.doutc(w_n352_8[2]),.din(w_n352_2[1]));
	jspl3 jspl3_w_n352_9(.douta(w_n352_9[0]),.doutb(w_n352_9[1]),.doutc(w_n352_9[2]),.din(w_n352_2[2]));
	jspl3 jspl3_w_n352_10(.douta(w_n352_10[0]),.doutb(w_n352_10[1]),.doutc(w_n352_10[2]),.din(w_n352_3[0]));
	jspl3 jspl3_w_n352_11(.douta(w_n352_11[0]),.doutb(w_n352_11[1]),.doutc(w_n352_11[2]),.din(w_n352_3[1]));
	jspl3 jspl3_w_n352_12(.douta(w_n352_12[0]),.doutb(w_n352_12[1]),.doutc(w_n352_12[2]),.din(w_n352_3[2]));
	jspl3 jspl3_w_n352_13(.douta(w_n352_13[0]),.doutb(w_n352_13[1]),.doutc(w_n352_13[2]),.din(w_n352_4[0]));
	jspl3 jspl3_w_n352_14(.douta(w_n352_14[0]),.doutb(w_n352_14[1]),.doutc(w_n352_14[2]),.din(w_n352_4[1]));
	jspl3 jspl3_w_n352_15(.douta(w_n352_15[0]),.doutb(w_n352_15[1]),.doutc(w_n352_15[2]),.din(w_n352_4[2]));
	jspl3 jspl3_w_n352_16(.douta(w_n352_16[0]),.doutb(w_n352_16[1]),.doutc(w_n352_16[2]),.din(w_n352_5[0]));
	jspl3 jspl3_w_n352_17(.douta(w_n352_17[0]),.doutb(w_n352_17[1]),.doutc(w_n352_17[2]),.din(w_n352_5[1]));
	jspl3 jspl3_w_n352_18(.douta(w_n352_18[0]),.doutb(w_n352_18[1]),.doutc(w_n352_18[2]),.din(w_n352_5[2]));
	jspl3 jspl3_w_n352_19(.douta(w_n352_19[0]),.doutb(w_n352_19[1]),.doutc(w_n352_19[2]),.din(w_n352_6[0]));
	jspl3 jspl3_w_n352_20(.douta(w_n352_20[0]),.doutb(w_n352_20[1]),.doutc(w_n352_20[2]),.din(w_n352_6[1]));
	jspl3 jspl3_w_n352_21(.douta(w_n352_21[0]),.doutb(w_n352_21[1]),.doutc(w_n352_21[2]),.din(w_n352_6[2]));
	jspl3 jspl3_w_n352_22(.douta(w_n352_22[0]),.doutb(w_n352_22[1]),.doutc(w_n352_22[2]),.din(w_n352_7[0]));
	jspl3 jspl3_w_n352_23(.douta(w_n352_23[0]),.doutb(w_n352_23[1]),.doutc(w_n352_23[2]),.din(w_n352_7[1]));
	jspl3 jspl3_w_n352_24(.douta(w_n352_24[0]),.doutb(w_n352_24[1]),.doutc(w_n352_24[2]),.din(w_n352_7[2]));
	jspl3 jspl3_w_n352_25(.douta(w_n352_25[0]),.doutb(w_n352_25[1]),.doutc(w_n352_25[2]),.din(w_n352_8[0]));
	jspl3 jspl3_w_n352_26(.douta(w_n352_26[0]),.doutb(w_n352_26[1]),.doutc(w_n352_26[2]),.din(w_n352_8[1]));
	jspl3 jspl3_w_n352_27(.douta(w_n352_27[0]),.doutb(w_n352_27[1]),.doutc(w_n352_27[2]),.din(w_n352_8[2]));
	jspl3 jspl3_w_n352_28(.douta(w_n352_28[0]),.doutb(w_n352_28[1]),.doutc(w_n352_28[2]),.din(w_n352_9[0]));
	jspl3 jspl3_w_n352_29(.douta(w_n352_29[0]),.doutb(w_n352_29[1]),.doutc(w_n352_29[2]),.din(w_n352_9[1]));
	jspl3 jspl3_w_n352_30(.douta(w_n352_30[0]),.doutb(w_n352_30[1]),.doutc(w_n352_30[2]),.din(w_n352_9[2]));
	jspl3 jspl3_w_n352_31(.douta(w_n352_31[0]),.doutb(w_n352_31[1]),.doutc(w_n352_31[2]),.din(w_n352_10[0]));
	jspl3 jspl3_w_n352_32(.douta(w_n352_32[0]),.doutb(w_n352_32[1]),.doutc(w_n352_32[2]),.din(w_n352_10[1]));
	jspl3 jspl3_w_n352_33(.douta(w_n352_33[0]),.doutb(w_n352_33[1]),.doutc(w_n352_33[2]),.din(w_n352_10[2]));
	jspl3 jspl3_w_n352_34(.douta(w_n352_34[0]),.doutb(w_n352_34[1]),.doutc(w_n352_34[2]),.din(w_n352_11[0]));
	jspl3 jspl3_w_n352_35(.douta(w_n352_35[0]),.doutb(w_n352_35[1]),.doutc(w_n352_35[2]),.din(w_n352_11[1]));
	jspl3 jspl3_w_n352_36(.douta(w_n352_36[0]),.doutb(w_n352_36[1]),.doutc(w_n352_36[2]),.din(w_n352_11[2]));
	jspl3 jspl3_w_n352_37(.douta(w_n352_37[0]),.doutb(w_n352_37[1]),.doutc(w_n352_37[2]),.din(w_n352_12[0]));
	jspl3 jspl3_w_n352_38(.douta(w_n352_38[0]),.doutb(w_n352_38[1]),.doutc(w_n352_38[2]),.din(w_n352_12[1]));
	jspl3 jspl3_w_n352_39(.douta(w_n352_39[0]),.doutb(w_n352_39[1]),.doutc(w_n352_39[2]),.din(w_n352_12[2]));
	jspl3 jspl3_w_n352_40(.douta(w_n352_40[0]),.doutb(w_n352_40[1]),.doutc(w_n352_40[2]),.din(w_n352_13[0]));
	jspl3 jspl3_w_n352_41(.douta(w_n352_41[0]),.doutb(w_n352_41[1]),.doutc(w_n352_41[2]),.din(w_n352_13[1]));
	jspl3 jspl3_w_n352_42(.douta(w_n352_42[0]),.doutb(w_n352_42[1]),.doutc(w_n352_42[2]),.din(w_n352_13[2]));
	jspl3 jspl3_w_n352_43(.douta(w_n352_43[0]),.doutb(w_n352_43[1]),.doutc(w_n352_43[2]),.din(w_n352_14[0]));
	jspl3 jspl3_w_n352_44(.douta(w_n352_44[0]),.doutb(w_n352_44[1]),.doutc(w_n352_44[2]),.din(w_n352_14[1]));
	jspl3 jspl3_w_n352_45(.douta(w_n352_45[0]),.doutb(w_n352_45[1]),.doutc(w_n352_45[2]),.din(w_n352_14[2]));
	jspl3 jspl3_w_n352_46(.douta(w_n352_46[0]),.doutb(w_n352_46[1]),.doutc(w_n352_46[2]),.din(w_n352_15[0]));
	jspl3 jspl3_w_n352_47(.douta(w_n352_47[0]),.doutb(w_n352_47[1]),.doutc(w_n352_47[2]),.din(w_n352_15[1]));
	jspl3 jspl3_w_n352_48(.douta(w_n352_48[0]),.doutb(w_n352_48[1]),.doutc(w_n352_48[2]),.din(w_n352_15[2]));
	jspl3 jspl3_w_n352_49(.douta(w_n352_49[0]),.doutb(w_n352_49[1]),.doutc(w_n352_49[2]),.din(w_n352_16[0]));
	jspl3 jspl3_w_n352_50(.douta(w_n352_50[0]),.doutb(w_n352_50[1]),.doutc(w_n352_50[2]),.din(w_n352_16[1]));
	jspl3 jspl3_w_n352_51(.douta(w_n352_51[0]),.doutb(w_n352_51[1]),.doutc(w_n352_51[2]),.din(w_n352_16[2]));
	jspl3 jspl3_w_n352_52(.douta(w_n352_52[0]),.doutb(w_n352_52[1]),.doutc(w_n352_52[2]),.din(w_n352_17[0]));
	jspl3 jspl3_w_n352_53(.douta(w_n352_53[0]),.doutb(w_n352_53[1]),.doutc(w_n352_53[2]),.din(w_n352_17[1]));
	jspl3 jspl3_w_n352_54(.douta(w_n352_54[0]),.doutb(w_n352_54[1]),.doutc(w_n352_54[2]),.din(w_n352_17[2]));
	jspl3 jspl3_w_n352_55(.douta(w_n352_55[0]),.doutb(w_n352_55[1]),.doutc(w_n352_55[2]),.din(w_n352_18[0]));
	jspl3 jspl3_w_n352_56(.douta(w_n352_56[0]),.doutb(w_n352_56[1]),.doutc(w_n352_56[2]),.din(w_n352_18[1]));
	jspl3 jspl3_w_n352_57(.douta(w_n352_57[0]),.doutb(w_n352_57[1]),.doutc(w_n352_57[2]),.din(w_n352_18[2]));
	jspl3 jspl3_w_n352_58(.douta(w_n352_58[0]),.doutb(w_n352_58[1]),.doutc(w_n352_58[2]),.din(w_n352_19[0]));
	jspl3 jspl3_w_n352_59(.douta(w_n352_59[0]),.doutb(w_n352_59[1]),.doutc(w_n352_59[2]),.din(w_n352_19[1]));
	jspl3 jspl3_w_n352_60(.douta(w_n352_60[0]),.doutb(w_n352_60[1]),.doutc(w_n352_60[2]),.din(w_n352_19[2]));
	jspl3 jspl3_w_n352_61(.douta(w_n352_61[0]),.doutb(w_n352_61[1]),.doutc(w_n352_61[2]),.din(w_n352_20[0]));
	jspl3 jspl3_w_n352_62(.douta(w_n352_62[0]),.doutb(w_n352_62[1]),.doutc(w_n352_62[2]),.din(w_n352_20[1]));
	jspl3 jspl3_w_n352_63(.douta(w_n352_63[0]),.doutb(w_n352_63[1]),.doutc(w_n352_63[2]),.din(w_n352_20[2]));
	jspl3 jspl3_w_n352_64(.douta(w_n352_64[0]),.doutb(w_n352_64[1]),.doutc(w_n352_64[2]),.din(w_n352_21[0]));
	jspl3 jspl3_w_n352_65(.douta(w_n352_65[0]),.doutb(w_n352_65[1]),.doutc(w_n352_65[2]),.din(w_n352_21[1]));
	jspl3 jspl3_w_n352_66(.douta(w_n352_66[0]),.doutb(w_n352_66[1]),.doutc(w_n352_66[2]),.din(w_n352_21[2]));
	jspl3 jspl3_w_n352_67(.douta(w_n352_67[0]),.doutb(w_n352_67[1]),.doutc(w_n352_67[2]),.din(w_n352_22[0]));
	jspl3 jspl3_w_n352_68(.douta(w_n352_68[0]),.doutb(w_n352_68[1]),.doutc(w_n352_68[2]),.din(w_n352_22[1]));
	jspl3 jspl3_w_n352_69(.douta(w_n352_69[0]),.doutb(w_n352_69[1]),.doutc(w_n352_69[2]),.din(w_n352_22[2]));
	jspl3 jspl3_w_n352_70(.douta(w_n352_70[0]),.doutb(w_n352_70[1]),.doutc(w_n352_70[2]),.din(w_n352_23[0]));
	jspl3 jspl3_w_n352_71(.douta(w_n352_71[0]),.doutb(w_n352_71[1]),.doutc(w_n352_71[2]),.din(w_n352_23[1]));
	jspl3 jspl3_w_n352_72(.douta(w_n352_72[0]),.doutb(w_n352_72[1]),.doutc(w_n352_72[2]),.din(w_n352_23[2]));
	jspl3 jspl3_w_n352_73(.douta(w_n352_73[0]),.doutb(w_n352_73[1]),.doutc(w_n352_73[2]),.din(w_n352_24[0]));
	jspl jspl_w_n352_74(.douta(w_n352_74[0]),.doutb(w_n352_74[1]),.din(w_n352_24[1]));
	jspl3 jspl3_w_n354_0(.douta(w_n354_0[0]),.doutb(w_n354_0[1]),.doutc(w_n354_0[2]),.din(n354));
	jspl3 jspl3_w_n354_1(.douta(w_n354_1[0]),.doutb(w_n354_1[1]),.doutc(w_n354_1[2]),.din(w_n354_0[0]));
	jspl jspl_w_n355_0(.douta(w_n355_0[0]),.doutb(w_n355_0[1]),.din(n355));
	jspl3 jspl3_w_n356_0(.douta(w_n356_0[0]),.doutb(w_n356_0[1]),.doutc(w_n356_0[2]),.din(n356));
	jspl jspl_w_n357_0(.douta(w_n357_0[0]),.doutb(w_n357_0[1]),.din(n357));
	jspl3 jspl3_w_n359_0(.douta(w_n359_0[0]),.doutb(w_n359_0[1]),.doutc(w_n359_0[2]),.din(n359));
	jspl jspl_w_n360_0(.douta(w_n360_0[0]),.doutb(w_n360_0[1]),.din(n360));
	jspl3 jspl3_w_n367_0(.douta(w_n367_0[0]),.doutb(w_n367_0[1]),.doutc(w_n367_0[2]),.din(n367));
	jspl jspl_w_n368_0(.douta(w_n368_0[0]),.doutb(w_n368_0[1]),.din(n368));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(n371));
	jspl3 jspl3_w_n373_0(.douta(w_n373_0[0]),.doutb(w_n373_0[1]),.doutc(w_n373_0[2]),.din(n373));
	jspl3 jspl3_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.doutc(w_n375_0[2]),.din(n375));
	jspl jspl_w_n376_0(.douta(w_n376_0[0]),.doutb(w_n376_0[1]),.din(n376));
	jspl3 jspl3_w_n380_0(.douta(w_n380_0[0]),.doutb(w_n380_0[1]),.doutc(w_n380_0[2]),.din(n380));
	jspl3 jspl3_w_n383_0(.douta(w_n383_0[0]),.doutb(w_n383_0[1]),.doutc(w_n383_0[2]),.din(n383));
	jspl3 jspl3_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.doutc(w_n386_0[2]),.din(n386));
	jspl jspl_w_n386_1(.douta(w_n386_1[0]),.doutb(w_n386_1[1]),.din(w_n386_0[0]));
	jspl3 jspl3_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.doutc(w_n387_0[2]),.din(n387));
	jspl jspl_w_n388_0(.douta(w_n388_0[0]),.doutb(w_n388_0[1]),.din(n388));
	jspl jspl_w_n389_0(.douta(w_n389_0[0]),.doutb(w_n389_0[1]),.din(n389));
	jspl jspl_w_n390_0(.douta(w_n390_0[0]),.doutb(w_n390_0[1]),.din(n390));
	jspl jspl_w_n393_0(.douta(w_n393_0[0]),.doutb(w_n393_0[1]),.din(n393));
	jspl jspl_w_n395_0(.douta(w_n395_0[0]),.doutb(w_n395_0[1]),.din(n395));
	jspl jspl_w_n407_0(.douta(w_n407_0[0]),.doutb(w_n407_0[1]),.din(n407));
	jspl jspl_w_n418_0(.douta(w_n418_0[0]),.doutb(w_n418_0[1]),.din(n418));
	jspl jspl_w_n419_0(.douta(w_n419_0[0]),.doutb(w_n419_0[1]),.din(n419));
	jspl3 jspl3_w_n422_0(.douta(w_n422_0[0]),.doutb(w_n422_0[1]),.doutc(w_n422_0[2]),.din(n422));
	jspl jspl_w_n423_0(.douta(w_n423_0[0]),.doutb(w_n423_0[1]),.din(n423));
	jspl3 jspl3_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.doutc(w_n425_0[2]),.din(n425));
	jspl jspl_w_n425_1(.douta(w_n425_1[0]),.doutb(w_n425_1[1]),.din(w_n425_0[0]));
	jspl jspl_w_n426_0(.douta(w_n426_0[0]),.doutb(w_n426_0[1]),.din(n426));
	jspl3 jspl3_w_n427_0(.douta(w_n427_0[0]),.doutb(w_n427_0[1]),.doutc(w_n427_0[2]),.din(n427));
	jspl jspl_w_n428_0(.douta(w_n428_0[0]),.doutb(w_n428_0[1]),.din(n428));
	jspl3 jspl3_w_n429_0(.douta(w_n429_0[0]),.doutb(w_n429_0[1]),.doutc(w_n429_0[2]),.din(n429));
	jspl jspl_w_n430_0(.douta(w_n430_0[0]),.doutb(w_n430_0[1]),.din(n430));
	jspl jspl_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.din(n435));
	jspl jspl_w_n440_0(.douta(w_n440_0[0]),.doutb(w_n440_0[1]),.din(n440));
	jspl jspl_w_n441_0(.douta(w_n441_0[0]),.doutb(w_n441_0[1]),.din(n441));
	jspl3 jspl3_w_n443_0(.douta(w_n443_0[0]),.doutb(w_n443_0[1]),.doutc(w_n443_0[2]),.din(n443));
	jspl3 jspl3_w_n443_1(.douta(w_n443_1[0]),.doutb(w_n443_1[1]),.doutc(w_n443_1[2]),.din(w_n443_0[0]));
	jspl3 jspl3_w_n443_2(.douta(w_n443_2[0]),.doutb(w_n443_2[1]),.doutc(w_n443_2[2]),.din(w_n443_0[1]));
	jspl3 jspl3_w_n443_3(.douta(w_n443_3[0]),.doutb(w_n443_3[1]),.doutc(w_n443_3[2]),.din(w_n443_0[2]));
	jspl3 jspl3_w_n443_4(.douta(w_n443_4[0]),.doutb(w_n443_4[1]),.doutc(w_n443_4[2]),.din(w_n443_1[0]));
	jspl3 jspl3_w_n443_5(.douta(w_n443_5[0]),.doutb(w_n443_5[1]),.doutc(w_n443_5[2]),.din(w_n443_1[1]));
	jspl3 jspl3_w_n443_6(.douta(w_n443_6[0]),.doutb(w_n443_6[1]),.doutc(w_n443_6[2]),.din(w_n443_1[2]));
	jspl3 jspl3_w_n443_7(.douta(w_n443_7[0]),.doutb(w_n443_7[1]),.doutc(w_n443_7[2]),.din(w_n443_2[0]));
	jspl3 jspl3_w_n443_8(.douta(w_n443_8[0]),.doutb(w_n443_8[1]),.doutc(w_n443_8[2]),.din(w_n443_2[1]));
	jspl3 jspl3_w_n443_9(.douta(w_n443_9[0]),.doutb(w_n443_9[1]),.doutc(w_n443_9[2]),.din(w_n443_2[2]));
	jspl3 jspl3_w_n443_10(.douta(w_n443_10[0]),.doutb(w_n443_10[1]),.doutc(w_n443_10[2]),.din(w_n443_3[0]));
	jspl3 jspl3_w_n443_11(.douta(w_n443_11[0]),.doutb(w_n443_11[1]),.doutc(w_n443_11[2]),.din(w_n443_3[1]));
	jspl3 jspl3_w_n443_12(.douta(w_n443_12[0]),.doutb(w_n443_12[1]),.doutc(w_n443_12[2]),.din(w_n443_3[2]));
	jspl3 jspl3_w_n443_13(.douta(w_n443_13[0]),.doutb(w_n443_13[1]),.doutc(w_n443_13[2]),.din(w_n443_4[0]));
	jspl3 jspl3_w_n443_14(.douta(w_n443_14[0]),.doutb(w_n443_14[1]),.doutc(w_n443_14[2]),.din(w_n443_4[1]));
	jspl3 jspl3_w_n443_15(.douta(w_n443_15[0]),.doutb(w_n443_15[1]),.doutc(w_n443_15[2]),.din(w_n443_4[2]));
	jspl3 jspl3_w_n443_16(.douta(w_n443_16[0]),.doutb(w_n443_16[1]),.doutc(w_n443_16[2]),.din(w_n443_5[0]));
	jspl3 jspl3_w_n443_17(.douta(w_n443_17[0]),.doutb(w_n443_17[1]),.doutc(w_n443_17[2]),.din(w_n443_5[1]));
	jspl3 jspl3_w_n443_18(.douta(w_n443_18[0]),.doutb(w_n443_18[1]),.doutc(w_n443_18[2]),.din(w_n443_5[2]));
	jspl3 jspl3_w_n443_19(.douta(w_n443_19[0]),.doutb(w_n443_19[1]),.doutc(w_n443_19[2]),.din(w_n443_6[0]));
	jspl3 jspl3_w_n443_20(.douta(w_n443_20[0]),.doutb(w_n443_20[1]),.doutc(w_n443_20[2]),.din(w_n443_6[1]));
	jspl3 jspl3_w_n443_21(.douta(w_n443_21[0]),.doutb(w_n443_21[1]),.doutc(w_n443_21[2]),.din(w_n443_6[2]));
	jspl3 jspl3_w_n443_22(.douta(w_n443_22[0]),.doutb(w_n443_22[1]),.doutc(w_n443_22[2]),.din(w_n443_7[0]));
	jspl3 jspl3_w_n443_23(.douta(w_n443_23[0]),.doutb(w_n443_23[1]),.doutc(w_n443_23[2]),.din(w_n443_7[1]));
	jspl3 jspl3_w_n443_24(.douta(w_n443_24[0]),.doutb(w_n443_24[1]),.doutc(w_n443_24[2]),.din(w_n443_7[2]));
	jspl3 jspl3_w_n443_25(.douta(w_n443_25[0]),.doutb(w_n443_25[1]),.doutc(w_n443_25[2]),.din(w_n443_8[0]));
	jspl3 jspl3_w_n443_26(.douta(w_n443_26[0]),.doutb(w_n443_26[1]),.doutc(w_n443_26[2]),.din(w_n443_8[1]));
	jspl3 jspl3_w_n443_27(.douta(w_n443_27[0]),.doutb(w_n443_27[1]),.doutc(w_n443_27[2]),.din(w_n443_8[2]));
	jspl3 jspl3_w_n443_28(.douta(w_n443_28[0]),.doutb(w_n443_28[1]),.doutc(w_n443_28[2]),.din(w_n443_9[0]));
	jspl3 jspl3_w_n443_29(.douta(w_n443_29[0]),.doutb(w_n443_29[1]),.doutc(w_n443_29[2]),.din(w_n443_9[1]));
	jspl3 jspl3_w_n443_30(.douta(w_n443_30[0]),.doutb(w_n443_30[1]),.doutc(w_n443_30[2]),.din(w_n443_9[2]));
	jspl3 jspl3_w_n443_31(.douta(w_n443_31[0]),.doutb(w_n443_31[1]),.doutc(w_n443_31[2]),.din(w_n443_10[0]));
	jspl3 jspl3_w_n443_32(.douta(w_n443_32[0]),.doutb(w_n443_32[1]),.doutc(w_n443_32[2]),.din(w_n443_10[1]));
	jspl3 jspl3_w_n443_33(.douta(w_n443_33[0]),.doutb(w_n443_33[1]),.doutc(w_n443_33[2]),.din(w_n443_10[2]));
	jspl3 jspl3_w_n443_34(.douta(w_n443_34[0]),.doutb(w_n443_34[1]),.doutc(w_n443_34[2]),.din(w_n443_11[0]));
	jspl3 jspl3_w_n443_35(.douta(w_n443_35[0]),.doutb(w_n443_35[1]),.doutc(w_n443_35[2]),.din(w_n443_11[1]));
	jspl3 jspl3_w_n443_36(.douta(w_n443_36[0]),.doutb(w_n443_36[1]),.doutc(w_n443_36[2]),.din(w_n443_11[2]));
	jspl3 jspl3_w_n443_37(.douta(w_n443_37[0]),.doutb(w_n443_37[1]),.doutc(w_n443_37[2]),.din(w_n443_12[0]));
	jspl3 jspl3_w_n443_38(.douta(w_n443_38[0]),.doutb(w_n443_38[1]),.doutc(w_n443_38[2]),.din(w_n443_12[1]));
	jspl3 jspl3_w_n443_39(.douta(w_n443_39[0]),.doutb(w_n443_39[1]),.doutc(w_n443_39[2]),.din(w_n443_12[2]));
	jspl3 jspl3_w_n443_40(.douta(w_n443_40[0]),.doutb(w_n443_40[1]),.doutc(w_n443_40[2]),.din(w_n443_13[0]));
	jspl3 jspl3_w_n443_41(.douta(w_n443_41[0]),.doutb(w_n443_41[1]),.doutc(w_n443_41[2]),.din(w_n443_13[1]));
	jspl3 jspl3_w_n443_42(.douta(w_n443_42[0]),.doutb(w_n443_42[1]),.doutc(w_n443_42[2]),.din(w_n443_13[2]));
	jspl3 jspl3_w_n443_43(.douta(w_n443_43[0]),.doutb(w_n443_43[1]),.doutc(w_n443_43[2]),.din(w_n443_14[0]));
	jspl3 jspl3_w_n443_44(.douta(w_n443_44[0]),.doutb(w_n443_44[1]),.doutc(w_n443_44[2]),.din(w_n443_14[1]));
	jspl3 jspl3_w_n443_45(.douta(w_n443_45[0]),.doutb(w_n443_45[1]),.doutc(w_n443_45[2]),.din(w_n443_14[2]));
	jspl3 jspl3_w_n443_46(.douta(w_n443_46[0]),.doutb(w_n443_46[1]),.doutc(w_n443_46[2]),.din(w_n443_15[0]));
	jspl3 jspl3_w_n443_47(.douta(w_n443_47[0]),.doutb(w_n443_47[1]),.doutc(w_n443_47[2]),.din(w_n443_15[1]));
	jspl3 jspl3_w_n443_48(.douta(w_n443_48[0]),.doutb(w_n443_48[1]),.doutc(w_n443_48[2]),.din(w_n443_15[2]));
	jspl3 jspl3_w_n443_49(.douta(w_n443_49[0]),.doutb(w_n443_49[1]),.doutc(w_n443_49[2]),.din(w_n443_16[0]));
	jspl3 jspl3_w_n443_50(.douta(w_n443_50[0]),.doutb(w_n443_50[1]),.doutc(w_n443_50[2]),.din(w_n443_16[1]));
	jspl3 jspl3_w_n443_51(.douta(w_n443_51[0]),.doutb(w_n443_51[1]),.doutc(w_n443_51[2]),.din(w_n443_16[2]));
	jspl3 jspl3_w_n443_52(.douta(w_n443_52[0]),.doutb(w_n443_52[1]),.doutc(w_n443_52[2]),.din(w_n443_17[0]));
	jspl3 jspl3_w_n443_53(.douta(w_n443_53[0]),.doutb(w_n443_53[1]),.doutc(w_n443_53[2]),.din(w_n443_17[1]));
	jspl3 jspl3_w_n443_54(.douta(w_n443_54[0]),.doutb(w_n443_54[1]),.doutc(w_n443_54[2]),.din(w_n443_17[2]));
	jspl3 jspl3_w_n443_55(.douta(w_n443_55[0]),.doutb(w_n443_55[1]),.doutc(w_n443_55[2]),.din(w_n443_18[0]));
	jspl3 jspl3_w_n443_56(.douta(w_n443_56[0]),.doutb(w_n443_56[1]),.doutc(w_n443_56[2]),.din(w_n443_18[1]));
	jspl3 jspl3_w_n443_57(.douta(w_n443_57[0]),.doutb(w_n443_57[1]),.doutc(w_n443_57[2]),.din(w_n443_18[2]));
	jspl3 jspl3_w_n443_58(.douta(w_n443_58[0]),.doutb(w_n443_58[1]),.doutc(w_n443_58[2]),.din(w_n443_19[0]));
	jspl3 jspl3_w_n443_59(.douta(w_n443_59[0]),.doutb(w_n443_59[1]),.doutc(w_n443_59[2]),.din(w_n443_19[1]));
	jspl3 jspl3_w_n443_60(.douta(w_n443_60[0]),.doutb(w_n443_60[1]),.doutc(w_n443_60[2]),.din(w_n443_19[2]));
	jspl3 jspl3_w_n443_61(.douta(w_n443_61[0]),.doutb(w_n443_61[1]),.doutc(w_n443_61[2]),.din(w_n443_20[0]));
	jspl3 jspl3_w_n443_62(.douta(w_n443_62[0]),.doutb(w_n443_62[1]),.doutc(w_n443_62[2]),.din(w_n443_20[1]));
	jspl3 jspl3_w_n443_63(.douta(w_n443_63[0]),.doutb(w_n443_63[1]),.doutc(w_n443_63[2]),.din(w_n443_20[2]));
	jspl3 jspl3_w_n443_64(.douta(w_n443_64[0]),.doutb(w_n443_64[1]),.doutc(w_n443_64[2]),.din(w_n443_21[0]));
	jspl3 jspl3_w_n443_65(.douta(w_n443_65[0]),.doutb(w_n443_65[1]),.doutc(w_n443_65[2]),.din(w_n443_21[1]));
	jspl3 jspl3_w_n443_66(.douta(w_n443_66[0]),.doutb(w_n443_66[1]),.doutc(w_n443_66[2]),.din(w_n443_21[2]));
	jspl3 jspl3_w_n443_67(.douta(w_n443_67[0]),.doutb(w_n443_67[1]),.doutc(w_n443_67[2]),.din(w_n443_22[0]));
	jspl3 jspl3_w_n443_68(.douta(w_n443_68[0]),.doutb(w_n443_68[1]),.doutc(w_n443_68[2]),.din(w_n443_22[1]));
	jspl3 jspl3_w_n443_69(.douta(w_n443_69[0]),.doutb(w_n443_69[1]),.doutc(w_n443_69[2]),.din(w_n443_22[2]));
	jspl3 jspl3_w_n443_70(.douta(w_n443_70[0]),.doutb(w_n443_70[1]),.doutc(w_n443_70[2]),.din(w_n443_23[0]));
	jspl3 jspl3_w_n443_71(.douta(w_n443_71[0]),.doutb(w_n443_71[1]),.doutc(w_n443_71[2]),.din(w_n443_23[1]));
	jspl3 jspl3_w_n443_72(.douta(w_n443_72[0]),.doutb(w_n443_72[1]),.doutc(w_n443_72[2]),.din(w_n443_23[2]));
	jspl jspl_w_n443_73(.douta(w_n443_73[0]),.doutb(w_n443_73[1]),.din(w_n443_24[0]));
	jspl3 jspl3_w_n447_0(.douta(w_n447_0[0]),.doutb(w_n447_0[1]),.doutc(w_n447_0[2]),.din(n447));
	jspl jspl_w_n448_0(.douta(w_n448_0[0]),.doutb(w_n448_0[1]),.din(n448));
	jspl jspl_w_n450_0(.douta(w_n450_0[0]),.doutb(w_n450_0[1]),.din(n450));
	jspl jspl_w_n452_0(.douta(w_n452_0[0]),.doutb(w_n452_0[1]),.din(n452));
	jspl jspl_w_n453_0(.douta(w_n453_0[0]),.doutb(w_n453_0[1]),.din(n453));
	jspl3 jspl3_w_n455_0(.douta(w_n455_0[0]),.doutb(w_n455_0[1]),.doutc(w_n455_0[2]),.din(n455));
	jspl jspl_w_n456_0(.douta(w_n456_0[0]),.doutb(w_n456_0[1]),.din(n456));
	jspl jspl_w_n460_0(.douta(w_n460_0[0]),.doutb(w_n460_0[1]),.din(n460));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_n462_0[1]),.doutc(w_n462_0[2]),.din(n462));
	jspl jspl_w_n463_0(.douta(w_n463_0[0]),.doutb(w_n463_0[1]),.din(n463));
	jspl jspl_w_n474_0(.douta(w_n474_0[0]),.doutb(w_n474_0[1]),.din(n474));
	jspl jspl_w_n481_0(.douta(w_n481_0[0]),.doutb(w_n481_0[1]),.din(n481));
	jspl3 jspl3_w_n487_0(.douta(w_n487_0[0]),.doutb(w_n487_0[1]),.doutc(w_n487_0[2]),.din(n487));
	jspl jspl_w_n489_0(.douta(w_n489_0[0]),.doutb(w_n489_0[1]),.din(n489));
	jspl jspl_w_n490_0(.douta(w_n490_0[0]),.doutb(w_n490_0[1]),.din(n490));
	jspl jspl_w_n493_0(.douta(w_n493_0[0]),.doutb(w_n493_0[1]),.din(n493));
	jspl jspl_w_n499_0(.douta(w_n499_0[0]),.doutb(w_n499_0[1]),.din(n499));
	jspl3 jspl3_w_n500_0(.douta(w_n500_0[0]),.doutb(w_n500_0[1]),.doutc(w_n500_0[2]),.din(n500));
	jspl jspl_w_n504_0(.douta(w_n504_0[0]),.doutb(w_n504_0[1]),.din(n504));
	jspl jspl_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.din(n507));
	jspl jspl_w_n511_0(.douta(w_n511_0[0]),.doutb(w_n511_0[1]),.din(n511));
	jspl3 jspl3_w_n515_0(.douta(w_n515_0[0]),.doutb(w_n515_0[1]),.doutc(w_n515_0[2]),.din(n515));
	jspl3 jspl3_w_n515_1(.douta(w_n515_1[0]),.doutb(w_n515_1[1]),.doutc(w_n515_1[2]),.din(w_n515_0[0]));
	jspl3 jspl3_w_n515_2(.douta(w_n515_2[0]),.doutb(w_n515_2[1]),.doutc(w_n515_2[2]),.din(w_n515_0[1]));
	jspl3 jspl3_w_n515_3(.douta(w_n515_3[0]),.doutb(w_n515_3[1]),.doutc(w_n515_3[2]),.din(w_n515_0[2]));
	jspl3 jspl3_w_n515_4(.douta(w_n515_4[0]),.doutb(w_n515_4[1]),.doutc(w_n515_4[2]),.din(w_n515_1[0]));
	jspl3 jspl3_w_n515_5(.douta(w_n515_5[0]),.doutb(w_n515_5[1]),.doutc(w_n515_5[2]),.din(w_n515_1[1]));
	jspl3 jspl3_w_n515_6(.douta(w_n515_6[0]),.doutb(w_n515_6[1]),.doutc(w_n515_6[2]),.din(w_n515_1[2]));
	jspl3 jspl3_w_n515_7(.douta(w_n515_7[0]),.doutb(w_n515_7[1]),.doutc(w_n515_7[2]),.din(w_n515_2[0]));
	jspl3 jspl3_w_n515_8(.douta(w_n515_8[0]),.doutb(w_n515_8[1]),.doutc(w_n515_8[2]),.din(w_n515_2[1]));
	jspl3 jspl3_w_n515_9(.douta(w_n515_9[0]),.doutb(w_n515_9[1]),.doutc(w_n515_9[2]),.din(w_n515_2[2]));
	jspl3 jspl3_w_n515_10(.douta(w_n515_10[0]),.doutb(w_n515_10[1]),.doutc(w_n515_10[2]),.din(w_n515_3[0]));
	jspl3 jspl3_w_n515_11(.douta(w_n515_11[0]),.doutb(w_n515_11[1]),.doutc(w_n515_11[2]),.din(w_n515_3[1]));
	jspl3 jspl3_w_n515_12(.douta(w_n515_12[0]),.doutb(w_n515_12[1]),.doutc(w_n515_12[2]),.din(w_n515_3[2]));
	jspl3 jspl3_w_n515_13(.douta(w_n515_13[0]),.doutb(w_n515_13[1]),.doutc(w_n515_13[2]),.din(w_n515_4[0]));
	jspl3 jspl3_w_n515_14(.douta(w_n515_14[0]),.doutb(w_n515_14[1]),.doutc(w_n515_14[2]),.din(w_n515_4[1]));
	jspl3 jspl3_w_n515_15(.douta(w_n515_15[0]),.doutb(w_n515_15[1]),.doutc(w_n515_15[2]),.din(w_n515_4[2]));
	jspl3 jspl3_w_n515_16(.douta(w_n515_16[0]),.doutb(w_n515_16[1]),.doutc(w_n515_16[2]),.din(w_n515_5[0]));
	jspl3 jspl3_w_n515_17(.douta(w_n515_17[0]),.doutb(w_n515_17[1]),.doutc(w_n515_17[2]),.din(w_n515_5[1]));
	jspl3 jspl3_w_n515_18(.douta(w_n515_18[0]),.doutb(w_n515_18[1]),.doutc(w_n515_18[2]),.din(w_n515_5[2]));
	jspl3 jspl3_w_n515_19(.douta(w_n515_19[0]),.doutb(w_n515_19[1]),.doutc(w_n515_19[2]),.din(w_n515_6[0]));
	jspl3 jspl3_w_n515_20(.douta(w_n515_20[0]),.doutb(w_n515_20[1]),.doutc(w_n515_20[2]),.din(w_n515_6[1]));
	jspl3 jspl3_w_n515_21(.douta(w_n515_21[0]),.doutb(w_n515_21[1]),.doutc(w_n515_21[2]),.din(w_n515_6[2]));
	jspl3 jspl3_w_n515_22(.douta(w_n515_22[0]),.doutb(w_n515_22[1]),.doutc(w_n515_22[2]),.din(w_n515_7[0]));
	jspl3 jspl3_w_n515_23(.douta(w_n515_23[0]),.doutb(w_n515_23[1]),.doutc(w_n515_23[2]),.din(w_n515_7[1]));
	jspl3 jspl3_w_n515_24(.douta(w_n515_24[0]),.doutb(w_n515_24[1]),.doutc(w_n515_24[2]),.din(w_n515_7[2]));
	jspl3 jspl3_w_n515_25(.douta(w_n515_25[0]),.doutb(w_n515_25[1]),.doutc(w_n515_25[2]),.din(w_n515_8[0]));
	jspl3 jspl3_w_n515_26(.douta(w_n515_26[0]),.doutb(w_n515_26[1]),.doutc(w_n515_26[2]),.din(w_n515_8[1]));
	jspl3 jspl3_w_n515_27(.douta(w_n515_27[0]),.doutb(w_n515_27[1]),.doutc(w_n515_27[2]),.din(w_n515_8[2]));
	jspl3 jspl3_w_n515_28(.douta(w_n515_28[0]),.doutb(w_n515_28[1]),.doutc(w_n515_28[2]),.din(w_n515_9[0]));
	jspl3 jspl3_w_n515_29(.douta(w_n515_29[0]),.doutb(w_n515_29[1]),.doutc(w_n515_29[2]),.din(w_n515_9[1]));
	jspl3 jspl3_w_n515_30(.douta(w_n515_30[0]),.doutb(w_n515_30[1]),.doutc(w_n515_30[2]),.din(w_n515_9[2]));
	jspl3 jspl3_w_n515_31(.douta(w_n515_31[0]),.doutb(w_n515_31[1]),.doutc(w_n515_31[2]),.din(w_n515_10[0]));
	jspl3 jspl3_w_n515_32(.douta(w_n515_32[0]),.doutb(w_n515_32[1]),.doutc(w_n515_32[2]),.din(w_n515_10[1]));
	jspl3 jspl3_w_n515_33(.douta(w_n515_33[0]),.doutb(w_n515_33[1]),.doutc(w_n515_33[2]),.din(w_n515_10[2]));
	jspl3 jspl3_w_n515_34(.douta(w_n515_34[0]),.doutb(w_n515_34[1]),.doutc(w_n515_34[2]),.din(w_n515_11[0]));
	jspl3 jspl3_w_n515_35(.douta(w_n515_35[0]),.doutb(w_n515_35[1]),.doutc(w_n515_35[2]),.din(w_n515_11[1]));
	jspl3 jspl3_w_n515_36(.douta(w_n515_36[0]),.doutb(w_n515_36[1]),.doutc(w_n515_36[2]),.din(w_n515_11[2]));
	jspl3 jspl3_w_n515_37(.douta(w_n515_37[0]),.doutb(w_n515_37[1]),.doutc(w_n515_37[2]),.din(w_n515_12[0]));
	jspl3 jspl3_w_n515_38(.douta(w_n515_38[0]),.doutb(w_n515_38[1]),.doutc(w_n515_38[2]),.din(w_n515_12[1]));
	jspl3 jspl3_w_n515_39(.douta(w_n515_39[0]),.doutb(w_n515_39[1]),.doutc(w_n515_39[2]),.din(w_n515_12[2]));
	jspl3 jspl3_w_n515_40(.douta(w_n515_40[0]),.doutb(w_n515_40[1]),.doutc(w_n515_40[2]),.din(w_n515_13[0]));
	jspl3 jspl3_w_n515_41(.douta(w_n515_41[0]),.doutb(w_n515_41[1]),.doutc(w_n515_41[2]),.din(w_n515_13[1]));
	jspl3 jspl3_w_n515_42(.douta(w_n515_42[0]),.doutb(w_n515_42[1]),.doutc(w_n515_42[2]),.din(w_n515_13[2]));
	jspl3 jspl3_w_n515_43(.douta(w_n515_43[0]),.doutb(w_n515_43[1]),.doutc(w_n515_43[2]),.din(w_n515_14[0]));
	jspl3 jspl3_w_n515_44(.douta(w_n515_44[0]),.doutb(w_n515_44[1]),.doutc(w_n515_44[2]),.din(w_n515_14[1]));
	jspl3 jspl3_w_n515_45(.douta(w_n515_45[0]),.doutb(w_n515_45[1]),.doutc(w_n515_45[2]),.din(w_n515_14[2]));
	jspl3 jspl3_w_n515_46(.douta(w_n515_46[0]),.doutb(w_n515_46[1]),.doutc(w_n515_46[2]),.din(w_n515_15[0]));
	jspl3 jspl3_w_n515_47(.douta(w_n515_47[0]),.doutb(w_n515_47[1]),.doutc(w_n515_47[2]),.din(w_n515_15[1]));
	jspl3 jspl3_w_n515_48(.douta(w_n515_48[0]),.doutb(w_n515_48[1]),.doutc(w_n515_48[2]),.din(w_n515_15[2]));
	jspl3 jspl3_w_n515_49(.douta(w_n515_49[0]),.doutb(w_n515_49[1]),.doutc(w_n515_49[2]),.din(w_n515_16[0]));
	jspl3 jspl3_w_n515_50(.douta(w_n515_50[0]),.doutb(w_n515_50[1]),.doutc(w_n515_50[2]),.din(w_n515_16[1]));
	jspl3 jspl3_w_n515_51(.douta(w_n515_51[0]),.doutb(w_n515_51[1]),.doutc(w_n515_51[2]),.din(w_n515_16[2]));
	jspl3 jspl3_w_n515_52(.douta(w_n515_52[0]),.doutb(w_n515_52[1]),.doutc(w_n515_52[2]),.din(w_n515_17[0]));
	jspl3 jspl3_w_n515_53(.douta(w_n515_53[0]),.doutb(w_n515_53[1]),.doutc(w_n515_53[2]),.din(w_n515_17[1]));
	jspl3 jspl3_w_n515_54(.douta(w_n515_54[0]),.doutb(w_n515_54[1]),.doutc(w_n515_54[2]),.din(w_n515_17[2]));
	jspl3 jspl3_w_n515_55(.douta(w_n515_55[0]),.doutb(w_n515_55[1]),.doutc(w_n515_55[2]),.din(w_n515_18[0]));
	jspl3 jspl3_w_n515_56(.douta(w_n515_56[0]),.doutb(w_n515_56[1]),.doutc(w_n515_56[2]),.din(w_n515_18[1]));
	jspl3 jspl3_w_n515_57(.douta(w_n515_57[0]),.doutb(w_n515_57[1]),.doutc(w_n515_57[2]),.din(w_n515_18[2]));
	jspl3 jspl3_w_n515_58(.douta(w_n515_58[0]),.doutb(w_n515_58[1]),.doutc(w_n515_58[2]),.din(w_n515_19[0]));
	jspl3 jspl3_w_n515_59(.douta(w_n515_59[0]),.doutb(w_n515_59[1]),.doutc(w_n515_59[2]),.din(w_n515_19[1]));
	jspl3 jspl3_w_n515_60(.douta(w_n515_60[0]),.doutb(w_n515_60[1]),.doutc(w_n515_60[2]),.din(w_n515_19[2]));
	jspl3 jspl3_w_n515_61(.douta(w_n515_61[0]),.doutb(w_n515_61[1]),.doutc(w_n515_61[2]),.din(w_n515_20[0]));
	jspl3 jspl3_w_n515_62(.douta(w_n515_62[0]),.doutb(w_n515_62[1]),.doutc(w_n515_62[2]),.din(w_n515_20[1]));
	jspl3 jspl3_w_n515_63(.douta(w_n515_63[0]),.doutb(w_n515_63[1]),.doutc(w_n515_63[2]),.din(w_n515_20[2]));
	jspl3 jspl3_w_n515_64(.douta(w_n515_64[0]),.doutb(w_n515_64[1]),.doutc(w_n515_64[2]),.din(w_n515_21[0]));
	jspl3 jspl3_w_n515_65(.douta(w_n515_65[0]),.doutb(w_n515_65[1]),.doutc(w_n515_65[2]),.din(w_n515_21[1]));
	jspl3 jspl3_w_n515_66(.douta(w_n515_66[0]),.doutb(w_n515_66[1]),.doutc(w_n515_66[2]),.din(w_n515_21[2]));
	jspl3 jspl3_w_n515_67(.douta(w_n515_67[0]),.doutb(w_n515_67[1]),.doutc(w_n515_67[2]),.din(w_n515_22[0]));
	jspl3 jspl3_w_n515_68(.douta(w_n515_68[0]),.doutb(w_n515_68[1]),.doutc(w_n515_68[2]),.din(w_n515_22[1]));
	jspl3 jspl3_w_n515_69(.douta(w_n515_69[0]),.doutb(w_n515_69[1]),.doutc(w_n515_69[2]),.din(w_n515_22[2]));
	jspl3 jspl3_w_n515_70(.douta(w_n515_70[0]),.doutb(w_n515_70[1]),.doutc(w_n515_70[2]),.din(w_n515_23[0]));
	jspl3 jspl3_w_n515_71(.douta(w_n515_71[0]),.doutb(w_n515_71[1]),.doutc(w_n515_71[2]),.din(w_n515_23[1]));
	jspl3 jspl3_w_n515_72(.douta(w_n515_72[0]),.doutb(w_n515_72[1]),.doutc(w_n515_72[2]),.din(w_n515_23[2]));
	jspl jspl_w_n515_73(.douta(w_n515_73[0]),.doutb(w_n515_73[1]),.din(w_n515_24[0]));
	jspl3 jspl3_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.doutc(w_n518_0[2]),.din(n518));
	jspl3 jspl3_w_n519_0(.douta(w_n519_0[0]),.doutb(w_n519_0[1]),.doutc(w_n519_0[2]),.din(n519));
	jspl3 jspl3_w_n521_0(.douta(w_n521_0[0]),.doutb(w_n521_0[1]),.doutc(w_n521_0[2]),.din(n521));
	jspl3 jspl3_w_n521_1(.douta(w_n521_1[0]),.doutb(w_n521_1[1]),.doutc(w_n521_1[2]),.din(w_n521_0[0]));
	jspl jspl_w_n522_0(.douta(w_n522_0[0]),.doutb(w_n522_0[1]),.din(n522));
	jspl3 jspl3_w_n523_0(.douta(w_n523_0[0]),.doutb(w_n523_0[1]),.doutc(w_n523_0[2]),.din(n523));
	jspl jspl_w_n524_0(.douta(w_n524_0[0]),.doutb(w_n524_0[1]),.din(n524));
	jspl3 jspl3_w_n526_0(.douta(w_n526_0[0]),.doutb(w_n526_0[1]),.doutc(w_n526_0[2]),.din(n526));
	jspl jspl_w_n527_0(.douta(w_n527_0[0]),.doutb(w_n527_0[1]),.din(n527));
	jspl3 jspl3_w_n534_0(.douta(w_n534_0[0]),.doutb(w_n534_0[1]),.doutc(w_n534_0[2]),.din(n534));
	jspl jspl_w_n535_0(.douta(w_n535_0[0]),.doutb(w_n535_0[1]),.din(n535));
	jspl jspl_w_n538_0(.douta(w_n538_0[0]),.doutb(w_n538_0[1]),.din(n538));
	jspl jspl_w_n539_0(.douta(w_n539_0[0]),.doutb(w_n539_0[1]),.din(n539));
	jspl3 jspl3_w_n544_0(.douta(w_n544_0[0]),.doutb(w_n544_0[1]),.doutc(w_n544_0[2]),.din(n544));
	jspl3 jspl3_w_n546_0(.douta(w_n546_0[0]),.doutb(w_n546_0[1]),.doutc(w_n546_0[2]),.din(n546));
	jspl jspl_w_n547_0(.douta(w_n547_0[0]),.doutb(w_n547_0[1]),.din(n547));
	jspl3 jspl3_w_n551_0(.douta(w_n551_0[0]),.doutb(w_n551_0[1]),.doutc(w_n551_0[2]),.din(n551));
	jspl3 jspl3_w_n554_0(.douta(w_n554_0[0]),.doutb(w_n554_0[1]),.doutc(w_n554_0[2]),.din(n554));
	jspl jspl_w_n555_0(.douta(w_n555_0[0]),.doutb(w_n555_0[1]),.din(n555));
	jspl3 jspl3_w_n559_0(.douta(w_n559_0[0]),.doutb(w_n559_0[1]),.doutc(w_n559_0[2]),.din(n559));
	jspl3 jspl3_w_n561_0(.douta(w_n561_0[0]),.doutb(w_n561_0[1]),.doutc(w_n561_0[2]),.din(n561));
	jspl jspl_w_n562_0(.douta(w_n562_0[0]),.doutb(w_n562_0[1]),.din(n562));
	jspl3 jspl3_w_n566_0(.douta(w_n566_0[0]),.doutb(w_n566_0[1]),.doutc(w_n566_0[2]),.din(n566));
	jspl3 jspl3_w_n569_0(.douta(w_n569_0[0]),.doutb(w_n569_0[1]),.doutc(w_n569_0[2]),.din(n569));
	jspl jspl_w_n570_0(.douta(w_n570_0[0]),.doutb(w_n570_0[1]),.din(n570));
	jspl jspl_w_n572_0(.douta(w_n572_0[0]),.doutb(w_n572_0[1]),.din(n572));
	jspl jspl_w_n575_0(.douta(w_n575_0[0]),.doutb(w_n575_0[1]),.din(n575));
	jspl jspl_w_n576_0(.douta(w_n576_0[0]),.doutb(w_n576_0[1]),.din(n576));
	jspl jspl_w_n581_0(.douta(w_n581_0[0]),.doutb(w_n581_0[1]),.din(n581));
	jspl jspl_w_n582_0(.douta(w_n582_0[0]),.doutb(w_n582_0[1]),.din(n582));
	jspl3 jspl3_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.doutc(w_n588_0[2]),.din(n588));
	jspl3 jspl3_w_n589_0(.douta(w_n589_0[0]),.doutb(w_n589_0[1]),.doutc(w_n589_0[2]),.din(n589));
	jspl jspl_w_n589_1(.douta(w_n589_1[0]),.doutb(w_n589_1[1]),.din(w_n589_0[0]));
	jspl jspl_w_n590_0(.douta(w_n590_0[0]),.doutb(w_n590_0[1]),.din(n590));
	jspl3 jspl3_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.doutc(w_n591_0[2]),.din(n591));
	jspl jspl_w_n592_0(.douta(w_n592_0[0]),.doutb(w_n592_0[1]),.din(n592));
	jspl3 jspl3_w_n594_0(.douta(w_n594_0[0]),.doutb(w_n594_0[1]),.doutc(w_n594_0[2]),.din(n594));
	jspl jspl_w_n595_0(.douta(w_n595_0[0]),.doutb(w_n595_0[1]),.din(n595));
	jspl jspl_w_n610_0(.douta(w_n610_0[0]),.doutb(w_n610_0[1]),.din(n610));
	jspl jspl_w_n626_0(.douta(w_n626_0[0]),.doutb(w_n626_0[1]),.din(n626));
	jspl jspl_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.din(n627));
	jspl jspl_w_n630_0(.douta(w_n630_0[0]),.doutb(w_n630_0[1]),.din(n630));
	jspl3 jspl3_w_n632_0(.douta(w_n632_0[0]),.doutb(w_n632_0[1]),.doutc(w_n632_0[2]),.din(n632));
	jspl3 jspl3_w_n635_0(.douta(w_n635_0[0]),.doutb(w_n635_0[1]),.doutc(w_n635_0[2]),.din(n635));
	jspl3 jspl3_w_n635_1(.douta(w_n635_1[0]),.doutb(w_n635_1[1]),.doutc(w_n635_1[2]),.din(w_n635_0[0]));
	jspl3 jspl3_w_n635_2(.douta(w_n635_2[0]),.doutb(w_n635_2[1]),.doutc(w_n635_2[2]),.din(w_n635_0[1]));
	jspl3 jspl3_w_n635_3(.douta(w_n635_3[0]),.doutb(w_n635_3[1]),.doutc(w_n635_3[2]),.din(w_n635_0[2]));
	jspl3 jspl3_w_n635_4(.douta(w_n635_4[0]),.doutb(w_n635_4[1]),.doutc(w_n635_4[2]),.din(w_n635_1[0]));
	jspl3 jspl3_w_n635_5(.douta(w_n635_5[0]),.doutb(w_n635_5[1]),.doutc(w_n635_5[2]),.din(w_n635_1[1]));
	jspl3 jspl3_w_n635_6(.douta(w_n635_6[0]),.doutb(w_n635_6[1]),.doutc(w_n635_6[2]),.din(w_n635_1[2]));
	jspl3 jspl3_w_n635_7(.douta(w_n635_7[0]),.doutb(w_n635_7[1]),.doutc(w_n635_7[2]),.din(w_n635_2[0]));
	jspl3 jspl3_w_n635_8(.douta(w_n635_8[0]),.doutb(w_n635_8[1]),.doutc(w_n635_8[2]),.din(w_n635_2[1]));
	jspl3 jspl3_w_n635_9(.douta(w_n635_9[0]),.doutb(w_n635_9[1]),.doutc(w_n635_9[2]),.din(w_n635_2[2]));
	jspl3 jspl3_w_n635_10(.douta(w_n635_10[0]),.doutb(w_n635_10[1]),.doutc(w_n635_10[2]),.din(w_n635_3[0]));
	jspl3 jspl3_w_n635_11(.douta(w_n635_11[0]),.doutb(w_n635_11[1]),.doutc(w_n635_11[2]),.din(w_n635_3[1]));
	jspl3 jspl3_w_n635_12(.douta(w_n635_12[0]),.doutb(w_n635_12[1]),.doutc(w_n635_12[2]),.din(w_n635_3[2]));
	jspl3 jspl3_w_n635_13(.douta(w_n635_13[0]),.doutb(w_n635_13[1]),.doutc(w_n635_13[2]),.din(w_n635_4[0]));
	jspl3 jspl3_w_n635_14(.douta(w_n635_14[0]),.doutb(w_n635_14[1]),.doutc(w_n635_14[2]),.din(w_n635_4[1]));
	jspl3 jspl3_w_n635_15(.douta(w_n635_15[0]),.doutb(w_n635_15[1]),.doutc(w_n635_15[2]),.din(w_n635_4[2]));
	jspl3 jspl3_w_n635_16(.douta(w_n635_16[0]),.doutb(w_n635_16[1]),.doutc(w_n635_16[2]),.din(w_n635_5[0]));
	jspl3 jspl3_w_n635_17(.douta(w_n635_17[0]),.doutb(w_n635_17[1]),.doutc(w_n635_17[2]),.din(w_n635_5[1]));
	jspl3 jspl3_w_n635_18(.douta(w_n635_18[0]),.doutb(w_n635_18[1]),.doutc(w_n635_18[2]),.din(w_n635_5[2]));
	jspl3 jspl3_w_n635_19(.douta(w_n635_19[0]),.doutb(w_n635_19[1]),.doutc(w_n635_19[2]),.din(w_n635_6[0]));
	jspl3 jspl3_w_n635_20(.douta(w_n635_20[0]),.doutb(w_n635_20[1]),.doutc(w_n635_20[2]),.din(w_n635_6[1]));
	jspl3 jspl3_w_n635_21(.douta(w_n635_21[0]),.doutb(w_n635_21[1]),.doutc(w_n635_21[2]),.din(w_n635_6[2]));
	jspl3 jspl3_w_n635_22(.douta(w_n635_22[0]),.doutb(w_n635_22[1]),.doutc(w_n635_22[2]),.din(w_n635_7[0]));
	jspl3 jspl3_w_n635_23(.douta(w_n635_23[0]),.doutb(w_n635_23[1]),.doutc(w_n635_23[2]),.din(w_n635_7[1]));
	jspl3 jspl3_w_n635_24(.douta(w_n635_24[0]),.doutb(w_n635_24[1]),.doutc(w_n635_24[2]),.din(w_n635_7[2]));
	jspl3 jspl3_w_n635_25(.douta(w_n635_25[0]),.doutb(w_n635_25[1]),.doutc(w_n635_25[2]),.din(w_n635_8[0]));
	jspl3 jspl3_w_n635_26(.douta(w_n635_26[0]),.doutb(w_n635_26[1]),.doutc(w_n635_26[2]),.din(w_n635_8[1]));
	jspl3 jspl3_w_n635_27(.douta(w_n635_27[0]),.doutb(w_n635_27[1]),.doutc(w_n635_27[2]),.din(w_n635_8[2]));
	jspl3 jspl3_w_n635_28(.douta(w_n635_28[0]),.doutb(w_n635_28[1]),.doutc(w_n635_28[2]),.din(w_n635_9[0]));
	jspl3 jspl3_w_n635_29(.douta(w_n635_29[0]),.doutb(w_n635_29[1]),.doutc(w_n635_29[2]),.din(w_n635_9[1]));
	jspl3 jspl3_w_n635_30(.douta(w_n635_30[0]),.doutb(w_n635_30[1]),.doutc(w_n635_30[2]),.din(w_n635_9[2]));
	jspl3 jspl3_w_n635_31(.douta(w_n635_31[0]),.doutb(w_n635_31[1]),.doutc(w_n635_31[2]),.din(w_n635_10[0]));
	jspl3 jspl3_w_n635_32(.douta(w_n635_32[0]),.doutb(w_n635_32[1]),.doutc(w_n635_32[2]),.din(w_n635_10[1]));
	jspl3 jspl3_w_n635_33(.douta(w_n635_33[0]),.doutb(w_n635_33[1]),.doutc(w_n635_33[2]),.din(w_n635_10[2]));
	jspl3 jspl3_w_n635_34(.douta(w_n635_34[0]),.doutb(w_n635_34[1]),.doutc(w_n635_34[2]),.din(w_n635_11[0]));
	jspl3 jspl3_w_n635_35(.douta(w_n635_35[0]),.doutb(w_n635_35[1]),.doutc(w_n635_35[2]),.din(w_n635_11[1]));
	jspl3 jspl3_w_n635_36(.douta(w_n635_36[0]),.doutb(w_n635_36[1]),.doutc(w_n635_36[2]),.din(w_n635_11[2]));
	jspl3 jspl3_w_n635_37(.douta(w_n635_37[0]),.doutb(w_n635_37[1]),.doutc(w_n635_37[2]),.din(w_n635_12[0]));
	jspl3 jspl3_w_n635_38(.douta(w_n635_38[0]),.doutb(w_n635_38[1]),.doutc(w_n635_38[2]),.din(w_n635_12[1]));
	jspl3 jspl3_w_n635_39(.douta(w_n635_39[0]),.doutb(w_n635_39[1]),.doutc(w_n635_39[2]),.din(w_n635_12[2]));
	jspl3 jspl3_w_n635_40(.douta(w_n635_40[0]),.doutb(w_n635_40[1]),.doutc(w_n635_40[2]),.din(w_n635_13[0]));
	jspl3 jspl3_w_n635_41(.douta(w_n635_41[0]),.doutb(w_n635_41[1]),.doutc(w_n635_41[2]),.din(w_n635_13[1]));
	jspl3 jspl3_w_n635_42(.douta(w_n635_42[0]),.doutb(w_n635_42[1]),.doutc(w_n635_42[2]),.din(w_n635_13[2]));
	jspl3 jspl3_w_n635_43(.douta(w_n635_43[0]),.doutb(w_n635_43[1]),.doutc(w_n635_43[2]),.din(w_n635_14[0]));
	jspl3 jspl3_w_n635_44(.douta(w_n635_44[0]),.doutb(w_n635_44[1]),.doutc(w_n635_44[2]),.din(w_n635_14[1]));
	jspl3 jspl3_w_n635_45(.douta(w_n635_45[0]),.doutb(w_n635_45[1]),.doutc(w_n635_45[2]),.din(w_n635_14[2]));
	jspl3 jspl3_w_n635_46(.douta(w_n635_46[0]),.doutb(w_n635_46[1]),.doutc(w_n635_46[2]),.din(w_n635_15[0]));
	jspl3 jspl3_w_n635_47(.douta(w_n635_47[0]),.doutb(w_n635_47[1]),.doutc(w_n635_47[2]),.din(w_n635_15[1]));
	jspl3 jspl3_w_n635_48(.douta(w_n635_48[0]),.doutb(w_n635_48[1]),.doutc(w_n635_48[2]),.din(w_n635_15[2]));
	jspl3 jspl3_w_n635_49(.douta(w_n635_49[0]),.doutb(w_n635_49[1]),.doutc(w_n635_49[2]),.din(w_n635_16[0]));
	jspl3 jspl3_w_n635_50(.douta(w_n635_50[0]),.doutb(w_n635_50[1]),.doutc(w_n635_50[2]),.din(w_n635_16[1]));
	jspl3 jspl3_w_n635_51(.douta(w_n635_51[0]),.doutb(w_n635_51[1]),.doutc(w_n635_51[2]),.din(w_n635_16[2]));
	jspl3 jspl3_w_n635_52(.douta(w_n635_52[0]),.doutb(w_n635_52[1]),.doutc(w_n635_52[2]),.din(w_n635_17[0]));
	jspl3 jspl3_w_n635_53(.douta(w_n635_53[0]),.doutb(w_n635_53[1]),.doutc(w_n635_53[2]),.din(w_n635_17[1]));
	jspl3 jspl3_w_n635_54(.douta(w_n635_54[0]),.doutb(w_n635_54[1]),.doutc(w_n635_54[2]),.din(w_n635_17[2]));
	jspl3 jspl3_w_n635_55(.douta(w_n635_55[0]),.doutb(w_n635_55[1]),.doutc(w_n635_55[2]),.din(w_n635_18[0]));
	jspl3 jspl3_w_n635_56(.douta(w_n635_56[0]),.doutb(w_n635_56[1]),.doutc(w_n635_56[2]),.din(w_n635_18[1]));
	jspl3 jspl3_w_n635_57(.douta(w_n635_57[0]),.doutb(w_n635_57[1]),.doutc(w_n635_57[2]),.din(w_n635_18[2]));
	jspl3 jspl3_w_n635_58(.douta(w_n635_58[0]),.doutb(w_n635_58[1]),.doutc(w_n635_58[2]),.din(w_n635_19[0]));
	jspl3 jspl3_w_n635_59(.douta(w_n635_59[0]),.doutb(w_n635_59[1]),.doutc(w_n635_59[2]),.din(w_n635_19[1]));
	jspl3 jspl3_w_n635_60(.douta(w_n635_60[0]),.doutb(w_n635_60[1]),.doutc(w_n635_60[2]),.din(w_n635_19[2]));
	jspl3 jspl3_w_n635_61(.douta(w_n635_61[0]),.doutb(w_n635_61[1]),.doutc(w_n635_61[2]),.din(w_n635_20[0]));
	jspl3 jspl3_w_n635_62(.douta(w_n635_62[0]),.doutb(w_n635_62[1]),.doutc(w_n635_62[2]),.din(w_n635_20[1]));
	jspl3 jspl3_w_n635_63(.douta(w_n635_63[0]),.doutb(w_n635_63[1]),.doutc(w_n635_63[2]),.din(w_n635_20[2]));
	jspl3 jspl3_w_n635_64(.douta(w_n635_64[0]),.doutb(w_n635_64[1]),.doutc(w_n635_64[2]),.din(w_n635_21[0]));
	jspl3 jspl3_w_n635_65(.douta(w_n635_65[0]),.doutb(w_n635_65[1]),.doutc(w_n635_65[2]),.din(w_n635_21[1]));
	jspl3 jspl3_w_n635_66(.douta(w_n635_66[0]),.doutb(w_n635_66[1]),.doutc(w_n635_66[2]),.din(w_n635_21[2]));
	jspl3 jspl3_w_n635_67(.douta(w_n635_67[0]),.doutb(w_n635_67[1]),.doutc(w_n635_67[2]),.din(w_n635_22[0]));
	jspl3 jspl3_w_n635_68(.douta(w_n635_68[0]),.doutb(w_n635_68[1]),.doutc(w_n635_68[2]),.din(w_n635_22[1]));
	jspl3 jspl3_w_n635_69(.douta(w_n635_69[0]),.doutb(w_n635_69[1]),.doutc(w_n635_69[2]),.din(w_n635_22[2]));
	jspl3 jspl3_w_n635_70(.douta(w_n635_70[0]),.doutb(w_n635_70[1]),.doutc(w_n635_70[2]),.din(w_n635_23[0]));
	jspl3 jspl3_w_n639_0(.douta(w_n639_0[0]),.doutb(w_n639_0[1]),.doutc(w_n639_0[2]),.din(n639));
	jspl jspl_w_n640_0(.douta(w_n640_0[0]),.doutb(w_n640_0[1]),.din(n640));
	jspl jspl_w_n642_0(.douta(w_n642_0[0]),.doutb(w_n642_0[1]),.din(n642));
	jspl jspl_w_n647_0(.douta(w_n647_0[0]),.doutb(w_n647_0[1]),.din(n647));
	jspl jspl_w_n648_0(.douta(w_n648_0[0]),.doutb(w_n648_0[1]),.din(n648));
	jspl3 jspl3_w_n650_0(.douta(w_n650_0[0]),.doutb(w_n650_0[1]),.doutc(w_n650_0[2]),.din(n650));
	jspl jspl_w_n651_0(.douta(w_n651_0[0]),.doutb(w_n651_0[1]),.din(n651));
	jspl jspl_w_n655_0(.douta(w_n655_0[0]),.doutb(w_n655_0[1]),.din(n655));
	jspl3 jspl3_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.doutc(w_n657_0[2]),.din(n657));
	jspl jspl_w_n658_0(.douta(w_n658_0[0]),.doutb(w_n658_0[1]),.din(n658));
	jspl jspl_w_n662_0(.douta(w_n662_0[0]),.doutb(w_n662_0[1]),.din(n662));
	jspl jspl_w_n663_0(.douta(w_n663_0[0]),.doutb(w_n663_0[1]),.din(n663));
	jspl3 jspl3_w_n665_0(.douta(w_n665_0[0]),.doutb(w_n665_0[1]),.doutc(w_n665_0[2]),.din(n665));
	jspl jspl_w_n666_0(.douta(w_n666_0[0]),.doutb(w_n666_0[1]),.din(n666));
	jspl jspl_w_n670_0(.douta(w_n670_0[0]),.doutb(w_n670_0[1]),.din(n670));
	jspl3 jspl3_w_n672_0(.douta(w_n672_0[0]),.doutb(w_n672_0[1]),.doutc(w_n672_0[2]),.din(n672));
	jspl jspl_w_n673_0(.douta(w_n673_0[0]),.doutb(w_n673_0[1]),.din(n673));
	jspl jspl_w_n677_0(.douta(w_n677_0[0]),.doutb(w_n677_0[1]),.din(n677));
	jspl jspl_w_n678_0(.douta(w_n678_0[0]),.doutb(w_n678_0[1]),.din(n678));
	jspl jspl_w_n680_0(.douta(w_n680_0[0]),.doutb(w_n680_0[1]),.din(n680));
	jspl3 jspl3_w_n681_0(.douta(w_n681_0[0]),.doutb(w_n681_0[1]),.doutc(w_n681_0[2]),.din(n681));
	jspl jspl_w_n681_1(.douta(w_n681_1[0]),.doutb(w_n681_1[1]),.din(w_n681_0[0]));
	jspl3 jspl3_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.doutc(w_n682_0[2]),.din(n682));
	jspl jspl_w_n686_0(.douta(w_n686_0[0]),.doutb(w_n686_0[1]),.din(n686));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_n687_0[1]),.din(n687));
	jspl jspl_w_n701_0(.douta(w_n701_0[0]),.doutb(w_n701_0[1]),.din(n701));
	jspl jspl_w_n708_0(.douta(w_n708_0[0]),.doutb(w_n708_0[1]),.din(n708));
	jspl jspl_w_n715_0(.douta(w_n715_0[0]),.doutb(w_n715_0[1]),.din(n715));
	jspl jspl_w_n720_0(.douta(w_n720_0[0]),.doutb(w_n720_0[1]),.din(n720));
	jspl jspl_w_n721_0(.douta(w_n721_0[0]),.doutb(w_n721_0[1]),.din(n721));
	jspl jspl_w_n723_0(.douta(w_n723_0[0]),.doutb(w_n723_0[1]),.din(n723));
	jspl jspl_w_n725_0(.douta(w_n725_0[0]),.doutb(w_n725_0[1]),.din(n725));
	jspl jspl_w_n726_0(.douta(w_n726_0[0]),.doutb(w_n726_0[1]),.din(n726));
	jspl jspl_w_n728_0(.douta(w_n728_0[0]),.doutb(w_n728_0[1]),.din(n728));
	jspl3 jspl3_w_n730_0(.douta(w_n730_0[0]),.doutb(w_n730_0[1]),.doutc(w_n730_0[2]),.din(n730));
	jspl3 jspl3_w_n730_1(.douta(w_n730_1[0]),.doutb(w_n730_1[1]),.doutc(w_n730_1[2]),.din(w_n730_0[0]));
	jspl jspl_w_n731_0(.douta(w_n731_0[0]),.doutb(w_n731_0[1]),.din(n731));
	jspl3 jspl3_w_n732_0(.douta(w_n732_0[0]),.doutb(w_n732_0[1]),.doutc(w_n732_0[2]),.din(n732));
	jspl jspl_w_n733_0(.douta(w_n733_0[0]),.doutb(w_n733_0[1]),.din(n733));
	jspl jspl_w_n736_0(.douta(w_n736_0[0]),.doutb(w_n736_0[1]),.din(n736));
	jspl jspl_w_n742_0(.douta(w_n742_0[0]),.doutb(w_n742_0[1]),.din(n742));
	jspl3 jspl3_w_n743_0(.douta(w_n743_0[0]),.doutb(w_n743_0[1]),.doutc(w_n743_0[2]),.din(n743));
	jspl3 jspl3_w_n743_1(.douta(w_n743_1[0]),.doutb(w_n743_1[1]),.doutc(w_n743_1[2]),.din(w_n743_0[0]));
	jspl3 jspl3_w_n743_2(.douta(w_n743_2[0]),.doutb(w_n743_2[1]),.doutc(w_n743_2[2]),.din(w_n743_0[1]));
	jspl3 jspl3_w_n743_3(.douta(w_n743_3[0]),.doutb(w_n743_3[1]),.doutc(w_n743_3[2]),.din(w_n743_0[2]));
	jspl3 jspl3_w_n743_4(.douta(w_n743_4[0]),.doutb(w_n743_4[1]),.doutc(w_n743_4[2]),.din(w_n743_1[0]));
	jspl3 jspl3_w_n743_5(.douta(w_n743_5[0]),.doutb(w_n743_5[1]),.doutc(w_n743_5[2]),.din(w_n743_1[1]));
	jspl3 jspl3_w_n743_6(.douta(w_n743_6[0]),.doutb(w_n743_6[1]),.doutc(w_n743_6[2]),.din(w_n743_1[2]));
	jspl3 jspl3_w_n743_7(.douta(w_n743_7[0]),.doutb(w_n743_7[1]),.doutc(w_n743_7[2]),.din(w_n743_2[0]));
	jspl3 jspl3_w_n743_8(.douta(w_n743_8[0]),.doutb(w_n743_8[1]),.doutc(w_n743_8[2]),.din(w_n743_2[1]));
	jspl3 jspl3_w_n743_9(.douta(w_n743_9[0]),.doutb(w_n743_9[1]),.doutc(w_n743_9[2]),.din(w_n743_2[2]));
	jspl3 jspl3_w_n743_10(.douta(w_n743_10[0]),.doutb(w_n743_10[1]),.doutc(w_n743_10[2]),.din(w_n743_3[0]));
	jspl3 jspl3_w_n743_11(.douta(w_n743_11[0]),.doutb(w_n743_11[1]),.doutc(w_n743_11[2]),.din(w_n743_3[1]));
	jspl3 jspl3_w_n743_12(.douta(w_n743_12[0]),.doutb(w_n743_12[1]),.doutc(w_n743_12[2]),.din(w_n743_3[2]));
	jspl3 jspl3_w_n743_13(.douta(w_n743_13[0]),.doutb(w_n743_13[1]),.doutc(w_n743_13[2]),.din(w_n743_4[0]));
	jspl3 jspl3_w_n743_14(.douta(w_n743_14[0]),.doutb(w_n743_14[1]),.doutc(w_n743_14[2]),.din(w_n743_4[1]));
	jspl3 jspl3_w_n743_15(.douta(w_n743_15[0]),.doutb(w_n743_15[1]),.doutc(w_n743_15[2]),.din(w_n743_4[2]));
	jspl3 jspl3_w_n743_16(.douta(w_n743_16[0]),.doutb(w_n743_16[1]),.doutc(w_n743_16[2]),.din(w_n743_5[0]));
	jspl3 jspl3_w_n743_17(.douta(w_n743_17[0]),.doutb(w_n743_17[1]),.doutc(w_n743_17[2]),.din(w_n743_5[1]));
	jspl3 jspl3_w_n743_18(.douta(w_n743_18[0]),.doutb(w_n743_18[1]),.doutc(w_n743_18[2]),.din(w_n743_5[2]));
	jspl3 jspl3_w_n743_19(.douta(w_n743_19[0]),.doutb(w_n743_19[1]),.doutc(w_n743_19[2]),.din(w_n743_6[0]));
	jspl3 jspl3_w_n743_20(.douta(w_n743_20[0]),.doutb(w_n743_20[1]),.doutc(w_n743_20[2]),.din(w_n743_6[1]));
	jspl3 jspl3_w_n743_21(.douta(w_n743_21[0]),.doutb(w_n743_21[1]),.doutc(w_n743_21[2]),.din(w_n743_6[2]));
	jspl3 jspl3_w_n743_22(.douta(w_n743_22[0]),.doutb(w_n743_22[1]),.doutc(w_n743_22[2]),.din(w_n743_7[0]));
	jspl3 jspl3_w_n743_23(.douta(w_n743_23[0]),.doutb(w_n743_23[1]),.doutc(w_n743_23[2]),.din(w_n743_7[1]));
	jspl3 jspl3_w_n743_24(.douta(w_n743_24[0]),.doutb(w_n743_24[1]),.doutc(w_n743_24[2]),.din(w_n743_7[2]));
	jspl3 jspl3_w_n743_25(.douta(w_n743_25[0]),.doutb(w_n743_25[1]),.doutc(w_n743_25[2]),.din(w_n743_8[0]));
	jspl3 jspl3_w_n743_26(.douta(w_n743_26[0]),.doutb(w_n743_26[1]),.doutc(w_n743_26[2]),.din(w_n743_8[1]));
	jspl3 jspl3_w_n743_27(.douta(w_n743_27[0]),.doutb(w_n743_27[1]),.doutc(w_n743_27[2]),.din(w_n743_8[2]));
	jspl3 jspl3_w_n743_28(.douta(w_n743_28[0]),.doutb(w_n743_28[1]),.doutc(w_n743_28[2]),.din(w_n743_9[0]));
	jspl3 jspl3_w_n743_29(.douta(w_n743_29[0]),.doutb(w_n743_29[1]),.doutc(w_n743_29[2]),.din(w_n743_9[1]));
	jspl3 jspl3_w_n743_30(.douta(w_n743_30[0]),.doutb(w_n743_30[1]),.doutc(w_n743_30[2]),.din(w_n743_9[2]));
	jspl3 jspl3_w_n743_31(.douta(w_n743_31[0]),.doutb(w_n743_31[1]),.doutc(w_n743_31[2]),.din(w_n743_10[0]));
	jspl3 jspl3_w_n743_32(.douta(w_n743_32[0]),.doutb(w_n743_32[1]),.doutc(w_n743_32[2]),.din(w_n743_10[1]));
	jspl3 jspl3_w_n743_33(.douta(w_n743_33[0]),.doutb(w_n743_33[1]),.doutc(w_n743_33[2]),.din(w_n743_10[2]));
	jspl3 jspl3_w_n743_34(.douta(w_n743_34[0]),.doutb(w_n743_34[1]),.doutc(w_n743_34[2]),.din(w_n743_11[0]));
	jspl3 jspl3_w_n743_35(.douta(w_n743_35[0]),.doutb(w_n743_35[1]),.doutc(w_n743_35[2]),.din(w_n743_11[1]));
	jspl3 jspl3_w_n743_36(.douta(w_n743_36[0]),.doutb(w_n743_36[1]),.doutc(w_n743_36[2]),.din(w_n743_11[2]));
	jspl3 jspl3_w_n743_37(.douta(w_n743_37[0]),.doutb(w_n743_37[1]),.doutc(w_n743_37[2]),.din(w_n743_12[0]));
	jspl3 jspl3_w_n743_38(.douta(w_n743_38[0]),.doutb(w_n743_38[1]),.doutc(w_n743_38[2]),.din(w_n743_12[1]));
	jspl3 jspl3_w_n743_39(.douta(w_n743_39[0]),.doutb(w_n743_39[1]),.doutc(w_n743_39[2]),.din(w_n743_12[2]));
	jspl3 jspl3_w_n743_40(.douta(w_n743_40[0]),.doutb(w_n743_40[1]),.doutc(w_n743_40[2]),.din(w_n743_13[0]));
	jspl3 jspl3_w_n743_41(.douta(w_n743_41[0]),.doutb(w_n743_41[1]),.doutc(w_n743_41[2]),.din(w_n743_13[1]));
	jspl3 jspl3_w_n743_42(.douta(w_n743_42[0]),.doutb(w_n743_42[1]),.doutc(w_n743_42[2]),.din(w_n743_13[2]));
	jspl3 jspl3_w_n743_43(.douta(w_n743_43[0]),.doutb(w_n743_43[1]),.doutc(w_n743_43[2]),.din(w_n743_14[0]));
	jspl3 jspl3_w_n743_44(.douta(w_n743_44[0]),.doutb(w_n743_44[1]),.doutc(w_n743_44[2]),.din(w_n743_14[1]));
	jspl3 jspl3_w_n743_45(.douta(w_n743_45[0]),.doutb(w_n743_45[1]),.doutc(w_n743_45[2]),.din(w_n743_14[2]));
	jspl3 jspl3_w_n743_46(.douta(w_n743_46[0]),.doutb(w_n743_46[1]),.doutc(w_n743_46[2]),.din(w_n743_15[0]));
	jspl3 jspl3_w_n743_47(.douta(w_n743_47[0]),.doutb(w_n743_47[1]),.doutc(w_n743_47[2]),.din(w_n743_15[1]));
	jspl3 jspl3_w_n743_48(.douta(w_n743_48[0]),.doutb(w_n743_48[1]),.doutc(w_n743_48[2]),.din(w_n743_15[2]));
	jspl3 jspl3_w_n743_49(.douta(w_n743_49[0]),.doutb(w_n743_49[1]),.doutc(w_n743_49[2]),.din(w_n743_16[0]));
	jspl3 jspl3_w_n743_50(.douta(w_n743_50[0]),.doutb(w_n743_50[1]),.doutc(w_n743_50[2]),.din(w_n743_16[1]));
	jspl3 jspl3_w_n743_51(.douta(w_n743_51[0]),.doutb(w_n743_51[1]),.doutc(w_n743_51[2]),.din(w_n743_16[2]));
	jspl3 jspl3_w_n743_52(.douta(w_n743_52[0]),.doutb(w_n743_52[1]),.doutc(w_n743_52[2]),.din(w_n743_17[0]));
	jspl3 jspl3_w_n743_53(.douta(w_n743_53[0]),.doutb(w_n743_53[1]),.doutc(w_n743_53[2]),.din(w_n743_17[1]));
	jspl3 jspl3_w_n743_54(.douta(w_n743_54[0]),.doutb(w_n743_54[1]),.doutc(w_n743_54[2]),.din(w_n743_17[2]));
	jspl3 jspl3_w_n743_55(.douta(w_n743_55[0]),.doutb(w_n743_55[1]),.doutc(w_n743_55[2]),.din(w_n743_18[0]));
	jspl3 jspl3_w_n743_56(.douta(w_n743_56[0]),.doutb(w_n743_56[1]),.doutc(w_n743_56[2]),.din(w_n743_18[1]));
	jspl3 jspl3_w_n743_57(.douta(w_n743_57[0]),.doutb(w_n743_57[1]),.doutc(w_n743_57[2]),.din(w_n743_18[2]));
	jspl3 jspl3_w_n743_58(.douta(w_n743_58[0]),.doutb(w_n743_58[1]),.doutc(w_n743_58[2]),.din(w_n743_19[0]));
	jspl3 jspl3_w_n743_59(.douta(w_n743_59[0]),.doutb(w_n743_59[1]),.doutc(w_n743_59[2]),.din(w_n743_19[1]));
	jspl3 jspl3_w_n743_60(.douta(w_n743_60[0]),.doutb(w_n743_60[1]),.doutc(w_n743_60[2]),.din(w_n743_19[2]));
	jspl3 jspl3_w_n743_61(.douta(w_n743_61[0]),.doutb(w_n743_61[1]),.doutc(w_n743_61[2]),.din(w_n743_20[0]));
	jspl3 jspl3_w_n743_62(.douta(w_n743_62[0]),.doutb(w_n743_62[1]),.doutc(w_n743_62[2]),.din(w_n743_20[1]));
	jspl3 jspl3_w_n743_63(.douta(w_n743_63[0]),.doutb(w_n743_63[1]),.doutc(w_n743_63[2]),.din(w_n743_20[2]));
	jspl3 jspl3_w_n743_64(.douta(w_n743_64[0]),.doutb(w_n743_64[1]),.doutc(w_n743_64[2]),.din(w_n743_21[0]));
	jspl3 jspl3_w_n743_65(.douta(w_n743_65[0]),.doutb(w_n743_65[1]),.doutc(w_n743_65[2]),.din(w_n743_21[1]));
	jspl3 jspl3_w_n743_66(.douta(w_n743_66[0]),.doutb(w_n743_66[1]),.doutc(w_n743_66[2]),.din(w_n743_21[2]));
	jspl3 jspl3_w_n743_67(.douta(w_n743_67[0]),.doutb(w_n743_67[1]),.doutc(w_n743_67[2]),.din(w_n743_22[0]));
	jspl3 jspl3_w_n743_68(.douta(w_n743_68[0]),.doutb(w_n743_68[1]),.doutc(w_n743_68[2]),.din(w_n743_22[1]));
	jspl3 jspl3_w_n743_69(.douta(w_n743_69[0]),.doutb(w_n743_69[1]),.doutc(w_n743_69[2]),.din(w_n743_22[2]));
	jspl3 jspl3_w_n743_70(.douta(w_n743_70[0]),.doutb(w_n743_70[1]),.doutc(w_n743_70[2]),.din(w_n743_23[0]));
	jspl3 jspl3_w_n745_0(.douta(w_n745_0[0]),.doutb(w_n745_0[1]),.doutc(w_n745_0[2]),.din(n745));
	jspl jspl_w_n746_0(.douta(w_n746_0[0]),.doutb(w_n746_0[1]),.din(n746));
	jspl3 jspl3_w_n753_0(.douta(w_n753_0[0]),.doutb(w_n753_0[1]),.doutc(w_n753_0[2]),.din(n753));
	jspl jspl_w_n754_0(.douta(w_n754_0[0]),.doutb(w_n754_0[1]),.din(n754));
	jspl jspl_w_n757_0(.douta(w_n757_0[0]),.doutb(w_n757_0[1]),.din(n757));
	jspl jspl_w_n762_0(.douta(w_n762_0[0]),.doutb(w_n762_0[1]),.din(n762));
	jspl3 jspl3_w_n764_0(.douta(w_n764_0[0]),.doutb(w_n764_0[1]),.doutc(w_n764_0[2]),.din(n764));
	jspl jspl_w_n765_0(.douta(w_n765_0[0]),.doutb(w_n765_0[1]),.din(n765));
	jspl3 jspl3_w_n769_0(.douta(w_n769_0[0]),.doutb(w_n769_0[1]),.doutc(w_n769_0[2]),.din(n769));
	jspl3 jspl3_w_n772_0(.douta(w_n772_0[0]),.doutb(w_n772_0[1]),.doutc(w_n772_0[2]),.din(n772));
	jspl jspl_w_n773_0(.douta(w_n773_0[0]),.doutb(w_n773_0[1]),.din(n773));
	jspl3 jspl3_w_n777_0(.douta(w_n777_0[0]),.doutb(w_n777_0[1]),.doutc(w_n777_0[2]),.din(n777));
	jspl3 jspl3_w_n779_0(.douta(w_n779_0[0]),.doutb(w_n779_0[1]),.doutc(w_n779_0[2]),.din(n779));
	jspl jspl_w_n780_0(.douta(w_n780_0[0]),.doutb(w_n780_0[1]),.din(n780));
	jspl3 jspl3_w_n784_0(.douta(w_n784_0[0]),.doutb(w_n784_0[1]),.doutc(w_n784_0[2]),.din(n784));
	jspl3 jspl3_w_n787_0(.douta(w_n787_0[0]),.doutb(w_n787_0[1]),.doutc(w_n787_0[2]),.din(n787));
	jspl jspl_w_n788_0(.douta(w_n788_0[0]),.doutb(w_n788_0[1]),.din(n788));
	jspl3 jspl3_w_n792_0(.douta(w_n792_0[0]),.doutb(w_n792_0[1]),.doutc(w_n792_0[2]),.din(n792));
	jspl3 jspl3_w_n794_0(.douta(w_n794_0[0]),.doutb(w_n794_0[1]),.doutc(w_n794_0[2]),.din(n794));
	jspl jspl_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.din(n795));
	jspl3 jspl3_w_n799_0(.douta(w_n799_0[0]),.doutb(w_n799_0[1]),.doutc(w_n799_0[2]),.din(n799));
	jspl3 jspl3_w_n802_0(.douta(w_n802_0[0]),.doutb(w_n802_0[1]),.doutc(w_n802_0[2]),.din(n802));
	jspl3 jspl3_w_n805_0(.douta(w_n805_0[0]),.doutb(w_n805_0[1]),.doutc(w_n805_0[2]),.din(n805));
	jspl jspl_w_n805_1(.douta(w_n805_1[0]),.doutb(w_n805_1[1]),.din(w_n805_0[0]));
	jspl3 jspl3_w_n806_0(.douta(w_n806_0[0]),.doutb(w_n806_0[1]),.doutc(w_n806_0[2]),.din(n806));
	jspl jspl_w_n808_0(.douta(w_n808_0[0]),.doutb(w_n808_0[1]),.din(n808));
	jspl jspl_w_n809_0(.douta(w_n809_0[0]),.doutb(w_n809_0[1]),.din(n809));
	jspl jspl_w_n816_0(.douta(w_n816_0[0]),.doutb(w_n816_0[1]),.din(n816));
	jspl jspl_w_n817_0(.douta(w_n817_0[0]),.doutb(w_n817_0[1]),.din(n817));
	jspl jspl_w_n819_0(.douta(w_n819_0[0]),.doutb(w_n819_0[1]),.din(n819));
	jspl jspl_w_n834_0(.douta(w_n834_0[0]),.doutb(w_n834_0[1]),.din(n834));
	jspl jspl_w_n838_0(.douta(w_n838_0[0]),.doutb(w_n838_0[1]),.din(n838));
	jspl jspl_w_n859_0(.douta(w_n859_0[0]),.doutb(w_n859_0[1]),.din(n859));
	jspl jspl_w_n860_0(.douta(w_n860_0[0]),.doutb(w_n860_0[1]),.din(n860));
	jspl3 jspl3_w_n863_0(.douta(w_n863_0[0]),.doutb(w_n863_0[1]),.doutc(w_n863_0[2]),.din(n863));
	jspl jspl_w_n864_0(.douta(w_n864_0[0]),.doutb(w_n864_0[1]),.din(n864));
	jspl3 jspl3_w_n865_0(.douta(w_n865_0[0]),.doutb(w_n865_0[1]),.doutc(w_n865_0[2]),.din(n865));
	jspl jspl_w_n865_1(.douta(w_n865_1[0]),.doutb(w_n865_1[1]),.din(w_n865_0[0]));
	jspl jspl_w_n866_0(.douta(w_n866_0[0]),.doutb(w_n866_0[1]),.din(n866));
	jspl3 jspl3_w_n867_0(.douta(w_n867_0[0]),.doutb(w_n867_0[1]),.doutc(w_n867_0[2]),.din(n867));
	jspl jspl_w_n868_0(.douta(w_n868_0[0]),.doutb(w_n868_0[1]),.din(n868));
	jspl3 jspl3_w_n870_0(.douta(w_n870_0[0]),.doutb(w_n870_0[1]),.doutc(w_n870_0[2]),.din(n870));
	jspl jspl_w_n871_0(.douta(w_n871_0[0]),.doutb(w_n871_0[1]),.din(n871));
	jspl3 jspl3_w_n876_0(.douta(w_n876_0[0]),.doutb(w_n876_0[1]),.doutc(w_n876_0[2]),.din(n876));
	jspl jspl_w_n876_1(.douta(w_n876_1[0]),.doutb(w_n876_1[1]),.din(w_n876_0[0]));
	jspl jspl_w_n881_0(.douta(w_n881_0[0]),.doutb(w_n881_0[1]),.din(n881));
	jspl jspl_w_n882_0(.douta(w_n882_0[0]),.doutb(w_n882_0[1]),.din(n882));
	jspl3 jspl3_w_n884_0(.douta(w_n884_0[0]),.doutb(w_n884_0[1]),.doutc(w_n884_0[2]),.din(n884));
	jspl3 jspl3_w_n884_1(.douta(w_n884_1[0]),.doutb(w_n884_1[1]),.doutc(w_n884_1[2]),.din(w_n884_0[0]));
	jspl3 jspl3_w_n884_2(.douta(w_n884_2[0]),.doutb(w_n884_2[1]),.doutc(w_n884_2[2]),.din(w_n884_0[1]));
	jspl3 jspl3_w_n884_3(.douta(w_n884_3[0]),.doutb(w_n884_3[1]),.doutc(w_n884_3[2]),.din(w_n884_0[2]));
	jspl3 jspl3_w_n884_4(.douta(w_n884_4[0]),.doutb(w_n884_4[1]),.doutc(w_n884_4[2]),.din(w_n884_1[0]));
	jspl3 jspl3_w_n884_5(.douta(w_n884_5[0]),.doutb(w_n884_5[1]),.doutc(w_n884_5[2]),.din(w_n884_1[1]));
	jspl3 jspl3_w_n884_6(.douta(w_n884_6[0]),.doutb(w_n884_6[1]),.doutc(w_n884_6[2]),.din(w_n884_1[2]));
	jspl3 jspl3_w_n884_7(.douta(w_n884_7[0]),.doutb(w_n884_7[1]),.doutc(w_n884_7[2]),.din(w_n884_2[0]));
	jspl3 jspl3_w_n884_8(.douta(w_n884_8[0]),.doutb(w_n884_8[1]),.doutc(w_n884_8[2]),.din(w_n884_2[1]));
	jspl3 jspl3_w_n884_9(.douta(w_n884_9[0]),.doutb(w_n884_9[1]),.doutc(w_n884_9[2]),.din(w_n884_2[2]));
	jspl3 jspl3_w_n884_10(.douta(w_n884_10[0]),.doutb(w_n884_10[1]),.doutc(w_n884_10[2]),.din(w_n884_3[0]));
	jspl3 jspl3_w_n884_11(.douta(w_n884_11[0]),.doutb(w_n884_11[1]),.doutc(w_n884_11[2]),.din(w_n884_3[1]));
	jspl3 jspl3_w_n884_12(.douta(w_n884_12[0]),.doutb(w_n884_12[1]),.doutc(w_n884_12[2]),.din(w_n884_3[2]));
	jspl3 jspl3_w_n884_13(.douta(w_n884_13[0]),.doutb(w_n884_13[1]),.doutc(w_n884_13[2]),.din(w_n884_4[0]));
	jspl3 jspl3_w_n884_14(.douta(w_n884_14[0]),.doutb(w_n884_14[1]),.doutc(w_n884_14[2]),.din(w_n884_4[1]));
	jspl3 jspl3_w_n884_15(.douta(w_n884_15[0]),.doutb(w_n884_15[1]),.doutc(w_n884_15[2]),.din(w_n884_4[2]));
	jspl3 jspl3_w_n884_16(.douta(w_n884_16[0]),.doutb(w_n884_16[1]),.doutc(w_n884_16[2]),.din(w_n884_5[0]));
	jspl3 jspl3_w_n884_17(.douta(w_n884_17[0]),.doutb(w_n884_17[1]),.doutc(w_n884_17[2]),.din(w_n884_5[1]));
	jspl3 jspl3_w_n884_18(.douta(w_n884_18[0]),.doutb(w_n884_18[1]),.doutc(w_n884_18[2]),.din(w_n884_5[2]));
	jspl3 jspl3_w_n884_19(.douta(w_n884_19[0]),.doutb(w_n884_19[1]),.doutc(w_n884_19[2]),.din(w_n884_6[0]));
	jspl3 jspl3_w_n884_20(.douta(w_n884_20[0]),.doutb(w_n884_20[1]),.doutc(w_n884_20[2]),.din(w_n884_6[1]));
	jspl3 jspl3_w_n884_21(.douta(w_n884_21[0]),.doutb(w_n884_21[1]),.doutc(w_n884_21[2]),.din(w_n884_6[2]));
	jspl3 jspl3_w_n884_22(.douta(w_n884_22[0]),.doutb(w_n884_22[1]),.doutc(w_n884_22[2]),.din(w_n884_7[0]));
	jspl3 jspl3_w_n884_23(.douta(w_n884_23[0]),.doutb(w_n884_23[1]),.doutc(w_n884_23[2]),.din(w_n884_7[1]));
	jspl3 jspl3_w_n884_24(.douta(w_n884_24[0]),.doutb(w_n884_24[1]),.doutc(w_n884_24[2]),.din(w_n884_7[2]));
	jspl3 jspl3_w_n884_25(.douta(w_n884_25[0]),.doutb(w_n884_25[1]),.doutc(w_n884_25[2]),.din(w_n884_8[0]));
	jspl3 jspl3_w_n884_26(.douta(w_n884_26[0]),.doutb(w_n884_26[1]),.doutc(w_n884_26[2]),.din(w_n884_8[1]));
	jspl3 jspl3_w_n884_27(.douta(w_n884_27[0]),.doutb(w_n884_27[1]),.doutc(w_n884_27[2]),.din(w_n884_8[2]));
	jspl3 jspl3_w_n884_28(.douta(w_n884_28[0]),.doutb(w_n884_28[1]),.doutc(w_n884_28[2]),.din(w_n884_9[0]));
	jspl3 jspl3_w_n884_29(.douta(w_n884_29[0]),.doutb(w_n884_29[1]),.doutc(w_n884_29[2]),.din(w_n884_9[1]));
	jspl3 jspl3_w_n884_30(.douta(w_n884_30[0]),.doutb(w_n884_30[1]),.doutc(w_n884_30[2]),.din(w_n884_9[2]));
	jspl3 jspl3_w_n884_31(.douta(w_n884_31[0]),.doutb(w_n884_31[1]),.doutc(w_n884_31[2]),.din(w_n884_10[0]));
	jspl3 jspl3_w_n884_32(.douta(w_n884_32[0]),.doutb(w_n884_32[1]),.doutc(w_n884_32[2]),.din(w_n884_10[1]));
	jspl3 jspl3_w_n884_33(.douta(w_n884_33[0]),.doutb(w_n884_33[1]),.doutc(w_n884_33[2]),.din(w_n884_10[2]));
	jspl3 jspl3_w_n884_34(.douta(w_n884_34[0]),.doutb(w_n884_34[1]),.doutc(w_n884_34[2]),.din(w_n884_11[0]));
	jspl3 jspl3_w_n884_35(.douta(w_n884_35[0]),.doutb(w_n884_35[1]),.doutc(w_n884_35[2]),.din(w_n884_11[1]));
	jspl3 jspl3_w_n884_36(.douta(w_n884_36[0]),.doutb(w_n884_36[1]),.doutc(w_n884_36[2]),.din(w_n884_11[2]));
	jspl3 jspl3_w_n884_37(.douta(w_n884_37[0]),.doutb(w_n884_37[1]),.doutc(w_n884_37[2]),.din(w_n884_12[0]));
	jspl3 jspl3_w_n884_38(.douta(w_n884_38[0]),.doutb(w_n884_38[1]),.doutc(w_n884_38[2]),.din(w_n884_12[1]));
	jspl3 jspl3_w_n884_39(.douta(w_n884_39[0]),.doutb(w_n884_39[1]),.doutc(w_n884_39[2]),.din(w_n884_12[2]));
	jspl3 jspl3_w_n884_40(.douta(w_n884_40[0]),.doutb(w_n884_40[1]),.doutc(w_n884_40[2]),.din(w_n884_13[0]));
	jspl3 jspl3_w_n884_41(.douta(w_n884_41[0]),.doutb(w_n884_41[1]),.doutc(w_n884_41[2]),.din(w_n884_13[1]));
	jspl3 jspl3_w_n884_42(.douta(w_n884_42[0]),.doutb(w_n884_42[1]),.doutc(w_n884_42[2]),.din(w_n884_13[2]));
	jspl3 jspl3_w_n884_43(.douta(w_n884_43[0]),.doutb(w_n884_43[1]),.doutc(w_n884_43[2]),.din(w_n884_14[0]));
	jspl3 jspl3_w_n884_44(.douta(w_n884_44[0]),.doutb(w_n884_44[1]),.doutc(w_n884_44[2]),.din(w_n884_14[1]));
	jspl3 jspl3_w_n884_45(.douta(w_n884_45[0]),.doutb(w_n884_45[1]),.doutc(w_n884_45[2]),.din(w_n884_14[2]));
	jspl3 jspl3_w_n884_46(.douta(w_n884_46[0]),.doutb(w_n884_46[1]),.doutc(w_n884_46[2]),.din(w_n884_15[0]));
	jspl3 jspl3_w_n884_47(.douta(w_n884_47[0]),.doutb(w_n884_47[1]),.doutc(w_n884_47[2]),.din(w_n884_15[1]));
	jspl3 jspl3_w_n884_48(.douta(w_n884_48[0]),.doutb(w_n884_48[1]),.doutc(w_n884_48[2]),.din(w_n884_15[2]));
	jspl3 jspl3_w_n884_49(.douta(w_n884_49[0]),.doutb(w_n884_49[1]),.doutc(w_n884_49[2]),.din(w_n884_16[0]));
	jspl3 jspl3_w_n884_50(.douta(w_n884_50[0]),.doutb(w_n884_50[1]),.doutc(w_n884_50[2]),.din(w_n884_16[1]));
	jspl3 jspl3_w_n884_51(.douta(w_n884_51[0]),.doutb(w_n884_51[1]),.doutc(w_n884_51[2]),.din(w_n884_16[2]));
	jspl3 jspl3_w_n884_52(.douta(w_n884_52[0]),.doutb(w_n884_52[1]),.doutc(w_n884_52[2]),.din(w_n884_17[0]));
	jspl3 jspl3_w_n884_53(.douta(w_n884_53[0]),.doutb(w_n884_53[1]),.doutc(w_n884_53[2]),.din(w_n884_17[1]));
	jspl3 jspl3_w_n884_54(.douta(w_n884_54[0]),.doutb(w_n884_54[1]),.doutc(w_n884_54[2]),.din(w_n884_17[2]));
	jspl3 jspl3_w_n884_55(.douta(w_n884_55[0]),.doutb(w_n884_55[1]),.doutc(w_n884_55[2]),.din(w_n884_18[0]));
	jspl3 jspl3_w_n884_56(.douta(w_n884_56[0]),.doutb(w_n884_56[1]),.doutc(w_n884_56[2]),.din(w_n884_18[1]));
	jspl3 jspl3_w_n884_57(.douta(w_n884_57[0]),.doutb(w_n884_57[1]),.doutc(w_n884_57[2]),.din(w_n884_18[2]));
	jspl3 jspl3_w_n884_58(.douta(w_n884_58[0]),.doutb(w_n884_58[1]),.doutc(w_n884_58[2]),.din(w_n884_19[0]));
	jspl3 jspl3_w_n884_59(.douta(w_n884_59[0]),.doutb(w_n884_59[1]),.doutc(w_n884_59[2]),.din(w_n884_19[1]));
	jspl3 jspl3_w_n884_60(.douta(w_n884_60[0]),.doutb(w_n884_60[1]),.doutc(w_n884_60[2]),.din(w_n884_19[2]));
	jspl3 jspl3_w_n884_61(.douta(w_n884_61[0]),.doutb(w_n884_61[1]),.doutc(w_n884_61[2]),.din(w_n884_20[0]));
	jspl3 jspl3_w_n884_62(.douta(w_n884_62[0]),.doutb(w_n884_62[1]),.doutc(w_n884_62[2]),.din(w_n884_20[1]));
	jspl3 jspl3_w_n884_63(.douta(w_n884_63[0]),.doutb(w_n884_63[1]),.doutc(w_n884_63[2]),.din(w_n884_20[2]));
	jspl3 jspl3_w_n884_64(.douta(w_n884_64[0]),.doutb(w_n884_64[1]),.doutc(w_n884_64[2]),.din(w_n884_21[0]));
	jspl3 jspl3_w_n884_65(.douta(w_n884_65[0]),.doutb(w_n884_65[1]),.doutc(w_n884_65[2]),.din(w_n884_21[1]));
	jspl3 jspl3_w_n884_66(.douta(w_n884_66[0]),.doutb(w_n884_66[1]),.doutc(w_n884_66[2]),.din(w_n884_21[2]));
	jspl3 jspl3_w_n884_67(.douta(w_n884_67[0]),.doutb(w_n884_67[1]),.doutc(w_n884_67[2]),.din(w_n884_22[0]));
	jspl jspl_w_n886_0(.douta(w_n886_0[0]),.doutb(w_n886_0[1]),.din(n886));
	jspl3 jspl3_w_n888_0(.douta(w_n888_0[0]),.doutb(w_n888_0[1]),.doutc(w_n888_0[2]),.din(n888));
	jspl jspl_w_n889_0(.douta(w_n889_0[0]),.doutb(w_n889_0[1]),.din(n889));
	jspl jspl_w_n891_0(.douta(w_n891_0[0]),.doutb(w_n891_0[1]),.din(n891));
	jspl jspl_w_n896_0(.douta(w_n896_0[0]),.doutb(w_n896_0[1]),.din(n896));
	jspl jspl_w_n897_0(.douta(w_n897_0[0]),.doutb(w_n897_0[1]),.din(n897));
	jspl3 jspl3_w_n899_0(.douta(w_n899_0[0]),.doutb(w_n899_0[1]),.doutc(w_n899_0[2]),.din(n899));
	jspl jspl_w_n900_0(.douta(w_n900_0[0]),.doutb(w_n900_0[1]),.din(n900));
	jspl jspl_w_n904_0(.douta(w_n904_0[0]),.doutb(w_n904_0[1]),.din(n904));
	jspl3 jspl3_w_n906_0(.douta(w_n906_0[0]),.doutb(w_n906_0[1]),.doutc(w_n906_0[2]),.din(n906));
	jspl jspl_w_n907_0(.douta(w_n907_0[0]),.doutb(w_n907_0[1]),.din(n907));
	jspl jspl_w_n911_0(.douta(w_n911_0[0]),.doutb(w_n911_0[1]),.din(n911));
	jspl3 jspl3_w_n913_0(.douta(w_n913_0[0]),.doutb(w_n913_0[1]),.doutc(w_n913_0[2]),.din(n913));
	jspl jspl_w_n914_0(.douta(w_n914_0[0]),.doutb(w_n914_0[1]),.din(n914));
	jspl jspl_w_n918_0(.douta(w_n918_0[0]),.doutb(w_n918_0[1]),.din(n918));
	jspl3 jspl3_w_n920_0(.douta(w_n920_0[0]),.doutb(w_n920_0[1]),.doutc(w_n920_0[2]),.din(n920));
	jspl jspl_w_n921_0(.douta(w_n921_0[0]),.doutb(w_n921_0[1]),.din(n921));
	jspl jspl_w_n925_0(.douta(w_n925_0[0]),.doutb(w_n925_0[1]),.din(n925));
	jspl jspl_w_n926_0(.douta(w_n926_0[0]),.doutb(w_n926_0[1]),.din(n926));
	jspl3 jspl3_w_n928_0(.douta(w_n928_0[0]),.doutb(w_n928_0[1]),.doutc(w_n928_0[2]),.din(n928));
	jspl jspl_w_n929_0(.douta(w_n929_0[0]),.doutb(w_n929_0[1]),.din(n929));
	jspl jspl_w_n933_0(.douta(w_n933_0[0]),.doutb(w_n933_0[1]),.din(n933));
	jspl3 jspl3_w_n935_0(.douta(w_n935_0[0]),.doutb(w_n935_0[1]),.doutc(w_n935_0[2]),.din(n935));
	jspl jspl_w_n936_0(.douta(w_n936_0[0]),.doutb(w_n936_0[1]),.din(n936));
	jspl jspl_w_n958_0(.douta(w_n958_0[0]),.doutb(w_n958_0[1]),.din(n958));
	jspl jspl_w_n962_0(.douta(w_n962_0[0]),.doutb(w_n962_0[1]),.din(n962));
	jspl jspl_w_n966_0(.douta(w_n966_0[0]),.doutb(w_n966_0[1]),.din(n966));
	jspl jspl_w_n973_0(.douta(w_n973_0[0]),.doutb(w_n973_0[1]),.din(n973));
	jspl jspl_w_n979_0(.douta(w_n979_0[0]),.doutb(w_n979_0[1]),.din(n979));
	jspl jspl_w_n981_0(.douta(w_n981_0[0]),.doutb(w_n981_0[1]),.din(n981));
	jspl jspl_w_n982_0(.douta(w_n982_0[0]),.doutb(w_n982_0[1]),.din(n982));
	jspl jspl_w_n985_0(.douta(w_n985_0[0]),.doutb(w_n985_0[1]),.din(n985));
	jspl jspl_w_n989_0(.douta(w_n989_0[0]),.doutb(w_n989_0[1]),.din(n989));
	jspl jspl_w_n991_0(.douta(w_n991_0[0]),.doutb(w_n991_0[1]),.din(n991));
	jspl3 jspl3_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.doutc(w_n992_0[2]),.din(n992));
	jspl jspl_w_n997_0(.douta(w_n997_0[0]),.doutb(w_n997_0[1]),.din(n997));
	jspl jspl_w_n1000_0(.douta(w_n1000_0[0]),.doutb(w_n1000_0[1]),.din(n1000));
	jspl jspl_w_n1004_0(.douta(w_n1004_0[0]),.doutb(w_n1004_0[1]),.din(n1004));
	jspl3 jspl3_w_n1008_0(.douta(w_n1008_0[0]),.doutb(w_n1008_0[1]),.doutc(w_n1008_0[2]),.din(n1008));
	jspl3 jspl3_w_n1008_1(.douta(w_n1008_1[0]),.doutb(w_n1008_1[1]),.doutc(w_n1008_1[2]),.din(w_n1008_0[0]));
	jspl3 jspl3_w_n1008_2(.douta(w_n1008_2[0]),.doutb(w_n1008_2[1]),.doutc(w_n1008_2[2]),.din(w_n1008_0[1]));
	jspl3 jspl3_w_n1008_3(.douta(w_n1008_3[0]),.doutb(w_n1008_3[1]),.doutc(w_n1008_3[2]),.din(w_n1008_0[2]));
	jspl3 jspl3_w_n1008_4(.douta(w_n1008_4[0]),.doutb(w_n1008_4[1]),.doutc(w_n1008_4[2]),.din(w_n1008_1[0]));
	jspl3 jspl3_w_n1008_5(.douta(w_n1008_5[0]),.doutb(w_n1008_5[1]),.doutc(w_n1008_5[2]),.din(w_n1008_1[1]));
	jspl3 jspl3_w_n1008_6(.douta(w_n1008_6[0]),.doutb(w_n1008_6[1]),.doutc(w_n1008_6[2]),.din(w_n1008_1[2]));
	jspl3 jspl3_w_n1008_7(.douta(w_n1008_7[0]),.doutb(w_n1008_7[1]),.doutc(w_n1008_7[2]),.din(w_n1008_2[0]));
	jspl3 jspl3_w_n1008_8(.douta(w_n1008_8[0]),.doutb(w_n1008_8[1]),.doutc(w_n1008_8[2]),.din(w_n1008_2[1]));
	jspl3 jspl3_w_n1008_9(.douta(w_n1008_9[0]),.doutb(w_n1008_9[1]),.doutc(w_n1008_9[2]),.din(w_n1008_2[2]));
	jspl3 jspl3_w_n1008_10(.douta(w_n1008_10[0]),.doutb(w_n1008_10[1]),.doutc(w_n1008_10[2]),.din(w_n1008_3[0]));
	jspl3 jspl3_w_n1008_11(.douta(w_n1008_11[0]),.doutb(w_n1008_11[1]),.doutc(w_n1008_11[2]),.din(w_n1008_3[1]));
	jspl3 jspl3_w_n1008_12(.douta(w_n1008_12[0]),.doutb(w_n1008_12[1]),.doutc(w_n1008_12[2]),.din(w_n1008_3[2]));
	jspl3 jspl3_w_n1008_13(.douta(w_n1008_13[0]),.doutb(w_n1008_13[1]),.doutc(w_n1008_13[2]),.din(w_n1008_4[0]));
	jspl3 jspl3_w_n1008_14(.douta(w_n1008_14[0]),.doutb(w_n1008_14[1]),.doutc(w_n1008_14[2]),.din(w_n1008_4[1]));
	jspl3 jspl3_w_n1008_15(.douta(w_n1008_15[0]),.doutb(w_n1008_15[1]),.doutc(w_n1008_15[2]),.din(w_n1008_4[2]));
	jspl3 jspl3_w_n1008_16(.douta(w_n1008_16[0]),.doutb(w_n1008_16[1]),.doutc(w_n1008_16[2]),.din(w_n1008_5[0]));
	jspl3 jspl3_w_n1008_17(.douta(w_n1008_17[0]),.doutb(w_n1008_17[1]),.doutc(w_n1008_17[2]),.din(w_n1008_5[1]));
	jspl3 jspl3_w_n1008_18(.douta(w_n1008_18[0]),.doutb(w_n1008_18[1]),.doutc(w_n1008_18[2]),.din(w_n1008_5[2]));
	jspl3 jspl3_w_n1008_19(.douta(w_n1008_19[0]),.doutb(w_n1008_19[1]),.doutc(w_n1008_19[2]),.din(w_n1008_6[0]));
	jspl3 jspl3_w_n1008_20(.douta(w_n1008_20[0]),.doutb(w_n1008_20[1]),.doutc(w_n1008_20[2]),.din(w_n1008_6[1]));
	jspl3 jspl3_w_n1008_21(.douta(w_n1008_21[0]),.doutb(w_n1008_21[1]),.doutc(w_n1008_21[2]),.din(w_n1008_6[2]));
	jspl3 jspl3_w_n1008_22(.douta(w_n1008_22[0]),.doutb(w_n1008_22[1]),.doutc(w_n1008_22[2]),.din(w_n1008_7[0]));
	jspl3 jspl3_w_n1008_23(.douta(w_n1008_23[0]),.doutb(w_n1008_23[1]),.doutc(w_n1008_23[2]),.din(w_n1008_7[1]));
	jspl3 jspl3_w_n1008_24(.douta(w_n1008_24[0]),.doutb(w_n1008_24[1]),.doutc(w_n1008_24[2]),.din(w_n1008_7[2]));
	jspl3 jspl3_w_n1008_25(.douta(w_n1008_25[0]),.doutb(w_n1008_25[1]),.doutc(w_n1008_25[2]),.din(w_n1008_8[0]));
	jspl3 jspl3_w_n1008_26(.douta(w_n1008_26[0]),.doutb(w_n1008_26[1]),.doutc(w_n1008_26[2]),.din(w_n1008_8[1]));
	jspl3 jspl3_w_n1008_27(.douta(w_n1008_27[0]),.doutb(w_n1008_27[1]),.doutc(w_n1008_27[2]),.din(w_n1008_8[2]));
	jspl3 jspl3_w_n1008_28(.douta(w_n1008_28[0]),.doutb(w_n1008_28[1]),.doutc(w_n1008_28[2]),.din(w_n1008_9[0]));
	jspl3 jspl3_w_n1008_29(.douta(w_n1008_29[0]),.doutb(w_n1008_29[1]),.doutc(w_n1008_29[2]),.din(w_n1008_9[1]));
	jspl3 jspl3_w_n1008_30(.douta(w_n1008_30[0]),.doutb(w_n1008_30[1]),.doutc(w_n1008_30[2]),.din(w_n1008_9[2]));
	jspl3 jspl3_w_n1008_31(.douta(w_n1008_31[0]),.doutb(w_n1008_31[1]),.doutc(w_n1008_31[2]),.din(w_n1008_10[0]));
	jspl3 jspl3_w_n1008_32(.douta(w_n1008_32[0]),.doutb(w_n1008_32[1]),.doutc(w_n1008_32[2]),.din(w_n1008_10[1]));
	jspl3 jspl3_w_n1008_33(.douta(w_n1008_33[0]),.doutb(w_n1008_33[1]),.doutc(w_n1008_33[2]),.din(w_n1008_10[2]));
	jspl3 jspl3_w_n1008_34(.douta(w_n1008_34[0]),.doutb(w_n1008_34[1]),.doutc(w_n1008_34[2]),.din(w_n1008_11[0]));
	jspl3 jspl3_w_n1008_35(.douta(w_n1008_35[0]),.doutb(w_n1008_35[1]),.doutc(w_n1008_35[2]),.din(w_n1008_11[1]));
	jspl3 jspl3_w_n1008_36(.douta(w_n1008_36[0]),.doutb(w_n1008_36[1]),.doutc(w_n1008_36[2]),.din(w_n1008_11[2]));
	jspl3 jspl3_w_n1008_37(.douta(w_n1008_37[0]),.doutb(w_n1008_37[1]),.doutc(w_n1008_37[2]),.din(w_n1008_12[0]));
	jspl3 jspl3_w_n1008_38(.douta(w_n1008_38[0]),.doutb(w_n1008_38[1]),.doutc(w_n1008_38[2]),.din(w_n1008_12[1]));
	jspl3 jspl3_w_n1008_39(.douta(w_n1008_39[0]),.doutb(w_n1008_39[1]),.doutc(w_n1008_39[2]),.din(w_n1008_12[2]));
	jspl3 jspl3_w_n1008_40(.douta(w_n1008_40[0]),.doutb(w_n1008_40[1]),.doutc(w_n1008_40[2]),.din(w_n1008_13[0]));
	jspl3 jspl3_w_n1008_41(.douta(w_n1008_41[0]),.doutb(w_n1008_41[1]),.doutc(w_n1008_41[2]),.din(w_n1008_13[1]));
	jspl3 jspl3_w_n1008_42(.douta(w_n1008_42[0]),.doutb(w_n1008_42[1]),.doutc(w_n1008_42[2]),.din(w_n1008_13[2]));
	jspl3 jspl3_w_n1008_43(.douta(w_n1008_43[0]),.doutb(w_n1008_43[1]),.doutc(w_n1008_43[2]),.din(w_n1008_14[0]));
	jspl3 jspl3_w_n1008_44(.douta(w_n1008_44[0]),.doutb(w_n1008_44[1]),.doutc(w_n1008_44[2]),.din(w_n1008_14[1]));
	jspl3 jspl3_w_n1008_45(.douta(w_n1008_45[0]),.doutb(w_n1008_45[1]),.doutc(w_n1008_45[2]),.din(w_n1008_14[2]));
	jspl3 jspl3_w_n1008_46(.douta(w_n1008_46[0]),.doutb(w_n1008_46[1]),.doutc(w_n1008_46[2]),.din(w_n1008_15[0]));
	jspl3 jspl3_w_n1008_47(.douta(w_n1008_47[0]),.doutb(w_n1008_47[1]),.doutc(w_n1008_47[2]),.din(w_n1008_15[1]));
	jspl3 jspl3_w_n1008_48(.douta(w_n1008_48[0]),.doutb(w_n1008_48[1]),.doutc(w_n1008_48[2]),.din(w_n1008_15[2]));
	jspl3 jspl3_w_n1008_49(.douta(w_n1008_49[0]),.doutb(w_n1008_49[1]),.doutc(w_n1008_49[2]),.din(w_n1008_16[0]));
	jspl3 jspl3_w_n1008_50(.douta(w_n1008_50[0]),.doutb(w_n1008_50[1]),.doutc(w_n1008_50[2]),.din(w_n1008_16[1]));
	jspl3 jspl3_w_n1008_51(.douta(w_n1008_51[0]),.doutb(w_n1008_51[1]),.doutc(w_n1008_51[2]),.din(w_n1008_16[2]));
	jspl3 jspl3_w_n1008_52(.douta(w_n1008_52[0]),.doutb(w_n1008_52[1]),.doutc(w_n1008_52[2]),.din(w_n1008_17[0]));
	jspl3 jspl3_w_n1008_53(.douta(w_n1008_53[0]),.doutb(w_n1008_53[1]),.doutc(w_n1008_53[2]),.din(w_n1008_17[1]));
	jspl3 jspl3_w_n1008_54(.douta(w_n1008_54[0]),.doutb(w_n1008_54[1]),.doutc(w_n1008_54[2]),.din(w_n1008_17[2]));
	jspl3 jspl3_w_n1008_55(.douta(w_n1008_55[0]),.doutb(w_n1008_55[1]),.doutc(w_n1008_55[2]),.din(w_n1008_18[0]));
	jspl3 jspl3_w_n1008_56(.douta(w_n1008_56[0]),.doutb(w_n1008_56[1]),.doutc(w_n1008_56[2]),.din(w_n1008_18[1]));
	jspl3 jspl3_w_n1008_57(.douta(w_n1008_57[0]),.doutb(w_n1008_57[1]),.doutc(w_n1008_57[2]),.din(w_n1008_18[2]));
	jspl3 jspl3_w_n1008_58(.douta(w_n1008_58[0]),.doutb(w_n1008_58[1]),.doutc(w_n1008_58[2]),.din(w_n1008_19[0]));
	jspl3 jspl3_w_n1008_59(.douta(w_n1008_59[0]),.doutb(w_n1008_59[1]),.doutc(w_n1008_59[2]),.din(w_n1008_19[1]));
	jspl3 jspl3_w_n1008_60(.douta(w_n1008_60[0]),.doutb(w_n1008_60[1]),.doutc(w_n1008_60[2]),.din(w_n1008_19[2]));
	jspl3 jspl3_w_n1008_61(.douta(w_n1008_61[0]),.doutb(w_n1008_61[1]),.doutc(w_n1008_61[2]),.din(w_n1008_20[0]));
	jspl3 jspl3_w_n1008_62(.douta(w_n1008_62[0]),.doutb(w_n1008_62[1]),.doutc(w_n1008_62[2]),.din(w_n1008_20[1]));
	jspl3 jspl3_w_n1008_63(.douta(w_n1008_63[0]),.doutb(w_n1008_63[1]),.doutc(w_n1008_63[2]),.din(w_n1008_20[2]));
	jspl3 jspl3_w_n1008_64(.douta(w_n1008_64[0]),.doutb(w_n1008_64[1]),.doutc(w_n1008_64[2]),.din(w_n1008_21[0]));
	jspl3 jspl3_w_n1008_65(.douta(w_n1008_65[0]),.doutb(w_n1008_65[1]),.doutc(w_n1008_65[2]),.din(w_n1008_21[1]));
	jspl3 jspl3_w_n1008_66(.douta(w_n1008_66[0]),.doutb(w_n1008_66[1]),.doutc(w_n1008_66[2]),.din(w_n1008_21[2]));
	jspl3 jspl3_w_n1008_67(.douta(w_n1008_67[0]),.doutb(w_n1008_67[1]),.doutc(w_n1008_67[2]),.din(w_n1008_22[0]));
	jspl3 jspl3_w_n1008_68(.douta(w_n1008_68[0]),.doutb(w_n1008_68[1]),.doutc(w_n1008_68[2]),.din(w_n1008_22[1]));
	jspl3 jspl3_w_n1008_69(.douta(w_n1008_69[0]),.doutb(w_n1008_69[1]),.doutc(w_n1008_69[2]),.din(w_n1008_22[2]));
	jspl jspl_w_n1008_70(.douta(w_n1008_70[0]),.doutb(w_n1008_70[1]),.din(w_n1008_23[0]));
	jspl3 jspl3_w_n1010_0(.douta(w_n1010_0[0]),.doutb(w_n1010_0[1]),.doutc(w_n1010_0[2]),.din(n1010));
	jspl3 jspl3_w_n1010_1(.douta(w_n1010_1[0]),.doutb(w_n1010_1[1]),.doutc(w_n1010_1[2]),.din(w_n1010_0[0]));
	jspl jspl_w_n1011_0(.douta(w_n1011_0[0]),.doutb(w_n1011_0[1]),.din(n1011));
	jspl3 jspl3_w_n1012_0(.douta(w_n1012_0[0]),.doutb(w_n1012_0[1]),.doutc(w_n1012_0[2]),.din(n1012));
	jspl jspl_w_n1013_0(.douta(w_n1013_0[0]),.doutb(w_n1013_0[1]),.din(n1013));
	jspl3 jspl3_w_n1015_0(.douta(w_n1015_0[0]),.doutb(w_n1015_0[1]),.doutc(w_n1015_0[2]),.din(n1015));
	jspl jspl_w_n1016_0(.douta(w_n1016_0[0]),.doutb(w_n1016_0[1]),.din(n1016));
	jspl3 jspl3_w_n1023_0(.douta(w_n1023_0[0]),.doutb(w_n1023_0[1]),.doutc(w_n1023_0[2]),.din(n1023));
	jspl jspl_w_n1024_0(.douta(w_n1024_0[0]),.doutb(w_n1024_0[1]),.din(n1024));
	jspl jspl_w_n1027_0(.douta(w_n1027_0[0]),.doutb(w_n1027_0[1]),.din(n1027));
	jspl jspl_w_n1028_0(.douta(w_n1028_0[0]),.doutb(w_n1028_0[1]),.din(n1028));
	jspl3 jspl3_w_n1033_0(.douta(w_n1033_0[0]),.doutb(w_n1033_0[1]),.doutc(w_n1033_0[2]),.din(n1033));
	jspl3 jspl3_w_n1035_0(.douta(w_n1035_0[0]),.doutb(w_n1035_0[1]),.doutc(w_n1035_0[2]),.din(n1035));
	jspl jspl_w_n1036_0(.douta(w_n1036_0[0]),.doutb(w_n1036_0[1]),.din(n1036));
	jspl3 jspl3_w_n1040_0(.douta(w_n1040_0[0]),.doutb(w_n1040_0[1]),.doutc(w_n1040_0[2]),.din(n1040));
	jspl3 jspl3_w_n1042_0(.douta(w_n1042_0[0]),.doutb(w_n1042_0[1]),.doutc(w_n1042_0[2]),.din(n1042));
	jspl jspl_w_n1043_0(.douta(w_n1043_0[0]),.doutb(w_n1043_0[1]),.din(n1043));
	jspl3 jspl3_w_n1047_0(.douta(w_n1047_0[0]),.doutb(w_n1047_0[1]),.doutc(w_n1047_0[2]),.din(n1047));
	jspl3 jspl3_w_n1049_0(.douta(w_n1049_0[0]),.doutb(w_n1049_0[1]),.doutc(w_n1049_0[2]),.din(n1049));
	jspl jspl_w_n1050_0(.douta(w_n1050_0[0]),.doutb(w_n1050_0[1]),.din(n1050));
	jspl3 jspl3_w_n1054_0(.douta(w_n1054_0[0]),.doutb(w_n1054_0[1]),.doutc(w_n1054_0[2]),.din(n1054));
	jspl3 jspl3_w_n1057_0(.douta(w_n1057_0[0]),.doutb(w_n1057_0[1]),.doutc(w_n1057_0[2]),.din(n1057));
	jspl jspl_w_n1058_0(.douta(w_n1058_0[0]),.doutb(w_n1058_0[1]),.din(n1058));
	jspl3 jspl3_w_n1062_0(.douta(w_n1062_0[0]),.doutb(w_n1062_0[1]),.doutc(w_n1062_0[2]),.din(n1062));
	jspl3 jspl3_w_n1065_0(.douta(w_n1065_0[0]),.doutb(w_n1065_0[1]),.doutc(w_n1065_0[2]),.din(n1065));
	jspl jspl_w_n1066_0(.douta(w_n1066_0[0]),.doutb(w_n1066_0[1]),.din(n1066));
	jspl3 jspl3_w_n1070_0(.douta(w_n1070_0[0]),.doutb(w_n1070_0[1]),.doutc(w_n1070_0[2]),.din(n1070));
	jspl3 jspl3_w_n1073_0(.douta(w_n1073_0[0]),.doutb(w_n1073_0[1]),.doutc(w_n1073_0[2]),.din(n1073));
	jspl jspl_w_n1074_0(.douta(w_n1074_0[0]),.doutb(w_n1074_0[1]),.din(n1074));
	jspl3 jspl3_w_n1078_0(.douta(w_n1078_0[0]),.doutb(w_n1078_0[1]),.doutc(w_n1078_0[2]),.din(n1078));
	jspl3 jspl3_w_n1080_0(.douta(w_n1080_0[0]),.doutb(w_n1080_0[1]),.doutc(w_n1080_0[2]),.din(n1080));
	jspl jspl_w_n1081_0(.douta(w_n1081_0[0]),.doutb(w_n1081_0[1]),.din(n1081));
	jspl jspl_w_n1085_0(.douta(w_n1085_0[0]),.doutb(w_n1085_0[1]),.din(n1085));
	jspl jspl_w_n1086_0(.douta(w_n1086_0[0]),.doutb(w_n1086_0[1]),.din(n1086));
	jspl3 jspl3_w_n1088_0(.douta(w_n1088_0[0]),.doutb(w_n1088_0[1]),.doutc(w_n1088_0[2]),.din(n1088));
	jspl jspl_w_n1088_1(.douta(w_n1088_1[0]),.doutb(w_n1088_1[1]),.din(w_n1088_0[0]));
	jspl3 jspl3_w_n1091_0(.douta(w_n1091_0[0]),.doutb(w_n1091_0[1]),.doutc(w_n1091_0[2]),.din(n1091));
	jspl jspl_w_n1091_1(.douta(w_n1091_1[0]),.doutb(w_n1091_1[1]),.din(w_n1091_0[0]));
	jspl jspl_w_n1092_0(.douta(w_n1092_0[0]),.doutb(w_n1092_0[1]),.din(n1092));
	jspl jspl_w_n1096_0(.douta(w_n1096_0[0]),.doutb(w_n1096_0[1]),.din(n1096));
	jspl jspl_w_n1097_0(.douta(w_n1097_0[0]),.doutb(w_n1097_0[1]),.din(n1097));
	jspl jspl_w_n1101_0(.douta(w_n1101_0[0]),.doutb(w_n1101_0[1]),.din(n1101));
	jspl jspl_w_n1104_0(.douta(w_n1104_0[0]),.doutb(w_n1104_0[1]),.din(n1104));
	jspl3 jspl3_w_n1108_0(.douta(w_n1108_0[0]),.doutb(w_n1108_0[1]),.doutc(w_n1108_0[2]),.din(n1108));
	jspl jspl_w_n1108_1(.douta(w_n1108_1[0]),.doutb(w_n1108_1[1]),.din(w_n1108_0[0]));
	jspl jspl_w_n1109_0(.douta(w_n1109_0[0]),.doutb(w_n1109_0[1]),.din(n1109));
	jspl3 jspl3_w_n1110_0(.douta(w_n1110_0[0]),.doutb(w_n1110_0[1]),.doutc(w_n1110_0[2]),.din(n1110));
	jspl jspl_w_n1111_0(.douta(w_n1111_0[0]),.doutb(w_n1111_0[1]),.din(n1111));
	jspl3 jspl3_w_n1113_0(.douta(w_n1113_0[0]),.doutb(w_n1113_0[1]),.doutc(w_n1113_0[2]),.din(n1113));
	jspl jspl_w_n1114_0(.douta(w_n1114_0[0]),.doutb(w_n1114_0[1]),.din(n1114));
	jspl jspl_w_n1119_0(.douta(w_n1119_0[0]),.doutb(w_n1119_0[1]),.din(n1119));
	jspl jspl_w_n1134_0(.douta(w_n1134_0[0]),.doutb(w_n1134_0[1]),.din(n1134));
	jspl jspl_w_n1169_0(.douta(w_n1169_0[0]),.doutb(w_n1169_0[1]),.din(n1169));
	jspl jspl_w_n1172_0(.douta(w_n1172_0[0]),.doutb(w_n1172_0[1]),.din(n1172));
	jspl3 jspl3_w_n1173_0(.douta(w_n1173_0[0]),.doutb(w_n1173_0[1]),.doutc(w_n1173_0[2]),.din(n1173));
	jspl3 jspl3_w_n1173_1(.douta(w_n1173_1[0]),.doutb(w_n1173_1[1]),.doutc(w_n1173_1[2]),.din(w_n1173_0[0]));
	jspl3 jspl3_w_n1173_2(.douta(w_n1173_2[0]),.doutb(w_n1173_2[1]),.doutc(w_n1173_2[2]),.din(w_n1173_0[1]));
	jspl3 jspl3_w_n1173_3(.douta(w_n1173_3[0]),.doutb(w_n1173_3[1]),.doutc(w_n1173_3[2]),.din(w_n1173_0[2]));
	jspl3 jspl3_w_n1173_4(.douta(w_n1173_4[0]),.doutb(w_n1173_4[1]),.doutc(w_n1173_4[2]),.din(w_n1173_1[0]));
	jspl3 jspl3_w_n1173_5(.douta(w_n1173_5[0]),.doutb(w_n1173_5[1]),.doutc(w_n1173_5[2]),.din(w_n1173_1[1]));
	jspl3 jspl3_w_n1173_6(.douta(w_n1173_6[0]),.doutb(w_n1173_6[1]),.doutc(w_n1173_6[2]),.din(w_n1173_1[2]));
	jspl3 jspl3_w_n1173_7(.douta(w_n1173_7[0]),.doutb(w_n1173_7[1]),.doutc(w_n1173_7[2]),.din(w_n1173_2[0]));
	jspl3 jspl3_w_n1173_8(.douta(w_n1173_8[0]),.doutb(w_n1173_8[1]),.doutc(w_n1173_8[2]),.din(w_n1173_2[1]));
	jspl3 jspl3_w_n1173_9(.douta(w_n1173_9[0]),.doutb(w_n1173_9[1]),.doutc(w_n1173_9[2]),.din(w_n1173_2[2]));
	jspl3 jspl3_w_n1173_10(.douta(w_n1173_10[0]),.doutb(w_n1173_10[1]),.doutc(w_n1173_10[2]),.din(w_n1173_3[0]));
	jspl3 jspl3_w_n1173_11(.douta(w_n1173_11[0]),.doutb(w_n1173_11[1]),.doutc(w_n1173_11[2]),.din(w_n1173_3[1]));
	jspl3 jspl3_w_n1173_12(.douta(w_n1173_12[0]),.doutb(w_n1173_12[1]),.doutc(w_n1173_12[2]),.din(w_n1173_3[2]));
	jspl3 jspl3_w_n1173_13(.douta(w_n1173_13[0]),.doutb(w_n1173_13[1]),.doutc(w_n1173_13[2]),.din(w_n1173_4[0]));
	jspl3 jspl3_w_n1173_14(.douta(w_n1173_14[0]),.doutb(w_n1173_14[1]),.doutc(w_n1173_14[2]),.din(w_n1173_4[1]));
	jspl3 jspl3_w_n1173_15(.douta(w_n1173_15[0]),.doutb(w_n1173_15[1]),.doutc(w_n1173_15[2]),.din(w_n1173_4[2]));
	jspl3 jspl3_w_n1173_16(.douta(w_n1173_16[0]),.doutb(w_n1173_16[1]),.doutc(w_n1173_16[2]),.din(w_n1173_5[0]));
	jspl3 jspl3_w_n1173_17(.douta(w_n1173_17[0]),.doutb(w_n1173_17[1]),.doutc(w_n1173_17[2]),.din(w_n1173_5[1]));
	jspl3 jspl3_w_n1173_18(.douta(w_n1173_18[0]),.doutb(w_n1173_18[1]),.doutc(w_n1173_18[2]),.din(w_n1173_5[2]));
	jspl3 jspl3_w_n1173_19(.douta(w_n1173_19[0]),.doutb(w_n1173_19[1]),.doutc(w_n1173_19[2]),.din(w_n1173_6[0]));
	jspl3 jspl3_w_n1173_20(.douta(w_n1173_20[0]),.doutb(w_n1173_20[1]),.doutc(w_n1173_20[2]),.din(w_n1173_6[1]));
	jspl3 jspl3_w_n1173_21(.douta(w_n1173_21[0]),.doutb(w_n1173_21[1]),.doutc(w_n1173_21[2]),.din(w_n1173_6[2]));
	jspl3 jspl3_w_n1173_22(.douta(w_n1173_22[0]),.doutb(w_n1173_22[1]),.doutc(w_n1173_22[2]),.din(w_n1173_7[0]));
	jspl3 jspl3_w_n1173_23(.douta(w_n1173_23[0]),.doutb(w_n1173_23[1]),.doutc(w_n1173_23[2]),.din(w_n1173_7[1]));
	jspl3 jspl3_w_n1173_24(.douta(w_n1173_24[0]),.doutb(w_n1173_24[1]),.doutc(w_n1173_24[2]),.din(w_n1173_7[2]));
	jspl3 jspl3_w_n1173_25(.douta(w_n1173_25[0]),.doutb(w_n1173_25[1]),.doutc(w_n1173_25[2]),.din(w_n1173_8[0]));
	jspl3 jspl3_w_n1173_26(.douta(w_n1173_26[0]),.doutb(w_n1173_26[1]),.doutc(w_n1173_26[2]),.din(w_n1173_8[1]));
	jspl3 jspl3_w_n1173_27(.douta(w_n1173_27[0]),.doutb(w_n1173_27[1]),.doutc(w_n1173_27[2]),.din(w_n1173_8[2]));
	jspl3 jspl3_w_n1173_28(.douta(w_n1173_28[0]),.doutb(w_n1173_28[1]),.doutc(w_n1173_28[2]),.din(w_n1173_9[0]));
	jspl3 jspl3_w_n1173_29(.douta(w_n1173_29[0]),.doutb(w_n1173_29[1]),.doutc(w_n1173_29[2]),.din(w_n1173_9[1]));
	jspl3 jspl3_w_n1173_30(.douta(w_n1173_30[0]),.doutb(w_n1173_30[1]),.doutc(w_n1173_30[2]),.din(w_n1173_9[2]));
	jspl3 jspl3_w_n1173_31(.douta(w_n1173_31[0]),.doutb(w_n1173_31[1]),.doutc(w_n1173_31[2]),.din(w_n1173_10[0]));
	jspl3 jspl3_w_n1173_32(.douta(w_n1173_32[0]),.doutb(w_n1173_32[1]),.doutc(w_n1173_32[2]),.din(w_n1173_10[1]));
	jspl3 jspl3_w_n1173_33(.douta(w_n1173_33[0]),.doutb(w_n1173_33[1]),.doutc(w_n1173_33[2]),.din(w_n1173_10[2]));
	jspl3 jspl3_w_n1173_34(.douta(w_n1173_34[0]),.doutb(w_n1173_34[1]),.doutc(w_n1173_34[2]),.din(w_n1173_11[0]));
	jspl3 jspl3_w_n1173_35(.douta(w_n1173_35[0]),.doutb(w_n1173_35[1]),.doutc(w_n1173_35[2]),.din(w_n1173_11[1]));
	jspl3 jspl3_w_n1173_36(.douta(w_n1173_36[0]),.doutb(w_n1173_36[1]),.doutc(w_n1173_36[2]),.din(w_n1173_11[2]));
	jspl3 jspl3_w_n1173_37(.douta(w_n1173_37[0]),.doutb(w_n1173_37[1]),.doutc(w_n1173_37[2]),.din(w_n1173_12[0]));
	jspl3 jspl3_w_n1173_38(.douta(w_n1173_38[0]),.doutb(w_n1173_38[1]),.doutc(w_n1173_38[2]),.din(w_n1173_12[1]));
	jspl3 jspl3_w_n1173_39(.douta(w_n1173_39[0]),.doutb(w_n1173_39[1]),.doutc(w_n1173_39[2]),.din(w_n1173_12[2]));
	jspl3 jspl3_w_n1173_40(.douta(w_n1173_40[0]),.doutb(w_n1173_40[1]),.doutc(w_n1173_40[2]),.din(w_n1173_13[0]));
	jspl3 jspl3_w_n1173_41(.douta(w_n1173_41[0]),.doutb(w_n1173_41[1]),.doutc(w_n1173_41[2]),.din(w_n1173_13[1]));
	jspl3 jspl3_w_n1173_42(.douta(w_n1173_42[0]),.doutb(w_n1173_42[1]),.doutc(w_n1173_42[2]),.din(w_n1173_13[2]));
	jspl3 jspl3_w_n1173_43(.douta(w_n1173_43[0]),.doutb(w_n1173_43[1]),.doutc(w_n1173_43[2]),.din(w_n1173_14[0]));
	jspl3 jspl3_w_n1173_44(.douta(w_n1173_44[0]),.doutb(w_n1173_44[1]),.doutc(w_n1173_44[2]),.din(w_n1173_14[1]));
	jspl3 jspl3_w_n1173_45(.douta(w_n1173_45[0]),.doutb(w_n1173_45[1]),.doutc(w_n1173_45[2]),.din(w_n1173_14[2]));
	jspl3 jspl3_w_n1173_46(.douta(w_n1173_46[0]),.doutb(w_n1173_46[1]),.doutc(w_n1173_46[2]),.din(w_n1173_15[0]));
	jspl3 jspl3_w_n1173_47(.douta(w_n1173_47[0]),.doutb(w_n1173_47[1]),.doutc(w_n1173_47[2]),.din(w_n1173_15[1]));
	jspl3 jspl3_w_n1173_48(.douta(w_n1173_48[0]),.doutb(w_n1173_48[1]),.doutc(w_n1173_48[2]),.din(w_n1173_15[2]));
	jspl3 jspl3_w_n1173_49(.douta(w_n1173_49[0]),.doutb(w_n1173_49[1]),.doutc(w_n1173_49[2]),.din(w_n1173_16[0]));
	jspl3 jspl3_w_n1173_50(.douta(w_n1173_50[0]),.doutb(w_n1173_50[1]),.doutc(w_n1173_50[2]),.din(w_n1173_16[1]));
	jspl3 jspl3_w_n1173_51(.douta(w_n1173_51[0]),.doutb(w_n1173_51[1]),.doutc(w_n1173_51[2]),.din(w_n1173_16[2]));
	jspl3 jspl3_w_n1173_52(.douta(w_n1173_52[0]),.doutb(w_n1173_52[1]),.doutc(w_n1173_52[2]),.din(w_n1173_17[0]));
	jspl3 jspl3_w_n1173_53(.douta(w_n1173_53[0]),.doutb(w_n1173_53[1]),.doutc(w_n1173_53[2]),.din(w_n1173_17[1]));
	jspl3 jspl3_w_n1173_54(.douta(w_n1173_54[0]),.doutb(w_n1173_54[1]),.doutc(w_n1173_54[2]),.din(w_n1173_17[2]));
	jspl3 jspl3_w_n1173_55(.douta(w_n1173_55[0]),.doutb(w_n1173_55[1]),.doutc(w_n1173_55[2]),.din(w_n1173_18[0]));
	jspl3 jspl3_w_n1173_56(.douta(w_n1173_56[0]),.doutb(w_n1173_56[1]),.doutc(w_n1173_56[2]),.din(w_n1173_18[1]));
	jspl3 jspl3_w_n1173_57(.douta(w_n1173_57[0]),.doutb(w_n1173_57[1]),.doutc(w_n1173_57[2]),.din(w_n1173_18[2]));
	jspl3 jspl3_w_n1173_58(.douta(w_n1173_58[0]),.doutb(w_n1173_58[1]),.doutc(w_n1173_58[2]),.din(w_n1173_19[0]));
	jspl3 jspl3_w_n1173_59(.douta(w_n1173_59[0]),.doutb(w_n1173_59[1]),.doutc(w_n1173_59[2]),.din(w_n1173_19[1]));
	jspl3 jspl3_w_n1173_60(.douta(w_n1173_60[0]),.doutb(w_n1173_60[1]),.doutc(w_n1173_60[2]),.din(w_n1173_19[2]));
	jspl3 jspl3_w_n1173_61(.douta(w_n1173_61[0]),.doutb(w_n1173_61[1]),.doutc(w_n1173_61[2]),.din(w_n1173_20[0]));
	jspl3 jspl3_w_n1173_62(.douta(w_n1173_62[0]),.doutb(w_n1173_62[1]),.doutc(w_n1173_62[2]),.din(w_n1173_20[1]));
	jspl3 jspl3_w_n1173_63(.douta(w_n1173_63[0]),.doutb(w_n1173_63[1]),.doutc(w_n1173_63[2]),.din(w_n1173_20[2]));
	jspl3 jspl3_w_n1173_64(.douta(w_n1173_64[0]),.doutb(w_n1173_64[1]),.doutc(w_n1173_64[2]),.din(w_n1173_21[0]));
	jspl jspl_w_n1175_0(.douta(w_n1175_0[0]),.doutb(w_n1175_0[1]),.din(n1175));
	jspl3 jspl3_w_n1177_0(.douta(w_n1177_0[0]),.doutb(w_n1177_0[1]),.doutc(w_n1177_0[2]),.din(n1177));
	jspl jspl_w_n1178_0(.douta(w_n1178_0[0]),.doutb(w_n1178_0[1]),.din(n1178));
	jspl jspl_w_n1180_0(.douta(w_n1180_0[0]),.doutb(w_n1180_0[1]),.din(n1180));
	jspl jspl_w_n1185_0(.douta(w_n1185_0[0]),.doutb(w_n1185_0[1]),.din(n1185));
	jspl jspl_w_n1186_0(.douta(w_n1186_0[0]),.doutb(w_n1186_0[1]),.din(n1186));
	jspl3 jspl3_w_n1188_0(.douta(w_n1188_0[0]),.doutb(w_n1188_0[1]),.doutc(w_n1188_0[2]),.din(n1188));
	jspl jspl_w_n1189_0(.douta(w_n1189_0[0]),.doutb(w_n1189_0[1]),.din(n1189));
	jspl jspl_w_n1193_0(.douta(w_n1193_0[0]),.doutb(w_n1193_0[1]),.din(n1193));
	jspl3 jspl3_w_n1195_0(.douta(w_n1195_0[0]),.doutb(w_n1195_0[1]),.doutc(w_n1195_0[2]),.din(n1195));
	jspl jspl_w_n1196_0(.douta(w_n1196_0[0]),.doutb(w_n1196_0[1]),.din(n1196));
	jspl jspl_w_n1200_0(.douta(w_n1200_0[0]),.doutb(w_n1200_0[1]),.din(n1200));
	jspl jspl_w_n1201_0(.douta(w_n1201_0[0]),.doutb(w_n1201_0[1]),.din(n1201));
	jspl3 jspl3_w_n1203_0(.douta(w_n1203_0[0]),.doutb(w_n1203_0[1]),.doutc(w_n1203_0[2]),.din(n1203));
	jspl jspl_w_n1204_0(.douta(w_n1204_0[0]),.doutb(w_n1204_0[1]),.din(n1204));
	jspl jspl_w_n1208_0(.douta(w_n1208_0[0]),.doutb(w_n1208_0[1]),.din(n1208));
	jspl jspl_w_n1209_0(.douta(w_n1209_0[0]),.doutb(w_n1209_0[1]),.din(n1209));
	jspl3 jspl3_w_n1211_0(.douta(w_n1211_0[0]),.doutb(w_n1211_0[1]),.doutc(w_n1211_0[2]),.din(n1211));
	jspl jspl_w_n1212_0(.douta(w_n1212_0[0]),.doutb(w_n1212_0[1]),.din(n1212));
	jspl jspl_w_n1216_0(.douta(w_n1216_0[0]),.doutb(w_n1216_0[1]),.din(n1216));
	jspl jspl_w_n1217_0(.douta(w_n1217_0[0]),.doutb(w_n1217_0[1]),.din(n1217));
	jspl3 jspl3_w_n1219_0(.douta(w_n1219_0[0]),.doutb(w_n1219_0[1]),.doutc(w_n1219_0[2]),.din(n1219));
	jspl jspl_w_n1220_0(.douta(w_n1220_0[0]),.doutb(w_n1220_0[1]),.din(n1220));
	jspl jspl_w_n1224_0(.douta(w_n1224_0[0]),.doutb(w_n1224_0[1]),.din(n1224));
	jspl3 jspl3_w_n1226_0(.douta(w_n1226_0[0]),.doutb(w_n1226_0[1]),.doutc(w_n1226_0[2]),.din(n1226));
	jspl jspl_w_n1227_0(.douta(w_n1227_0[0]),.doutb(w_n1227_0[1]),.din(n1227));
	jspl jspl_w_n1231_0(.douta(w_n1231_0[0]),.doutb(w_n1231_0[1]),.din(n1231));
	jspl3 jspl3_w_n1233_0(.douta(w_n1233_0[0]),.doutb(w_n1233_0[1]),.doutc(w_n1233_0[2]),.din(n1233));
	jspl jspl_w_n1234_0(.douta(w_n1234_0[0]),.doutb(w_n1234_0[1]),.din(n1234));
	jspl jspl_w_n1238_0(.douta(w_n1238_0[0]),.doutb(w_n1238_0[1]),.din(n1238));
	jspl3 jspl3_w_n1240_0(.douta(w_n1240_0[0]),.doutb(w_n1240_0[1]),.doutc(w_n1240_0[2]),.din(n1240));
	jspl jspl_w_n1241_0(.douta(w_n1241_0[0]),.doutb(w_n1241_0[1]),.din(n1241));
	jspl jspl_w_n1245_0(.douta(w_n1245_0[0]),.doutb(w_n1245_0[1]),.din(n1245));
	jspl jspl_w_n1246_0(.douta(w_n1246_0[0]),.doutb(w_n1246_0[1]),.din(n1246));
	jspl jspl_w_n1248_0(.douta(w_n1248_0[0]),.doutb(w_n1248_0[1]),.din(n1248));
	jspl jspl_w_n1251_0(.douta(w_n1251_0[0]),.doutb(w_n1251_0[1]),.din(n1251));
	jspl jspl_w_n1252_0(.douta(w_n1252_0[0]),.doutb(w_n1252_0[1]),.din(n1252));
	jspl3 jspl3_w_n1253_0(.douta(w_n1253_0[0]),.doutb(w_n1253_0[1]),.doutc(w_n1253_0[2]),.din(n1253));
	jspl jspl_w_n1253_1(.douta(w_n1253_1[0]),.doutb(w_n1253_1[1]),.din(w_n1253_0[0]));
	jspl3 jspl3_w_n1254_0(.douta(w_n1254_0[0]),.doutb(w_n1254_0[1]),.doutc(w_n1254_0[2]),.din(n1254));
	jspl jspl_w_n1279_0(.douta(w_n1279_0[0]),.doutb(w_n1279_0[1]),.din(n1279));
	jspl jspl_w_n1292_0(.douta(w_n1292_0[0]),.doutb(w_n1292_0[1]),.din(n1292));
	jspl jspl_w_n1296_0(.douta(w_n1296_0[0]),.doutb(w_n1296_0[1]),.din(n1296));
	jspl jspl_w_n1300_0(.douta(w_n1300_0[0]),.doutb(w_n1300_0[1]),.din(n1300));
	jspl jspl_w_n1305_0(.douta(w_n1305_0[0]),.doutb(w_n1305_0[1]),.din(n1305));
	jspl jspl_w_n1306_0(.douta(w_n1306_0[0]),.doutb(w_n1306_0[1]),.din(n1306));
	jspl jspl_w_n1307_0(.douta(w_n1307_0[0]),.doutb(w_n1307_0[1]),.din(n1307));
	jspl jspl_w_n1309_0(.douta(w_n1309_0[0]),.doutb(w_n1309_0[1]),.din(n1309));
	jspl jspl_w_n1311_0(.douta(w_n1311_0[0]),.doutb(w_n1311_0[1]),.din(n1311));
	jspl jspl_w_n1314_0(.douta(w_n1314_0[0]),.doutb(w_n1314_0[1]),.din(n1314));
	jspl jspl_w_n1315_0(.douta(w_n1315_0[0]),.doutb(w_n1315_0[1]),.din(n1315));
	jspl jspl_w_n1316_0(.douta(w_n1316_0[0]),.doutb(w_n1316_0[1]),.din(n1316));
	jspl3 jspl3_w_n1319_0(.douta(w_n1319_0[0]),.doutb(w_n1319_0[1]),.doutc(w_n1319_0[2]),.din(n1319));
	jspl3 jspl3_w_n1319_1(.douta(w_n1319_1[0]),.doutb(w_n1319_1[1]),.doutc(w_n1319_1[2]),.din(w_n1319_0[0]));
	jspl jspl_w_n1320_0(.douta(w_n1320_0[0]),.doutb(w_n1320_0[1]),.din(n1320));
	jspl3 jspl3_w_n1321_0(.douta(w_n1321_0[0]),.doutb(w_n1321_0[1]),.doutc(w_n1321_0[2]),.din(n1321));
	jspl jspl_w_n1322_0(.douta(w_n1322_0[0]),.doutb(w_n1322_0[1]),.din(n1322));
	jspl jspl_w_n1325_0(.douta(w_n1325_0[0]),.doutb(w_n1325_0[1]),.din(n1325));
	jspl jspl_w_n1330_0(.douta(w_n1330_0[0]),.doutb(w_n1330_0[1]),.din(n1330));
	jspl3 jspl3_w_n1332_0(.douta(w_n1332_0[0]),.doutb(w_n1332_0[1]),.doutc(w_n1332_0[2]),.din(n1332));
	jspl3 jspl3_w_n1332_1(.douta(w_n1332_1[0]),.doutb(w_n1332_1[1]),.doutc(w_n1332_1[2]),.din(w_n1332_0[0]));
	jspl3 jspl3_w_n1332_2(.douta(w_n1332_2[0]),.doutb(w_n1332_2[1]),.doutc(w_n1332_2[2]),.din(w_n1332_0[1]));
	jspl3 jspl3_w_n1332_3(.douta(w_n1332_3[0]),.doutb(w_n1332_3[1]),.doutc(w_n1332_3[2]),.din(w_n1332_0[2]));
	jspl3 jspl3_w_n1332_4(.douta(w_n1332_4[0]),.doutb(w_n1332_4[1]),.doutc(w_n1332_4[2]),.din(w_n1332_1[0]));
	jspl3 jspl3_w_n1332_5(.douta(w_n1332_5[0]),.doutb(w_n1332_5[1]),.doutc(w_n1332_5[2]),.din(w_n1332_1[1]));
	jspl3 jspl3_w_n1332_6(.douta(w_n1332_6[0]),.doutb(w_n1332_6[1]),.doutc(w_n1332_6[2]),.din(w_n1332_1[2]));
	jspl3 jspl3_w_n1332_7(.douta(w_n1332_7[0]),.doutb(w_n1332_7[1]),.doutc(w_n1332_7[2]),.din(w_n1332_2[0]));
	jspl3 jspl3_w_n1332_8(.douta(w_n1332_8[0]),.doutb(w_n1332_8[1]),.doutc(w_n1332_8[2]),.din(w_n1332_2[1]));
	jspl3 jspl3_w_n1332_9(.douta(w_n1332_9[0]),.doutb(w_n1332_9[1]),.doutc(w_n1332_9[2]),.din(w_n1332_2[2]));
	jspl3 jspl3_w_n1332_10(.douta(w_n1332_10[0]),.doutb(w_n1332_10[1]),.doutc(w_n1332_10[2]),.din(w_n1332_3[0]));
	jspl3 jspl3_w_n1332_11(.douta(w_n1332_11[0]),.doutb(w_n1332_11[1]),.doutc(w_n1332_11[2]),.din(w_n1332_3[1]));
	jspl3 jspl3_w_n1332_12(.douta(w_n1332_12[0]),.doutb(w_n1332_12[1]),.doutc(w_n1332_12[2]),.din(w_n1332_3[2]));
	jspl3 jspl3_w_n1332_13(.douta(w_n1332_13[0]),.doutb(w_n1332_13[1]),.doutc(w_n1332_13[2]),.din(w_n1332_4[0]));
	jspl3 jspl3_w_n1332_14(.douta(w_n1332_14[0]),.doutb(w_n1332_14[1]),.doutc(w_n1332_14[2]),.din(w_n1332_4[1]));
	jspl3 jspl3_w_n1332_15(.douta(w_n1332_15[0]),.doutb(w_n1332_15[1]),.doutc(w_n1332_15[2]),.din(w_n1332_4[2]));
	jspl3 jspl3_w_n1332_16(.douta(w_n1332_16[0]),.doutb(w_n1332_16[1]),.doutc(w_n1332_16[2]),.din(w_n1332_5[0]));
	jspl3 jspl3_w_n1332_17(.douta(w_n1332_17[0]),.doutb(w_n1332_17[1]),.doutc(w_n1332_17[2]),.din(w_n1332_5[1]));
	jspl3 jspl3_w_n1332_18(.douta(w_n1332_18[0]),.doutb(w_n1332_18[1]),.doutc(w_n1332_18[2]),.din(w_n1332_5[2]));
	jspl3 jspl3_w_n1332_19(.douta(w_n1332_19[0]),.doutb(w_n1332_19[1]),.doutc(w_n1332_19[2]),.din(w_n1332_6[0]));
	jspl3 jspl3_w_n1332_20(.douta(w_n1332_20[0]),.doutb(w_n1332_20[1]),.doutc(w_n1332_20[2]),.din(w_n1332_6[1]));
	jspl3 jspl3_w_n1332_21(.douta(w_n1332_21[0]),.doutb(w_n1332_21[1]),.doutc(w_n1332_21[2]),.din(w_n1332_6[2]));
	jspl3 jspl3_w_n1332_22(.douta(w_n1332_22[0]),.doutb(w_n1332_22[1]),.doutc(w_n1332_22[2]),.din(w_n1332_7[0]));
	jspl3 jspl3_w_n1332_23(.douta(w_n1332_23[0]),.doutb(w_n1332_23[1]),.doutc(w_n1332_23[2]),.din(w_n1332_7[1]));
	jspl3 jspl3_w_n1332_24(.douta(w_n1332_24[0]),.doutb(w_n1332_24[1]),.doutc(w_n1332_24[2]),.din(w_n1332_7[2]));
	jspl3 jspl3_w_n1332_25(.douta(w_n1332_25[0]),.doutb(w_n1332_25[1]),.doutc(w_n1332_25[2]),.din(w_n1332_8[0]));
	jspl3 jspl3_w_n1332_26(.douta(w_n1332_26[0]),.doutb(w_n1332_26[1]),.doutc(w_n1332_26[2]),.din(w_n1332_8[1]));
	jspl3 jspl3_w_n1332_27(.douta(w_n1332_27[0]),.doutb(w_n1332_27[1]),.doutc(w_n1332_27[2]),.din(w_n1332_8[2]));
	jspl3 jspl3_w_n1332_28(.douta(w_n1332_28[0]),.doutb(w_n1332_28[1]),.doutc(w_n1332_28[2]),.din(w_n1332_9[0]));
	jspl3 jspl3_w_n1332_29(.douta(w_n1332_29[0]),.doutb(w_n1332_29[1]),.doutc(w_n1332_29[2]),.din(w_n1332_9[1]));
	jspl3 jspl3_w_n1332_30(.douta(w_n1332_30[0]),.doutb(w_n1332_30[1]),.doutc(w_n1332_30[2]),.din(w_n1332_9[2]));
	jspl3 jspl3_w_n1332_31(.douta(w_n1332_31[0]),.doutb(w_n1332_31[1]),.doutc(w_n1332_31[2]),.din(w_n1332_10[0]));
	jspl3 jspl3_w_n1332_32(.douta(w_n1332_32[0]),.doutb(w_n1332_32[1]),.doutc(w_n1332_32[2]),.din(w_n1332_10[1]));
	jspl3 jspl3_w_n1332_33(.douta(w_n1332_33[0]),.doutb(w_n1332_33[1]),.doutc(w_n1332_33[2]),.din(w_n1332_10[2]));
	jspl3 jspl3_w_n1332_34(.douta(w_n1332_34[0]),.doutb(w_n1332_34[1]),.doutc(w_n1332_34[2]),.din(w_n1332_11[0]));
	jspl3 jspl3_w_n1332_35(.douta(w_n1332_35[0]),.doutb(w_n1332_35[1]),.doutc(w_n1332_35[2]),.din(w_n1332_11[1]));
	jspl3 jspl3_w_n1332_36(.douta(w_n1332_36[0]),.doutb(w_n1332_36[1]),.doutc(w_n1332_36[2]),.din(w_n1332_11[2]));
	jspl3 jspl3_w_n1332_37(.douta(w_n1332_37[0]),.doutb(w_n1332_37[1]),.doutc(w_n1332_37[2]),.din(w_n1332_12[0]));
	jspl3 jspl3_w_n1332_38(.douta(w_n1332_38[0]),.doutb(w_n1332_38[1]),.doutc(w_n1332_38[2]),.din(w_n1332_12[1]));
	jspl3 jspl3_w_n1332_39(.douta(w_n1332_39[0]),.doutb(w_n1332_39[1]),.doutc(w_n1332_39[2]),.din(w_n1332_12[2]));
	jspl3 jspl3_w_n1332_40(.douta(w_n1332_40[0]),.doutb(w_n1332_40[1]),.doutc(w_n1332_40[2]),.din(w_n1332_13[0]));
	jspl3 jspl3_w_n1332_41(.douta(w_n1332_41[0]),.doutb(w_n1332_41[1]),.doutc(w_n1332_41[2]),.din(w_n1332_13[1]));
	jspl3 jspl3_w_n1332_42(.douta(w_n1332_42[0]),.doutb(w_n1332_42[1]),.doutc(w_n1332_42[2]),.din(w_n1332_13[2]));
	jspl3 jspl3_w_n1332_43(.douta(w_n1332_43[0]),.doutb(w_n1332_43[1]),.doutc(w_n1332_43[2]),.din(w_n1332_14[0]));
	jspl3 jspl3_w_n1332_44(.douta(w_n1332_44[0]),.doutb(w_n1332_44[1]),.doutc(w_n1332_44[2]),.din(w_n1332_14[1]));
	jspl3 jspl3_w_n1332_45(.douta(w_n1332_45[0]),.doutb(w_n1332_45[1]),.doutc(w_n1332_45[2]),.din(w_n1332_14[2]));
	jspl3 jspl3_w_n1332_46(.douta(w_n1332_46[0]),.doutb(w_n1332_46[1]),.doutc(w_n1332_46[2]),.din(w_n1332_15[0]));
	jspl3 jspl3_w_n1332_47(.douta(w_n1332_47[0]),.doutb(w_n1332_47[1]),.doutc(w_n1332_47[2]),.din(w_n1332_15[1]));
	jspl3 jspl3_w_n1332_48(.douta(w_n1332_48[0]),.doutb(w_n1332_48[1]),.doutc(w_n1332_48[2]),.din(w_n1332_15[2]));
	jspl3 jspl3_w_n1332_49(.douta(w_n1332_49[0]),.doutb(w_n1332_49[1]),.doutc(w_n1332_49[2]),.din(w_n1332_16[0]));
	jspl3 jspl3_w_n1332_50(.douta(w_n1332_50[0]),.doutb(w_n1332_50[1]),.doutc(w_n1332_50[2]),.din(w_n1332_16[1]));
	jspl3 jspl3_w_n1332_51(.douta(w_n1332_51[0]),.doutb(w_n1332_51[1]),.doutc(w_n1332_51[2]),.din(w_n1332_16[2]));
	jspl3 jspl3_w_n1332_52(.douta(w_n1332_52[0]),.doutb(w_n1332_52[1]),.doutc(w_n1332_52[2]),.din(w_n1332_17[0]));
	jspl3 jspl3_w_n1332_53(.douta(w_n1332_53[0]),.doutb(w_n1332_53[1]),.doutc(w_n1332_53[2]),.din(w_n1332_17[1]));
	jspl3 jspl3_w_n1332_54(.douta(w_n1332_54[0]),.doutb(w_n1332_54[1]),.doutc(w_n1332_54[2]),.din(w_n1332_17[2]));
	jspl3 jspl3_w_n1332_55(.douta(w_n1332_55[0]),.doutb(w_n1332_55[1]),.doutc(w_n1332_55[2]),.din(w_n1332_18[0]));
	jspl3 jspl3_w_n1332_56(.douta(w_n1332_56[0]),.doutb(w_n1332_56[1]),.doutc(w_n1332_56[2]),.din(w_n1332_18[1]));
	jspl3 jspl3_w_n1332_57(.douta(w_n1332_57[0]),.doutb(w_n1332_57[1]),.doutc(w_n1332_57[2]),.din(w_n1332_18[2]));
	jspl3 jspl3_w_n1332_58(.douta(w_n1332_58[0]),.doutb(w_n1332_58[1]),.doutc(w_n1332_58[2]),.din(w_n1332_19[0]));
	jspl3 jspl3_w_n1332_59(.douta(w_n1332_59[0]),.doutb(w_n1332_59[1]),.doutc(w_n1332_59[2]),.din(w_n1332_19[1]));
	jspl3 jspl3_w_n1332_60(.douta(w_n1332_60[0]),.doutb(w_n1332_60[1]),.doutc(w_n1332_60[2]),.din(w_n1332_19[2]));
	jspl3 jspl3_w_n1332_61(.douta(w_n1332_61[0]),.doutb(w_n1332_61[1]),.doutc(w_n1332_61[2]),.din(w_n1332_20[0]));
	jspl3 jspl3_w_n1332_62(.douta(w_n1332_62[0]),.doutb(w_n1332_62[1]),.doutc(w_n1332_62[2]),.din(w_n1332_20[1]));
	jspl3 jspl3_w_n1332_63(.douta(w_n1332_63[0]),.doutb(w_n1332_63[1]),.doutc(w_n1332_63[2]),.din(w_n1332_20[2]));
	jspl3 jspl3_w_n1332_64(.douta(w_n1332_64[0]),.doutb(w_n1332_64[1]),.doutc(w_n1332_64[2]),.din(w_n1332_21[0]));
	jspl3 jspl3_w_n1332_65(.douta(w_n1332_65[0]),.doutb(w_n1332_65[1]),.doutc(w_n1332_65[2]),.din(w_n1332_21[1]));
	jspl3 jspl3_w_n1332_66(.douta(w_n1332_66[0]),.doutb(w_n1332_66[1]),.doutc(w_n1332_66[2]),.din(w_n1332_21[2]));
	jspl3 jspl3_w_n1332_67(.douta(w_n1332_67[0]),.doutb(w_n1332_67[1]),.doutc(w_n1332_67[2]),.din(w_n1332_22[0]));
	jspl3 jspl3_w_n1334_0(.douta(w_n1334_0[0]),.doutb(w_n1334_0[1]),.doutc(w_n1334_0[2]),.din(n1334));
	jspl jspl_w_n1335_0(.douta(w_n1335_0[0]),.doutb(w_n1335_0[1]),.din(n1335));
	jspl3 jspl3_w_n1342_0(.douta(w_n1342_0[0]),.doutb(w_n1342_0[1]),.doutc(w_n1342_0[2]),.din(n1342));
	jspl jspl_w_n1343_0(.douta(w_n1343_0[0]),.doutb(w_n1343_0[1]),.din(n1343));
	jspl jspl_w_n1346_0(.douta(w_n1346_0[0]),.doutb(w_n1346_0[1]),.din(n1346));
	jspl3 jspl3_w_n1351_0(.douta(w_n1351_0[0]),.doutb(w_n1351_0[1]),.doutc(w_n1351_0[2]),.din(n1351));
	jspl3 jspl3_w_n1353_0(.douta(w_n1353_0[0]),.doutb(w_n1353_0[1]),.doutc(w_n1353_0[2]),.din(n1353));
	jspl jspl_w_n1354_0(.douta(w_n1354_0[0]),.doutb(w_n1354_0[1]),.din(n1354));
	jspl3 jspl3_w_n1358_0(.douta(w_n1358_0[0]),.doutb(w_n1358_0[1]),.doutc(w_n1358_0[2]),.din(n1358));
	jspl3 jspl3_w_n1360_0(.douta(w_n1360_0[0]),.doutb(w_n1360_0[1]),.doutc(w_n1360_0[2]),.din(n1360));
	jspl jspl_w_n1361_0(.douta(w_n1361_0[0]),.doutb(w_n1361_0[1]),.din(n1361));
	jspl3 jspl3_w_n1365_0(.douta(w_n1365_0[0]),.doutb(w_n1365_0[1]),.doutc(w_n1365_0[2]),.din(n1365));
	jspl3 jspl3_w_n1367_0(.douta(w_n1367_0[0]),.doutb(w_n1367_0[1]),.doutc(w_n1367_0[2]),.din(n1367));
	jspl jspl_w_n1368_0(.douta(w_n1368_0[0]),.doutb(w_n1368_0[1]),.din(n1368));
	jspl3 jspl3_w_n1372_0(.douta(w_n1372_0[0]),.doutb(w_n1372_0[1]),.doutc(w_n1372_0[2]),.din(n1372));
	jspl3 jspl3_w_n1375_0(.douta(w_n1375_0[0]),.doutb(w_n1375_0[1]),.doutc(w_n1375_0[2]),.din(n1375));
	jspl jspl_w_n1376_0(.douta(w_n1376_0[0]),.doutb(w_n1376_0[1]),.din(n1376));
	jspl3 jspl3_w_n1380_0(.douta(w_n1380_0[0]),.doutb(w_n1380_0[1]),.doutc(w_n1380_0[2]),.din(n1380));
	jspl3 jspl3_w_n1382_0(.douta(w_n1382_0[0]),.doutb(w_n1382_0[1]),.doutc(w_n1382_0[2]),.din(n1382));
	jspl jspl_w_n1383_0(.douta(w_n1383_0[0]),.doutb(w_n1383_0[1]),.din(n1383));
	jspl3 jspl3_w_n1387_0(.douta(w_n1387_0[0]),.doutb(w_n1387_0[1]),.doutc(w_n1387_0[2]),.din(n1387));
	jspl3 jspl3_w_n1389_0(.douta(w_n1389_0[0]),.doutb(w_n1389_0[1]),.doutc(w_n1389_0[2]),.din(n1389));
	jspl jspl_w_n1390_0(.douta(w_n1390_0[0]),.doutb(w_n1390_0[1]),.din(n1390));
	jspl3 jspl3_w_n1394_0(.douta(w_n1394_0[0]),.doutb(w_n1394_0[1]),.doutc(w_n1394_0[2]),.din(n1394));
	jspl3 jspl3_w_n1396_0(.douta(w_n1396_0[0]),.doutb(w_n1396_0[1]),.doutc(w_n1396_0[2]),.din(n1396));
	jspl jspl_w_n1397_0(.douta(w_n1397_0[0]),.doutb(w_n1397_0[1]),.din(n1397));
	jspl3 jspl3_w_n1401_0(.douta(w_n1401_0[0]),.doutb(w_n1401_0[1]),.doutc(w_n1401_0[2]),.din(n1401));
	jspl3 jspl3_w_n1404_0(.douta(w_n1404_0[0]),.doutb(w_n1404_0[1]),.doutc(w_n1404_0[2]),.din(n1404));
	jspl jspl_w_n1405_0(.douta(w_n1405_0[0]),.doutb(w_n1405_0[1]),.din(n1405));
	jspl3 jspl3_w_n1409_0(.douta(w_n1409_0[0]),.doutb(w_n1409_0[1]),.doutc(w_n1409_0[2]),.din(n1409));
	jspl3 jspl3_w_n1412_0(.douta(w_n1412_0[0]),.doutb(w_n1412_0[1]),.doutc(w_n1412_0[2]),.din(n1412));
	jspl jspl_w_n1413_0(.douta(w_n1413_0[0]),.doutb(w_n1413_0[1]),.din(n1413));
	jspl jspl_w_n1417_0(.douta(w_n1417_0[0]),.doutb(w_n1417_0[1]),.din(n1417));
	jspl jspl_w_n1418_0(.douta(w_n1418_0[0]),.doutb(w_n1418_0[1]),.din(n1418));
	jspl3 jspl3_w_n1420_0(.douta(w_n1420_0[0]),.doutb(w_n1420_0[1]),.doutc(w_n1420_0[2]),.din(n1420));
	jspl jspl_w_n1420_1(.douta(w_n1420_1[0]),.doutb(w_n1420_1[1]),.din(w_n1420_0[0]));
	jspl3 jspl3_w_n1423_0(.douta(w_n1423_0[0]),.doutb(w_n1423_0[1]),.doutc(w_n1423_0[2]),.din(n1423));
	jspl3 jspl3_w_n1423_1(.douta(w_n1423_1[0]),.doutb(w_n1423_1[1]),.doutc(w_n1423_1[2]),.din(w_n1423_0[0]));
	jspl jspl_w_n1424_0(.douta(w_n1424_0[0]),.doutb(w_n1424_0[1]),.din(n1424));
	jspl jspl_w_n1426_0(.douta(w_n1426_0[0]),.doutb(w_n1426_0[1]),.din(n1426));
	jspl jspl_w_n1434_0(.douta(w_n1434_0[0]),.doutb(w_n1434_0[1]),.din(n1434));
	jspl jspl_w_n1435_0(.douta(w_n1435_0[0]),.doutb(w_n1435_0[1]),.din(n1435));
	jspl3 jspl3_w_n1440_0(.douta(w_n1440_0[0]),.doutb(w_n1440_0[1]),.doutc(w_n1440_0[2]),.din(n1440));
	jspl jspl_w_n1440_1(.douta(w_n1440_1[0]),.doutb(w_n1440_1[1]),.din(w_n1440_0[0]));
	jspl jspl_w_n1441_0(.douta(w_n1441_0[0]),.doutb(w_n1441_0[1]),.din(n1441));
	jspl3 jspl3_w_n1442_0(.douta(w_n1442_0[0]),.doutb(w_n1442_0[1]),.doutc(w_n1442_0[2]),.din(n1442));
	jspl jspl_w_n1443_0(.douta(w_n1443_0[0]),.doutb(w_n1443_0[1]),.din(n1443));
	jspl3 jspl3_w_n1445_0(.douta(w_n1445_0[0]),.doutb(w_n1445_0[1]),.doutc(w_n1445_0[2]),.din(n1445));
	jspl jspl_w_n1446_0(.douta(w_n1446_0[0]),.doutb(w_n1446_0[1]),.din(n1446));
	jspl jspl_w_n1451_0(.douta(w_n1451_0[0]),.doutb(w_n1451_0[1]),.din(n1451));
	jspl jspl_w_n1470_0(.douta(w_n1470_0[0]),.doutb(w_n1470_0[1]),.din(n1470));
	jspl jspl_w_n1513_0(.douta(w_n1513_0[0]),.doutb(w_n1513_0[1]),.din(n1513));
	jspl jspl_w_n1514_0(.douta(w_n1514_0[0]),.doutb(w_n1514_0[1]),.din(n1514));
	jspl3 jspl3_w_n1516_0(.douta(w_n1516_0[0]),.doutb(w_n1516_0[1]),.doutc(w_n1516_0[2]),.din(n1516));
	jspl3 jspl3_w_n1516_1(.douta(w_n1516_1[0]),.doutb(w_n1516_1[1]),.doutc(w_n1516_1[2]),.din(w_n1516_0[0]));
	jspl3 jspl3_w_n1516_2(.douta(w_n1516_2[0]),.doutb(w_n1516_2[1]),.doutc(w_n1516_2[2]),.din(w_n1516_0[1]));
	jspl3 jspl3_w_n1516_3(.douta(w_n1516_3[0]),.doutb(w_n1516_3[1]),.doutc(w_n1516_3[2]),.din(w_n1516_0[2]));
	jspl3 jspl3_w_n1516_4(.douta(w_n1516_4[0]),.doutb(w_n1516_4[1]),.doutc(w_n1516_4[2]),.din(w_n1516_1[0]));
	jspl3 jspl3_w_n1516_5(.douta(w_n1516_5[0]),.doutb(w_n1516_5[1]),.doutc(w_n1516_5[2]),.din(w_n1516_1[1]));
	jspl3 jspl3_w_n1516_6(.douta(w_n1516_6[0]),.doutb(w_n1516_6[1]),.doutc(w_n1516_6[2]),.din(w_n1516_1[2]));
	jspl3 jspl3_w_n1516_7(.douta(w_n1516_7[0]),.doutb(w_n1516_7[1]),.doutc(w_n1516_7[2]),.din(w_n1516_2[0]));
	jspl3 jspl3_w_n1516_8(.douta(w_n1516_8[0]),.doutb(w_n1516_8[1]),.doutc(w_n1516_8[2]),.din(w_n1516_2[1]));
	jspl3 jspl3_w_n1516_9(.douta(w_n1516_9[0]),.doutb(w_n1516_9[1]),.doutc(w_n1516_9[2]),.din(w_n1516_2[2]));
	jspl3 jspl3_w_n1516_10(.douta(w_n1516_10[0]),.doutb(w_n1516_10[1]),.doutc(w_n1516_10[2]),.din(w_n1516_3[0]));
	jspl3 jspl3_w_n1516_11(.douta(w_n1516_11[0]),.doutb(w_n1516_11[1]),.doutc(w_n1516_11[2]),.din(w_n1516_3[1]));
	jspl3 jspl3_w_n1516_12(.douta(w_n1516_12[0]),.doutb(w_n1516_12[1]),.doutc(w_n1516_12[2]),.din(w_n1516_3[2]));
	jspl3 jspl3_w_n1516_13(.douta(w_n1516_13[0]),.doutb(w_n1516_13[1]),.doutc(w_n1516_13[2]),.din(w_n1516_4[0]));
	jspl3 jspl3_w_n1516_14(.douta(w_n1516_14[0]),.doutb(w_n1516_14[1]),.doutc(w_n1516_14[2]),.din(w_n1516_4[1]));
	jspl3 jspl3_w_n1516_15(.douta(w_n1516_15[0]),.doutb(w_n1516_15[1]),.doutc(w_n1516_15[2]),.din(w_n1516_4[2]));
	jspl3 jspl3_w_n1516_16(.douta(w_n1516_16[0]),.doutb(w_n1516_16[1]),.doutc(w_n1516_16[2]),.din(w_n1516_5[0]));
	jspl3 jspl3_w_n1516_17(.douta(w_n1516_17[0]),.doutb(w_n1516_17[1]),.doutc(w_n1516_17[2]),.din(w_n1516_5[1]));
	jspl3 jspl3_w_n1516_18(.douta(w_n1516_18[0]),.doutb(w_n1516_18[1]),.doutc(w_n1516_18[2]),.din(w_n1516_5[2]));
	jspl3 jspl3_w_n1516_19(.douta(w_n1516_19[0]),.doutb(w_n1516_19[1]),.doutc(w_n1516_19[2]),.din(w_n1516_6[0]));
	jspl3 jspl3_w_n1516_20(.douta(w_n1516_20[0]),.doutb(w_n1516_20[1]),.doutc(w_n1516_20[2]),.din(w_n1516_6[1]));
	jspl3 jspl3_w_n1516_21(.douta(w_n1516_21[0]),.doutb(w_n1516_21[1]),.doutc(w_n1516_21[2]),.din(w_n1516_6[2]));
	jspl3 jspl3_w_n1516_22(.douta(w_n1516_22[0]),.doutb(w_n1516_22[1]),.doutc(w_n1516_22[2]),.din(w_n1516_7[0]));
	jspl3 jspl3_w_n1516_23(.douta(w_n1516_23[0]),.doutb(w_n1516_23[1]),.doutc(w_n1516_23[2]),.din(w_n1516_7[1]));
	jspl3 jspl3_w_n1516_24(.douta(w_n1516_24[0]),.doutb(w_n1516_24[1]),.doutc(w_n1516_24[2]),.din(w_n1516_7[2]));
	jspl3 jspl3_w_n1516_25(.douta(w_n1516_25[0]),.doutb(w_n1516_25[1]),.doutc(w_n1516_25[2]),.din(w_n1516_8[0]));
	jspl3 jspl3_w_n1516_26(.douta(w_n1516_26[0]),.doutb(w_n1516_26[1]),.doutc(w_n1516_26[2]),.din(w_n1516_8[1]));
	jspl3 jspl3_w_n1516_27(.douta(w_n1516_27[0]),.doutb(w_n1516_27[1]),.doutc(w_n1516_27[2]),.din(w_n1516_8[2]));
	jspl3 jspl3_w_n1516_28(.douta(w_n1516_28[0]),.doutb(w_n1516_28[1]),.doutc(w_n1516_28[2]),.din(w_n1516_9[0]));
	jspl3 jspl3_w_n1516_29(.douta(w_n1516_29[0]),.doutb(w_n1516_29[1]),.doutc(w_n1516_29[2]),.din(w_n1516_9[1]));
	jspl3 jspl3_w_n1516_30(.douta(w_n1516_30[0]),.doutb(w_n1516_30[1]),.doutc(w_n1516_30[2]),.din(w_n1516_9[2]));
	jspl3 jspl3_w_n1516_31(.douta(w_n1516_31[0]),.doutb(w_n1516_31[1]),.doutc(w_n1516_31[2]),.din(w_n1516_10[0]));
	jspl3 jspl3_w_n1516_32(.douta(w_n1516_32[0]),.doutb(w_n1516_32[1]),.doutc(w_n1516_32[2]),.din(w_n1516_10[1]));
	jspl3 jspl3_w_n1516_33(.douta(w_n1516_33[0]),.doutb(w_n1516_33[1]),.doutc(w_n1516_33[2]),.din(w_n1516_10[2]));
	jspl3 jspl3_w_n1516_34(.douta(w_n1516_34[0]),.doutb(w_n1516_34[1]),.doutc(w_n1516_34[2]),.din(w_n1516_11[0]));
	jspl3 jspl3_w_n1516_35(.douta(w_n1516_35[0]),.doutb(w_n1516_35[1]),.doutc(w_n1516_35[2]),.din(w_n1516_11[1]));
	jspl3 jspl3_w_n1516_36(.douta(w_n1516_36[0]),.doutb(w_n1516_36[1]),.doutc(w_n1516_36[2]),.din(w_n1516_11[2]));
	jspl3 jspl3_w_n1516_37(.douta(w_n1516_37[0]),.doutb(w_n1516_37[1]),.doutc(w_n1516_37[2]),.din(w_n1516_12[0]));
	jspl3 jspl3_w_n1516_38(.douta(w_n1516_38[0]),.doutb(w_n1516_38[1]),.doutc(w_n1516_38[2]),.din(w_n1516_12[1]));
	jspl3 jspl3_w_n1516_39(.douta(w_n1516_39[0]),.doutb(w_n1516_39[1]),.doutc(w_n1516_39[2]),.din(w_n1516_12[2]));
	jspl3 jspl3_w_n1516_40(.douta(w_n1516_40[0]),.doutb(w_n1516_40[1]),.doutc(w_n1516_40[2]),.din(w_n1516_13[0]));
	jspl3 jspl3_w_n1516_41(.douta(w_n1516_41[0]),.doutb(w_n1516_41[1]),.doutc(w_n1516_41[2]),.din(w_n1516_13[1]));
	jspl3 jspl3_w_n1516_42(.douta(w_n1516_42[0]),.doutb(w_n1516_42[1]),.doutc(w_n1516_42[2]),.din(w_n1516_13[2]));
	jspl3 jspl3_w_n1516_43(.douta(w_n1516_43[0]),.doutb(w_n1516_43[1]),.doutc(w_n1516_43[2]),.din(w_n1516_14[0]));
	jspl3 jspl3_w_n1516_44(.douta(w_n1516_44[0]),.doutb(w_n1516_44[1]),.doutc(w_n1516_44[2]),.din(w_n1516_14[1]));
	jspl3 jspl3_w_n1516_45(.douta(w_n1516_45[0]),.doutb(w_n1516_45[1]),.doutc(w_n1516_45[2]),.din(w_n1516_14[2]));
	jspl3 jspl3_w_n1516_46(.douta(w_n1516_46[0]),.doutb(w_n1516_46[1]),.doutc(w_n1516_46[2]),.din(w_n1516_15[0]));
	jspl3 jspl3_w_n1516_47(.douta(w_n1516_47[0]),.doutb(w_n1516_47[1]),.doutc(w_n1516_47[2]),.din(w_n1516_15[1]));
	jspl3 jspl3_w_n1516_48(.douta(w_n1516_48[0]),.doutb(w_n1516_48[1]),.doutc(w_n1516_48[2]),.din(w_n1516_15[2]));
	jspl3 jspl3_w_n1516_49(.douta(w_n1516_49[0]),.doutb(w_n1516_49[1]),.doutc(w_n1516_49[2]),.din(w_n1516_16[0]));
	jspl3 jspl3_w_n1516_50(.douta(w_n1516_50[0]),.doutb(w_n1516_50[1]),.doutc(w_n1516_50[2]),.din(w_n1516_16[1]));
	jspl3 jspl3_w_n1516_51(.douta(w_n1516_51[0]),.doutb(w_n1516_51[1]),.doutc(w_n1516_51[2]),.din(w_n1516_16[2]));
	jspl3 jspl3_w_n1516_52(.douta(w_n1516_52[0]),.doutb(w_n1516_52[1]),.doutc(w_n1516_52[2]),.din(w_n1516_17[0]));
	jspl3 jspl3_w_n1516_53(.douta(w_n1516_53[0]),.doutb(w_n1516_53[1]),.doutc(w_n1516_53[2]),.din(w_n1516_17[1]));
	jspl3 jspl3_w_n1516_54(.douta(w_n1516_54[0]),.doutb(w_n1516_54[1]),.doutc(w_n1516_54[2]),.din(w_n1516_17[2]));
	jspl3 jspl3_w_n1516_55(.douta(w_n1516_55[0]),.doutb(w_n1516_55[1]),.doutc(w_n1516_55[2]),.din(w_n1516_18[0]));
	jspl3 jspl3_w_n1516_56(.douta(w_n1516_56[0]),.doutb(w_n1516_56[1]),.doutc(w_n1516_56[2]),.din(w_n1516_18[1]));
	jspl3 jspl3_w_n1516_57(.douta(w_n1516_57[0]),.doutb(w_n1516_57[1]),.doutc(w_n1516_57[2]),.din(w_n1516_18[2]));
	jspl3 jspl3_w_n1516_58(.douta(w_n1516_58[0]),.doutb(w_n1516_58[1]),.doutc(w_n1516_58[2]),.din(w_n1516_19[0]));
	jspl3 jspl3_w_n1516_59(.douta(w_n1516_59[0]),.doutb(w_n1516_59[1]),.doutc(w_n1516_59[2]),.din(w_n1516_19[1]));
	jspl3 jspl3_w_n1516_60(.douta(w_n1516_60[0]),.doutb(w_n1516_60[1]),.doutc(w_n1516_60[2]),.din(w_n1516_19[2]));
	jspl3 jspl3_w_n1516_61(.douta(w_n1516_61[0]),.doutb(w_n1516_61[1]),.doutc(w_n1516_61[2]),.din(w_n1516_20[0]));
	jspl3 jspl3_w_n1516_62(.douta(w_n1516_62[0]),.doutb(w_n1516_62[1]),.doutc(w_n1516_62[2]),.din(w_n1516_20[1]));
	jspl jspl_w_n1518_0(.douta(w_n1518_0[0]),.doutb(w_n1518_0[1]),.din(n1518));
	jspl3 jspl3_w_n1520_0(.douta(w_n1520_0[0]),.doutb(w_n1520_0[1]),.doutc(w_n1520_0[2]),.din(n1520));
	jspl jspl_w_n1521_0(.douta(w_n1521_0[0]),.doutb(w_n1521_0[1]),.din(n1521));
	jspl jspl_w_n1523_0(.douta(w_n1523_0[0]),.doutb(w_n1523_0[1]),.din(n1523));
	jspl3 jspl3_w_n1528_0(.douta(w_n1528_0[0]),.doutb(w_n1528_0[1]),.doutc(w_n1528_0[2]),.din(n1528));
	jspl3 jspl3_w_n1531_0(.douta(w_n1531_0[0]),.doutb(w_n1531_0[1]),.doutc(w_n1531_0[2]),.din(n1531));
	jspl jspl_w_n1532_0(.douta(w_n1532_0[0]),.doutb(w_n1532_0[1]),.din(n1532));
	jspl jspl_w_n1536_0(.douta(w_n1536_0[0]),.doutb(w_n1536_0[1]),.din(n1536));
	jspl3 jspl3_w_n1538_0(.douta(w_n1538_0[0]),.doutb(w_n1538_0[1]),.doutc(w_n1538_0[2]),.din(n1538));
	jspl jspl_w_n1539_0(.douta(w_n1539_0[0]),.doutb(w_n1539_0[1]),.din(n1539));
	jspl jspl_w_n1543_0(.douta(w_n1543_0[0]),.doutb(w_n1543_0[1]),.din(n1543));
	jspl jspl_w_n1544_0(.douta(w_n1544_0[0]),.doutb(w_n1544_0[1]),.din(n1544));
	jspl3 jspl3_w_n1546_0(.douta(w_n1546_0[0]),.doutb(w_n1546_0[1]),.doutc(w_n1546_0[2]),.din(n1546));
	jspl jspl_w_n1547_0(.douta(w_n1547_0[0]),.doutb(w_n1547_0[1]),.din(n1547));
	jspl jspl_w_n1551_0(.douta(w_n1551_0[0]),.doutb(w_n1551_0[1]),.din(n1551));
	jspl jspl_w_n1552_0(.douta(w_n1552_0[0]),.doutb(w_n1552_0[1]),.din(n1552));
	jspl3 jspl3_w_n1554_0(.douta(w_n1554_0[0]),.doutb(w_n1554_0[1]),.doutc(w_n1554_0[2]),.din(n1554));
	jspl jspl_w_n1555_0(.douta(w_n1555_0[0]),.doutb(w_n1555_0[1]),.din(n1555));
	jspl jspl_w_n1559_0(.douta(w_n1559_0[0]),.doutb(w_n1559_0[1]),.din(n1559));
	jspl jspl_w_n1560_0(.douta(w_n1560_0[0]),.doutb(w_n1560_0[1]),.din(n1560));
	jspl3 jspl3_w_n1562_0(.douta(w_n1562_0[0]),.doutb(w_n1562_0[1]),.doutc(w_n1562_0[2]),.din(n1562));
	jspl jspl_w_n1563_0(.douta(w_n1563_0[0]),.doutb(w_n1563_0[1]),.din(n1563));
	jspl jspl_w_n1567_0(.douta(w_n1567_0[0]),.doutb(w_n1567_0[1]),.din(n1567));
	jspl3 jspl3_w_n1569_0(.douta(w_n1569_0[0]),.doutb(w_n1569_0[1]),.doutc(w_n1569_0[2]),.din(n1569));
	jspl jspl_w_n1570_0(.douta(w_n1570_0[0]),.doutb(w_n1570_0[1]),.din(n1570));
	jspl jspl_w_n1574_0(.douta(w_n1574_0[0]),.doutb(w_n1574_0[1]),.din(n1574));
	jspl jspl_w_n1575_0(.douta(w_n1575_0[0]),.doutb(w_n1575_0[1]),.din(n1575));
	jspl3 jspl3_w_n1577_0(.douta(w_n1577_0[0]),.doutb(w_n1577_0[1]),.doutc(w_n1577_0[2]),.din(n1577));
	jspl jspl_w_n1578_0(.douta(w_n1578_0[0]),.doutb(w_n1578_0[1]),.din(n1578));
	jspl jspl_w_n1582_0(.douta(w_n1582_0[0]),.doutb(w_n1582_0[1]),.din(n1582));
	jspl jspl_w_n1583_0(.douta(w_n1583_0[0]),.doutb(w_n1583_0[1]),.din(n1583));
	jspl3 jspl3_w_n1585_0(.douta(w_n1585_0[0]),.doutb(w_n1585_0[1]),.doutc(w_n1585_0[2]),.din(n1585));
	jspl jspl_w_n1586_0(.douta(w_n1586_0[0]),.doutb(w_n1586_0[1]),.din(n1586));
	jspl jspl_w_n1590_0(.douta(w_n1590_0[0]),.doutb(w_n1590_0[1]),.din(n1590));
	jspl jspl_w_n1591_0(.douta(w_n1591_0[0]),.doutb(w_n1591_0[1]),.din(n1591));
	jspl3 jspl3_w_n1593_0(.douta(w_n1593_0[0]),.doutb(w_n1593_0[1]),.doutc(w_n1593_0[2]),.din(n1593));
	jspl jspl_w_n1594_0(.douta(w_n1594_0[0]),.doutb(w_n1594_0[1]),.din(n1594));
	jspl jspl_w_n1598_0(.douta(w_n1598_0[0]),.doutb(w_n1598_0[1]),.din(n1598));
	jspl3 jspl3_w_n1600_0(.douta(w_n1600_0[0]),.doutb(w_n1600_0[1]),.doutc(w_n1600_0[2]),.din(n1600));
	jspl jspl_w_n1601_0(.douta(w_n1601_0[0]),.doutb(w_n1601_0[1]),.din(n1601));
	jspl jspl_w_n1627_0(.douta(w_n1627_0[0]),.doutb(w_n1627_0[1]),.din(n1627));
	jspl jspl_w_n1640_0(.douta(w_n1640_0[0]),.doutb(w_n1640_0[1]),.din(n1640));
	jspl jspl_w_n1653_0(.douta(w_n1653_0[0]),.doutb(w_n1653_0[1]),.din(n1653));
	jspl3 jspl3_w_n1659_0(.douta(w_n1659_0[0]),.doutb(w_n1659_0[1]),.doutc(w_n1659_0[2]),.din(n1659));
	jspl3 jspl3_w_n1662_0(.douta(w_n1662_0[0]),.doutb(w_n1662_0[1]),.doutc(w_n1662_0[2]),.din(n1662));
	jspl3 jspl3_w_n1665_0(.douta(w_n1665_0[0]),.doutb(w_n1665_0[1]),.doutc(w_n1665_0[2]),.din(n1665));
	jspl jspl_w_n1665_1(.douta(w_n1665_1[0]),.doutb(w_n1665_1[1]),.din(w_n1665_0[0]));
	jspl jspl_w_n1666_0(.douta(w_n1666_0[0]),.doutb(w_n1666_0[1]),.din(n1666));
	jspl jspl_w_n1667_0(.douta(w_n1667_0[0]),.doutb(w_n1667_0[1]),.din(n1667));
	jspl jspl_w_n1669_0(.douta(w_n1669_0[0]),.doutb(w_n1669_0[1]),.din(n1669));
	jspl jspl_w_n1671_0(.douta(w_n1671_0[0]),.doutb(w_n1671_0[1]),.din(n1671));
	jspl jspl_w_n1672_0(.douta(w_n1672_0[0]),.doutb(w_n1672_0[1]),.din(n1672));
	jspl3 jspl3_w_n1673_0(.douta(w_n1673_0[0]),.doutb(w_n1673_0[1]),.doutc(w_n1673_0[2]),.din(n1673));
	jspl jspl_w_n1677_0(.douta(w_n1677_0[0]),.doutb(w_n1677_0[1]),.din(n1677));
	jspl jspl_w_n1678_0(.douta(w_n1678_0[0]),.doutb(w_n1678_0[1]),.din(n1678));
	jspl3 jspl3_w_n1681_0(.douta(w_n1681_0[0]),.doutb(w_n1681_0[1]),.doutc(w_n1681_0[2]),.din(n1681));
	jspl3 jspl3_w_n1681_1(.douta(w_n1681_1[0]),.doutb(w_n1681_1[1]),.doutc(w_n1681_1[2]),.din(w_n1681_0[0]));
	jspl jspl_w_n1682_0(.douta(w_n1682_0[0]),.doutb(w_n1682_0[1]),.din(n1682));
	jspl3 jspl3_w_n1683_0(.douta(w_n1683_0[0]),.doutb(w_n1683_0[1]),.doutc(w_n1683_0[2]),.din(n1683));
	jspl jspl_w_n1684_0(.douta(w_n1684_0[0]),.doutb(w_n1684_0[1]),.din(n1684));
	jspl jspl_w_n1688_0(.douta(w_n1688_0[0]),.doutb(w_n1688_0[1]),.din(n1688));
	jspl jspl_w_n1689_0(.douta(w_n1689_0[0]),.doutb(w_n1689_0[1]),.din(n1689));
	jspl jspl_w_n1690_0(.douta(w_n1690_0[0]),.doutb(w_n1690_0[1]),.din(n1690));
	jspl3 jspl3_w_n1695_0(.douta(w_n1695_0[0]),.doutb(w_n1695_0[1]),.doutc(w_n1695_0[2]),.din(n1695));
	jspl3 jspl3_w_n1699_0(.douta(w_n1699_0[0]),.doutb(w_n1699_0[1]),.doutc(w_n1699_0[2]),.din(n1699));
	jspl3 jspl3_w_n1699_1(.douta(w_n1699_1[0]),.doutb(w_n1699_1[1]),.doutc(w_n1699_1[2]),.din(w_n1699_0[0]));
	jspl3 jspl3_w_n1699_2(.douta(w_n1699_2[0]),.doutb(w_n1699_2[1]),.doutc(w_n1699_2[2]),.din(w_n1699_0[1]));
	jspl3 jspl3_w_n1699_3(.douta(w_n1699_3[0]),.doutb(w_n1699_3[1]),.doutc(w_n1699_3[2]),.din(w_n1699_0[2]));
	jspl3 jspl3_w_n1699_4(.douta(w_n1699_4[0]),.doutb(w_n1699_4[1]),.doutc(w_n1699_4[2]),.din(w_n1699_1[0]));
	jspl3 jspl3_w_n1699_5(.douta(w_n1699_5[0]),.doutb(w_n1699_5[1]),.doutc(w_n1699_5[2]),.din(w_n1699_1[1]));
	jspl3 jspl3_w_n1699_6(.douta(w_n1699_6[0]),.doutb(w_n1699_6[1]),.doutc(w_n1699_6[2]),.din(w_n1699_1[2]));
	jspl3 jspl3_w_n1699_7(.douta(w_n1699_7[0]),.doutb(w_n1699_7[1]),.doutc(w_n1699_7[2]),.din(w_n1699_2[0]));
	jspl3 jspl3_w_n1699_8(.douta(w_n1699_8[0]),.doutb(w_n1699_8[1]),.doutc(w_n1699_8[2]),.din(w_n1699_2[1]));
	jspl3 jspl3_w_n1699_9(.douta(w_n1699_9[0]),.doutb(w_n1699_9[1]),.doutc(w_n1699_9[2]),.din(w_n1699_2[2]));
	jspl3 jspl3_w_n1699_10(.douta(w_n1699_10[0]),.doutb(w_n1699_10[1]),.doutc(w_n1699_10[2]),.din(w_n1699_3[0]));
	jspl3 jspl3_w_n1699_11(.douta(w_n1699_11[0]),.doutb(w_n1699_11[1]),.doutc(w_n1699_11[2]),.din(w_n1699_3[1]));
	jspl3 jspl3_w_n1699_12(.douta(w_n1699_12[0]),.doutb(w_n1699_12[1]),.doutc(w_n1699_12[2]),.din(w_n1699_3[2]));
	jspl3 jspl3_w_n1699_13(.douta(w_n1699_13[0]),.doutb(w_n1699_13[1]),.doutc(w_n1699_13[2]),.din(w_n1699_4[0]));
	jspl3 jspl3_w_n1699_14(.douta(w_n1699_14[0]),.doutb(w_n1699_14[1]),.doutc(w_n1699_14[2]),.din(w_n1699_4[1]));
	jspl3 jspl3_w_n1699_15(.douta(w_n1699_15[0]),.doutb(w_n1699_15[1]),.doutc(w_n1699_15[2]),.din(w_n1699_4[2]));
	jspl3 jspl3_w_n1699_16(.douta(w_n1699_16[0]),.doutb(w_n1699_16[1]),.doutc(w_n1699_16[2]),.din(w_n1699_5[0]));
	jspl3 jspl3_w_n1699_17(.douta(w_n1699_17[0]),.doutb(w_n1699_17[1]),.doutc(w_n1699_17[2]),.din(w_n1699_5[1]));
	jspl3 jspl3_w_n1699_18(.douta(w_n1699_18[0]),.doutb(w_n1699_18[1]),.doutc(w_n1699_18[2]),.din(w_n1699_5[2]));
	jspl3 jspl3_w_n1699_19(.douta(w_n1699_19[0]),.doutb(w_n1699_19[1]),.doutc(w_n1699_19[2]),.din(w_n1699_6[0]));
	jspl3 jspl3_w_n1699_20(.douta(w_n1699_20[0]),.doutb(w_n1699_20[1]),.doutc(w_n1699_20[2]),.din(w_n1699_6[1]));
	jspl3 jspl3_w_n1699_21(.douta(w_n1699_21[0]),.doutb(w_n1699_21[1]),.doutc(w_n1699_21[2]),.din(w_n1699_6[2]));
	jspl3 jspl3_w_n1699_22(.douta(w_n1699_22[0]),.doutb(w_n1699_22[1]),.doutc(w_n1699_22[2]),.din(w_n1699_7[0]));
	jspl3 jspl3_w_n1699_23(.douta(w_n1699_23[0]),.doutb(w_n1699_23[1]),.doutc(w_n1699_23[2]),.din(w_n1699_7[1]));
	jspl3 jspl3_w_n1699_24(.douta(w_n1699_24[0]),.doutb(w_n1699_24[1]),.doutc(w_n1699_24[2]),.din(w_n1699_7[2]));
	jspl3 jspl3_w_n1699_25(.douta(w_n1699_25[0]),.doutb(w_n1699_25[1]),.doutc(w_n1699_25[2]),.din(w_n1699_8[0]));
	jspl3 jspl3_w_n1699_26(.douta(w_n1699_26[0]),.doutb(w_n1699_26[1]),.doutc(w_n1699_26[2]),.din(w_n1699_8[1]));
	jspl3 jspl3_w_n1699_27(.douta(w_n1699_27[0]),.doutb(w_n1699_27[1]),.doutc(w_n1699_27[2]),.din(w_n1699_8[2]));
	jspl3 jspl3_w_n1699_28(.douta(w_n1699_28[0]),.doutb(w_n1699_28[1]),.doutc(w_n1699_28[2]),.din(w_n1699_9[0]));
	jspl3 jspl3_w_n1699_29(.douta(w_n1699_29[0]),.doutb(w_n1699_29[1]),.doutc(w_n1699_29[2]),.din(w_n1699_9[1]));
	jspl3 jspl3_w_n1699_30(.douta(w_n1699_30[0]),.doutb(w_n1699_30[1]),.doutc(w_n1699_30[2]),.din(w_n1699_9[2]));
	jspl3 jspl3_w_n1699_31(.douta(w_n1699_31[0]),.doutb(w_n1699_31[1]),.doutc(w_n1699_31[2]),.din(w_n1699_10[0]));
	jspl3 jspl3_w_n1699_32(.douta(w_n1699_32[0]),.doutb(w_n1699_32[1]),.doutc(w_n1699_32[2]),.din(w_n1699_10[1]));
	jspl3 jspl3_w_n1699_33(.douta(w_n1699_33[0]),.doutb(w_n1699_33[1]),.doutc(w_n1699_33[2]),.din(w_n1699_10[2]));
	jspl3 jspl3_w_n1699_34(.douta(w_n1699_34[0]),.doutb(w_n1699_34[1]),.doutc(w_n1699_34[2]),.din(w_n1699_11[0]));
	jspl3 jspl3_w_n1699_35(.douta(w_n1699_35[0]),.doutb(w_n1699_35[1]),.doutc(w_n1699_35[2]),.din(w_n1699_11[1]));
	jspl3 jspl3_w_n1699_36(.douta(w_n1699_36[0]),.doutb(w_n1699_36[1]),.doutc(w_n1699_36[2]),.din(w_n1699_11[2]));
	jspl3 jspl3_w_n1699_37(.douta(w_n1699_37[0]),.doutb(w_n1699_37[1]),.doutc(w_n1699_37[2]),.din(w_n1699_12[0]));
	jspl3 jspl3_w_n1699_38(.douta(w_n1699_38[0]),.doutb(w_n1699_38[1]),.doutc(w_n1699_38[2]),.din(w_n1699_12[1]));
	jspl3 jspl3_w_n1699_39(.douta(w_n1699_39[0]),.doutb(w_n1699_39[1]),.doutc(w_n1699_39[2]),.din(w_n1699_12[2]));
	jspl3 jspl3_w_n1699_40(.douta(w_n1699_40[0]),.doutb(w_n1699_40[1]),.doutc(w_n1699_40[2]),.din(w_n1699_13[0]));
	jspl3 jspl3_w_n1699_41(.douta(w_n1699_41[0]),.doutb(w_n1699_41[1]),.doutc(w_n1699_41[2]),.din(w_n1699_13[1]));
	jspl3 jspl3_w_n1699_42(.douta(w_n1699_42[0]),.doutb(w_n1699_42[1]),.doutc(w_n1699_42[2]),.din(w_n1699_13[2]));
	jspl3 jspl3_w_n1699_43(.douta(w_n1699_43[0]),.doutb(w_n1699_43[1]),.doutc(w_n1699_43[2]),.din(w_n1699_14[0]));
	jspl3 jspl3_w_n1699_44(.douta(w_n1699_44[0]),.doutb(w_n1699_44[1]),.doutc(w_n1699_44[2]),.din(w_n1699_14[1]));
	jspl3 jspl3_w_n1699_45(.douta(w_n1699_45[0]),.doutb(w_n1699_45[1]),.doutc(w_n1699_45[2]),.din(w_n1699_14[2]));
	jspl3 jspl3_w_n1699_46(.douta(w_n1699_46[0]),.doutb(w_n1699_46[1]),.doutc(w_n1699_46[2]),.din(w_n1699_15[0]));
	jspl3 jspl3_w_n1699_47(.douta(w_n1699_47[0]),.doutb(w_n1699_47[1]),.doutc(w_n1699_47[2]),.din(w_n1699_15[1]));
	jspl3 jspl3_w_n1699_48(.douta(w_n1699_48[0]),.doutb(w_n1699_48[1]),.doutc(w_n1699_48[2]),.din(w_n1699_15[2]));
	jspl3 jspl3_w_n1699_49(.douta(w_n1699_49[0]),.doutb(w_n1699_49[1]),.doutc(w_n1699_49[2]),.din(w_n1699_16[0]));
	jspl3 jspl3_w_n1699_50(.douta(w_n1699_50[0]),.doutb(w_n1699_50[1]),.doutc(w_n1699_50[2]),.din(w_n1699_16[1]));
	jspl3 jspl3_w_n1699_51(.douta(w_n1699_51[0]),.doutb(w_n1699_51[1]),.doutc(w_n1699_51[2]),.din(w_n1699_16[2]));
	jspl3 jspl3_w_n1699_52(.douta(w_n1699_52[0]),.doutb(w_n1699_52[1]),.doutc(w_n1699_52[2]),.din(w_n1699_17[0]));
	jspl3 jspl3_w_n1699_53(.douta(w_n1699_53[0]),.doutb(w_n1699_53[1]),.doutc(w_n1699_53[2]),.din(w_n1699_17[1]));
	jspl3 jspl3_w_n1699_54(.douta(w_n1699_54[0]),.doutb(w_n1699_54[1]),.doutc(w_n1699_54[2]),.din(w_n1699_17[2]));
	jspl3 jspl3_w_n1699_55(.douta(w_n1699_55[0]),.doutb(w_n1699_55[1]),.doutc(w_n1699_55[2]),.din(w_n1699_18[0]));
	jspl3 jspl3_w_n1699_56(.douta(w_n1699_56[0]),.doutb(w_n1699_56[1]),.doutc(w_n1699_56[2]),.din(w_n1699_18[1]));
	jspl3 jspl3_w_n1699_57(.douta(w_n1699_57[0]),.doutb(w_n1699_57[1]),.doutc(w_n1699_57[2]),.din(w_n1699_18[2]));
	jspl3 jspl3_w_n1699_58(.douta(w_n1699_58[0]),.doutb(w_n1699_58[1]),.doutc(w_n1699_58[2]),.din(w_n1699_19[0]));
	jspl3 jspl3_w_n1699_59(.douta(w_n1699_59[0]),.doutb(w_n1699_59[1]),.doutc(w_n1699_59[2]),.din(w_n1699_19[1]));
	jspl3 jspl3_w_n1699_60(.douta(w_n1699_60[0]),.doutb(w_n1699_60[1]),.doutc(w_n1699_60[2]),.din(w_n1699_19[2]));
	jspl3 jspl3_w_n1699_61(.douta(w_n1699_61[0]),.doutb(w_n1699_61[1]),.doutc(w_n1699_61[2]),.din(w_n1699_20[0]));
	jspl3 jspl3_w_n1699_62(.douta(w_n1699_62[0]),.doutb(w_n1699_62[1]),.doutc(w_n1699_62[2]),.din(w_n1699_20[1]));
	jspl3 jspl3_w_n1699_63(.douta(w_n1699_63[0]),.doutb(w_n1699_63[1]),.doutc(w_n1699_63[2]),.din(w_n1699_20[2]));
	jspl3 jspl3_w_n1699_64(.douta(w_n1699_64[0]),.doutb(w_n1699_64[1]),.doutc(w_n1699_64[2]),.din(w_n1699_21[0]));
	jspl3 jspl3_w_n1699_65(.douta(w_n1699_65[0]),.doutb(w_n1699_65[1]),.doutc(w_n1699_65[2]),.din(w_n1699_21[1]));
	jspl3 jspl3_w_n1699_66(.douta(w_n1699_66[0]),.doutb(w_n1699_66[1]),.doutc(w_n1699_66[2]),.din(w_n1699_21[2]));
	jspl jspl_w_n1699_67(.douta(w_n1699_67[0]),.doutb(w_n1699_67[1]),.din(w_n1699_22[0]));
	jspl3 jspl3_w_n1701_0(.douta(w_n1701_0[0]),.doutb(w_n1701_0[1]),.doutc(w_n1701_0[2]),.din(n1701));
	jspl jspl_w_n1702_0(.douta(w_n1702_0[0]),.doutb(w_n1702_0[1]),.din(n1702));
	jspl3 jspl3_w_n1709_0(.douta(w_n1709_0[0]),.doutb(w_n1709_0[1]),.doutc(w_n1709_0[2]),.din(n1709));
	jspl jspl_w_n1710_0(.douta(w_n1710_0[0]),.doutb(w_n1710_0[1]),.din(n1710));
	jspl jspl_w_n1713_0(.douta(w_n1713_0[0]),.doutb(w_n1713_0[1]),.din(n1713));
	jspl3 jspl3_w_n1718_0(.douta(w_n1718_0[0]),.doutb(w_n1718_0[1]),.doutc(w_n1718_0[2]),.din(n1718));
	jspl3 jspl3_w_n1720_0(.douta(w_n1720_0[0]),.doutb(w_n1720_0[1]),.doutc(w_n1720_0[2]),.din(n1720));
	jspl jspl_w_n1721_0(.douta(w_n1721_0[0]),.doutb(w_n1721_0[1]),.din(n1721));
	jspl3 jspl3_w_n1725_0(.douta(w_n1725_0[0]),.doutb(w_n1725_0[1]),.doutc(w_n1725_0[2]),.din(n1725));
	jspl3 jspl3_w_n1727_0(.douta(w_n1727_0[0]),.doutb(w_n1727_0[1]),.doutc(w_n1727_0[2]),.din(n1727));
	jspl jspl_w_n1728_0(.douta(w_n1728_0[0]),.doutb(w_n1728_0[1]),.din(n1728));
	jspl3 jspl3_w_n1732_0(.douta(w_n1732_0[0]),.doutb(w_n1732_0[1]),.doutc(w_n1732_0[2]),.din(n1732));
	jspl3 jspl3_w_n1735_0(.douta(w_n1735_0[0]),.doutb(w_n1735_0[1]),.doutc(w_n1735_0[2]),.din(n1735));
	jspl jspl_w_n1736_0(.douta(w_n1736_0[0]),.doutb(w_n1736_0[1]),.din(n1736));
	jspl3 jspl3_w_n1740_0(.douta(w_n1740_0[0]),.doutb(w_n1740_0[1]),.doutc(w_n1740_0[2]),.din(n1740));
	jspl3 jspl3_w_n1743_0(.douta(w_n1743_0[0]),.doutb(w_n1743_0[1]),.doutc(w_n1743_0[2]),.din(n1743));
	jspl jspl_w_n1744_0(.douta(w_n1744_0[0]),.doutb(w_n1744_0[1]),.din(n1744));
	jspl3 jspl3_w_n1748_0(.douta(w_n1748_0[0]),.doutb(w_n1748_0[1]),.doutc(w_n1748_0[2]),.din(n1748));
	jspl3 jspl3_w_n1750_0(.douta(w_n1750_0[0]),.doutb(w_n1750_0[1]),.doutc(w_n1750_0[2]),.din(n1750));
	jspl jspl_w_n1751_0(.douta(w_n1751_0[0]),.doutb(w_n1751_0[1]),.din(n1751));
	jspl3 jspl3_w_n1755_0(.douta(w_n1755_0[0]),.doutb(w_n1755_0[1]),.doutc(w_n1755_0[2]),.din(n1755));
	jspl3 jspl3_w_n1757_0(.douta(w_n1757_0[0]),.doutb(w_n1757_0[1]),.doutc(w_n1757_0[2]),.din(n1757));
	jspl jspl_w_n1758_0(.douta(w_n1758_0[0]),.doutb(w_n1758_0[1]),.din(n1758));
	jspl3 jspl3_w_n1762_0(.douta(w_n1762_0[0]),.doutb(w_n1762_0[1]),.doutc(w_n1762_0[2]),.din(n1762));
	jspl3 jspl3_w_n1764_0(.douta(w_n1764_0[0]),.doutb(w_n1764_0[1]),.doutc(w_n1764_0[2]),.din(n1764));
	jspl jspl_w_n1765_0(.douta(w_n1765_0[0]),.doutb(w_n1765_0[1]),.din(n1765));
	jspl3 jspl3_w_n1769_0(.douta(w_n1769_0[0]),.doutb(w_n1769_0[1]),.doutc(w_n1769_0[2]),.din(n1769));
	jspl3 jspl3_w_n1772_0(.douta(w_n1772_0[0]),.doutb(w_n1772_0[1]),.doutc(w_n1772_0[2]),.din(n1772));
	jspl jspl_w_n1773_0(.douta(w_n1773_0[0]),.doutb(w_n1773_0[1]),.din(n1773));
	jspl3 jspl3_w_n1777_0(.douta(w_n1777_0[0]),.doutb(w_n1777_0[1]),.doutc(w_n1777_0[2]),.din(n1777));
	jspl3 jspl3_w_n1779_0(.douta(w_n1779_0[0]),.doutb(w_n1779_0[1]),.doutc(w_n1779_0[2]),.din(n1779));
	jspl jspl_w_n1780_0(.douta(w_n1780_0[0]),.doutb(w_n1780_0[1]),.din(n1780));
	jspl3 jspl3_w_n1784_0(.douta(w_n1784_0[0]),.doutb(w_n1784_0[1]),.doutc(w_n1784_0[2]),.din(n1784));
	jspl3 jspl3_w_n1786_0(.douta(w_n1786_0[0]),.doutb(w_n1786_0[1]),.doutc(w_n1786_0[2]),.din(n1786));
	jspl jspl_w_n1787_0(.douta(w_n1787_0[0]),.doutb(w_n1787_0[1]),.din(n1787));
	jspl3 jspl3_w_n1791_0(.douta(w_n1791_0[0]),.doutb(w_n1791_0[1]),.doutc(w_n1791_0[2]),.din(n1791));
	jspl3 jspl3_w_n1793_0(.douta(w_n1793_0[0]),.doutb(w_n1793_0[1]),.doutc(w_n1793_0[2]),.din(n1793));
	jspl jspl_w_n1794_0(.douta(w_n1794_0[0]),.doutb(w_n1794_0[1]),.din(n1794));
	jspl3 jspl3_w_n1798_0(.douta(w_n1798_0[0]),.doutb(w_n1798_0[1]),.doutc(w_n1798_0[2]),.din(n1798));
	jspl3 jspl3_w_n1801_0(.douta(w_n1801_0[0]),.doutb(w_n1801_0[1]),.doutc(w_n1801_0[2]),.din(n1801));
	jspl3 jspl3_w_n1804_0(.douta(w_n1804_0[0]),.doutb(w_n1804_0[1]),.doutc(w_n1804_0[2]),.din(n1804));
	jspl jspl_w_n1804_1(.douta(w_n1804_1[0]),.doutb(w_n1804_1[1]),.din(w_n1804_0[0]));
	jspl3 jspl3_w_n1805_0(.douta(w_n1805_0[0]),.doutb(w_n1805_0[1]),.doutc(w_n1805_0[2]),.din(n1805));
	jspl jspl_w_n1809_0(.douta(w_n1809_0[0]),.doutb(w_n1809_0[1]),.din(n1809));
	jspl jspl_w_n1810_0(.douta(w_n1810_0[0]),.doutb(w_n1810_0[1]),.din(n1810));
	jspl jspl_w_n1812_0(.douta(w_n1812_0[0]),.doutb(w_n1812_0[1]),.din(n1812));
	jspl jspl_w_n1813_0(.douta(w_n1813_0[0]),.doutb(w_n1813_0[1]),.din(n1813));
	jspl jspl_w_n1817_0(.douta(w_n1817_0[0]),.doutb(w_n1817_0[1]),.din(n1817));
	jspl jspl_w_n1819_0(.douta(w_n1819_0[0]),.doutb(w_n1819_0[1]),.din(n1819));
	jspl jspl_w_n1839_0(.douta(w_n1839_0[0]),.doutb(w_n1839_0[1]),.din(n1839));
	jspl jspl_w_n1887_0(.douta(w_n1887_0[0]),.doutb(w_n1887_0[1]),.din(n1887));
	jspl jspl_w_n1888_0(.douta(w_n1888_0[0]),.doutb(w_n1888_0[1]),.din(n1888));
	jspl3 jspl3_w_n1891_0(.douta(w_n1891_0[0]),.doutb(w_n1891_0[1]),.doutc(w_n1891_0[2]),.din(n1891));
	jspl3 jspl3_w_n1894_0(.douta(w_n1894_0[0]),.doutb(w_n1894_0[1]),.doutc(w_n1894_0[2]),.din(n1894));
	jspl jspl_w_n1894_1(.douta(w_n1894_1[0]),.doutb(w_n1894_1[1]),.din(w_n1894_0[0]));
	jspl jspl_w_n1895_0(.douta(w_n1895_0[0]),.doutb(w_n1895_0[1]),.din(n1895));
	jspl3 jspl3_w_n1896_0(.douta(w_n1896_0[0]),.doutb(w_n1896_0[1]),.doutc(w_n1896_0[2]),.din(n1896));
	jspl jspl_w_n1897_0(.douta(w_n1897_0[0]),.doutb(w_n1897_0[1]),.din(n1897));
	jspl3 jspl3_w_n1898_0(.douta(w_n1898_0[0]),.doutb(w_n1898_0[1]),.doutc(w_n1898_0[2]),.din(n1898));
	jspl jspl_w_n1899_0(.douta(w_n1899_0[0]),.doutb(w_n1899_0[1]),.din(n1899));
	jspl3 jspl3_w_n1904_0(.douta(w_n1904_0[0]),.doutb(w_n1904_0[1]),.doutc(w_n1904_0[2]),.din(n1904));
	jspl jspl_w_n1904_1(.douta(w_n1904_1[0]),.doutb(w_n1904_1[1]),.din(w_n1904_0[0]));
	jspl jspl_w_n1908_0(.douta(w_n1908_0[0]),.doutb(w_n1908_0[1]),.din(n1908));
	jspl jspl_w_n1911_0(.douta(w_n1911_0[0]),.doutb(w_n1911_0[1]),.din(n1911));
	jspl3 jspl3_w_n1912_0(.douta(w_n1912_0[0]),.doutb(w_n1912_0[1]),.doutc(w_n1912_0[2]),.din(n1912));
	jspl3 jspl3_w_n1912_1(.douta(w_n1912_1[0]),.doutb(w_n1912_1[1]),.doutc(w_n1912_1[2]),.din(w_n1912_0[0]));
	jspl3 jspl3_w_n1912_2(.douta(w_n1912_2[0]),.doutb(w_n1912_2[1]),.doutc(w_n1912_2[2]),.din(w_n1912_0[1]));
	jspl3 jspl3_w_n1912_3(.douta(w_n1912_3[0]),.doutb(w_n1912_3[1]),.doutc(w_n1912_3[2]),.din(w_n1912_0[2]));
	jspl3 jspl3_w_n1912_4(.douta(w_n1912_4[0]),.doutb(w_n1912_4[1]),.doutc(w_n1912_4[2]),.din(w_n1912_1[0]));
	jspl3 jspl3_w_n1912_5(.douta(w_n1912_5[0]),.doutb(w_n1912_5[1]),.doutc(w_n1912_5[2]),.din(w_n1912_1[1]));
	jspl3 jspl3_w_n1912_6(.douta(w_n1912_6[0]),.doutb(w_n1912_6[1]),.doutc(w_n1912_6[2]),.din(w_n1912_1[2]));
	jspl3 jspl3_w_n1912_7(.douta(w_n1912_7[0]),.doutb(w_n1912_7[1]),.doutc(w_n1912_7[2]),.din(w_n1912_2[0]));
	jspl3 jspl3_w_n1912_8(.douta(w_n1912_8[0]),.doutb(w_n1912_8[1]),.doutc(w_n1912_8[2]),.din(w_n1912_2[1]));
	jspl3 jspl3_w_n1912_9(.douta(w_n1912_9[0]),.doutb(w_n1912_9[1]),.doutc(w_n1912_9[2]),.din(w_n1912_2[2]));
	jspl3 jspl3_w_n1912_10(.douta(w_n1912_10[0]),.doutb(w_n1912_10[1]),.doutc(w_n1912_10[2]),.din(w_n1912_3[0]));
	jspl3 jspl3_w_n1912_11(.douta(w_n1912_11[0]),.doutb(w_n1912_11[1]),.doutc(w_n1912_11[2]),.din(w_n1912_3[1]));
	jspl3 jspl3_w_n1912_12(.douta(w_n1912_12[0]),.doutb(w_n1912_12[1]),.doutc(w_n1912_12[2]),.din(w_n1912_3[2]));
	jspl3 jspl3_w_n1912_13(.douta(w_n1912_13[0]),.doutb(w_n1912_13[1]),.doutc(w_n1912_13[2]),.din(w_n1912_4[0]));
	jspl3 jspl3_w_n1912_14(.douta(w_n1912_14[0]),.doutb(w_n1912_14[1]),.doutc(w_n1912_14[2]),.din(w_n1912_4[1]));
	jspl3 jspl3_w_n1912_15(.douta(w_n1912_15[0]),.doutb(w_n1912_15[1]),.doutc(w_n1912_15[2]),.din(w_n1912_4[2]));
	jspl3 jspl3_w_n1912_16(.douta(w_n1912_16[0]),.doutb(w_n1912_16[1]),.doutc(w_n1912_16[2]),.din(w_n1912_5[0]));
	jspl3 jspl3_w_n1912_17(.douta(w_n1912_17[0]),.doutb(w_n1912_17[1]),.doutc(w_n1912_17[2]),.din(w_n1912_5[1]));
	jspl3 jspl3_w_n1912_18(.douta(w_n1912_18[0]),.doutb(w_n1912_18[1]),.doutc(w_n1912_18[2]),.din(w_n1912_5[2]));
	jspl3 jspl3_w_n1912_19(.douta(w_n1912_19[0]),.doutb(w_n1912_19[1]),.doutc(w_n1912_19[2]),.din(w_n1912_6[0]));
	jspl3 jspl3_w_n1912_20(.douta(w_n1912_20[0]),.doutb(w_n1912_20[1]),.doutc(w_n1912_20[2]),.din(w_n1912_6[1]));
	jspl3 jspl3_w_n1912_21(.douta(w_n1912_21[0]),.doutb(w_n1912_21[1]),.doutc(w_n1912_21[2]),.din(w_n1912_6[2]));
	jspl3 jspl3_w_n1912_22(.douta(w_n1912_22[0]),.doutb(w_n1912_22[1]),.doutc(w_n1912_22[2]),.din(w_n1912_7[0]));
	jspl3 jspl3_w_n1912_23(.douta(w_n1912_23[0]),.doutb(w_n1912_23[1]),.doutc(w_n1912_23[2]),.din(w_n1912_7[1]));
	jspl3 jspl3_w_n1912_24(.douta(w_n1912_24[0]),.doutb(w_n1912_24[1]),.doutc(w_n1912_24[2]),.din(w_n1912_7[2]));
	jspl3 jspl3_w_n1912_25(.douta(w_n1912_25[0]),.doutb(w_n1912_25[1]),.doutc(w_n1912_25[2]),.din(w_n1912_8[0]));
	jspl3 jspl3_w_n1912_26(.douta(w_n1912_26[0]),.doutb(w_n1912_26[1]),.doutc(w_n1912_26[2]),.din(w_n1912_8[1]));
	jspl3 jspl3_w_n1912_27(.douta(w_n1912_27[0]),.doutb(w_n1912_27[1]),.doutc(w_n1912_27[2]),.din(w_n1912_8[2]));
	jspl3 jspl3_w_n1912_28(.douta(w_n1912_28[0]),.doutb(w_n1912_28[1]),.doutc(w_n1912_28[2]),.din(w_n1912_9[0]));
	jspl3 jspl3_w_n1912_29(.douta(w_n1912_29[0]),.doutb(w_n1912_29[1]),.doutc(w_n1912_29[2]),.din(w_n1912_9[1]));
	jspl3 jspl3_w_n1912_30(.douta(w_n1912_30[0]),.doutb(w_n1912_30[1]),.doutc(w_n1912_30[2]),.din(w_n1912_9[2]));
	jspl3 jspl3_w_n1912_31(.douta(w_n1912_31[0]),.doutb(w_n1912_31[1]),.doutc(w_n1912_31[2]),.din(w_n1912_10[0]));
	jspl3 jspl3_w_n1912_32(.douta(w_n1912_32[0]),.doutb(w_n1912_32[1]),.doutc(w_n1912_32[2]),.din(w_n1912_10[1]));
	jspl3 jspl3_w_n1912_33(.douta(w_n1912_33[0]),.doutb(w_n1912_33[1]),.doutc(w_n1912_33[2]),.din(w_n1912_10[2]));
	jspl3 jspl3_w_n1912_34(.douta(w_n1912_34[0]),.doutb(w_n1912_34[1]),.doutc(w_n1912_34[2]),.din(w_n1912_11[0]));
	jspl3 jspl3_w_n1912_35(.douta(w_n1912_35[0]),.doutb(w_n1912_35[1]),.doutc(w_n1912_35[2]),.din(w_n1912_11[1]));
	jspl3 jspl3_w_n1912_36(.douta(w_n1912_36[0]),.doutb(w_n1912_36[1]),.doutc(w_n1912_36[2]),.din(w_n1912_11[2]));
	jspl3 jspl3_w_n1912_37(.douta(w_n1912_37[0]),.doutb(w_n1912_37[1]),.doutc(w_n1912_37[2]),.din(w_n1912_12[0]));
	jspl3 jspl3_w_n1912_38(.douta(w_n1912_38[0]),.doutb(w_n1912_38[1]),.doutc(w_n1912_38[2]),.din(w_n1912_12[1]));
	jspl3 jspl3_w_n1912_39(.douta(w_n1912_39[0]),.doutb(w_n1912_39[1]),.doutc(w_n1912_39[2]),.din(w_n1912_12[2]));
	jspl3 jspl3_w_n1912_40(.douta(w_n1912_40[0]),.doutb(w_n1912_40[1]),.doutc(w_n1912_40[2]),.din(w_n1912_13[0]));
	jspl3 jspl3_w_n1912_41(.douta(w_n1912_41[0]),.doutb(w_n1912_41[1]),.doutc(w_n1912_41[2]),.din(w_n1912_13[1]));
	jspl3 jspl3_w_n1912_42(.douta(w_n1912_42[0]),.doutb(w_n1912_42[1]),.doutc(w_n1912_42[2]),.din(w_n1912_13[2]));
	jspl3 jspl3_w_n1912_43(.douta(w_n1912_43[0]),.doutb(w_n1912_43[1]),.doutc(w_n1912_43[2]),.din(w_n1912_14[0]));
	jspl3 jspl3_w_n1912_44(.douta(w_n1912_44[0]),.doutb(w_n1912_44[1]),.doutc(w_n1912_44[2]),.din(w_n1912_14[1]));
	jspl3 jspl3_w_n1912_45(.douta(w_n1912_45[0]),.doutb(w_n1912_45[1]),.doutc(w_n1912_45[2]),.din(w_n1912_14[2]));
	jspl3 jspl3_w_n1912_46(.douta(w_n1912_46[0]),.doutb(w_n1912_46[1]),.doutc(w_n1912_46[2]),.din(w_n1912_15[0]));
	jspl3 jspl3_w_n1912_47(.douta(w_n1912_47[0]),.doutb(w_n1912_47[1]),.doutc(w_n1912_47[2]),.din(w_n1912_15[1]));
	jspl3 jspl3_w_n1912_48(.douta(w_n1912_48[0]),.doutb(w_n1912_48[1]),.doutc(w_n1912_48[2]),.din(w_n1912_15[2]));
	jspl3 jspl3_w_n1912_49(.douta(w_n1912_49[0]),.doutb(w_n1912_49[1]),.doutc(w_n1912_49[2]),.din(w_n1912_16[0]));
	jspl3 jspl3_w_n1912_50(.douta(w_n1912_50[0]),.doutb(w_n1912_50[1]),.doutc(w_n1912_50[2]),.din(w_n1912_16[1]));
	jspl3 jspl3_w_n1912_51(.douta(w_n1912_51[0]),.doutb(w_n1912_51[1]),.doutc(w_n1912_51[2]),.din(w_n1912_16[2]));
	jspl3 jspl3_w_n1912_52(.douta(w_n1912_52[0]),.doutb(w_n1912_52[1]),.doutc(w_n1912_52[2]),.din(w_n1912_17[0]));
	jspl3 jspl3_w_n1912_53(.douta(w_n1912_53[0]),.doutb(w_n1912_53[1]),.doutc(w_n1912_53[2]),.din(w_n1912_17[1]));
	jspl3 jspl3_w_n1912_54(.douta(w_n1912_54[0]),.doutb(w_n1912_54[1]),.doutc(w_n1912_54[2]),.din(w_n1912_17[2]));
	jspl3 jspl3_w_n1912_55(.douta(w_n1912_55[0]),.doutb(w_n1912_55[1]),.doutc(w_n1912_55[2]),.din(w_n1912_18[0]));
	jspl3 jspl3_w_n1912_56(.douta(w_n1912_56[0]),.doutb(w_n1912_56[1]),.doutc(w_n1912_56[2]),.din(w_n1912_18[1]));
	jspl3 jspl3_w_n1912_57(.douta(w_n1912_57[0]),.doutb(w_n1912_57[1]),.doutc(w_n1912_57[2]),.din(w_n1912_18[2]));
	jspl3 jspl3_w_n1912_58(.douta(w_n1912_58[0]),.doutb(w_n1912_58[1]),.doutc(w_n1912_58[2]),.din(w_n1912_19[0]));
	jspl3 jspl3_w_n1912_59(.douta(w_n1912_59[0]),.doutb(w_n1912_59[1]),.doutc(w_n1912_59[2]),.din(w_n1912_19[1]));
	jspl jspl_w_n1912_60(.douta(w_n1912_60[0]),.doutb(w_n1912_60[1]),.din(w_n1912_19[2]));
	jspl3 jspl3_w_n1916_0(.douta(w_n1916_0[0]),.doutb(w_n1916_0[1]),.doutc(w_n1916_0[2]),.din(n1916));
	jspl jspl_w_n1917_0(.douta(w_n1917_0[0]),.doutb(w_n1917_0[1]),.din(n1917));
	jspl jspl_w_n1919_0(.douta(w_n1919_0[0]),.doutb(w_n1919_0[1]),.din(n1919));
	jspl jspl_w_n1924_0(.douta(w_n1924_0[0]),.doutb(w_n1924_0[1]),.din(n1924));
	jspl jspl_w_n1925_0(.douta(w_n1925_0[0]),.doutb(w_n1925_0[1]),.din(n1925));
	jspl3 jspl3_w_n1927_0(.douta(w_n1927_0[0]),.doutb(w_n1927_0[1]),.doutc(w_n1927_0[2]),.din(n1927));
	jspl jspl_w_n1928_0(.douta(w_n1928_0[0]),.doutb(w_n1928_0[1]),.din(n1928));
	jspl jspl_w_n1932_0(.douta(w_n1932_0[0]),.doutb(w_n1932_0[1]),.din(n1932));
	jspl3 jspl3_w_n1934_0(.douta(w_n1934_0[0]),.doutb(w_n1934_0[1]),.doutc(w_n1934_0[2]),.din(n1934));
	jspl jspl_w_n1935_0(.douta(w_n1935_0[0]),.doutb(w_n1935_0[1]),.din(n1935));
	jspl jspl_w_n1939_0(.douta(w_n1939_0[0]),.doutb(w_n1939_0[1]),.din(n1939));
	jspl jspl_w_n1940_0(.douta(w_n1940_0[0]),.doutb(w_n1940_0[1]),.din(n1940));
	jspl3 jspl3_w_n1942_0(.douta(w_n1942_0[0]),.doutb(w_n1942_0[1]),.doutc(w_n1942_0[2]),.din(n1942));
	jspl jspl_w_n1943_0(.douta(w_n1943_0[0]),.doutb(w_n1943_0[1]),.din(n1943));
	jspl jspl_w_n1947_0(.douta(w_n1947_0[0]),.doutb(w_n1947_0[1]),.din(n1947));
	jspl jspl_w_n1948_0(.douta(w_n1948_0[0]),.doutb(w_n1948_0[1]),.din(n1948));
	jspl3 jspl3_w_n1950_0(.douta(w_n1950_0[0]),.doutb(w_n1950_0[1]),.doutc(w_n1950_0[2]),.din(n1950));
	jspl jspl_w_n1951_0(.douta(w_n1951_0[0]),.doutb(w_n1951_0[1]),.din(n1951));
	jspl jspl_w_n1955_0(.douta(w_n1955_0[0]),.doutb(w_n1955_0[1]),.din(n1955));
	jspl3 jspl3_w_n1957_0(.douta(w_n1957_0[0]),.doutb(w_n1957_0[1]),.doutc(w_n1957_0[2]),.din(n1957));
	jspl jspl_w_n1958_0(.douta(w_n1958_0[0]),.doutb(w_n1958_0[1]),.din(n1958));
	jspl jspl_w_n1962_0(.douta(w_n1962_0[0]),.doutb(w_n1962_0[1]),.din(n1962));
	jspl3 jspl3_w_n1964_0(.douta(w_n1964_0[0]),.doutb(w_n1964_0[1]),.doutc(w_n1964_0[2]),.din(n1964));
	jspl jspl_w_n1965_0(.douta(w_n1965_0[0]),.doutb(w_n1965_0[1]),.din(n1965));
	jspl jspl_w_n1969_0(.douta(w_n1969_0[0]),.doutb(w_n1969_0[1]),.din(n1969));
	jspl jspl_w_n1970_0(.douta(w_n1970_0[0]),.doutb(w_n1970_0[1]),.din(n1970));
	jspl3 jspl3_w_n1972_0(.douta(w_n1972_0[0]),.doutb(w_n1972_0[1]),.doutc(w_n1972_0[2]),.din(n1972));
	jspl jspl_w_n1973_0(.douta(w_n1973_0[0]),.doutb(w_n1973_0[1]),.din(n1973));
	jspl jspl_w_n1977_0(.douta(w_n1977_0[0]),.doutb(w_n1977_0[1]),.din(n1977));
	jspl jspl_w_n1978_0(.douta(w_n1978_0[0]),.doutb(w_n1978_0[1]),.din(n1978));
	jspl3 jspl3_w_n1980_0(.douta(w_n1980_0[0]),.doutb(w_n1980_0[1]),.doutc(w_n1980_0[2]),.din(n1980));
	jspl jspl_w_n1981_0(.douta(w_n1981_0[0]),.doutb(w_n1981_0[1]),.din(n1981));
	jspl3 jspl3_w_n1985_0(.douta(w_n1985_0[0]),.doutb(w_n1985_0[1]),.doutc(w_n1985_0[2]),.din(n1985));
	jspl3 jspl3_w_n1988_0(.douta(w_n1988_0[0]),.doutb(w_n1988_0[1]),.doutc(w_n1988_0[2]),.din(n1988));
	jspl jspl_w_n1989_0(.douta(w_n1989_0[0]),.doutb(w_n1989_0[1]),.din(n1989));
	jspl jspl_w_n1993_0(.douta(w_n1993_0[0]),.doutb(w_n1993_0[1]),.din(n1993));
	jspl3 jspl3_w_n1995_0(.douta(w_n1995_0[0]),.doutb(w_n1995_0[1]),.doutc(w_n1995_0[2]),.din(n1995));
	jspl jspl_w_n1996_0(.douta(w_n1996_0[0]),.doutb(w_n1996_0[1]),.din(n1996));
	jspl jspl_w_n2000_0(.douta(w_n2000_0[0]),.doutb(w_n2000_0[1]),.din(n2000));
	jspl jspl_w_n2001_0(.douta(w_n2001_0[0]),.doutb(w_n2001_0[1]),.din(n2001));
	jspl3 jspl3_w_n2003_0(.douta(w_n2003_0[0]),.doutb(w_n2003_0[1]),.doutc(w_n2003_0[2]),.din(n2003));
	jspl jspl_w_n2004_0(.douta(w_n2004_0[0]),.doutb(w_n2004_0[1]),.din(n2004));
	jspl jspl_w_n2008_0(.douta(w_n2008_0[0]),.doutb(w_n2008_0[1]),.din(n2008));
	jspl jspl_w_n2009_0(.douta(w_n2009_0[0]),.doutb(w_n2009_0[1]),.din(n2009));
	jspl3 jspl3_w_n2011_0(.douta(w_n2011_0[0]),.doutb(w_n2011_0[1]),.doutc(w_n2011_0[2]),.din(n2011));
	jspl jspl_w_n2012_0(.douta(w_n2012_0[0]),.doutb(w_n2012_0[1]),.din(n2012));
	jspl jspl_w_n2033_0(.douta(w_n2033_0[0]),.doutb(w_n2033_0[1]),.din(n2033));
	jspl jspl_w_n2040_0(.douta(w_n2040_0[0]),.doutb(w_n2040_0[1]),.din(n2040));
	jspl jspl_w_n2050_0(.douta(w_n2050_0[0]),.doutb(w_n2050_0[1]),.din(n2050));
	jspl jspl_w_n2054_0(.douta(w_n2054_0[0]),.doutb(w_n2054_0[1]),.din(n2054));
	jspl jspl_w_n2067_0(.douta(w_n2067_0[0]),.doutb(w_n2067_0[1]),.din(n2067));
	jspl jspl_w_n2079_0(.douta(w_n2079_0[0]),.doutb(w_n2079_0[1]),.din(n2079));
	jspl jspl_w_n2081_0(.douta(w_n2081_0[0]),.doutb(w_n2081_0[1]),.din(n2081));
	jspl jspl_w_n2082_0(.douta(w_n2082_0[0]),.doutb(w_n2082_0[1]),.din(n2082));
	jspl jspl_w_n2085_0(.douta(w_n2085_0[0]),.doutb(w_n2085_0[1]),.din(n2085));
	jspl jspl_w_n2089_0(.douta(w_n2089_0[0]),.doutb(w_n2089_0[1]),.din(n2089));
	jspl jspl_w_n2091_0(.douta(w_n2091_0[0]),.doutb(w_n2091_0[1]),.din(n2091));
	jspl3 jspl3_w_n2092_0(.douta(w_n2092_0[0]),.doutb(w_n2092_0[1]),.doutc(w_n2092_0[2]),.din(n2092));
	jspl jspl_w_n2097_0(.douta(w_n2097_0[0]),.doutb(w_n2097_0[1]),.din(n2097));
	jspl jspl_w_n2100_0(.douta(w_n2100_0[0]),.doutb(w_n2100_0[1]),.din(n2100));
	jspl jspl_w_n2104_0(.douta(w_n2104_0[0]),.doutb(w_n2104_0[1]),.din(n2104));
	jspl3 jspl3_w_n2108_0(.douta(w_n2108_0[0]),.doutb(w_n2108_0[1]),.doutc(w_n2108_0[2]),.din(n2108));
	jspl3 jspl3_w_n2108_1(.douta(w_n2108_1[0]),.doutb(w_n2108_1[1]),.doutc(w_n2108_1[2]),.din(w_n2108_0[0]));
	jspl3 jspl3_w_n2108_2(.douta(w_n2108_2[0]),.doutb(w_n2108_2[1]),.doutc(w_n2108_2[2]),.din(w_n2108_0[1]));
	jspl3 jspl3_w_n2108_3(.douta(w_n2108_3[0]),.doutb(w_n2108_3[1]),.doutc(w_n2108_3[2]),.din(w_n2108_0[2]));
	jspl3 jspl3_w_n2108_4(.douta(w_n2108_4[0]),.doutb(w_n2108_4[1]),.doutc(w_n2108_4[2]),.din(w_n2108_1[0]));
	jspl3 jspl3_w_n2108_5(.douta(w_n2108_5[0]),.doutb(w_n2108_5[1]),.doutc(w_n2108_5[2]),.din(w_n2108_1[1]));
	jspl3 jspl3_w_n2108_6(.douta(w_n2108_6[0]),.doutb(w_n2108_6[1]),.doutc(w_n2108_6[2]),.din(w_n2108_1[2]));
	jspl3 jspl3_w_n2108_7(.douta(w_n2108_7[0]),.doutb(w_n2108_7[1]),.doutc(w_n2108_7[2]),.din(w_n2108_2[0]));
	jspl3 jspl3_w_n2108_8(.douta(w_n2108_8[0]),.doutb(w_n2108_8[1]),.doutc(w_n2108_8[2]),.din(w_n2108_2[1]));
	jspl3 jspl3_w_n2108_9(.douta(w_n2108_9[0]),.doutb(w_n2108_9[1]),.doutc(w_n2108_9[2]),.din(w_n2108_2[2]));
	jspl3 jspl3_w_n2108_10(.douta(w_n2108_10[0]),.doutb(w_n2108_10[1]),.doutc(w_n2108_10[2]),.din(w_n2108_3[0]));
	jspl3 jspl3_w_n2108_11(.douta(w_n2108_11[0]),.doutb(w_n2108_11[1]),.doutc(w_n2108_11[2]),.din(w_n2108_3[1]));
	jspl3 jspl3_w_n2108_12(.douta(w_n2108_12[0]),.doutb(w_n2108_12[1]),.doutc(w_n2108_12[2]),.din(w_n2108_3[2]));
	jspl3 jspl3_w_n2108_13(.douta(w_n2108_13[0]),.doutb(w_n2108_13[1]),.doutc(w_n2108_13[2]),.din(w_n2108_4[0]));
	jspl3 jspl3_w_n2108_14(.douta(w_n2108_14[0]),.doutb(w_n2108_14[1]),.doutc(w_n2108_14[2]),.din(w_n2108_4[1]));
	jspl3 jspl3_w_n2108_15(.douta(w_n2108_15[0]),.doutb(w_n2108_15[1]),.doutc(w_n2108_15[2]),.din(w_n2108_4[2]));
	jspl3 jspl3_w_n2108_16(.douta(w_n2108_16[0]),.doutb(w_n2108_16[1]),.doutc(w_n2108_16[2]),.din(w_n2108_5[0]));
	jspl3 jspl3_w_n2108_17(.douta(w_n2108_17[0]),.doutb(w_n2108_17[1]),.doutc(w_n2108_17[2]),.din(w_n2108_5[1]));
	jspl3 jspl3_w_n2108_18(.douta(w_n2108_18[0]),.doutb(w_n2108_18[1]),.doutc(w_n2108_18[2]),.din(w_n2108_5[2]));
	jspl3 jspl3_w_n2108_19(.douta(w_n2108_19[0]),.doutb(w_n2108_19[1]),.doutc(w_n2108_19[2]),.din(w_n2108_6[0]));
	jspl3 jspl3_w_n2108_20(.douta(w_n2108_20[0]),.doutb(w_n2108_20[1]),.doutc(w_n2108_20[2]),.din(w_n2108_6[1]));
	jspl3 jspl3_w_n2108_21(.douta(w_n2108_21[0]),.doutb(w_n2108_21[1]),.doutc(w_n2108_21[2]),.din(w_n2108_6[2]));
	jspl3 jspl3_w_n2108_22(.douta(w_n2108_22[0]),.doutb(w_n2108_22[1]),.doutc(w_n2108_22[2]),.din(w_n2108_7[0]));
	jspl3 jspl3_w_n2108_23(.douta(w_n2108_23[0]),.doutb(w_n2108_23[1]),.doutc(w_n2108_23[2]),.din(w_n2108_7[1]));
	jspl3 jspl3_w_n2108_24(.douta(w_n2108_24[0]),.doutb(w_n2108_24[1]),.doutc(w_n2108_24[2]),.din(w_n2108_7[2]));
	jspl3 jspl3_w_n2108_25(.douta(w_n2108_25[0]),.doutb(w_n2108_25[1]),.doutc(w_n2108_25[2]),.din(w_n2108_8[0]));
	jspl3 jspl3_w_n2108_26(.douta(w_n2108_26[0]),.doutb(w_n2108_26[1]),.doutc(w_n2108_26[2]),.din(w_n2108_8[1]));
	jspl3 jspl3_w_n2108_27(.douta(w_n2108_27[0]),.doutb(w_n2108_27[1]),.doutc(w_n2108_27[2]),.din(w_n2108_8[2]));
	jspl3 jspl3_w_n2108_28(.douta(w_n2108_28[0]),.doutb(w_n2108_28[1]),.doutc(w_n2108_28[2]),.din(w_n2108_9[0]));
	jspl3 jspl3_w_n2108_29(.douta(w_n2108_29[0]),.doutb(w_n2108_29[1]),.doutc(w_n2108_29[2]),.din(w_n2108_9[1]));
	jspl3 jspl3_w_n2108_30(.douta(w_n2108_30[0]),.doutb(w_n2108_30[1]),.doutc(w_n2108_30[2]),.din(w_n2108_9[2]));
	jspl3 jspl3_w_n2108_31(.douta(w_n2108_31[0]),.doutb(w_n2108_31[1]),.doutc(w_n2108_31[2]),.din(w_n2108_10[0]));
	jspl3 jspl3_w_n2108_32(.douta(w_n2108_32[0]),.doutb(w_n2108_32[1]),.doutc(w_n2108_32[2]),.din(w_n2108_10[1]));
	jspl3 jspl3_w_n2108_33(.douta(w_n2108_33[0]),.doutb(w_n2108_33[1]),.doutc(w_n2108_33[2]),.din(w_n2108_10[2]));
	jspl3 jspl3_w_n2108_34(.douta(w_n2108_34[0]),.doutb(w_n2108_34[1]),.doutc(w_n2108_34[2]),.din(w_n2108_11[0]));
	jspl3 jspl3_w_n2108_35(.douta(w_n2108_35[0]),.doutb(w_n2108_35[1]),.doutc(w_n2108_35[2]),.din(w_n2108_11[1]));
	jspl3 jspl3_w_n2108_36(.douta(w_n2108_36[0]),.doutb(w_n2108_36[1]),.doutc(w_n2108_36[2]),.din(w_n2108_11[2]));
	jspl3 jspl3_w_n2108_37(.douta(w_n2108_37[0]),.doutb(w_n2108_37[1]),.doutc(w_n2108_37[2]),.din(w_n2108_12[0]));
	jspl3 jspl3_w_n2108_38(.douta(w_n2108_38[0]),.doutb(w_n2108_38[1]),.doutc(w_n2108_38[2]),.din(w_n2108_12[1]));
	jspl3 jspl3_w_n2108_39(.douta(w_n2108_39[0]),.doutb(w_n2108_39[1]),.doutc(w_n2108_39[2]),.din(w_n2108_12[2]));
	jspl3 jspl3_w_n2108_40(.douta(w_n2108_40[0]),.doutb(w_n2108_40[1]),.doutc(w_n2108_40[2]),.din(w_n2108_13[0]));
	jspl3 jspl3_w_n2108_41(.douta(w_n2108_41[0]),.doutb(w_n2108_41[1]),.doutc(w_n2108_41[2]),.din(w_n2108_13[1]));
	jspl3 jspl3_w_n2108_42(.douta(w_n2108_42[0]),.doutb(w_n2108_42[1]),.doutc(w_n2108_42[2]),.din(w_n2108_13[2]));
	jspl3 jspl3_w_n2108_43(.douta(w_n2108_43[0]),.doutb(w_n2108_43[1]),.doutc(w_n2108_43[2]),.din(w_n2108_14[0]));
	jspl3 jspl3_w_n2108_44(.douta(w_n2108_44[0]),.doutb(w_n2108_44[1]),.doutc(w_n2108_44[2]),.din(w_n2108_14[1]));
	jspl3 jspl3_w_n2108_45(.douta(w_n2108_45[0]),.doutb(w_n2108_45[1]),.doutc(w_n2108_45[2]),.din(w_n2108_14[2]));
	jspl3 jspl3_w_n2108_46(.douta(w_n2108_46[0]),.doutb(w_n2108_46[1]),.doutc(w_n2108_46[2]),.din(w_n2108_15[0]));
	jspl3 jspl3_w_n2108_47(.douta(w_n2108_47[0]),.doutb(w_n2108_47[1]),.doutc(w_n2108_47[2]),.din(w_n2108_15[1]));
	jspl3 jspl3_w_n2108_48(.douta(w_n2108_48[0]),.doutb(w_n2108_48[1]),.doutc(w_n2108_48[2]),.din(w_n2108_15[2]));
	jspl3 jspl3_w_n2108_49(.douta(w_n2108_49[0]),.doutb(w_n2108_49[1]),.doutc(w_n2108_49[2]),.din(w_n2108_16[0]));
	jspl3 jspl3_w_n2108_50(.douta(w_n2108_50[0]),.doutb(w_n2108_50[1]),.doutc(w_n2108_50[2]),.din(w_n2108_16[1]));
	jspl3 jspl3_w_n2108_51(.douta(w_n2108_51[0]),.doutb(w_n2108_51[1]),.doutc(w_n2108_51[2]),.din(w_n2108_16[2]));
	jspl3 jspl3_w_n2108_52(.douta(w_n2108_52[0]),.doutb(w_n2108_52[1]),.doutc(w_n2108_52[2]),.din(w_n2108_17[0]));
	jspl3 jspl3_w_n2108_53(.douta(w_n2108_53[0]),.doutb(w_n2108_53[1]),.doutc(w_n2108_53[2]),.din(w_n2108_17[1]));
	jspl3 jspl3_w_n2108_54(.douta(w_n2108_54[0]),.doutb(w_n2108_54[1]),.doutc(w_n2108_54[2]),.din(w_n2108_17[2]));
	jspl3 jspl3_w_n2108_55(.douta(w_n2108_55[0]),.doutb(w_n2108_55[1]),.doutc(w_n2108_55[2]),.din(w_n2108_18[0]));
	jspl3 jspl3_w_n2108_56(.douta(w_n2108_56[0]),.doutb(w_n2108_56[1]),.doutc(w_n2108_56[2]),.din(w_n2108_18[1]));
	jspl3 jspl3_w_n2108_57(.douta(w_n2108_57[0]),.doutb(w_n2108_57[1]),.doutc(w_n2108_57[2]),.din(w_n2108_18[2]));
	jspl3 jspl3_w_n2108_58(.douta(w_n2108_58[0]),.doutb(w_n2108_58[1]),.doutc(w_n2108_58[2]),.din(w_n2108_19[0]));
	jspl3 jspl3_w_n2108_59(.douta(w_n2108_59[0]),.doutb(w_n2108_59[1]),.doutc(w_n2108_59[2]),.din(w_n2108_19[1]));
	jspl3 jspl3_w_n2108_60(.douta(w_n2108_60[0]),.doutb(w_n2108_60[1]),.doutc(w_n2108_60[2]),.din(w_n2108_19[2]));
	jspl3 jspl3_w_n2108_61(.douta(w_n2108_61[0]),.doutb(w_n2108_61[1]),.doutc(w_n2108_61[2]),.din(w_n2108_20[0]));
	jspl3 jspl3_w_n2108_62(.douta(w_n2108_62[0]),.doutb(w_n2108_62[1]),.doutc(w_n2108_62[2]),.din(w_n2108_20[1]));
	jspl3 jspl3_w_n2108_63(.douta(w_n2108_63[0]),.doutb(w_n2108_63[1]),.doutc(w_n2108_63[2]),.din(w_n2108_20[2]));
	jspl3 jspl3_w_n2108_64(.douta(w_n2108_64[0]),.doutb(w_n2108_64[1]),.doutc(w_n2108_64[2]),.din(w_n2108_21[0]));
	jspl jspl_w_n2108_65(.douta(w_n2108_65[0]),.doutb(w_n2108_65[1]),.din(w_n2108_21[1]));
	jspl3 jspl3_w_n2110_0(.douta(w_n2110_0[0]),.doutb(w_n2110_0[1]),.doutc(w_n2110_0[2]),.din(n2110));
	jspl3 jspl3_w_n2110_1(.douta(w_n2110_1[0]),.doutb(w_n2110_1[1]),.doutc(w_n2110_1[2]),.din(w_n2110_0[0]));
	jspl jspl_w_n2111_0(.douta(w_n2111_0[0]),.doutb(w_n2111_0[1]),.din(n2111));
	jspl3 jspl3_w_n2112_0(.douta(w_n2112_0[0]),.doutb(w_n2112_0[1]),.doutc(w_n2112_0[2]),.din(n2112));
	jspl jspl_w_n2113_0(.douta(w_n2113_0[0]),.doutb(w_n2113_0[1]),.din(n2113));
	jspl3 jspl3_w_n2115_0(.douta(w_n2115_0[0]),.doutb(w_n2115_0[1]),.doutc(w_n2115_0[2]),.din(n2115));
	jspl jspl_w_n2116_0(.douta(w_n2116_0[0]),.doutb(w_n2116_0[1]),.din(n2116));
	jspl3 jspl3_w_n2123_0(.douta(w_n2123_0[0]),.doutb(w_n2123_0[1]),.doutc(w_n2123_0[2]),.din(n2123));
	jspl jspl_w_n2124_0(.douta(w_n2124_0[0]),.doutb(w_n2124_0[1]),.din(n2124));
	jspl jspl_w_n2127_0(.douta(w_n2127_0[0]),.doutb(w_n2127_0[1]),.din(n2127));
	jspl jspl_w_n2128_0(.douta(w_n2128_0[0]),.doutb(w_n2128_0[1]),.din(n2128));
	jspl3 jspl3_w_n2133_0(.douta(w_n2133_0[0]),.doutb(w_n2133_0[1]),.doutc(w_n2133_0[2]),.din(n2133));
	jspl3 jspl3_w_n2135_0(.douta(w_n2135_0[0]),.doutb(w_n2135_0[1]),.doutc(w_n2135_0[2]),.din(n2135));
	jspl jspl_w_n2136_0(.douta(w_n2136_0[0]),.doutb(w_n2136_0[1]),.din(n2136));
	jspl3 jspl3_w_n2140_0(.douta(w_n2140_0[0]),.doutb(w_n2140_0[1]),.doutc(w_n2140_0[2]),.din(n2140));
	jspl3 jspl3_w_n2143_0(.douta(w_n2143_0[0]),.doutb(w_n2143_0[1]),.doutc(w_n2143_0[2]),.din(n2143));
	jspl jspl_w_n2144_0(.douta(w_n2144_0[0]),.doutb(w_n2144_0[1]),.din(n2144));
	jspl3 jspl3_w_n2148_0(.douta(w_n2148_0[0]),.doutb(w_n2148_0[1]),.doutc(w_n2148_0[2]),.din(n2148));
	jspl3 jspl3_w_n2150_0(.douta(w_n2150_0[0]),.doutb(w_n2150_0[1]),.doutc(w_n2150_0[2]),.din(n2150));
	jspl jspl_w_n2151_0(.douta(w_n2151_0[0]),.doutb(w_n2151_0[1]),.din(n2151));
	jspl3 jspl3_w_n2155_0(.douta(w_n2155_0[0]),.doutb(w_n2155_0[1]),.doutc(w_n2155_0[2]),.din(n2155));
	jspl3 jspl3_w_n2158_0(.douta(w_n2158_0[0]),.doutb(w_n2158_0[1]),.doutc(w_n2158_0[2]),.din(n2158));
	jspl jspl_w_n2159_0(.douta(w_n2159_0[0]),.doutb(w_n2159_0[1]),.din(n2159));
	jspl3 jspl3_w_n2163_0(.douta(w_n2163_0[0]),.doutb(w_n2163_0[1]),.doutc(w_n2163_0[2]),.din(n2163));
	jspl3 jspl3_w_n2165_0(.douta(w_n2165_0[0]),.doutb(w_n2165_0[1]),.doutc(w_n2165_0[2]),.din(n2165));
	jspl jspl_w_n2166_0(.douta(w_n2166_0[0]),.doutb(w_n2166_0[1]),.din(n2166));
	jspl3 jspl3_w_n2170_0(.douta(w_n2170_0[0]),.doutb(w_n2170_0[1]),.doutc(w_n2170_0[2]),.din(n2170));
	jspl3 jspl3_w_n2172_0(.douta(w_n2172_0[0]),.doutb(w_n2172_0[1]),.doutc(w_n2172_0[2]),.din(n2172));
	jspl jspl_w_n2173_0(.douta(w_n2173_0[0]),.doutb(w_n2173_0[1]),.din(n2173));
	jspl3 jspl3_w_n2177_0(.douta(w_n2177_0[0]),.doutb(w_n2177_0[1]),.doutc(w_n2177_0[2]),.din(n2177));
	jspl3 jspl3_w_n2180_0(.douta(w_n2180_0[0]),.doutb(w_n2180_0[1]),.doutc(w_n2180_0[2]),.din(n2180));
	jspl jspl_w_n2181_0(.douta(w_n2181_0[0]),.doutb(w_n2181_0[1]),.din(n2181));
	jspl3 jspl3_w_n2185_0(.douta(w_n2185_0[0]),.doutb(w_n2185_0[1]),.doutc(w_n2185_0[2]),.din(n2185));
	jspl3 jspl3_w_n2188_0(.douta(w_n2188_0[0]),.doutb(w_n2188_0[1]),.doutc(w_n2188_0[2]),.din(n2188));
	jspl jspl_w_n2189_0(.douta(w_n2189_0[0]),.doutb(w_n2189_0[1]),.din(n2189));
	jspl3 jspl3_w_n2193_0(.douta(w_n2193_0[0]),.doutb(w_n2193_0[1]),.doutc(w_n2193_0[2]),.din(n2193));
	jspl3 jspl3_w_n2195_0(.douta(w_n2195_0[0]),.doutb(w_n2195_0[1]),.doutc(w_n2195_0[2]),.din(n2195));
	jspl jspl_w_n2196_0(.douta(w_n2196_0[0]),.doutb(w_n2196_0[1]),.din(n2196));
	jspl jspl_w_n2200_0(.douta(w_n2200_0[0]),.doutb(w_n2200_0[1]),.din(n2200));
	jspl3 jspl3_w_n2202_0(.douta(w_n2202_0[0]),.doutb(w_n2202_0[1]),.doutc(w_n2202_0[2]),.din(n2202));
	jspl jspl_w_n2203_0(.douta(w_n2203_0[0]),.doutb(w_n2203_0[1]),.din(n2203));
	jspl3 jspl3_w_n2207_0(.douta(w_n2207_0[0]),.doutb(w_n2207_0[1]),.doutc(w_n2207_0[2]),.din(n2207));
	jspl3 jspl3_w_n2210_0(.douta(w_n2210_0[0]),.doutb(w_n2210_0[1]),.doutc(w_n2210_0[2]),.din(n2210));
	jspl jspl_w_n2211_0(.douta(w_n2211_0[0]),.doutb(w_n2211_0[1]),.din(n2211));
	jspl3 jspl3_w_n2215_0(.douta(w_n2215_0[0]),.doutb(w_n2215_0[1]),.doutc(w_n2215_0[2]),.din(n2215));
	jspl3 jspl3_w_n2218_0(.douta(w_n2218_0[0]),.doutb(w_n2218_0[1]),.doutc(w_n2218_0[2]),.din(n2218));
	jspl jspl_w_n2219_0(.douta(w_n2219_0[0]),.doutb(w_n2219_0[1]),.din(n2219));
	jspl3 jspl3_w_n2223_0(.douta(w_n2223_0[0]),.doutb(w_n2223_0[1]),.doutc(w_n2223_0[2]),.din(n2223));
	jspl3 jspl3_w_n2225_0(.douta(w_n2225_0[0]),.doutb(w_n2225_0[1]),.doutc(w_n2225_0[2]),.din(n2225));
	jspl jspl_w_n2226_0(.douta(w_n2226_0[0]),.doutb(w_n2226_0[1]),.din(n2226));
	jspl3 jspl3_w_n2230_0(.douta(w_n2230_0[0]),.doutb(w_n2230_0[1]),.doutc(w_n2230_0[2]),.din(n2230));
	jspl3 jspl3_w_n2232_0(.douta(w_n2232_0[0]),.doutb(w_n2232_0[1]),.doutc(w_n2232_0[2]),.din(n2232));
	jspl3 jspl3_w_n2235_0(.douta(w_n2235_0[0]),.doutb(w_n2235_0[1]),.doutc(w_n2235_0[2]),.din(n2235));
	jspl jspl_w_n2235_1(.douta(w_n2235_1[0]),.doutb(w_n2235_1[1]),.din(w_n2235_0[0]));
	jspl3 jspl3_w_n2236_0(.douta(w_n2236_0[0]),.doutb(w_n2236_0[1]),.doutc(w_n2236_0[2]),.din(n2236));
	jspl jspl_w_n2238_0(.douta(w_n2238_0[0]),.doutb(w_n2238_0[1]),.din(n2238));
	jspl jspl_w_n2240_0(.douta(w_n2240_0[0]),.doutb(w_n2240_0[1]),.din(n2240));
	jspl jspl_w_n2246_0(.douta(w_n2246_0[0]),.doutb(w_n2246_0[1]),.din(n2246));
	jspl jspl_w_n2247_0(.douta(w_n2247_0[0]),.doutb(w_n2247_0[1]),.din(n2247));
	jspl jspl_w_n2249_0(.douta(w_n2249_0[0]),.doutb(w_n2249_0[1]),.din(n2249));
	jspl3 jspl3_w_n2252_0(.douta(w_n2252_0[0]),.doutb(w_n2252_0[1]),.doutc(w_n2252_0[2]),.din(n2252));
	jspl jspl_w_n2252_1(.douta(w_n2252_1[0]),.doutb(w_n2252_1[1]),.din(w_n2252_0[0]));
	jspl jspl_w_n2253_0(.douta(w_n2253_0[0]),.doutb(w_n2253_0[1]),.din(n2253));
	jspl3 jspl3_w_n2254_0(.douta(w_n2254_0[0]),.doutb(w_n2254_0[1]),.doutc(w_n2254_0[2]),.din(n2254));
	jspl jspl_w_n2255_0(.douta(w_n2255_0[0]),.doutb(w_n2255_0[1]),.din(n2255));
	jspl3 jspl3_w_n2257_0(.douta(w_n2257_0[0]),.doutb(w_n2257_0[1]),.doutc(w_n2257_0[2]),.din(n2257));
	jspl jspl_w_n2258_0(.douta(w_n2258_0[0]),.doutb(w_n2258_0[1]),.din(n2258));
	jspl3 jspl3_w_n2263_0(.douta(w_n2263_0[0]),.doutb(w_n2263_0[1]),.doutc(w_n2263_0[2]),.din(n2263));
	jspl jspl_w_n2263_1(.douta(w_n2263_1[0]),.doutb(w_n2263_1[1]),.din(w_n2263_0[0]));
	jspl jspl_w_n2285_0(.douta(w_n2285_0[0]),.doutb(w_n2285_0[1]),.din(n2285));
	jspl jspl_w_n2321_0(.douta(w_n2321_0[0]),.doutb(w_n2321_0[1]),.din(n2321));
	jspl jspl_w_n2339_0(.douta(w_n2339_0[0]),.doutb(w_n2339_0[1]),.din(n2339));
	jspl jspl_w_n2342_0(.douta(w_n2342_0[0]),.doutb(w_n2342_0[1]),.din(n2342));
	jspl jspl_w_n2343_0(.douta(w_n2343_0[0]),.doutb(w_n2343_0[1]),.din(n2343));
	jspl3 jspl3_w_n2345_0(.douta(w_n2345_0[0]),.doutb(w_n2345_0[1]),.doutc(w_n2345_0[2]),.din(n2345));
	jspl3 jspl3_w_n2345_1(.douta(w_n2345_1[0]),.doutb(w_n2345_1[1]),.doutc(w_n2345_1[2]),.din(w_n2345_0[0]));
	jspl3 jspl3_w_n2345_2(.douta(w_n2345_2[0]),.doutb(w_n2345_2[1]),.doutc(w_n2345_2[2]),.din(w_n2345_0[1]));
	jspl3 jspl3_w_n2345_3(.douta(w_n2345_3[0]),.doutb(w_n2345_3[1]),.doutc(w_n2345_3[2]),.din(w_n2345_0[2]));
	jspl3 jspl3_w_n2345_4(.douta(w_n2345_4[0]),.doutb(w_n2345_4[1]),.doutc(w_n2345_4[2]),.din(w_n2345_1[0]));
	jspl3 jspl3_w_n2345_5(.douta(w_n2345_5[0]),.doutb(w_n2345_5[1]),.doutc(w_n2345_5[2]),.din(w_n2345_1[1]));
	jspl3 jspl3_w_n2345_6(.douta(w_n2345_6[0]),.doutb(w_n2345_6[1]),.doutc(w_n2345_6[2]),.din(w_n2345_1[2]));
	jspl3 jspl3_w_n2345_7(.douta(w_n2345_7[0]),.doutb(w_n2345_7[1]),.doutc(w_n2345_7[2]),.din(w_n2345_2[0]));
	jspl3 jspl3_w_n2345_8(.douta(w_n2345_8[0]),.doutb(w_n2345_8[1]),.doutc(w_n2345_8[2]),.din(w_n2345_2[1]));
	jspl3 jspl3_w_n2345_9(.douta(w_n2345_9[0]),.doutb(w_n2345_9[1]),.doutc(w_n2345_9[2]),.din(w_n2345_2[2]));
	jspl3 jspl3_w_n2345_10(.douta(w_n2345_10[0]),.doutb(w_n2345_10[1]),.doutc(w_n2345_10[2]),.din(w_n2345_3[0]));
	jspl3 jspl3_w_n2345_11(.douta(w_n2345_11[0]),.doutb(w_n2345_11[1]),.doutc(w_n2345_11[2]),.din(w_n2345_3[1]));
	jspl3 jspl3_w_n2345_12(.douta(w_n2345_12[0]),.doutb(w_n2345_12[1]),.doutc(w_n2345_12[2]),.din(w_n2345_3[2]));
	jspl3 jspl3_w_n2345_13(.douta(w_n2345_13[0]),.doutb(w_n2345_13[1]),.doutc(w_n2345_13[2]),.din(w_n2345_4[0]));
	jspl3 jspl3_w_n2345_14(.douta(w_n2345_14[0]),.doutb(w_n2345_14[1]),.doutc(w_n2345_14[2]),.din(w_n2345_4[1]));
	jspl3 jspl3_w_n2345_15(.douta(w_n2345_15[0]),.doutb(w_n2345_15[1]),.doutc(w_n2345_15[2]),.din(w_n2345_4[2]));
	jspl3 jspl3_w_n2345_16(.douta(w_n2345_16[0]),.doutb(w_n2345_16[1]),.doutc(w_n2345_16[2]),.din(w_n2345_5[0]));
	jspl3 jspl3_w_n2345_17(.douta(w_n2345_17[0]),.doutb(w_n2345_17[1]),.doutc(w_n2345_17[2]),.din(w_n2345_5[1]));
	jspl3 jspl3_w_n2345_18(.douta(w_n2345_18[0]),.doutb(w_n2345_18[1]),.doutc(w_n2345_18[2]),.din(w_n2345_5[2]));
	jspl3 jspl3_w_n2345_19(.douta(w_n2345_19[0]),.doutb(w_n2345_19[1]),.doutc(w_n2345_19[2]),.din(w_n2345_6[0]));
	jspl3 jspl3_w_n2345_20(.douta(w_n2345_20[0]),.doutb(w_n2345_20[1]),.doutc(w_n2345_20[2]),.din(w_n2345_6[1]));
	jspl3 jspl3_w_n2345_21(.douta(w_n2345_21[0]),.doutb(w_n2345_21[1]),.doutc(w_n2345_21[2]),.din(w_n2345_6[2]));
	jspl3 jspl3_w_n2345_22(.douta(w_n2345_22[0]),.doutb(w_n2345_22[1]),.doutc(w_n2345_22[2]),.din(w_n2345_7[0]));
	jspl3 jspl3_w_n2345_23(.douta(w_n2345_23[0]),.doutb(w_n2345_23[1]),.doutc(w_n2345_23[2]),.din(w_n2345_7[1]));
	jspl3 jspl3_w_n2345_24(.douta(w_n2345_24[0]),.doutb(w_n2345_24[1]),.doutc(w_n2345_24[2]),.din(w_n2345_7[2]));
	jspl3 jspl3_w_n2345_25(.douta(w_n2345_25[0]),.doutb(w_n2345_25[1]),.doutc(w_n2345_25[2]),.din(w_n2345_8[0]));
	jspl3 jspl3_w_n2345_26(.douta(w_n2345_26[0]),.doutb(w_n2345_26[1]),.doutc(w_n2345_26[2]),.din(w_n2345_8[1]));
	jspl3 jspl3_w_n2345_27(.douta(w_n2345_27[0]),.doutb(w_n2345_27[1]),.doutc(w_n2345_27[2]),.din(w_n2345_8[2]));
	jspl3 jspl3_w_n2345_28(.douta(w_n2345_28[0]),.doutb(w_n2345_28[1]),.doutc(w_n2345_28[2]),.din(w_n2345_9[0]));
	jspl3 jspl3_w_n2345_29(.douta(w_n2345_29[0]),.doutb(w_n2345_29[1]),.doutc(w_n2345_29[2]),.din(w_n2345_9[1]));
	jspl3 jspl3_w_n2345_30(.douta(w_n2345_30[0]),.doutb(w_n2345_30[1]),.doutc(w_n2345_30[2]),.din(w_n2345_9[2]));
	jspl3 jspl3_w_n2345_31(.douta(w_n2345_31[0]),.doutb(w_n2345_31[1]),.doutc(w_n2345_31[2]),.din(w_n2345_10[0]));
	jspl3 jspl3_w_n2345_32(.douta(w_n2345_32[0]),.doutb(w_n2345_32[1]),.doutc(w_n2345_32[2]),.din(w_n2345_10[1]));
	jspl3 jspl3_w_n2345_33(.douta(w_n2345_33[0]),.doutb(w_n2345_33[1]),.doutc(w_n2345_33[2]),.din(w_n2345_10[2]));
	jspl3 jspl3_w_n2345_34(.douta(w_n2345_34[0]),.doutb(w_n2345_34[1]),.doutc(w_n2345_34[2]),.din(w_n2345_11[0]));
	jspl3 jspl3_w_n2345_35(.douta(w_n2345_35[0]),.doutb(w_n2345_35[1]),.doutc(w_n2345_35[2]),.din(w_n2345_11[1]));
	jspl3 jspl3_w_n2345_36(.douta(w_n2345_36[0]),.doutb(w_n2345_36[1]),.doutc(w_n2345_36[2]),.din(w_n2345_11[2]));
	jspl3 jspl3_w_n2345_37(.douta(w_n2345_37[0]),.doutb(w_n2345_37[1]),.doutc(w_n2345_37[2]),.din(w_n2345_12[0]));
	jspl3 jspl3_w_n2345_38(.douta(w_n2345_38[0]),.doutb(w_n2345_38[1]),.doutc(w_n2345_38[2]),.din(w_n2345_12[1]));
	jspl3 jspl3_w_n2345_39(.douta(w_n2345_39[0]),.doutb(w_n2345_39[1]),.doutc(w_n2345_39[2]),.din(w_n2345_12[2]));
	jspl3 jspl3_w_n2345_40(.douta(w_n2345_40[0]),.doutb(w_n2345_40[1]),.doutc(w_n2345_40[2]),.din(w_n2345_13[0]));
	jspl3 jspl3_w_n2345_41(.douta(w_n2345_41[0]),.doutb(w_n2345_41[1]),.doutc(w_n2345_41[2]),.din(w_n2345_13[1]));
	jspl3 jspl3_w_n2345_42(.douta(w_n2345_42[0]),.doutb(w_n2345_42[1]),.doutc(w_n2345_42[2]),.din(w_n2345_13[2]));
	jspl3 jspl3_w_n2345_43(.douta(w_n2345_43[0]),.doutb(w_n2345_43[1]),.doutc(w_n2345_43[2]),.din(w_n2345_14[0]));
	jspl3 jspl3_w_n2345_44(.douta(w_n2345_44[0]),.doutb(w_n2345_44[1]),.doutc(w_n2345_44[2]),.din(w_n2345_14[1]));
	jspl3 jspl3_w_n2345_45(.douta(w_n2345_45[0]),.doutb(w_n2345_45[1]),.doutc(w_n2345_45[2]),.din(w_n2345_14[2]));
	jspl3 jspl3_w_n2345_46(.douta(w_n2345_46[0]),.doutb(w_n2345_46[1]),.doutc(w_n2345_46[2]),.din(w_n2345_15[0]));
	jspl3 jspl3_w_n2345_47(.douta(w_n2345_47[0]),.doutb(w_n2345_47[1]),.doutc(w_n2345_47[2]),.din(w_n2345_15[1]));
	jspl3 jspl3_w_n2345_48(.douta(w_n2345_48[0]),.doutb(w_n2345_48[1]),.doutc(w_n2345_48[2]),.din(w_n2345_15[2]));
	jspl3 jspl3_w_n2345_49(.douta(w_n2345_49[0]),.doutb(w_n2345_49[1]),.doutc(w_n2345_49[2]),.din(w_n2345_16[0]));
	jspl3 jspl3_w_n2345_50(.douta(w_n2345_50[0]),.doutb(w_n2345_50[1]),.doutc(w_n2345_50[2]),.din(w_n2345_16[1]));
	jspl3 jspl3_w_n2345_51(.douta(w_n2345_51[0]),.doutb(w_n2345_51[1]),.doutc(w_n2345_51[2]),.din(w_n2345_16[2]));
	jspl3 jspl3_w_n2345_52(.douta(w_n2345_52[0]),.doutb(w_n2345_52[1]),.doutc(w_n2345_52[2]),.din(w_n2345_17[0]));
	jspl3 jspl3_w_n2345_53(.douta(w_n2345_53[0]),.doutb(w_n2345_53[1]),.doutc(w_n2345_53[2]),.din(w_n2345_17[1]));
	jspl3 jspl3_w_n2345_54(.douta(w_n2345_54[0]),.doutb(w_n2345_54[1]),.doutc(w_n2345_54[2]),.din(w_n2345_17[2]));
	jspl3 jspl3_w_n2345_55(.douta(w_n2345_55[0]),.doutb(w_n2345_55[1]),.doutc(w_n2345_55[2]),.din(w_n2345_18[0]));
	jspl3 jspl3_w_n2345_56(.douta(w_n2345_56[0]),.doutb(w_n2345_56[1]),.doutc(w_n2345_56[2]),.din(w_n2345_18[1]));
	jspl3 jspl3_w_n2345_57(.douta(w_n2345_57[0]),.doutb(w_n2345_57[1]),.doutc(w_n2345_57[2]),.din(w_n2345_18[2]));
	jspl3 jspl3_w_n2349_0(.douta(w_n2349_0[0]),.doutb(w_n2349_0[1]),.doutc(w_n2349_0[2]),.din(n2349));
	jspl jspl_w_n2350_0(.douta(w_n2350_0[0]),.doutb(w_n2350_0[1]),.din(n2350));
	jspl jspl_w_n2352_0(.douta(w_n2352_0[0]),.doutb(w_n2352_0[1]),.din(n2352));
	jspl jspl_w_n2357_0(.douta(w_n2357_0[0]),.doutb(w_n2357_0[1]),.din(n2357));
	jspl jspl_w_n2358_0(.douta(w_n2358_0[0]),.doutb(w_n2358_0[1]),.din(n2358));
	jspl3 jspl3_w_n2360_0(.douta(w_n2360_0[0]),.doutb(w_n2360_0[1]),.doutc(w_n2360_0[2]),.din(n2360));
	jspl jspl_w_n2361_0(.douta(w_n2361_0[0]),.doutb(w_n2361_0[1]),.din(n2361));
	jspl jspl_w_n2365_0(.douta(w_n2365_0[0]),.doutb(w_n2365_0[1]),.din(n2365));
	jspl3 jspl3_w_n2367_0(.douta(w_n2367_0[0]),.doutb(w_n2367_0[1]),.doutc(w_n2367_0[2]),.din(n2367));
	jspl jspl_w_n2368_0(.douta(w_n2368_0[0]),.doutb(w_n2368_0[1]),.din(n2368));
	jspl jspl_w_n2372_0(.douta(w_n2372_0[0]),.doutb(w_n2372_0[1]),.din(n2372));
	jspl jspl_w_n2373_0(.douta(w_n2373_0[0]),.doutb(w_n2373_0[1]),.din(n2373));
	jspl3 jspl3_w_n2375_0(.douta(w_n2375_0[0]),.doutb(w_n2375_0[1]),.doutc(w_n2375_0[2]),.din(n2375));
	jspl jspl_w_n2376_0(.douta(w_n2376_0[0]),.doutb(w_n2376_0[1]),.din(n2376));
	jspl jspl_w_n2380_0(.douta(w_n2380_0[0]),.doutb(w_n2380_0[1]),.din(n2380));
	jspl3 jspl3_w_n2382_0(.douta(w_n2382_0[0]),.doutb(w_n2382_0[1]),.doutc(w_n2382_0[2]),.din(n2382));
	jspl jspl_w_n2383_0(.douta(w_n2383_0[0]),.doutb(w_n2383_0[1]),.din(n2383));
	jspl jspl_w_n2387_0(.douta(w_n2387_0[0]),.doutb(w_n2387_0[1]),.din(n2387));
	jspl jspl_w_n2388_0(.douta(w_n2388_0[0]),.doutb(w_n2388_0[1]),.din(n2388));
	jspl3 jspl3_w_n2390_0(.douta(w_n2390_0[0]),.doutb(w_n2390_0[1]),.doutc(w_n2390_0[2]),.din(n2390));
	jspl jspl_w_n2391_0(.douta(w_n2391_0[0]),.doutb(w_n2391_0[1]),.din(n2391));
	jspl jspl_w_n2395_0(.douta(w_n2395_0[0]),.doutb(w_n2395_0[1]),.din(n2395));
	jspl3 jspl3_w_n2397_0(.douta(w_n2397_0[0]),.doutb(w_n2397_0[1]),.doutc(w_n2397_0[2]),.din(n2397));
	jspl jspl_w_n2398_0(.douta(w_n2398_0[0]),.doutb(w_n2398_0[1]),.din(n2398));
	jspl jspl_w_n2402_0(.douta(w_n2402_0[0]),.doutb(w_n2402_0[1]),.din(n2402));
	jspl jspl_w_n2403_0(.douta(w_n2403_0[0]),.doutb(w_n2403_0[1]),.din(n2403));
	jspl3 jspl3_w_n2405_0(.douta(w_n2405_0[0]),.doutb(w_n2405_0[1]),.doutc(w_n2405_0[2]),.din(n2405));
	jspl jspl_w_n2406_0(.douta(w_n2406_0[0]),.doutb(w_n2406_0[1]),.din(n2406));
	jspl jspl_w_n2410_0(.douta(w_n2410_0[0]),.doutb(w_n2410_0[1]),.din(n2410));
	jspl jspl_w_n2411_0(.douta(w_n2411_0[0]),.doutb(w_n2411_0[1]),.din(n2411));
	jspl3 jspl3_w_n2413_0(.douta(w_n2413_0[0]),.doutb(w_n2413_0[1]),.doutc(w_n2413_0[2]),.din(n2413));
	jspl jspl_w_n2414_0(.douta(w_n2414_0[0]),.doutb(w_n2414_0[1]),.din(n2414));
	jspl jspl_w_n2418_0(.douta(w_n2418_0[0]),.doutb(w_n2418_0[1]),.din(n2418));
	jspl3 jspl3_w_n2420_0(.douta(w_n2420_0[0]),.doutb(w_n2420_0[1]),.doutc(w_n2420_0[2]),.din(n2420));
	jspl jspl_w_n2421_0(.douta(w_n2421_0[0]),.doutb(w_n2421_0[1]),.din(n2421));
	jspl jspl_w_n2425_0(.douta(w_n2425_0[0]),.doutb(w_n2425_0[1]),.din(n2425));
	jspl3 jspl3_w_n2427_0(.douta(w_n2427_0[0]),.doutb(w_n2427_0[1]),.doutc(w_n2427_0[2]),.din(n2427));
	jspl jspl_w_n2428_0(.douta(w_n2428_0[0]),.doutb(w_n2428_0[1]),.din(n2428));
	jspl jspl_w_n2432_0(.douta(w_n2432_0[0]),.doutb(w_n2432_0[1]),.din(n2432));
	jspl jspl_w_n2433_0(.douta(w_n2433_0[0]),.doutb(w_n2433_0[1]),.din(n2433));
	jspl3 jspl3_w_n2435_0(.douta(w_n2435_0[0]),.doutb(w_n2435_0[1]),.doutc(w_n2435_0[2]),.din(n2435));
	jspl jspl_w_n2436_0(.douta(w_n2436_0[0]),.doutb(w_n2436_0[1]),.din(n2436));
	jspl jspl_w_n2440_0(.douta(w_n2440_0[0]),.doutb(w_n2440_0[1]),.din(n2440));
	jspl3 jspl3_w_n2442_0(.douta(w_n2442_0[0]),.doutb(w_n2442_0[1]),.doutc(w_n2442_0[2]),.din(n2442));
	jspl jspl_w_n2443_0(.douta(w_n2443_0[0]),.doutb(w_n2443_0[1]),.din(n2443));
	jspl jspl_w_n2447_0(.douta(w_n2447_0[0]),.doutb(w_n2447_0[1]),.din(n2447));
	jspl3 jspl3_w_n2449_0(.douta(w_n2449_0[0]),.doutb(w_n2449_0[1]),.doutc(w_n2449_0[2]),.din(n2449));
	jspl jspl_w_n2450_0(.douta(w_n2450_0[0]),.doutb(w_n2450_0[1]),.din(n2450));
	jspl jspl_w_n2454_0(.douta(w_n2454_0[0]),.doutb(w_n2454_0[1]),.din(n2454));
	jspl3 jspl3_w_n2456_0(.douta(w_n2456_0[0]),.doutb(w_n2456_0[1]),.doutc(w_n2456_0[2]),.din(n2456));
	jspl jspl_w_n2457_0(.douta(w_n2457_0[0]),.doutb(w_n2457_0[1]),.din(n2457));
	jspl3 jspl3_w_n2461_0(.douta(w_n2461_0[0]),.doutb(w_n2461_0[1]),.doutc(w_n2461_0[2]),.din(n2461));
	jspl jspl_w_n2464_0(.douta(w_n2464_0[0]),.doutb(w_n2464_0[1]),.din(n2464));
	jspl jspl_w_n2467_0(.douta(w_n2467_0[0]),.doutb(w_n2467_0[1]),.din(n2467));
	jspl jspl_w_n2468_0(.douta(w_n2468_0[0]),.doutb(w_n2468_0[1]),.din(n2468));
	jspl3 jspl3_w_n2469_0(.douta(w_n2469_0[0]),.doutb(w_n2469_0[1]),.doutc(w_n2469_0[2]),.din(n2469));
	jspl jspl_w_n2469_1(.douta(w_n2469_1[0]),.doutb(w_n2469_1[1]),.din(w_n2469_0[0]));
	jspl3 jspl3_w_n2470_0(.douta(w_n2470_0[0]),.doutb(w_n2470_0[1]),.doutc(w_n2470_0[2]),.din(n2470));
	jspl jspl_w_n2474_0(.douta(w_n2474_0[0]),.doutb(w_n2474_0[1]),.din(n2474));
	jspl jspl_w_n2475_0(.douta(w_n2475_0[0]),.doutb(w_n2475_0[1]),.din(n2475));
	jspl jspl_w_n2476_0(.douta(w_n2476_0[0]),.doutb(w_n2476_0[1]),.din(n2476));
	jspl jspl_w_n2499_0(.douta(w_n2499_0[0]),.doutb(w_n2499_0[1]),.din(n2499));
	jspl jspl_w_n2506_0(.douta(w_n2506_0[0]),.doutb(w_n2506_0[1]),.din(n2506));
	jspl jspl_w_n2513_0(.douta(w_n2513_0[0]),.doutb(w_n2513_0[1]),.din(n2513));
	jspl jspl_w_n2520_0(.douta(w_n2520_0[0]),.doutb(w_n2520_0[1]),.din(n2520));
	jspl jspl_w_n2530_0(.douta(w_n2530_0[0]),.doutb(w_n2530_0[1]),.din(n2530));
	jspl jspl_w_n2534_0(.douta(w_n2534_0[0]),.doutb(w_n2534_0[1]),.din(n2534));
	jspl jspl_w_n2541_0(.douta(w_n2541_0[0]),.doutb(w_n2541_0[1]),.din(n2541));
	jspl jspl_w_n2545_0(.douta(w_n2545_0[0]),.doutb(w_n2545_0[1]),.din(n2545));
	jspl jspl_w_n2549_0(.douta(w_n2549_0[0]),.doutb(w_n2549_0[1]),.din(n2549));
	jspl jspl_w_n2554_0(.douta(w_n2554_0[0]),.doutb(w_n2554_0[1]),.din(n2554));
	jspl jspl_w_n2555_0(.douta(w_n2555_0[0]),.doutb(w_n2555_0[1]),.din(n2555));
	jspl jspl_w_n2558_0(.douta(w_n2558_0[0]),.doutb(w_n2558_0[1]),.din(n2558));
	jspl jspl_w_n2559_0(.douta(w_n2559_0[0]),.doutb(w_n2559_0[1]),.din(n2559));
	jspl jspl_w_n2561_0(.douta(w_n2561_0[0]),.doutb(w_n2561_0[1]),.din(n2561));
	jspl jspl_w_n2565_0(.douta(w_n2565_0[0]),.doutb(w_n2565_0[1]),.din(n2565));
	jspl jspl_w_n2571_0(.douta(w_n2571_0[0]),.doutb(w_n2571_0[1]),.din(n2571));
	jspl3 jspl3_w_n2572_0(.douta(w_n2572_0[0]),.doutb(w_n2572_0[1]),.doutc(w_n2572_0[2]),.din(n2572));
	jspl3 jspl3_w_n2572_1(.douta(w_n2572_1[0]),.doutb(w_n2572_1[1]),.doutc(w_n2572_1[2]),.din(w_n2572_0[0]));
	jspl3 jspl3_w_n2572_2(.douta(w_n2572_2[0]),.doutb(w_n2572_2[1]),.doutc(w_n2572_2[2]),.din(w_n2572_0[1]));
	jspl3 jspl3_w_n2572_3(.douta(w_n2572_3[0]),.doutb(w_n2572_3[1]),.doutc(w_n2572_3[2]),.din(w_n2572_0[2]));
	jspl3 jspl3_w_n2572_4(.douta(w_n2572_4[0]),.doutb(w_n2572_4[1]),.doutc(w_n2572_4[2]),.din(w_n2572_1[0]));
	jspl3 jspl3_w_n2572_5(.douta(w_n2572_5[0]),.doutb(w_n2572_5[1]),.doutc(w_n2572_5[2]),.din(w_n2572_1[1]));
	jspl3 jspl3_w_n2572_6(.douta(w_n2572_6[0]),.doutb(w_n2572_6[1]),.doutc(w_n2572_6[2]),.din(w_n2572_1[2]));
	jspl3 jspl3_w_n2572_7(.douta(w_n2572_7[0]),.doutb(w_n2572_7[1]),.doutc(w_n2572_7[2]),.din(w_n2572_2[0]));
	jspl3 jspl3_w_n2572_8(.douta(w_n2572_8[0]),.doutb(w_n2572_8[1]),.doutc(w_n2572_8[2]),.din(w_n2572_2[1]));
	jspl3 jspl3_w_n2572_9(.douta(w_n2572_9[0]),.doutb(w_n2572_9[1]),.doutc(w_n2572_9[2]),.din(w_n2572_2[2]));
	jspl3 jspl3_w_n2572_10(.douta(w_n2572_10[0]),.doutb(w_n2572_10[1]),.doutc(w_n2572_10[2]),.din(w_n2572_3[0]));
	jspl3 jspl3_w_n2572_11(.douta(w_n2572_11[0]),.doutb(w_n2572_11[1]),.doutc(w_n2572_11[2]),.din(w_n2572_3[1]));
	jspl3 jspl3_w_n2572_12(.douta(w_n2572_12[0]),.doutb(w_n2572_12[1]),.doutc(w_n2572_12[2]),.din(w_n2572_3[2]));
	jspl3 jspl3_w_n2572_13(.douta(w_n2572_13[0]),.doutb(w_n2572_13[1]),.doutc(w_n2572_13[2]),.din(w_n2572_4[0]));
	jspl3 jspl3_w_n2572_14(.douta(w_n2572_14[0]),.doutb(w_n2572_14[1]),.doutc(w_n2572_14[2]),.din(w_n2572_4[1]));
	jspl3 jspl3_w_n2572_15(.douta(w_n2572_15[0]),.doutb(w_n2572_15[1]),.doutc(w_n2572_15[2]),.din(w_n2572_4[2]));
	jspl3 jspl3_w_n2572_16(.douta(w_n2572_16[0]),.doutb(w_n2572_16[1]),.doutc(w_n2572_16[2]),.din(w_n2572_5[0]));
	jspl3 jspl3_w_n2572_17(.douta(w_n2572_17[0]),.doutb(w_n2572_17[1]),.doutc(w_n2572_17[2]),.din(w_n2572_5[1]));
	jspl3 jspl3_w_n2572_18(.douta(w_n2572_18[0]),.doutb(w_n2572_18[1]),.doutc(w_n2572_18[2]),.din(w_n2572_5[2]));
	jspl3 jspl3_w_n2572_19(.douta(w_n2572_19[0]),.doutb(w_n2572_19[1]),.doutc(w_n2572_19[2]),.din(w_n2572_6[0]));
	jspl3 jspl3_w_n2572_20(.douta(w_n2572_20[0]),.doutb(w_n2572_20[1]),.doutc(w_n2572_20[2]),.din(w_n2572_6[1]));
	jspl3 jspl3_w_n2572_21(.douta(w_n2572_21[0]),.doutb(w_n2572_21[1]),.doutc(w_n2572_21[2]),.din(w_n2572_6[2]));
	jspl3 jspl3_w_n2572_22(.douta(w_n2572_22[0]),.doutb(w_n2572_22[1]),.doutc(w_n2572_22[2]),.din(w_n2572_7[0]));
	jspl3 jspl3_w_n2572_23(.douta(w_n2572_23[0]),.doutb(w_n2572_23[1]),.doutc(w_n2572_23[2]),.din(w_n2572_7[1]));
	jspl3 jspl3_w_n2572_24(.douta(w_n2572_24[0]),.doutb(w_n2572_24[1]),.doutc(w_n2572_24[2]),.din(w_n2572_7[2]));
	jspl3 jspl3_w_n2572_25(.douta(w_n2572_25[0]),.doutb(w_n2572_25[1]),.doutc(w_n2572_25[2]),.din(w_n2572_8[0]));
	jspl3 jspl3_w_n2572_26(.douta(w_n2572_26[0]),.doutb(w_n2572_26[1]),.doutc(w_n2572_26[2]),.din(w_n2572_8[1]));
	jspl3 jspl3_w_n2572_27(.douta(w_n2572_27[0]),.doutb(w_n2572_27[1]),.doutc(w_n2572_27[2]),.din(w_n2572_8[2]));
	jspl3 jspl3_w_n2572_28(.douta(w_n2572_28[0]),.doutb(w_n2572_28[1]),.doutc(w_n2572_28[2]),.din(w_n2572_9[0]));
	jspl3 jspl3_w_n2572_29(.douta(w_n2572_29[0]),.doutb(w_n2572_29[1]),.doutc(w_n2572_29[2]),.din(w_n2572_9[1]));
	jspl3 jspl3_w_n2572_30(.douta(w_n2572_30[0]),.doutb(w_n2572_30[1]),.doutc(w_n2572_30[2]),.din(w_n2572_9[2]));
	jspl3 jspl3_w_n2572_31(.douta(w_n2572_31[0]),.doutb(w_n2572_31[1]),.doutc(w_n2572_31[2]),.din(w_n2572_10[0]));
	jspl3 jspl3_w_n2572_32(.douta(w_n2572_32[0]),.doutb(w_n2572_32[1]),.doutc(w_n2572_32[2]),.din(w_n2572_10[1]));
	jspl3 jspl3_w_n2572_33(.douta(w_n2572_33[0]),.doutb(w_n2572_33[1]),.doutc(w_n2572_33[2]),.din(w_n2572_10[2]));
	jspl3 jspl3_w_n2572_34(.douta(w_n2572_34[0]),.doutb(w_n2572_34[1]),.doutc(w_n2572_34[2]),.din(w_n2572_11[0]));
	jspl3 jspl3_w_n2572_35(.douta(w_n2572_35[0]),.doutb(w_n2572_35[1]),.doutc(w_n2572_35[2]),.din(w_n2572_11[1]));
	jspl3 jspl3_w_n2572_36(.douta(w_n2572_36[0]),.doutb(w_n2572_36[1]),.doutc(w_n2572_36[2]),.din(w_n2572_11[2]));
	jspl3 jspl3_w_n2572_37(.douta(w_n2572_37[0]),.doutb(w_n2572_37[1]),.doutc(w_n2572_37[2]),.din(w_n2572_12[0]));
	jspl3 jspl3_w_n2572_38(.douta(w_n2572_38[0]),.doutb(w_n2572_38[1]),.doutc(w_n2572_38[2]),.din(w_n2572_12[1]));
	jspl3 jspl3_w_n2572_39(.douta(w_n2572_39[0]),.doutb(w_n2572_39[1]),.doutc(w_n2572_39[2]),.din(w_n2572_12[2]));
	jspl3 jspl3_w_n2572_40(.douta(w_n2572_40[0]),.doutb(w_n2572_40[1]),.doutc(w_n2572_40[2]),.din(w_n2572_13[0]));
	jspl3 jspl3_w_n2572_41(.douta(w_n2572_41[0]),.doutb(w_n2572_41[1]),.doutc(w_n2572_41[2]),.din(w_n2572_13[1]));
	jspl3 jspl3_w_n2572_42(.douta(w_n2572_42[0]),.doutb(w_n2572_42[1]),.doutc(w_n2572_42[2]),.din(w_n2572_13[2]));
	jspl3 jspl3_w_n2572_43(.douta(w_n2572_43[0]),.doutb(w_n2572_43[1]),.doutc(w_n2572_43[2]),.din(w_n2572_14[0]));
	jspl3 jspl3_w_n2572_44(.douta(w_n2572_44[0]),.doutb(w_n2572_44[1]),.doutc(w_n2572_44[2]),.din(w_n2572_14[1]));
	jspl3 jspl3_w_n2572_45(.douta(w_n2572_45[0]),.doutb(w_n2572_45[1]),.doutc(w_n2572_45[2]),.din(w_n2572_14[2]));
	jspl3 jspl3_w_n2572_46(.douta(w_n2572_46[0]),.doutb(w_n2572_46[1]),.doutc(w_n2572_46[2]),.din(w_n2572_15[0]));
	jspl3 jspl3_w_n2572_47(.douta(w_n2572_47[0]),.doutb(w_n2572_47[1]),.doutc(w_n2572_47[2]),.din(w_n2572_15[1]));
	jspl3 jspl3_w_n2572_48(.douta(w_n2572_48[0]),.doutb(w_n2572_48[1]),.doutc(w_n2572_48[2]),.din(w_n2572_15[2]));
	jspl3 jspl3_w_n2572_49(.douta(w_n2572_49[0]),.doutb(w_n2572_49[1]),.doutc(w_n2572_49[2]),.din(w_n2572_16[0]));
	jspl3 jspl3_w_n2572_50(.douta(w_n2572_50[0]),.doutb(w_n2572_50[1]),.doutc(w_n2572_50[2]),.din(w_n2572_16[1]));
	jspl3 jspl3_w_n2572_51(.douta(w_n2572_51[0]),.doutb(w_n2572_51[1]),.doutc(w_n2572_51[2]),.din(w_n2572_16[2]));
	jspl3 jspl3_w_n2572_52(.douta(w_n2572_52[0]),.doutb(w_n2572_52[1]),.doutc(w_n2572_52[2]),.din(w_n2572_17[0]));
	jspl3 jspl3_w_n2572_53(.douta(w_n2572_53[0]),.doutb(w_n2572_53[1]),.doutc(w_n2572_53[2]),.din(w_n2572_17[1]));
	jspl3 jspl3_w_n2572_54(.douta(w_n2572_54[0]),.doutb(w_n2572_54[1]),.doutc(w_n2572_54[2]),.din(w_n2572_17[2]));
	jspl3 jspl3_w_n2572_55(.douta(w_n2572_55[0]),.doutb(w_n2572_55[1]),.doutc(w_n2572_55[2]),.din(w_n2572_18[0]));
	jspl3 jspl3_w_n2572_56(.douta(w_n2572_56[0]),.doutb(w_n2572_56[1]),.doutc(w_n2572_56[2]),.din(w_n2572_18[1]));
	jspl3 jspl3_w_n2572_57(.douta(w_n2572_57[0]),.doutb(w_n2572_57[1]),.doutc(w_n2572_57[2]),.din(w_n2572_18[2]));
	jspl3 jspl3_w_n2572_58(.douta(w_n2572_58[0]),.doutb(w_n2572_58[1]),.doutc(w_n2572_58[2]),.din(w_n2572_19[0]));
	jspl3 jspl3_w_n2572_59(.douta(w_n2572_59[0]),.doutb(w_n2572_59[1]),.doutc(w_n2572_59[2]),.din(w_n2572_19[1]));
	jspl3 jspl3_w_n2572_60(.douta(w_n2572_60[0]),.doutb(w_n2572_60[1]),.doutc(w_n2572_60[2]),.din(w_n2572_19[2]));
	jspl3 jspl3_w_n2572_61(.douta(w_n2572_61[0]),.doutb(w_n2572_61[1]),.doutc(w_n2572_61[2]),.din(w_n2572_20[0]));
	jspl3 jspl3_w_n2572_62(.douta(w_n2572_62[0]),.doutb(w_n2572_62[1]),.doutc(w_n2572_62[2]),.din(w_n2572_20[1]));
	jspl jspl_w_n2572_63(.douta(w_n2572_63[0]),.doutb(w_n2572_63[1]),.din(w_n2572_20[2]));
	jspl jspl_w_n2575_0(.douta(w_n2575_0[0]),.doutb(w_n2575_0[1]),.din(n2575));
	jspl3 jspl3_w_n2576_0(.douta(w_n2576_0[0]),.doutb(w_n2576_0[1]),.doutc(w_n2576_0[2]),.din(n2576));
	jspl3 jspl3_w_n2578_0(.douta(w_n2578_0[0]),.doutb(w_n2578_0[1]),.doutc(w_n2578_0[2]),.din(n2578));
	jspl3 jspl3_w_n2578_1(.douta(w_n2578_1[0]),.doutb(w_n2578_1[1]),.doutc(w_n2578_1[2]),.din(w_n2578_0[0]));
	jspl jspl_w_n2579_0(.douta(w_n2579_0[0]),.doutb(w_n2579_0[1]),.din(n2579));
	jspl3 jspl3_w_n2580_0(.douta(w_n2580_0[0]),.doutb(w_n2580_0[1]),.doutc(w_n2580_0[2]),.din(n2580));
	jspl jspl_w_n2581_0(.douta(w_n2581_0[0]),.doutb(w_n2581_0[1]),.din(n2581));
	jspl3 jspl3_w_n2583_0(.douta(w_n2583_0[0]),.doutb(w_n2583_0[1]),.doutc(w_n2583_0[2]),.din(n2583));
	jspl jspl_w_n2584_0(.douta(w_n2584_0[0]),.doutb(w_n2584_0[1]),.din(n2584));
	jspl3 jspl3_w_n2591_0(.douta(w_n2591_0[0]),.doutb(w_n2591_0[1]),.doutc(w_n2591_0[2]),.din(n2591));
	jspl jspl_w_n2592_0(.douta(w_n2592_0[0]),.doutb(w_n2592_0[1]),.din(n2592));
	jspl jspl_w_n2595_0(.douta(w_n2595_0[0]),.doutb(w_n2595_0[1]),.din(n2595));
	jspl3 jspl3_w_n2600_0(.douta(w_n2600_0[0]),.doutb(w_n2600_0[1]),.doutc(w_n2600_0[2]),.din(n2600));
	jspl3 jspl3_w_n2602_0(.douta(w_n2602_0[0]),.doutb(w_n2602_0[1]),.doutc(w_n2602_0[2]),.din(n2602));
	jspl jspl_w_n2603_0(.douta(w_n2603_0[0]),.doutb(w_n2603_0[1]),.din(n2603));
	jspl3 jspl3_w_n2607_0(.douta(w_n2607_0[0]),.doutb(w_n2607_0[1]),.doutc(w_n2607_0[2]),.din(n2607));
	jspl3 jspl3_w_n2610_0(.douta(w_n2610_0[0]),.doutb(w_n2610_0[1]),.doutc(w_n2610_0[2]),.din(n2610));
	jspl jspl_w_n2611_0(.douta(w_n2611_0[0]),.doutb(w_n2611_0[1]),.din(n2611));
	jspl3 jspl3_w_n2615_0(.douta(w_n2615_0[0]),.doutb(w_n2615_0[1]),.doutc(w_n2615_0[2]),.din(n2615));
	jspl3 jspl3_w_n2617_0(.douta(w_n2617_0[0]),.doutb(w_n2617_0[1]),.doutc(w_n2617_0[2]),.din(n2617));
	jspl jspl_w_n2618_0(.douta(w_n2618_0[0]),.doutb(w_n2618_0[1]),.din(n2618));
	jspl3 jspl3_w_n2622_0(.douta(w_n2622_0[0]),.doutb(w_n2622_0[1]),.doutc(w_n2622_0[2]),.din(n2622));
	jspl3 jspl3_w_n2625_0(.douta(w_n2625_0[0]),.doutb(w_n2625_0[1]),.doutc(w_n2625_0[2]),.din(n2625));
	jspl jspl_w_n2626_0(.douta(w_n2626_0[0]),.doutb(w_n2626_0[1]),.din(n2626));
	jspl3 jspl3_w_n2630_0(.douta(w_n2630_0[0]),.doutb(w_n2630_0[1]),.doutc(w_n2630_0[2]),.din(n2630));
	jspl3 jspl3_w_n2632_0(.douta(w_n2632_0[0]),.doutb(w_n2632_0[1]),.doutc(w_n2632_0[2]),.din(n2632));
	jspl jspl_w_n2633_0(.douta(w_n2633_0[0]),.doutb(w_n2633_0[1]),.din(n2633));
	jspl3 jspl3_w_n2637_0(.douta(w_n2637_0[0]),.doutb(w_n2637_0[1]),.doutc(w_n2637_0[2]),.din(n2637));
	jspl3 jspl3_w_n2640_0(.douta(w_n2640_0[0]),.doutb(w_n2640_0[1]),.doutc(w_n2640_0[2]),.din(n2640));
	jspl jspl_w_n2641_0(.douta(w_n2641_0[0]),.doutb(w_n2641_0[1]),.din(n2641));
	jspl3 jspl3_w_n2645_0(.douta(w_n2645_0[0]),.doutb(w_n2645_0[1]),.doutc(w_n2645_0[2]),.din(n2645));
	jspl3 jspl3_w_n2647_0(.douta(w_n2647_0[0]),.doutb(w_n2647_0[1]),.doutc(w_n2647_0[2]),.din(n2647));
	jspl jspl_w_n2648_0(.douta(w_n2648_0[0]),.doutb(w_n2648_0[1]),.din(n2648));
	jspl3 jspl3_w_n2652_0(.douta(w_n2652_0[0]),.doutb(w_n2652_0[1]),.doutc(w_n2652_0[2]),.din(n2652));
	jspl3 jspl3_w_n2655_0(.douta(w_n2655_0[0]),.doutb(w_n2655_0[1]),.doutc(w_n2655_0[2]),.din(n2655));
	jspl jspl_w_n2656_0(.douta(w_n2656_0[0]),.doutb(w_n2656_0[1]),.din(n2656));
	jspl3 jspl3_w_n2660_0(.douta(w_n2660_0[0]),.doutb(w_n2660_0[1]),.doutc(w_n2660_0[2]),.din(n2660));
	jspl3 jspl3_w_n2662_0(.douta(w_n2662_0[0]),.doutb(w_n2662_0[1]),.doutc(w_n2662_0[2]),.din(n2662));
	jspl jspl_w_n2663_0(.douta(w_n2663_0[0]),.doutb(w_n2663_0[1]),.din(n2663));
	jspl3 jspl3_w_n2667_0(.douta(w_n2667_0[0]),.doutb(w_n2667_0[1]),.doutc(w_n2667_0[2]),.din(n2667));
	jspl3 jspl3_w_n2669_0(.douta(w_n2669_0[0]),.doutb(w_n2669_0[1]),.doutc(w_n2669_0[2]),.din(n2669));
	jspl jspl_w_n2670_0(.douta(w_n2670_0[0]),.doutb(w_n2670_0[1]),.din(n2670));
	jspl3 jspl3_w_n2674_0(.douta(w_n2674_0[0]),.doutb(w_n2674_0[1]),.doutc(w_n2674_0[2]),.din(n2674));
	jspl3 jspl3_w_n2677_0(.douta(w_n2677_0[0]),.doutb(w_n2677_0[1]),.doutc(w_n2677_0[2]),.din(n2677));
	jspl jspl_w_n2678_0(.douta(w_n2678_0[0]),.doutb(w_n2678_0[1]),.din(n2678));
	jspl3 jspl3_w_n2682_0(.douta(w_n2682_0[0]),.doutb(w_n2682_0[1]),.doutc(w_n2682_0[2]),.din(n2682));
	jspl3 jspl3_w_n2685_0(.douta(w_n2685_0[0]),.doutb(w_n2685_0[1]),.doutc(w_n2685_0[2]),.din(n2685));
	jspl jspl_w_n2686_0(.douta(w_n2686_0[0]),.doutb(w_n2686_0[1]),.din(n2686));
	jspl3 jspl3_w_n2690_0(.douta(w_n2690_0[0]),.doutb(w_n2690_0[1]),.doutc(w_n2690_0[2]),.din(n2690));
	jspl3 jspl3_w_n2692_0(.douta(w_n2692_0[0]),.doutb(w_n2692_0[1]),.doutc(w_n2692_0[2]),.din(n2692));
	jspl jspl_w_n2693_0(.douta(w_n2693_0[0]),.doutb(w_n2693_0[1]),.din(n2693));
	jspl3 jspl3_w_n2697_0(.douta(w_n2697_0[0]),.doutb(w_n2697_0[1]),.doutc(w_n2697_0[2]),.din(n2697));
	jspl3 jspl3_w_n2700_0(.douta(w_n2700_0[0]),.doutb(w_n2700_0[1]),.doutc(w_n2700_0[2]),.din(n2700));
	jspl jspl_w_n2701_0(.douta(w_n2701_0[0]),.doutb(w_n2701_0[1]),.din(n2701));
	jspl3 jspl3_w_n2705_0(.douta(w_n2705_0[0]),.doutb(w_n2705_0[1]),.doutc(w_n2705_0[2]),.din(n2705));
	jspl3 jspl3_w_n2708_0(.douta(w_n2708_0[0]),.doutb(w_n2708_0[1]),.doutc(w_n2708_0[2]),.din(n2708));
	jspl jspl_w_n2709_0(.douta(w_n2709_0[0]),.doutb(w_n2709_0[1]),.din(n2709));
	jspl jspl_w_n2713_0(.douta(w_n2713_0[0]),.doutb(w_n2713_0[1]),.din(n2713));
	jspl jspl_w_n2714_0(.douta(w_n2714_0[0]),.doutb(w_n2714_0[1]),.din(n2714));
	jspl3 jspl3_w_n2716_0(.douta(w_n2716_0[0]),.doutb(w_n2716_0[1]),.doutc(w_n2716_0[2]),.din(n2716));
	jspl3 jspl3_w_n2717_0(.douta(w_n2717_0[0]),.doutb(w_n2717_0[1]),.doutc(w_n2717_0[2]),.din(n2717));
	jspl jspl_w_n2719_0(.douta(w_n2719_0[0]),.doutb(w_n2719_0[1]),.din(n2719));
	jspl jspl_w_n2720_0(.douta(w_n2720_0[0]),.doutb(w_n2720_0[1]),.din(n2720));
	jspl jspl_w_n2727_0(.douta(w_n2727_0[0]),.doutb(w_n2727_0[1]),.din(n2727));
	jspl jspl_w_n2728_0(.douta(w_n2728_0[0]),.doutb(w_n2728_0[1]),.din(n2728));
	jspl jspl_w_n2730_0(.douta(w_n2730_0[0]),.doutb(w_n2730_0[1]),.din(n2730));
	jspl3 jspl3_w_n2734_0(.douta(w_n2734_0[0]),.doutb(w_n2734_0[1]),.doutc(w_n2734_0[2]),.din(n2734));
	jspl jspl_w_n2734_1(.douta(w_n2734_1[0]),.doutb(w_n2734_1[1]),.din(w_n2734_0[0]));
	jspl jspl_w_n2735_0(.douta(w_n2735_0[0]),.doutb(w_n2735_0[1]),.din(n2735));
	jspl3 jspl3_w_n2736_0(.douta(w_n2736_0[0]),.doutb(w_n2736_0[1]),.doutc(w_n2736_0[2]),.din(n2736));
	jspl jspl_w_n2737_0(.douta(w_n2737_0[0]),.doutb(w_n2737_0[1]),.din(n2737));
	jspl3 jspl3_w_n2738_0(.douta(w_n2738_0[0]),.doutb(w_n2738_0[1]),.doutc(w_n2738_0[2]),.din(n2738));
	jspl jspl_w_n2739_0(.douta(w_n2739_0[0]),.doutb(w_n2739_0[1]),.din(n2739));
	jspl3 jspl3_w_n2744_0(.douta(w_n2744_0[0]),.doutb(w_n2744_0[1]),.doutc(w_n2744_0[2]),.din(n2744));
	jspl jspl_w_n2744_1(.douta(w_n2744_1[0]),.doutb(w_n2744_1[1]),.din(w_n2744_0[0]));
	jspl jspl_w_n2769_0(.douta(w_n2769_0[0]),.doutb(w_n2769_0[1]),.din(n2769));
	jspl jspl_w_n2827_0(.douta(w_n2827_0[0]),.doutb(w_n2827_0[1]),.din(n2827));
	jspl jspl_w_n2830_0(.douta(w_n2830_0[0]),.doutb(w_n2830_0[1]),.din(n2830));
	jspl jspl_w_n2831_0(.douta(w_n2831_0[0]),.doutb(w_n2831_0[1]),.din(n2831));
	jspl3 jspl3_w_n2833_0(.douta(w_n2833_0[0]),.doutb(w_n2833_0[1]),.doutc(w_n2833_0[2]),.din(n2833));
	jspl3 jspl3_w_n2833_1(.douta(w_n2833_1[0]),.doutb(w_n2833_1[1]),.doutc(w_n2833_1[2]),.din(w_n2833_0[0]));
	jspl3 jspl3_w_n2833_2(.douta(w_n2833_2[0]),.doutb(w_n2833_2[1]),.doutc(w_n2833_2[2]),.din(w_n2833_0[1]));
	jspl3 jspl3_w_n2833_3(.douta(w_n2833_3[0]),.doutb(w_n2833_3[1]),.doutc(w_n2833_3[2]),.din(w_n2833_0[2]));
	jspl3 jspl3_w_n2833_4(.douta(w_n2833_4[0]),.doutb(w_n2833_4[1]),.doutc(w_n2833_4[2]),.din(w_n2833_1[0]));
	jspl3 jspl3_w_n2833_5(.douta(w_n2833_5[0]),.doutb(w_n2833_5[1]),.doutc(w_n2833_5[2]),.din(w_n2833_1[1]));
	jspl3 jspl3_w_n2833_6(.douta(w_n2833_6[0]),.doutb(w_n2833_6[1]),.doutc(w_n2833_6[2]),.din(w_n2833_1[2]));
	jspl3 jspl3_w_n2833_7(.douta(w_n2833_7[0]),.doutb(w_n2833_7[1]),.doutc(w_n2833_7[2]),.din(w_n2833_2[0]));
	jspl3 jspl3_w_n2833_8(.douta(w_n2833_8[0]),.doutb(w_n2833_8[1]),.doutc(w_n2833_8[2]),.din(w_n2833_2[1]));
	jspl3 jspl3_w_n2833_9(.douta(w_n2833_9[0]),.doutb(w_n2833_9[1]),.doutc(w_n2833_9[2]),.din(w_n2833_2[2]));
	jspl3 jspl3_w_n2833_10(.douta(w_n2833_10[0]),.doutb(w_n2833_10[1]),.doutc(w_n2833_10[2]),.din(w_n2833_3[0]));
	jspl3 jspl3_w_n2833_11(.douta(w_n2833_11[0]),.doutb(w_n2833_11[1]),.doutc(w_n2833_11[2]),.din(w_n2833_3[1]));
	jspl3 jspl3_w_n2833_12(.douta(w_n2833_12[0]),.doutb(w_n2833_12[1]),.doutc(w_n2833_12[2]),.din(w_n2833_3[2]));
	jspl3 jspl3_w_n2833_13(.douta(w_n2833_13[0]),.doutb(w_n2833_13[1]),.doutc(w_n2833_13[2]),.din(w_n2833_4[0]));
	jspl3 jspl3_w_n2833_14(.douta(w_n2833_14[0]),.doutb(w_n2833_14[1]),.doutc(w_n2833_14[2]),.din(w_n2833_4[1]));
	jspl3 jspl3_w_n2833_15(.douta(w_n2833_15[0]),.doutb(w_n2833_15[1]),.doutc(w_n2833_15[2]),.din(w_n2833_4[2]));
	jspl3 jspl3_w_n2833_16(.douta(w_n2833_16[0]),.doutb(w_n2833_16[1]),.doutc(w_n2833_16[2]),.din(w_n2833_5[0]));
	jspl3 jspl3_w_n2833_17(.douta(w_n2833_17[0]),.doutb(w_n2833_17[1]),.doutc(w_n2833_17[2]),.din(w_n2833_5[1]));
	jspl3 jspl3_w_n2833_18(.douta(w_n2833_18[0]),.doutb(w_n2833_18[1]),.doutc(w_n2833_18[2]),.din(w_n2833_5[2]));
	jspl3 jspl3_w_n2833_19(.douta(w_n2833_19[0]),.doutb(w_n2833_19[1]),.doutc(w_n2833_19[2]),.din(w_n2833_6[0]));
	jspl3 jspl3_w_n2833_20(.douta(w_n2833_20[0]),.doutb(w_n2833_20[1]),.doutc(w_n2833_20[2]),.din(w_n2833_6[1]));
	jspl3 jspl3_w_n2833_21(.douta(w_n2833_21[0]),.doutb(w_n2833_21[1]),.doutc(w_n2833_21[2]),.din(w_n2833_6[2]));
	jspl3 jspl3_w_n2833_22(.douta(w_n2833_22[0]),.doutb(w_n2833_22[1]),.doutc(w_n2833_22[2]),.din(w_n2833_7[0]));
	jspl3 jspl3_w_n2833_23(.douta(w_n2833_23[0]),.doutb(w_n2833_23[1]),.doutc(w_n2833_23[2]),.din(w_n2833_7[1]));
	jspl3 jspl3_w_n2833_24(.douta(w_n2833_24[0]),.doutb(w_n2833_24[1]),.doutc(w_n2833_24[2]),.din(w_n2833_7[2]));
	jspl3 jspl3_w_n2833_25(.douta(w_n2833_25[0]),.doutb(w_n2833_25[1]),.doutc(w_n2833_25[2]),.din(w_n2833_8[0]));
	jspl3 jspl3_w_n2833_26(.douta(w_n2833_26[0]),.doutb(w_n2833_26[1]),.doutc(w_n2833_26[2]),.din(w_n2833_8[1]));
	jspl3 jspl3_w_n2833_27(.douta(w_n2833_27[0]),.doutb(w_n2833_27[1]),.doutc(w_n2833_27[2]),.din(w_n2833_8[2]));
	jspl3 jspl3_w_n2833_28(.douta(w_n2833_28[0]),.doutb(w_n2833_28[1]),.doutc(w_n2833_28[2]),.din(w_n2833_9[0]));
	jspl3 jspl3_w_n2833_29(.douta(w_n2833_29[0]),.doutb(w_n2833_29[1]),.doutc(w_n2833_29[2]),.din(w_n2833_9[1]));
	jspl3 jspl3_w_n2833_30(.douta(w_n2833_30[0]),.doutb(w_n2833_30[1]),.doutc(w_n2833_30[2]),.din(w_n2833_9[2]));
	jspl3 jspl3_w_n2833_31(.douta(w_n2833_31[0]),.doutb(w_n2833_31[1]),.doutc(w_n2833_31[2]),.din(w_n2833_10[0]));
	jspl3 jspl3_w_n2833_32(.douta(w_n2833_32[0]),.doutb(w_n2833_32[1]),.doutc(w_n2833_32[2]),.din(w_n2833_10[1]));
	jspl3 jspl3_w_n2833_33(.douta(w_n2833_33[0]),.doutb(w_n2833_33[1]),.doutc(w_n2833_33[2]),.din(w_n2833_10[2]));
	jspl3 jspl3_w_n2833_34(.douta(w_n2833_34[0]),.doutb(w_n2833_34[1]),.doutc(w_n2833_34[2]),.din(w_n2833_11[0]));
	jspl3 jspl3_w_n2833_35(.douta(w_n2833_35[0]),.doutb(w_n2833_35[1]),.doutc(w_n2833_35[2]),.din(w_n2833_11[1]));
	jspl3 jspl3_w_n2833_36(.douta(w_n2833_36[0]),.doutb(w_n2833_36[1]),.doutc(w_n2833_36[2]),.din(w_n2833_11[2]));
	jspl3 jspl3_w_n2833_37(.douta(w_n2833_37[0]),.doutb(w_n2833_37[1]),.doutc(w_n2833_37[2]),.din(w_n2833_12[0]));
	jspl3 jspl3_w_n2833_38(.douta(w_n2833_38[0]),.doutb(w_n2833_38[1]),.doutc(w_n2833_38[2]),.din(w_n2833_12[1]));
	jspl3 jspl3_w_n2833_39(.douta(w_n2833_39[0]),.doutb(w_n2833_39[1]),.doutc(w_n2833_39[2]),.din(w_n2833_12[2]));
	jspl3 jspl3_w_n2833_40(.douta(w_n2833_40[0]),.doutb(w_n2833_40[1]),.doutc(w_n2833_40[2]),.din(w_n2833_13[0]));
	jspl3 jspl3_w_n2833_41(.douta(w_n2833_41[0]),.doutb(w_n2833_41[1]),.doutc(w_n2833_41[2]),.din(w_n2833_13[1]));
	jspl3 jspl3_w_n2833_42(.douta(w_n2833_42[0]),.doutb(w_n2833_42[1]),.doutc(w_n2833_42[2]),.din(w_n2833_13[2]));
	jspl3 jspl3_w_n2833_43(.douta(w_n2833_43[0]),.doutb(w_n2833_43[1]),.doutc(w_n2833_43[2]),.din(w_n2833_14[0]));
	jspl3 jspl3_w_n2833_44(.douta(w_n2833_44[0]),.doutb(w_n2833_44[1]),.doutc(w_n2833_44[2]),.din(w_n2833_14[1]));
	jspl3 jspl3_w_n2833_45(.douta(w_n2833_45[0]),.doutb(w_n2833_45[1]),.doutc(w_n2833_45[2]),.din(w_n2833_14[2]));
	jspl3 jspl3_w_n2833_46(.douta(w_n2833_46[0]),.doutb(w_n2833_46[1]),.doutc(w_n2833_46[2]),.din(w_n2833_15[0]));
	jspl3 jspl3_w_n2833_47(.douta(w_n2833_47[0]),.doutb(w_n2833_47[1]),.doutc(w_n2833_47[2]),.din(w_n2833_15[1]));
	jspl3 jspl3_w_n2833_48(.douta(w_n2833_48[0]),.doutb(w_n2833_48[1]),.doutc(w_n2833_48[2]),.din(w_n2833_15[2]));
	jspl3 jspl3_w_n2833_49(.douta(w_n2833_49[0]),.doutb(w_n2833_49[1]),.doutc(w_n2833_49[2]),.din(w_n2833_16[0]));
	jspl3 jspl3_w_n2833_50(.douta(w_n2833_50[0]),.doutb(w_n2833_50[1]),.doutc(w_n2833_50[2]),.din(w_n2833_16[1]));
	jspl3 jspl3_w_n2833_51(.douta(w_n2833_51[0]),.doutb(w_n2833_51[1]),.doutc(w_n2833_51[2]),.din(w_n2833_16[2]));
	jspl3 jspl3_w_n2833_52(.douta(w_n2833_52[0]),.doutb(w_n2833_52[1]),.doutc(w_n2833_52[2]),.din(w_n2833_17[0]));
	jspl3 jspl3_w_n2833_53(.douta(w_n2833_53[0]),.doutb(w_n2833_53[1]),.doutc(w_n2833_53[2]),.din(w_n2833_17[1]));
	jspl3 jspl3_w_n2833_54(.douta(w_n2833_54[0]),.doutb(w_n2833_54[1]),.doutc(w_n2833_54[2]),.din(w_n2833_17[2]));
	jspl jspl_w_n2833_55(.douta(w_n2833_55[0]),.doutb(w_n2833_55[1]),.din(w_n2833_18[0]));
	jspl jspl_w_n2835_0(.douta(w_n2835_0[0]),.doutb(w_n2835_0[1]),.din(n2835));
	jspl3 jspl3_w_n2837_0(.douta(w_n2837_0[0]),.doutb(w_n2837_0[1]),.doutc(w_n2837_0[2]),.din(n2837));
	jspl jspl_w_n2838_0(.douta(w_n2838_0[0]),.doutb(w_n2838_0[1]),.din(n2838));
	jspl jspl_w_n2840_0(.douta(w_n2840_0[0]),.doutb(w_n2840_0[1]),.din(n2840));
	jspl jspl_w_n2845_0(.douta(w_n2845_0[0]),.doutb(w_n2845_0[1]),.din(n2845));
	jspl jspl_w_n2846_0(.douta(w_n2846_0[0]),.doutb(w_n2846_0[1]),.din(n2846));
	jspl3 jspl3_w_n2848_0(.douta(w_n2848_0[0]),.doutb(w_n2848_0[1]),.doutc(w_n2848_0[2]),.din(n2848));
	jspl jspl_w_n2849_0(.douta(w_n2849_0[0]),.doutb(w_n2849_0[1]),.din(n2849));
	jspl jspl_w_n2853_0(.douta(w_n2853_0[0]),.doutb(w_n2853_0[1]),.din(n2853));
	jspl3 jspl3_w_n2855_0(.douta(w_n2855_0[0]),.doutb(w_n2855_0[1]),.doutc(w_n2855_0[2]),.din(n2855));
	jspl jspl_w_n2856_0(.douta(w_n2856_0[0]),.doutb(w_n2856_0[1]),.din(n2856));
	jspl jspl_w_n2860_0(.douta(w_n2860_0[0]),.doutb(w_n2860_0[1]),.din(n2860));
	jspl jspl_w_n2861_0(.douta(w_n2861_0[0]),.doutb(w_n2861_0[1]),.din(n2861));
	jspl3 jspl3_w_n2863_0(.douta(w_n2863_0[0]),.doutb(w_n2863_0[1]),.doutc(w_n2863_0[2]),.din(n2863));
	jspl jspl_w_n2864_0(.douta(w_n2864_0[0]),.doutb(w_n2864_0[1]),.din(n2864));
	jspl jspl_w_n2868_0(.douta(w_n2868_0[0]),.doutb(w_n2868_0[1]),.din(n2868));
	jspl3 jspl3_w_n2870_0(.douta(w_n2870_0[0]),.doutb(w_n2870_0[1]),.doutc(w_n2870_0[2]),.din(n2870));
	jspl jspl_w_n2871_0(.douta(w_n2871_0[0]),.doutb(w_n2871_0[1]),.din(n2871));
	jspl jspl_w_n2875_0(.douta(w_n2875_0[0]),.doutb(w_n2875_0[1]),.din(n2875));
	jspl jspl_w_n2876_0(.douta(w_n2876_0[0]),.doutb(w_n2876_0[1]),.din(n2876));
	jspl3 jspl3_w_n2878_0(.douta(w_n2878_0[0]),.doutb(w_n2878_0[1]),.doutc(w_n2878_0[2]),.din(n2878));
	jspl jspl_w_n2879_0(.douta(w_n2879_0[0]),.doutb(w_n2879_0[1]),.din(n2879));
	jspl jspl_w_n2883_0(.douta(w_n2883_0[0]),.doutb(w_n2883_0[1]),.din(n2883));
	jspl3 jspl3_w_n2885_0(.douta(w_n2885_0[0]),.doutb(w_n2885_0[1]),.doutc(w_n2885_0[2]),.din(n2885));
	jspl jspl_w_n2886_0(.douta(w_n2886_0[0]),.doutb(w_n2886_0[1]),.din(n2886));
	jspl jspl_w_n2890_0(.douta(w_n2890_0[0]),.doutb(w_n2890_0[1]),.din(n2890));
	jspl jspl_w_n2891_0(.douta(w_n2891_0[0]),.doutb(w_n2891_0[1]),.din(n2891));
	jspl3 jspl3_w_n2893_0(.douta(w_n2893_0[0]),.doutb(w_n2893_0[1]),.doutc(w_n2893_0[2]),.din(n2893));
	jspl jspl_w_n2894_0(.douta(w_n2894_0[0]),.doutb(w_n2894_0[1]),.din(n2894));
	jspl jspl_w_n2898_0(.douta(w_n2898_0[0]),.doutb(w_n2898_0[1]),.din(n2898));
	jspl3 jspl3_w_n2900_0(.douta(w_n2900_0[0]),.doutb(w_n2900_0[1]),.doutc(w_n2900_0[2]),.din(n2900));
	jspl jspl_w_n2901_0(.douta(w_n2901_0[0]),.doutb(w_n2901_0[1]),.din(n2901));
	jspl jspl_w_n2905_0(.douta(w_n2905_0[0]),.doutb(w_n2905_0[1]),.din(n2905));
	jspl jspl_w_n2906_0(.douta(w_n2906_0[0]),.doutb(w_n2906_0[1]),.din(n2906));
	jspl3 jspl3_w_n2908_0(.douta(w_n2908_0[0]),.doutb(w_n2908_0[1]),.doutc(w_n2908_0[2]),.din(n2908));
	jspl jspl_w_n2909_0(.douta(w_n2909_0[0]),.doutb(w_n2909_0[1]),.din(n2909));
	jspl jspl_w_n2913_0(.douta(w_n2913_0[0]),.doutb(w_n2913_0[1]),.din(n2913));
	jspl3 jspl3_w_n2915_0(.douta(w_n2915_0[0]),.doutb(w_n2915_0[1]),.doutc(w_n2915_0[2]),.din(n2915));
	jspl jspl_w_n2916_0(.douta(w_n2916_0[0]),.doutb(w_n2916_0[1]),.din(n2916));
	jspl jspl_w_n2920_0(.douta(w_n2920_0[0]),.doutb(w_n2920_0[1]),.din(n2920));
	jspl jspl_w_n2921_0(.douta(w_n2921_0[0]),.doutb(w_n2921_0[1]),.din(n2921));
	jspl3 jspl3_w_n2923_0(.douta(w_n2923_0[0]),.doutb(w_n2923_0[1]),.doutc(w_n2923_0[2]),.din(n2923));
	jspl jspl_w_n2924_0(.douta(w_n2924_0[0]),.doutb(w_n2924_0[1]),.din(n2924));
	jspl jspl_w_n2928_0(.douta(w_n2928_0[0]),.doutb(w_n2928_0[1]),.din(n2928));
	jspl jspl_w_n2929_0(.douta(w_n2929_0[0]),.doutb(w_n2929_0[1]),.din(n2929));
	jspl3 jspl3_w_n2931_0(.douta(w_n2931_0[0]),.doutb(w_n2931_0[1]),.doutc(w_n2931_0[2]),.din(n2931));
	jspl jspl_w_n2932_0(.douta(w_n2932_0[0]),.doutb(w_n2932_0[1]),.din(n2932));
	jspl jspl_w_n2936_0(.douta(w_n2936_0[0]),.doutb(w_n2936_0[1]),.din(n2936));
	jspl3 jspl3_w_n2938_0(.douta(w_n2938_0[0]),.doutb(w_n2938_0[1]),.doutc(w_n2938_0[2]),.din(n2938));
	jspl jspl_w_n2939_0(.douta(w_n2939_0[0]),.doutb(w_n2939_0[1]),.din(n2939));
	jspl jspl_w_n2943_0(.douta(w_n2943_0[0]),.doutb(w_n2943_0[1]),.din(n2943));
	jspl3 jspl3_w_n2945_0(.douta(w_n2945_0[0]),.doutb(w_n2945_0[1]),.doutc(w_n2945_0[2]),.din(n2945));
	jspl jspl_w_n2946_0(.douta(w_n2946_0[0]),.doutb(w_n2946_0[1]),.din(n2946));
	jspl jspl_w_n2950_0(.douta(w_n2950_0[0]),.doutb(w_n2950_0[1]),.din(n2950));
	jspl jspl_w_n2951_0(.douta(w_n2951_0[0]),.doutb(w_n2951_0[1]),.din(n2951));
	jspl3 jspl3_w_n2953_0(.douta(w_n2953_0[0]),.doutb(w_n2953_0[1]),.doutc(w_n2953_0[2]),.din(n2953));
	jspl jspl_w_n2954_0(.douta(w_n2954_0[0]),.doutb(w_n2954_0[1]),.din(n2954));
	jspl jspl_w_n2958_0(.douta(w_n2958_0[0]),.doutb(w_n2958_0[1]),.din(n2958));
	jspl3 jspl3_w_n2960_0(.douta(w_n2960_0[0]),.doutb(w_n2960_0[1]),.doutc(w_n2960_0[2]),.din(n2960));
	jspl jspl_w_n2961_0(.douta(w_n2961_0[0]),.doutb(w_n2961_0[1]),.din(n2961));
	jspl3 jspl3_w_n2965_0(.douta(w_n2965_0[0]),.doutb(w_n2965_0[1]),.doutc(w_n2965_0[2]),.din(n2965));
	jspl jspl_w_n2967_0(.douta(w_n2967_0[0]),.doutb(w_n2967_0[1]),.din(n2967));
	jspl3 jspl3_w_n2970_0(.douta(w_n2970_0[0]),.doutb(w_n2970_0[1]),.doutc(w_n2970_0[2]),.din(n2970));
	jspl jspl_w_n2971_0(.douta(w_n2971_0[0]),.doutb(w_n2971_0[1]),.din(n2971));
	jspl3 jspl3_w_n2972_0(.douta(w_n2972_0[0]),.doutb(w_n2972_0[1]),.doutc(w_n2972_0[2]),.din(n2972));
	jspl3 jspl3_w_n2973_0(.douta(w_n2973_0[0]),.doutb(w_n2973_0[1]),.doutc(w_n2973_0[2]),.din(n2973));
	jspl jspl_w_n2977_0(.douta(w_n2977_0[0]),.doutb(w_n2977_0[1]),.din(n2977));
	jspl jspl_w_n2978_0(.douta(w_n2978_0[0]),.doutb(w_n2978_0[1]),.din(n2978));
	jspl jspl_w_n2979_0(.douta(w_n2979_0[0]),.doutb(w_n2979_0[1]),.din(n2979));
	jspl jspl_w_n3011_0(.douta(w_n3011_0[0]),.doutb(w_n3011_0[1]),.din(n3011));
	jspl jspl_w_n3018_0(.douta(w_n3018_0[0]),.doutb(w_n3018_0[1]),.din(n3018));
	jspl jspl_w_n3025_0(.douta(w_n3025_0[0]),.doutb(w_n3025_0[1]),.din(n3025));
	jspl jspl_w_n3032_0(.douta(w_n3032_0[0]),.doutb(w_n3032_0[1]),.din(n3032));
	jspl jspl_w_n3039_0(.douta(w_n3039_0[0]),.doutb(w_n3039_0[1]),.din(n3039));
	jspl jspl_w_n3049_0(.douta(w_n3049_0[0]),.doutb(w_n3049_0[1]),.din(n3049));
	jspl jspl_w_n3053_0(.douta(w_n3053_0[0]),.doutb(w_n3053_0[1]),.din(n3053));
	jspl jspl_w_n3060_0(.douta(w_n3060_0[0]),.doutb(w_n3060_0[1]),.din(n3060));
	jspl jspl_w_n3066_0(.douta(w_n3066_0[0]),.doutb(w_n3066_0[1]),.din(n3066));
	jspl jspl_w_n3067_0(.douta(w_n3067_0[0]),.doutb(w_n3067_0[1]),.din(n3067));
	jspl jspl_w_n3070_0(.douta(w_n3070_0[0]),.doutb(w_n3070_0[1]),.din(n3070));
	jspl jspl_w_n3071_0(.douta(w_n3071_0[0]),.doutb(w_n3071_0[1]),.din(n3071));
	jspl jspl_w_n3073_0(.douta(w_n3073_0[0]),.doutb(w_n3073_0[1]),.din(n3073));
	jspl3 jspl3_w_n3075_0(.douta(w_n3075_0[0]),.doutb(w_n3075_0[1]),.doutc(w_n3075_0[2]),.din(n3075));
	jspl3 jspl3_w_n3075_1(.douta(w_n3075_1[0]),.doutb(w_n3075_1[1]),.doutc(w_n3075_1[2]),.din(w_n3075_0[0]));
	jspl jspl_w_n3076_0(.douta(w_n3076_0[0]),.doutb(w_n3076_0[1]),.din(n3076));
	jspl3 jspl3_w_n3077_0(.douta(w_n3077_0[0]),.doutb(w_n3077_0[1]),.doutc(w_n3077_0[2]),.din(n3077));
	jspl jspl_w_n3078_0(.douta(w_n3078_0[0]),.doutb(w_n3078_0[1]),.din(n3078));
	jspl jspl_w_n3082_0(.douta(w_n3082_0[0]),.doutb(w_n3082_0[1]),.din(n3082));
	jspl jspl_w_n3088_0(.douta(w_n3088_0[0]),.doutb(w_n3088_0[1]),.din(n3088));
	jspl3 jspl3_w_n3089_0(.douta(w_n3089_0[0]),.doutb(w_n3089_0[1]),.doutc(w_n3089_0[2]),.din(n3089));
	jspl3 jspl3_w_n3089_1(.douta(w_n3089_1[0]),.doutb(w_n3089_1[1]),.doutc(w_n3089_1[2]),.din(w_n3089_0[0]));
	jspl3 jspl3_w_n3089_2(.douta(w_n3089_2[0]),.doutb(w_n3089_2[1]),.doutc(w_n3089_2[2]),.din(w_n3089_0[1]));
	jspl3 jspl3_w_n3089_3(.douta(w_n3089_3[0]),.doutb(w_n3089_3[1]),.doutc(w_n3089_3[2]),.din(w_n3089_0[2]));
	jspl3 jspl3_w_n3089_4(.douta(w_n3089_4[0]),.doutb(w_n3089_4[1]),.doutc(w_n3089_4[2]),.din(w_n3089_1[0]));
	jspl3 jspl3_w_n3089_5(.douta(w_n3089_5[0]),.doutb(w_n3089_5[1]),.doutc(w_n3089_5[2]),.din(w_n3089_1[1]));
	jspl3 jspl3_w_n3089_6(.douta(w_n3089_6[0]),.doutb(w_n3089_6[1]),.doutc(w_n3089_6[2]),.din(w_n3089_1[2]));
	jspl3 jspl3_w_n3089_7(.douta(w_n3089_7[0]),.doutb(w_n3089_7[1]),.doutc(w_n3089_7[2]),.din(w_n3089_2[0]));
	jspl3 jspl3_w_n3089_8(.douta(w_n3089_8[0]),.doutb(w_n3089_8[1]),.doutc(w_n3089_8[2]),.din(w_n3089_2[1]));
	jspl3 jspl3_w_n3089_9(.douta(w_n3089_9[0]),.doutb(w_n3089_9[1]),.doutc(w_n3089_9[2]),.din(w_n3089_2[2]));
	jspl3 jspl3_w_n3089_10(.douta(w_n3089_10[0]),.doutb(w_n3089_10[1]),.doutc(w_n3089_10[2]),.din(w_n3089_3[0]));
	jspl3 jspl3_w_n3089_11(.douta(w_n3089_11[0]),.doutb(w_n3089_11[1]),.doutc(w_n3089_11[2]),.din(w_n3089_3[1]));
	jspl3 jspl3_w_n3089_12(.douta(w_n3089_12[0]),.doutb(w_n3089_12[1]),.doutc(w_n3089_12[2]),.din(w_n3089_3[2]));
	jspl3 jspl3_w_n3089_13(.douta(w_n3089_13[0]),.doutb(w_n3089_13[1]),.doutc(w_n3089_13[2]),.din(w_n3089_4[0]));
	jspl3 jspl3_w_n3089_14(.douta(w_n3089_14[0]),.doutb(w_n3089_14[1]),.doutc(w_n3089_14[2]),.din(w_n3089_4[1]));
	jspl3 jspl3_w_n3089_15(.douta(w_n3089_15[0]),.doutb(w_n3089_15[1]),.doutc(w_n3089_15[2]),.din(w_n3089_4[2]));
	jspl3 jspl3_w_n3089_16(.douta(w_n3089_16[0]),.doutb(w_n3089_16[1]),.doutc(w_n3089_16[2]),.din(w_n3089_5[0]));
	jspl3 jspl3_w_n3089_17(.douta(w_n3089_17[0]),.doutb(w_n3089_17[1]),.doutc(w_n3089_17[2]),.din(w_n3089_5[1]));
	jspl3 jspl3_w_n3089_18(.douta(w_n3089_18[0]),.doutb(w_n3089_18[1]),.doutc(w_n3089_18[2]),.din(w_n3089_5[2]));
	jspl3 jspl3_w_n3089_19(.douta(w_n3089_19[0]),.doutb(w_n3089_19[1]),.doutc(w_n3089_19[2]),.din(w_n3089_6[0]));
	jspl3 jspl3_w_n3089_20(.douta(w_n3089_20[0]),.doutb(w_n3089_20[1]),.doutc(w_n3089_20[2]),.din(w_n3089_6[1]));
	jspl3 jspl3_w_n3089_21(.douta(w_n3089_21[0]),.doutb(w_n3089_21[1]),.doutc(w_n3089_21[2]),.din(w_n3089_6[2]));
	jspl3 jspl3_w_n3089_22(.douta(w_n3089_22[0]),.doutb(w_n3089_22[1]),.doutc(w_n3089_22[2]),.din(w_n3089_7[0]));
	jspl3 jspl3_w_n3089_23(.douta(w_n3089_23[0]),.doutb(w_n3089_23[1]),.doutc(w_n3089_23[2]),.din(w_n3089_7[1]));
	jspl3 jspl3_w_n3089_24(.douta(w_n3089_24[0]),.doutb(w_n3089_24[1]),.doutc(w_n3089_24[2]),.din(w_n3089_7[2]));
	jspl3 jspl3_w_n3089_25(.douta(w_n3089_25[0]),.doutb(w_n3089_25[1]),.doutc(w_n3089_25[2]),.din(w_n3089_8[0]));
	jspl3 jspl3_w_n3089_26(.douta(w_n3089_26[0]),.doutb(w_n3089_26[1]),.doutc(w_n3089_26[2]),.din(w_n3089_8[1]));
	jspl3 jspl3_w_n3089_27(.douta(w_n3089_27[0]),.doutb(w_n3089_27[1]),.doutc(w_n3089_27[2]),.din(w_n3089_8[2]));
	jspl3 jspl3_w_n3089_28(.douta(w_n3089_28[0]),.doutb(w_n3089_28[1]),.doutc(w_n3089_28[2]),.din(w_n3089_9[0]));
	jspl3 jspl3_w_n3089_29(.douta(w_n3089_29[0]),.doutb(w_n3089_29[1]),.doutc(w_n3089_29[2]),.din(w_n3089_9[1]));
	jspl3 jspl3_w_n3089_30(.douta(w_n3089_30[0]),.doutb(w_n3089_30[1]),.doutc(w_n3089_30[2]),.din(w_n3089_9[2]));
	jspl3 jspl3_w_n3089_31(.douta(w_n3089_31[0]),.doutb(w_n3089_31[1]),.doutc(w_n3089_31[2]),.din(w_n3089_10[0]));
	jspl3 jspl3_w_n3089_32(.douta(w_n3089_32[0]),.doutb(w_n3089_32[1]),.doutc(w_n3089_32[2]),.din(w_n3089_10[1]));
	jspl3 jspl3_w_n3089_33(.douta(w_n3089_33[0]),.doutb(w_n3089_33[1]),.doutc(w_n3089_33[2]),.din(w_n3089_10[2]));
	jspl3 jspl3_w_n3089_34(.douta(w_n3089_34[0]),.doutb(w_n3089_34[1]),.doutc(w_n3089_34[2]),.din(w_n3089_11[0]));
	jspl3 jspl3_w_n3089_35(.douta(w_n3089_35[0]),.doutb(w_n3089_35[1]),.doutc(w_n3089_35[2]),.din(w_n3089_11[1]));
	jspl3 jspl3_w_n3089_36(.douta(w_n3089_36[0]),.doutb(w_n3089_36[1]),.doutc(w_n3089_36[2]),.din(w_n3089_11[2]));
	jspl3 jspl3_w_n3089_37(.douta(w_n3089_37[0]),.doutb(w_n3089_37[1]),.doutc(w_n3089_37[2]),.din(w_n3089_12[0]));
	jspl3 jspl3_w_n3089_38(.douta(w_n3089_38[0]),.doutb(w_n3089_38[1]),.doutc(w_n3089_38[2]),.din(w_n3089_12[1]));
	jspl3 jspl3_w_n3089_39(.douta(w_n3089_39[0]),.doutb(w_n3089_39[1]),.doutc(w_n3089_39[2]),.din(w_n3089_12[2]));
	jspl3 jspl3_w_n3089_40(.douta(w_n3089_40[0]),.doutb(w_n3089_40[1]),.doutc(w_n3089_40[2]),.din(w_n3089_13[0]));
	jspl3 jspl3_w_n3089_41(.douta(w_n3089_41[0]),.doutb(w_n3089_41[1]),.doutc(w_n3089_41[2]),.din(w_n3089_13[1]));
	jspl3 jspl3_w_n3089_42(.douta(w_n3089_42[0]),.doutb(w_n3089_42[1]),.doutc(w_n3089_42[2]),.din(w_n3089_13[2]));
	jspl3 jspl3_w_n3089_43(.douta(w_n3089_43[0]),.doutb(w_n3089_43[1]),.doutc(w_n3089_43[2]),.din(w_n3089_14[0]));
	jspl3 jspl3_w_n3089_44(.douta(w_n3089_44[0]),.doutb(w_n3089_44[1]),.doutc(w_n3089_44[2]),.din(w_n3089_14[1]));
	jspl3 jspl3_w_n3089_45(.douta(w_n3089_45[0]),.doutb(w_n3089_45[1]),.doutc(w_n3089_45[2]),.din(w_n3089_14[2]));
	jspl3 jspl3_w_n3089_46(.douta(w_n3089_46[0]),.doutb(w_n3089_46[1]),.doutc(w_n3089_46[2]),.din(w_n3089_15[0]));
	jspl3 jspl3_w_n3089_47(.douta(w_n3089_47[0]),.doutb(w_n3089_47[1]),.doutc(w_n3089_47[2]),.din(w_n3089_15[1]));
	jspl3 jspl3_w_n3089_48(.douta(w_n3089_48[0]),.doutb(w_n3089_48[1]),.doutc(w_n3089_48[2]),.din(w_n3089_15[2]));
	jspl3 jspl3_w_n3089_49(.douta(w_n3089_49[0]),.doutb(w_n3089_49[1]),.doutc(w_n3089_49[2]),.din(w_n3089_16[0]));
	jspl3 jspl3_w_n3089_50(.douta(w_n3089_50[0]),.doutb(w_n3089_50[1]),.doutc(w_n3089_50[2]),.din(w_n3089_16[1]));
	jspl3 jspl3_w_n3089_51(.douta(w_n3089_51[0]),.doutb(w_n3089_51[1]),.doutc(w_n3089_51[2]),.din(w_n3089_16[2]));
	jspl3 jspl3_w_n3089_52(.douta(w_n3089_52[0]),.doutb(w_n3089_52[1]),.doutc(w_n3089_52[2]),.din(w_n3089_17[0]));
	jspl3 jspl3_w_n3089_53(.douta(w_n3089_53[0]),.doutb(w_n3089_53[1]),.doutc(w_n3089_53[2]),.din(w_n3089_17[1]));
	jspl3 jspl3_w_n3089_54(.douta(w_n3089_54[0]),.doutb(w_n3089_54[1]),.doutc(w_n3089_54[2]),.din(w_n3089_17[2]));
	jspl3 jspl3_w_n3089_55(.douta(w_n3089_55[0]),.doutb(w_n3089_55[1]),.doutc(w_n3089_55[2]),.din(w_n3089_18[0]));
	jspl3 jspl3_w_n3089_56(.douta(w_n3089_56[0]),.doutb(w_n3089_56[1]),.doutc(w_n3089_56[2]),.din(w_n3089_18[1]));
	jspl3 jspl3_w_n3089_57(.douta(w_n3089_57[0]),.doutb(w_n3089_57[1]),.doutc(w_n3089_57[2]),.din(w_n3089_18[2]));
	jspl3 jspl3_w_n3089_58(.douta(w_n3089_58[0]),.doutb(w_n3089_58[1]),.doutc(w_n3089_58[2]),.din(w_n3089_19[0]));
	jspl3 jspl3_w_n3089_59(.douta(w_n3089_59[0]),.doutb(w_n3089_59[1]),.doutc(w_n3089_59[2]),.din(w_n3089_19[1]));
	jspl3 jspl3_w_n3089_60(.douta(w_n3089_60[0]),.doutb(w_n3089_60[1]),.doutc(w_n3089_60[2]),.din(w_n3089_19[2]));
	jspl3 jspl3_w_n3089_61(.douta(w_n3089_61[0]),.doutb(w_n3089_61[1]),.doutc(w_n3089_61[2]),.din(w_n3089_20[0]));
	jspl jspl_w_n3089_62(.douta(w_n3089_62[0]),.doutb(w_n3089_62[1]),.din(w_n3089_20[1]));
	jspl3 jspl3_w_n3091_0(.douta(w_n3091_0[0]),.doutb(w_n3091_0[1]),.doutc(w_n3091_0[2]),.din(n3091));
	jspl jspl_w_n3092_0(.douta(w_n3092_0[0]),.doutb(w_n3092_0[1]),.din(n3092));
	jspl3 jspl3_w_n3099_0(.douta(w_n3099_0[0]),.doutb(w_n3099_0[1]),.doutc(w_n3099_0[2]),.din(n3099));
	jspl jspl_w_n3100_0(.douta(w_n3100_0[0]),.doutb(w_n3100_0[1]),.din(n3100));
	jspl jspl_w_n3103_0(.douta(w_n3103_0[0]),.doutb(w_n3103_0[1]),.din(n3103));
	jspl jspl_w_n3108_0(.douta(w_n3108_0[0]),.doutb(w_n3108_0[1]),.din(n3108));
	jspl3 jspl3_w_n3110_0(.douta(w_n3110_0[0]),.doutb(w_n3110_0[1]),.doutc(w_n3110_0[2]),.din(n3110));
	jspl jspl_w_n3111_0(.douta(w_n3111_0[0]),.doutb(w_n3111_0[1]),.din(n3111));
	jspl3 jspl3_w_n3115_0(.douta(w_n3115_0[0]),.doutb(w_n3115_0[1]),.doutc(w_n3115_0[2]),.din(n3115));
	jspl3 jspl3_w_n3117_0(.douta(w_n3117_0[0]),.doutb(w_n3117_0[1]),.doutc(w_n3117_0[2]),.din(n3117));
	jspl jspl_w_n3118_0(.douta(w_n3118_0[0]),.doutb(w_n3118_0[1]),.din(n3118));
	jspl3 jspl3_w_n3122_0(.douta(w_n3122_0[0]),.doutb(w_n3122_0[1]),.doutc(w_n3122_0[2]),.din(n3122));
	jspl3 jspl3_w_n3124_0(.douta(w_n3124_0[0]),.doutb(w_n3124_0[1]),.doutc(w_n3124_0[2]),.din(n3124));
	jspl jspl_w_n3125_0(.douta(w_n3125_0[0]),.doutb(w_n3125_0[1]),.din(n3125));
	jspl3 jspl3_w_n3129_0(.douta(w_n3129_0[0]),.doutb(w_n3129_0[1]),.doutc(w_n3129_0[2]),.din(n3129));
	jspl3 jspl3_w_n3132_0(.douta(w_n3132_0[0]),.doutb(w_n3132_0[1]),.doutc(w_n3132_0[2]),.din(n3132));
	jspl jspl_w_n3133_0(.douta(w_n3133_0[0]),.doutb(w_n3133_0[1]),.din(n3133));
	jspl3 jspl3_w_n3137_0(.douta(w_n3137_0[0]),.doutb(w_n3137_0[1]),.doutc(w_n3137_0[2]),.din(n3137));
	jspl3 jspl3_w_n3139_0(.douta(w_n3139_0[0]),.doutb(w_n3139_0[1]),.doutc(w_n3139_0[2]),.din(n3139));
	jspl jspl_w_n3140_0(.douta(w_n3140_0[0]),.doutb(w_n3140_0[1]),.din(n3140));
	jspl3 jspl3_w_n3144_0(.douta(w_n3144_0[0]),.doutb(w_n3144_0[1]),.doutc(w_n3144_0[2]),.din(n3144));
	jspl3 jspl3_w_n3147_0(.douta(w_n3147_0[0]),.doutb(w_n3147_0[1]),.doutc(w_n3147_0[2]),.din(n3147));
	jspl jspl_w_n3148_0(.douta(w_n3148_0[0]),.doutb(w_n3148_0[1]),.din(n3148));
	jspl3 jspl3_w_n3152_0(.douta(w_n3152_0[0]),.doutb(w_n3152_0[1]),.doutc(w_n3152_0[2]),.din(n3152));
	jspl3 jspl3_w_n3154_0(.douta(w_n3154_0[0]),.doutb(w_n3154_0[1]),.doutc(w_n3154_0[2]),.din(n3154));
	jspl jspl_w_n3155_0(.douta(w_n3155_0[0]),.doutb(w_n3155_0[1]),.din(n3155));
	jspl3 jspl3_w_n3159_0(.douta(w_n3159_0[0]),.doutb(w_n3159_0[1]),.doutc(w_n3159_0[2]),.din(n3159));
	jspl3 jspl3_w_n3162_0(.douta(w_n3162_0[0]),.doutb(w_n3162_0[1]),.doutc(w_n3162_0[2]),.din(n3162));
	jspl jspl_w_n3163_0(.douta(w_n3163_0[0]),.doutb(w_n3163_0[1]),.din(n3163));
	jspl3 jspl3_w_n3167_0(.douta(w_n3167_0[0]),.doutb(w_n3167_0[1]),.doutc(w_n3167_0[2]),.din(n3167));
	jspl3 jspl3_w_n3169_0(.douta(w_n3169_0[0]),.doutb(w_n3169_0[1]),.doutc(w_n3169_0[2]),.din(n3169));
	jspl jspl_w_n3170_0(.douta(w_n3170_0[0]),.doutb(w_n3170_0[1]),.din(n3170));
	jspl3 jspl3_w_n3174_0(.douta(w_n3174_0[0]),.doutb(w_n3174_0[1]),.doutc(w_n3174_0[2]),.din(n3174));
	jspl3 jspl3_w_n3177_0(.douta(w_n3177_0[0]),.doutb(w_n3177_0[1]),.doutc(w_n3177_0[2]),.din(n3177));
	jspl jspl_w_n3178_0(.douta(w_n3178_0[0]),.doutb(w_n3178_0[1]),.din(n3178));
	jspl3 jspl3_w_n3182_0(.douta(w_n3182_0[0]),.doutb(w_n3182_0[1]),.doutc(w_n3182_0[2]),.din(n3182));
	jspl3 jspl3_w_n3184_0(.douta(w_n3184_0[0]),.doutb(w_n3184_0[1]),.doutc(w_n3184_0[2]),.din(n3184));
	jspl jspl_w_n3185_0(.douta(w_n3185_0[0]),.doutb(w_n3185_0[1]),.din(n3185));
	jspl3 jspl3_w_n3189_0(.douta(w_n3189_0[0]),.doutb(w_n3189_0[1]),.doutc(w_n3189_0[2]),.din(n3189));
	jspl3 jspl3_w_n3192_0(.douta(w_n3192_0[0]),.doutb(w_n3192_0[1]),.doutc(w_n3192_0[2]),.din(n3192));
	jspl jspl_w_n3193_0(.douta(w_n3193_0[0]),.doutb(w_n3193_0[1]),.din(n3193));
	jspl3 jspl3_w_n3197_0(.douta(w_n3197_0[0]),.doutb(w_n3197_0[1]),.doutc(w_n3197_0[2]),.din(n3197));
	jspl3 jspl3_w_n3199_0(.douta(w_n3199_0[0]),.doutb(w_n3199_0[1]),.doutc(w_n3199_0[2]),.din(n3199));
	jspl jspl_w_n3200_0(.douta(w_n3200_0[0]),.doutb(w_n3200_0[1]),.din(n3200));
	jspl3 jspl3_w_n3204_0(.douta(w_n3204_0[0]),.doutb(w_n3204_0[1]),.doutc(w_n3204_0[2]),.din(n3204));
	jspl3 jspl3_w_n3206_0(.douta(w_n3206_0[0]),.doutb(w_n3206_0[1]),.doutc(w_n3206_0[2]),.din(n3206));
	jspl jspl_w_n3207_0(.douta(w_n3207_0[0]),.doutb(w_n3207_0[1]),.din(n3207));
	jspl3 jspl3_w_n3211_0(.douta(w_n3211_0[0]),.doutb(w_n3211_0[1]),.doutc(w_n3211_0[2]),.din(n3211));
	jspl3 jspl3_w_n3214_0(.douta(w_n3214_0[0]),.doutb(w_n3214_0[1]),.doutc(w_n3214_0[2]),.din(n3214));
	jspl jspl_w_n3215_0(.douta(w_n3215_0[0]),.doutb(w_n3215_0[1]),.din(n3215));
	jspl3 jspl3_w_n3219_0(.douta(w_n3219_0[0]),.doutb(w_n3219_0[1]),.doutc(w_n3219_0[2]),.din(n3219));
	jspl3 jspl3_w_n3222_0(.douta(w_n3222_0[0]),.doutb(w_n3222_0[1]),.doutc(w_n3222_0[2]),.din(n3222));
	jspl jspl_w_n3223_0(.douta(w_n3223_0[0]),.doutb(w_n3223_0[1]),.din(n3223));
	jspl3 jspl3_w_n3227_0(.douta(w_n3227_0[0]),.doutb(w_n3227_0[1]),.doutc(w_n3227_0[2]),.din(n3227));
	jspl3 jspl3_w_n3229_0(.douta(w_n3229_0[0]),.doutb(w_n3229_0[1]),.doutc(w_n3229_0[2]),.din(n3229));
	jspl jspl_w_n3230_0(.douta(w_n3230_0[0]),.doutb(w_n3230_0[1]),.din(n3230));
	jspl jspl_w_n3234_0(.douta(w_n3234_0[0]),.doutb(w_n3234_0[1]),.din(n3234));
	jspl jspl_w_n3235_0(.douta(w_n3235_0[0]),.doutb(w_n3235_0[1]),.din(n3235));
	jspl3 jspl3_w_n3237_0(.douta(w_n3237_0[0]),.doutb(w_n3237_0[1]),.doutc(w_n3237_0[2]),.din(n3237));
	jspl jspl_w_n3237_1(.douta(w_n3237_1[0]),.doutb(w_n3237_1[1]),.din(w_n3237_0[0]));
	jspl3 jspl3_w_n3240_0(.douta(w_n3240_0[0]),.doutb(w_n3240_0[1]),.doutc(w_n3240_0[2]),.din(n3240));
	jspl jspl_w_n3240_1(.douta(w_n3240_1[0]),.doutb(w_n3240_1[1]),.din(w_n3240_0[0]));
	jspl jspl_w_n3241_0(.douta(w_n3241_0[0]),.doutb(w_n3241_0[1]),.din(n3241));
	jspl jspl_w_n3245_0(.douta(w_n3245_0[0]),.doutb(w_n3245_0[1]),.din(n3245));
	jspl jspl_w_n3246_0(.douta(w_n3246_0[0]),.doutb(w_n3246_0[1]),.din(n3246));
	jspl jspl_w_n3250_0(.douta(w_n3250_0[0]),.doutb(w_n3250_0[1]),.din(n3250));
	jspl jspl_w_n3253_0(.douta(w_n3253_0[0]),.doutb(w_n3253_0[1]),.din(n3253));
	jspl3 jspl3_w_n3258_0(.douta(w_n3258_0[0]),.doutb(w_n3258_0[1]),.doutc(w_n3258_0[2]),.din(n3258));
	jspl jspl_w_n3258_1(.douta(w_n3258_1[0]),.doutb(w_n3258_1[1]),.din(w_n3258_0[0]));
	jspl jspl_w_n3259_0(.douta(w_n3259_0[0]),.doutb(w_n3259_0[1]),.din(n3259));
	jspl3 jspl3_w_n3260_0(.douta(w_n3260_0[0]),.doutb(w_n3260_0[1]),.doutc(w_n3260_0[2]),.din(n3260));
	jspl jspl_w_n3261_0(.douta(w_n3261_0[0]),.doutb(w_n3261_0[1]),.din(n3261));
	jspl3 jspl3_w_n3262_0(.douta(w_n3262_0[0]),.doutb(w_n3262_0[1]),.doutc(w_n3262_0[2]),.din(n3262));
	jspl jspl_w_n3263_0(.douta(w_n3263_0[0]),.doutb(w_n3263_0[1]),.din(n3263));
	jspl jspl_w_n3268_0(.douta(w_n3268_0[0]),.doutb(w_n3268_0[1]),.din(n3268));
	jspl jspl_w_n3293_0(.douta(w_n3293_0[0]),.doutb(w_n3293_0[1]),.din(n3293));
	jspl jspl_w_n3297_0(.douta(w_n3297_0[0]),.doutb(w_n3297_0[1]),.din(n3297));
	jspl jspl_w_n3364_0(.douta(w_n3364_0[0]),.doutb(w_n3364_0[1]),.din(n3364));
	jspl jspl_w_n3367_0(.douta(w_n3367_0[0]),.doutb(w_n3367_0[1]),.din(n3367));
	jspl3 jspl3_w_n3368_0(.douta(w_n3368_0[0]),.doutb(w_n3368_0[1]),.doutc(w_n3368_0[2]),.din(n3368));
	jspl3 jspl3_w_n3368_1(.douta(w_n3368_1[0]),.doutb(w_n3368_1[1]),.doutc(w_n3368_1[2]),.din(w_n3368_0[0]));
	jspl3 jspl3_w_n3368_2(.douta(w_n3368_2[0]),.doutb(w_n3368_2[1]),.doutc(w_n3368_2[2]),.din(w_n3368_0[1]));
	jspl3 jspl3_w_n3368_3(.douta(w_n3368_3[0]),.doutb(w_n3368_3[1]),.doutc(w_n3368_3[2]),.din(w_n3368_0[2]));
	jspl3 jspl3_w_n3368_4(.douta(w_n3368_4[0]),.doutb(w_n3368_4[1]),.doutc(w_n3368_4[2]),.din(w_n3368_1[0]));
	jspl3 jspl3_w_n3368_5(.douta(w_n3368_5[0]),.doutb(w_n3368_5[1]),.doutc(w_n3368_5[2]),.din(w_n3368_1[1]));
	jspl3 jspl3_w_n3368_6(.douta(w_n3368_6[0]),.doutb(w_n3368_6[1]),.doutc(w_n3368_6[2]),.din(w_n3368_1[2]));
	jspl3 jspl3_w_n3368_7(.douta(w_n3368_7[0]),.doutb(w_n3368_7[1]),.doutc(w_n3368_7[2]),.din(w_n3368_2[0]));
	jspl3 jspl3_w_n3368_8(.douta(w_n3368_8[0]),.doutb(w_n3368_8[1]),.doutc(w_n3368_8[2]),.din(w_n3368_2[1]));
	jspl3 jspl3_w_n3368_9(.douta(w_n3368_9[0]),.doutb(w_n3368_9[1]),.doutc(w_n3368_9[2]),.din(w_n3368_2[2]));
	jspl3 jspl3_w_n3368_10(.douta(w_n3368_10[0]),.doutb(w_n3368_10[1]),.doutc(w_n3368_10[2]),.din(w_n3368_3[0]));
	jspl3 jspl3_w_n3368_11(.douta(w_n3368_11[0]),.doutb(w_n3368_11[1]),.doutc(w_n3368_11[2]),.din(w_n3368_3[1]));
	jspl3 jspl3_w_n3368_12(.douta(w_n3368_12[0]),.doutb(w_n3368_12[1]),.doutc(w_n3368_12[2]),.din(w_n3368_3[2]));
	jspl3 jspl3_w_n3368_13(.douta(w_n3368_13[0]),.doutb(w_n3368_13[1]),.doutc(w_n3368_13[2]),.din(w_n3368_4[0]));
	jspl3 jspl3_w_n3368_14(.douta(w_n3368_14[0]),.doutb(w_n3368_14[1]),.doutc(w_n3368_14[2]),.din(w_n3368_4[1]));
	jspl3 jspl3_w_n3368_15(.douta(w_n3368_15[0]),.doutb(w_n3368_15[1]),.doutc(w_n3368_15[2]),.din(w_n3368_4[2]));
	jspl3 jspl3_w_n3368_16(.douta(w_n3368_16[0]),.doutb(w_n3368_16[1]),.doutc(w_n3368_16[2]),.din(w_n3368_5[0]));
	jspl3 jspl3_w_n3368_17(.douta(w_n3368_17[0]),.doutb(w_n3368_17[1]),.doutc(w_n3368_17[2]),.din(w_n3368_5[1]));
	jspl3 jspl3_w_n3368_18(.douta(w_n3368_18[0]),.doutb(w_n3368_18[1]),.doutc(w_n3368_18[2]),.din(w_n3368_5[2]));
	jspl3 jspl3_w_n3368_19(.douta(w_n3368_19[0]),.doutb(w_n3368_19[1]),.doutc(w_n3368_19[2]),.din(w_n3368_6[0]));
	jspl3 jspl3_w_n3368_20(.douta(w_n3368_20[0]),.doutb(w_n3368_20[1]),.doutc(w_n3368_20[2]),.din(w_n3368_6[1]));
	jspl3 jspl3_w_n3368_21(.douta(w_n3368_21[0]),.doutb(w_n3368_21[1]),.doutc(w_n3368_21[2]),.din(w_n3368_6[2]));
	jspl3 jspl3_w_n3368_22(.douta(w_n3368_22[0]),.doutb(w_n3368_22[1]),.doutc(w_n3368_22[2]),.din(w_n3368_7[0]));
	jspl3 jspl3_w_n3368_23(.douta(w_n3368_23[0]),.doutb(w_n3368_23[1]),.doutc(w_n3368_23[2]),.din(w_n3368_7[1]));
	jspl3 jspl3_w_n3368_24(.douta(w_n3368_24[0]),.doutb(w_n3368_24[1]),.doutc(w_n3368_24[2]),.din(w_n3368_7[2]));
	jspl3 jspl3_w_n3368_25(.douta(w_n3368_25[0]),.doutb(w_n3368_25[1]),.doutc(w_n3368_25[2]),.din(w_n3368_8[0]));
	jspl3 jspl3_w_n3368_26(.douta(w_n3368_26[0]),.doutb(w_n3368_26[1]),.doutc(w_n3368_26[2]),.din(w_n3368_8[1]));
	jspl3 jspl3_w_n3368_27(.douta(w_n3368_27[0]),.doutb(w_n3368_27[1]),.doutc(w_n3368_27[2]),.din(w_n3368_8[2]));
	jspl3 jspl3_w_n3368_28(.douta(w_n3368_28[0]),.doutb(w_n3368_28[1]),.doutc(w_n3368_28[2]),.din(w_n3368_9[0]));
	jspl3 jspl3_w_n3368_29(.douta(w_n3368_29[0]),.doutb(w_n3368_29[1]),.doutc(w_n3368_29[2]),.din(w_n3368_9[1]));
	jspl3 jspl3_w_n3368_30(.douta(w_n3368_30[0]),.doutb(w_n3368_30[1]),.doutc(w_n3368_30[2]),.din(w_n3368_9[2]));
	jspl3 jspl3_w_n3368_31(.douta(w_n3368_31[0]),.doutb(w_n3368_31[1]),.doutc(w_n3368_31[2]),.din(w_n3368_10[0]));
	jspl3 jspl3_w_n3368_32(.douta(w_n3368_32[0]),.doutb(w_n3368_32[1]),.doutc(w_n3368_32[2]),.din(w_n3368_10[1]));
	jspl3 jspl3_w_n3368_33(.douta(w_n3368_33[0]),.doutb(w_n3368_33[1]),.doutc(w_n3368_33[2]),.din(w_n3368_10[2]));
	jspl3 jspl3_w_n3368_34(.douta(w_n3368_34[0]),.doutb(w_n3368_34[1]),.doutc(w_n3368_34[2]),.din(w_n3368_11[0]));
	jspl3 jspl3_w_n3368_35(.douta(w_n3368_35[0]),.doutb(w_n3368_35[1]),.doutc(w_n3368_35[2]),.din(w_n3368_11[1]));
	jspl3 jspl3_w_n3368_36(.douta(w_n3368_36[0]),.doutb(w_n3368_36[1]),.doutc(w_n3368_36[2]),.din(w_n3368_11[2]));
	jspl3 jspl3_w_n3368_37(.douta(w_n3368_37[0]),.doutb(w_n3368_37[1]),.doutc(w_n3368_37[2]),.din(w_n3368_12[0]));
	jspl3 jspl3_w_n3368_38(.douta(w_n3368_38[0]),.doutb(w_n3368_38[1]),.doutc(w_n3368_38[2]),.din(w_n3368_12[1]));
	jspl3 jspl3_w_n3368_39(.douta(w_n3368_39[0]),.doutb(w_n3368_39[1]),.doutc(w_n3368_39[2]),.din(w_n3368_12[2]));
	jspl3 jspl3_w_n3368_40(.douta(w_n3368_40[0]),.doutb(w_n3368_40[1]),.doutc(w_n3368_40[2]),.din(w_n3368_13[0]));
	jspl3 jspl3_w_n3368_41(.douta(w_n3368_41[0]),.doutb(w_n3368_41[1]),.doutc(w_n3368_41[2]),.din(w_n3368_13[1]));
	jspl3 jspl3_w_n3368_42(.douta(w_n3368_42[0]),.doutb(w_n3368_42[1]),.doutc(w_n3368_42[2]),.din(w_n3368_13[2]));
	jspl3 jspl3_w_n3368_43(.douta(w_n3368_43[0]),.doutb(w_n3368_43[1]),.doutc(w_n3368_43[2]),.din(w_n3368_14[0]));
	jspl3 jspl3_w_n3368_44(.douta(w_n3368_44[0]),.doutb(w_n3368_44[1]),.doutc(w_n3368_44[2]),.din(w_n3368_14[1]));
	jspl3 jspl3_w_n3368_45(.douta(w_n3368_45[0]),.doutb(w_n3368_45[1]),.doutc(w_n3368_45[2]),.din(w_n3368_14[2]));
	jspl3 jspl3_w_n3368_46(.douta(w_n3368_46[0]),.doutb(w_n3368_46[1]),.doutc(w_n3368_46[2]),.din(w_n3368_15[0]));
	jspl3 jspl3_w_n3368_47(.douta(w_n3368_47[0]),.doutb(w_n3368_47[1]),.doutc(w_n3368_47[2]),.din(w_n3368_15[1]));
	jspl3 jspl3_w_n3368_48(.douta(w_n3368_48[0]),.doutb(w_n3368_48[1]),.doutc(w_n3368_48[2]),.din(w_n3368_15[2]));
	jspl3 jspl3_w_n3368_49(.douta(w_n3368_49[0]),.doutb(w_n3368_49[1]),.doutc(w_n3368_49[2]),.din(w_n3368_16[0]));
	jspl3 jspl3_w_n3368_50(.douta(w_n3368_50[0]),.doutb(w_n3368_50[1]),.doutc(w_n3368_50[2]),.din(w_n3368_16[1]));
	jspl3 jspl3_w_n3368_51(.douta(w_n3368_51[0]),.doutb(w_n3368_51[1]),.doutc(w_n3368_51[2]),.din(w_n3368_16[2]));
	jspl jspl_w_n3368_52(.douta(w_n3368_52[0]),.doutb(w_n3368_52[1]),.din(w_n3368_17[0]));
	jspl3 jspl3_w_n3372_0(.douta(w_n3372_0[0]),.doutb(w_n3372_0[1]),.doutc(w_n3372_0[2]),.din(n3372));
	jspl jspl_w_n3373_0(.douta(w_n3373_0[0]),.doutb(w_n3373_0[1]),.din(n3373));
	jspl jspl_w_n3375_0(.douta(w_n3375_0[0]),.doutb(w_n3375_0[1]),.din(n3375));
	jspl jspl_w_n3380_0(.douta(w_n3380_0[0]),.doutb(w_n3380_0[1]),.din(n3380));
	jspl jspl_w_n3381_0(.douta(w_n3381_0[0]),.doutb(w_n3381_0[1]),.din(n3381));
	jspl3 jspl3_w_n3383_0(.douta(w_n3383_0[0]),.doutb(w_n3383_0[1]),.doutc(w_n3383_0[2]),.din(n3383));
	jspl jspl_w_n3384_0(.douta(w_n3384_0[0]),.doutb(w_n3384_0[1]),.din(n3384));
	jspl jspl_w_n3388_0(.douta(w_n3388_0[0]),.doutb(w_n3388_0[1]),.din(n3388));
	jspl3 jspl3_w_n3390_0(.douta(w_n3390_0[0]),.doutb(w_n3390_0[1]),.doutc(w_n3390_0[2]),.din(n3390));
	jspl jspl_w_n3391_0(.douta(w_n3391_0[0]),.doutb(w_n3391_0[1]),.din(n3391));
	jspl jspl_w_n3395_0(.douta(w_n3395_0[0]),.doutb(w_n3395_0[1]),.din(n3395));
	jspl3 jspl3_w_n3397_0(.douta(w_n3397_0[0]),.doutb(w_n3397_0[1]),.doutc(w_n3397_0[2]),.din(n3397));
	jspl jspl_w_n3398_0(.douta(w_n3398_0[0]),.doutb(w_n3398_0[1]),.din(n3398));
	jspl jspl_w_n3402_0(.douta(w_n3402_0[0]),.doutb(w_n3402_0[1]),.din(n3402));
	jspl jspl_w_n3403_0(.douta(w_n3403_0[0]),.doutb(w_n3403_0[1]),.din(n3403));
	jspl3 jspl3_w_n3405_0(.douta(w_n3405_0[0]),.doutb(w_n3405_0[1]),.doutc(w_n3405_0[2]),.din(n3405));
	jspl jspl_w_n3406_0(.douta(w_n3406_0[0]),.doutb(w_n3406_0[1]),.din(n3406));
	jspl jspl_w_n3410_0(.douta(w_n3410_0[0]),.doutb(w_n3410_0[1]),.din(n3410));
	jspl jspl_w_n3411_0(.douta(w_n3411_0[0]),.doutb(w_n3411_0[1]),.din(n3411));
	jspl3 jspl3_w_n3413_0(.douta(w_n3413_0[0]),.doutb(w_n3413_0[1]),.doutc(w_n3413_0[2]),.din(n3413));
	jspl jspl_w_n3414_0(.douta(w_n3414_0[0]),.doutb(w_n3414_0[1]),.din(n3414));
	jspl jspl_w_n3418_0(.douta(w_n3418_0[0]),.doutb(w_n3418_0[1]),.din(n3418));
	jspl3 jspl3_w_n3420_0(.douta(w_n3420_0[0]),.doutb(w_n3420_0[1]),.doutc(w_n3420_0[2]),.din(n3420));
	jspl jspl_w_n3421_0(.douta(w_n3421_0[0]),.doutb(w_n3421_0[1]),.din(n3421));
	jspl jspl_w_n3425_0(.douta(w_n3425_0[0]),.doutb(w_n3425_0[1]),.din(n3425));
	jspl jspl_w_n3426_0(.douta(w_n3426_0[0]),.doutb(w_n3426_0[1]),.din(n3426));
	jspl3 jspl3_w_n3428_0(.douta(w_n3428_0[0]),.doutb(w_n3428_0[1]),.doutc(w_n3428_0[2]),.din(n3428));
	jspl jspl_w_n3429_0(.douta(w_n3429_0[0]),.doutb(w_n3429_0[1]),.din(n3429));
	jspl jspl_w_n3433_0(.douta(w_n3433_0[0]),.doutb(w_n3433_0[1]),.din(n3433));
	jspl3 jspl3_w_n3435_0(.douta(w_n3435_0[0]),.doutb(w_n3435_0[1]),.doutc(w_n3435_0[2]),.din(n3435));
	jspl jspl_w_n3436_0(.douta(w_n3436_0[0]),.doutb(w_n3436_0[1]),.din(n3436));
	jspl jspl_w_n3440_0(.douta(w_n3440_0[0]),.doutb(w_n3440_0[1]),.din(n3440));
	jspl jspl_w_n3441_0(.douta(w_n3441_0[0]),.doutb(w_n3441_0[1]),.din(n3441));
	jspl3 jspl3_w_n3443_0(.douta(w_n3443_0[0]),.doutb(w_n3443_0[1]),.doutc(w_n3443_0[2]),.din(n3443));
	jspl jspl_w_n3444_0(.douta(w_n3444_0[0]),.doutb(w_n3444_0[1]),.din(n3444));
	jspl jspl_w_n3448_0(.douta(w_n3448_0[0]),.doutb(w_n3448_0[1]),.din(n3448));
	jspl3 jspl3_w_n3450_0(.douta(w_n3450_0[0]),.doutb(w_n3450_0[1]),.doutc(w_n3450_0[2]),.din(n3450));
	jspl jspl_w_n3451_0(.douta(w_n3451_0[0]),.doutb(w_n3451_0[1]),.din(n3451));
	jspl jspl_w_n3455_0(.douta(w_n3455_0[0]),.doutb(w_n3455_0[1]),.din(n3455));
	jspl jspl_w_n3456_0(.douta(w_n3456_0[0]),.doutb(w_n3456_0[1]),.din(n3456));
	jspl3 jspl3_w_n3458_0(.douta(w_n3458_0[0]),.doutb(w_n3458_0[1]),.doutc(w_n3458_0[2]),.din(n3458));
	jspl jspl_w_n3459_0(.douta(w_n3459_0[0]),.doutb(w_n3459_0[1]),.din(n3459));
	jspl jspl_w_n3463_0(.douta(w_n3463_0[0]),.doutb(w_n3463_0[1]),.din(n3463));
	jspl3 jspl3_w_n3465_0(.douta(w_n3465_0[0]),.doutb(w_n3465_0[1]),.doutc(w_n3465_0[2]),.din(n3465));
	jspl jspl_w_n3466_0(.douta(w_n3466_0[0]),.doutb(w_n3466_0[1]),.din(n3466));
	jspl jspl_w_n3470_0(.douta(w_n3470_0[0]),.doutb(w_n3470_0[1]),.din(n3470));
	jspl jspl_w_n3471_0(.douta(w_n3471_0[0]),.doutb(w_n3471_0[1]),.din(n3471));
	jspl3 jspl3_w_n3473_0(.douta(w_n3473_0[0]),.doutb(w_n3473_0[1]),.doutc(w_n3473_0[2]),.din(n3473));
	jspl jspl_w_n3474_0(.douta(w_n3474_0[0]),.doutb(w_n3474_0[1]),.din(n3474));
	jspl jspl_w_n3478_0(.douta(w_n3478_0[0]),.doutb(w_n3478_0[1]),.din(n3478));
	jspl3 jspl3_w_n3480_0(.douta(w_n3480_0[0]),.doutb(w_n3480_0[1]),.doutc(w_n3480_0[2]),.din(n3480));
	jspl jspl_w_n3481_0(.douta(w_n3481_0[0]),.doutb(w_n3481_0[1]),.din(n3481));
	jspl jspl_w_n3485_0(.douta(w_n3485_0[0]),.doutb(w_n3485_0[1]),.din(n3485));
	jspl jspl_w_n3486_0(.douta(w_n3486_0[0]),.doutb(w_n3486_0[1]),.din(n3486));
	jspl3 jspl3_w_n3488_0(.douta(w_n3488_0[0]),.doutb(w_n3488_0[1]),.doutc(w_n3488_0[2]),.din(n3488));
	jspl jspl_w_n3489_0(.douta(w_n3489_0[0]),.doutb(w_n3489_0[1]),.din(n3489));
	jspl jspl_w_n3493_0(.douta(w_n3493_0[0]),.doutb(w_n3493_0[1]),.din(n3493));
	jspl jspl_w_n3494_0(.douta(w_n3494_0[0]),.doutb(w_n3494_0[1]),.din(n3494));
	jspl3 jspl3_w_n3496_0(.douta(w_n3496_0[0]),.doutb(w_n3496_0[1]),.doutc(w_n3496_0[2]),.din(n3496));
	jspl jspl_w_n3497_0(.douta(w_n3497_0[0]),.doutb(w_n3497_0[1]),.din(n3497));
	jspl jspl_w_n3501_0(.douta(w_n3501_0[0]),.doutb(w_n3501_0[1]),.din(n3501));
	jspl3 jspl3_w_n3503_0(.douta(w_n3503_0[0]),.doutb(w_n3503_0[1]),.doutc(w_n3503_0[2]),.din(n3503));
	jspl jspl_w_n3504_0(.douta(w_n3504_0[0]),.doutb(w_n3504_0[1]),.din(n3504));
	jspl jspl_w_n3508_0(.douta(w_n3508_0[0]),.doutb(w_n3508_0[1]),.din(n3508));
	jspl3 jspl3_w_n3510_0(.douta(w_n3510_0[0]),.doutb(w_n3510_0[1]),.doutc(w_n3510_0[2]),.din(n3510));
	jspl jspl_w_n3511_0(.douta(w_n3511_0[0]),.doutb(w_n3511_0[1]),.din(n3511));
	jspl3 jspl3_w_n3515_0(.douta(w_n3515_0[0]),.doutb(w_n3515_0[1]),.doutc(w_n3515_0[2]),.din(n3515));
	jspl jspl_w_n3518_0(.douta(w_n3518_0[0]),.doutb(w_n3518_0[1]),.din(n3518));
	jspl3 jspl3_w_n3521_0(.douta(w_n3521_0[0]),.doutb(w_n3521_0[1]),.doutc(w_n3521_0[2]),.din(n3521));
	jspl jspl_w_n3522_0(.douta(w_n3522_0[0]),.doutb(w_n3522_0[1]),.din(n3522));
	jspl3 jspl3_w_n3523_0(.douta(w_n3523_0[0]),.doutb(w_n3523_0[1]),.doutc(w_n3523_0[2]),.din(n3523));
	jspl jspl_w_n3523_1(.douta(w_n3523_1[0]),.doutb(w_n3523_1[1]),.din(w_n3523_0[0]));
	jspl3 jspl3_w_n3524_0(.douta(w_n3524_0[0]),.doutb(w_n3524_0[1]),.doutc(w_n3524_0[2]),.din(n3524));
	jspl jspl_w_n3552_0(.douta(w_n3552_0[0]),.doutb(w_n3552_0[1]),.din(n3552));
	jspl jspl_w_n3559_0(.douta(w_n3559_0[0]),.doutb(w_n3559_0[1]),.din(n3559));
	jspl jspl_w_n3563_0(.douta(w_n3563_0[0]),.doutb(w_n3563_0[1]),.din(n3563));
	jspl jspl_w_n3573_0(.douta(w_n3573_0[0]),.doutb(w_n3573_0[1]),.din(n3573));
	jspl jspl_w_n3580_0(.douta(w_n3580_0[0]),.doutb(w_n3580_0[1]),.din(n3580));
	jspl jspl_w_n3587_0(.douta(w_n3587_0[0]),.doutb(w_n3587_0[1]),.din(n3587));
	jspl jspl_w_n3594_0(.douta(w_n3594_0[0]),.doutb(w_n3594_0[1]),.din(n3594));
	jspl jspl_w_n3601_0(.douta(w_n3601_0[0]),.doutb(w_n3601_0[1]),.din(n3601));
	jspl jspl_w_n3611_0(.douta(w_n3611_0[0]),.doutb(w_n3611_0[1]),.din(n3611));
	jspl jspl_w_n3615_0(.douta(w_n3615_0[0]),.doutb(w_n3615_0[1]),.din(n3615));
	jspl jspl_w_n3620_0(.douta(w_n3620_0[0]),.doutb(w_n3620_0[1]),.din(n3620));
	jspl jspl_w_n3621_0(.douta(w_n3621_0[0]),.doutb(w_n3621_0[1]),.din(n3621));
	jspl jspl_w_n3622_0(.douta(w_n3622_0[0]),.doutb(w_n3622_0[1]),.din(n3622));
	jspl jspl_w_n3624_0(.douta(w_n3624_0[0]),.doutb(w_n3624_0[1]),.din(n3624));
	jspl jspl_w_n3626_0(.douta(w_n3626_0[0]),.doutb(w_n3626_0[1]),.din(n3626));
	jspl jspl_w_n3629_0(.douta(w_n3629_0[0]),.doutb(w_n3629_0[1]),.din(n3629));
	jspl jspl_w_n3630_0(.douta(w_n3630_0[0]),.doutb(w_n3630_0[1]),.din(n3630));
	jspl jspl_w_n3631_0(.douta(w_n3631_0[0]),.doutb(w_n3631_0[1]),.din(n3631));
	jspl jspl_w_n3635_0(.douta(w_n3635_0[0]),.doutb(w_n3635_0[1]),.din(n3635));
	jspl jspl_w_n3640_0(.douta(w_n3640_0[0]),.doutb(w_n3640_0[1]),.din(n3640));
	jspl3 jspl3_w_n3642_0(.douta(w_n3642_0[0]),.doutb(w_n3642_0[1]),.doutc(w_n3642_0[2]),.din(n3642));
	jspl3 jspl3_w_n3642_1(.douta(w_n3642_1[0]),.doutb(w_n3642_1[1]),.doutc(w_n3642_1[2]),.din(w_n3642_0[0]));
	jspl3 jspl3_w_n3642_2(.douta(w_n3642_2[0]),.doutb(w_n3642_2[1]),.doutc(w_n3642_2[2]),.din(w_n3642_0[1]));
	jspl3 jspl3_w_n3642_3(.douta(w_n3642_3[0]),.doutb(w_n3642_3[1]),.doutc(w_n3642_3[2]),.din(w_n3642_0[2]));
	jspl3 jspl3_w_n3642_4(.douta(w_n3642_4[0]),.doutb(w_n3642_4[1]),.doutc(w_n3642_4[2]),.din(w_n3642_1[0]));
	jspl3 jspl3_w_n3642_5(.douta(w_n3642_5[0]),.doutb(w_n3642_5[1]),.doutc(w_n3642_5[2]),.din(w_n3642_1[1]));
	jspl3 jspl3_w_n3642_6(.douta(w_n3642_6[0]),.doutb(w_n3642_6[1]),.doutc(w_n3642_6[2]),.din(w_n3642_1[2]));
	jspl3 jspl3_w_n3642_7(.douta(w_n3642_7[0]),.doutb(w_n3642_7[1]),.doutc(w_n3642_7[2]),.din(w_n3642_2[0]));
	jspl3 jspl3_w_n3642_8(.douta(w_n3642_8[0]),.doutb(w_n3642_8[1]),.doutc(w_n3642_8[2]),.din(w_n3642_2[1]));
	jspl3 jspl3_w_n3642_9(.douta(w_n3642_9[0]),.doutb(w_n3642_9[1]),.doutc(w_n3642_9[2]),.din(w_n3642_2[2]));
	jspl3 jspl3_w_n3642_10(.douta(w_n3642_10[0]),.doutb(w_n3642_10[1]),.doutc(w_n3642_10[2]),.din(w_n3642_3[0]));
	jspl3 jspl3_w_n3642_11(.douta(w_n3642_11[0]),.doutb(w_n3642_11[1]),.doutc(w_n3642_11[2]),.din(w_n3642_3[1]));
	jspl3 jspl3_w_n3642_12(.douta(w_n3642_12[0]),.doutb(w_n3642_12[1]),.doutc(w_n3642_12[2]),.din(w_n3642_3[2]));
	jspl3 jspl3_w_n3642_13(.douta(w_n3642_13[0]),.doutb(w_n3642_13[1]),.doutc(w_n3642_13[2]),.din(w_n3642_4[0]));
	jspl3 jspl3_w_n3642_14(.douta(w_n3642_14[0]),.doutb(w_n3642_14[1]),.doutc(w_n3642_14[2]),.din(w_n3642_4[1]));
	jspl3 jspl3_w_n3642_15(.douta(w_n3642_15[0]),.doutb(w_n3642_15[1]),.doutc(w_n3642_15[2]),.din(w_n3642_4[2]));
	jspl3 jspl3_w_n3642_16(.douta(w_n3642_16[0]),.doutb(w_n3642_16[1]),.doutc(w_n3642_16[2]),.din(w_n3642_5[0]));
	jspl3 jspl3_w_n3642_17(.douta(w_n3642_17[0]),.doutb(w_n3642_17[1]),.doutc(w_n3642_17[2]),.din(w_n3642_5[1]));
	jspl3 jspl3_w_n3642_18(.douta(w_n3642_18[0]),.doutb(w_n3642_18[1]),.doutc(w_n3642_18[2]),.din(w_n3642_5[2]));
	jspl3 jspl3_w_n3642_19(.douta(w_n3642_19[0]),.doutb(w_n3642_19[1]),.doutc(w_n3642_19[2]),.din(w_n3642_6[0]));
	jspl3 jspl3_w_n3642_20(.douta(w_n3642_20[0]),.doutb(w_n3642_20[1]),.doutc(w_n3642_20[2]),.din(w_n3642_6[1]));
	jspl3 jspl3_w_n3642_21(.douta(w_n3642_21[0]),.doutb(w_n3642_21[1]),.doutc(w_n3642_21[2]),.din(w_n3642_6[2]));
	jspl3 jspl3_w_n3642_22(.douta(w_n3642_22[0]),.doutb(w_n3642_22[1]),.doutc(w_n3642_22[2]),.din(w_n3642_7[0]));
	jspl3 jspl3_w_n3642_23(.douta(w_n3642_23[0]),.doutb(w_n3642_23[1]),.doutc(w_n3642_23[2]),.din(w_n3642_7[1]));
	jspl3 jspl3_w_n3642_24(.douta(w_n3642_24[0]),.doutb(w_n3642_24[1]),.doutc(w_n3642_24[2]),.din(w_n3642_7[2]));
	jspl3 jspl3_w_n3642_25(.douta(w_n3642_25[0]),.doutb(w_n3642_25[1]),.doutc(w_n3642_25[2]),.din(w_n3642_8[0]));
	jspl3 jspl3_w_n3642_26(.douta(w_n3642_26[0]),.doutb(w_n3642_26[1]),.doutc(w_n3642_26[2]),.din(w_n3642_8[1]));
	jspl3 jspl3_w_n3642_27(.douta(w_n3642_27[0]),.doutb(w_n3642_27[1]),.doutc(w_n3642_27[2]),.din(w_n3642_8[2]));
	jspl3 jspl3_w_n3642_28(.douta(w_n3642_28[0]),.doutb(w_n3642_28[1]),.doutc(w_n3642_28[2]),.din(w_n3642_9[0]));
	jspl3 jspl3_w_n3642_29(.douta(w_n3642_29[0]),.doutb(w_n3642_29[1]),.doutc(w_n3642_29[2]),.din(w_n3642_9[1]));
	jspl3 jspl3_w_n3642_30(.douta(w_n3642_30[0]),.doutb(w_n3642_30[1]),.doutc(w_n3642_30[2]),.din(w_n3642_9[2]));
	jspl3 jspl3_w_n3642_31(.douta(w_n3642_31[0]),.doutb(w_n3642_31[1]),.doutc(w_n3642_31[2]),.din(w_n3642_10[0]));
	jspl3 jspl3_w_n3642_32(.douta(w_n3642_32[0]),.doutb(w_n3642_32[1]),.doutc(w_n3642_32[2]),.din(w_n3642_10[1]));
	jspl3 jspl3_w_n3642_33(.douta(w_n3642_33[0]),.doutb(w_n3642_33[1]),.doutc(w_n3642_33[2]),.din(w_n3642_10[2]));
	jspl3 jspl3_w_n3642_34(.douta(w_n3642_34[0]),.doutb(w_n3642_34[1]),.doutc(w_n3642_34[2]),.din(w_n3642_11[0]));
	jspl3 jspl3_w_n3642_35(.douta(w_n3642_35[0]),.doutb(w_n3642_35[1]),.doutc(w_n3642_35[2]),.din(w_n3642_11[1]));
	jspl3 jspl3_w_n3642_36(.douta(w_n3642_36[0]),.doutb(w_n3642_36[1]),.doutc(w_n3642_36[2]),.din(w_n3642_11[2]));
	jspl3 jspl3_w_n3642_37(.douta(w_n3642_37[0]),.doutb(w_n3642_37[1]),.doutc(w_n3642_37[2]),.din(w_n3642_12[0]));
	jspl3 jspl3_w_n3642_38(.douta(w_n3642_38[0]),.doutb(w_n3642_38[1]),.doutc(w_n3642_38[2]),.din(w_n3642_12[1]));
	jspl3 jspl3_w_n3642_39(.douta(w_n3642_39[0]),.doutb(w_n3642_39[1]),.doutc(w_n3642_39[2]),.din(w_n3642_12[2]));
	jspl3 jspl3_w_n3642_40(.douta(w_n3642_40[0]),.doutb(w_n3642_40[1]),.doutc(w_n3642_40[2]),.din(w_n3642_13[0]));
	jspl3 jspl3_w_n3642_41(.douta(w_n3642_41[0]),.doutb(w_n3642_41[1]),.doutc(w_n3642_41[2]),.din(w_n3642_13[1]));
	jspl3 jspl3_w_n3642_42(.douta(w_n3642_42[0]),.doutb(w_n3642_42[1]),.doutc(w_n3642_42[2]),.din(w_n3642_13[2]));
	jspl3 jspl3_w_n3642_43(.douta(w_n3642_43[0]),.doutb(w_n3642_43[1]),.doutc(w_n3642_43[2]),.din(w_n3642_14[0]));
	jspl3 jspl3_w_n3642_44(.douta(w_n3642_44[0]),.doutb(w_n3642_44[1]),.doutc(w_n3642_44[2]),.din(w_n3642_14[1]));
	jspl3 jspl3_w_n3642_45(.douta(w_n3642_45[0]),.doutb(w_n3642_45[1]),.doutc(w_n3642_45[2]),.din(w_n3642_14[2]));
	jspl3 jspl3_w_n3642_46(.douta(w_n3642_46[0]),.doutb(w_n3642_46[1]),.doutc(w_n3642_46[2]),.din(w_n3642_15[0]));
	jspl3 jspl3_w_n3642_47(.douta(w_n3642_47[0]),.doutb(w_n3642_47[1]),.doutc(w_n3642_47[2]),.din(w_n3642_15[1]));
	jspl3 jspl3_w_n3642_48(.douta(w_n3642_48[0]),.doutb(w_n3642_48[1]),.doutc(w_n3642_48[2]),.din(w_n3642_15[2]));
	jspl3 jspl3_w_n3642_49(.douta(w_n3642_49[0]),.doutb(w_n3642_49[1]),.doutc(w_n3642_49[2]),.din(w_n3642_16[0]));
	jspl3 jspl3_w_n3642_50(.douta(w_n3642_50[0]),.doutb(w_n3642_50[1]),.doutc(w_n3642_50[2]),.din(w_n3642_16[1]));
	jspl3 jspl3_w_n3642_51(.douta(w_n3642_51[0]),.doutb(w_n3642_51[1]),.doutc(w_n3642_51[2]),.din(w_n3642_16[2]));
	jspl3 jspl3_w_n3642_52(.douta(w_n3642_52[0]),.doutb(w_n3642_52[1]),.doutc(w_n3642_52[2]),.din(w_n3642_17[0]));
	jspl3 jspl3_w_n3642_53(.douta(w_n3642_53[0]),.doutb(w_n3642_53[1]),.doutc(w_n3642_53[2]),.din(w_n3642_17[1]));
	jspl3 jspl3_w_n3642_54(.douta(w_n3642_54[0]),.doutb(w_n3642_54[1]),.doutc(w_n3642_54[2]),.din(w_n3642_17[2]));
	jspl3 jspl3_w_n3642_55(.douta(w_n3642_55[0]),.doutb(w_n3642_55[1]),.doutc(w_n3642_55[2]),.din(w_n3642_18[0]));
	jspl3 jspl3_w_n3642_56(.douta(w_n3642_56[0]),.doutb(w_n3642_56[1]),.doutc(w_n3642_56[2]),.din(w_n3642_18[1]));
	jspl3 jspl3_w_n3642_57(.douta(w_n3642_57[0]),.doutb(w_n3642_57[1]),.doutc(w_n3642_57[2]),.din(w_n3642_18[2]));
	jspl3 jspl3_w_n3642_58(.douta(w_n3642_58[0]),.doutb(w_n3642_58[1]),.doutc(w_n3642_58[2]),.din(w_n3642_19[0]));
	jspl3 jspl3_w_n3642_59(.douta(w_n3642_59[0]),.doutb(w_n3642_59[1]),.doutc(w_n3642_59[2]),.din(w_n3642_19[1]));
	jspl3 jspl3_w_n3642_60(.douta(w_n3642_60[0]),.doutb(w_n3642_60[1]),.doutc(w_n3642_60[2]),.din(w_n3642_19[2]));
	jspl jspl_w_n3645_0(.douta(w_n3645_0[0]),.doutb(w_n3645_0[1]),.din(n3645));
	jspl3 jspl3_w_n3646_0(.douta(w_n3646_0[0]),.doutb(w_n3646_0[1]),.doutc(w_n3646_0[2]),.din(n3646));
	jspl jspl_w_n3646_1(.douta(w_n3646_1[0]),.doutb(w_n3646_1[1]),.din(w_n3646_0[0]));
	jspl3 jspl3_w_n3648_0(.douta(w_n3648_0[0]),.doutb(w_n3648_0[1]),.doutc(w_n3648_0[2]),.din(n3648));
	jspl3 jspl3_w_n3648_1(.douta(w_n3648_1[0]),.doutb(w_n3648_1[1]),.doutc(w_n3648_1[2]),.din(w_n3648_0[0]));
	jspl jspl_w_n3649_0(.douta(w_n3649_0[0]),.doutb(w_n3649_0[1]),.din(n3649));
	jspl3 jspl3_w_n3650_0(.douta(w_n3650_0[0]),.doutb(w_n3650_0[1]),.doutc(w_n3650_0[2]),.din(n3650));
	jspl jspl_w_n3651_0(.douta(w_n3651_0[0]),.doutb(w_n3651_0[1]),.din(n3651));
	jspl3 jspl3_w_n3653_0(.douta(w_n3653_0[0]),.doutb(w_n3653_0[1]),.doutc(w_n3653_0[2]),.din(n3653));
	jspl jspl_w_n3654_0(.douta(w_n3654_0[0]),.doutb(w_n3654_0[1]),.din(n3654));
	jspl3 jspl3_w_n3661_0(.douta(w_n3661_0[0]),.doutb(w_n3661_0[1]),.doutc(w_n3661_0[2]),.din(n3661));
	jspl jspl_w_n3662_0(.douta(w_n3662_0[0]),.doutb(w_n3662_0[1]),.din(n3662));
	jspl jspl_w_n3665_0(.douta(w_n3665_0[0]),.doutb(w_n3665_0[1]),.din(n3665));
	jspl3 jspl3_w_n3670_0(.douta(w_n3670_0[0]),.doutb(w_n3670_0[1]),.doutc(w_n3670_0[2]),.din(n3670));
	jspl3 jspl3_w_n3672_0(.douta(w_n3672_0[0]),.doutb(w_n3672_0[1]),.doutc(w_n3672_0[2]),.din(n3672));
	jspl jspl_w_n3673_0(.douta(w_n3673_0[0]),.doutb(w_n3673_0[1]),.din(n3673));
	jspl3 jspl3_w_n3677_0(.douta(w_n3677_0[0]),.doutb(w_n3677_0[1]),.doutc(w_n3677_0[2]),.din(n3677));
	jspl3 jspl3_w_n3680_0(.douta(w_n3680_0[0]),.doutb(w_n3680_0[1]),.doutc(w_n3680_0[2]),.din(n3680));
	jspl jspl_w_n3681_0(.douta(w_n3681_0[0]),.doutb(w_n3681_0[1]),.din(n3681));
	jspl3 jspl3_w_n3685_0(.douta(w_n3685_0[0]),.doutb(w_n3685_0[1]),.doutc(w_n3685_0[2]),.din(n3685));
	jspl3 jspl3_w_n3687_0(.douta(w_n3687_0[0]),.doutb(w_n3687_0[1]),.doutc(w_n3687_0[2]),.din(n3687));
	jspl jspl_w_n3688_0(.douta(w_n3688_0[0]),.doutb(w_n3688_0[1]),.din(n3688));
	jspl3 jspl3_w_n3692_0(.douta(w_n3692_0[0]),.doutb(w_n3692_0[1]),.doutc(w_n3692_0[2]),.din(n3692));
	jspl3 jspl3_w_n3695_0(.douta(w_n3695_0[0]),.doutb(w_n3695_0[1]),.doutc(w_n3695_0[2]),.din(n3695));
	jspl jspl_w_n3696_0(.douta(w_n3696_0[0]),.doutb(w_n3696_0[1]),.din(n3696));
	jspl3 jspl3_w_n3700_0(.douta(w_n3700_0[0]),.doutb(w_n3700_0[1]),.doutc(w_n3700_0[2]),.din(n3700));
	jspl3 jspl3_w_n3703_0(.douta(w_n3703_0[0]),.doutb(w_n3703_0[1]),.doutc(w_n3703_0[2]),.din(n3703));
	jspl jspl_w_n3704_0(.douta(w_n3704_0[0]),.doutb(w_n3704_0[1]),.din(n3704));
	jspl3 jspl3_w_n3708_0(.douta(w_n3708_0[0]),.doutb(w_n3708_0[1]),.doutc(w_n3708_0[2]),.din(n3708));
	jspl3 jspl3_w_n3710_0(.douta(w_n3710_0[0]),.doutb(w_n3710_0[1]),.doutc(w_n3710_0[2]),.din(n3710));
	jspl jspl_w_n3711_0(.douta(w_n3711_0[0]),.doutb(w_n3711_0[1]),.din(n3711));
	jspl3 jspl3_w_n3715_0(.douta(w_n3715_0[0]),.doutb(w_n3715_0[1]),.doutc(w_n3715_0[2]),.din(n3715));
	jspl3 jspl3_w_n3717_0(.douta(w_n3717_0[0]),.doutb(w_n3717_0[1]),.doutc(w_n3717_0[2]),.din(n3717));
	jspl jspl_w_n3718_0(.douta(w_n3718_0[0]),.doutb(w_n3718_0[1]),.din(n3718));
	jspl3 jspl3_w_n3722_0(.douta(w_n3722_0[0]),.doutb(w_n3722_0[1]),.doutc(w_n3722_0[2]),.din(n3722));
	jspl3 jspl3_w_n3725_0(.douta(w_n3725_0[0]),.doutb(w_n3725_0[1]),.doutc(w_n3725_0[2]),.din(n3725));
	jspl jspl_w_n3726_0(.douta(w_n3726_0[0]),.doutb(w_n3726_0[1]),.din(n3726));
	jspl3 jspl3_w_n3730_0(.douta(w_n3730_0[0]),.doutb(w_n3730_0[1]),.doutc(w_n3730_0[2]),.din(n3730));
	jspl3 jspl3_w_n3732_0(.douta(w_n3732_0[0]),.doutb(w_n3732_0[1]),.doutc(w_n3732_0[2]),.din(n3732));
	jspl jspl_w_n3733_0(.douta(w_n3733_0[0]),.doutb(w_n3733_0[1]),.din(n3733));
	jspl3 jspl3_w_n3737_0(.douta(w_n3737_0[0]),.doutb(w_n3737_0[1]),.doutc(w_n3737_0[2]),.din(n3737));
	jspl3 jspl3_w_n3740_0(.douta(w_n3740_0[0]),.doutb(w_n3740_0[1]),.doutc(w_n3740_0[2]),.din(n3740));
	jspl jspl_w_n3741_0(.douta(w_n3741_0[0]),.doutb(w_n3741_0[1]),.din(n3741));
	jspl3 jspl3_w_n3745_0(.douta(w_n3745_0[0]),.doutb(w_n3745_0[1]),.doutc(w_n3745_0[2]),.din(n3745));
	jspl3 jspl3_w_n3747_0(.douta(w_n3747_0[0]),.doutb(w_n3747_0[1]),.doutc(w_n3747_0[2]),.din(n3747));
	jspl jspl_w_n3748_0(.douta(w_n3748_0[0]),.doutb(w_n3748_0[1]),.din(n3748));
	jspl3 jspl3_w_n3752_0(.douta(w_n3752_0[0]),.doutb(w_n3752_0[1]),.doutc(w_n3752_0[2]),.din(n3752));
	jspl3 jspl3_w_n3755_0(.douta(w_n3755_0[0]),.doutb(w_n3755_0[1]),.doutc(w_n3755_0[2]),.din(n3755));
	jspl jspl_w_n3756_0(.douta(w_n3756_0[0]),.doutb(w_n3756_0[1]),.din(n3756));
	jspl3 jspl3_w_n3760_0(.douta(w_n3760_0[0]),.doutb(w_n3760_0[1]),.doutc(w_n3760_0[2]),.din(n3760));
	jspl3 jspl3_w_n3762_0(.douta(w_n3762_0[0]),.doutb(w_n3762_0[1]),.doutc(w_n3762_0[2]),.din(n3762));
	jspl jspl_w_n3763_0(.douta(w_n3763_0[0]),.doutb(w_n3763_0[1]),.din(n3763));
	jspl3 jspl3_w_n3767_0(.douta(w_n3767_0[0]),.doutb(w_n3767_0[1]),.doutc(w_n3767_0[2]),.din(n3767));
	jspl3 jspl3_w_n3770_0(.douta(w_n3770_0[0]),.doutb(w_n3770_0[1]),.doutc(w_n3770_0[2]),.din(n3770));
	jspl jspl_w_n3771_0(.douta(w_n3771_0[0]),.doutb(w_n3771_0[1]),.din(n3771));
	jspl3 jspl3_w_n3775_0(.douta(w_n3775_0[0]),.doutb(w_n3775_0[1]),.doutc(w_n3775_0[2]),.din(n3775));
	jspl3 jspl3_w_n3777_0(.douta(w_n3777_0[0]),.doutb(w_n3777_0[1]),.doutc(w_n3777_0[2]),.din(n3777));
	jspl jspl_w_n3778_0(.douta(w_n3778_0[0]),.doutb(w_n3778_0[1]),.din(n3778));
	jspl3 jspl3_w_n3782_0(.douta(w_n3782_0[0]),.doutb(w_n3782_0[1]),.doutc(w_n3782_0[2]),.din(n3782));
	jspl3 jspl3_w_n3785_0(.douta(w_n3785_0[0]),.doutb(w_n3785_0[1]),.doutc(w_n3785_0[2]),.din(n3785));
	jspl jspl_w_n3786_0(.douta(w_n3786_0[0]),.doutb(w_n3786_0[1]),.din(n3786));
	jspl3 jspl3_w_n3790_0(.douta(w_n3790_0[0]),.doutb(w_n3790_0[1]),.doutc(w_n3790_0[2]),.din(n3790));
	jspl3 jspl3_w_n3792_0(.douta(w_n3792_0[0]),.doutb(w_n3792_0[1]),.doutc(w_n3792_0[2]),.din(n3792));
	jspl jspl_w_n3793_0(.douta(w_n3793_0[0]),.doutb(w_n3793_0[1]),.din(n3793));
	jspl3 jspl3_w_n3797_0(.douta(w_n3797_0[0]),.doutb(w_n3797_0[1]),.doutc(w_n3797_0[2]),.din(n3797));
	jspl3 jspl3_w_n3799_0(.douta(w_n3799_0[0]),.doutb(w_n3799_0[1]),.doutc(w_n3799_0[2]),.din(n3799));
	jspl jspl_w_n3800_0(.douta(w_n3800_0[0]),.doutb(w_n3800_0[1]),.din(n3800));
	jspl3 jspl3_w_n3804_0(.douta(w_n3804_0[0]),.doutb(w_n3804_0[1]),.doutc(w_n3804_0[2]),.din(n3804));
	jspl3 jspl3_w_n3807_0(.douta(w_n3807_0[0]),.doutb(w_n3807_0[1]),.doutc(w_n3807_0[2]),.din(n3807));
	jspl jspl_w_n3808_0(.douta(w_n3808_0[0]),.doutb(w_n3808_0[1]),.din(n3808));
	jspl3 jspl3_w_n3812_0(.douta(w_n3812_0[0]),.doutb(w_n3812_0[1]),.doutc(w_n3812_0[2]),.din(n3812));
	jspl3 jspl3_w_n3815_0(.douta(w_n3815_0[0]),.doutb(w_n3815_0[1]),.doutc(w_n3815_0[2]),.din(n3815));
	jspl jspl_w_n3815_1(.douta(w_n3815_1[0]),.doutb(w_n3815_1[1]),.din(w_n3815_0[0]));
	jspl jspl_w_n3816_0(.douta(w_n3816_0[0]),.doutb(w_n3816_0[1]),.din(n3816));
	jspl jspl_w_n3820_0(.douta(w_n3820_0[0]),.doutb(w_n3820_0[1]),.din(n3820));
	jspl jspl_w_n3821_0(.douta(w_n3821_0[0]),.doutb(w_n3821_0[1]),.din(n3821));
	jspl jspl_w_n3823_0(.douta(w_n3823_0[0]),.doutb(w_n3823_0[1]),.din(n3823));
	jspl jspl_w_n3828_0(.douta(w_n3828_0[0]),.doutb(w_n3828_0[1]),.din(n3828));
	jspl3 jspl3_w_n3834_0(.douta(w_n3834_0[0]),.doutb(w_n3834_0[1]),.doutc(w_n3834_0[2]),.din(n3834));
	jspl3 jspl3_w_n3835_0(.douta(w_n3835_0[0]),.doutb(w_n3835_0[1]),.doutc(w_n3835_0[2]),.din(n3835));
	jspl3 jspl3_w_n3837_0(.douta(w_n3837_0[0]),.doutb(w_n3837_0[1]),.doutc(w_n3837_0[2]),.din(n3837));
	jspl jspl_w_n3837_1(.douta(w_n3837_1[0]),.doutb(w_n3837_1[1]),.din(w_n3837_0[0]));
	jspl jspl_w_n3838_0(.douta(w_n3838_0[0]),.doutb(w_n3838_0[1]),.din(n3838));
	jspl3 jspl3_w_n3839_0(.douta(w_n3839_0[0]),.doutb(w_n3839_0[1]),.doutc(w_n3839_0[2]),.din(n3839));
	jspl jspl_w_n3840_0(.douta(w_n3840_0[0]),.doutb(w_n3840_0[1]),.din(n3840));
	jspl3 jspl3_w_n3841_0(.douta(w_n3841_0[0]),.doutb(w_n3841_0[1]),.doutc(w_n3841_0[2]),.din(n3841));
	jspl jspl_w_n3842_0(.douta(w_n3842_0[0]),.doutb(w_n3842_0[1]),.din(n3842));
	jspl jspl_w_n3847_0(.douta(w_n3847_0[0]),.doutb(w_n3847_0[1]),.din(n3847));
	jspl jspl_w_n3875_0(.douta(w_n3875_0[0]),.doutb(w_n3875_0[1]),.din(n3875));
	jspl jspl_w_n3951_0(.douta(w_n3951_0[0]),.doutb(w_n3951_0[1]),.din(n3951));
	jspl jspl_w_n3954_0(.douta(w_n3954_0[0]),.doutb(w_n3954_0[1]),.din(n3954));
	jspl3 jspl3_w_n3955_0(.douta(w_n3955_0[0]),.doutb(w_n3955_0[1]),.doutc(w_n3955_0[2]),.din(n3955));
	jspl3 jspl3_w_n3955_1(.douta(w_n3955_1[0]),.doutb(w_n3955_1[1]),.doutc(w_n3955_1[2]),.din(w_n3955_0[0]));
	jspl3 jspl3_w_n3955_2(.douta(w_n3955_2[0]),.doutb(w_n3955_2[1]),.doutc(w_n3955_2[2]),.din(w_n3955_0[1]));
	jspl3 jspl3_w_n3955_3(.douta(w_n3955_3[0]),.doutb(w_n3955_3[1]),.doutc(w_n3955_3[2]),.din(w_n3955_0[2]));
	jspl3 jspl3_w_n3955_4(.douta(w_n3955_4[0]),.doutb(w_n3955_4[1]),.doutc(w_n3955_4[2]),.din(w_n3955_1[0]));
	jspl3 jspl3_w_n3955_5(.douta(w_n3955_5[0]),.doutb(w_n3955_5[1]),.doutc(w_n3955_5[2]),.din(w_n3955_1[1]));
	jspl3 jspl3_w_n3955_6(.douta(w_n3955_6[0]),.doutb(w_n3955_6[1]),.doutc(w_n3955_6[2]),.din(w_n3955_1[2]));
	jspl3 jspl3_w_n3955_7(.douta(w_n3955_7[0]),.doutb(w_n3955_7[1]),.doutc(w_n3955_7[2]),.din(w_n3955_2[0]));
	jspl3 jspl3_w_n3955_8(.douta(w_n3955_8[0]),.doutb(w_n3955_8[1]),.doutc(w_n3955_8[2]),.din(w_n3955_2[1]));
	jspl3 jspl3_w_n3955_9(.douta(w_n3955_9[0]),.doutb(w_n3955_9[1]),.doutc(w_n3955_9[2]),.din(w_n3955_2[2]));
	jspl3 jspl3_w_n3955_10(.douta(w_n3955_10[0]),.doutb(w_n3955_10[1]),.doutc(w_n3955_10[2]),.din(w_n3955_3[0]));
	jspl3 jspl3_w_n3955_11(.douta(w_n3955_11[0]),.doutb(w_n3955_11[1]),.doutc(w_n3955_11[2]),.din(w_n3955_3[1]));
	jspl3 jspl3_w_n3955_12(.douta(w_n3955_12[0]),.doutb(w_n3955_12[1]),.doutc(w_n3955_12[2]),.din(w_n3955_3[2]));
	jspl3 jspl3_w_n3955_13(.douta(w_n3955_13[0]),.doutb(w_n3955_13[1]),.doutc(w_n3955_13[2]),.din(w_n3955_4[0]));
	jspl3 jspl3_w_n3955_14(.douta(w_n3955_14[0]),.doutb(w_n3955_14[1]),.doutc(w_n3955_14[2]),.din(w_n3955_4[1]));
	jspl3 jspl3_w_n3955_15(.douta(w_n3955_15[0]),.doutb(w_n3955_15[1]),.doutc(w_n3955_15[2]),.din(w_n3955_4[2]));
	jspl3 jspl3_w_n3955_16(.douta(w_n3955_16[0]),.doutb(w_n3955_16[1]),.doutc(w_n3955_16[2]),.din(w_n3955_5[0]));
	jspl3 jspl3_w_n3955_17(.douta(w_n3955_17[0]),.doutb(w_n3955_17[1]),.doutc(w_n3955_17[2]),.din(w_n3955_5[1]));
	jspl3 jspl3_w_n3955_18(.douta(w_n3955_18[0]),.doutb(w_n3955_18[1]),.doutc(w_n3955_18[2]),.din(w_n3955_5[2]));
	jspl3 jspl3_w_n3955_19(.douta(w_n3955_19[0]),.doutb(w_n3955_19[1]),.doutc(w_n3955_19[2]),.din(w_n3955_6[0]));
	jspl3 jspl3_w_n3955_20(.douta(w_n3955_20[0]),.doutb(w_n3955_20[1]),.doutc(w_n3955_20[2]),.din(w_n3955_6[1]));
	jspl3 jspl3_w_n3955_21(.douta(w_n3955_21[0]),.doutb(w_n3955_21[1]),.doutc(w_n3955_21[2]),.din(w_n3955_6[2]));
	jspl3 jspl3_w_n3955_22(.douta(w_n3955_22[0]),.doutb(w_n3955_22[1]),.doutc(w_n3955_22[2]),.din(w_n3955_7[0]));
	jspl3 jspl3_w_n3955_23(.douta(w_n3955_23[0]),.doutb(w_n3955_23[1]),.doutc(w_n3955_23[2]),.din(w_n3955_7[1]));
	jspl3 jspl3_w_n3955_24(.douta(w_n3955_24[0]),.doutb(w_n3955_24[1]),.doutc(w_n3955_24[2]),.din(w_n3955_7[2]));
	jspl3 jspl3_w_n3955_25(.douta(w_n3955_25[0]),.doutb(w_n3955_25[1]),.doutc(w_n3955_25[2]),.din(w_n3955_8[0]));
	jspl3 jspl3_w_n3955_26(.douta(w_n3955_26[0]),.doutb(w_n3955_26[1]),.doutc(w_n3955_26[2]),.din(w_n3955_8[1]));
	jspl3 jspl3_w_n3955_27(.douta(w_n3955_27[0]),.doutb(w_n3955_27[1]),.doutc(w_n3955_27[2]),.din(w_n3955_8[2]));
	jspl3 jspl3_w_n3955_28(.douta(w_n3955_28[0]),.doutb(w_n3955_28[1]),.doutc(w_n3955_28[2]),.din(w_n3955_9[0]));
	jspl3 jspl3_w_n3955_29(.douta(w_n3955_29[0]),.doutb(w_n3955_29[1]),.doutc(w_n3955_29[2]),.din(w_n3955_9[1]));
	jspl3 jspl3_w_n3955_30(.douta(w_n3955_30[0]),.doutb(w_n3955_30[1]),.doutc(w_n3955_30[2]),.din(w_n3955_9[2]));
	jspl3 jspl3_w_n3955_31(.douta(w_n3955_31[0]),.doutb(w_n3955_31[1]),.doutc(w_n3955_31[2]),.din(w_n3955_10[0]));
	jspl3 jspl3_w_n3955_32(.douta(w_n3955_32[0]),.doutb(w_n3955_32[1]),.doutc(w_n3955_32[2]),.din(w_n3955_10[1]));
	jspl3 jspl3_w_n3955_33(.douta(w_n3955_33[0]),.doutb(w_n3955_33[1]),.doutc(w_n3955_33[2]),.din(w_n3955_10[2]));
	jspl3 jspl3_w_n3955_34(.douta(w_n3955_34[0]),.doutb(w_n3955_34[1]),.doutc(w_n3955_34[2]),.din(w_n3955_11[0]));
	jspl3 jspl3_w_n3955_35(.douta(w_n3955_35[0]),.doutb(w_n3955_35[1]),.doutc(w_n3955_35[2]),.din(w_n3955_11[1]));
	jspl3 jspl3_w_n3955_36(.douta(w_n3955_36[0]),.doutb(w_n3955_36[1]),.doutc(w_n3955_36[2]),.din(w_n3955_11[2]));
	jspl3 jspl3_w_n3955_37(.douta(w_n3955_37[0]),.doutb(w_n3955_37[1]),.doutc(w_n3955_37[2]),.din(w_n3955_12[0]));
	jspl3 jspl3_w_n3955_38(.douta(w_n3955_38[0]),.doutb(w_n3955_38[1]),.doutc(w_n3955_38[2]),.din(w_n3955_12[1]));
	jspl3 jspl3_w_n3955_39(.douta(w_n3955_39[0]),.doutb(w_n3955_39[1]),.doutc(w_n3955_39[2]),.din(w_n3955_12[2]));
	jspl3 jspl3_w_n3955_40(.douta(w_n3955_40[0]),.doutb(w_n3955_40[1]),.doutc(w_n3955_40[2]),.din(w_n3955_13[0]));
	jspl3 jspl3_w_n3955_41(.douta(w_n3955_41[0]),.doutb(w_n3955_41[1]),.doutc(w_n3955_41[2]),.din(w_n3955_13[1]));
	jspl3 jspl3_w_n3955_42(.douta(w_n3955_42[0]),.doutb(w_n3955_42[1]),.doutc(w_n3955_42[2]),.din(w_n3955_13[2]));
	jspl3 jspl3_w_n3955_43(.douta(w_n3955_43[0]),.doutb(w_n3955_43[1]),.doutc(w_n3955_43[2]),.din(w_n3955_14[0]));
	jspl3 jspl3_w_n3955_44(.douta(w_n3955_44[0]),.doutb(w_n3955_44[1]),.doutc(w_n3955_44[2]),.din(w_n3955_14[1]));
	jspl3 jspl3_w_n3955_45(.douta(w_n3955_45[0]),.doutb(w_n3955_45[1]),.doutc(w_n3955_45[2]),.din(w_n3955_14[2]));
	jspl3 jspl3_w_n3955_46(.douta(w_n3955_46[0]),.doutb(w_n3955_46[1]),.doutc(w_n3955_46[2]),.din(w_n3955_15[0]));
	jspl3 jspl3_w_n3955_47(.douta(w_n3955_47[0]),.doutb(w_n3955_47[1]),.doutc(w_n3955_47[2]),.din(w_n3955_15[1]));
	jspl3 jspl3_w_n3955_48(.douta(w_n3955_48[0]),.doutb(w_n3955_48[1]),.doutc(w_n3955_48[2]),.din(w_n3955_15[2]));
	jspl3 jspl3_w_n3955_49(.douta(w_n3955_49[0]),.doutb(w_n3955_49[1]),.doutc(w_n3955_49[2]),.din(w_n3955_16[0]));
	jspl jspl_w_n3955_50(.douta(w_n3955_50[0]),.doutb(w_n3955_50[1]),.din(w_n3955_16[1]));
	jspl jspl_w_n3957_0(.douta(w_n3957_0[0]),.doutb(w_n3957_0[1]),.din(n3957));
	jspl3 jspl3_w_n3959_0(.douta(w_n3959_0[0]),.doutb(w_n3959_0[1]),.doutc(w_n3959_0[2]),.din(n3959));
	jspl jspl_w_n3960_0(.douta(w_n3960_0[0]),.doutb(w_n3960_0[1]),.din(n3960));
	jspl jspl_w_n3962_0(.douta(w_n3962_0[0]),.doutb(w_n3962_0[1]),.din(n3962));
	jspl jspl_w_n3967_0(.douta(w_n3967_0[0]),.doutb(w_n3967_0[1]),.din(n3967));
	jspl jspl_w_n3968_0(.douta(w_n3968_0[0]),.doutb(w_n3968_0[1]),.din(n3968));
	jspl3 jspl3_w_n3970_0(.douta(w_n3970_0[0]),.doutb(w_n3970_0[1]),.doutc(w_n3970_0[2]),.din(n3970));
	jspl jspl_w_n3971_0(.douta(w_n3971_0[0]),.doutb(w_n3971_0[1]),.din(n3971));
	jspl jspl_w_n3975_0(.douta(w_n3975_0[0]),.doutb(w_n3975_0[1]),.din(n3975));
	jspl3 jspl3_w_n3977_0(.douta(w_n3977_0[0]),.doutb(w_n3977_0[1]),.doutc(w_n3977_0[2]),.din(n3977));
	jspl jspl_w_n3978_0(.douta(w_n3978_0[0]),.doutb(w_n3978_0[1]),.din(n3978));
	jspl jspl_w_n3982_0(.douta(w_n3982_0[0]),.doutb(w_n3982_0[1]),.din(n3982));
	jspl jspl_w_n3983_0(.douta(w_n3983_0[0]),.doutb(w_n3983_0[1]),.din(n3983));
	jspl3 jspl3_w_n3985_0(.douta(w_n3985_0[0]),.doutb(w_n3985_0[1]),.doutc(w_n3985_0[2]),.din(n3985));
	jspl jspl_w_n3986_0(.douta(w_n3986_0[0]),.doutb(w_n3986_0[1]),.din(n3986));
	jspl jspl_w_n3990_0(.douta(w_n3990_0[0]),.doutb(w_n3990_0[1]),.din(n3990));
	jspl3 jspl3_w_n3992_0(.douta(w_n3992_0[0]),.doutb(w_n3992_0[1]),.doutc(w_n3992_0[2]),.din(n3992));
	jspl jspl_w_n3993_0(.douta(w_n3993_0[0]),.doutb(w_n3993_0[1]),.din(n3993));
	jspl jspl_w_n3997_0(.douta(w_n3997_0[0]),.doutb(w_n3997_0[1]),.din(n3997));
	jspl jspl_w_n3998_0(.douta(w_n3998_0[0]),.doutb(w_n3998_0[1]),.din(n3998));
	jspl3 jspl3_w_n4000_0(.douta(w_n4000_0[0]),.doutb(w_n4000_0[1]),.doutc(w_n4000_0[2]),.din(n4000));
	jspl jspl_w_n4001_0(.douta(w_n4001_0[0]),.doutb(w_n4001_0[1]),.din(n4001));
	jspl jspl_w_n4005_0(.douta(w_n4005_0[0]),.doutb(w_n4005_0[1]),.din(n4005));
	jspl3 jspl3_w_n4007_0(.douta(w_n4007_0[0]),.doutb(w_n4007_0[1]),.doutc(w_n4007_0[2]),.din(n4007));
	jspl jspl_w_n4008_0(.douta(w_n4008_0[0]),.doutb(w_n4008_0[1]),.din(n4008));
	jspl jspl_w_n4012_0(.douta(w_n4012_0[0]),.doutb(w_n4012_0[1]),.din(n4012));
	jspl3 jspl3_w_n4014_0(.douta(w_n4014_0[0]),.doutb(w_n4014_0[1]),.doutc(w_n4014_0[2]),.din(n4014));
	jspl jspl_w_n4015_0(.douta(w_n4015_0[0]),.doutb(w_n4015_0[1]),.din(n4015));
	jspl jspl_w_n4019_0(.douta(w_n4019_0[0]),.doutb(w_n4019_0[1]),.din(n4019));
	jspl jspl_w_n4020_0(.douta(w_n4020_0[0]),.doutb(w_n4020_0[1]),.din(n4020));
	jspl3 jspl3_w_n4022_0(.douta(w_n4022_0[0]),.doutb(w_n4022_0[1]),.doutc(w_n4022_0[2]),.din(n4022));
	jspl jspl_w_n4023_0(.douta(w_n4023_0[0]),.doutb(w_n4023_0[1]),.din(n4023));
	jspl jspl_w_n4027_0(.douta(w_n4027_0[0]),.doutb(w_n4027_0[1]),.din(n4027));
	jspl jspl_w_n4028_0(.douta(w_n4028_0[0]),.doutb(w_n4028_0[1]),.din(n4028));
	jspl3 jspl3_w_n4030_0(.douta(w_n4030_0[0]),.doutb(w_n4030_0[1]),.doutc(w_n4030_0[2]),.din(n4030));
	jspl jspl_w_n4031_0(.douta(w_n4031_0[0]),.doutb(w_n4031_0[1]),.din(n4031));
	jspl jspl_w_n4035_0(.douta(w_n4035_0[0]),.doutb(w_n4035_0[1]),.din(n4035));
	jspl3 jspl3_w_n4037_0(.douta(w_n4037_0[0]),.doutb(w_n4037_0[1]),.doutc(w_n4037_0[2]),.din(n4037));
	jspl jspl_w_n4038_0(.douta(w_n4038_0[0]),.doutb(w_n4038_0[1]),.din(n4038));
	jspl jspl_w_n4042_0(.douta(w_n4042_0[0]),.doutb(w_n4042_0[1]),.din(n4042));
	jspl jspl_w_n4043_0(.douta(w_n4043_0[0]),.doutb(w_n4043_0[1]),.din(n4043));
	jspl3 jspl3_w_n4045_0(.douta(w_n4045_0[0]),.doutb(w_n4045_0[1]),.doutc(w_n4045_0[2]),.din(n4045));
	jspl jspl_w_n4046_0(.douta(w_n4046_0[0]),.doutb(w_n4046_0[1]),.din(n4046));
	jspl jspl_w_n4050_0(.douta(w_n4050_0[0]),.doutb(w_n4050_0[1]),.din(n4050));
	jspl3 jspl3_w_n4052_0(.douta(w_n4052_0[0]),.doutb(w_n4052_0[1]),.doutc(w_n4052_0[2]),.din(n4052));
	jspl jspl_w_n4053_0(.douta(w_n4053_0[0]),.doutb(w_n4053_0[1]),.din(n4053));
	jspl jspl_w_n4057_0(.douta(w_n4057_0[0]),.doutb(w_n4057_0[1]),.din(n4057));
	jspl jspl_w_n4058_0(.douta(w_n4058_0[0]),.doutb(w_n4058_0[1]),.din(n4058));
	jspl3 jspl3_w_n4060_0(.douta(w_n4060_0[0]),.doutb(w_n4060_0[1]),.doutc(w_n4060_0[2]),.din(n4060));
	jspl jspl_w_n4061_0(.douta(w_n4061_0[0]),.doutb(w_n4061_0[1]),.din(n4061));
	jspl jspl_w_n4065_0(.douta(w_n4065_0[0]),.doutb(w_n4065_0[1]),.din(n4065));
	jspl3 jspl3_w_n4067_0(.douta(w_n4067_0[0]),.doutb(w_n4067_0[1]),.doutc(w_n4067_0[2]),.din(n4067));
	jspl jspl_w_n4068_0(.douta(w_n4068_0[0]),.doutb(w_n4068_0[1]),.din(n4068));
	jspl jspl_w_n4072_0(.douta(w_n4072_0[0]),.doutb(w_n4072_0[1]),.din(n4072));
	jspl jspl_w_n4073_0(.douta(w_n4073_0[0]),.doutb(w_n4073_0[1]),.din(n4073));
	jspl3 jspl3_w_n4075_0(.douta(w_n4075_0[0]),.doutb(w_n4075_0[1]),.doutc(w_n4075_0[2]),.din(n4075));
	jspl jspl_w_n4076_0(.douta(w_n4076_0[0]),.doutb(w_n4076_0[1]),.din(n4076));
	jspl jspl_w_n4080_0(.douta(w_n4080_0[0]),.doutb(w_n4080_0[1]),.din(n4080));
	jspl3 jspl3_w_n4082_0(.douta(w_n4082_0[0]),.doutb(w_n4082_0[1]),.doutc(w_n4082_0[2]),.din(n4082));
	jspl jspl_w_n4083_0(.douta(w_n4083_0[0]),.doutb(w_n4083_0[1]),.din(n4083));
	jspl jspl_w_n4087_0(.douta(w_n4087_0[0]),.doutb(w_n4087_0[1]),.din(n4087));
	jspl jspl_w_n4088_0(.douta(w_n4088_0[0]),.doutb(w_n4088_0[1]),.din(n4088));
	jspl3 jspl3_w_n4090_0(.douta(w_n4090_0[0]),.doutb(w_n4090_0[1]),.doutc(w_n4090_0[2]),.din(n4090));
	jspl jspl_w_n4091_0(.douta(w_n4091_0[0]),.doutb(w_n4091_0[1]),.din(n4091));
	jspl jspl_w_n4095_0(.douta(w_n4095_0[0]),.doutb(w_n4095_0[1]),.din(n4095));
	jspl3 jspl3_w_n4097_0(.douta(w_n4097_0[0]),.doutb(w_n4097_0[1]),.doutc(w_n4097_0[2]),.din(n4097));
	jspl jspl_w_n4098_0(.douta(w_n4098_0[0]),.doutb(w_n4098_0[1]),.din(n4098));
	jspl jspl_w_n4102_0(.douta(w_n4102_0[0]),.doutb(w_n4102_0[1]),.din(n4102));
	jspl jspl_w_n4103_0(.douta(w_n4103_0[0]),.doutb(w_n4103_0[1]),.din(n4103));
	jspl3 jspl3_w_n4105_0(.douta(w_n4105_0[0]),.doutb(w_n4105_0[1]),.doutc(w_n4105_0[2]),.din(n4105));
	jspl jspl_w_n4106_0(.douta(w_n4106_0[0]),.doutb(w_n4106_0[1]),.din(n4106));
	jspl jspl_w_n4110_0(.douta(w_n4110_0[0]),.doutb(w_n4110_0[1]),.din(n4110));
	jspl jspl_w_n4111_0(.douta(w_n4111_0[0]),.doutb(w_n4111_0[1]),.din(n4111));
	jspl3 jspl3_w_n4113_0(.douta(w_n4113_0[0]),.doutb(w_n4113_0[1]),.doutc(w_n4113_0[2]),.din(n4113));
	jspl jspl_w_n4114_0(.douta(w_n4114_0[0]),.doutb(w_n4114_0[1]),.din(n4114));
	jspl jspl_w_n4150_0(.douta(w_n4150_0[0]),.doutb(w_n4150_0[1]),.din(n4150));
	jspl jspl_w_n4157_0(.douta(w_n4157_0[0]),.doutb(w_n4157_0[1]),.din(n4157));
	jspl jspl_w_n4164_0(.douta(w_n4164_0[0]),.doutb(w_n4164_0[1]),.din(n4164));
	jspl jspl_w_n4168_0(.douta(w_n4168_0[0]),.doutb(w_n4168_0[1]),.din(n4168));
	jspl jspl_w_n4178_0(.douta(w_n4178_0[0]),.doutb(w_n4178_0[1]),.din(n4178));
	jspl jspl_w_n4185_0(.douta(w_n4185_0[0]),.doutb(w_n4185_0[1]),.din(n4185));
	jspl jspl_w_n4192_0(.douta(w_n4192_0[0]),.doutb(w_n4192_0[1]),.din(n4192));
	jspl jspl_w_n4199_0(.douta(w_n4199_0[0]),.doutb(w_n4199_0[1]),.din(n4199));
	jspl jspl_w_n4206_0(.douta(w_n4206_0[0]),.doutb(w_n4206_0[1]),.din(n4206));
	jspl jspl_w_n4218_0(.douta(w_n4218_0[0]),.doutb(w_n4218_0[1]),.din(n4218));
	jspl jspl_w_n4219_0(.douta(w_n4219_0[0]),.doutb(w_n4219_0[1]),.din(n4219));
	jspl3 jspl3_w_n4221_0(.douta(w_n4221_0[0]),.doutb(w_n4221_0[1]),.doutc(w_n4221_0[2]),.din(n4221));
	jspl jspl_w_n4222_0(.douta(w_n4222_0[0]),.doutb(w_n4222_0[1]),.din(n4222));
	jspl jspl_w_n4223_0(.douta(w_n4223_0[0]),.doutb(w_n4223_0[1]),.din(n4223));
	jspl jspl_w_n4225_0(.douta(w_n4225_0[0]),.doutb(w_n4225_0[1]),.din(n4225));
	jspl jspl_w_n4227_0(.douta(w_n4227_0[0]),.doutb(w_n4227_0[1]),.din(n4227));
	jspl jspl_w_n4228_0(.douta(w_n4228_0[0]),.doutb(w_n4228_0[1]),.din(n4228));
	jspl3 jspl3_w_n4229_0(.douta(w_n4229_0[0]),.doutb(w_n4229_0[1]),.doutc(w_n4229_0[2]),.din(n4229));
	jspl jspl_w_n4233_0(.douta(w_n4233_0[0]),.doutb(w_n4233_0[1]),.din(n4233));
	jspl jspl_w_n4234_0(.douta(w_n4234_0[0]),.doutb(w_n4234_0[1]),.din(n4234));
	jspl jspl_w_n4239_0(.douta(w_n4239_0[0]),.doutb(w_n4239_0[1]),.din(n4239));
	jspl jspl_w_n4240_0(.douta(w_n4240_0[0]),.doutb(w_n4240_0[1]),.din(n4240));
	jspl3 jspl3_w_n4245_0(.douta(w_n4245_0[0]),.doutb(w_n4245_0[1]),.doutc(w_n4245_0[2]),.din(n4245));
	jspl3 jspl3_w_n4249_0(.douta(w_n4249_0[0]),.doutb(w_n4249_0[1]),.doutc(w_n4249_0[2]),.din(n4249));
	jspl3 jspl3_w_n4249_1(.douta(w_n4249_1[0]),.doutb(w_n4249_1[1]),.doutc(w_n4249_1[2]),.din(w_n4249_0[0]));
	jspl3 jspl3_w_n4249_2(.douta(w_n4249_2[0]),.doutb(w_n4249_2[1]),.doutc(w_n4249_2[2]),.din(w_n4249_0[1]));
	jspl3 jspl3_w_n4249_3(.douta(w_n4249_3[0]),.doutb(w_n4249_3[1]),.doutc(w_n4249_3[2]),.din(w_n4249_0[2]));
	jspl3 jspl3_w_n4249_4(.douta(w_n4249_4[0]),.doutb(w_n4249_4[1]),.doutc(w_n4249_4[2]),.din(w_n4249_1[0]));
	jspl3 jspl3_w_n4249_5(.douta(w_n4249_5[0]),.doutb(w_n4249_5[1]),.doutc(w_n4249_5[2]),.din(w_n4249_1[1]));
	jspl3 jspl3_w_n4249_6(.douta(w_n4249_6[0]),.doutb(w_n4249_6[1]),.doutc(w_n4249_6[2]),.din(w_n4249_1[2]));
	jspl3 jspl3_w_n4249_7(.douta(w_n4249_7[0]),.doutb(w_n4249_7[1]),.doutc(w_n4249_7[2]),.din(w_n4249_2[0]));
	jspl3 jspl3_w_n4249_8(.douta(w_n4249_8[0]),.doutb(w_n4249_8[1]),.doutc(w_n4249_8[2]),.din(w_n4249_2[1]));
	jspl3 jspl3_w_n4249_9(.douta(w_n4249_9[0]),.doutb(w_n4249_9[1]),.doutc(w_n4249_9[2]),.din(w_n4249_2[2]));
	jspl3 jspl3_w_n4249_10(.douta(w_n4249_10[0]),.doutb(w_n4249_10[1]),.doutc(w_n4249_10[2]),.din(w_n4249_3[0]));
	jspl3 jspl3_w_n4249_11(.douta(w_n4249_11[0]),.doutb(w_n4249_11[1]),.doutc(w_n4249_11[2]),.din(w_n4249_3[1]));
	jspl3 jspl3_w_n4249_12(.douta(w_n4249_12[0]),.doutb(w_n4249_12[1]),.doutc(w_n4249_12[2]),.din(w_n4249_3[2]));
	jspl3 jspl3_w_n4249_13(.douta(w_n4249_13[0]),.doutb(w_n4249_13[1]),.doutc(w_n4249_13[2]),.din(w_n4249_4[0]));
	jspl3 jspl3_w_n4249_14(.douta(w_n4249_14[0]),.doutb(w_n4249_14[1]),.doutc(w_n4249_14[2]),.din(w_n4249_4[1]));
	jspl3 jspl3_w_n4249_15(.douta(w_n4249_15[0]),.doutb(w_n4249_15[1]),.doutc(w_n4249_15[2]),.din(w_n4249_4[2]));
	jspl3 jspl3_w_n4249_16(.douta(w_n4249_16[0]),.doutb(w_n4249_16[1]),.doutc(w_n4249_16[2]),.din(w_n4249_5[0]));
	jspl3 jspl3_w_n4249_17(.douta(w_n4249_17[0]),.doutb(w_n4249_17[1]),.doutc(w_n4249_17[2]),.din(w_n4249_5[1]));
	jspl3 jspl3_w_n4249_18(.douta(w_n4249_18[0]),.doutb(w_n4249_18[1]),.doutc(w_n4249_18[2]),.din(w_n4249_5[2]));
	jspl3 jspl3_w_n4249_19(.douta(w_n4249_19[0]),.doutb(w_n4249_19[1]),.doutc(w_n4249_19[2]),.din(w_n4249_6[0]));
	jspl3 jspl3_w_n4249_20(.douta(w_n4249_20[0]),.doutb(w_n4249_20[1]),.doutc(w_n4249_20[2]),.din(w_n4249_6[1]));
	jspl3 jspl3_w_n4249_21(.douta(w_n4249_21[0]),.doutb(w_n4249_21[1]),.doutc(w_n4249_21[2]),.din(w_n4249_6[2]));
	jspl3 jspl3_w_n4249_22(.douta(w_n4249_22[0]),.doutb(w_n4249_22[1]),.doutc(w_n4249_22[2]),.din(w_n4249_7[0]));
	jspl3 jspl3_w_n4249_23(.douta(w_n4249_23[0]),.doutb(w_n4249_23[1]),.doutc(w_n4249_23[2]),.din(w_n4249_7[1]));
	jspl3 jspl3_w_n4249_24(.douta(w_n4249_24[0]),.doutb(w_n4249_24[1]),.doutc(w_n4249_24[2]),.din(w_n4249_7[2]));
	jspl3 jspl3_w_n4249_25(.douta(w_n4249_25[0]),.doutb(w_n4249_25[1]),.doutc(w_n4249_25[2]),.din(w_n4249_8[0]));
	jspl3 jspl3_w_n4249_26(.douta(w_n4249_26[0]),.doutb(w_n4249_26[1]),.doutc(w_n4249_26[2]),.din(w_n4249_8[1]));
	jspl3 jspl3_w_n4249_27(.douta(w_n4249_27[0]),.doutb(w_n4249_27[1]),.doutc(w_n4249_27[2]),.din(w_n4249_8[2]));
	jspl3 jspl3_w_n4249_28(.douta(w_n4249_28[0]),.doutb(w_n4249_28[1]),.doutc(w_n4249_28[2]),.din(w_n4249_9[0]));
	jspl3 jspl3_w_n4249_29(.douta(w_n4249_29[0]),.doutb(w_n4249_29[1]),.doutc(w_n4249_29[2]),.din(w_n4249_9[1]));
	jspl3 jspl3_w_n4249_30(.douta(w_n4249_30[0]),.doutb(w_n4249_30[1]),.doutc(w_n4249_30[2]),.din(w_n4249_9[2]));
	jspl3 jspl3_w_n4249_31(.douta(w_n4249_31[0]),.doutb(w_n4249_31[1]),.doutc(w_n4249_31[2]),.din(w_n4249_10[0]));
	jspl3 jspl3_w_n4249_32(.douta(w_n4249_32[0]),.doutb(w_n4249_32[1]),.doutc(w_n4249_32[2]),.din(w_n4249_10[1]));
	jspl3 jspl3_w_n4249_33(.douta(w_n4249_33[0]),.doutb(w_n4249_33[1]),.doutc(w_n4249_33[2]),.din(w_n4249_10[2]));
	jspl3 jspl3_w_n4249_34(.douta(w_n4249_34[0]),.doutb(w_n4249_34[1]),.doutc(w_n4249_34[2]),.din(w_n4249_11[0]));
	jspl3 jspl3_w_n4249_35(.douta(w_n4249_35[0]),.doutb(w_n4249_35[1]),.doutc(w_n4249_35[2]),.din(w_n4249_11[1]));
	jspl3 jspl3_w_n4249_36(.douta(w_n4249_36[0]),.doutb(w_n4249_36[1]),.doutc(w_n4249_36[2]),.din(w_n4249_11[2]));
	jspl3 jspl3_w_n4249_37(.douta(w_n4249_37[0]),.doutb(w_n4249_37[1]),.doutc(w_n4249_37[2]),.din(w_n4249_12[0]));
	jspl3 jspl3_w_n4249_38(.douta(w_n4249_38[0]),.doutb(w_n4249_38[1]),.doutc(w_n4249_38[2]),.din(w_n4249_12[1]));
	jspl3 jspl3_w_n4249_39(.douta(w_n4249_39[0]),.doutb(w_n4249_39[1]),.doutc(w_n4249_39[2]),.din(w_n4249_12[2]));
	jspl3 jspl3_w_n4249_40(.douta(w_n4249_40[0]),.doutb(w_n4249_40[1]),.doutc(w_n4249_40[2]),.din(w_n4249_13[0]));
	jspl3 jspl3_w_n4249_41(.douta(w_n4249_41[0]),.doutb(w_n4249_41[1]),.doutc(w_n4249_41[2]),.din(w_n4249_13[1]));
	jspl3 jspl3_w_n4249_42(.douta(w_n4249_42[0]),.doutb(w_n4249_42[1]),.doutc(w_n4249_42[2]),.din(w_n4249_13[2]));
	jspl3 jspl3_w_n4249_43(.douta(w_n4249_43[0]),.doutb(w_n4249_43[1]),.doutc(w_n4249_43[2]),.din(w_n4249_14[0]));
	jspl3 jspl3_w_n4249_44(.douta(w_n4249_44[0]),.doutb(w_n4249_44[1]),.doutc(w_n4249_44[2]),.din(w_n4249_14[1]));
	jspl3 jspl3_w_n4249_45(.douta(w_n4249_45[0]),.doutb(w_n4249_45[1]),.doutc(w_n4249_45[2]),.din(w_n4249_14[2]));
	jspl3 jspl3_w_n4249_46(.douta(w_n4249_46[0]),.doutb(w_n4249_46[1]),.doutc(w_n4249_46[2]),.din(w_n4249_15[0]));
	jspl3 jspl3_w_n4249_47(.douta(w_n4249_47[0]),.doutb(w_n4249_47[1]),.doutc(w_n4249_47[2]),.din(w_n4249_15[1]));
	jspl3 jspl3_w_n4249_48(.douta(w_n4249_48[0]),.doutb(w_n4249_48[1]),.doutc(w_n4249_48[2]),.din(w_n4249_15[2]));
	jspl3 jspl3_w_n4249_49(.douta(w_n4249_49[0]),.doutb(w_n4249_49[1]),.doutc(w_n4249_49[2]),.din(w_n4249_16[0]));
	jspl3 jspl3_w_n4249_50(.douta(w_n4249_50[0]),.doutb(w_n4249_50[1]),.doutc(w_n4249_50[2]),.din(w_n4249_16[1]));
	jspl3 jspl3_w_n4249_51(.douta(w_n4249_51[0]),.doutb(w_n4249_51[1]),.doutc(w_n4249_51[2]),.din(w_n4249_16[2]));
	jspl3 jspl3_w_n4249_52(.douta(w_n4249_52[0]),.doutb(w_n4249_52[1]),.doutc(w_n4249_52[2]),.din(w_n4249_17[0]));
	jspl3 jspl3_w_n4249_53(.douta(w_n4249_53[0]),.doutb(w_n4249_53[1]),.doutc(w_n4249_53[2]),.din(w_n4249_17[1]));
	jspl3 jspl3_w_n4249_54(.douta(w_n4249_54[0]),.doutb(w_n4249_54[1]),.doutc(w_n4249_54[2]),.din(w_n4249_17[2]));
	jspl3 jspl3_w_n4249_55(.douta(w_n4249_55[0]),.doutb(w_n4249_55[1]),.doutc(w_n4249_55[2]),.din(w_n4249_18[0]));
	jspl3 jspl3_w_n4249_56(.douta(w_n4249_56[0]),.doutb(w_n4249_56[1]),.doutc(w_n4249_56[2]),.din(w_n4249_18[1]));
	jspl3 jspl3_w_n4249_57(.douta(w_n4249_57[0]),.doutb(w_n4249_57[1]),.doutc(w_n4249_57[2]),.din(w_n4249_18[2]));
	jspl3 jspl3_w_n4249_58(.douta(w_n4249_58[0]),.doutb(w_n4249_58[1]),.doutc(w_n4249_58[2]),.din(w_n4249_19[0]));
	jspl3 jspl3_w_n4249_59(.douta(w_n4249_59[0]),.doutb(w_n4249_59[1]),.doutc(w_n4249_59[2]),.din(w_n4249_19[1]));
	jspl jspl_w_n4252_0(.douta(w_n4252_0[0]),.doutb(w_n4252_0[1]),.din(n4252));
	jspl3 jspl3_w_n4253_0(.douta(w_n4253_0[0]),.doutb(w_n4253_0[1]),.doutc(w_n4253_0[2]),.din(n4253));
	jspl3 jspl3_w_n4255_0(.douta(w_n4255_0[0]),.doutb(w_n4255_0[1]),.doutc(w_n4255_0[2]),.din(n4255));
	jspl3 jspl3_w_n4255_1(.douta(w_n4255_1[0]),.doutb(w_n4255_1[1]),.doutc(w_n4255_1[2]),.din(w_n4255_0[0]));
	jspl jspl_w_n4256_0(.douta(w_n4256_0[0]),.doutb(w_n4256_0[1]),.din(n4256));
	jspl3 jspl3_w_n4257_0(.douta(w_n4257_0[0]),.doutb(w_n4257_0[1]),.doutc(w_n4257_0[2]),.din(n4257));
	jspl jspl_w_n4258_0(.douta(w_n4258_0[0]),.doutb(w_n4258_0[1]),.din(n4258));
	jspl3 jspl3_w_n4260_0(.douta(w_n4260_0[0]),.doutb(w_n4260_0[1]),.doutc(w_n4260_0[2]),.din(n4260));
	jspl jspl_w_n4261_0(.douta(w_n4261_0[0]),.doutb(w_n4261_0[1]),.din(n4261));
	jspl jspl_w_n4266_0(.douta(w_n4266_0[0]),.doutb(w_n4266_0[1]),.din(n4266));
	jspl3 jspl3_w_n4268_0(.douta(w_n4268_0[0]),.doutb(w_n4268_0[1]),.doutc(w_n4268_0[2]),.din(n4268));
	jspl jspl_w_n4269_0(.douta(w_n4269_0[0]),.doutb(w_n4269_0[1]),.din(n4269));
	jspl jspl_w_n4272_0(.douta(w_n4272_0[0]),.doutb(w_n4272_0[1]),.din(n4272));
	jspl3 jspl3_w_n4277_0(.douta(w_n4277_0[0]),.doutb(w_n4277_0[1]),.doutc(w_n4277_0[2]),.din(n4277));
	jspl3 jspl3_w_n4279_0(.douta(w_n4279_0[0]),.doutb(w_n4279_0[1]),.doutc(w_n4279_0[2]),.din(n4279));
	jspl jspl_w_n4280_0(.douta(w_n4280_0[0]),.doutb(w_n4280_0[1]),.din(n4280));
	jspl3 jspl3_w_n4284_0(.douta(w_n4284_0[0]),.doutb(w_n4284_0[1]),.doutc(w_n4284_0[2]),.din(n4284));
	jspl3 jspl3_w_n4286_0(.douta(w_n4286_0[0]),.doutb(w_n4286_0[1]),.doutc(w_n4286_0[2]),.din(n4286));
	jspl jspl_w_n4287_0(.douta(w_n4287_0[0]),.doutb(w_n4287_0[1]),.din(n4287));
	jspl3 jspl3_w_n4291_0(.douta(w_n4291_0[0]),.doutb(w_n4291_0[1]),.doutc(w_n4291_0[2]),.din(n4291));
	jspl3 jspl3_w_n4293_0(.douta(w_n4293_0[0]),.doutb(w_n4293_0[1]),.doutc(w_n4293_0[2]),.din(n4293));
	jspl jspl_w_n4294_0(.douta(w_n4294_0[0]),.doutb(w_n4294_0[1]),.din(n4294));
	jspl3 jspl3_w_n4298_0(.douta(w_n4298_0[0]),.doutb(w_n4298_0[1]),.doutc(w_n4298_0[2]),.din(n4298));
	jspl3 jspl3_w_n4301_0(.douta(w_n4301_0[0]),.doutb(w_n4301_0[1]),.doutc(w_n4301_0[2]),.din(n4301));
	jspl jspl_w_n4302_0(.douta(w_n4302_0[0]),.doutb(w_n4302_0[1]),.din(n4302));
	jspl3 jspl3_w_n4306_0(.douta(w_n4306_0[0]),.doutb(w_n4306_0[1]),.doutc(w_n4306_0[2]),.din(n4306));
	jspl3 jspl3_w_n4308_0(.douta(w_n4308_0[0]),.doutb(w_n4308_0[1]),.doutc(w_n4308_0[2]),.din(n4308));
	jspl jspl_w_n4309_0(.douta(w_n4309_0[0]),.doutb(w_n4309_0[1]),.din(n4309));
	jspl3 jspl3_w_n4313_0(.douta(w_n4313_0[0]),.doutb(w_n4313_0[1]),.doutc(w_n4313_0[2]),.din(n4313));
	jspl3 jspl3_w_n4316_0(.douta(w_n4316_0[0]),.doutb(w_n4316_0[1]),.doutc(w_n4316_0[2]),.din(n4316));
	jspl jspl_w_n4317_0(.douta(w_n4317_0[0]),.doutb(w_n4317_0[1]),.din(n4317));
	jspl3 jspl3_w_n4321_0(.douta(w_n4321_0[0]),.doutb(w_n4321_0[1]),.doutc(w_n4321_0[2]),.din(n4321));
	jspl3 jspl3_w_n4323_0(.douta(w_n4323_0[0]),.doutb(w_n4323_0[1]),.doutc(w_n4323_0[2]),.din(n4323));
	jspl jspl_w_n4324_0(.douta(w_n4324_0[0]),.doutb(w_n4324_0[1]),.din(n4324));
	jspl3 jspl3_w_n4328_0(.douta(w_n4328_0[0]),.doutb(w_n4328_0[1]),.doutc(w_n4328_0[2]),.din(n4328));
	jspl3 jspl3_w_n4331_0(.douta(w_n4331_0[0]),.doutb(w_n4331_0[1]),.doutc(w_n4331_0[2]),.din(n4331));
	jspl jspl_w_n4332_0(.douta(w_n4332_0[0]),.doutb(w_n4332_0[1]),.din(n4332));
	jspl3 jspl3_w_n4336_0(.douta(w_n4336_0[0]),.doutb(w_n4336_0[1]),.doutc(w_n4336_0[2]),.din(n4336));
	jspl3 jspl3_w_n4339_0(.douta(w_n4339_0[0]),.doutb(w_n4339_0[1]),.doutc(w_n4339_0[2]),.din(n4339));
	jspl jspl_w_n4340_0(.douta(w_n4340_0[0]),.doutb(w_n4340_0[1]),.din(n4340));
	jspl3 jspl3_w_n4344_0(.douta(w_n4344_0[0]),.doutb(w_n4344_0[1]),.doutc(w_n4344_0[2]),.din(n4344));
	jspl3 jspl3_w_n4346_0(.douta(w_n4346_0[0]),.doutb(w_n4346_0[1]),.doutc(w_n4346_0[2]),.din(n4346));
	jspl jspl_w_n4347_0(.douta(w_n4347_0[0]),.doutb(w_n4347_0[1]),.din(n4347));
	jspl3 jspl3_w_n4351_0(.douta(w_n4351_0[0]),.doutb(w_n4351_0[1]),.doutc(w_n4351_0[2]),.din(n4351));
	jspl3 jspl3_w_n4353_0(.douta(w_n4353_0[0]),.doutb(w_n4353_0[1]),.doutc(w_n4353_0[2]),.din(n4353));
	jspl jspl_w_n4354_0(.douta(w_n4354_0[0]),.doutb(w_n4354_0[1]),.din(n4354));
	jspl3 jspl3_w_n4358_0(.douta(w_n4358_0[0]),.doutb(w_n4358_0[1]),.doutc(w_n4358_0[2]),.din(n4358));
	jspl3 jspl3_w_n4361_0(.douta(w_n4361_0[0]),.doutb(w_n4361_0[1]),.doutc(w_n4361_0[2]),.din(n4361));
	jspl jspl_w_n4362_0(.douta(w_n4362_0[0]),.doutb(w_n4362_0[1]),.din(n4362));
	jspl3 jspl3_w_n4366_0(.douta(w_n4366_0[0]),.doutb(w_n4366_0[1]),.doutc(w_n4366_0[2]),.din(n4366));
	jspl3 jspl3_w_n4368_0(.douta(w_n4368_0[0]),.doutb(w_n4368_0[1]),.doutc(w_n4368_0[2]),.din(n4368));
	jspl jspl_w_n4369_0(.douta(w_n4369_0[0]),.doutb(w_n4369_0[1]),.din(n4369));
	jspl3 jspl3_w_n4373_0(.douta(w_n4373_0[0]),.doutb(w_n4373_0[1]),.doutc(w_n4373_0[2]),.din(n4373));
	jspl3 jspl3_w_n4376_0(.douta(w_n4376_0[0]),.doutb(w_n4376_0[1]),.doutc(w_n4376_0[2]),.din(n4376));
	jspl jspl_w_n4377_0(.douta(w_n4377_0[0]),.doutb(w_n4377_0[1]),.din(n4377));
	jspl3 jspl3_w_n4381_0(.douta(w_n4381_0[0]),.doutb(w_n4381_0[1]),.doutc(w_n4381_0[2]),.din(n4381));
	jspl3 jspl3_w_n4383_0(.douta(w_n4383_0[0]),.doutb(w_n4383_0[1]),.doutc(w_n4383_0[2]),.din(n4383));
	jspl jspl_w_n4384_0(.douta(w_n4384_0[0]),.doutb(w_n4384_0[1]),.din(n4384));
	jspl3 jspl3_w_n4388_0(.douta(w_n4388_0[0]),.doutb(w_n4388_0[1]),.doutc(w_n4388_0[2]),.din(n4388));
	jspl3 jspl3_w_n4391_0(.douta(w_n4391_0[0]),.doutb(w_n4391_0[1]),.doutc(w_n4391_0[2]),.din(n4391));
	jspl jspl_w_n4392_0(.douta(w_n4392_0[0]),.doutb(w_n4392_0[1]),.din(n4392));
	jspl3 jspl3_w_n4396_0(.douta(w_n4396_0[0]),.doutb(w_n4396_0[1]),.doutc(w_n4396_0[2]),.din(n4396));
	jspl3 jspl3_w_n4398_0(.douta(w_n4398_0[0]),.doutb(w_n4398_0[1]),.doutc(w_n4398_0[2]),.din(n4398));
	jspl jspl_w_n4399_0(.douta(w_n4399_0[0]),.doutb(w_n4399_0[1]),.din(n4399));
	jspl3 jspl3_w_n4403_0(.douta(w_n4403_0[0]),.doutb(w_n4403_0[1]),.doutc(w_n4403_0[2]),.din(n4403));
	jspl3 jspl3_w_n4406_0(.douta(w_n4406_0[0]),.doutb(w_n4406_0[1]),.doutc(w_n4406_0[2]),.din(n4406));
	jspl jspl_w_n4407_0(.douta(w_n4407_0[0]),.doutb(w_n4407_0[1]),.din(n4407));
	jspl3 jspl3_w_n4411_0(.douta(w_n4411_0[0]),.doutb(w_n4411_0[1]),.doutc(w_n4411_0[2]),.din(n4411));
	jspl3 jspl3_w_n4413_0(.douta(w_n4413_0[0]),.doutb(w_n4413_0[1]),.doutc(w_n4413_0[2]),.din(n4413));
	jspl jspl_w_n4414_0(.douta(w_n4414_0[0]),.doutb(w_n4414_0[1]),.din(n4414));
	jspl3 jspl3_w_n4418_0(.douta(w_n4418_0[0]),.doutb(w_n4418_0[1]),.doutc(w_n4418_0[2]),.din(n4418));
	jspl3 jspl3_w_n4421_0(.douta(w_n4421_0[0]),.doutb(w_n4421_0[1]),.doutc(w_n4421_0[2]),.din(n4421));
	jspl jspl_w_n4422_0(.douta(w_n4422_0[0]),.doutb(w_n4422_0[1]),.din(n4422));
	jspl3 jspl3_w_n4426_0(.douta(w_n4426_0[0]),.doutb(w_n4426_0[1]),.doutc(w_n4426_0[2]),.din(n4426));
	jspl3 jspl3_w_n4428_0(.douta(w_n4428_0[0]),.doutb(w_n4428_0[1]),.doutc(w_n4428_0[2]),.din(n4428));
	jspl jspl_w_n4429_0(.douta(w_n4429_0[0]),.doutb(w_n4429_0[1]),.din(n4429));
	jspl jspl_w_n4433_0(.douta(w_n4433_0[0]),.doutb(w_n4433_0[1]),.din(n4433));
	jspl3 jspl3_w_n4435_0(.douta(w_n4435_0[0]),.doutb(w_n4435_0[1]),.doutc(w_n4435_0[2]),.din(n4435));
	jspl jspl_w_n4436_0(.douta(w_n4436_0[0]),.doutb(w_n4436_0[1]),.din(n4436));
	jspl jspl_w_n4437_0(.douta(w_n4437_0[0]),.doutb(w_n4437_0[1]),.din(n4437));
	jspl3 jspl3_w_n4442_0(.douta(w_n4442_0[0]),.doutb(w_n4442_0[1]),.doutc(w_n4442_0[2]),.din(n4442));
	jspl jspl_w_n4447_0(.douta(w_n4447_0[0]),.doutb(w_n4447_0[1]),.din(n4447));
	jspl jspl_w_n4450_0(.douta(w_n4450_0[0]),.doutb(w_n4450_0[1]),.din(n4450));
	jspl jspl_w_n4452_0(.douta(w_n4452_0[0]),.doutb(w_n4452_0[1]),.din(n4452));
	jspl3 jspl3_w_n4455_0(.douta(w_n4455_0[0]),.doutb(w_n4455_0[1]),.doutc(w_n4455_0[2]),.din(n4455));
	jspl3 jspl3_w_n4457_0(.douta(w_n4457_0[0]),.doutb(w_n4457_0[1]),.doutc(w_n4457_0[2]),.din(n4457));
	jspl jspl_w_n4457_1(.douta(w_n4457_1[0]),.doutb(w_n4457_1[1]),.din(w_n4457_0[0]));
	jspl jspl_w_n4458_0(.douta(w_n4458_0[0]),.doutb(w_n4458_0[1]),.din(n4458));
	jspl3 jspl3_w_n4459_0(.douta(w_n4459_0[0]),.doutb(w_n4459_0[1]),.doutc(w_n4459_0[2]),.din(n4459));
	jspl jspl_w_n4460_0(.douta(w_n4460_0[0]),.doutb(w_n4460_0[1]),.din(n4460));
	jspl3 jspl3_w_n4461_0(.douta(w_n4461_0[0]),.doutb(w_n4461_0[1]),.doutc(w_n4461_0[2]),.din(n4461));
	jspl jspl_w_n4462_0(.douta(w_n4462_0[0]),.doutb(w_n4462_0[1]),.din(n4462));
	jspl jspl_w_n4576_0(.douta(w_n4576_0[0]),.doutb(w_n4576_0[1]),.din(n4576));
	jspl jspl_w_n4580_0(.douta(w_n4580_0[0]),.doutb(w_n4580_0[1]),.din(n4580));
	jspl3 jspl3_w_n4582_0(.douta(w_n4582_0[0]),.doutb(w_n4582_0[1]),.doutc(w_n4582_0[2]),.din(n4582));
	jspl3 jspl3_w_n4582_1(.douta(w_n4582_1[0]),.doutb(w_n4582_1[1]),.doutc(w_n4582_1[2]),.din(w_n4582_0[0]));
	jspl3 jspl3_w_n4582_2(.douta(w_n4582_2[0]),.doutb(w_n4582_2[1]),.doutc(w_n4582_2[2]),.din(w_n4582_0[1]));
	jspl3 jspl3_w_n4582_3(.douta(w_n4582_3[0]),.doutb(w_n4582_3[1]),.doutc(w_n4582_3[2]),.din(w_n4582_0[2]));
	jspl3 jspl3_w_n4582_4(.douta(w_n4582_4[0]),.doutb(w_n4582_4[1]),.doutc(w_n4582_4[2]),.din(w_n4582_1[0]));
	jspl3 jspl3_w_n4582_5(.douta(w_n4582_5[0]),.doutb(w_n4582_5[1]),.doutc(w_n4582_5[2]),.din(w_n4582_1[1]));
	jspl3 jspl3_w_n4582_6(.douta(w_n4582_6[0]),.doutb(w_n4582_6[1]),.doutc(w_n4582_6[2]),.din(w_n4582_1[2]));
	jspl3 jspl3_w_n4582_7(.douta(w_n4582_7[0]),.doutb(w_n4582_7[1]),.doutc(w_n4582_7[2]),.din(w_n4582_2[0]));
	jspl3 jspl3_w_n4582_8(.douta(w_n4582_8[0]),.doutb(w_n4582_8[1]),.doutc(w_n4582_8[2]),.din(w_n4582_2[1]));
	jspl3 jspl3_w_n4582_9(.douta(w_n4582_9[0]),.doutb(w_n4582_9[1]),.doutc(w_n4582_9[2]),.din(w_n4582_2[2]));
	jspl3 jspl3_w_n4582_10(.douta(w_n4582_10[0]),.doutb(w_n4582_10[1]),.doutc(w_n4582_10[2]),.din(w_n4582_3[0]));
	jspl3 jspl3_w_n4582_11(.douta(w_n4582_11[0]),.doutb(w_n4582_11[1]),.doutc(w_n4582_11[2]),.din(w_n4582_3[1]));
	jspl3 jspl3_w_n4582_12(.douta(w_n4582_12[0]),.doutb(w_n4582_12[1]),.doutc(w_n4582_12[2]),.din(w_n4582_3[2]));
	jspl3 jspl3_w_n4582_13(.douta(w_n4582_13[0]),.doutb(w_n4582_13[1]),.doutc(w_n4582_13[2]),.din(w_n4582_4[0]));
	jspl3 jspl3_w_n4582_14(.douta(w_n4582_14[0]),.doutb(w_n4582_14[1]),.doutc(w_n4582_14[2]),.din(w_n4582_4[1]));
	jspl3 jspl3_w_n4582_15(.douta(w_n4582_15[0]),.doutb(w_n4582_15[1]),.doutc(w_n4582_15[2]),.din(w_n4582_4[2]));
	jspl3 jspl3_w_n4582_16(.douta(w_n4582_16[0]),.doutb(w_n4582_16[1]),.doutc(w_n4582_16[2]),.din(w_n4582_5[0]));
	jspl3 jspl3_w_n4582_17(.douta(w_n4582_17[0]),.doutb(w_n4582_17[1]),.doutc(w_n4582_17[2]),.din(w_n4582_5[1]));
	jspl3 jspl3_w_n4582_18(.douta(w_n4582_18[0]),.doutb(w_n4582_18[1]),.doutc(w_n4582_18[2]),.din(w_n4582_5[2]));
	jspl3 jspl3_w_n4582_19(.douta(w_n4582_19[0]),.doutb(w_n4582_19[1]),.doutc(w_n4582_19[2]),.din(w_n4582_6[0]));
	jspl3 jspl3_w_n4582_20(.douta(w_n4582_20[0]),.doutb(w_n4582_20[1]),.doutc(w_n4582_20[2]),.din(w_n4582_6[1]));
	jspl3 jspl3_w_n4582_21(.douta(w_n4582_21[0]),.doutb(w_n4582_21[1]),.doutc(w_n4582_21[2]),.din(w_n4582_6[2]));
	jspl3 jspl3_w_n4582_22(.douta(w_n4582_22[0]),.doutb(w_n4582_22[1]),.doutc(w_n4582_22[2]),.din(w_n4582_7[0]));
	jspl3 jspl3_w_n4582_23(.douta(w_n4582_23[0]),.doutb(w_n4582_23[1]),.doutc(w_n4582_23[2]),.din(w_n4582_7[1]));
	jspl3 jspl3_w_n4582_24(.douta(w_n4582_24[0]),.doutb(w_n4582_24[1]),.doutc(w_n4582_24[2]),.din(w_n4582_7[2]));
	jspl3 jspl3_w_n4582_25(.douta(w_n4582_25[0]),.doutb(w_n4582_25[1]),.doutc(w_n4582_25[2]),.din(w_n4582_8[0]));
	jspl3 jspl3_w_n4582_26(.douta(w_n4582_26[0]),.doutb(w_n4582_26[1]),.doutc(w_n4582_26[2]),.din(w_n4582_8[1]));
	jspl3 jspl3_w_n4582_27(.douta(w_n4582_27[0]),.doutb(w_n4582_27[1]),.doutc(w_n4582_27[2]),.din(w_n4582_8[2]));
	jspl3 jspl3_w_n4582_28(.douta(w_n4582_28[0]),.doutb(w_n4582_28[1]),.doutc(w_n4582_28[2]),.din(w_n4582_9[0]));
	jspl3 jspl3_w_n4582_29(.douta(w_n4582_29[0]),.doutb(w_n4582_29[1]),.doutc(w_n4582_29[2]),.din(w_n4582_9[1]));
	jspl3 jspl3_w_n4582_30(.douta(w_n4582_30[0]),.doutb(w_n4582_30[1]),.doutc(w_n4582_30[2]),.din(w_n4582_9[2]));
	jspl3 jspl3_w_n4582_31(.douta(w_n4582_31[0]),.doutb(w_n4582_31[1]),.doutc(w_n4582_31[2]),.din(w_n4582_10[0]));
	jspl3 jspl3_w_n4582_32(.douta(w_n4582_32[0]),.doutb(w_n4582_32[1]),.doutc(w_n4582_32[2]),.din(w_n4582_10[1]));
	jspl3 jspl3_w_n4582_33(.douta(w_n4582_33[0]),.doutb(w_n4582_33[1]),.doutc(w_n4582_33[2]),.din(w_n4582_10[2]));
	jspl3 jspl3_w_n4582_34(.douta(w_n4582_34[0]),.doutb(w_n4582_34[1]),.doutc(w_n4582_34[2]),.din(w_n4582_11[0]));
	jspl3 jspl3_w_n4582_35(.douta(w_n4582_35[0]),.doutb(w_n4582_35[1]),.doutc(w_n4582_35[2]),.din(w_n4582_11[1]));
	jspl3 jspl3_w_n4582_36(.douta(w_n4582_36[0]),.doutb(w_n4582_36[1]),.doutc(w_n4582_36[2]),.din(w_n4582_11[2]));
	jspl3 jspl3_w_n4582_37(.douta(w_n4582_37[0]),.doutb(w_n4582_37[1]),.doutc(w_n4582_37[2]),.din(w_n4582_12[0]));
	jspl3 jspl3_w_n4582_38(.douta(w_n4582_38[0]),.doutb(w_n4582_38[1]),.doutc(w_n4582_38[2]),.din(w_n4582_12[1]));
	jspl3 jspl3_w_n4582_39(.douta(w_n4582_39[0]),.doutb(w_n4582_39[1]),.doutc(w_n4582_39[2]),.din(w_n4582_12[2]));
	jspl3 jspl3_w_n4582_40(.douta(w_n4582_40[0]),.doutb(w_n4582_40[1]),.doutc(w_n4582_40[2]),.din(w_n4582_13[0]));
	jspl3 jspl3_w_n4582_41(.douta(w_n4582_41[0]),.doutb(w_n4582_41[1]),.doutc(w_n4582_41[2]),.din(w_n4582_13[1]));
	jspl3 jspl3_w_n4582_42(.douta(w_n4582_42[0]),.doutb(w_n4582_42[1]),.doutc(w_n4582_42[2]),.din(w_n4582_13[2]));
	jspl3 jspl3_w_n4582_43(.douta(w_n4582_43[0]),.doutb(w_n4582_43[1]),.doutc(w_n4582_43[2]),.din(w_n4582_14[0]));
	jspl3 jspl3_w_n4582_44(.douta(w_n4582_44[0]),.doutb(w_n4582_44[1]),.doutc(w_n4582_44[2]),.din(w_n4582_14[1]));
	jspl3 jspl3_w_n4582_45(.douta(w_n4582_45[0]),.doutb(w_n4582_45[1]),.doutc(w_n4582_45[2]),.din(w_n4582_14[2]));
	jspl3 jspl3_w_n4582_46(.douta(w_n4582_46[0]),.doutb(w_n4582_46[1]),.doutc(w_n4582_46[2]),.din(w_n4582_15[0]));
	jspl3 jspl3_w_n4582_47(.douta(w_n4582_47[0]),.doutb(w_n4582_47[1]),.doutc(w_n4582_47[2]),.din(w_n4582_15[1]));
	jspl jspl_w_n4582_48(.douta(w_n4582_48[0]),.doutb(w_n4582_48[1]),.din(w_n4582_15[2]));
	jspl3 jspl3_w_n4586_0(.douta(w_n4586_0[0]),.doutb(w_n4586_0[1]),.doutc(w_n4586_0[2]),.din(n4586));
	jspl jspl_w_n4587_0(.douta(w_n4587_0[0]),.doutb(w_n4587_0[1]),.din(n4587));
	jspl jspl_w_n4589_0(.douta(w_n4589_0[0]),.doutb(w_n4589_0[1]),.din(n4589));
	jspl jspl_w_n4590_0(.douta(w_n4590_0[0]),.doutb(w_n4590_0[1]),.din(n4590));
	jspl3 jspl3_w_n4595_0(.douta(w_n4595_0[0]),.doutb(w_n4595_0[1]),.doutc(w_n4595_0[2]),.din(n4595));
	jspl3 jspl3_w_n4598_0(.douta(w_n4598_0[0]),.doutb(w_n4598_0[1]),.doutc(w_n4598_0[2]),.din(n4598));
	jspl jspl_w_n4599_0(.douta(w_n4599_0[0]),.doutb(w_n4599_0[1]),.din(n4599));
	jspl jspl_w_n4603_0(.douta(w_n4603_0[0]),.doutb(w_n4603_0[1]),.din(n4603));
	jspl jspl_w_n4604_0(.douta(w_n4604_0[0]),.doutb(w_n4604_0[1]),.din(n4604));
	jspl3 jspl3_w_n4606_0(.douta(w_n4606_0[0]),.doutb(w_n4606_0[1]),.doutc(w_n4606_0[2]),.din(n4606));
	jspl jspl_w_n4607_0(.douta(w_n4607_0[0]),.doutb(w_n4607_0[1]),.din(n4607));
	jspl jspl_w_n4611_0(.douta(w_n4611_0[0]),.doutb(w_n4611_0[1]),.din(n4611));
	jspl jspl_w_n4612_0(.douta(w_n4612_0[0]),.doutb(w_n4612_0[1]),.din(n4612));
	jspl3 jspl3_w_n4614_0(.douta(w_n4614_0[0]),.doutb(w_n4614_0[1]),.doutc(w_n4614_0[2]),.din(n4614));
	jspl jspl_w_n4615_0(.douta(w_n4615_0[0]),.doutb(w_n4615_0[1]),.din(n4615));
	jspl jspl_w_n4619_0(.douta(w_n4619_0[0]),.doutb(w_n4619_0[1]),.din(n4619));
	jspl jspl_w_n4620_0(.douta(w_n4620_0[0]),.doutb(w_n4620_0[1]),.din(n4620));
	jspl3 jspl3_w_n4622_0(.douta(w_n4622_0[0]),.doutb(w_n4622_0[1]),.doutc(w_n4622_0[2]),.din(n4622));
	jspl jspl_w_n4623_0(.douta(w_n4623_0[0]),.doutb(w_n4623_0[1]),.din(n4623));
	jspl jspl_w_n4627_0(.douta(w_n4627_0[0]),.doutb(w_n4627_0[1]),.din(n4627));
	jspl jspl_w_n4628_0(.douta(w_n4628_0[0]),.doutb(w_n4628_0[1]),.din(n4628));
	jspl3 jspl3_w_n4630_0(.douta(w_n4630_0[0]),.doutb(w_n4630_0[1]),.doutc(w_n4630_0[2]),.din(n4630));
	jspl jspl_w_n4631_0(.douta(w_n4631_0[0]),.doutb(w_n4631_0[1]),.din(n4631));
	jspl jspl_w_n4635_0(.douta(w_n4635_0[0]),.doutb(w_n4635_0[1]),.din(n4635));
	jspl3 jspl3_w_n4637_0(.douta(w_n4637_0[0]),.doutb(w_n4637_0[1]),.doutc(w_n4637_0[2]),.din(n4637));
	jspl jspl_w_n4638_0(.douta(w_n4638_0[0]),.doutb(w_n4638_0[1]),.din(n4638));
	jspl jspl_w_n4642_0(.douta(w_n4642_0[0]),.doutb(w_n4642_0[1]),.din(n4642));
	jspl jspl_w_n4643_0(.douta(w_n4643_0[0]),.doutb(w_n4643_0[1]),.din(n4643));
	jspl3 jspl3_w_n4645_0(.douta(w_n4645_0[0]),.doutb(w_n4645_0[1]),.doutc(w_n4645_0[2]),.din(n4645));
	jspl jspl_w_n4646_0(.douta(w_n4646_0[0]),.doutb(w_n4646_0[1]),.din(n4646));
	jspl jspl_w_n4650_0(.douta(w_n4650_0[0]),.doutb(w_n4650_0[1]),.din(n4650));
	jspl3 jspl3_w_n4652_0(.douta(w_n4652_0[0]),.doutb(w_n4652_0[1]),.doutc(w_n4652_0[2]),.din(n4652));
	jspl jspl_w_n4653_0(.douta(w_n4653_0[0]),.doutb(w_n4653_0[1]),.din(n4653));
	jspl jspl_w_n4657_0(.douta(w_n4657_0[0]),.doutb(w_n4657_0[1]),.din(n4657));
	jspl jspl_w_n4658_0(.douta(w_n4658_0[0]),.doutb(w_n4658_0[1]),.din(n4658));
	jspl3 jspl3_w_n4660_0(.douta(w_n4660_0[0]),.doutb(w_n4660_0[1]),.doutc(w_n4660_0[2]),.din(n4660));
	jspl jspl_w_n4661_0(.douta(w_n4661_0[0]),.doutb(w_n4661_0[1]),.din(n4661));
	jspl jspl_w_n4665_0(.douta(w_n4665_0[0]),.doutb(w_n4665_0[1]),.din(n4665));
	jspl3 jspl3_w_n4667_0(.douta(w_n4667_0[0]),.doutb(w_n4667_0[1]),.doutc(w_n4667_0[2]),.din(n4667));
	jspl jspl_w_n4668_0(.douta(w_n4668_0[0]),.doutb(w_n4668_0[1]),.din(n4668));
	jspl jspl_w_n4672_0(.douta(w_n4672_0[0]),.doutb(w_n4672_0[1]),.din(n4672));
	jspl3 jspl3_w_n4674_0(.douta(w_n4674_0[0]),.doutb(w_n4674_0[1]),.doutc(w_n4674_0[2]),.din(n4674));
	jspl jspl_w_n4675_0(.douta(w_n4675_0[0]),.doutb(w_n4675_0[1]),.din(n4675));
	jspl jspl_w_n4679_0(.douta(w_n4679_0[0]),.doutb(w_n4679_0[1]),.din(n4679));
	jspl jspl_w_n4680_0(.douta(w_n4680_0[0]),.doutb(w_n4680_0[1]),.din(n4680));
	jspl3 jspl3_w_n4682_0(.douta(w_n4682_0[0]),.doutb(w_n4682_0[1]),.doutc(w_n4682_0[2]),.din(n4682));
	jspl jspl_w_n4683_0(.douta(w_n4683_0[0]),.doutb(w_n4683_0[1]),.din(n4683));
	jspl jspl_w_n4687_0(.douta(w_n4687_0[0]),.doutb(w_n4687_0[1]),.din(n4687));
	jspl jspl_w_n4688_0(.douta(w_n4688_0[0]),.doutb(w_n4688_0[1]),.din(n4688));
	jspl3 jspl3_w_n4690_0(.douta(w_n4690_0[0]),.doutb(w_n4690_0[1]),.doutc(w_n4690_0[2]),.din(n4690));
	jspl jspl_w_n4691_0(.douta(w_n4691_0[0]),.doutb(w_n4691_0[1]),.din(n4691));
	jspl jspl_w_n4695_0(.douta(w_n4695_0[0]),.doutb(w_n4695_0[1]),.din(n4695));
	jspl3 jspl3_w_n4697_0(.douta(w_n4697_0[0]),.doutb(w_n4697_0[1]),.doutc(w_n4697_0[2]),.din(n4697));
	jspl jspl_w_n4698_0(.douta(w_n4698_0[0]),.doutb(w_n4698_0[1]),.din(n4698));
	jspl jspl_w_n4702_0(.douta(w_n4702_0[0]),.doutb(w_n4702_0[1]),.din(n4702));
	jspl jspl_w_n4703_0(.douta(w_n4703_0[0]),.doutb(w_n4703_0[1]),.din(n4703));
	jspl3 jspl3_w_n4705_0(.douta(w_n4705_0[0]),.doutb(w_n4705_0[1]),.doutc(w_n4705_0[2]),.din(n4705));
	jspl jspl_w_n4706_0(.douta(w_n4706_0[0]),.doutb(w_n4706_0[1]),.din(n4706));
	jspl jspl_w_n4710_0(.douta(w_n4710_0[0]),.doutb(w_n4710_0[1]),.din(n4710));
	jspl3 jspl3_w_n4712_0(.douta(w_n4712_0[0]),.doutb(w_n4712_0[1]),.doutc(w_n4712_0[2]),.din(n4712));
	jspl jspl_w_n4713_0(.douta(w_n4713_0[0]),.doutb(w_n4713_0[1]),.din(n4713));
	jspl jspl_w_n4717_0(.douta(w_n4717_0[0]),.doutb(w_n4717_0[1]),.din(n4717));
	jspl jspl_w_n4718_0(.douta(w_n4718_0[0]),.doutb(w_n4718_0[1]),.din(n4718));
	jspl3 jspl3_w_n4720_0(.douta(w_n4720_0[0]),.doutb(w_n4720_0[1]),.doutc(w_n4720_0[2]),.din(n4720));
	jspl jspl_w_n4721_0(.douta(w_n4721_0[0]),.doutb(w_n4721_0[1]),.din(n4721));
	jspl jspl_w_n4725_0(.douta(w_n4725_0[0]),.doutb(w_n4725_0[1]),.din(n4725));
	jspl3 jspl3_w_n4727_0(.douta(w_n4727_0[0]),.doutb(w_n4727_0[1]),.doutc(w_n4727_0[2]),.din(n4727));
	jspl jspl_w_n4728_0(.douta(w_n4728_0[0]),.doutb(w_n4728_0[1]),.din(n4728));
	jspl jspl_w_n4732_0(.douta(w_n4732_0[0]),.doutb(w_n4732_0[1]),.din(n4732));
	jspl jspl_w_n4733_0(.douta(w_n4733_0[0]),.doutb(w_n4733_0[1]),.din(n4733));
	jspl3 jspl3_w_n4735_0(.douta(w_n4735_0[0]),.doutb(w_n4735_0[1]),.doutc(w_n4735_0[2]),.din(n4735));
	jspl jspl_w_n4736_0(.douta(w_n4736_0[0]),.doutb(w_n4736_0[1]),.din(n4736));
	jspl jspl_w_n4740_0(.douta(w_n4740_0[0]),.doutb(w_n4740_0[1]),.din(n4740));
	jspl3 jspl3_w_n4742_0(.douta(w_n4742_0[0]),.doutb(w_n4742_0[1]),.doutc(w_n4742_0[2]),.din(n4742));
	jspl jspl_w_n4743_0(.douta(w_n4743_0[0]),.doutb(w_n4743_0[1]),.din(n4743));
	jspl jspl_w_n4747_0(.douta(w_n4747_0[0]),.doutb(w_n4747_0[1]),.din(n4747));
	jspl jspl_w_n4748_0(.douta(w_n4748_0[0]),.doutb(w_n4748_0[1]),.din(n4748));
	jspl3 jspl3_w_n4750_0(.douta(w_n4750_0[0]),.doutb(w_n4750_0[1]),.doutc(w_n4750_0[2]),.din(n4750));
	jspl jspl_w_n4751_0(.douta(w_n4751_0[0]),.doutb(w_n4751_0[1]),.din(n4751));
	jspl jspl_w_n4755_0(.douta(w_n4755_0[0]),.doutb(w_n4755_0[1]),.din(n4755));
	jspl3 jspl3_w_n4757_0(.douta(w_n4757_0[0]),.doutb(w_n4757_0[1]),.doutc(w_n4757_0[2]),.din(n4757));
	jspl jspl_w_n4758_0(.douta(w_n4758_0[0]),.doutb(w_n4758_0[1]),.din(n4758));
	jspl3 jspl3_w_n4762_0(.douta(w_n4762_0[0]),.doutb(w_n4762_0[1]),.doutc(w_n4762_0[2]),.din(n4762));
	jspl jspl_w_n4765_0(.douta(w_n4765_0[0]),.doutb(w_n4765_0[1]),.din(n4765));
	jspl3 jspl3_w_n4766_0(.douta(w_n4766_0[0]),.doutb(w_n4766_0[1]),.doutc(w_n4766_0[2]),.din(n4766));
	jspl jspl_w_n4766_1(.douta(w_n4766_1[0]),.doutb(w_n4766_1[1]),.din(w_n4766_0[0]));
	jspl3 jspl3_w_n4767_0(.douta(w_n4767_0[0]),.doutb(w_n4767_0[1]),.doutc(w_n4767_0[2]),.din(n4767));
	jspl jspl_w_n4771_0(.douta(w_n4771_0[0]),.doutb(w_n4771_0[1]),.din(n4771));
	jspl jspl_w_n4772_0(.douta(w_n4772_0[0]),.doutb(w_n4772_0[1]),.din(n4772));
	jspl jspl_w_n4804_0(.douta(w_n4804_0[0]),.doutb(w_n4804_0[1]),.din(n4804));
	jspl jspl_w_n4823_0(.douta(w_n4823_0[0]),.doutb(w_n4823_0[1]),.din(n4823));
	jspl jspl_w_n4830_0(.douta(w_n4830_0[0]),.doutb(w_n4830_0[1]),.din(n4830));
	jspl jspl_w_n4837_0(.douta(w_n4837_0[0]),.doutb(w_n4837_0[1]),.din(n4837));
	jspl jspl_w_n4841_0(.douta(w_n4841_0[0]),.doutb(w_n4841_0[1]),.din(n4841));
	jspl jspl_w_n4851_0(.douta(w_n4851_0[0]),.doutb(w_n4851_0[1]),.din(n4851));
	jspl jspl_w_n4858_0(.douta(w_n4858_0[0]),.doutb(w_n4858_0[1]),.din(n4858));
	jspl jspl_w_n4865_0(.douta(w_n4865_0[0]),.doutb(w_n4865_0[1]),.din(n4865));
	jspl jspl_w_n4872_0(.douta(w_n4872_0[0]),.doutb(w_n4872_0[1]),.din(n4872));
	jspl jspl_w_n4879_0(.douta(w_n4879_0[0]),.doutb(w_n4879_0[1]),.din(n4879));
	jspl jspl_w_n4884_0(.douta(w_n4884_0[0]),.doutb(w_n4884_0[1]),.din(n4884));
	jspl jspl_w_n4885_0(.douta(w_n4885_0[0]),.doutb(w_n4885_0[1]),.din(n4885));
	jspl jspl_w_n4887_0(.douta(w_n4887_0[0]),.doutb(w_n4887_0[1]),.din(n4887));
	jspl jspl_w_n4889_0(.douta(w_n4889_0[0]),.doutb(w_n4889_0[1]),.din(n4889));
	jspl jspl_w_n4890_0(.douta(w_n4890_0[0]),.doutb(w_n4890_0[1]),.din(n4890));
	jspl jspl_w_n4892_0(.douta(w_n4892_0[0]),.doutb(w_n4892_0[1]),.din(n4892));
	jspl jspl_w_n4895_0(.douta(w_n4895_0[0]),.doutb(w_n4895_0[1]),.din(n4895));
	jspl jspl_w_n4901_0(.douta(w_n4901_0[0]),.doutb(w_n4901_0[1]),.din(n4901));
	jspl3 jspl3_w_n4902_0(.douta(w_n4902_0[0]),.doutb(w_n4902_0[1]),.doutc(w_n4902_0[2]),.din(n4902));
	jspl3 jspl3_w_n4902_1(.douta(w_n4902_1[0]),.doutb(w_n4902_1[1]),.doutc(w_n4902_1[2]),.din(w_n4902_0[0]));
	jspl3 jspl3_w_n4902_2(.douta(w_n4902_2[0]),.doutb(w_n4902_2[1]),.doutc(w_n4902_2[2]),.din(w_n4902_0[1]));
	jspl3 jspl3_w_n4902_3(.douta(w_n4902_3[0]),.doutb(w_n4902_3[1]),.doutc(w_n4902_3[2]),.din(w_n4902_0[2]));
	jspl3 jspl3_w_n4902_4(.douta(w_n4902_4[0]),.doutb(w_n4902_4[1]),.doutc(w_n4902_4[2]),.din(w_n4902_1[0]));
	jspl3 jspl3_w_n4902_5(.douta(w_n4902_5[0]),.doutb(w_n4902_5[1]),.doutc(w_n4902_5[2]),.din(w_n4902_1[1]));
	jspl3 jspl3_w_n4902_6(.douta(w_n4902_6[0]),.doutb(w_n4902_6[1]),.doutc(w_n4902_6[2]),.din(w_n4902_1[2]));
	jspl3 jspl3_w_n4902_7(.douta(w_n4902_7[0]),.doutb(w_n4902_7[1]),.doutc(w_n4902_7[2]),.din(w_n4902_2[0]));
	jspl3 jspl3_w_n4902_8(.douta(w_n4902_8[0]),.doutb(w_n4902_8[1]),.doutc(w_n4902_8[2]),.din(w_n4902_2[1]));
	jspl3 jspl3_w_n4902_9(.douta(w_n4902_9[0]),.doutb(w_n4902_9[1]),.doutc(w_n4902_9[2]),.din(w_n4902_2[2]));
	jspl3 jspl3_w_n4902_10(.douta(w_n4902_10[0]),.doutb(w_n4902_10[1]),.doutc(w_n4902_10[2]),.din(w_n4902_3[0]));
	jspl3 jspl3_w_n4902_11(.douta(w_n4902_11[0]),.doutb(w_n4902_11[1]),.doutc(w_n4902_11[2]),.din(w_n4902_3[1]));
	jspl3 jspl3_w_n4902_12(.douta(w_n4902_12[0]),.doutb(w_n4902_12[1]),.doutc(w_n4902_12[2]),.din(w_n4902_3[2]));
	jspl3 jspl3_w_n4902_13(.douta(w_n4902_13[0]),.doutb(w_n4902_13[1]),.doutc(w_n4902_13[2]),.din(w_n4902_4[0]));
	jspl3 jspl3_w_n4902_14(.douta(w_n4902_14[0]),.doutb(w_n4902_14[1]),.doutc(w_n4902_14[2]),.din(w_n4902_4[1]));
	jspl3 jspl3_w_n4902_15(.douta(w_n4902_15[0]),.doutb(w_n4902_15[1]),.doutc(w_n4902_15[2]),.din(w_n4902_4[2]));
	jspl3 jspl3_w_n4902_16(.douta(w_n4902_16[0]),.doutb(w_n4902_16[1]),.doutc(w_n4902_16[2]),.din(w_n4902_5[0]));
	jspl3 jspl3_w_n4902_17(.douta(w_n4902_17[0]),.doutb(w_n4902_17[1]),.doutc(w_n4902_17[2]),.din(w_n4902_5[1]));
	jspl3 jspl3_w_n4902_18(.douta(w_n4902_18[0]),.doutb(w_n4902_18[1]),.doutc(w_n4902_18[2]),.din(w_n4902_5[2]));
	jspl3 jspl3_w_n4902_19(.douta(w_n4902_19[0]),.doutb(w_n4902_19[1]),.doutc(w_n4902_19[2]),.din(w_n4902_6[0]));
	jspl3 jspl3_w_n4902_20(.douta(w_n4902_20[0]),.doutb(w_n4902_20[1]),.doutc(w_n4902_20[2]),.din(w_n4902_6[1]));
	jspl3 jspl3_w_n4902_21(.douta(w_n4902_21[0]),.doutb(w_n4902_21[1]),.doutc(w_n4902_21[2]),.din(w_n4902_6[2]));
	jspl3 jspl3_w_n4902_22(.douta(w_n4902_22[0]),.doutb(w_n4902_22[1]),.doutc(w_n4902_22[2]),.din(w_n4902_7[0]));
	jspl3 jspl3_w_n4902_23(.douta(w_n4902_23[0]),.doutb(w_n4902_23[1]),.doutc(w_n4902_23[2]),.din(w_n4902_7[1]));
	jspl3 jspl3_w_n4902_24(.douta(w_n4902_24[0]),.doutb(w_n4902_24[1]),.doutc(w_n4902_24[2]),.din(w_n4902_7[2]));
	jspl3 jspl3_w_n4902_25(.douta(w_n4902_25[0]),.doutb(w_n4902_25[1]),.doutc(w_n4902_25[2]),.din(w_n4902_8[0]));
	jspl3 jspl3_w_n4902_26(.douta(w_n4902_26[0]),.doutb(w_n4902_26[1]),.doutc(w_n4902_26[2]),.din(w_n4902_8[1]));
	jspl3 jspl3_w_n4902_27(.douta(w_n4902_27[0]),.doutb(w_n4902_27[1]),.doutc(w_n4902_27[2]),.din(w_n4902_8[2]));
	jspl3 jspl3_w_n4902_28(.douta(w_n4902_28[0]),.doutb(w_n4902_28[1]),.doutc(w_n4902_28[2]),.din(w_n4902_9[0]));
	jspl3 jspl3_w_n4902_29(.douta(w_n4902_29[0]),.doutb(w_n4902_29[1]),.doutc(w_n4902_29[2]),.din(w_n4902_9[1]));
	jspl3 jspl3_w_n4902_30(.douta(w_n4902_30[0]),.doutb(w_n4902_30[1]),.doutc(w_n4902_30[2]),.din(w_n4902_9[2]));
	jspl3 jspl3_w_n4902_31(.douta(w_n4902_31[0]),.doutb(w_n4902_31[1]),.doutc(w_n4902_31[2]),.din(w_n4902_10[0]));
	jspl3 jspl3_w_n4902_32(.douta(w_n4902_32[0]),.doutb(w_n4902_32[1]),.doutc(w_n4902_32[2]),.din(w_n4902_10[1]));
	jspl3 jspl3_w_n4902_33(.douta(w_n4902_33[0]),.doutb(w_n4902_33[1]),.doutc(w_n4902_33[2]),.din(w_n4902_10[2]));
	jspl3 jspl3_w_n4902_34(.douta(w_n4902_34[0]),.doutb(w_n4902_34[1]),.doutc(w_n4902_34[2]),.din(w_n4902_11[0]));
	jspl3 jspl3_w_n4902_35(.douta(w_n4902_35[0]),.doutb(w_n4902_35[1]),.doutc(w_n4902_35[2]),.din(w_n4902_11[1]));
	jspl3 jspl3_w_n4902_36(.douta(w_n4902_36[0]),.doutb(w_n4902_36[1]),.doutc(w_n4902_36[2]),.din(w_n4902_11[2]));
	jspl3 jspl3_w_n4902_37(.douta(w_n4902_37[0]),.doutb(w_n4902_37[1]),.doutc(w_n4902_37[2]),.din(w_n4902_12[0]));
	jspl3 jspl3_w_n4902_38(.douta(w_n4902_38[0]),.doutb(w_n4902_38[1]),.doutc(w_n4902_38[2]),.din(w_n4902_12[1]));
	jspl3 jspl3_w_n4902_39(.douta(w_n4902_39[0]),.doutb(w_n4902_39[1]),.doutc(w_n4902_39[2]),.din(w_n4902_12[2]));
	jspl3 jspl3_w_n4902_40(.douta(w_n4902_40[0]),.doutb(w_n4902_40[1]),.doutc(w_n4902_40[2]),.din(w_n4902_13[0]));
	jspl3 jspl3_w_n4902_41(.douta(w_n4902_41[0]),.doutb(w_n4902_41[1]),.doutc(w_n4902_41[2]),.din(w_n4902_13[1]));
	jspl3 jspl3_w_n4902_42(.douta(w_n4902_42[0]),.doutb(w_n4902_42[1]),.doutc(w_n4902_42[2]),.din(w_n4902_13[2]));
	jspl3 jspl3_w_n4902_43(.douta(w_n4902_43[0]),.doutb(w_n4902_43[1]),.doutc(w_n4902_43[2]),.din(w_n4902_14[0]));
	jspl3 jspl3_w_n4902_44(.douta(w_n4902_44[0]),.doutb(w_n4902_44[1]),.doutc(w_n4902_44[2]),.din(w_n4902_14[1]));
	jspl3 jspl3_w_n4902_45(.douta(w_n4902_45[0]),.doutb(w_n4902_45[1]),.doutc(w_n4902_45[2]),.din(w_n4902_14[2]));
	jspl3 jspl3_w_n4902_46(.douta(w_n4902_46[0]),.doutb(w_n4902_46[1]),.doutc(w_n4902_46[2]),.din(w_n4902_15[0]));
	jspl3 jspl3_w_n4902_47(.douta(w_n4902_47[0]),.doutb(w_n4902_47[1]),.doutc(w_n4902_47[2]),.din(w_n4902_15[1]));
	jspl3 jspl3_w_n4902_48(.douta(w_n4902_48[0]),.doutb(w_n4902_48[1]),.doutc(w_n4902_48[2]),.din(w_n4902_15[2]));
	jspl3 jspl3_w_n4902_49(.douta(w_n4902_49[0]),.doutb(w_n4902_49[1]),.doutc(w_n4902_49[2]),.din(w_n4902_16[0]));
	jspl3 jspl3_w_n4902_50(.douta(w_n4902_50[0]),.doutb(w_n4902_50[1]),.doutc(w_n4902_50[2]),.din(w_n4902_16[1]));
	jspl3 jspl3_w_n4902_51(.douta(w_n4902_51[0]),.doutb(w_n4902_51[1]),.doutc(w_n4902_51[2]),.din(w_n4902_16[2]));
	jspl3 jspl3_w_n4902_52(.douta(w_n4902_52[0]),.doutb(w_n4902_52[1]),.doutc(w_n4902_52[2]),.din(w_n4902_17[0]));
	jspl3 jspl3_w_n4902_53(.douta(w_n4902_53[0]),.doutb(w_n4902_53[1]),.doutc(w_n4902_53[2]),.din(w_n4902_17[1]));
	jspl3 jspl3_w_n4902_54(.douta(w_n4902_54[0]),.doutb(w_n4902_54[1]),.doutc(w_n4902_54[2]),.din(w_n4902_17[2]));
	jspl3 jspl3_w_n4902_55(.douta(w_n4902_55[0]),.doutb(w_n4902_55[1]),.doutc(w_n4902_55[2]),.din(w_n4902_18[0]));
	jspl3 jspl3_w_n4902_56(.douta(w_n4902_56[0]),.doutb(w_n4902_56[1]),.doutc(w_n4902_56[2]),.din(w_n4902_18[1]));
	jspl jspl_w_n4902_57(.douta(w_n4902_57[0]),.doutb(w_n4902_57[1]),.din(w_n4902_18[2]));
	jspl jspl_w_n4905_0(.douta(w_n4905_0[0]),.doutb(w_n4905_0[1]),.din(n4905));
	jspl3 jspl3_w_n4906_0(.douta(w_n4906_0[0]),.doutb(w_n4906_0[1]),.doutc(w_n4906_0[2]),.din(n4906));
	jspl3 jspl3_w_n4908_0(.douta(w_n4908_0[0]),.doutb(w_n4908_0[1]),.doutc(w_n4908_0[2]),.din(n4908));
	jspl3 jspl3_w_n4908_1(.douta(w_n4908_1[0]),.doutb(w_n4908_1[1]),.doutc(w_n4908_1[2]),.din(w_n4908_0[0]));
	jspl jspl_w_n4909_0(.douta(w_n4909_0[0]),.doutb(w_n4909_0[1]),.din(n4909));
	jspl3 jspl3_w_n4910_0(.douta(w_n4910_0[0]),.doutb(w_n4910_0[1]),.doutc(w_n4910_0[2]),.din(n4910));
	jspl jspl_w_n4911_0(.douta(w_n4911_0[0]),.doutb(w_n4911_0[1]),.din(n4911));
	jspl3 jspl3_w_n4913_0(.douta(w_n4913_0[0]),.doutb(w_n4913_0[1]),.doutc(w_n4913_0[2]),.din(n4913));
	jspl jspl_w_n4914_0(.douta(w_n4914_0[0]),.doutb(w_n4914_0[1]),.din(n4914));
	jspl3 jspl3_w_n4921_0(.douta(w_n4921_0[0]),.doutb(w_n4921_0[1]),.doutc(w_n4921_0[2]),.din(n4921));
	jspl jspl_w_n4922_0(.douta(w_n4922_0[0]),.doutb(w_n4922_0[1]),.din(n4922));
	jspl jspl_w_n4925_0(.douta(w_n4925_0[0]),.doutb(w_n4925_0[1]),.din(n4925));
	jspl3 jspl3_w_n4930_0(.douta(w_n4930_0[0]),.doutb(w_n4930_0[1]),.doutc(w_n4930_0[2]),.din(n4930));
	jspl3 jspl3_w_n4932_0(.douta(w_n4932_0[0]),.doutb(w_n4932_0[1]),.doutc(w_n4932_0[2]),.din(n4932));
	jspl jspl_w_n4933_0(.douta(w_n4933_0[0]),.doutb(w_n4933_0[1]),.din(n4933));
	jspl3 jspl3_w_n4937_0(.douta(w_n4937_0[0]),.doutb(w_n4937_0[1]),.doutc(w_n4937_0[2]),.din(n4937));
	jspl3 jspl3_w_n4940_0(.douta(w_n4940_0[0]),.doutb(w_n4940_0[1]),.doutc(w_n4940_0[2]),.din(n4940));
	jspl jspl_w_n4941_0(.douta(w_n4941_0[0]),.doutb(w_n4941_0[1]),.din(n4941));
	jspl3 jspl3_w_n4945_0(.douta(w_n4945_0[0]),.doutb(w_n4945_0[1]),.doutc(w_n4945_0[2]),.din(n4945));
	jspl3 jspl3_w_n4948_0(.douta(w_n4948_0[0]),.doutb(w_n4948_0[1]),.doutc(w_n4948_0[2]),.din(n4948));
	jspl jspl_w_n4949_0(.douta(w_n4949_0[0]),.doutb(w_n4949_0[1]),.din(n4949));
	jspl jspl_w_n4953_0(.douta(w_n4953_0[0]),.doutb(w_n4953_0[1]),.din(n4953));
	jspl3 jspl3_w_n4955_0(.douta(w_n4955_0[0]),.doutb(w_n4955_0[1]),.doutc(w_n4955_0[2]),.din(n4955));
	jspl jspl_w_n4956_0(.douta(w_n4956_0[0]),.doutb(w_n4956_0[1]),.din(n4956));
	jspl3 jspl3_w_n4960_0(.douta(w_n4960_0[0]),.doutb(w_n4960_0[1]),.doutc(w_n4960_0[2]),.din(n4960));
	jspl3 jspl3_w_n4962_0(.douta(w_n4962_0[0]),.doutb(w_n4962_0[1]),.doutc(w_n4962_0[2]),.din(n4962));
	jspl jspl_w_n4963_0(.douta(w_n4963_0[0]),.doutb(w_n4963_0[1]),.din(n4963));
	jspl3 jspl3_w_n4967_0(.douta(w_n4967_0[0]),.doutb(w_n4967_0[1]),.doutc(w_n4967_0[2]),.din(n4967));
	jspl3 jspl3_w_n4969_0(.douta(w_n4969_0[0]),.doutb(w_n4969_0[1]),.doutc(w_n4969_0[2]),.din(n4969));
	jspl jspl_w_n4970_0(.douta(w_n4970_0[0]),.doutb(w_n4970_0[1]),.din(n4970));
	jspl3 jspl3_w_n4974_0(.douta(w_n4974_0[0]),.doutb(w_n4974_0[1]),.doutc(w_n4974_0[2]),.din(n4974));
	jspl3 jspl3_w_n4976_0(.douta(w_n4976_0[0]),.doutb(w_n4976_0[1]),.doutc(w_n4976_0[2]),.din(n4976));
	jspl jspl_w_n4977_0(.douta(w_n4977_0[0]),.doutb(w_n4977_0[1]),.din(n4977));
	jspl3 jspl3_w_n4981_0(.douta(w_n4981_0[0]),.doutb(w_n4981_0[1]),.doutc(w_n4981_0[2]),.din(n4981));
	jspl3 jspl3_w_n4984_0(.douta(w_n4984_0[0]),.doutb(w_n4984_0[1]),.doutc(w_n4984_0[2]),.din(n4984));
	jspl jspl_w_n4985_0(.douta(w_n4985_0[0]),.doutb(w_n4985_0[1]),.din(n4985));
	jspl3 jspl3_w_n4989_0(.douta(w_n4989_0[0]),.doutb(w_n4989_0[1]),.doutc(w_n4989_0[2]),.din(n4989));
	jspl3 jspl3_w_n4991_0(.douta(w_n4991_0[0]),.doutb(w_n4991_0[1]),.doutc(w_n4991_0[2]),.din(n4991));
	jspl jspl_w_n4992_0(.douta(w_n4992_0[0]),.doutb(w_n4992_0[1]),.din(n4992));
	jspl3 jspl3_w_n4996_0(.douta(w_n4996_0[0]),.doutb(w_n4996_0[1]),.doutc(w_n4996_0[2]),.din(n4996));
	jspl3 jspl3_w_n4999_0(.douta(w_n4999_0[0]),.doutb(w_n4999_0[1]),.doutc(w_n4999_0[2]),.din(n4999));
	jspl jspl_w_n5000_0(.douta(w_n5000_0[0]),.doutb(w_n5000_0[1]),.din(n5000));
	jspl3 jspl3_w_n5004_0(.douta(w_n5004_0[0]),.doutb(w_n5004_0[1]),.doutc(w_n5004_0[2]),.din(n5004));
	jspl3 jspl3_w_n5006_0(.douta(w_n5006_0[0]),.doutb(w_n5006_0[1]),.doutc(w_n5006_0[2]),.din(n5006));
	jspl jspl_w_n5007_0(.douta(w_n5007_0[0]),.doutb(w_n5007_0[1]),.din(n5007));
	jspl3 jspl3_w_n5011_0(.douta(w_n5011_0[0]),.doutb(w_n5011_0[1]),.doutc(w_n5011_0[2]),.din(n5011));
	jspl3 jspl3_w_n5014_0(.douta(w_n5014_0[0]),.doutb(w_n5014_0[1]),.doutc(w_n5014_0[2]),.din(n5014));
	jspl jspl_w_n5015_0(.douta(w_n5015_0[0]),.doutb(w_n5015_0[1]),.din(n5015));
	jspl3 jspl3_w_n5019_0(.douta(w_n5019_0[0]),.doutb(w_n5019_0[1]),.doutc(w_n5019_0[2]),.din(n5019));
	jspl3 jspl3_w_n5022_0(.douta(w_n5022_0[0]),.doutb(w_n5022_0[1]),.doutc(w_n5022_0[2]),.din(n5022));
	jspl jspl_w_n5023_0(.douta(w_n5023_0[0]),.doutb(w_n5023_0[1]),.din(n5023));
	jspl3 jspl3_w_n5027_0(.douta(w_n5027_0[0]),.doutb(w_n5027_0[1]),.doutc(w_n5027_0[2]),.din(n5027));
	jspl3 jspl3_w_n5029_0(.douta(w_n5029_0[0]),.doutb(w_n5029_0[1]),.doutc(w_n5029_0[2]),.din(n5029));
	jspl jspl_w_n5030_0(.douta(w_n5030_0[0]),.doutb(w_n5030_0[1]),.din(n5030));
	jspl3 jspl3_w_n5034_0(.douta(w_n5034_0[0]),.doutb(w_n5034_0[1]),.doutc(w_n5034_0[2]),.din(n5034));
	jspl3 jspl3_w_n5036_0(.douta(w_n5036_0[0]),.doutb(w_n5036_0[1]),.doutc(w_n5036_0[2]),.din(n5036));
	jspl jspl_w_n5037_0(.douta(w_n5037_0[0]),.doutb(w_n5037_0[1]),.din(n5037));
	jspl3 jspl3_w_n5041_0(.douta(w_n5041_0[0]),.doutb(w_n5041_0[1]),.doutc(w_n5041_0[2]),.din(n5041));
	jspl3 jspl3_w_n5044_0(.douta(w_n5044_0[0]),.doutb(w_n5044_0[1]),.doutc(w_n5044_0[2]),.din(n5044));
	jspl jspl_w_n5045_0(.douta(w_n5045_0[0]),.doutb(w_n5045_0[1]),.din(n5045));
	jspl3 jspl3_w_n5049_0(.douta(w_n5049_0[0]),.doutb(w_n5049_0[1]),.doutc(w_n5049_0[2]),.din(n5049));
	jspl3 jspl3_w_n5051_0(.douta(w_n5051_0[0]),.doutb(w_n5051_0[1]),.doutc(w_n5051_0[2]),.din(n5051));
	jspl jspl_w_n5052_0(.douta(w_n5052_0[0]),.doutb(w_n5052_0[1]),.din(n5052));
	jspl3 jspl3_w_n5056_0(.douta(w_n5056_0[0]),.doutb(w_n5056_0[1]),.doutc(w_n5056_0[2]),.din(n5056));
	jspl3 jspl3_w_n5059_0(.douta(w_n5059_0[0]),.doutb(w_n5059_0[1]),.doutc(w_n5059_0[2]),.din(n5059));
	jspl jspl_w_n5060_0(.douta(w_n5060_0[0]),.doutb(w_n5060_0[1]),.din(n5060));
	jspl3 jspl3_w_n5064_0(.douta(w_n5064_0[0]),.doutb(w_n5064_0[1]),.doutc(w_n5064_0[2]),.din(n5064));
	jspl3 jspl3_w_n5066_0(.douta(w_n5066_0[0]),.doutb(w_n5066_0[1]),.doutc(w_n5066_0[2]),.din(n5066));
	jspl jspl_w_n5067_0(.douta(w_n5067_0[0]),.doutb(w_n5067_0[1]),.din(n5067));
	jspl jspl_w_n5071_0(.douta(w_n5071_0[0]),.doutb(w_n5071_0[1]),.din(n5071));
	jspl jspl_w_n5072_0(.douta(w_n5072_0[0]),.doutb(w_n5072_0[1]),.din(n5072));
	jspl3 jspl3_w_n5074_0(.douta(w_n5074_0[0]),.doutb(w_n5074_0[1]),.doutc(w_n5074_0[2]),.din(n5074));
	jspl jspl_w_n5075_0(.douta(w_n5075_0[0]),.doutb(w_n5075_0[1]),.din(n5075));
	jspl3 jspl3_w_n5079_0(.douta(w_n5079_0[0]),.doutb(w_n5079_0[1]),.doutc(w_n5079_0[2]),.din(n5079));
	jspl3 jspl3_w_n5081_0(.douta(w_n5081_0[0]),.doutb(w_n5081_0[1]),.doutc(w_n5081_0[2]),.din(n5081));
	jspl jspl_w_n5082_0(.douta(w_n5082_0[0]),.doutb(w_n5082_0[1]),.din(n5082));
	jspl3 jspl3_w_n5086_0(.douta(w_n5086_0[0]),.doutb(w_n5086_0[1]),.doutc(w_n5086_0[2]),.din(n5086));
	jspl3 jspl3_w_n5089_0(.douta(w_n5089_0[0]),.doutb(w_n5089_0[1]),.doutc(w_n5089_0[2]),.din(n5089));
	jspl jspl_w_n5090_0(.douta(w_n5090_0[0]),.doutb(w_n5090_0[1]),.din(n5090));
	jspl3 jspl3_w_n5094_0(.douta(w_n5094_0[0]),.doutb(w_n5094_0[1]),.doutc(w_n5094_0[2]),.din(n5094));
	jspl3 jspl3_w_n5096_0(.douta(w_n5096_0[0]),.doutb(w_n5096_0[1]),.doutc(w_n5096_0[2]),.din(n5096));
	jspl jspl_w_n5097_0(.douta(w_n5097_0[0]),.doutb(w_n5097_0[1]),.din(n5097));
	jspl jspl_w_n5101_0(.douta(w_n5101_0[0]),.doutb(w_n5101_0[1]),.din(n5101));
	jspl jspl_w_n5102_0(.douta(w_n5102_0[0]),.doutb(w_n5102_0[1]),.din(n5102));
	jspl3 jspl3_w_n5104_0(.douta(w_n5104_0[0]),.doutb(w_n5104_0[1]),.doutc(w_n5104_0[2]),.din(n5104));
	jspl3 jspl3_w_n5105_0(.douta(w_n5105_0[0]),.doutb(w_n5105_0[1]),.doutc(w_n5105_0[2]),.din(n5105));
	jspl jspl_w_n5107_0(.douta(w_n5107_0[0]),.doutb(w_n5107_0[1]),.din(n5107));
	jspl jspl_w_n5108_0(.douta(w_n5108_0[0]),.doutb(w_n5108_0[1]),.din(n5108));
	jspl jspl_w_n5115_0(.douta(w_n5115_0[0]),.doutb(w_n5115_0[1]),.din(n5115));
	jspl jspl_w_n5116_0(.douta(w_n5116_0[0]),.doutb(w_n5116_0[1]),.din(n5116));
	jspl jspl_w_n5118_0(.douta(w_n5118_0[0]),.doutb(w_n5118_0[1]),.din(n5118));
	jspl3 jspl3_w_n5121_0(.douta(w_n5121_0[0]),.doutb(w_n5121_0[1]),.doutc(w_n5121_0[2]),.din(n5121));
	jspl jspl_w_n5121_1(.douta(w_n5121_1[0]),.doutb(w_n5121_1[1]),.din(w_n5121_0[0]));
	jspl jspl_w_n5122_0(.douta(w_n5122_0[0]),.doutb(w_n5122_0[1]),.din(n5122));
	jspl3 jspl3_w_n5123_0(.douta(w_n5123_0[0]),.doutb(w_n5123_0[1]),.doutc(w_n5123_0[2]),.din(n5123));
	jspl jspl_w_n5124_0(.douta(w_n5124_0[0]),.doutb(w_n5124_0[1]),.din(n5124));
	jspl3 jspl3_w_n5126_0(.douta(w_n5126_0[0]),.doutb(w_n5126_0[1]),.doutc(w_n5126_0[2]),.din(n5126));
	jspl jspl_w_n5127_0(.douta(w_n5127_0[0]),.doutb(w_n5127_0[1]),.din(n5127));
	jspl3 jspl3_w_n5132_0(.douta(w_n5132_0[0]),.doutb(w_n5132_0[1]),.doutc(w_n5132_0[2]),.din(n5132));
	jspl jspl_w_n5132_1(.douta(w_n5132_1[0]),.doutb(w_n5132_1[1]),.din(w_n5132_0[0]));
	jspl jspl_w_n5165_0(.douta(w_n5165_0[0]),.doutb(w_n5165_0[1]),.din(n5165));
	jspl jspl_w_n5179_0(.douta(w_n5179_0[0]),.doutb(w_n5179_0[1]),.din(n5179));
	jspl jspl_w_n5253_0(.douta(w_n5253_0[0]),.doutb(w_n5253_0[1]),.din(n5253));
	jspl jspl_w_n5256_0(.douta(w_n5256_0[0]),.doutb(w_n5256_0[1]),.din(n5256));
	jspl jspl_w_n5257_0(.douta(w_n5257_0[0]),.doutb(w_n5257_0[1]),.din(n5257));
	jspl3 jspl3_w_n5259_0(.douta(w_n5259_0[0]),.doutb(w_n5259_0[1]),.doutc(w_n5259_0[2]),.din(n5259));
	jspl3 jspl3_w_n5259_1(.douta(w_n5259_1[0]),.doutb(w_n5259_1[1]),.doutc(w_n5259_1[2]),.din(w_n5259_0[0]));
	jspl3 jspl3_w_n5259_2(.douta(w_n5259_2[0]),.doutb(w_n5259_2[1]),.doutc(w_n5259_2[2]),.din(w_n5259_0[1]));
	jspl3 jspl3_w_n5259_3(.douta(w_n5259_3[0]),.doutb(w_n5259_3[1]),.doutc(w_n5259_3[2]),.din(w_n5259_0[2]));
	jspl3 jspl3_w_n5259_4(.douta(w_n5259_4[0]),.doutb(w_n5259_4[1]),.doutc(w_n5259_4[2]),.din(w_n5259_1[0]));
	jspl3 jspl3_w_n5259_5(.douta(w_n5259_5[0]),.doutb(w_n5259_5[1]),.doutc(w_n5259_5[2]),.din(w_n5259_1[1]));
	jspl3 jspl3_w_n5259_6(.douta(w_n5259_6[0]),.doutb(w_n5259_6[1]),.doutc(w_n5259_6[2]),.din(w_n5259_1[2]));
	jspl3 jspl3_w_n5259_7(.douta(w_n5259_7[0]),.doutb(w_n5259_7[1]),.doutc(w_n5259_7[2]),.din(w_n5259_2[0]));
	jspl3 jspl3_w_n5259_8(.douta(w_n5259_8[0]),.doutb(w_n5259_8[1]),.doutc(w_n5259_8[2]),.din(w_n5259_2[1]));
	jspl3 jspl3_w_n5259_9(.douta(w_n5259_9[0]),.doutb(w_n5259_9[1]),.doutc(w_n5259_9[2]),.din(w_n5259_2[2]));
	jspl3 jspl3_w_n5259_10(.douta(w_n5259_10[0]),.doutb(w_n5259_10[1]),.doutc(w_n5259_10[2]),.din(w_n5259_3[0]));
	jspl3 jspl3_w_n5259_11(.douta(w_n5259_11[0]),.doutb(w_n5259_11[1]),.doutc(w_n5259_11[2]),.din(w_n5259_3[1]));
	jspl3 jspl3_w_n5259_12(.douta(w_n5259_12[0]),.doutb(w_n5259_12[1]),.doutc(w_n5259_12[2]),.din(w_n5259_3[2]));
	jspl3 jspl3_w_n5259_13(.douta(w_n5259_13[0]),.doutb(w_n5259_13[1]),.doutc(w_n5259_13[2]),.din(w_n5259_4[0]));
	jspl3 jspl3_w_n5259_14(.douta(w_n5259_14[0]),.doutb(w_n5259_14[1]),.doutc(w_n5259_14[2]),.din(w_n5259_4[1]));
	jspl3 jspl3_w_n5259_15(.douta(w_n5259_15[0]),.doutb(w_n5259_15[1]),.doutc(w_n5259_15[2]),.din(w_n5259_4[2]));
	jspl3 jspl3_w_n5259_16(.douta(w_n5259_16[0]),.doutb(w_n5259_16[1]),.doutc(w_n5259_16[2]),.din(w_n5259_5[0]));
	jspl3 jspl3_w_n5259_17(.douta(w_n5259_17[0]),.doutb(w_n5259_17[1]),.doutc(w_n5259_17[2]),.din(w_n5259_5[1]));
	jspl3 jspl3_w_n5259_18(.douta(w_n5259_18[0]),.doutb(w_n5259_18[1]),.doutc(w_n5259_18[2]),.din(w_n5259_5[2]));
	jspl3 jspl3_w_n5259_19(.douta(w_n5259_19[0]),.doutb(w_n5259_19[1]),.doutc(w_n5259_19[2]),.din(w_n5259_6[0]));
	jspl3 jspl3_w_n5259_20(.douta(w_n5259_20[0]),.doutb(w_n5259_20[1]),.doutc(w_n5259_20[2]),.din(w_n5259_6[1]));
	jspl3 jspl3_w_n5259_21(.douta(w_n5259_21[0]),.doutb(w_n5259_21[1]),.doutc(w_n5259_21[2]),.din(w_n5259_6[2]));
	jspl3 jspl3_w_n5259_22(.douta(w_n5259_22[0]),.doutb(w_n5259_22[1]),.doutc(w_n5259_22[2]),.din(w_n5259_7[0]));
	jspl3 jspl3_w_n5259_23(.douta(w_n5259_23[0]),.doutb(w_n5259_23[1]),.doutc(w_n5259_23[2]),.din(w_n5259_7[1]));
	jspl3 jspl3_w_n5259_24(.douta(w_n5259_24[0]),.doutb(w_n5259_24[1]),.doutc(w_n5259_24[2]),.din(w_n5259_7[2]));
	jspl3 jspl3_w_n5259_25(.douta(w_n5259_25[0]),.doutb(w_n5259_25[1]),.doutc(w_n5259_25[2]),.din(w_n5259_8[0]));
	jspl3 jspl3_w_n5259_26(.douta(w_n5259_26[0]),.doutb(w_n5259_26[1]),.doutc(w_n5259_26[2]),.din(w_n5259_8[1]));
	jspl3 jspl3_w_n5259_27(.douta(w_n5259_27[0]),.doutb(w_n5259_27[1]),.doutc(w_n5259_27[2]),.din(w_n5259_8[2]));
	jspl3 jspl3_w_n5259_28(.douta(w_n5259_28[0]),.doutb(w_n5259_28[1]),.doutc(w_n5259_28[2]),.din(w_n5259_9[0]));
	jspl3 jspl3_w_n5259_29(.douta(w_n5259_29[0]),.doutb(w_n5259_29[1]),.doutc(w_n5259_29[2]),.din(w_n5259_9[1]));
	jspl3 jspl3_w_n5259_30(.douta(w_n5259_30[0]),.doutb(w_n5259_30[1]),.doutc(w_n5259_30[2]),.din(w_n5259_9[2]));
	jspl3 jspl3_w_n5259_31(.douta(w_n5259_31[0]),.doutb(w_n5259_31[1]),.doutc(w_n5259_31[2]),.din(w_n5259_10[0]));
	jspl3 jspl3_w_n5259_32(.douta(w_n5259_32[0]),.doutb(w_n5259_32[1]),.doutc(w_n5259_32[2]),.din(w_n5259_10[1]));
	jspl3 jspl3_w_n5259_33(.douta(w_n5259_33[0]),.doutb(w_n5259_33[1]),.doutc(w_n5259_33[2]),.din(w_n5259_10[2]));
	jspl3 jspl3_w_n5259_34(.douta(w_n5259_34[0]),.doutb(w_n5259_34[1]),.doutc(w_n5259_34[2]),.din(w_n5259_11[0]));
	jspl3 jspl3_w_n5259_35(.douta(w_n5259_35[0]),.doutb(w_n5259_35[1]),.doutc(w_n5259_35[2]),.din(w_n5259_11[1]));
	jspl3 jspl3_w_n5259_36(.douta(w_n5259_36[0]),.doutb(w_n5259_36[1]),.doutc(w_n5259_36[2]),.din(w_n5259_11[2]));
	jspl3 jspl3_w_n5259_37(.douta(w_n5259_37[0]),.doutb(w_n5259_37[1]),.doutc(w_n5259_37[2]),.din(w_n5259_12[0]));
	jspl3 jspl3_w_n5259_38(.douta(w_n5259_38[0]),.doutb(w_n5259_38[1]),.doutc(w_n5259_38[2]),.din(w_n5259_12[1]));
	jspl3 jspl3_w_n5259_39(.douta(w_n5259_39[0]),.doutb(w_n5259_39[1]),.doutc(w_n5259_39[2]),.din(w_n5259_12[2]));
	jspl3 jspl3_w_n5259_40(.douta(w_n5259_40[0]),.doutb(w_n5259_40[1]),.doutc(w_n5259_40[2]),.din(w_n5259_13[0]));
	jspl3 jspl3_w_n5259_41(.douta(w_n5259_41[0]),.doutb(w_n5259_41[1]),.doutc(w_n5259_41[2]),.din(w_n5259_13[1]));
	jspl3 jspl3_w_n5259_42(.douta(w_n5259_42[0]),.doutb(w_n5259_42[1]),.doutc(w_n5259_42[2]),.din(w_n5259_13[2]));
	jspl3 jspl3_w_n5259_43(.douta(w_n5259_43[0]),.doutb(w_n5259_43[1]),.doutc(w_n5259_43[2]),.din(w_n5259_14[0]));
	jspl3 jspl3_w_n5259_44(.douta(w_n5259_44[0]),.doutb(w_n5259_44[1]),.doutc(w_n5259_44[2]),.din(w_n5259_14[1]));
	jspl jspl_w_n5259_45(.douta(w_n5259_45[0]),.doutb(w_n5259_45[1]),.din(w_n5259_14[2]));
	jspl3 jspl3_w_n5263_0(.douta(w_n5263_0[0]),.doutb(w_n5263_0[1]),.doutc(w_n5263_0[2]),.din(n5263));
	jspl jspl_w_n5264_0(.douta(w_n5264_0[0]),.doutb(w_n5264_0[1]),.din(n5264));
	jspl jspl_w_n5266_0(.douta(w_n5266_0[0]),.doutb(w_n5266_0[1]),.din(n5266));
	jspl jspl_w_n5271_0(.douta(w_n5271_0[0]),.doutb(w_n5271_0[1]),.din(n5271));
	jspl jspl_w_n5272_0(.douta(w_n5272_0[0]),.doutb(w_n5272_0[1]),.din(n5272));
	jspl3 jspl3_w_n5274_0(.douta(w_n5274_0[0]),.doutb(w_n5274_0[1]),.doutc(w_n5274_0[2]),.din(n5274));
	jspl jspl_w_n5275_0(.douta(w_n5275_0[0]),.doutb(w_n5275_0[1]),.din(n5275));
	jspl jspl_w_n5279_0(.douta(w_n5279_0[0]),.doutb(w_n5279_0[1]),.din(n5279));
	jspl3 jspl3_w_n5281_0(.douta(w_n5281_0[0]),.doutb(w_n5281_0[1]),.doutc(w_n5281_0[2]),.din(n5281));
	jspl jspl_w_n5282_0(.douta(w_n5282_0[0]),.doutb(w_n5282_0[1]),.din(n5282));
	jspl jspl_w_n5286_0(.douta(w_n5286_0[0]),.doutb(w_n5286_0[1]),.din(n5286));
	jspl jspl_w_n5287_0(.douta(w_n5287_0[0]),.doutb(w_n5287_0[1]),.din(n5287));
	jspl3 jspl3_w_n5289_0(.douta(w_n5289_0[0]),.doutb(w_n5289_0[1]),.doutc(w_n5289_0[2]),.din(n5289));
	jspl jspl_w_n5290_0(.douta(w_n5290_0[0]),.doutb(w_n5290_0[1]),.din(n5290));
	jspl jspl_w_n5294_0(.douta(w_n5294_0[0]),.doutb(w_n5294_0[1]),.din(n5294));
	jspl3 jspl3_w_n5296_0(.douta(w_n5296_0[0]),.doutb(w_n5296_0[1]),.doutc(w_n5296_0[2]),.din(n5296));
	jspl jspl_w_n5297_0(.douta(w_n5297_0[0]),.doutb(w_n5297_0[1]),.din(n5297));
	jspl jspl_w_n5301_0(.douta(w_n5301_0[0]),.doutb(w_n5301_0[1]),.din(n5301));
	jspl3 jspl3_w_n5303_0(.douta(w_n5303_0[0]),.doutb(w_n5303_0[1]),.doutc(w_n5303_0[2]),.din(n5303));
	jspl jspl_w_n5304_0(.douta(w_n5304_0[0]),.doutb(w_n5304_0[1]),.din(n5304));
	jspl jspl_w_n5308_0(.douta(w_n5308_0[0]),.doutb(w_n5308_0[1]),.din(n5308));
	jspl3 jspl3_w_n5310_0(.douta(w_n5310_0[0]),.doutb(w_n5310_0[1]),.doutc(w_n5310_0[2]),.din(n5310));
	jspl jspl_w_n5311_0(.douta(w_n5311_0[0]),.doutb(w_n5311_0[1]),.din(n5311));
	jspl jspl_w_n5315_0(.douta(w_n5315_0[0]),.doutb(w_n5315_0[1]),.din(n5315));
	jspl jspl_w_n5316_0(.douta(w_n5316_0[0]),.doutb(w_n5316_0[1]),.din(n5316));
	jspl3 jspl3_w_n5318_0(.douta(w_n5318_0[0]),.doutb(w_n5318_0[1]),.doutc(w_n5318_0[2]),.din(n5318));
	jspl jspl_w_n5319_0(.douta(w_n5319_0[0]),.doutb(w_n5319_0[1]),.din(n5319));
	jspl jspl_w_n5323_0(.douta(w_n5323_0[0]),.doutb(w_n5323_0[1]),.din(n5323));
	jspl jspl_w_n5324_0(.douta(w_n5324_0[0]),.doutb(w_n5324_0[1]),.din(n5324));
	jspl3 jspl3_w_n5326_0(.douta(w_n5326_0[0]),.doutb(w_n5326_0[1]),.doutc(w_n5326_0[2]),.din(n5326));
	jspl jspl_w_n5327_0(.douta(w_n5327_0[0]),.doutb(w_n5327_0[1]),.din(n5327));
	jspl jspl_w_n5331_0(.douta(w_n5331_0[0]),.doutb(w_n5331_0[1]),.din(n5331));
	jspl jspl_w_n5332_0(.douta(w_n5332_0[0]),.doutb(w_n5332_0[1]),.din(n5332));
	jspl3 jspl3_w_n5334_0(.douta(w_n5334_0[0]),.doutb(w_n5334_0[1]),.doutc(w_n5334_0[2]),.din(n5334));
	jspl jspl_w_n5335_0(.douta(w_n5335_0[0]),.doutb(w_n5335_0[1]),.din(n5335));
	jspl jspl_w_n5339_0(.douta(w_n5339_0[0]),.doutb(w_n5339_0[1]),.din(n5339));
	jspl3 jspl3_w_n5341_0(.douta(w_n5341_0[0]),.doutb(w_n5341_0[1]),.doutc(w_n5341_0[2]),.din(n5341));
	jspl jspl_w_n5342_0(.douta(w_n5342_0[0]),.doutb(w_n5342_0[1]),.din(n5342));
	jspl jspl_w_n5346_0(.douta(w_n5346_0[0]),.doutb(w_n5346_0[1]),.din(n5346));
	jspl jspl_w_n5347_0(.douta(w_n5347_0[0]),.doutb(w_n5347_0[1]),.din(n5347));
	jspl3 jspl3_w_n5349_0(.douta(w_n5349_0[0]),.doutb(w_n5349_0[1]),.doutc(w_n5349_0[2]),.din(n5349));
	jspl jspl_w_n5350_0(.douta(w_n5350_0[0]),.doutb(w_n5350_0[1]),.din(n5350));
	jspl jspl_w_n5354_0(.douta(w_n5354_0[0]),.doutb(w_n5354_0[1]),.din(n5354));
	jspl3 jspl3_w_n5356_0(.douta(w_n5356_0[0]),.doutb(w_n5356_0[1]),.doutc(w_n5356_0[2]),.din(n5356));
	jspl jspl_w_n5357_0(.douta(w_n5357_0[0]),.doutb(w_n5357_0[1]),.din(n5357));
	jspl jspl_w_n5361_0(.douta(w_n5361_0[0]),.doutb(w_n5361_0[1]),.din(n5361));
	jspl jspl_w_n5362_0(.douta(w_n5362_0[0]),.doutb(w_n5362_0[1]),.din(n5362));
	jspl3 jspl3_w_n5364_0(.douta(w_n5364_0[0]),.doutb(w_n5364_0[1]),.doutc(w_n5364_0[2]),.din(n5364));
	jspl jspl_w_n5365_0(.douta(w_n5365_0[0]),.doutb(w_n5365_0[1]),.din(n5365));
	jspl jspl_w_n5369_0(.douta(w_n5369_0[0]),.doutb(w_n5369_0[1]),.din(n5369));
	jspl3 jspl3_w_n5371_0(.douta(w_n5371_0[0]),.doutb(w_n5371_0[1]),.doutc(w_n5371_0[2]),.din(n5371));
	jspl jspl_w_n5372_0(.douta(w_n5372_0[0]),.doutb(w_n5372_0[1]),.din(n5372));
	jspl jspl_w_n5376_0(.douta(w_n5376_0[0]),.doutb(w_n5376_0[1]),.din(n5376));
	jspl3 jspl3_w_n5378_0(.douta(w_n5378_0[0]),.doutb(w_n5378_0[1]),.doutc(w_n5378_0[2]),.din(n5378));
	jspl jspl_w_n5379_0(.douta(w_n5379_0[0]),.doutb(w_n5379_0[1]),.din(n5379));
	jspl jspl_w_n5383_0(.douta(w_n5383_0[0]),.doutb(w_n5383_0[1]),.din(n5383));
	jspl jspl_w_n5384_0(.douta(w_n5384_0[0]),.doutb(w_n5384_0[1]),.din(n5384));
	jspl3 jspl3_w_n5386_0(.douta(w_n5386_0[0]),.doutb(w_n5386_0[1]),.doutc(w_n5386_0[2]),.din(n5386));
	jspl jspl_w_n5387_0(.douta(w_n5387_0[0]),.doutb(w_n5387_0[1]),.din(n5387));
	jspl jspl_w_n5391_0(.douta(w_n5391_0[0]),.doutb(w_n5391_0[1]),.din(n5391));
	jspl jspl_w_n5392_0(.douta(w_n5392_0[0]),.doutb(w_n5392_0[1]),.din(n5392));
	jspl3 jspl3_w_n5394_0(.douta(w_n5394_0[0]),.doutb(w_n5394_0[1]),.doutc(w_n5394_0[2]),.din(n5394));
	jspl jspl_w_n5395_0(.douta(w_n5395_0[0]),.doutb(w_n5395_0[1]),.din(n5395));
	jspl jspl_w_n5399_0(.douta(w_n5399_0[0]),.doutb(w_n5399_0[1]),.din(n5399));
	jspl3 jspl3_w_n5401_0(.douta(w_n5401_0[0]),.doutb(w_n5401_0[1]),.doutc(w_n5401_0[2]),.din(n5401));
	jspl jspl_w_n5402_0(.douta(w_n5402_0[0]),.doutb(w_n5402_0[1]),.din(n5402));
	jspl jspl_w_n5406_0(.douta(w_n5406_0[0]),.doutb(w_n5406_0[1]),.din(n5406));
	jspl jspl_w_n5407_0(.douta(w_n5407_0[0]),.doutb(w_n5407_0[1]),.din(n5407));
	jspl3 jspl3_w_n5409_0(.douta(w_n5409_0[0]),.doutb(w_n5409_0[1]),.doutc(w_n5409_0[2]),.din(n5409));
	jspl jspl_w_n5410_0(.douta(w_n5410_0[0]),.doutb(w_n5410_0[1]),.din(n5410));
	jspl jspl_w_n5414_0(.douta(w_n5414_0[0]),.doutb(w_n5414_0[1]),.din(n5414));
	jspl3 jspl3_w_n5416_0(.douta(w_n5416_0[0]),.doutb(w_n5416_0[1]),.doutc(w_n5416_0[2]),.din(n5416));
	jspl jspl_w_n5417_0(.douta(w_n5417_0[0]),.doutb(w_n5417_0[1]),.din(n5417));
	jspl jspl_w_n5421_0(.douta(w_n5421_0[0]),.doutb(w_n5421_0[1]),.din(n5421));
	jspl jspl_w_n5422_0(.douta(w_n5422_0[0]),.doutb(w_n5422_0[1]),.din(n5422));
	jspl3 jspl3_w_n5424_0(.douta(w_n5424_0[0]),.doutb(w_n5424_0[1]),.doutc(w_n5424_0[2]),.din(n5424));
	jspl jspl_w_n5425_0(.douta(w_n5425_0[0]),.doutb(w_n5425_0[1]),.din(n5425));
	jspl jspl_w_n5429_0(.douta(w_n5429_0[0]),.doutb(w_n5429_0[1]),.din(n5429));
	jspl jspl_w_n5430_0(.douta(w_n5430_0[0]),.doutb(w_n5430_0[1]),.din(n5430));
	jspl3 jspl3_w_n5432_0(.douta(w_n5432_0[0]),.doutb(w_n5432_0[1]),.doutc(w_n5432_0[2]),.din(n5432));
	jspl jspl_w_n5433_0(.douta(w_n5433_0[0]),.doutb(w_n5433_0[1]),.din(n5433));
	jspl jspl_w_n5437_0(.douta(w_n5437_0[0]),.doutb(w_n5437_0[1]),.din(n5437));
	jspl jspl_w_n5438_0(.douta(w_n5438_0[0]),.doutb(w_n5438_0[1]),.din(n5438));
	jspl3 jspl3_w_n5440_0(.douta(w_n5440_0[0]),.doutb(w_n5440_0[1]),.doutc(w_n5440_0[2]),.din(n5440));
	jspl jspl_w_n5441_0(.douta(w_n5441_0[0]),.doutb(w_n5441_0[1]),.din(n5441));
	jspl jspl_w_n5445_0(.douta(w_n5445_0[0]),.doutb(w_n5445_0[1]),.din(n5445));
	jspl3 jspl3_w_n5447_0(.douta(w_n5447_0[0]),.doutb(w_n5447_0[1]),.doutc(w_n5447_0[2]),.din(n5447));
	jspl jspl_w_n5448_0(.douta(w_n5448_0[0]),.doutb(w_n5448_0[1]),.din(n5448));
	jspl3 jspl3_w_n5452_0(.douta(w_n5452_0[0]),.doutb(w_n5452_0[1]),.doutc(w_n5452_0[2]),.din(n5452));
	jspl3 jspl3_w_n5455_0(.douta(w_n5455_0[0]),.doutb(w_n5455_0[1]),.doutc(w_n5455_0[2]),.din(n5455));
	jspl jspl_w_n5458_0(.douta(w_n5458_0[0]),.doutb(w_n5458_0[1]),.din(n5458));
	jspl3 jspl3_w_n5459_0(.douta(w_n5459_0[0]),.doutb(w_n5459_0[1]),.doutc(w_n5459_0[2]),.din(n5459));
	jspl jspl_w_n5460_0(.douta(w_n5460_0[0]),.doutb(w_n5460_0[1]),.din(n5460));
	jspl jspl_w_n5461_0(.douta(w_n5461_0[0]),.doutb(w_n5461_0[1]),.din(n5461));
	jspl jspl_w_n5465_0(.douta(w_n5465_0[0]),.doutb(w_n5465_0[1]),.din(n5465));
	jspl jspl_w_n5466_0(.douta(w_n5466_0[0]),.doutb(w_n5466_0[1]),.din(n5466));
	jspl jspl_w_n5467_0(.douta(w_n5467_0[0]),.doutb(w_n5467_0[1]),.din(n5467));
	jspl jspl_w_n5500_0(.douta(w_n5500_0[0]),.doutb(w_n5500_0[1]),.din(n5500));
	jspl jspl_w_n5507_0(.douta(w_n5507_0[0]),.doutb(w_n5507_0[1]),.din(n5507));
	jspl jspl_w_n5514_0(.douta(w_n5514_0[0]),.doutb(w_n5514_0[1]),.din(n5514));
	jspl jspl_w_n5518_0(.douta(w_n5518_0[0]),.doutb(w_n5518_0[1]),.din(n5518));
	jspl jspl_w_n5522_0(.douta(w_n5522_0[0]),.doutb(w_n5522_0[1]),.din(n5522));
	jspl jspl_w_n5535_0(.douta(w_n5535_0[0]),.doutb(w_n5535_0[1]),.din(n5535));
	jspl jspl_w_n5542_0(.douta(w_n5542_0[0]),.doutb(w_n5542_0[1]),.din(n5542));
	jspl jspl_w_n5549_0(.douta(w_n5549_0[0]),.doutb(w_n5549_0[1]),.din(n5549));
	jspl jspl_w_n5553_0(.douta(w_n5553_0[0]),.doutb(w_n5553_0[1]),.din(n5553));
	jspl jspl_w_n5563_0(.douta(w_n5563_0[0]),.doutb(w_n5563_0[1]),.din(n5563));
	jspl jspl_w_n5570_0(.douta(w_n5570_0[0]),.doutb(w_n5570_0[1]),.din(n5570));
	jspl jspl_w_n5583_0(.douta(w_n5583_0[0]),.doutb(w_n5583_0[1]),.din(n5583));
	jspl jspl_w_n5588_0(.douta(w_n5588_0[0]),.doutb(w_n5588_0[1]),.din(n5588));
	jspl jspl_w_n5592_0(.douta(w_n5592_0[0]),.doutb(w_n5592_0[1]),.din(n5592));
	jspl jspl_w_n5593_0(.douta(w_n5593_0[0]),.doutb(w_n5593_0[1]),.din(n5593));
	jspl jspl_w_n5605_0(.douta(w_n5605_0[0]),.doutb(w_n5605_0[1]),.din(n5605));
	jspl3 jspl3_w_n5606_0(.douta(w_n5606_0[0]),.doutb(w_n5606_0[1]),.doutc(w_n5606_0[2]),.din(n5606));
	jspl3 jspl3_w_n5606_1(.douta(w_n5606_1[0]),.doutb(w_n5606_1[1]),.doutc(w_n5606_1[2]),.din(w_n5606_0[0]));
	jspl3 jspl3_w_n5606_2(.douta(w_n5606_2[0]),.doutb(w_n5606_2[1]),.doutc(w_n5606_2[2]),.din(w_n5606_0[1]));
	jspl3 jspl3_w_n5606_3(.douta(w_n5606_3[0]),.doutb(w_n5606_3[1]),.doutc(w_n5606_3[2]),.din(w_n5606_0[2]));
	jspl3 jspl3_w_n5606_4(.douta(w_n5606_4[0]),.doutb(w_n5606_4[1]),.doutc(w_n5606_4[2]),.din(w_n5606_1[0]));
	jspl3 jspl3_w_n5606_5(.douta(w_n5606_5[0]),.doutb(w_n5606_5[1]),.doutc(w_n5606_5[2]),.din(w_n5606_1[1]));
	jspl3 jspl3_w_n5606_6(.douta(w_n5606_6[0]),.doutb(w_n5606_6[1]),.doutc(w_n5606_6[2]),.din(w_n5606_1[2]));
	jspl3 jspl3_w_n5606_7(.douta(w_n5606_7[0]),.doutb(w_n5606_7[1]),.doutc(w_n5606_7[2]),.din(w_n5606_2[0]));
	jspl3 jspl3_w_n5606_8(.douta(w_n5606_8[0]),.doutb(w_n5606_8[1]),.doutc(w_n5606_8[2]),.din(w_n5606_2[1]));
	jspl3 jspl3_w_n5606_9(.douta(w_n5606_9[0]),.doutb(w_n5606_9[1]),.doutc(w_n5606_9[2]),.din(w_n5606_2[2]));
	jspl3 jspl3_w_n5606_10(.douta(w_n5606_10[0]),.doutb(w_n5606_10[1]),.doutc(w_n5606_10[2]),.din(w_n5606_3[0]));
	jspl3 jspl3_w_n5606_11(.douta(w_n5606_11[0]),.doutb(w_n5606_11[1]),.doutc(w_n5606_11[2]),.din(w_n5606_3[1]));
	jspl3 jspl3_w_n5606_12(.douta(w_n5606_12[0]),.doutb(w_n5606_12[1]),.doutc(w_n5606_12[2]),.din(w_n5606_3[2]));
	jspl3 jspl3_w_n5606_13(.douta(w_n5606_13[0]),.doutb(w_n5606_13[1]),.doutc(w_n5606_13[2]),.din(w_n5606_4[0]));
	jspl3 jspl3_w_n5606_14(.douta(w_n5606_14[0]),.doutb(w_n5606_14[1]),.doutc(w_n5606_14[2]),.din(w_n5606_4[1]));
	jspl3 jspl3_w_n5606_15(.douta(w_n5606_15[0]),.doutb(w_n5606_15[1]),.doutc(w_n5606_15[2]),.din(w_n5606_4[2]));
	jspl3 jspl3_w_n5606_16(.douta(w_n5606_16[0]),.doutb(w_n5606_16[1]),.doutc(w_n5606_16[2]),.din(w_n5606_5[0]));
	jspl3 jspl3_w_n5606_17(.douta(w_n5606_17[0]),.doutb(w_n5606_17[1]),.doutc(w_n5606_17[2]),.din(w_n5606_5[1]));
	jspl3 jspl3_w_n5606_18(.douta(w_n5606_18[0]),.doutb(w_n5606_18[1]),.doutc(w_n5606_18[2]),.din(w_n5606_5[2]));
	jspl3 jspl3_w_n5606_19(.douta(w_n5606_19[0]),.doutb(w_n5606_19[1]),.doutc(w_n5606_19[2]),.din(w_n5606_6[0]));
	jspl3 jspl3_w_n5606_20(.douta(w_n5606_20[0]),.doutb(w_n5606_20[1]),.doutc(w_n5606_20[2]),.din(w_n5606_6[1]));
	jspl3 jspl3_w_n5606_21(.douta(w_n5606_21[0]),.doutb(w_n5606_21[1]),.doutc(w_n5606_21[2]),.din(w_n5606_6[2]));
	jspl3 jspl3_w_n5606_22(.douta(w_n5606_22[0]),.doutb(w_n5606_22[1]),.doutc(w_n5606_22[2]),.din(w_n5606_7[0]));
	jspl3 jspl3_w_n5606_23(.douta(w_n5606_23[0]),.doutb(w_n5606_23[1]),.doutc(w_n5606_23[2]),.din(w_n5606_7[1]));
	jspl3 jspl3_w_n5606_24(.douta(w_n5606_24[0]),.doutb(w_n5606_24[1]),.doutc(w_n5606_24[2]),.din(w_n5606_7[2]));
	jspl3 jspl3_w_n5606_25(.douta(w_n5606_25[0]),.doutb(w_n5606_25[1]),.doutc(w_n5606_25[2]),.din(w_n5606_8[0]));
	jspl3 jspl3_w_n5606_26(.douta(w_n5606_26[0]),.doutb(w_n5606_26[1]),.doutc(w_n5606_26[2]),.din(w_n5606_8[1]));
	jspl3 jspl3_w_n5606_27(.douta(w_n5606_27[0]),.doutb(w_n5606_27[1]),.doutc(w_n5606_27[2]),.din(w_n5606_8[2]));
	jspl3 jspl3_w_n5606_28(.douta(w_n5606_28[0]),.doutb(w_n5606_28[1]),.doutc(w_n5606_28[2]),.din(w_n5606_9[0]));
	jspl3 jspl3_w_n5606_29(.douta(w_n5606_29[0]),.doutb(w_n5606_29[1]),.doutc(w_n5606_29[2]),.din(w_n5606_9[1]));
	jspl3 jspl3_w_n5606_30(.douta(w_n5606_30[0]),.doutb(w_n5606_30[1]),.doutc(w_n5606_30[2]),.din(w_n5606_9[2]));
	jspl3 jspl3_w_n5606_31(.douta(w_n5606_31[0]),.doutb(w_n5606_31[1]),.doutc(w_n5606_31[2]),.din(w_n5606_10[0]));
	jspl3 jspl3_w_n5606_32(.douta(w_n5606_32[0]),.doutb(w_n5606_32[1]),.doutc(w_n5606_32[2]),.din(w_n5606_10[1]));
	jspl3 jspl3_w_n5606_33(.douta(w_n5606_33[0]),.doutb(w_n5606_33[1]),.doutc(w_n5606_33[2]),.din(w_n5606_10[2]));
	jspl3 jspl3_w_n5606_34(.douta(w_n5606_34[0]),.doutb(w_n5606_34[1]),.doutc(w_n5606_34[2]),.din(w_n5606_11[0]));
	jspl3 jspl3_w_n5606_35(.douta(w_n5606_35[0]),.doutb(w_n5606_35[1]),.doutc(w_n5606_35[2]),.din(w_n5606_11[1]));
	jspl3 jspl3_w_n5606_36(.douta(w_n5606_36[0]),.doutb(w_n5606_36[1]),.doutc(w_n5606_36[2]),.din(w_n5606_11[2]));
	jspl3 jspl3_w_n5606_37(.douta(w_n5606_37[0]),.doutb(w_n5606_37[1]),.doutc(w_n5606_37[2]),.din(w_n5606_12[0]));
	jspl3 jspl3_w_n5606_38(.douta(w_n5606_38[0]),.doutb(w_n5606_38[1]),.doutc(w_n5606_38[2]),.din(w_n5606_12[1]));
	jspl3 jspl3_w_n5606_39(.douta(w_n5606_39[0]),.doutb(w_n5606_39[1]),.doutc(w_n5606_39[2]),.din(w_n5606_12[2]));
	jspl3 jspl3_w_n5606_40(.douta(w_n5606_40[0]),.doutb(w_n5606_40[1]),.doutc(w_n5606_40[2]),.din(w_n5606_13[0]));
	jspl3 jspl3_w_n5606_41(.douta(w_n5606_41[0]),.doutb(w_n5606_41[1]),.doutc(w_n5606_41[2]),.din(w_n5606_13[1]));
	jspl3 jspl3_w_n5606_42(.douta(w_n5606_42[0]),.doutb(w_n5606_42[1]),.doutc(w_n5606_42[2]),.din(w_n5606_13[2]));
	jspl3 jspl3_w_n5606_43(.douta(w_n5606_43[0]),.doutb(w_n5606_43[1]),.doutc(w_n5606_43[2]),.din(w_n5606_14[0]));
	jspl3 jspl3_w_n5606_44(.douta(w_n5606_44[0]),.doutb(w_n5606_44[1]),.doutc(w_n5606_44[2]),.din(w_n5606_14[1]));
	jspl3 jspl3_w_n5606_45(.douta(w_n5606_45[0]),.doutb(w_n5606_45[1]),.doutc(w_n5606_45[2]),.din(w_n5606_14[2]));
	jspl3 jspl3_w_n5606_46(.douta(w_n5606_46[0]),.doutb(w_n5606_46[1]),.doutc(w_n5606_46[2]),.din(w_n5606_15[0]));
	jspl3 jspl3_w_n5606_47(.douta(w_n5606_47[0]),.doutb(w_n5606_47[1]),.doutc(w_n5606_47[2]),.din(w_n5606_15[1]));
	jspl3 jspl3_w_n5606_48(.douta(w_n5606_48[0]),.doutb(w_n5606_48[1]),.doutc(w_n5606_48[2]),.din(w_n5606_15[2]));
	jspl3 jspl3_w_n5606_49(.douta(w_n5606_49[0]),.doutb(w_n5606_49[1]),.doutc(w_n5606_49[2]),.din(w_n5606_16[0]));
	jspl3 jspl3_w_n5606_50(.douta(w_n5606_50[0]),.doutb(w_n5606_50[1]),.doutc(w_n5606_50[2]),.din(w_n5606_16[1]));
	jspl3 jspl3_w_n5606_51(.douta(w_n5606_51[0]),.doutb(w_n5606_51[1]),.doutc(w_n5606_51[2]),.din(w_n5606_16[2]));
	jspl3 jspl3_w_n5606_52(.douta(w_n5606_52[0]),.doutb(w_n5606_52[1]),.doutc(w_n5606_52[2]),.din(w_n5606_17[0]));
	jspl3 jspl3_w_n5606_53(.douta(w_n5606_53[0]),.doutb(w_n5606_53[1]),.doutc(w_n5606_53[2]),.din(w_n5606_17[1]));
	jspl3 jspl3_w_n5606_54(.douta(w_n5606_54[0]),.doutb(w_n5606_54[1]),.doutc(w_n5606_54[2]),.din(w_n5606_17[2]));
	jspl3 jspl3_w_n5606_55(.douta(w_n5606_55[0]),.doutb(w_n5606_55[1]),.doutc(w_n5606_55[2]),.din(w_n5606_18[0]));
	jspl jspl_w_n5609_0(.douta(w_n5609_0[0]),.doutb(w_n5609_0[1]),.din(n5609));
	jspl3 jspl3_w_n5610_0(.douta(w_n5610_0[0]),.doutb(w_n5610_0[1]),.doutc(w_n5610_0[2]),.din(n5610));
	jspl3 jspl3_w_n5612_0(.douta(w_n5612_0[0]),.doutb(w_n5612_0[1]),.doutc(w_n5612_0[2]),.din(n5612));
	jspl3 jspl3_w_n5612_1(.douta(w_n5612_1[0]),.doutb(w_n5612_1[1]),.doutc(w_n5612_1[2]),.din(w_n5612_0[0]));
	jspl jspl_w_n5613_0(.douta(w_n5613_0[0]),.doutb(w_n5613_0[1]),.din(n5613));
	jspl3 jspl3_w_n5614_0(.douta(w_n5614_0[0]),.doutb(w_n5614_0[1]),.doutc(w_n5614_0[2]),.din(n5614));
	jspl jspl_w_n5615_0(.douta(w_n5615_0[0]),.doutb(w_n5615_0[1]),.din(n5615));
	jspl3 jspl3_w_n5617_0(.douta(w_n5617_0[0]),.doutb(w_n5617_0[1]),.doutc(w_n5617_0[2]),.din(n5617));
	jspl jspl_w_n5618_0(.douta(w_n5618_0[0]),.doutb(w_n5618_0[1]),.din(n5618));
	jspl3 jspl3_w_n5625_0(.douta(w_n5625_0[0]),.doutb(w_n5625_0[1]),.doutc(w_n5625_0[2]),.din(n5625));
	jspl jspl_w_n5626_0(.douta(w_n5626_0[0]),.doutb(w_n5626_0[1]),.din(n5626));
	jspl jspl_w_n5629_0(.douta(w_n5629_0[0]),.doutb(w_n5629_0[1]),.din(n5629));
	jspl3 jspl3_w_n5634_0(.douta(w_n5634_0[0]),.doutb(w_n5634_0[1]),.doutc(w_n5634_0[2]),.din(n5634));
	jspl3 jspl3_w_n5636_0(.douta(w_n5636_0[0]),.doutb(w_n5636_0[1]),.doutc(w_n5636_0[2]),.din(n5636));
	jspl jspl_w_n5637_0(.douta(w_n5637_0[0]),.doutb(w_n5637_0[1]),.din(n5637));
	jspl3 jspl3_w_n5641_0(.douta(w_n5641_0[0]),.doutb(w_n5641_0[1]),.doutc(w_n5641_0[2]),.din(n5641));
	jspl3 jspl3_w_n5644_0(.douta(w_n5644_0[0]),.doutb(w_n5644_0[1]),.doutc(w_n5644_0[2]),.din(n5644));
	jspl jspl_w_n5645_0(.douta(w_n5645_0[0]),.doutb(w_n5645_0[1]),.din(n5645));
	jspl3 jspl3_w_n5649_0(.douta(w_n5649_0[0]),.doutb(w_n5649_0[1]),.doutc(w_n5649_0[2]),.din(n5649));
	jspl3 jspl3_w_n5651_0(.douta(w_n5651_0[0]),.doutb(w_n5651_0[1]),.doutc(w_n5651_0[2]),.din(n5651));
	jspl jspl_w_n5652_0(.douta(w_n5652_0[0]),.doutb(w_n5652_0[1]),.din(n5652));
	jspl3 jspl3_w_n5656_0(.douta(w_n5656_0[0]),.doutb(w_n5656_0[1]),.doutc(w_n5656_0[2]),.din(n5656));
	jspl3 jspl3_w_n5659_0(.douta(w_n5659_0[0]),.doutb(w_n5659_0[1]),.doutc(w_n5659_0[2]),.din(n5659));
	jspl jspl_w_n5660_0(.douta(w_n5660_0[0]),.doutb(w_n5660_0[1]),.din(n5660));
	jspl3 jspl3_w_n5664_0(.douta(w_n5664_0[0]),.doutb(w_n5664_0[1]),.doutc(w_n5664_0[2]),.din(n5664));
	jspl3 jspl3_w_n5666_0(.douta(w_n5666_0[0]),.doutb(w_n5666_0[1]),.doutc(w_n5666_0[2]),.din(n5666));
	jspl jspl_w_n5667_0(.douta(w_n5667_0[0]),.doutb(w_n5667_0[1]),.din(n5667));
	jspl3 jspl3_w_n5671_0(.douta(w_n5671_0[0]),.doutb(w_n5671_0[1]),.doutc(w_n5671_0[2]),.din(n5671));
	jspl3 jspl3_w_n5674_0(.douta(w_n5674_0[0]),.doutb(w_n5674_0[1]),.doutc(w_n5674_0[2]),.din(n5674));
	jspl jspl_w_n5675_0(.douta(w_n5675_0[0]),.doutb(w_n5675_0[1]),.din(n5675));
	jspl3 jspl3_w_n5679_0(.douta(w_n5679_0[0]),.doutb(w_n5679_0[1]),.doutc(w_n5679_0[2]),.din(n5679));
	jspl3 jspl3_w_n5682_0(.douta(w_n5682_0[0]),.doutb(w_n5682_0[1]),.doutc(w_n5682_0[2]),.din(n5682));
	jspl jspl_w_n5683_0(.douta(w_n5683_0[0]),.doutb(w_n5683_0[1]),.din(n5683));
	jspl3 jspl3_w_n5687_0(.douta(w_n5687_0[0]),.doutb(w_n5687_0[1]),.doutc(w_n5687_0[2]),.din(n5687));
	jspl3 jspl3_w_n5690_0(.douta(w_n5690_0[0]),.doutb(w_n5690_0[1]),.doutc(w_n5690_0[2]),.din(n5690));
	jspl jspl_w_n5691_0(.douta(w_n5691_0[0]),.doutb(w_n5691_0[1]),.din(n5691));
	jspl3 jspl3_w_n5695_0(.douta(w_n5695_0[0]),.doutb(w_n5695_0[1]),.doutc(w_n5695_0[2]),.din(n5695));
	jspl3 jspl3_w_n5697_0(.douta(w_n5697_0[0]),.doutb(w_n5697_0[1]),.doutc(w_n5697_0[2]),.din(n5697));
	jspl jspl_w_n5698_0(.douta(w_n5698_0[0]),.doutb(w_n5698_0[1]),.din(n5698));
	jspl3 jspl3_w_n5702_0(.douta(w_n5702_0[0]),.doutb(w_n5702_0[1]),.doutc(w_n5702_0[2]),.din(n5702));
	jspl3 jspl3_w_n5704_0(.douta(w_n5704_0[0]),.doutb(w_n5704_0[1]),.doutc(w_n5704_0[2]),.din(n5704));
	jspl jspl_w_n5705_0(.douta(w_n5705_0[0]),.doutb(w_n5705_0[1]),.din(n5705));
	jspl3 jspl3_w_n5709_0(.douta(w_n5709_0[0]),.doutb(w_n5709_0[1]),.doutc(w_n5709_0[2]),.din(n5709));
	jspl3 jspl3_w_n5711_0(.douta(w_n5711_0[0]),.doutb(w_n5711_0[1]),.doutc(w_n5711_0[2]),.din(n5711));
	jspl jspl_w_n5712_0(.douta(w_n5712_0[0]),.doutb(w_n5712_0[1]),.din(n5712));
	jspl3 jspl3_w_n5716_0(.douta(w_n5716_0[0]),.doutb(w_n5716_0[1]),.doutc(w_n5716_0[2]),.din(n5716));
	jspl3 jspl3_w_n5719_0(.douta(w_n5719_0[0]),.doutb(w_n5719_0[1]),.doutc(w_n5719_0[2]),.din(n5719));
	jspl jspl_w_n5720_0(.douta(w_n5720_0[0]),.doutb(w_n5720_0[1]),.din(n5720));
	jspl3 jspl3_w_n5724_0(.douta(w_n5724_0[0]),.doutb(w_n5724_0[1]),.doutc(w_n5724_0[2]),.din(n5724));
	jspl3 jspl3_w_n5726_0(.douta(w_n5726_0[0]),.doutb(w_n5726_0[1]),.doutc(w_n5726_0[2]),.din(n5726));
	jspl jspl_w_n5727_0(.douta(w_n5727_0[0]),.doutb(w_n5727_0[1]),.din(n5727));
	jspl3 jspl3_w_n5731_0(.douta(w_n5731_0[0]),.doutb(w_n5731_0[1]),.doutc(w_n5731_0[2]),.din(n5731));
	jspl3 jspl3_w_n5734_0(.douta(w_n5734_0[0]),.doutb(w_n5734_0[1]),.doutc(w_n5734_0[2]),.din(n5734));
	jspl jspl_w_n5735_0(.douta(w_n5735_0[0]),.doutb(w_n5735_0[1]),.din(n5735));
	jspl3 jspl3_w_n5739_0(.douta(w_n5739_0[0]),.doutb(w_n5739_0[1]),.doutc(w_n5739_0[2]),.din(n5739));
	jspl3 jspl3_w_n5741_0(.douta(w_n5741_0[0]),.doutb(w_n5741_0[1]),.doutc(w_n5741_0[2]),.din(n5741));
	jspl jspl_w_n5742_0(.douta(w_n5742_0[0]),.doutb(w_n5742_0[1]),.din(n5742));
	jspl3 jspl3_w_n5746_0(.douta(w_n5746_0[0]),.doutb(w_n5746_0[1]),.doutc(w_n5746_0[2]),.din(n5746));
	jspl3 jspl3_w_n5749_0(.douta(w_n5749_0[0]),.doutb(w_n5749_0[1]),.doutc(w_n5749_0[2]),.din(n5749));
	jspl jspl_w_n5750_0(.douta(w_n5750_0[0]),.doutb(w_n5750_0[1]),.din(n5750));
	jspl3 jspl3_w_n5754_0(.douta(w_n5754_0[0]),.doutb(w_n5754_0[1]),.doutc(w_n5754_0[2]),.din(n5754));
	jspl3 jspl3_w_n5757_0(.douta(w_n5757_0[0]),.doutb(w_n5757_0[1]),.doutc(w_n5757_0[2]),.din(n5757));
	jspl jspl_w_n5758_0(.douta(w_n5758_0[0]),.doutb(w_n5758_0[1]),.din(n5758));
	jspl3 jspl3_w_n5762_0(.douta(w_n5762_0[0]),.doutb(w_n5762_0[1]),.doutc(w_n5762_0[2]),.din(n5762));
	jspl3 jspl3_w_n5764_0(.douta(w_n5764_0[0]),.doutb(w_n5764_0[1]),.doutc(w_n5764_0[2]),.din(n5764));
	jspl jspl_w_n5765_0(.douta(w_n5765_0[0]),.doutb(w_n5765_0[1]),.din(n5765));
	jspl3 jspl3_w_n5769_0(.douta(w_n5769_0[0]),.doutb(w_n5769_0[1]),.doutc(w_n5769_0[2]),.din(n5769));
	jspl3 jspl3_w_n5771_0(.douta(w_n5771_0[0]),.doutb(w_n5771_0[1]),.doutc(w_n5771_0[2]),.din(n5771));
	jspl jspl_w_n5772_0(.douta(w_n5772_0[0]),.doutb(w_n5772_0[1]),.din(n5772));
	jspl3 jspl3_w_n5776_0(.douta(w_n5776_0[0]),.doutb(w_n5776_0[1]),.doutc(w_n5776_0[2]),.din(n5776));
	jspl3 jspl3_w_n5779_0(.douta(w_n5779_0[0]),.doutb(w_n5779_0[1]),.doutc(w_n5779_0[2]),.din(n5779));
	jspl jspl_w_n5780_0(.douta(w_n5780_0[0]),.doutb(w_n5780_0[1]),.din(n5780));
	jspl3 jspl3_w_n5784_0(.douta(w_n5784_0[0]),.doutb(w_n5784_0[1]),.doutc(w_n5784_0[2]),.din(n5784));
	jspl3 jspl3_w_n5786_0(.douta(w_n5786_0[0]),.doutb(w_n5786_0[1]),.doutc(w_n5786_0[2]),.din(n5786));
	jspl jspl_w_n5787_0(.douta(w_n5787_0[0]),.doutb(w_n5787_0[1]),.din(n5787));
	jspl3 jspl3_w_n5791_0(.douta(w_n5791_0[0]),.doutb(w_n5791_0[1]),.doutc(w_n5791_0[2]),.din(n5791));
	jspl3 jspl3_w_n5794_0(.douta(w_n5794_0[0]),.doutb(w_n5794_0[1]),.doutc(w_n5794_0[2]),.din(n5794));
	jspl jspl_w_n5795_0(.douta(w_n5795_0[0]),.doutb(w_n5795_0[1]),.din(n5795));
	jspl3 jspl3_w_n5799_0(.douta(w_n5799_0[0]),.doutb(w_n5799_0[1]),.doutc(w_n5799_0[2]),.din(n5799));
	jspl3 jspl3_w_n5801_0(.douta(w_n5801_0[0]),.doutb(w_n5801_0[1]),.doutc(w_n5801_0[2]),.din(n5801));
	jspl jspl_w_n5802_0(.douta(w_n5802_0[0]),.doutb(w_n5802_0[1]),.din(n5802));
	jspl3 jspl3_w_n5806_0(.douta(w_n5806_0[0]),.doutb(w_n5806_0[1]),.doutc(w_n5806_0[2]),.din(n5806));
	jspl3 jspl3_w_n5808_0(.douta(w_n5808_0[0]),.doutb(w_n5808_0[1]),.doutc(w_n5808_0[2]),.din(n5808));
	jspl jspl_w_n5809_0(.douta(w_n5809_0[0]),.doutb(w_n5809_0[1]),.din(n5809));
	jspl3 jspl3_w_n5813_0(.douta(w_n5813_0[0]),.doutb(w_n5813_0[1]),.doutc(w_n5813_0[2]),.din(n5813));
	jspl3 jspl3_w_n5815_0(.douta(w_n5815_0[0]),.doutb(w_n5815_0[1]),.doutc(w_n5815_0[2]),.din(n5815));
	jspl jspl_w_n5816_0(.douta(w_n5816_0[0]),.doutb(w_n5816_0[1]),.din(n5816));
	jspl3 jspl3_w_n5820_0(.douta(w_n5820_0[0]),.doutb(w_n5820_0[1]),.doutc(w_n5820_0[2]),.din(n5820));
	jspl3 jspl3_w_n5823_0(.douta(w_n5823_0[0]),.doutb(w_n5823_0[1]),.doutc(w_n5823_0[2]),.din(n5823));
	jspl jspl_w_n5823_1(.douta(w_n5823_1[0]),.doutb(w_n5823_1[1]),.din(w_n5823_0[0]));
	jspl jspl_w_n5824_0(.douta(w_n5824_0[0]),.doutb(w_n5824_0[1]),.din(n5824));
	jspl jspl_w_n5827_0(.douta(w_n5827_0[0]),.doutb(w_n5827_0[1]),.din(n5827));
	jspl jspl_w_n5829_0(.douta(w_n5829_0[0]),.doutb(w_n5829_0[1]),.din(n5829));
	jspl jspl_w_n5834_0(.douta(w_n5834_0[0]),.doutb(w_n5834_0[1]),.din(n5834));
	jspl jspl_w_n5835_0(.douta(w_n5835_0[0]),.doutb(w_n5835_0[1]),.din(n5835));
	jspl3 jspl3_w_n5842_0(.douta(w_n5842_0[0]),.doutb(w_n5842_0[1]),.doutc(w_n5842_0[2]),.din(n5842));
	jspl3 jspl3_w_n5843_0(.douta(w_n5843_0[0]),.doutb(w_n5843_0[1]),.doutc(w_n5843_0[2]),.din(n5843));
	jspl jspl_w_n5843_1(.douta(w_n5843_1[0]),.doutb(w_n5843_1[1]),.din(w_n5843_0[0]));
	jspl jspl_w_n5844_0(.douta(w_n5844_0[0]),.doutb(w_n5844_0[1]),.din(n5844));
	jspl3 jspl3_w_n5845_0(.douta(w_n5845_0[0]),.doutb(w_n5845_0[1]),.doutc(w_n5845_0[2]),.din(n5845));
	jspl jspl_w_n5846_0(.douta(w_n5846_0[0]),.doutb(w_n5846_0[1]),.din(n5846));
	jspl3 jspl3_w_n5848_0(.douta(w_n5848_0[0]),.doutb(w_n5848_0[1]),.doutc(w_n5848_0[2]),.din(n5848));
	jspl jspl_w_n5849_0(.douta(w_n5849_0[0]),.doutb(w_n5849_0[1]),.din(n5849));
	jspl jspl_w_n5854_0(.douta(w_n5854_0[0]),.doutb(w_n5854_0[1]),.din(n5854));
	jspl jspl_w_n5888_0(.douta(w_n5888_0[0]),.doutb(w_n5888_0[1]),.din(n5888));
	jspl jspl_w_n5986_0(.douta(w_n5986_0[0]),.doutb(w_n5986_0[1]),.din(n5986));
	jspl jspl_w_n5987_0(.douta(w_n5987_0[0]),.doutb(w_n5987_0[1]),.din(n5987));
	jspl3 jspl3_w_n5989_0(.douta(w_n5989_0[0]),.doutb(w_n5989_0[1]),.doutc(w_n5989_0[2]),.din(n5989));
	jspl3 jspl3_w_n5989_1(.douta(w_n5989_1[0]),.doutb(w_n5989_1[1]),.doutc(w_n5989_1[2]),.din(w_n5989_0[0]));
	jspl3 jspl3_w_n5989_2(.douta(w_n5989_2[0]),.doutb(w_n5989_2[1]),.doutc(w_n5989_2[2]),.din(w_n5989_0[1]));
	jspl3 jspl3_w_n5989_3(.douta(w_n5989_3[0]),.doutb(w_n5989_3[1]),.doutc(w_n5989_3[2]),.din(w_n5989_0[2]));
	jspl3 jspl3_w_n5989_4(.douta(w_n5989_4[0]),.doutb(w_n5989_4[1]),.doutc(w_n5989_4[2]),.din(w_n5989_1[0]));
	jspl3 jspl3_w_n5989_5(.douta(w_n5989_5[0]),.doutb(w_n5989_5[1]),.doutc(w_n5989_5[2]),.din(w_n5989_1[1]));
	jspl3 jspl3_w_n5989_6(.douta(w_n5989_6[0]),.doutb(w_n5989_6[1]),.doutc(w_n5989_6[2]),.din(w_n5989_1[2]));
	jspl3 jspl3_w_n5989_7(.douta(w_n5989_7[0]),.doutb(w_n5989_7[1]),.doutc(w_n5989_7[2]),.din(w_n5989_2[0]));
	jspl3 jspl3_w_n5989_8(.douta(w_n5989_8[0]),.doutb(w_n5989_8[1]),.doutc(w_n5989_8[2]),.din(w_n5989_2[1]));
	jspl3 jspl3_w_n5989_9(.douta(w_n5989_9[0]),.doutb(w_n5989_9[1]),.doutc(w_n5989_9[2]),.din(w_n5989_2[2]));
	jspl3 jspl3_w_n5989_10(.douta(w_n5989_10[0]),.doutb(w_n5989_10[1]),.doutc(w_n5989_10[2]),.din(w_n5989_3[0]));
	jspl3 jspl3_w_n5989_11(.douta(w_n5989_11[0]),.doutb(w_n5989_11[1]),.doutc(w_n5989_11[2]),.din(w_n5989_3[1]));
	jspl3 jspl3_w_n5989_12(.douta(w_n5989_12[0]),.doutb(w_n5989_12[1]),.doutc(w_n5989_12[2]),.din(w_n5989_3[2]));
	jspl3 jspl3_w_n5989_13(.douta(w_n5989_13[0]),.doutb(w_n5989_13[1]),.doutc(w_n5989_13[2]),.din(w_n5989_4[0]));
	jspl3 jspl3_w_n5989_14(.douta(w_n5989_14[0]),.doutb(w_n5989_14[1]),.doutc(w_n5989_14[2]),.din(w_n5989_4[1]));
	jspl3 jspl3_w_n5989_15(.douta(w_n5989_15[0]),.doutb(w_n5989_15[1]),.doutc(w_n5989_15[2]),.din(w_n5989_4[2]));
	jspl3 jspl3_w_n5989_16(.douta(w_n5989_16[0]),.doutb(w_n5989_16[1]),.doutc(w_n5989_16[2]),.din(w_n5989_5[0]));
	jspl3 jspl3_w_n5989_17(.douta(w_n5989_17[0]),.doutb(w_n5989_17[1]),.doutc(w_n5989_17[2]),.din(w_n5989_5[1]));
	jspl3 jspl3_w_n5989_18(.douta(w_n5989_18[0]),.doutb(w_n5989_18[1]),.doutc(w_n5989_18[2]),.din(w_n5989_5[2]));
	jspl3 jspl3_w_n5989_19(.douta(w_n5989_19[0]),.doutb(w_n5989_19[1]),.doutc(w_n5989_19[2]),.din(w_n5989_6[0]));
	jspl3 jspl3_w_n5989_20(.douta(w_n5989_20[0]),.doutb(w_n5989_20[1]),.doutc(w_n5989_20[2]),.din(w_n5989_6[1]));
	jspl3 jspl3_w_n5989_21(.douta(w_n5989_21[0]),.doutb(w_n5989_21[1]),.doutc(w_n5989_21[2]),.din(w_n5989_6[2]));
	jspl3 jspl3_w_n5989_22(.douta(w_n5989_22[0]),.doutb(w_n5989_22[1]),.doutc(w_n5989_22[2]),.din(w_n5989_7[0]));
	jspl3 jspl3_w_n5989_23(.douta(w_n5989_23[0]),.doutb(w_n5989_23[1]),.doutc(w_n5989_23[2]),.din(w_n5989_7[1]));
	jspl3 jspl3_w_n5989_24(.douta(w_n5989_24[0]),.doutb(w_n5989_24[1]),.doutc(w_n5989_24[2]),.din(w_n5989_7[2]));
	jspl3 jspl3_w_n5989_25(.douta(w_n5989_25[0]),.doutb(w_n5989_25[1]),.doutc(w_n5989_25[2]),.din(w_n5989_8[0]));
	jspl3 jspl3_w_n5989_26(.douta(w_n5989_26[0]),.doutb(w_n5989_26[1]),.doutc(w_n5989_26[2]),.din(w_n5989_8[1]));
	jspl3 jspl3_w_n5989_27(.douta(w_n5989_27[0]),.doutb(w_n5989_27[1]),.doutc(w_n5989_27[2]),.din(w_n5989_8[2]));
	jspl3 jspl3_w_n5989_28(.douta(w_n5989_28[0]),.doutb(w_n5989_28[1]),.doutc(w_n5989_28[2]),.din(w_n5989_9[0]));
	jspl3 jspl3_w_n5989_29(.douta(w_n5989_29[0]),.doutb(w_n5989_29[1]),.doutc(w_n5989_29[2]),.din(w_n5989_9[1]));
	jspl3 jspl3_w_n5989_30(.douta(w_n5989_30[0]),.doutb(w_n5989_30[1]),.doutc(w_n5989_30[2]),.din(w_n5989_9[2]));
	jspl3 jspl3_w_n5989_31(.douta(w_n5989_31[0]),.doutb(w_n5989_31[1]),.doutc(w_n5989_31[2]),.din(w_n5989_10[0]));
	jspl3 jspl3_w_n5989_32(.douta(w_n5989_32[0]),.doutb(w_n5989_32[1]),.doutc(w_n5989_32[2]),.din(w_n5989_10[1]));
	jspl3 jspl3_w_n5989_33(.douta(w_n5989_33[0]),.doutb(w_n5989_33[1]),.doutc(w_n5989_33[2]),.din(w_n5989_10[2]));
	jspl3 jspl3_w_n5989_34(.douta(w_n5989_34[0]),.doutb(w_n5989_34[1]),.doutc(w_n5989_34[2]),.din(w_n5989_11[0]));
	jspl3 jspl3_w_n5989_35(.douta(w_n5989_35[0]),.doutb(w_n5989_35[1]),.doutc(w_n5989_35[2]),.din(w_n5989_11[1]));
	jspl3 jspl3_w_n5989_36(.douta(w_n5989_36[0]),.doutb(w_n5989_36[1]),.doutc(w_n5989_36[2]),.din(w_n5989_11[2]));
	jspl3 jspl3_w_n5989_37(.douta(w_n5989_37[0]),.doutb(w_n5989_37[1]),.doutc(w_n5989_37[2]),.din(w_n5989_12[0]));
	jspl3 jspl3_w_n5989_38(.douta(w_n5989_38[0]),.doutb(w_n5989_38[1]),.doutc(w_n5989_38[2]),.din(w_n5989_12[1]));
	jspl3 jspl3_w_n5989_39(.douta(w_n5989_39[0]),.doutb(w_n5989_39[1]),.doutc(w_n5989_39[2]),.din(w_n5989_12[2]));
	jspl3 jspl3_w_n5989_40(.douta(w_n5989_40[0]),.doutb(w_n5989_40[1]),.doutc(w_n5989_40[2]),.din(w_n5989_13[0]));
	jspl3 jspl3_w_n5989_41(.douta(w_n5989_41[0]),.doutb(w_n5989_41[1]),.doutc(w_n5989_41[2]),.din(w_n5989_13[1]));
	jspl jspl_w_n5989_42(.douta(w_n5989_42[0]),.doutb(w_n5989_42[1]),.din(w_n5989_13[2]));
	jspl3 jspl3_w_n5993_0(.douta(w_n5993_0[0]),.doutb(w_n5993_0[1]),.doutc(w_n5993_0[2]),.din(n5993));
	jspl jspl_w_n5994_0(.douta(w_n5994_0[0]),.doutb(w_n5994_0[1]),.din(n5994));
	jspl jspl_w_n5996_0(.douta(w_n5996_0[0]),.doutb(w_n5996_0[1]),.din(n5996));
	jspl jspl_w_n6001_0(.douta(w_n6001_0[0]),.doutb(w_n6001_0[1]),.din(n6001));
	jspl jspl_w_n6002_0(.douta(w_n6002_0[0]),.doutb(w_n6002_0[1]),.din(n6002));
	jspl3 jspl3_w_n6004_0(.douta(w_n6004_0[0]),.doutb(w_n6004_0[1]),.doutc(w_n6004_0[2]),.din(n6004));
	jspl jspl_w_n6005_0(.douta(w_n6005_0[0]),.doutb(w_n6005_0[1]),.din(n6005));
	jspl jspl_w_n6009_0(.douta(w_n6009_0[0]),.doutb(w_n6009_0[1]),.din(n6009));
	jspl3 jspl3_w_n6011_0(.douta(w_n6011_0[0]),.doutb(w_n6011_0[1]),.doutc(w_n6011_0[2]),.din(n6011));
	jspl jspl_w_n6012_0(.douta(w_n6012_0[0]),.doutb(w_n6012_0[1]),.din(n6012));
	jspl jspl_w_n6016_0(.douta(w_n6016_0[0]),.doutb(w_n6016_0[1]),.din(n6016));
	jspl jspl_w_n6017_0(.douta(w_n6017_0[0]),.doutb(w_n6017_0[1]),.din(n6017));
	jspl3 jspl3_w_n6019_0(.douta(w_n6019_0[0]),.doutb(w_n6019_0[1]),.doutc(w_n6019_0[2]),.din(n6019));
	jspl jspl_w_n6020_0(.douta(w_n6020_0[0]),.doutb(w_n6020_0[1]),.din(n6020));
	jspl jspl_w_n6024_0(.douta(w_n6024_0[0]),.doutb(w_n6024_0[1]),.din(n6024));
	jspl3 jspl3_w_n6026_0(.douta(w_n6026_0[0]),.doutb(w_n6026_0[1]),.doutc(w_n6026_0[2]),.din(n6026));
	jspl jspl_w_n6027_0(.douta(w_n6027_0[0]),.doutb(w_n6027_0[1]),.din(n6027));
	jspl jspl_w_n6031_0(.douta(w_n6031_0[0]),.doutb(w_n6031_0[1]),.din(n6031));
	jspl jspl_w_n6032_0(.douta(w_n6032_0[0]),.doutb(w_n6032_0[1]),.din(n6032));
	jspl3 jspl3_w_n6034_0(.douta(w_n6034_0[0]),.doutb(w_n6034_0[1]),.doutc(w_n6034_0[2]),.din(n6034));
	jspl jspl_w_n6035_0(.douta(w_n6035_0[0]),.doutb(w_n6035_0[1]),.din(n6035));
	jspl jspl_w_n6039_0(.douta(w_n6039_0[0]),.doutb(w_n6039_0[1]),.din(n6039));
	jspl3 jspl3_w_n6041_0(.douta(w_n6041_0[0]),.doutb(w_n6041_0[1]),.doutc(w_n6041_0[2]),.din(n6041));
	jspl jspl_w_n6042_0(.douta(w_n6042_0[0]),.doutb(w_n6042_0[1]),.din(n6042));
	jspl jspl_w_n6046_0(.douta(w_n6046_0[0]),.doutb(w_n6046_0[1]),.din(n6046));
	jspl jspl_w_n6047_0(.douta(w_n6047_0[0]),.doutb(w_n6047_0[1]),.din(n6047));
	jspl3 jspl3_w_n6049_0(.douta(w_n6049_0[0]),.doutb(w_n6049_0[1]),.doutc(w_n6049_0[2]),.din(n6049));
	jspl jspl_w_n6050_0(.douta(w_n6050_0[0]),.doutb(w_n6050_0[1]),.din(n6050));
	jspl jspl_w_n6054_0(.douta(w_n6054_0[0]),.doutb(w_n6054_0[1]),.din(n6054));
	jspl3 jspl3_w_n6056_0(.douta(w_n6056_0[0]),.doutb(w_n6056_0[1]),.doutc(w_n6056_0[2]),.din(n6056));
	jspl jspl_w_n6057_0(.douta(w_n6057_0[0]),.doutb(w_n6057_0[1]),.din(n6057));
	jspl jspl_w_n6061_0(.douta(w_n6061_0[0]),.doutb(w_n6061_0[1]),.din(n6061));
	jspl3 jspl3_w_n6063_0(.douta(w_n6063_0[0]),.doutb(w_n6063_0[1]),.doutc(w_n6063_0[2]),.din(n6063));
	jspl jspl_w_n6064_0(.douta(w_n6064_0[0]),.doutb(w_n6064_0[1]),.din(n6064));
	jspl jspl_w_n6068_0(.douta(w_n6068_0[0]),.doutb(w_n6068_0[1]),.din(n6068));
	jspl3 jspl3_w_n6070_0(.douta(w_n6070_0[0]),.doutb(w_n6070_0[1]),.doutc(w_n6070_0[2]),.din(n6070));
	jspl jspl_w_n6071_0(.douta(w_n6071_0[0]),.doutb(w_n6071_0[1]),.din(n6071));
	jspl jspl_w_n6075_0(.douta(w_n6075_0[0]),.doutb(w_n6075_0[1]),.din(n6075));
	jspl jspl_w_n6076_0(.douta(w_n6076_0[0]),.doutb(w_n6076_0[1]),.din(n6076));
	jspl3 jspl3_w_n6078_0(.douta(w_n6078_0[0]),.doutb(w_n6078_0[1]),.doutc(w_n6078_0[2]),.din(n6078));
	jspl jspl_w_n6079_0(.douta(w_n6079_0[0]),.doutb(w_n6079_0[1]),.din(n6079));
	jspl jspl_w_n6083_0(.douta(w_n6083_0[0]),.doutb(w_n6083_0[1]),.din(n6083));
	jspl jspl_w_n6084_0(.douta(w_n6084_0[0]),.doutb(w_n6084_0[1]),.din(n6084));
	jspl3 jspl3_w_n6086_0(.douta(w_n6086_0[0]),.doutb(w_n6086_0[1]),.doutc(w_n6086_0[2]),.din(n6086));
	jspl jspl_w_n6087_0(.douta(w_n6087_0[0]),.doutb(w_n6087_0[1]),.din(n6087));
	jspl jspl_w_n6091_0(.douta(w_n6091_0[0]),.doutb(w_n6091_0[1]),.din(n6091));
	jspl jspl_w_n6092_0(.douta(w_n6092_0[0]),.doutb(w_n6092_0[1]),.din(n6092));
	jspl3 jspl3_w_n6094_0(.douta(w_n6094_0[0]),.doutb(w_n6094_0[1]),.doutc(w_n6094_0[2]),.din(n6094));
	jspl jspl_w_n6095_0(.douta(w_n6095_0[0]),.doutb(w_n6095_0[1]),.din(n6095));
	jspl jspl_w_n6099_0(.douta(w_n6099_0[0]),.doutb(w_n6099_0[1]),.din(n6099));
	jspl3 jspl3_w_n6101_0(.douta(w_n6101_0[0]),.doutb(w_n6101_0[1]),.doutc(w_n6101_0[2]),.din(n6101));
	jspl jspl_w_n6102_0(.douta(w_n6102_0[0]),.doutb(w_n6102_0[1]),.din(n6102));
	jspl jspl_w_n6106_0(.douta(w_n6106_0[0]),.doutb(w_n6106_0[1]),.din(n6106));
	jspl jspl_w_n6107_0(.douta(w_n6107_0[0]),.doutb(w_n6107_0[1]),.din(n6107));
	jspl3 jspl3_w_n6109_0(.douta(w_n6109_0[0]),.doutb(w_n6109_0[1]),.doutc(w_n6109_0[2]),.din(n6109));
	jspl jspl_w_n6110_0(.douta(w_n6110_0[0]),.doutb(w_n6110_0[1]),.din(n6110));
	jspl jspl_w_n6114_0(.douta(w_n6114_0[0]),.doutb(w_n6114_0[1]),.din(n6114));
	jspl3 jspl3_w_n6116_0(.douta(w_n6116_0[0]),.doutb(w_n6116_0[1]),.doutc(w_n6116_0[2]),.din(n6116));
	jspl jspl_w_n6117_0(.douta(w_n6117_0[0]),.doutb(w_n6117_0[1]),.din(n6117));
	jspl jspl_w_n6121_0(.douta(w_n6121_0[0]),.doutb(w_n6121_0[1]),.din(n6121));
	jspl jspl_w_n6122_0(.douta(w_n6122_0[0]),.doutb(w_n6122_0[1]),.din(n6122));
	jspl3 jspl3_w_n6124_0(.douta(w_n6124_0[0]),.doutb(w_n6124_0[1]),.doutc(w_n6124_0[2]),.din(n6124));
	jspl jspl_w_n6125_0(.douta(w_n6125_0[0]),.doutb(w_n6125_0[1]),.din(n6125));
	jspl jspl_w_n6129_0(.douta(w_n6129_0[0]),.doutb(w_n6129_0[1]),.din(n6129));
	jspl3 jspl3_w_n6131_0(.douta(w_n6131_0[0]),.doutb(w_n6131_0[1]),.doutc(w_n6131_0[2]),.din(n6131));
	jspl jspl_w_n6132_0(.douta(w_n6132_0[0]),.doutb(w_n6132_0[1]),.din(n6132));
	jspl jspl_w_n6136_0(.douta(w_n6136_0[0]),.doutb(w_n6136_0[1]),.din(n6136));
	jspl3 jspl3_w_n6138_0(.douta(w_n6138_0[0]),.doutb(w_n6138_0[1]),.doutc(w_n6138_0[2]),.din(n6138));
	jspl jspl_w_n6139_0(.douta(w_n6139_0[0]),.doutb(w_n6139_0[1]),.din(n6139));
	jspl jspl_w_n6143_0(.douta(w_n6143_0[0]),.doutb(w_n6143_0[1]),.din(n6143));
	jspl jspl_w_n6144_0(.douta(w_n6144_0[0]),.doutb(w_n6144_0[1]),.din(n6144));
	jspl3 jspl3_w_n6146_0(.douta(w_n6146_0[0]),.doutb(w_n6146_0[1]),.doutc(w_n6146_0[2]),.din(n6146));
	jspl jspl_w_n6147_0(.douta(w_n6147_0[0]),.doutb(w_n6147_0[1]),.din(n6147));
	jspl jspl_w_n6151_0(.douta(w_n6151_0[0]),.doutb(w_n6151_0[1]),.din(n6151));
	jspl jspl_w_n6152_0(.douta(w_n6152_0[0]),.doutb(w_n6152_0[1]),.din(n6152));
	jspl3 jspl3_w_n6154_0(.douta(w_n6154_0[0]),.doutb(w_n6154_0[1]),.doutc(w_n6154_0[2]),.din(n6154));
	jspl jspl_w_n6155_0(.douta(w_n6155_0[0]),.doutb(w_n6155_0[1]),.din(n6155));
	jspl jspl_w_n6159_0(.douta(w_n6159_0[0]),.doutb(w_n6159_0[1]),.din(n6159));
	jspl3 jspl3_w_n6161_0(.douta(w_n6161_0[0]),.doutb(w_n6161_0[1]),.doutc(w_n6161_0[2]),.din(n6161));
	jspl jspl_w_n6162_0(.douta(w_n6162_0[0]),.doutb(w_n6162_0[1]),.din(n6162));
	jspl3 jspl3_w_n6166_0(.douta(w_n6166_0[0]),.doutb(w_n6166_0[1]),.doutc(w_n6166_0[2]),.din(n6166));
	jspl3 jspl3_w_n6169_0(.douta(w_n6169_0[0]),.doutb(w_n6169_0[1]),.doutc(w_n6169_0[2]),.din(n6169));
	jspl jspl_w_n6170_0(.douta(w_n6170_0[0]),.doutb(w_n6170_0[1]),.din(n6170));
	jspl jspl_w_n6174_0(.douta(w_n6174_0[0]),.doutb(w_n6174_0[1]),.din(n6174));
	jspl3 jspl3_w_n6176_0(.douta(w_n6176_0[0]),.doutb(w_n6176_0[1]),.doutc(w_n6176_0[2]),.din(n6176));
	jspl jspl_w_n6177_0(.douta(w_n6177_0[0]),.doutb(w_n6177_0[1]),.din(n6177));
	jspl jspl_w_n6181_0(.douta(w_n6181_0[0]),.doutb(w_n6181_0[1]),.din(n6181));
	jspl jspl_w_n6182_0(.douta(w_n6182_0[0]),.doutb(w_n6182_0[1]),.din(n6182));
	jspl3 jspl3_w_n6184_0(.douta(w_n6184_0[0]),.doutb(w_n6184_0[1]),.doutc(w_n6184_0[2]),.din(n6184));
	jspl jspl_w_n6185_0(.douta(w_n6185_0[0]),.doutb(w_n6185_0[1]),.din(n6185));
	jspl jspl_w_n6189_0(.douta(w_n6189_0[0]),.doutb(w_n6189_0[1]),.din(n6189));
	jspl jspl_w_n6190_0(.douta(w_n6190_0[0]),.doutb(w_n6190_0[1]),.din(n6190));
	jspl3 jspl3_w_n6192_0(.douta(w_n6192_0[0]),.doutb(w_n6192_0[1]),.doutc(w_n6192_0[2]),.din(n6192));
	jspl jspl_w_n6193_0(.douta(w_n6193_0[0]),.doutb(w_n6193_0[1]),.din(n6193));
	jspl3 jspl3_w_n6197_0(.douta(w_n6197_0[0]),.doutb(w_n6197_0[1]),.doutc(w_n6197_0[2]),.din(n6197));
	jspl jspl_w_n6200_0(.douta(w_n6200_0[0]),.doutb(w_n6200_0[1]),.din(n6200));
	jspl3 jspl3_w_n6201_0(.douta(w_n6201_0[0]),.doutb(w_n6201_0[1]),.doutc(w_n6201_0[2]),.din(n6201));
	jspl jspl_w_n6201_1(.douta(w_n6201_1[0]),.doutb(w_n6201_1[1]),.din(w_n6201_0[0]));
	jspl3 jspl3_w_n6202_0(.douta(w_n6202_0[0]),.doutb(w_n6202_0[1]),.doutc(w_n6202_0[2]),.din(n6202));
	jspl jspl_w_n6204_0(.douta(w_n6204_0[0]),.doutb(w_n6204_0[1]),.din(n6204));
	jspl jspl_w_n6239_0(.douta(w_n6239_0[0]),.doutb(w_n6239_0[1]),.din(n6239));
	jspl jspl_w_n6246_0(.douta(w_n6246_0[0]),.doutb(w_n6246_0[1]),.din(n6246));
	jspl jspl_w_n6253_0(.douta(w_n6253_0[0]),.doutb(w_n6253_0[1]),.din(n6253));
	jspl jspl_w_n6260_0(.douta(w_n6260_0[0]),.doutb(w_n6260_0[1]),.din(n6260));
	jspl jspl_w_n6267_0(.douta(w_n6267_0[0]),.doutb(w_n6267_0[1]),.din(n6267));
	jspl jspl_w_n6271_0(.douta(w_n6271_0[0]),.doutb(w_n6271_0[1]),.din(n6271));
	jspl jspl_w_n6275_0(.douta(w_n6275_0[0]),.doutb(w_n6275_0[1]),.din(n6275));
	jspl jspl_w_n6288_0(.douta(w_n6288_0[0]),.doutb(w_n6288_0[1]),.din(n6288));
	jspl jspl_w_n6295_0(.douta(w_n6295_0[0]),.doutb(w_n6295_0[1]),.din(n6295));
	jspl jspl_w_n6302_0(.douta(w_n6302_0[0]),.doutb(w_n6302_0[1]),.din(n6302));
	jspl jspl_w_n6306_0(.douta(w_n6306_0[0]),.doutb(w_n6306_0[1]),.din(n6306));
	jspl jspl_w_n6316_0(.douta(w_n6316_0[0]),.doutb(w_n6316_0[1]),.din(n6316));
	jspl jspl_w_n6323_0(.douta(w_n6323_0[0]),.doutb(w_n6323_0[1]),.din(n6323));
	jspl jspl_w_n6334_0(.douta(w_n6334_0[0]),.doutb(w_n6334_0[1]),.din(n6334));
	jspl jspl_w_n6335_0(.douta(w_n6335_0[0]),.doutb(w_n6335_0[1]),.din(n6335));
	jspl jspl_w_n6336_0(.douta(w_n6336_0[0]),.doutb(w_n6336_0[1]),.din(n6336));
	jspl jspl_w_n6338_0(.douta(w_n6338_0[0]),.doutb(w_n6338_0[1]),.din(n6338));
	jspl jspl_w_n6340_0(.douta(w_n6340_0[0]),.doutb(w_n6340_0[1]),.din(n6340));
	jspl jspl_w_n6343_0(.douta(w_n6343_0[0]),.doutb(w_n6343_0[1]),.din(n6343));
	jspl jspl_w_n6344_0(.douta(w_n6344_0[0]),.doutb(w_n6344_0[1]),.din(n6344));
	jspl jspl_w_n6345_0(.douta(w_n6345_0[0]),.doutb(w_n6345_0[1]),.din(n6345));
	jspl jspl_w_n6348_0(.douta(w_n6348_0[0]),.doutb(w_n6348_0[1]),.din(n6348));
	jspl jspl_w_n6349_0(.douta(w_n6349_0[0]),.doutb(w_n6349_0[1]),.din(n6349));
	jspl jspl_w_n6355_0(.douta(w_n6355_0[0]),.doutb(w_n6355_0[1]),.din(n6355));
	jspl3 jspl3_w_n6357_0(.douta(w_n6357_0[0]),.doutb(w_n6357_0[1]),.doutc(w_n6357_0[2]),.din(n6357));
	jspl3 jspl3_w_n6357_1(.douta(w_n6357_1[0]),.doutb(w_n6357_1[1]),.doutc(w_n6357_1[2]),.din(w_n6357_0[0]));
	jspl3 jspl3_w_n6357_2(.douta(w_n6357_2[0]),.doutb(w_n6357_2[1]),.doutc(w_n6357_2[2]),.din(w_n6357_0[1]));
	jspl3 jspl3_w_n6357_3(.douta(w_n6357_3[0]),.doutb(w_n6357_3[1]),.doutc(w_n6357_3[2]),.din(w_n6357_0[2]));
	jspl3 jspl3_w_n6357_4(.douta(w_n6357_4[0]),.doutb(w_n6357_4[1]),.doutc(w_n6357_4[2]),.din(w_n6357_1[0]));
	jspl3 jspl3_w_n6357_5(.douta(w_n6357_5[0]),.doutb(w_n6357_5[1]),.doutc(w_n6357_5[2]),.din(w_n6357_1[1]));
	jspl3 jspl3_w_n6357_6(.douta(w_n6357_6[0]),.doutb(w_n6357_6[1]),.doutc(w_n6357_6[2]),.din(w_n6357_1[2]));
	jspl3 jspl3_w_n6357_7(.douta(w_n6357_7[0]),.doutb(w_n6357_7[1]),.doutc(w_n6357_7[2]),.din(w_n6357_2[0]));
	jspl3 jspl3_w_n6357_8(.douta(w_n6357_8[0]),.doutb(w_n6357_8[1]),.doutc(w_n6357_8[2]),.din(w_n6357_2[1]));
	jspl3 jspl3_w_n6357_9(.douta(w_n6357_9[0]),.doutb(w_n6357_9[1]),.doutc(w_n6357_9[2]),.din(w_n6357_2[2]));
	jspl3 jspl3_w_n6357_10(.douta(w_n6357_10[0]),.doutb(w_n6357_10[1]),.doutc(w_n6357_10[2]),.din(w_n6357_3[0]));
	jspl3 jspl3_w_n6357_11(.douta(w_n6357_11[0]),.doutb(w_n6357_11[1]),.doutc(w_n6357_11[2]),.din(w_n6357_3[1]));
	jspl3 jspl3_w_n6357_12(.douta(w_n6357_12[0]),.doutb(w_n6357_12[1]),.doutc(w_n6357_12[2]),.din(w_n6357_3[2]));
	jspl3 jspl3_w_n6357_13(.douta(w_n6357_13[0]),.doutb(w_n6357_13[1]),.doutc(w_n6357_13[2]),.din(w_n6357_4[0]));
	jspl3 jspl3_w_n6357_14(.douta(w_n6357_14[0]),.doutb(w_n6357_14[1]),.doutc(w_n6357_14[2]),.din(w_n6357_4[1]));
	jspl3 jspl3_w_n6357_15(.douta(w_n6357_15[0]),.doutb(w_n6357_15[1]),.doutc(w_n6357_15[2]),.din(w_n6357_4[2]));
	jspl3 jspl3_w_n6357_16(.douta(w_n6357_16[0]),.doutb(w_n6357_16[1]),.doutc(w_n6357_16[2]),.din(w_n6357_5[0]));
	jspl3 jspl3_w_n6357_17(.douta(w_n6357_17[0]),.doutb(w_n6357_17[1]),.doutc(w_n6357_17[2]),.din(w_n6357_5[1]));
	jspl3 jspl3_w_n6357_18(.douta(w_n6357_18[0]),.doutb(w_n6357_18[1]),.doutc(w_n6357_18[2]),.din(w_n6357_5[2]));
	jspl3 jspl3_w_n6357_19(.douta(w_n6357_19[0]),.doutb(w_n6357_19[1]),.doutc(w_n6357_19[2]),.din(w_n6357_6[0]));
	jspl3 jspl3_w_n6357_20(.douta(w_n6357_20[0]),.doutb(w_n6357_20[1]),.doutc(w_n6357_20[2]),.din(w_n6357_6[1]));
	jspl3 jspl3_w_n6357_21(.douta(w_n6357_21[0]),.doutb(w_n6357_21[1]),.doutc(w_n6357_21[2]),.din(w_n6357_6[2]));
	jspl3 jspl3_w_n6357_22(.douta(w_n6357_22[0]),.doutb(w_n6357_22[1]),.doutc(w_n6357_22[2]),.din(w_n6357_7[0]));
	jspl3 jspl3_w_n6357_23(.douta(w_n6357_23[0]),.doutb(w_n6357_23[1]),.doutc(w_n6357_23[2]),.din(w_n6357_7[1]));
	jspl3 jspl3_w_n6357_24(.douta(w_n6357_24[0]),.doutb(w_n6357_24[1]),.doutc(w_n6357_24[2]),.din(w_n6357_7[2]));
	jspl3 jspl3_w_n6357_25(.douta(w_n6357_25[0]),.doutb(w_n6357_25[1]),.doutc(w_n6357_25[2]),.din(w_n6357_8[0]));
	jspl3 jspl3_w_n6357_26(.douta(w_n6357_26[0]),.doutb(w_n6357_26[1]),.doutc(w_n6357_26[2]),.din(w_n6357_8[1]));
	jspl3 jspl3_w_n6357_27(.douta(w_n6357_27[0]),.doutb(w_n6357_27[1]),.doutc(w_n6357_27[2]),.din(w_n6357_8[2]));
	jspl3 jspl3_w_n6357_28(.douta(w_n6357_28[0]),.doutb(w_n6357_28[1]),.doutc(w_n6357_28[2]),.din(w_n6357_9[0]));
	jspl3 jspl3_w_n6357_29(.douta(w_n6357_29[0]),.doutb(w_n6357_29[1]),.doutc(w_n6357_29[2]),.din(w_n6357_9[1]));
	jspl3 jspl3_w_n6357_30(.douta(w_n6357_30[0]),.doutb(w_n6357_30[1]),.doutc(w_n6357_30[2]),.din(w_n6357_9[2]));
	jspl3 jspl3_w_n6357_31(.douta(w_n6357_31[0]),.doutb(w_n6357_31[1]),.doutc(w_n6357_31[2]),.din(w_n6357_10[0]));
	jspl3 jspl3_w_n6357_32(.douta(w_n6357_32[0]),.doutb(w_n6357_32[1]),.doutc(w_n6357_32[2]),.din(w_n6357_10[1]));
	jspl3 jspl3_w_n6357_33(.douta(w_n6357_33[0]),.doutb(w_n6357_33[1]),.doutc(w_n6357_33[2]),.din(w_n6357_10[2]));
	jspl3 jspl3_w_n6357_34(.douta(w_n6357_34[0]),.doutb(w_n6357_34[1]),.doutc(w_n6357_34[2]),.din(w_n6357_11[0]));
	jspl3 jspl3_w_n6357_35(.douta(w_n6357_35[0]),.doutb(w_n6357_35[1]),.doutc(w_n6357_35[2]),.din(w_n6357_11[1]));
	jspl3 jspl3_w_n6357_36(.douta(w_n6357_36[0]),.doutb(w_n6357_36[1]),.doutc(w_n6357_36[2]),.din(w_n6357_11[2]));
	jspl3 jspl3_w_n6357_37(.douta(w_n6357_37[0]),.doutb(w_n6357_37[1]),.doutc(w_n6357_37[2]),.din(w_n6357_12[0]));
	jspl3 jspl3_w_n6357_38(.douta(w_n6357_38[0]),.doutb(w_n6357_38[1]),.doutc(w_n6357_38[2]),.din(w_n6357_12[1]));
	jspl3 jspl3_w_n6357_39(.douta(w_n6357_39[0]),.doutb(w_n6357_39[1]),.doutc(w_n6357_39[2]),.din(w_n6357_12[2]));
	jspl3 jspl3_w_n6357_40(.douta(w_n6357_40[0]),.doutb(w_n6357_40[1]),.doutc(w_n6357_40[2]),.din(w_n6357_13[0]));
	jspl3 jspl3_w_n6357_41(.douta(w_n6357_41[0]),.doutb(w_n6357_41[1]),.doutc(w_n6357_41[2]),.din(w_n6357_13[1]));
	jspl3 jspl3_w_n6357_42(.douta(w_n6357_42[0]),.doutb(w_n6357_42[1]),.doutc(w_n6357_42[2]),.din(w_n6357_13[2]));
	jspl3 jspl3_w_n6357_43(.douta(w_n6357_43[0]),.doutb(w_n6357_43[1]),.doutc(w_n6357_43[2]),.din(w_n6357_14[0]));
	jspl3 jspl3_w_n6357_44(.douta(w_n6357_44[0]),.doutb(w_n6357_44[1]),.doutc(w_n6357_44[2]),.din(w_n6357_14[1]));
	jspl3 jspl3_w_n6357_45(.douta(w_n6357_45[0]),.doutb(w_n6357_45[1]),.doutc(w_n6357_45[2]),.din(w_n6357_14[2]));
	jspl3 jspl3_w_n6357_46(.douta(w_n6357_46[0]),.doutb(w_n6357_46[1]),.doutc(w_n6357_46[2]),.din(w_n6357_15[0]));
	jspl3 jspl3_w_n6357_47(.douta(w_n6357_47[0]),.doutb(w_n6357_47[1]),.doutc(w_n6357_47[2]),.din(w_n6357_15[1]));
	jspl3 jspl3_w_n6357_48(.douta(w_n6357_48[0]),.doutb(w_n6357_48[1]),.doutc(w_n6357_48[2]),.din(w_n6357_15[2]));
	jspl3 jspl3_w_n6357_49(.douta(w_n6357_49[0]),.doutb(w_n6357_49[1]),.doutc(w_n6357_49[2]),.din(w_n6357_16[0]));
	jspl3 jspl3_w_n6357_50(.douta(w_n6357_50[0]),.doutb(w_n6357_50[1]),.doutc(w_n6357_50[2]),.din(w_n6357_16[1]));
	jspl3 jspl3_w_n6357_51(.douta(w_n6357_51[0]),.doutb(w_n6357_51[1]),.doutc(w_n6357_51[2]),.din(w_n6357_16[2]));
	jspl3 jspl3_w_n6357_52(.douta(w_n6357_52[0]),.doutb(w_n6357_52[1]),.doutc(w_n6357_52[2]),.din(w_n6357_17[0]));
	jspl3 jspl3_w_n6357_53(.douta(w_n6357_53[0]),.doutb(w_n6357_53[1]),.doutc(w_n6357_53[2]),.din(w_n6357_17[1]));
	jspl3 jspl3_w_n6357_54(.douta(w_n6357_54[0]),.doutb(w_n6357_54[1]),.doutc(w_n6357_54[2]),.din(w_n6357_17[2]));
	jspl jspl_w_n6360_0(.douta(w_n6360_0[0]),.doutb(w_n6360_0[1]),.din(n6360));
	jspl3 jspl3_w_n6361_0(.douta(w_n6361_0[0]),.doutb(w_n6361_0[1]),.doutc(w_n6361_0[2]),.din(n6361));
	jspl3 jspl3_w_n6362_0(.douta(w_n6362_0[0]),.doutb(w_n6362_0[1]),.doutc(w_n6362_0[2]),.din(n6362));
	jspl3 jspl3_w_n6362_1(.douta(w_n6362_1[0]),.doutb(w_n6362_1[1]),.doutc(w_n6362_1[2]),.din(w_n6362_0[0]));
	jspl jspl_w_n6363_0(.douta(w_n6363_0[0]),.doutb(w_n6363_0[1]),.din(n6363));
	jspl3 jspl3_w_n6364_0(.douta(w_n6364_0[0]),.doutb(w_n6364_0[1]),.doutc(w_n6364_0[2]),.din(n6364));
	jspl jspl_w_n6365_0(.douta(w_n6365_0[0]),.doutb(w_n6365_0[1]),.din(n6365));
	jspl3 jspl3_w_n6368_0(.douta(w_n6368_0[0]),.doutb(w_n6368_0[1]),.doutc(w_n6368_0[2]),.din(n6368));
	jspl jspl_w_n6369_0(.douta(w_n6369_0[0]),.doutb(w_n6369_0[1]),.din(n6369));
	jspl3 jspl3_w_n6376_0(.douta(w_n6376_0[0]),.doutb(w_n6376_0[1]),.doutc(w_n6376_0[2]),.din(n6376));
	jspl jspl_w_n6377_0(.douta(w_n6377_0[0]),.doutb(w_n6377_0[1]),.din(n6377));
	jspl jspl_w_n6380_0(.douta(w_n6380_0[0]),.doutb(w_n6380_0[1]),.din(n6380));
	jspl jspl_w_n6385_0(.douta(w_n6385_0[0]),.doutb(w_n6385_0[1]),.din(n6385));
	jspl3 jspl3_w_n6387_0(.douta(w_n6387_0[0]),.doutb(w_n6387_0[1]),.doutc(w_n6387_0[2]),.din(n6387));
	jspl jspl_w_n6388_0(.douta(w_n6388_0[0]),.doutb(w_n6388_0[1]),.din(n6388));
	jspl3 jspl3_w_n6392_0(.douta(w_n6392_0[0]),.doutb(w_n6392_0[1]),.doutc(w_n6392_0[2]),.din(n6392));
	jspl3 jspl3_w_n6395_0(.douta(w_n6395_0[0]),.doutb(w_n6395_0[1]),.doutc(w_n6395_0[2]),.din(n6395));
	jspl jspl_w_n6396_0(.douta(w_n6396_0[0]),.doutb(w_n6396_0[1]),.din(n6396));
	jspl3 jspl3_w_n6400_0(.douta(w_n6400_0[0]),.doutb(w_n6400_0[1]),.doutc(w_n6400_0[2]),.din(n6400));
	jspl3 jspl3_w_n6402_0(.douta(w_n6402_0[0]),.doutb(w_n6402_0[1]),.doutc(w_n6402_0[2]),.din(n6402));
	jspl jspl_w_n6403_0(.douta(w_n6403_0[0]),.doutb(w_n6403_0[1]),.din(n6403));
	jspl3 jspl3_w_n6407_0(.douta(w_n6407_0[0]),.doutb(w_n6407_0[1]),.doutc(w_n6407_0[2]),.din(n6407));
	jspl3 jspl3_w_n6410_0(.douta(w_n6410_0[0]),.doutb(w_n6410_0[1]),.doutc(w_n6410_0[2]),.din(n6410));
	jspl jspl_w_n6411_0(.douta(w_n6411_0[0]),.doutb(w_n6411_0[1]),.din(n6411));
	jspl3 jspl3_w_n6415_0(.douta(w_n6415_0[0]),.doutb(w_n6415_0[1]),.doutc(w_n6415_0[2]),.din(n6415));
	jspl3 jspl3_w_n6417_0(.douta(w_n6417_0[0]),.doutb(w_n6417_0[1]),.doutc(w_n6417_0[2]),.din(n6417));
	jspl jspl_w_n6418_0(.douta(w_n6418_0[0]),.doutb(w_n6418_0[1]),.din(n6418));
	jspl3 jspl3_w_n6422_0(.douta(w_n6422_0[0]),.doutb(w_n6422_0[1]),.doutc(w_n6422_0[2]),.din(n6422));
	jspl3 jspl3_w_n6425_0(.douta(w_n6425_0[0]),.doutb(w_n6425_0[1]),.doutc(w_n6425_0[2]),.din(n6425));
	jspl jspl_w_n6426_0(.douta(w_n6426_0[0]),.doutb(w_n6426_0[1]),.din(n6426));
	jspl3 jspl3_w_n6430_0(.douta(w_n6430_0[0]),.doutb(w_n6430_0[1]),.doutc(w_n6430_0[2]),.din(n6430));
	jspl3 jspl3_w_n6432_0(.douta(w_n6432_0[0]),.doutb(w_n6432_0[1]),.doutc(w_n6432_0[2]),.din(n6432));
	jspl jspl_w_n6433_0(.douta(w_n6433_0[0]),.doutb(w_n6433_0[1]),.din(n6433));
	jspl3 jspl3_w_n6437_0(.douta(w_n6437_0[0]),.doutb(w_n6437_0[1]),.doutc(w_n6437_0[2]),.din(n6437));
	jspl3 jspl3_w_n6440_0(.douta(w_n6440_0[0]),.doutb(w_n6440_0[1]),.doutc(w_n6440_0[2]),.din(n6440));
	jspl jspl_w_n6441_0(.douta(w_n6441_0[0]),.doutb(w_n6441_0[1]),.din(n6441));
	jspl3 jspl3_w_n6445_0(.douta(w_n6445_0[0]),.doutb(w_n6445_0[1]),.doutc(w_n6445_0[2]),.din(n6445));
	jspl3 jspl3_w_n6447_0(.douta(w_n6447_0[0]),.doutb(w_n6447_0[1]),.doutc(w_n6447_0[2]),.din(n6447));
	jspl jspl_w_n6448_0(.douta(w_n6448_0[0]),.doutb(w_n6448_0[1]),.din(n6448));
	jspl3 jspl3_w_n6452_0(.douta(w_n6452_0[0]),.doutb(w_n6452_0[1]),.doutc(w_n6452_0[2]),.din(n6452));
	jspl3 jspl3_w_n6455_0(.douta(w_n6455_0[0]),.doutb(w_n6455_0[1]),.doutc(w_n6455_0[2]),.din(n6455));
	jspl jspl_w_n6456_0(.douta(w_n6456_0[0]),.doutb(w_n6456_0[1]),.din(n6456));
	jspl3 jspl3_w_n6460_0(.douta(w_n6460_0[0]),.doutb(w_n6460_0[1]),.doutc(w_n6460_0[2]),.din(n6460));
	jspl3 jspl3_w_n6463_0(.douta(w_n6463_0[0]),.doutb(w_n6463_0[1]),.doutc(w_n6463_0[2]),.din(n6463));
	jspl jspl_w_n6464_0(.douta(w_n6464_0[0]),.doutb(w_n6464_0[1]),.din(n6464));
	jspl3 jspl3_w_n6468_0(.douta(w_n6468_0[0]),.doutb(w_n6468_0[1]),.doutc(w_n6468_0[2]),.din(n6468));
	jspl3 jspl3_w_n6471_0(.douta(w_n6471_0[0]),.doutb(w_n6471_0[1]),.doutc(w_n6471_0[2]),.din(n6471));
	jspl jspl_w_n6472_0(.douta(w_n6472_0[0]),.doutb(w_n6472_0[1]),.din(n6472));
	jspl3 jspl3_w_n6476_0(.douta(w_n6476_0[0]),.doutb(w_n6476_0[1]),.doutc(w_n6476_0[2]),.din(n6476));
	jspl3 jspl3_w_n6478_0(.douta(w_n6478_0[0]),.doutb(w_n6478_0[1]),.doutc(w_n6478_0[2]),.din(n6478));
	jspl jspl_w_n6479_0(.douta(w_n6479_0[0]),.doutb(w_n6479_0[1]),.din(n6479));
	jspl3 jspl3_w_n6483_0(.douta(w_n6483_0[0]),.doutb(w_n6483_0[1]),.doutc(w_n6483_0[2]),.din(n6483));
	jspl3 jspl3_w_n6485_0(.douta(w_n6485_0[0]),.doutb(w_n6485_0[1]),.doutc(w_n6485_0[2]),.din(n6485));
	jspl jspl_w_n6486_0(.douta(w_n6486_0[0]),.doutb(w_n6486_0[1]),.din(n6486));
	jspl3 jspl3_w_n6490_0(.douta(w_n6490_0[0]),.doutb(w_n6490_0[1]),.doutc(w_n6490_0[2]),.din(n6490));
	jspl3 jspl3_w_n6492_0(.douta(w_n6492_0[0]),.doutb(w_n6492_0[1]),.doutc(w_n6492_0[2]),.din(n6492));
	jspl jspl_w_n6493_0(.douta(w_n6493_0[0]),.doutb(w_n6493_0[1]),.din(n6493));
	jspl3 jspl3_w_n6497_0(.douta(w_n6497_0[0]),.doutb(w_n6497_0[1]),.doutc(w_n6497_0[2]),.din(n6497));
	jspl3 jspl3_w_n6500_0(.douta(w_n6500_0[0]),.doutb(w_n6500_0[1]),.doutc(w_n6500_0[2]),.din(n6500));
	jspl jspl_w_n6501_0(.douta(w_n6501_0[0]),.doutb(w_n6501_0[1]),.din(n6501));
	jspl3 jspl3_w_n6505_0(.douta(w_n6505_0[0]),.doutb(w_n6505_0[1]),.doutc(w_n6505_0[2]),.din(n6505));
	jspl3 jspl3_w_n6507_0(.douta(w_n6507_0[0]),.doutb(w_n6507_0[1]),.doutc(w_n6507_0[2]),.din(n6507));
	jspl jspl_w_n6508_0(.douta(w_n6508_0[0]),.doutb(w_n6508_0[1]),.din(n6508));
	jspl3 jspl3_w_n6512_0(.douta(w_n6512_0[0]),.doutb(w_n6512_0[1]),.doutc(w_n6512_0[2]),.din(n6512));
	jspl3 jspl3_w_n6515_0(.douta(w_n6515_0[0]),.doutb(w_n6515_0[1]),.doutc(w_n6515_0[2]),.din(n6515));
	jspl jspl_w_n6516_0(.douta(w_n6516_0[0]),.doutb(w_n6516_0[1]),.din(n6516));
	jspl3 jspl3_w_n6520_0(.douta(w_n6520_0[0]),.doutb(w_n6520_0[1]),.doutc(w_n6520_0[2]),.din(n6520));
	jspl3 jspl3_w_n6522_0(.douta(w_n6522_0[0]),.doutb(w_n6522_0[1]),.doutc(w_n6522_0[2]),.din(n6522));
	jspl jspl_w_n6523_0(.douta(w_n6523_0[0]),.doutb(w_n6523_0[1]),.din(n6523));
	jspl3 jspl3_w_n6527_0(.douta(w_n6527_0[0]),.doutb(w_n6527_0[1]),.doutc(w_n6527_0[2]),.din(n6527));
	jspl3 jspl3_w_n6530_0(.douta(w_n6530_0[0]),.doutb(w_n6530_0[1]),.doutc(w_n6530_0[2]),.din(n6530));
	jspl jspl_w_n6531_0(.douta(w_n6531_0[0]),.doutb(w_n6531_0[1]),.din(n6531));
	jspl3 jspl3_w_n6535_0(.douta(w_n6535_0[0]),.doutb(w_n6535_0[1]),.doutc(w_n6535_0[2]),.din(n6535));
	jspl3 jspl3_w_n6538_0(.douta(w_n6538_0[0]),.doutb(w_n6538_0[1]),.doutc(w_n6538_0[2]),.din(n6538));
	jspl jspl_w_n6539_0(.douta(w_n6539_0[0]),.doutb(w_n6539_0[1]),.din(n6539));
	jspl3 jspl3_w_n6543_0(.douta(w_n6543_0[0]),.doutb(w_n6543_0[1]),.doutc(w_n6543_0[2]),.din(n6543));
	jspl3 jspl3_w_n6545_0(.douta(w_n6545_0[0]),.doutb(w_n6545_0[1]),.doutc(w_n6545_0[2]),.din(n6545));
	jspl jspl_w_n6546_0(.douta(w_n6546_0[0]),.doutb(w_n6546_0[1]),.din(n6546));
	jspl3 jspl3_w_n6550_0(.douta(w_n6550_0[0]),.doutb(w_n6550_0[1]),.doutc(w_n6550_0[2]),.din(n6550));
	jspl3 jspl3_w_n6552_0(.douta(w_n6552_0[0]),.doutb(w_n6552_0[1]),.doutc(w_n6552_0[2]),.din(n6552));
	jspl jspl_w_n6553_0(.douta(w_n6553_0[0]),.doutb(w_n6553_0[1]),.din(n6553));
	jspl jspl_w_n6557_0(.douta(w_n6557_0[0]),.doutb(w_n6557_0[1]),.din(n6557));
	jspl jspl_w_n6558_0(.douta(w_n6558_0[0]),.doutb(w_n6558_0[1]),.din(n6558));
	jspl3 jspl3_w_n6560_0(.douta(w_n6560_0[0]),.doutb(w_n6560_0[1]),.doutc(w_n6560_0[2]),.din(n6560));
	jspl jspl_w_n6561_0(.douta(w_n6561_0[0]),.doutb(w_n6561_0[1]),.din(n6561));
	jspl3 jspl3_w_n6565_0(.douta(w_n6565_0[0]),.doutb(w_n6565_0[1]),.doutc(w_n6565_0[2]),.din(n6565));
	jspl3 jspl3_w_n6568_0(.douta(w_n6568_0[0]),.doutb(w_n6568_0[1]),.doutc(w_n6568_0[2]),.din(n6568));
	jspl jspl_w_n6569_0(.douta(w_n6569_0[0]),.doutb(w_n6569_0[1]),.din(n6569));
	jspl3 jspl3_w_n6573_0(.douta(w_n6573_0[0]),.doutb(w_n6573_0[1]),.doutc(w_n6573_0[2]),.din(n6573));
	jspl3 jspl3_w_n6576_0(.douta(w_n6576_0[0]),.doutb(w_n6576_0[1]),.doutc(w_n6576_0[2]),.din(n6576));
	jspl jspl_w_n6577_0(.douta(w_n6577_0[0]),.doutb(w_n6577_0[1]),.din(n6577));
	jspl3 jspl3_w_n6581_0(.douta(w_n6581_0[0]),.doutb(w_n6581_0[1]),.doutc(w_n6581_0[2]),.din(n6581));
	jspl3 jspl3_w_n6583_0(.douta(w_n6583_0[0]),.doutb(w_n6583_0[1]),.doutc(w_n6583_0[2]),.din(n6583));
	jspl jspl_w_n6584_0(.douta(w_n6584_0[0]),.doutb(w_n6584_0[1]),.din(n6584));
	jspl3 jspl3_w_n6588_0(.douta(w_n6588_0[0]),.doutb(w_n6588_0[1]),.doutc(w_n6588_0[2]),.din(n6588));
	jspl3 jspl3_w_n6590_0(.douta(w_n6590_0[0]),.doutb(w_n6590_0[1]),.doutc(w_n6590_0[2]),.din(n6590));
	jspl jspl_w_n6591_0(.douta(w_n6591_0[0]),.doutb(w_n6591_0[1]),.din(n6591));
	jspl3 jspl3_w_n6596_0(.douta(w_n6596_0[0]),.doutb(w_n6596_0[1]),.doutc(w_n6596_0[2]),.din(n6596));
	jspl jspl_w_n6601_0(.douta(w_n6601_0[0]),.doutb(w_n6601_0[1]),.din(n6601));
	jspl jspl_w_n6604_0(.douta(w_n6604_0[0]),.doutb(w_n6604_0[1]),.din(n6604));
	jspl3 jspl3_w_n6606_0(.douta(w_n6606_0[0]),.doutb(w_n6606_0[1]),.doutc(w_n6606_0[2]),.din(n6606));
	jspl3 jspl3_w_n6606_1(.douta(w_n6606_1[0]),.doutb(w_n6606_1[1]),.doutc(w_n6606_1[2]),.din(w_n6606_0[0]));
	jspl jspl_w_n6607_0(.douta(w_n6607_0[0]),.doutb(w_n6607_0[1]),.din(n6607));
	jspl3 jspl3_w_n6608_0(.douta(w_n6608_0[0]),.doutb(w_n6608_0[1]),.doutc(w_n6608_0[2]),.din(n6608));
	jspl jspl_w_n6609_0(.douta(w_n6609_0[0]),.doutb(w_n6609_0[1]),.din(n6609));
	jspl3 jspl3_w_n6611_0(.douta(w_n6611_0[0]),.doutb(w_n6611_0[1]),.doutc(w_n6611_0[2]),.din(n6611));
	jspl jspl_w_n6612_0(.douta(w_n6612_0[0]),.doutb(w_n6612_0[1]),.din(n6612));
	jspl jspl_w_n6652_0(.douta(w_n6652_0[0]),.doutb(w_n6652_0[1]),.din(n6652));
	jspl jspl_w_n6656_0(.douta(w_n6656_0[0]),.doutb(w_n6656_0[1]),.din(n6656));
	jspl jspl_w_n6753_0(.douta(w_n6753_0[0]),.doutb(w_n6753_0[1]),.din(n6753));
	jspl jspl_w_n6756_0(.douta(w_n6756_0[0]),.doutb(w_n6756_0[1]),.din(n6756));
	jspl3 jspl3_w_n6758_0(.douta(w_n6758_0[0]),.doutb(w_n6758_0[1]),.doutc(w_n6758_0[2]),.din(n6758));
	jspl3 jspl3_w_n6758_1(.douta(w_n6758_1[0]),.doutb(w_n6758_1[1]),.doutc(w_n6758_1[2]),.din(w_n6758_0[0]));
	jspl3 jspl3_w_n6758_2(.douta(w_n6758_2[0]),.doutb(w_n6758_2[1]),.doutc(w_n6758_2[2]),.din(w_n6758_0[1]));
	jspl3 jspl3_w_n6758_3(.douta(w_n6758_3[0]),.doutb(w_n6758_3[1]),.doutc(w_n6758_3[2]),.din(w_n6758_0[2]));
	jspl3 jspl3_w_n6758_4(.douta(w_n6758_4[0]),.doutb(w_n6758_4[1]),.doutc(w_n6758_4[2]),.din(w_n6758_1[0]));
	jspl3 jspl3_w_n6758_5(.douta(w_n6758_5[0]),.doutb(w_n6758_5[1]),.doutc(w_n6758_5[2]),.din(w_n6758_1[1]));
	jspl3 jspl3_w_n6758_6(.douta(w_n6758_6[0]),.doutb(w_n6758_6[1]),.doutc(w_n6758_6[2]),.din(w_n6758_1[2]));
	jspl3 jspl3_w_n6758_7(.douta(w_n6758_7[0]),.doutb(w_n6758_7[1]),.doutc(w_n6758_7[2]),.din(w_n6758_2[0]));
	jspl3 jspl3_w_n6758_8(.douta(w_n6758_8[0]),.doutb(w_n6758_8[1]),.doutc(w_n6758_8[2]),.din(w_n6758_2[1]));
	jspl3 jspl3_w_n6758_9(.douta(w_n6758_9[0]),.doutb(w_n6758_9[1]),.doutc(w_n6758_9[2]),.din(w_n6758_2[2]));
	jspl3 jspl3_w_n6758_10(.douta(w_n6758_10[0]),.doutb(w_n6758_10[1]),.doutc(w_n6758_10[2]),.din(w_n6758_3[0]));
	jspl3 jspl3_w_n6758_11(.douta(w_n6758_11[0]),.doutb(w_n6758_11[1]),.doutc(w_n6758_11[2]),.din(w_n6758_3[1]));
	jspl3 jspl3_w_n6758_12(.douta(w_n6758_12[0]),.doutb(w_n6758_12[1]),.doutc(w_n6758_12[2]),.din(w_n6758_3[2]));
	jspl3 jspl3_w_n6758_13(.douta(w_n6758_13[0]),.doutb(w_n6758_13[1]),.doutc(w_n6758_13[2]),.din(w_n6758_4[0]));
	jspl3 jspl3_w_n6758_14(.douta(w_n6758_14[0]),.doutb(w_n6758_14[1]),.doutc(w_n6758_14[2]),.din(w_n6758_4[1]));
	jspl3 jspl3_w_n6758_15(.douta(w_n6758_15[0]),.doutb(w_n6758_15[1]),.doutc(w_n6758_15[2]),.din(w_n6758_4[2]));
	jspl3 jspl3_w_n6758_16(.douta(w_n6758_16[0]),.doutb(w_n6758_16[1]),.doutc(w_n6758_16[2]),.din(w_n6758_5[0]));
	jspl3 jspl3_w_n6758_17(.douta(w_n6758_17[0]),.doutb(w_n6758_17[1]),.doutc(w_n6758_17[2]),.din(w_n6758_5[1]));
	jspl3 jspl3_w_n6758_18(.douta(w_n6758_18[0]),.doutb(w_n6758_18[1]),.doutc(w_n6758_18[2]),.din(w_n6758_5[2]));
	jspl3 jspl3_w_n6758_19(.douta(w_n6758_19[0]),.doutb(w_n6758_19[1]),.doutc(w_n6758_19[2]),.din(w_n6758_6[0]));
	jspl3 jspl3_w_n6758_20(.douta(w_n6758_20[0]),.doutb(w_n6758_20[1]),.doutc(w_n6758_20[2]),.din(w_n6758_6[1]));
	jspl3 jspl3_w_n6758_21(.douta(w_n6758_21[0]),.doutb(w_n6758_21[1]),.doutc(w_n6758_21[2]),.din(w_n6758_6[2]));
	jspl3 jspl3_w_n6758_22(.douta(w_n6758_22[0]),.doutb(w_n6758_22[1]),.doutc(w_n6758_22[2]),.din(w_n6758_7[0]));
	jspl3 jspl3_w_n6758_23(.douta(w_n6758_23[0]),.doutb(w_n6758_23[1]),.doutc(w_n6758_23[2]),.din(w_n6758_7[1]));
	jspl3 jspl3_w_n6758_24(.douta(w_n6758_24[0]),.doutb(w_n6758_24[1]),.doutc(w_n6758_24[2]),.din(w_n6758_7[2]));
	jspl3 jspl3_w_n6758_25(.douta(w_n6758_25[0]),.doutb(w_n6758_25[1]),.doutc(w_n6758_25[2]),.din(w_n6758_8[0]));
	jspl3 jspl3_w_n6758_26(.douta(w_n6758_26[0]),.doutb(w_n6758_26[1]),.doutc(w_n6758_26[2]),.din(w_n6758_8[1]));
	jspl3 jspl3_w_n6758_27(.douta(w_n6758_27[0]),.doutb(w_n6758_27[1]),.doutc(w_n6758_27[2]),.din(w_n6758_8[2]));
	jspl3 jspl3_w_n6758_28(.douta(w_n6758_28[0]),.doutb(w_n6758_28[1]),.doutc(w_n6758_28[2]),.din(w_n6758_9[0]));
	jspl3 jspl3_w_n6758_29(.douta(w_n6758_29[0]),.doutb(w_n6758_29[1]),.doutc(w_n6758_29[2]),.din(w_n6758_9[1]));
	jspl3 jspl3_w_n6758_30(.douta(w_n6758_30[0]),.doutb(w_n6758_30[1]),.doutc(w_n6758_30[2]),.din(w_n6758_9[2]));
	jspl3 jspl3_w_n6758_31(.douta(w_n6758_31[0]),.doutb(w_n6758_31[1]),.doutc(w_n6758_31[2]),.din(w_n6758_10[0]));
	jspl3 jspl3_w_n6758_32(.douta(w_n6758_32[0]),.doutb(w_n6758_32[1]),.doutc(w_n6758_32[2]),.din(w_n6758_10[1]));
	jspl3 jspl3_w_n6758_33(.douta(w_n6758_33[0]),.doutb(w_n6758_33[1]),.doutc(w_n6758_33[2]),.din(w_n6758_10[2]));
	jspl3 jspl3_w_n6758_34(.douta(w_n6758_34[0]),.doutb(w_n6758_34[1]),.doutc(w_n6758_34[2]),.din(w_n6758_11[0]));
	jspl3 jspl3_w_n6758_35(.douta(w_n6758_35[0]),.doutb(w_n6758_35[1]),.doutc(w_n6758_35[2]),.din(w_n6758_11[1]));
	jspl3 jspl3_w_n6758_36(.douta(w_n6758_36[0]),.doutb(w_n6758_36[1]),.doutc(w_n6758_36[2]),.din(w_n6758_11[2]));
	jspl3 jspl3_w_n6758_37(.douta(w_n6758_37[0]),.doutb(w_n6758_37[1]),.doutc(w_n6758_37[2]),.din(w_n6758_12[0]));
	jspl3 jspl3_w_n6758_38(.douta(w_n6758_38[0]),.doutb(w_n6758_38[1]),.doutc(w_n6758_38[2]),.din(w_n6758_12[1]));
	jspl3 jspl3_w_n6758_39(.douta(w_n6758_39[0]),.doutb(w_n6758_39[1]),.doutc(w_n6758_39[2]),.din(w_n6758_12[2]));
	jspl3 jspl3_w_n6758_40(.douta(w_n6758_40[0]),.doutb(w_n6758_40[1]),.doutc(w_n6758_40[2]),.din(w_n6758_13[0]));
	jspl3 jspl3_w_n6762_0(.douta(w_n6762_0[0]),.doutb(w_n6762_0[1]),.doutc(w_n6762_0[2]),.din(n6762));
	jspl jspl_w_n6763_0(.douta(w_n6763_0[0]),.doutb(w_n6763_0[1]),.din(n6763));
	jspl jspl_w_n6765_0(.douta(w_n6765_0[0]),.doutb(w_n6765_0[1]),.din(n6765));
	jspl jspl_w_n6766_0(.douta(w_n6766_0[0]),.doutb(w_n6766_0[1]),.din(n6766));
	jspl jspl_w_n6771_0(.douta(w_n6771_0[0]),.doutb(w_n6771_0[1]),.din(n6771));
	jspl jspl_w_n6772_0(.douta(w_n6772_0[0]),.doutb(w_n6772_0[1]),.din(n6772));
	jspl3 jspl3_w_n6774_0(.douta(w_n6774_0[0]),.doutb(w_n6774_0[1]),.doutc(w_n6774_0[2]),.din(n6774));
	jspl jspl_w_n6775_0(.douta(w_n6775_0[0]),.doutb(w_n6775_0[1]),.din(n6775));
	jspl jspl_w_n6779_0(.douta(w_n6779_0[0]),.doutb(w_n6779_0[1]),.din(n6779));
	jspl3 jspl3_w_n6781_0(.douta(w_n6781_0[0]),.doutb(w_n6781_0[1]),.doutc(w_n6781_0[2]),.din(n6781));
	jspl jspl_w_n6782_0(.douta(w_n6782_0[0]),.doutb(w_n6782_0[1]),.din(n6782));
	jspl jspl_w_n6786_0(.douta(w_n6786_0[0]),.doutb(w_n6786_0[1]),.din(n6786));
	jspl3 jspl3_w_n6788_0(.douta(w_n6788_0[0]),.doutb(w_n6788_0[1]),.doutc(w_n6788_0[2]),.din(n6788));
	jspl jspl_w_n6789_0(.douta(w_n6789_0[0]),.doutb(w_n6789_0[1]),.din(n6789));
	jspl jspl_w_n6793_0(.douta(w_n6793_0[0]),.doutb(w_n6793_0[1]),.din(n6793));
	jspl3 jspl3_w_n6795_0(.douta(w_n6795_0[0]),.doutb(w_n6795_0[1]),.doutc(w_n6795_0[2]),.din(n6795));
	jspl jspl_w_n6796_0(.douta(w_n6796_0[0]),.doutb(w_n6796_0[1]),.din(n6796));
	jspl jspl_w_n6800_0(.douta(w_n6800_0[0]),.doutb(w_n6800_0[1]),.din(n6800));
	jspl jspl_w_n6801_0(.douta(w_n6801_0[0]),.doutb(w_n6801_0[1]),.din(n6801));
	jspl3 jspl3_w_n6803_0(.douta(w_n6803_0[0]),.doutb(w_n6803_0[1]),.doutc(w_n6803_0[2]),.din(n6803));
	jspl jspl_w_n6804_0(.douta(w_n6804_0[0]),.doutb(w_n6804_0[1]),.din(n6804));
	jspl jspl_w_n6808_0(.douta(w_n6808_0[0]),.doutb(w_n6808_0[1]),.din(n6808));
	jspl3 jspl3_w_n6810_0(.douta(w_n6810_0[0]),.doutb(w_n6810_0[1]),.doutc(w_n6810_0[2]),.din(n6810));
	jspl jspl_w_n6811_0(.douta(w_n6811_0[0]),.doutb(w_n6811_0[1]),.din(n6811));
	jspl jspl_w_n6815_0(.douta(w_n6815_0[0]),.doutb(w_n6815_0[1]),.din(n6815));
	jspl jspl_w_n6816_0(.douta(w_n6816_0[0]),.doutb(w_n6816_0[1]),.din(n6816));
	jspl3 jspl3_w_n6818_0(.douta(w_n6818_0[0]),.doutb(w_n6818_0[1]),.doutc(w_n6818_0[2]),.din(n6818));
	jspl jspl_w_n6819_0(.douta(w_n6819_0[0]),.doutb(w_n6819_0[1]),.din(n6819));
	jspl jspl_w_n6823_0(.douta(w_n6823_0[0]),.doutb(w_n6823_0[1]),.din(n6823));
	jspl3 jspl3_w_n6825_0(.douta(w_n6825_0[0]),.doutb(w_n6825_0[1]),.doutc(w_n6825_0[2]),.din(n6825));
	jspl jspl_w_n6826_0(.douta(w_n6826_0[0]),.doutb(w_n6826_0[1]),.din(n6826));
	jspl jspl_w_n6830_0(.douta(w_n6830_0[0]),.doutb(w_n6830_0[1]),.din(n6830));
	jspl jspl_w_n6831_0(.douta(w_n6831_0[0]),.doutb(w_n6831_0[1]),.din(n6831));
	jspl3 jspl3_w_n6833_0(.douta(w_n6833_0[0]),.doutb(w_n6833_0[1]),.doutc(w_n6833_0[2]),.din(n6833));
	jspl jspl_w_n6834_0(.douta(w_n6834_0[0]),.doutb(w_n6834_0[1]),.din(n6834));
	jspl jspl_w_n6838_0(.douta(w_n6838_0[0]),.doutb(w_n6838_0[1]),.din(n6838));
	jspl3 jspl3_w_n6840_0(.douta(w_n6840_0[0]),.doutb(w_n6840_0[1]),.doutc(w_n6840_0[2]),.din(n6840));
	jspl jspl_w_n6841_0(.douta(w_n6841_0[0]),.doutb(w_n6841_0[1]),.din(n6841));
	jspl jspl_w_n6845_0(.douta(w_n6845_0[0]),.doutb(w_n6845_0[1]),.din(n6845));
	jspl jspl_w_n6846_0(.douta(w_n6846_0[0]),.doutb(w_n6846_0[1]),.din(n6846));
	jspl3 jspl3_w_n6848_0(.douta(w_n6848_0[0]),.doutb(w_n6848_0[1]),.doutc(w_n6848_0[2]),.din(n6848));
	jspl jspl_w_n6849_0(.douta(w_n6849_0[0]),.doutb(w_n6849_0[1]),.din(n6849));
	jspl jspl_w_n6853_0(.douta(w_n6853_0[0]),.doutb(w_n6853_0[1]),.din(n6853));
	jspl3 jspl3_w_n6855_0(.douta(w_n6855_0[0]),.doutb(w_n6855_0[1]),.doutc(w_n6855_0[2]),.din(n6855));
	jspl jspl_w_n6856_0(.douta(w_n6856_0[0]),.doutb(w_n6856_0[1]),.din(n6856));
	jspl jspl_w_n6860_0(.douta(w_n6860_0[0]),.doutb(w_n6860_0[1]),.din(n6860));
	jspl3 jspl3_w_n6862_0(.douta(w_n6862_0[0]),.doutb(w_n6862_0[1]),.doutc(w_n6862_0[2]),.din(n6862));
	jspl jspl_w_n6863_0(.douta(w_n6863_0[0]),.doutb(w_n6863_0[1]),.din(n6863));
	jspl jspl_w_n6867_0(.douta(w_n6867_0[0]),.doutb(w_n6867_0[1]),.din(n6867));
	jspl3 jspl3_w_n6869_0(.douta(w_n6869_0[0]),.doutb(w_n6869_0[1]),.doutc(w_n6869_0[2]),.din(n6869));
	jspl jspl_w_n6870_0(.douta(w_n6870_0[0]),.doutb(w_n6870_0[1]),.din(n6870));
	jspl jspl_w_n6874_0(.douta(w_n6874_0[0]),.doutb(w_n6874_0[1]),.din(n6874));
	jspl jspl_w_n6875_0(.douta(w_n6875_0[0]),.doutb(w_n6875_0[1]),.din(n6875));
	jspl3 jspl3_w_n6877_0(.douta(w_n6877_0[0]),.doutb(w_n6877_0[1]),.doutc(w_n6877_0[2]),.din(n6877));
	jspl jspl_w_n6878_0(.douta(w_n6878_0[0]),.doutb(w_n6878_0[1]),.din(n6878));
	jspl jspl_w_n6882_0(.douta(w_n6882_0[0]),.doutb(w_n6882_0[1]),.din(n6882));
	jspl jspl_w_n6883_0(.douta(w_n6883_0[0]),.doutb(w_n6883_0[1]),.din(n6883));
	jspl3 jspl3_w_n6885_0(.douta(w_n6885_0[0]),.doutb(w_n6885_0[1]),.doutc(w_n6885_0[2]),.din(n6885));
	jspl jspl_w_n6886_0(.douta(w_n6886_0[0]),.doutb(w_n6886_0[1]),.din(n6886));
	jspl jspl_w_n6890_0(.douta(w_n6890_0[0]),.doutb(w_n6890_0[1]),.din(n6890));
	jspl jspl_w_n6891_0(.douta(w_n6891_0[0]),.doutb(w_n6891_0[1]),.din(n6891));
	jspl3 jspl3_w_n6893_0(.douta(w_n6893_0[0]),.doutb(w_n6893_0[1]),.doutc(w_n6893_0[2]),.din(n6893));
	jspl jspl_w_n6894_0(.douta(w_n6894_0[0]),.doutb(w_n6894_0[1]),.din(n6894));
	jspl jspl_w_n6898_0(.douta(w_n6898_0[0]),.doutb(w_n6898_0[1]),.din(n6898));
	jspl3 jspl3_w_n6900_0(.douta(w_n6900_0[0]),.doutb(w_n6900_0[1]),.doutc(w_n6900_0[2]),.din(n6900));
	jspl jspl_w_n6901_0(.douta(w_n6901_0[0]),.doutb(w_n6901_0[1]),.din(n6901));
	jspl jspl_w_n6905_0(.douta(w_n6905_0[0]),.doutb(w_n6905_0[1]),.din(n6905));
	jspl jspl_w_n6906_0(.douta(w_n6906_0[0]),.doutb(w_n6906_0[1]),.din(n6906));
	jspl3 jspl3_w_n6908_0(.douta(w_n6908_0[0]),.doutb(w_n6908_0[1]),.doutc(w_n6908_0[2]),.din(n6908));
	jspl jspl_w_n6909_0(.douta(w_n6909_0[0]),.doutb(w_n6909_0[1]),.din(n6909));
	jspl jspl_w_n6913_0(.douta(w_n6913_0[0]),.doutb(w_n6913_0[1]),.din(n6913));
	jspl3 jspl3_w_n6915_0(.douta(w_n6915_0[0]),.doutb(w_n6915_0[1]),.doutc(w_n6915_0[2]),.din(n6915));
	jspl jspl_w_n6916_0(.douta(w_n6916_0[0]),.doutb(w_n6916_0[1]),.din(n6916));
	jspl jspl_w_n6920_0(.douta(w_n6920_0[0]),.doutb(w_n6920_0[1]),.din(n6920));
	jspl jspl_w_n6921_0(.douta(w_n6921_0[0]),.doutb(w_n6921_0[1]),.din(n6921));
	jspl3 jspl3_w_n6923_0(.douta(w_n6923_0[0]),.doutb(w_n6923_0[1]),.doutc(w_n6923_0[2]),.din(n6923));
	jspl jspl_w_n6924_0(.douta(w_n6924_0[0]),.doutb(w_n6924_0[1]),.din(n6924));
	jspl jspl_w_n6928_0(.douta(w_n6928_0[0]),.doutb(w_n6928_0[1]),.din(n6928));
	jspl3 jspl3_w_n6930_0(.douta(w_n6930_0[0]),.doutb(w_n6930_0[1]),.doutc(w_n6930_0[2]),.din(n6930));
	jspl jspl_w_n6931_0(.douta(w_n6931_0[0]),.doutb(w_n6931_0[1]),.din(n6931));
	jspl jspl_w_n6935_0(.douta(w_n6935_0[0]),.doutb(w_n6935_0[1]),.din(n6935));
	jspl3 jspl3_w_n6937_0(.douta(w_n6937_0[0]),.doutb(w_n6937_0[1]),.doutc(w_n6937_0[2]),.din(n6937));
	jspl jspl_w_n6938_0(.douta(w_n6938_0[0]),.doutb(w_n6938_0[1]),.din(n6938));
	jspl jspl_w_n6942_0(.douta(w_n6942_0[0]),.doutb(w_n6942_0[1]),.din(n6942));
	jspl jspl_w_n6943_0(.douta(w_n6943_0[0]),.doutb(w_n6943_0[1]),.din(n6943));
	jspl3 jspl3_w_n6945_0(.douta(w_n6945_0[0]),.doutb(w_n6945_0[1]),.doutc(w_n6945_0[2]),.din(n6945));
	jspl jspl_w_n6946_0(.douta(w_n6946_0[0]),.doutb(w_n6946_0[1]),.din(n6946));
	jspl jspl_w_n6950_0(.douta(w_n6950_0[0]),.doutb(w_n6950_0[1]),.din(n6950));
	jspl jspl_w_n6951_0(.douta(w_n6951_0[0]),.doutb(w_n6951_0[1]),.din(n6951));
	jspl3 jspl3_w_n6953_0(.douta(w_n6953_0[0]),.doutb(w_n6953_0[1]),.doutc(w_n6953_0[2]),.din(n6953));
	jspl jspl_w_n6954_0(.douta(w_n6954_0[0]),.doutb(w_n6954_0[1]),.din(n6954));
	jspl jspl_w_n6958_0(.douta(w_n6958_0[0]),.doutb(w_n6958_0[1]),.din(n6958));
	jspl jspl_w_n6959_0(.douta(w_n6959_0[0]),.doutb(w_n6959_0[1]),.din(n6959));
	jspl3 jspl3_w_n6961_0(.douta(w_n6961_0[0]),.doutb(w_n6961_0[1]),.doutc(w_n6961_0[2]),.din(n6961));
	jspl jspl_w_n6962_0(.douta(w_n6962_0[0]),.doutb(w_n6962_0[1]),.din(n6962));
	jspl jspl_w_n6966_0(.douta(w_n6966_0[0]),.doutb(w_n6966_0[1]),.din(n6966));
	jspl3 jspl3_w_n6968_0(.douta(w_n6968_0[0]),.doutb(w_n6968_0[1]),.doutc(w_n6968_0[2]),.din(n6968));
	jspl jspl_w_n6969_0(.douta(w_n6969_0[0]),.doutb(w_n6969_0[1]),.din(n6969));
	jspl jspl_w_n6973_0(.douta(w_n6973_0[0]),.doutb(w_n6973_0[1]),.din(n6973));
	jspl3 jspl3_w_n6975_0(.douta(w_n6975_0[0]),.doutb(w_n6975_0[1]),.doutc(w_n6975_0[2]),.din(n6975));
	jspl jspl_w_n6976_0(.douta(w_n6976_0[0]),.doutb(w_n6976_0[1]),.din(n6976));
	jspl jspl_w_n6980_0(.douta(w_n6980_0[0]),.doutb(w_n6980_0[1]),.din(n6980));
	jspl jspl_w_n6981_0(.douta(w_n6981_0[0]),.doutb(w_n6981_0[1]),.din(n6981));
	jspl jspl_w_n6983_0(.douta(w_n6983_0[0]),.doutb(w_n6983_0[1]),.din(n6983));
	jspl3 jspl3_w_n6986_0(.douta(w_n6986_0[0]),.doutb(w_n6986_0[1]),.doutc(w_n6986_0[2]),.din(n6986));
	jspl jspl_w_n6987_0(.douta(w_n6987_0[0]),.doutb(w_n6987_0[1]),.din(n6987));
	jspl3 jspl3_w_n6988_0(.douta(w_n6988_0[0]),.doutb(w_n6988_0[1]),.doutc(w_n6988_0[2]),.din(n6988));
	jspl jspl_w_n6988_1(.douta(w_n6988_1[0]),.doutb(w_n6988_1[1]),.din(w_n6988_0[0]));
	jspl3 jspl3_w_n6989_0(.douta(w_n6989_0[0]),.doutb(w_n6989_0[1]),.doutc(w_n6989_0[2]),.din(n6989));
	jspl jspl_w_n6993_0(.douta(w_n6993_0[0]),.doutb(w_n6993_0[1]),.din(n6993));
	jspl jspl_w_n6994_0(.douta(w_n6994_0[0]),.doutb(w_n6994_0[1]),.din(n6994));
	jspl jspl_w_n7031_0(.douta(w_n7031_0[0]),.doutb(w_n7031_0[1]),.din(n7031));
	jspl jspl_w_n7038_0(.douta(w_n7038_0[0]),.doutb(w_n7038_0[1]),.din(n7038));
	jspl jspl_w_n7042_0(.douta(w_n7042_0[0]),.doutb(w_n7042_0[1]),.din(n7042));
	jspl jspl_w_n7046_0(.douta(w_n7046_0[0]),.doutb(w_n7046_0[1]),.din(n7046));
	jspl jspl_w_n7053_0(.douta(w_n7053_0[0]),.doutb(w_n7053_0[1]),.din(n7053));
	jspl jspl_w_n7060_0(.douta(w_n7060_0[0]),.doutb(w_n7060_0[1]),.din(n7060));
	jspl jspl_w_n7067_0(.douta(w_n7067_0[0]),.doutb(w_n7067_0[1]),.din(n7067));
	jspl jspl_w_n7074_0(.douta(w_n7074_0[0]),.doutb(w_n7074_0[1]),.din(n7074));
	jspl jspl_w_n7078_0(.douta(w_n7078_0[0]),.doutb(w_n7078_0[1]),.din(n7078));
	jspl jspl_w_n7082_0(.douta(w_n7082_0[0]),.doutb(w_n7082_0[1]),.din(n7082));
	jspl jspl_w_n7095_0(.douta(w_n7095_0[0]),.doutb(w_n7095_0[1]),.din(n7095));
	jspl jspl_w_n7102_0(.douta(w_n7102_0[0]),.doutb(w_n7102_0[1]),.din(n7102));
	jspl jspl_w_n7109_0(.douta(w_n7109_0[0]),.doutb(w_n7109_0[1]),.din(n7109));
	jspl jspl_w_n7113_0(.douta(w_n7113_0[0]),.doutb(w_n7113_0[1]),.din(n7113));
	jspl jspl_w_n7126_0(.douta(w_n7126_0[0]),.doutb(w_n7126_0[1]),.din(n7126));
	jspl jspl_w_n7130_0(.douta(w_n7130_0[0]),.doutb(w_n7130_0[1]),.din(n7130));
	jspl jspl_w_n7135_0(.douta(w_n7135_0[0]),.doutb(w_n7135_0[1]),.din(n7135));
	jspl jspl_w_n7136_0(.douta(w_n7136_0[0]),.doutb(w_n7136_0[1]),.din(n7136));
	jspl jspl_w_n7138_0(.douta(w_n7138_0[0]),.doutb(w_n7138_0[1]),.din(n7138));
	jspl jspl_w_n7140_0(.douta(w_n7140_0[0]),.doutb(w_n7140_0[1]),.din(n7140));
	jspl jspl_w_n7141_0(.douta(w_n7141_0[0]),.doutb(w_n7141_0[1]),.din(n7141));
	jspl jspl_w_n7143_0(.douta(w_n7143_0[0]),.doutb(w_n7143_0[1]),.din(n7143));
	jspl jspl_w_n7145_0(.douta(w_n7145_0[0]),.doutb(w_n7145_0[1]),.din(n7145));
	jspl jspl_w_n7146_0(.douta(w_n7146_0[0]),.doutb(w_n7146_0[1]),.din(n7146));
	jspl jspl_w_n7153_0(.douta(w_n7153_0[0]),.doutb(w_n7153_0[1]),.din(n7153));
	jspl3 jspl3_w_n7154_0(.douta(w_n7154_0[0]),.doutb(w_n7154_0[1]),.doutc(w_n7154_0[2]),.din(n7154));
	jspl3 jspl3_w_n7154_1(.douta(w_n7154_1[0]),.doutb(w_n7154_1[1]),.doutc(w_n7154_1[2]),.din(w_n7154_0[0]));
	jspl3 jspl3_w_n7154_2(.douta(w_n7154_2[0]),.doutb(w_n7154_2[1]),.doutc(w_n7154_2[2]),.din(w_n7154_0[1]));
	jspl3 jspl3_w_n7154_3(.douta(w_n7154_3[0]),.doutb(w_n7154_3[1]),.doutc(w_n7154_3[2]),.din(w_n7154_0[2]));
	jspl3 jspl3_w_n7154_4(.douta(w_n7154_4[0]),.doutb(w_n7154_4[1]),.doutc(w_n7154_4[2]),.din(w_n7154_1[0]));
	jspl3 jspl3_w_n7154_5(.douta(w_n7154_5[0]),.doutb(w_n7154_5[1]),.doutc(w_n7154_5[2]),.din(w_n7154_1[1]));
	jspl3 jspl3_w_n7154_6(.douta(w_n7154_6[0]),.doutb(w_n7154_6[1]),.doutc(w_n7154_6[2]),.din(w_n7154_1[2]));
	jspl3 jspl3_w_n7154_7(.douta(w_n7154_7[0]),.doutb(w_n7154_7[1]),.doutc(w_n7154_7[2]),.din(w_n7154_2[0]));
	jspl3 jspl3_w_n7154_8(.douta(w_n7154_8[0]),.doutb(w_n7154_8[1]),.doutc(w_n7154_8[2]),.din(w_n7154_2[1]));
	jspl3 jspl3_w_n7154_9(.douta(w_n7154_9[0]),.doutb(w_n7154_9[1]),.doutc(w_n7154_9[2]),.din(w_n7154_2[2]));
	jspl3 jspl3_w_n7154_10(.douta(w_n7154_10[0]),.doutb(w_n7154_10[1]),.doutc(w_n7154_10[2]),.din(w_n7154_3[0]));
	jspl3 jspl3_w_n7154_11(.douta(w_n7154_11[0]),.doutb(w_n7154_11[1]),.doutc(w_n7154_11[2]),.din(w_n7154_3[1]));
	jspl3 jspl3_w_n7154_12(.douta(w_n7154_12[0]),.doutb(w_n7154_12[1]),.doutc(w_n7154_12[2]),.din(w_n7154_3[2]));
	jspl3 jspl3_w_n7154_13(.douta(w_n7154_13[0]),.doutb(w_n7154_13[1]),.doutc(w_n7154_13[2]),.din(w_n7154_4[0]));
	jspl3 jspl3_w_n7154_14(.douta(w_n7154_14[0]),.doutb(w_n7154_14[1]),.doutc(w_n7154_14[2]),.din(w_n7154_4[1]));
	jspl3 jspl3_w_n7154_15(.douta(w_n7154_15[0]),.doutb(w_n7154_15[1]),.doutc(w_n7154_15[2]),.din(w_n7154_4[2]));
	jspl3 jspl3_w_n7154_16(.douta(w_n7154_16[0]),.doutb(w_n7154_16[1]),.doutc(w_n7154_16[2]),.din(w_n7154_5[0]));
	jspl3 jspl3_w_n7154_17(.douta(w_n7154_17[0]),.doutb(w_n7154_17[1]),.doutc(w_n7154_17[2]),.din(w_n7154_5[1]));
	jspl3 jspl3_w_n7154_18(.douta(w_n7154_18[0]),.doutb(w_n7154_18[1]),.doutc(w_n7154_18[2]),.din(w_n7154_5[2]));
	jspl3 jspl3_w_n7154_19(.douta(w_n7154_19[0]),.doutb(w_n7154_19[1]),.doutc(w_n7154_19[2]),.din(w_n7154_6[0]));
	jspl3 jspl3_w_n7154_20(.douta(w_n7154_20[0]),.doutb(w_n7154_20[1]),.doutc(w_n7154_20[2]),.din(w_n7154_6[1]));
	jspl3 jspl3_w_n7154_21(.douta(w_n7154_21[0]),.doutb(w_n7154_21[1]),.doutc(w_n7154_21[2]),.din(w_n7154_6[2]));
	jspl3 jspl3_w_n7154_22(.douta(w_n7154_22[0]),.doutb(w_n7154_22[1]),.doutc(w_n7154_22[2]),.din(w_n7154_7[0]));
	jspl3 jspl3_w_n7154_23(.douta(w_n7154_23[0]),.doutb(w_n7154_23[1]),.doutc(w_n7154_23[2]),.din(w_n7154_7[1]));
	jspl3 jspl3_w_n7154_24(.douta(w_n7154_24[0]),.doutb(w_n7154_24[1]),.doutc(w_n7154_24[2]),.din(w_n7154_7[2]));
	jspl3 jspl3_w_n7154_25(.douta(w_n7154_25[0]),.doutb(w_n7154_25[1]),.doutc(w_n7154_25[2]),.din(w_n7154_8[0]));
	jspl3 jspl3_w_n7154_26(.douta(w_n7154_26[0]),.doutb(w_n7154_26[1]),.doutc(w_n7154_26[2]),.din(w_n7154_8[1]));
	jspl3 jspl3_w_n7154_27(.douta(w_n7154_27[0]),.doutb(w_n7154_27[1]),.doutc(w_n7154_27[2]),.din(w_n7154_8[2]));
	jspl3 jspl3_w_n7154_28(.douta(w_n7154_28[0]),.doutb(w_n7154_28[1]),.doutc(w_n7154_28[2]),.din(w_n7154_9[0]));
	jspl3 jspl3_w_n7154_29(.douta(w_n7154_29[0]),.doutb(w_n7154_29[1]),.doutc(w_n7154_29[2]),.din(w_n7154_9[1]));
	jspl3 jspl3_w_n7154_30(.douta(w_n7154_30[0]),.doutb(w_n7154_30[1]),.doutc(w_n7154_30[2]),.din(w_n7154_9[2]));
	jspl3 jspl3_w_n7154_31(.douta(w_n7154_31[0]),.doutb(w_n7154_31[1]),.doutc(w_n7154_31[2]),.din(w_n7154_10[0]));
	jspl3 jspl3_w_n7154_32(.douta(w_n7154_32[0]),.doutb(w_n7154_32[1]),.doutc(w_n7154_32[2]),.din(w_n7154_10[1]));
	jspl3 jspl3_w_n7154_33(.douta(w_n7154_33[0]),.doutb(w_n7154_33[1]),.doutc(w_n7154_33[2]),.din(w_n7154_10[2]));
	jspl3 jspl3_w_n7154_34(.douta(w_n7154_34[0]),.doutb(w_n7154_34[1]),.doutc(w_n7154_34[2]),.din(w_n7154_11[0]));
	jspl3 jspl3_w_n7154_35(.douta(w_n7154_35[0]),.doutb(w_n7154_35[1]),.doutc(w_n7154_35[2]),.din(w_n7154_11[1]));
	jspl3 jspl3_w_n7154_36(.douta(w_n7154_36[0]),.doutb(w_n7154_36[1]),.doutc(w_n7154_36[2]),.din(w_n7154_11[2]));
	jspl3 jspl3_w_n7154_37(.douta(w_n7154_37[0]),.doutb(w_n7154_37[1]),.doutc(w_n7154_37[2]),.din(w_n7154_12[0]));
	jspl3 jspl3_w_n7154_38(.douta(w_n7154_38[0]),.doutb(w_n7154_38[1]),.doutc(w_n7154_38[2]),.din(w_n7154_12[1]));
	jspl3 jspl3_w_n7154_39(.douta(w_n7154_39[0]),.doutb(w_n7154_39[1]),.doutc(w_n7154_39[2]),.din(w_n7154_12[2]));
	jspl3 jspl3_w_n7154_40(.douta(w_n7154_40[0]),.doutb(w_n7154_40[1]),.doutc(w_n7154_40[2]),.din(w_n7154_13[0]));
	jspl3 jspl3_w_n7154_41(.douta(w_n7154_41[0]),.doutb(w_n7154_41[1]),.doutc(w_n7154_41[2]),.din(w_n7154_13[1]));
	jspl3 jspl3_w_n7154_42(.douta(w_n7154_42[0]),.doutb(w_n7154_42[1]),.doutc(w_n7154_42[2]),.din(w_n7154_13[2]));
	jspl3 jspl3_w_n7154_43(.douta(w_n7154_43[0]),.doutb(w_n7154_43[1]),.doutc(w_n7154_43[2]),.din(w_n7154_14[0]));
	jspl3 jspl3_w_n7154_44(.douta(w_n7154_44[0]),.doutb(w_n7154_44[1]),.doutc(w_n7154_44[2]),.din(w_n7154_14[1]));
	jspl3 jspl3_w_n7154_45(.douta(w_n7154_45[0]),.doutb(w_n7154_45[1]),.doutc(w_n7154_45[2]),.din(w_n7154_14[2]));
	jspl3 jspl3_w_n7154_46(.douta(w_n7154_46[0]),.doutb(w_n7154_46[1]),.doutc(w_n7154_46[2]),.din(w_n7154_15[0]));
	jspl3 jspl3_w_n7154_47(.douta(w_n7154_47[0]),.doutb(w_n7154_47[1]),.doutc(w_n7154_47[2]),.din(w_n7154_15[1]));
	jspl3 jspl3_w_n7154_48(.douta(w_n7154_48[0]),.doutb(w_n7154_48[1]),.doutc(w_n7154_48[2]),.din(w_n7154_15[2]));
	jspl3 jspl3_w_n7154_49(.douta(w_n7154_49[0]),.doutb(w_n7154_49[1]),.doutc(w_n7154_49[2]),.din(w_n7154_16[0]));
	jspl3 jspl3_w_n7154_50(.douta(w_n7154_50[0]),.doutb(w_n7154_50[1]),.doutc(w_n7154_50[2]),.din(w_n7154_16[1]));
	jspl3 jspl3_w_n7154_51(.douta(w_n7154_51[0]),.doutb(w_n7154_51[1]),.doutc(w_n7154_51[2]),.din(w_n7154_16[2]));
	jspl3 jspl3_w_n7154_52(.douta(w_n7154_52[0]),.doutb(w_n7154_52[1]),.doutc(w_n7154_52[2]),.din(w_n7154_17[0]));
	jspl3 jspl3_w_n7154_53(.douta(w_n7154_53[0]),.doutb(w_n7154_53[1]),.doutc(w_n7154_53[2]),.din(w_n7154_17[1]));
	jspl3 jspl3_w_n7156_0(.douta(w_n7156_0[0]),.doutb(w_n7156_0[1]),.doutc(w_n7156_0[2]),.din(n7156));
	jspl3 jspl3_w_n7156_1(.douta(w_n7156_1[0]),.doutb(w_n7156_1[1]),.doutc(w_n7156_1[2]),.din(w_n7156_0[0]));
	jspl jspl_w_n7157_0(.douta(w_n7157_0[0]),.doutb(w_n7157_0[1]),.din(n7157));
	jspl3 jspl3_w_n7158_0(.douta(w_n7158_0[0]),.doutb(w_n7158_0[1]),.doutc(w_n7158_0[2]),.din(n7158));
	jspl jspl_w_n7159_0(.douta(w_n7159_0[0]),.doutb(w_n7159_0[1]),.din(n7159));
	jspl3 jspl3_w_n7161_0(.douta(w_n7161_0[0]),.doutb(w_n7161_0[1]),.doutc(w_n7161_0[2]),.din(n7161));
	jspl jspl_w_n7162_0(.douta(w_n7162_0[0]),.doutb(w_n7162_0[1]),.din(n7162));
	jspl3 jspl3_w_n7169_0(.douta(w_n7169_0[0]),.doutb(w_n7169_0[1]),.doutc(w_n7169_0[2]),.din(n7169));
	jspl jspl_w_n7170_0(.douta(w_n7170_0[0]),.doutb(w_n7170_0[1]),.din(n7170));
	jspl jspl_w_n7173_0(.douta(w_n7173_0[0]),.doutb(w_n7173_0[1]),.din(n7173));
	jspl3 jspl3_w_n7178_0(.douta(w_n7178_0[0]),.doutb(w_n7178_0[1]),.doutc(w_n7178_0[2]),.din(n7178));
	jspl3 jspl3_w_n7180_0(.douta(w_n7180_0[0]),.doutb(w_n7180_0[1]),.doutc(w_n7180_0[2]),.din(n7180));
	jspl jspl_w_n7181_0(.douta(w_n7181_0[0]),.doutb(w_n7181_0[1]),.din(n7181));
	jspl3 jspl3_w_n7185_0(.douta(w_n7185_0[0]),.doutb(w_n7185_0[1]),.doutc(w_n7185_0[2]),.din(n7185));
	jspl3 jspl3_w_n7188_0(.douta(w_n7188_0[0]),.doutb(w_n7188_0[1]),.doutc(w_n7188_0[2]),.din(n7188));
	jspl jspl_w_n7189_0(.douta(w_n7189_0[0]),.doutb(w_n7189_0[1]),.din(n7189));
	jspl3 jspl3_w_n7193_0(.douta(w_n7193_0[0]),.doutb(w_n7193_0[1]),.doutc(w_n7193_0[2]),.din(n7193));
	jspl3 jspl3_w_n7195_0(.douta(w_n7195_0[0]),.doutb(w_n7195_0[1]),.doutc(w_n7195_0[2]),.din(n7195));
	jspl jspl_w_n7196_0(.douta(w_n7196_0[0]),.doutb(w_n7196_0[1]),.din(n7196));
	jspl3 jspl3_w_n7200_0(.douta(w_n7200_0[0]),.doutb(w_n7200_0[1]),.doutc(w_n7200_0[2]),.din(n7200));
	jspl3 jspl3_w_n7203_0(.douta(w_n7203_0[0]),.doutb(w_n7203_0[1]),.doutc(w_n7203_0[2]),.din(n7203));
	jspl jspl_w_n7204_0(.douta(w_n7204_0[0]),.doutb(w_n7204_0[1]),.din(n7204));
	jspl3 jspl3_w_n7208_0(.douta(w_n7208_0[0]),.doutb(w_n7208_0[1]),.doutc(w_n7208_0[2]),.din(n7208));
	jspl3 jspl3_w_n7211_0(.douta(w_n7211_0[0]),.doutb(w_n7211_0[1]),.doutc(w_n7211_0[2]),.din(n7211));
	jspl jspl_w_n7212_0(.douta(w_n7212_0[0]),.doutb(w_n7212_0[1]),.din(n7212));
	jspl3 jspl3_w_n7216_0(.douta(w_n7216_0[0]),.doutb(w_n7216_0[1]),.doutc(w_n7216_0[2]),.din(n7216));
	jspl3 jspl3_w_n7219_0(.douta(w_n7219_0[0]),.doutb(w_n7219_0[1]),.doutc(w_n7219_0[2]),.din(n7219));
	jspl jspl_w_n7220_0(.douta(w_n7220_0[0]),.doutb(w_n7220_0[1]),.din(n7220));
	jspl3 jspl3_w_n7224_0(.douta(w_n7224_0[0]),.doutb(w_n7224_0[1]),.doutc(w_n7224_0[2]),.din(n7224));
	jspl3 jspl3_w_n7226_0(.douta(w_n7226_0[0]),.doutb(w_n7226_0[1]),.doutc(w_n7226_0[2]),.din(n7226));
	jspl jspl_w_n7227_0(.douta(w_n7227_0[0]),.doutb(w_n7227_0[1]),.din(n7227));
	jspl3 jspl3_w_n7231_0(.douta(w_n7231_0[0]),.doutb(w_n7231_0[1]),.doutc(w_n7231_0[2]),.din(n7231));
	jspl3 jspl3_w_n7234_0(.douta(w_n7234_0[0]),.doutb(w_n7234_0[1]),.doutc(w_n7234_0[2]),.din(n7234));
	jspl jspl_w_n7235_0(.douta(w_n7235_0[0]),.doutb(w_n7235_0[1]),.din(n7235));
	jspl3 jspl3_w_n7239_0(.douta(w_n7239_0[0]),.doutb(w_n7239_0[1]),.doutc(w_n7239_0[2]),.din(n7239));
	jspl3 jspl3_w_n7241_0(.douta(w_n7241_0[0]),.doutb(w_n7241_0[1]),.doutc(w_n7241_0[2]),.din(n7241));
	jspl jspl_w_n7242_0(.douta(w_n7242_0[0]),.doutb(w_n7242_0[1]),.din(n7242));
	jspl3 jspl3_w_n7246_0(.douta(w_n7246_0[0]),.doutb(w_n7246_0[1]),.doutc(w_n7246_0[2]),.din(n7246));
	jspl3 jspl3_w_n7249_0(.douta(w_n7249_0[0]),.doutb(w_n7249_0[1]),.doutc(w_n7249_0[2]),.din(n7249));
	jspl jspl_w_n7250_0(.douta(w_n7250_0[0]),.doutb(w_n7250_0[1]),.din(n7250));
	jspl3 jspl3_w_n7254_0(.douta(w_n7254_0[0]),.doutb(w_n7254_0[1]),.doutc(w_n7254_0[2]),.din(n7254));
	jspl3 jspl3_w_n7256_0(.douta(w_n7256_0[0]),.doutb(w_n7256_0[1]),.doutc(w_n7256_0[2]),.din(n7256));
	jspl jspl_w_n7257_0(.douta(w_n7257_0[0]),.doutb(w_n7257_0[1]),.din(n7257));
	jspl3 jspl3_w_n7261_0(.douta(w_n7261_0[0]),.doutb(w_n7261_0[1]),.doutc(w_n7261_0[2]),.din(n7261));
	jspl3 jspl3_w_n7264_0(.douta(w_n7264_0[0]),.doutb(w_n7264_0[1]),.doutc(w_n7264_0[2]),.din(n7264));
	jspl jspl_w_n7265_0(.douta(w_n7265_0[0]),.doutb(w_n7265_0[1]),.din(n7265));
	jspl3 jspl3_w_n7269_0(.douta(w_n7269_0[0]),.doutb(w_n7269_0[1]),.doutc(w_n7269_0[2]),.din(n7269));
	jspl3 jspl3_w_n7271_0(.douta(w_n7271_0[0]),.doutb(w_n7271_0[1]),.doutc(w_n7271_0[2]),.din(n7271));
	jspl jspl_w_n7272_0(.douta(w_n7272_0[0]),.doutb(w_n7272_0[1]),.din(n7272));
	jspl3 jspl3_w_n7276_0(.douta(w_n7276_0[0]),.doutb(w_n7276_0[1]),.doutc(w_n7276_0[2]),.din(n7276));
	jspl3 jspl3_w_n7279_0(.douta(w_n7279_0[0]),.doutb(w_n7279_0[1]),.doutc(w_n7279_0[2]),.din(n7279));
	jspl jspl_w_n7280_0(.douta(w_n7280_0[0]),.doutb(w_n7280_0[1]),.din(n7280));
	jspl3 jspl3_w_n7284_0(.douta(w_n7284_0[0]),.doutb(w_n7284_0[1]),.doutc(w_n7284_0[2]),.din(n7284));
	jspl3 jspl3_w_n7287_0(.douta(w_n7287_0[0]),.doutb(w_n7287_0[1]),.doutc(w_n7287_0[2]),.din(n7287));
	jspl jspl_w_n7288_0(.douta(w_n7288_0[0]),.doutb(w_n7288_0[1]),.din(n7288));
	jspl3 jspl3_w_n7292_0(.douta(w_n7292_0[0]),.doutb(w_n7292_0[1]),.doutc(w_n7292_0[2]),.din(n7292));
	jspl3 jspl3_w_n7295_0(.douta(w_n7295_0[0]),.doutb(w_n7295_0[1]),.doutc(w_n7295_0[2]),.din(n7295));
	jspl jspl_w_n7296_0(.douta(w_n7296_0[0]),.doutb(w_n7296_0[1]),.din(n7296));
	jspl3 jspl3_w_n7300_0(.douta(w_n7300_0[0]),.doutb(w_n7300_0[1]),.doutc(w_n7300_0[2]),.din(n7300));
	jspl3 jspl3_w_n7302_0(.douta(w_n7302_0[0]),.doutb(w_n7302_0[1]),.doutc(w_n7302_0[2]),.din(n7302));
	jspl jspl_w_n7303_0(.douta(w_n7303_0[0]),.doutb(w_n7303_0[1]),.din(n7303));
	jspl3 jspl3_w_n7307_0(.douta(w_n7307_0[0]),.doutb(w_n7307_0[1]),.doutc(w_n7307_0[2]),.din(n7307));
	jspl3 jspl3_w_n7309_0(.douta(w_n7309_0[0]),.doutb(w_n7309_0[1]),.doutc(w_n7309_0[2]),.din(n7309));
	jspl jspl_w_n7310_0(.douta(w_n7310_0[0]),.doutb(w_n7310_0[1]),.din(n7310));
	jspl3 jspl3_w_n7314_0(.douta(w_n7314_0[0]),.doutb(w_n7314_0[1]),.doutc(w_n7314_0[2]),.din(n7314));
	jspl3 jspl3_w_n7316_0(.douta(w_n7316_0[0]),.doutb(w_n7316_0[1]),.doutc(w_n7316_0[2]),.din(n7316));
	jspl jspl_w_n7317_0(.douta(w_n7317_0[0]),.doutb(w_n7317_0[1]),.din(n7317));
	jspl3 jspl3_w_n7321_0(.douta(w_n7321_0[0]),.doutb(w_n7321_0[1]),.doutc(w_n7321_0[2]),.din(n7321));
	jspl3 jspl3_w_n7324_0(.douta(w_n7324_0[0]),.doutb(w_n7324_0[1]),.doutc(w_n7324_0[2]),.din(n7324));
	jspl jspl_w_n7325_0(.douta(w_n7325_0[0]),.doutb(w_n7325_0[1]),.din(n7325));
	jspl3 jspl3_w_n7329_0(.douta(w_n7329_0[0]),.doutb(w_n7329_0[1]),.doutc(w_n7329_0[2]),.din(n7329));
	jspl3 jspl3_w_n7331_0(.douta(w_n7331_0[0]),.doutb(w_n7331_0[1]),.doutc(w_n7331_0[2]),.din(n7331));
	jspl jspl_w_n7332_0(.douta(w_n7332_0[0]),.doutb(w_n7332_0[1]),.din(n7332));
	jspl3 jspl3_w_n7336_0(.douta(w_n7336_0[0]),.doutb(w_n7336_0[1]),.doutc(w_n7336_0[2]),.din(n7336));
	jspl3 jspl3_w_n7339_0(.douta(w_n7339_0[0]),.doutb(w_n7339_0[1]),.doutc(w_n7339_0[2]),.din(n7339));
	jspl jspl_w_n7340_0(.douta(w_n7340_0[0]),.doutb(w_n7340_0[1]),.din(n7340));
	jspl3 jspl3_w_n7344_0(.douta(w_n7344_0[0]),.doutb(w_n7344_0[1]),.doutc(w_n7344_0[2]),.din(n7344));
	jspl3 jspl3_w_n7346_0(.douta(w_n7346_0[0]),.doutb(w_n7346_0[1]),.doutc(w_n7346_0[2]),.din(n7346));
	jspl jspl_w_n7347_0(.douta(w_n7347_0[0]),.doutb(w_n7347_0[1]),.din(n7347));
	jspl3 jspl3_w_n7351_0(.douta(w_n7351_0[0]),.doutb(w_n7351_0[1]),.doutc(w_n7351_0[2]),.din(n7351));
	jspl3 jspl3_w_n7354_0(.douta(w_n7354_0[0]),.doutb(w_n7354_0[1]),.doutc(w_n7354_0[2]),.din(n7354));
	jspl jspl_w_n7355_0(.douta(w_n7355_0[0]),.doutb(w_n7355_0[1]),.din(n7355));
	jspl3 jspl3_w_n7359_0(.douta(w_n7359_0[0]),.doutb(w_n7359_0[1]),.doutc(w_n7359_0[2]),.din(n7359));
	jspl3 jspl3_w_n7362_0(.douta(w_n7362_0[0]),.doutb(w_n7362_0[1]),.doutc(w_n7362_0[2]),.din(n7362));
	jspl jspl_w_n7363_0(.douta(w_n7363_0[0]),.doutb(w_n7363_0[1]),.din(n7363));
	jspl3 jspl3_w_n7367_0(.douta(w_n7367_0[0]),.doutb(w_n7367_0[1]),.doutc(w_n7367_0[2]),.din(n7367));
	jspl3 jspl3_w_n7369_0(.douta(w_n7369_0[0]),.doutb(w_n7369_0[1]),.doutc(w_n7369_0[2]),.din(n7369));
	jspl jspl_w_n7370_0(.douta(w_n7370_0[0]),.doutb(w_n7370_0[1]),.din(n7370));
	jspl3 jspl3_w_n7374_0(.douta(w_n7374_0[0]),.doutb(w_n7374_0[1]),.doutc(w_n7374_0[2]),.din(n7374));
	jspl3 jspl3_w_n7376_0(.douta(w_n7376_0[0]),.doutb(w_n7376_0[1]),.doutc(w_n7376_0[2]),.din(n7376));
	jspl jspl_w_n7377_0(.douta(w_n7377_0[0]),.doutb(w_n7377_0[1]),.din(n7377));
	jspl3 jspl3_w_n7381_0(.douta(w_n7381_0[0]),.doutb(w_n7381_0[1]),.doutc(w_n7381_0[2]),.din(n7381));
	jspl3 jspl3_w_n7383_0(.douta(w_n7383_0[0]),.doutb(w_n7383_0[1]),.doutc(w_n7383_0[2]),.din(n7383));
	jspl jspl_w_n7384_0(.douta(w_n7384_0[0]),.doutb(w_n7384_0[1]),.din(n7384));
	jspl3 jspl3_w_n7388_0(.douta(w_n7388_0[0]),.doutb(w_n7388_0[1]),.doutc(w_n7388_0[2]),.din(n7388));
	jspl3 jspl3_w_n7391_0(.douta(w_n7391_0[0]),.doutb(w_n7391_0[1]),.doutc(w_n7391_0[2]),.din(n7391));
	jspl jspl_w_n7392_0(.douta(w_n7392_0[0]),.doutb(w_n7392_0[1]),.din(n7392));
	jspl3 jspl3_w_n7396_0(.douta(w_n7396_0[0]),.doutb(w_n7396_0[1]),.doutc(w_n7396_0[2]),.din(n7396));
	jspl3 jspl3_w_n7399_0(.douta(w_n7399_0[0]),.doutb(w_n7399_0[1]),.doutc(w_n7399_0[2]),.din(n7399));
	jspl3 jspl3_w_n7402_0(.douta(w_n7402_0[0]),.doutb(w_n7402_0[1]),.doutc(w_n7402_0[2]),.din(n7402));
	jspl jspl_w_n7402_1(.douta(w_n7402_1[0]),.doutb(w_n7402_1[1]),.din(w_n7402_0[0]));
	jspl jspl_w_n7403_0(.douta(w_n7403_0[0]),.doutb(w_n7403_0[1]),.din(n7403));
	jspl jspl_w_n7406_0(.douta(w_n7406_0[0]),.doutb(w_n7406_0[1]),.din(n7406));
	jspl3 jspl3_w_n7408_0(.douta(w_n7408_0[0]),.doutb(w_n7408_0[1]),.doutc(w_n7408_0[2]),.din(n7408));
	jspl jspl_w_n7408_1(.douta(w_n7408_1[0]),.doutb(w_n7408_1[1]),.din(w_n7408_0[0]));
	jspl jspl_w_n7413_0(.douta(w_n7413_0[0]),.doutb(w_n7413_0[1]),.din(n7413));
	jspl jspl_w_n7415_0(.douta(w_n7415_0[0]),.doutb(w_n7415_0[1]),.din(n7415));
	jspl3 jspl3_w_n7419_0(.douta(w_n7419_0[0]),.doutb(w_n7419_0[1]),.doutc(w_n7419_0[2]),.din(n7419));
	jspl3 jspl3_w_n7421_0(.douta(w_n7421_0[0]),.doutb(w_n7421_0[1]),.doutc(w_n7421_0[2]),.din(n7421));
	jspl3 jspl3_w_n7421_1(.douta(w_n7421_1[0]),.doutb(w_n7421_1[1]),.doutc(w_n7421_1[2]),.din(w_n7421_0[0]));
	jspl jspl_w_n7422_0(.douta(w_n7422_0[0]),.doutb(w_n7422_0[1]),.din(n7422));
	jspl3 jspl3_w_n7423_0(.douta(w_n7423_0[0]),.doutb(w_n7423_0[1]),.doutc(w_n7423_0[2]),.din(n7423));
	jspl jspl_w_n7424_0(.douta(w_n7424_0[0]),.doutb(w_n7424_0[1]),.din(n7424));
	jspl3 jspl3_w_n7425_0(.douta(w_n7425_0[0]),.doutb(w_n7425_0[1]),.doutc(w_n7425_0[2]),.din(n7425));
	jspl jspl_w_n7426_0(.douta(w_n7426_0[0]),.doutb(w_n7426_0[1]),.din(n7426));
	jspl jspl_w_n7465_0(.douta(w_n7465_0[0]),.doutb(w_n7465_0[1]),.din(n7465));
	jspl jspl_w_n7576_0(.douta(w_n7576_0[0]),.doutb(w_n7576_0[1]),.din(n7576));
	jspl3 jspl3_w_n7581_0(.douta(w_n7581_0[0]),.doutb(w_n7581_0[1]),.doutc(w_n7581_0[2]),.din(n7581));
	jspl3 jspl3_w_n7581_1(.douta(w_n7581_1[0]),.doutb(w_n7581_1[1]),.doutc(w_n7581_1[2]),.din(w_n7581_0[0]));
	jspl3 jspl3_w_n7581_2(.douta(w_n7581_2[0]),.doutb(w_n7581_2[1]),.doutc(w_n7581_2[2]),.din(w_n7581_0[1]));
	jspl3 jspl3_w_n7581_3(.douta(w_n7581_3[0]),.doutb(w_n7581_3[1]),.doutc(w_n7581_3[2]),.din(w_n7581_0[2]));
	jspl3 jspl3_w_n7581_4(.douta(w_n7581_4[0]),.doutb(w_n7581_4[1]),.doutc(w_n7581_4[2]),.din(w_n7581_1[0]));
	jspl3 jspl3_w_n7581_5(.douta(w_n7581_5[0]),.doutb(w_n7581_5[1]),.doutc(w_n7581_5[2]),.din(w_n7581_1[1]));
	jspl3 jspl3_w_n7581_6(.douta(w_n7581_6[0]),.doutb(w_n7581_6[1]),.doutc(w_n7581_6[2]),.din(w_n7581_1[2]));
	jspl3 jspl3_w_n7581_7(.douta(w_n7581_7[0]),.doutb(w_n7581_7[1]),.doutc(w_n7581_7[2]),.din(w_n7581_2[0]));
	jspl3 jspl3_w_n7581_8(.douta(w_n7581_8[0]),.doutb(w_n7581_8[1]),.doutc(w_n7581_8[2]),.din(w_n7581_2[1]));
	jspl3 jspl3_w_n7581_9(.douta(w_n7581_9[0]),.doutb(w_n7581_9[1]),.doutc(w_n7581_9[2]),.din(w_n7581_2[2]));
	jspl3 jspl3_w_n7581_10(.douta(w_n7581_10[0]),.doutb(w_n7581_10[1]),.doutc(w_n7581_10[2]),.din(w_n7581_3[0]));
	jspl3 jspl3_w_n7581_11(.douta(w_n7581_11[0]),.doutb(w_n7581_11[1]),.doutc(w_n7581_11[2]),.din(w_n7581_3[1]));
	jspl3 jspl3_w_n7581_12(.douta(w_n7581_12[0]),.doutb(w_n7581_12[1]),.doutc(w_n7581_12[2]),.din(w_n7581_3[2]));
	jspl3 jspl3_w_n7581_13(.douta(w_n7581_13[0]),.doutb(w_n7581_13[1]),.doutc(w_n7581_13[2]),.din(w_n7581_4[0]));
	jspl3 jspl3_w_n7581_14(.douta(w_n7581_14[0]),.doutb(w_n7581_14[1]),.doutc(w_n7581_14[2]),.din(w_n7581_4[1]));
	jspl3 jspl3_w_n7581_15(.douta(w_n7581_15[0]),.doutb(w_n7581_15[1]),.doutc(w_n7581_15[2]),.din(w_n7581_4[2]));
	jspl3 jspl3_w_n7581_16(.douta(w_n7581_16[0]),.doutb(w_n7581_16[1]),.doutc(w_n7581_16[2]),.din(w_n7581_5[0]));
	jspl3 jspl3_w_n7581_17(.douta(w_n7581_17[0]),.doutb(w_n7581_17[1]),.doutc(w_n7581_17[2]),.din(w_n7581_5[1]));
	jspl3 jspl3_w_n7581_18(.douta(w_n7581_18[0]),.doutb(w_n7581_18[1]),.doutc(w_n7581_18[2]),.din(w_n7581_5[2]));
	jspl3 jspl3_w_n7581_19(.douta(w_n7581_19[0]),.doutb(w_n7581_19[1]),.doutc(w_n7581_19[2]),.din(w_n7581_6[0]));
	jspl3 jspl3_w_n7581_20(.douta(w_n7581_20[0]),.doutb(w_n7581_20[1]),.doutc(w_n7581_20[2]),.din(w_n7581_6[1]));
	jspl3 jspl3_w_n7581_21(.douta(w_n7581_21[0]),.doutb(w_n7581_21[1]),.doutc(w_n7581_21[2]),.din(w_n7581_6[2]));
	jspl3 jspl3_w_n7581_22(.douta(w_n7581_22[0]),.doutb(w_n7581_22[1]),.doutc(w_n7581_22[2]),.din(w_n7581_7[0]));
	jspl3 jspl3_w_n7581_23(.douta(w_n7581_23[0]),.doutb(w_n7581_23[1]),.doutc(w_n7581_23[2]),.din(w_n7581_7[1]));
	jspl3 jspl3_w_n7581_24(.douta(w_n7581_24[0]),.doutb(w_n7581_24[1]),.doutc(w_n7581_24[2]),.din(w_n7581_7[2]));
	jspl3 jspl3_w_n7581_25(.douta(w_n7581_25[0]),.doutb(w_n7581_25[1]),.doutc(w_n7581_25[2]),.din(w_n7581_8[0]));
	jspl3 jspl3_w_n7581_26(.douta(w_n7581_26[0]),.doutb(w_n7581_26[1]),.doutc(w_n7581_26[2]),.din(w_n7581_8[1]));
	jspl3 jspl3_w_n7581_27(.douta(w_n7581_27[0]),.doutb(w_n7581_27[1]),.doutc(w_n7581_27[2]),.din(w_n7581_8[2]));
	jspl3 jspl3_w_n7581_28(.douta(w_n7581_28[0]),.doutb(w_n7581_28[1]),.doutc(w_n7581_28[2]),.din(w_n7581_9[0]));
	jspl3 jspl3_w_n7581_29(.douta(w_n7581_29[0]),.doutb(w_n7581_29[1]),.doutc(w_n7581_29[2]),.din(w_n7581_9[1]));
	jspl3 jspl3_w_n7581_30(.douta(w_n7581_30[0]),.doutb(w_n7581_30[1]),.doutc(w_n7581_30[2]),.din(w_n7581_9[2]));
	jspl3 jspl3_w_n7581_31(.douta(w_n7581_31[0]),.doutb(w_n7581_31[1]),.doutc(w_n7581_31[2]),.din(w_n7581_10[0]));
	jspl3 jspl3_w_n7581_32(.douta(w_n7581_32[0]),.doutb(w_n7581_32[1]),.doutc(w_n7581_32[2]),.din(w_n7581_10[1]));
	jspl3 jspl3_w_n7581_33(.douta(w_n7581_33[0]),.doutb(w_n7581_33[1]),.doutc(w_n7581_33[2]),.din(w_n7581_10[2]));
	jspl3 jspl3_w_n7581_34(.douta(w_n7581_34[0]),.doutb(w_n7581_34[1]),.doutc(w_n7581_34[2]),.din(w_n7581_11[0]));
	jspl3 jspl3_w_n7581_35(.douta(w_n7581_35[0]),.doutb(w_n7581_35[1]),.doutc(w_n7581_35[2]),.din(w_n7581_11[1]));
	jspl3 jspl3_w_n7581_36(.douta(w_n7581_36[0]),.doutb(w_n7581_36[1]),.doutc(w_n7581_36[2]),.din(w_n7581_11[2]));
	jspl3 jspl3_w_n7581_37(.douta(w_n7581_37[0]),.doutb(w_n7581_37[1]),.doutc(w_n7581_37[2]),.din(w_n7581_12[0]));
	jspl jspl_w_n7581_38(.douta(w_n7581_38[0]),.doutb(w_n7581_38[1]),.din(w_n7581_12[1]));
	jspl jspl_w_n7582_0(.douta(w_n7582_0[0]),.doutb(w_n7582_0[1]),.din(n7582));
	jspl jspl_w_n7583_0(.douta(w_n7583_0[0]),.doutb(w_n7583_0[1]),.din(n7583));
	jspl3 jspl3_w_n7585_0(.douta(w_n7585_0[0]),.doutb(w_n7585_0[1]),.doutc(w_n7585_0[2]),.din(n7585));
	jspl jspl_w_n7586_0(.douta(w_n7586_0[0]),.doutb(w_n7586_0[1]),.din(n7586));
	jspl jspl_w_n7592_0(.douta(w_n7592_0[0]),.doutb(w_n7592_0[1]),.din(n7592));
	jspl jspl_w_n7593_0(.douta(w_n7593_0[0]),.doutb(w_n7593_0[1]),.din(n7593));
	jspl3 jspl3_w_n7595_0(.douta(w_n7595_0[0]),.doutb(w_n7595_0[1]),.doutc(w_n7595_0[2]),.din(n7595));
	jspl jspl_w_n7596_0(.douta(w_n7596_0[0]),.doutb(w_n7596_0[1]),.din(n7596));
	jspl jspl_w_n7599_0(.douta(w_n7599_0[0]),.doutb(w_n7599_0[1]),.din(n7599));
	jspl3 jspl3_w_n7602_0(.douta(w_n7602_0[0]),.doutb(w_n7602_0[1]),.doutc(w_n7602_0[2]),.din(n7602));
	jspl jspl_w_n7603_0(.douta(w_n7603_0[0]),.doutb(w_n7603_0[1]),.din(n7603));
	jspl jspl_w_n7607_0(.douta(w_n7607_0[0]),.doutb(w_n7607_0[1]),.din(n7607));
	jspl jspl_w_n7608_0(.douta(w_n7608_0[0]),.doutb(w_n7608_0[1]),.din(n7608));
	jspl3 jspl3_w_n7610_0(.douta(w_n7610_0[0]),.doutb(w_n7610_0[1]),.doutc(w_n7610_0[2]),.din(n7610));
	jspl jspl_w_n7611_0(.douta(w_n7611_0[0]),.doutb(w_n7611_0[1]),.din(n7611));
	jspl jspl_w_n7615_0(.douta(w_n7615_0[0]),.doutb(w_n7615_0[1]),.din(n7615));
	jspl3 jspl3_w_n7617_0(.douta(w_n7617_0[0]),.doutb(w_n7617_0[1]),.doutc(w_n7617_0[2]),.din(n7617));
	jspl jspl_w_n7618_0(.douta(w_n7618_0[0]),.doutb(w_n7618_0[1]),.din(n7618));
	jspl jspl_w_n7622_0(.douta(w_n7622_0[0]),.doutb(w_n7622_0[1]),.din(n7622));
	jspl jspl_w_n7623_0(.douta(w_n7623_0[0]),.doutb(w_n7623_0[1]),.din(n7623));
	jspl3 jspl3_w_n7625_0(.douta(w_n7625_0[0]),.doutb(w_n7625_0[1]),.doutc(w_n7625_0[2]),.din(n7625));
	jspl jspl_w_n7626_0(.douta(w_n7626_0[0]),.doutb(w_n7626_0[1]),.din(n7626));
	jspl jspl_w_n7630_0(.douta(w_n7630_0[0]),.doutb(w_n7630_0[1]),.din(n7630));
	jspl3 jspl3_w_n7632_0(.douta(w_n7632_0[0]),.doutb(w_n7632_0[1]),.doutc(w_n7632_0[2]),.din(n7632));
	jspl jspl_w_n7633_0(.douta(w_n7633_0[0]),.doutb(w_n7633_0[1]),.din(n7633));
	jspl jspl_w_n7637_0(.douta(w_n7637_0[0]),.doutb(w_n7637_0[1]),.din(n7637));
	jspl3 jspl3_w_n7639_0(.douta(w_n7639_0[0]),.doutb(w_n7639_0[1]),.doutc(w_n7639_0[2]),.din(n7639));
	jspl jspl_w_n7640_0(.douta(w_n7640_0[0]),.doutb(w_n7640_0[1]),.din(n7640));
	jspl jspl_w_n7644_0(.douta(w_n7644_0[0]),.doutb(w_n7644_0[1]),.din(n7644));
	jspl3 jspl3_w_n7646_0(.douta(w_n7646_0[0]),.doutb(w_n7646_0[1]),.doutc(w_n7646_0[2]),.din(n7646));
	jspl jspl_w_n7647_0(.douta(w_n7647_0[0]),.doutb(w_n7647_0[1]),.din(n7647));
	jspl jspl_w_n7651_0(.douta(w_n7651_0[0]),.doutb(w_n7651_0[1]),.din(n7651));
	jspl jspl_w_n7652_0(.douta(w_n7652_0[0]),.doutb(w_n7652_0[1]),.din(n7652));
	jspl3 jspl3_w_n7654_0(.douta(w_n7654_0[0]),.doutb(w_n7654_0[1]),.doutc(w_n7654_0[2]),.din(n7654));
	jspl jspl_w_n7655_0(.douta(w_n7655_0[0]),.doutb(w_n7655_0[1]),.din(n7655));
	jspl jspl_w_n7659_0(.douta(w_n7659_0[0]),.doutb(w_n7659_0[1]),.din(n7659));
	jspl3 jspl3_w_n7661_0(.douta(w_n7661_0[0]),.doutb(w_n7661_0[1]),.doutc(w_n7661_0[2]),.din(n7661));
	jspl jspl_w_n7662_0(.douta(w_n7662_0[0]),.doutb(w_n7662_0[1]),.din(n7662));
	jspl jspl_w_n7666_0(.douta(w_n7666_0[0]),.doutb(w_n7666_0[1]),.din(n7666));
	jspl jspl_w_n7667_0(.douta(w_n7667_0[0]),.doutb(w_n7667_0[1]),.din(n7667));
	jspl3 jspl3_w_n7669_0(.douta(w_n7669_0[0]),.doutb(w_n7669_0[1]),.doutc(w_n7669_0[2]),.din(n7669));
	jspl jspl_w_n7670_0(.douta(w_n7670_0[0]),.doutb(w_n7670_0[1]),.din(n7670));
	jspl jspl_w_n7674_0(.douta(w_n7674_0[0]),.doutb(w_n7674_0[1]),.din(n7674));
	jspl3 jspl3_w_n7676_0(.douta(w_n7676_0[0]),.doutb(w_n7676_0[1]),.doutc(w_n7676_0[2]),.din(n7676));
	jspl jspl_w_n7677_0(.douta(w_n7677_0[0]),.doutb(w_n7677_0[1]),.din(n7677));
	jspl jspl_w_n7681_0(.douta(w_n7681_0[0]),.doutb(w_n7681_0[1]),.din(n7681));
	jspl jspl_w_n7682_0(.douta(w_n7682_0[0]),.doutb(w_n7682_0[1]),.din(n7682));
	jspl3 jspl3_w_n7684_0(.douta(w_n7684_0[0]),.doutb(w_n7684_0[1]),.doutc(w_n7684_0[2]),.din(n7684));
	jspl jspl_w_n7685_0(.douta(w_n7685_0[0]),.doutb(w_n7685_0[1]),.din(n7685));
	jspl jspl_w_n7689_0(.douta(w_n7689_0[0]),.doutb(w_n7689_0[1]),.din(n7689));
	jspl3 jspl3_w_n7691_0(.douta(w_n7691_0[0]),.doutb(w_n7691_0[1]),.doutc(w_n7691_0[2]),.din(n7691));
	jspl jspl_w_n7692_0(.douta(w_n7692_0[0]),.doutb(w_n7692_0[1]),.din(n7692));
	jspl jspl_w_n7696_0(.douta(w_n7696_0[0]),.doutb(w_n7696_0[1]),.din(n7696));
	jspl jspl_w_n7697_0(.douta(w_n7697_0[0]),.doutb(w_n7697_0[1]),.din(n7697));
	jspl3 jspl3_w_n7699_0(.douta(w_n7699_0[0]),.doutb(w_n7699_0[1]),.doutc(w_n7699_0[2]),.din(n7699));
	jspl jspl_w_n7700_0(.douta(w_n7700_0[0]),.doutb(w_n7700_0[1]),.din(n7700));
	jspl jspl_w_n7704_0(.douta(w_n7704_0[0]),.doutb(w_n7704_0[1]),.din(n7704));
	jspl3 jspl3_w_n7706_0(.douta(w_n7706_0[0]),.doutb(w_n7706_0[1]),.doutc(w_n7706_0[2]),.din(n7706));
	jspl jspl_w_n7707_0(.douta(w_n7707_0[0]),.doutb(w_n7707_0[1]),.din(n7707));
	jspl jspl_w_n7711_0(.douta(w_n7711_0[0]),.doutb(w_n7711_0[1]),.din(n7711));
	jspl3 jspl3_w_n7713_0(.douta(w_n7713_0[0]),.doutb(w_n7713_0[1]),.doutc(w_n7713_0[2]),.din(n7713));
	jspl jspl_w_n7714_0(.douta(w_n7714_0[0]),.doutb(w_n7714_0[1]),.din(n7714));
	jspl jspl_w_n7718_0(.douta(w_n7718_0[0]),.doutb(w_n7718_0[1]),.din(n7718));
	jspl3 jspl3_w_n7720_0(.douta(w_n7720_0[0]),.doutb(w_n7720_0[1]),.doutc(w_n7720_0[2]),.din(n7720));
	jspl jspl_w_n7721_0(.douta(w_n7721_0[0]),.doutb(w_n7721_0[1]),.din(n7721));
	jspl jspl_w_n7725_0(.douta(w_n7725_0[0]),.doutb(w_n7725_0[1]),.din(n7725));
	jspl jspl_w_n7726_0(.douta(w_n7726_0[0]),.doutb(w_n7726_0[1]),.din(n7726));
	jspl3 jspl3_w_n7728_0(.douta(w_n7728_0[0]),.doutb(w_n7728_0[1]),.doutc(w_n7728_0[2]),.din(n7728));
	jspl jspl_w_n7729_0(.douta(w_n7729_0[0]),.doutb(w_n7729_0[1]),.din(n7729));
	jspl jspl_w_n7733_0(.douta(w_n7733_0[0]),.doutb(w_n7733_0[1]),.din(n7733));
	jspl jspl_w_n7734_0(.douta(w_n7734_0[0]),.doutb(w_n7734_0[1]),.din(n7734));
	jspl3 jspl3_w_n7736_0(.douta(w_n7736_0[0]),.doutb(w_n7736_0[1]),.doutc(w_n7736_0[2]),.din(n7736));
	jspl jspl_w_n7737_0(.douta(w_n7737_0[0]),.doutb(w_n7737_0[1]),.din(n7737));
	jspl jspl_w_n7741_0(.douta(w_n7741_0[0]),.doutb(w_n7741_0[1]),.din(n7741));
	jspl jspl_w_n7742_0(.douta(w_n7742_0[0]),.doutb(w_n7742_0[1]),.din(n7742));
	jspl3 jspl3_w_n7744_0(.douta(w_n7744_0[0]),.doutb(w_n7744_0[1]),.doutc(w_n7744_0[2]),.din(n7744));
	jspl jspl_w_n7745_0(.douta(w_n7745_0[0]),.doutb(w_n7745_0[1]),.din(n7745));
	jspl jspl_w_n7749_0(.douta(w_n7749_0[0]),.doutb(w_n7749_0[1]),.din(n7749));
	jspl3 jspl3_w_n7751_0(.douta(w_n7751_0[0]),.doutb(w_n7751_0[1]),.doutc(w_n7751_0[2]),.din(n7751));
	jspl jspl_w_n7752_0(.douta(w_n7752_0[0]),.doutb(w_n7752_0[1]),.din(n7752));
	jspl jspl_w_n7756_0(.douta(w_n7756_0[0]),.doutb(w_n7756_0[1]),.din(n7756));
	jspl jspl_w_n7757_0(.douta(w_n7757_0[0]),.doutb(w_n7757_0[1]),.din(n7757));
	jspl3 jspl3_w_n7759_0(.douta(w_n7759_0[0]),.doutb(w_n7759_0[1]),.doutc(w_n7759_0[2]),.din(n7759));
	jspl jspl_w_n7760_0(.douta(w_n7760_0[0]),.doutb(w_n7760_0[1]),.din(n7760));
	jspl jspl_w_n7764_0(.douta(w_n7764_0[0]),.doutb(w_n7764_0[1]),.din(n7764));
	jspl3 jspl3_w_n7766_0(.douta(w_n7766_0[0]),.doutb(w_n7766_0[1]),.doutc(w_n7766_0[2]),.din(n7766));
	jspl jspl_w_n7767_0(.douta(w_n7767_0[0]),.doutb(w_n7767_0[1]),.din(n7767));
	jspl jspl_w_n7771_0(.douta(w_n7771_0[0]),.doutb(w_n7771_0[1]),.din(n7771));
	jspl jspl_w_n7772_0(.douta(w_n7772_0[0]),.doutb(w_n7772_0[1]),.din(n7772));
	jspl3 jspl3_w_n7774_0(.douta(w_n7774_0[0]),.doutb(w_n7774_0[1]),.doutc(w_n7774_0[2]),.din(n7774));
	jspl jspl_w_n7775_0(.douta(w_n7775_0[0]),.doutb(w_n7775_0[1]),.din(n7775));
	jspl jspl_w_n7779_0(.douta(w_n7779_0[0]),.doutb(w_n7779_0[1]),.din(n7779));
	jspl3 jspl3_w_n7781_0(.douta(w_n7781_0[0]),.doutb(w_n7781_0[1]),.doutc(w_n7781_0[2]),.din(n7781));
	jspl jspl_w_n7782_0(.douta(w_n7782_0[0]),.doutb(w_n7782_0[1]),.din(n7782));
	jspl jspl_w_n7786_0(.douta(w_n7786_0[0]),.doutb(w_n7786_0[1]),.din(n7786));
	jspl3 jspl3_w_n7788_0(.douta(w_n7788_0[0]),.doutb(w_n7788_0[1]),.doutc(w_n7788_0[2]),.din(n7788));
	jspl jspl_w_n7789_0(.douta(w_n7789_0[0]),.doutb(w_n7789_0[1]),.din(n7789));
	jspl jspl_w_n7793_0(.douta(w_n7793_0[0]),.doutb(w_n7793_0[1]),.din(n7793));
	jspl jspl_w_n7794_0(.douta(w_n7794_0[0]),.doutb(w_n7794_0[1]),.din(n7794));
	jspl3 jspl3_w_n7796_0(.douta(w_n7796_0[0]),.doutb(w_n7796_0[1]),.doutc(w_n7796_0[2]),.din(n7796));
	jspl jspl_w_n7797_0(.douta(w_n7797_0[0]),.doutb(w_n7797_0[1]),.din(n7797));
	jspl jspl_w_n7801_0(.douta(w_n7801_0[0]),.doutb(w_n7801_0[1]),.din(n7801));
	jspl jspl_w_n7802_0(.douta(w_n7802_0[0]),.doutb(w_n7802_0[1]),.din(n7802));
	jspl3 jspl3_w_n7804_0(.douta(w_n7804_0[0]),.doutb(w_n7804_0[1]),.doutc(w_n7804_0[2]),.din(n7804));
	jspl jspl_w_n7805_0(.douta(w_n7805_0[0]),.doutb(w_n7805_0[1]),.din(n7805));
	jspl jspl_w_n7809_0(.douta(w_n7809_0[0]),.doutb(w_n7809_0[1]),.din(n7809));
	jspl jspl_w_n7810_0(.douta(w_n7810_0[0]),.doutb(w_n7810_0[1]),.din(n7810));
	jspl3 jspl3_w_n7812_0(.douta(w_n7812_0[0]),.doutb(w_n7812_0[1]),.doutc(w_n7812_0[2]),.din(n7812));
	jspl jspl_w_n7813_0(.douta(w_n7813_0[0]),.doutb(w_n7813_0[1]),.din(n7813));
	jspl3 jspl3_w_n7817_0(.douta(w_n7817_0[0]),.doutb(w_n7817_0[1]),.doutc(w_n7817_0[2]),.din(n7817));
	jspl jspl_w_n7819_0(.douta(w_n7819_0[0]),.doutb(w_n7819_0[1]),.din(n7819));
	jspl3 jspl3_w_n7820_0(.douta(w_n7820_0[0]),.doutb(w_n7820_0[1]),.doutc(w_n7820_0[2]),.din(n7820));
	jspl jspl_w_n7820_1(.douta(w_n7820_1[0]),.doutb(w_n7820_1[1]),.din(w_n7820_0[0]));
	jspl3 jspl3_w_n7821_0(.douta(w_n7821_0[0]),.doutb(w_n7821_0[1]),.doutc(w_n7821_0[2]),.din(n7821));
	jspl jspl_w_n7826_0(.douta(w_n7826_0[0]),.doutb(w_n7826_0[1]),.din(n7826));
	jspl jspl_w_n7827_0(.douta(w_n7827_0[0]),.doutb(w_n7827_0[1]),.din(n7827));
	jspl jspl_w_n7828_0(.douta(w_n7828_0[0]),.doutb(w_n7828_0[1]),.din(n7828));
	jspl jspl_w_n7859_0(.douta(w_n7859_0[0]),.doutb(w_n7859_0[1]),.din(n7859));
	jspl jspl_w_n7882_0(.douta(w_n7882_0[0]),.doutb(w_n7882_0[1]),.din(n7882));
	jspl jspl_w_n7889_0(.douta(w_n7889_0[0]),.doutb(w_n7889_0[1]),.din(n7889));
	jspl jspl_w_n7893_0(.douta(w_n7893_0[0]),.doutb(w_n7893_0[1]),.din(n7893));
	jspl jspl_w_n7897_0(.douta(w_n7897_0[0]),.doutb(w_n7897_0[1]),.din(n7897));
	jspl jspl_w_n7904_0(.douta(w_n7904_0[0]),.doutb(w_n7904_0[1]),.din(n7904));
	jspl jspl_w_n7911_0(.douta(w_n7911_0[0]),.doutb(w_n7911_0[1]),.din(n7911));
	jspl jspl_w_n7918_0(.douta(w_n7918_0[0]),.doutb(w_n7918_0[1]),.din(n7918));
	jspl jspl_w_n7925_0(.douta(w_n7925_0[0]),.doutb(w_n7925_0[1]),.din(n7925));
	jspl jspl_w_n7929_0(.douta(w_n7929_0[0]),.doutb(w_n7929_0[1]),.din(n7929));
	jspl jspl_w_n7933_0(.douta(w_n7933_0[0]),.doutb(w_n7933_0[1]),.din(n7933));
	jspl jspl_w_n7946_0(.douta(w_n7946_0[0]),.doutb(w_n7946_0[1]),.din(n7946));
	jspl jspl_w_n7953_0(.douta(w_n7953_0[0]),.doutb(w_n7953_0[1]),.din(n7953));
	jspl jspl_w_n7960_0(.douta(w_n7960_0[0]),.doutb(w_n7960_0[1]),.din(n7960));
	jspl jspl_w_n7964_0(.douta(w_n7964_0[0]),.doutb(w_n7964_0[1]),.din(n7964));
	jspl jspl_w_n7979_0(.douta(w_n7979_0[0]),.doutb(w_n7979_0[1]),.din(n7979));
	jspl jspl_w_n7980_0(.douta(w_n7980_0[0]),.doutb(w_n7980_0[1]),.din(n7980));
	jspl jspl_w_n7982_0(.douta(w_n7982_0[0]),.doutb(w_n7982_0[1]),.din(n7982));
	jspl jspl_w_n7984_0(.douta(w_n7984_0[0]),.doutb(w_n7984_0[1]),.din(n7984));
	jspl jspl_w_n7985_0(.douta(w_n7985_0[0]),.doutb(w_n7985_0[1]),.din(n7985));
	jspl jspl_w_n7987_0(.douta(w_n7987_0[0]),.doutb(w_n7987_0[1]),.din(n7987));
	jspl jspl_w_n7989_0(.douta(w_n7989_0[0]),.doutb(w_n7989_0[1]),.din(n7989));
	jspl jspl_w_n7990_0(.douta(w_n7990_0[0]),.doutb(w_n7990_0[1]),.din(n7990));
	jspl3 jspl3_w_n7991_0(.douta(w_n7991_0[0]),.doutb(w_n7991_0[1]),.doutc(w_n7991_0[2]),.din(n7991));
	jspl3 jspl3_w_n7991_1(.douta(w_n7991_1[0]),.doutb(w_n7991_1[1]),.doutc(w_n7991_1[2]),.din(w_n7991_0[0]));
	jspl jspl_w_n7992_0(.douta(w_n7992_0[0]),.doutb(w_n7992_0[1]),.din(n7992));
	jspl3 jspl3_w_n7993_0(.douta(w_n7993_0[0]),.doutb(w_n7993_0[1]),.doutc(w_n7993_0[2]),.din(n7993));
	jspl jspl_w_n7994_0(.douta(w_n7994_0[0]),.doutb(w_n7994_0[1]),.din(n7994));
	jspl jspl_w_n8002_0(.douta(w_n8002_0[0]),.doutb(w_n8002_0[1]),.din(n8002));
	jspl3 jspl3_w_n8003_0(.douta(w_n8003_0[0]),.doutb(w_n8003_0[1]),.doutc(w_n8003_0[2]),.din(n8003));
	jspl3 jspl3_w_n8003_1(.douta(w_n8003_1[0]),.doutb(w_n8003_1[1]),.doutc(w_n8003_1[2]),.din(w_n8003_0[0]));
	jspl3 jspl3_w_n8003_2(.douta(w_n8003_2[0]),.doutb(w_n8003_2[1]),.doutc(w_n8003_2[2]),.din(w_n8003_0[1]));
	jspl3 jspl3_w_n8003_3(.douta(w_n8003_3[0]),.doutb(w_n8003_3[1]),.doutc(w_n8003_3[2]),.din(w_n8003_0[2]));
	jspl3 jspl3_w_n8003_4(.douta(w_n8003_4[0]),.doutb(w_n8003_4[1]),.doutc(w_n8003_4[2]),.din(w_n8003_1[0]));
	jspl3 jspl3_w_n8003_5(.douta(w_n8003_5[0]),.doutb(w_n8003_5[1]),.doutc(w_n8003_5[2]),.din(w_n8003_1[1]));
	jspl3 jspl3_w_n8003_6(.douta(w_n8003_6[0]),.doutb(w_n8003_6[1]),.doutc(w_n8003_6[2]),.din(w_n8003_1[2]));
	jspl3 jspl3_w_n8003_7(.douta(w_n8003_7[0]),.doutb(w_n8003_7[1]),.doutc(w_n8003_7[2]),.din(w_n8003_2[0]));
	jspl3 jspl3_w_n8003_8(.douta(w_n8003_8[0]),.doutb(w_n8003_8[1]),.doutc(w_n8003_8[2]),.din(w_n8003_2[1]));
	jspl3 jspl3_w_n8003_9(.douta(w_n8003_9[0]),.doutb(w_n8003_9[1]),.doutc(w_n8003_9[2]),.din(w_n8003_2[2]));
	jspl3 jspl3_w_n8003_10(.douta(w_n8003_10[0]),.doutb(w_n8003_10[1]),.doutc(w_n8003_10[2]),.din(w_n8003_3[0]));
	jspl3 jspl3_w_n8003_11(.douta(w_n8003_11[0]),.doutb(w_n8003_11[1]),.doutc(w_n8003_11[2]),.din(w_n8003_3[1]));
	jspl3 jspl3_w_n8003_12(.douta(w_n8003_12[0]),.doutb(w_n8003_12[1]),.doutc(w_n8003_12[2]),.din(w_n8003_3[2]));
	jspl3 jspl3_w_n8003_13(.douta(w_n8003_13[0]),.doutb(w_n8003_13[1]),.doutc(w_n8003_13[2]),.din(w_n8003_4[0]));
	jspl3 jspl3_w_n8003_14(.douta(w_n8003_14[0]),.doutb(w_n8003_14[1]),.doutc(w_n8003_14[2]),.din(w_n8003_4[1]));
	jspl3 jspl3_w_n8003_15(.douta(w_n8003_15[0]),.doutb(w_n8003_15[1]),.doutc(w_n8003_15[2]),.din(w_n8003_4[2]));
	jspl3 jspl3_w_n8003_16(.douta(w_n8003_16[0]),.doutb(w_n8003_16[1]),.doutc(w_n8003_16[2]),.din(w_n8003_5[0]));
	jspl3 jspl3_w_n8003_17(.douta(w_n8003_17[0]),.doutb(w_n8003_17[1]),.doutc(w_n8003_17[2]),.din(w_n8003_5[1]));
	jspl3 jspl3_w_n8003_18(.douta(w_n8003_18[0]),.doutb(w_n8003_18[1]),.doutc(w_n8003_18[2]),.din(w_n8003_5[2]));
	jspl3 jspl3_w_n8003_19(.douta(w_n8003_19[0]),.doutb(w_n8003_19[1]),.doutc(w_n8003_19[2]),.din(w_n8003_6[0]));
	jspl3 jspl3_w_n8003_20(.douta(w_n8003_20[0]),.doutb(w_n8003_20[1]),.doutc(w_n8003_20[2]),.din(w_n8003_6[1]));
	jspl3 jspl3_w_n8003_21(.douta(w_n8003_21[0]),.doutb(w_n8003_21[1]),.doutc(w_n8003_21[2]),.din(w_n8003_6[2]));
	jspl3 jspl3_w_n8003_22(.douta(w_n8003_22[0]),.doutb(w_n8003_22[1]),.doutc(w_n8003_22[2]),.din(w_n8003_7[0]));
	jspl3 jspl3_w_n8003_23(.douta(w_n8003_23[0]),.doutb(w_n8003_23[1]),.doutc(w_n8003_23[2]),.din(w_n8003_7[1]));
	jspl3 jspl3_w_n8003_24(.douta(w_n8003_24[0]),.doutb(w_n8003_24[1]),.doutc(w_n8003_24[2]),.din(w_n8003_7[2]));
	jspl3 jspl3_w_n8003_25(.douta(w_n8003_25[0]),.doutb(w_n8003_25[1]),.doutc(w_n8003_25[2]),.din(w_n8003_8[0]));
	jspl3 jspl3_w_n8003_26(.douta(w_n8003_26[0]),.doutb(w_n8003_26[1]),.doutc(w_n8003_26[2]),.din(w_n8003_8[1]));
	jspl3 jspl3_w_n8003_27(.douta(w_n8003_27[0]),.doutb(w_n8003_27[1]),.doutc(w_n8003_27[2]),.din(w_n8003_8[2]));
	jspl3 jspl3_w_n8003_28(.douta(w_n8003_28[0]),.doutb(w_n8003_28[1]),.doutc(w_n8003_28[2]),.din(w_n8003_9[0]));
	jspl3 jspl3_w_n8003_29(.douta(w_n8003_29[0]),.doutb(w_n8003_29[1]),.doutc(w_n8003_29[2]),.din(w_n8003_9[1]));
	jspl3 jspl3_w_n8003_30(.douta(w_n8003_30[0]),.doutb(w_n8003_30[1]),.doutc(w_n8003_30[2]),.din(w_n8003_9[2]));
	jspl3 jspl3_w_n8003_31(.douta(w_n8003_31[0]),.doutb(w_n8003_31[1]),.doutc(w_n8003_31[2]),.din(w_n8003_10[0]));
	jspl3 jspl3_w_n8003_32(.douta(w_n8003_32[0]),.doutb(w_n8003_32[1]),.doutc(w_n8003_32[2]),.din(w_n8003_10[1]));
	jspl3 jspl3_w_n8003_33(.douta(w_n8003_33[0]),.doutb(w_n8003_33[1]),.doutc(w_n8003_33[2]),.din(w_n8003_10[2]));
	jspl3 jspl3_w_n8003_34(.douta(w_n8003_34[0]),.doutb(w_n8003_34[1]),.doutc(w_n8003_34[2]),.din(w_n8003_11[0]));
	jspl3 jspl3_w_n8003_35(.douta(w_n8003_35[0]),.doutb(w_n8003_35[1]),.doutc(w_n8003_35[2]),.din(w_n8003_11[1]));
	jspl3 jspl3_w_n8003_36(.douta(w_n8003_36[0]),.doutb(w_n8003_36[1]),.doutc(w_n8003_36[2]),.din(w_n8003_11[2]));
	jspl3 jspl3_w_n8003_37(.douta(w_n8003_37[0]),.doutb(w_n8003_37[1]),.doutc(w_n8003_37[2]),.din(w_n8003_12[0]));
	jspl3 jspl3_w_n8003_38(.douta(w_n8003_38[0]),.doutb(w_n8003_38[1]),.doutc(w_n8003_38[2]),.din(w_n8003_12[1]));
	jspl3 jspl3_w_n8003_39(.douta(w_n8003_39[0]),.doutb(w_n8003_39[1]),.doutc(w_n8003_39[2]),.din(w_n8003_12[2]));
	jspl3 jspl3_w_n8003_40(.douta(w_n8003_40[0]),.doutb(w_n8003_40[1]),.doutc(w_n8003_40[2]),.din(w_n8003_13[0]));
	jspl3 jspl3_w_n8003_41(.douta(w_n8003_41[0]),.doutb(w_n8003_41[1]),.doutc(w_n8003_41[2]),.din(w_n8003_13[1]));
	jspl3 jspl3_w_n8003_42(.douta(w_n8003_42[0]),.doutb(w_n8003_42[1]),.doutc(w_n8003_42[2]),.din(w_n8003_13[2]));
	jspl3 jspl3_w_n8003_43(.douta(w_n8003_43[0]),.doutb(w_n8003_43[1]),.doutc(w_n8003_43[2]),.din(w_n8003_14[0]));
	jspl3 jspl3_w_n8003_44(.douta(w_n8003_44[0]),.doutb(w_n8003_44[1]),.doutc(w_n8003_44[2]),.din(w_n8003_14[1]));
	jspl3 jspl3_w_n8003_45(.douta(w_n8003_45[0]),.doutb(w_n8003_45[1]),.doutc(w_n8003_45[2]),.din(w_n8003_14[2]));
	jspl3 jspl3_w_n8003_46(.douta(w_n8003_46[0]),.doutb(w_n8003_46[1]),.doutc(w_n8003_46[2]),.din(w_n8003_15[0]));
	jspl3 jspl3_w_n8003_47(.douta(w_n8003_47[0]),.doutb(w_n8003_47[1]),.doutc(w_n8003_47[2]),.din(w_n8003_15[1]));
	jspl3 jspl3_w_n8003_48(.douta(w_n8003_48[0]),.doutb(w_n8003_48[1]),.doutc(w_n8003_48[2]),.din(w_n8003_15[2]));
	jspl3 jspl3_w_n8003_49(.douta(w_n8003_49[0]),.doutb(w_n8003_49[1]),.doutc(w_n8003_49[2]),.din(w_n8003_16[0]));
	jspl3 jspl3_w_n8003_50(.douta(w_n8003_50[0]),.doutb(w_n8003_50[1]),.doutc(w_n8003_50[2]),.din(w_n8003_16[1]));
	jspl3 jspl3_w_n8003_51(.douta(w_n8003_51[0]),.doutb(w_n8003_51[1]),.doutc(w_n8003_51[2]),.din(w_n8003_16[2]));
	jspl jspl_w_n8003_52(.douta(w_n8003_52[0]),.doutb(w_n8003_52[1]),.din(w_n8003_17[0]));
	jspl3 jspl3_w_n8005_0(.douta(w_n8005_0[0]),.doutb(w_n8005_0[1]),.doutc(w_n8005_0[2]),.din(n8005));
	jspl jspl_w_n8006_0(.douta(w_n8006_0[0]),.doutb(w_n8006_0[1]),.din(n8006));
	jspl3 jspl3_w_n8013_0(.douta(w_n8013_0[0]),.doutb(w_n8013_0[1]),.doutc(w_n8013_0[2]),.din(n8013));
	jspl jspl_w_n8014_0(.douta(w_n8014_0[0]),.doutb(w_n8014_0[1]),.din(n8014));
	jspl jspl_w_n8017_0(.douta(w_n8017_0[0]),.doutb(w_n8017_0[1]),.din(n8017));
	jspl3 jspl3_w_n8022_0(.douta(w_n8022_0[0]),.doutb(w_n8022_0[1]),.doutc(w_n8022_0[2]),.din(n8022));
	jspl3 jspl3_w_n8024_0(.douta(w_n8024_0[0]),.doutb(w_n8024_0[1]),.doutc(w_n8024_0[2]),.din(n8024));
	jspl jspl_w_n8025_0(.douta(w_n8025_0[0]),.doutb(w_n8025_0[1]),.din(n8025));
	jspl3 jspl3_w_n8029_0(.douta(w_n8029_0[0]),.doutb(w_n8029_0[1]),.doutc(w_n8029_0[2]),.din(n8029));
	jspl3 jspl3_w_n8031_0(.douta(w_n8031_0[0]),.doutb(w_n8031_0[1]),.doutc(w_n8031_0[2]),.din(n8031));
	jspl jspl_w_n8032_0(.douta(w_n8032_0[0]),.doutb(w_n8032_0[1]),.din(n8032));
	jspl3 jspl3_w_n8036_0(.douta(w_n8036_0[0]),.doutb(w_n8036_0[1]),.doutc(w_n8036_0[2]),.din(n8036));
	jspl3 jspl3_w_n8038_0(.douta(w_n8038_0[0]),.doutb(w_n8038_0[1]),.doutc(w_n8038_0[2]),.din(n8038));
	jspl jspl_w_n8039_0(.douta(w_n8039_0[0]),.doutb(w_n8039_0[1]),.din(n8039));
	jspl3 jspl3_w_n8042_0(.douta(w_n8042_0[0]),.doutb(w_n8042_0[1]),.doutc(w_n8042_0[2]),.din(n8042));
	jspl3 jspl3_w_n8046_0(.douta(w_n8046_0[0]),.doutb(w_n8046_0[1]),.doutc(w_n8046_0[2]),.din(n8046));
	jspl jspl_w_n8047_0(.douta(w_n8047_0[0]),.doutb(w_n8047_0[1]),.din(n8047));
	jspl3 jspl3_w_n8051_0(.douta(w_n8051_0[0]),.doutb(w_n8051_0[1]),.doutc(w_n8051_0[2]),.din(n8051));
	jspl3 jspl3_w_n8053_0(.douta(w_n8053_0[0]),.doutb(w_n8053_0[1]),.doutc(w_n8053_0[2]),.din(n8053));
	jspl jspl_w_n8054_0(.douta(w_n8054_0[0]),.doutb(w_n8054_0[1]),.din(n8054));
	jspl3 jspl3_w_n8058_0(.douta(w_n8058_0[0]),.doutb(w_n8058_0[1]),.doutc(w_n8058_0[2]),.din(n8058));
	jspl3 jspl3_w_n8061_0(.douta(w_n8061_0[0]),.doutb(w_n8061_0[1]),.doutc(w_n8061_0[2]),.din(n8061));
	jspl jspl_w_n8062_0(.douta(w_n8062_0[0]),.doutb(w_n8062_0[1]),.din(n8062));
	jspl3 jspl3_w_n8066_0(.douta(w_n8066_0[0]),.doutb(w_n8066_0[1]),.doutc(w_n8066_0[2]),.din(n8066));
	jspl3 jspl3_w_n8068_0(.douta(w_n8068_0[0]),.doutb(w_n8068_0[1]),.doutc(w_n8068_0[2]),.din(n8068));
	jspl jspl_w_n8069_0(.douta(w_n8069_0[0]),.doutb(w_n8069_0[1]),.din(n8069));
	jspl3 jspl3_w_n8073_0(.douta(w_n8073_0[0]),.doutb(w_n8073_0[1]),.doutc(w_n8073_0[2]),.din(n8073));
	jspl3 jspl3_w_n8076_0(.douta(w_n8076_0[0]),.doutb(w_n8076_0[1]),.doutc(w_n8076_0[2]),.din(n8076));
	jspl jspl_w_n8077_0(.douta(w_n8077_0[0]),.doutb(w_n8077_0[1]),.din(n8077));
	jspl3 jspl3_w_n8081_0(.douta(w_n8081_0[0]),.doutb(w_n8081_0[1]),.doutc(w_n8081_0[2]),.din(n8081));
	jspl3 jspl3_w_n8084_0(.douta(w_n8084_0[0]),.doutb(w_n8084_0[1]),.doutc(w_n8084_0[2]),.din(n8084));
	jspl jspl_w_n8085_0(.douta(w_n8085_0[0]),.doutb(w_n8085_0[1]),.din(n8085));
	jspl3 jspl3_w_n8089_0(.douta(w_n8089_0[0]),.doutb(w_n8089_0[1]),.doutc(w_n8089_0[2]),.din(n8089));
	jspl3 jspl3_w_n8092_0(.douta(w_n8092_0[0]),.doutb(w_n8092_0[1]),.doutc(w_n8092_0[2]),.din(n8092));
	jspl jspl_w_n8093_0(.douta(w_n8093_0[0]),.doutb(w_n8093_0[1]),.din(n8093));
	jspl3 jspl3_w_n8097_0(.douta(w_n8097_0[0]),.doutb(w_n8097_0[1]),.doutc(w_n8097_0[2]),.din(n8097));
	jspl3 jspl3_w_n8099_0(.douta(w_n8099_0[0]),.doutb(w_n8099_0[1]),.doutc(w_n8099_0[2]),.din(n8099));
	jspl jspl_w_n8100_0(.douta(w_n8100_0[0]),.doutb(w_n8100_0[1]),.din(n8100));
	jspl3 jspl3_w_n8104_0(.douta(w_n8104_0[0]),.doutb(w_n8104_0[1]),.doutc(w_n8104_0[2]),.din(n8104));
	jspl3 jspl3_w_n8107_0(.douta(w_n8107_0[0]),.doutb(w_n8107_0[1]),.doutc(w_n8107_0[2]),.din(n8107));
	jspl jspl_w_n8108_0(.douta(w_n8108_0[0]),.doutb(w_n8108_0[1]),.din(n8108));
	jspl3 jspl3_w_n8112_0(.douta(w_n8112_0[0]),.doutb(w_n8112_0[1]),.doutc(w_n8112_0[2]),.din(n8112));
	jspl3 jspl3_w_n8114_0(.douta(w_n8114_0[0]),.doutb(w_n8114_0[1]),.doutc(w_n8114_0[2]),.din(n8114));
	jspl jspl_w_n8115_0(.douta(w_n8115_0[0]),.doutb(w_n8115_0[1]),.din(n8115));
	jspl3 jspl3_w_n8119_0(.douta(w_n8119_0[0]),.doutb(w_n8119_0[1]),.doutc(w_n8119_0[2]),.din(n8119));
	jspl3 jspl3_w_n8122_0(.douta(w_n8122_0[0]),.doutb(w_n8122_0[1]),.doutc(w_n8122_0[2]),.din(n8122));
	jspl jspl_w_n8123_0(.douta(w_n8123_0[0]),.doutb(w_n8123_0[1]),.din(n8123));
	jspl3 jspl3_w_n8127_0(.douta(w_n8127_0[0]),.doutb(w_n8127_0[1]),.doutc(w_n8127_0[2]),.din(n8127));
	jspl3 jspl3_w_n8129_0(.douta(w_n8129_0[0]),.doutb(w_n8129_0[1]),.doutc(w_n8129_0[2]),.din(n8129));
	jspl jspl_w_n8130_0(.douta(w_n8130_0[0]),.doutb(w_n8130_0[1]),.din(n8130));
	jspl3 jspl3_w_n8134_0(.douta(w_n8134_0[0]),.doutb(w_n8134_0[1]),.doutc(w_n8134_0[2]),.din(n8134));
	jspl3 jspl3_w_n8137_0(.douta(w_n8137_0[0]),.doutb(w_n8137_0[1]),.doutc(w_n8137_0[2]),.din(n8137));
	jspl jspl_w_n8138_0(.douta(w_n8138_0[0]),.doutb(w_n8138_0[1]),.din(n8138));
	jspl3 jspl3_w_n8142_0(.douta(w_n8142_0[0]),.doutb(w_n8142_0[1]),.doutc(w_n8142_0[2]),.din(n8142));
	jspl3 jspl3_w_n8144_0(.douta(w_n8144_0[0]),.doutb(w_n8144_0[1]),.doutc(w_n8144_0[2]),.din(n8144));
	jspl jspl_w_n8145_0(.douta(w_n8145_0[0]),.doutb(w_n8145_0[1]),.din(n8145));
	jspl3 jspl3_w_n8149_0(.douta(w_n8149_0[0]),.doutb(w_n8149_0[1]),.doutc(w_n8149_0[2]),.din(n8149));
	jspl3 jspl3_w_n8152_0(.douta(w_n8152_0[0]),.doutb(w_n8152_0[1]),.doutc(w_n8152_0[2]),.din(n8152));
	jspl jspl_w_n8153_0(.douta(w_n8153_0[0]),.doutb(w_n8153_0[1]),.din(n8153));
	jspl3 jspl3_w_n8157_0(.douta(w_n8157_0[0]),.doutb(w_n8157_0[1]),.doutc(w_n8157_0[2]),.din(n8157));
	jspl3 jspl3_w_n8160_0(.douta(w_n8160_0[0]),.doutb(w_n8160_0[1]),.doutc(w_n8160_0[2]),.din(n8160));
	jspl jspl_w_n8161_0(.douta(w_n8161_0[0]),.doutb(w_n8161_0[1]),.din(n8161));
	jspl3 jspl3_w_n8165_0(.douta(w_n8165_0[0]),.doutb(w_n8165_0[1]),.doutc(w_n8165_0[2]),.din(n8165));
	jspl3 jspl3_w_n8168_0(.douta(w_n8168_0[0]),.doutb(w_n8168_0[1]),.doutc(w_n8168_0[2]),.din(n8168));
	jspl jspl_w_n8169_0(.douta(w_n8169_0[0]),.doutb(w_n8169_0[1]),.din(n8169));
	jspl3 jspl3_w_n8173_0(.douta(w_n8173_0[0]),.doutb(w_n8173_0[1]),.doutc(w_n8173_0[2]),.din(n8173));
	jspl3 jspl3_w_n8175_0(.douta(w_n8175_0[0]),.doutb(w_n8175_0[1]),.doutc(w_n8175_0[2]),.din(n8175));
	jspl jspl_w_n8176_0(.douta(w_n8176_0[0]),.doutb(w_n8176_0[1]),.din(n8176));
	jspl3 jspl3_w_n8180_0(.douta(w_n8180_0[0]),.doutb(w_n8180_0[1]),.doutc(w_n8180_0[2]),.din(n8180));
	jspl3 jspl3_w_n8182_0(.douta(w_n8182_0[0]),.doutb(w_n8182_0[1]),.doutc(w_n8182_0[2]),.din(n8182));
	jspl jspl_w_n8183_0(.douta(w_n8183_0[0]),.doutb(w_n8183_0[1]),.din(n8183));
	jspl3 jspl3_w_n8187_0(.douta(w_n8187_0[0]),.doutb(w_n8187_0[1]),.doutc(w_n8187_0[2]),.din(n8187));
	jspl3 jspl3_w_n8189_0(.douta(w_n8189_0[0]),.doutb(w_n8189_0[1]),.doutc(w_n8189_0[2]),.din(n8189));
	jspl jspl_w_n8190_0(.douta(w_n8190_0[0]),.doutb(w_n8190_0[1]),.din(n8190));
	jspl3 jspl3_w_n8194_0(.douta(w_n8194_0[0]),.doutb(w_n8194_0[1]),.doutc(w_n8194_0[2]),.din(n8194));
	jspl3 jspl3_w_n8197_0(.douta(w_n8197_0[0]),.doutb(w_n8197_0[1]),.doutc(w_n8197_0[2]),.din(n8197));
	jspl jspl_w_n8198_0(.douta(w_n8198_0[0]),.doutb(w_n8198_0[1]),.din(n8198));
	jspl3 jspl3_w_n8202_0(.douta(w_n8202_0[0]),.doutb(w_n8202_0[1]),.doutc(w_n8202_0[2]),.din(n8202));
	jspl3 jspl3_w_n8204_0(.douta(w_n8204_0[0]),.doutb(w_n8204_0[1]),.doutc(w_n8204_0[2]),.din(n8204));
	jspl jspl_w_n8205_0(.douta(w_n8205_0[0]),.doutb(w_n8205_0[1]),.din(n8205));
	jspl3 jspl3_w_n8209_0(.douta(w_n8209_0[0]),.doutb(w_n8209_0[1]),.doutc(w_n8209_0[2]),.din(n8209));
	jspl3 jspl3_w_n8212_0(.douta(w_n8212_0[0]),.doutb(w_n8212_0[1]),.doutc(w_n8212_0[2]),.din(n8212));
	jspl jspl_w_n8213_0(.douta(w_n8213_0[0]),.doutb(w_n8213_0[1]),.din(n8213));
	jspl3 jspl3_w_n8217_0(.douta(w_n8217_0[0]),.doutb(w_n8217_0[1]),.doutc(w_n8217_0[2]),.din(n8217));
	jspl3 jspl3_w_n8219_0(.douta(w_n8219_0[0]),.doutb(w_n8219_0[1]),.doutc(w_n8219_0[2]),.din(n8219));
	jspl jspl_w_n8220_0(.douta(w_n8220_0[0]),.doutb(w_n8220_0[1]),.din(n8220));
	jspl3 jspl3_w_n8224_0(.douta(w_n8224_0[0]),.doutb(w_n8224_0[1]),.doutc(w_n8224_0[2]),.din(n8224));
	jspl3 jspl3_w_n8227_0(.douta(w_n8227_0[0]),.doutb(w_n8227_0[1]),.doutc(w_n8227_0[2]),.din(n8227));
	jspl jspl_w_n8228_0(.douta(w_n8228_0[0]),.doutb(w_n8228_0[1]),.din(n8228));
	jspl3 jspl3_w_n8232_0(.douta(w_n8232_0[0]),.doutb(w_n8232_0[1]),.doutc(w_n8232_0[2]),.din(n8232));
	jspl3 jspl3_w_n8235_0(.douta(w_n8235_0[0]),.doutb(w_n8235_0[1]),.doutc(w_n8235_0[2]),.din(n8235));
	jspl jspl_w_n8236_0(.douta(w_n8236_0[0]),.doutb(w_n8236_0[1]),.din(n8236));
	jspl3 jspl3_w_n8240_0(.douta(w_n8240_0[0]),.doutb(w_n8240_0[1]),.doutc(w_n8240_0[2]),.din(n8240));
	jspl3 jspl3_w_n8242_0(.douta(w_n8242_0[0]),.doutb(w_n8242_0[1]),.doutc(w_n8242_0[2]),.din(n8242));
	jspl jspl_w_n8243_0(.douta(w_n8243_0[0]),.doutb(w_n8243_0[1]),.din(n8243));
	jspl3 jspl3_w_n8247_0(.douta(w_n8247_0[0]),.doutb(w_n8247_0[1]),.doutc(w_n8247_0[2]),.din(n8247));
	jspl3 jspl3_w_n8249_0(.douta(w_n8249_0[0]),.doutb(w_n8249_0[1]),.doutc(w_n8249_0[2]),.din(n8249));
	jspl jspl_w_n8250_0(.douta(w_n8250_0[0]),.doutb(w_n8250_0[1]),.din(n8250));
	jspl jspl_w_n8254_0(.douta(w_n8254_0[0]),.doutb(w_n8254_0[1]),.din(n8254));
	jspl3 jspl3_w_n8256_0(.douta(w_n8256_0[0]),.doutb(w_n8256_0[1]),.doutc(w_n8256_0[2]),.din(n8256));
	jspl3 jspl3_w_n8259_0(.douta(w_n8259_0[0]),.doutb(w_n8259_0[1]),.doutc(w_n8259_0[2]),.din(n8259));
	jspl jspl_w_n8260_0(.douta(w_n8260_0[0]),.doutb(w_n8260_0[1]),.din(n8260));
	jspl jspl_w_n8263_0(.douta(w_n8263_0[0]),.doutb(w_n8263_0[1]),.din(n8263));
	jspl3 jspl3_w_n8265_0(.douta(w_n8265_0[0]),.doutb(w_n8265_0[1]),.doutc(w_n8265_0[2]),.din(n8265));
	jspl jspl_w_n8265_1(.douta(w_n8265_1[0]),.doutb(w_n8265_1[1]),.din(w_n8265_0[0]));
	jspl jspl_w_n8270_0(.douta(w_n8270_0[0]),.doutb(w_n8270_0[1]),.din(n8270));
	jspl jspl_w_n8272_0(.douta(w_n8272_0[0]),.doutb(w_n8272_0[1]),.din(n8272));
	jspl jspl_w_n8274_0(.douta(w_n8274_0[0]),.doutb(w_n8274_0[1]),.din(n8274));
	jspl3 jspl3_w_n8277_0(.douta(w_n8277_0[0]),.doutb(w_n8277_0[1]),.doutc(w_n8277_0[2]),.din(n8277));
	jspl3 jspl3_w_n8279_0(.douta(w_n8279_0[0]),.doutb(w_n8279_0[1]),.doutc(w_n8279_0[2]),.din(n8279));
	jspl jspl_w_n8279_1(.douta(w_n8279_1[0]),.doutb(w_n8279_1[1]),.din(w_n8279_0[0]));
	jspl jspl_w_n8280_0(.douta(w_n8280_0[0]),.doutb(w_n8280_0[1]),.din(n8280));
	jspl3 jspl3_w_n8281_0(.douta(w_n8281_0[0]),.doutb(w_n8281_0[1]),.doutc(w_n8281_0[2]),.din(n8281));
	jspl jspl_w_n8282_0(.douta(w_n8282_0[0]),.doutb(w_n8282_0[1]),.din(n8282));
	jspl3 jspl3_w_n8283_0(.douta(w_n8283_0[0]),.doutb(w_n8283_0[1]),.doutc(w_n8283_0[2]),.din(n8283));
	jspl jspl_w_n8284_0(.douta(w_n8284_0[0]),.doutb(w_n8284_0[1]),.din(n8284));
	jspl jspl_w_n8328_0(.douta(w_n8328_0[0]),.doutb(w_n8328_0[1]),.din(n8328));
	jspl jspl_w_n8444_0(.douta(w_n8444_0[0]),.doutb(w_n8444_0[1]),.din(n8444));
	jspl3 jspl3_w_n8449_0(.douta(w_n8449_0[0]),.doutb(w_n8449_0[1]),.doutc(w_n8449_0[2]),.din(n8449));
	jspl3 jspl3_w_n8449_1(.douta(w_n8449_1[0]),.doutb(w_n8449_1[1]),.doutc(w_n8449_1[2]),.din(w_n8449_0[0]));
	jspl3 jspl3_w_n8449_2(.douta(w_n8449_2[0]),.doutb(w_n8449_2[1]),.doutc(w_n8449_2[2]),.din(w_n8449_0[1]));
	jspl3 jspl3_w_n8449_3(.douta(w_n8449_3[0]),.doutb(w_n8449_3[1]),.doutc(w_n8449_3[2]),.din(w_n8449_0[2]));
	jspl3 jspl3_w_n8449_4(.douta(w_n8449_4[0]),.doutb(w_n8449_4[1]),.doutc(w_n8449_4[2]),.din(w_n8449_1[0]));
	jspl3 jspl3_w_n8449_5(.douta(w_n8449_5[0]),.doutb(w_n8449_5[1]),.doutc(w_n8449_5[2]),.din(w_n8449_1[1]));
	jspl3 jspl3_w_n8449_6(.douta(w_n8449_6[0]),.doutb(w_n8449_6[1]),.doutc(w_n8449_6[2]),.din(w_n8449_1[2]));
	jspl3 jspl3_w_n8449_7(.douta(w_n8449_7[0]),.doutb(w_n8449_7[1]),.doutc(w_n8449_7[2]),.din(w_n8449_2[0]));
	jspl3 jspl3_w_n8449_8(.douta(w_n8449_8[0]),.doutb(w_n8449_8[1]),.doutc(w_n8449_8[2]),.din(w_n8449_2[1]));
	jspl3 jspl3_w_n8449_9(.douta(w_n8449_9[0]),.doutb(w_n8449_9[1]),.doutc(w_n8449_9[2]),.din(w_n8449_2[2]));
	jspl3 jspl3_w_n8449_10(.douta(w_n8449_10[0]),.doutb(w_n8449_10[1]),.doutc(w_n8449_10[2]),.din(w_n8449_3[0]));
	jspl3 jspl3_w_n8449_11(.douta(w_n8449_11[0]),.doutb(w_n8449_11[1]),.doutc(w_n8449_11[2]),.din(w_n8449_3[1]));
	jspl3 jspl3_w_n8449_12(.douta(w_n8449_12[0]),.doutb(w_n8449_12[1]),.doutc(w_n8449_12[2]),.din(w_n8449_3[2]));
	jspl3 jspl3_w_n8449_13(.douta(w_n8449_13[0]),.doutb(w_n8449_13[1]),.doutc(w_n8449_13[2]),.din(w_n8449_4[0]));
	jspl3 jspl3_w_n8449_14(.douta(w_n8449_14[0]),.doutb(w_n8449_14[1]),.doutc(w_n8449_14[2]),.din(w_n8449_4[1]));
	jspl3 jspl3_w_n8449_15(.douta(w_n8449_15[0]),.doutb(w_n8449_15[1]),.doutc(w_n8449_15[2]),.din(w_n8449_4[2]));
	jspl3 jspl3_w_n8449_16(.douta(w_n8449_16[0]),.doutb(w_n8449_16[1]),.doutc(w_n8449_16[2]),.din(w_n8449_5[0]));
	jspl3 jspl3_w_n8449_17(.douta(w_n8449_17[0]),.doutb(w_n8449_17[1]),.doutc(w_n8449_17[2]),.din(w_n8449_5[1]));
	jspl3 jspl3_w_n8449_18(.douta(w_n8449_18[0]),.doutb(w_n8449_18[1]),.doutc(w_n8449_18[2]),.din(w_n8449_5[2]));
	jspl3 jspl3_w_n8449_19(.douta(w_n8449_19[0]),.doutb(w_n8449_19[1]),.doutc(w_n8449_19[2]),.din(w_n8449_6[0]));
	jspl3 jspl3_w_n8449_20(.douta(w_n8449_20[0]),.doutb(w_n8449_20[1]),.doutc(w_n8449_20[2]),.din(w_n8449_6[1]));
	jspl3 jspl3_w_n8449_21(.douta(w_n8449_21[0]),.doutb(w_n8449_21[1]),.doutc(w_n8449_21[2]),.din(w_n8449_6[2]));
	jspl3 jspl3_w_n8449_22(.douta(w_n8449_22[0]),.doutb(w_n8449_22[1]),.doutc(w_n8449_22[2]),.din(w_n8449_7[0]));
	jspl3 jspl3_w_n8449_23(.douta(w_n8449_23[0]),.doutb(w_n8449_23[1]),.doutc(w_n8449_23[2]),.din(w_n8449_7[1]));
	jspl3 jspl3_w_n8449_24(.douta(w_n8449_24[0]),.doutb(w_n8449_24[1]),.doutc(w_n8449_24[2]),.din(w_n8449_7[2]));
	jspl3 jspl3_w_n8449_25(.douta(w_n8449_25[0]),.doutb(w_n8449_25[1]),.doutc(w_n8449_25[2]),.din(w_n8449_8[0]));
	jspl3 jspl3_w_n8449_26(.douta(w_n8449_26[0]),.doutb(w_n8449_26[1]),.doutc(w_n8449_26[2]),.din(w_n8449_8[1]));
	jspl3 jspl3_w_n8449_27(.douta(w_n8449_27[0]),.doutb(w_n8449_27[1]),.doutc(w_n8449_27[2]),.din(w_n8449_8[2]));
	jspl3 jspl3_w_n8449_28(.douta(w_n8449_28[0]),.doutb(w_n8449_28[1]),.doutc(w_n8449_28[2]),.din(w_n8449_9[0]));
	jspl3 jspl3_w_n8449_29(.douta(w_n8449_29[0]),.doutb(w_n8449_29[1]),.doutc(w_n8449_29[2]),.din(w_n8449_9[1]));
	jspl3 jspl3_w_n8449_30(.douta(w_n8449_30[0]),.doutb(w_n8449_30[1]),.doutc(w_n8449_30[2]),.din(w_n8449_9[2]));
	jspl3 jspl3_w_n8449_31(.douta(w_n8449_31[0]),.doutb(w_n8449_31[1]),.doutc(w_n8449_31[2]),.din(w_n8449_10[0]));
	jspl3 jspl3_w_n8449_32(.douta(w_n8449_32[0]),.doutb(w_n8449_32[1]),.doutc(w_n8449_32[2]),.din(w_n8449_10[1]));
	jspl3 jspl3_w_n8449_33(.douta(w_n8449_33[0]),.doutb(w_n8449_33[1]),.doutc(w_n8449_33[2]),.din(w_n8449_10[2]));
	jspl3 jspl3_w_n8449_34(.douta(w_n8449_34[0]),.doutb(w_n8449_34[1]),.doutc(w_n8449_34[2]),.din(w_n8449_11[0]));
	jspl jspl_w_n8449_35(.douta(w_n8449_35[0]),.doutb(w_n8449_35[1]),.din(w_n8449_11[1]));
	jspl jspl_w_n8450_0(.douta(w_n8450_0[0]),.doutb(w_n8450_0[1]),.din(n8450));
	jspl3 jspl3_w_n8453_0(.douta(w_n8453_0[0]),.doutb(w_n8453_0[1]),.doutc(w_n8453_0[2]),.din(n8453));
	jspl jspl_w_n8454_0(.douta(w_n8454_0[0]),.doutb(w_n8454_0[1]),.din(n8454));
	jspl jspl_w_n8460_0(.douta(w_n8460_0[0]),.doutb(w_n8460_0[1]),.din(n8460));
	jspl jspl_w_n8461_0(.douta(w_n8461_0[0]),.doutb(w_n8461_0[1]),.din(n8461));
	jspl3 jspl3_w_n8463_0(.douta(w_n8463_0[0]),.doutb(w_n8463_0[1]),.doutc(w_n8463_0[2]),.din(n8463));
	jspl jspl_w_n8464_0(.douta(w_n8464_0[0]),.doutb(w_n8464_0[1]),.din(n8464));
	jspl3 jspl3_w_n8468_0(.douta(w_n8468_0[0]),.doutb(w_n8468_0[1]),.doutc(w_n8468_0[2]),.din(n8468));
	jspl3 jspl3_w_n8470_0(.douta(w_n8470_0[0]),.doutb(w_n8470_0[1]),.doutc(w_n8470_0[2]),.din(n8470));
	jspl jspl_w_n8471_0(.douta(w_n8471_0[0]),.doutb(w_n8471_0[1]),.din(n8471));
	jspl jspl_w_n8475_0(.douta(w_n8475_0[0]),.doutb(w_n8475_0[1]),.din(n8475));
	jspl jspl_w_n8476_0(.douta(w_n8476_0[0]),.doutb(w_n8476_0[1]),.din(n8476));
	jspl3 jspl3_w_n8478_0(.douta(w_n8478_0[0]),.doutb(w_n8478_0[1]),.doutc(w_n8478_0[2]),.din(n8478));
	jspl jspl_w_n8479_0(.douta(w_n8479_0[0]),.doutb(w_n8479_0[1]),.din(n8479));
	jspl jspl_w_n8483_0(.douta(w_n8483_0[0]),.doutb(w_n8483_0[1]),.din(n8483));
	jspl jspl_w_n8484_0(.douta(w_n8484_0[0]),.doutb(w_n8484_0[1]),.din(n8484));
	jspl3 jspl3_w_n8486_0(.douta(w_n8486_0[0]),.doutb(w_n8486_0[1]),.doutc(w_n8486_0[2]),.din(n8486));
	jspl jspl_w_n8487_0(.douta(w_n8487_0[0]),.doutb(w_n8487_0[1]),.din(n8487));
	jspl jspl_w_n8491_0(.douta(w_n8491_0[0]),.doutb(w_n8491_0[1]),.din(n8491));
	jspl jspl_w_n8492_0(.douta(w_n8492_0[0]),.doutb(w_n8492_0[1]),.din(n8492));
	jspl3 jspl3_w_n8494_0(.douta(w_n8494_0[0]),.doutb(w_n8494_0[1]),.doutc(w_n8494_0[2]),.din(n8494));
	jspl jspl_w_n8495_0(.douta(w_n8495_0[0]),.doutb(w_n8495_0[1]),.din(n8495));
	jspl jspl_w_n8498_0(.douta(w_n8498_0[0]),.doutb(w_n8498_0[1]),.din(n8498));
	jspl3 jspl3_w_n8501_0(.douta(w_n8501_0[0]),.doutb(w_n8501_0[1]),.doutc(w_n8501_0[2]),.din(n8501));
	jspl jspl_w_n8502_0(.douta(w_n8502_0[0]),.doutb(w_n8502_0[1]),.din(n8502));
	jspl jspl_w_n8506_0(.douta(w_n8506_0[0]),.doutb(w_n8506_0[1]),.din(n8506));
	jspl jspl_w_n8507_0(.douta(w_n8507_0[0]),.doutb(w_n8507_0[1]),.din(n8507));
	jspl3 jspl3_w_n8509_0(.douta(w_n8509_0[0]),.doutb(w_n8509_0[1]),.doutc(w_n8509_0[2]),.din(n8509));
	jspl jspl_w_n8510_0(.douta(w_n8510_0[0]),.doutb(w_n8510_0[1]),.din(n8510));
	jspl jspl_w_n8514_0(.douta(w_n8514_0[0]),.doutb(w_n8514_0[1]),.din(n8514));
	jspl3 jspl3_w_n8516_0(.douta(w_n8516_0[0]),.doutb(w_n8516_0[1]),.doutc(w_n8516_0[2]),.din(n8516));
	jspl jspl_w_n8517_0(.douta(w_n8517_0[0]),.doutb(w_n8517_0[1]),.din(n8517));
	jspl jspl_w_n8521_0(.douta(w_n8521_0[0]),.doutb(w_n8521_0[1]),.din(n8521));
	jspl jspl_w_n8522_0(.douta(w_n8522_0[0]),.doutb(w_n8522_0[1]),.din(n8522));
	jspl3 jspl3_w_n8524_0(.douta(w_n8524_0[0]),.doutb(w_n8524_0[1]),.doutc(w_n8524_0[2]),.din(n8524));
	jspl jspl_w_n8525_0(.douta(w_n8525_0[0]),.doutb(w_n8525_0[1]),.din(n8525));
	jspl jspl_w_n8529_0(.douta(w_n8529_0[0]),.doutb(w_n8529_0[1]),.din(n8529));
	jspl3 jspl3_w_n8531_0(.douta(w_n8531_0[0]),.doutb(w_n8531_0[1]),.doutc(w_n8531_0[2]),.din(n8531));
	jspl jspl_w_n8532_0(.douta(w_n8532_0[0]),.doutb(w_n8532_0[1]),.din(n8532));
	jspl jspl_w_n8536_0(.douta(w_n8536_0[0]),.doutb(w_n8536_0[1]),.din(n8536));
	jspl3 jspl3_w_n8538_0(.douta(w_n8538_0[0]),.doutb(w_n8538_0[1]),.doutc(w_n8538_0[2]),.din(n8538));
	jspl jspl_w_n8539_0(.douta(w_n8539_0[0]),.doutb(w_n8539_0[1]),.din(n8539));
	jspl jspl_w_n8543_0(.douta(w_n8543_0[0]),.doutb(w_n8543_0[1]),.din(n8543));
	jspl3 jspl3_w_n8545_0(.douta(w_n8545_0[0]),.doutb(w_n8545_0[1]),.doutc(w_n8545_0[2]),.din(n8545));
	jspl jspl_w_n8546_0(.douta(w_n8546_0[0]),.doutb(w_n8546_0[1]),.din(n8546));
	jspl jspl_w_n8550_0(.douta(w_n8550_0[0]),.doutb(w_n8550_0[1]),.din(n8550));
	jspl jspl_w_n8551_0(.douta(w_n8551_0[0]),.doutb(w_n8551_0[1]),.din(n8551));
	jspl3 jspl3_w_n8553_0(.douta(w_n8553_0[0]),.doutb(w_n8553_0[1]),.doutc(w_n8553_0[2]),.din(n8553));
	jspl jspl_w_n8554_0(.douta(w_n8554_0[0]),.doutb(w_n8554_0[1]),.din(n8554));
	jspl jspl_w_n8558_0(.douta(w_n8558_0[0]),.doutb(w_n8558_0[1]),.din(n8558));
	jspl3 jspl3_w_n8560_0(.douta(w_n8560_0[0]),.doutb(w_n8560_0[1]),.doutc(w_n8560_0[2]),.din(n8560));
	jspl jspl_w_n8561_0(.douta(w_n8561_0[0]),.doutb(w_n8561_0[1]),.din(n8561));
	jspl jspl_w_n8565_0(.douta(w_n8565_0[0]),.doutb(w_n8565_0[1]),.din(n8565));
	jspl jspl_w_n8566_0(.douta(w_n8566_0[0]),.doutb(w_n8566_0[1]),.din(n8566));
	jspl3 jspl3_w_n8568_0(.douta(w_n8568_0[0]),.doutb(w_n8568_0[1]),.doutc(w_n8568_0[2]),.din(n8568));
	jspl jspl_w_n8569_0(.douta(w_n8569_0[0]),.doutb(w_n8569_0[1]),.din(n8569));
	jspl jspl_w_n8573_0(.douta(w_n8573_0[0]),.doutb(w_n8573_0[1]),.din(n8573));
	jspl3 jspl3_w_n8575_0(.douta(w_n8575_0[0]),.doutb(w_n8575_0[1]),.doutc(w_n8575_0[2]),.din(n8575));
	jspl jspl_w_n8576_0(.douta(w_n8576_0[0]),.doutb(w_n8576_0[1]),.din(n8576));
	jspl jspl_w_n8580_0(.douta(w_n8580_0[0]),.doutb(w_n8580_0[1]),.din(n8580));
	jspl jspl_w_n8581_0(.douta(w_n8581_0[0]),.doutb(w_n8581_0[1]),.din(n8581));
	jspl3 jspl3_w_n8583_0(.douta(w_n8583_0[0]),.doutb(w_n8583_0[1]),.doutc(w_n8583_0[2]),.din(n8583));
	jspl jspl_w_n8584_0(.douta(w_n8584_0[0]),.doutb(w_n8584_0[1]),.din(n8584));
	jspl jspl_w_n8588_0(.douta(w_n8588_0[0]),.doutb(w_n8588_0[1]),.din(n8588));
	jspl3 jspl3_w_n8590_0(.douta(w_n8590_0[0]),.doutb(w_n8590_0[1]),.doutc(w_n8590_0[2]),.din(n8590));
	jspl jspl_w_n8591_0(.douta(w_n8591_0[0]),.doutb(w_n8591_0[1]),.din(n8591));
	jspl jspl_w_n8595_0(.douta(w_n8595_0[0]),.doutb(w_n8595_0[1]),.din(n8595));
	jspl jspl_w_n8596_0(.douta(w_n8596_0[0]),.doutb(w_n8596_0[1]),.din(n8596));
	jspl3 jspl3_w_n8598_0(.douta(w_n8598_0[0]),.doutb(w_n8598_0[1]),.doutc(w_n8598_0[2]),.din(n8598));
	jspl jspl_w_n8599_0(.douta(w_n8599_0[0]),.doutb(w_n8599_0[1]),.din(n8599));
	jspl jspl_w_n8603_0(.douta(w_n8603_0[0]),.doutb(w_n8603_0[1]),.din(n8603));
	jspl3 jspl3_w_n8605_0(.douta(w_n8605_0[0]),.doutb(w_n8605_0[1]),.doutc(w_n8605_0[2]),.din(n8605));
	jspl jspl_w_n8606_0(.douta(w_n8606_0[0]),.doutb(w_n8606_0[1]),.din(n8606));
	jspl jspl_w_n8610_0(.douta(w_n8610_0[0]),.doutb(w_n8610_0[1]),.din(n8610));
	jspl3 jspl3_w_n8612_0(.douta(w_n8612_0[0]),.doutb(w_n8612_0[1]),.doutc(w_n8612_0[2]),.din(n8612));
	jspl jspl_w_n8613_0(.douta(w_n8613_0[0]),.doutb(w_n8613_0[1]),.din(n8613));
	jspl jspl_w_n8617_0(.douta(w_n8617_0[0]),.doutb(w_n8617_0[1]),.din(n8617));
	jspl3 jspl3_w_n8619_0(.douta(w_n8619_0[0]),.doutb(w_n8619_0[1]),.doutc(w_n8619_0[2]),.din(n8619));
	jspl jspl_w_n8620_0(.douta(w_n8620_0[0]),.doutb(w_n8620_0[1]),.din(n8620));
	jspl jspl_w_n8624_0(.douta(w_n8624_0[0]),.doutb(w_n8624_0[1]),.din(n8624));
	jspl jspl_w_n8625_0(.douta(w_n8625_0[0]),.doutb(w_n8625_0[1]),.din(n8625));
	jspl3 jspl3_w_n8627_0(.douta(w_n8627_0[0]),.doutb(w_n8627_0[1]),.doutc(w_n8627_0[2]),.din(n8627));
	jspl jspl_w_n8628_0(.douta(w_n8628_0[0]),.doutb(w_n8628_0[1]),.din(n8628));
	jspl jspl_w_n8632_0(.douta(w_n8632_0[0]),.doutb(w_n8632_0[1]),.din(n8632));
	jspl jspl_w_n8633_0(.douta(w_n8633_0[0]),.doutb(w_n8633_0[1]),.din(n8633));
	jspl3 jspl3_w_n8635_0(.douta(w_n8635_0[0]),.doutb(w_n8635_0[1]),.doutc(w_n8635_0[2]),.din(n8635));
	jspl jspl_w_n8636_0(.douta(w_n8636_0[0]),.doutb(w_n8636_0[1]),.din(n8636));
	jspl jspl_w_n8640_0(.douta(w_n8640_0[0]),.doutb(w_n8640_0[1]),.din(n8640));
	jspl jspl_w_n8641_0(.douta(w_n8641_0[0]),.doutb(w_n8641_0[1]),.din(n8641));
	jspl3 jspl3_w_n8643_0(.douta(w_n8643_0[0]),.doutb(w_n8643_0[1]),.doutc(w_n8643_0[2]),.din(n8643));
	jspl jspl_w_n8644_0(.douta(w_n8644_0[0]),.doutb(w_n8644_0[1]),.din(n8644));
	jspl jspl_w_n8648_0(.douta(w_n8648_0[0]),.doutb(w_n8648_0[1]),.din(n8648));
	jspl3 jspl3_w_n8650_0(.douta(w_n8650_0[0]),.doutb(w_n8650_0[1]),.doutc(w_n8650_0[2]),.din(n8650));
	jspl jspl_w_n8651_0(.douta(w_n8651_0[0]),.doutb(w_n8651_0[1]),.din(n8651));
	jspl jspl_w_n8655_0(.douta(w_n8655_0[0]),.doutb(w_n8655_0[1]),.din(n8655));
	jspl jspl_w_n8656_0(.douta(w_n8656_0[0]),.doutb(w_n8656_0[1]),.din(n8656));
	jspl3 jspl3_w_n8658_0(.douta(w_n8658_0[0]),.doutb(w_n8658_0[1]),.doutc(w_n8658_0[2]),.din(n8658));
	jspl jspl_w_n8659_0(.douta(w_n8659_0[0]),.doutb(w_n8659_0[1]),.din(n8659));
	jspl jspl_w_n8663_0(.douta(w_n8663_0[0]),.doutb(w_n8663_0[1]),.din(n8663));
	jspl3 jspl3_w_n8665_0(.douta(w_n8665_0[0]),.doutb(w_n8665_0[1]),.doutc(w_n8665_0[2]),.din(n8665));
	jspl jspl_w_n8666_0(.douta(w_n8666_0[0]),.doutb(w_n8666_0[1]),.din(n8666));
	jspl jspl_w_n8670_0(.douta(w_n8670_0[0]),.doutb(w_n8670_0[1]),.din(n8670));
	jspl jspl_w_n8671_0(.douta(w_n8671_0[0]),.doutb(w_n8671_0[1]),.din(n8671));
	jspl3 jspl3_w_n8673_0(.douta(w_n8673_0[0]),.doutb(w_n8673_0[1]),.doutc(w_n8673_0[2]),.din(n8673));
	jspl jspl_w_n8674_0(.douta(w_n8674_0[0]),.doutb(w_n8674_0[1]),.din(n8674));
	jspl jspl_w_n8678_0(.douta(w_n8678_0[0]),.doutb(w_n8678_0[1]),.din(n8678));
	jspl3 jspl3_w_n8680_0(.douta(w_n8680_0[0]),.doutb(w_n8680_0[1]),.doutc(w_n8680_0[2]),.din(n8680));
	jspl jspl_w_n8681_0(.douta(w_n8681_0[0]),.doutb(w_n8681_0[1]),.din(n8681));
	jspl jspl_w_n8685_0(.douta(w_n8685_0[0]),.doutb(w_n8685_0[1]),.din(n8685));
	jspl3 jspl3_w_n8687_0(.douta(w_n8687_0[0]),.doutb(w_n8687_0[1]),.doutc(w_n8687_0[2]),.din(n8687));
	jspl jspl_w_n8688_0(.douta(w_n8688_0[0]),.doutb(w_n8688_0[1]),.din(n8688));
	jspl jspl_w_n8692_0(.douta(w_n8692_0[0]),.doutb(w_n8692_0[1]),.din(n8692));
	jspl jspl_w_n8693_0(.douta(w_n8693_0[0]),.doutb(w_n8693_0[1]),.din(n8693));
	jspl3 jspl3_w_n8695_0(.douta(w_n8695_0[0]),.doutb(w_n8695_0[1]),.doutc(w_n8695_0[2]),.din(n8695));
	jspl jspl_w_n8696_0(.douta(w_n8696_0[0]),.doutb(w_n8696_0[1]),.din(n8696));
	jspl3 jspl3_w_n8700_0(.douta(w_n8700_0[0]),.doutb(w_n8700_0[1]),.doutc(w_n8700_0[2]),.din(n8700));
	jspl jspl_w_n8703_0(.douta(w_n8703_0[0]),.doutb(w_n8703_0[1]),.din(n8703));
	jspl3 jspl3_w_n8704_0(.douta(w_n8704_0[0]),.doutb(w_n8704_0[1]),.doutc(w_n8704_0[2]),.din(n8704));
	jspl3 jspl3_w_n8705_0(.douta(w_n8705_0[0]),.doutb(w_n8705_0[1]),.doutc(w_n8705_0[2]),.din(n8705));
	jspl jspl_w_n8707_0(.douta(w_n8707_0[0]),.doutb(w_n8707_0[1]),.din(n8707));
	jspl jspl_w_n8736_0(.douta(w_n8736_0[0]),.doutb(w_n8736_0[1]),.din(n8736));
	jspl jspl_w_n8750_0(.douta(w_n8750_0[0]),.doutb(w_n8750_0[1]),.din(n8750));
	jspl jspl_w_n8776_0(.douta(w_n8776_0[0]),.doutb(w_n8776_0[1]),.din(n8776));
	jspl jspl_w_n8783_0(.douta(w_n8783_0[0]),.doutb(w_n8783_0[1]),.din(n8783));
	jspl jspl_w_n8787_0(.douta(w_n8787_0[0]),.doutb(w_n8787_0[1]),.din(n8787));
	jspl jspl_w_n8791_0(.douta(w_n8791_0[0]),.doutb(w_n8791_0[1]),.din(n8791));
	jspl jspl_w_n8798_0(.douta(w_n8798_0[0]),.doutb(w_n8798_0[1]),.din(n8798));
	jspl jspl_w_n8805_0(.douta(w_n8805_0[0]),.doutb(w_n8805_0[1]),.din(n8805));
	jspl jspl_w_n8812_0(.douta(w_n8812_0[0]),.doutb(w_n8812_0[1]),.din(n8812));
	jspl jspl_w_n8819_0(.douta(w_n8819_0[0]),.doutb(w_n8819_0[1]),.din(n8819));
	jspl jspl_w_n8823_0(.douta(w_n8823_0[0]),.doutb(w_n8823_0[1]),.din(n8823));
	jspl jspl_w_n8827_0(.douta(w_n8827_0[0]),.doutb(w_n8827_0[1]),.din(n8827));
	jspl jspl_w_n8840_0(.douta(w_n8840_0[0]),.doutb(w_n8840_0[1]),.din(n8840));
	jspl jspl_w_n8847_0(.douta(w_n8847_0[0]),.doutb(w_n8847_0[1]),.din(n8847));
	jspl jspl_w_n8854_0(.douta(w_n8854_0[0]),.doutb(w_n8854_0[1]),.din(n8854));
	jspl jspl_w_n8858_0(.douta(w_n8858_0[0]),.doutb(w_n8858_0[1]),.din(n8858));
	jspl jspl_w_n8866_0(.douta(w_n8866_0[0]),.doutb(w_n8866_0[1]),.din(n8866));
	jspl jspl_w_n8867_0(.douta(w_n8867_0[0]),.doutb(w_n8867_0[1]),.din(n8867));
	jspl jspl_w_n8868_0(.douta(w_n8868_0[0]),.doutb(w_n8868_0[1]),.din(n8868));
	jspl jspl_w_n8871_0(.douta(w_n8871_0[0]),.doutb(w_n8871_0[1]),.din(n8871));
	jspl jspl_w_n8874_0(.douta(w_n8874_0[0]),.doutb(w_n8874_0[1]),.din(n8874));
	jspl jspl_w_n8876_0(.douta(w_n8876_0[0]),.doutb(w_n8876_0[1]),.din(n8876));
	jspl jspl_w_n8877_0(.douta(w_n8877_0[0]),.doutb(w_n8877_0[1]),.din(n8877));
	jspl jspl_w_n8878_0(.douta(w_n8878_0[0]),.doutb(w_n8878_0[1]),.din(n8878));
	jspl jspl_w_n8882_0(.douta(w_n8882_0[0]),.doutb(w_n8882_0[1]),.din(n8882));
	jspl jspl_w_n8888_0(.douta(w_n8888_0[0]),.doutb(w_n8888_0[1]),.din(n8888));
	jspl3 jspl3_w_n8890_0(.douta(w_n8890_0[0]),.doutb(w_n8890_0[1]),.doutc(w_n8890_0[2]),.din(n8890));
	jspl3 jspl3_w_n8890_1(.douta(w_n8890_1[0]),.doutb(w_n8890_1[1]),.doutc(w_n8890_1[2]),.din(w_n8890_0[0]));
	jspl3 jspl3_w_n8890_2(.douta(w_n8890_2[0]),.doutb(w_n8890_2[1]),.doutc(w_n8890_2[2]),.din(w_n8890_0[1]));
	jspl3 jspl3_w_n8890_3(.douta(w_n8890_3[0]),.doutb(w_n8890_3[1]),.doutc(w_n8890_3[2]),.din(w_n8890_0[2]));
	jspl3 jspl3_w_n8890_4(.douta(w_n8890_4[0]),.doutb(w_n8890_4[1]),.doutc(w_n8890_4[2]),.din(w_n8890_1[0]));
	jspl3 jspl3_w_n8890_5(.douta(w_n8890_5[0]),.doutb(w_n8890_5[1]),.doutc(w_n8890_5[2]),.din(w_n8890_1[1]));
	jspl3 jspl3_w_n8890_6(.douta(w_n8890_6[0]),.doutb(w_n8890_6[1]),.doutc(w_n8890_6[2]),.din(w_n8890_1[2]));
	jspl3 jspl3_w_n8890_7(.douta(w_n8890_7[0]),.doutb(w_n8890_7[1]),.doutc(w_n8890_7[2]),.din(w_n8890_2[0]));
	jspl3 jspl3_w_n8890_8(.douta(w_n8890_8[0]),.doutb(w_n8890_8[1]),.doutc(w_n8890_8[2]),.din(w_n8890_2[1]));
	jspl3 jspl3_w_n8890_9(.douta(w_n8890_9[0]),.doutb(w_n8890_9[1]),.doutc(w_n8890_9[2]),.din(w_n8890_2[2]));
	jspl3 jspl3_w_n8890_10(.douta(w_n8890_10[0]),.doutb(w_n8890_10[1]),.doutc(w_n8890_10[2]),.din(w_n8890_3[0]));
	jspl3 jspl3_w_n8890_11(.douta(w_n8890_11[0]),.doutb(w_n8890_11[1]),.doutc(w_n8890_11[2]),.din(w_n8890_3[1]));
	jspl3 jspl3_w_n8890_12(.douta(w_n8890_12[0]),.doutb(w_n8890_12[1]),.doutc(w_n8890_12[2]),.din(w_n8890_3[2]));
	jspl3 jspl3_w_n8890_13(.douta(w_n8890_13[0]),.doutb(w_n8890_13[1]),.doutc(w_n8890_13[2]),.din(w_n8890_4[0]));
	jspl3 jspl3_w_n8890_14(.douta(w_n8890_14[0]),.doutb(w_n8890_14[1]),.doutc(w_n8890_14[2]),.din(w_n8890_4[1]));
	jspl3 jspl3_w_n8890_15(.douta(w_n8890_15[0]),.doutb(w_n8890_15[1]),.doutc(w_n8890_15[2]),.din(w_n8890_4[2]));
	jspl3 jspl3_w_n8890_16(.douta(w_n8890_16[0]),.doutb(w_n8890_16[1]),.doutc(w_n8890_16[2]),.din(w_n8890_5[0]));
	jspl3 jspl3_w_n8890_17(.douta(w_n8890_17[0]),.doutb(w_n8890_17[1]),.doutc(w_n8890_17[2]),.din(w_n8890_5[1]));
	jspl3 jspl3_w_n8890_18(.douta(w_n8890_18[0]),.doutb(w_n8890_18[1]),.doutc(w_n8890_18[2]),.din(w_n8890_5[2]));
	jspl3 jspl3_w_n8890_19(.douta(w_n8890_19[0]),.doutb(w_n8890_19[1]),.doutc(w_n8890_19[2]),.din(w_n8890_6[0]));
	jspl3 jspl3_w_n8890_20(.douta(w_n8890_20[0]),.doutb(w_n8890_20[1]),.doutc(w_n8890_20[2]),.din(w_n8890_6[1]));
	jspl3 jspl3_w_n8890_21(.douta(w_n8890_21[0]),.doutb(w_n8890_21[1]),.doutc(w_n8890_21[2]),.din(w_n8890_6[2]));
	jspl3 jspl3_w_n8890_22(.douta(w_n8890_22[0]),.doutb(w_n8890_22[1]),.doutc(w_n8890_22[2]),.din(w_n8890_7[0]));
	jspl3 jspl3_w_n8890_23(.douta(w_n8890_23[0]),.doutb(w_n8890_23[1]),.doutc(w_n8890_23[2]),.din(w_n8890_7[1]));
	jspl3 jspl3_w_n8890_24(.douta(w_n8890_24[0]),.doutb(w_n8890_24[1]),.doutc(w_n8890_24[2]),.din(w_n8890_7[2]));
	jspl3 jspl3_w_n8890_25(.douta(w_n8890_25[0]),.doutb(w_n8890_25[1]),.doutc(w_n8890_25[2]),.din(w_n8890_8[0]));
	jspl3 jspl3_w_n8890_26(.douta(w_n8890_26[0]),.doutb(w_n8890_26[1]),.doutc(w_n8890_26[2]),.din(w_n8890_8[1]));
	jspl3 jspl3_w_n8890_27(.douta(w_n8890_27[0]),.doutb(w_n8890_27[1]),.doutc(w_n8890_27[2]),.din(w_n8890_8[2]));
	jspl3 jspl3_w_n8890_28(.douta(w_n8890_28[0]),.doutb(w_n8890_28[1]),.doutc(w_n8890_28[2]),.din(w_n8890_9[0]));
	jspl3 jspl3_w_n8890_29(.douta(w_n8890_29[0]),.doutb(w_n8890_29[1]),.doutc(w_n8890_29[2]),.din(w_n8890_9[1]));
	jspl3 jspl3_w_n8890_30(.douta(w_n8890_30[0]),.doutb(w_n8890_30[1]),.doutc(w_n8890_30[2]),.din(w_n8890_9[2]));
	jspl3 jspl3_w_n8890_31(.douta(w_n8890_31[0]),.doutb(w_n8890_31[1]),.doutc(w_n8890_31[2]),.din(w_n8890_10[0]));
	jspl3 jspl3_w_n8890_32(.douta(w_n8890_32[0]),.doutb(w_n8890_32[1]),.doutc(w_n8890_32[2]),.din(w_n8890_10[1]));
	jspl3 jspl3_w_n8890_33(.douta(w_n8890_33[0]),.doutb(w_n8890_33[1]),.doutc(w_n8890_33[2]),.din(w_n8890_10[2]));
	jspl3 jspl3_w_n8890_34(.douta(w_n8890_34[0]),.doutb(w_n8890_34[1]),.doutc(w_n8890_34[2]),.din(w_n8890_11[0]));
	jspl3 jspl3_w_n8890_35(.douta(w_n8890_35[0]),.doutb(w_n8890_35[1]),.doutc(w_n8890_35[2]),.din(w_n8890_11[1]));
	jspl3 jspl3_w_n8890_36(.douta(w_n8890_36[0]),.doutb(w_n8890_36[1]),.doutc(w_n8890_36[2]),.din(w_n8890_11[2]));
	jspl3 jspl3_w_n8890_37(.douta(w_n8890_37[0]),.doutb(w_n8890_37[1]),.doutc(w_n8890_37[2]),.din(w_n8890_12[0]));
	jspl3 jspl3_w_n8890_38(.douta(w_n8890_38[0]),.doutb(w_n8890_38[1]),.doutc(w_n8890_38[2]),.din(w_n8890_12[1]));
	jspl3 jspl3_w_n8890_39(.douta(w_n8890_39[0]),.doutb(w_n8890_39[1]),.doutc(w_n8890_39[2]),.din(w_n8890_12[2]));
	jspl3 jspl3_w_n8890_40(.douta(w_n8890_40[0]),.doutb(w_n8890_40[1]),.doutc(w_n8890_40[2]),.din(w_n8890_13[0]));
	jspl3 jspl3_w_n8890_41(.douta(w_n8890_41[0]),.doutb(w_n8890_41[1]),.doutc(w_n8890_41[2]),.din(w_n8890_13[1]));
	jspl3 jspl3_w_n8890_42(.douta(w_n8890_42[0]),.doutb(w_n8890_42[1]),.doutc(w_n8890_42[2]),.din(w_n8890_13[2]));
	jspl3 jspl3_w_n8890_43(.douta(w_n8890_43[0]),.doutb(w_n8890_43[1]),.doutc(w_n8890_43[2]),.din(w_n8890_14[0]));
	jspl3 jspl3_w_n8890_44(.douta(w_n8890_44[0]),.doutb(w_n8890_44[1]),.doutc(w_n8890_44[2]),.din(w_n8890_14[1]));
	jspl3 jspl3_w_n8890_45(.douta(w_n8890_45[0]),.doutb(w_n8890_45[1]),.doutc(w_n8890_45[2]),.din(w_n8890_14[2]));
	jspl3 jspl3_w_n8890_46(.douta(w_n8890_46[0]),.doutb(w_n8890_46[1]),.doutc(w_n8890_46[2]),.din(w_n8890_15[0]));
	jspl3 jspl3_w_n8890_47(.douta(w_n8890_47[0]),.doutb(w_n8890_47[1]),.doutc(w_n8890_47[2]),.din(w_n8890_15[1]));
	jspl3 jspl3_w_n8890_48(.douta(w_n8890_48[0]),.doutb(w_n8890_48[1]),.doutc(w_n8890_48[2]),.din(w_n8890_15[2]));
	jspl3 jspl3_w_n8890_49(.douta(w_n8890_49[0]),.doutb(w_n8890_49[1]),.doutc(w_n8890_49[2]),.din(w_n8890_16[0]));
	jspl jspl_w_n8890_50(.douta(w_n8890_50[0]),.doutb(w_n8890_50[1]),.din(w_n8890_16[1]));
	jspl jspl_w_n8893_0(.douta(w_n8893_0[0]),.doutb(w_n8893_0[1]),.din(n8893));
	jspl3 jspl3_w_n8894_0(.douta(w_n8894_0[0]),.doutb(w_n8894_0[1]),.doutc(w_n8894_0[2]),.din(n8894));
	jspl jspl_w_n8894_1(.douta(w_n8894_1[0]),.doutb(w_n8894_1[1]),.din(w_n8894_0[0]));
	jspl3 jspl3_w_n8895_0(.douta(w_n8895_0[0]),.doutb(w_n8895_0[1]),.doutc(w_n8895_0[2]),.din(n8895));
	jspl3 jspl3_w_n8895_1(.douta(w_n8895_1[0]),.doutb(w_n8895_1[1]),.doutc(w_n8895_1[2]),.din(w_n8895_0[0]));
	jspl jspl_w_n8896_0(.douta(w_n8896_0[0]),.doutb(w_n8896_0[1]),.din(n8896));
	jspl3 jspl3_w_n8897_0(.douta(w_n8897_0[0]),.doutb(w_n8897_0[1]),.doutc(w_n8897_0[2]),.din(n8897));
	jspl jspl_w_n8898_0(.douta(w_n8898_0[0]),.doutb(w_n8898_0[1]),.din(n8898));
	jspl3 jspl3_w_n8901_0(.douta(w_n8901_0[0]),.doutb(w_n8901_0[1]),.doutc(w_n8901_0[2]),.din(n8901));
	jspl jspl_w_n8902_0(.douta(w_n8902_0[0]),.doutb(w_n8902_0[1]),.din(n8902));
	jspl3 jspl3_w_n8909_0(.douta(w_n8909_0[0]),.doutb(w_n8909_0[1]),.doutc(w_n8909_0[2]),.din(n8909));
	jspl jspl_w_n8910_0(.douta(w_n8910_0[0]),.doutb(w_n8910_0[1]),.din(n8910));
	jspl jspl_w_n8913_0(.douta(w_n8913_0[0]),.doutb(w_n8913_0[1]),.din(n8913));
	jspl3 jspl3_w_n8918_0(.douta(w_n8918_0[0]),.doutb(w_n8918_0[1]),.doutc(w_n8918_0[2]),.din(n8918));
	jspl3 jspl3_w_n8920_0(.douta(w_n8920_0[0]),.doutb(w_n8920_0[1]),.doutc(w_n8920_0[2]),.din(n8920));
	jspl jspl_w_n8921_0(.douta(w_n8921_0[0]),.doutb(w_n8921_0[1]),.din(n8921));
	jspl3 jspl3_w_n8925_0(.douta(w_n8925_0[0]),.doutb(w_n8925_0[1]),.doutc(w_n8925_0[2]),.din(n8925));
	jspl3 jspl3_w_n8928_0(.douta(w_n8928_0[0]),.doutb(w_n8928_0[1]),.doutc(w_n8928_0[2]),.din(n8928));
	jspl jspl_w_n8929_0(.douta(w_n8929_0[0]),.doutb(w_n8929_0[1]),.din(n8929));
	jspl3 jspl3_w_n8933_0(.douta(w_n8933_0[0]),.doutb(w_n8933_0[1]),.doutc(w_n8933_0[2]),.din(n8933));
	jspl3 jspl3_w_n8935_0(.douta(w_n8935_0[0]),.doutb(w_n8935_0[1]),.doutc(w_n8935_0[2]),.din(n8935));
	jspl jspl_w_n8936_0(.douta(w_n8936_0[0]),.doutb(w_n8936_0[1]),.din(n8936));
	jspl3 jspl3_w_n8940_0(.douta(w_n8940_0[0]),.doutb(w_n8940_0[1]),.doutc(w_n8940_0[2]),.din(n8940));
	jspl3 jspl3_w_n8942_0(.douta(w_n8942_0[0]),.doutb(w_n8942_0[1]),.doutc(w_n8942_0[2]),.din(n8942));
	jspl jspl_w_n8943_0(.douta(w_n8943_0[0]),.doutb(w_n8943_0[1]),.din(n8943));
	jspl3 jspl3_w_n8947_0(.douta(w_n8947_0[0]),.doutb(w_n8947_0[1]),.doutc(w_n8947_0[2]),.din(n8947));
	jspl3 jspl3_w_n8949_0(.douta(w_n8949_0[0]),.doutb(w_n8949_0[1]),.doutc(w_n8949_0[2]),.din(n8949));
	jspl jspl_w_n8950_0(.douta(w_n8950_0[0]),.doutb(w_n8950_0[1]),.din(n8950));
	jspl3 jspl3_w_n8954_0(.douta(w_n8954_0[0]),.doutb(w_n8954_0[1]),.doutc(w_n8954_0[2]),.din(n8954));
	jspl3 jspl3_w_n8956_0(.douta(w_n8956_0[0]),.doutb(w_n8956_0[1]),.doutc(w_n8956_0[2]),.din(n8956));
	jspl jspl_w_n8957_0(.douta(w_n8957_0[0]),.doutb(w_n8957_0[1]),.din(n8957));
	jspl3 jspl3_w_n8961_0(.douta(w_n8961_0[0]),.doutb(w_n8961_0[1]),.doutc(w_n8961_0[2]),.din(n8961));
	jspl3 jspl3_w_n8963_0(.douta(w_n8963_0[0]),.doutb(w_n8963_0[1]),.doutc(w_n8963_0[2]),.din(n8963));
	jspl jspl_w_n8964_0(.douta(w_n8964_0[0]),.doutb(w_n8964_0[1]),.din(n8964));
	jspl3 jspl3_w_n8967_0(.douta(w_n8967_0[0]),.doutb(w_n8967_0[1]),.doutc(w_n8967_0[2]),.din(n8967));
	jspl3 jspl3_w_n8971_0(.douta(w_n8971_0[0]),.doutb(w_n8971_0[1]),.doutc(w_n8971_0[2]),.din(n8971));
	jspl jspl_w_n8972_0(.douta(w_n8972_0[0]),.doutb(w_n8972_0[1]),.din(n8972));
	jspl3 jspl3_w_n8976_0(.douta(w_n8976_0[0]),.doutb(w_n8976_0[1]),.doutc(w_n8976_0[2]),.din(n8976));
	jspl3 jspl3_w_n8978_0(.douta(w_n8978_0[0]),.doutb(w_n8978_0[1]),.doutc(w_n8978_0[2]),.din(n8978));
	jspl jspl_w_n8979_0(.douta(w_n8979_0[0]),.doutb(w_n8979_0[1]),.din(n8979));
	jspl3 jspl3_w_n8983_0(.douta(w_n8983_0[0]),.doutb(w_n8983_0[1]),.doutc(w_n8983_0[2]),.din(n8983));
	jspl3 jspl3_w_n8986_0(.douta(w_n8986_0[0]),.doutb(w_n8986_0[1]),.doutc(w_n8986_0[2]),.din(n8986));
	jspl jspl_w_n8987_0(.douta(w_n8987_0[0]),.doutb(w_n8987_0[1]),.din(n8987));
	jspl3 jspl3_w_n8991_0(.douta(w_n8991_0[0]),.doutb(w_n8991_0[1]),.doutc(w_n8991_0[2]),.din(n8991));
	jspl3 jspl3_w_n8993_0(.douta(w_n8993_0[0]),.doutb(w_n8993_0[1]),.doutc(w_n8993_0[2]),.din(n8993));
	jspl jspl_w_n8994_0(.douta(w_n8994_0[0]),.doutb(w_n8994_0[1]),.din(n8994));
	jspl3 jspl3_w_n8998_0(.douta(w_n8998_0[0]),.doutb(w_n8998_0[1]),.doutc(w_n8998_0[2]),.din(n8998));
	jspl3 jspl3_w_n9001_0(.douta(w_n9001_0[0]),.doutb(w_n9001_0[1]),.doutc(w_n9001_0[2]),.din(n9001));
	jspl jspl_w_n9002_0(.douta(w_n9002_0[0]),.doutb(w_n9002_0[1]),.din(n9002));
	jspl3 jspl3_w_n9006_0(.douta(w_n9006_0[0]),.doutb(w_n9006_0[1]),.doutc(w_n9006_0[2]),.din(n9006));
	jspl3 jspl3_w_n9009_0(.douta(w_n9009_0[0]),.doutb(w_n9009_0[1]),.doutc(w_n9009_0[2]),.din(n9009));
	jspl jspl_w_n9010_0(.douta(w_n9010_0[0]),.doutb(w_n9010_0[1]),.din(n9010));
	jspl jspl_w_n9014_0(.douta(w_n9014_0[0]),.doutb(w_n9014_0[1]),.din(n9014));
	jspl jspl_w_n9015_0(.douta(w_n9015_0[0]),.doutb(w_n9015_0[1]),.din(n9015));
	jspl3 jspl3_w_n9017_0(.douta(w_n9017_0[0]),.doutb(w_n9017_0[1]),.doutc(w_n9017_0[2]),.din(n9017));
	jspl jspl_w_n9018_0(.douta(w_n9018_0[0]),.doutb(w_n9018_0[1]),.din(n9018));
	jspl3 jspl3_w_n9022_0(.douta(w_n9022_0[0]),.doutb(w_n9022_0[1]),.doutc(w_n9022_0[2]),.din(n9022));
	jspl3 jspl3_w_n9024_0(.douta(w_n9024_0[0]),.doutb(w_n9024_0[1]),.doutc(w_n9024_0[2]),.din(n9024));
	jspl jspl_w_n9025_0(.douta(w_n9025_0[0]),.doutb(w_n9025_0[1]),.din(n9025));
	jspl3 jspl3_w_n9029_0(.douta(w_n9029_0[0]),.doutb(w_n9029_0[1]),.doutc(w_n9029_0[2]),.din(n9029));
	jspl3 jspl3_w_n9032_0(.douta(w_n9032_0[0]),.doutb(w_n9032_0[1]),.doutc(w_n9032_0[2]),.din(n9032));
	jspl jspl_w_n9033_0(.douta(w_n9033_0[0]),.doutb(w_n9033_0[1]),.din(n9033));
	jspl3 jspl3_w_n9037_0(.douta(w_n9037_0[0]),.doutb(w_n9037_0[1]),.doutc(w_n9037_0[2]),.din(n9037));
	jspl3 jspl3_w_n9039_0(.douta(w_n9039_0[0]),.doutb(w_n9039_0[1]),.doutc(w_n9039_0[2]),.din(n9039));
	jspl jspl_w_n9040_0(.douta(w_n9040_0[0]),.doutb(w_n9040_0[1]),.din(n9040));
	jspl3 jspl3_w_n9044_0(.douta(w_n9044_0[0]),.doutb(w_n9044_0[1]),.doutc(w_n9044_0[2]),.din(n9044));
	jspl3 jspl3_w_n9047_0(.douta(w_n9047_0[0]),.doutb(w_n9047_0[1]),.doutc(w_n9047_0[2]),.din(n9047));
	jspl jspl_w_n9048_0(.douta(w_n9048_0[0]),.doutb(w_n9048_0[1]),.din(n9048));
	jspl3 jspl3_w_n9052_0(.douta(w_n9052_0[0]),.doutb(w_n9052_0[1]),.doutc(w_n9052_0[2]),.din(n9052));
	jspl3 jspl3_w_n9054_0(.douta(w_n9054_0[0]),.doutb(w_n9054_0[1]),.doutc(w_n9054_0[2]),.din(n9054));
	jspl jspl_w_n9055_0(.douta(w_n9055_0[0]),.doutb(w_n9055_0[1]),.din(n9055));
	jspl3 jspl3_w_n9059_0(.douta(w_n9059_0[0]),.doutb(w_n9059_0[1]),.doutc(w_n9059_0[2]),.din(n9059));
	jspl3 jspl3_w_n9062_0(.douta(w_n9062_0[0]),.doutb(w_n9062_0[1]),.doutc(w_n9062_0[2]),.din(n9062));
	jspl jspl_w_n9063_0(.douta(w_n9063_0[0]),.doutb(w_n9063_0[1]),.din(n9063));
	jspl3 jspl3_w_n9067_0(.douta(w_n9067_0[0]),.doutb(w_n9067_0[1]),.doutc(w_n9067_0[2]),.din(n9067));
	jspl3 jspl3_w_n9069_0(.douta(w_n9069_0[0]),.doutb(w_n9069_0[1]),.doutc(w_n9069_0[2]),.din(n9069));
	jspl jspl_w_n9070_0(.douta(w_n9070_0[0]),.doutb(w_n9070_0[1]),.din(n9070));
	jspl3 jspl3_w_n9074_0(.douta(w_n9074_0[0]),.doutb(w_n9074_0[1]),.doutc(w_n9074_0[2]),.din(n9074));
	jspl3 jspl3_w_n9077_0(.douta(w_n9077_0[0]),.doutb(w_n9077_0[1]),.doutc(w_n9077_0[2]),.din(n9077));
	jspl jspl_w_n9078_0(.douta(w_n9078_0[0]),.doutb(w_n9078_0[1]),.din(n9078));
	jspl3 jspl3_w_n9082_0(.douta(w_n9082_0[0]),.doutb(w_n9082_0[1]),.doutc(w_n9082_0[2]),.din(n9082));
	jspl3 jspl3_w_n9085_0(.douta(w_n9085_0[0]),.doutb(w_n9085_0[1]),.doutc(w_n9085_0[2]),.din(n9085));
	jspl jspl_w_n9086_0(.douta(w_n9086_0[0]),.doutb(w_n9086_0[1]),.din(n9086));
	jspl3 jspl3_w_n9090_0(.douta(w_n9090_0[0]),.doutb(w_n9090_0[1]),.doutc(w_n9090_0[2]),.din(n9090));
	jspl3 jspl3_w_n9093_0(.douta(w_n9093_0[0]),.doutb(w_n9093_0[1]),.doutc(w_n9093_0[2]),.din(n9093));
	jspl jspl_w_n9094_0(.douta(w_n9094_0[0]),.doutb(w_n9094_0[1]),.din(n9094));
	jspl3 jspl3_w_n9098_0(.douta(w_n9098_0[0]),.doutb(w_n9098_0[1]),.doutc(w_n9098_0[2]),.din(n9098));
	jspl3 jspl3_w_n9100_0(.douta(w_n9100_0[0]),.doutb(w_n9100_0[1]),.doutc(w_n9100_0[2]),.din(n9100));
	jspl jspl_w_n9101_0(.douta(w_n9101_0[0]),.doutb(w_n9101_0[1]),.din(n9101));
	jspl3 jspl3_w_n9105_0(.douta(w_n9105_0[0]),.doutb(w_n9105_0[1]),.doutc(w_n9105_0[2]),.din(n9105));
	jspl3 jspl3_w_n9107_0(.douta(w_n9107_0[0]),.doutb(w_n9107_0[1]),.doutc(w_n9107_0[2]),.din(n9107));
	jspl jspl_w_n9108_0(.douta(w_n9108_0[0]),.doutb(w_n9108_0[1]),.din(n9108));
	jspl3 jspl3_w_n9112_0(.douta(w_n9112_0[0]),.doutb(w_n9112_0[1]),.doutc(w_n9112_0[2]),.din(n9112));
	jspl3 jspl3_w_n9114_0(.douta(w_n9114_0[0]),.doutb(w_n9114_0[1]),.doutc(w_n9114_0[2]),.din(n9114));
	jspl jspl_w_n9115_0(.douta(w_n9115_0[0]),.doutb(w_n9115_0[1]),.din(n9115));
	jspl3 jspl3_w_n9119_0(.douta(w_n9119_0[0]),.doutb(w_n9119_0[1]),.doutc(w_n9119_0[2]),.din(n9119));
	jspl3 jspl3_w_n9122_0(.douta(w_n9122_0[0]),.doutb(w_n9122_0[1]),.doutc(w_n9122_0[2]),.din(n9122));
	jspl jspl_w_n9123_0(.douta(w_n9123_0[0]),.doutb(w_n9123_0[1]),.din(n9123));
	jspl3 jspl3_w_n9127_0(.douta(w_n9127_0[0]),.doutb(w_n9127_0[1]),.doutc(w_n9127_0[2]),.din(n9127));
	jspl3 jspl3_w_n9129_0(.douta(w_n9129_0[0]),.doutb(w_n9129_0[1]),.doutc(w_n9129_0[2]),.din(n9129));
	jspl jspl_w_n9130_0(.douta(w_n9130_0[0]),.doutb(w_n9130_0[1]),.din(n9130));
	jspl jspl_w_n9134_0(.douta(w_n9134_0[0]),.doutb(w_n9134_0[1]),.din(n9134));
	jspl jspl_w_n9135_0(.douta(w_n9135_0[0]),.doutb(w_n9135_0[1]),.din(n9135));
	jspl3 jspl3_w_n9137_0(.douta(w_n9137_0[0]),.doutb(w_n9137_0[1]),.doutc(w_n9137_0[2]),.din(n9137));
	jspl jspl_w_n9138_0(.douta(w_n9138_0[0]),.doutb(w_n9138_0[1]),.din(n9138));
	jspl3 jspl3_w_n9142_0(.douta(w_n9142_0[0]),.doutb(w_n9142_0[1]),.doutc(w_n9142_0[2]),.din(n9142));
	jspl3 jspl3_w_n9144_0(.douta(w_n9144_0[0]),.doutb(w_n9144_0[1]),.doutc(w_n9144_0[2]),.din(n9144));
	jspl jspl_w_n9145_0(.douta(w_n9145_0[0]),.doutb(w_n9145_0[1]),.din(n9145));
	jspl3 jspl3_w_n9149_0(.douta(w_n9149_0[0]),.doutb(w_n9149_0[1]),.doutc(w_n9149_0[2]),.din(n9149));
	jspl3 jspl3_w_n9152_0(.douta(w_n9152_0[0]),.doutb(w_n9152_0[1]),.doutc(w_n9152_0[2]),.din(n9152));
	jspl jspl_w_n9153_0(.douta(w_n9153_0[0]),.doutb(w_n9153_0[1]),.din(n9153));
	jspl3 jspl3_w_n9157_0(.douta(w_n9157_0[0]),.doutb(w_n9157_0[1]),.doutc(w_n9157_0[2]),.din(n9157));
	jspl3 jspl3_w_n9160_0(.douta(w_n9160_0[0]),.doutb(w_n9160_0[1]),.doutc(w_n9160_0[2]),.din(n9160));
	jspl jspl_w_n9161_0(.douta(w_n9161_0[0]),.doutb(w_n9161_0[1]),.din(n9161));
	jspl jspl_w_n9165_0(.douta(w_n9165_0[0]),.doutb(w_n9165_0[1]),.din(n9165));
	jspl3 jspl3_w_n9167_0(.douta(w_n9167_0[0]),.doutb(w_n9167_0[1]),.doutc(w_n9167_0[2]),.din(n9167));
	jspl jspl_w_n9167_1(.douta(w_n9167_1[0]),.doutb(w_n9167_1[1]),.din(w_n9167_0[0]));
	jspl jspl_w_n9168_0(.douta(w_n9168_0[0]),.doutb(w_n9168_0[1]),.din(n9168));
	jspl jspl_w_n9172_0(.douta(w_n9172_0[0]),.doutb(w_n9172_0[1]),.din(n9172));
	jspl jspl_w_n9173_0(.douta(w_n9173_0[0]),.doutb(w_n9173_0[1]),.din(n9173));
	jspl jspl_w_n9177_0(.douta(w_n9177_0[0]),.doutb(w_n9177_0[1]),.din(n9177));
	jspl jspl_w_n9180_0(.douta(w_n9180_0[0]),.doutb(w_n9180_0[1]),.din(n9180));
	jspl jspl_w_n9184_0(.douta(w_n9184_0[0]),.doutb(w_n9184_0[1]),.din(n9184));
	jspl3 jspl3_w_n9187_0(.douta(w_n9187_0[0]),.doutb(w_n9187_0[1]),.doutc(w_n9187_0[2]),.din(n9187));
	jspl3 jspl3_w_n9188_0(.douta(w_n9188_0[0]),.doutb(w_n9188_0[1]),.doutc(w_n9188_0[2]),.din(n9188));
	jspl3 jspl3_w_n9188_1(.douta(w_n9188_1[0]),.doutb(w_n9188_1[1]),.doutc(w_n9188_1[2]),.din(w_n9188_0[0]));
	jspl jspl_w_n9189_0(.douta(w_n9189_0[0]),.doutb(w_n9189_0[1]),.din(n9189));
	jspl3 jspl3_w_n9190_0(.douta(w_n9190_0[0]),.doutb(w_n9190_0[1]),.doutc(w_n9190_0[2]),.din(n9190));
	jspl jspl_w_n9191_0(.douta(w_n9191_0[0]),.doutb(w_n9191_0[1]),.din(n9191));
	jspl3 jspl3_w_n9193_0(.douta(w_n9193_0[0]),.doutb(w_n9193_0[1]),.doutc(w_n9193_0[2]),.din(n9193));
	jspl jspl_w_n9194_0(.douta(w_n9194_0[0]),.doutb(w_n9194_0[1]),.din(n9194));
	jspl jspl_w_n9199_0(.douta(w_n9199_0[0]),.doutb(w_n9199_0[1]),.din(n9199));
	jspl jspl_w_n9240_0(.douta(w_n9240_0[0]),.doutb(w_n9240_0[1]),.din(n9240));
	jspl jspl_w_n9365_0(.douta(w_n9365_0[0]),.doutb(w_n9365_0[1]),.din(n9365));
	jspl jspl_w_n9368_0(.douta(w_n9368_0[0]),.doutb(w_n9368_0[1]),.din(n9368));
	jspl3 jspl3_w_n9369_0(.douta(w_n9369_0[0]),.doutb(w_n9369_0[1]),.doutc(w_n9369_0[2]),.din(n9369));
	jspl3 jspl3_w_n9369_1(.douta(w_n9369_1[0]),.doutb(w_n9369_1[1]),.doutc(w_n9369_1[2]),.din(w_n9369_0[0]));
	jspl3 jspl3_w_n9369_2(.douta(w_n9369_2[0]),.doutb(w_n9369_2[1]),.doutc(w_n9369_2[2]),.din(w_n9369_0[1]));
	jspl3 jspl3_w_n9369_3(.douta(w_n9369_3[0]),.doutb(w_n9369_3[1]),.doutc(w_n9369_3[2]),.din(w_n9369_0[2]));
	jspl3 jspl3_w_n9369_4(.douta(w_n9369_4[0]),.doutb(w_n9369_4[1]),.doutc(w_n9369_4[2]),.din(w_n9369_1[0]));
	jspl3 jspl3_w_n9369_5(.douta(w_n9369_5[0]),.doutb(w_n9369_5[1]),.doutc(w_n9369_5[2]),.din(w_n9369_1[1]));
	jspl3 jspl3_w_n9369_6(.douta(w_n9369_6[0]),.doutb(w_n9369_6[1]),.doutc(w_n9369_6[2]),.din(w_n9369_1[2]));
	jspl3 jspl3_w_n9369_7(.douta(w_n9369_7[0]),.doutb(w_n9369_7[1]),.doutc(w_n9369_7[2]),.din(w_n9369_2[0]));
	jspl3 jspl3_w_n9369_8(.douta(w_n9369_8[0]),.doutb(w_n9369_8[1]),.doutc(w_n9369_8[2]),.din(w_n9369_2[1]));
	jspl3 jspl3_w_n9369_9(.douta(w_n9369_9[0]),.doutb(w_n9369_9[1]),.doutc(w_n9369_9[2]),.din(w_n9369_2[2]));
	jspl3 jspl3_w_n9369_10(.douta(w_n9369_10[0]),.doutb(w_n9369_10[1]),.doutc(w_n9369_10[2]),.din(w_n9369_3[0]));
	jspl3 jspl3_w_n9369_11(.douta(w_n9369_11[0]),.doutb(w_n9369_11[1]),.doutc(w_n9369_11[2]),.din(w_n9369_3[1]));
	jspl3 jspl3_w_n9369_12(.douta(w_n9369_12[0]),.doutb(w_n9369_12[1]),.doutc(w_n9369_12[2]),.din(w_n9369_3[2]));
	jspl3 jspl3_w_n9369_13(.douta(w_n9369_13[0]),.doutb(w_n9369_13[1]),.doutc(w_n9369_13[2]),.din(w_n9369_4[0]));
	jspl3 jspl3_w_n9369_14(.douta(w_n9369_14[0]),.doutb(w_n9369_14[1]),.doutc(w_n9369_14[2]),.din(w_n9369_4[1]));
	jspl3 jspl3_w_n9369_15(.douta(w_n9369_15[0]),.doutb(w_n9369_15[1]),.doutc(w_n9369_15[2]),.din(w_n9369_4[2]));
	jspl3 jspl3_w_n9369_16(.douta(w_n9369_16[0]),.doutb(w_n9369_16[1]),.doutc(w_n9369_16[2]),.din(w_n9369_5[0]));
	jspl3 jspl3_w_n9369_17(.douta(w_n9369_17[0]),.doutb(w_n9369_17[1]),.doutc(w_n9369_17[2]),.din(w_n9369_5[1]));
	jspl3 jspl3_w_n9369_18(.douta(w_n9369_18[0]),.doutb(w_n9369_18[1]),.doutc(w_n9369_18[2]),.din(w_n9369_5[2]));
	jspl3 jspl3_w_n9369_19(.douta(w_n9369_19[0]),.doutb(w_n9369_19[1]),.doutc(w_n9369_19[2]),.din(w_n9369_6[0]));
	jspl3 jspl3_w_n9369_20(.douta(w_n9369_20[0]),.doutb(w_n9369_20[1]),.doutc(w_n9369_20[2]),.din(w_n9369_6[1]));
	jspl3 jspl3_w_n9369_21(.douta(w_n9369_21[0]),.doutb(w_n9369_21[1]),.doutc(w_n9369_21[2]),.din(w_n9369_6[2]));
	jspl3 jspl3_w_n9369_22(.douta(w_n9369_22[0]),.doutb(w_n9369_22[1]),.doutc(w_n9369_22[2]),.din(w_n9369_7[0]));
	jspl3 jspl3_w_n9369_23(.douta(w_n9369_23[0]),.doutb(w_n9369_23[1]),.doutc(w_n9369_23[2]),.din(w_n9369_7[1]));
	jspl3 jspl3_w_n9369_24(.douta(w_n9369_24[0]),.doutb(w_n9369_24[1]),.doutc(w_n9369_24[2]),.din(w_n9369_7[2]));
	jspl3 jspl3_w_n9369_25(.douta(w_n9369_25[0]),.doutb(w_n9369_25[1]),.doutc(w_n9369_25[2]),.din(w_n9369_8[0]));
	jspl3 jspl3_w_n9369_26(.douta(w_n9369_26[0]),.doutb(w_n9369_26[1]),.doutc(w_n9369_26[2]),.din(w_n9369_8[1]));
	jspl3 jspl3_w_n9369_27(.douta(w_n9369_27[0]),.doutb(w_n9369_27[1]),.doutc(w_n9369_27[2]),.din(w_n9369_8[2]));
	jspl3 jspl3_w_n9369_28(.douta(w_n9369_28[0]),.doutb(w_n9369_28[1]),.doutc(w_n9369_28[2]),.din(w_n9369_9[0]));
	jspl3 jspl3_w_n9369_29(.douta(w_n9369_29[0]),.doutb(w_n9369_29[1]),.doutc(w_n9369_29[2]),.din(w_n9369_9[1]));
	jspl3 jspl3_w_n9369_30(.douta(w_n9369_30[0]),.doutb(w_n9369_30[1]),.doutc(w_n9369_30[2]),.din(w_n9369_9[2]));
	jspl3 jspl3_w_n9369_31(.douta(w_n9369_31[0]),.doutb(w_n9369_31[1]),.doutc(w_n9369_31[2]),.din(w_n9369_10[0]));
	jspl3 jspl3_w_n9369_32(.douta(w_n9369_32[0]),.doutb(w_n9369_32[1]),.doutc(w_n9369_32[2]),.din(w_n9369_10[1]));
	jspl jspl_w_n9369_33(.douta(w_n9369_33[0]),.doutb(w_n9369_33[1]),.din(w_n9369_10[2]));
	jspl3 jspl3_w_n9373_0(.douta(w_n9373_0[0]),.doutb(w_n9373_0[1]),.doutc(w_n9373_0[2]),.din(n9373));
	jspl jspl_w_n9374_0(.douta(w_n9374_0[0]),.doutb(w_n9374_0[1]),.din(n9374));
	jspl jspl_w_n9376_0(.douta(w_n9376_0[0]),.doutb(w_n9376_0[1]),.din(n9376));
	jspl jspl_w_n9381_0(.douta(w_n9381_0[0]),.doutb(w_n9381_0[1]),.din(n9381));
	jspl jspl_w_n9382_0(.douta(w_n9382_0[0]),.doutb(w_n9382_0[1]),.din(n9382));
	jspl3 jspl3_w_n9384_0(.douta(w_n9384_0[0]),.doutb(w_n9384_0[1]),.doutc(w_n9384_0[2]),.din(n9384));
	jspl jspl_w_n9385_0(.douta(w_n9385_0[0]),.doutb(w_n9385_0[1]),.din(n9385));
	jspl3 jspl3_w_n9389_0(.douta(w_n9389_0[0]),.doutb(w_n9389_0[1]),.doutc(w_n9389_0[2]),.din(n9389));
	jspl3 jspl3_w_n9391_0(.douta(w_n9391_0[0]),.doutb(w_n9391_0[1]),.doutc(w_n9391_0[2]),.din(n9391));
	jspl jspl_w_n9392_0(.douta(w_n9392_0[0]),.doutb(w_n9392_0[1]),.din(n9392));
	jspl jspl_w_n9396_0(.douta(w_n9396_0[0]),.doutb(w_n9396_0[1]),.din(n9396));
	jspl jspl_w_n9397_0(.douta(w_n9397_0[0]),.doutb(w_n9397_0[1]),.din(n9397));
	jspl3 jspl3_w_n9399_0(.douta(w_n9399_0[0]),.doutb(w_n9399_0[1]),.doutc(w_n9399_0[2]),.din(n9399));
	jspl jspl_w_n9400_0(.douta(w_n9400_0[0]),.doutb(w_n9400_0[1]),.din(n9400));
	jspl jspl_w_n9404_0(.douta(w_n9404_0[0]),.doutb(w_n9404_0[1]),.din(n9404));
	jspl3 jspl3_w_n9406_0(.douta(w_n9406_0[0]),.doutb(w_n9406_0[1]),.doutc(w_n9406_0[2]),.din(n9406));
	jspl jspl_w_n9407_0(.douta(w_n9407_0[0]),.doutb(w_n9407_0[1]),.din(n9407));
	jspl jspl_w_n9411_0(.douta(w_n9411_0[0]),.doutb(w_n9411_0[1]),.din(n9411));
	jspl jspl_w_n9412_0(.douta(w_n9412_0[0]),.doutb(w_n9412_0[1]),.din(n9412));
	jspl3 jspl3_w_n9414_0(.douta(w_n9414_0[0]),.doutb(w_n9414_0[1]),.doutc(w_n9414_0[2]),.din(n9414));
	jspl jspl_w_n9415_0(.douta(w_n9415_0[0]),.doutb(w_n9415_0[1]),.din(n9415));
	jspl jspl_w_n9419_0(.douta(w_n9419_0[0]),.doutb(w_n9419_0[1]),.din(n9419));
	jspl jspl_w_n9420_0(.douta(w_n9420_0[0]),.doutb(w_n9420_0[1]),.din(n9420));
	jspl3 jspl3_w_n9422_0(.douta(w_n9422_0[0]),.doutb(w_n9422_0[1]),.doutc(w_n9422_0[2]),.din(n9422));
	jspl jspl_w_n9423_0(.douta(w_n9423_0[0]),.doutb(w_n9423_0[1]),.din(n9423));
	jspl jspl_w_n9427_0(.douta(w_n9427_0[0]),.doutb(w_n9427_0[1]),.din(n9427));
	jspl jspl_w_n9428_0(.douta(w_n9428_0[0]),.doutb(w_n9428_0[1]),.din(n9428));
	jspl3 jspl3_w_n9430_0(.douta(w_n9430_0[0]),.doutb(w_n9430_0[1]),.doutc(w_n9430_0[2]),.din(n9430));
	jspl jspl_w_n9431_0(.douta(w_n9431_0[0]),.doutb(w_n9431_0[1]),.din(n9431));
	jspl jspl_w_n9435_0(.douta(w_n9435_0[0]),.doutb(w_n9435_0[1]),.din(n9435));
	jspl jspl_w_n9436_0(.douta(w_n9436_0[0]),.doutb(w_n9436_0[1]),.din(n9436));
	jspl3 jspl3_w_n9438_0(.douta(w_n9438_0[0]),.doutb(w_n9438_0[1]),.doutc(w_n9438_0[2]),.din(n9438));
	jspl jspl_w_n9439_0(.douta(w_n9439_0[0]),.doutb(w_n9439_0[1]),.din(n9439));
	jspl jspl_w_n9443_0(.douta(w_n9443_0[0]),.doutb(w_n9443_0[1]),.din(n9443));
	jspl jspl_w_n9444_0(.douta(w_n9444_0[0]),.doutb(w_n9444_0[1]),.din(n9444));
	jspl3 jspl3_w_n9446_0(.douta(w_n9446_0[0]),.doutb(w_n9446_0[1]),.doutc(w_n9446_0[2]),.din(n9446));
	jspl jspl_w_n9447_0(.douta(w_n9447_0[0]),.doutb(w_n9447_0[1]),.din(n9447));
	jspl jspl_w_n9450_0(.douta(w_n9450_0[0]),.doutb(w_n9450_0[1]),.din(n9450));
	jspl3 jspl3_w_n9453_0(.douta(w_n9453_0[0]),.doutb(w_n9453_0[1]),.doutc(w_n9453_0[2]),.din(n9453));
	jspl jspl_w_n9454_0(.douta(w_n9454_0[0]),.doutb(w_n9454_0[1]),.din(n9454));
	jspl jspl_w_n9458_0(.douta(w_n9458_0[0]),.doutb(w_n9458_0[1]),.din(n9458));
	jspl jspl_w_n9459_0(.douta(w_n9459_0[0]),.doutb(w_n9459_0[1]),.din(n9459));
	jspl3 jspl3_w_n9461_0(.douta(w_n9461_0[0]),.doutb(w_n9461_0[1]),.doutc(w_n9461_0[2]),.din(n9461));
	jspl jspl_w_n9462_0(.douta(w_n9462_0[0]),.doutb(w_n9462_0[1]),.din(n9462));
	jspl jspl_w_n9466_0(.douta(w_n9466_0[0]),.doutb(w_n9466_0[1]),.din(n9466));
	jspl3 jspl3_w_n9468_0(.douta(w_n9468_0[0]),.doutb(w_n9468_0[1]),.doutc(w_n9468_0[2]),.din(n9468));
	jspl jspl_w_n9469_0(.douta(w_n9469_0[0]),.doutb(w_n9469_0[1]),.din(n9469));
	jspl jspl_w_n9473_0(.douta(w_n9473_0[0]),.doutb(w_n9473_0[1]),.din(n9473));
	jspl jspl_w_n9474_0(.douta(w_n9474_0[0]),.doutb(w_n9474_0[1]),.din(n9474));
	jspl3 jspl3_w_n9476_0(.douta(w_n9476_0[0]),.doutb(w_n9476_0[1]),.doutc(w_n9476_0[2]),.din(n9476));
	jspl jspl_w_n9477_0(.douta(w_n9477_0[0]),.doutb(w_n9477_0[1]),.din(n9477));
	jspl jspl_w_n9481_0(.douta(w_n9481_0[0]),.doutb(w_n9481_0[1]),.din(n9481));
	jspl3 jspl3_w_n9483_0(.douta(w_n9483_0[0]),.doutb(w_n9483_0[1]),.doutc(w_n9483_0[2]),.din(n9483));
	jspl jspl_w_n9484_0(.douta(w_n9484_0[0]),.doutb(w_n9484_0[1]),.din(n9484));
	jspl3 jspl3_w_n9488_0(.douta(w_n9488_0[0]),.doutb(w_n9488_0[1]),.doutc(w_n9488_0[2]),.din(n9488));
	jspl3 jspl3_w_n9490_0(.douta(w_n9490_0[0]),.doutb(w_n9490_0[1]),.doutc(w_n9490_0[2]),.din(n9490));
	jspl jspl_w_n9491_0(.douta(w_n9491_0[0]),.doutb(w_n9491_0[1]),.din(n9491));
	jspl jspl_w_n9495_0(.douta(w_n9495_0[0]),.doutb(w_n9495_0[1]),.din(n9495));
	jspl jspl_w_n9496_0(.douta(w_n9496_0[0]),.doutb(w_n9496_0[1]),.din(n9496));
	jspl3 jspl3_w_n9498_0(.douta(w_n9498_0[0]),.doutb(w_n9498_0[1]),.doutc(w_n9498_0[2]),.din(n9498));
	jspl jspl_w_n9499_0(.douta(w_n9499_0[0]),.doutb(w_n9499_0[1]),.din(n9499));
	jspl jspl_w_n9503_0(.douta(w_n9503_0[0]),.doutb(w_n9503_0[1]),.din(n9503));
	jspl jspl_w_n9504_0(.douta(w_n9504_0[0]),.doutb(w_n9504_0[1]),.din(n9504));
	jspl3 jspl3_w_n9506_0(.douta(w_n9506_0[0]),.doutb(w_n9506_0[1]),.doutc(w_n9506_0[2]),.din(n9506));
	jspl jspl_w_n9507_0(.douta(w_n9507_0[0]),.doutb(w_n9507_0[1]),.din(n9507));
	jspl jspl_w_n9511_0(.douta(w_n9511_0[0]),.doutb(w_n9511_0[1]),.din(n9511));
	jspl3 jspl3_w_n9513_0(.douta(w_n9513_0[0]),.doutb(w_n9513_0[1]),.doutc(w_n9513_0[2]),.din(n9513));
	jspl jspl_w_n9514_0(.douta(w_n9514_0[0]),.doutb(w_n9514_0[1]),.din(n9514));
	jspl jspl_w_n9518_0(.douta(w_n9518_0[0]),.doutb(w_n9518_0[1]),.din(n9518));
	jspl jspl_w_n9519_0(.douta(w_n9519_0[0]),.doutb(w_n9519_0[1]),.din(n9519));
	jspl3 jspl3_w_n9521_0(.douta(w_n9521_0[0]),.doutb(w_n9521_0[1]),.doutc(w_n9521_0[2]),.din(n9521));
	jspl jspl_w_n9522_0(.douta(w_n9522_0[0]),.doutb(w_n9522_0[1]),.din(n9522));
	jspl jspl_w_n9526_0(.douta(w_n9526_0[0]),.doutb(w_n9526_0[1]),.din(n9526));
	jspl3 jspl3_w_n9528_0(.douta(w_n9528_0[0]),.doutb(w_n9528_0[1]),.doutc(w_n9528_0[2]),.din(n9528));
	jspl jspl_w_n9529_0(.douta(w_n9529_0[0]),.doutb(w_n9529_0[1]),.din(n9529));
	jspl jspl_w_n9533_0(.douta(w_n9533_0[0]),.doutb(w_n9533_0[1]),.din(n9533));
	jspl jspl_w_n9534_0(.douta(w_n9534_0[0]),.doutb(w_n9534_0[1]),.din(n9534));
	jspl3 jspl3_w_n9536_0(.douta(w_n9536_0[0]),.doutb(w_n9536_0[1]),.doutc(w_n9536_0[2]),.din(n9536));
	jspl jspl_w_n9537_0(.douta(w_n9537_0[0]),.doutb(w_n9537_0[1]),.din(n9537));
	jspl jspl_w_n9541_0(.douta(w_n9541_0[0]),.doutb(w_n9541_0[1]),.din(n9541));
	jspl3 jspl3_w_n9543_0(.douta(w_n9543_0[0]),.doutb(w_n9543_0[1]),.doutc(w_n9543_0[2]),.din(n9543));
	jspl jspl_w_n9544_0(.douta(w_n9544_0[0]),.doutb(w_n9544_0[1]),.din(n9544));
	jspl jspl_w_n9548_0(.douta(w_n9548_0[0]),.doutb(w_n9548_0[1]),.din(n9548));
	jspl jspl_w_n9549_0(.douta(w_n9549_0[0]),.doutb(w_n9549_0[1]),.din(n9549));
	jspl3 jspl3_w_n9551_0(.douta(w_n9551_0[0]),.doutb(w_n9551_0[1]),.doutc(w_n9551_0[2]),.din(n9551));
	jspl jspl_w_n9552_0(.douta(w_n9552_0[0]),.doutb(w_n9552_0[1]),.din(n9552));
	jspl jspl_w_n9556_0(.douta(w_n9556_0[0]),.doutb(w_n9556_0[1]),.din(n9556));
	jspl3 jspl3_w_n9558_0(.douta(w_n9558_0[0]),.doutb(w_n9558_0[1]),.doutc(w_n9558_0[2]),.din(n9558));
	jspl jspl_w_n9559_0(.douta(w_n9559_0[0]),.doutb(w_n9559_0[1]),.din(n9559));
	jspl jspl_w_n9563_0(.douta(w_n9563_0[0]),.doutb(w_n9563_0[1]),.din(n9563));
	jspl3 jspl3_w_n9565_0(.douta(w_n9565_0[0]),.doutb(w_n9565_0[1]),.doutc(w_n9565_0[2]),.din(n9565));
	jspl jspl_w_n9566_0(.douta(w_n9566_0[0]),.doutb(w_n9566_0[1]),.din(n9566));
	jspl jspl_w_n9570_0(.douta(w_n9570_0[0]),.doutb(w_n9570_0[1]),.din(n9570));
	jspl3 jspl3_w_n9572_0(.douta(w_n9572_0[0]),.doutb(w_n9572_0[1]),.doutc(w_n9572_0[2]),.din(n9572));
	jspl jspl_w_n9573_0(.douta(w_n9573_0[0]),.doutb(w_n9573_0[1]),.din(n9573));
	jspl jspl_w_n9577_0(.douta(w_n9577_0[0]),.doutb(w_n9577_0[1]),.din(n9577));
	jspl jspl_w_n9578_0(.douta(w_n9578_0[0]),.doutb(w_n9578_0[1]),.din(n9578));
	jspl3 jspl3_w_n9580_0(.douta(w_n9580_0[0]),.doutb(w_n9580_0[1]),.doutc(w_n9580_0[2]),.din(n9580));
	jspl jspl_w_n9581_0(.douta(w_n9581_0[0]),.doutb(w_n9581_0[1]),.din(n9581));
	jspl jspl_w_n9585_0(.douta(w_n9585_0[0]),.doutb(w_n9585_0[1]),.din(n9585));
	jspl jspl_w_n9586_0(.douta(w_n9586_0[0]),.doutb(w_n9586_0[1]),.din(n9586));
	jspl3 jspl3_w_n9588_0(.douta(w_n9588_0[0]),.doutb(w_n9588_0[1]),.doutc(w_n9588_0[2]),.din(n9588));
	jspl jspl_w_n9589_0(.douta(w_n9589_0[0]),.doutb(w_n9589_0[1]),.din(n9589));
	jspl jspl_w_n9593_0(.douta(w_n9593_0[0]),.doutb(w_n9593_0[1]),.din(n9593));
	jspl jspl_w_n9594_0(.douta(w_n9594_0[0]),.doutb(w_n9594_0[1]),.din(n9594));
	jspl3 jspl3_w_n9596_0(.douta(w_n9596_0[0]),.doutb(w_n9596_0[1]),.doutc(w_n9596_0[2]),.din(n9596));
	jspl jspl_w_n9597_0(.douta(w_n9597_0[0]),.doutb(w_n9597_0[1]),.din(n9597));
	jspl jspl_w_n9601_0(.douta(w_n9601_0[0]),.doutb(w_n9601_0[1]),.din(n9601));
	jspl3 jspl3_w_n9603_0(.douta(w_n9603_0[0]),.doutb(w_n9603_0[1]),.doutc(w_n9603_0[2]),.din(n9603));
	jspl jspl_w_n9604_0(.douta(w_n9604_0[0]),.doutb(w_n9604_0[1]),.din(n9604));
	jspl jspl_w_n9608_0(.douta(w_n9608_0[0]),.doutb(w_n9608_0[1]),.din(n9608));
	jspl jspl_w_n9609_0(.douta(w_n9609_0[0]),.doutb(w_n9609_0[1]),.din(n9609));
	jspl3 jspl3_w_n9611_0(.douta(w_n9611_0[0]),.doutb(w_n9611_0[1]),.doutc(w_n9611_0[2]),.din(n9611));
	jspl jspl_w_n9612_0(.douta(w_n9612_0[0]),.doutb(w_n9612_0[1]),.din(n9612));
	jspl jspl_w_n9616_0(.douta(w_n9616_0[0]),.doutb(w_n9616_0[1]),.din(n9616));
	jspl jspl_w_n9617_0(.douta(w_n9617_0[0]),.doutb(w_n9617_0[1]),.din(n9617));
	jspl3 jspl3_w_n9619_0(.douta(w_n9619_0[0]),.doutb(w_n9619_0[1]),.doutc(w_n9619_0[2]),.din(n9619));
	jspl jspl_w_n9620_0(.douta(w_n9620_0[0]),.doutb(w_n9620_0[1]),.din(n9620));
	jspl jspl_w_n9624_0(.douta(w_n9624_0[0]),.doutb(w_n9624_0[1]),.din(n9624));
	jspl jspl_w_n9625_0(.douta(w_n9625_0[0]),.doutb(w_n9625_0[1]),.din(n9625));
	jspl3 jspl3_w_n9627_0(.douta(w_n9627_0[0]),.doutb(w_n9627_0[1]),.doutc(w_n9627_0[2]),.din(n9627));
	jspl jspl_w_n9628_0(.douta(w_n9628_0[0]),.doutb(w_n9628_0[1]),.din(n9628));
	jspl jspl_w_n9632_0(.douta(w_n9632_0[0]),.doutb(w_n9632_0[1]),.din(n9632));
	jspl3 jspl3_w_n9634_0(.douta(w_n9634_0[0]),.doutb(w_n9634_0[1]),.doutc(w_n9634_0[2]),.din(n9634));
	jspl jspl_w_n9635_0(.douta(w_n9635_0[0]),.doutb(w_n9635_0[1]),.din(n9635));
	jspl3 jspl3_w_n9639_0(.douta(w_n9639_0[0]),.doutb(w_n9639_0[1]),.doutc(w_n9639_0[2]),.din(n9639));
	jspl jspl_w_n9641_0(.douta(w_n9641_0[0]),.doutb(w_n9641_0[1]),.din(n9641));
	jspl3 jspl3_w_n9642_0(.douta(w_n9642_0[0]),.doutb(w_n9642_0[1]),.doutc(w_n9642_0[2]),.din(n9642));
	jspl jspl_w_n9642_1(.douta(w_n9642_1[0]),.doutb(w_n9642_1[1]),.din(w_n9642_0[0]));
	jspl3 jspl3_w_n9643_0(.douta(w_n9643_0[0]),.doutb(w_n9643_0[1]),.doutc(w_n9643_0[2]),.din(n9643));
	jspl jspl_w_n9646_0(.douta(w_n9646_0[0]),.doutb(w_n9646_0[1]),.din(n9646));
	jspl jspl_w_n9647_0(.douta(w_n9647_0[0]),.doutb(w_n9647_0[1]),.din(n9647));
	jspl jspl_w_n9648_0(.douta(w_n9648_0[0]),.doutb(w_n9648_0[1]),.din(n9648));
	jspl jspl_w_n9649_0(.douta(w_n9649_0[0]),.doutb(w_n9649_0[1]),.din(n9649));
	jspl jspl_w_n9676_0(.douta(w_n9676_0[0]),.doutb(w_n9676_0[1]),.din(n9676));
	jspl jspl_w_n9693_0(.douta(w_n9693_0[0]),.doutb(w_n9693_0[1]),.din(n9693));
	jspl jspl_w_n9707_0(.douta(w_n9707_0[0]),.doutb(w_n9707_0[1]),.din(n9707));
	jspl jspl_w_n9732_0(.douta(w_n9732_0[0]),.doutb(w_n9732_0[1]),.din(n9732));
	jspl jspl_w_n9739_0(.douta(w_n9739_0[0]),.doutb(w_n9739_0[1]),.din(n9739));
	jspl jspl_w_n9753_0(.douta(w_n9753_0[0]),.doutb(w_n9753_0[1]),.din(n9753));
	jspl jspl_w_n9760_0(.douta(w_n9760_0[0]),.doutb(w_n9760_0[1]),.din(n9760));
	jspl jspl_w_n9767_0(.douta(w_n9767_0[0]),.doutb(w_n9767_0[1]),.din(n9767));
	jspl jspl_w_n9774_0(.douta(w_n9774_0[0]),.doutb(w_n9774_0[1]),.din(n9774));
	jspl jspl_w_n9778_0(.douta(w_n9778_0[0]),.doutb(w_n9778_0[1]),.din(n9778));
	jspl jspl_w_n9782_0(.douta(w_n9782_0[0]),.doutb(w_n9782_0[1]),.din(n9782));
	jspl jspl_w_n9795_0(.douta(w_n9795_0[0]),.doutb(w_n9795_0[1]),.din(n9795));
	jspl jspl_w_n9808_0(.douta(w_n9808_0[0]),.doutb(w_n9808_0[1]),.din(n9808));
	jspl jspl_w_n9814_0(.douta(w_n9814_0[0]),.doutb(w_n9814_0[1]),.din(n9814));
	jspl jspl_w_n9815_0(.douta(w_n9815_0[0]),.doutb(w_n9815_0[1]),.din(n9815));
	jspl jspl_w_n9816_0(.douta(w_n9816_0[0]),.doutb(w_n9816_0[1]),.din(n9816));
	jspl jspl_w_n9819_0(.douta(w_n9819_0[0]),.doutb(w_n9819_0[1]),.din(n9819));
	jspl jspl_w_n9820_0(.douta(w_n9820_0[0]),.doutb(w_n9820_0[1]),.din(n9820));
	jspl jspl_w_n9822_0(.douta(w_n9822_0[0]),.doutb(w_n9822_0[1]),.din(n9822));
	jspl jspl_w_n9824_0(.douta(w_n9824_0[0]),.doutb(w_n9824_0[1]),.din(n9824));
	jspl jspl_w_n9825_0(.douta(w_n9825_0[0]),.doutb(w_n9825_0[1]),.din(n9825));
	jspl jspl_w_n9831_0(.douta(w_n9831_0[0]),.doutb(w_n9831_0[1]),.din(n9831));
	jspl3 jspl3_w_n9832_0(.douta(w_n9832_0[0]),.doutb(w_n9832_0[1]),.doutc(w_n9832_0[2]),.din(n9832));
	jspl3 jspl3_w_n9832_1(.douta(w_n9832_1[0]),.doutb(w_n9832_1[1]),.doutc(w_n9832_1[2]),.din(w_n9832_0[0]));
	jspl3 jspl3_w_n9832_2(.douta(w_n9832_2[0]),.doutb(w_n9832_2[1]),.doutc(w_n9832_2[2]),.din(w_n9832_0[1]));
	jspl3 jspl3_w_n9832_3(.douta(w_n9832_3[0]),.doutb(w_n9832_3[1]),.doutc(w_n9832_3[2]),.din(w_n9832_0[2]));
	jspl3 jspl3_w_n9832_4(.douta(w_n9832_4[0]),.doutb(w_n9832_4[1]),.doutc(w_n9832_4[2]),.din(w_n9832_1[0]));
	jspl3 jspl3_w_n9832_5(.douta(w_n9832_5[0]),.doutb(w_n9832_5[1]),.doutc(w_n9832_5[2]),.din(w_n9832_1[1]));
	jspl3 jspl3_w_n9832_6(.douta(w_n9832_6[0]),.doutb(w_n9832_6[1]),.doutc(w_n9832_6[2]),.din(w_n9832_1[2]));
	jspl3 jspl3_w_n9832_7(.douta(w_n9832_7[0]),.doutb(w_n9832_7[1]),.doutc(w_n9832_7[2]),.din(w_n9832_2[0]));
	jspl3 jspl3_w_n9832_8(.douta(w_n9832_8[0]),.doutb(w_n9832_8[1]),.doutc(w_n9832_8[2]),.din(w_n9832_2[1]));
	jspl3 jspl3_w_n9832_9(.douta(w_n9832_9[0]),.doutb(w_n9832_9[1]),.doutc(w_n9832_9[2]),.din(w_n9832_2[2]));
	jspl3 jspl3_w_n9832_10(.douta(w_n9832_10[0]),.doutb(w_n9832_10[1]),.doutc(w_n9832_10[2]),.din(w_n9832_3[0]));
	jspl3 jspl3_w_n9832_11(.douta(w_n9832_11[0]),.doutb(w_n9832_11[1]),.doutc(w_n9832_11[2]),.din(w_n9832_3[1]));
	jspl3 jspl3_w_n9832_12(.douta(w_n9832_12[0]),.doutb(w_n9832_12[1]),.doutc(w_n9832_12[2]),.din(w_n9832_3[2]));
	jspl3 jspl3_w_n9832_13(.douta(w_n9832_13[0]),.doutb(w_n9832_13[1]),.doutc(w_n9832_13[2]),.din(w_n9832_4[0]));
	jspl3 jspl3_w_n9832_14(.douta(w_n9832_14[0]),.doutb(w_n9832_14[1]),.doutc(w_n9832_14[2]),.din(w_n9832_4[1]));
	jspl3 jspl3_w_n9832_15(.douta(w_n9832_15[0]),.doutb(w_n9832_15[1]),.doutc(w_n9832_15[2]),.din(w_n9832_4[2]));
	jspl3 jspl3_w_n9832_16(.douta(w_n9832_16[0]),.doutb(w_n9832_16[1]),.doutc(w_n9832_16[2]),.din(w_n9832_5[0]));
	jspl3 jspl3_w_n9832_17(.douta(w_n9832_17[0]),.doutb(w_n9832_17[1]),.doutc(w_n9832_17[2]),.din(w_n9832_5[1]));
	jspl3 jspl3_w_n9832_18(.douta(w_n9832_18[0]),.doutb(w_n9832_18[1]),.doutc(w_n9832_18[2]),.din(w_n9832_5[2]));
	jspl3 jspl3_w_n9832_19(.douta(w_n9832_19[0]),.doutb(w_n9832_19[1]),.doutc(w_n9832_19[2]),.din(w_n9832_6[0]));
	jspl3 jspl3_w_n9832_20(.douta(w_n9832_20[0]),.doutb(w_n9832_20[1]),.doutc(w_n9832_20[2]),.din(w_n9832_6[1]));
	jspl3 jspl3_w_n9832_21(.douta(w_n9832_21[0]),.doutb(w_n9832_21[1]),.doutc(w_n9832_21[2]),.din(w_n9832_6[2]));
	jspl3 jspl3_w_n9832_22(.douta(w_n9832_22[0]),.doutb(w_n9832_22[1]),.doutc(w_n9832_22[2]),.din(w_n9832_7[0]));
	jspl3 jspl3_w_n9832_23(.douta(w_n9832_23[0]),.doutb(w_n9832_23[1]),.doutc(w_n9832_23[2]),.din(w_n9832_7[1]));
	jspl3 jspl3_w_n9832_24(.douta(w_n9832_24[0]),.doutb(w_n9832_24[1]),.doutc(w_n9832_24[2]),.din(w_n9832_7[2]));
	jspl3 jspl3_w_n9832_25(.douta(w_n9832_25[0]),.doutb(w_n9832_25[1]),.doutc(w_n9832_25[2]),.din(w_n9832_8[0]));
	jspl3 jspl3_w_n9832_26(.douta(w_n9832_26[0]),.doutb(w_n9832_26[1]),.doutc(w_n9832_26[2]),.din(w_n9832_8[1]));
	jspl3 jspl3_w_n9832_27(.douta(w_n9832_27[0]),.doutb(w_n9832_27[1]),.doutc(w_n9832_27[2]),.din(w_n9832_8[2]));
	jspl3 jspl3_w_n9832_28(.douta(w_n9832_28[0]),.doutb(w_n9832_28[1]),.doutc(w_n9832_28[2]),.din(w_n9832_9[0]));
	jspl3 jspl3_w_n9832_29(.douta(w_n9832_29[0]),.doutb(w_n9832_29[1]),.doutc(w_n9832_29[2]),.din(w_n9832_9[1]));
	jspl3 jspl3_w_n9832_30(.douta(w_n9832_30[0]),.doutb(w_n9832_30[1]),.doutc(w_n9832_30[2]),.din(w_n9832_9[2]));
	jspl3 jspl3_w_n9832_31(.douta(w_n9832_31[0]),.doutb(w_n9832_31[1]),.doutc(w_n9832_31[2]),.din(w_n9832_10[0]));
	jspl3 jspl3_w_n9832_32(.douta(w_n9832_32[0]),.doutb(w_n9832_32[1]),.doutc(w_n9832_32[2]),.din(w_n9832_10[1]));
	jspl3 jspl3_w_n9832_33(.douta(w_n9832_33[0]),.doutb(w_n9832_33[1]),.doutc(w_n9832_33[2]),.din(w_n9832_10[2]));
	jspl3 jspl3_w_n9832_34(.douta(w_n9832_34[0]),.doutb(w_n9832_34[1]),.doutc(w_n9832_34[2]),.din(w_n9832_11[0]));
	jspl3 jspl3_w_n9832_35(.douta(w_n9832_35[0]),.doutb(w_n9832_35[1]),.doutc(w_n9832_35[2]),.din(w_n9832_11[1]));
	jspl3 jspl3_w_n9832_36(.douta(w_n9832_36[0]),.doutb(w_n9832_36[1]),.doutc(w_n9832_36[2]),.din(w_n9832_11[2]));
	jspl3 jspl3_w_n9832_37(.douta(w_n9832_37[0]),.doutb(w_n9832_37[1]),.doutc(w_n9832_37[2]),.din(w_n9832_12[0]));
	jspl3 jspl3_w_n9832_38(.douta(w_n9832_38[0]),.doutb(w_n9832_38[1]),.doutc(w_n9832_38[2]),.din(w_n9832_12[1]));
	jspl3 jspl3_w_n9832_39(.douta(w_n9832_39[0]),.doutb(w_n9832_39[1]),.doutc(w_n9832_39[2]),.din(w_n9832_12[2]));
	jspl3 jspl3_w_n9832_40(.douta(w_n9832_40[0]),.doutb(w_n9832_40[1]),.doutc(w_n9832_40[2]),.din(w_n9832_13[0]));
	jspl3 jspl3_w_n9832_41(.douta(w_n9832_41[0]),.doutb(w_n9832_41[1]),.doutc(w_n9832_41[2]),.din(w_n9832_13[1]));
	jspl3 jspl3_w_n9832_42(.douta(w_n9832_42[0]),.doutb(w_n9832_42[1]),.doutc(w_n9832_42[2]),.din(w_n9832_13[2]));
	jspl3 jspl3_w_n9832_43(.douta(w_n9832_43[0]),.doutb(w_n9832_43[1]),.doutc(w_n9832_43[2]),.din(w_n9832_14[0]));
	jspl3 jspl3_w_n9832_44(.douta(w_n9832_44[0]),.doutb(w_n9832_44[1]),.doutc(w_n9832_44[2]),.din(w_n9832_14[1]));
	jspl3 jspl3_w_n9832_45(.douta(w_n9832_45[0]),.doutb(w_n9832_45[1]),.doutc(w_n9832_45[2]),.din(w_n9832_14[2]));
	jspl3 jspl3_w_n9832_46(.douta(w_n9832_46[0]),.doutb(w_n9832_46[1]),.doutc(w_n9832_46[2]),.din(w_n9832_15[0]));
	jspl3 jspl3_w_n9832_47(.douta(w_n9832_47[0]),.doutb(w_n9832_47[1]),.doutc(w_n9832_47[2]),.din(w_n9832_15[1]));
	jspl3 jspl3_w_n9832_48(.douta(w_n9832_48[0]),.doutb(w_n9832_48[1]),.doutc(w_n9832_48[2]),.din(w_n9832_15[2]));
	jspl jspl_w_n9832_49(.douta(w_n9832_49[0]),.doutb(w_n9832_49[1]),.din(w_n9832_16[0]));
	jspl3 jspl3_w_n9834_0(.douta(w_n9834_0[0]),.doutb(w_n9834_0[1]),.doutc(w_n9834_0[2]),.din(n9834));
	jspl3 jspl3_w_n9834_1(.douta(w_n9834_1[0]),.doutb(w_n9834_1[1]),.doutc(w_n9834_1[2]),.din(w_n9834_0[0]));
	jspl jspl_w_n9835_0(.douta(w_n9835_0[0]),.doutb(w_n9835_0[1]),.din(n9835));
	jspl3 jspl3_w_n9836_0(.douta(w_n9836_0[0]),.doutb(w_n9836_0[1]),.doutc(w_n9836_0[2]),.din(n9836));
	jspl jspl_w_n9837_0(.douta(w_n9837_0[0]),.doutb(w_n9837_0[1]),.din(n9837));
	jspl3 jspl3_w_n9839_0(.douta(w_n9839_0[0]),.doutb(w_n9839_0[1]),.doutc(w_n9839_0[2]),.din(n9839));
	jspl jspl_w_n9840_0(.douta(w_n9840_0[0]),.doutb(w_n9840_0[1]),.din(n9840));
	jspl3 jspl3_w_n9847_0(.douta(w_n9847_0[0]),.doutb(w_n9847_0[1]),.doutc(w_n9847_0[2]),.din(n9847));
	jspl jspl_w_n9848_0(.douta(w_n9848_0[0]),.doutb(w_n9848_0[1]),.din(n9848));
	jspl jspl_w_n9851_0(.douta(w_n9851_0[0]),.doutb(w_n9851_0[1]),.din(n9851));
	jspl3 jspl3_w_n9856_0(.douta(w_n9856_0[0]),.doutb(w_n9856_0[1]),.doutc(w_n9856_0[2]),.din(n9856));
	jspl3 jspl3_w_n9858_0(.douta(w_n9858_0[0]),.doutb(w_n9858_0[1]),.doutc(w_n9858_0[2]),.din(n9858));
	jspl jspl_w_n9859_0(.douta(w_n9859_0[0]),.doutb(w_n9859_0[1]),.din(n9859));
	jspl3 jspl3_w_n9863_0(.douta(w_n9863_0[0]),.doutb(w_n9863_0[1]),.doutc(w_n9863_0[2]),.din(n9863));
	jspl3 jspl3_w_n9866_0(.douta(w_n9866_0[0]),.doutb(w_n9866_0[1]),.doutc(w_n9866_0[2]),.din(n9866));
	jspl jspl_w_n9867_0(.douta(w_n9867_0[0]),.doutb(w_n9867_0[1]),.din(n9867));
	jspl3 jspl3_w_n9871_0(.douta(w_n9871_0[0]),.doutb(w_n9871_0[1]),.doutc(w_n9871_0[2]),.din(n9871));
	jspl3 jspl3_w_n9873_0(.douta(w_n9873_0[0]),.doutb(w_n9873_0[1]),.doutc(w_n9873_0[2]),.din(n9873));
	jspl jspl_w_n9874_0(.douta(w_n9874_0[0]),.doutb(w_n9874_0[1]),.din(n9874));
	jspl3 jspl3_w_n9878_0(.douta(w_n9878_0[0]),.doutb(w_n9878_0[1]),.doutc(w_n9878_0[2]),.din(n9878));
	jspl3 jspl3_w_n9880_0(.douta(w_n9880_0[0]),.doutb(w_n9880_0[1]),.doutc(w_n9880_0[2]),.din(n9880));
	jspl jspl_w_n9881_0(.douta(w_n9881_0[0]),.doutb(w_n9881_0[1]),.din(n9881));
	jspl3 jspl3_w_n9885_0(.douta(w_n9885_0[0]),.doutb(w_n9885_0[1]),.doutc(w_n9885_0[2]),.din(n9885));
	jspl3 jspl3_w_n9887_0(.douta(w_n9887_0[0]),.doutb(w_n9887_0[1]),.doutc(w_n9887_0[2]),.din(n9887));
	jspl jspl_w_n9888_0(.douta(w_n9888_0[0]),.doutb(w_n9888_0[1]),.din(n9888));
	jspl3 jspl3_w_n9892_0(.douta(w_n9892_0[0]),.doutb(w_n9892_0[1]),.doutc(w_n9892_0[2]),.din(n9892));
	jspl3 jspl3_w_n9895_0(.douta(w_n9895_0[0]),.doutb(w_n9895_0[1]),.doutc(w_n9895_0[2]),.din(n9895));
	jspl jspl_w_n9896_0(.douta(w_n9896_0[0]),.doutb(w_n9896_0[1]),.din(n9896));
	jspl3 jspl3_w_n9900_0(.douta(w_n9900_0[0]),.doutb(w_n9900_0[1]),.doutc(w_n9900_0[2]),.din(n9900));
	jspl3 jspl3_w_n9902_0(.douta(w_n9902_0[0]),.doutb(w_n9902_0[1]),.doutc(w_n9902_0[2]),.din(n9902));
	jspl jspl_w_n9903_0(.douta(w_n9903_0[0]),.doutb(w_n9903_0[1]),.din(n9903));
	jspl3 jspl3_w_n9907_0(.douta(w_n9907_0[0]),.doutb(w_n9907_0[1]),.doutc(w_n9907_0[2]),.din(n9907));
	jspl3 jspl3_w_n9909_0(.douta(w_n9909_0[0]),.doutb(w_n9909_0[1]),.doutc(w_n9909_0[2]),.din(n9909));
	jspl jspl_w_n9910_0(.douta(w_n9910_0[0]),.doutb(w_n9910_0[1]),.din(n9910));
	jspl3 jspl3_w_n9914_0(.douta(w_n9914_0[0]),.doutb(w_n9914_0[1]),.doutc(w_n9914_0[2]),.din(n9914));
	jspl3 jspl3_w_n9916_0(.douta(w_n9916_0[0]),.doutb(w_n9916_0[1]),.doutc(w_n9916_0[2]),.din(n9916));
	jspl jspl_w_n9917_0(.douta(w_n9917_0[0]),.doutb(w_n9917_0[1]),.din(n9917));
	jspl3 jspl3_w_n9921_0(.douta(w_n9921_0[0]),.doutb(w_n9921_0[1]),.doutc(w_n9921_0[2]),.din(n9921));
	jspl3 jspl3_w_n9923_0(.douta(w_n9923_0[0]),.doutb(w_n9923_0[1]),.doutc(w_n9923_0[2]),.din(n9923));
	jspl jspl_w_n9924_0(.douta(w_n9924_0[0]),.doutb(w_n9924_0[1]),.din(n9924));
	jspl3 jspl3_w_n9928_0(.douta(w_n9928_0[0]),.doutb(w_n9928_0[1]),.doutc(w_n9928_0[2]),.din(n9928));
	jspl3 jspl3_w_n9930_0(.douta(w_n9930_0[0]),.doutb(w_n9930_0[1]),.doutc(w_n9930_0[2]),.din(n9930));
	jspl jspl_w_n9931_0(.douta(w_n9931_0[0]),.doutb(w_n9931_0[1]),.din(n9931));
	jspl3 jspl3_w_n9934_0(.douta(w_n9934_0[0]),.doutb(w_n9934_0[1]),.doutc(w_n9934_0[2]),.din(n9934));
	jspl3 jspl3_w_n9938_0(.douta(w_n9938_0[0]),.doutb(w_n9938_0[1]),.doutc(w_n9938_0[2]),.din(n9938));
	jspl jspl_w_n9939_0(.douta(w_n9939_0[0]),.doutb(w_n9939_0[1]),.din(n9939));
	jspl3 jspl3_w_n9943_0(.douta(w_n9943_0[0]),.doutb(w_n9943_0[1]),.doutc(w_n9943_0[2]),.din(n9943));
	jspl3 jspl3_w_n9945_0(.douta(w_n9945_0[0]),.doutb(w_n9945_0[1]),.doutc(w_n9945_0[2]),.din(n9945));
	jspl jspl_w_n9946_0(.douta(w_n9946_0[0]),.doutb(w_n9946_0[1]),.din(n9946));
	jspl3 jspl3_w_n9950_0(.douta(w_n9950_0[0]),.doutb(w_n9950_0[1]),.doutc(w_n9950_0[2]),.din(n9950));
	jspl3 jspl3_w_n9953_0(.douta(w_n9953_0[0]),.doutb(w_n9953_0[1]),.doutc(w_n9953_0[2]),.din(n9953));
	jspl jspl_w_n9954_0(.douta(w_n9954_0[0]),.doutb(w_n9954_0[1]),.din(n9954));
	jspl3 jspl3_w_n9958_0(.douta(w_n9958_0[0]),.doutb(w_n9958_0[1]),.doutc(w_n9958_0[2]),.din(n9958));
	jspl3 jspl3_w_n9960_0(.douta(w_n9960_0[0]),.doutb(w_n9960_0[1]),.doutc(w_n9960_0[2]),.din(n9960));
	jspl jspl_w_n9961_0(.douta(w_n9961_0[0]),.doutb(w_n9961_0[1]),.din(n9961));
	jspl3 jspl3_w_n9965_0(.douta(w_n9965_0[0]),.doutb(w_n9965_0[1]),.doutc(w_n9965_0[2]),.din(n9965));
	jspl3 jspl3_w_n9968_0(.douta(w_n9968_0[0]),.doutb(w_n9968_0[1]),.doutc(w_n9968_0[2]),.din(n9968));
	jspl jspl_w_n9969_0(.douta(w_n9969_0[0]),.doutb(w_n9969_0[1]),.din(n9969));
	jspl3 jspl3_w_n9973_0(.douta(w_n9973_0[0]),.doutb(w_n9973_0[1]),.doutc(w_n9973_0[2]),.din(n9973));
	jspl3 jspl3_w_n9975_0(.douta(w_n9975_0[0]),.doutb(w_n9975_0[1]),.doutc(w_n9975_0[2]),.din(n9975));
	jspl jspl_w_n9976_0(.douta(w_n9976_0[0]),.doutb(w_n9976_0[1]),.din(n9976));
	jspl3 jspl3_w_n9980_0(.douta(w_n9980_0[0]),.doutb(w_n9980_0[1]),.doutc(w_n9980_0[2]),.din(n9980));
	jspl3 jspl3_w_n9982_0(.douta(w_n9982_0[0]),.doutb(w_n9982_0[1]),.doutc(w_n9982_0[2]),.din(n9982));
	jspl jspl_w_n9983_0(.douta(w_n9983_0[0]),.doutb(w_n9983_0[1]),.din(n9983));
	jspl3 jspl3_w_n9987_0(.douta(w_n9987_0[0]),.doutb(w_n9987_0[1]),.doutc(w_n9987_0[2]),.din(n9987));
	jspl3 jspl3_w_n9989_0(.douta(w_n9989_0[0]),.doutb(w_n9989_0[1]),.doutc(w_n9989_0[2]),.din(n9989));
	jspl jspl_w_n9990_0(.douta(w_n9990_0[0]),.doutb(w_n9990_0[1]),.din(n9990));
	jspl3 jspl3_w_n9994_0(.douta(w_n9994_0[0]),.doutb(w_n9994_0[1]),.doutc(w_n9994_0[2]),.din(n9994));
	jspl3 jspl3_w_n9997_0(.douta(w_n9997_0[0]),.doutb(w_n9997_0[1]),.doutc(w_n9997_0[2]),.din(n9997));
	jspl jspl_w_n9998_0(.douta(w_n9998_0[0]),.doutb(w_n9998_0[1]),.din(n9998));
	jspl3 jspl3_w_n10002_0(.douta(w_n10002_0[0]),.doutb(w_n10002_0[1]),.doutc(w_n10002_0[2]),.din(n10002));
	jspl3 jspl3_w_n10004_0(.douta(w_n10004_0[0]),.doutb(w_n10004_0[1]),.doutc(w_n10004_0[2]),.din(n10004));
	jspl jspl_w_n10005_0(.douta(w_n10005_0[0]),.doutb(w_n10005_0[1]),.din(n10005));
	jspl3 jspl3_w_n10009_0(.douta(w_n10009_0[0]),.doutb(w_n10009_0[1]),.doutc(w_n10009_0[2]),.din(n10009));
	jspl3 jspl3_w_n10012_0(.douta(w_n10012_0[0]),.doutb(w_n10012_0[1]),.doutc(w_n10012_0[2]),.din(n10012));
	jspl jspl_w_n10013_0(.douta(w_n10013_0[0]),.doutb(w_n10013_0[1]),.din(n10013));
	jspl3 jspl3_w_n10017_0(.douta(w_n10017_0[0]),.doutb(w_n10017_0[1]),.doutc(w_n10017_0[2]),.din(n10017));
	jspl3 jspl3_w_n10019_0(.douta(w_n10019_0[0]),.doutb(w_n10019_0[1]),.doutc(w_n10019_0[2]),.din(n10019));
	jspl jspl_w_n10020_0(.douta(w_n10020_0[0]),.doutb(w_n10020_0[1]),.din(n10020));
	jspl3 jspl3_w_n10024_0(.douta(w_n10024_0[0]),.doutb(w_n10024_0[1]),.doutc(w_n10024_0[2]),.din(n10024));
	jspl3 jspl3_w_n10027_0(.douta(w_n10027_0[0]),.doutb(w_n10027_0[1]),.doutc(w_n10027_0[2]),.din(n10027));
	jspl jspl_w_n10028_0(.douta(w_n10028_0[0]),.doutb(w_n10028_0[1]),.din(n10028));
	jspl3 jspl3_w_n10032_0(.douta(w_n10032_0[0]),.doutb(w_n10032_0[1]),.doutc(w_n10032_0[2]),.din(n10032));
	jspl3 jspl3_w_n10034_0(.douta(w_n10034_0[0]),.doutb(w_n10034_0[1]),.doutc(w_n10034_0[2]),.din(n10034));
	jspl jspl_w_n10035_0(.douta(w_n10035_0[0]),.doutb(w_n10035_0[1]),.din(n10035));
	jspl3 jspl3_w_n10039_0(.douta(w_n10039_0[0]),.doutb(w_n10039_0[1]),.doutc(w_n10039_0[2]),.din(n10039));
	jspl3 jspl3_w_n10042_0(.douta(w_n10042_0[0]),.doutb(w_n10042_0[1]),.doutc(w_n10042_0[2]),.din(n10042));
	jspl jspl_w_n10043_0(.douta(w_n10043_0[0]),.doutb(w_n10043_0[1]),.din(n10043));
	jspl3 jspl3_w_n10047_0(.douta(w_n10047_0[0]),.doutb(w_n10047_0[1]),.doutc(w_n10047_0[2]),.din(n10047));
	jspl3 jspl3_w_n10050_0(.douta(w_n10050_0[0]),.doutb(w_n10050_0[1]),.doutc(w_n10050_0[2]),.din(n10050));
	jspl jspl_w_n10051_0(.douta(w_n10051_0[0]),.doutb(w_n10051_0[1]),.din(n10051));
	jspl3 jspl3_w_n10055_0(.douta(w_n10055_0[0]),.doutb(w_n10055_0[1]),.doutc(w_n10055_0[2]),.din(n10055));
	jspl3 jspl3_w_n10058_0(.douta(w_n10058_0[0]),.doutb(w_n10058_0[1]),.doutc(w_n10058_0[2]),.din(n10058));
	jspl jspl_w_n10059_0(.douta(w_n10059_0[0]),.doutb(w_n10059_0[1]),.din(n10059));
	jspl3 jspl3_w_n10063_0(.douta(w_n10063_0[0]),.doutb(w_n10063_0[1]),.doutc(w_n10063_0[2]),.din(n10063));
	jspl3 jspl3_w_n10065_0(.douta(w_n10065_0[0]),.doutb(w_n10065_0[1]),.doutc(w_n10065_0[2]),.din(n10065));
	jspl jspl_w_n10066_0(.douta(w_n10066_0[0]),.doutb(w_n10066_0[1]),.din(n10066));
	jspl3 jspl3_w_n10070_0(.douta(w_n10070_0[0]),.doutb(w_n10070_0[1]),.doutc(w_n10070_0[2]),.din(n10070));
	jspl3 jspl3_w_n10072_0(.douta(w_n10072_0[0]),.doutb(w_n10072_0[1]),.doutc(w_n10072_0[2]),.din(n10072));
	jspl jspl_w_n10073_0(.douta(w_n10073_0[0]),.doutb(w_n10073_0[1]),.din(n10073));
	jspl3 jspl3_w_n10077_0(.douta(w_n10077_0[0]),.doutb(w_n10077_0[1]),.doutc(w_n10077_0[2]),.din(n10077));
	jspl3 jspl3_w_n10079_0(.douta(w_n10079_0[0]),.doutb(w_n10079_0[1]),.doutc(w_n10079_0[2]),.din(n10079));
	jspl jspl_w_n10080_0(.douta(w_n10080_0[0]),.doutb(w_n10080_0[1]),.din(n10080));
	jspl3 jspl3_w_n10084_0(.douta(w_n10084_0[0]),.doutb(w_n10084_0[1]),.doutc(w_n10084_0[2]),.din(n10084));
	jspl3 jspl3_w_n10087_0(.douta(w_n10087_0[0]),.doutb(w_n10087_0[1]),.doutc(w_n10087_0[2]),.din(n10087));
	jspl jspl_w_n10088_0(.douta(w_n10088_0[0]),.doutb(w_n10088_0[1]),.din(n10088));
	jspl3 jspl3_w_n10092_0(.douta(w_n10092_0[0]),.doutb(w_n10092_0[1]),.doutc(w_n10092_0[2]),.din(n10092));
	jspl3 jspl3_w_n10094_0(.douta(w_n10094_0[0]),.doutb(w_n10094_0[1]),.doutc(w_n10094_0[2]),.din(n10094));
	jspl jspl_w_n10095_0(.douta(w_n10095_0[0]),.doutb(w_n10095_0[1]),.din(n10095));
	jspl3 jspl3_w_n10099_0(.douta(w_n10099_0[0]),.doutb(w_n10099_0[1]),.doutc(w_n10099_0[2]),.din(n10099));
	jspl3 jspl3_w_n10101_0(.douta(w_n10101_0[0]),.doutb(w_n10101_0[1]),.doutc(w_n10101_0[2]),.din(n10101));
	jspl jspl_w_n10102_0(.douta(w_n10102_0[0]),.doutb(w_n10102_0[1]),.din(n10102));
	jspl3 jspl3_w_n10106_0(.douta(w_n10106_0[0]),.doutb(w_n10106_0[1]),.doutc(w_n10106_0[2]),.din(n10106));
	jspl3 jspl3_w_n10108_0(.douta(w_n10108_0[0]),.doutb(w_n10108_0[1]),.doutc(w_n10108_0[2]),.din(n10108));
	jspl jspl_w_n10109_0(.douta(w_n10109_0[0]),.doutb(w_n10109_0[1]),.din(n10109));
	jspl jspl_w_n10113_0(.douta(w_n10113_0[0]),.doutb(w_n10113_0[1]),.din(n10113));
	jspl jspl_w_n10114_0(.douta(w_n10114_0[0]),.doutb(w_n10114_0[1]),.din(n10114));
	jspl3 jspl3_w_n10116_0(.douta(w_n10116_0[0]),.doutb(w_n10116_0[1]),.doutc(w_n10116_0[2]),.din(n10116));
	jspl3 jspl3_w_n10119_0(.douta(w_n10119_0[0]),.doutb(w_n10119_0[1]),.doutc(w_n10119_0[2]),.din(n10119));
	jspl jspl_w_n10119_1(.douta(w_n10119_1[0]),.doutb(w_n10119_1[1]),.din(w_n10119_0[0]));
	jspl jspl_w_n10120_0(.douta(w_n10120_0[0]),.doutb(w_n10120_0[1]),.din(n10120));
	jspl jspl_w_n10123_0(.douta(w_n10123_0[0]),.doutb(w_n10123_0[1]),.din(n10123));
	jspl3 jspl3_w_n10125_0(.douta(w_n10125_0[0]),.doutb(w_n10125_0[1]),.doutc(w_n10125_0[2]),.din(n10125));
	jspl jspl_w_n10125_1(.douta(w_n10125_1[0]),.doutb(w_n10125_1[1]),.din(w_n10125_0[0]));
	jspl jspl_w_n10130_0(.douta(w_n10130_0[0]),.doutb(w_n10130_0[1]),.din(n10130));
	jspl jspl_w_n10132_0(.douta(w_n10132_0[0]),.doutb(w_n10132_0[1]),.din(n10132));
	jspl3 jspl3_w_n10134_0(.douta(w_n10134_0[0]),.doutb(w_n10134_0[1]),.doutc(w_n10134_0[2]),.din(n10134));
	jspl jspl_w_n10134_1(.douta(w_n10134_1[0]),.doutb(w_n10134_1[1]),.din(w_n10134_0[0]));
	jspl jspl_w_n10135_0(.douta(w_n10135_0[0]),.doutb(w_n10135_0[1]),.din(n10135));
	jspl3 jspl3_w_n10136_0(.douta(w_n10136_0[0]),.doutb(w_n10136_0[1]),.doutc(w_n10136_0[2]),.din(n10136));
	jspl jspl_w_n10137_0(.douta(w_n10137_0[0]),.doutb(w_n10137_0[1]),.din(n10137));
	jspl3 jspl3_w_n10139_0(.douta(w_n10139_0[0]),.doutb(w_n10139_0[1]),.doutc(w_n10139_0[2]),.din(n10139));
	jspl jspl_w_n10140_0(.douta(w_n10140_0[0]),.doutb(w_n10140_0[1]),.din(n10140));
	jspl jspl_w_n10188_0(.douta(w_n10188_0[0]),.doutb(w_n10188_0[1]),.din(n10188));
	jspl jspl_w_n10323_0(.douta(w_n10323_0[0]),.doutb(w_n10323_0[1]),.din(n10323));
	jspl3 jspl3_w_n10328_0(.douta(w_n10328_0[0]),.doutb(w_n10328_0[1]),.doutc(w_n10328_0[2]),.din(n10328));
	jspl3 jspl3_w_n10328_1(.douta(w_n10328_1[0]),.doutb(w_n10328_1[1]),.doutc(w_n10328_1[2]),.din(w_n10328_0[0]));
	jspl3 jspl3_w_n10328_2(.douta(w_n10328_2[0]),.doutb(w_n10328_2[1]),.doutc(w_n10328_2[2]),.din(w_n10328_0[1]));
	jspl3 jspl3_w_n10328_3(.douta(w_n10328_3[0]),.doutb(w_n10328_3[1]),.doutc(w_n10328_3[2]),.din(w_n10328_0[2]));
	jspl3 jspl3_w_n10328_4(.douta(w_n10328_4[0]),.doutb(w_n10328_4[1]),.doutc(w_n10328_4[2]),.din(w_n10328_1[0]));
	jspl3 jspl3_w_n10328_5(.douta(w_n10328_5[0]),.doutb(w_n10328_5[1]),.doutc(w_n10328_5[2]),.din(w_n10328_1[1]));
	jspl3 jspl3_w_n10328_6(.douta(w_n10328_6[0]),.doutb(w_n10328_6[1]),.doutc(w_n10328_6[2]),.din(w_n10328_1[2]));
	jspl3 jspl3_w_n10328_7(.douta(w_n10328_7[0]),.doutb(w_n10328_7[1]),.doutc(w_n10328_7[2]),.din(w_n10328_2[0]));
	jspl3 jspl3_w_n10328_8(.douta(w_n10328_8[0]),.doutb(w_n10328_8[1]),.doutc(w_n10328_8[2]),.din(w_n10328_2[1]));
	jspl3 jspl3_w_n10328_9(.douta(w_n10328_9[0]),.doutb(w_n10328_9[1]),.doutc(w_n10328_9[2]),.din(w_n10328_2[2]));
	jspl3 jspl3_w_n10328_10(.douta(w_n10328_10[0]),.doutb(w_n10328_10[1]),.doutc(w_n10328_10[2]),.din(w_n10328_3[0]));
	jspl3 jspl3_w_n10328_11(.douta(w_n10328_11[0]),.doutb(w_n10328_11[1]),.doutc(w_n10328_11[2]),.din(w_n10328_3[1]));
	jspl3 jspl3_w_n10328_12(.douta(w_n10328_12[0]),.doutb(w_n10328_12[1]),.doutc(w_n10328_12[2]),.din(w_n10328_3[2]));
	jspl3 jspl3_w_n10328_13(.douta(w_n10328_13[0]),.doutb(w_n10328_13[1]),.doutc(w_n10328_13[2]),.din(w_n10328_4[0]));
	jspl3 jspl3_w_n10328_14(.douta(w_n10328_14[0]),.doutb(w_n10328_14[1]),.doutc(w_n10328_14[2]),.din(w_n10328_4[1]));
	jspl3 jspl3_w_n10328_15(.douta(w_n10328_15[0]),.doutb(w_n10328_15[1]),.doutc(w_n10328_15[2]),.din(w_n10328_4[2]));
	jspl3 jspl3_w_n10328_16(.douta(w_n10328_16[0]),.doutb(w_n10328_16[1]),.doutc(w_n10328_16[2]),.din(w_n10328_5[0]));
	jspl3 jspl3_w_n10328_17(.douta(w_n10328_17[0]),.doutb(w_n10328_17[1]),.doutc(w_n10328_17[2]),.din(w_n10328_5[1]));
	jspl3 jspl3_w_n10328_18(.douta(w_n10328_18[0]),.doutb(w_n10328_18[1]),.doutc(w_n10328_18[2]),.din(w_n10328_5[2]));
	jspl3 jspl3_w_n10328_19(.douta(w_n10328_19[0]),.doutb(w_n10328_19[1]),.doutc(w_n10328_19[2]),.din(w_n10328_6[0]));
	jspl3 jspl3_w_n10328_20(.douta(w_n10328_20[0]),.doutb(w_n10328_20[1]),.doutc(w_n10328_20[2]),.din(w_n10328_6[1]));
	jspl3 jspl3_w_n10328_21(.douta(w_n10328_21[0]),.doutb(w_n10328_21[1]),.doutc(w_n10328_21[2]),.din(w_n10328_6[2]));
	jspl3 jspl3_w_n10328_22(.douta(w_n10328_22[0]),.doutb(w_n10328_22[1]),.doutc(w_n10328_22[2]),.din(w_n10328_7[0]));
	jspl3 jspl3_w_n10328_23(.douta(w_n10328_23[0]),.doutb(w_n10328_23[1]),.doutc(w_n10328_23[2]),.din(w_n10328_7[1]));
	jspl3 jspl3_w_n10328_24(.douta(w_n10328_24[0]),.doutb(w_n10328_24[1]),.doutc(w_n10328_24[2]),.din(w_n10328_7[2]));
	jspl3 jspl3_w_n10328_25(.douta(w_n10328_25[0]),.doutb(w_n10328_25[1]),.doutc(w_n10328_25[2]),.din(w_n10328_8[0]));
	jspl3 jspl3_w_n10328_26(.douta(w_n10328_26[0]),.doutb(w_n10328_26[1]),.doutc(w_n10328_26[2]),.din(w_n10328_8[1]));
	jspl3 jspl3_w_n10328_27(.douta(w_n10328_27[0]),.doutb(w_n10328_27[1]),.doutc(w_n10328_27[2]),.din(w_n10328_8[2]));
	jspl3 jspl3_w_n10328_28(.douta(w_n10328_28[0]),.doutb(w_n10328_28[1]),.doutc(w_n10328_28[2]),.din(w_n10328_9[0]));
	jspl3 jspl3_w_n10328_29(.douta(w_n10328_29[0]),.doutb(w_n10328_29[1]),.doutc(w_n10328_29[2]),.din(w_n10328_9[1]));
	jspl3 jspl3_w_n10328_30(.douta(w_n10328_30[0]),.doutb(w_n10328_30[1]),.doutc(w_n10328_30[2]),.din(w_n10328_9[2]));
	jspl jspl_w_n10329_0(.douta(w_n10329_0[0]),.doutb(w_n10329_0[1]),.din(n10329));
	jspl jspl_w_n10330_0(.douta(w_n10330_0[0]),.doutb(w_n10330_0[1]),.din(n10330));
	jspl3 jspl3_w_n10332_0(.douta(w_n10332_0[0]),.doutb(w_n10332_0[1]),.doutc(w_n10332_0[2]),.din(n10332));
	jspl jspl_w_n10333_0(.douta(w_n10333_0[0]),.doutb(w_n10333_0[1]),.din(n10333));
	jspl jspl_w_n10339_0(.douta(w_n10339_0[0]),.doutb(w_n10339_0[1]),.din(n10339));
	jspl jspl_w_n10340_0(.douta(w_n10340_0[0]),.doutb(w_n10340_0[1]),.din(n10340));
	jspl3 jspl3_w_n10342_0(.douta(w_n10342_0[0]),.doutb(w_n10342_0[1]),.doutc(w_n10342_0[2]),.din(n10342));
	jspl jspl_w_n10343_0(.douta(w_n10343_0[0]),.doutb(w_n10343_0[1]),.din(n10343));
	jspl jspl_w_n10347_0(.douta(w_n10347_0[0]),.doutb(w_n10347_0[1]),.din(n10347));
	jspl3 jspl3_w_n10349_0(.douta(w_n10349_0[0]),.doutb(w_n10349_0[1]),.doutc(w_n10349_0[2]),.din(n10349));
	jspl jspl_w_n10350_0(.douta(w_n10350_0[0]),.doutb(w_n10350_0[1]),.din(n10350));
	jspl jspl_w_n10354_0(.douta(w_n10354_0[0]),.doutb(w_n10354_0[1]),.din(n10354));
	jspl jspl_w_n10355_0(.douta(w_n10355_0[0]),.doutb(w_n10355_0[1]),.din(n10355));
	jspl3 jspl3_w_n10357_0(.douta(w_n10357_0[0]),.doutb(w_n10357_0[1]),.doutc(w_n10357_0[2]),.din(n10357));
	jspl jspl_w_n10358_0(.douta(w_n10358_0[0]),.doutb(w_n10358_0[1]),.din(n10358));
	jspl jspl_w_n10362_0(.douta(w_n10362_0[0]),.doutb(w_n10362_0[1]),.din(n10362));
	jspl3 jspl3_w_n10364_0(.douta(w_n10364_0[0]),.doutb(w_n10364_0[1]),.doutc(w_n10364_0[2]),.din(n10364));
	jspl jspl_w_n10365_0(.douta(w_n10365_0[0]),.doutb(w_n10365_0[1]),.din(n10365));
	jspl jspl_w_n10369_0(.douta(w_n10369_0[0]),.doutb(w_n10369_0[1]),.din(n10369));
	jspl jspl_w_n10370_0(.douta(w_n10370_0[0]),.doutb(w_n10370_0[1]),.din(n10370));
	jspl3 jspl3_w_n10372_0(.douta(w_n10372_0[0]),.doutb(w_n10372_0[1]),.doutc(w_n10372_0[2]),.din(n10372));
	jspl jspl_w_n10373_0(.douta(w_n10373_0[0]),.doutb(w_n10373_0[1]),.din(n10373));
	jspl jspl_w_n10377_0(.douta(w_n10377_0[0]),.doutb(w_n10377_0[1]),.din(n10377));
	jspl jspl_w_n10378_0(.douta(w_n10378_0[0]),.doutb(w_n10378_0[1]),.din(n10378));
	jspl3 jspl3_w_n10380_0(.douta(w_n10380_0[0]),.doutb(w_n10380_0[1]),.doutc(w_n10380_0[2]),.din(n10380));
	jspl jspl_w_n10381_0(.douta(w_n10381_0[0]),.doutb(w_n10381_0[1]),.din(n10381));
	jspl jspl_w_n10385_0(.douta(w_n10385_0[0]),.doutb(w_n10385_0[1]),.din(n10385));
	jspl jspl_w_n10386_0(.douta(w_n10386_0[0]),.doutb(w_n10386_0[1]),.din(n10386));
	jspl3 jspl3_w_n10388_0(.douta(w_n10388_0[0]),.doutb(w_n10388_0[1]),.doutc(w_n10388_0[2]),.din(n10388));
	jspl jspl_w_n10389_0(.douta(w_n10389_0[0]),.doutb(w_n10389_0[1]),.din(n10389));
	jspl jspl_w_n10393_0(.douta(w_n10393_0[0]),.doutb(w_n10393_0[1]),.din(n10393));
	jspl3 jspl3_w_n10395_0(.douta(w_n10395_0[0]),.doutb(w_n10395_0[1]),.doutc(w_n10395_0[2]),.din(n10395));
	jspl jspl_w_n10396_0(.douta(w_n10396_0[0]),.doutb(w_n10396_0[1]),.din(n10396));
	jspl jspl_w_n10400_0(.douta(w_n10400_0[0]),.doutb(w_n10400_0[1]),.din(n10400));
	jspl jspl_w_n10401_0(.douta(w_n10401_0[0]),.doutb(w_n10401_0[1]),.din(n10401));
	jspl3 jspl3_w_n10403_0(.douta(w_n10403_0[0]),.doutb(w_n10403_0[1]),.doutc(w_n10403_0[2]),.din(n10403));
	jspl jspl_w_n10404_0(.douta(w_n10404_0[0]),.doutb(w_n10404_0[1]),.din(n10404));
	jspl jspl_w_n10408_0(.douta(w_n10408_0[0]),.doutb(w_n10408_0[1]),.din(n10408));
	jspl jspl_w_n10409_0(.douta(w_n10409_0[0]),.doutb(w_n10409_0[1]),.din(n10409));
	jspl3 jspl3_w_n10411_0(.douta(w_n10411_0[0]),.doutb(w_n10411_0[1]),.doutc(w_n10411_0[2]),.din(n10411));
	jspl jspl_w_n10412_0(.douta(w_n10412_0[0]),.doutb(w_n10412_0[1]),.din(n10412));
	jspl jspl_w_n10416_0(.douta(w_n10416_0[0]),.doutb(w_n10416_0[1]),.din(n10416));
	jspl jspl_w_n10417_0(.douta(w_n10417_0[0]),.doutb(w_n10417_0[1]),.din(n10417));
	jspl3 jspl3_w_n10419_0(.douta(w_n10419_0[0]),.doutb(w_n10419_0[1]),.doutc(w_n10419_0[2]),.din(n10419));
	jspl jspl_w_n10420_0(.douta(w_n10420_0[0]),.doutb(w_n10420_0[1]),.din(n10420));
	jspl jspl_w_n10424_0(.douta(w_n10424_0[0]),.doutb(w_n10424_0[1]),.din(n10424));
	jspl jspl_w_n10425_0(.douta(w_n10425_0[0]),.doutb(w_n10425_0[1]),.din(n10425));
	jspl3 jspl3_w_n10427_0(.douta(w_n10427_0[0]),.doutb(w_n10427_0[1]),.doutc(w_n10427_0[2]),.din(n10427));
	jspl jspl_w_n10428_0(.douta(w_n10428_0[0]),.doutb(w_n10428_0[1]),.din(n10428));
	jspl jspl_w_n10432_0(.douta(w_n10432_0[0]),.doutb(w_n10432_0[1]),.din(n10432));
	jspl jspl_w_n10433_0(.douta(w_n10433_0[0]),.doutb(w_n10433_0[1]),.din(n10433));
	jspl3 jspl3_w_n10435_0(.douta(w_n10435_0[0]),.doutb(w_n10435_0[1]),.doutc(w_n10435_0[2]),.din(n10435));
	jspl jspl_w_n10436_0(.douta(w_n10436_0[0]),.doutb(w_n10436_0[1]),.din(n10436));
	jspl jspl_w_n10439_0(.douta(w_n10439_0[0]),.doutb(w_n10439_0[1]),.din(n10439));
	jspl3 jspl3_w_n10442_0(.douta(w_n10442_0[0]),.doutb(w_n10442_0[1]),.doutc(w_n10442_0[2]),.din(n10442));
	jspl jspl_w_n10443_0(.douta(w_n10443_0[0]),.doutb(w_n10443_0[1]),.din(n10443));
	jspl jspl_w_n10447_0(.douta(w_n10447_0[0]),.doutb(w_n10447_0[1]),.din(n10447));
	jspl jspl_w_n10448_0(.douta(w_n10448_0[0]),.doutb(w_n10448_0[1]),.din(n10448));
	jspl3 jspl3_w_n10450_0(.douta(w_n10450_0[0]),.doutb(w_n10450_0[1]),.doutc(w_n10450_0[2]),.din(n10450));
	jspl jspl_w_n10451_0(.douta(w_n10451_0[0]),.doutb(w_n10451_0[1]),.din(n10451));
	jspl jspl_w_n10455_0(.douta(w_n10455_0[0]),.doutb(w_n10455_0[1]),.din(n10455));
	jspl3 jspl3_w_n10457_0(.douta(w_n10457_0[0]),.doutb(w_n10457_0[1]),.doutc(w_n10457_0[2]),.din(n10457));
	jspl jspl_w_n10458_0(.douta(w_n10458_0[0]),.doutb(w_n10458_0[1]),.din(n10458));
	jspl jspl_w_n10462_0(.douta(w_n10462_0[0]),.doutb(w_n10462_0[1]),.din(n10462));
	jspl jspl_w_n10463_0(.douta(w_n10463_0[0]),.doutb(w_n10463_0[1]),.din(n10463));
	jspl3 jspl3_w_n10465_0(.douta(w_n10465_0[0]),.doutb(w_n10465_0[1]),.doutc(w_n10465_0[2]),.din(n10465));
	jspl jspl_w_n10466_0(.douta(w_n10466_0[0]),.doutb(w_n10466_0[1]),.din(n10466));
	jspl jspl_w_n10470_0(.douta(w_n10470_0[0]),.doutb(w_n10470_0[1]),.din(n10470));
	jspl3 jspl3_w_n10472_0(.douta(w_n10472_0[0]),.doutb(w_n10472_0[1]),.doutc(w_n10472_0[2]),.din(n10472));
	jspl jspl_w_n10473_0(.douta(w_n10473_0[0]),.doutb(w_n10473_0[1]),.din(n10473));
	jspl jspl_w_n10477_0(.douta(w_n10477_0[0]),.doutb(w_n10477_0[1]),.din(n10477));
	jspl jspl_w_n10478_0(.douta(w_n10478_0[0]),.doutb(w_n10478_0[1]),.din(n10478));
	jspl3 jspl3_w_n10480_0(.douta(w_n10480_0[0]),.doutb(w_n10480_0[1]),.doutc(w_n10480_0[2]),.din(n10480));
	jspl jspl_w_n10481_0(.douta(w_n10481_0[0]),.doutb(w_n10481_0[1]),.din(n10481));
	jspl jspl_w_n10485_0(.douta(w_n10485_0[0]),.doutb(w_n10485_0[1]),.din(n10485));
	jspl jspl_w_n10486_0(.douta(w_n10486_0[0]),.doutb(w_n10486_0[1]),.din(n10486));
	jspl3 jspl3_w_n10488_0(.douta(w_n10488_0[0]),.doutb(w_n10488_0[1]),.doutc(w_n10488_0[2]),.din(n10488));
	jspl jspl_w_n10489_0(.douta(w_n10489_0[0]),.doutb(w_n10489_0[1]),.din(n10489));
	jspl jspl_w_n10493_0(.douta(w_n10493_0[0]),.doutb(w_n10493_0[1]),.din(n10493));
	jspl jspl_w_n10494_0(.douta(w_n10494_0[0]),.doutb(w_n10494_0[1]),.din(n10494));
	jspl3 jspl3_w_n10496_0(.douta(w_n10496_0[0]),.doutb(w_n10496_0[1]),.doutc(w_n10496_0[2]),.din(n10496));
	jspl jspl_w_n10497_0(.douta(w_n10497_0[0]),.doutb(w_n10497_0[1]),.din(n10497));
	jspl jspl_w_n10501_0(.douta(w_n10501_0[0]),.doutb(w_n10501_0[1]),.din(n10501));
	jspl3 jspl3_w_n10503_0(.douta(w_n10503_0[0]),.doutb(w_n10503_0[1]),.doutc(w_n10503_0[2]),.din(n10503));
	jspl jspl_w_n10504_0(.douta(w_n10504_0[0]),.doutb(w_n10504_0[1]),.din(n10504));
	jspl jspl_w_n10508_0(.douta(w_n10508_0[0]),.doutb(w_n10508_0[1]),.din(n10508));
	jspl jspl_w_n10509_0(.douta(w_n10509_0[0]),.doutb(w_n10509_0[1]),.din(n10509));
	jspl3 jspl3_w_n10511_0(.douta(w_n10511_0[0]),.doutb(w_n10511_0[1]),.doutc(w_n10511_0[2]),.din(n10511));
	jspl jspl_w_n10512_0(.douta(w_n10512_0[0]),.doutb(w_n10512_0[1]),.din(n10512));
	jspl jspl_w_n10516_0(.douta(w_n10516_0[0]),.doutb(w_n10516_0[1]),.din(n10516));
	jspl3 jspl3_w_n10518_0(.douta(w_n10518_0[0]),.doutb(w_n10518_0[1]),.doutc(w_n10518_0[2]),.din(n10518));
	jspl jspl_w_n10519_0(.douta(w_n10519_0[0]),.doutb(w_n10519_0[1]),.din(n10519));
	jspl jspl_w_n10523_0(.douta(w_n10523_0[0]),.doutb(w_n10523_0[1]),.din(n10523));
	jspl jspl_w_n10524_0(.douta(w_n10524_0[0]),.doutb(w_n10524_0[1]),.din(n10524));
	jspl3 jspl3_w_n10526_0(.douta(w_n10526_0[0]),.doutb(w_n10526_0[1]),.doutc(w_n10526_0[2]),.din(n10526));
	jspl jspl_w_n10527_0(.douta(w_n10527_0[0]),.doutb(w_n10527_0[1]),.din(n10527));
	jspl jspl_w_n10531_0(.douta(w_n10531_0[0]),.doutb(w_n10531_0[1]),.din(n10531));
	jspl3 jspl3_w_n10533_0(.douta(w_n10533_0[0]),.doutb(w_n10533_0[1]),.doutc(w_n10533_0[2]),.din(n10533));
	jspl jspl_w_n10534_0(.douta(w_n10534_0[0]),.doutb(w_n10534_0[1]),.din(n10534));
	jspl jspl_w_n10538_0(.douta(w_n10538_0[0]),.doutb(w_n10538_0[1]),.din(n10538));
	jspl jspl_w_n10539_0(.douta(w_n10539_0[0]),.doutb(w_n10539_0[1]),.din(n10539));
	jspl3 jspl3_w_n10541_0(.douta(w_n10541_0[0]),.doutb(w_n10541_0[1]),.doutc(w_n10541_0[2]),.din(n10541));
	jspl jspl_w_n10542_0(.douta(w_n10542_0[0]),.doutb(w_n10542_0[1]),.din(n10542));
	jspl jspl_w_n10546_0(.douta(w_n10546_0[0]),.doutb(w_n10546_0[1]),.din(n10546));
	jspl3 jspl3_w_n10548_0(.douta(w_n10548_0[0]),.doutb(w_n10548_0[1]),.doutc(w_n10548_0[2]),.din(n10548));
	jspl jspl_w_n10549_0(.douta(w_n10549_0[0]),.doutb(w_n10549_0[1]),.din(n10549));
	jspl jspl_w_n10553_0(.douta(w_n10553_0[0]),.doutb(w_n10553_0[1]),.din(n10553));
	jspl3 jspl3_w_n10555_0(.douta(w_n10555_0[0]),.doutb(w_n10555_0[1]),.doutc(w_n10555_0[2]),.din(n10555));
	jspl jspl_w_n10556_0(.douta(w_n10556_0[0]),.doutb(w_n10556_0[1]),.din(n10556));
	jspl jspl_w_n10560_0(.douta(w_n10560_0[0]),.doutb(w_n10560_0[1]),.din(n10560));
	jspl3 jspl3_w_n10562_0(.douta(w_n10562_0[0]),.doutb(w_n10562_0[1]),.doutc(w_n10562_0[2]),.din(n10562));
	jspl jspl_w_n10563_0(.douta(w_n10563_0[0]),.doutb(w_n10563_0[1]),.din(n10563));
	jspl jspl_w_n10567_0(.douta(w_n10567_0[0]),.doutb(w_n10567_0[1]),.din(n10567));
	jspl jspl_w_n10568_0(.douta(w_n10568_0[0]),.doutb(w_n10568_0[1]),.din(n10568));
	jspl3 jspl3_w_n10570_0(.douta(w_n10570_0[0]),.doutb(w_n10570_0[1]),.doutc(w_n10570_0[2]),.din(n10570));
	jspl jspl_w_n10571_0(.douta(w_n10571_0[0]),.doutb(w_n10571_0[1]),.din(n10571));
	jspl jspl_w_n10575_0(.douta(w_n10575_0[0]),.doutb(w_n10575_0[1]),.din(n10575));
	jspl jspl_w_n10576_0(.douta(w_n10576_0[0]),.doutb(w_n10576_0[1]),.din(n10576));
	jspl3 jspl3_w_n10578_0(.douta(w_n10578_0[0]),.doutb(w_n10578_0[1]),.doutc(w_n10578_0[2]),.din(n10578));
	jspl jspl_w_n10579_0(.douta(w_n10579_0[0]),.doutb(w_n10579_0[1]),.din(n10579));
	jspl jspl_w_n10583_0(.douta(w_n10583_0[0]),.doutb(w_n10583_0[1]),.din(n10583));
	jspl jspl_w_n10584_0(.douta(w_n10584_0[0]),.doutb(w_n10584_0[1]),.din(n10584));
	jspl3 jspl3_w_n10586_0(.douta(w_n10586_0[0]),.doutb(w_n10586_0[1]),.doutc(w_n10586_0[2]),.din(n10586));
	jspl jspl_w_n10587_0(.douta(w_n10587_0[0]),.doutb(w_n10587_0[1]),.din(n10587));
	jspl jspl_w_n10591_0(.douta(w_n10591_0[0]),.doutb(w_n10591_0[1]),.din(n10591));
	jspl3 jspl3_w_n10593_0(.douta(w_n10593_0[0]),.doutb(w_n10593_0[1]),.doutc(w_n10593_0[2]),.din(n10593));
	jspl jspl_w_n10594_0(.douta(w_n10594_0[0]),.doutb(w_n10594_0[1]),.din(n10594));
	jspl jspl_w_n10598_0(.douta(w_n10598_0[0]),.doutb(w_n10598_0[1]),.din(n10598));
	jspl jspl_w_n10599_0(.douta(w_n10599_0[0]),.doutb(w_n10599_0[1]),.din(n10599));
	jspl3 jspl3_w_n10601_0(.douta(w_n10601_0[0]),.doutb(w_n10601_0[1]),.doutc(w_n10601_0[2]),.din(n10601));
	jspl jspl_w_n10602_0(.douta(w_n10602_0[0]),.doutb(w_n10602_0[1]),.din(n10602));
	jspl jspl_w_n10606_0(.douta(w_n10606_0[0]),.doutb(w_n10606_0[1]),.din(n10606));
	jspl jspl_w_n10607_0(.douta(w_n10607_0[0]),.doutb(w_n10607_0[1]),.din(n10607));
	jspl3 jspl3_w_n10609_0(.douta(w_n10609_0[0]),.doutb(w_n10609_0[1]),.doutc(w_n10609_0[2]),.din(n10609));
	jspl jspl_w_n10610_0(.douta(w_n10610_0[0]),.doutb(w_n10610_0[1]),.din(n10610));
	jspl jspl_w_n10635_0(.douta(w_n10635_0[0]),.doutb(w_n10635_0[1]),.din(n10635));
	jspl jspl_w_n10664_0(.douta(w_n10664_0[0]),.doutb(w_n10664_0[1]),.din(n10664));
	jspl jspl_w_n10671_0(.douta(w_n10671_0[0]),.doutb(w_n10671_0[1]),.din(n10671));
	jspl jspl_w_n10684_0(.douta(w_n10684_0[0]),.doutb(w_n10684_0[1]),.din(n10684));
	jspl jspl_w_n10709_0(.douta(w_n10709_0[0]),.doutb(w_n10709_0[1]),.din(n10709));
	jspl jspl_w_n10716_0(.douta(w_n10716_0[0]),.doutb(w_n10716_0[1]),.din(n10716));
	jspl jspl_w_n10729_0(.douta(w_n10729_0[0]),.doutb(w_n10729_0[1]),.din(n10729));
	jspl jspl_w_n10736_0(.douta(w_n10736_0[0]),.doutb(w_n10736_0[1]),.din(n10736));
	jspl jspl_w_n10743_0(.douta(w_n10743_0[0]),.doutb(w_n10743_0[1]),.din(n10743));
	jspl jspl_w_n10750_0(.douta(w_n10750_0[0]),.doutb(w_n10750_0[1]),.din(n10750));
	jspl jspl_w_n10754_0(.douta(w_n10754_0[0]),.doutb(w_n10754_0[1]),.din(n10754));
	jspl jspl_w_n10758_0(.douta(w_n10758_0[0]),.doutb(w_n10758_0[1]),.din(n10758));
	jspl jspl_w_n10771_0(.douta(w_n10771_0[0]),.doutb(w_n10771_0[1]),.din(n10771));
	jspl jspl_w_n10783_0(.douta(w_n10783_0[0]),.doutb(w_n10783_0[1]),.din(n10783));
	jspl3 jspl3_w_n10785_0(.douta(w_n10785_0[0]),.doutb(w_n10785_0[1]),.doutc(w_n10785_0[2]),.din(n10785));
	jspl3 jspl3_w_n10788_0(.douta(w_n10788_0[0]),.doutb(w_n10788_0[1]),.doutc(w_n10788_0[2]),.din(n10788));
	jspl jspl_w_n10788_1(.douta(w_n10788_1[0]),.doutb(w_n10788_1[1]),.din(w_n10788_0[0]));
	jspl jspl_w_n10789_0(.douta(w_n10789_0[0]),.doutb(w_n10789_0[1]),.din(n10789));
	jspl jspl_w_n10791_0(.douta(w_n10791_0[0]),.doutb(w_n10791_0[1]),.din(n10791));
	jspl jspl_w_n10793_0(.douta(w_n10793_0[0]),.doutb(w_n10793_0[1]),.din(n10793));
	jspl jspl_w_n10794_0(.douta(w_n10794_0[0]),.doutb(w_n10794_0[1]),.din(n10794));
	jspl3 jspl3_w_n10795_0(.douta(w_n10795_0[0]),.doutb(w_n10795_0[1]),.doutc(w_n10795_0[2]),.din(n10795));
	jspl jspl_w_n10801_0(.douta(w_n10801_0[0]),.doutb(w_n10801_0[1]),.din(n10801));
	jspl jspl_w_n10802_0(.douta(w_n10802_0[0]),.doutb(w_n10802_0[1]),.din(n10802));
	jspl3 jspl3_w_n10805_0(.douta(w_n10805_0[0]),.doutb(w_n10805_0[1]),.doutc(w_n10805_0[2]),.din(n10805));
	jspl3 jspl3_w_n10805_1(.douta(w_n10805_1[0]),.doutb(w_n10805_1[1]),.doutc(w_n10805_1[2]),.din(w_n10805_0[0]));
	jspl jspl_w_n10806_0(.douta(w_n10806_0[0]),.doutb(w_n10806_0[1]),.din(n10806));
	jspl3 jspl3_w_n10807_0(.douta(w_n10807_0[0]),.doutb(w_n10807_0[1]),.doutc(w_n10807_0[2]),.din(n10807));
	jspl jspl_w_n10808_0(.douta(w_n10808_0[0]),.doutb(w_n10808_0[1]),.din(n10808));
	jspl jspl_w_n10811_0(.douta(w_n10811_0[0]),.doutb(w_n10811_0[1]),.din(n10811));
	jspl jspl_w_n10813_0(.douta(w_n10813_0[0]),.doutb(w_n10813_0[1]),.din(n10813));
	jspl jspl_w_n10814_0(.douta(w_n10814_0[0]),.doutb(w_n10814_0[1]),.din(n10814));
	jspl jspl_w_n10815_0(.douta(w_n10815_0[0]),.doutb(w_n10815_0[1]),.din(n10815));
	jspl3 jspl3_w_n10820_0(.douta(w_n10820_0[0]),.doutb(w_n10820_0[1]),.doutc(w_n10820_0[2]),.din(n10820));
	jspl3 jspl3_w_n10824_0(.douta(w_n10824_0[0]),.doutb(w_n10824_0[1]),.doutc(w_n10824_0[2]),.din(n10824));
	jspl3 jspl3_w_n10824_1(.douta(w_n10824_1[0]),.doutb(w_n10824_1[1]),.doutc(w_n10824_1[2]),.din(w_n10824_0[0]));
	jspl3 jspl3_w_n10824_2(.douta(w_n10824_2[0]),.doutb(w_n10824_2[1]),.doutc(w_n10824_2[2]),.din(w_n10824_0[1]));
	jspl3 jspl3_w_n10824_3(.douta(w_n10824_3[0]),.doutb(w_n10824_3[1]),.doutc(w_n10824_3[2]),.din(w_n10824_0[2]));
	jspl3 jspl3_w_n10824_4(.douta(w_n10824_4[0]),.doutb(w_n10824_4[1]),.doutc(w_n10824_4[2]),.din(w_n10824_1[0]));
	jspl3 jspl3_w_n10824_5(.douta(w_n10824_5[0]),.doutb(w_n10824_5[1]),.doutc(w_n10824_5[2]),.din(w_n10824_1[1]));
	jspl3 jspl3_w_n10824_6(.douta(w_n10824_6[0]),.doutb(w_n10824_6[1]),.doutc(w_n10824_6[2]),.din(w_n10824_1[2]));
	jspl3 jspl3_w_n10824_7(.douta(w_n10824_7[0]),.doutb(w_n10824_7[1]),.doutc(w_n10824_7[2]),.din(w_n10824_2[0]));
	jspl3 jspl3_w_n10824_8(.douta(w_n10824_8[0]),.doutb(w_n10824_8[1]),.doutc(w_n10824_8[2]),.din(w_n10824_2[1]));
	jspl3 jspl3_w_n10824_9(.douta(w_n10824_9[0]),.doutb(w_n10824_9[1]),.doutc(w_n10824_9[2]),.din(w_n10824_2[2]));
	jspl3 jspl3_w_n10824_10(.douta(w_n10824_10[0]),.doutb(w_n10824_10[1]),.doutc(w_n10824_10[2]),.din(w_n10824_3[0]));
	jspl3 jspl3_w_n10824_11(.douta(w_n10824_11[0]),.doutb(w_n10824_11[1]),.doutc(w_n10824_11[2]),.din(w_n10824_3[1]));
	jspl3 jspl3_w_n10824_12(.douta(w_n10824_12[0]),.doutb(w_n10824_12[1]),.doutc(w_n10824_12[2]),.din(w_n10824_3[2]));
	jspl3 jspl3_w_n10824_13(.douta(w_n10824_13[0]),.doutb(w_n10824_13[1]),.doutc(w_n10824_13[2]),.din(w_n10824_4[0]));
	jspl3 jspl3_w_n10824_14(.douta(w_n10824_14[0]),.doutb(w_n10824_14[1]),.doutc(w_n10824_14[2]),.din(w_n10824_4[1]));
	jspl3 jspl3_w_n10824_15(.douta(w_n10824_15[0]),.doutb(w_n10824_15[1]),.doutc(w_n10824_15[2]),.din(w_n10824_4[2]));
	jspl3 jspl3_w_n10824_16(.douta(w_n10824_16[0]),.doutb(w_n10824_16[1]),.doutc(w_n10824_16[2]),.din(w_n10824_5[0]));
	jspl3 jspl3_w_n10824_17(.douta(w_n10824_17[0]),.doutb(w_n10824_17[1]),.doutc(w_n10824_17[2]),.din(w_n10824_5[1]));
	jspl3 jspl3_w_n10824_18(.douta(w_n10824_18[0]),.doutb(w_n10824_18[1]),.doutc(w_n10824_18[2]),.din(w_n10824_5[2]));
	jspl3 jspl3_w_n10824_19(.douta(w_n10824_19[0]),.doutb(w_n10824_19[1]),.doutc(w_n10824_19[2]),.din(w_n10824_6[0]));
	jspl3 jspl3_w_n10824_20(.douta(w_n10824_20[0]),.doutb(w_n10824_20[1]),.doutc(w_n10824_20[2]),.din(w_n10824_6[1]));
	jspl3 jspl3_w_n10824_21(.douta(w_n10824_21[0]),.doutb(w_n10824_21[1]),.doutc(w_n10824_21[2]),.din(w_n10824_6[2]));
	jspl3 jspl3_w_n10824_22(.douta(w_n10824_22[0]),.doutb(w_n10824_22[1]),.doutc(w_n10824_22[2]),.din(w_n10824_7[0]));
	jspl3 jspl3_w_n10824_23(.douta(w_n10824_23[0]),.doutb(w_n10824_23[1]),.doutc(w_n10824_23[2]),.din(w_n10824_7[1]));
	jspl3 jspl3_w_n10824_24(.douta(w_n10824_24[0]),.doutb(w_n10824_24[1]),.doutc(w_n10824_24[2]),.din(w_n10824_7[2]));
	jspl3 jspl3_w_n10824_25(.douta(w_n10824_25[0]),.doutb(w_n10824_25[1]),.doutc(w_n10824_25[2]),.din(w_n10824_8[0]));
	jspl3 jspl3_w_n10824_26(.douta(w_n10824_26[0]),.doutb(w_n10824_26[1]),.doutc(w_n10824_26[2]),.din(w_n10824_8[1]));
	jspl3 jspl3_w_n10824_27(.douta(w_n10824_27[0]),.doutb(w_n10824_27[1]),.doutc(w_n10824_27[2]),.din(w_n10824_8[2]));
	jspl3 jspl3_w_n10824_28(.douta(w_n10824_28[0]),.doutb(w_n10824_28[1]),.doutc(w_n10824_28[2]),.din(w_n10824_9[0]));
	jspl3 jspl3_w_n10824_29(.douta(w_n10824_29[0]),.doutb(w_n10824_29[1]),.doutc(w_n10824_29[2]),.din(w_n10824_9[1]));
	jspl3 jspl3_w_n10824_30(.douta(w_n10824_30[0]),.doutb(w_n10824_30[1]),.doutc(w_n10824_30[2]),.din(w_n10824_9[2]));
	jspl3 jspl3_w_n10824_31(.douta(w_n10824_31[0]),.doutb(w_n10824_31[1]),.doutc(w_n10824_31[2]),.din(w_n10824_10[0]));
	jspl3 jspl3_w_n10824_32(.douta(w_n10824_32[0]),.doutb(w_n10824_32[1]),.doutc(w_n10824_32[2]),.din(w_n10824_10[1]));
	jspl3 jspl3_w_n10824_33(.douta(w_n10824_33[0]),.doutb(w_n10824_33[1]),.doutc(w_n10824_33[2]),.din(w_n10824_10[2]));
	jspl3 jspl3_w_n10824_34(.douta(w_n10824_34[0]),.doutb(w_n10824_34[1]),.doutc(w_n10824_34[2]),.din(w_n10824_11[0]));
	jspl3 jspl3_w_n10824_35(.douta(w_n10824_35[0]),.doutb(w_n10824_35[1]),.doutc(w_n10824_35[2]),.din(w_n10824_11[1]));
	jspl3 jspl3_w_n10824_36(.douta(w_n10824_36[0]),.doutb(w_n10824_36[1]),.doutc(w_n10824_36[2]),.din(w_n10824_11[2]));
	jspl3 jspl3_w_n10824_37(.douta(w_n10824_37[0]),.doutb(w_n10824_37[1]),.doutc(w_n10824_37[2]),.din(w_n10824_12[0]));
	jspl3 jspl3_w_n10824_38(.douta(w_n10824_38[0]),.doutb(w_n10824_38[1]),.doutc(w_n10824_38[2]),.din(w_n10824_12[1]));
	jspl3 jspl3_w_n10824_39(.douta(w_n10824_39[0]),.doutb(w_n10824_39[1]),.doutc(w_n10824_39[2]),.din(w_n10824_12[2]));
	jspl3 jspl3_w_n10824_40(.douta(w_n10824_40[0]),.doutb(w_n10824_40[1]),.doutc(w_n10824_40[2]),.din(w_n10824_13[0]));
	jspl3 jspl3_w_n10824_41(.douta(w_n10824_41[0]),.doutb(w_n10824_41[1]),.doutc(w_n10824_41[2]),.din(w_n10824_13[1]));
	jspl3 jspl3_w_n10824_42(.douta(w_n10824_42[0]),.doutb(w_n10824_42[1]),.doutc(w_n10824_42[2]),.din(w_n10824_13[2]));
	jspl3 jspl3_w_n10824_43(.douta(w_n10824_43[0]),.doutb(w_n10824_43[1]),.doutc(w_n10824_43[2]),.din(w_n10824_14[0]));
	jspl3 jspl3_w_n10824_44(.douta(w_n10824_44[0]),.doutb(w_n10824_44[1]),.doutc(w_n10824_44[2]),.din(w_n10824_14[1]));
	jspl3 jspl3_w_n10824_45(.douta(w_n10824_45[0]),.doutb(w_n10824_45[1]),.doutc(w_n10824_45[2]),.din(w_n10824_14[2]));
	jspl3 jspl3_w_n10824_46(.douta(w_n10824_46[0]),.doutb(w_n10824_46[1]),.doutc(w_n10824_46[2]),.din(w_n10824_15[0]));
	jspl3 jspl3_w_n10824_47(.douta(w_n10824_47[0]),.doutb(w_n10824_47[1]),.doutc(w_n10824_47[2]),.din(w_n10824_15[1]));
	jspl3 jspl3_w_n10826_0(.douta(w_n10826_0[0]),.doutb(w_n10826_0[1]),.doutc(w_n10826_0[2]),.din(n10826));
	jspl jspl_w_n10827_0(.douta(w_n10827_0[0]),.doutb(w_n10827_0[1]),.din(n10827));
	jspl3 jspl3_w_n10834_0(.douta(w_n10834_0[0]),.doutb(w_n10834_0[1]),.doutc(w_n10834_0[2]),.din(n10834));
	jspl jspl_w_n10835_0(.douta(w_n10835_0[0]),.doutb(w_n10835_0[1]),.din(n10835));
	jspl jspl_w_n10838_0(.douta(w_n10838_0[0]),.doutb(w_n10838_0[1]),.din(n10838));
	jspl3 jspl3_w_n10843_0(.douta(w_n10843_0[0]),.doutb(w_n10843_0[1]),.doutc(w_n10843_0[2]),.din(n10843));
	jspl3 jspl3_w_n10845_0(.douta(w_n10845_0[0]),.doutb(w_n10845_0[1]),.doutc(w_n10845_0[2]),.din(n10845));
	jspl jspl_w_n10846_0(.douta(w_n10846_0[0]),.doutb(w_n10846_0[1]),.din(n10846));
	jspl3 jspl3_w_n10850_0(.douta(w_n10850_0[0]),.doutb(w_n10850_0[1]),.doutc(w_n10850_0[2]),.din(n10850));
	jspl3 jspl3_w_n10852_0(.douta(w_n10852_0[0]),.doutb(w_n10852_0[1]),.doutc(w_n10852_0[2]),.din(n10852));
	jspl jspl_w_n10853_0(.douta(w_n10853_0[0]),.doutb(w_n10853_0[1]),.din(n10853));
	jspl3 jspl3_w_n10857_0(.douta(w_n10857_0[0]),.doutb(w_n10857_0[1]),.doutc(w_n10857_0[2]),.din(n10857));
	jspl3 jspl3_w_n10859_0(.douta(w_n10859_0[0]),.doutb(w_n10859_0[1]),.doutc(w_n10859_0[2]),.din(n10859));
	jspl jspl_w_n10860_0(.douta(w_n10860_0[0]),.doutb(w_n10860_0[1]),.din(n10860));
	jspl3 jspl3_w_n10864_0(.douta(w_n10864_0[0]),.doutb(w_n10864_0[1]),.doutc(w_n10864_0[2]),.din(n10864));
	jspl3 jspl3_w_n10867_0(.douta(w_n10867_0[0]),.doutb(w_n10867_0[1]),.doutc(w_n10867_0[2]),.din(n10867));
	jspl jspl_w_n10868_0(.douta(w_n10868_0[0]),.doutb(w_n10868_0[1]),.din(n10868));
	jspl3 jspl3_w_n10872_0(.douta(w_n10872_0[0]),.doutb(w_n10872_0[1]),.doutc(w_n10872_0[2]),.din(n10872));
	jspl3 jspl3_w_n10874_0(.douta(w_n10874_0[0]),.doutb(w_n10874_0[1]),.doutc(w_n10874_0[2]),.din(n10874));
	jspl jspl_w_n10875_0(.douta(w_n10875_0[0]),.doutb(w_n10875_0[1]),.din(n10875));
	jspl3 jspl3_w_n10879_0(.douta(w_n10879_0[0]),.doutb(w_n10879_0[1]),.doutc(w_n10879_0[2]),.din(n10879));
	jspl3 jspl3_w_n10882_0(.douta(w_n10882_0[0]),.doutb(w_n10882_0[1]),.doutc(w_n10882_0[2]),.din(n10882));
	jspl jspl_w_n10883_0(.douta(w_n10883_0[0]),.doutb(w_n10883_0[1]),.din(n10883));
	jspl3 jspl3_w_n10887_0(.douta(w_n10887_0[0]),.doutb(w_n10887_0[1]),.doutc(w_n10887_0[2]),.din(n10887));
	jspl3 jspl3_w_n10889_0(.douta(w_n10889_0[0]),.doutb(w_n10889_0[1]),.doutc(w_n10889_0[2]),.din(n10889));
	jspl jspl_w_n10890_0(.douta(w_n10890_0[0]),.doutb(w_n10890_0[1]),.din(n10890));
	jspl3 jspl3_w_n10894_0(.douta(w_n10894_0[0]),.doutb(w_n10894_0[1]),.doutc(w_n10894_0[2]),.din(n10894));
	jspl3 jspl3_w_n10896_0(.douta(w_n10896_0[0]),.doutb(w_n10896_0[1]),.doutc(w_n10896_0[2]),.din(n10896));
	jspl jspl_w_n10897_0(.douta(w_n10897_0[0]),.doutb(w_n10897_0[1]),.din(n10897));
	jspl3 jspl3_w_n10901_0(.douta(w_n10901_0[0]),.doutb(w_n10901_0[1]),.doutc(w_n10901_0[2]),.din(n10901));
	jspl3 jspl3_w_n10903_0(.douta(w_n10903_0[0]),.doutb(w_n10903_0[1]),.doutc(w_n10903_0[2]),.din(n10903));
	jspl jspl_w_n10904_0(.douta(w_n10904_0[0]),.doutb(w_n10904_0[1]),.din(n10904));
	jspl3 jspl3_w_n10908_0(.douta(w_n10908_0[0]),.doutb(w_n10908_0[1]),.doutc(w_n10908_0[2]),.din(n10908));
	jspl3 jspl3_w_n10911_0(.douta(w_n10911_0[0]),.doutb(w_n10911_0[1]),.doutc(w_n10911_0[2]),.din(n10911));
	jspl jspl_w_n10912_0(.douta(w_n10912_0[0]),.doutb(w_n10912_0[1]),.din(n10912));
	jspl3 jspl3_w_n10916_0(.douta(w_n10916_0[0]),.doutb(w_n10916_0[1]),.doutc(w_n10916_0[2]),.din(n10916));
	jspl3 jspl3_w_n10918_0(.douta(w_n10918_0[0]),.doutb(w_n10918_0[1]),.doutc(w_n10918_0[2]),.din(n10918));
	jspl jspl_w_n10919_0(.douta(w_n10919_0[0]),.doutb(w_n10919_0[1]),.din(n10919));
	jspl3 jspl3_w_n10923_0(.douta(w_n10923_0[0]),.doutb(w_n10923_0[1]),.doutc(w_n10923_0[2]),.din(n10923));
	jspl3 jspl3_w_n10925_0(.douta(w_n10925_0[0]),.doutb(w_n10925_0[1]),.doutc(w_n10925_0[2]),.din(n10925));
	jspl jspl_w_n10926_0(.douta(w_n10926_0[0]),.doutb(w_n10926_0[1]),.din(n10926));
	jspl3 jspl3_w_n10930_0(.douta(w_n10930_0[0]),.doutb(w_n10930_0[1]),.doutc(w_n10930_0[2]),.din(n10930));
	jspl3 jspl3_w_n10932_0(.douta(w_n10932_0[0]),.doutb(w_n10932_0[1]),.doutc(w_n10932_0[2]),.din(n10932));
	jspl jspl_w_n10933_0(.douta(w_n10933_0[0]),.doutb(w_n10933_0[1]),.din(n10933));
	jspl3 jspl3_w_n10937_0(.douta(w_n10937_0[0]),.doutb(w_n10937_0[1]),.doutc(w_n10937_0[2]),.din(n10937));
	jspl3 jspl3_w_n10939_0(.douta(w_n10939_0[0]),.doutb(w_n10939_0[1]),.doutc(w_n10939_0[2]),.din(n10939));
	jspl jspl_w_n10940_0(.douta(w_n10940_0[0]),.doutb(w_n10940_0[1]),.din(n10940));
	jspl3 jspl3_w_n10944_0(.douta(w_n10944_0[0]),.doutb(w_n10944_0[1]),.doutc(w_n10944_0[2]),.din(n10944));
	jspl3 jspl3_w_n10946_0(.douta(w_n10946_0[0]),.doutb(w_n10946_0[1]),.doutc(w_n10946_0[2]),.din(n10946));
	jspl jspl_w_n10947_0(.douta(w_n10947_0[0]),.doutb(w_n10947_0[1]),.din(n10947));
	jspl3 jspl3_w_n10950_0(.douta(w_n10950_0[0]),.doutb(w_n10950_0[1]),.doutc(w_n10950_0[2]),.din(n10950));
	jspl3 jspl3_w_n10954_0(.douta(w_n10954_0[0]),.doutb(w_n10954_0[1]),.doutc(w_n10954_0[2]),.din(n10954));
	jspl jspl_w_n10955_0(.douta(w_n10955_0[0]),.doutb(w_n10955_0[1]),.din(n10955));
	jspl3 jspl3_w_n10959_0(.douta(w_n10959_0[0]),.doutb(w_n10959_0[1]),.doutc(w_n10959_0[2]),.din(n10959));
	jspl3 jspl3_w_n10961_0(.douta(w_n10961_0[0]),.doutb(w_n10961_0[1]),.doutc(w_n10961_0[2]),.din(n10961));
	jspl jspl_w_n10962_0(.douta(w_n10962_0[0]),.doutb(w_n10962_0[1]),.din(n10962));
	jspl3 jspl3_w_n10966_0(.douta(w_n10966_0[0]),.doutb(w_n10966_0[1]),.doutc(w_n10966_0[2]),.din(n10966));
	jspl3 jspl3_w_n10969_0(.douta(w_n10969_0[0]),.doutb(w_n10969_0[1]),.doutc(w_n10969_0[2]),.din(n10969));
	jspl jspl_w_n10970_0(.douta(w_n10970_0[0]),.doutb(w_n10970_0[1]),.din(n10970));
	jspl3 jspl3_w_n10974_0(.douta(w_n10974_0[0]),.doutb(w_n10974_0[1]),.doutc(w_n10974_0[2]),.din(n10974));
	jspl3 jspl3_w_n10976_0(.douta(w_n10976_0[0]),.doutb(w_n10976_0[1]),.doutc(w_n10976_0[2]),.din(n10976));
	jspl jspl_w_n10977_0(.douta(w_n10977_0[0]),.doutb(w_n10977_0[1]),.din(n10977));
	jspl3 jspl3_w_n10981_0(.douta(w_n10981_0[0]),.doutb(w_n10981_0[1]),.doutc(w_n10981_0[2]),.din(n10981));
	jspl3 jspl3_w_n10984_0(.douta(w_n10984_0[0]),.doutb(w_n10984_0[1]),.doutc(w_n10984_0[2]),.din(n10984));
	jspl jspl_w_n10985_0(.douta(w_n10985_0[0]),.doutb(w_n10985_0[1]),.din(n10985));
	jspl3 jspl3_w_n10989_0(.douta(w_n10989_0[0]),.doutb(w_n10989_0[1]),.doutc(w_n10989_0[2]),.din(n10989));
	jspl3 jspl3_w_n10991_0(.douta(w_n10991_0[0]),.doutb(w_n10991_0[1]),.doutc(w_n10991_0[2]),.din(n10991));
	jspl jspl_w_n10992_0(.douta(w_n10992_0[0]),.doutb(w_n10992_0[1]),.din(n10992));
	jspl3 jspl3_w_n10996_0(.douta(w_n10996_0[0]),.doutb(w_n10996_0[1]),.doutc(w_n10996_0[2]),.din(n10996));
	jspl3 jspl3_w_n10998_0(.douta(w_n10998_0[0]),.doutb(w_n10998_0[1]),.doutc(w_n10998_0[2]),.din(n10998));
	jspl jspl_w_n10999_0(.douta(w_n10999_0[0]),.doutb(w_n10999_0[1]),.din(n10999));
	jspl3 jspl3_w_n11003_0(.douta(w_n11003_0[0]),.doutb(w_n11003_0[1]),.doutc(w_n11003_0[2]),.din(n11003));
	jspl3 jspl3_w_n11005_0(.douta(w_n11005_0[0]),.doutb(w_n11005_0[1]),.doutc(w_n11005_0[2]),.din(n11005));
	jspl jspl_w_n11006_0(.douta(w_n11006_0[0]),.doutb(w_n11006_0[1]),.din(n11006));
	jspl3 jspl3_w_n11010_0(.douta(w_n11010_0[0]),.doutb(w_n11010_0[1]),.doutc(w_n11010_0[2]),.din(n11010));
	jspl3 jspl3_w_n11013_0(.douta(w_n11013_0[0]),.doutb(w_n11013_0[1]),.doutc(w_n11013_0[2]),.din(n11013));
	jspl jspl_w_n11014_0(.douta(w_n11014_0[0]),.doutb(w_n11014_0[1]),.din(n11014));
	jspl3 jspl3_w_n11018_0(.douta(w_n11018_0[0]),.doutb(w_n11018_0[1]),.doutc(w_n11018_0[2]),.din(n11018));
	jspl3 jspl3_w_n11020_0(.douta(w_n11020_0[0]),.doutb(w_n11020_0[1]),.doutc(w_n11020_0[2]),.din(n11020));
	jspl jspl_w_n11021_0(.douta(w_n11021_0[0]),.doutb(w_n11021_0[1]),.din(n11021));
	jspl3 jspl3_w_n11025_0(.douta(w_n11025_0[0]),.doutb(w_n11025_0[1]),.doutc(w_n11025_0[2]),.din(n11025));
	jspl3 jspl3_w_n11028_0(.douta(w_n11028_0[0]),.doutb(w_n11028_0[1]),.doutc(w_n11028_0[2]),.din(n11028));
	jspl jspl_w_n11029_0(.douta(w_n11029_0[0]),.doutb(w_n11029_0[1]),.din(n11029));
	jspl3 jspl3_w_n11033_0(.douta(w_n11033_0[0]),.doutb(w_n11033_0[1]),.doutc(w_n11033_0[2]),.din(n11033));
	jspl3 jspl3_w_n11035_0(.douta(w_n11035_0[0]),.doutb(w_n11035_0[1]),.doutc(w_n11035_0[2]),.din(n11035));
	jspl jspl_w_n11036_0(.douta(w_n11036_0[0]),.doutb(w_n11036_0[1]),.din(n11036));
	jspl3 jspl3_w_n11040_0(.douta(w_n11040_0[0]),.doutb(w_n11040_0[1]),.doutc(w_n11040_0[2]),.din(n11040));
	jspl3 jspl3_w_n11043_0(.douta(w_n11043_0[0]),.doutb(w_n11043_0[1]),.doutc(w_n11043_0[2]),.din(n11043));
	jspl jspl_w_n11044_0(.douta(w_n11044_0[0]),.doutb(w_n11044_0[1]),.din(n11044));
	jspl3 jspl3_w_n11048_0(.douta(w_n11048_0[0]),.doutb(w_n11048_0[1]),.doutc(w_n11048_0[2]),.din(n11048));
	jspl3 jspl3_w_n11050_0(.douta(w_n11050_0[0]),.doutb(w_n11050_0[1]),.doutc(w_n11050_0[2]),.din(n11050));
	jspl jspl_w_n11051_0(.douta(w_n11051_0[0]),.doutb(w_n11051_0[1]),.din(n11051));
	jspl3 jspl3_w_n11055_0(.douta(w_n11055_0[0]),.doutb(w_n11055_0[1]),.doutc(w_n11055_0[2]),.din(n11055));
	jspl3 jspl3_w_n11058_0(.douta(w_n11058_0[0]),.doutb(w_n11058_0[1]),.doutc(w_n11058_0[2]),.din(n11058));
	jspl jspl_w_n11059_0(.douta(w_n11059_0[0]),.doutb(w_n11059_0[1]),.din(n11059));
	jspl3 jspl3_w_n11063_0(.douta(w_n11063_0[0]),.doutb(w_n11063_0[1]),.doutc(w_n11063_0[2]),.din(n11063));
	jspl3 jspl3_w_n11066_0(.douta(w_n11066_0[0]),.doutb(w_n11066_0[1]),.doutc(w_n11066_0[2]),.din(n11066));
	jspl jspl_w_n11067_0(.douta(w_n11067_0[0]),.doutb(w_n11067_0[1]),.din(n11067));
	jspl3 jspl3_w_n11071_0(.douta(w_n11071_0[0]),.doutb(w_n11071_0[1]),.doutc(w_n11071_0[2]),.din(n11071));
	jspl3 jspl3_w_n11074_0(.douta(w_n11074_0[0]),.doutb(w_n11074_0[1]),.doutc(w_n11074_0[2]),.din(n11074));
	jspl jspl_w_n11075_0(.douta(w_n11075_0[0]),.doutb(w_n11075_0[1]),.din(n11075));
	jspl3 jspl3_w_n11079_0(.douta(w_n11079_0[0]),.doutb(w_n11079_0[1]),.doutc(w_n11079_0[2]),.din(n11079));
	jspl3 jspl3_w_n11081_0(.douta(w_n11081_0[0]),.doutb(w_n11081_0[1]),.doutc(w_n11081_0[2]),.din(n11081));
	jspl jspl_w_n11082_0(.douta(w_n11082_0[0]),.doutb(w_n11082_0[1]),.din(n11082));
	jspl3 jspl3_w_n11086_0(.douta(w_n11086_0[0]),.doutb(w_n11086_0[1]),.doutc(w_n11086_0[2]),.din(n11086));
	jspl3 jspl3_w_n11088_0(.douta(w_n11088_0[0]),.doutb(w_n11088_0[1]),.doutc(w_n11088_0[2]),.din(n11088));
	jspl jspl_w_n11089_0(.douta(w_n11089_0[0]),.doutb(w_n11089_0[1]),.din(n11089));
	jspl3 jspl3_w_n11093_0(.douta(w_n11093_0[0]),.doutb(w_n11093_0[1]),.doutc(w_n11093_0[2]),.din(n11093));
	jspl3 jspl3_w_n11095_0(.douta(w_n11095_0[0]),.doutb(w_n11095_0[1]),.doutc(w_n11095_0[2]),.din(n11095));
	jspl jspl_w_n11096_0(.douta(w_n11096_0[0]),.doutb(w_n11096_0[1]),.din(n11096));
	jspl3 jspl3_w_n11100_0(.douta(w_n11100_0[0]),.doutb(w_n11100_0[1]),.doutc(w_n11100_0[2]),.din(n11100));
	jspl3 jspl3_w_n11103_0(.douta(w_n11103_0[0]),.doutb(w_n11103_0[1]),.doutc(w_n11103_0[2]),.din(n11103));
	jspl jspl_w_n11104_0(.douta(w_n11104_0[0]),.doutb(w_n11104_0[1]),.din(n11104));
	jspl3 jspl3_w_n11108_0(.douta(w_n11108_0[0]),.doutb(w_n11108_0[1]),.doutc(w_n11108_0[2]),.din(n11108));
	jspl3 jspl3_w_n11110_0(.douta(w_n11110_0[0]),.doutb(w_n11110_0[1]),.doutc(w_n11110_0[2]),.din(n11110));
	jspl jspl_w_n11111_0(.douta(w_n11111_0[0]),.doutb(w_n11111_0[1]),.din(n11111));
	jspl jspl_w_n11115_0(.douta(w_n11115_0[0]),.doutb(w_n11115_0[1]),.din(n11115));
	jspl3 jspl3_w_n11117_0(.douta(w_n11117_0[0]),.doutb(w_n11117_0[1]),.doutc(w_n11117_0[2]),.din(n11117));
	jspl jspl_w_n11117_1(.douta(w_n11117_1[0]),.doutb(w_n11117_1[1]),.din(w_n11117_0[0]));
	jspl3 jspl3_w_n11120_0(.douta(w_n11120_0[0]),.doutb(w_n11120_0[1]),.doutc(w_n11120_0[2]),.din(n11120));
	jspl jspl_w_n11120_1(.douta(w_n11120_1[0]),.doutb(w_n11120_1[1]),.din(w_n11120_0[0]));
	jspl jspl_w_n11121_0(.douta(w_n11121_0[0]),.doutb(w_n11121_0[1]),.din(n11121));
	jspl jspl_w_n11125_0(.douta(w_n11125_0[0]),.doutb(w_n11125_0[1]),.din(n11125));
	jspl jspl_w_n11126_0(.douta(w_n11126_0[0]),.doutb(w_n11126_0[1]),.din(n11126));
	jspl jspl_w_n11128_0(.douta(w_n11128_0[0]),.doutb(w_n11128_0[1]),.din(n11128));
	jspl jspl_w_n11133_0(.douta(w_n11133_0[0]),.doutb(w_n11133_0[1]),.din(n11133));
	jspl jspl_w_n11137_0(.douta(w_n11137_0[0]),.doutb(w_n11137_0[1]),.din(n11137));
	jspl3 jspl3_w_n11140_0(.douta(w_n11140_0[0]),.doutb(w_n11140_0[1]),.doutc(w_n11140_0[2]),.din(n11140));
	jspl3 jspl3_w_n11142_0(.douta(w_n11142_0[0]),.doutb(w_n11142_0[1]),.doutc(w_n11142_0[2]),.din(n11142));
	jspl jspl_w_n11142_1(.douta(w_n11142_1[0]),.doutb(w_n11142_1[1]),.din(w_n11142_0[0]));
	jspl jspl_w_n11143_0(.douta(w_n11143_0[0]),.doutb(w_n11143_0[1]),.din(n11143));
	jspl3 jspl3_w_n11144_0(.douta(w_n11144_0[0]),.doutb(w_n11144_0[1]),.doutc(w_n11144_0[2]),.din(n11144));
	jspl jspl_w_n11145_0(.douta(w_n11145_0[0]),.doutb(w_n11145_0[1]),.din(n11145));
	jspl3 jspl3_w_n11146_0(.douta(w_n11146_0[0]),.doutb(w_n11146_0[1]),.doutc(w_n11146_0[2]),.din(n11146));
	jspl jspl_w_n11147_0(.douta(w_n11147_0[0]),.doutb(w_n11147_0[1]),.din(n11147));
	jspl jspl_w_n11152_0(.douta(w_n11152_0[0]),.doutb(w_n11152_0[1]),.din(n11152));
	jspl jspl_w_n11198_0(.douta(w_n11198_0[0]),.doutb(w_n11198_0[1]),.din(n11198));
	jspl jspl_w_n11343_0(.douta(w_n11343_0[0]),.doutb(w_n11343_0[1]),.din(n11343));
	jspl jspl_w_n11346_0(.douta(w_n11346_0[0]),.doutb(w_n11346_0[1]),.din(n11346));
	jspl3 jspl3_w_n11347_0(.douta(w_n11347_0[0]),.doutb(w_n11347_0[1]),.doutc(w_n11347_0[2]),.din(n11347));
	jspl3 jspl3_w_n11347_1(.douta(w_n11347_1[0]),.doutb(w_n11347_1[1]),.doutc(w_n11347_1[2]),.din(w_n11347_0[0]));
	jspl3 jspl3_w_n11347_2(.douta(w_n11347_2[0]),.doutb(w_n11347_2[1]),.doutc(w_n11347_2[2]),.din(w_n11347_0[1]));
	jspl3 jspl3_w_n11347_3(.douta(w_n11347_3[0]),.doutb(w_n11347_3[1]),.doutc(w_n11347_3[2]),.din(w_n11347_0[2]));
	jspl3 jspl3_w_n11347_4(.douta(w_n11347_4[0]),.doutb(w_n11347_4[1]),.doutc(w_n11347_4[2]),.din(w_n11347_1[0]));
	jspl3 jspl3_w_n11347_5(.douta(w_n11347_5[0]),.doutb(w_n11347_5[1]),.doutc(w_n11347_5[2]),.din(w_n11347_1[1]));
	jspl3 jspl3_w_n11347_6(.douta(w_n11347_6[0]),.doutb(w_n11347_6[1]),.doutc(w_n11347_6[2]),.din(w_n11347_1[2]));
	jspl3 jspl3_w_n11347_7(.douta(w_n11347_7[0]),.doutb(w_n11347_7[1]),.doutc(w_n11347_7[2]),.din(w_n11347_2[0]));
	jspl3 jspl3_w_n11347_8(.douta(w_n11347_8[0]),.doutb(w_n11347_8[1]),.doutc(w_n11347_8[2]),.din(w_n11347_2[1]));
	jspl3 jspl3_w_n11347_9(.douta(w_n11347_9[0]),.doutb(w_n11347_9[1]),.doutc(w_n11347_9[2]),.din(w_n11347_2[2]));
	jspl3 jspl3_w_n11347_10(.douta(w_n11347_10[0]),.doutb(w_n11347_10[1]),.doutc(w_n11347_10[2]),.din(w_n11347_3[0]));
	jspl3 jspl3_w_n11347_11(.douta(w_n11347_11[0]),.doutb(w_n11347_11[1]),.doutc(w_n11347_11[2]),.din(w_n11347_3[1]));
	jspl3 jspl3_w_n11347_12(.douta(w_n11347_12[0]),.doutb(w_n11347_12[1]),.doutc(w_n11347_12[2]),.din(w_n11347_3[2]));
	jspl3 jspl3_w_n11347_13(.douta(w_n11347_13[0]),.doutb(w_n11347_13[1]),.doutc(w_n11347_13[2]),.din(w_n11347_4[0]));
	jspl3 jspl3_w_n11347_14(.douta(w_n11347_14[0]),.doutb(w_n11347_14[1]),.doutc(w_n11347_14[2]),.din(w_n11347_4[1]));
	jspl3 jspl3_w_n11347_15(.douta(w_n11347_15[0]),.doutb(w_n11347_15[1]),.doutc(w_n11347_15[2]),.din(w_n11347_4[2]));
	jspl3 jspl3_w_n11347_16(.douta(w_n11347_16[0]),.doutb(w_n11347_16[1]),.doutc(w_n11347_16[2]),.din(w_n11347_5[0]));
	jspl3 jspl3_w_n11347_17(.douta(w_n11347_17[0]),.doutb(w_n11347_17[1]),.doutc(w_n11347_17[2]),.din(w_n11347_5[1]));
	jspl3 jspl3_w_n11347_18(.douta(w_n11347_18[0]),.doutb(w_n11347_18[1]),.doutc(w_n11347_18[2]),.din(w_n11347_5[2]));
	jspl3 jspl3_w_n11347_19(.douta(w_n11347_19[0]),.doutb(w_n11347_19[1]),.doutc(w_n11347_19[2]),.din(w_n11347_6[0]));
	jspl3 jspl3_w_n11347_20(.douta(w_n11347_20[0]),.doutb(w_n11347_20[1]),.doutc(w_n11347_20[2]),.din(w_n11347_6[1]));
	jspl3 jspl3_w_n11347_21(.douta(w_n11347_21[0]),.doutb(w_n11347_21[1]),.doutc(w_n11347_21[2]),.din(w_n11347_6[2]));
	jspl3 jspl3_w_n11347_22(.douta(w_n11347_22[0]),.doutb(w_n11347_22[1]),.doutc(w_n11347_22[2]),.din(w_n11347_7[0]));
	jspl3 jspl3_w_n11347_23(.douta(w_n11347_23[0]),.doutb(w_n11347_23[1]),.doutc(w_n11347_23[2]),.din(w_n11347_7[1]));
	jspl3 jspl3_w_n11347_24(.douta(w_n11347_24[0]),.doutb(w_n11347_24[1]),.doutc(w_n11347_24[2]),.din(w_n11347_7[2]));
	jspl3 jspl3_w_n11347_25(.douta(w_n11347_25[0]),.doutb(w_n11347_25[1]),.doutc(w_n11347_25[2]),.din(w_n11347_8[0]));
	jspl3 jspl3_w_n11347_26(.douta(w_n11347_26[0]),.doutb(w_n11347_26[1]),.doutc(w_n11347_26[2]),.din(w_n11347_8[1]));
	jspl jspl_w_n11347_27(.douta(w_n11347_27[0]),.doutb(w_n11347_27[1]),.din(w_n11347_8[2]));
	jspl3 jspl3_w_n11351_0(.douta(w_n11351_0[0]),.doutb(w_n11351_0[1]),.doutc(w_n11351_0[2]),.din(n11351));
	jspl jspl_w_n11352_0(.douta(w_n11352_0[0]),.doutb(w_n11352_0[1]),.din(n11352));
	jspl jspl_w_n11354_0(.douta(w_n11354_0[0]),.doutb(w_n11354_0[1]),.din(n11354));
	jspl jspl_w_n11359_0(.douta(w_n11359_0[0]),.doutb(w_n11359_0[1]),.din(n11359));
	jspl jspl_w_n11360_0(.douta(w_n11360_0[0]),.doutb(w_n11360_0[1]),.din(n11360));
	jspl3 jspl3_w_n11362_0(.douta(w_n11362_0[0]),.doutb(w_n11362_0[1]),.doutc(w_n11362_0[2]),.din(n11362));
	jspl jspl_w_n11363_0(.douta(w_n11363_0[0]),.doutb(w_n11363_0[1]),.din(n11363));
	jspl jspl_w_n11367_0(.douta(w_n11367_0[0]),.doutb(w_n11367_0[1]),.din(n11367));
	jspl3 jspl3_w_n11369_0(.douta(w_n11369_0[0]),.doutb(w_n11369_0[1]),.doutc(w_n11369_0[2]),.din(n11369));
	jspl jspl_w_n11370_0(.douta(w_n11370_0[0]),.doutb(w_n11370_0[1]),.din(n11370));
	jspl jspl_w_n11374_0(.douta(w_n11374_0[0]),.doutb(w_n11374_0[1]),.din(n11374));
	jspl jspl_w_n11375_0(.douta(w_n11375_0[0]),.doutb(w_n11375_0[1]),.din(n11375));
	jspl3 jspl3_w_n11377_0(.douta(w_n11377_0[0]),.doutb(w_n11377_0[1]),.doutc(w_n11377_0[2]),.din(n11377));
	jspl jspl_w_n11378_0(.douta(w_n11378_0[0]),.doutb(w_n11378_0[1]),.din(n11378));
	jspl jspl_w_n11382_0(.douta(w_n11382_0[0]),.doutb(w_n11382_0[1]),.din(n11382));
	jspl jspl_w_n11383_0(.douta(w_n11383_0[0]),.doutb(w_n11383_0[1]),.din(n11383));
	jspl3 jspl3_w_n11385_0(.douta(w_n11385_0[0]),.doutb(w_n11385_0[1]),.doutc(w_n11385_0[2]),.din(n11385));
	jspl jspl_w_n11386_0(.douta(w_n11386_0[0]),.doutb(w_n11386_0[1]),.din(n11386));
	jspl jspl_w_n11390_0(.douta(w_n11390_0[0]),.doutb(w_n11390_0[1]),.din(n11390));
	jspl jspl_w_n11391_0(.douta(w_n11391_0[0]),.doutb(w_n11391_0[1]),.din(n11391));
	jspl3 jspl3_w_n11393_0(.douta(w_n11393_0[0]),.doutb(w_n11393_0[1]),.doutc(w_n11393_0[2]),.din(n11393));
	jspl jspl_w_n11394_0(.douta(w_n11394_0[0]),.doutb(w_n11394_0[1]),.din(n11394));
	jspl jspl_w_n11398_0(.douta(w_n11398_0[0]),.doutb(w_n11398_0[1]),.din(n11398));
	jspl3 jspl3_w_n11400_0(.douta(w_n11400_0[0]),.doutb(w_n11400_0[1]),.doutc(w_n11400_0[2]),.din(n11400));
	jspl jspl_w_n11401_0(.douta(w_n11401_0[0]),.doutb(w_n11401_0[1]),.din(n11401));
	jspl jspl_w_n11405_0(.douta(w_n11405_0[0]),.doutb(w_n11405_0[1]),.din(n11405));
	jspl jspl_w_n11406_0(.douta(w_n11406_0[0]),.doutb(w_n11406_0[1]),.din(n11406));
	jspl3 jspl3_w_n11408_0(.douta(w_n11408_0[0]),.doutb(w_n11408_0[1]),.doutc(w_n11408_0[2]),.din(n11408));
	jspl jspl_w_n11409_0(.douta(w_n11409_0[0]),.doutb(w_n11409_0[1]),.din(n11409));
	jspl jspl_w_n11413_0(.douta(w_n11413_0[0]),.doutb(w_n11413_0[1]),.din(n11413));
	jspl3 jspl3_w_n11415_0(.douta(w_n11415_0[0]),.doutb(w_n11415_0[1]),.doutc(w_n11415_0[2]),.din(n11415));
	jspl jspl_w_n11416_0(.douta(w_n11416_0[0]),.doutb(w_n11416_0[1]),.din(n11416));
	jspl jspl_w_n11420_0(.douta(w_n11420_0[0]),.doutb(w_n11420_0[1]),.din(n11420));
	jspl jspl_w_n11421_0(.douta(w_n11421_0[0]),.doutb(w_n11421_0[1]),.din(n11421));
	jspl3 jspl3_w_n11423_0(.douta(w_n11423_0[0]),.doutb(w_n11423_0[1]),.doutc(w_n11423_0[2]),.din(n11423));
	jspl jspl_w_n11424_0(.douta(w_n11424_0[0]),.doutb(w_n11424_0[1]),.din(n11424));
	jspl jspl_w_n11428_0(.douta(w_n11428_0[0]),.doutb(w_n11428_0[1]),.din(n11428));
	jspl jspl_w_n11429_0(.douta(w_n11429_0[0]),.doutb(w_n11429_0[1]),.din(n11429));
	jspl3 jspl3_w_n11431_0(.douta(w_n11431_0[0]),.doutb(w_n11431_0[1]),.doutc(w_n11431_0[2]),.din(n11431));
	jspl jspl_w_n11432_0(.douta(w_n11432_0[0]),.doutb(w_n11432_0[1]),.din(n11432));
	jspl jspl_w_n11436_0(.douta(w_n11436_0[0]),.doutb(w_n11436_0[1]),.din(n11436));
	jspl jspl_w_n11437_0(.douta(w_n11437_0[0]),.doutb(w_n11437_0[1]),.din(n11437));
	jspl3 jspl3_w_n11439_0(.douta(w_n11439_0[0]),.doutb(w_n11439_0[1]),.doutc(w_n11439_0[2]),.din(n11439));
	jspl jspl_w_n11440_0(.douta(w_n11440_0[0]),.doutb(w_n11440_0[1]),.din(n11440));
	jspl jspl_w_n11444_0(.douta(w_n11444_0[0]),.doutb(w_n11444_0[1]),.din(n11444));
	jspl3 jspl3_w_n11446_0(.douta(w_n11446_0[0]),.doutb(w_n11446_0[1]),.doutc(w_n11446_0[2]),.din(n11446));
	jspl jspl_w_n11447_0(.douta(w_n11447_0[0]),.doutb(w_n11447_0[1]),.din(n11447));
	jspl jspl_w_n11451_0(.douta(w_n11451_0[0]),.doutb(w_n11451_0[1]),.din(n11451));
	jspl jspl_w_n11452_0(.douta(w_n11452_0[0]),.doutb(w_n11452_0[1]),.din(n11452));
	jspl3 jspl3_w_n11454_0(.douta(w_n11454_0[0]),.doutb(w_n11454_0[1]),.doutc(w_n11454_0[2]),.din(n11454));
	jspl jspl_w_n11455_0(.douta(w_n11455_0[0]),.doutb(w_n11455_0[1]),.din(n11455));
	jspl jspl_w_n11459_0(.douta(w_n11459_0[0]),.doutb(w_n11459_0[1]),.din(n11459));
	jspl jspl_w_n11460_0(.douta(w_n11460_0[0]),.doutb(w_n11460_0[1]),.din(n11460));
	jspl3 jspl3_w_n11462_0(.douta(w_n11462_0[0]),.doutb(w_n11462_0[1]),.doutc(w_n11462_0[2]),.din(n11462));
	jspl jspl_w_n11463_0(.douta(w_n11463_0[0]),.doutb(w_n11463_0[1]),.din(n11463));
	jspl jspl_w_n11467_0(.douta(w_n11467_0[0]),.doutb(w_n11467_0[1]),.din(n11467));
	jspl jspl_w_n11468_0(.douta(w_n11468_0[0]),.doutb(w_n11468_0[1]),.din(n11468));
	jspl3 jspl3_w_n11470_0(.douta(w_n11470_0[0]),.doutb(w_n11470_0[1]),.doutc(w_n11470_0[2]),.din(n11470));
	jspl jspl_w_n11471_0(.douta(w_n11471_0[0]),.doutb(w_n11471_0[1]),.din(n11471));
	jspl jspl_w_n11475_0(.douta(w_n11475_0[0]),.doutb(w_n11475_0[1]),.din(n11475));
	jspl jspl_w_n11476_0(.douta(w_n11476_0[0]),.doutb(w_n11476_0[1]),.din(n11476));
	jspl3 jspl3_w_n11478_0(.douta(w_n11478_0[0]),.doutb(w_n11478_0[1]),.doutc(w_n11478_0[2]),.din(n11478));
	jspl jspl_w_n11479_0(.douta(w_n11479_0[0]),.doutb(w_n11479_0[1]),.din(n11479));
	jspl jspl_w_n11483_0(.douta(w_n11483_0[0]),.doutb(w_n11483_0[1]),.din(n11483));
	jspl jspl_w_n11484_0(.douta(w_n11484_0[0]),.doutb(w_n11484_0[1]),.din(n11484));
	jspl3 jspl3_w_n11486_0(.douta(w_n11486_0[0]),.doutb(w_n11486_0[1]),.doutc(w_n11486_0[2]),.din(n11486));
	jspl jspl_w_n11487_0(.douta(w_n11487_0[0]),.doutb(w_n11487_0[1]),.din(n11487));
	jspl jspl_w_n11490_0(.douta(w_n11490_0[0]),.doutb(w_n11490_0[1]),.din(n11490));
	jspl3 jspl3_w_n11493_0(.douta(w_n11493_0[0]),.doutb(w_n11493_0[1]),.doutc(w_n11493_0[2]),.din(n11493));
	jspl jspl_w_n11494_0(.douta(w_n11494_0[0]),.doutb(w_n11494_0[1]),.din(n11494));
	jspl jspl_w_n11498_0(.douta(w_n11498_0[0]),.doutb(w_n11498_0[1]),.din(n11498));
	jspl jspl_w_n11499_0(.douta(w_n11499_0[0]),.doutb(w_n11499_0[1]),.din(n11499));
	jspl3 jspl3_w_n11501_0(.douta(w_n11501_0[0]),.doutb(w_n11501_0[1]),.doutc(w_n11501_0[2]),.din(n11501));
	jspl jspl_w_n11502_0(.douta(w_n11502_0[0]),.doutb(w_n11502_0[1]),.din(n11502));
	jspl jspl_w_n11506_0(.douta(w_n11506_0[0]),.doutb(w_n11506_0[1]),.din(n11506));
	jspl3 jspl3_w_n11508_0(.douta(w_n11508_0[0]),.doutb(w_n11508_0[1]),.doutc(w_n11508_0[2]),.din(n11508));
	jspl jspl_w_n11509_0(.douta(w_n11509_0[0]),.doutb(w_n11509_0[1]),.din(n11509));
	jspl jspl_w_n11513_0(.douta(w_n11513_0[0]),.doutb(w_n11513_0[1]),.din(n11513));
	jspl jspl_w_n11514_0(.douta(w_n11514_0[0]),.doutb(w_n11514_0[1]),.din(n11514));
	jspl3 jspl3_w_n11516_0(.douta(w_n11516_0[0]),.doutb(w_n11516_0[1]),.doutc(w_n11516_0[2]),.din(n11516));
	jspl jspl_w_n11517_0(.douta(w_n11517_0[0]),.doutb(w_n11517_0[1]),.din(n11517));
	jspl jspl_w_n11521_0(.douta(w_n11521_0[0]),.doutb(w_n11521_0[1]),.din(n11521));
	jspl3 jspl3_w_n11523_0(.douta(w_n11523_0[0]),.doutb(w_n11523_0[1]),.doutc(w_n11523_0[2]),.din(n11523));
	jspl jspl_w_n11524_0(.douta(w_n11524_0[0]),.doutb(w_n11524_0[1]),.din(n11524));
	jspl jspl_w_n11528_0(.douta(w_n11528_0[0]),.doutb(w_n11528_0[1]),.din(n11528));
	jspl jspl_w_n11529_0(.douta(w_n11529_0[0]),.doutb(w_n11529_0[1]),.din(n11529));
	jspl3 jspl3_w_n11531_0(.douta(w_n11531_0[0]),.doutb(w_n11531_0[1]),.doutc(w_n11531_0[2]),.din(n11531));
	jspl jspl_w_n11532_0(.douta(w_n11532_0[0]),.doutb(w_n11532_0[1]),.din(n11532));
	jspl jspl_w_n11536_0(.douta(w_n11536_0[0]),.doutb(w_n11536_0[1]),.din(n11536));
	jspl jspl_w_n11537_0(.douta(w_n11537_0[0]),.doutb(w_n11537_0[1]),.din(n11537));
	jspl3 jspl3_w_n11539_0(.douta(w_n11539_0[0]),.doutb(w_n11539_0[1]),.doutc(w_n11539_0[2]),.din(n11539));
	jspl jspl_w_n11540_0(.douta(w_n11540_0[0]),.doutb(w_n11540_0[1]),.din(n11540));
	jspl jspl_w_n11544_0(.douta(w_n11544_0[0]),.doutb(w_n11544_0[1]),.din(n11544));
	jspl jspl_w_n11545_0(.douta(w_n11545_0[0]),.doutb(w_n11545_0[1]),.din(n11545));
	jspl3 jspl3_w_n11547_0(.douta(w_n11547_0[0]),.doutb(w_n11547_0[1]),.doutc(w_n11547_0[2]),.din(n11547));
	jspl jspl_w_n11548_0(.douta(w_n11548_0[0]),.doutb(w_n11548_0[1]),.din(n11548));
	jspl jspl_w_n11552_0(.douta(w_n11552_0[0]),.doutb(w_n11552_0[1]),.din(n11552));
	jspl3 jspl3_w_n11554_0(.douta(w_n11554_0[0]),.doutb(w_n11554_0[1]),.doutc(w_n11554_0[2]),.din(n11554));
	jspl jspl_w_n11555_0(.douta(w_n11555_0[0]),.doutb(w_n11555_0[1]),.din(n11555));
	jspl jspl_w_n11559_0(.douta(w_n11559_0[0]),.doutb(w_n11559_0[1]),.din(n11559));
	jspl jspl_w_n11560_0(.douta(w_n11560_0[0]),.doutb(w_n11560_0[1]),.din(n11560));
	jspl3 jspl3_w_n11562_0(.douta(w_n11562_0[0]),.doutb(w_n11562_0[1]),.doutc(w_n11562_0[2]),.din(n11562));
	jspl jspl_w_n11563_0(.douta(w_n11563_0[0]),.doutb(w_n11563_0[1]),.din(n11563));
	jspl jspl_w_n11567_0(.douta(w_n11567_0[0]),.doutb(w_n11567_0[1]),.din(n11567));
	jspl3 jspl3_w_n11569_0(.douta(w_n11569_0[0]),.doutb(w_n11569_0[1]),.doutc(w_n11569_0[2]),.din(n11569));
	jspl jspl_w_n11570_0(.douta(w_n11570_0[0]),.doutb(w_n11570_0[1]),.din(n11570));
	jspl jspl_w_n11574_0(.douta(w_n11574_0[0]),.doutb(w_n11574_0[1]),.din(n11574));
	jspl jspl_w_n11575_0(.douta(w_n11575_0[0]),.doutb(w_n11575_0[1]),.din(n11575));
	jspl3 jspl3_w_n11577_0(.douta(w_n11577_0[0]),.doutb(w_n11577_0[1]),.doutc(w_n11577_0[2]),.din(n11577));
	jspl jspl_w_n11578_0(.douta(w_n11578_0[0]),.doutb(w_n11578_0[1]),.din(n11578));
	jspl jspl_w_n11582_0(.douta(w_n11582_0[0]),.doutb(w_n11582_0[1]),.din(n11582));
	jspl3 jspl3_w_n11584_0(.douta(w_n11584_0[0]),.doutb(w_n11584_0[1]),.doutc(w_n11584_0[2]),.din(n11584));
	jspl jspl_w_n11585_0(.douta(w_n11585_0[0]),.doutb(w_n11585_0[1]),.din(n11585));
	jspl jspl_w_n11589_0(.douta(w_n11589_0[0]),.doutb(w_n11589_0[1]),.din(n11589));
	jspl jspl_w_n11590_0(.douta(w_n11590_0[0]),.doutb(w_n11590_0[1]),.din(n11590));
	jspl3 jspl3_w_n11592_0(.douta(w_n11592_0[0]),.doutb(w_n11592_0[1]),.doutc(w_n11592_0[2]),.din(n11592));
	jspl jspl_w_n11593_0(.douta(w_n11593_0[0]),.doutb(w_n11593_0[1]),.din(n11593));
	jspl jspl_w_n11597_0(.douta(w_n11597_0[0]),.doutb(w_n11597_0[1]),.din(n11597));
	jspl3 jspl3_w_n11599_0(.douta(w_n11599_0[0]),.doutb(w_n11599_0[1]),.doutc(w_n11599_0[2]),.din(n11599));
	jspl jspl_w_n11600_0(.douta(w_n11600_0[0]),.doutb(w_n11600_0[1]),.din(n11600));
	jspl jspl_w_n11604_0(.douta(w_n11604_0[0]),.doutb(w_n11604_0[1]),.din(n11604));
	jspl3 jspl3_w_n11606_0(.douta(w_n11606_0[0]),.doutb(w_n11606_0[1]),.doutc(w_n11606_0[2]),.din(n11606));
	jspl jspl_w_n11607_0(.douta(w_n11607_0[0]),.doutb(w_n11607_0[1]),.din(n11607));
	jspl jspl_w_n11611_0(.douta(w_n11611_0[0]),.doutb(w_n11611_0[1]),.din(n11611));
	jspl3 jspl3_w_n11613_0(.douta(w_n11613_0[0]),.doutb(w_n11613_0[1]),.doutc(w_n11613_0[2]),.din(n11613));
	jspl jspl_w_n11614_0(.douta(w_n11614_0[0]),.doutb(w_n11614_0[1]),.din(n11614));
	jspl jspl_w_n11618_0(.douta(w_n11618_0[0]),.doutb(w_n11618_0[1]),.din(n11618));
	jspl jspl_w_n11619_0(.douta(w_n11619_0[0]),.doutb(w_n11619_0[1]),.din(n11619));
	jspl3 jspl3_w_n11621_0(.douta(w_n11621_0[0]),.doutb(w_n11621_0[1]),.doutc(w_n11621_0[2]),.din(n11621));
	jspl jspl_w_n11622_0(.douta(w_n11622_0[0]),.doutb(w_n11622_0[1]),.din(n11622));
	jspl jspl_w_n11626_0(.douta(w_n11626_0[0]),.doutb(w_n11626_0[1]),.din(n11626));
	jspl jspl_w_n11627_0(.douta(w_n11627_0[0]),.doutb(w_n11627_0[1]),.din(n11627));
	jspl3 jspl3_w_n11629_0(.douta(w_n11629_0[0]),.doutb(w_n11629_0[1]),.doutc(w_n11629_0[2]),.din(n11629));
	jspl jspl_w_n11630_0(.douta(w_n11630_0[0]),.doutb(w_n11630_0[1]),.din(n11630));
	jspl jspl_w_n11634_0(.douta(w_n11634_0[0]),.doutb(w_n11634_0[1]),.din(n11634));
	jspl jspl_w_n11635_0(.douta(w_n11635_0[0]),.doutb(w_n11635_0[1]),.din(n11635));
	jspl3 jspl3_w_n11637_0(.douta(w_n11637_0[0]),.doutb(w_n11637_0[1]),.doutc(w_n11637_0[2]),.din(n11637));
	jspl jspl_w_n11638_0(.douta(w_n11638_0[0]),.doutb(w_n11638_0[1]),.din(n11638));
	jspl jspl_w_n11642_0(.douta(w_n11642_0[0]),.doutb(w_n11642_0[1]),.din(n11642));
	jspl3 jspl3_w_n11644_0(.douta(w_n11644_0[0]),.doutb(w_n11644_0[1]),.doutc(w_n11644_0[2]),.din(n11644));
	jspl jspl_w_n11645_0(.douta(w_n11645_0[0]),.doutb(w_n11645_0[1]),.din(n11645));
	jspl3 jspl3_w_n11649_0(.douta(w_n11649_0[0]),.doutb(w_n11649_0[1]),.doutc(w_n11649_0[2]),.din(n11649));
	jspl jspl_w_n11652_0(.douta(w_n11652_0[0]),.doutb(w_n11652_0[1]),.din(n11652));
	jspl3 jspl3_w_n11653_0(.douta(w_n11653_0[0]),.doutb(w_n11653_0[1]),.doutc(w_n11653_0[2]),.din(n11653));
	jspl jspl_w_n11653_1(.douta(w_n11653_1[0]),.doutb(w_n11653_1[1]),.din(w_n11653_0[0]));
	jspl3 jspl3_w_n11654_0(.douta(w_n11654_0[0]),.doutb(w_n11654_0[1]),.doutc(w_n11654_0[2]),.din(n11654));
	jspl jspl_w_n11679_0(.douta(w_n11679_0[0]),.doutb(w_n11679_0[1]),.din(n11679));
	jspl jspl_w_n11704_0(.douta(w_n11704_0[0]),.doutb(w_n11704_0[1]),.din(n11704));
	jspl jspl_w_n11711_0(.douta(w_n11711_0[0]),.doutb(w_n11711_0[1]),.din(n11711));
	jspl jspl_w_n11724_0(.douta(w_n11724_0[0]),.doutb(w_n11724_0[1]),.din(n11724));
	jspl jspl_w_n11731_0(.douta(w_n11731_0[0]),.doutb(w_n11731_0[1]),.din(n11731));
	jspl jspl_w_n11744_0(.douta(w_n11744_0[0]),.doutb(w_n11744_0[1]),.din(n11744));
	jspl jspl_w_n11769_0(.douta(w_n11769_0[0]),.doutb(w_n11769_0[1]),.din(n11769));
	jspl jspl_w_n11776_0(.douta(w_n11776_0[0]),.doutb(w_n11776_0[1]),.din(n11776));
	jspl jspl_w_n11789_0(.douta(w_n11789_0[0]),.doutb(w_n11789_0[1]),.din(n11789));
	jspl jspl_w_n11796_0(.douta(w_n11796_0[0]),.doutb(w_n11796_0[1]),.din(n11796));
	jspl jspl_w_n11803_0(.douta(w_n11803_0[0]),.doutb(w_n11803_0[1]),.din(n11803));
	jspl jspl_w_n11810_0(.douta(w_n11810_0[0]),.doutb(w_n11810_0[1]),.din(n11810));
	jspl jspl_w_n11814_0(.douta(w_n11814_0[0]),.doutb(w_n11814_0[1]),.din(n11814));
	jspl jspl_w_n11818_0(.douta(w_n11818_0[0]),.doutb(w_n11818_0[1]),.din(n11818));
	jspl jspl_w_n11831_0(.douta(w_n11831_0[0]),.doutb(w_n11831_0[1]),.din(n11831));
	jspl jspl_w_n11836_0(.douta(w_n11836_0[0]),.doutb(w_n11836_0[1]),.din(n11836));
	jspl jspl_w_n11837_0(.douta(w_n11837_0[0]),.doutb(w_n11837_0[1]),.din(n11837));
	jspl jspl_w_n11838_0(.douta(w_n11838_0[0]),.doutb(w_n11838_0[1]),.din(n11838));
	jspl jspl_w_n11840_0(.douta(w_n11840_0[0]),.doutb(w_n11840_0[1]),.din(n11840));
	jspl jspl_w_n11842_0(.douta(w_n11842_0[0]),.doutb(w_n11842_0[1]),.din(n11842));
	jspl jspl_w_n11845_0(.douta(w_n11845_0[0]),.doutb(w_n11845_0[1]),.din(n11845));
	jspl jspl_w_n11846_0(.douta(w_n11846_0[0]),.doutb(w_n11846_0[1]),.din(n11846));
	jspl jspl_w_n11847_0(.douta(w_n11847_0[0]),.doutb(w_n11847_0[1]),.din(n11847));
	jspl jspl_w_n11851_0(.douta(w_n11851_0[0]),.doutb(w_n11851_0[1]),.din(n11851));
	jspl jspl_w_n11856_0(.douta(w_n11856_0[0]),.doutb(w_n11856_0[1]),.din(n11856));
	jspl3 jspl3_w_n11858_0(.douta(w_n11858_0[0]),.doutb(w_n11858_0[1]),.doutc(w_n11858_0[2]),.din(n11858));
	jspl3 jspl3_w_n11858_1(.douta(w_n11858_1[0]),.doutb(w_n11858_1[1]),.doutc(w_n11858_1[2]),.din(w_n11858_0[0]));
	jspl3 jspl3_w_n11858_2(.douta(w_n11858_2[0]),.doutb(w_n11858_2[1]),.doutc(w_n11858_2[2]),.din(w_n11858_0[1]));
	jspl3 jspl3_w_n11858_3(.douta(w_n11858_3[0]),.doutb(w_n11858_3[1]),.doutc(w_n11858_3[2]),.din(w_n11858_0[2]));
	jspl3 jspl3_w_n11858_4(.douta(w_n11858_4[0]),.doutb(w_n11858_4[1]),.doutc(w_n11858_4[2]),.din(w_n11858_1[0]));
	jspl3 jspl3_w_n11858_5(.douta(w_n11858_5[0]),.doutb(w_n11858_5[1]),.doutc(w_n11858_5[2]),.din(w_n11858_1[1]));
	jspl3 jspl3_w_n11858_6(.douta(w_n11858_6[0]),.doutb(w_n11858_6[1]),.doutc(w_n11858_6[2]),.din(w_n11858_1[2]));
	jspl3 jspl3_w_n11858_7(.douta(w_n11858_7[0]),.doutb(w_n11858_7[1]),.doutc(w_n11858_7[2]),.din(w_n11858_2[0]));
	jspl3 jspl3_w_n11858_8(.douta(w_n11858_8[0]),.doutb(w_n11858_8[1]),.doutc(w_n11858_8[2]),.din(w_n11858_2[1]));
	jspl3 jspl3_w_n11858_9(.douta(w_n11858_9[0]),.doutb(w_n11858_9[1]),.doutc(w_n11858_9[2]),.din(w_n11858_2[2]));
	jspl3 jspl3_w_n11858_10(.douta(w_n11858_10[0]),.doutb(w_n11858_10[1]),.doutc(w_n11858_10[2]),.din(w_n11858_3[0]));
	jspl3 jspl3_w_n11858_11(.douta(w_n11858_11[0]),.doutb(w_n11858_11[1]),.doutc(w_n11858_11[2]),.din(w_n11858_3[1]));
	jspl3 jspl3_w_n11858_12(.douta(w_n11858_12[0]),.doutb(w_n11858_12[1]),.doutc(w_n11858_12[2]),.din(w_n11858_3[2]));
	jspl3 jspl3_w_n11858_13(.douta(w_n11858_13[0]),.doutb(w_n11858_13[1]),.doutc(w_n11858_13[2]),.din(w_n11858_4[0]));
	jspl3 jspl3_w_n11858_14(.douta(w_n11858_14[0]),.doutb(w_n11858_14[1]),.doutc(w_n11858_14[2]),.din(w_n11858_4[1]));
	jspl3 jspl3_w_n11858_15(.douta(w_n11858_15[0]),.doutb(w_n11858_15[1]),.doutc(w_n11858_15[2]),.din(w_n11858_4[2]));
	jspl3 jspl3_w_n11858_16(.douta(w_n11858_16[0]),.doutb(w_n11858_16[1]),.doutc(w_n11858_16[2]),.din(w_n11858_5[0]));
	jspl3 jspl3_w_n11858_17(.douta(w_n11858_17[0]),.doutb(w_n11858_17[1]),.doutc(w_n11858_17[2]),.din(w_n11858_5[1]));
	jspl3 jspl3_w_n11858_18(.douta(w_n11858_18[0]),.doutb(w_n11858_18[1]),.doutc(w_n11858_18[2]),.din(w_n11858_5[2]));
	jspl3 jspl3_w_n11858_19(.douta(w_n11858_19[0]),.doutb(w_n11858_19[1]),.doutc(w_n11858_19[2]),.din(w_n11858_6[0]));
	jspl3 jspl3_w_n11858_20(.douta(w_n11858_20[0]),.doutb(w_n11858_20[1]),.doutc(w_n11858_20[2]),.din(w_n11858_6[1]));
	jspl3 jspl3_w_n11858_21(.douta(w_n11858_21[0]),.doutb(w_n11858_21[1]),.doutc(w_n11858_21[2]),.din(w_n11858_6[2]));
	jspl3 jspl3_w_n11858_22(.douta(w_n11858_22[0]),.doutb(w_n11858_22[1]),.doutc(w_n11858_22[2]),.din(w_n11858_7[0]));
	jspl3 jspl3_w_n11858_23(.douta(w_n11858_23[0]),.doutb(w_n11858_23[1]),.doutc(w_n11858_23[2]),.din(w_n11858_7[1]));
	jspl3 jspl3_w_n11858_24(.douta(w_n11858_24[0]),.doutb(w_n11858_24[1]),.doutc(w_n11858_24[2]),.din(w_n11858_7[2]));
	jspl3 jspl3_w_n11858_25(.douta(w_n11858_25[0]),.doutb(w_n11858_25[1]),.doutc(w_n11858_25[2]),.din(w_n11858_8[0]));
	jspl3 jspl3_w_n11858_26(.douta(w_n11858_26[0]),.doutb(w_n11858_26[1]),.doutc(w_n11858_26[2]),.din(w_n11858_8[1]));
	jspl3 jspl3_w_n11858_27(.douta(w_n11858_27[0]),.doutb(w_n11858_27[1]),.doutc(w_n11858_27[2]),.din(w_n11858_8[2]));
	jspl3 jspl3_w_n11858_28(.douta(w_n11858_28[0]),.doutb(w_n11858_28[1]),.doutc(w_n11858_28[2]),.din(w_n11858_9[0]));
	jspl3 jspl3_w_n11858_29(.douta(w_n11858_29[0]),.doutb(w_n11858_29[1]),.doutc(w_n11858_29[2]),.din(w_n11858_9[1]));
	jspl3 jspl3_w_n11858_30(.douta(w_n11858_30[0]),.doutb(w_n11858_30[1]),.doutc(w_n11858_30[2]),.din(w_n11858_9[2]));
	jspl3 jspl3_w_n11858_31(.douta(w_n11858_31[0]),.doutb(w_n11858_31[1]),.doutc(w_n11858_31[2]),.din(w_n11858_10[0]));
	jspl3 jspl3_w_n11858_32(.douta(w_n11858_32[0]),.doutb(w_n11858_32[1]),.doutc(w_n11858_32[2]),.din(w_n11858_10[1]));
	jspl3 jspl3_w_n11858_33(.douta(w_n11858_33[0]),.doutb(w_n11858_33[1]),.doutc(w_n11858_33[2]),.din(w_n11858_10[2]));
	jspl3 jspl3_w_n11858_34(.douta(w_n11858_34[0]),.doutb(w_n11858_34[1]),.doutc(w_n11858_34[2]),.din(w_n11858_11[0]));
	jspl3 jspl3_w_n11858_35(.douta(w_n11858_35[0]),.doutb(w_n11858_35[1]),.doutc(w_n11858_35[2]),.din(w_n11858_11[1]));
	jspl3 jspl3_w_n11858_36(.douta(w_n11858_36[0]),.doutb(w_n11858_36[1]),.doutc(w_n11858_36[2]),.din(w_n11858_11[2]));
	jspl3 jspl3_w_n11858_37(.douta(w_n11858_37[0]),.doutb(w_n11858_37[1]),.doutc(w_n11858_37[2]),.din(w_n11858_12[0]));
	jspl3 jspl3_w_n11858_38(.douta(w_n11858_38[0]),.doutb(w_n11858_38[1]),.doutc(w_n11858_38[2]),.din(w_n11858_12[1]));
	jspl3 jspl3_w_n11858_39(.douta(w_n11858_39[0]),.doutb(w_n11858_39[1]),.doutc(w_n11858_39[2]),.din(w_n11858_12[2]));
	jspl3 jspl3_w_n11858_40(.douta(w_n11858_40[0]),.doutb(w_n11858_40[1]),.doutc(w_n11858_40[2]),.din(w_n11858_13[0]));
	jspl3 jspl3_w_n11858_41(.douta(w_n11858_41[0]),.doutb(w_n11858_41[1]),.doutc(w_n11858_41[2]),.din(w_n11858_13[1]));
	jspl3 jspl3_w_n11858_42(.douta(w_n11858_42[0]),.doutb(w_n11858_42[1]),.doutc(w_n11858_42[2]),.din(w_n11858_13[2]));
	jspl3 jspl3_w_n11858_43(.douta(w_n11858_43[0]),.doutb(w_n11858_43[1]),.doutc(w_n11858_43[2]),.din(w_n11858_14[0]));
	jspl3 jspl3_w_n11858_44(.douta(w_n11858_44[0]),.doutb(w_n11858_44[1]),.doutc(w_n11858_44[2]),.din(w_n11858_14[1]));
	jspl jspl_w_n11858_45(.douta(w_n11858_45[0]),.doutb(w_n11858_45[1]),.din(w_n11858_14[2]));
	jspl jspl_w_n11861_0(.douta(w_n11861_0[0]),.doutb(w_n11861_0[1]),.din(n11861));
	jspl3 jspl3_w_n11862_0(.douta(w_n11862_0[0]),.doutb(w_n11862_0[1]),.doutc(w_n11862_0[2]),.din(n11862));
	jspl3 jspl3_w_n11864_0(.douta(w_n11864_0[0]),.doutb(w_n11864_0[1]),.doutc(w_n11864_0[2]),.din(n11864));
	jspl3 jspl3_w_n11864_1(.douta(w_n11864_1[0]),.doutb(w_n11864_1[1]),.doutc(w_n11864_1[2]),.din(w_n11864_0[0]));
	jspl jspl_w_n11865_0(.douta(w_n11865_0[0]),.doutb(w_n11865_0[1]),.din(n11865));
	jspl3 jspl3_w_n11866_0(.douta(w_n11866_0[0]),.doutb(w_n11866_0[1]),.doutc(w_n11866_0[2]),.din(n11866));
	jspl jspl_w_n11867_0(.douta(w_n11867_0[0]),.doutb(w_n11867_0[1]),.din(n11867));
	jspl3 jspl3_w_n11869_0(.douta(w_n11869_0[0]),.doutb(w_n11869_0[1]),.doutc(w_n11869_0[2]),.din(n11869));
	jspl jspl_w_n11870_0(.douta(w_n11870_0[0]),.doutb(w_n11870_0[1]),.din(n11870));
	jspl3 jspl3_w_n11877_0(.douta(w_n11877_0[0]),.doutb(w_n11877_0[1]),.doutc(w_n11877_0[2]),.din(n11877));
	jspl jspl_w_n11878_0(.douta(w_n11878_0[0]),.doutb(w_n11878_0[1]),.din(n11878));
	jspl jspl_w_n11881_0(.douta(w_n11881_0[0]),.doutb(w_n11881_0[1]),.din(n11881));
	jspl3 jspl3_w_n11886_0(.douta(w_n11886_0[0]),.doutb(w_n11886_0[1]),.doutc(w_n11886_0[2]),.din(n11886));
	jspl3 jspl3_w_n11888_0(.douta(w_n11888_0[0]),.doutb(w_n11888_0[1]),.doutc(w_n11888_0[2]),.din(n11888));
	jspl jspl_w_n11889_0(.douta(w_n11889_0[0]),.doutb(w_n11889_0[1]),.din(n11889));
	jspl3 jspl3_w_n11893_0(.douta(w_n11893_0[0]),.doutb(w_n11893_0[1]),.doutc(w_n11893_0[2]),.din(n11893));
	jspl3 jspl3_w_n11896_0(.douta(w_n11896_0[0]),.doutb(w_n11896_0[1]),.doutc(w_n11896_0[2]),.din(n11896));
	jspl jspl_w_n11897_0(.douta(w_n11897_0[0]),.doutb(w_n11897_0[1]),.din(n11897));
	jspl3 jspl3_w_n11901_0(.douta(w_n11901_0[0]),.doutb(w_n11901_0[1]),.doutc(w_n11901_0[2]),.din(n11901));
	jspl3 jspl3_w_n11903_0(.douta(w_n11903_0[0]),.doutb(w_n11903_0[1]),.doutc(w_n11903_0[2]),.din(n11903));
	jspl jspl_w_n11904_0(.douta(w_n11904_0[0]),.doutb(w_n11904_0[1]),.din(n11904));
	jspl3 jspl3_w_n11908_0(.douta(w_n11908_0[0]),.doutb(w_n11908_0[1]),.doutc(w_n11908_0[2]),.din(n11908));
	jspl3 jspl3_w_n11911_0(.douta(w_n11911_0[0]),.doutb(w_n11911_0[1]),.doutc(w_n11911_0[2]),.din(n11911));
	jspl jspl_w_n11912_0(.douta(w_n11912_0[0]),.doutb(w_n11912_0[1]),.din(n11912));
	jspl3 jspl3_w_n11916_0(.douta(w_n11916_0[0]),.doutb(w_n11916_0[1]),.doutc(w_n11916_0[2]),.din(n11916));
	jspl3 jspl3_w_n11918_0(.douta(w_n11918_0[0]),.doutb(w_n11918_0[1]),.doutc(w_n11918_0[2]),.din(n11918));
	jspl jspl_w_n11919_0(.douta(w_n11919_0[0]),.doutb(w_n11919_0[1]),.din(n11919));
	jspl3 jspl3_w_n11923_0(.douta(w_n11923_0[0]),.doutb(w_n11923_0[1]),.doutc(w_n11923_0[2]),.din(n11923));
	jspl3 jspl3_w_n11925_0(.douta(w_n11925_0[0]),.doutb(w_n11925_0[1]),.doutc(w_n11925_0[2]),.din(n11925));
	jspl jspl_w_n11926_0(.douta(w_n11926_0[0]),.doutb(w_n11926_0[1]),.din(n11926));
	jspl3 jspl3_w_n11930_0(.douta(w_n11930_0[0]),.doutb(w_n11930_0[1]),.doutc(w_n11930_0[2]),.din(n11930));
	jspl3 jspl3_w_n11932_0(.douta(w_n11932_0[0]),.doutb(w_n11932_0[1]),.doutc(w_n11932_0[2]),.din(n11932));
	jspl jspl_w_n11933_0(.douta(w_n11933_0[0]),.doutb(w_n11933_0[1]),.din(n11933));
	jspl3 jspl3_w_n11937_0(.douta(w_n11937_0[0]),.doutb(w_n11937_0[1]),.doutc(w_n11937_0[2]),.din(n11937));
	jspl3 jspl3_w_n11940_0(.douta(w_n11940_0[0]),.doutb(w_n11940_0[1]),.doutc(w_n11940_0[2]),.din(n11940));
	jspl jspl_w_n11941_0(.douta(w_n11941_0[0]),.doutb(w_n11941_0[1]),.din(n11941));
	jspl3 jspl3_w_n11945_0(.douta(w_n11945_0[0]),.doutb(w_n11945_0[1]),.doutc(w_n11945_0[2]),.din(n11945));
	jspl3 jspl3_w_n11947_0(.douta(w_n11947_0[0]),.doutb(w_n11947_0[1]),.doutc(w_n11947_0[2]),.din(n11947));
	jspl jspl_w_n11948_0(.douta(w_n11948_0[0]),.doutb(w_n11948_0[1]),.din(n11948));
	jspl3 jspl3_w_n11952_0(.douta(w_n11952_0[0]),.doutb(w_n11952_0[1]),.doutc(w_n11952_0[2]),.din(n11952));
	jspl3 jspl3_w_n11955_0(.douta(w_n11955_0[0]),.doutb(w_n11955_0[1]),.doutc(w_n11955_0[2]),.din(n11955));
	jspl jspl_w_n11956_0(.douta(w_n11956_0[0]),.doutb(w_n11956_0[1]),.din(n11956));
	jspl3 jspl3_w_n11960_0(.douta(w_n11960_0[0]),.doutb(w_n11960_0[1]),.doutc(w_n11960_0[2]),.din(n11960));
	jspl3 jspl3_w_n11962_0(.douta(w_n11962_0[0]),.doutb(w_n11962_0[1]),.doutc(w_n11962_0[2]),.din(n11962));
	jspl jspl_w_n11963_0(.douta(w_n11963_0[0]),.doutb(w_n11963_0[1]),.din(n11963));
	jspl3 jspl3_w_n11967_0(.douta(w_n11967_0[0]),.doutb(w_n11967_0[1]),.doutc(w_n11967_0[2]),.din(n11967));
	jspl3 jspl3_w_n11969_0(.douta(w_n11969_0[0]),.doutb(w_n11969_0[1]),.doutc(w_n11969_0[2]),.din(n11969));
	jspl jspl_w_n11970_0(.douta(w_n11970_0[0]),.doutb(w_n11970_0[1]),.din(n11970));
	jspl3 jspl3_w_n11974_0(.douta(w_n11974_0[0]),.doutb(w_n11974_0[1]),.doutc(w_n11974_0[2]),.din(n11974));
	jspl3 jspl3_w_n11976_0(.douta(w_n11976_0[0]),.doutb(w_n11976_0[1]),.doutc(w_n11976_0[2]),.din(n11976));
	jspl jspl_w_n11977_0(.douta(w_n11977_0[0]),.doutb(w_n11977_0[1]),.din(n11977));
	jspl3 jspl3_w_n11981_0(.douta(w_n11981_0[0]),.doutb(w_n11981_0[1]),.doutc(w_n11981_0[2]),.din(n11981));
	jspl3 jspl3_w_n11984_0(.douta(w_n11984_0[0]),.doutb(w_n11984_0[1]),.doutc(w_n11984_0[2]),.din(n11984));
	jspl jspl_w_n11985_0(.douta(w_n11985_0[0]),.doutb(w_n11985_0[1]),.din(n11985));
	jspl3 jspl3_w_n11989_0(.douta(w_n11989_0[0]),.doutb(w_n11989_0[1]),.doutc(w_n11989_0[2]),.din(n11989));
	jspl3 jspl3_w_n11991_0(.douta(w_n11991_0[0]),.doutb(w_n11991_0[1]),.doutc(w_n11991_0[2]),.din(n11991));
	jspl jspl_w_n11992_0(.douta(w_n11992_0[0]),.doutb(w_n11992_0[1]),.din(n11992));
	jspl3 jspl3_w_n11996_0(.douta(w_n11996_0[0]),.doutb(w_n11996_0[1]),.doutc(w_n11996_0[2]),.din(n11996));
	jspl3 jspl3_w_n11998_0(.douta(w_n11998_0[0]),.doutb(w_n11998_0[1]),.doutc(w_n11998_0[2]),.din(n11998));
	jspl jspl_w_n11999_0(.douta(w_n11999_0[0]),.doutb(w_n11999_0[1]),.din(n11999));
	jspl3 jspl3_w_n12003_0(.douta(w_n12003_0[0]),.doutb(w_n12003_0[1]),.doutc(w_n12003_0[2]),.din(n12003));
	jspl3 jspl3_w_n12005_0(.douta(w_n12005_0[0]),.doutb(w_n12005_0[1]),.doutc(w_n12005_0[2]),.din(n12005));
	jspl jspl_w_n12006_0(.douta(w_n12006_0[0]),.doutb(w_n12006_0[1]),.din(n12006));
	jspl3 jspl3_w_n12010_0(.douta(w_n12010_0[0]),.doutb(w_n12010_0[1]),.doutc(w_n12010_0[2]),.din(n12010));
	jspl3 jspl3_w_n12012_0(.douta(w_n12012_0[0]),.doutb(w_n12012_0[1]),.doutc(w_n12012_0[2]),.din(n12012));
	jspl jspl_w_n12013_0(.douta(w_n12013_0[0]),.doutb(w_n12013_0[1]),.din(n12013));
	jspl3 jspl3_w_n12017_0(.douta(w_n12017_0[0]),.doutb(w_n12017_0[1]),.doutc(w_n12017_0[2]),.din(n12017));
	jspl3 jspl3_w_n12019_0(.douta(w_n12019_0[0]),.doutb(w_n12019_0[1]),.doutc(w_n12019_0[2]),.din(n12019));
	jspl jspl_w_n12020_0(.douta(w_n12020_0[0]),.doutb(w_n12020_0[1]),.din(n12020));
	jspl3 jspl3_w_n12023_0(.douta(w_n12023_0[0]),.doutb(w_n12023_0[1]),.doutc(w_n12023_0[2]),.din(n12023));
	jspl3 jspl3_w_n12027_0(.douta(w_n12027_0[0]),.doutb(w_n12027_0[1]),.doutc(w_n12027_0[2]),.din(n12027));
	jspl jspl_w_n12028_0(.douta(w_n12028_0[0]),.doutb(w_n12028_0[1]),.din(n12028));
	jspl3 jspl3_w_n12032_0(.douta(w_n12032_0[0]),.doutb(w_n12032_0[1]),.doutc(w_n12032_0[2]),.din(n12032));
	jspl3 jspl3_w_n12034_0(.douta(w_n12034_0[0]),.doutb(w_n12034_0[1]),.doutc(w_n12034_0[2]),.din(n12034));
	jspl jspl_w_n12035_0(.douta(w_n12035_0[0]),.doutb(w_n12035_0[1]),.din(n12035));
	jspl3 jspl3_w_n12039_0(.douta(w_n12039_0[0]),.doutb(w_n12039_0[1]),.doutc(w_n12039_0[2]),.din(n12039));
	jspl3 jspl3_w_n12042_0(.douta(w_n12042_0[0]),.doutb(w_n12042_0[1]),.doutc(w_n12042_0[2]),.din(n12042));
	jspl jspl_w_n12043_0(.douta(w_n12043_0[0]),.doutb(w_n12043_0[1]),.din(n12043));
	jspl3 jspl3_w_n12047_0(.douta(w_n12047_0[0]),.doutb(w_n12047_0[1]),.doutc(w_n12047_0[2]),.din(n12047));
	jspl3 jspl3_w_n12049_0(.douta(w_n12049_0[0]),.doutb(w_n12049_0[1]),.doutc(w_n12049_0[2]),.din(n12049));
	jspl jspl_w_n12050_0(.douta(w_n12050_0[0]),.doutb(w_n12050_0[1]),.din(n12050));
	jspl3 jspl3_w_n12054_0(.douta(w_n12054_0[0]),.doutb(w_n12054_0[1]),.doutc(w_n12054_0[2]),.din(n12054));
	jspl3 jspl3_w_n12057_0(.douta(w_n12057_0[0]),.doutb(w_n12057_0[1]),.doutc(w_n12057_0[2]),.din(n12057));
	jspl jspl_w_n12058_0(.douta(w_n12058_0[0]),.doutb(w_n12058_0[1]),.din(n12058));
	jspl3 jspl3_w_n12062_0(.douta(w_n12062_0[0]),.doutb(w_n12062_0[1]),.doutc(w_n12062_0[2]),.din(n12062));
	jspl3 jspl3_w_n12064_0(.douta(w_n12064_0[0]),.doutb(w_n12064_0[1]),.doutc(w_n12064_0[2]),.din(n12064));
	jspl jspl_w_n12065_0(.douta(w_n12065_0[0]),.doutb(w_n12065_0[1]),.din(n12065));
	jspl3 jspl3_w_n12069_0(.douta(w_n12069_0[0]),.doutb(w_n12069_0[1]),.doutc(w_n12069_0[2]),.din(n12069));
	jspl3 jspl3_w_n12071_0(.douta(w_n12071_0[0]),.doutb(w_n12071_0[1]),.doutc(w_n12071_0[2]),.din(n12071));
	jspl jspl_w_n12072_0(.douta(w_n12072_0[0]),.doutb(w_n12072_0[1]),.din(n12072));
	jspl3 jspl3_w_n12076_0(.douta(w_n12076_0[0]),.doutb(w_n12076_0[1]),.doutc(w_n12076_0[2]),.din(n12076));
	jspl3 jspl3_w_n12078_0(.douta(w_n12078_0[0]),.doutb(w_n12078_0[1]),.doutc(w_n12078_0[2]),.din(n12078));
	jspl jspl_w_n12079_0(.douta(w_n12079_0[0]),.doutb(w_n12079_0[1]),.din(n12079));
	jspl3 jspl3_w_n12083_0(.douta(w_n12083_0[0]),.doutb(w_n12083_0[1]),.doutc(w_n12083_0[2]),.din(n12083));
	jspl3 jspl3_w_n12086_0(.douta(w_n12086_0[0]),.doutb(w_n12086_0[1]),.doutc(w_n12086_0[2]),.din(n12086));
	jspl jspl_w_n12087_0(.douta(w_n12087_0[0]),.doutb(w_n12087_0[1]),.din(n12087));
	jspl3 jspl3_w_n12091_0(.douta(w_n12091_0[0]),.doutb(w_n12091_0[1]),.doutc(w_n12091_0[2]),.din(n12091));
	jspl3 jspl3_w_n12093_0(.douta(w_n12093_0[0]),.doutb(w_n12093_0[1]),.doutc(w_n12093_0[2]),.din(n12093));
	jspl jspl_w_n12094_0(.douta(w_n12094_0[0]),.doutb(w_n12094_0[1]),.din(n12094));
	jspl3 jspl3_w_n12098_0(.douta(w_n12098_0[0]),.doutb(w_n12098_0[1]),.doutc(w_n12098_0[2]),.din(n12098));
	jspl3 jspl3_w_n12101_0(.douta(w_n12101_0[0]),.doutb(w_n12101_0[1]),.doutc(w_n12101_0[2]),.din(n12101));
	jspl jspl_w_n12102_0(.douta(w_n12102_0[0]),.doutb(w_n12102_0[1]),.din(n12102));
	jspl3 jspl3_w_n12106_0(.douta(w_n12106_0[0]),.doutb(w_n12106_0[1]),.doutc(w_n12106_0[2]),.din(n12106));
	jspl3 jspl3_w_n12108_0(.douta(w_n12108_0[0]),.doutb(w_n12108_0[1]),.doutc(w_n12108_0[2]),.din(n12108));
	jspl jspl_w_n12109_0(.douta(w_n12109_0[0]),.doutb(w_n12109_0[1]),.din(n12109));
	jspl3 jspl3_w_n12113_0(.douta(w_n12113_0[0]),.doutb(w_n12113_0[1]),.doutc(w_n12113_0[2]),.din(n12113));
	jspl3 jspl3_w_n12116_0(.douta(w_n12116_0[0]),.doutb(w_n12116_0[1]),.doutc(w_n12116_0[2]),.din(n12116));
	jspl jspl_w_n12117_0(.douta(w_n12117_0[0]),.doutb(w_n12117_0[1]),.din(n12117));
	jspl3 jspl3_w_n12121_0(.douta(w_n12121_0[0]),.doutb(w_n12121_0[1]),.doutc(w_n12121_0[2]),.din(n12121));
	jspl3 jspl3_w_n12123_0(.douta(w_n12123_0[0]),.doutb(w_n12123_0[1]),.doutc(w_n12123_0[2]),.din(n12123));
	jspl jspl_w_n12124_0(.douta(w_n12124_0[0]),.doutb(w_n12124_0[1]),.din(n12124));
	jspl3 jspl3_w_n12128_0(.douta(w_n12128_0[0]),.doutb(w_n12128_0[1]),.doutc(w_n12128_0[2]),.din(n12128));
	jspl3 jspl3_w_n12131_0(.douta(w_n12131_0[0]),.doutb(w_n12131_0[1]),.doutc(w_n12131_0[2]),.din(n12131));
	jspl jspl_w_n12132_0(.douta(w_n12132_0[0]),.doutb(w_n12132_0[1]),.din(n12132));
	jspl3 jspl3_w_n12136_0(.douta(w_n12136_0[0]),.doutb(w_n12136_0[1]),.doutc(w_n12136_0[2]),.din(n12136));
	jspl3 jspl3_w_n12139_0(.douta(w_n12139_0[0]),.doutb(w_n12139_0[1]),.doutc(w_n12139_0[2]),.din(n12139));
	jspl jspl_w_n12140_0(.douta(w_n12140_0[0]),.doutb(w_n12140_0[1]),.din(n12140));
	jspl3 jspl3_w_n12144_0(.douta(w_n12144_0[0]),.doutb(w_n12144_0[1]),.doutc(w_n12144_0[2]),.din(n12144));
	jspl3 jspl3_w_n12147_0(.douta(w_n12147_0[0]),.doutb(w_n12147_0[1]),.doutc(w_n12147_0[2]),.din(n12147));
	jspl jspl_w_n12148_0(.douta(w_n12148_0[0]),.doutb(w_n12148_0[1]),.din(n12148));
	jspl3 jspl3_w_n12152_0(.douta(w_n12152_0[0]),.doutb(w_n12152_0[1]),.doutc(w_n12152_0[2]),.din(n12152));
	jspl3 jspl3_w_n12154_0(.douta(w_n12154_0[0]),.doutb(w_n12154_0[1]),.doutc(w_n12154_0[2]),.din(n12154));
	jspl jspl_w_n12155_0(.douta(w_n12155_0[0]),.doutb(w_n12155_0[1]),.din(n12155));
	jspl3 jspl3_w_n12159_0(.douta(w_n12159_0[0]),.doutb(w_n12159_0[1]),.doutc(w_n12159_0[2]),.din(n12159));
	jspl3 jspl3_w_n12161_0(.douta(w_n12161_0[0]),.doutb(w_n12161_0[1]),.doutc(w_n12161_0[2]),.din(n12161));
	jspl jspl_w_n12162_0(.douta(w_n12162_0[0]),.doutb(w_n12162_0[1]),.din(n12162));
	jspl3 jspl3_w_n12166_0(.douta(w_n12166_0[0]),.doutb(w_n12166_0[1]),.doutc(w_n12166_0[2]),.din(n12166));
	jspl3 jspl3_w_n12168_0(.douta(w_n12168_0[0]),.doutb(w_n12168_0[1]),.doutc(w_n12168_0[2]),.din(n12168));
	jspl jspl_w_n12169_0(.douta(w_n12169_0[0]),.doutb(w_n12169_0[1]),.din(n12169));
	jspl3 jspl3_w_n12173_0(.douta(w_n12173_0[0]),.doutb(w_n12173_0[1]),.doutc(w_n12173_0[2]),.din(n12173));
	jspl3 jspl3_w_n12176_0(.douta(w_n12176_0[0]),.doutb(w_n12176_0[1]),.doutc(w_n12176_0[2]),.din(n12176));
	jspl3 jspl3_w_n12177_0(.douta(w_n12177_0[0]),.doutb(w_n12177_0[1]),.doutc(w_n12177_0[2]),.din(n12177));
	jspl jspl_w_n12179_0(.douta(w_n12179_0[0]),.doutb(w_n12179_0[1]),.din(n12179));
	jspl jspl_w_n12180_0(.douta(w_n12180_0[0]),.doutb(w_n12180_0[1]),.din(n12180));
	jspl jspl_w_n12187_0(.douta(w_n12187_0[0]),.doutb(w_n12187_0[1]),.din(n12187));
	jspl jspl_w_n12188_0(.douta(w_n12188_0[0]),.doutb(w_n12188_0[1]),.din(n12188));
	jspl jspl_w_n12190_0(.douta(w_n12190_0[0]),.doutb(w_n12190_0[1]),.din(n12190));
	jspl3 jspl3_w_n12195_0(.douta(w_n12195_0[0]),.doutb(w_n12195_0[1]),.doutc(w_n12195_0[2]),.din(n12195));
	jspl3 jspl3_w_n12196_0(.douta(w_n12196_0[0]),.doutb(w_n12196_0[1]),.doutc(w_n12196_0[2]),.din(n12196));
	jspl3 jspl3_w_n12196_1(.douta(w_n12196_1[0]),.doutb(w_n12196_1[1]),.doutc(w_n12196_1[2]),.din(w_n12196_0[0]));
	jspl jspl_w_n12197_0(.douta(w_n12197_0[0]),.doutb(w_n12197_0[1]),.din(n12197));
	jspl3 jspl3_w_n12198_0(.douta(w_n12198_0[0]),.doutb(w_n12198_0[1]),.doutc(w_n12198_0[2]),.din(n12198));
	jspl jspl_w_n12199_0(.douta(w_n12199_0[0]),.doutb(w_n12199_0[1]),.din(n12199));
	jspl3 jspl3_w_n12201_0(.douta(w_n12201_0[0]),.doutb(w_n12201_0[1]),.doutc(w_n12201_0[2]),.din(n12201));
	jspl jspl_w_n12202_0(.douta(w_n12202_0[0]),.doutb(w_n12202_0[1]),.din(n12202));
	jspl3 jspl3_w_n12207_0(.douta(w_n12207_0[0]),.doutb(w_n12207_0[1]),.doutc(w_n12207_0[2]),.din(n12207));
	jspl jspl_w_n12207_1(.douta(w_n12207_1[0]),.doutb(w_n12207_1[1]),.din(w_n12207_0[0]));
	jspl jspl_w_n12256_0(.douta(w_n12256_0[0]),.doutb(w_n12256_0[1]),.din(n12256));
	jspl jspl_w_n12404_0(.douta(w_n12404_0[0]),.doutb(w_n12404_0[1]),.din(n12404));
	jspl jspl_w_n12407_0(.douta(w_n12407_0[0]),.doutb(w_n12407_0[1]),.din(n12407));
	jspl jspl_w_n12408_0(.douta(w_n12408_0[0]),.doutb(w_n12408_0[1]),.din(n12408));
	jspl3 jspl3_w_n12410_0(.douta(w_n12410_0[0]),.doutb(w_n12410_0[1]),.doutc(w_n12410_0[2]),.din(n12410));
	jspl3 jspl3_w_n12410_1(.douta(w_n12410_1[0]),.doutb(w_n12410_1[1]),.doutc(w_n12410_1[2]),.din(w_n12410_0[0]));
	jspl3 jspl3_w_n12410_2(.douta(w_n12410_2[0]),.doutb(w_n12410_2[1]),.doutc(w_n12410_2[2]),.din(w_n12410_0[1]));
	jspl3 jspl3_w_n12410_3(.douta(w_n12410_3[0]),.doutb(w_n12410_3[1]),.doutc(w_n12410_3[2]),.din(w_n12410_0[2]));
	jspl3 jspl3_w_n12410_4(.douta(w_n12410_4[0]),.doutb(w_n12410_4[1]),.doutc(w_n12410_4[2]),.din(w_n12410_1[0]));
	jspl3 jspl3_w_n12410_5(.douta(w_n12410_5[0]),.doutb(w_n12410_5[1]),.doutc(w_n12410_5[2]),.din(w_n12410_1[1]));
	jspl3 jspl3_w_n12410_6(.douta(w_n12410_6[0]),.doutb(w_n12410_6[1]),.doutc(w_n12410_6[2]),.din(w_n12410_1[2]));
	jspl3 jspl3_w_n12410_7(.douta(w_n12410_7[0]),.doutb(w_n12410_7[1]),.doutc(w_n12410_7[2]),.din(w_n12410_2[0]));
	jspl3 jspl3_w_n12410_8(.douta(w_n12410_8[0]),.doutb(w_n12410_8[1]),.doutc(w_n12410_8[2]),.din(w_n12410_2[1]));
	jspl3 jspl3_w_n12410_9(.douta(w_n12410_9[0]),.doutb(w_n12410_9[1]),.doutc(w_n12410_9[2]),.din(w_n12410_2[2]));
	jspl3 jspl3_w_n12410_10(.douta(w_n12410_10[0]),.doutb(w_n12410_10[1]),.doutc(w_n12410_10[2]),.din(w_n12410_3[0]));
	jspl3 jspl3_w_n12410_11(.douta(w_n12410_11[0]),.doutb(w_n12410_11[1]),.doutc(w_n12410_11[2]),.din(w_n12410_3[1]));
	jspl3 jspl3_w_n12410_12(.douta(w_n12410_12[0]),.doutb(w_n12410_12[1]),.doutc(w_n12410_12[2]),.din(w_n12410_3[2]));
	jspl3 jspl3_w_n12410_13(.douta(w_n12410_13[0]),.doutb(w_n12410_13[1]),.doutc(w_n12410_13[2]),.din(w_n12410_4[0]));
	jspl3 jspl3_w_n12410_14(.douta(w_n12410_14[0]),.doutb(w_n12410_14[1]),.doutc(w_n12410_14[2]),.din(w_n12410_4[1]));
	jspl3 jspl3_w_n12410_15(.douta(w_n12410_15[0]),.doutb(w_n12410_15[1]),.doutc(w_n12410_15[2]),.din(w_n12410_4[2]));
	jspl3 jspl3_w_n12410_16(.douta(w_n12410_16[0]),.doutb(w_n12410_16[1]),.doutc(w_n12410_16[2]),.din(w_n12410_5[0]));
	jspl3 jspl3_w_n12410_17(.douta(w_n12410_17[0]),.doutb(w_n12410_17[1]),.doutc(w_n12410_17[2]),.din(w_n12410_5[1]));
	jspl3 jspl3_w_n12410_18(.douta(w_n12410_18[0]),.doutb(w_n12410_18[1]),.doutc(w_n12410_18[2]),.din(w_n12410_5[2]));
	jspl3 jspl3_w_n12410_19(.douta(w_n12410_19[0]),.doutb(w_n12410_19[1]),.doutc(w_n12410_19[2]),.din(w_n12410_6[0]));
	jspl3 jspl3_w_n12410_20(.douta(w_n12410_20[0]),.doutb(w_n12410_20[1]),.doutc(w_n12410_20[2]),.din(w_n12410_6[1]));
	jspl3 jspl3_w_n12410_21(.douta(w_n12410_21[0]),.doutb(w_n12410_21[1]),.doutc(w_n12410_21[2]),.din(w_n12410_6[2]));
	jspl3 jspl3_w_n12410_22(.douta(w_n12410_22[0]),.doutb(w_n12410_22[1]),.doutc(w_n12410_22[2]),.din(w_n12410_7[0]));
	jspl3 jspl3_w_n12410_23(.douta(w_n12410_23[0]),.doutb(w_n12410_23[1]),.doutc(w_n12410_23[2]),.din(w_n12410_7[1]));
	jspl3 jspl3_w_n12410_24(.douta(w_n12410_24[0]),.doutb(w_n12410_24[1]),.doutc(w_n12410_24[2]),.din(w_n12410_7[2]));
	jspl jspl_w_n12410_25(.douta(w_n12410_25[0]),.doutb(w_n12410_25[1]),.din(w_n12410_8[0]));
	jspl3 jspl3_w_n12414_0(.douta(w_n12414_0[0]),.doutb(w_n12414_0[1]),.doutc(w_n12414_0[2]),.din(n12414));
	jspl jspl_w_n12415_0(.douta(w_n12415_0[0]),.doutb(w_n12415_0[1]),.din(n12415));
	jspl jspl_w_n12417_0(.douta(w_n12417_0[0]),.doutb(w_n12417_0[1]),.din(n12417));
	jspl jspl_w_n12422_0(.douta(w_n12422_0[0]),.doutb(w_n12422_0[1]),.din(n12422));
	jspl jspl_w_n12423_0(.douta(w_n12423_0[0]),.doutb(w_n12423_0[1]),.din(n12423));
	jspl3 jspl3_w_n12425_0(.douta(w_n12425_0[0]),.doutb(w_n12425_0[1]),.doutc(w_n12425_0[2]),.din(n12425));
	jspl jspl_w_n12426_0(.douta(w_n12426_0[0]),.doutb(w_n12426_0[1]),.din(n12426));
	jspl jspl_w_n12430_0(.douta(w_n12430_0[0]),.doutb(w_n12430_0[1]),.din(n12430));
	jspl3 jspl3_w_n12432_0(.douta(w_n12432_0[0]),.doutb(w_n12432_0[1]),.doutc(w_n12432_0[2]),.din(n12432));
	jspl jspl_w_n12433_0(.douta(w_n12433_0[0]),.doutb(w_n12433_0[1]),.din(n12433));
	jspl jspl_w_n12437_0(.douta(w_n12437_0[0]),.doutb(w_n12437_0[1]),.din(n12437));
	jspl jspl_w_n12438_0(.douta(w_n12438_0[0]),.doutb(w_n12438_0[1]),.din(n12438));
	jspl3 jspl3_w_n12440_0(.douta(w_n12440_0[0]),.doutb(w_n12440_0[1]),.doutc(w_n12440_0[2]),.din(n12440));
	jspl jspl_w_n12441_0(.douta(w_n12441_0[0]),.doutb(w_n12441_0[1]),.din(n12441));
	jspl jspl_w_n12445_0(.douta(w_n12445_0[0]),.doutb(w_n12445_0[1]),.din(n12445));
	jspl3 jspl3_w_n12447_0(.douta(w_n12447_0[0]),.doutb(w_n12447_0[1]),.doutc(w_n12447_0[2]),.din(n12447));
	jspl jspl_w_n12448_0(.douta(w_n12448_0[0]),.doutb(w_n12448_0[1]),.din(n12448));
	jspl jspl_w_n12452_0(.douta(w_n12452_0[0]),.doutb(w_n12452_0[1]),.din(n12452));
	jspl jspl_w_n12453_0(.douta(w_n12453_0[0]),.doutb(w_n12453_0[1]),.din(n12453));
	jspl3 jspl3_w_n12455_0(.douta(w_n12455_0[0]),.doutb(w_n12455_0[1]),.doutc(w_n12455_0[2]),.din(n12455));
	jspl jspl_w_n12456_0(.douta(w_n12456_0[0]),.doutb(w_n12456_0[1]),.din(n12456));
	jspl jspl_w_n12460_0(.douta(w_n12460_0[0]),.doutb(w_n12460_0[1]),.din(n12460));
	jspl3 jspl3_w_n12462_0(.douta(w_n12462_0[0]),.doutb(w_n12462_0[1]),.doutc(w_n12462_0[2]),.din(n12462));
	jspl jspl_w_n12463_0(.douta(w_n12463_0[0]),.doutb(w_n12463_0[1]),.din(n12463));
	jspl jspl_w_n12467_0(.douta(w_n12467_0[0]),.doutb(w_n12467_0[1]),.din(n12467));
	jspl jspl_w_n12468_0(.douta(w_n12468_0[0]),.doutb(w_n12468_0[1]),.din(n12468));
	jspl3 jspl3_w_n12470_0(.douta(w_n12470_0[0]),.doutb(w_n12470_0[1]),.doutc(w_n12470_0[2]),.din(n12470));
	jspl jspl_w_n12471_0(.douta(w_n12471_0[0]),.doutb(w_n12471_0[1]),.din(n12471));
	jspl jspl_w_n12475_0(.douta(w_n12475_0[0]),.doutb(w_n12475_0[1]),.din(n12475));
	jspl jspl_w_n12476_0(.douta(w_n12476_0[0]),.doutb(w_n12476_0[1]),.din(n12476));
	jspl3 jspl3_w_n12478_0(.douta(w_n12478_0[0]),.doutb(w_n12478_0[1]),.doutc(w_n12478_0[2]),.din(n12478));
	jspl jspl_w_n12479_0(.douta(w_n12479_0[0]),.doutb(w_n12479_0[1]),.din(n12479));
	jspl jspl_w_n12483_0(.douta(w_n12483_0[0]),.doutb(w_n12483_0[1]),.din(n12483));
	jspl jspl_w_n12484_0(.douta(w_n12484_0[0]),.doutb(w_n12484_0[1]),.din(n12484));
	jspl3 jspl3_w_n12486_0(.douta(w_n12486_0[0]),.doutb(w_n12486_0[1]),.doutc(w_n12486_0[2]),.din(n12486));
	jspl jspl_w_n12487_0(.douta(w_n12487_0[0]),.doutb(w_n12487_0[1]),.din(n12487));
	jspl jspl_w_n12491_0(.douta(w_n12491_0[0]),.doutb(w_n12491_0[1]),.din(n12491));
	jspl3 jspl3_w_n12493_0(.douta(w_n12493_0[0]),.doutb(w_n12493_0[1]),.doutc(w_n12493_0[2]),.din(n12493));
	jspl jspl_w_n12494_0(.douta(w_n12494_0[0]),.doutb(w_n12494_0[1]),.din(n12494));
	jspl jspl_w_n12498_0(.douta(w_n12498_0[0]),.doutb(w_n12498_0[1]),.din(n12498));
	jspl jspl_w_n12499_0(.douta(w_n12499_0[0]),.doutb(w_n12499_0[1]),.din(n12499));
	jspl3 jspl3_w_n12501_0(.douta(w_n12501_0[0]),.doutb(w_n12501_0[1]),.doutc(w_n12501_0[2]),.din(n12501));
	jspl jspl_w_n12502_0(.douta(w_n12502_0[0]),.doutb(w_n12502_0[1]),.din(n12502));
	jspl jspl_w_n12506_0(.douta(w_n12506_0[0]),.doutb(w_n12506_0[1]),.din(n12506));
	jspl3 jspl3_w_n12508_0(.douta(w_n12508_0[0]),.doutb(w_n12508_0[1]),.doutc(w_n12508_0[2]),.din(n12508));
	jspl jspl_w_n12509_0(.douta(w_n12509_0[0]),.doutb(w_n12509_0[1]),.din(n12509));
	jspl jspl_w_n12513_0(.douta(w_n12513_0[0]),.doutb(w_n12513_0[1]),.din(n12513));
	jspl jspl_w_n12514_0(.douta(w_n12514_0[0]),.doutb(w_n12514_0[1]),.din(n12514));
	jspl3 jspl3_w_n12516_0(.douta(w_n12516_0[0]),.doutb(w_n12516_0[1]),.doutc(w_n12516_0[2]),.din(n12516));
	jspl jspl_w_n12517_0(.douta(w_n12517_0[0]),.doutb(w_n12517_0[1]),.din(n12517));
	jspl jspl_w_n12521_0(.douta(w_n12521_0[0]),.doutb(w_n12521_0[1]),.din(n12521));
	jspl jspl_w_n12522_0(.douta(w_n12522_0[0]),.doutb(w_n12522_0[1]),.din(n12522));
	jspl3 jspl3_w_n12524_0(.douta(w_n12524_0[0]),.doutb(w_n12524_0[1]),.doutc(w_n12524_0[2]),.din(n12524));
	jspl jspl_w_n12525_0(.douta(w_n12525_0[0]),.doutb(w_n12525_0[1]),.din(n12525));
	jspl jspl_w_n12529_0(.douta(w_n12529_0[0]),.doutb(w_n12529_0[1]),.din(n12529));
	jspl jspl_w_n12530_0(.douta(w_n12530_0[0]),.doutb(w_n12530_0[1]),.din(n12530));
	jspl3 jspl3_w_n12532_0(.douta(w_n12532_0[0]),.doutb(w_n12532_0[1]),.doutc(w_n12532_0[2]),.din(n12532));
	jspl jspl_w_n12533_0(.douta(w_n12533_0[0]),.doutb(w_n12533_0[1]),.din(n12533));
	jspl jspl_w_n12537_0(.douta(w_n12537_0[0]),.doutb(w_n12537_0[1]),.din(n12537));
	jspl3 jspl3_w_n12539_0(.douta(w_n12539_0[0]),.doutb(w_n12539_0[1]),.doutc(w_n12539_0[2]),.din(n12539));
	jspl jspl_w_n12540_0(.douta(w_n12540_0[0]),.doutb(w_n12540_0[1]),.din(n12540));
	jspl jspl_w_n12544_0(.douta(w_n12544_0[0]),.doutb(w_n12544_0[1]),.din(n12544));
	jspl jspl_w_n12545_0(.douta(w_n12545_0[0]),.doutb(w_n12545_0[1]),.din(n12545));
	jspl3 jspl3_w_n12547_0(.douta(w_n12547_0[0]),.doutb(w_n12547_0[1]),.doutc(w_n12547_0[2]),.din(n12547));
	jspl jspl_w_n12548_0(.douta(w_n12548_0[0]),.doutb(w_n12548_0[1]),.din(n12548));
	jspl jspl_w_n12552_0(.douta(w_n12552_0[0]),.doutb(w_n12552_0[1]),.din(n12552));
	jspl jspl_w_n12553_0(.douta(w_n12553_0[0]),.doutb(w_n12553_0[1]),.din(n12553));
	jspl3 jspl3_w_n12555_0(.douta(w_n12555_0[0]),.doutb(w_n12555_0[1]),.doutc(w_n12555_0[2]),.din(n12555));
	jspl jspl_w_n12556_0(.douta(w_n12556_0[0]),.doutb(w_n12556_0[1]),.din(n12556));
	jspl jspl_w_n12560_0(.douta(w_n12560_0[0]),.doutb(w_n12560_0[1]),.din(n12560));
	jspl jspl_w_n12561_0(.douta(w_n12561_0[0]),.doutb(w_n12561_0[1]),.din(n12561));
	jspl3 jspl3_w_n12563_0(.douta(w_n12563_0[0]),.doutb(w_n12563_0[1]),.doutc(w_n12563_0[2]),.din(n12563));
	jspl jspl_w_n12564_0(.douta(w_n12564_0[0]),.doutb(w_n12564_0[1]),.din(n12564));
	jspl jspl_w_n12568_0(.douta(w_n12568_0[0]),.doutb(w_n12568_0[1]),.din(n12568));
	jspl jspl_w_n12569_0(.douta(w_n12569_0[0]),.doutb(w_n12569_0[1]),.din(n12569));
	jspl3 jspl3_w_n12571_0(.douta(w_n12571_0[0]),.doutb(w_n12571_0[1]),.doutc(w_n12571_0[2]),.din(n12571));
	jspl jspl_w_n12572_0(.douta(w_n12572_0[0]),.doutb(w_n12572_0[1]),.din(n12572));
	jspl3 jspl3_w_n12576_0(.douta(w_n12576_0[0]),.doutb(w_n12576_0[1]),.doutc(w_n12576_0[2]),.din(n12576));
	jspl3 jspl3_w_n12579_0(.douta(w_n12579_0[0]),.doutb(w_n12579_0[1]),.doutc(w_n12579_0[2]),.din(n12579));
	jspl jspl_w_n12580_0(.douta(w_n12580_0[0]),.doutb(w_n12580_0[1]),.din(n12580));
	jspl jspl_w_n12583_0(.douta(w_n12583_0[0]),.doutb(w_n12583_0[1]),.din(n12583));
	jspl3 jspl3_w_n12586_0(.douta(w_n12586_0[0]),.doutb(w_n12586_0[1]),.doutc(w_n12586_0[2]),.din(n12586));
	jspl jspl_w_n12587_0(.douta(w_n12587_0[0]),.doutb(w_n12587_0[1]),.din(n12587));
	jspl jspl_w_n12591_0(.douta(w_n12591_0[0]),.doutb(w_n12591_0[1]),.din(n12591));
	jspl jspl_w_n12592_0(.douta(w_n12592_0[0]),.doutb(w_n12592_0[1]),.din(n12592));
	jspl3 jspl3_w_n12594_0(.douta(w_n12594_0[0]),.doutb(w_n12594_0[1]),.doutc(w_n12594_0[2]),.din(n12594));
	jspl jspl_w_n12595_0(.douta(w_n12595_0[0]),.doutb(w_n12595_0[1]),.din(n12595));
	jspl jspl_w_n12599_0(.douta(w_n12599_0[0]),.doutb(w_n12599_0[1]),.din(n12599));
	jspl3 jspl3_w_n12601_0(.douta(w_n12601_0[0]),.doutb(w_n12601_0[1]),.doutc(w_n12601_0[2]),.din(n12601));
	jspl jspl_w_n12602_0(.douta(w_n12602_0[0]),.doutb(w_n12602_0[1]),.din(n12602));
	jspl jspl_w_n12606_0(.douta(w_n12606_0[0]),.doutb(w_n12606_0[1]),.din(n12606));
	jspl jspl_w_n12607_0(.douta(w_n12607_0[0]),.doutb(w_n12607_0[1]),.din(n12607));
	jspl3 jspl3_w_n12609_0(.douta(w_n12609_0[0]),.doutb(w_n12609_0[1]),.doutc(w_n12609_0[2]),.din(n12609));
	jspl jspl_w_n12610_0(.douta(w_n12610_0[0]),.doutb(w_n12610_0[1]),.din(n12610));
	jspl jspl_w_n12614_0(.douta(w_n12614_0[0]),.doutb(w_n12614_0[1]),.din(n12614));
	jspl3 jspl3_w_n12616_0(.douta(w_n12616_0[0]),.doutb(w_n12616_0[1]),.doutc(w_n12616_0[2]),.din(n12616));
	jspl jspl_w_n12617_0(.douta(w_n12617_0[0]),.doutb(w_n12617_0[1]),.din(n12617));
	jspl jspl_w_n12621_0(.douta(w_n12621_0[0]),.doutb(w_n12621_0[1]),.din(n12621));
	jspl jspl_w_n12622_0(.douta(w_n12622_0[0]),.doutb(w_n12622_0[1]),.din(n12622));
	jspl3 jspl3_w_n12624_0(.douta(w_n12624_0[0]),.doutb(w_n12624_0[1]),.doutc(w_n12624_0[2]),.din(n12624));
	jspl jspl_w_n12625_0(.douta(w_n12625_0[0]),.doutb(w_n12625_0[1]),.din(n12625));
	jspl jspl_w_n12629_0(.douta(w_n12629_0[0]),.doutb(w_n12629_0[1]),.din(n12629));
	jspl jspl_w_n12630_0(.douta(w_n12630_0[0]),.doutb(w_n12630_0[1]),.din(n12630));
	jspl3 jspl3_w_n12632_0(.douta(w_n12632_0[0]),.doutb(w_n12632_0[1]),.doutc(w_n12632_0[2]),.din(n12632));
	jspl jspl_w_n12633_0(.douta(w_n12633_0[0]),.doutb(w_n12633_0[1]),.din(n12633));
	jspl jspl_w_n12637_0(.douta(w_n12637_0[0]),.doutb(w_n12637_0[1]),.din(n12637));
	jspl jspl_w_n12638_0(.douta(w_n12638_0[0]),.doutb(w_n12638_0[1]),.din(n12638));
	jspl3 jspl3_w_n12640_0(.douta(w_n12640_0[0]),.doutb(w_n12640_0[1]),.doutc(w_n12640_0[2]),.din(n12640));
	jspl jspl_w_n12641_0(.douta(w_n12641_0[0]),.doutb(w_n12641_0[1]),.din(n12641));
	jspl jspl_w_n12645_0(.douta(w_n12645_0[0]),.doutb(w_n12645_0[1]),.din(n12645));
	jspl3 jspl3_w_n12647_0(.douta(w_n12647_0[0]),.doutb(w_n12647_0[1]),.doutc(w_n12647_0[2]),.din(n12647));
	jspl jspl_w_n12648_0(.douta(w_n12648_0[0]),.doutb(w_n12648_0[1]),.din(n12648));
	jspl jspl_w_n12652_0(.douta(w_n12652_0[0]),.doutb(w_n12652_0[1]),.din(n12652));
	jspl jspl_w_n12653_0(.douta(w_n12653_0[0]),.doutb(w_n12653_0[1]),.din(n12653));
	jspl3 jspl3_w_n12655_0(.douta(w_n12655_0[0]),.doutb(w_n12655_0[1]),.doutc(w_n12655_0[2]),.din(n12655));
	jspl jspl_w_n12656_0(.douta(w_n12656_0[0]),.doutb(w_n12656_0[1]),.din(n12656));
	jspl jspl_w_n12660_0(.douta(w_n12660_0[0]),.doutb(w_n12660_0[1]),.din(n12660));
	jspl3 jspl3_w_n12662_0(.douta(w_n12662_0[0]),.doutb(w_n12662_0[1]),.doutc(w_n12662_0[2]),.din(n12662));
	jspl jspl_w_n12663_0(.douta(w_n12663_0[0]),.doutb(w_n12663_0[1]),.din(n12663));
	jspl jspl_w_n12667_0(.douta(w_n12667_0[0]),.doutb(w_n12667_0[1]),.din(n12667));
	jspl jspl_w_n12668_0(.douta(w_n12668_0[0]),.doutb(w_n12668_0[1]),.din(n12668));
	jspl3 jspl3_w_n12670_0(.douta(w_n12670_0[0]),.doutb(w_n12670_0[1]),.doutc(w_n12670_0[2]),.din(n12670));
	jspl jspl_w_n12671_0(.douta(w_n12671_0[0]),.doutb(w_n12671_0[1]),.din(n12671));
	jspl jspl_w_n12675_0(.douta(w_n12675_0[0]),.doutb(w_n12675_0[1]),.din(n12675));
	jspl3 jspl3_w_n12677_0(.douta(w_n12677_0[0]),.doutb(w_n12677_0[1]),.doutc(w_n12677_0[2]),.din(n12677));
	jspl jspl_w_n12678_0(.douta(w_n12678_0[0]),.doutb(w_n12678_0[1]),.din(n12678));
	jspl jspl_w_n12682_0(.douta(w_n12682_0[0]),.doutb(w_n12682_0[1]),.din(n12682));
	jspl jspl_w_n12683_0(.douta(w_n12683_0[0]),.doutb(w_n12683_0[1]),.din(n12683));
	jspl3 jspl3_w_n12685_0(.douta(w_n12685_0[0]),.doutb(w_n12685_0[1]),.doutc(w_n12685_0[2]),.din(n12685));
	jspl jspl_w_n12686_0(.douta(w_n12686_0[0]),.doutb(w_n12686_0[1]),.din(n12686));
	jspl jspl_w_n12690_0(.douta(w_n12690_0[0]),.doutb(w_n12690_0[1]),.din(n12690));
	jspl3 jspl3_w_n12692_0(.douta(w_n12692_0[0]),.doutb(w_n12692_0[1]),.doutc(w_n12692_0[2]),.din(n12692));
	jspl jspl_w_n12693_0(.douta(w_n12693_0[0]),.doutb(w_n12693_0[1]),.din(n12693));
	jspl jspl_w_n12697_0(.douta(w_n12697_0[0]),.doutb(w_n12697_0[1]),.din(n12697));
	jspl3 jspl3_w_n12699_0(.douta(w_n12699_0[0]),.doutb(w_n12699_0[1]),.doutc(w_n12699_0[2]),.din(n12699));
	jspl jspl_w_n12700_0(.douta(w_n12700_0[0]),.doutb(w_n12700_0[1]),.din(n12700));
	jspl jspl_w_n12704_0(.douta(w_n12704_0[0]),.doutb(w_n12704_0[1]),.din(n12704));
	jspl3 jspl3_w_n12706_0(.douta(w_n12706_0[0]),.doutb(w_n12706_0[1]),.doutc(w_n12706_0[2]),.din(n12706));
	jspl jspl_w_n12707_0(.douta(w_n12707_0[0]),.doutb(w_n12707_0[1]),.din(n12707));
	jspl jspl_w_n12711_0(.douta(w_n12711_0[0]),.doutb(w_n12711_0[1]),.din(n12711));
	jspl jspl_w_n12712_0(.douta(w_n12712_0[0]),.doutb(w_n12712_0[1]),.din(n12712));
	jspl3 jspl3_w_n12714_0(.douta(w_n12714_0[0]),.doutb(w_n12714_0[1]),.doutc(w_n12714_0[2]),.din(n12714));
	jspl jspl_w_n12715_0(.douta(w_n12715_0[0]),.doutb(w_n12715_0[1]),.din(n12715));
	jspl jspl_w_n12719_0(.douta(w_n12719_0[0]),.doutb(w_n12719_0[1]),.din(n12719));
	jspl jspl_w_n12720_0(.douta(w_n12720_0[0]),.doutb(w_n12720_0[1]),.din(n12720));
	jspl3 jspl3_w_n12722_0(.douta(w_n12722_0[0]),.doutb(w_n12722_0[1]),.doutc(w_n12722_0[2]),.din(n12722));
	jspl jspl_w_n12723_0(.douta(w_n12723_0[0]),.doutb(w_n12723_0[1]),.din(n12723));
	jspl3 jspl3_w_n12727_0(.douta(w_n12727_0[0]),.doutb(w_n12727_0[1]),.doutc(w_n12727_0[2]),.din(n12727));
	jspl jspl_w_n12730_0(.douta(w_n12730_0[0]),.doutb(w_n12730_0[1]),.din(n12730));
	jspl3 jspl3_w_n12731_0(.douta(w_n12731_0[0]),.doutb(w_n12731_0[1]),.doutc(w_n12731_0[2]),.din(n12731));
	jspl jspl_w_n12731_1(.douta(w_n12731_1[0]),.doutb(w_n12731_1[1]),.din(w_n12731_0[0]));
	jspl3 jspl3_w_n12732_0(.douta(w_n12732_0[0]),.doutb(w_n12732_0[1]),.doutc(w_n12732_0[2]),.din(n12732));
	jspl jspl_w_n12736_0(.douta(w_n12736_0[0]),.doutb(w_n12736_0[1]),.din(n12736));
	jspl jspl_w_n12737_0(.douta(w_n12737_0[0]),.doutb(w_n12737_0[1]),.din(n12737));
	jspl jspl_w_n12738_0(.douta(w_n12738_0[0]),.doutb(w_n12738_0[1]),.din(n12738));
	jspl jspl_w_n12739_0(.douta(w_n12739_0[0]),.doutb(w_n12739_0[1]),.din(n12739));
	jspl jspl_w_n12760_0(.douta(w_n12760_0[0]),.doutb(w_n12760_0[1]),.din(n12760));
	jspl jspl_w_n12789_0(.douta(w_n12789_0[0]),.doutb(w_n12789_0[1]),.din(n12789));
	jspl jspl_w_n12796_0(.douta(w_n12796_0[0]),.doutb(w_n12796_0[1]),.din(n12796));
	jspl jspl_w_n12803_0(.douta(w_n12803_0[0]),.doutb(w_n12803_0[1]),.din(n12803));
	jspl jspl_w_n12810_0(.douta(w_n12810_0[0]),.doutb(w_n12810_0[1]),.din(n12810));
	jspl jspl_w_n12823_0(.douta(w_n12823_0[0]),.doutb(w_n12823_0[1]),.din(n12823));
	jspl jspl_w_n12830_0(.douta(w_n12830_0[0]),.doutb(w_n12830_0[1]),.din(n12830));
	jspl jspl_w_n12843_0(.douta(w_n12843_0[0]),.doutb(w_n12843_0[1]),.din(n12843));
	jspl jspl_w_n12868_0(.douta(w_n12868_0[0]),.doutb(w_n12868_0[1]),.din(n12868));
	jspl jspl_w_n12875_0(.douta(w_n12875_0[0]),.doutb(w_n12875_0[1]),.din(n12875));
	jspl jspl_w_n12888_0(.douta(w_n12888_0[0]),.doutb(w_n12888_0[1]),.din(n12888));
	jspl jspl_w_n12895_0(.douta(w_n12895_0[0]),.doutb(w_n12895_0[1]),.din(n12895));
	jspl jspl_w_n12902_0(.douta(w_n12902_0[0]),.doutb(w_n12902_0[1]),.din(n12902));
	jspl jspl_w_n12909_0(.douta(w_n12909_0[0]),.doutb(w_n12909_0[1]),.din(n12909));
	jspl jspl_w_n12913_0(.douta(w_n12913_0[0]),.doutb(w_n12913_0[1]),.din(n12913));
	jspl jspl_w_n12917_0(.douta(w_n12917_0[0]),.doutb(w_n12917_0[1]),.din(n12917));
	jspl jspl_w_n12928_0(.douta(w_n12928_0[0]),.doutb(w_n12928_0[1]),.din(n12928));
	jspl jspl_w_n12929_0(.douta(w_n12929_0[0]),.doutb(w_n12929_0[1]),.din(n12929));
	jspl jspl_w_n12932_0(.douta(w_n12932_0[0]),.doutb(w_n12932_0[1]),.din(n12932));
	jspl jspl_w_n12933_0(.douta(w_n12933_0[0]),.doutb(w_n12933_0[1]),.din(n12933));
	jspl jspl_w_n12935_0(.douta(w_n12935_0[0]),.doutb(w_n12935_0[1]),.din(n12935));
	jspl jspl_w_n12937_0(.douta(w_n12937_0[0]),.doutb(w_n12937_0[1]),.din(n12937));
	jspl jspl_w_n12938_0(.douta(w_n12938_0[0]),.doutb(w_n12938_0[1]),.din(n12938));
	jspl jspl_w_n12946_0(.douta(w_n12946_0[0]),.doutb(w_n12946_0[1]),.din(n12946));
	jspl3 jspl3_w_n12947_0(.douta(w_n12947_0[0]),.doutb(w_n12947_0[1]),.doutc(w_n12947_0[2]),.din(n12947));
	jspl3 jspl3_w_n12947_1(.douta(w_n12947_1[0]),.doutb(w_n12947_1[1]),.doutc(w_n12947_1[2]),.din(w_n12947_0[0]));
	jspl3 jspl3_w_n12947_2(.douta(w_n12947_2[0]),.doutb(w_n12947_2[1]),.doutc(w_n12947_2[2]),.din(w_n12947_0[1]));
	jspl3 jspl3_w_n12947_3(.douta(w_n12947_3[0]),.doutb(w_n12947_3[1]),.doutc(w_n12947_3[2]),.din(w_n12947_0[2]));
	jspl3 jspl3_w_n12947_4(.douta(w_n12947_4[0]),.doutb(w_n12947_4[1]),.doutc(w_n12947_4[2]),.din(w_n12947_1[0]));
	jspl3 jspl3_w_n12947_5(.douta(w_n12947_5[0]),.doutb(w_n12947_5[1]),.doutc(w_n12947_5[2]),.din(w_n12947_1[1]));
	jspl3 jspl3_w_n12947_6(.douta(w_n12947_6[0]),.doutb(w_n12947_6[1]),.doutc(w_n12947_6[2]),.din(w_n12947_1[2]));
	jspl3 jspl3_w_n12947_7(.douta(w_n12947_7[0]),.doutb(w_n12947_7[1]),.doutc(w_n12947_7[2]),.din(w_n12947_2[0]));
	jspl3 jspl3_w_n12947_8(.douta(w_n12947_8[0]),.doutb(w_n12947_8[1]),.doutc(w_n12947_8[2]),.din(w_n12947_2[1]));
	jspl3 jspl3_w_n12947_9(.douta(w_n12947_9[0]),.doutb(w_n12947_9[1]),.doutc(w_n12947_9[2]),.din(w_n12947_2[2]));
	jspl3 jspl3_w_n12947_10(.douta(w_n12947_10[0]),.doutb(w_n12947_10[1]),.doutc(w_n12947_10[2]),.din(w_n12947_3[0]));
	jspl3 jspl3_w_n12947_11(.douta(w_n12947_11[0]),.doutb(w_n12947_11[1]),.doutc(w_n12947_11[2]),.din(w_n12947_3[1]));
	jspl3 jspl3_w_n12947_12(.douta(w_n12947_12[0]),.doutb(w_n12947_12[1]),.doutc(w_n12947_12[2]),.din(w_n12947_3[2]));
	jspl3 jspl3_w_n12947_13(.douta(w_n12947_13[0]),.doutb(w_n12947_13[1]),.doutc(w_n12947_13[2]),.din(w_n12947_4[0]));
	jspl3 jspl3_w_n12947_14(.douta(w_n12947_14[0]),.doutb(w_n12947_14[1]),.doutc(w_n12947_14[2]),.din(w_n12947_4[1]));
	jspl3 jspl3_w_n12947_15(.douta(w_n12947_15[0]),.doutb(w_n12947_15[1]),.doutc(w_n12947_15[2]),.din(w_n12947_4[2]));
	jspl3 jspl3_w_n12947_16(.douta(w_n12947_16[0]),.doutb(w_n12947_16[1]),.doutc(w_n12947_16[2]),.din(w_n12947_5[0]));
	jspl3 jspl3_w_n12947_17(.douta(w_n12947_17[0]),.doutb(w_n12947_17[1]),.doutc(w_n12947_17[2]),.din(w_n12947_5[1]));
	jspl3 jspl3_w_n12947_18(.douta(w_n12947_18[0]),.doutb(w_n12947_18[1]),.doutc(w_n12947_18[2]),.din(w_n12947_5[2]));
	jspl3 jspl3_w_n12947_19(.douta(w_n12947_19[0]),.doutb(w_n12947_19[1]),.doutc(w_n12947_19[2]),.din(w_n12947_6[0]));
	jspl3 jspl3_w_n12947_20(.douta(w_n12947_20[0]),.doutb(w_n12947_20[1]),.doutc(w_n12947_20[2]),.din(w_n12947_6[1]));
	jspl3 jspl3_w_n12947_21(.douta(w_n12947_21[0]),.doutb(w_n12947_21[1]),.doutc(w_n12947_21[2]),.din(w_n12947_6[2]));
	jspl3 jspl3_w_n12947_22(.douta(w_n12947_22[0]),.doutb(w_n12947_22[1]),.doutc(w_n12947_22[2]),.din(w_n12947_7[0]));
	jspl3 jspl3_w_n12947_23(.douta(w_n12947_23[0]),.doutb(w_n12947_23[1]),.doutc(w_n12947_23[2]),.din(w_n12947_7[1]));
	jspl3 jspl3_w_n12947_24(.douta(w_n12947_24[0]),.doutb(w_n12947_24[1]),.doutc(w_n12947_24[2]),.din(w_n12947_7[2]));
	jspl3 jspl3_w_n12947_25(.douta(w_n12947_25[0]),.doutb(w_n12947_25[1]),.doutc(w_n12947_25[2]),.din(w_n12947_8[0]));
	jspl3 jspl3_w_n12947_26(.douta(w_n12947_26[0]),.doutb(w_n12947_26[1]),.doutc(w_n12947_26[2]),.din(w_n12947_8[1]));
	jspl3 jspl3_w_n12947_27(.douta(w_n12947_27[0]),.doutb(w_n12947_27[1]),.doutc(w_n12947_27[2]),.din(w_n12947_8[2]));
	jspl3 jspl3_w_n12947_28(.douta(w_n12947_28[0]),.doutb(w_n12947_28[1]),.doutc(w_n12947_28[2]),.din(w_n12947_9[0]));
	jspl3 jspl3_w_n12947_29(.douta(w_n12947_29[0]),.doutb(w_n12947_29[1]),.doutc(w_n12947_29[2]),.din(w_n12947_9[1]));
	jspl3 jspl3_w_n12947_30(.douta(w_n12947_30[0]),.doutb(w_n12947_30[1]),.doutc(w_n12947_30[2]),.din(w_n12947_9[2]));
	jspl3 jspl3_w_n12947_31(.douta(w_n12947_31[0]),.doutb(w_n12947_31[1]),.doutc(w_n12947_31[2]),.din(w_n12947_10[0]));
	jspl3 jspl3_w_n12947_32(.douta(w_n12947_32[0]),.doutb(w_n12947_32[1]),.doutc(w_n12947_32[2]),.din(w_n12947_10[1]));
	jspl3 jspl3_w_n12947_33(.douta(w_n12947_33[0]),.doutb(w_n12947_33[1]),.doutc(w_n12947_33[2]),.din(w_n12947_10[2]));
	jspl3 jspl3_w_n12947_34(.douta(w_n12947_34[0]),.doutb(w_n12947_34[1]),.doutc(w_n12947_34[2]),.din(w_n12947_11[0]));
	jspl3 jspl3_w_n12947_35(.douta(w_n12947_35[0]),.doutb(w_n12947_35[1]),.doutc(w_n12947_35[2]),.din(w_n12947_11[1]));
	jspl3 jspl3_w_n12947_36(.douta(w_n12947_36[0]),.doutb(w_n12947_36[1]),.doutc(w_n12947_36[2]),.din(w_n12947_11[2]));
	jspl3 jspl3_w_n12947_37(.douta(w_n12947_37[0]),.doutb(w_n12947_37[1]),.doutc(w_n12947_37[2]),.din(w_n12947_12[0]));
	jspl3 jspl3_w_n12947_38(.douta(w_n12947_38[0]),.doutb(w_n12947_38[1]),.doutc(w_n12947_38[2]),.din(w_n12947_12[1]));
	jspl3 jspl3_w_n12947_39(.douta(w_n12947_39[0]),.doutb(w_n12947_39[1]),.doutc(w_n12947_39[2]),.din(w_n12947_12[2]));
	jspl3 jspl3_w_n12947_40(.douta(w_n12947_40[0]),.doutb(w_n12947_40[1]),.doutc(w_n12947_40[2]),.din(w_n12947_13[0]));
	jspl3 jspl3_w_n12947_41(.douta(w_n12947_41[0]),.doutb(w_n12947_41[1]),.doutc(w_n12947_41[2]),.din(w_n12947_13[1]));
	jspl3 jspl3_w_n12947_42(.douta(w_n12947_42[0]),.doutb(w_n12947_42[1]),.doutc(w_n12947_42[2]),.din(w_n12947_13[2]));
	jspl3 jspl3_w_n12947_43(.douta(w_n12947_43[0]),.doutb(w_n12947_43[1]),.doutc(w_n12947_43[2]),.din(w_n12947_14[0]));
	jspl3 jspl3_w_n12947_44(.douta(w_n12947_44[0]),.doutb(w_n12947_44[1]),.doutc(w_n12947_44[2]),.din(w_n12947_14[1]));
	jspl jspl_w_n12950_0(.douta(w_n12950_0[0]),.doutb(w_n12950_0[1]),.din(n12950));
	jspl3 jspl3_w_n12951_0(.douta(w_n12951_0[0]),.doutb(w_n12951_0[1]),.doutc(w_n12951_0[2]),.din(n12951));
	jspl3 jspl3_w_n12953_0(.douta(w_n12953_0[0]),.doutb(w_n12953_0[1]),.doutc(w_n12953_0[2]),.din(n12953));
	jspl3 jspl3_w_n12953_1(.douta(w_n12953_1[0]),.doutb(w_n12953_1[1]),.doutc(w_n12953_1[2]),.din(w_n12953_0[0]));
	jspl jspl_w_n12954_0(.douta(w_n12954_0[0]),.doutb(w_n12954_0[1]),.din(n12954));
	jspl3 jspl3_w_n12955_0(.douta(w_n12955_0[0]),.doutb(w_n12955_0[1]),.doutc(w_n12955_0[2]),.din(n12955));
	jspl jspl_w_n12956_0(.douta(w_n12956_0[0]),.doutb(w_n12956_0[1]),.din(n12956));
	jspl3 jspl3_w_n12958_0(.douta(w_n12958_0[0]),.doutb(w_n12958_0[1]),.doutc(w_n12958_0[2]),.din(n12958));
	jspl jspl_w_n12959_0(.douta(w_n12959_0[0]),.doutb(w_n12959_0[1]),.din(n12959));
	jspl jspl_w_n12964_0(.douta(w_n12964_0[0]),.doutb(w_n12964_0[1]),.din(n12964));
	jspl3 jspl3_w_n12966_0(.douta(w_n12966_0[0]),.doutb(w_n12966_0[1]),.doutc(w_n12966_0[2]),.din(n12966));
	jspl jspl_w_n12967_0(.douta(w_n12967_0[0]),.doutb(w_n12967_0[1]),.din(n12967));
	jspl jspl_w_n12970_0(.douta(w_n12970_0[0]),.doutb(w_n12970_0[1]),.din(n12970));
	jspl3 jspl3_w_n12975_0(.douta(w_n12975_0[0]),.doutb(w_n12975_0[1]),.doutc(w_n12975_0[2]),.din(n12975));
	jspl3 jspl3_w_n12977_0(.douta(w_n12977_0[0]),.doutb(w_n12977_0[1]),.doutc(w_n12977_0[2]),.din(n12977));
	jspl jspl_w_n12978_0(.douta(w_n12978_0[0]),.doutb(w_n12978_0[1]),.din(n12978));
	jspl3 jspl3_w_n12982_0(.douta(w_n12982_0[0]),.doutb(w_n12982_0[1]),.doutc(w_n12982_0[2]),.din(n12982));
	jspl3 jspl3_w_n12985_0(.douta(w_n12985_0[0]),.doutb(w_n12985_0[1]),.doutc(w_n12985_0[2]),.din(n12985));
	jspl jspl_w_n12986_0(.douta(w_n12986_0[0]),.doutb(w_n12986_0[1]),.din(n12986));
	jspl3 jspl3_w_n12990_0(.douta(w_n12990_0[0]),.doutb(w_n12990_0[1]),.doutc(w_n12990_0[2]),.din(n12990));
	jspl3 jspl3_w_n12992_0(.douta(w_n12992_0[0]),.doutb(w_n12992_0[1]),.doutc(w_n12992_0[2]),.din(n12992));
	jspl jspl_w_n12993_0(.douta(w_n12993_0[0]),.doutb(w_n12993_0[1]),.din(n12993));
	jspl3 jspl3_w_n12997_0(.douta(w_n12997_0[0]),.doutb(w_n12997_0[1]),.doutc(w_n12997_0[2]),.din(n12997));
	jspl3 jspl3_w_n13000_0(.douta(w_n13000_0[0]),.doutb(w_n13000_0[1]),.doutc(w_n13000_0[2]),.din(n13000));
	jspl jspl_w_n13001_0(.douta(w_n13001_0[0]),.doutb(w_n13001_0[1]),.din(n13001));
	jspl3 jspl3_w_n13005_0(.douta(w_n13005_0[0]),.doutb(w_n13005_0[1]),.doutc(w_n13005_0[2]),.din(n13005));
	jspl3 jspl3_w_n13007_0(.douta(w_n13007_0[0]),.doutb(w_n13007_0[1]),.doutc(w_n13007_0[2]),.din(n13007));
	jspl jspl_w_n13008_0(.douta(w_n13008_0[0]),.doutb(w_n13008_0[1]),.din(n13008));
	jspl3 jspl3_w_n13012_0(.douta(w_n13012_0[0]),.doutb(w_n13012_0[1]),.doutc(w_n13012_0[2]),.din(n13012));
	jspl3 jspl3_w_n13015_0(.douta(w_n13015_0[0]),.doutb(w_n13015_0[1]),.doutc(w_n13015_0[2]),.din(n13015));
	jspl jspl_w_n13016_0(.douta(w_n13016_0[0]),.doutb(w_n13016_0[1]),.din(n13016));
	jspl3 jspl3_w_n13020_0(.douta(w_n13020_0[0]),.doutb(w_n13020_0[1]),.doutc(w_n13020_0[2]),.din(n13020));
	jspl3 jspl3_w_n13022_0(.douta(w_n13022_0[0]),.doutb(w_n13022_0[1]),.doutc(w_n13022_0[2]),.din(n13022));
	jspl jspl_w_n13023_0(.douta(w_n13023_0[0]),.doutb(w_n13023_0[1]),.din(n13023));
	jspl3 jspl3_w_n13027_0(.douta(w_n13027_0[0]),.doutb(w_n13027_0[1]),.doutc(w_n13027_0[2]),.din(n13027));
	jspl3 jspl3_w_n13030_0(.douta(w_n13030_0[0]),.doutb(w_n13030_0[1]),.doutc(w_n13030_0[2]),.din(n13030));
	jspl jspl_w_n13031_0(.douta(w_n13031_0[0]),.doutb(w_n13031_0[1]),.din(n13031));
	jspl3 jspl3_w_n13035_0(.douta(w_n13035_0[0]),.doutb(w_n13035_0[1]),.doutc(w_n13035_0[2]),.din(n13035));
	jspl3 jspl3_w_n13037_0(.douta(w_n13037_0[0]),.doutb(w_n13037_0[1]),.doutc(w_n13037_0[2]),.din(n13037));
	jspl jspl_w_n13038_0(.douta(w_n13038_0[0]),.doutb(w_n13038_0[1]),.din(n13038));
	jspl3 jspl3_w_n13042_0(.douta(w_n13042_0[0]),.doutb(w_n13042_0[1]),.doutc(w_n13042_0[2]),.din(n13042));
	jspl3 jspl3_w_n13044_0(.douta(w_n13044_0[0]),.doutb(w_n13044_0[1]),.doutc(w_n13044_0[2]),.din(n13044));
	jspl jspl_w_n13045_0(.douta(w_n13045_0[0]),.doutb(w_n13045_0[1]),.din(n13045));
	jspl3 jspl3_w_n13049_0(.douta(w_n13049_0[0]),.doutb(w_n13049_0[1]),.doutc(w_n13049_0[2]),.din(n13049));
	jspl3 jspl3_w_n13051_0(.douta(w_n13051_0[0]),.doutb(w_n13051_0[1]),.doutc(w_n13051_0[2]),.din(n13051));
	jspl jspl_w_n13052_0(.douta(w_n13052_0[0]),.doutb(w_n13052_0[1]),.din(n13052));
	jspl3 jspl3_w_n13056_0(.douta(w_n13056_0[0]),.doutb(w_n13056_0[1]),.doutc(w_n13056_0[2]),.din(n13056));
	jspl3 jspl3_w_n13059_0(.douta(w_n13059_0[0]),.doutb(w_n13059_0[1]),.doutc(w_n13059_0[2]),.din(n13059));
	jspl jspl_w_n13060_0(.douta(w_n13060_0[0]),.doutb(w_n13060_0[1]),.din(n13060));
	jspl3 jspl3_w_n13064_0(.douta(w_n13064_0[0]),.doutb(w_n13064_0[1]),.doutc(w_n13064_0[2]),.din(n13064));
	jspl3 jspl3_w_n13066_0(.douta(w_n13066_0[0]),.doutb(w_n13066_0[1]),.doutc(w_n13066_0[2]),.din(n13066));
	jspl jspl_w_n13067_0(.douta(w_n13067_0[0]),.doutb(w_n13067_0[1]),.din(n13067));
	jspl3 jspl3_w_n13071_0(.douta(w_n13071_0[0]),.doutb(w_n13071_0[1]),.doutc(w_n13071_0[2]),.din(n13071));
	jspl3 jspl3_w_n13074_0(.douta(w_n13074_0[0]),.doutb(w_n13074_0[1]),.doutc(w_n13074_0[2]),.din(n13074));
	jspl jspl_w_n13075_0(.douta(w_n13075_0[0]),.doutb(w_n13075_0[1]),.din(n13075));
	jspl3 jspl3_w_n13079_0(.douta(w_n13079_0[0]),.doutb(w_n13079_0[1]),.doutc(w_n13079_0[2]),.din(n13079));
	jspl3 jspl3_w_n13081_0(.douta(w_n13081_0[0]),.doutb(w_n13081_0[1]),.doutc(w_n13081_0[2]),.din(n13081));
	jspl jspl_w_n13082_0(.douta(w_n13082_0[0]),.doutb(w_n13082_0[1]),.din(n13082));
	jspl3 jspl3_w_n13086_0(.douta(w_n13086_0[0]),.doutb(w_n13086_0[1]),.doutc(w_n13086_0[2]),.din(n13086));
	jspl3 jspl3_w_n13088_0(.douta(w_n13088_0[0]),.doutb(w_n13088_0[1]),.doutc(w_n13088_0[2]),.din(n13088));
	jspl jspl_w_n13089_0(.douta(w_n13089_0[0]),.doutb(w_n13089_0[1]),.din(n13089));
	jspl3 jspl3_w_n13093_0(.douta(w_n13093_0[0]),.doutb(w_n13093_0[1]),.doutc(w_n13093_0[2]),.din(n13093));
	jspl3 jspl3_w_n13095_0(.douta(w_n13095_0[0]),.doutb(w_n13095_0[1]),.doutc(w_n13095_0[2]),.din(n13095));
	jspl jspl_w_n13096_0(.douta(w_n13096_0[0]),.doutb(w_n13096_0[1]),.din(n13096));
	jspl3 jspl3_w_n13100_0(.douta(w_n13100_0[0]),.doutb(w_n13100_0[1]),.doutc(w_n13100_0[2]),.din(n13100));
	jspl3 jspl3_w_n13103_0(.douta(w_n13103_0[0]),.doutb(w_n13103_0[1]),.doutc(w_n13103_0[2]),.din(n13103));
	jspl jspl_w_n13104_0(.douta(w_n13104_0[0]),.doutb(w_n13104_0[1]),.din(n13104));
	jspl3 jspl3_w_n13108_0(.douta(w_n13108_0[0]),.doutb(w_n13108_0[1]),.doutc(w_n13108_0[2]),.din(n13108));
	jspl3 jspl3_w_n13110_0(.douta(w_n13110_0[0]),.doutb(w_n13110_0[1]),.doutc(w_n13110_0[2]),.din(n13110));
	jspl jspl_w_n13111_0(.douta(w_n13111_0[0]),.doutb(w_n13111_0[1]),.din(n13111));
	jspl3 jspl3_w_n13115_0(.douta(w_n13115_0[0]),.doutb(w_n13115_0[1]),.doutc(w_n13115_0[2]),.din(n13115));
	jspl3 jspl3_w_n13117_0(.douta(w_n13117_0[0]),.doutb(w_n13117_0[1]),.doutc(w_n13117_0[2]),.din(n13117));
	jspl jspl_w_n13118_0(.douta(w_n13118_0[0]),.doutb(w_n13118_0[1]),.din(n13118));
	jspl3 jspl3_w_n13122_0(.douta(w_n13122_0[0]),.doutb(w_n13122_0[1]),.doutc(w_n13122_0[2]),.din(n13122));
	jspl3 jspl3_w_n13124_0(.douta(w_n13124_0[0]),.doutb(w_n13124_0[1]),.doutc(w_n13124_0[2]),.din(n13124));
	jspl jspl_w_n13125_0(.douta(w_n13125_0[0]),.doutb(w_n13125_0[1]),.din(n13125));
	jspl3 jspl3_w_n13129_0(.douta(w_n13129_0[0]),.doutb(w_n13129_0[1]),.doutc(w_n13129_0[2]),.din(n13129));
	jspl3 jspl3_w_n13131_0(.douta(w_n13131_0[0]),.doutb(w_n13131_0[1]),.doutc(w_n13131_0[2]),.din(n13131));
	jspl jspl_w_n13132_0(.douta(w_n13132_0[0]),.doutb(w_n13132_0[1]),.din(n13132));
	jspl3 jspl3_w_n13136_0(.douta(w_n13136_0[0]),.doutb(w_n13136_0[1]),.doutc(w_n13136_0[2]),.din(n13136));
	jspl3 jspl3_w_n13139_0(.douta(w_n13139_0[0]),.doutb(w_n13139_0[1]),.doutc(w_n13139_0[2]),.din(n13139));
	jspl jspl_w_n13140_0(.douta(w_n13140_0[0]),.doutb(w_n13140_0[1]),.din(n13140));
	jspl3 jspl3_w_n13143_0(.douta(w_n13143_0[0]),.doutb(w_n13143_0[1]),.doutc(w_n13143_0[2]),.din(n13143));
	jspl3 jspl3_w_n13147_0(.douta(w_n13147_0[0]),.doutb(w_n13147_0[1]),.doutc(w_n13147_0[2]),.din(n13147));
	jspl jspl_w_n13148_0(.douta(w_n13148_0[0]),.doutb(w_n13148_0[1]),.din(n13148));
	jspl3 jspl3_w_n13152_0(.douta(w_n13152_0[0]),.doutb(w_n13152_0[1]),.doutc(w_n13152_0[2]),.din(n13152));
	jspl3 jspl3_w_n13154_0(.douta(w_n13154_0[0]),.doutb(w_n13154_0[1]),.doutc(w_n13154_0[2]),.din(n13154));
	jspl jspl_w_n13155_0(.douta(w_n13155_0[0]),.doutb(w_n13155_0[1]),.din(n13155));
	jspl3 jspl3_w_n13159_0(.douta(w_n13159_0[0]),.doutb(w_n13159_0[1]),.doutc(w_n13159_0[2]),.din(n13159));
	jspl3 jspl3_w_n13162_0(.douta(w_n13162_0[0]),.doutb(w_n13162_0[1]),.doutc(w_n13162_0[2]),.din(n13162));
	jspl jspl_w_n13163_0(.douta(w_n13163_0[0]),.doutb(w_n13163_0[1]),.din(n13163));
	jspl3 jspl3_w_n13167_0(.douta(w_n13167_0[0]),.doutb(w_n13167_0[1]),.doutc(w_n13167_0[2]),.din(n13167));
	jspl3 jspl3_w_n13169_0(.douta(w_n13169_0[0]),.doutb(w_n13169_0[1]),.doutc(w_n13169_0[2]),.din(n13169));
	jspl jspl_w_n13170_0(.douta(w_n13170_0[0]),.doutb(w_n13170_0[1]),.din(n13170));
	jspl3 jspl3_w_n13174_0(.douta(w_n13174_0[0]),.doutb(w_n13174_0[1]),.doutc(w_n13174_0[2]),.din(n13174));
	jspl3 jspl3_w_n13177_0(.douta(w_n13177_0[0]),.doutb(w_n13177_0[1]),.doutc(w_n13177_0[2]),.din(n13177));
	jspl jspl_w_n13178_0(.douta(w_n13178_0[0]),.doutb(w_n13178_0[1]),.din(n13178));
	jspl3 jspl3_w_n13182_0(.douta(w_n13182_0[0]),.doutb(w_n13182_0[1]),.doutc(w_n13182_0[2]),.din(n13182));
	jspl3 jspl3_w_n13184_0(.douta(w_n13184_0[0]),.doutb(w_n13184_0[1]),.doutc(w_n13184_0[2]),.din(n13184));
	jspl jspl_w_n13185_0(.douta(w_n13185_0[0]),.doutb(w_n13185_0[1]),.din(n13185));
	jspl3 jspl3_w_n13189_0(.douta(w_n13189_0[0]),.doutb(w_n13189_0[1]),.doutc(w_n13189_0[2]),.din(n13189));
	jspl3 jspl3_w_n13191_0(.douta(w_n13191_0[0]),.doutb(w_n13191_0[1]),.doutc(w_n13191_0[2]),.din(n13191));
	jspl jspl_w_n13192_0(.douta(w_n13192_0[0]),.doutb(w_n13192_0[1]),.din(n13192));
	jspl3 jspl3_w_n13196_0(.douta(w_n13196_0[0]),.doutb(w_n13196_0[1]),.doutc(w_n13196_0[2]),.din(n13196));
	jspl3 jspl3_w_n13198_0(.douta(w_n13198_0[0]),.doutb(w_n13198_0[1]),.doutc(w_n13198_0[2]),.din(n13198));
	jspl jspl_w_n13199_0(.douta(w_n13199_0[0]),.doutb(w_n13199_0[1]),.din(n13199));
	jspl3 jspl3_w_n13203_0(.douta(w_n13203_0[0]),.doutb(w_n13203_0[1]),.doutc(w_n13203_0[2]),.din(n13203));
	jspl3 jspl3_w_n13206_0(.douta(w_n13206_0[0]),.doutb(w_n13206_0[1]),.doutc(w_n13206_0[2]),.din(n13206));
	jspl jspl_w_n13207_0(.douta(w_n13207_0[0]),.doutb(w_n13207_0[1]),.din(n13207));
	jspl3 jspl3_w_n13211_0(.douta(w_n13211_0[0]),.doutb(w_n13211_0[1]),.doutc(w_n13211_0[2]),.din(n13211));
	jspl3 jspl3_w_n13213_0(.douta(w_n13213_0[0]),.doutb(w_n13213_0[1]),.doutc(w_n13213_0[2]),.din(n13213));
	jspl jspl_w_n13214_0(.douta(w_n13214_0[0]),.doutb(w_n13214_0[1]),.din(n13214));
	jspl3 jspl3_w_n13218_0(.douta(w_n13218_0[0]),.doutb(w_n13218_0[1]),.doutc(w_n13218_0[2]),.din(n13218));
	jspl3 jspl3_w_n13221_0(.douta(w_n13221_0[0]),.doutb(w_n13221_0[1]),.doutc(w_n13221_0[2]),.din(n13221));
	jspl jspl_w_n13222_0(.douta(w_n13222_0[0]),.doutb(w_n13222_0[1]),.din(n13222));
	jspl3 jspl3_w_n13226_0(.douta(w_n13226_0[0]),.doutb(w_n13226_0[1]),.doutc(w_n13226_0[2]),.din(n13226));
	jspl3 jspl3_w_n13228_0(.douta(w_n13228_0[0]),.doutb(w_n13228_0[1]),.doutc(w_n13228_0[2]),.din(n13228));
	jspl jspl_w_n13229_0(.douta(w_n13229_0[0]),.doutb(w_n13229_0[1]),.din(n13229));
	jspl3 jspl3_w_n13233_0(.douta(w_n13233_0[0]),.doutb(w_n13233_0[1]),.doutc(w_n13233_0[2]),.din(n13233));
	jspl3 jspl3_w_n13236_0(.douta(w_n13236_0[0]),.doutb(w_n13236_0[1]),.doutc(w_n13236_0[2]),.din(n13236));
	jspl jspl_w_n13237_0(.douta(w_n13237_0[0]),.doutb(w_n13237_0[1]),.din(n13237));
	jspl3 jspl3_w_n13241_0(.douta(w_n13241_0[0]),.doutb(w_n13241_0[1]),.doutc(w_n13241_0[2]),.din(n13241));
	jspl3 jspl3_w_n13243_0(.douta(w_n13243_0[0]),.doutb(w_n13243_0[1]),.doutc(w_n13243_0[2]),.din(n13243));
	jspl jspl_w_n13244_0(.douta(w_n13244_0[0]),.doutb(w_n13244_0[1]),.din(n13244));
	jspl3 jspl3_w_n13248_0(.douta(w_n13248_0[0]),.doutb(w_n13248_0[1]),.doutc(w_n13248_0[2]),.din(n13248));
	jspl3 jspl3_w_n13251_0(.douta(w_n13251_0[0]),.doutb(w_n13251_0[1]),.doutc(w_n13251_0[2]),.din(n13251));
	jspl jspl_w_n13252_0(.douta(w_n13252_0[0]),.doutb(w_n13252_0[1]),.din(n13252));
	jspl3 jspl3_w_n13256_0(.douta(w_n13256_0[0]),.doutb(w_n13256_0[1]),.doutc(w_n13256_0[2]),.din(n13256));
	jspl3 jspl3_w_n13259_0(.douta(w_n13259_0[0]),.doutb(w_n13259_0[1]),.doutc(w_n13259_0[2]),.din(n13259));
	jspl jspl_w_n13260_0(.douta(w_n13260_0[0]),.doutb(w_n13260_0[1]),.din(n13260));
	jspl3 jspl3_w_n13264_0(.douta(w_n13264_0[0]),.doutb(w_n13264_0[1]),.doutc(w_n13264_0[2]),.din(n13264));
	jspl3 jspl3_w_n13267_0(.douta(w_n13267_0[0]),.doutb(w_n13267_0[1]),.doutc(w_n13267_0[2]),.din(n13267));
	jspl jspl_w_n13268_0(.douta(w_n13268_0[0]),.doutb(w_n13268_0[1]),.din(n13268));
	jspl3 jspl3_w_n13272_0(.douta(w_n13272_0[0]),.doutb(w_n13272_0[1]),.doutc(w_n13272_0[2]),.din(n13272));
	jspl3 jspl3_w_n13274_0(.douta(w_n13274_0[0]),.doutb(w_n13274_0[1]),.doutc(w_n13274_0[2]),.din(n13274));
	jspl jspl_w_n13275_0(.douta(w_n13275_0[0]),.doutb(w_n13275_0[1]),.din(n13275));
	jspl3 jspl3_w_n13279_0(.douta(w_n13279_0[0]),.doutb(w_n13279_0[1]),.doutc(w_n13279_0[2]),.din(n13279));
	jspl3 jspl3_w_n13281_0(.douta(w_n13281_0[0]),.doutb(w_n13281_0[1]),.doutc(w_n13281_0[2]),.din(n13281));
	jspl jspl_w_n13282_0(.douta(w_n13282_0[0]),.doutb(w_n13282_0[1]),.din(n13282));
	jspl jspl_w_n13285_0(.douta(w_n13285_0[0]),.doutb(w_n13285_0[1]),.din(n13285));
	jspl3 jspl3_w_n13287_0(.douta(w_n13287_0[0]),.doutb(w_n13287_0[1]),.doutc(w_n13287_0[2]),.din(n13287));
	jspl jspl_w_n13287_1(.douta(w_n13287_1[0]),.doutb(w_n13287_1[1]),.din(w_n13287_0[0]));
	jspl jspl_w_n13292_0(.douta(w_n13292_0[0]),.doutb(w_n13292_0[1]),.din(n13292));
	jspl jspl_w_n13294_0(.douta(w_n13294_0[0]),.doutb(w_n13294_0[1]),.din(n13294));
	jspl3 jspl3_w_n13296_0(.douta(w_n13296_0[0]),.doutb(w_n13296_0[1]),.doutc(w_n13296_0[2]),.din(n13296));
	jspl jspl_w_n13296_1(.douta(w_n13296_1[0]),.doutb(w_n13296_1[1]),.din(w_n13296_0[0]));
	jspl jspl_w_n13297_0(.douta(w_n13297_0[0]),.doutb(w_n13297_0[1]),.din(n13297));
	jspl3 jspl3_w_n13298_0(.douta(w_n13298_0[0]),.doutb(w_n13298_0[1]),.doutc(w_n13298_0[2]),.din(n13298));
	jspl jspl_w_n13299_0(.douta(w_n13299_0[0]),.doutb(w_n13299_0[1]),.din(n13299));
	jspl3 jspl3_w_n13301_0(.douta(w_n13301_0[0]),.doutb(w_n13301_0[1]),.doutc(w_n13301_0[2]),.din(n13301));
	jspl jspl_w_n13302_0(.douta(w_n13302_0[0]),.doutb(w_n13302_0[1]),.din(n13302));
	jspl jspl_w_n13510_0(.douta(w_n13510_0[0]),.doutb(w_n13510_0[1]),.din(n13510));
	jspl3 jspl3_w_n13515_0(.douta(w_n13515_0[0]),.doutb(w_n13515_0[1]),.doutc(w_n13515_0[2]),.din(n13515));
	jspl3 jspl3_w_n13515_1(.douta(w_n13515_1[0]),.doutb(w_n13515_1[1]),.doutc(w_n13515_1[2]),.din(w_n13515_0[0]));
	jspl3 jspl3_w_n13515_2(.douta(w_n13515_2[0]),.doutb(w_n13515_2[1]),.doutc(w_n13515_2[2]),.din(w_n13515_0[1]));
	jspl3 jspl3_w_n13515_3(.douta(w_n13515_3[0]),.doutb(w_n13515_3[1]),.doutc(w_n13515_3[2]),.din(w_n13515_0[2]));
	jspl3 jspl3_w_n13515_4(.douta(w_n13515_4[0]),.doutb(w_n13515_4[1]),.doutc(w_n13515_4[2]),.din(w_n13515_1[0]));
	jspl3 jspl3_w_n13515_5(.douta(w_n13515_5[0]),.doutb(w_n13515_5[1]),.doutc(w_n13515_5[2]),.din(w_n13515_1[1]));
	jspl3 jspl3_w_n13515_6(.douta(w_n13515_6[0]),.doutb(w_n13515_6[1]),.doutc(w_n13515_6[2]),.din(w_n13515_1[2]));
	jspl3 jspl3_w_n13515_7(.douta(w_n13515_7[0]),.doutb(w_n13515_7[1]),.doutc(w_n13515_7[2]),.din(w_n13515_2[0]));
	jspl3 jspl3_w_n13515_8(.douta(w_n13515_8[0]),.doutb(w_n13515_8[1]),.doutc(w_n13515_8[2]),.din(w_n13515_2[1]));
	jspl3 jspl3_w_n13515_9(.douta(w_n13515_9[0]),.doutb(w_n13515_9[1]),.doutc(w_n13515_9[2]),.din(w_n13515_2[2]));
	jspl3 jspl3_w_n13515_10(.douta(w_n13515_10[0]),.doutb(w_n13515_10[1]),.doutc(w_n13515_10[2]),.din(w_n13515_3[0]));
	jspl3 jspl3_w_n13515_11(.douta(w_n13515_11[0]),.doutb(w_n13515_11[1]),.doutc(w_n13515_11[2]),.din(w_n13515_3[1]));
	jspl3 jspl3_w_n13515_12(.douta(w_n13515_12[0]),.doutb(w_n13515_12[1]),.doutc(w_n13515_12[2]),.din(w_n13515_3[2]));
	jspl3 jspl3_w_n13515_13(.douta(w_n13515_13[0]),.doutb(w_n13515_13[1]),.doutc(w_n13515_13[2]),.din(w_n13515_4[0]));
	jspl3 jspl3_w_n13515_14(.douta(w_n13515_14[0]),.doutb(w_n13515_14[1]),.doutc(w_n13515_14[2]),.din(w_n13515_4[1]));
	jspl3 jspl3_w_n13515_15(.douta(w_n13515_15[0]),.doutb(w_n13515_15[1]),.doutc(w_n13515_15[2]),.din(w_n13515_4[2]));
	jspl3 jspl3_w_n13515_16(.douta(w_n13515_16[0]),.doutb(w_n13515_16[1]),.doutc(w_n13515_16[2]),.din(w_n13515_5[0]));
	jspl3 jspl3_w_n13515_17(.douta(w_n13515_17[0]),.doutb(w_n13515_17[1]),.doutc(w_n13515_17[2]),.din(w_n13515_5[1]));
	jspl3 jspl3_w_n13515_18(.douta(w_n13515_18[0]),.doutb(w_n13515_18[1]),.doutc(w_n13515_18[2]),.din(w_n13515_5[2]));
	jspl3 jspl3_w_n13515_19(.douta(w_n13515_19[0]),.doutb(w_n13515_19[1]),.doutc(w_n13515_19[2]),.din(w_n13515_6[0]));
	jspl3 jspl3_w_n13515_20(.douta(w_n13515_20[0]),.doutb(w_n13515_20[1]),.doutc(w_n13515_20[2]),.din(w_n13515_6[1]));
	jspl3 jspl3_w_n13515_21(.douta(w_n13515_21[0]),.doutb(w_n13515_21[1]),.doutc(w_n13515_21[2]),.din(w_n13515_6[2]));
	jspl3 jspl3_w_n13515_22(.douta(w_n13515_22[0]),.doutb(w_n13515_22[1]),.doutc(w_n13515_22[2]),.din(w_n13515_7[0]));
	jspl jspl_w_n13515_23(.douta(w_n13515_23[0]),.doutb(w_n13515_23[1]),.din(w_n13515_7[1]));
	jspl jspl_w_n13516_0(.douta(w_n13516_0[0]),.doutb(w_n13516_0[1]),.din(n13516));
	jspl3 jspl3_w_n13519_0(.douta(w_n13519_0[0]),.doutb(w_n13519_0[1]),.doutc(w_n13519_0[2]),.din(n13519));
	jspl jspl_w_n13520_0(.douta(w_n13520_0[0]),.doutb(w_n13520_0[1]),.din(n13520));
	jspl jspl_w_n13526_0(.douta(w_n13526_0[0]),.doutb(w_n13526_0[1]),.din(n13526));
	jspl jspl_w_n13527_0(.douta(w_n13527_0[0]),.doutb(w_n13527_0[1]),.din(n13527));
	jspl3 jspl3_w_n13529_0(.douta(w_n13529_0[0]),.doutb(w_n13529_0[1]),.doutc(w_n13529_0[2]),.din(n13529));
	jspl jspl_w_n13530_0(.douta(w_n13530_0[0]),.doutb(w_n13530_0[1]),.din(n13530));
	jspl jspl_w_n13534_0(.douta(w_n13534_0[0]),.doutb(w_n13534_0[1]),.din(n13534));
	jspl jspl_w_n13535_0(.douta(w_n13535_0[0]),.doutb(w_n13535_0[1]),.din(n13535));
	jspl3 jspl3_w_n13537_0(.douta(w_n13537_0[0]),.doutb(w_n13537_0[1]),.doutc(w_n13537_0[2]),.din(n13537));
	jspl jspl_w_n13538_0(.douta(w_n13538_0[0]),.doutb(w_n13538_0[1]),.din(n13538));
	jspl jspl_w_n13542_0(.douta(w_n13542_0[0]),.doutb(w_n13542_0[1]),.din(n13542));
	jspl jspl_w_n13543_0(.douta(w_n13543_0[0]),.doutb(w_n13543_0[1]),.din(n13543));
	jspl3 jspl3_w_n13545_0(.douta(w_n13545_0[0]),.doutb(w_n13545_0[1]),.doutc(w_n13545_0[2]),.din(n13545));
	jspl jspl_w_n13546_0(.douta(w_n13546_0[0]),.doutb(w_n13546_0[1]),.din(n13546));
	jspl jspl_w_n13550_0(.douta(w_n13550_0[0]),.doutb(w_n13550_0[1]),.din(n13550));
	jspl3 jspl3_w_n13552_0(.douta(w_n13552_0[0]),.doutb(w_n13552_0[1]),.doutc(w_n13552_0[2]),.din(n13552));
	jspl jspl_w_n13553_0(.douta(w_n13553_0[0]),.doutb(w_n13553_0[1]),.din(n13553));
	jspl jspl_w_n13557_0(.douta(w_n13557_0[0]),.doutb(w_n13557_0[1]),.din(n13557));
	jspl jspl_w_n13558_0(.douta(w_n13558_0[0]),.doutb(w_n13558_0[1]),.din(n13558));
	jspl3 jspl3_w_n13560_0(.douta(w_n13560_0[0]),.doutb(w_n13560_0[1]),.doutc(w_n13560_0[2]),.din(n13560));
	jspl jspl_w_n13561_0(.douta(w_n13561_0[0]),.doutb(w_n13561_0[1]),.din(n13561));
	jspl jspl_w_n13565_0(.douta(w_n13565_0[0]),.doutb(w_n13565_0[1]),.din(n13565));
	jspl3 jspl3_w_n13567_0(.douta(w_n13567_0[0]),.doutb(w_n13567_0[1]),.doutc(w_n13567_0[2]),.din(n13567));
	jspl jspl_w_n13568_0(.douta(w_n13568_0[0]),.doutb(w_n13568_0[1]),.din(n13568));
	jspl jspl_w_n13572_0(.douta(w_n13572_0[0]),.doutb(w_n13572_0[1]),.din(n13572));
	jspl jspl_w_n13573_0(.douta(w_n13573_0[0]),.doutb(w_n13573_0[1]),.din(n13573));
	jspl3 jspl3_w_n13575_0(.douta(w_n13575_0[0]),.doutb(w_n13575_0[1]),.doutc(w_n13575_0[2]),.din(n13575));
	jspl jspl_w_n13576_0(.douta(w_n13576_0[0]),.doutb(w_n13576_0[1]),.din(n13576));
	jspl jspl_w_n13580_0(.douta(w_n13580_0[0]),.doutb(w_n13580_0[1]),.din(n13580));
	jspl3 jspl3_w_n13582_0(.douta(w_n13582_0[0]),.doutb(w_n13582_0[1]),.doutc(w_n13582_0[2]),.din(n13582));
	jspl jspl_w_n13583_0(.douta(w_n13583_0[0]),.doutb(w_n13583_0[1]),.din(n13583));
	jspl jspl_w_n13587_0(.douta(w_n13587_0[0]),.doutb(w_n13587_0[1]),.din(n13587));
	jspl jspl_w_n13588_0(.douta(w_n13588_0[0]),.doutb(w_n13588_0[1]),.din(n13588));
	jspl3 jspl3_w_n13590_0(.douta(w_n13590_0[0]),.doutb(w_n13590_0[1]),.doutc(w_n13590_0[2]),.din(n13590));
	jspl jspl_w_n13591_0(.douta(w_n13591_0[0]),.doutb(w_n13591_0[1]),.din(n13591));
	jspl jspl_w_n13595_0(.douta(w_n13595_0[0]),.doutb(w_n13595_0[1]),.din(n13595));
	jspl3 jspl3_w_n13597_0(.douta(w_n13597_0[0]),.doutb(w_n13597_0[1]),.doutc(w_n13597_0[2]),.din(n13597));
	jspl jspl_w_n13598_0(.douta(w_n13598_0[0]),.doutb(w_n13598_0[1]),.din(n13598));
	jspl jspl_w_n13602_0(.douta(w_n13602_0[0]),.doutb(w_n13602_0[1]),.din(n13602));
	jspl jspl_w_n13603_0(.douta(w_n13603_0[0]),.doutb(w_n13603_0[1]),.din(n13603));
	jspl3 jspl3_w_n13605_0(.douta(w_n13605_0[0]),.doutb(w_n13605_0[1]),.doutc(w_n13605_0[2]),.din(n13605));
	jspl jspl_w_n13606_0(.douta(w_n13606_0[0]),.doutb(w_n13606_0[1]),.din(n13606));
	jspl jspl_w_n13610_0(.douta(w_n13610_0[0]),.doutb(w_n13610_0[1]),.din(n13610));
	jspl jspl_w_n13611_0(.douta(w_n13611_0[0]),.doutb(w_n13611_0[1]),.din(n13611));
	jspl3 jspl3_w_n13613_0(.douta(w_n13613_0[0]),.doutb(w_n13613_0[1]),.doutc(w_n13613_0[2]),.din(n13613));
	jspl jspl_w_n13614_0(.douta(w_n13614_0[0]),.doutb(w_n13614_0[1]),.din(n13614));
	jspl jspl_w_n13618_0(.douta(w_n13618_0[0]),.doutb(w_n13618_0[1]),.din(n13618));
	jspl jspl_w_n13619_0(.douta(w_n13619_0[0]),.doutb(w_n13619_0[1]),.din(n13619));
	jspl3 jspl3_w_n13621_0(.douta(w_n13621_0[0]),.doutb(w_n13621_0[1]),.doutc(w_n13621_0[2]),.din(n13621));
	jspl jspl_w_n13622_0(.douta(w_n13622_0[0]),.doutb(w_n13622_0[1]),.din(n13622));
	jspl jspl_w_n13626_0(.douta(w_n13626_0[0]),.doutb(w_n13626_0[1]),.din(n13626));
	jspl3 jspl3_w_n13628_0(.douta(w_n13628_0[0]),.doutb(w_n13628_0[1]),.doutc(w_n13628_0[2]),.din(n13628));
	jspl jspl_w_n13629_0(.douta(w_n13629_0[0]),.doutb(w_n13629_0[1]),.din(n13629));
	jspl jspl_w_n13633_0(.douta(w_n13633_0[0]),.doutb(w_n13633_0[1]),.din(n13633));
	jspl jspl_w_n13634_0(.douta(w_n13634_0[0]),.doutb(w_n13634_0[1]),.din(n13634));
	jspl3 jspl3_w_n13636_0(.douta(w_n13636_0[0]),.doutb(w_n13636_0[1]),.doutc(w_n13636_0[2]),.din(n13636));
	jspl jspl_w_n13637_0(.douta(w_n13637_0[0]),.doutb(w_n13637_0[1]),.din(n13637));
	jspl jspl_w_n13641_0(.douta(w_n13641_0[0]),.doutb(w_n13641_0[1]),.din(n13641));
	jspl3 jspl3_w_n13643_0(.douta(w_n13643_0[0]),.doutb(w_n13643_0[1]),.doutc(w_n13643_0[2]),.din(n13643));
	jspl jspl_w_n13644_0(.douta(w_n13644_0[0]),.doutb(w_n13644_0[1]),.din(n13644));
	jspl jspl_w_n13648_0(.douta(w_n13648_0[0]),.doutb(w_n13648_0[1]),.din(n13648));
	jspl jspl_w_n13649_0(.douta(w_n13649_0[0]),.doutb(w_n13649_0[1]),.din(n13649));
	jspl3 jspl3_w_n13651_0(.douta(w_n13651_0[0]),.doutb(w_n13651_0[1]),.doutc(w_n13651_0[2]),.din(n13651));
	jspl jspl_w_n13652_0(.douta(w_n13652_0[0]),.doutb(w_n13652_0[1]),.din(n13652));
	jspl jspl_w_n13656_0(.douta(w_n13656_0[0]),.doutb(w_n13656_0[1]),.din(n13656));
	jspl jspl_w_n13657_0(.douta(w_n13657_0[0]),.doutb(w_n13657_0[1]),.din(n13657));
	jspl3 jspl3_w_n13659_0(.douta(w_n13659_0[0]),.doutb(w_n13659_0[1]),.doutc(w_n13659_0[2]),.din(n13659));
	jspl jspl_w_n13660_0(.douta(w_n13660_0[0]),.doutb(w_n13660_0[1]),.din(n13660));
	jspl jspl_w_n13664_0(.douta(w_n13664_0[0]),.doutb(w_n13664_0[1]),.din(n13664));
	jspl jspl_w_n13665_0(.douta(w_n13665_0[0]),.doutb(w_n13665_0[1]),.din(n13665));
	jspl3 jspl3_w_n13667_0(.douta(w_n13667_0[0]),.doutb(w_n13667_0[1]),.doutc(w_n13667_0[2]),.din(n13667));
	jspl jspl_w_n13668_0(.douta(w_n13668_0[0]),.doutb(w_n13668_0[1]),.din(n13668));
	jspl jspl_w_n13672_0(.douta(w_n13672_0[0]),.doutb(w_n13672_0[1]),.din(n13672));
	jspl3 jspl3_w_n13674_0(.douta(w_n13674_0[0]),.doutb(w_n13674_0[1]),.doutc(w_n13674_0[2]),.din(n13674));
	jspl jspl_w_n13675_0(.douta(w_n13675_0[0]),.doutb(w_n13675_0[1]),.din(n13675));
	jspl jspl_w_n13679_0(.douta(w_n13679_0[0]),.doutb(w_n13679_0[1]),.din(n13679));
	jspl jspl_w_n13680_0(.douta(w_n13680_0[0]),.doutb(w_n13680_0[1]),.din(n13680));
	jspl3 jspl3_w_n13682_0(.douta(w_n13682_0[0]),.doutb(w_n13682_0[1]),.doutc(w_n13682_0[2]),.din(n13682));
	jspl jspl_w_n13683_0(.douta(w_n13683_0[0]),.doutb(w_n13683_0[1]),.din(n13683));
	jspl jspl_w_n13687_0(.douta(w_n13687_0[0]),.doutb(w_n13687_0[1]),.din(n13687));
	jspl jspl_w_n13688_0(.douta(w_n13688_0[0]),.doutb(w_n13688_0[1]),.din(n13688));
	jspl3 jspl3_w_n13690_0(.douta(w_n13690_0[0]),.doutb(w_n13690_0[1]),.doutc(w_n13690_0[2]),.din(n13690));
	jspl jspl_w_n13691_0(.douta(w_n13691_0[0]),.doutb(w_n13691_0[1]),.din(n13691));
	jspl jspl_w_n13695_0(.douta(w_n13695_0[0]),.doutb(w_n13695_0[1]),.din(n13695));
	jspl jspl_w_n13696_0(.douta(w_n13696_0[0]),.doutb(w_n13696_0[1]),.din(n13696));
	jspl3 jspl3_w_n13698_0(.douta(w_n13698_0[0]),.doutb(w_n13698_0[1]),.doutc(w_n13698_0[2]),.din(n13698));
	jspl jspl_w_n13699_0(.douta(w_n13699_0[0]),.doutb(w_n13699_0[1]),.din(n13699));
	jspl jspl_w_n13703_0(.douta(w_n13703_0[0]),.doutb(w_n13703_0[1]),.din(n13703));
	jspl jspl_w_n13704_0(.douta(w_n13704_0[0]),.doutb(w_n13704_0[1]),.din(n13704));
	jspl3 jspl3_w_n13706_0(.douta(w_n13706_0[0]),.doutb(w_n13706_0[1]),.doutc(w_n13706_0[2]),.din(n13706));
	jspl jspl_w_n13707_0(.douta(w_n13707_0[0]),.doutb(w_n13707_0[1]),.din(n13707));
	jspl jspl_w_n13711_0(.douta(w_n13711_0[0]),.doutb(w_n13711_0[1]),.din(n13711));
	jspl3 jspl3_w_n13713_0(.douta(w_n13713_0[0]),.doutb(w_n13713_0[1]),.doutc(w_n13713_0[2]),.din(n13713));
	jspl jspl_w_n13714_0(.douta(w_n13714_0[0]),.doutb(w_n13714_0[1]),.din(n13714));
	jspl jspl_w_n13717_0(.douta(w_n13717_0[0]),.doutb(w_n13717_0[1]),.din(n13717));
	jspl3 jspl3_w_n13720_0(.douta(w_n13720_0[0]),.doutb(w_n13720_0[1]),.doutc(w_n13720_0[2]),.din(n13720));
	jspl jspl_w_n13721_0(.douta(w_n13721_0[0]),.doutb(w_n13721_0[1]),.din(n13721));
	jspl jspl_w_n13725_0(.douta(w_n13725_0[0]),.doutb(w_n13725_0[1]),.din(n13725));
	jspl jspl_w_n13726_0(.douta(w_n13726_0[0]),.doutb(w_n13726_0[1]),.din(n13726));
	jspl3 jspl3_w_n13728_0(.douta(w_n13728_0[0]),.doutb(w_n13728_0[1]),.doutc(w_n13728_0[2]),.din(n13728));
	jspl jspl_w_n13729_0(.douta(w_n13729_0[0]),.doutb(w_n13729_0[1]),.din(n13729));
	jspl jspl_w_n13733_0(.douta(w_n13733_0[0]),.doutb(w_n13733_0[1]),.din(n13733));
	jspl3 jspl3_w_n13735_0(.douta(w_n13735_0[0]),.doutb(w_n13735_0[1]),.doutc(w_n13735_0[2]),.din(n13735));
	jspl jspl_w_n13736_0(.douta(w_n13736_0[0]),.doutb(w_n13736_0[1]),.din(n13736));
	jspl jspl_w_n13740_0(.douta(w_n13740_0[0]),.doutb(w_n13740_0[1]),.din(n13740));
	jspl jspl_w_n13741_0(.douta(w_n13741_0[0]),.doutb(w_n13741_0[1]),.din(n13741));
	jspl3 jspl3_w_n13743_0(.douta(w_n13743_0[0]),.doutb(w_n13743_0[1]),.doutc(w_n13743_0[2]),.din(n13743));
	jspl jspl_w_n13744_0(.douta(w_n13744_0[0]),.doutb(w_n13744_0[1]),.din(n13744));
	jspl jspl_w_n13748_0(.douta(w_n13748_0[0]),.doutb(w_n13748_0[1]),.din(n13748));
	jspl3 jspl3_w_n13750_0(.douta(w_n13750_0[0]),.doutb(w_n13750_0[1]),.doutc(w_n13750_0[2]),.din(n13750));
	jspl jspl_w_n13751_0(.douta(w_n13751_0[0]),.doutb(w_n13751_0[1]),.din(n13751));
	jspl jspl_w_n13755_0(.douta(w_n13755_0[0]),.doutb(w_n13755_0[1]),.din(n13755));
	jspl jspl_w_n13756_0(.douta(w_n13756_0[0]),.doutb(w_n13756_0[1]),.din(n13756));
	jspl3 jspl3_w_n13758_0(.douta(w_n13758_0[0]),.doutb(w_n13758_0[1]),.doutc(w_n13758_0[2]),.din(n13758));
	jspl jspl_w_n13759_0(.douta(w_n13759_0[0]),.doutb(w_n13759_0[1]),.din(n13759));
	jspl jspl_w_n13763_0(.douta(w_n13763_0[0]),.doutb(w_n13763_0[1]),.din(n13763));
	jspl jspl_w_n13764_0(.douta(w_n13764_0[0]),.doutb(w_n13764_0[1]),.din(n13764));
	jspl3 jspl3_w_n13766_0(.douta(w_n13766_0[0]),.doutb(w_n13766_0[1]),.doutc(w_n13766_0[2]),.din(n13766));
	jspl jspl_w_n13767_0(.douta(w_n13767_0[0]),.doutb(w_n13767_0[1]),.din(n13767));
	jspl jspl_w_n13771_0(.douta(w_n13771_0[0]),.doutb(w_n13771_0[1]),.din(n13771));
	jspl jspl_w_n13772_0(.douta(w_n13772_0[0]),.doutb(w_n13772_0[1]),.din(n13772));
	jspl3 jspl3_w_n13774_0(.douta(w_n13774_0[0]),.doutb(w_n13774_0[1]),.doutc(w_n13774_0[2]),.din(n13774));
	jspl jspl_w_n13775_0(.douta(w_n13775_0[0]),.doutb(w_n13775_0[1]),.din(n13775));
	jspl jspl_w_n13779_0(.douta(w_n13779_0[0]),.doutb(w_n13779_0[1]),.din(n13779));
	jspl3 jspl3_w_n13781_0(.douta(w_n13781_0[0]),.doutb(w_n13781_0[1]),.doutc(w_n13781_0[2]),.din(n13781));
	jspl jspl_w_n13782_0(.douta(w_n13782_0[0]),.doutb(w_n13782_0[1]),.din(n13782));
	jspl jspl_w_n13786_0(.douta(w_n13786_0[0]),.doutb(w_n13786_0[1]),.din(n13786));
	jspl jspl_w_n13787_0(.douta(w_n13787_0[0]),.doutb(w_n13787_0[1]),.din(n13787));
	jspl3 jspl3_w_n13789_0(.douta(w_n13789_0[0]),.doutb(w_n13789_0[1]),.doutc(w_n13789_0[2]),.din(n13789));
	jspl jspl_w_n13790_0(.douta(w_n13790_0[0]),.doutb(w_n13790_0[1]),.din(n13790));
	jspl jspl_w_n13794_0(.douta(w_n13794_0[0]),.doutb(w_n13794_0[1]),.din(n13794));
	jspl3 jspl3_w_n13796_0(.douta(w_n13796_0[0]),.doutb(w_n13796_0[1]),.doutc(w_n13796_0[2]),.din(n13796));
	jspl jspl_w_n13797_0(.douta(w_n13797_0[0]),.doutb(w_n13797_0[1]),.din(n13797));
	jspl jspl_w_n13801_0(.douta(w_n13801_0[0]),.doutb(w_n13801_0[1]),.din(n13801));
	jspl jspl_w_n13802_0(.douta(w_n13802_0[0]),.doutb(w_n13802_0[1]),.din(n13802));
	jspl3 jspl3_w_n13804_0(.douta(w_n13804_0[0]),.doutb(w_n13804_0[1]),.doutc(w_n13804_0[2]),.din(n13804));
	jspl jspl_w_n13805_0(.douta(w_n13805_0[0]),.doutb(w_n13805_0[1]),.din(n13805));
	jspl jspl_w_n13809_0(.douta(w_n13809_0[0]),.doutb(w_n13809_0[1]),.din(n13809));
	jspl3 jspl3_w_n13811_0(.douta(w_n13811_0[0]),.doutb(w_n13811_0[1]),.doutc(w_n13811_0[2]),.din(n13811));
	jspl jspl_w_n13812_0(.douta(w_n13812_0[0]),.doutb(w_n13812_0[1]),.din(n13812));
	jspl jspl_w_n13816_0(.douta(w_n13816_0[0]),.doutb(w_n13816_0[1]),.din(n13816));
	jspl jspl_w_n13817_0(.douta(w_n13817_0[0]),.doutb(w_n13817_0[1]),.din(n13817));
	jspl3 jspl3_w_n13819_0(.douta(w_n13819_0[0]),.doutb(w_n13819_0[1]),.doutc(w_n13819_0[2]),.din(n13819));
	jspl jspl_w_n13820_0(.douta(w_n13820_0[0]),.doutb(w_n13820_0[1]),.din(n13820));
	jspl jspl_w_n13824_0(.douta(w_n13824_0[0]),.doutb(w_n13824_0[1]),.din(n13824));
	jspl3 jspl3_w_n13826_0(.douta(w_n13826_0[0]),.doutb(w_n13826_0[1]),.doutc(w_n13826_0[2]),.din(n13826));
	jspl jspl_w_n13827_0(.douta(w_n13827_0[0]),.doutb(w_n13827_0[1]),.din(n13827));
	jspl jspl_w_n13831_0(.douta(w_n13831_0[0]),.doutb(w_n13831_0[1]),.din(n13831));
	jspl3 jspl3_w_n13833_0(.douta(w_n13833_0[0]),.doutb(w_n13833_0[1]),.doutc(w_n13833_0[2]),.din(n13833));
	jspl jspl_w_n13834_0(.douta(w_n13834_0[0]),.doutb(w_n13834_0[1]),.din(n13834));
	jspl jspl_w_n13838_0(.douta(w_n13838_0[0]),.doutb(w_n13838_0[1]),.din(n13838));
	jspl3 jspl3_w_n13840_0(.douta(w_n13840_0[0]),.doutb(w_n13840_0[1]),.doutc(w_n13840_0[2]),.din(n13840));
	jspl jspl_w_n13841_0(.douta(w_n13841_0[0]),.doutb(w_n13841_0[1]),.din(n13841));
	jspl jspl_w_n13845_0(.douta(w_n13845_0[0]),.doutb(w_n13845_0[1]),.din(n13845));
	jspl jspl_w_n13846_0(.douta(w_n13846_0[0]),.doutb(w_n13846_0[1]),.din(n13846));
	jspl3 jspl3_w_n13848_0(.douta(w_n13848_0[0]),.doutb(w_n13848_0[1]),.doutc(w_n13848_0[2]),.din(n13848));
	jspl jspl_w_n13851_0(.douta(w_n13851_0[0]),.doutb(w_n13851_0[1]),.din(n13851));
	jspl3 jspl3_w_n13852_0(.douta(w_n13852_0[0]),.doutb(w_n13852_0[1]),.doutc(w_n13852_0[2]),.din(n13852));
	jspl jspl_w_n13853_0(.douta(w_n13853_0[0]),.doutb(w_n13853_0[1]),.din(n13853));
	jspl jspl_w_n13854_0(.douta(w_n13854_0[0]),.doutb(w_n13854_0[1]),.din(n13854));
	jspl jspl_w_n13859_0(.douta(w_n13859_0[0]),.doutb(w_n13859_0[1]),.din(n13859));
	jspl jspl_w_n13860_0(.douta(w_n13860_0[0]),.doutb(w_n13860_0[1]),.din(n13860));
	jspl jspl_w_n13879_0(.douta(w_n13879_0[0]),.doutb(w_n13879_0[1]),.din(n13879));
	jspl jspl_w_n13913_0(.douta(w_n13913_0[0]),.doutb(w_n13913_0[1]),.din(n13913));
	jspl jspl_w_n13926_0(.douta(w_n13926_0[0]),.doutb(w_n13926_0[1]),.din(n13926));
	jspl jspl_w_n13933_0(.douta(w_n13933_0[0]),.doutb(w_n13933_0[1]),.din(n13933));
	jspl jspl_w_n13940_0(.douta(w_n13940_0[0]),.doutb(w_n13940_0[1]),.din(n13940));
	jspl jspl_w_n13947_0(.douta(w_n13947_0[0]),.doutb(w_n13947_0[1]),.din(n13947));
	jspl jspl_w_n13960_0(.douta(w_n13960_0[0]),.doutb(w_n13960_0[1]),.din(n13960));
	jspl jspl_w_n13967_0(.douta(w_n13967_0[0]),.doutb(w_n13967_0[1]),.din(n13967));
	jspl jspl_w_n13980_0(.douta(w_n13980_0[0]),.doutb(w_n13980_0[1]),.din(n13980));
	jspl jspl_w_n13996_0(.douta(w_n13996_0[0]),.doutb(w_n13996_0[1]),.din(n13996));
	jspl jspl_w_n14006_0(.douta(w_n14006_0[0]),.doutb(w_n14006_0[1]),.din(n14006));
	jspl jspl_w_n14013_0(.douta(w_n14013_0[0]),.doutb(w_n14013_0[1]),.din(n14013));
	jspl jspl_w_n14026_0(.douta(w_n14026_0[0]),.doutb(w_n14026_0[1]),.din(n14026));
	jspl jspl_w_n14033_0(.douta(w_n14033_0[0]),.doutb(w_n14033_0[1]),.din(n14033));
	jspl jspl_w_n14040_0(.douta(w_n14040_0[0]),.doutb(w_n14040_0[1]),.din(n14040));
	jspl jspl_w_n14047_0(.douta(w_n14047_0[0]),.doutb(w_n14047_0[1]),.din(n14047));
	jspl jspl_w_n14051_0(.douta(w_n14051_0[0]),.doutb(w_n14051_0[1]),.din(n14051));
	jspl jspl_w_n14055_0(.douta(w_n14055_0[0]),.doutb(w_n14055_0[1]),.din(n14055));
	jspl jspl_w_n14060_0(.douta(w_n14060_0[0]),.doutb(w_n14060_0[1]),.din(n14060));
	jspl jspl_w_n14063_0(.douta(w_n14063_0[0]),.doutb(w_n14063_0[1]),.din(n14063));
	jspl jspl_w_n14065_0(.douta(w_n14065_0[0]),.doutb(w_n14065_0[1]),.din(n14065));
	jspl jspl_w_n14066_0(.douta(w_n14066_0[0]),.doutb(w_n14066_0[1]),.din(n14066));
	jspl jspl_w_n14077_0(.douta(w_n14077_0[0]),.doutb(w_n14077_0[1]),.din(n14077));
	jspl3 jspl3_w_n14078_0(.douta(w_n14078_0[0]),.doutb(w_n14078_0[1]),.doutc(w_n14078_0[2]),.din(n14078));
	jspl3 jspl3_w_n14078_1(.douta(w_n14078_1[0]),.doutb(w_n14078_1[1]),.doutc(w_n14078_1[2]),.din(w_n14078_0[0]));
	jspl3 jspl3_w_n14078_2(.douta(w_n14078_2[0]),.doutb(w_n14078_2[1]),.doutc(w_n14078_2[2]),.din(w_n14078_0[1]));
	jspl3 jspl3_w_n14078_3(.douta(w_n14078_3[0]),.doutb(w_n14078_3[1]),.doutc(w_n14078_3[2]),.din(w_n14078_0[2]));
	jspl3 jspl3_w_n14078_4(.douta(w_n14078_4[0]),.doutb(w_n14078_4[1]),.doutc(w_n14078_4[2]),.din(w_n14078_1[0]));
	jspl3 jspl3_w_n14078_5(.douta(w_n14078_5[0]),.doutb(w_n14078_5[1]),.doutc(w_n14078_5[2]),.din(w_n14078_1[1]));
	jspl3 jspl3_w_n14078_6(.douta(w_n14078_6[0]),.doutb(w_n14078_6[1]),.doutc(w_n14078_6[2]),.din(w_n14078_1[2]));
	jspl3 jspl3_w_n14078_7(.douta(w_n14078_7[0]),.doutb(w_n14078_7[1]),.doutc(w_n14078_7[2]),.din(w_n14078_2[0]));
	jspl3 jspl3_w_n14078_8(.douta(w_n14078_8[0]),.doutb(w_n14078_8[1]),.doutc(w_n14078_8[2]),.din(w_n14078_2[1]));
	jspl3 jspl3_w_n14078_9(.douta(w_n14078_9[0]),.doutb(w_n14078_9[1]),.doutc(w_n14078_9[2]),.din(w_n14078_2[2]));
	jspl3 jspl3_w_n14078_10(.douta(w_n14078_10[0]),.doutb(w_n14078_10[1]),.doutc(w_n14078_10[2]),.din(w_n14078_3[0]));
	jspl3 jspl3_w_n14078_11(.douta(w_n14078_11[0]),.doutb(w_n14078_11[1]),.doutc(w_n14078_11[2]),.din(w_n14078_3[1]));
	jspl3 jspl3_w_n14078_12(.douta(w_n14078_12[0]),.doutb(w_n14078_12[1]),.doutc(w_n14078_12[2]),.din(w_n14078_3[2]));
	jspl3 jspl3_w_n14078_13(.douta(w_n14078_13[0]),.doutb(w_n14078_13[1]),.doutc(w_n14078_13[2]),.din(w_n14078_4[0]));
	jspl3 jspl3_w_n14078_14(.douta(w_n14078_14[0]),.doutb(w_n14078_14[1]),.doutc(w_n14078_14[2]),.din(w_n14078_4[1]));
	jspl3 jspl3_w_n14078_15(.douta(w_n14078_15[0]),.doutb(w_n14078_15[1]),.doutc(w_n14078_15[2]),.din(w_n14078_4[2]));
	jspl3 jspl3_w_n14078_16(.douta(w_n14078_16[0]),.doutb(w_n14078_16[1]),.doutc(w_n14078_16[2]),.din(w_n14078_5[0]));
	jspl3 jspl3_w_n14078_17(.douta(w_n14078_17[0]),.doutb(w_n14078_17[1]),.doutc(w_n14078_17[2]),.din(w_n14078_5[1]));
	jspl3 jspl3_w_n14078_18(.douta(w_n14078_18[0]),.doutb(w_n14078_18[1]),.doutc(w_n14078_18[2]),.din(w_n14078_5[2]));
	jspl3 jspl3_w_n14078_19(.douta(w_n14078_19[0]),.doutb(w_n14078_19[1]),.doutc(w_n14078_19[2]),.din(w_n14078_6[0]));
	jspl3 jspl3_w_n14078_20(.douta(w_n14078_20[0]),.doutb(w_n14078_20[1]),.doutc(w_n14078_20[2]),.din(w_n14078_6[1]));
	jspl3 jspl3_w_n14078_21(.douta(w_n14078_21[0]),.doutb(w_n14078_21[1]),.doutc(w_n14078_21[2]),.din(w_n14078_6[2]));
	jspl3 jspl3_w_n14078_22(.douta(w_n14078_22[0]),.doutb(w_n14078_22[1]),.doutc(w_n14078_22[2]),.din(w_n14078_7[0]));
	jspl3 jspl3_w_n14078_23(.douta(w_n14078_23[0]),.doutb(w_n14078_23[1]),.doutc(w_n14078_23[2]),.din(w_n14078_7[1]));
	jspl3 jspl3_w_n14078_24(.douta(w_n14078_24[0]),.doutb(w_n14078_24[1]),.doutc(w_n14078_24[2]),.din(w_n14078_7[2]));
	jspl3 jspl3_w_n14078_25(.douta(w_n14078_25[0]),.doutb(w_n14078_25[1]),.doutc(w_n14078_25[2]),.din(w_n14078_8[0]));
	jspl3 jspl3_w_n14078_26(.douta(w_n14078_26[0]),.doutb(w_n14078_26[1]),.doutc(w_n14078_26[2]),.din(w_n14078_8[1]));
	jspl3 jspl3_w_n14078_27(.douta(w_n14078_27[0]),.doutb(w_n14078_27[1]),.doutc(w_n14078_27[2]),.din(w_n14078_8[2]));
	jspl3 jspl3_w_n14078_28(.douta(w_n14078_28[0]),.doutb(w_n14078_28[1]),.doutc(w_n14078_28[2]),.din(w_n14078_9[0]));
	jspl3 jspl3_w_n14078_29(.douta(w_n14078_29[0]),.doutb(w_n14078_29[1]),.doutc(w_n14078_29[2]),.din(w_n14078_9[1]));
	jspl3 jspl3_w_n14078_30(.douta(w_n14078_30[0]),.doutb(w_n14078_30[1]),.doutc(w_n14078_30[2]),.din(w_n14078_9[2]));
	jspl3 jspl3_w_n14078_31(.douta(w_n14078_31[0]),.doutb(w_n14078_31[1]),.doutc(w_n14078_31[2]),.din(w_n14078_10[0]));
	jspl3 jspl3_w_n14078_32(.douta(w_n14078_32[0]),.doutb(w_n14078_32[1]),.doutc(w_n14078_32[2]),.din(w_n14078_10[1]));
	jspl3 jspl3_w_n14078_33(.douta(w_n14078_33[0]),.doutb(w_n14078_33[1]),.doutc(w_n14078_33[2]),.din(w_n14078_10[2]));
	jspl3 jspl3_w_n14078_34(.douta(w_n14078_34[0]),.doutb(w_n14078_34[1]),.doutc(w_n14078_34[2]),.din(w_n14078_11[0]));
	jspl3 jspl3_w_n14078_35(.douta(w_n14078_35[0]),.doutb(w_n14078_35[1]),.doutc(w_n14078_35[2]),.din(w_n14078_11[1]));
	jspl3 jspl3_w_n14078_36(.douta(w_n14078_36[0]),.doutb(w_n14078_36[1]),.doutc(w_n14078_36[2]),.din(w_n14078_11[2]));
	jspl3 jspl3_w_n14078_37(.douta(w_n14078_37[0]),.doutb(w_n14078_37[1]),.doutc(w_n14078_37[2]),.din(w_n14078_12[0]));
	jspl3 jspl3_w_n14078_38(.douta(w_n14078_38[0]),.doutb(w_n14078_38[1]),.doutc(w_n14078_38[2]),.din(w_n14078_12[1]));
	jspl3 jspl3_w_n14078_39(.douta(w_n14078_39[0]),.doutb(w_n14078_39[1]),.doutc(w_n14078_39[2]),.din(w_n14078_12[2]));
	jspl3 jspl3_w_n14078_40(.douta(w_n14078_40[0]),.doutb(w_n14078_40[1]),.doutc(w_n14078_40[2]),.din(w_n14078_13[0]));
	jspl3 jspl3_w_n14078_41(.douta(w_n14078_41[0]),.doutb(w_n14078_41[1]),.doutc(w_n14078_41[2]),.din(w_n14078_13[1]));
	jspl jspl_w_n14078_42(.douta(w_n14078_42[0]),.doutb(w_n14078_42[1]),.din(w_n14078_13[2]));
	jspl3 jspl3_w_n14080_0(.douta(w_n14080_0[0]),.doutb(w_n14080_0[1]),.doutc(w_n14080_0[2]),.din(n14080));
	jspl3 jspl3_w_n14080_1(.douta(w_n14080_1[0]),.doutb(w_n14080_1[1]),.doutc(w_n14080_1[2]),.din(w_n14080_0[0]));
	jspl jspl_w_n14081_0(.douta(w_n14081_0[0]),.doutb(w_n14081_0[1]),.din(n14081));
	jspl3 jspl3_w_n14082_0(.douta(w_n14082_0[0]),.doutb(w_n14082_0[1]),.doutc(w_n14082_0[2]),.din(n14082));
	jspl jspl_w_n14083_0(.douta(w_n14083_0[0]),.doutb(w_n14083_0[1]),.din(n14083));
	jspl3 jspl3_w_n14085_0(.douta(w_n14085_0[0]),.doutb(w_n14085_0[1]),.doutc(w_n14085_0[2]),.din(n14085));
	jspl jspl_w_n14086_0(.douta(w_n14086_0[0]),.doutb(w_n14086_0[1]),.din(n14086));
	jspl3 jspl3_w_n14093_0(.douta(w_n14093_0[0]),.doutb(w_n14093_0[1]),.doutc(w_n14093_0[2]),.din(n14093));
	jspl jspl_w_n14094_0(.douta(w_n14094_0[0]),.doutb(w_n14094_0[1]),.din(n14094));
	jspl jspl_w_n14097_0(.douta(w_n14097_0[0]),.doutb(w_n14097_0[1]),.din(n14097));
	jspl3 jspl3_w_n14102_0(.douta(w_n14102_0[0]),.doutb(w_n14102_0[1]),.doutc(w_n14102_0[2]),.din(n14102));
	jspl3 jspl3_w_n14104_0(.douta(w_n14104_0[0]),.doutb(w_n14104_0[1]),.doutc(w_n14104_0[2]),.din(n14104));
	jspl jspl_w_n14105_0(.douta(w_n14105_0[0]),.doutb(w_n14105_0[1]),.din(n14105));
	jspl3 jspl3_w_n14109_0(.douta(w_n14109_0[0]),.doutb(w_n14109_0[1]),.doutc(w_n14109_0[2]),.din(n14109));
	jspl3 jspl3_w_n14112_0(.douta(w_n14112_0[0]),.doutb(w_n14112_0[1]),.doutc(w_n14112_0[2]),.din(n14112));
	jspl jspl_w_n14113_0(.douta(w_n14113_0[0]),.doutb(w_n14113_0[1]),.din(n14113));
	jspl3 jspl3_w_n14117_0(.douta(w_n14117_0[0]),.doutb(w_n14117_0[1]),.doutc(w_n14117_0[2]),.din(n14117));
	jspl3 jspl3_w_n14119_0(.douta(w_n14119_0[0]),.doutb(w_n14119_0[1]),.doutc(w_n14119_0[2]),.din(n14119));
	jspl jspl_w_n14120_0(.douta(w_n14120_0[0]),.doutb(w_n14120_0[1]),.din(n14120));
	jspl3 jspl3_w_n14124_0(.douta(w_n14124_0[0]),.doutb(w_n14124_0[1]),.doutc(w_n14124_0[2]),.din(n14124));
	jspl3 jspl3_w_n14126_0(.douta(w_n14126_0[0]),.doutb(w_n14126_0[1]),.doutc(w_n14126_0[2]),.din(n14126));
	jspl jspl_w_n14127_0(.douta(w_n14127_0[0]),.doutb(w_n14127_0[1]),.din(n14127));
	jspl3 jspl3_w_n14131_0(.douta(w_n14131_0[0]),.doutb(w_n14131_0[1]),.doutc(w_n14131_0[2]),.din(n14131));
	jspl3 jspl3_w_n14133_0(.douta(w_n14133_0[0]),.doutb(w_n14133_0[1]),.doutc(w_n14133_0[2]),.din(n14133));
	jspl jspl_w_n14134_0(.douta(w_n14134_0[0]),.doutb(w_n14134_0[1]),.din(n14134));
	jspl3 jspl3_w_n14138_0(.douta(w_n14138_0[0]),.doutb(w_n14138_0[1]),.doutc(w_n14138_0[2]),.din(n14138));
	jspl3 jspl3_w_n14141_0(.douta(w_n14141_0[0]),.doutb(w_n14141_0[1]),.doutc(w_n14141_0[2]),.din(n14141));
	jspl jspl_w_n14142_0(.douta(w_n14142_0[0]),.doutb(w_n14142_0[1]),.din(n14142));
	jspl3 jspl3_w_n14146_0(.douta(w_n14146_0[0]),.doutb(w_n14146_0[1]),.doutc(w_n14146_0[2]),.din(n14146));
	jspl3 jspl3_w_n14148_0(.douta(w_n14148_0[0]),.doutb(w_n14148_0[1]),.doutc(w_n14148_0[2]),.din(n14148));
	jspl jspl_w_n14149_0(.douta(w_n14149_0[0]),.doutb(w_n14149_0[1]),.din(n14149));
	jspl3 jspl3_w_n14153_0(.douta(w_n14153_0[0]),.doutb(w_n14153_0[1]),.doutc(w_n14153_0[2]),.din(n14153));
	jspl3 jspl3_w_n14156_0(.douta(w_n14156_0[0]),.doutb(w_n14156_0[1]),.doutc(w_n14156_0[2]),.din(n14156));
	jspl jspl_w_n14157_0(.douta(w_n14157_0[0]),.doutb(w_n14157_0[1]),.din(n14157));
	jspl3 jspl3_w_n14161_0(.douta(w_n14161_0[0]),.doutb(w_n14161_0[1]),.doutc(w_n14161_0[2]),.din(n14161));
	jspl3 jspl3_w_n14163_0(.douta(w_n14163_0[0]),.doutb(w_n14163_0[1]),.doutc(w_n14163_0[2]),.din(n14163));
	jspl jspl_w_n14164_0(.douta(w_n14164_0[0]),.doutb(w_n14164_0[1]),.din(n14164));
	jspl3 jspl3_w_n14168_0(.douta(w_n14168_0[0]),.doutb(w_n14168_0[1]),.doutc(w_n14168_0[2]),.din(n14168));
	jspl3 jspl3_w_n14171_0(.douta(w_n14171_0[0]),.doutb(w_n14171_0[1]),.doutc(w_n14171_0[2]),.din(n14171));
	jspl jspl_w_n14172_0(.douta(w_n14172_0[0]),.doutb(w_n14172_0[1]),.din(n14172));
	jspl3 jspl3_w_n14176_0(.douta(w_n14176_0[0]),.doutb(w_n14176_0[1]),.doutc(w_n14176_0[2]),.din(n14176));
	jspl3 jspl3_w_n14178_0(.douta(w_n14178_0[0]),.doutb(w_n14178_0[1]),.doutc(w_n14178_0[2]),.din(n14178));
	jspl jspl_w_n14179_0(.douta(w_n14179_0[0]),.doutb(w_n14179_0[1]),.din(n14179));
	jspl3 jspl3_w_n14183_0(.douta(w_n14183_0[0]),.doutb(w_n14183_0[1]),.doutc(w_n14183_0[2]),.din(n14183));
	jspl3 jspl3_w_n14186_0(.douta(w_n14186_0[0]),.doutb(w_n14186_0[1]),.doutc(w_n14186_0[2]),.din(n14186));
	jspl jspl_w_n14187_0(.douta(w_n14187_0[0]),.doutb(w_n14187_0[1]),.din(n14187));
	jspl3 jspl3_w_n14191_0(.douta(w_n14191_0[0]),.doutb(w_n14191_0[1]),.doutc(w_n14191_0[2]),.din(n14191));
	jspl3 jspl3_w_n14193_0(.douta(w_n14193_0[0]),.doutb(w_n14193_0[1]),.doutc(w_n14193_0[2]),.din(n14193));
	jspl jspl_w_n14194_0(.douta(w_n14194_0[0]),.doutb(w_n14194_0[1]),.din(n14194));
	jspl3 jspl3_w_n14198_0(.douta(w_n14198_0[0]),.doutb(w_n14198_0[1]),.doutc(w_n14198_0[2]),.din(n14198));
	jspl3 jspl3_w_n14200_0(.douta(w_n14200_0[0]),.doutb(w_n14200_0[1]),.doutc(w_n14200_0[2]),.din(n14200));
	jspl jspl_w_n14201_0(.douta(w_n14201_0[0]),.doutb(w_n14201_0[1]),.din(n14201));
	jspl3 jspl3_w_n14205_0(.douta(w_n14205_0[0]),.doutb(w_n14205_0[1]),.doutc(w_n14205_0[2]),.din(n14205));
	jspl3 jspl3_w_n14207_0(.douta(w_n14207_0[0]),.doutb(w_n14207_0[1]),.doutc(w_n14207_0[2]),.din(n14207));
	jspl jspl_w_n14208_0(.douta(w_n14208_0[0]),.doutb(w_n14208_0[1]),.din(n14208));
	jspl3 jspl3_w_n14212_0(.douta(w_n14212_0[0]),.doutb(w_n14212_0[1]),.doutc(w_n14212_0[2]),.din(n14212));
	jspl3 jspl3_w_n14215_0(.douta(w_n14215_0[0]),.doutb(w_n14215_0[1]),.doutc(w_n14215_0[2]),.din(n14215));
	jspl jspl_w_n14216_0(.douta(w_n14216_0[0]),.doutb(w_n14216_0[1]),.din(n14216));
	jspl3 jspl3_w_n14220_0(.douta(w_n14220_0[0]),.doutb(w_n14220_0[1]),.doutc(w_n14220_0[2]),.din(n14220));
	jspl3 jspl3_w_n14222_0(.douta(w_n14222_0[0]),.doutb(w_n14222_0[1]),.doutc(w_n14222_0[2]),.din(n14222));
	jspl jspl_w_n14223_0(.douta(w_n14223_0[0]),.doutb(w_n14223_0[1]),.din(n14223));
	jspl3 jspl3_w_n14227_0(.douta(w_n14227_0[0]),.doutb(w_n14227_0[1]),.doutc(w_n14227_0[2]),.din(n14227));
	jspl3 jspl3_w_n14230_0(.douta(w_n14230_0[0]),.doutb(w_n14230_0[1]),.doutc(w_n14230_0[2]),.din(n14230));
	jspl jspl_w_n14231_0(.douta(w_n14231_0[0]),.doutb(w_n14231_0[1]),.din(n14231));
	jspl3 jspl3_w_n14235_0(.douta(w_n14235_0[0]),.doutb(w_n14235_0[1]),.doutc(w_n14235_0[2]),.din(n14235));
	jspl3 jspl3_w_n14237_0(.douta(w_n14237_0[0]),.doutb(w_n14237_0[1]),.doutc(w_n14237_0[2]),.din(n14237));
	jspl jspl_w_n14238_0(.douta(w_n14238_0[0]),.doutb(w_n14238_0[1]),.din(n14238));
	jspl3 jspl3_w_n14242_0(.douta(w_n14242_0[0]),.doutb(w_n14242_0[1]),.doutc(w_n14242_0[2]),.din(n14242));
	jspl3 jspl3_w_n14244_0(.douta(w_n14244_0[0]),.doutb(w_n14244_0[1]),.doutc(w_n14244_0[2]),.din(n14244));
	jspl jspl_w_n14245_0(.douta(w_n14245_0[0]),.doutb(w_n14245_0[1]),.din(n14245));
	jspl3 jspl3_w_n14249_0(.douta(w_n14249_0[0]),.doutb(w_n14249_0[1]),.doutc(w_n14249_0[2]),.din(n14249));
	jspl3 jspl3_w_n14251_0(.douta(w_n14251_0[0]),.doutb(w_n14251_0[1]),.doutc(w_n14251_0[2]),.din(n14251));
	jspl jspl_w_n14252_0(.douta(w_n14252_0[0]),.doutb(w_n14252_0[1]),.din(n14252));
	jspl3 jspl3_w_n14256_0(.douta(w_n14256_0[0]),.doutb(w_n14256_0[1]),.doutc(w_n14256_0[2]),.din(n14256));
	jspl3 jspl3_w_n14259_0(.douta(w_n14259_0[0]),.doutb(w_n14259_0[1]),.doutc(w_n14259_0[2]),.din(n14259));
	jspl jspl_w_n14260_0(.douta(w_n14260_0[0]),.doutb(w_n14260_0[1]),.din(n14260));
	jspl3 jspl3_w_n14264_0(.douta(w_n14264_0[0]),.doutb(w_n14264_0[1]),.doutc(w_n14264_0[2]),.din(n14264));
	jspl3 jspl3_w_n14266_0(.douta(w_n14266_0[0]),.doutb(w_n14266_0[1]),.doutc(w_n14266_0[2]),.din(n14266));
	jspl jspl_w_n14267_0(.douta(w_n14267_0[0]),.doutb(w_n14267_0[1]),.din(n14267));
	jspl jspl_w_n14271_0(.douta(w_n14271_0[0]),.doutb(w_n14271_0[1]),.din(n14271));
	jspl3 jspl3_w_n14273_0(.douta(w_n14273_0[0]),.doutb(w_n14273_0[1]),.doutc(w_n14273_0[2]),.din(n14273));
	jspl jspl_w_n14274_0(.douta(w_n14274_0[0]),.doutb(w_n14274_0[1]),.din(n14274));
	jspl3 jspl3_w_n14278_0(.douta(w_n14278_0[0]),.doutb(w_n14278_0[1]),.doutc(w_n14278_0[2]),.din(n14278));
	jspl3 jspl3_w_n14280_0(.douta(w_n14280_0[0]),.doutb(w_n14280_0[1]),.doutc(w_n14280_0[2]),.din(n14280));
	jspl jspl_w_n14281_0(.douta(w_n14281_0[0]),.doutb(w_n14281_0[1]),.din(n14281));
	jspl3 jspl3_w_n14285_0(.douta(w_n14285_0[0]),.doutb(w_n14285_0[1]),.doutc(w_n14285_0[2]),.din(n14285));
	jspl3 jspl3_w_n14287_0(.douta(w_n14287_0[0]),.doutb(w_n14287_0[1]),.doutc(w_n14287_0[2]),.din(n14287));
	jspl jspl_w_n14288_0(.douta(w_n14288_0[0]),.doutb(w_n14288_0[1]),.din(n14288));
	jspl3 jspl3_w_n14292_0(.douta(w_n14292_0[0]),.doutb(w_n14292_0[1]),.doutc(w_n14292_0[2]),.din(n14292));
	jspl3 jspl3_w_n14295_0(.douta(w_n14295_0[0]),.doutb(w_n14295_0[1]),.doutc(w_n14295_0[2]),.din(n14295));
	jspl jspl_w_n14296_0(.douta(w_n14296_0[0]),.doutb(w_n14296_0[1]),.din(n14296));
	jspl3 jspl3_w_n14299_0(.douta(w_n14299_0[0]),.doutb(w_n14299_0[1]),.doutc(w_n14299_0[2]),.din(n14299));
	jspl3 jspl3_w_n14303_0(.douta(w_n14303_0[0]),.doutb(w_n14303_0[1]),.doutc(w_n14303_0[2]),.din(n14303));
	jspl jspl_w_n14304_0(.douta(w_n14304_0[0]),.doutb(w_n14304_0[1]),.din(n14304));
	jspl3 jspl3_w_n14308_0(.douta(w_n14308_0[0]),.doutb(w_n14308_0[1]),.doutc(w_n14308_0[2]),.din(n14308));
	jspl3 jspl3_w_n14310_0(.douta(w_n14310_0[0]),.doutb(w_n14310_0[1]),.doutc(w_n14310_0[2]),.din(n14310));
	jspl jspl_w_n14311_0(.douta(w_n14311_0[0]),.doutb(w_n14311_0[1]),.din(n14311));
	jspl3 jspl3_w_n14315_0(.douta(w_n14315_0[0]),.doutb(w_n14315_0[1]),.doutc(w_n14315_0[2]),.din(n14315));
	jspl3 jspl3_w_n14318_0(.douta(w_n14318_0[0]),.doutb(w_n14318_0[1]),.doutc(w_n14318_0[2]),.din(n14318));
	jspl jspl_w_n14319_0(.douta(w_n14319_0[0]),.doutb(w_n14319_0[1]),.din(n14319));
	jspl3 jspl3_w_n14323_0(.douta(w_n14323_0[0]),.doutb(w_n14323_0[1]),.doutc(w_n14323_0[2]),.din(n14323));
	jspl3 jspl3_w_n14325_0(.douta(w_n14325_0[0]),.doutb(w_n14325_0[1]),.doutc(w_n14325_0[2]),.din(n14325));
	jspl jspl_w_n14326_0(.douta(w_n14326_0[0]),.doutb(w_n14326_0[1]),.din(n14326));
	jspl3 jspl3_w_n14330_0(.douta(w_n14330_0[0]),.doutb(w_n14330_0[1]),.doutc(w_n14330_0[2]),.din(n14330));
	jspl3 jspl3_w_n14333_0(.douta(w_n14333_0[0]),.doutb(w_n14333_0[1]),.doutc(w_n14333_0[2]),.din(n14333));
	jspl jspl_w_n14334_0(.douta(w_n14334_0[0]),.doutb(w_n14334_0[1]),.din(n14334));
	jspl3 jspl3_w_n14338_0(.douta(w_n14338_0[0]),.doutb(w_n14338_0[1]),.doutc(w_n14338_0[2]),.din(n14338));
	jspl3 jspl3_w_n14340_0(.douta(w_n14340_0[0]),.doutb(w_n14340_0[1]),.doutc(w_n14340_0[2]),.din(n14340));
	jspl jspl_w_n14341_0(.douta(w_n14341_0[0]),.doutb(w_n14341_0[1]),.din(n14341));
	jspl3 jspl3_w_n14345_0(.douta(w_n14345_0[0]),.doutb(w_n14345_0[1]),.doutc(w_n14345_0[2]),.din(n14345));
	jspl3 jspl3_w_n14347_0(.douta(w_n14347_0[0]),.doutb(w_n14347_0[1]),.doutc(w_n14347_0[2]),.din(n14347));
	jspl jspl_w_n14348_0(.douta(w_n14348_0[0]),.doutb(w_n14348_0[1]),.din(n14348));
	jspl3 jspl3_w_n14352_0(.douta(w_n14352_0[0]),.doutb(w_n14352_0[1]),.doutc(w_n14352_0[2]),.din(n14352));
	jspl3 jspl3_w_n14354_0(.douta(w_n14354_0[0]),.doutb(w_n14354_0[1]),.doutc(w_n14354_0[2]),.din(n14354));
	jspl jspl_w_n14355_0(.douta(w_n14355_0[0]),.doutb(w_n14355_0[1]),.din(n14355));
	jspl3 jspl3_w_n14359_0(.douta(w_n14359_0[0]),.doutb(w_n14359_0[1]),.doutc(w_n14359_0[2]),.din(n14359));
	jspl3 jspl3_w_n14362_0(.douta(w_n14362_0[0]),.doutb(w_n14362_0[1]),.doutc(w_n14362_0[2]),.din(n14362));
	jspl jspl_w_n14363_0(.douta(w_n14363_0[0]),.doutb(w_n14363_0[1]),.din(n14363));
	jspl3 jspl3_w_n14367_0(.douta(w_n14367_0[0]),.doutb(w_n14367_0[1]),.doutc(w_n14367_0[2]),.din(n14367));
	jspl3 jspl3_w_n14369_0(.douta(w_n14369_0[0]),.doutb(w_n14369_0[1]),.doutc(w_n14369_0[2]),.din(n14369));
	jspl jspl_w_n14370_0(.douta(w_n14370_0[0]),.doutb(w_n14370_0[1]),.din(n14370));
	jspl3 jspl3_w_n14374_0(.douta(w_n14374_0[0]),.doutb(w_n14374_0[1]),.doutc(w_n14374_0[2]),.din(n14374));
	jspl3 jspl3_w_n14377_0(.douta(w_n14377_0[0]),.doutb(w_n14377_0[1]),.doutc(w_n14377_0[2]),.din(n14377));
	jspl jspl_w_n14378_0(.douta(w_n14378_0[0]),.doutb(w_n14378_0[1]),.din(n14378));
	jspl3 jspl3_w_n14382_0(.douta(w_n14382_0[0]),.doutb(w_n14382_0[1]),.doutc(w_n14382_0[2]),.din(n14382));
	jspl3 jspl3_w_n14384_0(.douta(w_n14384_0[0]),.doutb(w_n14384_0[1]),.doutc(w_n14384_0[2]),.din(n14384));
	jspl jspl_w_n14385_0(.douta(w_n14385_0[0]),.doutb(w_n14385_0[1]),.din(n14385));
	jspl3 jspl3_w_n14389_0(.douta(w_n14389_0[0]),.doutb(w_n14389_0[1]),.doutc(w_n14389_0[2]),.din(n14389));
	jspl3 jspl3_w_n14392_0(.douta(w_n14392_0[0]),.doutb(w_n14392_0[1]),.doutc(w_n14392_0[2]),.din(n14392));
	jspl jspl_w_n14393_0(.douta(w_n14393_0[0]),.doutb(w_n14393_0[1]),.din(n14393));
	jspl3 jspl3_w_n14397_0(.douta(w_n14397_0[0]),.doutb(w_n14397_0[1]),.doutc(w_n14397_0[2]),.din(n14397));
	jspl3 jspl3_w_n14399_0(.douta(w_n14399_0[0]),.doutb(w_n14399_0[1]),.doutc(w_n14399_0[2]),.din(n14399));
	jspl jspl_w_n14400_0(.douta(w_n14400_0[0]),.doutb(w_n14400_0[1]),.din(n14400));
	jspl3 jspl3_w_n14404_0(.douta(w_n14404_0[0]),.doutb(w_n14404_0[1]),.doutc(w_n14404_0[2]),.din(n14404));
	jspl3 jspl3_w_n14407_0(.douta(w_n14407_0[0]),.doutb(w_n14407_0[1]),.doutc(w_n14407_0[2]),.din(n14407));
	jspl jspl_w_n14408_0(.douta(w_n14408_0[0]),.doutb(w_n14408_0[1]),.din(n14408));
	jspl3 jspl3_w_n14412_0(.douta(w_n14412_0[0]),.doutb(w_n14412_0[1]),.doutc(w_n14412_0[2]),.din(n14412));
	jspl3 jspl3_w_n14415_0(.douta(w_n14415_0[0]),.doutb(w_n14415_0[1]),.doutc(w_n14415_0[2]),.din(n14415));
	jspl jspl_w_n14416_0(.douta(w_n14416_0[0]),.doutb(w_n14416_0[1]),.din(n14416));
	jspl jspl_w_n14420_0(.douta(w_n14420_0[0]),.doutb(w_n14420_0[1]),.din(n14420));
	jspl jspl_w_n14421_0(.douta(w_n14421_0[0]),.doutb(w_n14421_0[1]),.din(n14421));
	jspl3 jspl3_w_n14423_0(.douta(w_n14423_0[0]),.doutb(w_n14423_0[1]),.doutc(w_n14423_0[2]),.din(n14423));
	jspl jspl_w_n14423_1(.douta(w_n14423_1[0]),.doutb(w_n14423_1[1]),.din(w_n14423_0[0]));
	jspl3 jspl3_w_n14426_0(.douta(w_n14426_0[0]),.doutb(w_n14426_0[1]),.doutc(w_n14426_0[2]),.din(n14426));
	jspl3 jspl3_w_n14426_1(.douta(w_n14426_1[0]),.doutb(w_n14426_1[1]),.doutc(w_n14426_1[2]),.din(w_n14426_0[0]));
	jspl jspl_w_n14427_0(.douta(w_n14427_0[0]),.doutb(w_n14427_0[1]),.din(n14427));
	jspl jspl_w_n14430_0(.douta(w_n14430_0[0]),.doutb(w_n14430_0[1]),.din(n14430));
	jspl jspl_w_n14432_0(.douta(w_n14432_0[0]),.doutb(w_n14432_0[1]),.din(n14432));
	jspl jspl_w_n14437_0(.douta(w_n14437_0[0]),.doutb(w_n14437_0[1]),.din(n14437));
	jspl jspl_w_n14438_0(.douta(w_n14438_0[0]),.doutb(w_n14438_0[1]),.din(n14438));
	jspl3 jspl3_w_n14443_0(.douta(w_n14443_0[0]),.doutb(w_n14443_0[1]),.doutc(w_n14443_0[2]),.din(n14443));
	jspl jspl_w_n14443_1(.douta(w_n14443_1[0]),.doutb(w_n14443_1[1]),.din(w_n14443_0[0]));
	jspl jspl_w_n14444_0(.douta(w_n14444_0[0]),.doutb(w_n14444_0[1]),.din(n14444));
	jspl3 jspl3_w_n14445_0(.douta(w_n14445_0[0]),.doutb(w_n14445_0[1]),.doutc(w_n14445_0[2]),.din(n14445));
	jspl jspl_w_n14446_0(.douta(w_n14446_0[0]),.doutb(w_n14446_0[1]),.din(n14446));
	jspl3 jspl3_w_n14448_0(.douta(w_n14448_0[0]),.doutb(w_n14448_0[1]),.doutc(w_n14448_0[2]),.din(n14448));
	jspl jspl_w_n14449_0(.douta(w_n14449_0[0]),.doutb(w_n14449_0[1]),.din(n14449));
	jspl jspl_w_n14454_0(.douta(w_n14454_0[0]),.doutb(w_n14454_0[1]),.din(n14454));
	jspl jspl_w_n14506_0(.douta(w_n14506_0[0]),.doutb(w_n14506_0[1]),.din(n14506));
	jspl jspl_w_n14594_0(.douta(w_n14594_0[0]),.doutb(w_n14594_0[1]),.din(n14594));
	jspl jspl_w_n14671_0(.douta(w_n14671_0[0]),.doutb(w_n14671_0[1]),.din(n14671));
	jspl jspl_w_n14672_0(.douta(w_n14672_0[0]),.doutb(w_n14672_0[1]),.din(n14672));
	jspl3 jspl3_w_n14674_0(.douta(w_n14674_0[0]),.doutb(w_n14674_0[1]),.doutc(w_n14674_0[2]),.din(n14674));
	jspl3 jspl3_w_n14674_1(.douta(w_n14674_1[0]),.doutb(w_n14674_1[1]),.doutc(w_n14674_1[2]),.din(w_n14674_0[0]));
	jspl3 jspl3_w_n14674_2(.douta(w_n14674_2[0]),.doutb(w_n14674_2[1]),.doutc(w_n14674_2[2]),.din(w_n14674_0[1]));
	jspl3 jspl3_w_n14674_3(.douta(w_n14674_3[0]),.doutb(w_n14674_3[1]),.doutc(w_n14674_3[2]),.din(w_n14674_0[2]));
	jspl3 jspl3_w_n14674_4(.douta(w_n14674_4[0]),.doutb(w_n14674_4[1]),.doutc(w_n14674_4[2]),.din(w_n14674_1[0]));
	jspl3 jspl3_w_n14674_5(.douta(w_n14674_5[0]),.doutb(w_n14674_5[1]),.doutc(w_n14674_5[2]),.din(w_n14674_1[1]));
	jspl3 jspl3_w_n14674_6(.douta(w_n14674_6[0]),.doutb(w_n14674_6[1]),.doutc(w_n14674_6[2]),.din(w_n14674_1[2]));
	jspl3 jspl3_w_n14674_7(.douta(w_n14674_7[0]),.doutb(w_n14674_7[1]),.doutc(w_n14674_7[2]),.din(w_n14674_2[0]));
	jspl3 jspl3_w_n14674_8(.douta(w_n14674_8[0]),.doutb(w_n14674_8[1]),.doutc(w_n14674_8[2]),.din(w_n14674_2[1]));
	jspl3 jspl3_w_n14674_9(.douta(w_n14674_9[0]),.doutb(w_n14674_9[1]),.doutc(w_n14674_9[2]),.din(w_n14674_2[2]));
	jspl3 jspl3_w_n14674_10(.douta(w_n14674_10[0]),.doutb(w_n14674_10[1]),.doutc(w_n14674_10[2]),.din(w_n14674_3[0]));
	jspl3 jspl3_w_n14674_11(.douta(w_n14674_11[0]),.doutb(w_n14674_11[1]),.doutc(w_n14674_11[2]),.din(w_n14674_3[1]));
	jspl3 jspl3_w_n14674_12(.douta(w_n14674_12[0]),.doutb(w_n14674_12[1]),.doutc(w_n14674_12[2]),.din(w_n14674_3[2]));
	jspl3 jspl3_w_n14674_13(.douta(w_n14674_13[0]),.doutb(w_n14674_13[1]),.doutc(w_n14674_13[2]),.din(w_n14674_4[0]));
	jspl3 jspl3_w_n14674_14(.douta(w_n14674_14[0]),.doutb(w_n14674_14[1]),.doutc(w_n14674_14[2]),.din(w_n14674_4[1]));
	jspl3 jspl3_w_n14674_15(.douta(w_n14674_15[0]),.doutb(w_n14674_15[1]),.doutc(w_n14674_15[2]),.din(w_n14674_4[2]));
	jspl3 jspl3_w_n14674_16(.douta(w_n14674_16[0]),.doutb(w_n14674_16[1]),.doutc(w_n14674_16[2]),.din(w_n14674_5[0]));
	jspl3 jspl3_w_n14674_17(.douta(w_n14674_17[0]),.doutb(w_n14674_17[1]),.doutc(w_n14674_17[2]),.din(w_n14674_5[1]));
	jspl3 jspl3_w_n14674_18(.douta(w_n14674_18[0]),.doutb(w_n14674_18[1]),.doutc(w_n14674_18[2]),.din(w_n14674_5[2]));
	jspl3 jspl3_w_n14674_19(.douta(w_n14674_19[0]),.doutb(w_n14674_19[1]),.doutc(w_n14674_19[2]),.din(w_n14674_6[0]));
	jspl jspl_w_n14674_20(.douta(w_n14674_20[0]),.doutb(w_n14674_20[1]),.din(w_n14674_6[1]));
	jspl3 jspl3_w_n14678_0(.douta(w_n14678_0[0]),.doutb(w_n14678_0[1]),.doutc(w_n14678_0[2]),.din(n14678));
	jspl jspl_w_n14679_0(.douta(w_n14679_0[0]),.doutb(w_n14679_0[1]),.din(n14679));
	jspl jspl_w_n14681_0(.douta(w_n14681_0[0]),.doutb(w_n14681_0[1]),.din(n14681));
	jspl jspl_w_n14686_0(.douta(w_n14686_0[0]),.doutb(w_n14686_0[1]),.din(n14686));
	jspl jspl_w_n14687_0(.douta(w_n14687_0[0]),.doutb(w_n14687_0[1]),.din(n14687));
	jspl3 jspl3_w_n14689_0(.douta(w_n14689_0[0]),.doutb(w_n14689_0[1]),.doutc(w_n14689_0[2]),.din(n14689));
	jspl jspl_w_n14690_0(.douta(w_n14690_0[0]),.doutb(w_n14690_0[1]),.din(n14690));
	jspl jspl_w_n14694_0(.douta(w_n14694_0[0]),.doutb(w_n14694_0[1]),.din(n14694));
	jspl3 jspl3_w_n14696_0(.douta(w_n14696_0[0]),.doutb(w_n14696_0[1]),.doutc(w_n14696_0[2]),.din(n14696));
	jspl jspl_w_n14697_0(.douta(w_n14697_0[0]),.doutb(w_n14697_0[1]),.din(n14697));
	jspl jspl_w_n14701_0(.douta(w_n14701_0[0]),.doutb(w_n14701_0[1]),.din(n14701));
	jspl jspl_w_n14702_0(.douta(w_n14702_0[0]),.doutb(w_n14702_0[1]),.din(n14702));
	jspl3 jspl3_w_n14704_0(.douta(w_n14704_0[0]),.doutb(w_n14704_0[1]),.doutc(w_n14704_0[2]),.din(n14704));
	jspl jspl_w_n14705_0(.douta(w_n14705_0[0]),.doutb(w_n14705_0[1]),.din(n14705));
	jspl jspl_w_n14709_0(.douta(w_n14709_0[0]),.doutb(w_n14709_0[1]),.din(n14709));
	jspl3 jspl3_w_n14711_0(.douta(w_n14711_0[0]),.doutb(w_n14711_0[1]),.doutc(w_n14711_0[2]),.din(n14711));
	jspl jspl_w_n14712_0(.douta(w_n14712_0[0]),.doutb(w_n14712_0[1]),.din(n14712));
	jspl jspl_w_n14716_0(.douta(w_n14716_0[0]),.doutb(w_n14716_0[1]),.din(n14716));
	jspl jspl_w_n14717_0(.douta(w_n14717_0[0]),.doutb(w_n14717_0[1]),.din(n14717));
	jspl3 jspl3_w_n14719_0(.douta(w_n14719_0[0]),.doutb(w_n14719_0[1]),.doutc(w_n14719_0[2]),.din(n14719));
	jspl jspl_w_n14720_0(.douta(w_n14720_0[0]),.doutb(w_n14720_0[1]),.din(n14720));
	jspl jspl_w_n14724_0(.douta(w_n14724_0[0]),.doutb(w_n14724_0[1]),.din(n14724));
	jspl jspl_w_n14725_0(.douta(w_n14725_0[0]),.doutb(w_n14725_0[1]),.din(n14725));
	jspl3 jspl3_w_n14727_0(.douta(w_n14727_0[0]),.doutb(w_n14727_0[1]),.doutc(w_n14727_0[2]),.din(n14727));
	jspl jspl_w_n14728_0(.douta(w_n14728_0[0]),.doutb(w_n14728_0[1]),.din(n14728));
	jspl jspl_w_n14732_0(.douta(w_n14732_0[0]),.doutb(w_n14732_0[1]),.din(n14732));
	jspl jspl_w_n14733_0(.douta(w_n14733_0[0]),.doutb(w_n14733_0[1]),.din(n14733));
	jspl3 jspl3_w_n14735_0(.douta(w_n14735_0[0]),.doutb(w_n14735_0[1]),.doutc(w_n14735_0[2]),.din(n14735));
	jspl jspl_w_n14736_0(.douta(w_n14736_0[0]),.doutb(w_n14736_0[1]),.din(n14736));
	jspl jspl_w_n14740_0(.douta(w_n14740_0[0]),.doutb(w_n14740_0[1]),.din(n14740));
	jspl3 jspl3_w_n14742_0(.douta(w_n14742_0[0]),.doutb(w_n14742_0[1]),.doutc(w_n14742_0[2]),.din(n14742));
	jspl jspl_w_n14743_0(.douta(w_n14743_0[0]),.doutb(w_n14743_0[1]),.din(n14743));
	jspl jspl_w_n14747_0(.douta(w_n14747_0[0]),.doutb(w_n14747_0[1]),.din(n14747));
	jspl jspl_w_n14748_0(.douta(w_n14748_0[0]),.doutb(w_n14748_0[1]),.din(n14748));
	jspl3 jspl3_w_n14750_0(.douta(w_n14750_0[0]),.doutb(w_n14750_0[1]),.doutc(w_n14750_0[2]),.din(n14750));
	jspl jspl_w_n14751_0(.douta(w_n14751_0[0]),.doutb(w_n14751_0[1]),.din(n14751));
	jspl jspl_w_n14755_0(.douta(w_n14755_0[0]),.doutb(w_n14755_0[1]),.din(n14755));
	jspl3 jspl3_w_n14757_0(.douta(w_n14757_0[0]),.doutb(w_n14757_0[1]),.doutc(w_n14757_0[2]),.din(n14757));
	jspl jspl_w_n14758_0(.douta(w_n14758_0[0]),.doutb(w_n14758_0[1]),.din(n14758));
	jspl jspl_w_n14762_0(.douta(w_n14762_0[0]),.doutb(w_n14762_0[1]),.din(n14762));
	jspl jspl_w_n14763_0(.douta(w_n14763_0[0]),.doutb(w_n14763_0[1]),.din(n14763));
	jspl3 jspl3_w_n14765_0(.douta(w_n14765_0[0]),.doutb(w_n14765_0[1]),.doutc(w_n14765_0[2]),.din(n14765));
	jspl jspl_w_n14766_0(.douta(w_n14766_0[0]),.doutb(w_n14766_0[1]),.din(n14766));
	jspl jspl_w_n14770_0(.douta(w_n14770_0[0]),.doutb(w_n14770_0[1]),.din(n14770));
	jspl3 jspl3_w_n14772_0(.douta(w_n14772_0[0]),.doutb(w_n14772_0[1]),.doutc(w_n14772_0[2]),.din(n14772));
	jspl jspl_w_n14773_0(.douta(w_n14773_0[0]),.doutb(w_n14773_0[1]),.din(n14773));
	jspl jspl_w_n14777_0(.douta(w_n14777_0[0]),.doutb(w_n14777_0[1]),.din(n14777));
	jspl jspl_w_n14778_0(.douta(w_n14778_0[0]),.doutb(w_n14778_0[1]),.din(n14778));
	jspl3 jspl3_w_n14780_0(.douta(w_n14780_0[0]),.doutb(w_n14780_0[1]),.doutc(w_n14780_0[2]),.din(n14780));
	jspl jspl_w_n14781_0(.douta(w_n14781_0[0]),.doutb(w_n14781_0[1]),.din(n14781));
	jspl jspl_w_n14785_0(.douta(w_n14785_0[0]),.doutb(w_n14785_0[1]),.din(n14785));
	jspl3 jspl3_w_n14787_0(.douta(w_n14787_0[0]),.doutb(w_n14787_0[1]),.doutc(w_n14787_0[2]),.din(n14787));
	jspl jspl_w_n14788_0(.douta(w_n14788_0[0]),.doutb(w_n14788_0[1]),.din(n14788));
	jspl jspl_w_n14792_0(.douta(w_n14792_0[0]),.doutb(w_n14792_0[1]),.din(n14792));
	jspl jspl_w_n14793_0(.douta(w_n14793_0[0]),.doutb(w_n14793_0[1]),.din(n14793));
	jspl3 jspl3_w_n14795_0(.douta(w_n14795_0[0]),.doutb(w_n14795_0[1]),.doutc(w_n14795_0[2]),.din(n14795));
	jspl jspl_w_n14796_0(.douta(w_n14796_0[0]),.doutb(w_n14796_0[1]),.din(n14796));
	jspl jspl_w_n14800_0(.douta(w_n14800_0[0]),.doutb(w_n14800_0[1]),.din(n14800));
	jspl jspl_w_n14801_0(.douta(w_n14801_0[0]),.doutb(w_n14801_0[1]),.din(n14801));
	jspl3 jspl3_w_n14803_0(.douta(w_n14803_0[0]),.doutb(w_n14803_0[1]),.doutc(w_n14803_0[2]),.din(n14803));
	jspl jspl_w_n14804_0(.douta(w_n14804_0[0]),.doutb(w_n14804_0[1]),.din(n14804));
	jspl jspl_w_n14808_0(.douta(w_n14808_0[0]),.doutb(w_n14808_0[1]),.din(n14808));
	jspl jspl_w_n14809_0(.douta(w_n14809_0[0]),.doutb(w_n14809_0[1]),.din(n14809));
	jspl3 jspl3_w_n14811_0(.douta(w_n14811_0[0]),.doutb(w_n14811_0[1]),.doutc(w_n14811_0[2]),.din(n14811));
	jspl jspl_w_n14812_0(.douta(w_n14812_0[0]),.doutb(w_n14812_0[1]),.din(n14812));
	jspl jspl_w_n14816_0(.douta(w_n14816_0[0]),.doutb(w_n14816_0[1]),.din(n14816));
	jspl3 jspl3_w_n14818_0(.douta(w_n14818_0[0]),.doutb(w_n14818_0[1]),.doutc(w_n14818_0[2]),.din(n14818));
	jspl jspl_w_n14819_0(.douta(w_n14819_0[0]),.doutb(w_n14819_0[1]),.din(n14819));
	jspl jspl_w_n14823_0(.douta(w_n14823_0[0]),.doutb(w_n14823_0[1]),.din(n14823));
	jspl jspl_w_n14824_0(.douta(w_n14824_0[0]),.doutb(w_n14824_0[1]),.din(n14824));
	jspl3 jspl3_w_n14826_0(.douta(w_n14826_0[0]),.doutb(w_n14826_0[1]),.doutc(w_n14826_0[2]),.din(n14826));
	jspl jspl_w_n14827_0(.douta(w_n14827_0[0]),.doutb(w_n14827_0[1]),.din(n14827));
	jspl jspl_w_n14831_0(.douta(w_n14831_0[0]),.doutb(w_n14831_0[1]),.din(n14831));
	jspl3 jspl3_w_n14833_0(.douta(w_n14833_0[0]),.doutb(w_n14833_0[1]),.doutc(w_n14833_0[2]),.din(n14833));
	jspl jspl_w_n14834_0(.douta(w_n14834_0[0]),.doutb(w_n14834_0[1]),.din(n14834));
	jspl jspl_w_n14838_0(.douta(w_n14838_0[0]),.doutb(w_n14838_0[1]),.din(n14838));
	jspl jspl_w_n14839_0(.douta(w_n14839_0[0]),.doutb(w_n14839_0[1]),.din(n14839));
	jspl3 jspl3_w_n14841_0(.douta(w_n14841_0[0]),.doutb(w_n14841_0[1]),.doutc(w_n14841_0[2]),.din(n14841));
	jspl jspl_w_n14842_0(.douta(w_n14842_0[0]),.doutb(w_n14842_0[1]),.din(n14842));
	jspl jspl_w_n14846_0(.douta(w_n14846_0[0]),.doutb(w_n14846_0[1]),.din(n14846));
	jspl jspl_w_n14847_0(.douta(w_n14847_0[0]),.doutb(w_n14847_0[1]),.din(n14847));
	jspl3 jspl3_w_n14849_0(.douta(w_n14849_0[0]),.doutb(w_n14849_0[1]),.doutc(w_n14849_0[2]),.din(n14849));
	jspl jspl_w_n14850_0(.douta(w_n14850_0[0]),.doutb(w_n14850_0[1]),.din(n14850));
	jspl jspl_w_n14854_0(.douta(w_n14854_0[0]),.doutb(w_n14854_0[1]),.din(n14854));
	jspl jspl_w_n14855_0(.douta(w_n14855_0[0]),.doutb(w_n14855_0[1]),.din(n14855));
	jspl3 jspl3_w_n14857_0(.douta(w_n14857_0[0]),.doutb(w_n14857_0[1]),.doutc(w_n14857_0[2]),.din(n14857));
	jspl jspl_w_n14858_0(.douta(w_n14858_0[0]),.doutb(w_n14858_0[1]),.din(n14858));
	jspl jspl_w_n14862_0(.douta(w_n14862_0[0]),.doutb(w_n14862_0[1]),.din(n14862));
	jspl3 jspl3_w_n14864_0(.douta(w_n14864_0[0]),.doutb(w_n14864_0[1]),.doutc(w_n14864_0[2]),.din(n14864));
	jspl jspl_w_n14865_0(.douta(w_n14865_0[0]),.doutb(w_n14865_0[1]),.din(n14865));
	jspl jspl_w_n14869_0(.douta(w_n14869_0[0]),.doutb(w_n14869_0[1]),.din(n14869));
	jspl jspl_w_n14870_0(.douta(w_n14870_0[0]),.doutb(w_n14870_0[1]),.din(n14870));
	jspl3 jspl3_w_n14872_0(.douta(w_n14872_0[0]),.doutb(w_n14872_0[1]),.doutc(w_n14872_0[2]),.din(n14872));
	jspl jspl_w_n14873_0(.douta(w_n14873_0[0]),.doutb(w_n14873_0[1]),.din(n14873));
	jspl jspl_w_n14877_0(.douta(w_n14877_0[0]),.doutb(w_n14877_0[1]),.din(n14877));
	jspl3 jspl3_w_n14879_0(.douta(w_n14879_0[0]),.doutb(w_n14879_0[1]),.doutc(w_n14879_0[2]),.din(n14879));
	jspl jspl_w_n14880_0(.douta(w_n14880_0[0]),.doutb(w_n14880_0[1]),.din(n14880));
	jspl jspl_w_n14884_0(.douta(w_n14884_0[0]),.doutb(w_n14884_0[1]),.din(n14884));
	jspl jspl_w_n14885_0(.douta(w_n14885_0[0]),.doutb(w_n14885_0[1]),.din(n14885));
	jspl3 jspl3_w_n14887_0(.douta(w_n14887_0[0]),.doutb(w_n14887_0[1]),.doutc(w_n14887_0[2]),.din(n14887));
	jspl jspl_w_n14888_0(.douta(w_n14888_0[0]),.doutb(w_n14888_0[1]),.din(n14888));
	jspl jspl_w_n14892_0(.douta(w_n14892_0[0]),.doutb(w_n14892_0[1]),.din(n14892));
	jspl jspl_w_n14893_0(.douta(w_n14893_0[0]),.doutb(w_n14893_0[1]),.din(n14893));
	jspl3 jspl3_w_n14895_0(.douta(w_n14895_0[0]),.doutb(w_n14895_0[1]),.doutc(w_n14895_0[2]),.din(n14895));
	jspl jspl_w_n14896_0(.douta(w_n14896_0[0]),.doutb(w_n14896_0[1]),.din(n14896));
	jspl jspl_w_n14900_0(.douta(w_n14900_0[0]),.doutb(w_n14900_0[1]),.din(n14900));
	jspl3 jspl3_w_n14902_0(.douta(w_n14902_0[0]),.doutb(w_n14902_0[1]),.doutc(w_n14902_0[2]),.din(n14902));
	jspl jspl_w_n14903_0(.douta(w_n14903_0[0]),.doutb(w_n14903_0[1]),.din(n14903));
	jspl jspl_w_n14906_0(.douta(w_n14906_0[0]),.doutb(w_n14906_0[1]),.din(n14906));
	jspl3 jspl3_w_n14909_0(.douta(w_n14909_0[0]),.doutb(w_n14909_0[1]),.doutc(w_n14909_0[2]),.din(n14909));
	jspl jspl_w_n14910_0(.douta(w_n14910_0[0]),.doutb(w_n14910_0[1]),.din(n14910));
	jspl jspl_w_n14914_0(.douta(w_n14914_0[0]),.doutb(w_n14914_0[1]),.din(n14914));
	jspl jspl_w_n14915_0(.douta(w_n14915_0[0]),.doutb(w_n14915_0[1]),.din(n14915));
	jspl3 jspl3_w_n14917_0(.douta(w_n14917_0[0]),.doutb(w_n14917_0[1]),.doutc(w_n14917_0[2]),.din(n14917));
	jspl jspl_w_n14918_0(.douta(w_n14918_0[0]),.doutb(w_n14918_0[1]),.din(n14918));
	jspl jspl_w_n14922_0(.douta(w_n14922_0[0]),.doutb(w_n14922_0[1]),.din(n14922));
	jspl3 jspl3_w_n14924_0(.douta(w_n14924_0[0]),.doutb(w_n14924_0[1]),.doutc(w_n14924_0[2]),.din(n14924));
	jspl jspl_w_n14925_0(.douta(w_n14925_0[0]),.doutb(w_n14925_0[1]),.din(n14925));
	jspl jspl_w_n14929_0(.douta(w_n14929_0[0]),.doutb(w_n14929_0[1]),.din(n14929));
	jspl jspl_w_n14930_0(.douta(w_n14930_0[0]),.doutb(w_n14930_0[1]),.din(n14930));
	jspl3 jspl3_w_n14932_0(.douta(w_n14932_0[0]),.doutb(w_n14932_0[1]),.doutc(w_n14932_0[2]),.din(n14932));
	jspl jspl_w_n14933_0(.douta(w_n14933_0[0]),.doutb(w_n14933_0[1]),.din(n14933));
	jspl jspl_w_n14937_0(.douta(w_n14937_0[0]),.doutb(w_n14937_0[1]),.din(n14937));
	jspl3 jspl3_w_n14939_0(.douta(w_n14939_0[0]),.doutb(w_n14939_0[1]),.doutc(w_n14939_0[2]),.din(n14939));
	jspl jspl_w_n14940_0(.douta(w_n14940_0[0]),.doutb(w_n14940_0[1]),.din(n14940));
	jspl jspl_w_n14944_0(.douta(w_n14944_0[0]),.doutb(w_n14944_0[1]),.din(n14944));
	jspl jspl_w_n14945_0(.douta(w_n14945_0[0]),.doutb(w_n14945_0[1]),.din(n14945));
	jspl3 jspl3_w_n14947_0(.douta(w_n14947_0[0]),.doutb(w_n14947_0[1]),.doutc(w_n14947_0[2]),.din(n14947));
	jspl jspl_w_n14948_0(.douta(w_n14948_0[0]),.doutb(w_n14948_0[1]),.din(n14948));
	jspl jspl_w_n14952_0(.douta(w_n14952_0[0]),.doutb(w_n14952_0[1]),.din(n14952));
	jspl jspl_w_n14953_0(.douta(w_n14953_0[0]),.doutb(w_n14953_0[1]),.din(n14953));
	jspl3 jspl3_w_n14955_0(.douta(w_n14955_0[0]),.doutb(w_n14955_0[1]),.doutc(w_n14955_0[2]),.din(n14955));
	jspl jspl_w_n14956_0(.douta(w_n14956_0[0]),.doutb(w_n14956_0[1]),.din(n14956));
	jspl jspl_w_n14960_0(.douta(w_n14960_0[0]),.doutb(w_n14960_0[1]),.din(n14960));
	jspl jspl_w_n14961_0(.douta(w_n14961_0[0]),.doutb(w_n14961_0[1]),.din(n14961));
	jspl3 jspl3_w_n14963_0(.douta(w_n14963_0[0]),.doutb(w_n14963_0[1]),.doutc(w_n14963_0[2]),.din(n14963));
	jspl jspl_w_n14964_0(.douta(w_n14964_0[0]),.doutb(w_n14964_0[1]),.din(n14964));
	jspl jspl_w_n14968_0(.douta(w_n14968_0[0]),.doutb(w_n14968_0[1]),.din(n14968));
	jspl3 jspl3_w_n14970_0(.douta(w_n14970_0[0]),.doutb(w_n14970_0[1]),.doutc(w_n14970_0[2]),.din(n14970));
	jspl jspl_w_n14971_0(.douta(w_n14971_0[0]),.doutb(w_n14971_0[1]),.din(n14971));
	jspl jspl_w_n14975_0(.douta(w_n14975_0[0]),.doutb(w_n14975_0[1]),.din(n14975));
	jspl jspl_w_n14976_0(.douta(w_n14976_0[0]),.doutb(w_n14976_0[1]),.din(n14976));
	jspl3 jspl3_w_n14978_0(.douta(w_n14978_0[0]),.doutb(w_n14978_0[1]),.doutc(w_n14978_0[2]),.din(n14978));
	jspl jspl_w_n14979_0(.douta(w_n14979_0[0]),.doutb(w_n14979_0[1]),.din(n14979));
	jspl jspl_w_n14983_0(.douta(w_n14983_0[0]),.doutb(w_n14983_0[1]),.din(n14983));
	jspl3 jspl3_w_n14985_0(.douta(w_n14985_0[0]),.doutb(w_n14985_0[1]),.doutc(w_n14985_0[2]),.din(n14985));
	jspl jspl_w_n14986_0(.douta(w_n14986_0[0]),.doutb(w_n14986_0[1]),.din(n14986));
	jspl jspl_w_n14990_0(.douta(w_n14990_0[0]),.doutb(w_n14990_0[1]),.din(n14990));
	jspl jspl_w_n14991_0(.douta(w_n14991_0[0]),.doutb(w_n14991_0[1]),.din(n14991));
	jspl3 jspl3_w_n14993_0(.douta(w_n14993_0[0]),.doutb(w_n14993_0[1]),.doutc(w_n14993_0[2]),.din(n14993));
	jspl jspl_w_n14994_0(.douta(w_n14994_0[0]),.doutb(w_n14994_0[1]),.din(n14994));
	jspl jspl_w_n14998_0(.douta(w_n14998_0[0]),.doutb(w_n14998_0[1]),.din(n14998));
	jspl3 jspl3_w_n15000_0(.douta(w_n15000_0[0]),.doutb(w_n15000_0[1]),.doutc(w_n15000_0[2]),.din(n15000));
	jspl jspl_w_n15001_0(.douta(w_n15001_0[0]),.doutb(w_n15001_0[1]),.din(n15001));
	jspl jspl_w_n15005_0(.douta(w_n15005_0[0]),.doutb(w_n15005_0[1]),.din(n15005));
	jspl jspl_w_n15006_0(.douta(w_n15006_0[0]),.doutb(w_n15006_0[1]),.din(n15006));
	jspl3 jspl3_w_n15008_0(.douta(w_n15008_0[0]),.doutb(w_n15008_0[1]),.doutc(w_n15008_0[2]),.din(n15008));
	jspl jspl_w_n15009_0(.douta(w_n15009_0[0]),.doutb(w_n15009_0[1]),.din(n15009));
	jspl jspl_w_n15013_0(.douta(w_n15013_0[0]),.doutb(w_n15013_0[1]),.din(n15013));
	jspl3 jspl3_w_n15015_0(.douta(w_n15015_0[0]),.doutb(w_n15015_0[1]),.doutc(w_n15015_0[2]),.din(n15015));
	jspl jspl_w_n15016_0(.douta(w_n15016_0[0]),.doutb(w_n15016_0[1]),.din(n15016));
	jspl jspl_w_n15033_0(.douta(w_n15033_0[0]),.doutb(w_n15033_0[1]),.din(n15033));
	jspl jspl_w_n15070_0(.douta(w_n15070_0[0]),.doutb(w_n15070_0[1]),.din(n15070));
	jspl jspl_w_n15077_0(.douta(w_n15077_0[0]),.doutb(w_n15077_0[1]),.din(n15077));
	jspl jspl_w_n15084_0(.douta(w_n15084_0[0]),.doutb(w_n15084_0[1]),.din(n15084));
	jspl jspl_w_n15097_0(.douta(w_n15097_0[0]),.doutb(w_n15097_0[1]),.din(n15097));
	jspl jspl_w_n15104_0(.douta(w_n15104_0[0]),.doutb(w_n15104_0[1]),.din(n15104));
	jspl jspl_w_n15111_0(.douta(w_n15111_0[0]),.doutb(w_n15111_0[1]),.din(n15111));
	jspl jspl_w_n15118_0(.douta(w_n15118_0[0]),.doutb(w_n15118_0[1]),.din(n15118));
	jspl jspl_w_n15131_0(.douta(w_n15131_0[0]),.doutb(w_n15131_0[1]),.din(n15131));
	jspl jspl_w_n15138_0(.douta(w_n15138_0[0]),.doutb(w_n15138_0[1]),.din(n15138));
	jspl jspl_w_n15151_0(.douta(w_n15151_0[0]),.doutb(w_n15151_0[1]),.din(n15151));
	jspl jspl_w_n15158_0(.douta(w_n15158_0[0]),.doutb(w_n15158_0[1]),.din(n15158));
	jspl jspl_w_n15168_0(.douta(w_n15168_0[0]),.doutb(w_n15168_0[1]),.din(n15168));
	jspl jspl_w_n15178_0(.douta(w_n15178_0[0]),.doutb(w_n15178_0[1]),.din(n15178));
	jspl jspl_w_n15185_0(.douta(w_n15185_0[0]),.doutb(w_n15185_0[1]),.din(n15185));
	jspl jspl_w_n15198_0(.douta(w_n15198_0[0]),.doutb(w_n15198_0[1]),.din(n15198));
	jspl jspl_w_n15205_0(.douta(w_n15205_0[0]),.doutb(w_n15205_0[1]),.din(n15205));
	jspl jspl_w_n15212_0(.douta(w_n15212_0[0]),.doutb(w_n15212_0[1]),.din(n15212));
	jspl jspl_w_n15219_0(.douta(w_n15219_0[0]),.doutb(w_n15219_0[1]),.din(n15219));
	jspl jspl_w_n15225_0(.douta(w_n15225_0[0]),.doutb(w_n15225_0[1]),.din(n15225));
	jspl jspl_w_n15226_0(.douta(w_n15226_0[0]),.doutb(w_n15226_0[1]),.din(n15226));
	jspl3 jspl3_w_n15228_0(.douta(w_n15228_0[0]),.doutb(w_n15228_0[1]),.doutc(w_n15228_0[2]),.din(n15228));
	jspl3 jspl3_w_n15231_0(.douta(w_n15231_0[0]),.doutb(w_n15231_0[1]),.doutc(w_n15231_0[2]),.din(n15231));
	jspl jspl_w_n15231_1(.douta(w_n15231_1[0]),.doutb(w_n15231_1[1]),.din(w_n15231_0[0]));
	jspl jspl_w_n15232_0(.douta(w_n15232_0[0]),.doutb(w_n15232_0[1]),.din(n15232));
	jspl jspl_w_n15233_0(.douta(w_n15233_0[0]),.doutb(w_n15233_0[1]),.din(n15233));
	jspl jspl_w_n15235_0(.douta(w_n15235_0[0]),.doutb(w_n15235_0[1]),.din(n15235));
	jspl jspl_w_n15237_0(.douta(w_n15237_0[0]),.doutb(w_n15237_0[1]),.din(n15237));
	jspl jspl_w_n15238_0(.douta(w_n15238_0[0]),.doutb(w_n15238_0[1]),.din(n15238));
	jspl3 jspl3_w_n15239_0(.douta(w_n15239_0[0]),.doutb(w_n15239_0[1]),.doutc(w_n15239_0[2]),.din(n15239));
	jspl jspl_w_n15243_0(.douta(w_n15243_0[0]),.doutb(w_n15243_0[1]),.din(n15243));
	jspl jspl_w_n15244_0(.douta(w_n15244_0[0]),.doutb(w_n15244_0[1]),.din(n15244));
	jspl jspl_w_n15249_0(.douta(w_n15249_0[0]),.doutb(w_n15249_0[1]),.din(n15249));
	jspl jspl_w_n15250_0(.douta(w_n15250_0[0]),.doutb(w_n15250_0[1]),.din(n15250));
	jspl jspl_w_n15251_0(.douta(w_n15251_0[0]),.doutb(w_n15251_0[1]),.din(n15251));
	jspl3 jspl3_w_n15256_0(.douta(w_n15256_0[0]),.doutb(w_n15256_0[1]),.doutc(w_n15256_0[2]),.din(n15256));
	jspl3 jspl3_w_n15260_0(.douta(w_n15260_0[0]),.doutb(w_n15260_0[1]),.doutc(w_n15260_0[2]),.din(n15260));
	jspl3 jspl3_w_n15260_1(.douta(w_n15260_1[0]),.doutb(w_n15260_1[1]),.doutc(w_n15260_1[2]),.din(w_n15260_0[0]));
	jspl3 jspl3_w_n15260_2(.douta(w_n15260_2[0]),.doutb(w_n15260_2[1]),.doutc(w_n15260_2[2]),.din(w_n15260_0[1]));
	jspl3 jspl3_w_n15260_3(.douta(w_n15260_3[0]),.doutb(w_n15260_3[1]),.doutc(w_n15260_3[2]),.din(w_n15260_0[2]));
	jspl3 jspl3_w_n15260_4(.douta(w_n15260_4[0]),.doutb(w_n15260_4[1]),.doutc(w_n15260_4[2]),.din(w_n15260_1[0]));
	jspl3 jspl3_w_n15260_5(.douta(w_n15260_5[0]),.doutb(w_n15260_5[1]),.doutc(w_n15260_5[2]),.din(w_n15260_1[1]));
	jspl3 jspl3_w_n15260_6(.douta(w_n15260_6[0]),.doutb(w_n15260_6[1]),.doutc(w_n15260_6[2]),.din(w_n15260_1[2]));
	jspl3 jspl3_w_n15260_7(.douta(w_n15260_7[0]),.doutb(w_n15260_7[1]),.doutc(w_n15260_7[2]),.din(w_n15260_2[0]));
	jspl3 jspl3_w_n15260_8(.douta(w_n15260_8[0]),.doutb(w_n15260_8[1]),.doutc(w_n15260_8[2]),.din(w_n15260_2[1]));
	jspl3 jspl3_w_n15260_9(.douta(w_n15260_9[0]),.doutb(w_n15260_9[1]),.doutc(w_n15260_9[2]),.din(w_n15260_2[2]));
	jspl3 jspl3_w_n15260_10(.douta(w_n15260_10[0]),.doutb(w_n15260_10[1]),.doutc(w_n15260_10[2]),.din(w_n15260_3[0]));
	jspl3 jspl3_w_n15260_11(.douta(w_n15260_11[0]),.doutb(w_n15260_11[1]),.doutc(w_n15260_11[2]),.din(w_n15260_3[1]));
	jspl3 jspl3_w_n15260_12(.douta(w_n15260_12[0]),.doutb(w_n15260_12[1]),.doutc(w_n15260_12[2]),.din(w_n15260_3[2]));
	jspl3 jspl3_w_n15260_13(.douta(w_n15260_13[0]),.doutb(w_n15260_13[1]),.doutc(w_n15260_13[2]),.din(w_n15260_4[0]));
	jspl3 jspl3_w_n15260_14(.douta(w_n15260_14[0]),.doutb(w_n15260_14[1]),.doutc(w_n15260_14[2]),.din(w_n15260_4[1]));
	jspl3 jspl3_w_n15260_15(.douta(w_n15260_15[0]),.doutb(w_n15260_15[1]),.doutc(w_n15260_15[2]),.din(w_n15260_4[2]));
	jspl3 jspl3_w_n15260_16(.douta(w_n15260_16[0]),.doutb(w_n15260_16[1]),.doutc(w_n15260_16[2]),.din(w_n15260_5[0]));
	jspl3 jspl3_w_n15260_17(.douta(w_n15260_17[0]),.doutb(w_n15260_17[1]),.doutc(w_n15260_17[2]),.din(w_n15260_5[1]));
	jspl3 jspl3_w_n15260_18(.douta(w_n15260_18[0]),.doutb(w_n15260_18[1]),.doutc(w_n15260_18[2]),.din(w_n15260_5[2]));
	jspl3 jspl3_w_n15260_19(.douta(w_n15260_19[0]),.doutb(w_n15260_19[1]),.doutc(w_n15260_19[2]),.din(w_n15260_6[0]));
	jspl3 jspl3_w_n15260_20(.douta(w_n15260_20[0]),.doutb(w_n15260_20[1]),.doutc(w_n15260_20[2]),.din(w_n15260_6[1]));
	jspl3 jspl3_w_n15260_21(.douta(w_n15260_21[0]),.doutb(w_n15260_21[1]),.doutc(w_n15260_21[2]),.din(w_n15260_6[2]));
	jspl3 jspl3_w_n15260_22(.douta(w_n15260_22[0]),.doutb(w_n15260_22[1]),.doutc(w_n15260_22[2]),.din(w_n15260_7[0]));
	jspl3 jspl3_w_n15260_23(.douta(w_n15260_23[0]),.doutb(w_n15260_23[1]),.doutc(w_n15260_23[2]),.din(w_n15260_7[1]));
	jspl3 jspl3_w_n15260_24(.douta(w_n15260_24[0]),.doutb(w_n15260_24[1]),.doutc(w_n15260_24[2]),.din(w_n15260_7[2]));
	jspl3 jspl3_w_n15260_25(.douta(w_n15260_25[0]),.doutb(w_n15260_25[1]),.doutc(w_n15260_25[2]),.din(w_n15260_8[0]));
	jspl3 jspl3_w_n15260_26(.douta(w_n15260_26[0]),.doutb(w_n15260_26[1]),.doutc(w_n15260_26[2]),.din(w_n15260_8[1]));
	jspl3 jspl3_w_n15260_27(.douta(w_n15260_27[0]),.doutb(w_n15260_27[1]),.doutc(w_n15260_27[2]),.din(w_n15260_8[2]));
	jspl3 jspl3_w_n15260_28(.douta(w_n15260_28[0]),.doutb(w_n15260_28[1]),.doutc(w_n15260_28[2]),.din(w_n15260_9[0]));
	jspl3 jspl3_w_n15260_29(.douta(w_n15260_29[0]),.doutb(w_n15260_29[1]),.doutc(w_n15260_29[2]),.din(w_n15260_9[1]));
	jspl3 jspl3_w_n15260_30(.douta(w_n15260_30[0]),.doutb(w_n15260_30[1]),.doutc(w_n15260_30[2]),.din(w_n15260_9[2]));
	jspl3 jspl3_w_n15260_31(.douta(w_n15260_31[0]),.doutb(w_n15260_31[1]),.doutc(w_n15260_31[2]),.din(w_n15260_10[0]));
	jspl3 jspl3_w_n15260_32(.douta(w_n15260_32[0]),.doutb(w_n15260_32[1]),.doutc(w_n15260_32[2]),.din(w_n15260_10[1]));
	jspl3 jspl3_w_n15260_33(.douta(w_n15260_33[0]),.doutb(w_n15260_33[1]),.doutc(w_n15260_33[2]),.din(w_n15260_10[2]));
	jspl3 jspl3_w_n15260_34(.douta(w_n15260_34[0]),.doutb(w_n15260_34[1]),.doutc(w_n15260_34[2]),.din(w_n15260_11[0]));
	jspl3 jspl3_w_n15260_35(.douta(w_n15260_35[0]),.doutb(w_n15260_35[1]),.doutc(w_n15260_35[2]),.din(w_n15260_11[1]));
	jspl3 jspl3_w_n15260_36(.douta(w_n15260_36[0]),.doutb(w_n15260_36[1]),.doutc(w_n15260_36[2]),.din(w_n15260_11[2]));
	jspl3 jspl3_w_n15260_37(.douta(w_n15260_37[0]),.doutb(w_n15260_37[1]),.doutc(w_n15260_37[2]),.din(w_n15260_12[0]));
	jspl3 jspl3_w_n15260_38(.douta(w_n15260_38[0]),.doutb(w_n15260_38[1]),.doutc(w_n15260_38[2]),.din(w_n15260_12[1]));
	jspl3 jspl3_w_n15260_39(.douta(w_n15260_39[0]),.doutb(w_n15260_39[1]),.doutc(w_n15260_39[2]),.din(w_n15260_12[2]));
	jspl3 jspl3_w_n15260_40(.douta(w_n15260_40[0]),.doutb(w_n15260_40[1]),.doutc(w_n15260_40[2]),.din(w_n15260_13[0]));
	jspl3 jspl3_w_n15260_41(.douta(w_n15260_41[0]),.doutb(w_n15260_41[1]),.doutc(w_n15260_41[2]),.din(w_n15260_13[1]));
	jspl jspl_w_n15263_0(.douta(w_n15263_0[0]),.doutb(w_n15263_0[1]),.din(n15263));
	jspl3 jspl3_w_n15264_0(.douta(w_n15264_0[0]),.doutb(w_n15264_0[1]),.doutc(w_n15264_0[2]),.din(n15264));
	jspl3 jspl3_w_n15265_0(.douta(w_n15265_0[0]),.doutb(w_n15265_0[1]),.doutc(w_n15265_0[2]),.din(n15265));
	jspl3 jspl3_w_n15265_1(.douta(w_n15265_1[0]),.doutb(w_n15265_1[1]),.doutc(w_n15265_1[2]),.din(w_n15265_0[0]));
	jspl jspl_w_n15266_0(.douta(w_n15266_0[0]),.doutb(w_n15266_0[1]),.din(n15266));
	jspl3 jspl3_w_n15267_0(.douta(w_n15267_0[0]),.doutb(w_n15267_0[1]),.doutc(w_n15267_0[2]),.din(n15267));
	jspl jspl_w_n15268_0(.douta(w_n15268_0[0]),.doutb(w_n15268_0[1]),.din(n15268));
	jspl3 jspl3_w_n15271_0(.douta(w_n15271_0[0]),.doutb(w_n15271_0[1]),.doutc(w_n15271_0[2]),.din(n15271));
	jspl jspl_w_n15272_0(.douta(w_n15272_0[0]),.doutb(w_n15272_0[1]),.din(n15272));
	jspl3 jspl3_w_n15279_0(.douta(w_n15279_0[0]),.doutb(w_n15279_0[1]),.doutc(w_n15279_0[2]),.din(n15279));
	jspl jspl_w_n15280_0(.douta(w_n15280_0[0]),.doutb(w_n15280_0[1]),.din(n15280));
	jspl jspl_w_n15283_0(.douta(w_n15283_0[0]),.doutb(w_n15283_0[1]),.din(n15283));
	jspl jspl_w_n15288_0(.douta(w_n15288_0[0]),.doutb(w_n15288_0[1]),.din(n15288));
	jspl3 jspl3_w_n15290_0(.douta(w_n15290_0[0]),.doutb(w_n15290_0[1]),.doutc(w_n15290_0[2]),.din(n15290));
	jspl jspl_w_n15291_0(.douta(w_n15291_0[0]),.doutb(w_n15291_0[1]),.din(n15291));
	jspl3 jspl3_w_n15295_0(.douta(w_n15295_0[0]),.doutb(w_n15295_0[1]),.doutc(w_n15295_0[2]),.din(n15295));
	jspl3 jspl3_w_n15298_0(.douta(w_n15298_0[0]),.doutb(w_n15298_0[1]),.doutc(w_n15298_0[2]),.din(n15298));
	jspl jspl_w_n15299_0(.douta(w_n15299_0[0]),.doutb(w_n15299_0[1]),.din(n15299));
	jspl3 jspl3_w_n15303_0(.douta(w_n15303_0[0]),.doutb(w_n15303_0[1]),.doutc(w_n15303_0[2]),.din(n15303));
	jspl3 jspl3_w_n15305_0(.douta(w_n15305_0[0]),.doutb(w_n15305_0[1]),.doutc(w_n15305_0[2]),.din(n15305));
	jspl jspl_w_n15306_0(.douta(w_n15306_0[0]),.doutb(w_n15306_0[1]),.din(n15306));
	jspl3 jspl3_w_n15310_0(.douta(w_n15310_0[0]),.doutb(w_n15310_0[1]),.doutc(w_n15310_0[2]),.din(n15310));
	jspl3 jspl3_w_n15313_0(.douta(w_n15313_0[0]),.doutb(w_n15313_0[1]),.doutc(w_n15313_0[2]),.din(n15313));
	jspl jspl_w_n15314_0(.douta(w_n15314_0[0]),.doutb(w_n15314_0[1]),.din(n15314));
	jspl3 jspl3_w_n15318_0(.douta(w_n15318_0[0]),.doutb(w_n15318_0[1]),.doutc(w_n15318_0[2]),.din(n15318));
	jspl3 jspl3_w_n15320_0(.douta(w_n15320_0[0]),.doutb(w_n15320_0[1]),.doutc(w_n15320_0[2]),.din(n15320));
	jspl jspl_w_n15321_0(.douta(w_n15321_0[0]),.doutb(w_n15321_0[1]),.din(n15321));
	jspl3 jspl3_w_n15325_0(.douta(w_n15325_0[0]),.doutb(w_n15325_0[1]),.doutc(w_n15325_0[2]),.din(n15325));
	jspl3 jspl3_w_n15328_0(.douta(w_n15328_0[0]),.doutb(w_n15328_0[1]),.doutc(w_n15328_0[2]),.din(n15328));
	jspl jspl_w_n15329_0(.douta(w_n15329_0[0]),.doutb(w_n15329_0[1]),.din(n15329));
	jspl3 jspl3_w_n15333_0(.douta(w_n15333_0[0]),.doutb(w_n15333_0[1]),.doutc(w_n15333_0[2]),.din(n15333));
	jspl3 jspl3_w_n15335_0(.douta(w_n15335_0[0]),.doutb(w_n15335_0[1]),.doutc(w_n15335_0[2]),.din(n15335));
	jspl jspl_w_n15336_0(.douta(w_n15336_0[0]),.doutb(w_n15336_0[1]),.din(n15336));
	jspl3 jspl3_w_n15340_0(.douta(w_n15340_0[0]),.doutb(w_n15340_0[1]),.doutc(w_n15340_0[2]),.din(n15340));
	jspl3 jspl3_w_n15342_0(.douta(w_n15342_0[0]),.doutb(w_n15342_0[1]),.doutc(w_n15342_0[2]),.din(n15342));
	jspl jspl_w_n15343_0(.douta(w_n15343_0[0]),.doutb(w_n15343_0[1]),.din(n15343));
	jspl3 jspl3_w_n15347_0(.douta(w_n15347_0[0]),.doutb(w_n15347_0[1]),.doutc(w_n15347_0[2]),.din(n15347));
	jspl3 jspl3_w_n15349_0(.douta(w_n15349_0[0]),.doutb(w_n15349_0[1]),.doutc(w_n15349_0[2]),.din(n15349));
	jspl jspl_w_n15350_0(.douta(w_n15350_0[0]),.doutb(w_n15350_0[1]),.din(n15350));
	jspl3 jspl3_w_n15354_0(.douta(w_n15354_0[0]),.doutb(w_n15354_0[1]),.doutc(w_n15354_0[2]),.din(n15354));
	jspl3 jspl3_w_n15357_0(.douta(w_n15357_0[0]),.doutb(w_n15357_0[1]),.doutc(w_n15357_0[2]),.din(n15357));
	jspl jspl_w_n15358_0(.douta(w_n15358_0[0]),.doutb(w_n15358_0[1]),.din(n15358));
	jspl3 jspl3_w_n15362_0(.douta(w_n15362_0[0]),.doutb(w_n15362_0[1]),.doutc(w_n15362_0[2]),.din(n15362));
	jspl3 jspl3_w_n15364_0(.douta(w_n15364_0[0]),.doutb(w_n15364_0[1]),.doutc(w_n15364_0[2]),.din(n15364));
	jspl jspl_w_n15365_0(.douta(w_n15365_0[0]),.doutb(w_n15365_0[1]),.din(n15365));
	jspl3 jspl3_w_n15369_0(.douta(w_n15369_0[0]),.doutb(w_n15369_0[1]),.doutc(w_n15369_0[2]),.din(n15369));
	jspl3 jspl3_w_n15372_0(.douta(w_n15372_0[0]),.doutb(w_n15372_0[1]),.doutc(w_n15372_0[2]),.din(n15372));
	jspl jspl_w_n15373_0(.douta(w_n15373_0[0]),.doutb(w_n15373_0[1]),.din(n15373));
	jspl3 jspl3_w_n15377_0(.douta(w_n15377_0[0]),.doutb(w_n15377_0[1]),.doutc(w_n15377_0[2]),.din(n15377));
	jspl3 jspl3_w_n15379_0(.douta(w_n15379_0[0]),.doutb(w_n15379_0[1]),.doutc(w_n15379_0[2]),.din(n15379));
	jspl jspl_w_n15380_0(.douta(w_n15380_0[0]),.doutb(w_n15380_0[1]),.din(n15380));
	jspl3 jspl3_w_n15384_0(.douta(w_n15384_0[0]),.doutb(w_n15384_0[1]),.doutc(w_n15384_0[2]),.din(n15384));
	jspl3 jspl3_w_n15387_0(.douta(w_n15387_0[0]),.doutb(w_n15387_0[1]),.doutc(w_n15387_0[2]),.din(n15387));
	jspl jspl_w_n15388_0(.douta(w_n15388_0[0]),.doutb(w_n15388_0[1]),.din(n15388));
	jspl3 jspl3_w_n15392_0(.douta(w_n15392_0[0]),.doutb(w_n15392_0[1]),.doutc(w_n15392_0[2]),.din(n15392));
	jspl3 jspl3_w_n15394_0(.douta(w_n15394_0[0]),.doutb(w_n15394_0[1]),.doutc(w_n15394_0[2]),.din(n15394));
	jspl jspl_w_n15395_0(.douta(w_n15395_0[0]),.doutb(w_n15395_0[1]),.din(n15395));
	jspl3 jspl3_w_n15399_0(.douta(w_n15399_0[0]),.doutb(w_n15399_0[1]),.doutc(w_n15399_0[2]),.din(n15399));
	jspl3 jspl3_w_n15402_0(.douta(w_n15402_0[0]),.doutb(w_n15402_0[1]),.doutc(w_n15402_0[2]),.din(n15402));
	jspl jspl_w_n15403_0(.douta(w_n15403_0[0]),.doutb(w_n15403_0[1]),.din(n15403));
	jspl3 jspl3_w_n15407_0(.douta(w_n15407_0[0]),.doutb(w_n15407_0[1]),.doutc(w_n15407_0[2]),.din(n15407));
	jspl3 jspl3_w_n15409_0(.douta(w_n15409_0[0]),.doutb(w_n15409_0[1]),.doutc(w_n15409_0[2]),.din(n15409));
	jspl jspl_w_n15410_0(.douta(w_n15410_0[0]),.doutb(w_n15410_0[1]),.din(n15410));
	jspl3 jspl3_w_n15414_0(.douta(w_n15414_0[0]),.doutb(w_n15414_0[1]),.doutc(w_n15414_0[2]),.din(n15414));
	jspl3 jspl3_w_n15416_0(.douta(w_n15416_0[0]),.doutb(w_n15416_0[1]),.doutc(w_n15416_0[2]),.din(n15416));
	jspl jspl_w_n15417_0(.douta(w_n15417_0[0]),.doutb(w_n15417_0[1]),.din(n15417));
	jspl3 jspl3_w_n15421_0(.douta(w_n15421_0[0]),.doutb(w_n15421_0[1]),.doutc(w_n15421_0[2]),.din(n15421));
	jspl3 jspl3_w_n15423_0(.douta(w_n15423_0[0]),.doutb(w_n15423_0[1]),.doutc(w_n15423_0[2]),.din(n15423));
	jspl jspl_w_n15424_0(.douta(w_n15424_0[0]),.doutb(w_n15424_0[1]),.din(n15424));
	jspl3 jspl3_w_n15428_0(.douta(w_n15428_0[0]),.doutb(w_n15428_0[1]),.doutc(w_n15428_0[2]),.din(n15428));
	jspl3 jspl3_w_n15431_0(.douta(w_n15431_0[0]),.doutb(w_n15431_0[1]),.doutc(w_n15431_0[2]),.din(n15431));
	jspl jspl_w_n15432_0(.douta(w_n15432_0[0]),.doutb(w_n15432_0[1]),.din(n15432));
	jspl3 jspl3_w_n15436_0(.douta(w_n15436_0[0]),.doutb(w_n15436_0[1]),.doutc(w_n15436_0[2]),.din(n15436));
	jspl3 jspl3_w_n15438_0(.douta(w_n15438_0[0]),.doutb(w_n15438_0[1]),.doutc(w_n15438_0[2]),.din(n15438));
	jspl jspl_w_n15439_0(.douta(w_n15439_0[0]),.doutb(w_n15439_0[1]),.din(n15439));
	jspl3 jspl3_w_n15443_0(.douta(w_n15443_0[0]),.doutb(w_n15443_0[1]),.doutc(w_n15443_0[2]),.din(n15443));
	jspl3 jspl3_w_n15446_0(.douta(w_n15446_0[0]),.doutb(w_n15446_0[1]),.doutc(w_n15446_0[2]),.din(n15446));
	jspl jspl_w_n15447_0(.douta(w_n15447_0[0]),.doutb(w_n15447_0[1]),.din(n15447));
	jspl3 jspl3_w_n15451_0(.douta(w_n15451_0[0]),.doutb(w_n15451_0[1]),.doutc(w_n15451_0[2]),.din(n15451));
	jspl3 jspl3_w_n15453_0(.douta(w_n15453_0[0]),.doutb(w_n15453_0[1]),.doutc(w_n15453_0[2]),.din(n15453));
	jspl jspl_w_n15454_0(.douta(w_n15454_0[0]),.doutb(w_n15454_0[1]),.din(n15454));
	jspl3 jspl3_w_n15458_0(.douta(w_n15458_0[0]),.doutb(w_n15458_0[1]),.doutc(w_n15458_0[2]),.din(n15458));
	jspl3 jspl3_w_n15460_0(.douta(w_n15460_0[0]),.doutb(w_n15460_0[1]),.doutc(w_n15460_0[2]),.din(n15460));
	jspl jspl_w_n15461_0(.douta(w_n15461_0[0]),.doutb(w_n15461_0[1]),.din(n15461));
	jspl3 jspl3_w_n15465_0(.douta(w_n15465_0[0]),.doutb(w_n15465_0[1]),.doutc(w_n15465_0[2]),.din(n15465));
	jspl3 jspl3_w_n15467_0(.douta(w_n15467_0[0]),.doutb(w_n15467_0[1]),.doutc(w_n15467_0[2]),.din(n15467));
	jspl jspl_w_n15468_0(.douta(w_n15468_0[0]),.doutb(w_n15468_0[1]),.din(n15468));
	jspl3 jspl3_w_n15472_0(.douta(w_n15472_0[0]),.doutb(w_n15472_0[1]),.doutc(w_n15472_0[2]),.din(n15472));
	jspl3 jspl3_w_n15475_0(.douta(w_n15475_0[0]),.doutb(w_n15475_0[1]),.doutc(w_n15475_0[2]),.din(n15475));
	jspl jspl_w_n15476_0(.douta(w_n15476_0[0]),.doutb(w_n15476_0[1]),.din(n15476));
	jspl3 jspl3_w_n15480_0(.douta(w_n15480_0[0]),.doutb(w_n15480_0[1]),.doutc(w_n15480_0[2]),.din(n15480));
	jspl3 jspl3_w_n15482_0(.douta(w_n15482_0[0]),.doutb(w_n15482_0[1]),.doutc(w_n15482_0[2]),.din(n15482));
	jspl jspl_w_n15483_0(.douta(w_n15483_0[0]),.doutb(w_n15483_0[1]),.din(n15483));
	jspl3 jspl3_w_n15487_0(.douta(w_n15487_0[0]),.doutb(w_n15487_0[1]),.doutc(w_n15487_0[2]),.din(n15487));
	jspl3 jspl3_w_n15490_0(.douta(w_n15490_0[0]),.doutb(w_n15490_0[1]),.doutc(w_n15490_0[2]),.din(n15490));
	jspl jspl_w_n15491_0(.douta(w_n15491_0[0]),.doutb(w_n15491_0[1]),.din(n15491));
	jspl3 jspl3_w_n15495_0(.douta(w_n15495_0[0]),.doutb(w_n15495_0[1]),.doutc(w_n15495_0[2]),.din(n15495));
	jspl3 jspl3_w_n15497_0(.douta(w_n15497_0[0]),.doutb(w_n15497_0[1]),.doutc(w_n15497_0[2]),.din(n15497));
	jspl jspl_w_n15498_0(.douta(w_n15498_0[0]),.doutb(w_n15498_0[1]),.din(n15498));
	jspl3 jspl3_w_n15502_0(.douta(w_n15502_0[0]),.doutb(w_n15502_0[1]),.doutc(w_n15502_0[2]),.din(n15502));
	jspl3 jspl3_w_n15504_0(.douta(w_n15504_0[0]),.doutb(w_n15504_0[1]),.doutc(w_n15504_0[2]),.din(n15504));
	jspl jspl_w_n15505_0(.douta(w_n15505_0[0]),.doutb(w_n15505_0[1]),.din(n15505));
	jspl3 jspl3_w_n15509_0(.douta(w_n15509_0[0]),.doutb(w_n15509_0[1]),.doutc(w_n15509_0[2]),.din(n15509));
	jspl3 jspl3_w_n15512_0(.douta(w_n15512_0[0]),.doutb(w_n15512_0[1]),.doutc(w_n15512_0[2]),.din(n15512));
	jspl jspl_w_n15513_0(.douta(w_n15513_0[0]),.doutb(w_n15513_0[1]),.din(n15513));
	jspl3 jspl3_w_n15516_0(.douta(w_n15516_0[0]),.doutb(w_n15516_0[1]),.doutc(w_n15516_0[2]),.din(n15516));
	jspl3 jspl3_w_n15520_0(.douta(w_n15520_0[0]),.doutb(w_n15520_0[1]),.doutc(w_n15520_0[2]),.din(n15520));
	jspl jspl_w_n15521_0(.douta(w_n15521_0[0]),.doutb(w_n15521_0[1]),.din(n15521));
	jspl3 jspl3_w_n15525_0(.douta(w_n15525_0[0]),.doutb(w_n15525_0[1]),.doutc(w_n15525_0[2]),.din(n15525));
	jspl3 jspl3_w_n15527_0(.douta(w_n15527_0[0]),.doutb(w_n15527_0[1]),.doutc(w_n15527_0[2]),.din(n15527));
	jspl jspl_w_n15528_0(.douta(w_n15528_0[0]),.doutb(w_n15528_0[1]),.din(n15528));
	jspl3 jspl3_w_n15532_0(.douta(w_n15532_0[0]),.doutb(w_n15532_0[1]),.doutc(w_n15532_0[2]),.din(n15532));
	jspl3 jspl3_w_n15535_0(.douta(w_n15535_0[0]),.doutb(w_n15535_0[1]),.doutc(w_n15535_0[2]),.din(n15535));
	jspl jspl_w_n15536_0(.douta(w_n15536_0[0]),.doutb(w_n15536_0[1]),.din(n15536));
	jspl3 jspl3_w_n15540_0(.douta(w_n15540_0[0]),.doutb(w_n15540_0[1]),.doutc(w_n15540_0[2]),.din(n15540));
	jspl3 jspl3_w_n15542_0(.douta(w_n15542_0[0]),.doutb(w_n15542_0[1]),.doutc(w_n15542_0[2]),.din(n15542));
	jspl jspl_w_n15543_0(.douta(w_n15543_0[0]),.doutb(w_n15543_0[1]),.din(n15543));
	jspl3 jspl3_w_n15547_0(.douta(w_n15547_0[0]),.doutb(w_n15547_0[1]),.doutc(w_n15547_0[2]),.din(n15547));
	jspl3 jspl3_w_n15550_0(.douta(w_n15550_0[0]),.doutb(w_n15550_0[1]),.doutc(w_n15550_0[2]),.din(n15550));
	jspl jspl_w_n15551_0(.douta(w_n15551_0[0]),.doutb(w_n15551_0[1]),.din(n15551));
	jspl3 jspl3_w_n15555_0(.douta(w_n15555_0[0]),.doutb(w_n15555_0[1]),.doutc(w_n15555_0[2]),.din(n15555));
	jspl3 jspl3_w_n15557_0(.douta(w_n15557_0[0]),.doutb(w_n15557_0[1]),.doutc(w_n15557_0[2]),.din(n15557));
	jspl jspl_w_n15558_0(.douta(w_n15558_0[0]),.doutb(w_n15558_0[1]),.din(n15558));
	jspl3 jspl3_w_n15562_0(.douta(w_n15562_0[0]),.doutb(w_n15562_0[1]),.doutc(w_n15562_0[2]),.din(n15562));
	jspl3 jspl3_w_n15564_0(.douta(w_n15564_0[0]),.doutb(w_n15564_0[1]),.doutc(w_n15564_0[2]),.din(n15564));
	jspl jspl_w_n15565_0(.douta(w_n15565_0[0]),.doutb(w_n15565_0[1]),.din(n15565));
	jspl3 jspl3_w_n15569_0(.douta(w_n15569_0[0]),.doutb(w_n15569_0[1]),.doutc(w_n15569_0[2]),.din(n15569));
	jspl3 jspl3_w_n15571_0(.douta(w_n15571_0[0]),.doutb(w_n15571_0[1]),.doutc(w_n15571_0[2]),.din(n15571));
	jspl jspl_w_n15572_0(.douta(w_n15572_0[0]),.doutb(w_n15572_0[1]),.din(n15572));
	jspl3 jspl3_w_n15576_0(.douta(w_n15576_0[0]),.doutb(w_n15576_0[1]),.doutc(w_n15576_0[2]),.din(n15576));
	jspl3 jspl3_w_n15579_0(.douta(w_n15579_0[0]),.doutb(w_n15579_0[1]),.doutc(w_n15579_0[2]),.din(n15579));
	jspl jspl_w_n15580_0(.douta(w_n15580_0[0]),.doutb(w_n15580_0[1]),.din(n15580));
	jspl3 jspl3_w_n15584_0(.douta(w_n15584_0[0]),.doutb(w_n15584_0[1]),.doutc(w_n15584_0[2]),.din(n15584));
	jspl3 jspl3_w_n15586_0(.douta(w_n15586_0[0]),.doutb(w_n15586_0[1]),.doutc(w_n15586_0[2]),.din(n15586));
	jspl jspl_w_n15587_0(.douta(w_n15587_0[0]),.doutb(w_n15587_0[1]),.din(n15587));
	jspl3 jspl3_w_n15591_0(.douta(w_n15591_0[0]),.doutb(w_n15591_0[1]),.doutc(w_n15591_0[2]),.din(n15591));
	jspl3 jspl3_w_n15594_0(.douta(w_n15594_0[0]),.doutb(w_n15594_0[1]),.doutc(w_n15594_0[2]),.din(n15594));
	jspl jspl_w_n15595_0(.douta(w_n15595_0[0]),.doutb(w_n15595_0[1]),.din(n15595));
	jspl3 jspl3_w_n15599_0(.douta(w_n15599_0[0]),.doutb(w_n15599_0[1]),.doutc(w_n15599_0[2]),.din(n15599));
	jspl3 jspl3_w_n15601_0(.douta(w_n15601_0[0]),.doutb(w_n15601_0[1]),.doutc(w_n15601_0[2]),.din(n15601));
	jspl jspl_w_n15602_0(.douta(w_n15602_0[0]),.doutb(w_n15602_0[1]),.din(n15602));
	jspl3 jspl3_w_n15606_0(.douta(w_n15606_0[0]),.doutb(w_n15606_0[1]),.doutc(w_n15606_0[2]),.din(n15606));
	jspl3 jspl3_w_n15609_0(.douta(w_n15609_0[0]),.doutb(w_n15609_0[1]),.doutc(w_n15609_0[2]),.din(n15609));
	jspl jspl_w_n15610_0(.douta(w_n15610_0[0]),.doutb(w_n15610_0[1]),.din(n15610));
	jspl3 jspl3_w_n15614_0(.douta(w_n15614_0[0]),.doutb(w_n15614_0[1]),.doutc(w_n15614_0[2]),.din(n15614));
	jspl3 jspl3_w_n15616_0(.douta(w_n15616_0[0]),.doutb(w_n15616_0[1]),.doutc(w_n15616_0[2]),.din(n15616));
	jspl jspl_w_n15617_0(.douta(w_n15617_0[0]),.doutb(w_n15617_0[1]),.din(n15617));
	jspl jspl_w_n15621_0(.douta(w_n15621_0[0]),.doutb(w_n15621_0[1]),.din(n15621));
	jspl jspl_w_n15622_0(.douta(w_n15622_0[0]),.doutb(w_n15622_0[1]),.din(n15622));
	jspl3 jspl3_w_n15624_0(.douta(w_n15624_0[0]),.doutb(w_n15624_0[1]),.doutc(w_n15624_0[2]),.din(n15624));
	jspl jspl_w_n15625_0(.douta(w_n15625_0[0]),.doutb(w_n15625_0[1]),.din(n15625));
	jspl jspl_w_n15626_0(.douta(w_n15626_0[0]),.doutb(w_n15626_0[1]),.din(n15626));
	jspl3 jspl3_w_n15631_0(.douta(w_n15631_0[0]),.doutb(w_n15631_0[1]),.doutc(w_n15631_0[2]),.din(n15631));
	jspl jspl_w_n15636_0(.douta(w_n15636_0[0]),.doutb(w_n15636_0[1]),.din(n15636));
	jspl jspl_w_n15639_0(.douta(w_n15639_0[0]),.doutb(w_n15639_0[1]),.din(n15639));
	jspl3 jspl3_w_n15642_0(.douta(w_n15642_0[0]),.doutb(w_n15642_0[1]),.doutc(w_n15642_0[2]),.din(n15642));
	jspl jspl_w_n15642_1(.douta(w_n15642_1[0]),.doutb(w_n15642_1[1]),.din(w_n15642_0[0]));
	jspl jspl_w_n15643_0(.douta(w_n15643_0[0]),.doutb(w_n15643_0[1]),.din(n15643));
	jspl3 jspl3_w_n15644_0(.douta(w_n15644_0[0]),.doutb(w_n15644_0[1]),.doutc(w_n15644_0[2]),.din(n15644));
	jspl jspl_w_n15645_0(.douta(w_n15645_0[0]),.doutb(w_n15645_0[1]),.din(n15645));
	jspl3 jspl3_w_n15646_0(.douta(w_n15646_0[0]),.doutb(w_n15646_0[1]),.doutc(w_n15646_0[2]),.din(n15646));
	jspl jspl_w_n15647_0(.douta(w_n15647_0[0]),.doutb(w_n15647_0[1]),.din(n15647));
	jspl jspl_w_n15704_0(.douta(w_n15704_0[0]),.doutb(w_n15704_0[1]),.din(n15704));
	jspl jspl_w_n15708_0(.douta(w_n15708_0[0]),.doutb(w_n15708_0[1]),.din(n15708));
	jspl jspl_w_n15872_0(.douta(w_n15872_0[0]),.doutb(w_n15872_0[1]),.din(n15872));
	jspl jspl_w_n15876_0(.douta(w_n15876_0[0]),.doutb(w_n15876_0[1]),.din(n15876));
	jspl3 jspl3_w_n15878_0(.douta(w_n15878_0[0]),.doutb(w_n15878_0[1]),.doutc(w_n15878_0[2]),.din(n15878));
	jspl3 jspl3_w_n15878_1(.douta(w_n15878_1[0]),.doutb(w_n15878_1[1]),.doutc(w_n15878_1[2]),.din(w_n15878_0[0]));
	jspl3 jspl3_w_n15878_2(.douta(w_n15878_2[0]),.doutb(w_n15878_2[1]),.doutc(w_n15878_2[2]),.din(w_n15878_0[1]));
	jspl3 jspl3_w_n15878_3(.douta(w_n15878_3[0]),.doutb(w_n15878_3[1]),.doutc(w_n15878_3[2]),.din(w_n15878_0[2]));
	jspl3 jspl3_w_n15878_4(.douta(w_n15878_4[0]),.doutb(w_n15878_4[1]),.doutc(w_n15878_4[2]),.din(w_n15878_1[0]));
	jspl3 jspl3_w_n15878_5(.douta(w_n15878_5[0]),.doutb(w_n15878_5[1]),.doutc(w_n15878_5[2]),.din(w_n15878_1[1]));
	jspl3 jspl3_w_n15878_6(.douta(w_n15878_6[0]),.doutb(w_n15878_6[1]),.doutc(w_n15878_6[2]),.din(w_n15878_1[2]));
	jspl3 jspl3_w_n15878_7(.douta(w_n15878_7[0]),.doutb(w_n15878_7[1]),.doutc(w_n15878_7[2]),.din(w_n15878_2[0]));
	jspl3 jspl3_w_n15878_8(.douta(w_n15878_8[0]),.doutb(w_n15878_8[1]),.doutc(w_n15878_8[2]),.din(w_n15878_2[1]));
	jspl3 jspl3_w_n15878_9(.douta(w_n15878_9[0]),.doutb(w_n15878_9[1]),.doutc(w_n15878_9[2]),.din(w_n15878_2[2]));
	jspl3 jspl3_w_n15878_10(.douta(w_n15878_10[0]),.doutb(w_n15878_10[1]),.doutc(w_n15878_10[2]),.din(w_n15878_3[0]));
	jspl3 jspl3_w_n15878_11(.douta(w_n15878_11[0]),.doutb(w_n15878_11[1]),.doutc(w_n15878_11[2]),.din(w_n15878_3[1]));
	jspl3 jspl3_w_n15878_12(.douta(w_n15878_12[0]),.doutb(w_n15878_12[1]),.doutc(w_n15878_12[2]),.din(w_n15878_3[2]));
	jspl3 jspl3_w_n15878_13(.douta(w_n15878_13[0]),.doutb(w_n15878_13[1]),.doutc(w_n15878_13[2]),.din(w_n15878_4[0]));
	jspl3 jspl3_w_n15878_14(.douta(w_n15878_14[0]),.doutb(w_n15878_14[1]),.doutc(w_n15878_14[2]),.din(w_n15878_4[1]));
	jspl3 jspl3_w_n15878_15(.douta(w_n15878_15[0]),.doutb(w_n15878_15[1]),.doutc(w_n15878_15[2]),.din(w_n15878_4[2]));
	jspl3 jspl3_w_n15878_16(.douta(w_n15878_16[0]),.doutb(w_n15878_16[1]),.doutc(w_n15878_16[2]),.din(w_n15878_5[0]));
	jspl3 jspl3_w_n15878_17(.douta(w_n15878_17[0]),.doutb(w_n15878_17[1]),.doutc(w_n15878_17[2]),.din(w_n15878_5[1]));
	jspl jspl_w_n15878_18(.douta(w_n15878_18[0]),.doutb(w_n15878_18[1]),.din(w_n15878_5[2]));
	jspl3 jspl3_w_n15882_0(.douta(w_n15882_0[0]),.doutb(w_n15882_0[1]),.doutc(w_n15882_0[2]),.din(n15882));
	jspl jspl_w_n15883_0(.douta(w_n15883_0[0]),.doutb(w_n15883_0[1]),.din(n15883));
	jspl jspl_w_n15885_0(.douta(w_n15885_0[0]),.doutb(w_n15885_0[1]),.din(n15885));
	jspl jspl_w_n15886_0(.douta(w_n15886_0[0]),.doutb(w_n15886_0[1]),.din(n15886));
	jspl jspl_w_n15891_0(.douta(w_n15891_0[0]),.doutb(w_n15891_0[1]),.din(n15891));
	jspl jspl_w_n15892_0(.douta(w_n15892_0[0]),.doutb(w_n15892_0[1]),.din(n15892));
	jspl3 jspl3_w_n15894_0(.douta(w_n15894_0[0]),.doutb(w_n15894_0[1]),.doutc(w_n15894_0[2]),.din(n15894));
	jspl jspl_w_n15895_0(.douta(w_n15895_0[0]),.doutb(w_n15895_0[1]),.din(n15895));
	jspl3 jspl3_w_n15899_0(.douta(w_n15899_0[0]),.doutb(w_n15899_0[1]),.doutc(w_n15899_0[2]),.din(n15899));
	jspl3 jspl3_w_n15901_0(.douta(w_n15901_0[0]),.doutb(w_n15901_0[1]),.doutc(w_n15901_0[2]),.din(n15901));
	jspl jspl_w_n15902_0(.douta(w_n15902_0[0]),.doutb(w_n15902_0[1]),.din(n15902));
	jspl jspl_w_n15906_0(.douta(w_n15906_0[0]),.doutb(w_n15906_0[1]),.din(n15906));
	jspl3 jspl3_w_n15908_0(.douta(w_n15908_0[0]),.doutb(w_n15908_0[1]),.doutc(w_n15908_0[2]),.din(n15908));
	jspl jspl_w_n15909_0(.douta(w_n15909_0[0]),.doutb(w_n15909_0[1]),.din(n15909));
	jspl jspl_w_n15913_0(.douta(w_n15913_0[0]),.doutb(w_n15913_0[1]),.din(n15913));
	jspl3 jspl3_w_n15915_0(.douta(w_n15915_0[0]),.doutb(w_n15915_0[1]),.doutc(w_n15915_0[2]),.din(n15915));
	jspl jspl_w_n15916_0(.douta(w_n15916_0[0]),.doutb(w_n15916_0[1]),.din(n15916));
	jspl jspl_w_n15920_0(.douta(w_n15920_0[0]),.doutb(w_n15920_0[1]),.din(n15920));
	jspl jspl_w_n15921_0(.douta(w_n15921_0[0]),.doutb(w_n15921_0[1]),.din(n15921));
	jspl3 jspl3_w_n15923_0(.douta(w_n15923_0[0]),.doutb(w_n15923_0[1]),.doutc(w_n15923_0[2]),.din(n15923));
	jspl jspl_w_n15924_0(.douta(w_n15924_0[0]),.doutb(w_n15924_0[1]),.din(n15924));
	jspl jspl_w_n15928_0(.douta(w_n15928_0[0]),.doutb(w_n15928_0[1]),.din(n15928));
	jspl3 jspl3_w_n15930_0(.douta(w_n15930_0[0]),.doutb(w_n15930_0[1]),.doutc(w_n15930_0[2]),.din(n15930));
	jspl jspl_w_n15931_0(.douta(w_n15931_0[0]),.doutb(w_n15931_0[1]),.din(n15931));
	jspl jspl_w_n15935_0(.douta(w_n15935_0[0]),.doutb(w_n15935_0[1]),.din(n15935));
	jspl jspl_w_n15936_0(.douta(w_n15936_0[0]),.doutb(w_n15936_0[1]),.din(n15936));
	jspl3 jspl3_w_n15938_0(.douta(w_n15938_0[0]),.doutb(w_n15938_0[1]),.doutc(w_n15938_0[2]),.din(n15938));
	jspl jspl_w_n15939_0(.douta(w_n15939_0[0]),.doutb(w_n15939_0[1]),.din(n15939));
	jspl jspl_w_n15943_0(.douta(w_n15943_0[0]),.doutb(w_n15943_0[1]),.din(n15943));
	jspl3 jspl3_w_n15945_0(.douta(w_n15945_0[0]),.doutb(w_n15945_0[1]),.doutc(w_n15945_0[2]),.din(n15945));
	jspl jspl_w_n15946_0(.douta(w_n15946_0[0]),.doutb(w_n15946_0[1]),.din(n15946));
	jspl jspl_w_n15950_0(.douta(w_n15950_0[0]),.doutb(w_n15950_0[1]),.din(n15950));
	jspl jspl_w_n15951_0(.douta(w_n15951_0[0]),.doutb(w_n15951_0[1]),.din(n15951));
	jspl3 jspl3_w_n15953_0(.douta(w_n15953_0[0]),.doutb(w_n15953_0[1]),.doutc(w_n15953_0[2]),.din(n15953));
	jspl jspl_w_n15954_0(.douta(w_n15954_0[0]),.doutb(w_n15954_0[1]),.din(n15954));
	jspl jspl_w_n15958_0(.douta(w_n15958_0[0]),.doutb(w_n15958_0[1]),.din(n15958));
	jspl jspl_w_n15959_0(.douta(w_n15959_0[0]),.doutb(w_n15959_0[1]),.din(n15959));
	jspl3 jspl3_w_n15961_0(.douta(w_n15961_0[0]),.doutb(w_n15961_0[1]),.doutc(w_n15961_0[2]),.din(n15961));
	jspl jspl_w_n15962_0(.douta(w_n15962_0[0]),.doutb(w_n15962_0[1]),.din(n15962));
	jspl jspl_w_n15966_0(.douta(w_n15966_0[0]),.doutb(w_n15966_0[1]),.din(n15966));
	jspl jspl_w_n15967_0(.douta(w_n15967_0[0]),.doutb(w_n15967_0[1]),.din(n15967));
	jspl3 jspl3_w_n15969_0(.douta(w_n15969_0[0]),.doutb(w_n15969_0[1]),.doutc(w_n15969_0[2]),.din(n15969));
	jspl jspl_w_n15970_0(.douta(w_n15970_0[0]),.doutb(w_n15970_0[1]),.din(n15970));
	jspl jspl_w_n15974_0(.douta(w_n15974_0[0]),.doutb(w_n15974_0[1]),.din(n15974));
	jspl3 jspl3_w_n15976_0(.douta(w_n15976_0[0]),.doutb(w_n15976_0[1]),.doutc(w_n15976_0[2]),.din(n15976));
	jspl jspl_w_n15977_0(.douta(w_n15977_0[0]),.doutb(w_n15977_0[1]),.din(n15977));
	jspl jspl_w_n15981_0(.douta(w_n15981_0[0]),.doutb(w_n15981_0[1]),.din(n15981));
	jspl jspl_w_n15982_0(.douta(w_n15982_0[0]),.doutb(w_n15982_0[1]),.din(n15982));
	jspl3 jspl3_w_n15984_0(.douta(w_n15984_0[0]),.doutb(w_n15984_0[1]),.doutc(w_n15984_0[2]),.din(n15984));
	jspl jspl_w_n15985_0(.douta(w_n15985_0[0]),.doutb(w_n15985_0[1]),.din(n15985));
	jspl jspl_w_n15989_0(.douta(w_n15989_0[0]),.doutb(w_n15989_0[1]),.din(n15989));
	jspl3 jspl3_w_n15991_0(.douta(w_n15991_0[0]),.doutb(w_n15991_0[1]),.doutc(w_n15991_0[2]),.din(n15991));
	jspl jspl_w_n15992_0(.douta(w_n15992_0[0]),.doutb(w_n15992_0[1]),.din(n15992));
	jspl jspl_w_n15996_0(.douta(w_n15996_0[0]),.doutb(w_n15996_0[1]),.din(n15996));
	jspl jspl_w_n15997_0(.douta(w_n15997_0[0]),.doutb(w_n15997_0[1]),.din(n15997));
	jspl3 jspl3_w_n15999_0(.douta(w_n15999_0[0]),.doutb(w_n15999_0[1]),.doutc(w_n15999_0[2]),.din(n15999));
	jspl jspl_w_n16000_0(.douta(w_n16000_0[0]),.doutb(w_n16000_0[1]),.din(n16000));
	jspl jspl_w_n16004_0(.douta(w_n16004_0[0]),.doutb(w_n16004_0[1]),.din(n16004));
	jspl3 jspl3_w_n16006_0(.douta(w_n16006_0[0]),.doutb(w_n16006_0[1]),.doutc(w_n16006_0[2]),.din(n16006));
	jspl jspl_w_n16007_0(.douta(w_n16007_0[0]),.doutb(w_n16007_0[1]),.din(n16007));
	jspl jspl_w_n16011_0(.douta(w_n16011_0[0]),.doutb(w_n16011_0[1]),.din(n16011));
	jspl jspl_w_n16012_0(.douta(w_n16012_0[0]),.doutb(w_n16012_0[1]),.din(n16012));
	jspl3 jspl3_w_n16014_0(.douta(w_n16014_0[0]),.doutb(w_n16014_0[1]),.doutc(w_n16014_0[2]),.din(n16014));
	jspl jspl_w_n16015_0(.douta(w_n16015_0[0]),.doutb(w_n16015_0[1]),.din(n16015));
	jspl jspl_w_n16019_0(.douta(w_n16019_0[0]),.doutb(w_n16019_0[1]),.din(n16019));
	jspl3 jspl3_w_n16021_0(.douta(w_n16021_0[0]),.doutb(w_n16021_0[1]),.doutc(w_n16021_0[2]),.din(n16021));
	jspl jspl_w_n16022_0(.douta(w_n16022_0[0]),.doutb(w_n16022_0[1]),.din(n16022));
	jspl jspl_w_n16026_0(.douta(w_n16026_0[0]),.doutb(w_n16026_0[1]),.din(n16026));
	jspl jspl_w_n16027_0(.douta(w_n16027_0[0]),.doutb(w_n16027_0[1]),.din(n16027));
	jspl3 jspl3_w_n16029_0(.douta(w_n16029_0[0]),.doutb(w_n16029_0[1]),.doutc(w_n16029_0[2]),.din(n16029));
	jspl jspl_w_n16030_0(.douta(w_n16030_0[0]),.doutb(w_n16030_0[1]),.din(n16030));
	jspl jspl_w_n16034_0(.douta(w_n16034_0[0]),.doutb(w_n16034_0[1]),.din(n16034));
	jspl jspl_w_n16035_0(.douta(w_n16035_0[0]),.doutb(w_n16035_0[1]),.din(n16035));
	jspl3 jspl3_w_n16037_0(.douta(w_n16037_0[0]),.doutb(w_n16037_0[1]),.doutc(w_n16037_0[2]),.din(n16037));
	jspl jspl_w_n16038_0(.douta(w_n16038_0[0]),.doutb(w_n16038_0[1]),.din(n16038));
	jspl jspl_w_n16042_0(.douta(w_n16042_0[0]),.doutb(w_n16042_0[1]),.din(n16042));
	jspl jspl_w_n16043_0(.douta(w_n16043_0[0]),.doutb(w_n16043_0[1]),.din(n16043));
	jspl3 jspl3_w_n16045_0(.douta(w_n16045_0[0]),.doutb(w_n16045_0[1]),.doutc(w_n16045_0[2]),.din(n16045));
	jspl jspl_w_n16046_0(.douta(w_n16046_0[0]),.doutb(w_n16046_0[1]),.din(n16046));
	jspl jspl_w_n16050_0(.douta(w_n16050_0[0]),.doutb(w_n16050_0[1]),.din(n16050));
	jspl3 jspl3_w_n16052_0(.douta(w_n16052_0[0]),.doutb(w_n16052_0[1]),.doutc(w_n16052_0[2]),.din(n16052));
	jspl jspl_w_n16053_0(.douta(w_n16053_0[0]),.doutb(w_n16053_0[1]),.din(n16053));
	jspl jspl_w_n16057_0(.douta(w_n16057_0[0]),.doutb(w_n16057_0[1]),.din(n16057));
	jspl jspl_w_n16058_0(.douta(w_n16058_0[0]),.doutb(w_n16058_0[1]),.din(n16058));
	jspl3 jspl3_w_n16060_0(.douta(w_n16060_0[0]),.doutb(w_n16060_0[1]),.doutc(w_n16060_0[2]),.din(n16060));
	jspl jspl_w_n16061_0(.douta(w_n16061_0[0]),.doutb(w_n16061_0[1]),.din(n16061));
	jspl jspl_w_n16065_0(.douta(w_n16065_0[0]),.doutb(w_n16065_0[1]),.din(n16065));
	jspl3 jspl3_w_n16067_0(.douta(w_n16067_0[0]),.doutb(w_n16067_0[1]),.doutc(w_n16067_0[2]),.din(n16067));
	jspl jspl_w_n16068_0(.douta(w_n16068_0[0]),.doutb(w_n16068_0[1]),.din(n16068));
	jspl jspl_w_n16072_0(.douta(w_n16072_0[0]),.doutb(w_n16072_0[1]),.din(n16072));
	jspl jspl_w_n16073_0(.douta(w_n16073_0[0]),.doutb(w_n16073_0[1]),.din(n16073));
	jspl3 jspl3_w_n16075_0(.douta(w_n16075_0[0]),.doutb(w_n16075_0[1]),.doutc(w_n16075_0[2]),.din(n16075));
	jspl jspl_w_n16076_0(.douta(w_n16076_0[0]),.doutb(w_n16076_0[1]),.din(n16076));
	jspl jspl_w_n16080_0(.douta(w_n16080_0[0]),.doutb(w_n16080_0[1]),.din(n16080));
	jspl jspl_w_n16081_0(.douta(w_n16081_0[0]),.doutb(w_n16081_0[1]),.din(n16081));
	jspl3 jspl3_w_n16083_0(.douta(w_n16083_0[0]),.doutb(w_n16083_0[1]),.doutc(w_n16083_0[2]),.din(n16083));
	jspl jspl_w_n16084_0(.douta(w_n16084_0[0]),.doutb(w_n16084_0[1]),.din(n16084));
	jspl jspl_w_n16088_0(.douta(w_n16088_0[0]),.doutb(w_n16088_0[1]),.din(n16088));
	jspl jspl_w_n16089_0(.douta(w_n16089_0[0]),.doutb(w_n16089_0[1]),.din(n16089));
	jspl3 jspl3_w_n16091_0(.douta(w_n16091_0[0]),.doutb(w_n16091_0[1]),.doutc(w_n16091_0[2]),.din(n16091));
	jspl jspl_w_n16092_0(.douta(w_n16092_0[0]),.doutb(w_n16092_0[1]),.din(n16092));
	jspl jspl_w_n16096_0(.douta(w_n16096_0[0]),.doutb(w_n16096_0[1]),.din(n16096));
	jspl3 jspl3_w_n16098_0(.douta(w_n16098_0[0]),.doutb(w_n16098_0[1]),.doutc(w_n16098_0[2]),.din(n16098));
	jspl jspl_w_n16099_0(.douta(w_n16099_0[0]),.doutb(w_n16099_0[1]),.din(n16099));
	jspl jspl_w_n16103_0(.douta(w_n16103_0[0]),.doutb(w_n16103_0[1]),.din(n16103));
	jspl jspl_w_n16104_0(.douta(w_n16104_0[0]),.doutb(w_n16104_0[1]),.din(n16104));
	jspl3 jspl3_w_n16106_0(.douta(w_n16106_0[0]),.doutb(w_n16106_0[1]),.doutc(w_n16106_0[2]),.din(n16106));
	jspl jspl_w_n16107_0(.douta(w_n16107_0[0]),.doutb(w_n16107_0[1]),.din(n16107));
	jspl jspl_w_n16111_0(.douta(w_n16111_0[0]),.doutb(w_n16111_0[1]),.din(n16111));
	jspl3 jspl3_w_n16113_0(.douta(w_n16113_0[0]),.doutb(w_n16113_0[1]),.doutc(w_n16113_0[2]),.din(n16113));
	jspl jspl_w_n16114_0(.douta(w_n16114_0[0]),.doutb(w_n16114_0[1]),.din(n16114));
	jspl jspl_w_n16118_0(.douta(w_n16118_0[0]),.doutb(w_n16118_0[1]),.din(n16118));
	jspl jspl_w_n16119_0(.douta(w_n16119_0[0]),.doutb(w_n16119_0[1]),.din(n16119));
	jspl3 jspl3_w_n16121_0(.douta(w_n16121_0[0]),.doutb(w_n16121_0[1]),.doutc(w_n16121_0[2]),.din(n16121));
	jspl jspl_w_n16122_0(.douta(w_n16122_0[0]),.doutb(w_n16122_0[1]),.din(n16122));
	jspl jspl_w_n16126_0(.douta(w_n16126_0[0]),.doutb(w_n16126_0[1]),.din(n16126));
	jspl jspl_w_n16127_0(.douta(w_n16127_0[0]),.doutb(w_n16127_0[1]),.din(n16127));
	jspl3 jspl3_w_n16129_0(.douta(w_n16129_0[0]),.doutb(w_n16129_0[1]),.doutc(w_n16129_0[2]),.din(n16129));
	jspl jspl_w_n16130_0(.douta(w_n16130_0[0]),.doutb(w_n16130_0[1]),.din(n16130));
	jspl jspl_w_n16134_0(.douta(w_n16134_0[0]),.doutb(w_n16134_0[1]),.din(n16134));
	jspl3 jspl3_w_n16136_0(.douta(w_n16136_0[0]),.doutb(w_n16136_0[1]),.doutc(w_n16136_0[2]),.din(n16136));
	jspl jspl_w_n16137_0(.douta(w_n16137_0[0]),.doutb(w_n16137_0[1]),.din(n16137));
	jspl jspl_w_n16140_0(.douta(w_n16140_0[0]),.doutb(w_n16140_0[1]),.din(n16140));
	jspl3 jspl3_w_n16143_0(.douta(w_n16143_0[0]),.doutb(w_n16143_0[1]),.doutc(w_n16143_0[2]),.din(n16143));
	jspl jspl_w_n16144_0(.douta(w_n16144_0[0]),.doutb(w_n16144_0[1]),.din(n16144));
	jspl jspl_w_n16148_0(.douta(w_n16148_0[0]),.doutb(w_n16148_0[1]),.din(n16148));
	jspl jspl_w_n16149_0(.douta(w_n16149_0[0]),.doutb(w_n16149_0[1]),.din(n16149));
	jspl3 jspl3_w_n16151_0(.douta(w_n16151_0[0]),.doutb(w_n16151_0[1]),.doutc(w_n16151_0[2]),.din(n16151));
	jspl jspl_w_n16152_0(.douta(w_n16152_0[0]),.doutb(w_n16152_0[1]),.din(n16152));
	jspl jspl_w_n16156_0(.douta(w_n16156_0[0]),.doutb(w_n16156_0[1]),.din(n16156));
	jspl3 jspl3_w_n16158_0(.douta(w_n16158_0[0]),.doutb(w_n16158_0[1]),.doutc(w_n16158_0[2]),.din(n16158));
	jspl jspl_w_n16159_0(.douta(w_n16159_0[0]),.doutb(w_n16159_0[1]),.din(n16159));
	jspl jspl_w_n16163_0(.douta(w_n16163_0[0]),.doutb(w_n16163_0[1]),.din(n16163));
	jspl jspl_w_n16164_0(.douta(w_n16164_0[0]),.doutb(w_n16164_0[1]),.din(n16164));
	jspl3 jspl3_w_n16166_0(.douta(w_n16166_0[0]),.doutb(w_n16166_0[1]),.doutc(w_n16166_0[2]),.din(n16166));
	jspl jspl_w_n16167_0(.douta(w_n16167_0[0]),.doutb(w_n16167_0[1]),.din(n16167));
	jspl jspl_w_n16171_0(.douta(w_n16171_0[0]),.doutb(w_n16171_0[1]),.din(n16171));
	jspl3 jspl3_w_n16173_0(.douta(w_n16173_0[0]),.doutb(w_n16173_0[1]),.doutc(w_n16173_0[2]),.din(n16173));
	jspl jspl_w_n16174_0(.douta(w_n16174_0[0]),.doutb(w_n16174_0[1]),.din(n16174));
	jspl jspl_w_n16178_0(.douta(w_n16178_0[0]),.doutb(w_n16178_0[1]),.din(n16178));
	jspl jspl_w_n16179_0(.douta(w_n16179_0[0]),.doutb(w_n16179_0[1]),.din(n16179));
	jspl3 jspl3_w_n16181_0(.douta(w_n16181_0[0]),.doutb(w_n16181_0[1]),.doutc(w_n16181_0[2]),.din(n16181));
	jspl jspl_w_n16182_0(.douta(w_n16182_0[0]),.doutb(w_n16182_0[1]),.din(n16182));
	jspl jspl_w_n16186_0(.douta(w_n16186_0[0]),.doutb(w_n16186_0[1]),.din(n16186));
	jspl jspl_w_n16187_0(.douta(w_n16187_0[0]),.doutb(w_n16187_0[1]),.din(n16187));
	jspl3 jspl3_w_n16189_0(.douta(w_n16189_0[0]),.doutb(w_n16189_0[1]),.doutc(w_n16189_0[2]),.din(n16189));
	jspl jspl_w_n16190_0(.douta(w_n16190_0[0]),.doutb(w_n16190_0[1]),.din(n16190));
	jspl jspl_w_n16194_0(.douta(w_n16194_0[0]),.doutb(w_n16194_0[1]),.din(n16194));
	jspl jspl_w_n16195_0(.douta(w_n16195_0[0]),.doutb(w_n16195_0[1]),.din(n16195));
	jspl3 jspl3_w_n16197_0(.douta(w_n16197_0[0]),.doutb(w_n16197_0[1]),.doutc(w_n16197_0[2]),.din(n16197));
	jspl jspl_w_n16198_0(.douta(w_n16198_0[0]),.doutb(w_n16198_0[1]),.din(n16198));
	jspl jspl_w_n16202_0(.douta(w_n16202_0[0]),.doutb(w_n16202_0[1]),.din(n16202));
	jspl3 jspl3_w_n16204_0(.douta(w_n16204_0[0]),.doutb(w_n16204_0[1]),.doutc(w_n16204_0[2]),.din(n16204));
	jspl jspl_w_n16205_0(.douta(w_n16205_0[0]),.doutb(w_n16205_0[1]),.din(n16205));
	jspl jspl_w_n16209_0(.douta(w_n16209_0[0]),.doutb(w_n16209_0[1]),.din(n16209));
	jspl jspl_w_n16210_0(.douta(w_n16210_0[0]),.doutb(w_n16210_0[1]),.din(n16210));
	jspl3 jspl3_w_n16212_0(.douta(w_n16212_0[0]),.doutb(w_n16212_0[1]),.doutc(w_n16212_0[2]),.din(n16212));
	jspl jspl_w_n16213_0(.douta(w_n16213_0[0]),.doutb(w_n16213_0[1]),.din(n16213));
	jspl jspl_w_n16217_0(.douta(w_n16217_0[0]),.doutb(w_n16217_0[1]),.din(n16217));
	jspl3 jspl3_w_n16219_0(.douta(w_n16219_0[0]),.doutb(w_n16219_0[1]),.doutc(w_n16219_0[2]),.din(n16219));
	jspl jspl_w_n16220_0(.douta(w_n16220_0[0]),.doutb(w_n16220_0[1]),.din(n16220));
	jspl jspl_w_n16224_0(.douta(w_n16224_0[0]),.doutb(w_n16224_0[1]),.din(n16224));
	jspl jspl_w_n16225_0(.douta(w_n16225_0[0]),.doutb(w_n16225_0[1]),.din(n16225));
	jspl3 jspl3_w_n16227_0(.douta(w_n16227_0[0]),.doutb(w_n16227_0[1]),.doutc(w_n16227_0[2]),.din(n16227));
	jspl jspl_w_n16228_0(.douta(w_n16228_0[0]),.doutb(w_n16228_0[1]),.din(n16228));
	jspl jspl_w_n16232_0(.douta(w_n16232_0[0]),.doutb(w_n16232_0[1]),.din(n16232));
	jspl3 jspl3_w_n16234_0(.douta(w_n16234_0[0]),.doutb(w_n16234_0[1]),.doutc(w_n16234_0[2]),.din(n16234));
	jspl jspl_w_n16235_0(.douta(w_n16235_0[0]),.doutb(w_n16235_0[1]),.din(n16235));
	jspl jspl_w_n16250_0(.douta(w_n16250_0[0]),.doutb(w_n16250_0[1]),.din(n16250));
	jspl jspl_w_n16291_0(.douta(w_n16291_0[0]),.doutb(w_n16291_0[1]),.din(n16291));
	jspl jspl_w_n16302_0(.douta(w_n16302_0[0]),.doutb(w_n16302_0[1]),.din(n16302));
	jspl jspl_w_n16306_0(.douta(w_n16306_0[0]),.doutb(w_n16306_0[1]),.din(n16306));
	jspl jspl_w_n16313_0(.douta(w_n16313_0[0]),.doutb(w_n16313_0[1]),.din(n16313));
	jspl jspl_w_n16320_0(.douta(w_n16320_0[0]),.doutb(w_n16320_0[1]),.din(n16320));
	jspl jspl_w_n16333_0(.douta(w_n16333_0[0]),.doutb(w_n16333_0[1]),.din(n16333));
	jspl jspl_w_n16340_0(.douta(w_n16340_0[0]),.doutb(w_n16340_0[1]),.din(n16340));
	jspl jspl_w_n16347_0(.douta(w_n16347_0[0]),.doutb(w_n16347_0[1]),.din(n16347));
	jspl jspl_w_n16354_0(.douta(w_n16354_0[0]),.doutb(w_n16354_0[1]),.din(n16354));
	jspl jspl_w_n16367_0(.douta(w_n16367_0[0]),.doutb(w_n16367_0[1]),.din(n16367));
	jspl jspl_w_n16374_0(.douta(w_n16374_0[0]),.doutb(w_n16374_0[1]),.din(n16374));
	jspl jspl_w_n16387_0(.douta(w_n16387_0[0]),.doutb(w_n16387_0[1]),.din(n16387));
	jspl jspl_w_n16394_0(.douta(w_n16394_0[0]),.doutb(w_n16394_0[1]),.din(n16394));
	jspl jspl_w_n16404_0(.douta(w_n16404_0[0]),.doutb(w_n16404_0[1]),.din(n16404));
	jspl jspl_w_n16414_0(.douta(w_n16414_0[0]),.doutb(w_n16414_0[1]),.din(n16414));
	jspl jspl_w_n16421_0(.douta(w_n16421_0[0]),.doutb(w_n16421_0[1]),.din(n16421));
	jspl jspl_w_n16434_0(.douta(w_n16434_0[0]),.doutb(w_n16434_0[1]),.din(n16434));
	jspl jspl_w_n16441_0(.douta(w_n16441_0[0]),.doutb(w_n16441_0[1]),.din(n16441));
	jspl jspl_w_n16448_0(.douta(w_n16448_0[0]),.doutb(w_n16448_0[1]),.din(n16448));
	jspl3 jspl3_w_n16454_0(.douta(w_n16454_0[0]),.doutb(w_n16454_0[1]),.doutc(w_n16454_0[2]),.din(n16454));
	jspl3 jspl3_w_n16456_0(.douta(w_n16456_0[0]),.doutb(w_n16456_0[1]),.doutc(w_n16456_0[2]),.din(n16456));
	jspl3 jspl3_w_n16459_0(.douta(w_n16459_0[0]),.doutb(w_n16459_0[1]),.doutc(w_n16459_0[2]),.din(n16459));
	jspl jspl_w_n16460_0(.douta(w_n16460_0[0]),.doutb(w_n16460_0[1]),.din(n16460));
	jspl jspl_w_n16462_0(.douta(w_n16462_0[0]),.doutb(w_n16462_0[1]),.din(n16462));
	jspl jspl_w_n16464_0(.douta(w_n16464_0[0]),.doutb(w_n16464_0[1]),.din(n16464));
	jspl jspl_w_n16465_0(.douta(w_n16465_0[0]),.doutb(w_n16465_0[1]),.din(n16465));
	jspl3 jspl3_w_n16466_0(.douta(w_n16466_0[0]),.doutb(w_n16466_0[1]),.doutc(w_n16466_0[2]),.din(n16466));
	jspl jspl_w_n16471_0(.douta(w_n16471_0[0]),.doutb(w_n16471_0[1]),.din(n16471));
	jspl jspl_w_n16472_0(.douta(w_n16472_0[0]),.doutb(w_n16472_0[1]),.din(n16472));
	jspl jspl_w_n16478_0(.douta(w_n16478_0[0]),.doutb(w_n16478_0[1]),.din(n16478));
	jspl jspl_w_n16479_0(.douta(w_n16479_0[0]),.doutb(w_n16479_0[1]),.din(n16479));
	jspl jspl_w_n16480_0(.douta(w_n16480_0[0]),.doutb(w_n16480_0[1]),.din(n16480));
	jspl3 jspl3_w_n16485_0(.douta(w_n16485_0[0]),.doutb(w_n16485_0[1]),.doutc(w_n16485_0[2]),.din(n16485));
	jspl3 jspl3_w_n16489_0(.douta(w_n16489_0[0]),.doutb(w_n16489_0[1]),.doutc(w_n16489_0[2]),.din(n16489));
	jspl3 jspl3_w_n16489_1(.douta(w_n16489_1[0]),.doutb(w_n16489_1[1]),.doutc(w_n16489_1[2]),.din(w_n16489_0[0]));
	jspl3 jspl3_w_n16489_2(.douta(w_n16489_2[0]),.doutb(w_n16489_2[1]),.doutc(w_n16489_2[2]),.din(w_n16489_0[1]));
	jspl3 jspl3_w_n16489_3(.douta(w_n16489_3[0]),.doutb(w_n16489_3[1]),.doutc(w_n16489_3[2]),.din(w_n16489_0[2]));
	jspl3 jspl3_w_n16489_4(.douta(w_n16489_4[0]),.doutb(w_n16489_4[1]),.doutc(w_n16489_4[2]),.din(w_n16489_1[0]));
	jspl3 jspl3_w_n16489_5(.douta(w_n16489_5[0]),.doutb(w_n16489_5[1]),.doutc(w_n16489_5[2]),.din(w_n16489_1[1]));
	jspl3 jspl3_w_n16489_6(.douta(w_n16489_6[0]),.doutb(w_n16489_6[1]),.doutc(w_n16489_6[2]),.din(w_n16489_1[2]));
	jspl3 jspl3_w_n16489_7(.douta(w_n16489_7[0]),.doutb(w_n16489_7[1]),.doutc(w_n16489_7[2]),.din(w_n16489_2[0]));
	jspl3 jspl3_w_n16489_8(.douta(w_n16489_8[0]),.doutb(w_n16489_8[1]),.doutc(w_n16489_8[2]),.din(w_n16489_2[1]));
	jspl3 jspl3_w_n16489_9(.douta(w_n16489_9[0]),.doutb(w_n16489_9[1]),.doutc(w_n16489_9[2]),.din(w_n16489_2[2]));
	jspl3 jspl3_w_n16489_10(.douta(w_n16489_10[0]),.doutb(w_n16489_10[1]),.doutc(w_n16489_10[2]),.din(w_n16489_3[0]));
	jspl3 jspl3_w_n16489_11(.douta(w_n16489_11[0]),.doutb(w_n16489_11[1]),.doutc(w_n16489_11[2]),.din(w_n16489_3[1]));
	jspl3 jspl3_w_n16489_12(.douta(w_n16489_12[0]),.doutb(w_n16489_12[1]),.doutc(w_n16489_12[2]),.din(w_n16489_3[2]));
	jspl3 jspl3_w_n16489_13(.douta(w_n16489_13[0]),.doutb(w_n16489_13[1]),.doutc(w_n16489_13[2]),.din(w_n16489_4[0]));
	jspl3 jspl3_w_n16489_14(.douta(w_n16489_14[0]),.doutb(w_n16489_14[1]),.doutc(w_n16489_14[2]),.din(w_n16489_4[1]));
	jspl3 jspl3_w_n16489_15(.douta(w_n16489_15[0]),.doutb(w_n16489_15[1]),.doutc(w_n16489_15[2]),.din(w_n16489_4[2]));
	jspl3 jspl3_w_n16489_16(.douta(w_n16489_16[0]),.doutb(w_n16489_16[1]),.doutc(w_n16489_16[2]),.din(w_n16489_5[0]));
	jspl3 jspl3_w_n16489_17(.douta(w_n16489_17[0]),.doutb(w_n16489_17[1]),.doutc(w_n16489_17[2]),.din(w_n16489_5[1]));
	jspl3 jspl3_w_n16489_18(.douta(w_n16489_18[0]),.doutb(w_n16489_18[1]),.doutc(w_n16489_18[2]),.din(w_n16489_5[2]));
	jspl3 jspl3_w_n16489_19(.douta(w_n16489_19[0]),.doutb(w_n16489_19[1]),.doutc(w_n16489_19[2]),.din(w_n16489_6[0]));
	jspl3 jspl3_w_n16489_20(.douta(w_n16489_20[0]),.doutb(w_n16489_20[1]),.doutc(w_n16489_20[2]),.din(w_n16489_6[1]));
	jspl3 jspl3_w_n16489_21(.douta(w_n16489_21[0]),.doutb(w_n16489_21[1]),.doutc(w_n16489_21[2]),.din(w_n16489_6[2]));
	jspl3 jspl3_w_n16489_22(.douta(w_n16489_22[0]),.doutb(w_n16489_22[1]),.doutc(w_n16489_22[2]),.din(w_n16489_7[0]));
	jspl3 jspl3_w_n16489_23(.douta(w_n16489_23[0]),.doutb(w_n16489_23[1]),.doutc(w_n16489_23[2]),.din(w_n16489_7[1]));
	jspl3 jspl3_w_n16489_24(.douta(w_n16489_24[0]),.doutb(w_n16489_24[1]),.doutc(w_n16489_24[2]),.din(w_n16489_7[2]));
	jspl3 jspl3_w_n16489_25(.douta(w_n16489_25[0]),.doutb(w_n16489_25[1]),.doutc(w_n16489_25[2]),.din(w_n16489_8[0]));
	jspl3 jspl3_w_n16489_26(.douta(w_n16489_26[0]),.doutb(w_n16489_26[1]),.doutc(w_n16489_26[2]),.din(w_n16489_8[1]));
	jspl3 jspl3_w_n16489_27(.douta(w_n16489_27[0]),.doutb(w_n16489_27[1]),.doutc(w_n16489_27[2]),.din(w_n16489_8[2]));
	jspl3 jspl3_w_n16489_28(.douta(w_n16489_28[0]),.doutb(w_n16489_28[1]),.doutc(w_n16489_28[2]),.din(w_n16489_9[0]));
	jspl3 jspl3_w_n16489_29(.douta(w_n16489_29[0]),.doutb(w_n16489_29[1]),.doutc(w_n16489_29[2]),.din(w_n16489_9[1]));
	jspl3 jspl3_w_n16489_30(.douta(w_n16489_30[0]),.doutb(w_n16489_30[1]),.doutc(w_n16489_30[2]),.din(w_n16489_9[2]));
	jspl3 jspl3_w_n16489_31(.douta(w_n16489_31[0]),.doutb(w_n16489_31[1]),.doutc(w_n16489_31[2]),.din(w_n16489_10[0]));
	jspl3 jspl3_w_n16489_32(.douta(w_n16489_32[0]),.doutb(w_n16489_32[1]),.doutc(w_n16489_32[2]),.din(w_n16489_10[1]));
	jspl3 jspl3_w_n16489_33(.douta(w_n16489_33[0]),.doutb(w_n16489_33[1]),.doutc(w_n16489_33[2]),.din(w_n16489_10[2]));
	jspl3 jspl3_w_n16489_34(.douta(w_n16489_34[0]),.doutb(w_n16489_34[1]),.doutc(w_n16489_34[2]),.din(w_n16489_11[0]));
	jspl3 jspl3_w_n16489_35(.douta(w_n16489_35[0]),.doutb(w_n16489_35[1]),.doutc(w_n16489_35[2]),.din(w_n16489_11[1]));
	jspl3 jspl3_w_n16489_36(.douta(w_n16489_36[0]),.doutb(w_n16489_36[1]),.doutc(w_n16489_36[2]),.din(w_n16489_11[2]));
	jspl3 jspl3_w_n16489_37(.douta(w_n16489_37[0]),.doutb(w_n16489_37[1]),.doutc(w_n16489_37[2]),.din(w_n16489_12[0]));
	jspl3 jspl3_w_n16489_38(.douta(w_n16489_38[0]),.doutb(w_n16489_38[1]),.doutc(w_n16489_38[2]),.din(w_n16489_12[1]));
	jspl3 jspl3_w_n16489_39(.douta(w_n16489_39[0]),.doutb(w_n16489_39[1]),.doutc(w_n16489_39[2]),.din(w_n16489_12[2]));
	jspl jspl_w_n16492_0(.douta(w_n16492_0[0]),.doutb(w_n16492_0[1]),.din(n16492));
	jspl3 jspl3_w_n16493_0(.douta(w_n16493_0[0]),.doutb(w_n16493_0[1]),.doutc(w_n16493_0[2]),.din(n16493));
	jspl3 jspl3_w_n16494_0(.douta(w_n16494_0[0]),.doutb(w_n16494_0[1]),.doutc(w_n16494_0[2]),.din(n16494));
	jspl3 jspl3_w_n16494_1(.douta(w_n16494_1[0]),.doutb(w_n16494_1[1]),.doutc(w_n16494_1[2]),.din(w_n16494_0[0]));
	jspl jspl_w_n16495_0(.douta(w_n16495_0[0]),.doutb(w_n16495_0[1]),.din(n16495));
	jspl3 jspl3_w_n16496_0(.douta(w_n16496_0[0]),.doutb(w_n16496_0[1]),.doutc(w_n16496_0[2]),.din(n16496));
	jspl jspl_w_n16497_0(.douta(w_n16497_0[0]),.doutb(w_n16497_0[1]),.din(n16497));
	jspl3 jspl3_w_n16500_0(.douta(w_n16500_0[0]),.doutb(w_n16500_0[1]),.doutc(w_n16500_0[2]),.din(n16500));
	jspl jspl_w_n16501_0(.douta(w_n16501_0[0]),.doutb(w_n16501_0[1]),.din(n16501));
	jspl3 jspl3_w_n16508_0(.douta(w_n16508_0[0]),.doutb(w_n16508_0[1]),.doutc(w_n16508_0[2]),.din(n16508));
	jspl jspl_w_n16509_0(.douta(w_n16509_0[0]),.doutb(w_n16509_0[1]),.din(n16509));
	jspl jspl_w_n16512_0(.douta(w_n16512_0[0]),.doutb(w_n16512_0[1]),.din(n16512));
	jspl3 jspl3_w_n16517_0(.douta(w_n16517_0[0]),.doutb(w_n16517_0[1]),.doutc(w_n16517_0[2]),.din(n16517));
	jspl3 jspl3_w_n16519_0(.douta(w_n16519_0[0]),.doutb(w_n16519_0[1]),.doutc(w_n16519_0[2]),.din(n16519));
	jspl jspl_w_n16520_0(.douta(w_n16520_0[0]),.doutb(w_n16520_0[1]),.din(n16520));
	jspl3 jspl3_w_n16524_0(.douta(w_n16524_0[0]),.doutb(w_n16524_0[1]),.doutc(w_n16524_0[2]),.din(n16524));
	jspl3 jspl3_w_n16527_0(.douta(w_n16527_0[0]),.doutb(w_n16527_0[1]),.doutc(w_n16527_0[2]),.din(n16527));
	jspl jspl_w_n16528_0(.douta(w_n16528_0[0]),.doutb(w_n16528_0[1]),.din(n16528));
	jspl3 jspl3_w_n16532_0(.douta(w_n16532_0[0]),.doutb(w_n16532_0[1]),.doutc(w_n16532_0[2]),.din(n16532));
	jspl3 jspl3_w_n16534_0(.douta(w_n16534_0[0]),.doutb(w_n16534_0[1]),.doutc(w_n16534_0[2]),.din(n16534));
	jspl jspl_w_n16535_0(.douta(w_n16535_0[0]),.doutb(w_n16535_0[1]),.din(n16535));
	jspl3 jspl3_w_n16539_0(.douta(w_n16539_0[0]),.doutb(w_n16539_0[1]),.doutc(w_n16539_0[2]),.din(n16539));
	jspl3 jspl3_w_n16541_0(.douta(w_n16541_0[0]),.doutb(w_n16541_0[1]),.doutc(w_n16541_0[2]),.din(n16541));
	jspl jspl_w_n16542_0(.douta(w_n16542_0[0]),.doutb(w_n16542_0[1]),.din(n16542));
	jspl3 jspl3_w_n16546_0(.douta(w_n16546_0[0]),.doutb(w_n16546_0[1]),.doutc(w_n16546_0[2]),.din(n16546));
	jspl3 jspl3_w_n16549_0(.douta(w_n16549_0[0]),.doutb(w_n16549_0[1]),.doutc(w_n16549_0[2]),.din(n16549));
	jspl jspl_w_n16550_0(.douta(w_n16550_0[0]),.doutb(w_n16550_0[1]),.din(n16550));
	jspl3 jspl3_w_n16554_0(.douta(w_n16554_0[0]),.doutb(w_n16554_0[1]),.doutc(w_n16554_0[2]),.din(n16554));
	jspl3 jspl3_w_n16557_0(.douta(w_n16557_0[0]),.doutb(w_n16557_0[1]),.doutc(w_n16557_0[2]),.din(n16557));
	jspl jspl_w_n16558_0(.douta(w_n16558_0[0]),.doutb(w_n16558_0[1]),.din(n16558));
	jspl3 jspl3_w_n16562_0(.douta(w_n16562_0[0]),.doutb(w_n16562_0[1]),.doutc(w_n16562_0[2]),.din(n16562));
	jspl3 jspl3_w_n16564_0(.douta(w_n16564_0[0]),.doutb(w_n16564_0[1]),.doutc(w_n16564_0[2]),.din(n16564));
	jspl jspl_w_n16565_0(.douta(w_n16565_0[0]),.doutb(w_n16565_0[1]),.din(n16565));
	jspl3 jspl3_w_n16569_0(.douta(w_n16569_0[0]),.doutb(w_n16569_0[1]),.doutc(w_n16569_0[2]),.din(n16569));
	jspl3 jspl3_w_n16572_0(.douta(w_n16572_0[0]),.doutb(w_n16572_0[1]),.doutc(w_n16572_0[2]),.din(n16572));
	jspl jspl_w_n16573_0(.douta(w_n16573_0[0]),.doutb(w_n16573_0[1]),.din(n16573));
	jspl3 jspl3_w_n16577_0(.douta(w_n16577_0[0]),.doutb(w_n16577_0[1]),.doutc(w_n16577_0[2]),.din(n16577));
	jspl3 jspl3_w_n16579_0(.douta(w_n16579_0[0]),.doutb(w_n16579_0[1]),.doutc(w_n16579_0[2]),.din(n16579));
	jspl jspl_w_n16580_0(.douta(w_n16580_0[0]),.doutb(w_n16580_0[1]),.din(n16580));
	jspl3 jspl3_w_n16584_0(.douta(w_n16584_0[0]),.doutb(w_n16584_0[1]),.doutc(w_n16584_0[2]),.din(n16584));
	jspl3 jspl3_w_n16587_0(.douta(w_n16587_0[0]),.doutb(w_n16587_0[1]),.doutc(w_n16587_0[2]),.din(n16587));
	jspl jspl_w_n16588_0(.douta(w_n16588_0[0]),.doutb(w_n16588_0[1]),.din(n16588));
	jspl3 jspl3_w_n16592_0(.douta(w_n16592_0[0]),.doutb(w_n16592_0[1]),.doutc(w_n16592_0[2]),.din(n16592));
	jspl3 jspl3_w_n16594_0(.douta(w_n16594_0[0]),.doutb(w_n16594_0[1]),.doutc(w_n16594_0[2]),.din(n16594));
	jspl jspl_w_n16595_0(.douta(w_n16595_0[0]),.doutb(w_n16595_0[1]),.din(n16595));
	jspl3 jspl3_w_n16599_0(.douta(w_n16599_0[0]),.doutb(w_n16599_0[1]),.doutc(w_n16599_0[2]),.din(n16599));
	jspl3 jspl3_w_n16601_0(.douta(w_n16601_0[0]),.doutb(w_n16601_0[1]),.doutc(w_n16601_0[2]),.din(n16601));
	jspl jspl_w_n16602_0(.douta(w_n16602_0[0]),.doutb(w_n16602_0[1]),.din(n16602));
	jspl3 jspl3_w_n16606_0(.douta(w_n16606_0[0]),.doutb(w_n16606_0[1]),.doutc(w_n16606_0[2]),.din(n16606));
	jspl3 jspl3_w_n16608_0(.douta(w_n16608_0[0]),.doutb(w_n16608_0[1]),.doutc(w_n16608_0[2]),.din(n16608));
	jspl jspl_w_n16609_0(.douta(w_n16609_0[0]),.doutb(w_n16609_0[1]),.din(n16609));
	jspl3 jspl3_w_n16613_0(.douta(w_n16613_0[0]),.doutb(w_n16613_0[1]),.doutc(w_n16613_0[2]),.din(n16613));
	jspl3 jspl3_w_n16616_0(.douta(w_n16616_0[0]),.doutb(w_n16616_0[1]),.doutc(w_n16616_0[2]),.din(n16616));
	jspl jspl_w_n16617_0(.douta(w_n16617_0[0]),.doutb(w_n16617_0[1]),.din(n16617));
	jspl3 jspl3_w_n16621_0(.douta(w_n16621_0[0]),.doutb(w_n16621_0[1]),.doutc(w_n16621_0[2]),.din(n16621));
	jspl3 jspl3_w_n16623_0(.douta(w_n16623_0[0]),.doutb(w_n16623_0[1]),.doutc(w_n16623_0[2]),.din(n16623));
	jspl jspl_w_n16624_0(.douta(w_n16624_0[0]),.doutb(w_n16624_0[1]),.din(n16624));
	jspl3 jspl3_w_n16628_0(.douta(w_n16628_0[0]),.doutb(w_n16628_0[1]),.doutc(w_n16628_0[2]),.din(n16628));
	jspl3 jspl3_w_n16631_0(.douta(w_n16631_0[0]),.doutb(w_n16631_0[1]),.doutc(w_n16631_0[2]),.din(n16631));
	jspl jspl_w_n16632_0(.douta(w_n16632_0[0]),.doutb(w_n16632_0[1]),.din(n16632));
	jspl3 jspl3_w_n16636_0(.douta(w_n16636_0[0]),.doutb(w_n16636_0[1]),.doutc(w_n16636_0[2]),.din(n16636));
	jspl3 jspl3_w_n16638_0(.douta(w_n16638_0[0]),.doutb(w_n16638_0[1]),.doutc(w_n16638_0[2]),.din(n16638));
	jspl jspl_w_n16639_0(.douta(w_n16639_0[0]),.doutb(w_n16639_0[1]),.din(n16639));
	jspl3 jspl3_w_n16643_0(.douta(w_n16643_0[0]),.doutb(w_n16643_0[1]),.doutc(w_n16643_0[2]),.din(n16643));
	jspl3 jspl3_w_n16646_0(.douta(w_n16646_0[0]),.doutb(w_n16646_0[1]),.doutc(w_n16646_0[2]),.din(n16646));
	jspl jspl_w_n16647_0(.douta(w_n16647_0[0]),.doutb(w_n16647_0[1]),.din(n16647));
	jspl3 jspl3_w_n16651_0(.douta(w_n16651_0[0]),.doutb(w_n16651_0[1]),.doutc(w_n16651_0[2]),.din(n16651));
	jspl3 jspl3_w_n16653_0(.douta(w_n16653_0[0]),.doutb(w_n16653_0[1]),.doutc(w_n16653_0[2]),.din(n16653));
	jspl jspl_w_n16654_0(.douta(w_n16654_0[0]),.doutb(w_n16654_0[1]),.din(n16654));
	jspl3 jspl3_w_n16658_0(.douta(w_n16658_0[0]),.doutb(w_n16658_0[1]),.doutc(w_n16658_0[2]),.din(n16658));
	jspl3 jspl3_w_n16661_0(.douta(w_n16661_0[0]),.doutb(w_n16661_0[1]),.doutc(w_n16661_0[2]),.din(n16661));
	jspl jspl_w_n16662_0(.douta(w_n16662_0[0]),.doutb(w_n16662_0[1]),.din(n16662));
	jspl3 jspl3_w_n16666_0(.douta(w_n16666_0[0]),.doutb(w_n16666_0[1]),.doutc(w_n16666_0[2]),.din(n16666));
	jspl3 jspl3_w_n16668_0(.douta(w_n16668_0[0]),.doutb(w_n16668_0[1]),.doutc(w_n16668_0[2]),.din(n16668));
	jspl jspl_w_n16669_0(.douta(w_n16669_0[0]),.doutb(w_n16669_0[1]),.din(n16669));
	jspl3 jspl3_w_n16673_0(.douta(w_n16673_0[0]),.doutb(w_n16673_0[1]),.doutc(w_n16673_0[2]),.din(n16673));
	jspl3 jspl3_w_n16675_0(.douta(w_n16675_0[0]),.doutb(w_n16675_0[1]),.doutc(w_n16675_0[2]),.din(n16675));
	jspl jspl_w_n16676_0(.douta(w_n16676_0[0]),.doutb(w_n16676_0[1]),.din(n16676));
	jspl3 jspl3_w_n16680_0(.douta(w_n16680_0[0]),.doutb(w_n16680_0[1]),.doutc(w_n16680_0[2]),.din(n16680));
	jspl3 jspl3_w_n16682_0(.douta(w_n16682_0[0]),.doutb(w_n16682_0[1]),.doutc(w_n16682_0[2]),.din(n16682));
	jspl jspl_w_n16683_0(.douta(w_n16683_0[0]),.doutb(w_n16683_0[1]),.din(n16683));
	jspl3 jspl3_w_n16687_0(.douta(w_n16687_0[0]),.doutb(w_n16687_0[1]),.doutc(w_n16687_0[2]),.din(n16687));
	jspl3 jspl3_w_n16690_0(.douta(w_n16690_0[0]),.doutb(w_n16690_0[1]),.doutc(w_n16690_0[2]),.din(n16690));
	jspl jspl_w_n16691_0(.douta(w_n16691_0[0]),.doutb(w_n16691_0[1]),.din(n16691));
	jspl3 jspl3_w_n16695_0(.douta(w_n16695_0[0]),.doutb(w_n16695_0[1]),.doutc(w_n16695_0[2]),.din(n16695));
	jspl3 jspl3_w_n16697_0(.douta(w_n16697_0[0]),.doutb(w_n16697_0[1]),.doutc(w_n16697_0[2]),.din(n16697));
	jspl jspl_w_n16698_0(.douta(w_n16698_0[0]),.doutb(w_n16698_0[1]),.din(n16698));
	jspl3 jspl3_w_n16702_0(.douta(w_n16702_0[0]),.doutb(w_n16702_0[1]),.doutc(w_n16702_0[2]),.din(n16702));
	jspl3 jspl3_w_n16705_0(.douta(w_n16705_0[0]),.doutb(w_n16705_0[1]),.doutc(w_n16705_0[2]),.din(n16705));
	jspl jspl_w_n16706_0(.douta(w_n16706_0[0]),.doutb(w_n16706_0[1]),.din(n16706));
	jspl3 jspl3_w_n16710_0(.douta(w_n16710_0[0]),.doutb(w_n16710_0[1]),.doutc(w_n16710_0[2]),.din(n16710));
	jspl3 jspl3_w_n16712_0(.douta(w_n16712_0[0]),.doutb(w_n16712_0[1]),.doutc(w_n16712_0[2]),.din(n16712));
	jspl jspl_w_n16713_0(.douta(w_n16713_0[0]),.doutb(w_n16713_0[1]),.din(n16713));
	jspl3 jspl3_w_n16717_0(.douta(w_n16717_0[0]),.doutb(w_n16717_0[1]),.doutc(w_n16717_0[2]),.din(n16717));
	jspl3 jspl3_w_n16719_0(.douta(w_n16719_0[0]),.doutb(w_n16719_0[1]),.doutc(w_n16719_0[2]),.din(n16719));
	jspl jspl_w_n16720_0(.douta(w_n16720_0[0]),.doutb(w_n16720_0[1]),.din(n16720));
	jspl3 jspl3_w_n16724_0(.douta(w_n16724_0[0]),.doutb(w_n16724_0[1]),.doutc(w_n16724_0[2]),.din(n16724));
	jspl3 jspl3_w_n16726_0(.douta(w_n16726_0[0]),.doutb(w_n16726_0[1]),.doutc(w_n16726_0[2]),.din(n16726));
	jspl jspl_w_n16727_0(.douta(w_n16727_0[0]),.doutb(w_n16727_0[1]),.din(n16727));
	jspl3 jspl3_w_n16731_0(.douta(w_n16731_0[0]),.doutb(w_n16731_0[1]),.doutc(w_n16731_0[2]),.din(n16731));
	jspl3 jspl3_w_n16734_0(.douta(w_n16734_0[0]),.doutb(w_n16734_0[1]),.doutc(w_n16734_0[2]),.din(n16734));
	jspl jspl_w_n16735_0(.douta(w_n16735_0[0]),.doutb(w_n16735_0[1]),.din(n16735));
	jspl3 jspl3_w_n16739_0(.douta(w_n16739_0[0]),.doutb(w_n16739_0[1]),.doutc(w_n16739_0[2]),.din(n16739));
	jspl3 jspl3_w_n16741_0(.douta(w_n16741_0[0]),.doutb(w_n16741_0[1]),.doutc(w_n16741_0[2]),.din(n16741));
	jspl jspl_w_n16742_0(.douta(w_n16742_0[0]),.doutb(w_n16742_0[1]),.din(n16742));
	jspl3 jspl3_w_n16746_0(.douta(w_n16746_0[0]),.doutb(w_n16746_0[1]),.doutc(w_n16746_0[2]),.din(n16746));
	jspl3 jspl3_w_n16749_0(.douta(w_n16749_0[0]),.doutb(w_n16749_0[1]),.doutc(w_n16749_0[2]),.din(n16749));
	jspl jspl_w_n16750_0(.douta(w_n16750_0[0]),.doutb(w_n16750_0[1]),.din(n16750));
	jspl3 jspl3_w_n16754_0(.douta(w_n16754_0[0]),.doutb(w_n16754_0[1]),.doutc(w_n16754_0[2]),.din(n16754));
	jspl3 jspl3_w_n16756_0(.douta(w_n16756_0[0]),.doutb(w_n16756_0[1]),.doutc(w_n16756_0[2]),.din(n16756));
	jspl jspl_w_n16757_0(.douta(w_n16757_0[0]),.doutb(w_n16757_0[1]),.din(n16757));
	jspl3 jspl3_w_n16761_0(.douta(w_n16761_0[0]),.doutb(w_n16761_0[1]),.doutc(w_n16761_0[2]),.din(n16761));
	jspl3 jspl3_w_n16763_0(.douta(w_n16763_0[0]),.doutb(w_n16763_0[1]),.doutc(w_n16763_0[2]),.din(n16763));
	jspl jspl_w_n16764_0(.douta(w_n16764_0[0]),.doutb(w_n16764_0[1]),.din(n16764));
	jspl3 jspl3_w_n16768_0(.douta(w_n16768_0[0]),.doutb(w_n16768_0[1]),.doutc(w_n16768_0[2]),.din(n16768));
	jspl3 jspl3_w_n16771_0(.douta(w_n16771_0[0]),.doutb(w_n16771_0[1]),.doutc(w_n16771_0[2]),.din(n16771));
	jspl jspl_w_n16772_0(.douta(w_n16772_0[0]),.doutb(w_n16772_0[1]),.din(n16772));
	jspl3 jspl3_w_n16775_0(.douta(w_n16775_0[0]),.doutb(w_n16775_0[1]),.doutc(w_n16775_0[2]),.din(n16775));
	jspl3 jspl3_w_n16779_0(.douta(w_n16779_0[0]),.doutb(w_n16779_0[1]),.doutc(w_n16779_0[2]),.din(n16779));
	jspl jspl_w_n16780_0(.douta(w_n16780_0[0]),.doutb(w_n16780_0[1]),.din(n16780));
	jspl3 jspl3_w_n16784_0(.douta(w_n16784_0[0]),.doutb(w_n16784_0[1]),.doutc(w_n16784_0[2]),.din(n16784));
	jspl3 jspl3_w_n16786_0(.douta(w_n16786_0[0]),.doutb(w_n16786_0[1]),.doutc(w_n16786_0[2]),.din(n16786));
	jspl jspl_w_n16787_0(.douta(w_n16787_0[0]),.doutb(w_n16787_0[1]),.din(n16787));
	jspl3 jspl3_w_n16791_0(.douta(w_n16791_0[0]),.doutb(w_n16791_0[1]),.doutc(w_n16791_0[2]),.din(n16791));
	jspl3 jspl3_w_n16794_0(.douta(w_n16794_0[0]),.doutb(w_n16794_0[1]),.doutc(w_n16794_0[2]),.din(n16794));
	jspl jspl_w_n16795_0(.douta(w_n16795_0[0]),.doutb(w_n16795_0[1]),.din(n16795));
	jspl3 jspl3_w_n16799_0(.douta(w_n16799_0[0]),.doutb(w_n16799_0[1]),.doutc(w_n16799_0[2]),.din(n16799));
	jspl3 jspl3_w_n16801_0(.douta(w_n16801_0[0]),.doutb(w_n16801_0[1]),.doutc(w_n16801_0[2]),.din(n16801));
	jspl jspl_w_n16802_0(.douta(w_n16802_0[0]),.doutb(w_n16802_0[1]),.din(n16802));
	jspl3 jspl3_w_n16806_0(.douta(w_n16806_0[0]),.doutb(w_n16806_0[1]),.doutc(w_n16806_0[2]),.din(n16806));
	jspl3 jspl3_w_n16809_0(.douta(w_n16809_0[0]),.doutb(w_n16809_0[1]),.doutc(w_n16809_0[2]),.din(n16809));
	jspl jspl_w_n16810_0(.douta(w_n16810_0[0]),.doutb(w_n16810_0[1]),.din(n16810));
	jspl3 jspl3_w_n16814_0(.douta(w_n16814_0[0]),.doutb(w_n16814_0[1]),.doutc(w_n16814_0[2]),.din(n16814));
	jspl3 jspl3_w_n16816_0(.douta(w_n16816_0[0]),.doutb(w_n16816_0[1]),.doutc(w_n16816_0[2]),.din(n16816));
	jspl jspl_w_n16817_0(.douta(w_n16817_0[0]),.doutb(w_n16817_0[1]),.din(n16817));
	jspl3 jspl3_w_n16821_0(.douta(w_n16821_0[0]),.doutb(w_n16821_0[1]),.doutc(w_n16821_0[2]),.din(n16821));
	jspl3 jspl3_w_n16823_0(.douta(w_n16823_0[0]),.doutb(w_n16823_0[1]),.doutc(w_n16823_0[2]),.din(n16823));
	jspl jspl_w_n16824_0(.douta(w_n16824_0[0]),.doutb(w_n16824_0[1]),.din(n16824));
	jspl3 jspl3_w_n16828_0(.douta(w_n16828_0[0]),.doutb(w_n16828_0[1]),.doutc(w_n16828_0[2]),.din(n16828));
	jspl3 jspl3_w_n16830_0(.douta(w_n16830_0[0]),.doutb(w_n16830_0[1]),.doutc(w_n16830_0[2]),.din(n16830));
	jspl jspl_w_n16831_0(.douta(w_n16831_0[0]),.doutb(w_n16831_0[1]),.din(n16831));
	jspl3 jspl3_w_n16835_0(.douta(w_n16835_0[0]),.doutb(w_n16835_0[1]),.doutc(w_n16835_0[2]),.din(n16835));
	jspl3 jspl3_w_n16838_0(.douta(w_n16838_0[0]),.doutb(w_n16838_0[1]),.doutc(w_n16838_0[2]),.din(n16838));
	jspl jspl_w_n16839_0(.douta(w_n16839_0[0]),.doutb(w_n16839_0[1]),.din(n16839));
	jspl3 jspl3_w_n16843_0(.douta(w_n16843_0[0]),.doutb(w_n16843_0[1]),.doutc(w_n16843_0[2]),.din(n16843));
	jspl3 jspl3_w_n16845_0(.douta(w_n16845_0[0]),.doutb(w_n16845_0[1]),.doutc(w_n16845_0[2]),.din(n16845));
	jspl jspl_w_n16846_0(.douta(w_n16846_0[0]),.doutb(w_n16846_0[1]),.din(n16846));
	jspl3 jspl3_w_n16850_0(.douta(w_n16850_0[0]),.doutb(w_n16850_0[1]),.doutc(w_n16850_0[2]),.din(n16850));
	jspl3 jspl3_w_n16853_0(.douta(w_n16853_0[0]),.doutb(w_n16853_0[1]),.doutc(w_n16853_0[2]),.din(n16853));
	jspl jspl_w_n16854_0(.douta(w_n16854_0[0]),.doutb(w_n16854_0[1]),.din(n16854));
	jspl3 jspl3_w_n16858_0(.douta(w_n16858_0[0]),.doutb(w_n16858_0[1]),.doutc(w_n16858_0[2]),.din(n16858));
	jspl3 jspl3_w_n16860_0(.douta(w_n16860_0[0]),.doutb(w_n16860_0[1]),.doutc(w_n16860_0[2]),.din(n16860));
	jspl jspl_w_n16861_0(.douta(w_n16861_0[0]),.doutb(w_n16861_0[1]),.din(n16861));
	jspl jspl_w_n16865_0(.douta(w_n16865_0[0]),.doutb(w_n16865_0[1]),.din(n16865));
	jspl jspl_w_n16866_0(.douta(w_n16866_0[0]),.doutb(w_n16866_0[1]),.din(n16866));
	jspl3 jspl3_w_n16868_0(.douta(w_n16868_0[0]),.doutb(w_n16868_0[1]),.doutc(w_n16868_0[2]),.din(n16868));
	jspl3 jspl3_w_n16869_0(.douta(w_n16869_0[0]),.doutb(w_n16869_0[1]),.doutc(w_n16869_0[2]),.din(n16869));
	jspl jspl_w_n16871_0(.douta(w_n16871_0[0]),.doutb(w_n16871_0[1]),.din(n16871));
	jspl jspl_w_n16872_0(.douta(w_n16872_0[0]),.doutb(w_n16872_0[1]),.din(n16872));
	jspl jspl_w_n16879_0(.douta(w_n16879_0[0]),.doutb(w_n16879_0[1]),.din(n16879));
	jspl jspl_w_n16880_0(.douta(w_n16880_0[0]),.doutb(w_n16880_0[1]),.din(n16880));
	jspl jspl_w_n16882_0(.douta(w_n16882_0[0]),.doutb(w_n16882_0[1]),.din(n16882));
	jspl3 jspl3_w_n16885_0(.douta(w_n16885_0[0]),.doutb(w_n16885_0[1]),.doutc(w_n16885_0[2]),.din(n16885));
	jspl jspl_w_n16885_1(.douta(w_n16885_1[0]),.doutb(w_n16885_1[1]),.din(w_n16885_0[0]));
	jspl jspl_w_n16886_0(.douta(w_n16886_0[0]),.doutb(w_n16886_0[1]),.din(n16886));
	jspl3 jspl3_w_n16887_0(.douta(w_n16887_0[0]),.doutb(w_n16887_0[1]),.doutc(w_n16887_0[2]),.din(n16887));
	jspl jspl_w_n16888_0(.douta(w_n16888_0[0]),.doutb(w_n16888_0[1]),.din(n16888));
	jspl3 jspl3_w_n16890_0(.douta(w_n16890_0[0]),.doutb(w_n16890_0[1]),.doutc(w_n16890_0[2]),.din(n16890));
	jspl jspl_w_n16891_0(.douta(w_n16891_0[0]),.doutb(w_n16891_0[1]),.din(n16891));
	jspl3 jspl3_w_n16896_0(.douta(w_n16896_0[0]),.doutb(w_n16896_0[1]),.doutc(w_n16896_0[2]),.din(n16896));
	jspl jspl_w_n16896_1(.douta(w_n16896_1[0]),.doutb(w_n16896_1[1]),.din(w_n16896_0[0]));
	jspl jspl_w_n16952_0(.douta(w_n16952_0[0]),.doutb(w_n16952_0[1]),.din(n16952));
	jspl jspl_w_n17127_0(.douta(w_n17127_0[0]),.doutb(w_n17127_0[1]),.din(n17127));
	jspl jspl_w_n17131_0(.douta(w_n17131_0[0]),.doutb(w_n17131_0[1]),.din(n17131));
	jspl jspl_w_n17132_0(.douta(w_n17132_0[0]),.doutb(w_n17132_0[1]),.din(n17132));
	jspl3 jspl3_w_n17134_0(.douta(w_n17134_0[0]),.doutb(w_n17134_0[1]),.doutc(w_n17134_0[2]),.din(n17134));
	jspl3 jspl3_w_n17134_1(.douta(w_n17134_1[0]),.doutb(w_n17134_1[1]),.doutc(w_n17134_1[2]),.din(w_n17134_0[0]));
	jspl3 jspl3_w_n17134_2(.douta(w_n17134_2[0]),.doutb(w_n17134_2[1]),.doutc(w_n17134_2[2]),.din(w_n17134_0[1]));
	jspl3 jspl3_w_n17134_3(.douta(w_n17134_3[0]),.doutb(w_n17134_3[1]),.doutc(w_n17134_3[2]),.din(w_n17134_0[2]));
	jspl3 jspl3_w_n17134_4(.douta(w_n17134_4[0]),.doutb(w_n17134_4[1]),.doutc(w_n17134_4[2]),.din(w_n17134_1[0]));
	jspl3 jspl3_w_n17134_5(.douta(w_n17134_5[0]),.doutb(w_n17134_5[1]),.doutc(w_n17134_5[2]),.din(w_n17134_1[1]));
	jspl3 jspl3_w_n17134_6(.douta(w_n17134_6[0]),.doutb(w_n17134_6[1]),.doutc(w_n17134_6[2]),.din(w_n17134_1[2]));
	jspl3 jspl3_w_n17134_7(.douta(w_n17134_7[0]),.doutb(w_n17134_7[1]),.doutc(w_n17134_7[2]),.din(w_n17134_2[0]));
	jspl3 jspl3_w_n17134_8(.douta(w_n17134_8[0]),.doutb(w_n17134_8[1]),.doutc(w_n17134_8[2]),.din(w_n17134_2[1]));
	jspl3 jspl3_w_n17134_9(.douta(w_n17134_9[0]),.doutb(w_n17134_9[1]),.doutc(w_n17134_9[2]),.din(w_n17134_2[2]));
	jspl3 jspl3_w_n17134_10(.douta(w_n17134_10[0]),.doutb(w_n17134_10[1]),.doutc(w_n17134_10[2]),.din(w_n17134_3[0]));
	jspl3 jspl3_w_n17134_11(.douta(w_n17134_11[0]),.doutb(w_n17134_11[1]),.doutc(w_n17134_11[2]),.din(w_n17134_3[1]));
	jspl3 jspl3_w_n17134_12(.douta(w_n17134_12[0]),.doutb(w_n17134_12[1]),.doutc(w_n17134_12[2]),.din(w_n17134_3[2]));
	jspl3 jspl3_w_n17134_13(.douta(w_n17134_13[0]),.doutb(w_n17134_13[1]),.doutc(w_n17134_13[2]),.din(w_n17134_4[0]));
	jspl3 jspl3_w_n17134_14(.douta(w_n17134_14[0]),.doutb(w_n17134_14[1]),.doutc(w_n17134_14[2]),.din(w_n17134_4[1]));
	jspl jspl_w_n17134_15(.douta(w_n17134_15[0]),.doutb(w_n17134_15[1]),.din(w_n17134_4[2]));
	jspl3 jspl3_w_n17138_0(.douta(w_n17138_0[0]),.doutb(w_n17138_0[1]),.doutc(w_n17138_0[2]),.din(n17138));
	jspl jspl_w_n17139_0(.douta(w_n17139_0[0]),.doutb(w_n17139_0[1]),.din(n17139));
	jspl jspl_w_n17141_0(.douta(w_n17141_0[0]),.doutb(w_n17141_0[1]),.din(n17141));
	jspl jspl_w_n17146_0(.douta(w_n17146_0[0]),.doutb(w_n17146_0[1]),.din(n17146));
	jspl jspl_w_n17147_0(.douta(w_n17147_0[0]),.doutb(w_n17147_0[1]),.din(n17147));
	jspl3 jspl3_w_n17149_0(.douta(w_n17149_0[0]),.doutb(w_n17149_0[1]),.doutc(w_n17149_0[2]),.din(n17149));
	jspl jspl_w_n17150_0(.douta(w_n17150_0[0]),.doutb(w_n17150_0[1]),.din(n17150));
	jspl jspl_w_n17154_0(.douta(w_n17154_0[0]),.doutb(w_n17154_0[1]),.din(n17154));
	jspl3 jspl3_w_n17156_0(.douta(w_n17156_0[0]),.doutb(w_n17156_0[1]),.doutc(w_n17156_0[2]),.din(n17156));
	jspl jspl_w_n17157_0(.douta(w_n17157_0[0]),.doutb(w_n17157_0[1]),.din(n17157));
	jspl jspl_w_n17161_0(.douta(w_n17161_0[0]),.doutb(w_n17161_0[1]),.din(n17161));
	jspl jspl_w_n17162_0(.douta(w_n17162_0[0]),.doutb(w_n17162_0[1]),.din(n17162));
	jspl3 jspl3_w_n17164_0(.douta(w_n17164_0[0]),.doutb(w_n17164_0[1]),.doutc(w_n17164_0[2]),.din(n17164));
	jspl jspl_w_n17165_0(.douta(w_n17165_0[0]),.doutb(w_n17165_0[1]),.din(n17165));
	jspl jspl_w_n17169_0(.douta(w_n17169_0[0]),.doutb(w_n17169_0[1]),.din(n17169));
	jspl3 jspl3_w_n17171_0(.douta(w_n17171_0[0]),.doutb(w_n17171_0[1]),.doutc(w_n17171_0[2]),.din(n17171));
	jspl jspl_w_n17172_0(.douta(w_n17172_0[0]),.doutb(w_n17172_0[1]),.din(n17172));
	jspl jspl_w_n17176_0(.douta(w_n17176_0[0]),.doutb(w_n17176_0[1]),.din(n17176));
	jspl jspl_w_n17177_0(.douta(w_n17177_0[0]),.doutb(w_n17177_0[1]),.din(n17177));
	jspl3 jspl3_w_n17179_0(.douta(w_n17179_0[0]),.doutb(w_n17179_0[1]),.doutc(w_n17179_0[2]),.din(n17179));
	jspl jspl_w_n17180_0(.douta(w_n17180_0[0]),.doutb(w_n17180_0[1]),.din(n17180));
	jspl jspl_w_n17184_0(.douta(w_n17184_0[0]),.doutb(w_n17184_0[1]),.din(n17184));
	jspl jspl_w_n17185_0(.douta(w_n17185_0[0]),.doutb(w_n17185_0[1]),.din(n17185));
	jspl3 jspl3_w_n17187_0(.douta(w_n17187_0[0]),.doutb(w_n17187_0[1]),.doutc(w_n17187_0[2]),.din(n17187));
	jspl jspl_w_n17188_0(.douta(w_n17188_0[0]),.doutb(w_n17188_0[1]),.din(n17188));
	jspl jspl_w_n17192_0(.douta(w_n17192_0[0]),.doutb(w_n17192_0[1]),.din(n17192));
	jspl3 jspl3_w_n17194_0(.douta(w_n17194_0[0]),.doutb(w_n17194_0[1]),.doutc(w_n17194_0[2]),.din(n17194));
	jspl jspl_w_n17195_0(.douta(w_n17195_0[0]),.doutb(w_n17195_0[1]),.din(n17195));
	jspl jspl_w_n17199_0(.douta(w_n17199_0[0]),.doutb(w_n17199_0[1]),.din(n17199));
	jspl3 jspl3_w_n17201_0(.douta(w_n17201_0[0]),.doutb(w_n17201_0[1]),.doutc(w_n17201_0[2]),.din(n17201));
	jspl jspl_w_n17202_0(.douta(w_n17202_0[0]),.doutb(w_n17202_0[1]),.din(n17202));
	jspl jspl_w_n17206_0(.douta(w_n17206_0[0]),.doutb(w_n17206_0[1]),.din(n17206));
	jspl jspl_w_n17207_0(.douta(w_n17207_0[0]),.doutb(w_n17207_0[1]),.din(n17207));
	jspl3 jspl3_w_n17209_0(.douta(w_n17209_0[0]),.doutb(w_n17209_0[1]),.doutc(w_n17209_0[2]),.din(n17209));
	jspl jspl_w_n17210_0(.douta(w_n17210_0[0]),.doutb(w_n17210_0[1]),.din(n17210));
	jspl jspl_w_n17214_0(.douta(w_n17214_0[0]),.doutb(w_n17214_0[1]),.din(n17214));
	jspl3 jspl3_w_n17216_0(.douta(w_n17216_0[0]),.doutb(w_n17216_0[1]),.doutc(w_n17216_0[2]),.din(n17216));
	jspl jspl_w_n17217_0(.douta(w_n17217_0[0]),.doutb(w_n17217_0[1]),.din(n17217));
	jspl jspl_w_n17221_0(.douta(w_n17221_0[0]),.doutb(w_n17221_0[1]),.din(n17221));
	jspl jspl_w_n17222_0(.douta(w_n17222_0[0]),.doutb(w_n17222_0[1]),.din(n17222));
	jspl3 jspl3_w_n17224_0(.douta(w_n17224_0[0]),.doutb(w_n17224_0[1]),.doutc(w_n17224_0[2]),.din(n17224));
	jspl jspl_w_n17225_0(.douta(w_n17225_0[0]),.doutb(w_n17225_0[1]),.din(n17225));
	jspl jspl_w_n17229_0(.douta(w_n17229_0[0]),.doutb(w_n17229_0[1]),.din(n17229));
	jspl3 jspl3_w_n17231_0(.douta(w_n17231_0[0]),.doutb(w_n17231_0[1]),.doutc(w_n17231_0[2]),.din(n17231));
	jspl jspl_w_n17232_0(.douta(w_n17232_0[0]),.doutb(w_n17232_0[1]),.din(n17232));
	jspl jspl_w_n17236_0(.douta(w_n17236_0[0]),.doutb(w_n17236_0[1]),.din(n17236));
	jspl jspl_w_n17237_0(.douta(w_n17237_0[0]),.doutb(w_n17237_0[1]),.din(n17237));
	jspl3 jspl3_w_n17239_0(.douta(w_n17239_0[0]),.doutb(w_n17239_0[1]),.doutc(w_n17239_0[2]),.din(n17239));
	jspl jspl_w_n17240_0(.douta(w_n17240_0[0]),.doutb(w_n17240_0[1]),.din(n17240));
	jspl jspl_w_n17244_0(.douta(w_n17244_0[0]),.doutb(w_n17244_0[1]),.din(n17244));
	jspl jspl_w_n17245_0(.douta(w_n17245_0[0]),.doutb(w_n17245_0[1]),.din(n17245));
	jspl3 jspl3_w_n17247_0(.douta(w_n17247_0[0]),.doutb(w_n17247_0[1]),.doutc(w_n17247_0[2]),.din(n17247));
	jspl jspl_w_n17248_0(.douta(w_n17248_0[0]),.doutb(w_n17248_0[1]),.din(n17248));
	jspl jspl_w_n17252_0(.douta(w_n17252_0[0]),.doutb(w_n17252_0[1]),.din(n17252));
	jspl jspl_w_n17253_0(.douta(w_n17253_0[0]),.doutb(w_n17253_0[1]),.din(n17253));
	jspl3 jspl3_w_n17255_0(.douta(w_n17255_0[0]),.doutb(w_n17255_0[1]),.doutc(w_n17255_0[2]),.din(n17255));
	jspl jspl_w_n17256_0(.douta(w_n17256_0[0]),.doutb(w_n17256_0[1]),.din(n17256));
	jspl jspl_w_n17260_0(.douta(w_n17260_0[0]),.doutb(w_n17260_0[1]),.din(n17260));
	jspl3 jspl3_w_n17262_0(.douta(w_n17262_0[0]),.doutb(w_n17262_0[1]),.doutc(w_n17262_0[2]),.din(n17262));
	jspl jspl_w_n17263_0(.douta(w_n17263_0[0]),.doutb(w_n17263_0[1]),.din(n17263));
	jspl jspl_w_n17267_0(.douta(w_n17267_0[0]),.doutb(w_n17267_0[1]),.din(n17267));
	jspl jspl_w_n17268_0(.douta(w_n17268_0[0]),.doutb(w_n17268_0[1]),.din(n17268));
	jspl3 jspl3_w_n17270_0(.douta(w_n17270_0[0]),.doutb(w_n17270_0[1]),.doutc(w_n17270_0[2]),.din(n17270));
	jspl jspl_w_n17271_0(.douta(w_n17271_0[0]),.doutb(w_n17271_0[1]),.din(n17271));
	jspl jspl_w_n17275_0(.douta(w_n17275_0[0]),.doutb(w_n17275_0[1]),.din(n17275));
	jspl3 jspl3_w_n17277_0(.douta(w_n17277_0[0]),.doutb(w_n17277_0[1]),.doutc(w_n17277_0[2]),.din(n17277));
	jspl jspl_w_n17278_0(.douta(w_n17278_0[0]),.doutb(w_n17278_0[1]),.din(n17278));
	jspl jspl_w_n17282_0(.douta(w_n17282_0[0]),.doutb(w_n17282_0[1]),.din(n17282));
	jspl jspl_w_n17283_0(.douta(w_n17283_0[0]),.doutb(w_n17283_0[1]),.din(n17283));
	jspl3 jspl3_w_n17285_0(.douta(w_n17285_0[0]),.doutb(w_n17285_0[1]),.doutc(w_n17285_0[2]),.din(n17285));
	jspl jspl_w_n17286_0(.douta(w_n17286_0[0]),.doutb(w_n17286_0[1]),.din(n17286));
	jspl jspl_w_n17290_0(.douta(w_n17290_0[0]),.doutb(w_n17290_0[1]),.din(n17290));
	jspl3 jspl3_w_n17292_0(.douta(w_n17292_0[0]),.doutb(w_n17292_0[1]),.doutc(w_n17292_0[2]),.din(n17292));
	jspl jspl_w_n17293_0(.douta(w_n17293_0[0]),.doutb(w_n17293_0[1]),.din(n17293));
	jspl jspl_w_n17297_0(.douta(w_n17297_0[0]),.doutb(w_n17297_0[1]),.din(n17297));
	jspl jspl_w_n17298_0(.douta(w_n17298_0[0]),.doutb(w_n17298_0[1]),.din(n17298));
	jspl3 jspl3_w_n17300_0(.douta(w_n17300_0[0]),.doutb(w_n17300_0[1]),.doutc(w_n17300_0[2]),.din(n17300));
	jspl jspl_w_n17301_0(.douta(w_n17301_0[0]),.doutb(w_n17301_0[1]),.din(n17301));
	jspl jspl_w_n17305_0(.douta(w_n17305_0[0]),.doutb(w_n17305_0[1]),.din(n17305));
	jspl3 jspl3_w_n17307_0(.douta(w_n17307_0[0]),.doutb(w_n17307_0[1]),.doutc(w_n17307_0[2]),.din(n17307));
	jspl jspl_w_n17308_0(.douta(w_n17308_0[0]),.doutb(w_n17308_0[1]),.din(n17308));
	jspl jspl_w_n17312_0(.douta(w_n17312_0[0]),.doutb(w_n17312_0[1]),.din(n17312));
	jspl jspl_w_n17313_0(.douta(w_n17313_0[0]),.doutb(w_n17313_0[1]),.din(n17313));
	jspl3 jspl3_w_n17315_0(.douta(w_n17315_0[0]),.doutb(w_n17315_0[1]),.doutc(w_n17315_0[2]),.din(n17315));
	jspl jspl_w_n17316_0(.douta(w_n17316_0[0]),.doutb(w_n17316_0[1]),.din(n17316));
	jspl jspl_w_n17320_0(.douta(w_n17320_0[0]),.doutb(w_n17320_0[1]),.din(n17320));
	jspl jspl_w_n17321_0(.douta(w_n17321_0[0]),.doutb(w_n17321_0[1]),.din(n17321));
	jspl3 jspl3_w_n17323_0(.douta(w_n17323_0[0]),.doutb(w_n17323_0[1]),.doutc(w_n17323_0[2]),.din(n17323));
	jspl jspl_w_n17324_0(.douta(w_n17324_0[0]),.doutb(w_n17324_0[1]),.din(n17324));
	jspl jspl_w_n17328_0(.douta(w_n17328_0[0]),.doutb(w_n17328_0[1]),.din(n17328));
	jspl jspl_w_n17329_0(.douta(w_n17329_0[0]),.doutb(w_n17329_0[1]),.din(n17329));
	jspl3 jspl3_w_n17331_0(.douta(w_n17331_0[0]),.doutb(w_n17331_0[1]),.doutc(w_n17331_0[2]),.din(n17331));
	jspl jspl_w_n17332_0(.douta(w_n17332_0[0]),.doutb(w_n17332_0[1]),.din(n17332));
	jspl jspl_w_n17336_0(.douta(w_n17336_0[0]),.doutb(w_n17336_0[1]),.din(n17336));
	jspl3 jspl3_w_n17338_0(.douta(w_n17338_0[0]),.doutb(w_n17338_0[1]),.doutc(w_n17338_0[2]),.din(n17338));
	jspl jspl_w_n17339_0(.douta(w_n17339_0[0]),.doutb(w_n17339_0[1]),.din(n17339));
	jspl jspl_w_n17343_0(.douta(w_n17343_0[0]),.doutb(w_n17343_0[1]),.din(n17343));
	jspl jspl_w_n17344_0(.douta(w_n17344_0[0]),.doutb(w_n17344_0[1]),.din(n17344));
	jspl3 jspl3_w_n17346_0(.douta(w_n17346_0[0]),.doutb(w_n17346_0[1]),.doutc(w_n17346_0[2]),.din(n17346));
	jspl jspl_w_n17347_0(.douta(w_n17347_0[0]),.doutb(w_n17347_0[1]),.din(n17347));
	jspl jspl_w_n17351_0(.douta(w_n17351_0[0]),.doutb(w_n17351_0[1]),.din(n17351));
	jspl3 jspl3_w_n17353_0(.douta(w_n17353_0[0]),.doutb(w_n17353_0[1]),.doutc(w_n17353_0[2]),.din(n17353));
	jspl jspl_w_n17354_0(.douta(w_n17354_0[0]),.doutb(w_n17354_0[1]),.din(n17354));
	jspl jspl_w_n17358_0(.douta(w_n17358_0[0]),.doutb(w_n17358_0[1]),.din(n17358));
	jspl jspl_w_n17359_0(.douta(w_n17359_0[0]),.doutb(w_n17359_0[1]),.din(n17359));
	jspl3 jspl3_w_n17361_0(.douta(w_n17361_0[0]),.doutb(w_n17361_0[1]),.doutc(w_n17361_0[2]),.din(n17361));
	jspl jspl_w_n17362_0(.douta(w_n17362_0[0]),.doutb(w_n17362_0[1]),.din(n17362));
	jspl jspl_w_n17366_0(.douta(w_n17366_0[0]),.doutb(w_n17366_0[1]),.din(n17366));
	jspl jspl_w_n17367_0(.douta(w_n17367_0[0]),.doutb(w_n17367_0[1]),.din(n17367));
	jspl3 jspl3_w_n17369_0(.douta(w_n17369_0[0]),.doutb(w_n17369_0[1]),.doutc(w_n17369_0[2]),.din(n17369));
	jspl jspl_w_n17370_0(.douta(w_n17370_0[0]),.doutb(w_n17370_0[1]),.din(n17370));
	jspl jspl_w_n17374_0(.douta(w_n17374_0[0]),.doutb(w_n17374_0[1]),.din(n17374));
	jspl jspl_w_n17375_0(.douta(w_n17375_0[0]),.doutb(w_n17375_0[1]),.din(n17375));
	jspl3 jspl3_w_n17377_0(.douta(w_n17377_0[0]),.doutb(w_n17377_0[1]),.doutc(w_n17377_0[2]),.din(n17377));
	jspl jspl_w_n17378_0(.douta(w_n17378_0[0]),.doutb(w_n17378_0[1]),.din(n17378));
	jspl jspl_w_n17382_0(.douta(w_n17382_0[0]),.doutb(w_n17382_0[1]),.din(n17382));
	jspl3 jspl3_w_n17384_0(.douta(w_n17384_0[0]),.doutb(w_n17384_0[1]),.doutc(w_n17384_0[2]),.din(n17384));
	jspl jspl_w_n17385_0(.douta(w_n17385_0[0]),.doutb(w_n17385_0[1]),.din(n17385));
	jspl jspl_w_n17389_0(.douta(w_n17389_0[0]),.doutb(w_n17389_0[1]),.din(n17389));
	jspl jspl_w_n17390_0(.douta(w_n17390_0[0]),.doutb(w_n17390_0[1]),.din(n17390));
	jspl3 jspl3_w_n17392_0(.douta(w_n17392_0[0]),.doutb(w_n17392_0[1]),.doutc(w_n17392_0[2]),.din(n17392));
	jspl jspl_w_n17393_0(.douta(w_n17393_0[0]),.doutb(w_n17393_0[1]),.din(n17393));
	jspl jspl_w_n17397_0(.douta(w_n17397_0[0]),.doutb(w_n17397_0[1]),.din(n17397));
	jspl3 jspl3_w_n17399_0(.douta(w_n17399_0[0]),.doutb(w_n17399_0[1]),.doutc(w_n17399_0[2]),.din(n17399));
	jspl jspl_w_n17400_0(.douta(w_n17400_0[0]),.doutb(w_n17400_0[1]),.din(n17400));
	jspl jspl_w_n17404_0(.douta(w_n17404_0[0]),.doutb(w_n17404_0[1]),.din(n17404));
	jspl jspl_w_n17405_0(.douta(w_n17405_0[0]),.doutb(w_n17405_0[1]),.din(n17405));
	jspl3 jspl3_w_n17407_0(.douta(w_n17407_0[0]),.doutb(w_n17407_0[1]),.doutc(w_n17407_0[2]),.din(n17407));
	jspl jspl_w_n17408_0(.douta(w_n17408_0[0]),.doutb(w_n17408_0[1]),.din(n17408));
	jspl jspl_w_n17412_0(.douta(w_n17412_0[0]),.doutb(w_n17412_0[1]),.din(n17412));
	jspl jspl_w_n17413_0(.douta(w_n17413_0[0]),.doutb(w_n17413_0[1]),.din(n17413));
	jspl3 jspl3_w_n17415_0(.douta(w_n17415_0[0]),.doutb(w_n17415_0[1]),.doutc(w_n17415_0[2]),.din(n17415));
	jspl jspl_w_n17416_0(.douta(w_n17416_0[0]),.doutb(w_n17416_0[1]),.din(n17416));
	jspl jspl_w_n17420_0(.douta(w_n17420_0[0]),.doutb(w_n17420_0[1]),.din(n17420));
	jspl3 jspl3_w_n17422_0(.douta(w_n17422_0[0]),.doutb(w_n17422_0[1]),.doutc(w_n17422_0[2]),.din(n17422));
	jspl jspl_w_n17423_0(.douta(w_n17423_0[0]),.doutb(w_n17423_0[1]),.din(n17423));
	jspl jspl_w_n17426_0(.douta(w_n17426_0[0]),.doutb(w_n17426_0[1]),.din(n17426));
	jspl3 jspl3_w_n17429_0(.douta(w_n17429_0[0]),.doutb(w_n17429_0[1]),.doutc(w_n17429_0[2]),.din(n17429));
	jspl jspl_w_n17430_0(.douta(w_n17430_0[0]),.doutb(w_n17430_0[1]),.din(n17430));
	jspl jspl_w_n17434_0(.douta(w_n17434_0[0]),.doutb(w_n17434_0[1]),.din(n17434));
	jspl jspl_w_n17435_0(.douta(w_n17435_0[0]),.doutb(w_n17435_0[1]),.din(n17435));
	jspl3 jspl3_w_n17437_0(.douta(w_n17437_0[0]),.doutb(w_n17437_0[1]),.doutc(w_n17437_0[2]),.din(n17437));
	jspl jspl_w_n17438_0(.douta(w_n17438_0[0]),.doutb(w_n17438_0[1]),.din(n17438));
	jspl jspl_w_n17442_0(.douta(w_n17442_0[0]),.doutb(w_n17442_0[1]),.din(n17442));
	jspl3 jspl3_w_n17444_0(.douta(w_n17444_0[0]),.doutb(w_n17444_0[1]),.doutc(w_n17444_0[2]),.din(n17444));
	jspl jspl_w_n17445_0(.douta(w_n17445_0[0]),.doutb(w_n17445_0[1]),.din(n17445));
	jspl jspl_w_n17449_0(.douta(w_n17449_0[0]),.doutb(w_n17449_0[1]),.din(n17449));
	jspl jspl_w_n17450_0(.douta(w_n17450_0[0]),.doutb(w_n17450_0[1]),.din(n17450));
	jspl3 jspl3_w_n17452_0(.douta(w_n17452_0[0]),.doutb(w_n17452_0[1]),.doutc(w_n17452_0[2]),.din(n17452));
	jspl jspl_w_n17453_0(.douta(w_n17453_0[0]),.doutb(w_n17453_0[1]),.din(n17453));
	jspl jspl_w_n17457_0(.douta(w_n17457_0[0]),.doutb(w_n17457_0[1]),.din(n17457));
	jspl3 jspl3_w_n17459_0(.douta(w_n17459_0[0]),.doutb(w_n17459_0[1]),.doutc(w_n17459_0[2]),.din(n17459));
	jspl jspl_w_n17460_0(.douta(w_n17460_0[0]),.doutb(w_n17460_0[1]),.din(n17460));
	jspl jspl_w_n17464_0(.douta(w_n17464_0[0]),.doutb(w_n17464_0[1]),.din(n17464));
	jspl jspl_w_n17465_0(.douta(w_n17465_0[0]),.doutb(w_n17465_0[1]),.din(n17465));
	jspl3 jspl3_w_n17467_0(.douta(w_n17467_0[0]),.doutb(w_n17467_0[1]),.doutc(w_n17467_0[2]),.din(n17467));
	jspl jspl_w_n17468_0(.douta(w_n17468_0[0]),.doutb(w_n17468_0[1]),.din(n17468));
	jspl jspl_w_n17472_0(.douta(w_n17472_0[0]),.doutb(w_n17472_0[1]),.din(n17472));
	jspl jspl_w_n17473_0(.douta(w_n17473_0[0]),.doutb(w_n17473_0[1]),.din(n17473));
	jspl3 jspl3_w_n17475_0(.douta(w_n17475_0[0]),.doutb(w_n17475_0[1]),.doutc(w_n17475_0[2]),.din(n17475));
	jspl jspl_w_n17476_0(.douta(w_n17476_0[0]),.doutb(w_n17476_0[1]),.din(n17476));
	jspl jspl_w_n17480_0(.douta(w_n17480_0[0]),.doutb(w_n17480_0[1]),.din(n17480));
	jspl jspl_w_n17481_0(.douta(w_n17481_0[0]),.doutb(w_n17481_0[1]),.din(n17481));
	jspl3 jspl3_w_n17483_0(.douta(w_n17483_0[0]),.doutb(w_n17483_0[1]),.doutc(w_n17483_0[2]),.din(n17483));
	jspl jspl_w_n17484_0(.douta(w_n17484_0[0]),.doutb(w_n17484_0[1]),.din(n17484));
	jspl jspl_w_n17488_0(.douta(w_n17488_0[0]),.doutb(w_n17488_0[1]),.din(n17488));
	jspl3 jspl3_w_n17490_0(.douta(w_n17490_0[0]),.doutb(w_n17490_0[1]),.doutc(w_n17490_0[2]),.din(n17490));
	jspl jspl_w_n17491_0(.douta(w_n17491_0[0]),.doutb(w_n17491_0[1]),.din(n17491));
	jspl jspl_w_n17495_0(.douta(w_n17495_0[0]),.doutb(w_n17495_0[1]),.din(n17495));
	jspl jspl_w_n17496_0(.douta(w_n17496_0[0]),.doutb(w_n17496_0[1]),.din(n17496));
	jspl3 jspl3_w_n17498_0(.douta(w_n17498_0[0]),.doutb(w_n17498_0[1]),.doutc(w_n17498_0[2]),.din(n17498));
	jspl jspl_w_n17499_0(.douta(w_n17499_0[0]),.doutb(w_n17499_0[1]),.din(n17499));
	jspl jspl_w_n17503_0(.douta(w_n17503_0[0]),.doutb(w_n17503_0[1]),.din(n17503));
	jspl3 jspl3_w_n17505_0(.douta(w_n17505_0[0]),.doutb(w_n17505_0[1]),.doutc(w_n17505_0[2]),.din(n17505));
	jspl jspl_w_n17506_0(.douta(w_n17506_0[0]),.doutb(w_n17506_0[1]),.din(n17506));
	jspl3 jspl3_w_n17510_0(.douta(w_n17510_0[0]),.doutb(w_n17510_0[1]),.doutc(w_n17510_0[2]),.din(n17510));
	jspl jspl_w_n17513_0(.douta(w_n17513_0[0]),.doutb(w_n17513_0[1]),.din(n17513));
	jspl3 jspl3_w_n17516_0(.douta(w_n17516_0[0]),.doutb(w_n17516_0[1]),.doutc(w_n17516_0[2]),.din(n17516));
	jspl jspl_w_n17517_0(.douta(w_n17517_0[0]),.doutb(w_n17517_0[1]),.din(n17517));
	jspl3 jspl3_w_n17518_0(.douta(w_n17518_0[0]),.doutb(w_n17518_0[1]),.doutc(w_n17518_0[2]),.din(n17518));
	jspl jspl_w_n17518_1(.douta(w_n17518_1[0]),.doutb(w_n17518_1[1]),.din(w_n17518_0[0]));
	jspl3 jspl3_w_n17519_0(.douta(w_n17519_0[0]),.doutb(w_n17519_0[1]),.doutc(w_n17519_0[2]),.din(n17519));
	jspl jspl_w_n17523_0(.douta(w_n17523_0[0]),.doutb(w_n17523_0[1]),.din(n17523));
	jspl jspl_w_n17524_0(.douta(w_n17524_0[0]),.doutb(w_n17524_0[1]),.din(n17524));
	jspl jspl_w_n17525_0(.douta(w_n17525_0[0]),.doutb(w_n17525_0[1]),.din(n17525));
	jspl jspl_w_n17538_0(.douta(w_n17538_0[0]),.doutb(w_n17538_0[1]),.din(n17538));
	jspl jspl_w_n17583_0(.douta(w_n17583_0[0]),.doutb(w_n17583_0[1]),.din(n17583));
	jspl jspl_w_n17590_0(.douta(w_n17590_0[0]),.doutb(w_n17590_0[1]),.din(n17590));
	jspl jspl_w_n17597_0(.douta(w_n17597_0[0]),.doutb(w_n17597_0[1]),.din(n17597));
	jspl jspl_w_n17607_0(.douta(w_n17607_0[0]),.doutb(w_n17607_0[1]),.din(n17607));
	jspl jspl_w_n17611_0(.douta(w_n17611_0[0]),.doutb(w_n17611_0[1]),.din(n17611));
	jspl jspl_w_n17618_0(.douta(w_n17618_0[0]),.doutb(w_n17618_0[1]),.din(n17618));
	jspl jspl_w_n17625_0(.douta(w_n17625_0[0]),.doutb(w_n17625_0[1]),.din(n17625));
	jspl jspl_w_n17638_0(.douta(w_n17638_0[0]),.doutb(w_n17638_0[1]),.din(n17638));
	jspl jspl_w_n17645_0(.douta(w_n17645_0[0]),.doutb(w_n17645_0[1]),.din(n17645));
	jspl jspl_w_n17652_0(.douta(w_n17652_0[0]),.doutb(w_n17652_0[1]),.din(n17652));
	jspl jspl_w_n17659_0(.douta(w_n17659_0[0]),.doutb(w_n17659_0[1]),.din(n17659));
	jspl jspl_w_n17672_0(.douta(w_n17672_0[0]),.doutb(w_n17672_0[1]),.din(n17672));
	jspl jspl_w_n17679_0(.douta(w_n17679_0[0]),.doutb(w_n17679_0[1]),.din(n17679));
	jspl jspl_w_n17692_0(.douta(w_n17692_0[0]),.doutb(w_n17692_0[1]),.din(n17692));
	jspl jspl_w_n17699_0(.douta(w_n17699_0[0]),.doutb(w_n17699_0[1]),.din(n17699));
	jspl jspl_w_n17709_0(.douta(w_n17709_0[0]),.doutb(w_n17709_0[1]),.din(n17709));
	jspl jspl_w_n17719_0(.douta(w_n17719_0[0]),.doutb(w_n17719_0[1]),.din(n17719));
	jspl jspl_w_n17726_0(.douta(w_n17726_0[0]),.doutb(w_n17726_0[1]),.din(n17726));
	jspl jspl_w_n17739_0(.douta(w_n17739_0[0]),.doutb(w_n17739_0[1]),.din(n17739));
	jspl jspl_w_n17746_0(.douta(w_n17746_0[0]),.doutb(w_n17746_0[1]),.din(n17746));
	jspl jspl_w_n17751_0(.douta(w_n17751_0[0]),.doutb(w_n17751_0[1]),.din(n17751));
	jspl jspl_w_n17752_0(.douta(w_n17752_0[0]),.doutb(w_n17752_0[1]),.din(n17752));
	jspl jspl_w_n17755_0(.douta(w_n17755_0[0]),.doutb(w_n17755_0[1]),.din(n17755));
	jspl jspl_w_n17756_0(.douta(w_n17756_0[0]),.doutb(w_n17756_0[1]),.din(n17756));
	jspl jspl_w_n17758_0(.douta(w_n17758_0[0]),.doutb(w_n17758_0[1]),.din(n17758));
	jspl jspl_w_n17762_0(.douta(w_n17762_0[0]),.doutb(w_n17762_0[1]),.din(n17762));
	jspl jspl_w_n17768_0(.douta(w_n17768_0[0]),.doutb(w_n17768_0[1]),.din(n17768));
	jspl3 jspl3_w_n17769_0(.douta(w_n17769_0[0]),.doutb(w_n17769_0[1]),.doutc(w_n17769_0[2]),.din(n17769));
	jspl3 jspl3_w_n17769_1(.douta(w_n17769_1[0]),.doutb(w_n17769_1[1]),.doutc(w_n17769_1[2]),.din(w_n17769_0[0]));
	jspl3 jspl3_w_n17769_2(.douta(w_n17769_2[0]),.doutb(w_n17769_2[1]),.doutc(w_n17769_2[2]),.din(w_n17769_0[1]));
	jspl3 jspl3_w_n17769_3(.douta(w_n17769_3[0]),.doutb(w_n17769_3[1]),.doutc(w_n17769_3[2]),.din(w_n17769_0[2]));
	jspl3 jspl3_w_n17769_4(.douta(w_n17769_4[0]),.doutb(w_n17769_4[1]),.doutc(w_n17769_4[2]),.din(w_n17769_1[0]));
	jspl3 jspl3_w_n17769_5(.douta(w_n17769_5[0]),.doutb(w_n17769_5[1]),.doutc(w_n17769_5[2]),.din(w_n17769_1[1]));
	jspl3 jspl3_w_n17769_6(.douta(w_n17769_6[0]),.doutb(w_n17769_6[1]),.doutc(w_n17769_6[2]),.din(w_n17769_1[2]));
	jspl3 jspl3_w_n17769_7(.douta(w_n17769_7[0]),.doutb(w_n17769_7[1]),.doutc(w_n17769_7[2]),.din(w_n17769_2[0]));
	jspl3 jspl3_w_n17769_8(.douta(w_n17769_8[0]),.doutb(w_n17769_8[1]),.doutc(w_n17769_8[2]),.din(w_n17769_2[1]));
	jspl3 jspl3_w_n17769_9(.douta(w_n17769_9[0]),.doutb(w_n17769_9[1]),.doutc(w_n17769_9[2]),.din(w_n17769_2[2]));
	jspl3 jspl3_w_n17769_10(.douta(w_n17769_10[0]),.doutb(w_n17769_10[1]),.doutc(w_n17769_10[2]),.din(w_n17769_3[0]));
	jspl3 jspl3_w_n17769_11(.douta(w_n17769_11[0]),.doutb(w_n17769_11[1]),.doutc(w_n17769_11[2]),.din(w_n17769_3[1]));
	jspl3 jspl3_w_n17769_12(.douta(w_n17769_12[0]),.doutb(w_n17769_12[1]),.doutc(w_n17769_12[2]),.din(w_n17769_3[2]));
	jspl3 jspl3_w_n17769_13(.douta(w_n17769_13[0]),.doutb(w_n17769_13[1]),.doutc(w_n17769_13[2]),.din(w_n17769_4[0]));
	jspl3 jspl3_w_n17769_14(.douta(w_n17769_14[0]),.doutb(w_n17769_14[1]),.doutc(w_n17769_14[2]),.din(w_n17769_4[1]));
	jspl3 jspl3_w_n17769_15(.douta(w_n17769_15[0]),.doutb(w_n17769_15[1]),.doutc(w_n17769_15[2]),.din(w_n17769_4[2]));
	jspl3 jspl3_w_n17769_16(.douta(w_n17769_16[0]),.doutb(w_n17769_16[1]),.doutc(w_n17769_16[2]),.din(w_n17769_5[0]));
	jspl3 jspl3_w_n17769_17(.douta(w_n17769_17[0]),.doutb(w_n17769_17[1]),.doutc(w_n17769_17[2]),.din(w_n17769_5[1]));
	jspl3 jspl3_w_n17769_18(.douta(w_n17769_18[0]),.doutb(w_n17769_18[1]),.doutc(w_n17769_18[2]),.din(w_n17769_5[2]));
	jspl3 jspl3_w_n17769_19(.douta(w_n17769_19[0]),.doutb(w_n17769_19[1]),.doutc(w_n17769_19[2]),.din(w_n17769_6[0]));
	jspl3 jspl3_w_n17769_20(.douta(w_n17769_20[0]),.doutb(w_n17769_20[1]),.doutc(w_n17769_20[2]),.din(w_n17769_6[1]));
	jspl3 jspl3_w_n17769_21(.douta(w_n17769_21[0]),.doutb(w_n17769_21[1]),.doutc(w_n17769_21[2]),.din(w_n17769_6[2]));
	jspl3 jspl3_w_n17769_22(.douta(w_n17769_22[0]),.doutb(w_n17769_22[1]),.doutc(w_n17769_22[2]),.din(w_n17769_7[0]));
	jspl3 jspl3_w_n17769_23(.douta(w_n17769_23[0]),.doutb(w_n17769_23[1]),.doutc(w_n17769_23[2]),.din(w_n17769_7[1]));
	jspl3 jspl3_w_n17769_24(.douta(w_n17769_24[0]),.doutb(w_n17769_24[1]),.doutc(w_n17769_24[2]),.din(w_n17769_7[2]));
	jspl3 jspl3_w_n17769_25(.douta(w_n17769_25[0]),.doutb(w_n17769_25[1]),.doutc(w_n17769_25[2]),.din(w_n17769_8[0]));
	jspl3 jspl3_w_n17769_26(.douta(w_n17769_26[0]),.doutb(w_n17769_26[1]),.doutc(w_n17769_26[2]),.din(w_n17769_8[1]));
	jspl3 jspl3_w_n17769_27(.douta(w_n17769_27[0]),.doutb(w_n17769_27[1]),.doutc(w_n17769_27[2]),.din(w_n17769_8[2]));
	jspl3 jspl3_w_n17769_28(.douta(w_n17769_28[0]),.doutb(w_n17769_28[1]),.doutc(w_n17769_28[2]),.din(w_n17769_9[0]));
	jspl3 jspl3_w_n17769_29(.douta(w_n17769_29[0]),.doutb(w_n17769_29[1]),.doutc(w_n17769_29[2]),.din(w_n17769_9[1]));
	jspl3 jspl3_w_n17769_30(.douta(w_n17769_30[0]),.doutb(w_n17769_30[1]),.doutc(w_n17769_30[2]),.din(w_n17769_9[2]));
	jspl3 jspl3_w_n17769_31(.douta(w_n17769_31[0]),.doutb(w_n17769_31[1]),.doutc(w_n17769_31[2]),.din(w_n17769_10[0]));
	jspl3 jspl3_w_n17769_32(.douta(w_n17769_32[0]),.doutb(w_n17769_32[1]),.doutc(w_n17769_32[2]),.din(w_n17769_10[1]));
	jspl3 jspl3_w_n17769_33(.douta(w_n17769_33[0]),.doutb(w_n17769_33[1]),.doutc(w_n17769_33[2]),.din(w_n17769_10[2]));
	jspl3 jspl3_w_n17769_34(.douta(w_n17769_34[0]),.doutb(w_n17769_34[1]),.doutc(w_n17769_34[2]),.din(w_n17769_11[0]));
	jspl3 jspl3_w_n17769_35(.douta(w_n17769_35[0]),.doutb(w_n17769_35[1]),.doutc(w_n17769_35[2]),.din(w_n17769_11[1]));
	jspl3 jspl3_w_n17769_36(.douta(w_n17769_36[0]),.doutb(w_n17769_36[1]),.doutc(w_n17769_36[2]),.din(w_n17769_11[2]));
	jspl3 jspl3_w_n17769_37(.douta(w_n17769_37[0]),.doutb(w_n17769_37[1]),.doutc(w_n17769_37[2]),.din(w_n17769_12[0]));
	jspl jspl_w_n17769_38(.douta(w_n17769_38[0]),.doutb(w_n17769_38[1]),.din(w_n17769_12[1]));
	jspl jspl_w_n17772_0(.douta(w_n17772_0[0]),.doutb(w_n17772_0[1]),.din(n17772));
	jspl3 jspl3_w_n17773_0(.douta(w_n17773_0[0]),.doutb(w_n17773_0[1]),.doutc(w_n17773_0[2]),.din(n17773));
	jspl3 jspl3_w_n17774_0(.douta(w_n17774_0[0]),.doutb(w_n17774_0[1]),.doutc(w_n17774_0[2]),.din(n17774));
	jspl3 jspl3_w_n17774_1(.douta(w_n17774_1[0]),.doutb(w_n17774_1[1]),.doutc(w_n17774_1[2]),.din(w_n17774_0[0]));
	jspl jspl_w_n17775_0(.douta(w_n17775_0[0]),.doutb(w_n17775_0[1]),.din(n17775));
	jspl3 jspl3_w_n17776_0(.douta(w_n17776_0[0]),.doutb(w_n17776_0[1]),.doutc(w_n17776_0[2]),.din(n17776));
	jspl jspl_w_n17777_0(.douta(w_n17777_0[0]),.doutb(w_n17777_0[1]),.din(n17777));
	jspl3 jspl3_w_n17780_0(.douta(w_n17780_0[0]),.doutb(w_n17780_0[1]),.doutc(w_n17780_0[2]),.din(n17780));
	jspl jspl_w_n17781_0(.douta(w_n17781_0[0]),.doutb(w_n17781_0[1]),.din(n17781));
	jspl3 jspl3_w_n17788_0(.douta(w_n17788_0[0]),.doutb(w_n17788_0[1]),.doutc(w_n17788_0[2]),.din(n17788));
	jspl jspl_w_n17789_0(.douta(w_n17789_0[0]),.doutb(w_n17789_0[1]),.din(n17789));
	jspl jspl_w_n17792_0(.douta(w_n17792_0[0]),.doutb(w_n17792_0[1]),.din(n17792));
	jspl3 jspl3_w_n17797_0(.douta(w_n17797_0[0]),.doutb(w_n17797_0[1]),.doutc(w_n17797_0[2]),.din(n17797));
	jspl3 jspl3_w_n17799_0(.douta(w_n17799_0[0]),.doutb(w_n17799_0[1]),.doutc(w_n17799_0[2]),.din(n17799));
	jspl jspl_w_n17800_0(.douta(w_n17800_0[0]),.doutb(w_n17800_0[1]),.din(n17800));
	jspl3 jspl3_w_n17804_0(.douta(w_n17804_0[0]),.doutb(w_n17804_0[1]),.doutc(w_n17804_0[2]),.din(n17804));
	jspl3 jspl3_w_n17807_0(.douta(w_n17807_0[0]),.doutb(w_n17807_0[1]),.doutc(w_n17807_0[2]),.din(n17807));
	jspl jspl_w_n17808_0(.douta(w_n17808_0[0]),.doutb(w_n17808_0[1]),.din(n17808));
	jspl3 jspl3_w_n17812_0(.douta(w_n17812_0[0]),.doutb(w_n17812_0[1]),.doutc(w_n17812_0[2]),.din(n17812));
	jspl3 jspl3_w_n17814_0(.douta(w_n17814_0[0]),.doutb(w_n17814_0[1]),.doutc(w_n17814_0[2]),.din(n17814));
	jspl jspl_w_n17815_0(.douta(w_n17815_0[0]),.doutb(w_n17815_0[1]),.din(n17815));
	jspl3 jspl3_w_n17819_0(.douta(w_n17819_0[0]),.doutb(w_n17819_0[1]),.doutc(w_n17819_0[2]),.din(n17819));
	jspl3 jspl3_w_n17822_0(.douta(w_n17822_0[0]),.doutb(w_n17822_0[1]),.doutc(w_n17822_0[2]),.din(n17822));
	jspl jspl_w_n17823_0(.douta(w_n17823_0[0]),.doutb(w_n17823_0[1]),.din(n17823));
	jspl3 jspl3_w_n17827_0(.douta(w_n17827_0[0]),.doutb(w_n17827_0[1]),.doutc(w_n17827_0[2]),.din(n17827));
	jspl3 jspl3_w_n17829_0(.douta(w_n17829_0[0]),.doutb(w_n17829_0[1]),.doutc(w_n17829_0[2]),.din(n17829));
	jspl jspl_w_n17830_0(.douta(w_n17830_0[0]),.doutb(w_n17830_0[1]),.din(n17830));
	jspl3 jspl3_w_n17834_0(.douta(w_n17834_0[0]),.doutb(w_n17834_0[1]),.doutc(w_n17834_0[2]),.din(n17834));
	jspl3 jspl3_w_n17837_0(.douta(w_n17837_0[0]),.doutb(w_n17837_0[1]),.doutc(w_n17837_0[2]),.din(n17837));
	jspl jspl_w_n17838_0(.douta(w_n17838_0[0]),.doutb(w_n17838_0[1]),.din(n17838));
	jspl3 jspl3_w_n17842_0(.douta(w_n17842_0[0]),.doutb(w_n17842_0[1]),.doutc(w_n17842_0[2]),.din(n17842));
	jspl3 jspl3_w_n17844_0(.douta(w_n17844_0[0]),.doutb(w_n17844_0[1]),.doutc(w_n17844_0[2]),.din(n17844));
	jspl jspl_w_n17845_0(.douta(w_n17845_0[0]),.doutb(w_n17845_0[1]),.din(n17845));
	jspl3 jspl3_w_n17849_0(.douta(w_n17849_0[0]),.doutb(w_n17849_0[1]),.doutc(w_n17849_0[2]),.din(n17849));
	jspl3 jspl3_w_n17851_0(.douta(w_n17851_0[0]),.doutb(w_n17851_0[1]),.doutc(w_n17851_0[2]),.din(n17851));
	jspl jspl_w_n17852_0(.douta(w_n17852_0[0]),.doutb(w_n17852_0[1]),.din(n17852));
	jspl3 jspl3_w_n17856_0(.douta(w_n17856_0[0]),.doutb(w_n17856_0[1]),.doutc(w_n17856_0[2]),.din(n17856));
	jspl3 jspl3_w_n17859_0(.douta(w_n17859_0[0]),.doutb(w_n17859_0[1]),.doutc(w_n17859_0[2]),.din(n17859));
	jspl jspl_w_n17860_0(.douta(w_n17860_0[0]),.doutb(w_n17860_0[1]),.din(n17860));
	jspl3 jspl3_w_n17864_0(.douta(w_n17864_0[0]),.doutb(w_n17864_0[1]),.doutc(w_n17864_0[2]),.din(n17864));
	jspl3 jspl3_w_n17867_0(.douta(w_n17867_0[0]),.doutb(w_n17867_0[1]),.doutc(w_n17867_0[2]),.din(n17867));
	jspl jspl_w_n17868_0(.douta(w_n17868_0[0]),.doutb(w_n17868_0[1]),.din(n17868));
	jspl3 jspl3_w_n17872_0(.douta(w_n17872_0[0]),.doutb(w_n17872_0[1]),.doutc(w_n17872_0[2]),.din(n17872));
	jspl3 jspl3_w_n17874_0(.douta(w_n17874_0[0]),.doutb(w_n17874_0[1]),.doutc(w_n17874_0[2]),.din(n17874));
	jspl jspl_w_n17875_0(.douta(w_n17875_0[0]),.doutb(w_n17875_0[1]),.din(n17875));
	jspl3 jspl3_w_n17879_0(.douta(w_n17879_0[0]),.doutb(w_n17879_0[1]),.doutc(w_n17879_0[2]),.din(n17879));
	jspl3 jspl3_w_n17882_0(.douta(w_n17882_0[0]),.doutb(w_n17882_0[1]),.doutc(w_n17882_0[2]),.din(n17882));
	jspl jspl_w_n17883_0(.douta(w_n17883_0[0]),.doutb(w_n17883_0[1]),.din(n17883));
	jspl3 jspl3_w_n17887_0(.douta(w_n17887_0[0]),.doutb(w_n17887_0[1]),.doutc(w_n17887_0[2]),.din(n17887));
	jspl3 jspl3_w_n17889_0(.douta(w_n17889_0[0]),.doutb(w_n17889_0[1]),.doutc(w_n17889_0[2]),.din(n17889));
	jspl jspl_w_n17890_0(.douta(w_n17890_0[0]),.doutb(w_n17890_0[1]),.din(n17890));
	jspl3 jspl3_w_n17894_0(.douta(w_n17894_0[0]),.doutb(w_n17894_0[1]),.doutc(w_n17894_0[2]),.din(n17894));
	jspl3 jspl3_w_n17897_0(.douta(w_n17897_0[0]),.doutb(w_n17897_0[1]),.doutc(w_n17897_0[2]),.din(n17897));
	jspl jspl_w_n17898_0(.douta(w_n17898_0[0]),.doutb(w_n17898_0[1]),.din(n17898));
	jspl3 jspl3_w_n17902_0(.douta(w_n17902_0[0]),.doutb(w_n17902_0[1]),.doutc(w_n17902_0[2]),.din(n17902));
	jspl3 jspl3_w_n17904_0(.douta(w_n17904_0[0]),.doutb(w_n17904_0[1]),.doutc(w_n17904_0[2]),.din(n17904));
	jspl jspl_w_n17905_0(.douta(w_n17905_0[0]),.doutb(w_n17905_0[1]),.din(n17905));
	jspl3 jspl3_w_n17909_0(.douta(w_n17909_0[0]),.doutb(w_n17909_0[1]),.doutc(w_n17909_0[2]),.din(n17909));
	jspl3 jspl3_w_n17911_0(.douta(w_n17911_0[0]),.doutb(w_n17911_0[1]),.doutc(w_n17911_0[2]),.din(n17911));
	jspl jspl_w_n17912_0(.douta(w_n17912_0[0]),.doutb(w_n17912_0[1]),.din(n17912));
	jspl3 jspl3_w_n17916_0(.douta(w_n17916_0[0]),.doutb(w_n17916_0[1]),.doutc(w_n17916_0[2]),.din(n17916));
	jspl3 jspl3_w_n17918_0(.douta(w_n17918_0[0]),.doutb(w_n17918_0[1]),.doutc(w_n17918_0[2]),.din(n17918));
	jspl jspl_w_n17919_0(.douta(w_n17919_0[0]),.doutb(w_n17919_0[1]),.din(n17919));
	jspl3 jspl3_w_n17923_0(.douta(w_n17923_0[0]),.doutb(w_n17923_0[1]),.doutc(w_n17923_0[2]),.din(n17923));
	jspl3 jspl3_w_n17926_0(.douta(w_n17926_0[0]),.doutb(w_n17926_0[1]),.doutc(w_n17926_0[2]),.din(n17926));
	jspl jspl_w_n17927_0(.douta(w_n17927_0[0]),.doutb(w_n17927_0[1]),.din(n17927));
	jspl3 jspl3_w_n17931_0(.douta(w_n17931_0[0]),.doutb(w_n17931_0[1]),.doutc(w_n17931_0[2]),.din(n17931));
	jspl3 jspl3_w_n17933_0(.douta(w_n17933_0[0]),.doutb(w_n17933_0[1]),.doutc(w_n17933_0[2]),.din(n17933));
	jspl jspl_w_n17934_0(.douta(w_n17934_0[0]),.doutb(w_n17934_0[1]),.din(n17934));
	jspl3 jspl3_w_n17938_0(.douta(w_n17938_0[0]),.doutb(w_n17938_0[1]),.doutc(w_n17938_0[2]),.din(n17938));
	jspl3 jspl3_w_n17941_0(.douta(w_n17941_0[0]),.doutb(w_n17941_0[1]),.doutc(w_n17941_0[2]),.din(n17941));
	jspl jspl_w_n17942_0(.douta(w_n17942_0[0]),.doutb(w_n17942_0[1]),.din(n17942));
	jspl3 jspl3_w_n17946_0(.douta(w_n17946_0[0]),.doutb(w_n17946_0[1]),.doutc(w_n17946_0[2]),.din(n17946));
	jspl3 jspl3_w_n17948_0(.douta(w_n17948_0[0]),.doutb(w_n17948_0[1]),.doutc(w_n17948_0[2]),.din(n17948));
	jspl jspl_w_n17949_0(.douta(w_n17949_0[0]),.doutb(w_n17949_0[1]),.din(n17949));
	jspl3 jspl3_w_n17953_0(.douta(w_n17953_0[0]),.doutb(w_n17953_0[1]),.doutc(w_n17953_0[2]),.din(n17953));
	jspl3 jspl3_w_n17956_0(.douta(w_n17956_0[0]),.doutb(w_n17956_0[1]),.doutc(w_n17956_0[2]),.din(n17956));
	jspl jspl_w_n17957_0(.douta(w_n17957_0[0]),.doutb(w_n17957_0[1]),.din(n17957));
	jspl3 jspl3_w_n17961_0(.douta(w_n17961_0[0]),.doutb(w_n17961_0[1]),.doutc(w_n17961_0[2]),.din(n17961));
	jspl3 jspl3_w_n17963_0(.douta(w_n17963_0[0]),.doutb(w_n17963_0[1]),.doutc(w_n17963_0[2]),.din(n17963));
	jspl jspl_w_n17964_0(.douta(w_n17964_0[0]),.doutb(w_n17964_0[1]),.din(n17964));
	jspl3 jspl3_w_n17968_0(.douta(w_n17968_0[0]),.doutb(w_n17968_0[1]),.doutc(w_n17968_0[2]),.din(n17968));
	jspl3 jspl3_w_n17971_0(.douta(w_n17971_0[0]),.doutb(w_n17971_0[1]),.doutc(w_n17971_0[2]),.din(n17971));
	jspl jspl_w_n17972_0(.douta(w_n17972_0[0]),.doutb(w_n17972_0[1]),.din(n17972));
	jspl3 jspl3_w_n17976_0(.douta(w_n17976_0[0]),.doutb(w_n17976_0[1]),.doutc(w_n17976_0[2]),.din(n17976));
	jspl3 jspl3_w_n17978_0(.douta(w_n17978_0[0]),.doutb(w_n17978_0[1]),.doutc(w_n17978_0[2]),.din(n17978));
	jspl jspl_w_n17979_0(.douta(w_n17979_0[0]),.doutb(w_n17979_0[1]),.din(n17979));
	jspl3 jspl3_w_n17983_0(.douta(w_n17983_0[0]),.doutb(w_n17983_0[1]),.doutc(w_n17983_0[2]),.din(n17983));
	jspl3 jspl3_w_n17985_0(.douta(w_n17985_0[0]),.doutb(w_n17985_0[1]),.doutc(w_n17985_0[2]),.din(n17985));
	jspl jspl_w_n17986_0(.douta(w_n17986_0[0]),.doutb(w_n17986_0[1]),.din(n17986));
	jspl3 jspl3_w_n17990_0(.douta(w_n17990_0[0]),.doutb(w_n17990_0[1]),.doutc(w_n17990_0[2]),.din(n17990));
	jspl3 jspl3_w_n17992_0(.douta(w_n17992_0[0]),.doutb(w_n17992_0[1]),.doutc(w_n17992_0[2]),.din(n17992));
	jspl jspl_w_n17993_0(.douta(w_n17993_0[0]),.doutb(w_n17993_0[1]),.din(n17993));
	jspl3 jspl3_w_n17997_0(.douta(w_n17997_0[0]),.doutb(w_n17997_0[1]),.doutc(w_n17997_0[2]),.din(n17997));
	jspl3 jspl3_w_n18000_0(.douta(w_n18000_0[0]),.doutb(w_n18000_0[1]),.doutc(w_n18000_0[2]),.din(n18000));
	jspl jspl_w_n18001_0(.douta(w_n18001_0[0]),.doutb(w_n18001_0[1]),.din(n18001));
	jspl3 jspl3_w_n18005_0(.douta(w_n18005_0[0]),.doutb(w_n18005_0[1]),.doutc(w_n18005_0[2]),.din(n18005));
	jspl3 jspl3_w_n18007_0(.douta(w_n18007_0[0]),.doutb(w_n18007_0[1]),.doutc(w_n18007_0[2]),.din(n18007));
	jspl jspl_w_n18008_0(.douta(w_n18008_0[0]),.doutb(w_n18008_0[1]),.din(n18008));
	jspl jspl_w_n18012_0(.douta(w_n18012_0[0]),.doutb(w_n18012_0[1]),.din(n18012));
	jspl jspl_w_n18013_0(.douta(w_n18013_0[0]),.doutb(w_n18013_0[1]),.din(n18013));
	jspl3 jspl3_w_n18015_0(.douta(w_n18015_0[0]),.doutb(w_n18015_0[1]),.doutc(w_n18015_0[2]),.din(n18015));
	jspl jspl_w_n18016_0(.douta(w_n18016_0[0]),.doutb(w_n18016_0[1]),.din(n18016));
	jspl3 jspl3_w_n18020_0(.douta(w_n18020_0[0]),.doutb(w_n18020_0[1]),.doutc(w_n18020_0[2]),.din(n18020));
	jspl3 jspl3_w_n18022_0(.douta(w_n18022_0[0]),.doutb(w_n18022_0[1]),.doutc(w_n18022_0[2]),.din(n18022));
	jspl jspl_w_n18023_0(.douta(w_n18023_0[0]),.doutb(w_n18023_0[1]),.din(n18023));
	jspl3 jspl3_w_n18027_0(.douta(w_n18027_0[0]),.doutb(w_n18027_0[1]),.doutc(w_n18027_0[2]),.din(n18027));
	jspl3 jspl3_w_n18029_0(.douta(w_n18029_0[0]),.doutb(w_n18029_0[1]),.doutc(w_n18029_0[2]),.din(n18029));
	jspl jspl_w_n18030_0(.douta(w_n18030_0[0]),.doutb(w_n18030_0[1]),.din(n18030));
	jspl3 jspl3_w_n18034_0(.douta(w_n18034_0[0]),.doutb(w_n18034_0[1]),.doutc(w_n18034_0[2]),.din(n18034));
	jspl3 jspl3_w_n18036_0(.douta(w_n18036_0[0]),.doutb(w_n18036_0[1]),.doutc(w_n18036_0[2]),.din(n18036));
	jspl jspl_w_n18037_0(.douta(w_n18037_0[0]),.doutb(w_n18037_0[1]),.din(n18037));
	jspl3 jspl3_w_n18041_0(.douta(w_n18041_0[0]),.doutb(w_n18041_0[1]),.doutc(w_n18041_0[2]),.din(n18041));
	jspl3 jspl3_w_n18044_0(.douta(w_n18044_0[0]),.doutb(w_n18044_0[1]),.doutc(w_n18044_0[2]),.din(n18044));
	jspl jspl_w_n18045_0(.douta(w_n18045_0[0]),.doutb(w_n18045_0[1]),.din(n18045));
	jspl3 jspl3_w_n18049_0(.douta(w_n18049_0[0]),.doutb(w_n18049_0[1]),.doutc(w_n18049_0[2]),.din(n18049));
	jspl3 jspl3_w_n18051_0(.douta(w_n18051_0[0]),.doutb(w_n18051_0[1]),.doutc(w_n18051_0[2]),.din(n18051));
	jspl jspl_w_n18052_0(.douta(w_n18052_0[0]),.doutb(w_n18052_0[1]),.din(n18052));
	jspl3 jspl3_w_n18056_0(.douta(w_n18056_0[0]),.doutb(w_n18056_0[1]),.doutc(w_n18056_0[2]),.din(n18056));
	jspl3 jspl3_w_n18059_0(.douta(w_n18059_0[0]),.doutb(w_n18059_0[1]),.doutc(w_n18059_0[2]),.din(n18059));
	jspl jspl_w_n18060_0(.douta(w_n18060_0[0]),.doutb(w_n18060_0[1]),.din(n18060));
	jspl3 jspl3_w_n18064_0(.douta(w_n18064_0[0]),.doutb(w_n18064_0[1]),.doutc(w_n18064_0[2]),.din(n18064));
	jspl3 jspl3_w_n18066_0(.douta(w_n18066_0[0]),.doutb(w_n18066_0[1]),.doutc(w_n18066_0[2]),.din(n18066));
	jspl jspl_w_n18067_0(.douta(w_n18067_0[0]),.doutb(w_n18067_0[1]),.din(n18067));
	jspl3 jspl3_w_n18071_0(.douta(w_n18071_0[0]),.doutb(w_n18071_0[1]),.doutc(w_n18071_0[2]),.din(n18071));
	jspl3 jspl3_w_n18073_0(.douta(w_n18073_0[0]),.doutb(w_n18073_0[1]),.doutc(w_n18073_0[2]),.din(n18073));
	jspl jspl_w_n18074_0(.douta(w_n18074_0[0]),.doutb(w_n18074_0[1]),.din(n18074));
	jspl3 jspl3_w_n18078_0(.douta(w_n18078_0[0]),.doutb(w_n18078_0[1]),.doutc(w_n18078_0[2]),.din(n18078));
	jspl3 jspl3_w_n18081_0(.douta(w_n18081_0[0]),.doutb(w_n18081_0[1]),.doutc(w_n18081_0[2]),.din(n18081));
	jspl jspl_w_n18082_0(.douta(w_n18082_0[0]),.doutb(w_n18082_0[1]),.din(n18082));
	jspl3 jspl3_w_n18085_0(.douta(w_n18085_0[0]),.doutb(w_n18085_0[1]),.doutc(w_n18085_0[2]),.din(n18085));
	jspl3 jspl3_w_n18089_0(.douta(w_n18089_0[0]),.doutb(w_n18089_0[1]),.doutc(w_n18089_0[2]),.din(n18089));
	jspl jspl_w_n18090_0(.douta(w_n18090_0[0]),.doutb(w_n18090_0[1]),.din(n18090));
	jspl3 jspl3_w_n18094_0(.douta(w_n18094_0[0]),.doutb(w_n18094_0[1]),.doutc(w_n18094_0[2]),.din(n18094));
	jspl3 jspl3_w_n18096_0(.douta(w_n18096_0[0]),.doutb(w_n18096_0[1]),.doutc(w_n18096_0[2]),.din(n18096));
	jspl jspl_w_n18097_0(.douta(w_n18097_0[0]),.doutb(w_n18097_0[1]),.din(n18097));
	jspl3 jspl3_w_n18101_0(.douta(w_n18101_0[0]),.doutb(w_n18101_0[1]),.doutc(w_n18101_0[2]),.din(n18101));
	jspl3 jspl3_w_n18104_0(.douta(w_n18104_0[0]),.doutb(w_n18104_0[1]),.doutc(w_n18104_0[2]),.din(n18104));
	jspl jspl_w_n18105_0(.douta(w_n18105_0[0]),.doutb(w_n18105_0[1]),.din(n18105));
	jspl3 jspl3_w_n18109_0(.douta(w_n18109_0[0]),.doutb(w_n18109_0[1]),.doutc(w_n18109_0[2]),.din(n18109));
	jspl3 jspl3_w_n18111_0(.douta(w_n18111_0[0]),.doutb(w_n18111_0[1]),.doutc(w_n18111_0[2]),.din(n18111));
	jspl jspl_w_n18112_0(.douta(w_n18112_0[0]),.doutb(w_n18112_0[1]),.din(n18112));
	jspl3 jspl3_w_n18116_0(.douta(w_n18116_0[0]),.doutb(w_n18116_0[1]),.doutc(w_n18116_0[2]),.din(n18116));
	jspl3 jspl3_w_n18119_0(.douta(w_n18119_0[0]),.doutb(w_n18119_0[1]),.doutc(w_n18119_0[2]),.din(n18119));
	jspl jspl_w_n18120_0(.douta(w_n18120_0[0]),.doutb(w_n18120_0[1]),.din(n18120));
	jspl3 jspl3_w_n18124_0(.douta(w_n18124_0[0]),.doutb(w_n18124_0[1]),.doutc(w_n18124_0[2]),.din(n18124));
	jspl3 jspl3_w_n18126_0(.douta(w_n18126_0[0]),.doutb(w_n18126_0[1]),.doutc(w_n18126_0[2]),.din(n18126));
	jspl jspl_w_n18127_0(.douta(w_n18127_0[0]),.doutb(w_n18127_0[1]),.din(n18127));
	jspl3 jspl3_w_n18131_0(.douta(w_n18131_0[0]),.doutb(w_n18131_0[1]),.doutc(w_n18131_0[2]),.din(n18131));
	jspl3 jspl3_w_n18133_0(.douta(w_n18133_0[0]),.doutb(w_n18133_0[1]),.doutc(w_n18133_0[2]),.din(n18133));
	jspl jspl_w_n18134_0(.douta(w_n18134_0[0]),.doutb(w_n18134_0[1]),.din(n18134));
	jspl3 jspl3_w_n18138_0(.douta(w_n18138_0[0]),.doutb(w_n18138_0[1]),.doutc(w_n18138_0[2]),.din(n18138));
	jspl3 jspl3_w_n18140_0(.douta(w_n18140_0[0]),.doutb(w_n18140_0[1]),.doutc(w_n18140_0[2]),.din(n18140));
	jspl jspl_w_n18141_0(.douta(w_n18141_0[0]),.doutb(w_n18141_0[1]),.din(n18141));
	jspl3 jspl3_w_n18145_0(.douta(w_n18145_0[0]),.doutb(w_n18145_0[1]),.doutc(w_n18145_0[2]),.din(n18145));
	jspl3 jspl3_w_n18148_0(.douta(w_n18148_0[0]),.doutb(w_n18148_0[1]),.doutc(w_n18148_0[2]),.din(n18148));
	jspl jspl_w_n18149_0(.douta(w_n18149_0[0]),.doutb(w_n18149_0[1]),.din(n18149));
	jspl3 jspl3_w_n18153_0(.douta(w_n18153_0[0]),.doutb(w_n18153_0[1]),.doutc(w_n18153_0[2]),.din(n18153));
	jspl3 jspl3_w_n18155_0(.douta(w_n18155_0[0]),.doutb(w_n18155_0[1]),.doutc(w_n18155_0[2]),.din(n18155));
	jspl jspl_w_n18156_0(.douta(w_n18156_0[0]),.doutb(w_n18156_0[1]),.din(n18156));
	jspl3 jspl3_w_n18160_0(.douta(w_n18160_0[0]),.doutb(w_n18160_0[1]),.doutc(w_n18160_0[2]),.din(n18160));
	jspl3 jspl3_w_n18163_0(.douta(w_n18163_0[0]),.doutb(w_n18163_0[1]),.doutc(w_n18163_0[2]),.din(n18163));
	jspl3 jspl3_w_n18164_0(.douta(w_n18164_0[0]),.doutb(w_n18164_0[1]),.doutc(w_n18164_0[2]),.din(n18164));
	jspl jspl_w_n18168_0(.douta(w_n18168_0[0]),.doutb(w_n18168_0[1]),.din(n18168));
	jspl jspl_w_n18169_0(.douta(w_n18169_0[0]),.doutb(w_n18169_0[1]),.din(n18169));
	jspl jspl_w_n18171_0(.douta(w_n18171_0[0]),.doutb(w_n18171_0[1]),.din(n18171));
	jspl jspl_w_n18172_0(.douta(w_n18172_0[0]),.doutb(w_n18172_0[1]),.din(n18172));
	jspl jspl_w_n18176_0(.douta(w_n18176_0[0]),.doutb(w_n18176_0[1]),.din(n18176));
	jspl jspl_w_n18178_0(.douta(w_n18178_0[0]),.doutb(w_n18178_0[1]),.din(n18178));
	jspl3 jspl3_w_n18182_0(.douta(w_n18182_0[0]),.doutb(w_n18182_0[1]),.doutc(w_n18182_0[2]),.din(n18182));
	jspl jspl_w_n18182_1(.douta(w_n18182_1[0]),.doutb(w_n18182_1[1]),.din(w_n18182_0[0]));
	jspl jspl_w_n18183_0(.douta(w_n18183_0[0]),.doutb(w_n18183_0[1]),.din(n18183));
	jspl3 jspl3_w_n18185_0(.douta(w_n18185_0[0]),.doutb(w_n18185_0[1]),.doutc(w_n18185_0[2]),.din(n18185));
	jspl jspl_w_n18185_1(.douta(w_n18185_1[0]),.doutb(w_n18185_1[1]),.din(w_n18185_0[0]));
	jspl jspl_w_n18186_0(.douta(w_n18186_0[0]),.doutb(w_n18186_0[1]),.din(n18186));
	jspl3 jspl3_w_n18187_0(.douta(w_n18187_0[0]),.doutb(w_n18187_0[1]),.doutc(w_n18187_0[2]),.din(n18187));
	jspl jspl_w_n18188_0(.douta(w_n18188_0[0]),.doutb(w_n18188_0[1]),.din(n18188));
	jspl3 jspl3_w_n18189_0(.douta(w_n18189_0[0]),.doutb(w_n18189_0[1]),.doutc(w_n18189_0[2]),.din(n18189));
	jspl jspl_w_n18190_0(.douta(w_n18190_0[0]),.doutb(w_n18190_0[1]),.din(n18190));
	jspl3 jspl3_w_n18195_0(.douta(w_n18195_0[0]),.doutb(w_n18195_0[1]),.doutc(w_n18195_0[2]),.din(n18195));
	jspl jspl_w_n18253_0(.douta(w_n18253_0[0]),.doutb(w_n18253_0[1]),.din(n18253));
	jspl jspl_w_n18435_0(.douta(w_n18435_0[0]),.doutb(w_n18435_0[1]),.din(n18435));
	jspl jspl_w_n18438_0(.douta(w_n18438_0[0]),.doutb(w_n18438_0[1]),.din(n18438));
	jspl jspl_w_n18441_0(.douta(w_n18441_0[0]),.doutb(w_n18441_0[1]),.din(n18441));
	jspl3 jspl3_w_n18442_0(.douta(w_n18442_0[0]),.doutb(w_n18442_0[1]),.doutc(w_n18442_0[2]),.din(n18442));
	jspl3 jspl3_w_n18442_1(.douta(w_n18442_1[0]),.doutb(w_n18442_1[1]),.doutc(w_n18442_1[2]),.din(w_n18442_0[0]));
	jspl3 jspl3_w_n18442_2(.douta(w_n18442_2[0]),.doutb(w_n18442_2[1]),.doutc(w_n18442_2[2]),.din(w_n18442_0[1]));
	jspl3 jspl3_w_n18442_3(.douta(w_n18442_3[0]),.doutb(w_n18442_3[1]),.doutc(w_n18442_3[2]),.din(w_n18442_0[2]));
	jspl3 jspl3_w_n18442_4(.douta(w_n18442_4[0]),.doutb(w_n18442_4[1]),.doutc(w_n18442_4[2]),.din(w_n18442_1[0]));
	jspl3 jspl3_w_n18442_5(.douta(w_n18442_5[0]),.doutb(w_n18442_5[1]),.doutc(w_n18442_5[2]),.din(w_n18442_1[1]));
	jspl3 jspl3_w_n18442_6(.douta(w_n18442_6[0]),.doutb(w_n18442_6[1]),.doutc(w_n18442_6[2]),.din(w_n18442_1[2]));
	jspl3 jspl3_w_n18442_7(.douta(w_n18442_7[0]),.doutb(w_n18442_7[1]),.doutc(w_n18442_7[2]),.din(w_n18442_2[0]));
	jspl3 jspl3_w_n18442_8(.douta(w_n18442_8[0]),.doutb(w_n18442_8[1]),.doutc(w_n18442_8[2]),.din(w_n18442_2[1]));
	jspl3 jspl3_w_n18442_9(.douta(w_n18442_9[0]),.doutb(w_n18442_9[1]),.doutc(w_n18442_9[2]),.din(w_n18442_2[2]));
	jspl3 jspl3_w_n18442_10(.douta(w_n18442_10[0]),.doutb(w_n18442_10[1]),.doutc(w_n18442_10[2]),.din(w_n18442_3[0]));
	jspl3 jspl3_w_n18442_11(.douta(w_n18442_11[0]),.doutb(w_n18442_11[1]),.doutc(w_n18442_11[2]),.din(w_n18442_3[1]));
	jspl3 jspl3_w_n18442_12(.douta(w_n18442_12[0]),.doutb(w_n18442_12[1]),.doutc(w_n18442_12[2]),.din(w_n18442_3[2]));
	jspl3 jspl3_w_n18446_0(.douta(w_n18446_0[0]),.doutb(w_n18446_0[1]),.doutc(w_n18446_0[2]),.din(n18446));
	jspl jspl_w_n18447_0(.douta(w_n18447_0[0]),.doutb(w_n18447_0[1]),.din(n18447));
	jspl jspl_w_n18449_0(.douta(w_n18449_0[0]),.doutb(w_n18449_0[1]),.din(n18449));
	jspl jspl_w_n18454_0(.douta(w_n18454_0[0]),.doutb(w_n18454_0[1]),.din(n18454));
	jspl jspl_w_n18455_0(.douta(w_n18455_0[0]),.doutb(w_n18455_0[1]),.din(n18455));
	jspl3 jspl3_w_n18457_0(.douta(w_n18457_0[0]),.doutb(w_n18457_0[1]),.doutc(w_n18457_0[2]),.din(n18457));
	jspl jspl_w_n18458_0(.douta(w_n18458_0[0]),.doutb(w_n18458_0[1]),.din(n18458));
	jspl jspl_w_n18462_0(.douta(w_n18462_0[0]),.doutb(w_n18462_0[1]),.din(n18462));
	jspl3 jspl3_w_n18464_0(.douta(w_n18464_0[0]),.doutb(w_n18464_0[1]),.doutc(w_n18464_0[2]),.din(n18464));
	jspl jspl_w_n18465_0(.douta(w_n18465_0[0]),.doutb(w_n18465_0[1]),.din(n18465));
	jspl jspl_w_n18469_0(.douta(w_n18469_0[0]),.doutb(w_n18469_0[1]),.din(n18469));
	jspl jspl_w_n18470_0(.douta(w_n18470_0[0]),.doutb(w_n18470_0[1]),.din(n18470));
	jspl3 jspl3_w_n18472_0(.douta(w_n18472_0[0]),.doutb(w_n18472_0[1]),.doutc(w_n18472_0[2]),.din(n18472));
	jspl jspl_w_n18473_0(.douta(w_n18473_0[0]),.doutb(w_n18473_0[1]),.din(n18473));
	jspl jspl_w_n18477_0(.douta(w_n18477_0[0]),.doutb(w_n18477_0[1]),.din(n18477));
	jspl3 jspl3_w_n18479_0(.douta(w_n18479_0[0]),.doutb(w_n18479_0[1]),.doutc(w_n18479_0[2]),.din(n18479));
	jspl jspl_w_n18480_0(.douta(w_n18480_0[0]),.doutb(w_n18480_0[1]),.din(n18480));
	jspl jspl_w_n18484_0(.douta(w_n18484_0[0]),.doutb(w_n18484_0[1]),.din(n18484));
	jspl jspl_w_n18485_0(.douta(w_n18485_0[0]),.doutb(w_n18485_0[1]),.din(n18485));
	jspl3 jspl3_w_n18487_0(.douta(w_n18487_0[0]),.doutb(w_n18487_0[1]),.doutc(w_n18487_0[2]),.din(n18487));
	jspl jspl_w_n18488_0(.douta(w_n18488_0[0]),.doutb(w_n18488_0[1]),.din(n18488));
	jspl jspl_w_n18492_0(.douta(w_n18492_0[0]),.doutb(w_n18492_0[1]),.din(n18492));
	jspl3 jspl3_w_n18494_0(.douta(w_n18494_0[0]),.doutb(w_n18494_0[1]),.doutc(w_n18494_0[2]),.din(n18494));
	jspl jspl_w_n18495_0(.douta(w_n18495_0[0]),.doutb(w_n18495_0[1]),.din(n18495));
	jspl jspl_w_n18499_0(.douta(w_n18499_0[0]),.doutb(w_n18499_0[1]),.din(n18499));
	jspl jspl_w_n18500_0(.douta(w_n18500_0[0]),.doutb(w_n18500_0[1]),.din(n18500));
	jspl3 jspl3_w_n18502_0(.douta(w_n18502_0[0]),.doutb(w_n18502_0[1]),.doutc(w_n18502_0[2]),.din(n18502));
	jspl jspl_w_n18503_0(.douta(w_n18503_0[0]),.doutb(w_n18503_0[1]),.din(n18503));
	jspl jspl_w_n18507_0(.douta(w_n18507_0[0]),.doutb(w_n18507_0[1]),.din(n18507));
	jspl3 jspl3_w_n18509_0(.douta(w_n18509_0[0]),.doutb(w_n18509_0[1]),.doutc(w_n18509_0[2]),.din(n18509));
	jspl jspl_w_n18510_0(.douta(w_n18510_0[0]),.doutb(w_n18510_0[1]),.din(n18510));
	jspl jspl_w_n18514_0(.douta(w_n18514_0[0]),.doutb(w_n18514_0[1]),.din(n18514));
	jspl jspl_w_n18515_0(.douta(w_n18515_0[0]),.doutb(w_n18515_0[1]),.din(n18515));
	jspl3 jspl3_w_n18517_0(.douta(w_n18517_0[0]),.doutb(w_n18517_0[1]),.doutc(w_n18517_0[2]),.din(n18517));
	jspl jspl_w_n18518_0(.douta(w_n18518_0[0]),.doutb(w_n18518_0[1]),.din(n18518));
	jspl jspl_w_n18522_0(.douta(w_n18522_0[0]),.doutb(w_n18522_0[1]),.din(n18522));
	jspl jspl_w_n18523_0(.douta(w_n18523_0[0]),.doutb(w_n18523_0[1]),.din(n18523));
	jspl3 jspl3_w_n18525_0(.douta(w_n18525_0[0]),.doutb(w_n18525_0[1]),.doutc(w_n18525_0[2]),.din(n18525));
	jspl jspl_w_n18526_0(.douta(w_n18526_0[0]),.doutb(w_n18526_0[1]),.din(n18526));
	jspl jspl_w_n18530_0(.douta(w_n18530_0[0]),.doutb(w_n18530_0[1]),.din(n18530));
	jspl3 jspl3_w_n18532_0(.douta(w_n18532_0[0]),.doutb(w_n18532_0[1]),.doutc(w_n18532_0[2]),.din(n18532));
	jspl jspl_w_n18533_0(.douta(w_n18533_0[0]),.doutb(w_n18533_0[1]),.din(n18533));
	jspl jspl_w_n18537_0(.douta(w_n18537_0[0]),.doutb(w_n18537_0[1]),.din(n18537));
	jspl3 jspl3_w_n18539_0(.douta(w_n18539_0[0]),.doutb(w_n18539_0[1]),.doutc(w_n18539_0[2]),.din(n18539));
	jspl jspl_w_n18540_0(.douta(w_n18540_0[0]),.doutb(w_n18540_0[1]),.din(n18540));
	jspl jspl_w_n18544_0(.douta(w_n18544_0[0]),.doutb(w_n18544_0[1]),.din(n18544));
	jspl jspl_w_n18545_0(.douta(w_n18545_0[0]),.doutb(w_n18545_0[1]),.din(n18545));
	jspl3 jspl3_w_n18547_0(.douta(w_n18547_0[0]),.doutb(w_n18547_0[1]),.doutc(w_n18547_0[2]),.din(n18547));
	jspl jspl_w_n18548_0(.douta(w_n18548_0[0]),.doutb(w_n18548_0[1]),.din(n18548));
	jspl jspl_w_n18552_0(.douta(w_n18552_0[0]),.doutb(w_n18552_0[1]),.din(n18552));
	jspl3 jspl3_w_n18554_0(.douta(w_n18554_0[0]),.doutb(w_n18554_0[1]),.doutc(w_n18554_0[2]),.din(n18554));
	jspl jspl_w_n18555_0(.douta(w_n18555_0[0]),.doutb(w_n18555_0[1]),.din(n18555));
	jspl jspl_w_n18559_0(.douta(w_n18559_0[0]),.doutb(w_n18559_0[1]),.din(n18559));
	jspl jspl_w_n18560_0(.douta(w_n18560_0[0]),.doutb(w_n18560_0[1]),.din(n18560));
	jspl3 jspl3_w_n18562_0(.douta(w_n18562_0[0]),.doutb(w_n18562_0[1]),.doutc(w_n18562_0[2]),.din(n18562));
	jspl jspl_w_n18563_0(.douta(w_n18563_0[0]),.doutb(w_n18563_0[1]),.din(n18563));
	jspl jspl_w_n18567_0(.douta(w_n18567_0[0]),.doutb(w_n18567_0[1]),.din(n18567));
	jspl3 jspl3_w_n18569_0(.douta(w_n18569_0[0]),.doutb(w_n18569_0[1]),.doutc(w_n18569_0[2]),.din(n18569));
	jspl jspl_w_n18570_0(.douta(w_n18570_0[0]),.doutb(w_n18570_0[1]),.din(n18570));
	jspl jspl_w_n18574_0(.douta(w_n18574_0[0]),.doutb(w_n18574_0[1]),.din(n18574));
	jspl jspl_w_n18575_0(.douta(w_n18575_0[0]),.doutb(w_n18575_0[1]),.din(n18575));
	jspl3 jspl3_w_n18577_0(.douta(w_n18577_0[0]),.doutb(w_n18577_0[1]),.doutc(w_n18577_0[2]),.din(n18577));
	jspl jspl_w_n18578_0(.douta(w_n18578_0[0]),.doutb(w_n18578_0[1]),.din(n18578));
	jspl jspl_w_n18582_0(.douta(w_n18582_0[0]),.doutb(w_n18582_0[1]),.din(n18582));
	jspl jspl_w_n18583_0(.douta(w_n18583_0[0]),.doutb(w_n18583_0[1]),.din(n18583));
	jspl3 jspl3_w_n18585_0(.douta(w_n18585_0[0]),.doutb(w_n18585_0[1]),.doutc(w_n18585_0[2]),.din(n18585));
	jspl jspl_w_n18586_0(.douta(w_n18586_0[0]),.doutb(w_n18586_0[1]),.din(n18586));
	jspl jspl_w_n18590_0(.douta(w_n18590_0[0]),.doutb(w_n18590_0[1]),.din(n18590));
	jspl jspl_w_n18591_0(.douta(w_n18591_0[0]),.doutb(w_n18591_0[1]),.din(n18591));
	jspl3 jspl3_w_n18593_0(.douta(w_n18593_0[0]),.doutb(w_n18593_0[1]),.doutc(w_n18593_0[2]),.din(n18593));
	jspl jspl_w_n18594_0(.douta(w_n18594_0[0]),.doutb(w_n18594_0[1]),.din(n18594));
	jspl jspl_w_n18598_0(.douta(w_n18598_0[0]),.doutb(w_n18598_0[1]),.din(n18598));
	jspl3 jspl3_w_n18600_0(.douta(w_n18600_0[0]),.doutb(w_n18600_0[1]),.doutc(w_n18600_0[2]),.din(n18600));
	jspl jspl_w_n18601_0(.douta(w_n18601_0[0]),.doutb(w_n18601_0[1]),.din(n18601));
	jspl jspl_w_n18605_0(.douta(w_n18605_0[0]),.doutb(w_n18605_0[1]),.din(n18605));
	jspl jspl_w_n18606_0(.douta(w_n18606_0[0]),.doutb(w_n18606_0[1]),.din(n18606));
	jspl3 jspl3_w_n18608_0(.douta(w_n18608_0[0]),.doutb(w_n18608_0[1]),.doutc(w_n18608_0[2]),.din(n18608));
	jspl jspl_w_n18609_0(.douta(w_n18609_0[0]),.doutb(w_n18609_0[1]),.din(n18609));
	jspl jspl_w_n18613_0(.douta(w_n18613_0[0]),.doutb(w_n18613_0[1]),.din(n18613));
	jspl3 jspl3_w_n18615_0(.douta(w_n18615_0[0]),.doutb(w_n18615_0[1]),.doutc(w_n18615_0[2]),.din(n18615));
	jspl jspl_w_n18616_0(.douta(w_n18616_0[0]),.doutb(w_n18616_0[1]),.din(n18616));
	jspl jspl_w_n18620_0(.douta(w_n18620_0[0]),.doutb(w_n18620_0[1]),.din(n18620));
	jspl jspl_w_n18621_0(.douta(w_n18621_0[0]),.doutb(w_n18621_0[1]),.din(n18621));
	jspl3 jspl3_w_n18623_0(.douta(w_n18623_0[0]),.doutb(w_n18623_0[1]),.doutc(w_n18623_0[2]),.din(n18623));
	jspl jspl_w_n18624_0(.douta(w_n18624_0[0]),.doutb(w_n18624_0[1]),.din(n18624));
	jspl jspl_w_n18628_0(.douta(w_n18628_0[0]),.doutb(w_n18628_0[1]),.din(n18628));
	jspl3 jspl3_w_n18630_0(.douta(w_n18630_0[0]),.doutb(w_n18630_0[1]),.doutc(w_n18630_0[2]),.din(n18630));
	jspl jspl_w_n18631_0(.douta(w_n18631_0[0]),.doutb(w_n18631_0[1]),.din(n18631));
	jspl jspl_w_n18635_0(.douta(w_n18635_0[0]),.doutb(w_n18635_0[1]),.din(n18635));
	jspl jspl_w_n18636_0(.douta(w_n18636_0[0]),.doutb(w_n18636_0[1]),.din(n18636));
	jspl3 jspl3_w_n18638_0(.douta(w_n18638_0[0]),.doutb(w_n18638_0[1]),.doutc(w_n18638_0[2]),.din(n18638));
	jspl jspl_w_n18639_0(.douta(w_n18639_0[0]),.doutb(w_n18639_0[1]),.din(n18639));
	jspl jspl_w_n18643_0(.douta(w_n18643_0[0]),.doutb(w_n18643_0[1]),.din(n18643));
	jspl3 jspl3_w_n18645_0(.douta(w_n18645_0[0]),.doutb(w_n18645_0[1]),.doutc(w_n18645_0[2]),.din(n18645));
	jspl jspl_w_n18646_0(.douta(w_n18646_0[0]),.doutb(w_n18646_0[1]),.din(n18646));
	jspl jspl_w_n18650_0(.douta(w_n18650_0[0]),.doutb(w_n18650_0[1]),.din(n18650));
	jspl jspl_w_n18651_0(.douta(w_n18651_0[0]),.doutb(w_n18651_0[1]),.din(n18651));
	jspl3 jspl3_w_n18653_0(.douta(w_n18653_0[0]),.doutb(w_n18653_0[1]),.doutc(w_n18653_0[2]),.din(n18653));
	jspl jspl_w_n18654_0(.douta(w_n18654_0[0]),.doutb(w_n18654_0[1]),.din(n18654));
	jspl jspl_w_n18658_0(.douta(w_n18658_0[0]),.doutb(w_n18658_0[1]),.din(n18658));
	jspl jspl_w_n18659_0(.douta(w_n18659_0[0]),.doutb(w_n18659_0[1]),.din(n18659));
	jspl3 jspl3_w_n18661_0(.douta(w_n18661_0[0]),.doutb(w_n18661_0[1]),.doutc(w_n18661_0[2]),.din(n18661));
	jspl jspl_w_n18662_0(.douta(w_n18662_0[0]),.doutb(w_n18662_0[1]),.din(n18662));
	jspl jspl_w_n18666_0(.douta(w_n18666_0[0]),.doutb(w_n18666_0[1]),.din(n18666));
	jspl jspl_w_n18667_0(.douta(w_n18667_0[0]),.doutb(w_n18667_0[1]),.din(n18667));
	jspl3 jspl3_w_n18669_0(.douta(w_n18669_0[0]),.doutb(w_n18669_0[1]),.doutc(w_n18669_0[2]),.din(n18669));
	jspl jspl_w_n18670_0(.douta(w_n18670_0[0]),.doutb(w_n18670_0[1]),.din(n18670));
	jspl jspl_w_n18674_0(.douta(w_n18674_0[0]),.doutb(w_n18674_0[1]),.din(n18674));
	jspl3 jspl3_w_n18676_0(.douta(w_n18676_0[0]),.doutb(w_n18676_0[1]),.doutc(w_n18676_0[2]),.din(n18676));
	jspl jspl_w_n18677_0(.douta(w_n18677_0[0]),.doutb(w_n18677_0[1]),.din(n18677));
	jspl jspl_w_n18681_0(.douta(w_n18681_0[0]),.doutb(w_n18681_0[1]),.din(n18681));
	jspl jspl_w_n18682_0(.douta(w_n18682_0[0]),.doutb(w_n18682_0[1]),.din(n18682));
	jspl3 jspl3_w_n18684_0(.douta(w_n18684_0[0]),.doutb(w_n18684_0[1]),.doutc(w_n18684_0[2]),.din(n18684));
	jspl jspl_w_n18685_0(.douta(w_n18685_0[0]),.doutb(w_n18685_0[1]),.din(n18685));
	jspl jspl_w_n18689_0(.douta(w_n18689_0[0]),.doutb(w_n18689_0[1]),.din(n18689));
	jspl jspl_w_n18690_0(.douta(w_n18690_0[0]),.doutb(w_n18690_0[1]),.din(n18690));
	jspl3 jspl3_w_n18692_0(.douta(w_n18692_0[0]),.doutb(w_n18692_0[1]),.doutc(w_n18692_0[2]),.din(n18692));
	jspl jspl_w_n18693_0(.douta(w_n18693_0[0]),.doutb(w_n18693_0[1]),.din(n18693));
	jspl jspl_w_n18697_0(.douta(w_n18697_0[0]),.doutb(w_n18697_0[1]),.din(n18697));
	jspl jspl_w_n18698_0(.douta(w_n18698_0[0]),.doutb(w_n18698_0[1]),.din(n18698));
	jspl3 jspl3_w_n18700_0(.douta(w_n18700_0[0]),.doutb(w_n18700_0[1]),.doutc(w_n18700_0[2]),.din(n18700));
	jspl jspl_w_n18701_0(.douta(w_n18701_0[0]),.doutb(w_n18701_0[1]),.din(n18701));
	jspl jspl_w_n18705_0(.douta(w_n18705_0[0]),.doutb(w_n18705_0[1]),.din(n18705));
	jspl jspl_w_n18706_0(.douta(w_n18706_0[0]),.doutb(w_n18706_0[1]),.din(n18706));
	jspl3 jspl3_w_n18708_0(.douta(w_n18708_0[0]),.doutb(w_n18708_0[1]),.doutc(w_n18708_0[2]),.din(n18708));
	jspl jspl_w_n18709_0(.douta(w_n18709_0[0]),.doutb(w_n18709_0[1]),.din(n18709));
	jspl jspl_w_n18713_0(.douta(w_n18713_0[0]),.doutb(w_n18713_0[1]),.din(n18713));
	jspl jspl_w_n18714_0(.douta(w_n18714_0[0]),.doutb(w_n18714_0[1]),.din(n18714));
	jspl3 jspl3_w_n18716_0(.douta(w_n18716_0[0]),.doutb(w_n18716_0[1]),.doutc(w_n18716_0[2]),.din(n18716));
	jspl jspl_w_n18717_0(.douta(w_n18717_0[0]),.doutb(w_n18717_0[1]),.din(n18717));
	jspl jspl_w_n18721_0(.douta(w_n18721_0[0]),.doutb(w_n18721_0[1]),.din(n18721));
	jspl3 jspl3_w_n18723_0(.douta(w_n18723_0[0]),.doutb(w_n18723_0[1]),.doutc(w_n18723_0[2]),.din(n18723));
	jspl jspl_w_n18724_0(.douta(w_n18724_0[0]),.doutb(w_n18724_0[1]),.din(n18724));
	jspl jspl_w_n18728_0(.douta(w_n18728_0[0]),.doutb(w_n18728_0[1]),.din(n18728));
	jspl jspl_w_n18729_0(.douta(w_n18729_0[0]),.doutb(w_n18729_0[1]),.din(n18729));
	jspl3 jspl3_w_n18731_0(.douta(w_n18731_0[0]),.doutb(w_n18731_0[1]),.doutc(w_n18731_0[2]),.din(n18731));
	jspl jspl_w_n18732_0(.douta(w_n18732_0[0]),.doutb(w_n18732_0[1]),.din(n18732));
	jspl jspl_w_n18736_0(.douta(w_n18736_0[0]),.doutb(w_n18736_0[1]),.din(n18736));
	jspl3 jspl3_w_n18738_0(.douta(w_n18738_0[0]),.doutb(w_n18738_0[1]),.doutc(w_n18738_0[2]),.din(n18738));
	jspl jspl_w_n18739_0(.douta(w_n18739_0[0]),.doutb(w_n18739_0[1]),.din(n18739));
	jspl jspl_w_n18743_0(.douta(w_n18743_0[0]),.doutb(w_n18743_0[1]),.din(n18743));
	jspl jspl_w_n18744_0(.douta(w_n18744_0[0]),.doutb(w_n18744_0[1]),.din(n18744));
	jspl3 jspl3_w_n18746_0(.douta(w_n18746_0[0]),.doutb(w_n18746_0[1]),.doutc(w_n18746_0[2]),.din(n18746));
	jspl jspl_w_n18747_0(.douta(w_n18747_0[0]),.doutb(w_n18747_0[1]),.din(n18747));
	jspl jspl_w_n18751_0(.douta(w_n18751_0[0]),.doutb(w_n18751_0[1]),.din(n18751));
	jspl jspl_w_n18752_0(.douta(w_n18752_0[0]),.doutb(w_n18752_0[1]),.din(n18752));
	jspl3 jspl3_w_n18754_0(.douta(w_n18754_0[0]),.doutb(w_n18754_0[1]),.doutc(w_n18754_0[2]),.din(n18754));
	jspl jspl_w_n18755_0(.douta(w_n18755_0[0]),.doutb(w_n18755_0[1]),.din(n18755));
	jspl jspl_w_n18759_0(.douta(w_n18759_0[0]),.doutb(w_n18759_0[1]),.din(n18759));
	jspl3 jspl3_w_n18761_0(.douta(w_n18761_0[0]),.doutb(w_n18761_0[1]),.doutc(w_n18761_0[2]),.din(n18761));
	jspl jspl_w_n18762_0(.douta(w_n18762_0[0]),.doutb(w_n18762_0[1]),.din(n18762));
	jspl jspl_w_n18765_0(.douta(w_n18765_0[0]),.doutb(w_n18765_0[1]),.din(n18765));
	jspl3 jspl3_w_n18768_0(.douta(w_n18768_0[0]),.doutb(w_n18768_0[1]),.doutc(w_n18768_0[2]),.din(n18768));
	jspl jspl_w_n18769_0(.douta(w_n18769_0[0]),.doutb(w_n18769_0[1]),.din(n18769));
	jspl jspl_w_n18773_0(.douta(w_n18773_0[0]),.doutb(w_n18773_0[1]),.din(n18773));
	jspl jspl_w_n18774_0(.douta(w_n18774_0[0]),.doutb(w_n18774_0[1]),.din(n18774));
	jspl3 jspl3_w_n18776_0(.douta(w_n18776_0[0]),.doutb(w_n18776_0[1]),.doutc(w_n18776_0[2]),.din(n18776));
	jspl jspl_w_n18777_0(.douta(w_n18777_0[0]),.doutb(w_n18777_0[1]),.din(n18777));
	jspl jspl_w_n18781_0(.douta(w_n18781_0[0]),.doutb(w_n18781_0[1]),.din(n18781));
	jspl3 jspl3_w_n18783_0(.douta(w_n18783_0[0]),.doutb(w_n18783_0[1]),.doutc(w_n18783_0[2]),.din(n18783));
	jspl jspl_w_n18784_0(.douta(w_n18784_0[0]),.doutb(w_n18784_0[1]),.din(n18784));
	jspl jspl_w_n18788_0(.douta(w_n18788_0[0]),.doutb(w_n18788_0[1]),.din(n18788));
	jspl jspl_w_n18789_0(.douta(w_n18789_0[0]),.doutb(w_n18789_0[1]),.din(n18789));
	jspl3 jspl3_w_n18791_0(.douta(w_n18791_0[0]),.doutb(w_n18791_0[1]),.doutc(w_n18791_0[2]),.din(n18791));
	jspl jspl_w_n18792_0(.douta(w_n18792_0[0]),.doutb(w_n18792_0[1]),.din(n18792));
	jspl jspl_w_n18796_0(.douta(w_n18796_0[0]),.doutb(w_n18796_0[1]),.din(n18796));
	jspl3 jspl3_w_n18798_0(.douta(w_n18798_0[0]),.doutb(w_n18798_0[1]),.doutc(w_n18798_0[2]),.din(n18798));
	jspl jspl_w_n18799_0(.douta(w_n18799_0[0]),.doutb(w_n18799_0[1]),.din(n18799));
	jspl3 jspl3_w_n18803_0(.douta(w_n18803_0[0]),.doutb(w_n18803_0[1]),.doutc(w_n18803_0[2]),.din(n18803));
	jspl3 jspl3_w_n18806_0(.douta(w_n18806_0[0]),.doutb(w_n18806_0[1]),.doutc(w_n18806_0[2]),.din(n18806));
	jspl jspl_w_n18807_0(.douta(w_n18807_0[0]),.doutb(w_n18807_0[1]),.din(n18807));
	jspl jspl_w_n18811_0(.douta(w_n18811_0[0]),.doutb(w_n18811_0[1]),.din(n18811));
	jspl jspl_w_n18812_0(.douta(w_n18812_0[0]),.doutb(w_n18812_0[1]),.din(n18812));
	jspl3 jspl3_w_n18814_0(.douta(w_n18814_0[0]),.doutb(w_n18814_0[1]),.doutc(w_n18814_0[2]),.din(n18814));
	jspl jspl_w_n18815_0(.douta(w_n18815_0[0]),.doutb(w_n18815_0[1]),.din(n18815));
	jspl jspl_w_n18819_0(.douta(w_n18819_0[0]),.doutb(w_n18819_0[1]),.din(n18819));
	jspl jspl_w_n18820_0(.douta(w_n18820_0[0]),.doutb(w_n18820_0[1]),.din(n18820));
	jspl3 jspl3_w_n18822_0(.douta(w_n18822_0[0]),.doutb(w_n18822_0[1]),.doutc(w_n18822_0[2]),.din(n18822));
	jspl jspl_w_n18823_0(.douta(w_n18823_0[0]),.doutb(w_n18823_0[1]),.din(n18823));
	jspl jspl_w_n18827_0(.douta(w_n18827_0[0]),.doutb(w_n18827_0[1]),.din(n18827));
	jspl3 jspl3_w_n18829_0(.douta(w_n18829_0[0]),.doutb(w_n18829_0[1]),.doutc(w_n18829_0[2]),.din(n18829));
	jspl jspl_w_n18830_0(.douta(w_n18830_0[0]),.doutb(w_n18830_0[1]),.din(n18830));
	jspl jspl_w_n18841_0(.douta(w_n18841_0[0]),.doutb(w_n18841_0[1]),.din(n18841));
	jspl jspl_w_n18890_0(.douta(w_n18890_0[0]),.doutb(w_n18890_0[1]),.din(n18890));
	jspl jspl_w_n18897_0(.douta(w_n18897_0[0]),.doutb(w_n18897_0[1]),.din(n18897));
	jspl jspl_w_n18904_0(.douta(w_n18904_0[0]),.doutb(w_n18904_0[1]),.din(n18904));
	jspl jspl_w_n18911_0(.douta(w_n18911_0[0]),.doutb(w_n18911_0[1]),.din(n18911));
	jspl jspl_w_n18918_0(.douta(w_n18918_0[0]),.doutb(w_n18918_0[1]),.din(n18918));
	jspl jspl_w_n18928_0(.douta(w_n18928_0[0]),.doutb(w_n18928_0[1]),.din(n18928));
	jspl jspl_w_n18932_0(.douta(w_n18932_0[0]),.doutb(w_n18932_0[1]),.din(n18932));
	jspl jspl_w_n18939_0(.douta(w_n18939_0[0]),.doutb(w_n18939_0[1]),.din(n18939));
	jspl jspl_w_n18946_0(.douta(w_n18946_0[0]),.doutb(w_n18946_0[1]),.din(n18946));
	jspl jspl_w_n18959_0(.douta(w_n18959_0[0]),.doutb(w_n18959_0[1]),.din(n18959));
	jspl jspl_w_n18966_0(.douta(w_n18966_0[0]),.doutb(w_n18966_0[1]),.din(n18966));
	jspl jspl_w_n18973_0(.douta(w_n18973_0[0]),.doutb(w_n18973_0[1]),.din(n18973));
	jspl jspl_w_n18980_0(.douta(w_n18980_0[0]),.doutb(w_n18980_0[1]),.din(n18980));
	jspl jspl_w_n18993_0(.douta(w_n18993_0[0]),.doutb(w_n18993_0[1]),.din(n18993));
	jspl jspl_w_n19012_0(.douta(w_n19012_0[0]),.doutb(w_n19012_0[1]),.din(n19012));
	jspl jspl_w_n19019_0(.douta(w_n19019_0[0]),.doutb(w_n19019_0[1]),.din(n19019));
	jspl jspl_w_n19029_0(.douta(w_n19029_0[0]),.doutb(w_n19029_0[1]),.din(n19029));
	jspl jspl_w_n19039_0(.douta(w_n19039_0[0]),.doutb(w_n19039_0[1]),.din(n19039));
	jspl jspl_w_n19046_0(.douta(w_n19046_0[0]),.doutb(w_n19046_0[1]),.din(n19046));
	jspl jspl_w_n19059_0(.douta(w_n19059_0[0]),.doutb(w_n19059_0[1]),.din(n19059));
	jspl3 jspl3_w_n19065_0(.douta(w_n19065_0[0]),.doutb(w_n19065_0[1]),.doutc(w_n19065_0[2]),.din(n19065));
	jspl jspl_w_n19067_0(.douta(w_n19067_0[0]),.doutb(w_n19067_0[1]),.din(n19067));
	jspl jspl_w_n19068_0(.douta(w_n19068_0[0]),.doutb(w_n19068_0[1]),.din(n19068));
	jspl jspl_w_n19070_0(.douta(w_n19070_0[0]),.doutb(w_n19070_0[1]),.din(n19070));
	jspl jspl_w_n19072_0(.douta(w_n19072_0[0]),.doutb(w_n19072_0[1]),.din(n19072));
	jspl jspl_w_n19073_0(.douta(w_n19073_0[0]),.doutb(w_n19073_0[1]),.din(n19073));
	jspl3 jspl3_w_n19074_0(.douta(w_n19074_0[0]),.doutb(w_n19074_0[1]),.doutc(w_n19074_0[2]),.din(n19074));
	jspl jspl_w_n19079_0(.douta(w_n19079_0[0]),.doutb(w_n19079_0[1]),.din(n19079));
	jspl jspl_w_n19080_0(.douta(w_n19080_0[0]),.doutb(w_n19080_0[1]),.din(n19080));
	jspl3 jspl3_w_n19086_0(.douta(w_n19086_0[0]),.doutb(w_n19086_0[1]),.doutc(w_n19086_0[2]),.din(n19086));
	jspl jspl_w_n19087_0(.douta(w_n19087_0[0]),.doutb(w_n19087_0[1]),.din(n19087));
	jspl3 jspl3_w_n19096_0(.douta(w_n19096_0[0]),.doutb(w_n19096_0[1]),.doutc(w_n19096_0[2]),.din(n19096));
	jspl3 jspl3_w_n19096_1(.douta(w_n19096_1[0]),.doutb(w_n19096_1[1]),.doutc(w_n19096_1[2]),.din(w_n19096_0[0]));
	jspl3 jspl3_w_n19096_2(.douta(w_n19096_2[0]),.doutb(w_n19096_2[1]),.doutc(w_n19096_2[2]),.din(w_n19096_0[1]));
	jspl3 jspl3_w_n19096_3(.douta(w_n19096_3[0]),.doutb(w_n19096_3[1]),.doutc(w_n19096_3[2]),.din(w_n19096_0[2]));
	jspl3 jspl3_w_n19096_4(.douta(w_n19096_4[0]),.doutb(w_n19096_4[1]),.doutc(w_n19096_4[2]),.din(w_n19096_1[0]));
	jspl3 jspl3_w_n19096_5(.douta(w_n19096_5[0]),.doutb(w_n19096_5[1]),.doutc(w_n19096_5[2]),.din(w_n19096_1[1]));
	jspl3 jspl3_w_n19096_6(.douta(w_n19096_6[0]),.doutb(w_n19096_6[1]),.doutc(w_n19096_6[2]),.din(w_n19096_1[2]));
	jspl3 jspl3_w_n19096_7(.douta(w_n19096_7[0]),.doutb(w_n19096_7[1]),.doutc(w_n19096_7[2]),.din(w_n19096_2[0]));
	jspl3 jspl3_w_n19096_8(.douta(w_n19096_8[0]),.doutb(w_n19096_8[1]),.doutc(w_n19096_8[2]),.din(w_n19096_2[1]));
	jspl3 jspl3_w_n19096_9(.douta(w_n19096_9[0]),.doutb(w_n19096_9[1]),.doutc(w_n19096_9[2]),.din(w_n19096_2[2]));
	jspl3 jspl3_w_n19096_10(.douta(w_n19096_10[0]),.doutb(w_n19096_10[1]),.doutc(w_n19096_10[2]),.din(w_n19096_3[0]));
	jspl3 jspl3_w_n19096_11(.douta(w_n19096_11[0]),.doutb(w_n19096_11[1]),.doutc(w_n19096_11[2]),.din(w_n19096_3[1]));
	jspl3 jspl3_w_n19096_12(.douta(w_n19096_12[0]),.doutb(w_n19096_12[1]),.doutc(w_n19096_12[2]),.din(w_n19096_3[2]));
	jspl3 jspl3_w_n19096_13(.douta(w_n19096_13[0]),.doutb(w_n19096_13[1]),.doutc(w_n19096_13[2]),.din(w_n19096_4[0]));
	jspl3 jspl3_w_n19096_14(.douta(w_n19096_14[0]),.doutb(w_n19096_14[1]),.doutc(w_n19096_14[2]),.din(w_n19096_4[1]));
	jspl3 jspl3_w_n19096_15(.douta(w_n19096_15[0]),.doutb(w_n19096_15[1]),.doutc(w_n19096_15[2]),.din(w_n19096_4[2]));
	jspl3 jspl3_w_n19096_16(.douta(w_n19096_16[0]),.doutb(w_n19096_16[1]),.doutc(w_n19096_16[2]),.din(w_n19096_5[0]));
	jspl3 jspl3_w_n19096_17(.douta(w_n19096_17[0]),.doutb(w_n19096_17[1]),.doutc(w_n19096_17[2]),.din(w_n19096_5[1]));
	jspl3 jspl3_w_n19096_18(.douta(w_n19096_18[0]),.doutb(w_n19096_18[1]),.doutc(w_n19096_18[2]),.din(w_n19096_5[2]));
	jspl3 jspl3_w_n19096_19(.douta(w_n19096_19[0]),.doutb(w_n19096_19[1]),.doutc(w_n19096_19[2]),.din(w_n19096_6[0]));
	jspl3 jspl3_w_n19096_20(.douta(w_n19096_20[0]),.doutb(w_n19096_20[1]),.doutc(w_n19096_20[2]),.din(w_n19096_6[1]));
	jspl3 jspl3_w_n19096_21(.douta(w_n19096_21[0]),.doutb(w_n19096_21[1]),.doutc(w_n19096_21[2]),.din(w_n19096_6[2]));
	jspl3 jspl3_w_n19096_22(.douta(w_n19096_22[0]),.doutb(w_n19096_22[1]),.doutc(w_n19096_22[2]),.din(w_n19096_7[0]));
	jspl3 jspl3_w_n19096_23(.douta(w_n19096_23[0]),.doutb(w_n19096_23[1]),.doutc(w_n19096_23[2]),.din(w_n19096_7[1]));
	jspl3 jspl3_w_n19096_24(.douta(w_n19096_24[0]),.doutb(w_n19096_24[1]),.doutc(w_n19096_24[2]),.din(w_n19096_7[2]));
	jspl3 jspl3_w_n19096_25(.douta(w_n19096_25[0]),.doutb(w_n19096_25[1]),.doutc(w_n19096_25[2]),.din(w_n19096_8[0]));
	jspl3 jspl3_w_n19096_26(.douta(w_n19096_26[0]),.doutb(w_n19096_26[1]),.doutc(w_n19096_26[2]),.din(w_n19096_8[1]));
	jspl3 jspl3_w_n19096_27(.douta(w_n19096_27[0]),.doutb(w_n19096_27[1]),.doutc(w_n19096_27[2]),.din(w_n19096_8[2]));
	jspl3 jspl3_w_n19096_28(.douta(w_n19096_28[0]),.doutb(w_n19096_28[1]),.doutc(w_n19096_28[2]),.din(w_n19096_9[0]));
	jspl3 jspl3_w_n19096_29(.douta(w_n19096_29[0]),.doutb(w_n19096_29[1]),.doutc(w_n19096_29[2]),.din(w_n19096_9[1]));
	jspl3 jspl3_w_n19096_30(.douta(w_n19096_30[0]),.doutb(w_n19096_30[1]),.doutc(w_n19096_30[2]),.din(w_n19096_9[2]));
	jspl3 jspl3_w_n19096_31(.douta(w_n19096_31[0]),.doutb(w_n19096_31[1]),.doutc(w_n19096_31[2]),.din(w_n19096_10[0]));
	jspl3 jspl3_w_n19096_32(.douta(w_n19096_32[0]),.doutb(w_n19096_32[1]),.doutc(w_n19096_32[2]),.din(w_n19096_10[1]));
	jspl3 jspl3_w_n19096_33(.douta(w_n19096_33[0]),.doutb(w_n19096_33[1]),.doutc(w_n19096_33[2]),.din(w_n19096_10[2]));
	jspl3 jspl3_w_n19096_34(.douta(w_n19096_34[0]),.doutb(w_n19096_34[1]),.doutc(w_n19096_34[2]),.din(w_n19096_11[0]));
	jspl3 jspl3_w_n19096_35(.douta(w_n19096_35[0]),.doutb(w_n19096_35[1]),.doutc(w_n19096_35[2]),.din(w_n19096_11[1]));
	jspl jspl_w_n19096_36(.douta(w_n19096_36[0]),.doutb(w_n19096_36[1]),.din(w_n19096_11[2]));
	jspl3 jspl3_w_n19099_0(.douta(w_n19099_0[0]),.doutb(w_n19099_0[1]),.doutc(w_n19099_0[2]),.din(n19099));
	jspl3 jspl3_w_n19100_0(.douta(w_n19100_0[0]),.doutb(w_n19100_0[1]),.doutc(w_n19100_0[2]),.din(n19100));
	jspl3 jspl3_w_n19101_0(.douta(w_n19101_0[0]),.doutb(w_n19101_0[1]),.doutc(w_n19101_0[2]),.din(n19101));
	jspl3 jspl3_w_n19101_1(.douta(w_n19101_1[0]),.doutb(w_n19101_1[1]),.doutc(w_n19101_1[2]),.din(w_n19101_0[0]));
	jspl jspl_w_n19102_0(.douta(w_n19102_0[0]),.doutb(w_n19102_0[1]),.din(n19102));
	jspl3 jspl3_w_n19103_0(.douta(w_n19103_0[0]),.doutb(w_n19103_0[1]),.doutc(w_n19103_0[2]),.din(n19103));
	jspl jspl_w_n19104_0(.douta(w_n19104_0[0]),.doutb(w_n19104_0[1]),.din(n19104));
	jspl3 jspl3_w_n19107_0(.douta(w_n19107_0[0]),.doutb(w_n19107_0[1]),.doutc(w_n19107_0[2]),.din(n19107));
	jspl jspl_w_n19108_0(.douta(w_n19108_0[0]),.doutb(w_n19108_0[1]),.din(n19108));
	jspl jspl_w_n19113_0(.douta(w_n19113_0[0]),.doutb(w_n19113_0[1]),.din(n19113));
	jspl3 jspl3_w_n19115_0(.douta(w_n19115_0[0]),.doutb(w_n19115_0[1]),.doutc(w_n19115_0[2]),.din(n19115));
	jspl jspl_w_n19116_0(.douta(w_n19116_0[0]),.doutb(w_n19116_0[1]),.din(n19116));
	jspl jspl_w_n19119_0(.douta(w_n19119_0[0]),.doutb(w_n19119_0[1]),.din(n19119));
	jspl3 jspl3_w_n19124_0(.douta(w_n19124_0[0]),.doutb(w_n19124_0[1]),.doutc(w_n19124_0[2]),.din(n19124));
	jspl3 jspl3_w_n19126_0(.douta(w_n19126_0[0]),.doutb(w_n19126_0[1]),.doutc(w_n19126_0[2]),.din(n19126));
	jspl jspl_w_n19127_0(.douta(w_n19127_0[0]),.doutb(w_n19127_0[1]),.din(n19127));
	jspl3 jspl3_w_n19131_0(.douta(w_n19131_0[0]),.doutb(w_n19131_0[1]),.doutc(w_n19131_0[2]),.din(n19131));
	jspl3 jspl3_w_n19134_0(.douta(w_n19134_0[0]),.doutb(w_n19134_0[1]),.doutc(w_n19134_0[2]),.din(n19134));
	jspl jspl_w_n19135_0(.douta(w_n19135_0[0]),.doutb(w_n19135_0[1]),.din(n19135));
	jspl3 jspl3_w_n19139_0(.douta(w_n19139_0[0]),.doutb(w_n19139_0[1]),.doutc(w_n19139_0[2]),.din(n19139));
	jspl3 jspl3_w_n19141_0(.douta(w_n19141_0[0]),.doutb(w_n19141_0[1]),.doutc(w_n19141_0[2]),.din(n19141));
	jspl jspl_w_n19142_0(.douta(w_n19142_0[0]),.doutb(w_n19142_0[1]),.din(n19142));
	jspl3 jspl3_w_n19146_0(.douta(w_n19146_0[0]),.doutb(w_n19146_0[1]),.doutc(w_n19146_0[2]),.din(n19146));
	jspl3 jspl3_w_n19149_0(.douta(w_n19149_0[0]),.doutb(w_n19149_0[1]),.doutc(w_n19149_0[2]),.din(n19149));
	jspl jspl_w_n19150_0(.douta(w_n19150_0[0]),.doutb(w_n19150_0[1]),.din(n19150));
	jspl3 jspl3_w_n19154_0(.douta(w_n19154_0[0]),.doutb(w_n19154_0[1]),.doutc(w_n19154_0[2]),.din(n19154));
	jspl3 jspl3_w_n19156_0(.douta(w_n19156_0[0]),.doutb(w_n19156_0[1]),.doutc(w_n19156_0[2]),.din(n19156));
	jspl jspl_w_n19157_0(.douta(w_n19157_0[0]),.doutb(w_n19157_0[1]),.din(n19157));
	jspl3 jspl3_w_n19161_0(.douta(w_n19161_0[0]),.doutb(w_n19161_0[1]),.doutc(w_n19161_0[2]),.din(n19161));
	jspl3 jspl3_w_n19164_0(.douta(w_n19164_0[0]),.doutb(w_n19164_0[1]),.doutc(w_n19164_0[2]),.din(n19164));
	jspl jspl_w_n19165_0(.douta(w_n19165_0[0]),.doutb(w_n19165_0[1]),.din(n19165));
	jspl3 jspl3_w_n19169_0(.douta(w_n19169_0[0]),.doutb(w_n19169_0[1]),.doutc(w_n19169_0[2]),.din(n19169));
	jspl3 jspl3_w_n19171_0(.douta(w_n19171_0[0]),.doutb(w_n19171_0[1]),.doutc(w_n19171_0[2]),.din(n19171));
	jspl jspl_w_n19172_0(.douta(w_n19172_0[0]),.doutb(w_n19172_0[1]),.din(n19172));
	jspl3 jspl3_w_n19176_0(.douta(w_n19176_0[0]),.doutb(w_n19176_0[1]),.doutc(w_n19176_0[2]),.din(n19176));
	jspl3 jspl3_w_n19179_0(.douta(w_n19179_0[0]),.doutb(w_n19179_0[1]),.doutc(w_n19179_0[2]),.din(n19179));
	jspl jspl_w_n19180_0(.douta(w_n19180_0[0]),.doutb(w_n19180_0[1]),.din(n19180));
	jspl3 jspl3_w_n19184_0(.douta(w_n19184_0[0]),.doutb(w_n19184_0[1]),.doutc(w_n19184_0[2]),.din(n19184));
	jspl3 jspl3_w_n19186_0(.douta(w_n19186_0[0]),.doutb(w_n19186_0[1]),.doutc(w_n19186_0[2]),.din(n19186));
	jspl jspl_w_n19187_0(.douta(w_n19187_0[0]),.doutb(w_n19187_0[1]),.din(n19187));
	jspl3 jspl3_w_n19191_0(.douta(w_n19191_0[0]),.doutb(w_n19191_0[1]),.doutc(w_n19191_0[2]),.din(n19191));
	jspl3 jspl3_w_n19194_0(.douta(w_n19194_0[0]),.doutb(w_n19194_0[1]),.doutc(w_n19194_0[2]),.din(n19194));
	jspl jspl_w_n19195_0(.douta(w_n19195_0[0]),.doutb(w_n19195_0[1]),.din(n19195));
	jspl3 jspl3_w_n19199_0(.douta(w_n19199_0[0]),.doutb(w_n19199_0[1]),.doutc(w_n19199_0[2]),.din(n19199));
	jspl3 jspl3_w_n19201_0(.douta(w_n19201_0[0]),.doutb(w_n19201_0[1]),.doutc(w_n19201_0[2]),.din(n19201));
	jspl jspl_w_n19202_0(.douta(w_n19202_0[0]),.doutb(w_n19202_0[1]),.din(n19202));
	jspl3 jspl3_w_n19206_0(.douta(w_n19206_0[0]),.doutb(w_n19206_0[1]),.doutc(w_n19206_0[2]),.din(n19206));
	jspl3 jspl3_w_n19208_0(.douta(w_n19208_0[0]),.doutb(w_n19208_0[1]),.doutc(w_n19208_0[2]),.din(n19208));
	jspl jspl_w_n19209_0(.douta(w_n19209_0[0]),.doutb(w_n19209_0[1]),.din(n19209));
	jspl3 jspl3_w_n19213_0(.douta(w_n19213_0[0]),.doutb(w_n19213_0[1]),.doutc(w_n19213_0[2]),.din(n19213));
	jspl3 jspl3_w_n19216_0(.douta(w_n19216_0[0]),.doutb(w_n19216_0[1]),.doutc(w_n19216_0[2]),.din(n19216));
	jspl jspl_w_n19217_0(.douta(w_n19217_0[0]),.doutb(w_n19217_0[1]),.din(n19217));
	jspl3 jspl3_w_n19221_0(.douta(w_n19221_0[0]),.doutb(w_n19221_0[1]),.doutc(w_n19221_0[2]),.din(n19221));
	jspl3 jspl3_w_n19224_0(.douta(w_n19224_0[0]),.doutb(w_n19224_0[1]),.doutc(w_n19224_0[2]),.din(n19224));
	jspl jspl_w_n19225_0(.douta(w_n19225_0[0]),.doutb(w_n19225_0[1]),.din(n19225));
	jspl3 jspl3_w_n19229_0(.douta(w_n19229_0[0]),.doutb(w_n19229_0[1]),.doutc(w_n19229_0[2]),.din(n19229));
	jspl3 jspl3_w_n19231_0(.douta(w_n19231_0[0]),.doutb(w_n19231_0[1]),.doutc(w_n19231_0[2]),.din(n19231));
	jspl jspl_w_n19232_0(.douta(w_n19232_0[0]),.doutb(w_n19232_0[1]),.din(n19232));
	jspl3 jspl3_w_n19236_0(.douta(w_n19236_0[0]),.doutb(w_n19236_0[1]),.doutc(w_n19236_0[2]),.din(n19236));
	jspl3 jspl3_w_n19239_0(.douta(w_n19239_0[0]),.doutb(w_n19239_0[1]),.doutc(w_n19239_0[2]),.din(n19239));
	jspl jspl_w_n19240_0(.douta(w_n19240_0[0]),.doutb(w_n19240_0[1]),.din(n19240));
	jspl3 jspl3_w_n19244_0(.douta(w_n19244_0[0]),.doutb(w_n19244_0[1]),.doutc(w_n19244_0[2]),.din(n19244));
	jspl3 jspl3_w_n19246_0(.douta(w_n19246_0[0]),.doutb(w_n19246_0[1]),.doutc(w_n19246_0[2]),.din(n19246));
	jspl jspl_w_n19247_0(.douta(w_n19247_0[0]),.doutb(w_n19247_0[1]),.din(n19247));
	jspl3 jspl3_w_n19251_0(.douta(w_n19251_0[0]),.doutb(w_n19251_0[1]),.doutc(w_n19251_0[2]),.din(n19251));
	jspl3 jspl3_w_n19254_0(.douta(w_n19254_0[0]),.doutb(w_n19254_0[1]),.doutc(w_n19254_0[2]),.din(n19254));
	jspl jspl_w_n19255_0(.douta(w_n19255_0[0]),.doutb(w_n19255_0[1]),.din(n19255));
	jspl3 jspl3_w_n19259_0(.douta(w_n19259_0[0]),.doutb(w_n19259_0[1]),.doutc(w_n19259_0[2]),.din(n19259));
	jspl3 jspl3_w_n19261_0(.douta(w_n19261_0[0]),.doutb(w_n19261_0[1]),.doutc(w_n19261_0[2]),.din(n19261));
	jspl jspl_w_n19262_0(.douta(w_n19262_0[0]),.doutb(w_n19262_0[1]),.din(n19262));
	jspl3 jspl3_w_n19266_0(.douta(w_n19266_0[0]),.doutb(w_n19266_0[1]),.doutc(w_n19266_0[2]),.din(n19266));
	jspl3 jspl3_w_n19268_0(.douta(w_n19268_0[0]),.doutb(w_n19268_0[1]),.doutc(w_n19268_0[2]),.din(n19268));
	jspl jspl_w_n19269_0(.douta(w_n19269_0[0]),.doutb(w_n19269_0[1]),.din(n19269));
	jspl3 jspl3_w_n19273_0(.douta(w_n19273_0[0]),.doutb(w_n19273_0[1]),.doutc(w_n19273_0[2]),.din(n19273));
	jspl3 jspl3_w_n19275_0(.douta(w_n19275_0[0]),.doutb(w_n19275_0[1]),.doutc(w_n19275_0[2]),.din(n19275));
	jspl jspl_w_n19276_0(.douta(w_n19276_0[0]),.doutb(w_n19276_0[1]),.din(n19276));
	jspl3 jspl3_w_n19280_0(.douta(w_n19280_0[0]),.doutb(w_n19280_0[1]),.doutc(w_n19280_0[2]),.din(n19280));
	jspl3 jspl3_w_n19283_0(.douta(w_n19283_0[0]),.doutb(w_n19283_0[1]),.doutc(w_n19283_0[2]),.din(n19283));
	jspl jspl_w_n19284_0(.douta(w_n19284_0[0]),.doutb(w_n19284_0[1]),.din(n19284));
	jspl3 jspl3_w_n19288_0(.douta(w_n19288_0[0]),.doutb(w_n19288_0[1]),.doutc(w_n19288_0[2]),.din(n19288));
	jspl3 jspl3_w_n19290_0(.douta(w_n19290_0[0]),.doutb(w_n19290_0[1]),.doutc(w_n19290_0[2]),.din(n19290));
	jspl jspl_w_n19291_0(.douta(w_n19291_0[0]),.doutb(w_n19291_0[1]),.din(n19291));
	jspl3 jspl3_w_n19295_0(.douta(w_n19295_0[0]),.doutb(w_n19295_0[1]),.doutc(w_n19295_0[2]),.din(n19295));
	jspl3 jspl3_w_n19298_0(.douta(w_n19298_0[0]),.doutb(w_n19298_0[1]),.doutc(w_n19298_0[2]),.din(n19298));
	jspl jspl_w_n19299_0(.douta(w_n19299_0[0]),.doutb(w_n19299_0[1]),.din(n19299));
	jspl3 jspl3_w_n19303_0(.douta(w_n19303_0[0]),.doutb(w_n19303_0[1]),.doutc(w_n19303_0[2]),.din(n19303));
	jspl3 jspl3_w_n19305_0(.douta(w_n19305_0[0]),.doutb(w_n19305_0[1]),.doutc(w_n19305_0[2]),.din(n19305));
	jspl jspl_w_n19306_0(.douta(w_n19306_0[0]),.doutb(w_n19306_0[1]),.din(n19306));
	jspl3 jspl3_w_n19310_0(.douta(w_n19310_0[0]),.doutb(w_n19310_0[1]),.doutc(w_n19310_0[2]),.din(n19310));
	jspl3 jspl3_w_n19313_0(.douta(w_n19313_0[0]),.doutb(w_n19313_0[1]),.doutc(w_n19313_0[2]),.din(n19313));
	jspl jspl_w_n19314_0(.douta(w_n19314_0[0]),.doutb(w_n19314_0[1]),.din(n19314));
	jspl3 jspl3_w_n19318_0(.douta(w_n19318_0[0]),.doutb(w_n19318_0[1]),.doutc(w_n19318_0[2]),.din(n19318));
	jspl3 jspl3_w_n19320_0(.douta(w_n19320_0[0]),.doutb(w_n19320_0[1]),.doutc(w_n19320_0[2]),.din(n19320));
	jspl jspl_w_n19321_0(.douta(w_n19321_0[0]),.doutb(w_n19321_0[1]),.din(n19321));
	jspl3 jspl3_w_n19325_0(.douta(w_n19325_0[0]),.doutb(w_n19325_0[1]),.doutc(w_n19325_0[2]),.din(n19325));
	jspl3 jspl3_w_n19328_0(.douta(w_n19328_0[0]),.doutb(w_n19328_0[1]),.doutc(w_n19328_0[2]),.din(n19328));
	jspl jspl_w_n19329_0(.douta(w_n19329_0[0]),.doutb(w_n19329_0[1]),.din(n19329));
	jspl3 jspl3_w_n19333_0(.douta(w_n19333_0[0]),.doutb(w_n19333_0[1]),.doutc(w_n19333_0[2]),.din(n19333));
	jspl3 jspl3_w_n19335_0(.douta(w_n19335_0[0]),.doutb(w_n19335_0[1]),.doutc(w_n19335_0[2]),.din(n19335));
	jspl jspl_w_n19336_0(.douta(w_n19336_0[0]),.doutb(w_n19336_0[1]),.din(n19336));
	jspl3 jspl3_w_n19340_0(.douta(w_n19340_0[0]),.doutb(w_n19340_0[1]),.doutc(w_n19340_0[2]),.din(n19340));
	jspl3 jspl3_w_n19342_0(.douta(w_n19342_0[0]),.doutb(w_n19342_0[1]),.doutc(w_n19342_0[2]),.din(n19342));
	jspl jspl_w_n19343_0(.douta(w_n19343_0[0]),.doutb(w_n19343_0[1]),.din(n19343));
	jspl3 jspl3_w_n19347_0(.douta(w_n19347_0[0]),.doutb(w_n19347_0[1]),.doutc(w_n19347_0[2]),.din(n19347));
	jspl3 jspl3_w_n19349_0(.douta(w_n19349_0[0]),.doutb(w_n19349_0[1]),.doutc(w_n19349_0[2]),.din(n19349));
	jspl jspl_w_n19350_0(.douta(w_n19350_0[0]),.doutb(w_n19350_0[1]),.din(n19350));
	jspl3 jspl3_w_n19354_0(.douta(w_n19354_0[0]),.doutb(w_n19354_0[1]),.doutc(w_n19354_0[2]),.din(n19354));
	jspl3 jspl3_w_n19357_0(.douta(w_n19357_0[0]),.doutb(w_n19357_0[1]),.doutc(w_n19357_0[2]),.din(n19357));
	jspl jspl_w_n19358_0(.douta(w_n19358_0[0]),.doutb(w_n19358_0[1]),.din(n19358));
	jspl3 jspl3_w_n19362_0(.douta(w_n19362_0[0]),.doutb(w_n19362_0[1]),.doutc(w_n19362_0[2]),.din(n19362));
	jspl3 jspl3_w_n19364_0(.douta(w_n19364_0[0]),.doutb(w_n19364_0[1]),.doutc(w_n19364_0[2]),.din(n19364));
	jspl jspl_w_n19365_0(.douta(w_n19365_0[0]),.doutb(w_n19365_0[1]),.din(n19365));
	jspl3 jspl3_w_n19369_0(.douta(w_n19369_0[0]),.doutb(w_n19369_0[1]),.doutc(w_n19369_0[2]),.din(n19369));
	jspl3 jspl3_w_n19371_0(.douta(w_n19371_0[0]),.doutb(w_n19371_0[1]),.doutc(w_n19371_0[2]),.din(n19371));
	jspl jspl_w_n19372_0(.douta(w_n19372_0[0]),.doutb(w_n19372_0[1]),.din(n19372));
	jspl3 jspl3_w_n19376_0(.douta(w_n19376_0[0]),.doutb(w_n19376_0[1]),.doutc(w_n19376_0[2]),.din(n19376));
	jspl3 jspl3_w_n19378_0(.douta(w_n19378_0[0]),.doutb(w_n19378_0[1]),.doutc(w_n19378_0[2]),.din(n19378));
	jspl jspl_w_n19379_0(.douta(w_n19379_0[0]),.doutb(w_n19379_0[1]),.din(n19379));
	jspl3 jspl3_w_n19383_0(.douta(w_n19383_0[0]),.doutb(w_n19383_0[1]),.doutc(w_n19383_0[2]),.din(n19383));
	jspl3 jspl3_w_n19385_0(.douta(w_n19385_0[0]),.doutb(w_n19385_0[1]),.doutc(w_n19385_0[2]),.din(n19385));
	jspl jspl_w_n19386_0(.douta(w_n19386_0[0]),.doutb(w_n19386_0[1]),.din(n19386));
	jspl3 jspl3_w_n19390_0(.douta(w_n19390_0[0]),.doutb(w_n19390_0[1]),.doutc(w_n19390_0[2]),.din(n19390));
	jspl3 jspl3_w_n19392_0(.douta(w_n19392_0[0]),.doutb(w_n19392_0[1]),.doutc(w_n19392_0[2]),.din(n19392));
	jspl jspl_w_n19393_0(.douta(w_n19393_0[0]),.doutb(w_n19393_0[1]),.din(n19393));
	jspl3 jspl3_w_n19397_0(.douta(w_n19397_0[0]),.doutb(w_n19397_0[1]),.doutc(w_n19397_0[2]),.din(n19397));
	jspl3 jspl3_w_n19400_0(.douta(w_n19400_0[0]),.doutb(w_n19400_0[1]),.doutc(w_n19400_0[2]),.din(n19400));
	jspl jspl_w_n19401_0(.douta(w_n19401_0[0]),.doutb(w_n19401_0[1]),.din(n19401));
	jspl3 jspl3_w_n19405_0(.douta(w_n19405_0[0]),.doutb(w_n19405_0[1]),.doutc(w_n19405_0[2]),.din(n19405));
	jspl3 jspl3_w_n19407_0(.douta(w_n19407_0[0]),.doutb(w_n19407_0[1]),.doutc(w_n19407_0[2]),.din(n19407));
	jspl jspl_w_n19408_0(.douta(w_n19408_0[0]),.doutb(w_n19408_0[1]),.din(n19408));
	jspl3 jspl3_w_n19412_0(.douta(w_n19412_0[0]),.doutb(w_n19412_0[1]),.doutc(w_n19412_0[2]),.din(n19412));
	jspl3 jspl3_w_n19415_0(.douta(w_n19415_0[0]),.doutb(w_n19415_0[1]),.doutc(w_n19415_0[2]),.din(n19415));
	jspl jspl_w_n19416_0(.douta(w_n19416_0[0]),.doutb(w_n19416_0[1]),.din(n19416));
	jspl3 jspl3_w_n19420_0(.douta(w_n19420_0[0]),.doutb(w_n19420_0[1]),.doutc(w_n19420_0[2]),.din(n19420));
	jspl3 jspl3_w_n19422_0(.douta(w_n19422_0[0]),.doutb(w_n19422_0[1]),.doutc(w_n19422_0[2]),.din(n19422));
	jspl jspl_w_n19423_0(.douta(w_n19423_0[0]),.doutb(w_n19423_0[1]),.din(n19423));
	jspl3 jspl3_w_n19427_0(.douta(w_n19427_0[0]),.doutb(w_n19427_0[1]),.doutc(w_n19427_0[2]),.din(n19427));
	jspl3 jspl3_w_n19429_0(.douta(w_n19429_0[0]),.doutb(w_n19429_0[1]),.doutc(w_n19429_0[2]),.din(n19429));
	jspl jspl_w_n19430_0(.douta(w_n19430_0[0]),.doutb(w_n19430_0[1]),.din(n19430));
	jspl3 jspl3_w_n19434_0(.douta(w_n19434_0[0]),.doutb(w_n19434_0[1]),.doutc(w_n19434_0[2]),.din(n19434));
	jspl3 jspl3_w_n19437_0(.douta(w_n19437_0[0]),.doutb(w_n19437_0[1]),.doutc(w_n19437_0[2]),.din(n19437));
	jspl jspl_w_n19438_0(.douta(w_n19438_0[0]),.doutb(w_n19438_0[1]),.din(n19438));
	jspl3 jspl3_w_n19441_0(.douta(w_n19441_0[0]),.doutb(w_n19441_0[1]),.doutc(w_n19441_0[2]),.din(n19441));
	jspl3 jspl3_w_n19445_0(.douta(w_n19445_0[0]),.doutb(w_n19445_0[1]),.doutc(w_n19445_0[2]),.din(n19445));
	jspl jspl_w_n19446_0(.douta(w_n19446_0[0]),.doutb(w_n19446_0[1]),.din(n19446));
	jspl3 jspl3_w_n19450_0(.douta(w_n19450_0[0]),.doutb(w_n19450_0[1]),.doutc(w_n19450_0[2]),.din(n19450));
	jspl3 jspl3_w_n19452_0(.douta(w_n19452_0[0]),.doutb(w_n19452_0[1]),.doutc(w_n19452_0[2]),.din(n19452));
	jspl jspl_w_n19453_0(.douta(w_n19453_0[0]),.doutb(w_n19453_0[1]),.din(n19453));
	jspl3 jspl3_w_n19457_0(.douta(w_n19457_0[0]),.doutb(w_n19457_0[1]),.doutc(w_n19457_0[2]),.din(n19457));
	jspl3 jspl3_w_n19460_0(.douta(w_n19460_0[0]),.doutb(w_n19460_0[1]),.doutc(w_n19460_0[2]),.din(n19460));
	jspl jspl_w_n19461_0(.douta(w_n19461_0[0]),.doutb(w_n19461_0[1]),.din(n19461));
	jspl3 jspl3_w_n19465_0(.douta(w_n19465_0[0]),.doutb(w_n19465_0[1]),.doutc(w_n19465_0[2]),.din(n19465));
	jspl3 jspl3_w_n19467_0(.douta(w_n19467_0[0]),.doutb(w_n19467_0[1]),.doutc(w_n19467_0[2]),.din(n19467));
	jspl jspl_w_n19468_0(.douta(w_n19468_0[0]),.doutb(w_n19468_0[1]),.din(n19468));
	jspl jspl_w_n19472_0(.douta(w_n19472_0[0]),.doutb(w_n19472_0[1]),.din(n19472));
	jspl jspl_w_n19473_0(.douta(w_n19473_0[0]),.doutb(w_n19473_0[1]),.din(n19473));
	jspl3 jspl3_w_n19475_0(.douta(w_n19475_0[0]),.doutb(w_n19475_0[1]),.doutc(w_n19475_0[2]),.din(n19475));
	jspl jspl_w_n19476_0(.douta(w_n19476_0[0]),.doutb(w_n19476_0[1]),.din(n19476));
	jspl3 jspl3_w_n19480_0(.douta(w_n19480_0[0]),.doutb(w_n19480_0[1]),.doutc(w_n19480_0[2]),.din(n19480));
	jspl3 jspl3_w_n19483_0(.douta(w_n19483_0[0]),.doutb(w_n19483_0[1]),.doutc(w_n19483_0[2]),.din(n19483));
	jspl jspl_w_n19484_0(.douta(w_n19484_0[0]),.doutb(w_n19484_0[1]),.din(n19484));
	jspl3 jspl3_w_n19488_0(.douta(w_n19488_0[0]),.doutb(w_n19488_0[1]),.doutc(w_n19488_0[2]),.din(n19488));
	jspl3 jspl3_w_n19490_0(.douta(w_n19490_0[0]),.doutb(w_n19490_0[1]),.doutc(w_n19490_0[2]),.din(n19490));
	jspl jspl_w_n19491_0(.douta(w_n19491_0[0]),.doutb(w_n19491_0[1]),.din(n19491));
	jspl3 jspl3_w_n19495_0(.douta(w_n19495_0[0]),.doutb(w_n19495_0[1]),.doutc(w_n19495_0[2]),.din(n19495));
	jspl3 jspl3_w_n19497_0(.douta(w_n19497_0[0]),.doutb(w_n19497_0[1]),.doutc(w_n19497_0[2]),.din(n19497));
	jspl jspl_w_n19498_0(.douta(w_n19498_0[0]),.doutb(w_n19498_0[1]),.din(n19498));
	jspl3 jspl3_w_n19502_0(.douta(w_n19502_0[0]),.doutb(w_n19502_0[1]),.doutc(w_n19502_0[2]),.din(n19502));
	jspl3 jspl3_w_n19505_0(.douta(w_n19505_0[0]),.doutb(w_n19505_0[1]),.doutc(w_n19505_0[2]),.din(n19505));
	jspl jspl_w_n19506_0(.douta(w_n19506_0[0]),.doutb(w_n19506_0[1]),.din(n19506));
	jspl jspl_w_n19508_0(.douta(w_n19508_0[0]),.doutb(w_n19508_0[1]),.din(n19508));
	jspl jspl_w_n19511_0(.douta(w_n19511_0[0]),.doutb(w_n19511_0[1]),.din(n19511));
	jspl jspl_w_n19515_0(.douta(w_n19515_0[0]),.doutb(w_n19515_0[1]),.din(n19515));
	jspl3 jspl3_w_n19522_0(.douta(w_n19522_0[0]),.doutb(w_n19522_0[1]),.doutc(w_n19522_0[2]),.din(n19522));
	jspl3 jspl3_w_n19523_0(.douta(w_n19523_0[0]),.doutb(w_n19523_0[1]),.doutc(w_n19523_0[2]),.din(n19523));
	jspl3 jspl3_w_n19524_0(.douta(w_n19524_0[0]),.doutb(w_n19524_0[1]),.doutc(w_n19524_0[2]),.din(n19524));
	jspl jspl_w_n19524_1(.douta(w_n19524_1[0]),.doutb(w_n19524_1[1]),.din(w_n19524_0[0]));
	jspl jspl_w_n19525_0(.douta(w_n19525_0[0]),.doutb(w_n19525_0[1]),.din(n19525));
	jspl3 jspl3_w_n19526_0(.douta(w_n19526_0[0]),.doutb(w_n19526_0[1]),.doutc(w_n19526_0[2]),.din(n19526));
	jspl jspl_w_n19527_0(.douta(w_n19527_0[0]),.doutb(w_n19527_0[1]),.din(n19527));
	jspl3 jspl3_w_n19529_0(.douta(w_n19529_0[0]),.doutb(w_n19529_0[1]),.doutc(w_n19529_0[2]),.din(n19529));
	jspl jspl_w_n19530_0(.douta(w_n19530_0[0]),.doutb(w_n19530_0[1]),.din(n19530));
	jspl jspl_w_n19781_0(.douta(w_n19781_0[0]),.doutb(w_n19781_0[1]),.din(n19781));
	jspl jspl_w_n19782_0(.douta(w_n19782_0[0]),.doutb(w_n19782_0[1]),.din(n19782));
	jspl jspl_w_n19785_0(.douta(w_n19785_0[0]),.doutb(w_n19785_0[1]),.din(n19785));
	jspl jspl_w_n19786_0(.douta(w_n19786_0[0]),.doutb(w_n19786_0[1]),.din(n19786));
	jspl jspl_w_n19788_0(.douta(w_n19788_0[0]),.doutb(w_n19788_0[1]),.din(n19788));
	jspl3 jspl3_w_n19791_0(.douta(w_n19791_0[0]),.doutb(w_n19791_0[1]),.doutc(w_n19791_0[2]),.din(n19791));
	jspl3 jspl3_w_n19791_1(.douta(w_n19791_1[0]),.doutb(w_n19791_1[1]),.doutc(w_n19791_1[2]),.din(w_n19791_0[0]));
	jspl3 jspl3_w_n19791_2(.douta(w_n19791_2[0]),.doutb(w_n19791_2[1]),.doutc(w_n19791_2[2]),.din(w_n19791_0[1]));
	jspl3 jspl3_w_n19791_3(.douta(w_n19791_3[0]),.doutb(w_n19791_3[1]),.doutc(w_n19791_3[2]),.din(w_n19791_0[2]));
	jspl3 jspl3_w_n19791_4(.douta(w_n19791_4[0]),.doutb(w_n19791_4[1]),.doutc(w_n19791_4[2]),.din(w_n19791_1[0]));
	jspl3 jspl3_w_n19791_5(.douta(w_n19791_5[0]),.doutb(w_n19791_5[1]),.doutc(w_n19791_5[2]),.din(w_n19791_1[1]));
	jspl3 jspl3_w_n19791_6(.douta(w_n19791_6[0]),.doutb(w_n19791_6[1]),.doutc(w_n19791_6[2]),.din(w_n19791_1[2]));
	jspl3 jspl3_w_n19791_7(.douta(w_n19791_7[0]),.doutb(w_n19791_7[1]),.doutc(w_n19791_7[2]),.din(w_n19791_2[0]));
	jspl3 jspl3_w_n19791_8(.douta(w_n19791_8[0]),.doutb(w_n19791_8[1]),.doutc(w_n19791_8[2]),.din(w_n19791_2[1]));
	jspl3 jspl3_w_n19791_9(.douta(w_n19791_9[0]),.doutb(w_n19791_9[1]),.doutc(w_n19791_9[2]),.din(w_n19791_2[2]));
	jspl3 jspl3_w_n19791_10(.douta(w_n19791_10[0]),.doutb(w_n19791_10[1]),.doutc(w_n19791_10[2]),.din(w_n19791_3[0]));
	jspl3 jspl3_w_n19795_0(.douta(w_n19795_0[0]),.doutb(w_n19795_0[1]),.doutc(w_n19795_0[2]),.din(n19795));
	jspl jspl_w_n19796_0(.douta(w_n19796_0[0]),.doutb(w_n19796_0[1]),.din(n19796));
	jspl jspl_w_n19798_0(.douta(w_n19798_0[0]),.doutb(w_n19798_0[1]),.din(n19798));
	jspl jspl_w_n19802_0(.douta(w_n19802_0[0]),.doutb(w_n19802_0[1]),.din(n19802));
	jspl jspl_w_n19803_0(.douta(w_n19803_0[0]),.doutb(w_n19803_0[1]),.din(n19803));
	jspl3 jspl3_w_n19805_0(.douta(w_n19805_0[0]),.doutb(w_n19805_0[1]),.doutc(w_n19805_0[2]),.din(n19805));
	jspl jspl_w_n19806_0(.douta(w_n19806_0[0]),.doutb(w_n19806_0[1]),.din(n19806));
	jspl jspl_w_n19810_0(.douta(w_n19810_0[0]),.doutb(w_n19810_0[1]),.din(n19810));
	jspl jspl_w_n19811_0(.douta(w_n19811_0[0]),.doutb(w_n19811_0[1]),.din(n19811));
	jspl3 jspl3_w_n19813_0(.douta(w_n19813_0[0]),.doutb(w_n19813_0[1]),.doutc(w_n19813_0[2]),.din(n19813));
	jspl jspl_w_n19814_0(.douta(w_n19814_0[0]),.doutb(w_n19814_0[1]),.din(n19814));
	jspl jspl_w_n19818_0(.douta(w_n19818_0[0]),.doutb(w_n19818_0[1]),.din(n19818));
	jspl jspl_w_n19819_0(.douta(w_n19819_0[0]),.doutb(w_n19819_0[1]),.din(n19819));
	jspl3 jspl3_w_n19821_0(.douta(w_n19821_0[0]),.doutb(w_n19821_0[1]),.doutc(w_n19821_0[2]),.din(n19821));
	jspl jspl_w_n19822_0(.douta(w_n19822_0[0]),.doutb(w_n19822_0[1]),.din(n19822));
	jspl jspl_w_n19826_0(.douta(w_n19826_0[0]),.doutb(w_n19826_0[1]),.din(n19826));
	jspl3 jspl3_w_n19828_0(.douta(w_n19828_0[0]),.doutb(w_n19828_0[1]),.doutc(w_n19828_0[2]),.din(n19828));
	jspl jspl_w_n19829_0(.douta(w_n19829_0[0]),.doutb(w_n19829_0[1]),.din(n19829));
	jspl jspl_w_n19833_0(.douta(w_n19833_0[0]),.doutb(w_n19833_0[1]),.din(n19833));
	jspl jspl_w_n19834_0(.douta(w_n19834_0[0]),.doutb(w_n19834_0[1]),.din(n19834));
	jspl3 jspl3_w_n19836_0(.douta(w_n19836_0[0]),.doutb(w_n19836_0[1]),.doutc(w_n19836_0[2]),.din(n19836));
	jspl jspl_w_n19837_0(.douta(w_n19837_0[0]),.doutb(w_n19837_0[1]),.din(n19837));
	jspl jspl_w_n19841_0(.douta(w_n19841_0[0]),.doutb(w_n19841_0[1]),.din(n19841));
	jspl3 jspl3_w_n19843_0(.douta(w_n19843_0[0]),.doutb(w_n19843_0[1]),.doutc(w_n19843_0[2]),.din(n19843));
	jspl jspl_w_n19844_0(.douta(w_n19844_0[0]),.doutb(w_n19844_0[1]),.din(n19844));
	jspl jspl_w_n19848_0(.douta(w_n19848_0[0]),.doutb(w_n19848_0[1]),.din(n19848));
	jspl jspl_w_n19849_0(.douta(w_n19849_0[0]),.doutb(w_n19849_0[1]),.din(n19849));
	jspl3 jspl3_w_n19851_0(.douta(w_n19851_0[0]),.doutb(w_n19851_0[1]),.doutc(w_n19851_0[2]),.din(n19851));
	jspl jspl_w_n19852_0(.douta(w_n19852_0[0]),.doutb(w_n19852_0[1]),.din(n19852));
	jspl jspl_w_n19856_0(.douta(w_n19856_0[0]),.doutb(w_n19856_0[1]),.din(n19856));
	jspl3 jspl3_w_n19858_0(.douta(w_n19858_0[0]),.doutb(w_n19858_0[1]),.doutc(w_n19858_0[2]),.din(n19858));
	jspl jspl_w_n19859_0(.douta(w_n19859_0[0]),.doutb(w_n19859_0[1]),.din(n19859));
	jspl jspl_w_n19863_0(.douta(w_n19863_0[0]),.doutb(w_n19863_0[1]),.din(n19863));
	jspl jspl_w_n19864_0(.douta(w_n19864_0[0]),.doutb(w_n19864_0[1]),.din(n19864));
	jspl3 jspl3_w_n19866_0(.douta(w_n19866_0[0]),.doutb(w_n19866_0[1]),.doutc(w_n19866_0[2]),.din(n19866));
	jspl jspl_w_n19867_0(.douta(w_n19867_0[0]),.doutb(w_n19867_0[1]),.din(n19867));
	jspl jspl_w_n19871_0(.douta(w_n19871_0[0]),.doutb(w_n19871_0[1]),.din(n19871));
	jspl3 jspl3_w_n19873_0(.douta(w_n19873_0[0]),.doutb(w_n19873_0[1]),.doutc(w_n19873_0[2]),.din(n19873));
	jspl jspl_w_n19874_0(.douta(w_n19874_0[0]),.doutb(w_n19874_0[1]),.din(n19874));
	jspl jspl_w_n19878_0(.douta(w_n19878_0[0]),.doutb(w_n19878_0[1]),.din(n19878));
	jspl jspl_w_n19879_0(.douta(w_n19879_0[0]),.doutb(w_n19879_0[1]),.din(n19879));
	jspl3 jspl3_w_n19881_0(.douta(w_n19881_0[0]),.doutb(w_n19881_0[1]),.doutc(w_n19881_0[2]),.din(n19881));
	jspl jspl_w_n19882_0(.douta(w_n19882_0[0]),.doutb(w_n19882_0[1]),.din(n19882));
	jspl jspl_w_n19886_0(.douta(w_n19886_0[0]),.doutb(w_n19886_0[1]),.din(n19886));
	jspl3 jspl3_w_n19888_0(.douta(w_n19888_0[0]),.doutb(w_n19888_0[1]),.doutc(w_n19888_0[2]),.din(n19888));
	jspl jspl_w_n19889_0(.douta(w_n19889_0[0]),.doutb(w_n19889_0[1]),.din(n19889));
	jspl jspl_w_n19893_0(.douta(w_n19893_0[0]),.doutb(w_n19893_0[1]),.din(n19893));
	jspl jspl_w_n19894_0(.douta(w_n19894_0[0]),.doutb(w_n19894_0[1]),.din(n19894));
	jspl3 jspl3_w_n19896_0(.douta(w_n19896_0[0]),.doutb(w_n19896_0[1]),.doutc(w_n19896_0[2]),.din(n19896));
	jspl jspl_w_n19897_0(.douta(w_n19897_0[0]),.doutb(w_n19897_0[1]),.din(n19897));
	jspl jspl_w_n19901_0(.douta(w_n19901_0[0]),.doutb(w_n19901_0[1]),.din(n19901));
	jspl jspl_w_n19902_0(.douta(w_n19902_0[0]),.doutb(w_n19902_0[1]),.din(n19902));
	jspl3 jspl3_w_n19904_0(.douta(w_n19904_0[0]),.doutb(w_n19904_0[1]),.doutc(w_n19904_0[2]),.din(n19904));
	jspl jspl_w_n19905_0(.douta(w_n19905_0[0]),.doutb(w_n19905_0[1]),.din(n19905));
	jspl jspl_w_n19909_0(.douta(w_n19909_0[0]),.doutb(w_n19909_0[1]),.din(n19909));
	jspl3 jspl3_w_n19911_0(.douta(w_n19911_0[0]),.doutb(w_n19911_0[1]),.doutc(w_n19911_0[2]),.din(n19911));
	jspl jspl_w_n19912_0(.douta(w_n19912_0[0]),.doutb(w_n19912_0[1]),.din(n19912));
	jspl jspl_w_n19916_0(.douta(w_n19916_0[0]),.doutb(w_n19916_0[1]),.din(n19916));
	jspl3 jspl3_w_n19918_0(.douta(w_n19918_0[0]),.doutb(w_n19918_0[1]),.doutc(w_n19918_0[2]),.din(n19918));
	jspl jspl_w_n19919_0(.douta(w_n19919_0[0]),.doutb(w_n19919_0[1]),.din(n19919));
	jspl jspl_w_n19923_0(.douta(w_n19923_0[0]),.doutb(w_n19923_0[1]),.din(n19923));
	jspl jspl_w_n19924_0(.douta(w_n19924_0[0]),.doutb(w_n19924_0[1]),.din(n19924));
	jspl3 jspl3_w_n19926_0(.douta(w_n19926_0[0]),.doutb(w_n19926_0[1]),.doutc(w_n19926_0[2]),.din(n19926));
	jspl jspl_w_n19927_0(.douta(w_n19927_0[0]),.doutb(w_n19927_0[1]),.din(n19927));
	jspl jspl_w_n19931_0(.douta(w_n19931_0[0]),.doutb(w_n19931_0[1]),.din(n19931));
	jspl3 jspl3_w_n19933_0(.douta(w_n19933_0[0]),.doutb(w_n19933_0[1]),.doutc(w_n19933_0[2]),.din(n19933));
	jspl jspl_w_n19934_0(.douta(w_n19934_0[0]),.doutb(w_n19934_0[1]),.din(n19934));
	jspl jspl_w_n19938_0(.douta(w_n19938_0[0]),.doutb(w_n19938_0[1]),.din(n19938));
	jspl jspl_w_n19939_0(.douta(w_n19939_0[0]),.doutb(w_n19939_0[1]),.din(n19939));
	jspl3 jspl3_w_n19941_0(.douta(w_n19941_0[0]),.doutb(w_n19941_0[1]),.doutc(w_n19941_0[2]),.din(n19941));
	jspl jspl_w_n19942_0(.douta(w_n19942_0[0]),.doutb(w_n19942_0[1]),.din(n19942));
	jspl jspl_w_n19946_0(.douta(w_n19946_0[0]),.doutb(w_n19946_0[1]),.din(n19946));
	jspl3 jspl3_w_n19948_0(.douta(w_n19948_0[0]),.doutb(w_n19948_0[1]),.doutc(w_n19948_0[2]),.din(n19948));
	jspl jspl_w_n19949_0(.douta(w_n19949_0[0]),.doutb(w_n19949_0[1]),.din(n19949));
	jspl jspl_w_n19953_0(.douta(w_n19953_0[0]),.doutb(w_n19953_0[1]),.din(n19953));
	jspl jspl_w_n19954_0(.douta(w_n19954_0[0]),.doutb(w_n19954_0[1]),.din(n19954));
	jspl3 jspl3_w_n19956_0(.douta(w_n19956_0[0]),.doutb(w_n19956_0[1]),.doutc(w_n19956_0[2]),.din(n19956));
	jspl jspl_w_n19957_0(.douta(w_n19957_0[0]),.doutb(w_n19957_0[1]),.din(n19957));
	jspl jspl_w_n19961_0(.douta(w_n19961_0[0]),.doutb(w_n19961_0[1]),.din(n19961));
	jspl jspl_w_n19962_0(.douta(w_n19962_0[0]),.doutb(w_n19962_0[1]),.din(n19962));
	jspl3 jspl3_w_n19964_0(.douta(w_n19964_0[0]),.doutb(w_n19964_0[1]),.doutc(w_n19964_0[2]),.din(n19964));
	jspl jspl_w_n19965_0(.douta(w_n19965_0[0]),.doutb(w_n19965_0[1]),.din(n19965));
	jspl jspl_w_n19969_0(.douta(w_n19969_0[0]),.doutb(w_n19969_0[1]),.din(n19969));
	jspl jspl_w_n19970_0(.douta(w_n19970_0[0]),.doutb(w_n19970_0[1]),.din(n19970));
	jspl3 jspl3_w_n19972_0(.douta(w_n19972_0[0]),.doutb(w_n19972_0[1]),.doutc(w_n19972_0[2]),.din(n19972));
	jspl jspl_w_n19973_0(.douta(w_n19973_0[0]),.doutb(w_n19973_0[1]),.din(n19973));
	jspl jspl_w_n19977_0(.douta(w_n19977_0[0]),.doutb(w_n19977_0[1]),.din(n19977));
	jspl3 jspl3_w_n19979_0(.douta(w_n19979_0[0]),.doutb(w_n19979_0[1]),.doutc(w_n19979_0[2]),.din(n19979));
	jspl jspl_w_n19980_0(.douta(w_n19980_0[0]),.doutb(w_n19980_0[1]),.din(n19980));
	jspl jspl_w_n19984_0(.douta(w_n19984_0[0]),.doutb(w_n19984_0[1]),.din(n19984));
	jspl jspl_w_n19985_0(.douta(w_n19985_0[0]),.doutb(w_n19985_0[1]),.din(n19985));
	jspl3 jspl3_w_n19987_0(.douta(w_n19987_0[0]),.doutb(w_n19987_0[1]),.doutc(w_n19987_0[2]),.din(n19987));
	jspl jspl_w_n19988_0(.douta(w_n19988_0[0]),.doutb(w_n19988_0[1]),.din(n19988));
	jspl jspl_w_n19992_0(.douta(w_n19992_0[0]),.doutb(w_n19992_0[1]),.din(n19992));
	jspl3 jspl3_w_n19994_0(.douta(w_n19994_0[0]),.doutb(w_n19994_0[1]),.doutc(w_n19994_0[2]),.din(n19994));
	jspl jspl_w_n19995_0(.douta(w_n19995_0[0]),.doutb(w_n19995_0[1]),.din(n19995));
	jspl jspl_w_n19999_0(.douta(w_n19999_0[0]),.doutb(w_n19999_0[1]),.din(n19999));
	jspl jspl_w_n20000_0(.douta(w_n20000_0[0]),.doutb(w_n20000_0[1]),.din(n20000));
	jspl3 jspl3_w_n20002_0(.douta(w_n20002_0[0]),.doutb(w_n20002_0[1]),.doutc(w_n20002_0[2]),.din(n20002));
	jspl jspl_w_n20003_0(.douta(w_n20003_0[0]),.doutb(w_n20003_0[1]),.din(n20003));
	jspl jspl_w_n20007_0(.douta(w_n20007_0[0]),.doutb(w_n20007_0[1]),.din(n20007));
	jspl3 jspl3_w_n20009_0(.douta(w_n20009_0[0]),.doutb(w_n20009_0[1]),.doutc(w_n20009_0[2]),.din(n20009));
	jspl jspl_w_n20010_0(.douta(w_n20010_0[0]),.doutb(w_n20010_0[1]),.din(n20010));
	jspl jspl_w_n20014_0(.douta(w_n20014_0[0]),.doutb(w_n20014_0[1]),.din(n20014));
	jspl jspl_w_n20015_0(.douta(w_n20015_0[0]),.doutb(w_n20015_0[1]),.din(n20015));
	jspl3 jspl3_w_n20017_0(.douta(w_n20017_0[0]),.doutb(w_n20017_0[1]),.doutc(w_n20017_0[2]),.din(n20017));
	jspl jspl_w_n20018_0(.douta(w_n20018_0[0]),.doutb(w_n20018_0[1]),.din(n20018));
	jspl jspl_w_n20022_0(.douta(w_n20022_0[0]),.doutb(w_n20022_0[1]),.din(n20022));
	jspl3 jspl3_w_n20024_0(.douta(w_n20024_0[0]),.doutb(w_n20024_0[1]),.doutc(w_n20024_0[2]),.din(n20024));
	jspl jspl_w_n20025_0(.douta(w_n20025_0[0]),.doutb(w_n20025_0[1]),.din(n20025));
	jspl jspl_w_n20029_0(.douta(w_n20029_0[0]),.doutb(w_n20029_0[1]),.din(n20029));
	jspl jspl_w_n20030_0(.douta(w_n20030_0[0]),.doutb(w_n20030_0[1]),.din(n20030));
	jspl3 jspl3_w_n20032_0(.douta(w_n20032_0[0]),.doutb(w_n20032_0[1]),.doutc(w_n20032_0[2]),.din(n20032));
	jspl jspl_w_n20033_0(.douta(w_n20033_0[0]),.doutb(w_n20033_0[1]),.din(n20033));
	jspl jspl_w_n20037_0(.douta(w_n20037_0[0]),.doutb(w_n20037_0[1]),.din(n20037));
	jspl jspl_w_n20038_0(.douta(w_n20038_0[0]),.doutb(w_n20038_0[1]),.din(n20038));
	jspl3 jspl3_w_n20040_0(.douta(w_n20040_0[0]),.doutb(w_n20040_0[1]),.doutc(w_n20040_0[2]),.din(n20040));
	jspl jspl_w_n20041_0(.douta(w_n20041_0[0]),.doutb(w_n20041_0[1]),.din(n20041));
	jspl jspl_w_n20045_0(.douta(w_n20045_0[0]),.doutb(w_n20045_0[1]),.din(n20045));
	jspl jspl_w_n20046_0(.douta(w_n20046_0[0]),.doutb(w_n20046_0[1]),.din(n20046));
	jspl3 jspl3_w_n20048_0(.douta(w_n20048_0[0]),.doutb(w_n20048_0[1]),.doutc(w_n20048_0[2]),.din(n20048));
	jspl jspl_w_n20049_0(.douta(w_n20049_0[0]),.doutb(w_n20049_0[1]),.din(n20049));
	jspl jspl_w_n20053_0(.douta(w_n20053_0[0]),.doutb(w_n20053_0[1]),.din(n20053));
	jspl3 jspl3_w_n20055_0(.douta(w_n20055_0[0]),.doutb(w_n20055_0[1]),.doutc(w_n20055_0[2]),.din(n20055));
	jspl jspl_w_n20056_0(.douta(w_n20056_0[0]),.doutb(w_n20056_0[1]),.din(n20056));
	jspl jspl_w_n20060_0(.douta(w_n20060_0[0]),.doutb(w_n20060_0[1]),.din(n20060));
	jspl jspl_w_n20061_0(.douta(w_n20061_0[0]),.doutb(w_n20061_0[1]),.din(n20061));
	jspl3 jspl3_w_n20063_0(.douta(w_n20063_0[0]),.doutb(w_n20063_0[1]),.doutc(w_n20063_0[2]),.din(n20063));
	jspl jspl_w_n20064_0(.douta(w_n20064_0[0]),.doutb(w_n20064_0[1]),.din(n20064));
	jspl jspl_w_n20068_0(.douta(w_n20068_0[0]),.doutb(w_n20068_0[1]),.din(n20068));
	jspl jspl_w_n20069_0(.douta(w_n20069_0[0]),.doutb(w_n20069_0[1]),.din(n20069));
	jspl3 jspl3_w_n20071_0(.douta(w_n20071_0[0]),.doutb(w_n20071_0[1]),.doutc(w_n20071_0[2]),.din(n20071));
	jspl jspl_w_n20072_0(.douta(w_n20072_0[0]),.doutb(w_n20072_0[1]),.din(n20072));
	jspl jspl_w_n20076_0(.douta(w_n20076_0[0]),.doutb(w_n20076_0[1]),.din(n20076));
	jspl jspl_w_n20077_0(.douta(w_n20077_0[0]),.doutb(w_n20077_0[1]),.din(n20077));
	jspl3 jspl3_w_n20079_0(.douta(w_n20079_0[0]),.doutb(w_n20079_0[1]),.doutc(w_n20079_0[2]),.din(n20079));
	jspl jspl_w_n20080_0(.douta(w_n20080_0[0]),.doutb(w_n20080_0[1]),.din(n20080));
	jspl jspl_w_n20084_0(.douta(w_n20084_0[0]),.doutb(w_n20084_0[1]),.din(n20084));
	jspl jspl_w_n20085_0(.douta(w_n20085_0[0]),.doutb(w_n20085_0[1]),.din(n20085));
	jspl3 jspl3_w_n20087_0(.douta(w_n20087_0[0]),.doutb(w_n20087_0[1]),.doutc(w_n20087_0[2]),.din(n20087));
	jspl jspl_w_n20088_0(.douta(w_n20088_0[0]),.doutb(w_n20088_0[1]),.din(n20088));
	jspl jspl_w_n20092_0(.douta(w_n20092_0[0]),.doutb(w_n20092_0[1]),.din(n20092));
	jspl jspl_w_n20093_0(.douta(w_n20093_0[0]),.doutb(w_n20093_0[1]),.din(n20093));
	jspl3 jspl3_w_n20095_0(.douta(w_n20095_0[0]),.doutb(w_n20095_0[1]),.doutc(w_n20095_0[2]),.din(n20095));
	jspl jspl_w_n20096_0(.douta(w_n20096_0[0]),.doutb(w_n20096_0[1]),.din(n20096));
	jspl jspl_w_n20100_0(.douta(w_n20100_0[0]),.doutb(w_n20100_0[1]),.din(n20100));
	jspl3 jspl3_w_n20102_0(.douta(w_n20102_0[0]),.doutb(w_n20102_0[1]),.doutc(w_n20102_0[2]),.din(n20102));
	jspl jspl_w_n20103_0(.douta(w_n20103_0[0]),.doutb(w_n20103_0[1]),.din(n20103));
	jspl jspl_w_n20107_0(.douta(w_n20107_0[0]),.doutb(w_n20107_0[1]),.din(n20107));
	jspl jspl_w_n20108_0(.douta(w_n20108_0[0]),.doutb(w_n20108_0[1]),.din(n20108));
	jspl3 jspl3_w_n20110_0(.douta(w_n20110_0[0]),.doutb(w_n20110_0[1]),.doutc(w_n20110_0[2]),.din(n20110));
	jspl jspl_w_n20111_0(.douta(w_n20111_0[0]),.doutb(w_n20111_0[1]),.din(n20111));
	jspl jspl_w_n20115_0(.douta(w_n20115_0[0]),.doutb(w_n20115_0[1]),.din(n20115));
	jspl3 jspl3_w_n20117_0(.douta(w_n20117_0[0]),.doutb(w_n20117_0[1]),.doutc(w_n20117_0[2]),.din(n20117));
	jspl jspl_w_n20118_0(.douta(w_n20118_0[0]),.doutb(w_n20118_0[1]),.din(n20118));
	jspl jspl_w_n20122_0(.douta(w_n20122_0[0]),.doutb(w_n20122_0[1]),.din(n20122));
	jspl jspl_w_n20123_0(.douta(w_n20123_0[0]),.doutb(w_n20123_0[1]),.din(n20123));
	jspl3 jspl3_w_n20125_0(.douta(w_n20125_0[0]),.doutb(w_n20125_0[1]),.doutc(w_n20125_0[2]),.din(n20125));
	jspl jspl_w_n20126_0(.douta(w_n20126_0[0]),.doutb(w_n20126_0[1]),.din(n20126));
	jspl jspl_w_n20130_0(.douta(w_n20130_0[0]),.doutb(w_n20130_0[1]),.din(n20130));
	jspl jspl_w_n20131_0(.douta(w_n20131_0[0]),.doutb(w_n20131_0[1]),.din(n20131));
	jspl3 jspl3_w_n20133_0(.douta(w_n20133_0[0]),.doutb(w_n20133_0[1]),.doutc(w_n20133_0[2]),.din(n20133));
	jspl jspl_w_n20134_0(.douta(w_n20134_0[0]),.doutb(w_n20134_0[1]),.din(n20134));
	jspl jspl_w_n20138_0(.douta(w_n20138_0[0]),.doutb(w_n20138_0[1]),.din(n20138));
	jspl3 jspl3_w_n20140_0(.douta(w_n20140_0[0]),.doutb(w_n20140_0[1]),.doutc(w_n20140_0[2]),.din(n20140));
	jspl jspl_w_n20141_0(.douta(w_n20141_0[0]),.doutb(w_n20141_0[1]),.din(n20141));
	jspl jspl_w_n20144_0(.douta(w_n20144_0[0]),.doutb(w_n20144_0[1]),.din(n20144));
	jspl3 jspl3_w_n20147_0(.douta(w_n20147_0[0]),.doutb(w_n20147_0[1]),.doutc(w_n20147_0[2]),.din(n20147));
	jspl jspl_w_n20148_0(.douta(w_n20148_0[0]),.doutb(w_n20148_0[1]),.din(n20148));
	jspl jspl_w_n20152_0(.douta(w_n20152_0[0]),.doutb(w_n20152_0[1]),.din(n20152));
	jspl jspl_w_n20153_0(.douta(w_n20153_0[0]),.doutb(w_n20153_0[1]),.din(n20153));
	jspl3 jspl3_w_n20155_0(.douta(w_n20155_0[0]),.doutb(w_n20155_0[1]),.doutc(w_n20155_0[2]),.din(n20155));
	jspl jspl_w_n20156_0(.douta(w_n20156_0[0]),.doutb(w_n20156_0[1]),.din(n20156));
	jspl jspl_w_n20160_0(.douta(w_n20160_0[0]),.doutb(w_n20160_0[1]),.din(n20160));
	jspl3 jspl3_w_n20162_0(.douta(w_n20162_0[0]),.doutb(w_n20162_0[1]),.doutc(w_n20162_0[2]),.din(n20162));
	jspl jspl_w_n20163_0(.douta(w_n20163_0[0]),.doutb(w_n20163_0[1]),.din(n20163));
	jspl jspl_w_n20167_0(.douta(w_n20167_0[0]),.doutb(w_n20167_0[1]),.din(n20167));
	jspl jspl_w_n20168_0(.douta(w_n20168_0[0]),.doutb(w_n20168_0[1]),.din(n20168));
	jspl3 jspl3_w_n20170_0(.douta(w_n20170_0[0]),.doutb(w_n20170_0[1]),.doutc(w_n20170_0[2]),.din(n20170));
	jspl jspl_w_n20171_0(.douta(w_n20171_0[0]),.doutb(w_n20171_0[1]),.din(n20171));
	jspl jspl_w_n20175_0(.douta(w_n20175_0[0]),.doutb(w_n20175_0[1]),.din(n20175));
	jspl jspl_w_n20176_0(.douta(w_n20176_0[0]),.doutb(w_n20176_0[1]),.din(n20176));
	jspl3 jspl3_w_n20178_0(.douta(w_n20178_0[0]),.doutb(w_n20178_0[1]),.doutc(w_n20178_0[2]),.din(n20178));
	jspl jspl_w_n20179_0(.douta(w_n20179_0[0]),.doutb(w_n20179_0[1]),.din(n20179));
	jspl jspl_w_n20183_0(.douta(w_n20183_0[0]),.doutb(w_n20183_0[1]),.din(n20183));
	jspl3 jspl3_w_n20185_0(.douta(w_n20185_0[0]),.doutb(w_n20185_0[1]),.doutc(w_n20185_0[2]),.din(n20185));
	jspl jspl_w_n20186_0(.douta(w_n20186_0[0]),.doutb(w_n20186_0[1]),.din(n20186));
	jspl jspl_w_n20190_0(.douta(w_n20190_0[0]),.doutb(w_n20190_0[1]),.din(n20190));
	jspl jspl_w_n20191_0(.douta(w_n20191_0[0]),.doutb(w_n20191_0[1]),.din(n20191));
	jspl3 jspl3_w_n20193_0(.douta(w_n20193_0[0]),.doutb(w_n20193_0[1]),.doutc(w_n20193_0[2]),.din(n20193));
	jspl jspl_w_n20194_0(.douta(w_n20194_0[0]),.doutb(w_n20194_0[1]),.din(n20194));
	jspl jspl_w_n20203_0(.douta(w_n20203_0[0]),.doutb(w_n20203_0[1]),.din(n20203));
	jspl jspl_w_n20256_0(.douta(w_n20256_0[0]),.doutb(w_n20256_0[1]),.din(n20256));
	jspl jspl_w_n20269_0(.douta(w_n20269_0[0]),.doutb(w_n20269_0[1]),.din(n20269));
	jspl jspl_w_n20276_0(.douta(w_n20276_0[0]),.doutb(w_n20276_0[1]),.din(n20276));
	jspl jspl_w_n20283_0(.douta(w_n20283_0[0]),.doutb(w_n20283_0[1]),.din(n20283));
	jspl jspl_w_n20290_0(.douta(w_n20290_0[0]),.doutb(w_n20290_0[1]),.din(n20290));
	jspl jspl_w_n20297_0(.douta(w_n20297_0[0]),.doutb(w_n20297_0[1]),.din(n20297));
	jspl jspl_w_n20307_0(.douta(w_n20307_0[0]),.doutb(w_n20307_0[1]),.din(n20307));
	jspl jspl_w_n20311_0(.douta(w_n20311_0[0]),.doutb(w_n20311_0[1]),.din(n20311));
	jspl jspl_w_n20318_0(.douta(w_n20318_0[0]),.doutb(w_n20318_0[1]),.din(n20318));
	jspl jspl_w_n20325_0(.douta(w_n20325_0[0]),.doutb(w_n20325_0[1]),.din(n20325));
	jspl jspl_w_n20338_0(.douta(w_n20338_0[0]),.doutb(w_n20338_0[1]),.din(n20338));
	jspl jspl_w_n20345_0(.douta(w_n20345_0[0]),.doutb(w_n20345_0[1]),.din(n20345));
	jspl jspl_w_n20352_0(.douta(w_n20352_0[0]),.doutb(w_n20352_0[1]),.din(n20352));
	jspl jspl_w_n20359_0(.douta(w_n20359_0[0]),.doutb(w_n20359_0[1]),.din(n20359));
	jspl jspl_w_n20372_0(.douta(w_n20372_0[0]),.doutb(w_n20372_0[1]),.din(n20372));
	jspl jspl_w_n20391_0(.douta(w_n20391_0[0]),.doutb(w_n20391_0[1]),.din(n20391));
	jspl jspl_w_n20398_0(.douta(w_n20398_0[0]),.doutb(w_n20398_0[1]),.din(n20398));
	jspl jspl_w_n20408_0(.douta(w_n20408_0[0]),.doutb(w_n20408_0[1]),.din(n20408));
	jspl jspl_w_n20418_0(.douta(w_n20418_0[0]),.doutb(w_n20418_0[1]),.din(n20418));
	jspl jspl_w_n20428_0(.douta(w_n20428_0[0]),.doutb(w_n20428_0[1]),.din(n20428));
	jspl3 jspl3_w_n20437_0(.douta(w_n20437_0[0]),.doutb(w_n20437_0[1]),.doutc(w_n20437_0[2]),.din(n20437));
	jspl3 jspl3_w_n20439_0(.douta(w_n20439_0[0]),.doutb(w_n20439_0[1]),.doutc(w_n20439_0[2]),.din(n20439));
	jspl jspl_w_n20440_0(.douta(w_n20440_0[0]),.doutb(w_n20440_0[1]),.din(n20440));
	jspl jspl_w_n20442_0(.douta(w_n20442_0[0]),.doutb(w_n20442_0[1]),.din(n20442));
	jspl jspl_w_n20444_0(.douta(w_n20444_0[0]),.doutb(w_n20444_0[1]),.din(n20444));
	jspl jspl_w_n20445_0(.douta(w_n20445_0[0]),.doutb(w_n20445_0[1]),.din(n20445));
	jspl3 jspl3_w_n20446_0(.douta(w_n20446_0[0]),.doutb(w_n20446_0[1]),.doutc(w_n20446_0[2]),.din(n20446));
	jspl jspl_w_n20451_0(.douta(w_n20451_0[0]),.doutb(w_n20451_0[1]),.din(n20451));
	jspl jspl_w_n20452_0(.douta(w_n20452_0[0]),.doutb(w_n20452_0[1]),.din(n20452));
	jspl jspl_w_n20458_0(.douta(w_n20458_0[0]),.doutb(w_n20458_0[1]),.din(n20458));
	jspl jspl_w_n20459_0(.douta(w_n20459_0[0]),.doutb(w_n20459_0[1]),.din(n20459));
	jspl jspl_w_n20464_0(.douta(w_n20464_0[0]),.doutb(w_n20464_0[1]),.din(n20464));
	jspl3 jspl3_w_n20468_0(.douta(w_n20468_0[0]),.doutb(w_n20468_0[1]),.doutc(w_n20468_0[2]),.din(n20468));
	jspl3 jspl3_w_n20468_1(.douta(w_n20468_1[0]),.doutb(w_n20468_1[1]),.doutc(w_n20468_1[2]),.din(w_n20468_0[0]));
	jspl3 jspl3_w_n20468_2(.douta(w_n20468_2[0]),.doutb(w_n20468_2[1]),.doutc(w_n20468_2[2]),.din(w_n20468_0[1]));
	jspl3 jspl3_w_n20468_3(.douta(w_n20468_3[0]),.doutb(w_n20468_3[1]),.doutc(w_n20468_3[2]),.din(w_n20468_0[2]));
	jspl3 jspl3_w_n20468_4(.douta(w_n20468_4[0]),.doutb(w_n20468_4[1]),.doutc(w_n20468_4[2]),.din(w_n20468_1[0]));
	jspl3 jspl3_w_n20468_5(.douta(w_n20468_5[0]),.doutb(w_n20468_5[1]),.doutc(w_n20468_5[2]),.din(w_n20468_1[1]));
	jspl3 jspl3_w_n20468_6(.douta(w_n20468_6[0]),.doutb(w_n20468_6[1]),.doutc(w_n20468_6[2]),.din(w_n20468_1[2]));
	jspl3 jspl3_w_n20468_7(.douta(w_n20468_7[0]),.doutb(w_n20468_7[1]),.doutc(w_n20468_7[2]),.din(w_n20468_2[0]));
	jspl3 jspl3_w_n20468_8(.douta(w_n20468_8[0]),.doutb(w_n20468_8[1]),.doutc(w_n20468_8[2]),.din(w_n20468_2[1]));
	jspl3 jspl3_w_n20468_9(.douta(w_n20468_9[0]),.doutb(w_n20468_9[1]),.doutc(w_n20468_9[2]),.din(w_n20468_2[2]));
	jspl3 jspl3_w_n20468_10(.douta(w_n20468_10[0]),.doutb(w_n20468_10[1]),.doutc(w_n20468_10[2]),.din(w_n20468_3[0]));
	jspl3 jspl3_w_n20468_11(.douta(w_n20468_11[0]),.doutb(w_n20468_11[1]),.doutc(w_n20468_11[2]),.din(w_n20468_3[1]));
	jspl3 jspl3_w_n20468_12(.douta(w_n20468_12[0]),.doutb(w_n20468_12[1]),.doutc(w_n20468_12[2]),.din(w_n20468_3[2]));
	jspl3 jspl3_w_n20468_13(.douta(w_n20468_13[0]),.doutb(w_n20468_13[1]),.doutc(w_n20468_13[2]),.din(w_n20468_4[0]));
	jspl3 jspl3_w_n20468_14(.douta(w_n20468_14[0]),.doutb(w_n20468_14[1]),.doutc(w_n20468_14[2]),.din(w_n20468_4[1]));
	jspl3 jspl3_w_n20468_15(.douta(w_n20468_15[0]),.doutb(w_n20468_15[1]),.doutc(w_n20468_15[2]),.din(w_n20468_4[2]));
	jspl3 jspl3_w_n20468_16(.douta(w_n20468_16[0]),.doutb(w_n20468_16[1]),.doutc(w_n20468_16[2]),.din(w_n20468_5[0]));
	jspl3 jspl3_w_n20468_17(.douta(w_n20468_17[0]),.doutb(w_n20468_17[1]),.doutc(w_n20468_17[2]),.din(w_n20468_5[1]));
	jspl3 jspl3_w_n20468_18(.douta(w_n20468_18[0]),.doutb(w_n20468_18[1]),.doutc(w_n20468_18[2]),.din(w_n20468_5[2]));
	jspl3 jspl3_w_n20468_19(.douta(w_n20468_19[0]),.doutb(w_n20468_19[1]),.doutc(w_n20468_19[2]),.din(w_n20468_6[0]));
	jspl3 jspl3_w_n20468_20(.douta(w_n20468_20[0]),.doutb(w_n20468_20[1]),.doutc(w_n20468_20[2]),.din(w_n20468_6[1]));
	jspl3 jspl3_w_n20468_21(.douta(w_n20468_21[0]),.doutb(w_n20468_21[1]),.doutc(w_n20468_21[2]),.din(w_n20468_6[2]));
	jspl3 jspl3_w_n20468_22(.douta(w_n20468_22[0]),.doutb(w_n20468_22[1]),.doutc(w_n20468_22[2]),.din(w_n20468_7[0]));
	jspl3 jspl3_w_n20468_23(.douta(w_n20468_23[0]),.doutb(w_n20468_23[1]),.doutc(w_n20468_23[2]),.din(w_n20468_7[1]));
	jspl3 jspl3_w_n20468_24(.douta(w_n20468_24[0]),.doutb(w_n20468_24[1]),.doutc(w_n20468_24[2]),.din(w_n20468_7[2]));
	jspl3 jspl3_w_n20468_25(.douta(w_n20468_25[0]),.doutb(w_n20468_25[1]),.doutc(w_n20468_25[2]),.din(w_n20468_8[0]));
	jspl3 jspl3_w_n20468_26(.douta(w_n20468_26[0]),.doutb(w_n20468_26[1]),.doutc(w_n20468_26[2]),.din(w_n20468_8[1]));
	jspl3 jspl3_w_n20468_27(.douta(w_n20468_27[0]),.doutb(w_n20468_27[1]),.doutc(w_n20468_27[2]),.din(w_n20468_8[2]));
	jspl3 jspl3_w_n20468_28(.douta(w_n20468_28[0]),.doutb(w_n20468_28[1]),.doutc(w_n20468_28[2]),.din(w_n20468_9[0]));
	jspl3 jspl3_w_n20468_29(.douta(w_n20468_29[0]),.doutb(w_n20468_29[1]),.doutc(w_n20468_29[2]),.din(w_n20468_9[1]));
	jspl3 jspl3_w_n20468_30(.douta(w_n20468_30[0]),.doutb(w_n20468_30[1]),.doutc(w_n20468_30[2]),.din(w_n20468_9[2]));
	jspl3 jspl3_w_n20468_31(.douta(w_n20468_31[0]),.doutb(w_n20468_31[1]),.doutc(w_n20468_31[2]),.din(w_n20468_10[0]));
	jspl3 jspl3_w_n20468_32(.douta(w_n20468_32[0]),.doutb(w_n20468_32[1]),.doutc(w_n20468_32[2]),.din(w_n20468_10[1]));
	jspl3 jspl3_w_n20468_33(.douta(w_n20468_33[0]),.doutb(w_n20468_33[1]),.doutc(w_n20468_33[2]),.din(w_n20468_10[2]));
	jspl3 jspl3_w_n20468_34(.douta(w_n20468_34[0]),.doutb(w_n20468_34[1]),.doutc(w_n20468_34[2]),.din(w_n20468_11[0]));
	jspl3 jspl3_w_n20468_35(.douta(w_n20468_35[0]),.doutb(w_n20468_35[1]),.doutc(w_n20468_35[2]),.din(w_n20468_11[1]));
	jspl3 jspl3_w_n20471_0(.douta(w_n20471_0[0]),.doutb(w_n20471_0[1]),.doutc(w_n20471_0[2]),.din(n20471));
	jspl jspl_w_n20472_0(.douta(w_n20472_0[0]),.doutb(w_n20472_0[1]),.din(n20472));
	jspl3 jspl3_w_n20473_0(.douta(w_n20473_0[0]),.doutb(w_n20473_0[1]),.doutc(w_n20473_0[2]),.din(n20473));
	jspl3 jspl3_w_n20473_1(.douta(w_n20473_1[0]),.doutb(w_n20473_1[1]),.doutc(w_n20473_1[2]),.din(w_n20473_0[0]));
	jspl jspl_w_n20474_0(.douta(w_n20474_0[0]),.doutb(w_n20474_0[1]),.din(n20474));
	jspl3 jspl3_w_n20475_0(.douta(w_n20475_0[0]),.doutb(w_n20475_0[1]),.doutc(w_n20475_0[2]),.din(n20475));
	jspl jspl_w_n20476_0(.douta(w_n20476_0[0]),.doutb(w_n20476_0[1]),.din(n20476));
	jspl3 jspl3_w_n20479_0(.douta(w_n20479_0[0]),.doutb(w_n20479_0[1]),.doutc(w_n20479_0[2]),.din(n20479));
	jspl jspl_w_n20480_0(.douta(w_n20480_0[0]),.doutb(w_n20480_0[1]),.din(n20480));
	jspl3 jspl3_w_n20487_0(.douta(w_n20487_0[0]),.doutb(w_n20487_0[1]),.doutc(w_n20487_0[2]),.din(n20487));
	jspl jspl_w_n20488_0(.douta(w_n20488_0[0]),.doutb(w_n20488_0[1]),.din(n20488));
	jspl jspl_w_n20491_0(.douta(w_n20491_0[0]),.doutb(w_n20491_0[1]),.din(n20491));
	jspl3 jspl3_w_n20496_0(.douta(w_n20496_0[0]),.doutb(w_n20496_0[1]),.doutc(w_n20496_0[2]),.din(n20496));
	jspl3 jspl3_w_n20498_0(.douta(w_n20498_0[0]),.doutb(w_n20498_0[1]),.doutc(w_n20498_0[2]),.din(n20498));
	jspl jspl_w_n20499_0(.douta(w_n20499_0[0]),.doutb(w_n20499_0[1]),.din(n20499));
	jspl3 jspl3_w_n20503_0(.douta(w_n20503_0[0]),.doutb(w_n20503_0[1]),.doutc(w_n20503_0[2]),.din(n20503));
	jspl3 jspl3_w_n20506_0(.douta(w_n20506_0[0]),.doutb(w_n20506_0[1]),.doutc(w_n20506_0[2]),.din(n20506));
	jspl jspl_w_n20507_0(.douta(w_n20507_0[0]),.doutb(w_n20507_0[1]),.din(n20507));
	jspl3 jspl3_w_n20511_0(.douta(w_n20511_0[0]),.doutb(w_n20511_0[1]),.doutc(w_n20511_0[2]),.din(n20511));
	jspl3 jspl3_w_n20513_0(.douta(w_n20513_0[0]),.doutb(w_n20513_0[1]),.doutc(w_n20513_0[2]),.din(n20513));
	jspl jspl_w_n20514_0(.douta(w_n20514_0[0]),.doutb(w_n20514_0[1]),.din(n20514));
	jspl3 jspl3_w_n20518_0(.douta(w_n20518_0[0]),.doutb(w_n20518_0[1]),.doutc(w_n20518_0[2]),.din(n20518));
	jspl3 jspl3_w_n20520_0(.douta(w_n20520_0[0]),.doutb(w_n20520_0[1]),.doutc(w_n20520_0[2]),.din(n20520));
	jspl jspl_w_n20521_0(.douta(w_n20521_0[0]),.doutb(w_n20521_0[1]),.din(n20521));
	jspl3 jspl3_w_n20525_0(.douta(w_n20525_0[0]),.doutb(w_n20525_0[1]),.doutc(w_n20525_0[2]),.din(n20525));
	jspl3 jspl3_w_n20527_0(.douta(w_n20527_0[0]),.doutb(w_n20527_0[1]),.doutc(w_n20527_0[2]),.din(n20527));
	jspl jspl_w_n20528_0(.douta(w_n20528_0[0]),.doutb(w_n20528_0[1]),.din(n20528));
	jspl3 jspl3_w_n20532_0(.douta(w_n20532_0[0]),.doutb(w_n20532_0[1]),.doutc(w_n20532_0[2]),.din(n20532));
	jspl3 jspl3_w_n20535_0(.douta(w_n20535_0[0]),.doutb(w_n20535_0[1]),.doutc(w_n20535_0[2]),.din(n20535));
	jspl jspl_w_n20536_0(.douta(w_n20536_0[0]),.doutb(w_n20536_0[1]),.din(n20536));
	jspl3 jspl3_w_n20540_0(.douta(w_n20540_0[0]),.doutb(w_n20540_0[1]),.doutc(w_n20540_0[2]),.din(n20540));
	jspl3 jspl3_w_n20542_0(.douta(w_n20542_0[0]),.doutb(w_n20542_0[1]),.doutc(w_n20542_0[2]),.din(n20542));
	jspl jspl_w_n20543_0(.douta(w_n20543_0[0]),.doutb(w_n20543_0[1]),.din(n20543));
	jspl jspl_w_n20547_0(.douta(w_n20547_0[0]),.doutb(w_n20547_0[1]),.din(n20547));
	jspl jspl_w_n20548_0(.douta(w_n20548_0[0]),.doutb(w_n20548_0[1]),.din(n20548));
	jspl3 jspl3_w_n20550_0(.douta(w_n20550_0[0]),.doutb(w_n20550_0[1]),.doutc(w_n20550_0[2]),.din(n20550));
	jspl jspl_w_n20551_0(.douta(w_n20551_0[0]),.doutb(w_n20551_0[1]),.din(n20551));
	jspl3 jspl3_w_n20555_0(.douta(w_n20555_0[0]),.doutb(w_n20555_0[1]),.doutc(w_n20555_0[2]),.din(n20555));
	jspl3 jspl3_w_n20557_0(.douta(w_n20557_0[0]),.doutb(w_n20557_0[1]),.doutc(w_n20557_0[2]),.din(n20557));
	jspl jspl_w_n20558_0(.douta(w_n20558_0[0]),.doutb(w_n20558_0[1]),.din(n20558));
	jspl3 jspl3_w_n20562_0(.douta(w_n20562_0[0]),.doutb(w_n20562_0[1]),.doutc(w_n20562_0[2]),.din(n20562));
	jspl3 jspl3_w_n20565_0(.douta(w_n20565_0[0]),.doutb(w_n20565_0[1]),.doutc(w_n20565_0[2]),.din(n20565));
	jspl jspl_w_n20566_0(.douta(w_n20566_0[0]),.doutb(w_n20566_0[1]),.din(n20566));
	jspl3 jspl3_w_n20570_0(.douta(w_n20570_0[0]),.doutb(w_n20570_0[1]),.doutc(w_n20570_0[2]),.din(n20570));
	jspl3 jspl3_w_n20572_0(.douta(w_n20572_0[0]),.doutb(w_n20572_0[1]),.doutc(w_n20572_0[2]),.din(n20572));
	jspl jspl_w_n20573_0(.douta(w_n20573_0[0]),.doutb(w_n20573_0[1]),.din(n20573));
	jspl3 jspl3_w_n20577_0(.douta(w_n20577_0[0]),.doutb(w_n20577_0[1]),.doutc(w_n20577_0[2]),.din(n20577));
	jspl3 jspl3_w_n20580_0(.douta(w_n20580_0[0]),.doutb(w_n20580_0[1]),.doutc(w_n20580_0[2]),.din(n20580));
	jspl jspl_w_n20581_0(.douta(w_n20581_0[0]),.doutb(w_n20581_0[1]),.din(n20581));
	jspl3 jspl3_w_n20585_0(.douta(w_n20585_0[0]),.doutb(w_n20585_0[1]),.doutc(w_n20585_0[2]),.din(n20585));
	jspl3 jspl3_w_n20587_0(.douta(w_n20587_0[0]),.doutb(w_n20587_0[1]),.doutc(w_n20587_0[2]),.din(n20587));
	jspl jspl_w_n20588_0(.douta(w_n20588_0[0]),.doutb(w_n20588_0[1]),.din(n20588));
	jspl3 jspl3_w_n20592_0(.douta(w_n20592_0[0]),.doutb(w_n20592_0[1]),.doutc(w_n20592_0[2]),.din(n20592));
	jspl3 jspl3_w_n20595_0(.douta(w_n20595_0[0]),.doutb(w_n20595_0[1]),.doutc(w_n20595_0[2]),.din(n20595));
	jspl jspl_w_n20596_0(.douta(w_n20596_0[0]),.doutb(w_n20596_0[1]),.din(n20596));
	jspl3 jspl3_w_n20600_0(.douta(w_n20600_0[0]),.doutb(w_n20600_0[1]),.doutc(w_n20600_0[2]),.din(n20600));
	jspl3 jspl3_w_n20602_0(.douta(w_n20602_0[0]),.doutb(w_n20602_0[1]),.doutc(w_n20602_0[2]),.din(n20602));
	jspl jspl_w_n20603_0(.douta(w_n20603_0[0]),.doutb(w_n20603_0[1]),.din(n20603));
	jspl3 jspl3_w_n20607_0(.douta(w_n20607_0[0]),.doutb(w_n20607_0[1]),.doutc(w_n20607_0[2]),.din(n20607));
	jspl3 jspl3_w_n20609_0(.douta(w_n20609_0[0]),.doutb(w_n20609_0[1]),.doutc(w_n20609_0[2]),.din(n20609));
	jspl jspl_w_n20610_0(.douta(w_n20610_0[0]),.doutb(w_n20610_0[1]),.din(n20610));
	jspl3 jspl3_w_n20614_0(.douta(w_n20614_0[0]),.doutb(w_n20614_0[1]),.doutc(w_n20614_0[2]),.din(n20614));
	jspl3 jspl3_w_n20617_0(.douta(w_n20617_0[0]),.doutb(w_n20617_0[1]),.doutc(w_n20617_0[2]),.din(n20617));
	jspl jspl_w_n20618_0(.douta(w_n20618_0[0]),.doutb(w_n20618_0[1]),.din(n20618));
	jspl3 jspl3_w_n20622_0(.douta(w_n20622_0[0]),.doutb(w_n20622_0[1]),.doutc(w_n20622_0[2]),.din(n20622));
	jspl3 jspl3_w_n20625_0(.douta(w_n20625_0[0]),.doutb(w_n20625_0[1]),.doutc(w_n20625_0[2]),.din(n20625));
	jspl jspl_w_n20626_0(.douta(w_n20626_0[0]),.doutb(w_n20626_0[1]),.din(n20626));
	jspl3 jspl3_w_n20630_0(.douta(w_n20630_0[0]),.doutb(w_n20630_0[1]),.doutc(w_n20630_0[2]),.din(n20630));
	jspl3 jspl3_w_n20632_0(.douta(w_n20632_0[0]),.doutb(w_n20632_0[1]),.doutc(w_n20632_0[2]),.din(n20632));
	jspl jspl_w_n20633_0(.douta(w_n20633_0[0]),.doutb(w_n20633_0[1]),.din(n20633));
	jspl3 jspl3_w_n20637_0(.douta(w_n20637_0[0]),.doutb(w_n20637_0[1]),.doutc(w_n20637_0[2]),.din(n20637));
	jspl3 jspl3_w_n20640_0(.douta(w_n20640_0[0]),.doutb(w_n20640_0[1]),.doutc(w_n20640_0[2]),.din(n20640));
	jspl jspl_w_n20641_0(.douta(w_n20641_0[0]),.doutb(w_n20641_0[1]),.din(n20641));
	jspl3 jspl3_w_n20645_0(.douta(w_n20645_0[0]),.doutb(w_n20645_0[1]),.doutc(w_n20645_0[2]),.din(n20645));
	jspl3 jspl3_w_n20647_0(.douta(w_n20647_0[0]),.doutb(w_n20647_0[1]),.doutc(w_n20647_0[2]),.din(n20647));
	jspl jspl_w_n20648_0(.douta(w_n20648_0[0]),.doutb(w_n20648_0[1]),.din(n20648));
	jspl3 jspl3_w_n20652_0(.douta(w_n20652_0[0]),.doutb(w_n20652_0[1]),.doutc(w_n20652_0[2]),.din(n20652));
	jspl3 jspl3_w_n20655_0(.douta(w_n20655_0[0]),.doutb(w_n20655_0[1]),.doutc(w_n20655_0[2]),.din(n20655));
	jspl jspl_w_n20656_0(.douta(w_n20656_0[0]),.doutb(w_n20656_0[1]),.din(n20656));
	jspl3 jspl3_w_n20660_0(.douta(w_n20660_0[0]),.doutb(w_n20660_0[1]),.doutc(w_n20660_0[2]),.din(n20660));
	jspl3 jspl3_w_n20662_0(.douta(w_n20662_0[0]),.doutb(w_n20662_0[1]),.doutc(w_n20662_0[2]),.din(n20662));
	jspl jspl_w_n20663_0(.douta(w_n20663_0[0]),.doutb(w_n20663_0[1]),.din(n20663));
	jspl3 jspl3_w_n20667_0(.douta(w_n20667_0[0]),.doutb(w_n20667_0[1]),.doutc(w_n20667_0[2]),.din(n20667));
	jspl3 jspl3_w_n20669_0(.douta(w_n20669_0[0]),.doutb(w_n20669_0[1]),.doutc(w_n20669_0[2]),.din(n20669));
	jspl jspl_w_n20670_0(.douta(w_n20670_0[0]),.doutb(w_n20670_0[1]),.din(n20670));
	jspl3 jspl3_w_n20674_0(.douta(w_n20674_0[0]),.doutb(w_n20674_0[1]),.doutc(w_n20674_0[2]),.din(n20674));
	jspl3 jspl3_w_n20676_0(.douta(w_n20676_0[0]),.doutb(w_n20676_0[1]),.doutc(w_n20676_0[2]),.din(n20676));
	jspl jspl_w_n20677_0(.douta(w_n20677_0[0]),.doutb(w_n20677_0[1]),.din(n20677));
	jspl3 jspl3_w_n20681_0(.douta(w_n20681_0[0]),.doutb(w_n20681_0[1]),.doutc(w_n20681_0[2]),.din(n20681));
	jspl3 jspl3_w_n20684_0(.douta(w_n20684_0[0]),.doutb(w_n20684_0[1]),.doutc(w_n20684_0[2]),.din(n20684));
	jspl jspl_w_n20685_0(.douta(w_n20685_0[0]),.doutb(w_n20685_0[1]),.din(n20685));
	jspl3 jspl3_w_n20689_0(.douta(w_n20689_0[0]),.doutb(w_n20689_0[1]),.doutc(w_n20689_0[2]),.din(n20689));
	jspl3 jspl3_w_n20691_0(.douta(w_n20691_0[0]),.doutb(w_n20691_0[1]),.doutc(w_n20691_0[2]),.din(n20691));
	jspl jspl_w_n20692_0(.douta(w_n20692_0[0]),.doutb(w_n20692_0[1]),.din(n20692));
	jspl3 jspl3_w_n20696_0(.douta(w_n20696_0[0]),.doutb(w_n20696_0[1]),.doutc(w_n20696_0[2]),.din(n20696));
	jspl3 jspl3_w_n20699_0(.douta(w_n20699_0[0]),.doutb(w_n20699_0[1]),.doutc(w_n20699_0[2]),.din(n20699));
	jspl jspl_w_n20700_0(.douta(w_n20700_0[0]),.doutb(w_n20700_0[1]),.din(n20700));
	jspl3 jspl3_w_n20704_0(.douta(w_n20704_0[0]),.doutb(w_n20704_0[1]),.doutc(w_n20704_0[2]),.din(n20704));
	jspl3 jspl3_w_n20706_0(.douta(w_n20706_0[0]),.doutb(w_n20706_0[1]),.doutc(w_n20706_0[2]),.din(n20706));
	jspl jspl_w_n20707_0(.douta(w_n20707_0[0]),.doutb(w_n20707_0[1]),.din(n20707));
	jspl3 jspl3_w_n20711_0(.douta(w_n20711_0[0]),.doutb(w_n20711_0[1]),.doutc(w_n20711_0[2]),.din(n20711));
	jspl3 jspl3_w_n20714_0(.douta(w_n20714_0[0]),.doutb(w_n20714_0[1]),.doutc(w_n20714_0[2]),.din(n20714));
	jspl jspl_w_n20715_0(.douta(w_n20715_0[0]),.doutb(w_n20715_0[1]),.din(n20715));
	jspl3 jspl3_w_n20719_0(.douta(w_n20719_0[0]),.doutb(w_n20719_0[1]),.doutc(w_n20719_0[2]),.din(n20719));
	jspl3 jspl3_w_n20721_0(.douta(w_n20721_0[0]),.doutb(w_n20721_0[1]),.doutc(w_n20721_0[2]),.din(n20721));
	jspl jspl_w_n20722_0(.douta(w_n20722_0[0]),.doutb(w_n20722_0[1]),.din(n20722));
	jspl3 jspl3_w_n20726_0(.douta(w_n20726_0[0]),.doutb(w_n20726_0[1]),.doutc(w_n20726_0[2]),.din(n20726));
	jspl3 jspl3_w_n20729_0(.douta(w_n20729_0[0]),.doutb(w_n20729_0[1]),.doutc(w_n20729_0[2]),.din(n20729));
	jspl jspl_w_n20730_0(.douta(w_n20730_0[0]),.doutb(w_n20730_0[1]),.din(n20730));
	jspl3 jspl3_w_n20734_0(.douta(w_n20734_0[0]),.doutb(w_n20734_0[1]),.doutc(w_n20734_0[2]),.din(n20734));
	jspl3 jspl3_w_n20736_0(.douta(w_n20736_0[0]),.doutb(w_n20736_0[1]),.doutc(w_n20736_0[2]),.din(n20736));
	jspl jspl_w_n20737_0(.douta(w_n20737_0[0]),.doutb(w_n20737_0[1]),.din(n20737));
	jspl3 jspl3_w_n20741_0(.douta(w_n20741_0[0]),.doutb(w_n20741_0[1]),.doutc(w_n20741_0[2]),.din(n20741));
	jspl3 jspl3_w_n20743_0(.douta(w_n20743_0[0]),.doutb(w_n20743_0[1]),.doutc(w_n20743_0[2]),.din(n20743));
	jspl jspl_w_n20744_0(.douta(w_n20744_0[0]),.doutb(w_n20744_0[1]),.din(n20744));
	jspl3 jspl3_w_n20748_0(.douta(w_n20748_0[0]),.doutb(w_n20748_0[1]),.doutc(w_n20748_0[2]),.din(n20748));
	jspl3 jspl3_w_n20750_0(.douta(w_n20750_0[0]),.doutb(w_n20750_0[1]),.doutc(w_n20750_0[2]),.din(n20750));
	jspl jspl_w_n20751_0(.douta(w_n20751_0[0]),.doutb(w_n20751_0[1]),.din(n20751));
	jspl3 jspl3_w_n20755_0(.douta(w_n20755_0[0]),.doutb(w_n20755_0[1]),.doutc(w_n20755_0[2]),.din(n20755));
	jspl3 jspl3_w_n20758_0(.douta(w_n20758_0[0]),.doutb(w_n20758_0[1]),.doutc(w_n20758_0[2]),.din(n20758));
	jspl jspl_w_n20759_0(.douta(w_n20759_0[0]),.doutb(w_n20759_0[1]),.din(n20759));
	jspl3 jspl3_w_n20763_0(.douta(w_n20763_0[0]),.doutb(w_n20763_0[1]),.doutc(w_n20763_0[2]),.din(n20763));
	jspl3 jspl3_w_n20765_0(.douta(w_n20765_0[0]),.doutb(w_n20765_0[1]),.doutc(w_n20765_0[2]),.din(n20765));
	jspl jspl_w_n20766_0(.douta(w_n20766_0[0]),.doutb(w_n20766_0[1]),.din(n20766));
	jspl3 jspl3_w_n20770_0(.douta(w_n20770_0[0]),.doutb(w_n20770_0[1]),.doutc(w_n20770_0[2]),.din(n20770));
	jspl3 jspl3_w_n20772_0(.douta(w_n20772_0[0]),.doutb(w_n20772_0[1]),.doutc(w_n20772_0[2]),.din(n20772));
	jspl jspl_w_n20773_0(.douta(w_n20773_0[0]),.doutb(w_n20773_0[1]),.din(n20773));
	jspl3 jspl3_w_n20777_0(.douta(w_n20777_0[0]),.doutb(w_n20777_0[1]),.doutc(w_n20777_0[2]),.din(n20777));
	jspl3 jspl3_w_n20779_0(.douta(w_n20779_0[0]),.doutb(w_n20779_0[1]),.doutc(w_n20779_0[2]),.din(n20779));
	jspl jspl_w_n20780_0(.douta(w_n20780_0[0]),.doutb(w_n20780_0[1]),.din(n20780));
	jspl3 jspl3_w_n20784_0(.douta(w_n20784_0[0]),.doutb(w_n20784_0[1]),.doutc(w_n20784_0[2]),.din(n20784));
	jspl3 jspl3_w_n20786_0(.douta(w_n20786_0[0]),.doutb(w_n20786_0[1]),.doutc(w_n20786_0[2]),.din(n20786));
	jspl jspl_w_n20787_0(.douta(w_n20787_0[0]),.doutb(w_n20787_0[1]),.din(n20787));
	jspl3 jspl3_w_n20791_0(.douta(w_n20791_0[0]),.doutb(w_n20791_0[1]),.doutc(w_n20791_0[2]),.din(n20791));
	jspl3 jspl3_w_n20793_0(.douta(w_n20793_0[0]),.doutb(w_n20793_0[1]),.doutc(w_n20793_0[2]),.din(n20793));
	jspl jspl_w_n20794_0(.douta(w_n20794_0[0]),.doutb(w_n20794_0[1]),.din(n20794));
	jspl3 jspl3_w_n20798_0(.douta(w_n20798_0[0]),.doutb(w_n20798_0[1]),.doutc(w_n20798_0[2]),.din(n20798));
	jspl3 jspl3_w_n20801_0(.douta(w_n20801_0[0]),.doutb(w_n20801_0[1]),.doutc(w_n20801_0[2]),.din(n20801));
	jspl jspl_w_n20802_0(.douta(w_n20802_0[0]),.doutb(w_n20802_0[1]),.din(n20802));
	jspl3 jspl3_w_n20806_0(.douta(w_n20806_0[0]),.doutb(w_n20806_0[1]),.doutc(w_n20806_0[2]),.din(n20806));
	jspl3 jspl3_w_n20808_0(.douta(w_n20808_0[0]),.doutb(w_n20808_0[1]),.doutc(w_n20808_0[2]),.din(n20808));
	jspl jspl_w_n20809_0(.douta(w_n20809_0[0]),.doutb(w_n20809_0[1]),.din(n20809));
	jspl3 jspl3_w_n20813_0(.douta(w_n20813_0[0]),.doutb(w_n20813_0[1]),.doutc(w_n20813_0[2]),.din(n20813));
	jspl3 jspl3_w_n20816_0(.douta(w_n20816_0[0]),.doutb(w_n20816_0[1]),.doutc(w_n20816_0[2]),.din(n20816));
	jspl jspl_w_n20817_0(.douta(w_n20817_0[0]),.doutb(w_n20817_0[1]),.din(n20817));
	jspl3 jspl3_w_n20821_0(.douta(w_n20821_0[0]),.doutb(w_n20821_0[1]),.doutc(w_n20821_0[2]),.din(n20821));
	jspl3 jspl3_w_n20823_0(.douta(w_n20823_0[0]),.doutb(w_n20823_0[1]),.doutc(w_n20823_0[2]),.din(n20823));
	jspl jspl_w_n20824_0(.douta(w_n20824_0[0]),.doutb(w_n20824_0[1]),.din(n20824));
	jspl3 jspl3_w_n20828_0(.douta(w_n20828_0[0]),.doutb(w_n20828_0[1]),.doutc(w_n20828_0[2]),.din(n20828));
	jspl3 jspl3_w_n20830_0(.douta(w_n20830_0[0]),.doutb(w_n20830_0[1]),.doutc(w_n20830_0[2]),.din(n20830));
	jspl jspl_w_n20831_0(.douta(w_n20831_0[0]),.doutb(w_n20831_0[1]),.din(n20831));
	jspl3 jspl3_w_n20835_0(.douta(w_n20835_0[0]),.doutb(w_n20835_0[1]),.doutc(w_n20835_0[2]),.din(n20835));
	jspl3 jspl3_w_n20838_0(.douta(w_n20838_0[0]),.doutb(w_n20838_0[1]),.doutc(w_n20838_0[2]),.din(n20838));
	jspl jspl_w_n20839_0(.douta(w_n20839_0[0]),.doutb(w_n20839_0[1]),.din(n20839));
	jspl3 jspl3_w_n20842_0(.douta(w_n20842_0[0]),.doutb(w_n20842_0[1]),.doutc(w_n20842_0[2]),.din(n20842));
	jspl3 jspl3_w_n20846_0(.douta(w_n20846_0[0]),.doutb(w_n20846_0[1]),.doutc(w_n20846_0[2]),.din(n20846));
	jspl jspl_w_n20847_0(.douta(w_n20847_0[0]),.doutb(w_n20847_0[1]),.din(n20847));
	jspl3 jspl3_w_n20851_0(.douta(w_n20851_0[0]),.doutb(w_n20851_0[1]),.doutc(w_n20851_0[2]),.din(n20851));
	jspl3 jspl3_w_n20853_0(.douta(w_n20853_0[0]),.doutb(w_n20853_0[1]),.doutc(w_n20853_0[2]),.din(n20853));
	jspl jspl_w_n20854_0(.douta(w_n20854_0[0]),.doutb(w_n20854_0[1]),.din(n20854));
	jspl jspl_w_n20858_0(.douta(w_n20858_0[0]),.doutb(w_n20858_0[1]),.din(n20858));
	jspl jspl_w_n20859_0(.douta(w_n20859_0[0]),.doutb(w_n20859_0[1]),.din(n20859));
	jspl3 jspl3_w_n20861_0(.douta(w_n20861_0[0]),.doutb(w_n20861_0[1]),.doutc(w_n20861_0[2]),.din(n20861));
	jspl jspl_w_n20862_0(.douta(w_n20862_0[0]),.doutb(w_n20862_0[1]),.din(n20862));
	jspl3 jspl3_w_n20866_0(.douta(w_n20866_0[0]),.doutb(w_n20866_0[1]),.doutc(w_n20866_0[2]),.din(n20866));
	jspl3 jspl3_w_n20868_0(.douta(w_n20868_0[0]),.doutb(w_n20868_0[1]),.doutc(w_n20868_0[2]),.din(n20868));
	jspl jspl_w_n20869_0(.douta(w_n20869_0[0]),.doutb(w_n20869_0[1]),.din(n20869));
	jspl3 jspl3_w_n20873_0(.douta(w_n20873_0[0]),.doutb(w_n20873_0[1]),.doutc(w_n20873_0[2]),.din(n20873));
	jspl3 jspl3_w_n20875_0(.douta(w_n20875_0[0]),.doutb(w_n20875_0[1]),.doutc(w_n20875_0[2]),.din(n20875));
	jspl jspl_w_n20876_0(.douta(w_n20876_0[0]),.doutb(w_n20876_0[1]),.din(n20876));
	jspl3 jspl3_w_n20880_0(.douta(w_n20880_0[0]),.doutb(w_n20880_0[1]),.doutc(w_n20880_0[2]),.din(n20880));
	jspl3 jspl3_w_n20883_0(.douta(w_n20883_0[0]),.doutb(w_n20883_0[1]),.doutc(w_n20883_0[2]),.din(n20883));
	jspl jspl_w_n20884_0(.douta(w_n20884_0[0]),.doutb(w_n20884_0[1]),.din(n20884));
	jspl3 jspl3_w_n20888_0(.douta(w_n20888_0[0]),.doutb(w_n20888_0[1]),.doutc(w_n20888_0[2]),.din(n20888));
	jspl3 jspl3_w_n20890_0(.douta(w_n20890_0[0]),.doutb(w_n20890_0[1]),.doutc(w_n20890_0[2]),.din(n20890));
	jspl jspl_w_n20891_0(.douta(w_n20891_0[0]),.doutb(w_n20891_0[1]),.din(n20891));
	jspl jspl_w_n20893_0(.douta(w_n20893_0[0]),.doutb(w_n20893_0[1]),.din(n20893));
	jspl jspl_w_n20896_0(.douta(w_n20896_0[0]),.doutb(w_n20896_0[1]),.din(n20896));
	jspl jspl_w_n20897_0(.douta(w_n20897_0[0]),.doutb(w_n20897_0[1]),.din(n20897));
	jspl jspl_w_n20902_0(.douta(w_n20902_0[0]),.doutb(w_n20902_0[1]),.din(n20902));
	jspl jspl_w_n20903_0(.douta(w_n20903_0[0]),.doutb(w_n20903_0[1]),.din(n20903));
	jspl3 jspl3_w_n20907_0(.douta(w_n20907_0[0]),.doutb(w_n20907_0[1]),.doutc(w_n20907_0[2]),.din(n20907));
	jspl3 jspl3_w_n20907_1(.douta(w_n20907_1[0]),.doutb(w_n20907_1[1]),.doutc(w_n20907_1[2]),.din(w_n20907_0[0]));
	jspl jspl_w_n20908_0(.douta(w_n20908_0[0]),.doutb(w_n20908_0[1]),.din(n20908));
	jspl3 jspl3_w_n20909_0(.douta(w_n20909_0[0]),.doutb(w_n20909_0[1]),.doutc(w_n20909_0[2]),.din(n20909));
	jspl jspl_w_n20910_0(.douta(w_n20910_0[0]),.doutb(w_n20910_0[1]),.din(n20910));
	jspl3 jspl3_w_n20912_0(.douta(w_n20912_0[0]),.doutb(w_n20912_0[1]),.doutc(w_n20912_0[2]),.din(n20912));
	jspl jspl_w_n20913_0(.douta(w_n20913_0[0]),.doutb(w_n20913_0[1]),.din(n20913));
	jspl jspl_w_n20978_0(.douta(w_n20978_0[0]),.doutb(w_n20978_0[1]),.din(n20978));
	jspl jspl_w_n21175_0(.douta(w_n21175_0[0]),.doutb(w_n21175_0[1]),.din(n21175));
	jspl jspl_w_n21176_0(.douta(w_n21176_0[0]),.doutb(w_n21176_0[1]),.din(n21176));
	jspl jspl_w_n21179_0(.douta(w_n21179_0[0]),.doutb(w_n21179_0[1]),.din(n21179));
	jspl3 jspl3_w_n21181_0(.douta(w_n21181_0[0]),.doutb(w_n21181_0[1]),.doutc(w_n21181_0[2]),.din(n21181));
	jspl jspl_w_n21181_1(.douta(w_n21181_1[0]),.doutb(w_n21181_1[1]),.din(w_n21181_0[0]));
	jspl3 jspl3_w_n21184_0(.douta(w_n21184_0[0]),.doutb(w_n21184_0[1]),.doutc(w_n21184_0[2]),.din(n21184));
	jspl3 jspl3_w_n21184_1(.douta(w_n21184_1[0]),.doutb(w_n21184_1[1]),.doutc(w_n21184_1[2]),.din(w_n21184_0[0]));
	jspl3 jspl3_w_n21184_2(.douta(w_n21184_2[0]),.doutb(w_n21184_2[1]),.doutc(w_n21184_2[2]),.din(w_n21184_0[1]));
	jspl3 jspl3_w_n21184_3(.douta(w_n21184_3[0]),.doutb(w_n21184_3[1]),.doutc(w_n21184_3[2]),.din(w_n21184_0[2]));
	jspl3 jspl3_w_n21184_4(.douta(w_n21184_4[0]),.doutb(w_n21184_4[1]),.doutc(w_n21184_4[2]),.din(w_n21184_1[0]));
	jspl3 jspl3_w_n21184_5(.douta(w_n21184_5[0]),.doutb(w_n21184_5[1]),.doutc(w_n21184_5[2]),.din(w_n21184_1[1]));
	jspl3 jspl3_w_n21184_6(.douta(w_n21184_6[0]),.doutb(w_n21184_6[1]),.doutc(w_n21184_6[2]),.din(w_n21184_1[2]));
	jspl3 jspl3_w_n21184_7(.douta(w_n21184_7[0]),.doutb(w_n21184_7[1]),.doutc(w_n21184_7[2]),.din(w_n21184_2[0]));
	jspl3 jspl3_w_n21188_0(.douta(w_n21188_0[0]),.doutb(w_n21188_0[1]),.doutc(w_n21188_0[2]),.din(n21188));
	jspl jspl_w_n21189_0(.douta(w_n21189_0[0]),.doutb(w_n21189_0[1]),.din(n21189));
	jspl jspl_w_n21191_0(.douta(w_n21191_0[0]),.doutb(w_n21191_0[1]),.din(n21191));
	jspl jspl_w_n21196_0(.douta(w_n21196_0[0]),.doutb(w_n21196_0[1]),.din(n21196));
	jspl jspl_w_n21197_0(.douta(w_n21197_0[0]),.doutb(w_n21197_0[1]),.din(n21197));
	jspl3 jspl3_w_n21199_0(.douta(w_n21199_0[0]),.doutb(w_n21199_0[1]),.doutc(w_n21199_0[2]),.din(n21199));
	jspl jspl_w_n21200_0(.douta(w_n21200_0[0]),.doutb(w_n21200_0[1]),.din(n21200));
	jspl jspl_w_n21204_0(.douta(w_n21204_0[0]),.doutb(w_n21204_0[1]),.din(n21204));
	jspl3 jspl3_w_n21206_0(.douta(w_n21206_0[0]),.doutb(w_n21206_0[1]),.doutc(w_n21206_0[2]),.din(n21206));
	jspl jspl_w_n21207_0(.douta(w_n21207_0[0]),.doutb(w_n21207_0[1]),.din(n21207));
	jspl jspl_w_n21211_0(.douta(w_n21211_0[0]),.doutb(w_n21211_0[1]),.din(n21211));
	jspl jspl_w_n21212_0(.douta(w_n21212_0[0]),.doutb(w_n21212_0[1]),.din(n21212));
	jspl3 jspl3_w_n21214_0(.douta(w_n21214_0[0]),.doutb(w_n21214_0[1]),.doutc(w_n21214_0[2]),.din(n21214));
	jspl jspl_w_n21215_0(.douta(w_n21215_0[0]),.doutb(w_n21215_0[1]),.din(n21215));
	jspl jspl_w_n21219_0(.douta(w_n21219_0[0]),.doutb(w_n21219_0[1]),.din(n21219));
	jspl3 jspl3_w_n21221_0(.douta(w_n21221_0[0]),.doutb(w_n21221_0[1]),.doutc(w_n21221_0[2]),.din(n21221));
	jspl jspl_w_n21222_0(.douta(w_n21222_0[0]),.doutb(w_n21222_0[1]),.din(n21222));
	jspl jspl_w_n21226_0(.douta(w_n21226_0[0]),.doutb(w_n21226_0[1]),.din(n21226));
	jspl jspl_w_n21227_0(.douta(w_n21227_0[0]),.doutb(w_n21227_0[1]),.din(n21227));
	jspl3 jspl3_w_n21229_0(.douta(w_n21229_0[0]),.doutb(w_n21229_0[1]),.doutc(w_n21229_0[2]),.din(n21229));
	jspl jspl_w_n21230_0(.douta(w_n21230_0[0]),.doutb(w_n21230_0[1]),.din(n21230));
	jspl jspl_w_n21234_0(.douta(w_n21234_0[0]),.doutb(w_n21234_0[1]),.din(n21234));
	jspl jspl_w_n21235_0(.douta(w_n21235_0[0]),.doutb(w_n21235_0[1]),.din(n21235));
	jspl3 jspl3_w_n21237_0(.douta(w_n21237_0[0]),.doutb(w_n21237_0[1]),.doutc(w_n21237_0[2]),.din(n21237));
	jspl jspl_w_n21238_0(.douta(w_n21238_0[0]),.doutb(w_n21238_0[1]),.din(n21238));
	jspl jspl_w_n21242_0(.douta(w_n21242_0[0]),.doutb(w_n21242_0[1]),.din(n21242));
	jspl jspl_w_n21243_0(.douta(w_n21243_0[0]),.doutb(w_n21243_0[1]),.din(n21243));
	jspl3 jspl3_w_n21245_0(.douta(w_n21245_0[0]),.doutb(w_n21245_0[1]),.doutc(w_n21245_0[2]),.din(n21245));
	jspl jspl_w_n21246_0(.douta(w_n21246_0[0]),.doutb(w_n21246_0[1]),.din(n21246));
	jspl jspl_w_n21250_0(.douta(w_n21250_0[0]),.doutb(w_n21250_0[1]),.din(n21250));
	jspl3 jspl3_w_n21252_0(.douta(w_n21252_0[0]),.doutb(w_n21252_0[1]),.doutc(w_n21252_0[2]),.din(n21252));
	jspl jspl_w_n21253_0(.douta(w_n21253_0[0]),.doutb(w_n21253_0[1]),.din(n21253));
	jspl jspl_w_n21257_0(.douta(w_n21257_0[0]),.doutb(w_n21257_0[1]),.din(n21257));
	jspl jspl_w_n21258_0(.douta(w_n21258_0[0]),.doutb(w_n21258_0[1]),.din(n21258));
	jspl3 jspl3_w_n21260_0(.douta(w_n21260_0[0]),.doutb(w_n21260_0[1]),.doutc(w_n21260_0[2]),.din(n21260));
	jspl jspl_w_n21261_0(.douta(w_n21261_0[0]),.doutb(w_n21261_0[1]),.din(n21261));
	jspl jspl_w_n21265_0(.douta(w_n21265_0[0]),.doutb(w_n21265_0[1]),.din(n21265));
	jspl jspl_w_n21266_0(.douta(w_n21266_0[0]),.doutb(w_n21266_0[1]),.din(n21266));
	jspl3 jspl3_w_n21268_0(.douta(w_n21268_0[0]),.doutb(w_n21268_0[1]),.doutc(w_n21268_0[2]),.din(n21268));
	jspl jspl_w_n21269_0(.douta(w_n21269_0[0]),.doutb(w_n21269_0[1]),.din(n21269));
	jspl jspl_w_n21273_0(.douta(w_n21273_0[0]),.doutb(w_n21273_0[1]),.din(n21273));
	jspl jspl_w_n21274_0(.douta(w_n21274_0[0]),.doutb(w_n21274_0[1]),.din(n21274));
	jspl3 jspl3_w_n21276_0(.douta(w_n21276_0[0]),.doutb(w_n21276_0[1]),.doutc(w_n21276_0[2]),.din(n21276));
	jspl jspl_w_n21277_0(.douta(w_n21277_0[0]),.doutb(w_n21277_0[1]),.din(n21277));
	jspl jspl_w_n21281_0(.douta(w_n21281_0[0]),.doutb(w_n21281_0[1]),.din(n21281));
	jspl3 jspl3_w_n21283_0(.douta(w_n21283_0[0]),.doutb(w_n21283_0[1]),.doutc(w_n21283_0[2]),.din(n21283));
	jspl jspl_w_n21284_0(.douta(w_n21284_0[0]),.doutb(w_n21284_0[1]),.din(n21284));
	jspl jspl_w_n21288_0(.douta(w_n21288_0[0]),.doutb(w_n21288_0[1]),.din(n21288));
	jspl jspl_w_n21289_0(.douta(w_n21289_0[0]),.doutb(w_n21289_0[1]),.din(n21289));
	jspl3 jspl3_w_n21291_0(.douta(w_n21291_0[0]),.doutb(w_n21291_0[1]),.doutc(w_n21291_0[2]),.din(n21291));
	jspl jspl_w_n21292_0(.douta(w_n21292_0[0]),.doutb(w_n21292_0[1]),.din(n21292));
	jspl jspl_w_n21296_0(.douta(w_n21296_0[0]),.doutb(w_n21296_0[1]),.din(n21296));
	jspl3 jspl3_w_n21298_0(.douta(w_n21298_0[0]),.doutb(w_n21298_0[1]),.doutc(w_n21298_0[2]),.din(n21298));
	jspl jspl_w_n21299_0(.douta(w_n21299_0[0]),.doutb(w_n21299_0[1]),.din(n21299));
	jspl jspl_w_n21303_0(.douta(w_n21303_0[0]),.doutb(w_n21303_0[1]),.din(n21303));
	jspl jspl_w_n21304_0(.douta(w_n21304_0[0]),.doutb(w_n21304_0[1]),.din(n21304));
	jspl3 jspl3_w_n21306_0(.douta(w_n21306_0[0]),.doutb(w_n21306_0[1]),.doutc(w_n21306_0[2]),.din(n21306));
	jspl jspl_w_n21307_0(.douta(w_n21307_0[0]),.doutb(w_n21307_0[1]),.din(n21307));
	jspl jspl_w_n21311_0(.douta(w_n21311_0[0]),.doutb(w_n21311_0[1]),.din(n21311));
	jspl3 jspl3_w_n21313_0(.douta(w_n21313_0[0]),.doutb(w_n21313_0[1]),.doutc(w_n21313_0[2]),.din(n21313));
	jspl jspl_w_n21314_0(.douta(w_n21314_0[0]),.doutb(w_n21314_0[1]),.din(n21314));
	jspl jspl_w_n21318_0(.douta(w_n21318_0[0]),.doutb(w_n21318_0[1]),.din(n21318));
	jspl jspl_w_n21319_0(.douta(w_n21319_0[0]),.doutb(w_n21319_0[1]),.din(n21319));
	jspl3 jspl3_w_n21321_0(.douta(w_n21321_0[0]),.doutb(w_n21321_0[1]),.doutc(w_n21321_0[2]),.din(n21321));
	jspl jspl_w_n21322_0(.douta(w_n21322_0[0]),.doutb(w_n21322_0[1]),.din(n21322));
	jspl jspl_w_n21326_0(.douta(w_n21326_0[0]),.doutb(w_n21326_0[1]),.din(n21326));
	jspl jspl_w_n21327_0(.douta(w_n21327_0[0]),.doutb(w_n21327_0[1]),.din(n21327));
	jspl3 jspl3_w_n21329_0(.douta(w_n21329_0[0]),.doutb(w_n21329_0[1]),.doutc(w_n21329_0[2]),.din(n21329));
	jspl jspl_w_n21330_0(.douta(w_n21330_0[0]),.doutb(w_n21330_0[1]),.din(n21330));
	jspl jspl_w_n21334_0(.douta(w_n21334_0[0]),.doutb(w_n21334_0[1]),.din(n21334));
	jspl3 jspl3_w_n21336_0(.douta(w_n21336_0[0]),.doutb(w_n21336_0[1]),.doutc(w_n21336_0[2]),.din(n21336));
	jspl jspl_w_n21337_0(.douta(w_n21337_0[0]),.doutb(w_n21337_0[1]),.din(n21337));
	jspl jspl_w_n21341_0(.douta(w_n21341_0[0]),.doutb(w_n21341_0[1]),.din(n21341));
	jspl3 jspl3_w_n21343_0(.douta(w_n21343_0[0]),.doutb(w_n21343_0[1]),.doutc(w_n21343_0[2]),.din(n21343));
	jspl jspl_w_n21344_0(.douta(w_n21344_0[0]),.doutb(w_n21344_0[1]),.din(n21344));
	jspl jspl_w_n21348_0(.douta(w_n21348_0[0]),.doutb(w_n21348_0[1]),.din(n21348));
	jspl jspl_w_n21349_0(.douta(w_n21349_0[0]),.doutb(w_n21349_0[1]),.din(n21349));
	jspl3 jspl3_w_n21351_0(.douta(w_n21351_0[0]),.doutb(w_n21351_0[1]),.doutc(w_n21351_0[2]),.din(n21351));
	jspl jspl_w_n21352_0(.douta(w_n21352_0[0]),.doutb(w_n21352_0[1]),.din(n21352));
	jspl jspl_w_n21356_0(.douta(w_n21356_0[0]),.doutb(w_n21356_0[1]),.din(n21356));
	jspl3 jspl3_w_n21358_0(.douta(w_n21358_0[0]),.doutb(w_n21358_0[1]),.doutc(w_n21358_0[2]),.din(n21358));
	jspl jspl_w_n21359_0(.douta(w_n21359_0[0]),.doutb(w_n21359_0[1]),.din(n21359));
	jspl jspl_w_n21363_0(.douta(w_n21363_0[0]),.doutb(w_n21363_0[1]),.din(n21363));
	jspl jspl_w_n21364_0(.douta(w_n21364_0[0]),.doutb(w_n21364_0[1]),.din(n21364));
	jspl3 jspl3_w_n21366_0(.douta(w_n21366_0[0]),.doutb(w_n21366_0[1]),.doutc(w_n21366_0[2]),.din(n21366));
	jspl jspl_w_n21367_0(.douta(w_n21367_0[0]),.doutb(w_n21367_0[1]),.din(n21367));
	jspl jspl_w_n21371_0(.douta(w_n21371_0[0]),.doutb(w_n21371_0[1]),.din(n21371));
	jspl3 jspl3_w_n21373_0(.douta(w_n21373_0[0]),.doutb(w_n21373_0[1]),.doutc(w_n21373_0[2]),.din(n21373));
	jspl jspl_w_n21374_0(.douta(w_n21374_0[0]),.doutb(w_n21374_0[1]),.din(n21374));
	jspl jspl_w_n21378_0(.douta(w_n21378_0[0]),.doutb(w_n21378_0[1]),.din(n21378));
	jspl jspl_w_n21379_0(.douta(w_n21379_0[0]),.doutb(w_n21379_0[1]),.din(n21379));
	jspl3 jspl3_w_n21381_0(.douta(w_n21381_0[0]),.doutb(w_n21381_0[1]),.doutc(w_n21381_0[2]),.din(n21381));
	jspl jspl_w_n21382_0(.douta(w_n21382_0[0]),.doutb(w_n21382_0[1]),.din(n21382));
	jspl jspl_w_n21386_0(.douta(w_n21386_0[0]),.doutb(w_n21386_0[1]),.din(n21386));
	jspl jspl_w_n21387_0(.douta(w_n21387_0[0]),.doutb(w_n21387_0[1]),.din(n21387));
	jspl3 jspl3_w_n21389_0(.douta(w_n21389_0[0]),.doutb(w_n21389_0[1]),.doutc(w_n21389_0[2]),.din(n21389));
	jspl jspl_w_n21390_0(.douta(w_n21390_0[0]),.doutb(w_n21390_0[1]),.din(n21390));
	jspl jspl_w_n21394_0(.douta(w_n21394_0[0]),.doutb(w_n21394_0[1]),.din(n21394));
	jspl jspl_w_n21395_0(.douta(w_n21395_0[0]),.doutb(w_n21395_0[1]),.din(n21395));
	jspl3 jspl3_w_n21397_0(.douta(w_n21397_0[0]),.doutb(w_n21397_0[1]),.doutc(w_n21397_0[2]),.din(n21397));
	jspl jspl_w_n21398_0(.douta(w_n21398_0[0]),.doutb(w_n21398_0[1]),.din(n21398));
	jspl jspl_w_n21402_0(.douta(w_n21402_0[0]),.doutb(w_n21402_0[1]),.din(n21402));
	jspl3 jspl3_w_n21404_0(.douta(w_n21404_0[0]),.doutb(w_n21404_0[1]),.doutc(w_n21404_0[2]),.din(n21404));
	jspl jspl_w_n21405_0(.douta(w_n21405_0[0]),.doutb(w_n21405_0[1]),.din(n21405));
	jspl jspl_w_n21409_0(.douta(w_n21409_0[0]),.doutb(w_n21409_0[1]),.din(n21409));
	jspl jspl_w_n21410_0(.douta(w_n21410_0[0]),.doutb(w_n21410_0[1]),.din(n21410));
	jspl3 jspl3_w_n21412_0(.douta(w_n21412_0[0]),.doutb(w_n21412_0[1]),.doutc(w_n21412_0[2]),.din(n21412));
	jspl jspl_w_n21413_0(.douta(w_n21413_0[0]),.doutb(w_n21413_0[1]),.din(n21413));
	jspl jspl_w_n21417_0(.douta(w_n21417_0[0]),.doutb(w_n21417_0[1]),.din(n21417));
	jspl3 jspl3_w_n21419_0(.douta(w_n21419_0[0]),.doutb(w_n21419_0[1]),.doutc(w_n21419_0[2]),.din(n21419));
	jspl jspl_w_n21420_0(.douta(w_n21420_0[0]),.doutb(w_n21420_0[1]),.din(n21420));
	jspl jspl_w_n21424_0(.douta(w_n21424_0[0]),.doutb(w_n21424_0[1]),.din(n21424));
	jspl jspl_w_n21425_0(.douta(w_n21425_0[0]),.doutb(w_n21425_0[1]),.din(n21425));
	jspl3 jspl3_w_n21427_0(.douta(w_n21427_0[0]),.doutb(w_n21427_0[1]),.doutc(w_n21427_0[2]),.din(n21427));
	jspl jspl_w_n21428_0(.douta(w_n21428_0[0]),.doutb(w_n21428_0[1]),.din(n21428));
	jspl jspl_w_n21432_0(.douta(w_n21432_0[0]),.doutb(w_n21432_0[1]),.din(n21432));
	jspl3 jspl3_w_n21434_0(.douta(w_n21434_0[0]),.doutb(w_n21434_0[1]),.doutc(w_n21434_0[2]),.din(n21434));
	jspl jspl_w_n21435_0(.douta(w_n21435_0[0]),.doutb(w_n21435_0[1]),.din(n21435));
	jspl jspl_w_n21439_0(.douta(w_n21439_0[0]),.doutb(w_n21439_0[1]),.din(n21439));
	jspl jspl_w_n21440_0(.douta(w_n21440_0[0]),.doutb(w_n21440_0[1]),.din(n21440));
	jspl3 jspl3_w_n21442_0(.douta(w_n21442_0[0]),.doutb(w_n21442_0[1]),.doutc(w_n21442_0[2]),.din(n21442));
	jspl jspl_w_n21443_0(.douta(w_n21443_0[0]),.doutb(w_n21443_0[1]),.din(n21443));
	jspl jspl_w_n21447_0(.douta(w_n21447_0[0]),.doutb(w_n21447_0[1]),.din(n21447));
	jspl3 jspl3_w_n21449_0(.douta(w_n21449_0[0]),.doutb(w_n21449_0[1]),.doutc(w_n21449_0[2]),.din(n21449));
	jspl jspl_w_n21450_0(.douta(w_n21450_0[0]),.doutb(w_n21450_0[1]),.din(n21450));
	jspl jspl_w_n21454_0(.douta(w_n21454_0[0]),.doutb(w_n21454_0[1]),.din(n21454));
	jspl jspl_w_n21455_0(.douta(w_n21455_0[0]),.doutb(w_n21455_0[1]),.din(n21455));
	jspl3 jspl3_w_n21457_0(.douta(w_n21457_0[0]),.doutb(w_n21457_0[1]),.doutc(w_n21457_0[2]),.din(n21457));
	jspl jspl_w_n21458_0(.douta(w_n21458_0[0]),.doutb(w_n21458_0[1]),.din(n21458));
	jspl jspl_w_n21462_0(.douta(w_n21462_0[0]),.doutb(w_n21462_0[1]),.din(n21462));
	jspl jspl_w_n21463_0(.douta(w_n21463_0[0]),.doutb(w_n21463_0[1]),.din(n21463));
	jspl3 jspl3_w_n21465_0(.douta(w_n21465_0[0]),.doutb(w_n21465_0[1]),.doutc(w_n21465_0[2]),.din(n21465));
	jspl jspl_w_n21466_0(.douta(w_n21466_0[0]),.doutb(w_n21466_0[1]),.din(n21466));
	jspl jspl_w_n21470_0(.douta(w_n21470_0[0]),.doutb(w_n21470_0[1]),.din(n21470));
	jspl jspl_w_n21471_0(.douta(w_n21471_0[0]),.doutb(w_n21471_0[1]),.din(n21471));
	jspl3 jspl3_w_n21473_0(.douta(w_n21473_0[0]),.doutb(w_n21473_0[1]),.doutc(w_n21473_0[2]),.din(n21473));
	jspl jspl_w_n21474_0(.douta(w_n21474_0[0]),.doutb(w_n21474_0[1]),.din(n21474));
	jspl jspl_w_n21478_0(.douta(w_n21478_0[0]),.doutb(w_n21478_0[1]),.din(n21478));
	jspl3 jspl3_w_n21480_0(.douta(w_n21480_0[0]),.doutb(w_n21480_0[1]),.doutc(w_n21480_0[2]),.din(n21480));
	jspl jspl_w_n21481_0(.douta(w_n21481_0[0]),.doutb(w_n21481_0[1]),.din(n21481));
	jspl jspl_w_n21485_0(.douta(w_n21485_0[0]),.doutb(w_n21485_0[1]),.din(n21485));
	jspl jspl_w_n21486_0(.douta(w_n21486_0[0]),.doutb(w_n21486_0[1]),.din(n21486));
	jspl3 jspl3_w_n21488_0(.douta(w_n21488_0[0]),.doutb(w_n21488_0[1]),.doutc(w_n21488_0[2]),.din(n21488));
	jspl jspl_w_n21489_0(.douta(w_n21489_0[0]),.doutb(w_n21489_0[1]),.din(n21489));
	jspl jspl_w_n21493_0(.douta(w_n21493_0[0]),.doutb(w_n21493_0[1]),.din(n21493));
	jspl jspl_w_n21494_0(.douta(w_n21494_0[0]),.doutb(w_n21494_0[1]),.din(n21494));
	jspl3 jspl3_w_n21496_0(.douta(w_n21496_0[0]),.doutb(w_n21496_0[1]),.doutc(w_n21496_0[2]),.din(n21496));
	jspl jspl_w_n21497_0(.douta(w_n21497_0[0]),.doutb(w_n21497_0[1]),.din(n21497));
	jspl jspl_w_n21501_0(.douta(w_n21501_0[0]),.doutb(w_n21501_0[1]),.din(n21501));
	jspl jspl_w_n21502_0(.douta(w_n21502_0[0]),.doutb(w_n21502_0[1]),.din(n21502));
	jspl3 jspl3_w_n21504_0(.douta(w_n21504_0[0]),.doutb(w_n21504_0[1]),.doutc(w_n21504_0[2]),.din(n21504));
	jspl jspl_w_n21505_0(.douta(w_n21505_0[0]),.doutb(w_n21505_0[1]),.din(n21505));
	jspl jspl_w_n21509_0(.douta(w_n21509_0[0]),.doutb(w_n21509_0[1]),.din(n21509));
	jspl jspl_w_n21510_0(.douta(w_n21510_0[0]),.doutb(w_n21510_0[1]),.din(n21510));
	jspl3 jspl3_w_n21512_0(.douta(w_n21512_0[0]),.doutb(w_n21512_0[1]),.doutc(w_n21512_0[2]),.din(n21512));
	jspl jspl_w_n21513_0(.douta(w_n21513_0[0]),.doutb(w_n21513_0[1]),.din(n21513));
	jspl jspl_w_n21517_0(.douta(w_n21517_0[0]),.doutb(w_n21517_0[1]),.din(n21517));
	jspl jspl_w_n21518_0(.douta(w_n21518_0[0]),.doutb(w_n21518_0[1]),.din(n21518));
	jspl3 jspl3_w_n21520_0(.douta(w_n21520_0[0]),.doutb(w_n21520_0[1]),.doutc(w_n21520_0[2]),.din(n21520));
	jspl jspl_w_n21521_0(.douta(w_n21521_0[0]),.doutb(w_n21521_0[1]),.din(n21521));
	jspl jspl_w_n21525_0(.douta(w_n21525_0[0]),.doutb(w_n21525_0[1]),.din(n21525));
	jspl3 jspl3_w_n21527_0(.douta(w_n21527_0[0]),.doutb(w_n21527_0[1]),.doutc(w_n21527_0[2]),.din(n21527));
	jspl jspl_w_n21528_0(.douta(w_n21528_0[0]),.doutb(w_n21528_0[1]),.din(n21528));
	jspl jspl_w_n21532_0(.douta(w_n21532_0[0]),.doutb(w_n21532_0[1]),.din(n21532));
	jspl jspl_w_n21533_0(.douta(w_n21533_0[0]),.doutb(w_n21533_0[1]),.din(n21533));
	jspl3 jspl3_w_n21535_0(.douta(w_n21535_0[0]),.doutb(w_n21535_0[1]),.doutc(w_n21535_0[2]),.din(n21535));
	jspl jspl_w_n21536_0(.douta(w_n21536_0[0]),.doutb(w_n21536_0[1]),.din(n21536));
	jspl jspl_w_n21540_0(.douta(w_n21540_0[0]),.doutb(w_n21540_0[1]),.din(n21540));
	jspl3 jspl3_w_n21542_0(.douta(w_n21542_0[0]),.doutb(w_n21542_0[1]),.doutc(w_n21542_0[2]),.din(n21542));
	jspl jspl_w_n21543_0(.douta(w_n21543_0[0]),.doutb(w_n21543_0[1]),.din(n21543));
	jspl jspl_w_n21547_0(.douta(w_n21547_0[0]),.doutb(w_n21547_0[1]),.din(n21547));
	jspl jspl_w_n21548_0(.douta(w_n21548_0[0]),.doutb(w_n21548_0[1]),.din(n21548));
	jspl3 jspl3_w_n21550_0(.douta(w_n21550_0[0]),.doutb(w_n21550_0[1]),.doutc(w_n21550_0[2]),.din(n21550));
	jspl jspl_w_n21551_0(.douta(w_n21551_0[0]),.doutb(w_n21551_0[1]),.din(n21551));
	jspl jspl_w_n21555_0(.douta(w_n21555_0[0]),.doutb(w_n21555_0[1]),.din(n21555));
	jspl jspl_w_n21556_0(.douta(w_n21556_0[0]),.doutb(w_n21556_0[1]),.din(n21556));
	jspl3 jspl3_w_n21558_0(.douta(w_n21558_0[0]),.doutb(w_n21558_0[1]),.doutc(w_n21558_0[2]),.din(n21558));
	jspl jspl_w_n21559_0(.douta(w_n21559_0[0]),.doutb(w_n21559_0[1]),.din(n21559));
	jspl jspl_w_n21563_0(.douta(w_n21563_0[0]),.doutb(w_n21563_0[1]),.din(n21563));
	jspl3 jspl3_w_n21565_0(.douta(w_n21565_0[0]),.doutb(w_n21565_0[1]),.doutc(w_n21565_0[2]),.din(n21565));
	jspl jspl_w_n21566_0(.douta(w_n21566_0[0]),.doutb(w_n21566_0[1]),.din(n21566));
	jspl jspl_w_n21570_0(.douta(w_n21570_0[0]),.doutb(w_n21570_0[1]),.din(n21570));
	jspl3 jspl3_w_n21572_0(.douta(w_n21572_0[0]),.doutb(w_n21572_0[1]),.doutc(w_n21572_0[2]),.din(n21572));
	jspl jspl_w_n21573_0(.douta(w_n21573_0[0]),.doutb(w_n21573_0[1]),.din(n21573));
	jspl jspl_w_n21577_0(.douta(w_n21577_0[0]),.doutb(w_n21577_0[1]),.din(n21577));
	jspl jspl_w_n21578_0(.douta(w_n21578_0[0]),.doutb(w_n21578_0[1]),.din(n21578));
	jspl3 jspl3_w_n21580_0(.douta(w_n21580_0[0]),.doutb(w_n21580_0[1]),.doutc(w_n21580_0[2]),.din(n21580));
	jspl jspl_w_n21581_0(.douta(w_n21581_0[0]),.doutb(w_n21581_0[1]),.din(n21581));
	jspl jspl_w_n21585_0(.douta(w_n21585_0[0]),.doutb(w_n21585_0[1]),.din(n21585));
	jspl jspl_w_n21586_0(.douta(w_n21586_0[0]),.doutb(w_n21586_0[1]),.din(n21586));
	jspl3 jspl3_w_n21588_0(.douta(w_n21588_0[0]),.doutb(w_n21588_0[1]),.doutc(w_n21588_0[2]),.din(n21588));
	jspl jspl_w_n21589_0(.douta(w_n21589_0[0]),.doutb(w_n21589_0[1]),.din(n21589));
	jspl jspl_w_n21593_0(.douta(w_n21593_0[0]),.doutb(w_n21593_0[1]),.din(n21593));
	jspl jspl_w_n21594_0(.douta(w_n21594_0[0]),.doutb(w_n21594_0[1]),.din(n21594));
	jspl3 jspl3_w_n21596_0(.douta(w_n21596_0[0]),.doutb(w_n21596_0[1]),.doutc(w_n21596_0[2]),.din(n21596));
	jspl jspl_w_n21597_0(.douta(w_n21597_0[0]),.doutb(w_n21597_0[1]),.din(n21597));
	jspl3 jspl3_w_n21601_0(.douta(w_n21601_0[0]),.doutb(w_n21601_0[1]),.doutc(w_n21601_0[2]),.din(n21601));
	jspl3 jspl3_w_n21604_0(.douta(w_n21604_0[0]),.doutb(w_n21604_0[1]),.doutc(w_n21604_0[2]),.din(n21604));
	jspl jspl_w_n21605_0(.douta(w_n21605_0[0]),.doutb(w_n21605_0[1]),.din(n21605));
	jspl3 jspl3_w_n21609_0(.douta(w_n21609_0[0]),.doutb(w_n21609_0[1]),.doutc(w_n21609_0[2]),.din(n21609));
	jspl3 jspl3_w_n21611_0(.douta(w_n21611_0[0]),.doutb(w_n21611_0[1]),.doutc(w_n21611_0[2]),.din(n21611));
	jspl jspl_w_n21614_0(.douta(w_n21614_0[0]),.doutb(w_n21614_0[1]),.din(n21614));
	jspl3 jspl3_w_n21615_0(.douta(w_n21615_0[0]),.doutb(w_n21615_0[1]),.doutc(w_n21615_0[2]),.din(n21615));
	jspl jspl_w_n21616_0(.douta(w_n21616_0[0]),.doutb(w_n21616_0[1]),.din(n21616));
	jspl jspl_w_n21618_0(.douta(w_n21618_0[0]),.doutb(w_n21618_0[1]),.din(n21618));
	jspl jspl_w_n21681_0(.douta(w_n21681_0[0]),.doutb(w_n21681_0[1]),.din(n21681));
	jspl jspl_w_n21688_0(.douta(w_n21688_0[0]),.doutb(w_n21688_0[1]),.din(n21688));
	jspl jspl_w_n21695_0(.douta(w_n21695_0[0]),.doutb(w_n21695_0[1]),.din(n21695));
	jspl jspl_w_n21708_0(.douta(w_n21708_0[0]),.doutb(w_n21708_0[1]),.din(n21708));
	jspl jspl_w_n21721_0(.douta(w_n21721_0[0]),.doutb(w_n21721_0[1]),.din(n21721));
	jspl jspl_w_n21728_0(.douta(w_n21728_0[0]),.doutb(w_n21728_0[1]),.din(n21728));
	jspl jspl_w_n21735_0(.douta(w_n21735_0[0]),.doutb(w_n21735_0[1]),.din(n21735));
	jspl jspl_w_n21745_0(.douta(w_n21745_0[0]),.doutb(w_n21745_0[1]),.din(n21745));
	jspl jspl_w_n21749_0(.douta(w_n21749_0[0]),.doutb(w_n21749_0[1]),.din(n21749));
	jspl jspl_w_n21756_0(.douta(w_n21756_0[0]),.doutb(w_n21756_0[1]),.din(n21756));
	jspl jspl_w_n21763_0(.douta(w_n21763_0[0]),.doutb(w_n21763_0[1]),.din(n21763));
	jspl jspl_w_n21776_0(.douta(w_n21776_0[0]),.doutb(w_n21776_0[1]),.din(n21776));
	jspl jspl_w_n21783_0(.douta(w_n21783_0[0]),.doutb(w_n21783_0[1]),.din(n21783));
	jspl jspl_w_n21790_0(.douta(w_n21790_0[0]),.doutb(w_n21790_0[1]),.din(n21790));
	jspl jspl_w_n21797_0(.douta(w_n21797_0[0]),.doutb(w_n21797_0[1]),.din(n21797));
	jspl jspl_w_n21810_0(.douta(w_n21810_0[0]),.doutb(w_n21810_0[1]),.din(n21810));
	jspl jspl_w_n21829_0(.douta(w_n21829_0[0]),.doutb(w_n21829_0[1]),.din(n21829));
	jspl jspl_w_n21836_0(.douta(w_n21836_0[0]),.doutb(w_n21836_0[1]),.din(n21836));
	jspl jspl_w_n21846_0(.douta(w_n21846_0[0]),.doutb(w_n21846_0[1]),.din(n21846));
	jspl jspl_w_n21850_0(.douta(w_n21850_0[0]),.doutb(w_n21850_0[1]),.din(n21850));
	jspl jspl_w_n21868_0(.douta(w_n21868_0[0]),.doutb(w_n21868_0[1]),.din(n21868));
	jspl jspl_w_n21877_0(.douta(w_n21877_0[0]),.doutb(w_n21877_0[1]),.din(n21877));
	jspl3 jspl3_w_n21887_0(.douta(w_n21887_0[0]),.doutb(w_n21887_0[1]),.doutc(w_n21887_0[2]),.din(n21887));
	jspl3 jspl3_w_n21887_1(.douta(w_n21887_1[0]),.doutb(w_n21887_1[1]),.doutc(w_n21887_1[2]),.din(w_n21887_0[0]));
	jspl3 jspl3_w_n21887_2(.douta(w_n21887_2[0]),.doutb(w_n21887_2[1]),.doutc(w_n21887_2[2]),.din(w_n21887_0[1]));
	jspl3 jspl3_w_n21887_3(.douta(w_n21887_3[0]),.doutb(w_n21887_3[1]),.doutc(w_n21887_3[2]),.din(w_n21887_0[2]));
	jspl3 jspl3_w_n21887_4(.douta(w_n21887_4[0]),.doutb(w_n21887_4[1]),.doutc(w_n21887_4[2]),.din(w_n21887_1[0]));
	jspl3 jspl3_w_n21887_5(.douta(w_n21887_5[0]),.doutb(w_n21887_5[1]),.doutc(w_n21887_5[2]),.din(w_n21887_1[1]));
	jspl3 jspl3_w_n21887_6(.douta(w_n21887_6[0]),.doutb(w_n21887_6[1]),.doutc(w_n21887_6[2]),.din(w_n21887_1[2]));
	jspl3 jspl3_w_n21887_7(.douta(w_n21887_7[0]),.doutb(w_n21887_7[1]),.doutc(w_n21887_7[2]),.din(w_n21887_2[0]));
	jspl3 jspl3_w_n21887_8(.douta(w_n21887_8[0]),.doutb(w_n21887_8[1]),.doutc(w_n21887_8[2]),.din(w_n21887_2[1]));
	jspl3 jspl3_w_n21887_9(.douta(w_n21887_9[0]),.doutb(w_n21887_9[1]),.doutc(w_n21887_9[2]),.din(w_n21887_2[2]));
	jspl3 jspl3_w_n21887_10(.douta(w_n21887_10[0]),.doutb(w_n21887_10[1]),.doutc(w_n21887_10[2]),.din(w_n21887_3[0]));
	jspl3 jspl3_w_n21887_11(.douta(w_n21887_11[0]),.doutb(w_n21887_11[1]),.doutc(w_n21887_11[2]),.din(w_n21887_3[1]));
	jspl3 jspl3_w_n21887_12(.douta(w_n21887_12[0]),.doutb(w_n21887_12[1]),.doutc(w_n21887_12[2]),.din(w_n21887_3[2]));
	jspl3 jspl3_w_n21887_13(.douta(w_n21887_13[0]),.doutb(w_n21887_13[1]),.doutc(w_n21887_13[2]),.din(w_n21887_4[0]));
	jspl3 jspl3_w_n21887_14(.douta(w_n21887_14[0]),.doutb(w_n21887_14[1]),.doutc(w_n21887_14[2]),.din(w_n21887_4[1]));
	jspl3 jspl3_w_n21887_15(.douta(w_n21887_15[0]),.doutb(w_n21887_15[1]),.doutc(w_n21887_15[2]),.din(w_n21887_4[2]));
	jspl3 jspl3_w_n21887_16(.douta(w_n21887_16[0]),.doutb(w_n21887_16[1]),.doutc(w_n21887_16[2]),.din(w_n21887_5[0]));
	jspl3 jspl3_w_n21887_17(.douta(w_n21887_17[0]),.doutb(w_n21887_17[1]),.doutc(w_n21887_17[2]),.din(w_n21887_5[1]));
	jspl3 jspl3_w_n21887_18(.douta(w_n21887_18[0]),.doutb(w_n21887_18[1]),.doutc(w_n21887_18[2]),.din(w_n21887_5[2]));
	jspl3 jspl3_w_n21887_19(.douta(w_n21887_19[0]),.doutb(w_n21887_19[1]),.doutc(w_n21887_19[2]),.din(w_n21887_6[0]));
	jspl3 jspl3_w_n21887_20(.douta(w_n21887_20[0]),.doutb(w_n21887_20[1]),.doutc(w_n21887_20[2]),.din(w_n21887_6[1]));
	jspl3 jspl3_w_n21887_21(.douta(w_n21887_21[0]),.doutb(w_n21887_21[1]),.doutc(w_n21887_21[2]),.din(w_n21887_6[2]));
	jspl3 jspl3_w_n21887_22(.douta(w_n21887_22[0]),.doutb(w_n21887_22[1]),.doutc(w_n21887_22[2]),.din(w_n21887_7[0]));
	jspl3 jspl3_w_n21887_23(.douta(w_n21887_23[0]),.doutb(w_n21887_23[1]),.doutc(w_n21887_23[2]),.din(w_n21887_7[1]));
	jspl3 jspl3_w_n21887_24(.douta(w_n21887_24[0]),.doutb(w_n21887_24[1]),.doutc(w_n21887_24[2]),.din(w_n21887_7[2]));
	jspl3 jspl3_w_n21887_25(.douta(w_n21887_25[0]),.doutb(w_n21887_25[1]),.doutc(w_n21887_25[2]),.din(w_n21887_8[0]));
	jspl3 jspl3_w_n21887_26(.douta(w_n21887_26[0]),.doutb(w_n21887_26[1]),.doutc(w_n21887_26[2]),.din(w_n21887_8[1]));
	jspl3 jspl3_w_n21887_27(.douta(w_n21887_27[0]),.doutb(w_n21887_27[1]),.doutc(w_n21887_27[2]),.din(w_n21887_8[2]));
	jspl3 jspl3_w_n21887_28(.douta(w_n21887_28[0]),.doutb(w_n21887_28[1]),.doutc(w_n21887_28[2]),.din(w_n21887_9[0]));
	jspl3 jspl3_w_n21887_29(.douta(w_n21887_29[0]),.doutb(w_n21887_29[1]),.doutc(w_n21887_29[2]),.din(w_n21887_9[1]));
	jspl3 jspl3_w_n21887_30(.douta(w_n21887_30[0]),.doutb(w_n21887_30[1]),.doutc(w_n21887_30[2]),.din(w_n21887_9[2]));
	jspl3 jspl3_w_n21887_31(.douta(w_n21887_31[0]),.doutb(w_n21887_31[1]),.doutc(w_n21887_31[2]),.din(w_n21887_10[0]));
	jspl3 jspl3_w_n21887_32(.douta(w_n21887_32[0]),.doutb(w_n21887_32[1]),.doutc(w_n21887_32[2]),.din(w_n21887_10[1]));
	jspl3 jspl3_w_n21887_33(.douta(w_n21887_33[0]),.doutb(w_n21887_33[1]),.doutc(w_n21887_33[2]),.din(w_n21887_10[2]));
	jspl jspl_w_n21887_34(.douta(w_n21887_34[0]),.doutb(w_n21887_34[1]),.din(w_n21887_11[0]));
	jspl3 jspl3_w_n21889_0(.douta(w_n21889_0[0]),.doutb(w_n21889_0[1]),.doutc(w_n21889_0[2]),.din(n21889));
	jspl3 jspl3_w_n21889_1(.douta(w_n21889_1[0]),.doutb(w_n21889_1[1]),.doutc(w_n21889_1[2]),.din(w_n21889_0[0]));
	jspl jspl_w_n21890_0(.douta(w_n21890_0[0]),.doutb(w_n21890_0[1]),.din(n21890));
	jspl3 jspl3_w_n21891_0(.douta(w_n21891_0[0]),.doutb(w_n21891_0[1]),.doutc(w_n21891_0[2]),.din(n21891));
	jspl jspl_w_n21892_0(.douta(w_n21892_0[0]),.doutb(w_n21892_0[1]),.din(n21892));
	jspl3 jspl3_w_n21894_0(.douta(w_n21894_0[0]),.doutb(w_n21894_0[1]),.doutc(w_n21894_0[2]),.din(n21894));
	jspl jspl_w_n21895_0(.douta(w_n21895_0[0]),.doutb(w_n21895_0[1]),.din(n21895));
	jspl3 jspl3_w_n21902_0(.douta(w_n21902_0[0]),.doutb(w_n21902_0[1]),.doutc(w_n21902_0[2]),.din(n21902));
	jspl jspl_w_n21903_0(.douta(w_n21903_0[0]),.doutb(w_n21903_0[1]),.din(n21903));
	jspl jspl_w_n21906_0(.douta(w_n21906_0[0]),.doutb(w_n21906_0[1]),.din(n21906));
	jspl jspl_w_n21909_0(.douta(w_n21909_0[0]),.doutb(w_n21909_0[1]),.din(n21909));
	jspl3 jspl3_w_n21911_0(.douta(w_n21911_0[0]),.doutb(w_n21911_0[1]),.doutc(w_n21911_0[2]),.din(n21911));
	jspl jspl_w_n21912_0(.douta(w_n21912_0[0]),.doutb(w_n21912_0[1]),.din(n21912));
	jspl3 jspl3_w_n21916_0(.douta(w_n21916_0[0]),.doutb(w_n21916_0[1]),.doutc(w_n21916_0[2]),.din(n21916));
	jspl3 jspl3_w_n21919_0(.douta(w_n21919_0[0]),.doutb(w_n21919_0[1]),.doutc(w_n21919_0[2]),.din(n21919));
	jspl jspl_w_n21920_0(.douta(w_n21920_0[0]),.doutb(w_n21920_0[1]),.din(n21920));
	jspl3 jspl3_w_n21924_0(.douta(w_n21924_0[0]),.doutb(w_n21924_0[1]),.doutc(w_n21924_0[2]),.din(n21924));
	jspl3 jspl3_w_n21926_0(.douta(w_n21926_0[0]),.doutb(w_n21926_0[1]),.doutc(w_n21926_0[2]),.din(n21926));
	jspl jspl_w_n21927_0(.douta(w_n21927_0[0]),.doutb(w_n21927_0[1]),.din(n21927));
	jspl3 jspl3_w_n21931_0(.douta(w_n21931_0[0]),.doutb(w_n21931_0[1]),.doutc(w_n21931_0[2]),.din(n21931));
	jspl3 jspl3_w_n21934_0(.douta(w_n21934_0[0]),.doutb(w_n21934_0[1]),.doutc(w_n21934_0[2]),.din(n21934));
	jspl jspl_w_n21935_0(.douta(w_n21935_0[0]),.doutb(w_n21935_0[1]),.din(n21935));
	jspl3 jspl3_w_n21939_0(.douta(w_n21939_0[0]),.doutb(w_n21939_0[1]),.doutc(w_n21939_0[2]),.din(n21939));
	jspl3 jspl3_w_n21941_0(.douta(w_n21941_0[0]),.doutb(w_n21941_0[1]),.doutc(w_n21941_0[2]),.din(n21941));
	jspl jspl_w_n21942_0(.douta(w_n21942_0[0]),.doutb(w_n21942_0[1]),.din(n21942));
	jspl3 jspl3_w_n21946_0(.douta(w_n21946_0[0]),.doutb(w_n21946_0[1]),.doutc(w_n21946_0[2]),.din(n21946));
	jspl3 jspl3_w_n21949_0(.douta(w_n21949_0[0]),.doutb(w_n21949_0[1]),.doutc(w_n21949_0[2]),.din(n21949));
	jspl jspl_w_n21950_0(.douta(w_n21950_0[0]),.doutb(w_n21950_0[1]),.din(n21950));
	jspl3 jspl3_w_n21954_0(.douta(w_n21954_0[0]),.doutb(w_n21954_0[1]),.doutc(w_n21954_0[2]),.din(n21954));
	jspl3 jspl3_w_n21956_0(.douta(w_n21956_0[0]),.doutb(w_n21956_0[1]),.doutc(w_n21956_0[2]),.din(n21956));
	jspl jspl_w_n21957_0(.douta(w_n21957_0[0]),.doutb(w_n21957_0[1]),.din(n21957));
	jspl3 jspl3_w_n21961_0(.douta(w_n21961_0[0]),.doutb(w_n21961_0[1]),.doutc(w_n21961_0[2]),.din(n21961));
	jspl3 jspl3_w_n21963_0(.douta(w_n21963_0[0]),.doutb(w_n21963_0[1]),.doutc(w_n21963_0[2]),.din(n21963));
	jspl jspl_w_n21964_0(.douta(w_n21964_0[0]),.doutb(w_n21964_0[1]),.din(n21964));
	jspl3 jspl3_w_n21968_0(.douta(w_n21968_0[0]),.doutb(w_n21968_0[1]),.doutc(w_n21968_0[2]),.din(n21968));
	jspl3 jspl3_w_n21970_0(.douta(w_n21970_0[0]),.doutb(w_n21970_0[1]),.doutc(w_n21970_0[2]),.din(n21970));
	jspl jspl_w_n21971_0(.douta(w_n21971_0[0]),.doutb(w_n21971_0[1]),.din(n21971));
	jspl3 jspl3_w_n21975_0(.douta(w_n21975_0[0]),.doutb(w_n21975_0[1]),.doutc(w_n21975_0[2]),.din(n21975));
	jspl3 jspl3_w_n21978_0(.douta(w_n21978_0[0]),.doutb(w_n21978_0[1]),.doutc(w_n21978_0[2]),.din(n21978));
	jspl jspl_w_n21979_0(.douta(w_n21979_0[0]),.doutb(w_n21979_0[1]),.din(n21979));
	jspl3 jspl3_w_n21983_0(.douta(w_n21983_0[0]),.doutb(w_n21983_0[1]),.doutc(w_n21983_0[2]),.din(n21983));
	jspl3 jspl3_w_n21985_0(.douta(w_n21985_0[0]),.doutb(w_n21985_0[1]),.doutc(w_n21985_0[2]),.din(n21985));
	jspl jspl_w_n21986_0(.douta(w_n21986_0[0]),.doutb(w_n21986_0[1]),.din(n21986));
	jspl3 jspl3_w_n21990_0(.douta(w_n21990_0[0]),.doutb(w_n21990_0[1]),.doutc(w_n21990_0[2]),.din(n21990));
	jspl3 jspl3_w_n21992_0(.douta(w_n21992_0[0]),.doutb(w_n21992_0[1]),.doutc(w_n21992_0[2]),.din(n21992));
	jspl jspl_w_n21993_0(.douta(w_n21993_0[0]),.doutb(w_n21993_0[1]),.din(n21993));
	jspl3 jspl3_w_n21997_0(.douta(w_n21997_0[0]),.doutb(w_n21997_0[1]),.doutc(w_n21997_0[2]),.din(n21997));
	jspl3 jspl3_w_n21999_0(.douta(w_n21999_0[0]),.doutb(w_n21999_0[1]),.doutc(w_n21999_0[2]),.din(n21999));
	jspl jspl_w_n22000_0(.douta(w_n22000_0[0]),.doutb(w_n22000_0[1]),.din(n22000));
	jspl3 jspl3_w_n22004_0(.douta(w_n22004_0[0]),.doutb(w_n22004_0[1]),.doutc(w_n22004_0[2]),.din(n22004));
	jspl3 jspl3_w_n22007_0(.douta(w_n22007_0[0]),.doutb(w_n22007_0[1]),.doutc(w_n22007_0[2]),.din(n22007));
	jspl jspl_w_n22008_0(.douta(w_n22008_0[0]),.doutb(w_n22008_0[1]),.din(n22008));
	jspl3 jspl3_w_n22012_0(.douta(w_n22012_0[0]),.doutb(w_n22012_0[1]),.doutc(w_n22012_0[2]),.din(n22012));
	jspl3 jspl3_w_n22014_0(.douta(w_n22014_0[0]),.doutb(w_n22014_0[1]),.doutc(w_n22014_0[2]),.din(n22014));
	jspl jspl_w_n22015_0(.douta(w_n22015_0[0]),.doutb(w_n22015_0[1]),.din(n22015));
	jspl3 jspl3_w_n22019_0(.douta(w_n22019_0[0]),.doutb(w_n22019_0[1]),.doutc(w_n22019_0[2]),.din(n22019));
	jspl3 jspl3_w_n22022_0(.douta(w_n22022_0[0]),.doutb(w_n22022_0[1]),.doutc(w_n22022_0[2]),.din(n22022));
	jspl jspl_w_n22023_0(.douta(w_n22023_0[0]),.doutb(w_n22023_0[1]),.din(n22023));
	jspl3 jspl3_w_n22027_0(.douta(w_n22027_0[0]),.doutb(w_n22027_0[1]),.doutc(w_n22027_0[2]),.din(n22027));
	jspl3 jspl3_w_n22029_0(.douta(w_n22029_0[0]),.doutb(w_n22029_0[1]),.doutc(w_n22029_0[2]),.din(n22029));
	jspl jspl_w_n22030_0(.douta(w_n22030_0[0]),.doutb(w_n22030_0[1]),.din(n22030));
	jspl3 jspl3_w_n22034_0(.douta(w_n22034_0[0]),.doutb(w_n22034_0[1]),.doutc(w_n22034_0[2]),.din(n22034));
	jspl3 jspl3_w_n22037_0(.douta(w_n22037_0[0]),.doutb(w_n22037_0[1]),.doutc(w_n22037_0[2]),.din(n22037));
	jspl jspl_w_n22038_0(.douta(w_n22038_0[0]),.doutb(w_n22038_0[1]),.din(n22038));
	jspl3 jspl3_w_n22042_0(.douta(w_n22042_0[0]),.doutb(w_n22042_0[1]),.doutc(w_n22042_0[2]),.din(n22042));
	jspl3 jspl3_w_n22044_0(.douta(w_n22044_0[0]),.doutb(w_n22044_0[1]),.doutc(w_n22044_0[2]),.din(n22044));
	jspl jspl_w_n22045_0(.douta(w_n22045_0[0]),.doutb(w_n22045_0[1]),.din(n22045));
	jspl3 jspl3_w_n22049_0(.douta(w_n22049_0[0]),.doutb(w_n22049_0[1]),.doutc(w_n22049_0[2]),.din(n22049));
	jspl3 jspl3_w_n22051_0(.douta(w_n22051_0[0]),.doutb(w_n22051_0[1]),.doutc(w_n22051_0[2]),.din(n22051));
	jspl jspl_w_n22052_0(.douta(w_n22052_0[0]),.doutb(w_n22052_0[1]),.din(n22052));
	jspl3 jspl3_w_n22056_0(.douta(w_n22056_0[0]),.doutb(w_n22056_0[1]),.doutc(w_n22056_0[2]),.din(n22056));
	jspl3 jspl3_w_n22059_0(.douta(w_n22059_0[0]),.doutb(w_n22059_0[1]),.doutc(w_n22059_0[2]),.din(n22059));
	jspl jspl_w_n22060_0(.douta(w_n22060_0[0]),.doutb(w_n22060_0[1]),.din(n22060));
	jspl3 jspl3_w_n22064_0(.douta(w_n22064_0[0]),.doutb(w_n22064_0[1]),.doutc(w_n22064_0[2]),.din(n22064));
	jspl3 jspl3_w_n22067_0(.douta(w_n22067_0[0]),.doutb(w_n22067_0[1]),.doutc(w_n22067_0[2]),.din(n22067));
	jspl jspl_w_n22068_0(.douta(w_n22068_0[0]),.doutb(w_n22068_0[1]),.din(n22068));
	jspl3 jspl3_w_n22072_0(.douta(w_n22072_0[0]),.doutb(w_n22072_0[1]),.doutc(w_n22072_0[2]),.din(n22072));
	jspl3 jspl3_w_n22074_0(.douta(w_n22074_0[0]),.doutb(w_n22074_0[1]),.doutc(w_n22074_0[2]),.din(n22074));
	jspl jspl_w_n22075_0(.douta(w_n22075_0[0]),.doutb(w_n22075_0[1]),.din(n22075));
	jspl3 jspl3_w_n22079_0(.douta(w_n22079_0[0]),.doutb(w_n22079_0[1]),.doutc(w_n22079_0[2]),.din(n22079));
	jspl3 jspl3_w_n22082_0(.douta(w_n22082_0[0]),.doutb(w_n22082_0[1]),.doutc(w_n22082_0[2]),.din(n22082));
	jspl jspl_w_n22083_0(.douta(w_n22083_0[0]),.doutb(w_n22083_0[1]),.din(n22083));
	jspl3 jspl3_w_n22087_0(.douta(w_n22087_0[0]),.doutb(w_n22087_0[1]),.doutc(w_n22087_0[2]),.din(n22087));
	jspl3 jspl3_w_n22089_0(.douta(w_n22089_0[0]),.doutb(w_n22089_0[1]),.doutc(w_n22089_0[2]),.din(n22089));
	jspl jspl_w_n22090_0(.douta(w_n22090_0[0]),.doutb(w_n22090_0[1]),.din(n22090));
	jspl3 jspl3_w_n22094_0(.douta(w_n22094_0[0]),.doutb(w_n22094_0[1]),.doutc(w_n22094_0[2]),.din(n22094));
	jspl3 jspl3_w_n22097_0(.douta(w_n22097_0[0]),.doutb(w_n22097_0[1]),.doutc(w_n22097_0[2]),.din(n22097));
	jspl jspl_w_n22098_0(.douta(w_n22098_0[0]),.doutb(w_n22098_0[1]),.din(n22098));
	jspl3 jspl3_w_n22102_0(.douta(w_n22102_0[0]),.doutb(w_n22102_0[1]),.doutc(w_n22102_0[2]),.din(n22102));
	jspl3 jspl3_w_n22104_0(.douta(w_n22104_0[0]),.doutb(w_n22104_0[1]),.doutc(w_n22104_0[2]),.din(n22104));
	jspl jspl_w_n22105_0(.douta(w_n22105_0[0]),.doutb(w_n22105_0[1]),.din(n22105));
	jspl3 jspl3_w_n22109_0(.douta(w_n22109_0[0]),.doutb(w_n22109_0[1]),.doutc(w_n22109_0[2]),.din(n22109));
	jspl3 jspl3_w_n22111_0(.douta(w_n22111_0[0]),.doutb(w_n22111_0[1]),.doutc(w_n22111_0[2]),.din(n22111));
	jspl jspl_w_n22112_0(.douta(w_n22112_0[0]),.doutb(w_n22112_0[1]),.din(n22112));
	jspl3 jspl3_w_n22116_0(.douta(w_n22116_0[0]),.doutb(w_n22116_0[1]),.doutc(w_n22116_0[2]),.din(n22116));
	jspl3 jspl3_w_n22118_0(.douta(w_n22118_0[0]),.doutb(w_n22118_0[1]),.doutc(w_n22118_0[2]),.din(n22118));
	jspl jspl_w_n22119_0(.douta(w_n22119_0[0]),.doutb(w_n22119_0[1]),.din(n22119));
	jspl3 jspl3_w_n22123_0(.douta(w_n22123_0[0]),.doutb(w_n22123_0[1]),.doutc(w_n22123_0[2]),.din(n22123));
	jspl3 jspl3_w_n22126_0(.douta(w_n22126_0[0]),.doutb(w_n22126_0[1]),.doutc(w_n22126_0[2]),.din(n22126));
	jspl jspl_w_n22127_0(.douta(w_n22127_0[0]),.doutb(w_n22127_0[1]),.din(n22127));
	jspl3 jspl3_w_n22131_0(.douta(w_n22131_0[0]),.doutb(w_n22131_0[1]),.doutc(w_n22131_0[2]),.din(n22131));
	jspl3 jspl3_w_n22133_0(.douta(w_n22133_0[0]),.doutb(w_n22133_0[1]),.doutc(w_n22133_0[2]),.din(n22133));
	jspl jspl_w_n22134_0(.douta(w_n22134_0[0]),.doutb(w_n22134_0[1]),.din(n22134));
	jspl3 jspl3_w_n22138_0(.douta(w_n22138_0[0]),.doutb(w_n22138_0[1]),.doutc(w_n22138_0[2]),.din(n22138));
	jspl3 jspl3_w_n22141_0(.douta(w_n22141_0[0]),.doutb(w_n22141_0[1]),.doutc(w_n22141_0[2]),.din(n22141));
	jspl jspl_w_n22142_0(.douta(w_n22142_0[0]),.doutb(w_n22142_0[1]),.din(n22142));
	jspl3 jspl3_w_n22146_0(.douta(w_n22146_0[0]),.doutb(w_n22146_0[1]),.doutc(w_n22146_0[2]),.din(n22146));
	jspl3 jspl3_w_n22148_0(.douta(w_n22148_0[0]),.doutb(w_n22148_0[1]),.doutc(w_n22148_0[2]),.din(n22148));
	jspl jspl_w_n22149_0(.douta(w_n22149_0[0]),.doutb(w_n22149_0[1]),.din(n22149));
	jspl3 jspl3_w_n22153_0(.douta(w_n22153_0[0]),.doutb(w_n22153_0[1]),.doutc(w_n22153_0[2]),.din(n22153));
	jspl3 jspl3_w_n22156_0(.douta(w_n22156_0[0]),.doutb(w_n22156_0[1]),.doutc(w_n22156_0[2]),.din(n22156));
	jspl jspl_w_n22157_0(.douta(w_n22157_0[0]),.doutb(w_n22157_0[1]),.din(n22157));
	jspl3 jspl3_w_n22161_0(.douta(w_n22161_0[0]),.doutb(w_n22161_0[1]),.doutc(w_n22161_0[2]),.din(n22161));
	jspl3 jspl3_w_n22163_0(.douta(w_n22163_0[0]),.doutb(w_n22163_0[1]),.doutc(w_n22163_0[2]),.din(n22163));
	jspl jspl_w_n22164_0(.douta(w_n22164_0[0]),.doutb(w_n22164_0[1]),.din(n22164));
	jspl3 jspl3_w_n22168_0(.douta(w_n22168_0[0]),.doutb(w_n22168_0[1]),.doutc(w_n22168_0[2]),.din(n22168));
	jspl3 jspl3_w_n22171_0(.douta(w_n22171_0[0]),.doutb(w_n22171_0[1]),.doutc(w_n22171_0[2]),.din(n22171));
	jspl jspl_w_n22172_0(.douta(w_n22172_0[0]),.doutb(w_n22172_0[1]),.din(n22172));
	jspl3 jspl3_w_n22176_0(.douta(w_n22176_0[0]),.doutb(w_n22176_0[1]),.doutc(w_n22176_0[2]),.din(n22176));
	jspl3 jspl3_w_n22178_0(.douta(w_n22178_0[0]),.doutb(w_n22178_0[1]),.doutc(w_n22178_0[2]),.din(n22178));
	jspl jspl_w_n22179_0(.douta(w_n22179_0[0]),.doutb(w_n22179_0[1]),.din(n22179));
	jspl3 jspl3_w_n22183_0(.douta(w_n22183_0[0]),.doutb(w_n22183_0[1]),.doutc(w_n22183_0[2]),.din(n22183));
	jspl3 jspl3_w_n22185_0(.douta(w_n22185_0[0]),.doutb(w_n22185_0[1]),.doutc(w_n22185_0[2]),.din(n22185));
	jspl jspl_w_n22186_0(.douta(w_n22186_0[0]),.doutb(w_n22186_0[1]),.din(n22186));
	jspl3 jspl3_w_n22190_0(.douta(w_n22190_0[0]),.doutb(w_n22190_0[1]),.doutc(w_n22190_0[2]),.din(n22190));
	jspl3 jspl3_w_n22192_0(.douta(w_n22192_0[0]),.doutb(w_n22192_0[1]),.doutc(w_n22192_0[2]),.din(n22192));
	jspl jspl_w_n22193_0(.douta(w_n22193_0[0]),.doutb(w_n22193_0[1]),.din(n22193));
	jspl3 jspl3_w_n22197_0(.douta(w_n22197_0[0]),.doutb(w_n22197_0[1]),.doutc(w_n22197_0[2]),.din(n22197));
	jspl3 jspl3_w_n22200_0(.douta(w_n22200_0[0]),.doutb(w_n22200_0[1]),.doutc(w_n22200_0[2]),.din(n22200));
	jspl jspl_w_n22201_0(.douta(w_n22201_0[0]),.doutb(w_n22201_0[1]),.din(n22201));
	jspl3 jspl3_w_n22205_0(.douta(w_n22205_0[0]),.doutb(w_n22205_0[1]),.doutc(w_n22205_0[2]),.din(n22205));
	jspl3 jspl3_w_n22207_0(.douta(w_n22207_0[0]),.doutb(w_n22207_0[1]),.doutc(w_n22207_0[2]),.din(n22207));
	jspl jspl_w_n22208_0(.douta(w_n22208_0[0]),.doutb(w_n22208_0[1]),.din(n22208));
	jspl3 jspl3_w_n22212_0(.douta(w_n22212_0[0]),.doutb(w_n22212_0[1]),.doutc(w_n22212_0[2]),.din(n22212));
	jspl3 jspl3_w_n22214_0(.douta(w_n22214_0[0]),.doutb(w_n22214_0[1]),.doutc(w_n22214_0[2]),.din(n22214));
	jspl jspl_w_n22215_0(.douta(w_n22215_0[0]),.doutb(w_n22215_0[1]),.din(n22215));
	jspl3 jspl3_w_n22219_0(.douta(w_n22219_0[0]),.doutb(w_n22219_0[1]),.doutc(w_n22219_0[2]),.din(n22219));
	jspl3 jspl3_w_n22221_0(.douta(w_n22221_0[0]),.doutb(w_n22221_0[1]),.doutc(w_n22221_0[2]),.din(n22221));
	jspl jspl_w_n22222_0(.douta(w_n22222_0[0]),.doutb(w_n22222_0[1]),.din(n22222));
	jspl3 jspl3_w_n22226_0(.douta(w_n22226_0[0]),.doutb(w_n22226_0[1]),.doutc(w_n22226_0[2]),.din(n22226));
	jspl3 jspl3_w_n22228_0(.douta(w_n22228_0[0]),.doutb(w_n22228_0[1]),.doutc(w_n22228_0[2]),.din(n22228));
	jspl jspl_w_n22229_0(.douta(w_n22229_0[0]),.doutb(w_n22229_0[1]),.din(n22229));
	jspl3 jspl3_w_n22233_0(.douta(w_n22233_0[0]),.doutb(w_n22233_0[1]),.doutc(w_n22233_0[2]),.din(n22233));
	jspl3 jspl3_w_n22235_0(.douta(w_n22235_0[0]),.doutb(w_n22235_0[1]),.doutc(w_n22235_0[2]),.din(n22235));
	jspl jspl_w_n22236_0(.douta(w_n22236_0[0]),.doutb(w_n22236_0[1]),.din(n22236));
	jspl3 jspl3_w_n22240_0(.douta(w_n22240_0[0]),.doutb(w_n22240_0[1]),.doutc(w_n22240_0[2]),.din(n22240));
	jspl3 jspl3_w_n22243_0(.douta(w_n22243_0[0]),.doutb(w_n22243_0[1]),.doutc(w_n22243_0[2]),.din(n22243));
	jspl jspl_w_n22244_0(.douta(w_n22244_0[0]),.doutb(w_n22244_0[1]),.din(n22244));
	jspl3 jspl3_w_n22248_0(.douta(w_n22248_0[0]),.doutb(w_n22248_0[1]),.doutc(w_n22248_0[2]),.din(n22248));
	jspl3 jspl3_w_n22250_0(.douta(w_n22250_0[0]),.doutb(w_n22250_0[1]),.doutc(w_n22250_0[2]),.din(n22250));
	jspl jspl_w_n22251_0(.douta(w_n22251_0[0]),.doutb(w_n22251_0[1]),.din(n22251));
	jspl3 jspl3_w_n22255_0(.douta(w_n22255_0[0]),.doutb(w_n22255_0[1]),.doutc(w_n22255_0[2]),.din(n22255));
	jspl3 jspl3_w_n22258_0(.douta(w_n22258_0[0]),.doutb(w_n22258_0[1]),.doutc(w_n22258_0[2]),.din(n22258));
	jspl jspl_w_n22259_0(.douta(w_n22259_0[0]),.doutb(w_n22259_0[1]),.din(n22259));
	jspl3 jspl3_w_n22263_0(.douta(w_n22263_0[0]),.doutb(w_n22263_0[1]),.doutc(w_n22263_0[2]),.din(n22263));
	jspl3 jspl3_w_n22265_0(.douta(w_n22265_0[0]),.doutb(w_n22265_0[1]),.doutc(w_n22265_0[2]),.din(n22265));
	jspl jspl_w_n22266_0(.douta(w_n22266_0[0]),.doutb(w_n22266_0[1]),.din(n22266));
	jspl3 jspl3_w_n22270_0(.douta(w_n22270_0[0]),.doutb(w_n22270_0[1]),.doutc(w_n22270_0[2]),.din(n22270));
	jspl3 jspl3_w_n22272_0(.douta(w_n22272_0[0]),.doutb(w_n22272_0[1]),.doutc(w_n22272_0[2]),.din(n22272));
	jspl jspl_w_n22273_0(.douta(w_n22273_0[0]),.doutb(w_n22273_0[1]),.din(n22273));
	jspl3 jspl3_w_n22277_0(.douta(w_n22277_0[0]),.doutb(w_n22277_0[1]),.doutc(w_n22277_0[2]),.din(n22277));
	jspl3 jspl3_w_n22280_0(.douta(w_n22280_0[0]),.doutb(w_n22280_0[1]),.doutc(w_n22280_0[2]),.din(n22280));
	jspl jspl_w_n22281_0(.douta(w_n22281_0[0]),.doutb(w_n22281_0[1]),.din(n22281));
	jspl3 jspl3_w_n22285_0(.douta(w_n22285_0[0]),.doutb(w_n22285_0[1]),.doutc(w_n22285_0[2]),.din(n22285));
	jspl3 jspl3_w_n22288_0(.douta(w_n22288_0[0]),.doutb(w_n22288_0[1]),.doutc(w_n22288_0[2]),.din(n22288));
	jspl jspl_w_n22289_0(.douta(w_n22289_0[0]),.doutb(w_n22289_0[1]),.din(n22289));
	jspl3 jspl3_w_n22293_0(.douta(w_n22293_0[0]),.doutb(w_n22293_0[1]),.doutc(w_n22293_0[2]),.din(n22293));
	jspl3 jspl3_w_n22295_0(.douta(w_n22295_0[0]),.doutb(w_n22295_0[1]),.doutc(w_n22295_0[2]),.din(n22295));
	jspl jspl_w_n22296_0(.douta(w_n22296_0[0]),.doutb(w_n22296_0[1]),.din(n22296));
	jspl3 jspl3_w_n22300_0(.douta(w_n22300_0[0]),.doutb(w_n22300_0[1]),.doutc(w_n22300_0[2]),.din(n22300));
	jspl3 jspl3_w_n22302_0(.douta(w_n22302_0[0]),.doutb(w_n22302_0[1]),.doutc(w_n22302_0[2]),.din(n22302));
	jspl jspl_w_n22303_0(.douta(w_n22303_0[0]),.doutb(w_n22303_0[1]),.din(n22303));
	jspl3 jspl3_w_n22307_0(.douta(w_n22307_0[0]),.doutb(w_n22307_0[1]),.doutc(w_n22307_0[2]),.din(n22307));
	jspl3 jspl3_w_n22309_0(.douta(w_n22309_0[0]),.doutb(w_n22309_0[1]),.doutc(w_n22309_0[2]),.din(n22309));
	jspl jspl_w_n22310_0(.douta(w_n22310_0[0]),.doutb(w_n22310_0[1]),.din(n22310));
	jspl jspl_w_n22314_0(.douta(w_n22314_0[0]),.doutb(w_n22314_0[1]),.din(n22314));
	jspl jspl_w_n22315_0(.douta(w_n22315_0[0]),.doutb(w_n22315_0[1]),.din(n22315));
	jspl3 jspl3_w_n22317_0(.douta(w_n22317_0[0]),.doutb(w_n22317_0[1]),.doutc(w_n22317_0[2]),.din(n22317));
	jspl jspl_w_n22317_1(.douta(w_n22317_1[0]),.doutb(w_n22317_1[1]),.din(w_n22317_0[0]));
	jspl3 jspl3_w_n22320_0(.douta(w_n22320_0[0]),.doutb(w_n22320_0[1]),.doutc(w_n22320_0[2]),.din(n22320));
	jspl jspl_w_n22320_1(.douta(w_n22320_1[0]),.doutb(w_n22320_1[1]),.din(w_n22320_0[0]));
	jspl3 jspl3_w_n22321_0(.douta(w_n22321_0[0]),.doutb(w_n22321_0[1]),.doutc(w_n22321_0[2]),.din(n22321));
	jspl jspl_w_n22324_0(.douta(w_n22324_0[0]),.doutb(w_n22324_0[1]),.din(n22324));
	jspl jspl_w_n22325_0(.douta(w_n22325_0[0]),.doutb(w_n22325_0[1]),.din(n22325));
	jspl jspl_w_n22330_0(.douta(w_n22330_0[0]),.doutb(w_n22330_0[1]),.din(n22330));
	jspl jspl_w_n22332_0(.douta(w_n22332_0[0]),.doutb(w_n22332_0[1]),.din(n22332));
	jspl3 jspl3_w_n22334_0(.douta(w_n22334_0[0]),.doutb(w_n22334_0[1]),.doutc(w_n22334_0[2]),.din(n22334));
	jspl3 jspl3_w_n22334_1(.douta(w_n22334_1[0]),.doutb(w_n22334_1[1]),.doutc(w_n22334_1[2]),.din(w_n22334_0[0]));
	jspl jspl_w_n22335_0(.douta(w_n22335_0[0]),.doutb(w_n22335_0[1]),.din(n22335));
	jspl3 jspl3_w_n22336_0(.douta(w_n22336_0[0]),.doutb(w_n22336_0[1]),.doutc(w_n22336_0[2]),.din(n22336));
	jspl jspl_w_n22337_0(.douta(w_n22337_0[0]),.doutb(w_n22337_0[1]),.din(n22337));
	jspl3 jspl3_w_n22339_0(.douta(w_n22339_0[0]),.doutb(w_n22339_0[1]),.doutc(w_n22339_0[2]),.din(n22339));
	jspl jspl_w_n22340_0(.douta(w_n22340_0[0]),.doutb(w_n22340_0[1]),.din(n22340));
	jspl jspl_w_n22345_0(.douta(w_n22345_0[0]),.doutb(w_n22345_0[1]),.din(n22345));
	jspl jspl_w_n22408_0(.douta(w_n22408_0[0]),.doutb(w_n22408_0[1]),.din(n22408));
	jspl jspl_w_n22412_0(.douta(w_n22412_0[0]),.doutb(w_n22412_0[1]),.din(n22412));
	jspl jspl_w_n22615_0(.douta(w_n22615_0[0]),.doutb(w_n22615_0[1]),.din(n22615));
	jspl jspl_w_n22619_0(.douta(w_n22619_0[0]),.doutb(w_n22619_0[1]),.din(n22619));
	jspl3 jspl3_w_n22620_0(.douta(w_n22620_0[0]),.doutb(w_n22620_0[1]),.doutc(w_n22620_0[2]),.din(n22620));
	jspl3 jspl3_w_n22620_1(.douta(w_n22620_1[0]),.doutb(w_n22620_1[1]),.doutc(w_n22620_1[2]),.din(w_n22620_0[0]));
	jspl3 jspl3_w_n22620_2(.douta(w_n22620_2[0]),.doutb(w_n22620_2[1]),.doutc(w_n22620_2[2]),.din(w_n22620_0[1]));
	jspl3 jspl3_w_n22620_3(.douta(w_n22620_3[0]),.doutb(w_n22620_3[1]),.doutc(w_n22620_3[2]),.din(w_n22620_0[2]));
	jspl3 jspl3_w_n22620_4(.douta(w_n22620_4[0]),.doutb(w_n22620_4[1]),.doutc(w_n22620_4[2]),.din(w_n22620_1[0]));
	jspl jspl_w_n22621_0(.douta(w_n22621_0[0]),.doutb(w_n22621_0[1]),.din(n22621));
	jspl jspl_w_n22622_0(.douta(w_n22622_0[0]),.doutb(w_n22622_0[1]),.din(n22622));
	jspl3 jspl3_w_n22624_0(.douta(w_n22624_0[0]),.doutb(w_n22624_0[1]),.doutc(w_n22624_0[2]),.din(n22624));
	jspl jspl_w_n22625_0(.douta(w_n22625_0[0]),.doutb(w_n22625_0[1]),.din(n22625));
	jspl jspl_w_n22629_0(.douta(w_n22629_0[0]),.doutb(w_n22629_0[1]),.din(n22629));
	jspl jspl_w_n22630_0(.douta(w_n22630_0[0]),.doutb(w_n22630_0[1]),.din(n22630));
	jspl3 jspl3_w_n22632_0(.douta(w_n22632_0[0]),.doutb(w_n22632_0[1]),.doutc(w_n22632_0[2]),.din(n22632));
	jspl jspl_w_n22633_0(.douta(w_n22633_0[0]),.doutb(w_n22633_0[1]),.din(n22633));
	jspl jspl_w_n22637_0(.douta(w_n22637_0[0]),.doutb(w_n22637_0[1]),.din(n22637));
	jspl3 jspl3_w_n22639_0(.douta(w_n22639_0[0]),.doutb(w_n22639_0[1]),.doutc(w_n22639_0[2]),.din(n22639));
	jspl jspl_w_n22640_0(.douta(w_n22640_0[0]),.doutb(w_n22640_0[1]),.din(n22640));
	jspl jspl_w_n22644_0(.douta(w_n22644_0[0]),.doutb(w_n22644_0[1]),.din(n22644));
	jspl3 jspl3_w_n22646_0(.douta(w_n22646_0[0]),.doutb(w_n22646_0[1]),.doutc(w_n22646_0[2]),.din(n22646));
	jspl jspl_w_n22647_0(.douta(w_n22647_0[0]),.doutb(w_n22647_0[1]),.din(n22647));
	jspl jspl_w_n22651_0(.douta(w_n22651_0[0]),.doutb(w_n22651_0[1]),.din(n22651));
	jspl3 jspl3_w_n22653_0(.douta(w_n22653_0[0]),.doutb(w_n22653_0[1]),.doutc(w_n22653_0[2]),.din(n22653));
	jspl jspl_w_n22654_0(.douta(w_n22654_0[0]),.doutb(w_n22654_0[1]),.din(n22654));
	jspl jspl_w_n22658_0(.douta(w_n22658_0[0]),.doutb(w_n22658_0[1]),.din(n22658));
	jspl jspl_w_n22659_0(.douta(w_n22659_0[0]),.doutb(w_n22659_0[1]),.din(n22659));
	jspl3 jspl3_w_n22661_0(.douta(w_n22661_0[0]),.doutb(w_n22661_0[1]),.doutc(w_n22661_0[2]),.din(n22661));
	jspl jspl_w_n22662_0(.douta(w_n22662_0[0]),.doutb(w_n22662_0[1]),.din(n22662));
	jspl jspl_w_n22666_0(.douta(w_n22666_0[0]),.doutb(w_n22666_0[1]),.din(n22666));
	jspl3 jspl3_w_n22668_0(.douta(w_n22668_0[0]),.doutb(w_n22668_0[1]),.doutc(w_n22668_0[2]),.din(n22668));
	jspl jspl_w_n22669_0(.douta(w_n22669_0[0]),.doutb(w_n22669_0[1]),.din(n22669));
	jspl jspl_w_n22673_0(.douta(w_n22673_0[0]),.doutb(w_n22673_0[1]),.din(n22673));
	jspl jspl_w_n22674_0(.douta(w_n22674_0[0]),.doutb(w_n22674_0[1]),.din(n22674));
	jspl3 jspl3_w_n22676_0(.douta(w_n22676_0[0]),.doutb(w_n22676_0[1]),.doutc(w_n22676_0[2]),.din(n22676));
	jspl jspl_w_n22677_0(.douta(w_n22677_0[0]),.doutb(w_n22677_0[1]),.din(n22677));
	jspl jspl_w_n22681_0(.douta(w_n22681_0[0]),.doutb(w_n22681_0[1]),.din(n22681));
	jspl3 jspl3_w_n22683_0(.douta(w_n22683_0[0]),.doutb(w_n22683_0[1]),.doutc(w_n22683_0[2]),.din(n22683));
	jspl jspl_w_n22684_0(.douta(w_n22684_0[0]),.doutb(w_n22684_0[1]),.din(n22684));
	jspl jspl_w_n22688_0(.douta(w_n22688_0[0]),.doutb(w_n22688_0[1]),.din(n22688));
	jspl jspl_w_n22689_0(.douta(w_n22689_0[0]),.doutb(w_n22689_0[1]),.din(n22689));
	jspl3 jspl3_w_n22691_0(.douta(w_n22691_0[0]),.doutb(w_n22691_0[1]),.doutc(w_n22691_0[2]),.din(n22691));
	jspl jspl_w_n22692_0(.douta(w_n22692_0[0]),.doutb(w_n22692_0[1]),.din(n22692));
	jspl jspl_w_n22696_0(.douta(w_n22696_0[0]),.doutb(w_n22696_0[1]),.din(n22696));
	jspl jspl_w_n22697_0(.douta(w_n22697_0[0]),.doutb(w_n22697_0[1]),.din(n22697));
	jspl3 jspl3_w_n22699_0(.douta(w_n22699_0[0]),.doutb(w_n22699_0[1]),.doutc(w_n22699_0[2]),.din(n22699));
	jspl jspl_w_n22700_0(.douta(w_n22700_0[0]),.doutb(w_n22700_0[1]),.din(n22700));
	jspl jspl_w_n22704_0(.douta(w_n22704_0[0]),.doutb(w_n22704_0[1]),.din(n22704));
	jspl jspl_w_n22705_0(.douta(w_n22705_0[0]),.doutb(w_n22705_0[1]),.din(n22705));
	jspl3 jspl3_w_n22707_0(.douta(w_n22707_0[0]),.doutb(w_n22707_0[1]),.doutc(w_n22707_0[2]),.din(n22707));
	jspl jspl_w_n22708_0(.douta(w_n22708_0[0]),.doutb(w_n22708_0[1]),.din(n22708));
	jspl jspl_w_n22712_0(.douta(w_n22712_0[0]),.doutb(w_n22712_0[1]),.din(n22712));
	jspl3 jspl3_w_n22714_0(.douta(w_n22714_0[0]),.doutb(w_n22714_0[1]),.doutc(w_n22714_0[2]),.din(n22714));
	jspl jspl_w_n22715_0(.douta(w_n22715_0[0]),.doutb(w_n22715_0[1]),.din(n22715));
	jspl jspl_w_n22719_0(.douta(w_n22719_0[0]),.doutb(w_n22719_0[1]),.din(n22719));
	jspl jspl_w_n22720_0(.douta(w_n22720_0[0]),.doutb(w_n22720_0[1]),.din(n22720));
	jspl3 jspl3_w_n22722_0(.douta(w_n22722_0[0]),.doutb(w_n22722_0[1]),.doutc(w_n22722_0[2]),.din(n22722));
	jspl jspl_w_n22723_0(.douta(w_n22723_0[0]),.doutb(w_n22723_0[1]),.din(n22723));
	jspl jspl_w_n22727_0(.douta(w_n22727_0[0]),.doutb(w_n22727_0[1]),.din(n22727));
	jspl jspl_w_n22728_0(.douta(w_n22728_0[0]),.doutb(w_n22728_0[1]),.din(n22728));
	jspl3 jspl3_w_n22730_0(.douta(w_n22730_0[0]),.doutb(w_n22730_0[1]),.doutc(w_n22730_0[2]),.din(n22730));
	jspl jspl_w_n22731_0(.douta(w_n22731_0[0]),.doutb(w_n22731_0[1]),.din(n22731));
	jspl jspl_w_n22735_0(.douta(w_n22735_0[0]),.doutb(w_n22735_0[1]),.din(n22735));
	jspl jspl_w_n22736_0(.douta(w_n22736_0[0]),.doutb(w_n22736_0[1]),.din(n22736));
	jspl3 jspl3_w_n22738_0(.douta(w_n22738_0[0]),.doutb(w_n22738_0[1]),.doutc(w_n22738_0[2]),.din(n22738));
	jspl jspl_w_n22739_0(.douta(w_n22739_0[0]),.doutb(w_n22739_0[1]),.din(n22739));
	jspl jspl_w_n22743_0(.douta(w_n22743_0[0]),.doutb(w_n22743_0[1]),.din(n22743));
	jspl3 jspl3_w_n22745_0(.douta(w_n22745_0[0]),.doutb(w_n22745_0[1]),.doutc(w_n22745_0[2]),.din(n22745));
	jspl jspl_w_n22746_0(.douta(w_n22746_0[0]),.doutb(w_n22746_0[1]),.din(n22746));
	jspl jspl_w_n22750_0(.douta(w_n22750_0[0]),.doutb(w_n22750_0[1]),.din(n22750));
	jspl jspl_w_n22751_0(.douta(w_n22751_0[0]),.doutb(w_n22751_0[1]),.din(n22751));
	jspl3 jspl3_w_n22753_0(.douta(w_n22753_0[0]),.doutb(w_n22753_0[1]),.doutc(w_n22753_0[2]),.din(n22753));
	jspl jspl_w_n22754_0(.douta(w_n22754_0[0]),.doutb(w_n22754_0[1]),.din(n22754));
	jspl jspl_w_n22758_0(.douta(w_n22758_0[0]),.doutb(w_n22758_0[1]),.din(n22758));
	jspl3 jspl3_w_n22760_0(.douta(w_n22760_0[0]),.doutb(w_n22760_0[1]),.doutc(w_n22760_0[2]),.din(n22760));
	jspl jspl_w_n22761_0(.douta(w_n22761_0[0]),.doutb(w_n22761_0[1]),.din(n22761));
	jspl jspl_w_n22765_0(.douta(w_n22765_0[0]),.doutb(w_n22765_0[1]),.din(n22765));
	jspl jspl_w_n22766_0(.douta(w_n22766_0[0]),.doutb(w_n22766_0[1]),.din(n22766));
	jspl3 jspl3_w_n22768_0(.douta(w_n22768_0[0]),.doutb(w_n22768_0[1]),.doutc(w_n22768_0[2]),.din(n22768));
	jspl jspl_w_n22769_0(.douta(w_n22769_0[0]),.doutb(w_n22769_0[1]),.din(n22769));
	jspl jspl_w_n22773_0(.douta(w_n22773_0[0]),.doutb(w_n22773_0[1]),.din(n22773));
	jspl3 jspl3_w_n22775_0(.douta(w_n22775_0[0]),.doutb(w_n22775_0[1]),.doutc(w_n22775_0[2]),.din(n22775));
	jspl jspl_w_n22776_0(.douta(w_n22776_0[0]),.doutb(w_n22776_0[1]),.din(n22776));
	jspl jspl_w_n22780_0(.douta(w_n22780_0[0]),.doutb(w_n22780_0[1]),.din(n22780));
	jspl jspl_w_n22781_0(.douta(w_n22781_0[0]),.doutb(w_n22781_0[1]),.din(n22781));
	jspl3 jspl3_w_n22783_0(.douta(w_n22783_0[0]),.doutb(w_n22783_0[1]),.doutc(w_n22783_0[2]),.din(n22783));
	jspl jspl_w_n22784_0(.douta(w_n22784_0[0]),.doutb(w_n22784_0[1]),.din(n22784));
	jspl jspl_w_n22788_0(.douta(w_n22788_0[0]),.doutb(w_n22788_0[1]),.din(n22788));
	jspl jspl_w_n22789_0(.douta(w_n22789_0[0]),.doutb(w_n22789_0[1]),.din(n22789));
	jspl3 jspl3_w_n22791_0(.douta(w_n22791_0[0]),.doutb(w_n22791_0[1]),.doutc(w_n22791_0[2]),.din(n22791));
	jspl jspl_w_n22792_0(.douta(w_n22792_0[0]),.doutb(w_n22792_0[1]),.din(n22792));
	jspl jspl_w_n22796_0(.douta(w_n22796_0[0]),.doutb(w_n22796_0[1]),.din(n22796));
	jspl3 jspl3_w_n22798_0(.douta(w_n22798_0[0]),.doutb(w_n22798_0[1]),.doutc(w_n22798_0[2]),.din(n22798));
	jspl jspl_w_n22799_0(.douta(w_n22799_0[0]),.doutb(w_n22799_0[1]),.din(n22799));
	jspl jspl_w_n22803_0(.douta(w_n22803_0[0]),.doutb(w_n22803_0[1]),.din(n22803));
	jspl3 jspl3_w_n22805_0(.douta(w_n22805_0[0]),.doutb(w_n22805_0[1]),.doutc(w_n22805_0[2]),.din(n22805));
	jspl jspl_w_n22806_0(.douta(w_n22806_0[0]),.doutb(w_n22806_0[1]),.din(n22806));
	jspl jspl_w_n22810_0(.douta(w_n22810_0[0]),.doutb(w_n22810_0[1]),.din(n22810));
	jspl jspl_w_n22811_0(.douta(w_n22811_0[0]),.doutb(w_n22811_0[1]),.din(n22811));
	jspl3 jspl3_w_n22813_0(.douta(w_n22813_0[0]),.doutb(w_n22813_0[1]),.doutc(w_n22813_0[2]),.din(n22813));
	jspl jspl_w_n22814_0(.douta(w_n22814_0[0]),.doutb(w_n22814_0[1]),.din(n22814));
	jspl jspl_w_n22818_0(.douta(w_n22818_0[0]),.doutb(w_n22818_0[1]),.din(n22818));
	jspl3 jspl3_w_n22820_0(.douta(w_n22820_0[0]),.doutb(w_n22820_0[1]),.doutc(w_n22820_0[2]),.din(n22820));
	jspl jspl_w_n22821_0(.douta(w_n22821_0[0]),.doutb(w_n22821_0[1]),.din(n22821));
	jspl jspl_w_n22825_0(.douta(w_n22825_0[0]),.doutb(w_n22825_0[1]),.din(n22825));
	jspl jspl_w_n22826_0(.douta(w_n22826_0[0]),.doutb(w_n22826_0[1]),.din(n22826));
	jspl3 jspl3_w_n22828_0(.douta(w_n22828_0[0]),.doutb(w_n22828_0[1]),.doutc(w_n22828_0[2]),.din(n22828));
	jspl jspl_w_n22829_0(.douta(w_n22829_0[0]),.doutb(w_n22829_0[1]),.din(n22829));
	jspl jspl_w_n22833_0(.douta(w_n22833_0[0]),.doutb(w_n22833_0[1]),.din(n22833));
	jspl3 jspl3_w_n22835_0(.douta(w_n22835_0[0]),.doutb(w_n22835_0[1]),.doutc(w_n22835_0[2]),.din(n22835));
	jspl jspl_w_n22836_0(.douta(w_n22836_0[0]),.doutb(w_n22836_0[1]),.din(n22836));
	jspl jspl_w_n22840_0(.douta(w_n22840_0[0]),.doutb(w_n22840_0[1]),.din(n22840));
	jspl jspl_w_n22841_0(.douta(w_n22841_0[0]),.doutb(w_n22841_0[1]),.din(n22841));
	jspl3 jspl3_w_n22843_0(.douta(w_n22843_0[0]),.doutb(w_n22843_0[1]),.doutc(w_n22843_0[2]),.din(n22843));
	jspl jspl_w_n22844_0(.douta(w_n22844_0[0]),.doutb(w_n22844_0[1]),.din(n22844));
	jspl jspl_w_n22848_0(.douta(w_n22848_0[0]),.doutb(w_n22848_0[1]),.din(n22848));
	jspl jspl_w_n22849_0(.douta(w_n22849_0[0]),.doutb(w_n22849_0[1]),.din(n22849));
	jspl3 jspl3_w_n22851_0(.douta(w_n22851_0[0]),.doutb(w_n22851_0[1]),.doutc(w_n22851_0[2]),.din(n22851));
	jspl jspl_w_n22852_0(.douta(w_n22852_0[0]),.doutb(w_n22852_0[1]),.din(n22852));
	jspl jspl_w_n22856_0(.douta(w_n22856_0[0]),.doutb(w_n22856_0[1]),.din(n22856));
	jspl jspl_w_n22857_0(.douta(w_n22857_0[0]),.doutb(w_n22857_0[1]),.din(n22857));
	jspl3 jspl3_w_n22859_0(.douta(w_n22859_0[0]),.doutb(w_n22859_0[1]),.doutc(w_n22859_0[2]),.din(n22859));
	jspl jspl_w_n22860_0(.douta(w_n22860_0[0]),.doutb(w_n22860_0[1]),.din(n22860));
	jspl jspl_w_n22864_0(.douta(w_n22864_0[0]),.doutb(w_n22864_0[1]),.din(n22864));
	jspl3 jspl3_w_n22866_0(.douta(w_n22866_0[0]),.doutb(w_n22866_0[1]),.doutc(w_n22866_0[2]),.din(n22866));
	jspl jspl_w_n22867_0(.douta(w_n22867_0[0]),.doutb(w_n22867_0[1]),.din(n22867));
	jspl jspl_w_n22871_0(.douta(w_n22871_0[0]),.doutb(w_n22871_0[1]),.din(n22871));
	jspl jspl_w_n22872_0(.douta(w_n22872_0[0]),.doutb(w_n22872_0[1]),.din(n22872));
	jspl3 jspl3_w_n22874_0(.douta(w_n22874_0[0]),.doutb(w_n22874_0[1]),.doutc(w_n22874_0[2]),.din(n22874));
	jspl jspl_w_n22875_0(.douta(w_n22875_0[0]),.doutb(w_n22875_0[1]),.din(n22875));
	jspl jspl_w_n22879_0(.douta(w_n22879_0[0]),.doutb(w_n22879_0[1]),.din(n22879));
	jspl3 jspl3_w_n22881_0(.douta(w_n22881_0[0]),.doutb(w_n22881_0[1]),.doutc(w_n22881_0[2]),.din(n22881));
	jspl jspl_w_n22882_0(.douta(w_n22882_0[0]),.doutb(w_n22882_0[1]),.din(n22882));
	jspl jspl_w_n22886_0(.douta(w_n22886_0[0]),.doutb(w_n22886_0[1]),.din(n22886));
	jspl jspl_w_n22887_0(.douta(w_n22887_0[0]),.doutb(w_n22887_0[1]),.din(n22887));
	jspl3 jspl3_w_n22889_0(.douta(w_n22889_0[0]),.doutb(w_n22889_0[1]),.doutc(w_n22889_0[2]),.din(n22889));
	jspl jspl_w_n22890_0(.douta(w_n22890_0[0]),.doutb(w_n22890_0[1]),.din(n22890));
	jspl jspl_w_n22894_0(.douta(w_n22894_0[0]),.doutb(w_n22894_0[1]),.din(n22894));
	jspl3 jspl3_w_n22896_0(.douta(w_n22896_0[0]),.doutb(w_n22896_0[1]),.doutc(w_n22896_0[2]),.din(n22896));
	jspl jspl_w_n22897_0(.douta(w_n22897_0[0]),.doutb(w_n22897_0[1]),.din(n22897));
	jspl jspl_w_n22901_0(.douta(w_n22901_0[0]),.doutb(w_n22901_0[1]),.din(n22901));
	jspl jspl_w_n22902_0(.douta(w_n22902_0[0]),.doutb(w_n22902_0[1]),.din(n22902));
	jspl3 jspl3_w_n22904_0(.douta(w_n22904_0[0]),.doutb(w_n22904_0[1]),.doutc(w_n22904_0[2]),.din(n22904));
	jspl jspl_w_n22905_0(.douta(w_n22905_0[0]),.doutb(w_n22905_0[1]),.din(n22905));
	jspl jspl_w_n22909_0(.douta(w_n22909_0[0]),.doutb(w_n22909_0[1]),.din(n22909));
	jspl3 jspl3_w_n22911_0(.douta(w_n22911_0[0]),.doutb(w_n22911_0[1]),.doutc(w_n22911_0[2]),.din(n22911));
	jspl jspl_w_n22912_0(.douta(w_n22912_0[0]),.doutb(w_n22912_0[1]),.din(n22912));
	jspl jspl_w_n22916_0(.douta(w_n22916_0[0]),.doutb(w_n22916_0[1]),.din(n22916));
	jspl jspl_w_n22917_0(.douta(w_n22917_0[0]),.doutb(w_n22917_0[1]),.din(n22917));
	jspl3 jspl3_w_n22919_0(.douta(w_n22919_0[0]),.doutb(w_n22919_0[1]),.doutc(w_n22919_0[2]),.din(n22919));
	jspl jspl_w_n22920_0(.douta(w_n22920_0[0]),.doutb(w_n22920_0[1]),.din(n22920));
	jspl jspl_w_n22924_0(.douta(w_n22924_0[0]),.doutb(w_n22924_0[1]),.din(n22924));
	jspl jspl_w_n22925_0(.douta(w_n22925_0[0]),.doutb(w_n22925_0[1]),.din(n22925));
	jspl3 jspl3_w_n22927_0(.douta(w_n22927_0[0]),.doutb(w_n22927_0[1]),.doutc(w_n22927_0[2]),.din(n22927));
	jspl jspl_w_n22928_0(.douta(w_n22928_0[0]),.doutb(w_n22928_0[1]),.din(n22928));
	jspl jspl_w_n22932_0(.douta(w_n22932_0[0]),.doutb(w_n22932_0[1]),.din(n22932));
	jspl jspl_w_n22933_0(.douta(w_n22933_0[0]),.doutb(w_n22933_0[1]),.din(n22933));
	jspl3 jspl3_w_n22935_0(.douta(w_n22935_0[0]),.doutb(w_n22935_0[1]),.doutc(w_n22935_0[2]),.din(n22935));
	jspl jspl_w_n22936_0(.douta(w_n22936_0[0]),.doutb(w_n22936_0[1]),.din(n22936));
	jspl jspl_w_n22940_0(.douta(w_n22940_0[0]),.doutb(w_n22940_0[1]),.din(n22940));
	jspl3 jspl3_w_n22942_0(.douta(w_n22942_0[0]),.doutb(w_n22942_0[1]),.doutc(w_n22942_0[2]),.din(n22942));
	jspl jspl_w_n22943_0(.douta(w_n22943_0[0]),.doutb(w_n22943_0[1]),.din(n22943));
	jspl jspl_w_n22947_0(.douta(w_n22947_0[0]),.doutb(w_n22947_0[1]),.din(n22947));
	jspl jspl_w_n22948_0(.douta(w_n22948_0[0]),.doutb(w_n22948_0[1]),.din(n22948));
	jspl3 jspl3_w_n22950_0(.douta(w_n22950_0[0]),.doutb(w_n22950_0[1]),.doutc(w_n22950_0[2]),.din(n22950));
	jspl jspl_w_n22951_0(.douta(w_n22951_0[0]),.doutb(w_n22951_0[1]),.din(n22951));
	jspl jspl_w_n22955_0(.douta(w_n22955_0[0]),.doutb(w_n22955_0[1]),.din(n22955));
	jspl jspl_w_n22956_0(.douta(w_n22956_0[0]),.doutb(w_n22956_0[1]),.din(n22956));
	jspl3 jspl3_w_n22958_0(.douta(w_n22958_0[0]),.doutb(w_n22958_0[1]),.doutc(w_n22958_0[2]),.din(n22958));
	jspl jspl_w_n22959_0(.douta(w_n22959_0[0]),.doutb(w_n22959_0[1]),.din(n22959));
	jspl jspl_w_n22963_0(.douta(w_n22963_0[0]),.doutb(w_n22963_0[1]),.din(n22963));
	jspl jspl_w_n22964_0(.douta(w_n22964_0[0]),.doutb(w_n22964_0[1]),.din(n22964));
	jspl3 jspl3_w_n22966_0(.douta(w_n22966_0[0]),.doutb(w_n22966_0[1]),.doutc(w_n22966_0[2]),.din(n22966));
	jspl jspl_w_n22967_0(.douta(w_n22967_0[0]),.doutb(w_n22967_0[1]),.din(n22967));
	jspl jspl_w_n22971_0(.douta(w_n22971_0[0]),.doutb(w_n22971_0[1]),.din(n22971));
	jspl jspl_w_n22972_0(.douta(w_n22972_0[0]),.doutb(w_n22972_0[1]),.din(n22972));
	jspl3 jspl3_w_n22974_0(.douta(w_n22974_0[0]),.doutb(w_n22974_0[1]),.doutc(w_n22974_0[2]),.din(n22974));
	jspl jspl_w_n22975_0(.douta(w_n22975_0[0]),.doutb(w_n22975_0[1]),.din(n22975));
	jspl jspl_w_n22979_0(.douta(w_n22979_0[0]),.doutb(w_n22979_0[1]),.din(n22979));
	jspl jspl_w_n22980_0(.douta(w_n22980_0[0]),.doutb(w_n22980_0[1]),.din(n22980));
	jspl3 jspl3_w_n22982_0(.douta(w_n22982_0[0]),.doutb(w_n22982_0[1]),.doutc(w_n22982_0[2]),.din(n22982));
	jspl jspl_w_n22983_0(.douta(w_n22983_0[0]),.doutb(w_n22983_0[1]),.din(n22983));
	jspl jspl_w_n22987_0(.douta(w_n22987_0[0]),.doutb(w_n22987_0[1]),.din(n22987));
	jspl3 jspl3_w_n22989_0(.douta(w_n22989_0[0]),.doutb(w_n22989_0[1]),.doutc(w_n22989_0[2]),.din(n22989));
	jspl jspl_w_n22990_0(.douta(w_n22990_0[0]),.doutb(w_n22990_0[1]),.din(n22990));
	jspl jspl_w_n22994_0(.douta(w_n22994_0[0]),.doutb(w_n22994_0[1]),.din(n22994));
	jspl jspl_w_n22995_0(.douta(w_n22995_0[0]),.doutb(w_n22995_0[1]),.din(n22995));
	jspl3 jspl3_w_n22997_0(.douta(w_n22997_0[0]),.doutb(w_n22997_0[1]),.doutc(w_n22997_0[2]),.din(n22997));
	jspl jspl_w_n22998_0(.douta(w_n22998_0[0]),.doutb(w_n22998_0[1]),.din(n22998));
	jspl jspl_w_n23002_0(.douta(w_n23002_0[0]),.doutb(w_n23002_0[1]),.din(n23002));
	jspl3 jspl3_w_n23004_0(.douta(w_n23004_0[0]),.doutb(w_n23004_0[1]),.doutc(w_n23004_0[2]),.din(n23004));
	jspl jspl_w_n23005_0(.douta(w_n23005_0[0]),.doutb(w_n23005_0[1]),.din(n23005));
	jspl jspl_w_n23009_0(.douta(w_n23009_0[0]),.doutb(w_n23009_0[1]),.din(n23009));
	jspl jspl_w_n23010_0(.douta(w_n23010_0[0]),.doutb(w_n23010_0[1]),.din(n23010));
	jspl3 jspl3_w_n23012_0(.douta(w_n23012_0[0]),.doutb(w_n23012_0[1]),.doutc(w_n23012_0[2]),.din(n23012));
	jspl jspl_w_n23013_0(.douta(w_n23013_0[0]),.doutb(w_n23013_0[1]),.din(n23013));
	jspl jspl_w_n23017_0(.douta(w_n23017_0[0]),.doutb(w_n23017_0[1]),.din(n23017));
	jspl jspl_w_n23018_0(.douta(w_n23018_0[0]),.doutb(w_n23018_0[1]),.din(n23018));
	jspl3 jspl3_w_n23020_0(.douta(w_n23020_0[0]),.doutb(w_n23020_0[1]),.doutc(w_n23020_0[2]),.din(n23020));
	jspl jspl_w_n23021_0(.douta(w_n23021_0[0]),.doutb(w_n23021_0[1]),.din(n23021));
	jspl jspl_w_n23025_0(.douta(w_n23025_0[0]),.doutb(w_n23025_0[1]),.din(n23025));
	jspl3 jspl3_w_n23027_0(.douta(w_n23027_0[0]),.doutb(w_n23027_0[1]),.doutc(w_n23027_0[2]),.din(n23027));
	jspl jspl_w_n23028_0(.douta(w_n23028_0[0]),.doutb(w_n23028_0[1]),.din(n23028));
	jspl jspl_w_n23032_0(.douta(w_n23032_0[0]),.doutb(w_n23032_0[1]),.din(n23032));
	jspl3 jspl3_w_n23034_0(.douta(w_n23034_0[0]),.doutb(w_n23034_0[1]),.doutc(w_n23034_0[2]),.din(n23034));
	jspl jspl_w_n23035_0(.douta(w_n23035_0[0]),.doutb(w_n23035_0[1]),.din(n23035));
	jspl jspl_w_n23039_0(.douta(w_n23039_0[0]),.doutb(w_n23039_0[1]),.din(n23039));
	jspl jspl_w_n23040_0(.douta(w_n23040_0[0]),.doutb(w_n23040_0[1]),.din(n23040));
	jspl3 jspl3_w_n23042_0(.douta(w_n23042_0[0]),.doutb(w_n23042_0[1]),.doutc(w_n23042_0[2]),.din(n23042));
	jspl jspl_w_n23043_0(.douta(w_n23043_0[0]),.doutb(w_n23043_0[1]),.din(n23043));
	jspl jspl_w_n23047_0(.douta(w_n23047_0[0]),.doutb(w_n23047_0[1]),.din(n23047));
	jspl jspl_w_n23048_0(.douta(w_n23048_0[0]),.doutb(w_n23048_0[1]),.din(n23048));
	jspl3 jspl3_w_n23050_0(.douta(w_n23050_0[0]),.doutb(w_n23050_0[1]),.doutc(w_n23050_0[2]),.din(n23050));
	jspl jspl_w_n23051_0(.douta(w_n23051_0[0]),.doutb(w_n23051_0[1]),.din(n23051));
	jspl3 jspl3_w_n23055_0(.douta(w_n23055_0[0]),.doutb(w_n23055_0[1]),.doutc(w_n23055_0[2]),.din(n23055));
	jspl jspl_w_n23058_0(.douta(w_n23058_0[0]),.doutb(w_n23058_0[1]),.din(n23058));
	jspl jspl_w_n23061_0(.douta(w_n23061_0[0]),.doutb(w_n23061_0[1]),.din(n23061));
	jspl jspl_w_n23062_0(.douta(w_n23062_0[0]),.doutb(w_n23062_0[1]),.din(n23062));
	jspl3 jspl3_w_n23063_0(.douta(w_n23063_0[0]),.doutb(w_n23063_0[1]),.doutc(w_n23063_0[2]),.din(n23063));
	jspl jspl_w_n23063_1(.douta(w_n23063_1[0]),.doutb(w_n23063_1[1]),.din(w_n23063_0[0]));
	jspl jspl_w_n23064_0(.douta(w_n23064_0[0]),.doutb(w_n23064_0[1]),.din(n23064));
	jspl jspl_w_n23065_0(.douta(w_n23065_0[0]),.doutb(w_n23065_0[1]),.din(n23065));
	jspl jspl_w_n23138_0(.douta(w_n23138_0[0]),.doutb(w_n23138_0[1]),.din(n23138));
	jspl jspl_w_n23142_0(.douta(w_n23142_0[0]),.doutb(w_n23142_0[1]),.din(n23142));
	jspl jspl_w_n23146_0(.douta(w_n23146_0[0]),.doutb(w_n23146_0[1]),.din(n23146));
	jspl jspl_w_n23153_0(.douta(w_n23153_0[0]),.doutb(w_n23153_0[1]),.din(n23153));
	jspl jspl_w_n23160_0(.douta(w_n23160_0[0]),.doutb(w_n23160_0[1]),.din(n23160));
	jspl jspl_w_n23173_0(.douta(w_n23173_0[0]),.doutb(w_n23173_0[1]),.din(n23173));
	jspl jspl_w_n23186_0(.douta(w_n23186_0[0]),.doutb(w_n23186_0[1]),.din(n23186));
	jspl jspl_w_n23193_0(.douta(w_n23193_0[0]),.doutb(w_n23193_0[1]),.din(n23193));
	jspl jspl_w_n23200_0(.douta(w_n23200_0[0]),.doutb(w_n23200_0[1]),.din(n23200));
	jspl jspl_w_n23210_0(.douta(w_n23210_0[0]),.doutb(w_n23210_0[1]),.din(n23210));
	jspl jspl_w_n23214_0(.douta(w_n23214_0[0]),.doutb(w_n23214_0[1]),.din(n23214));
	jspl jspl_w_n23221_0(.douta(w_n23221_0[0]),.doutb(w_n23221_0[1]),.din(n23221));
	jspl jspl_w_n23228_0(.douta(w_n23228_0[0]),.doutb(w_n23228_0[1]),.din(n23228));
	jspl jspl_w_n23241_0(.douta(w_n23241_0[0]),.doutb(w_n23241_0[1]),.din(n23241));
	jspl jspl_w_n23248_0(.douta(w_n23248_0[0]),.doutb(w_n23248_0[1]),.din(n23248));
	jspl jspl_w_n23255_0(.douta(w_n23255_0[0]),.doutb(w_n23255_0[1]),.din(n23255));
	jspl jspl_w_n23262_0(.douta(w_n23262_0[0]),.doutb(w_n23262_0[1]),.din(n23262));
	jspl jspl_w_n23275_0(.douta(w_n23275_0[0]),.doutb(w_n23275_0[1]),.din(n23275));
	jspl jspl_w_n23294_0(.douta(w_n23294_0[0]),.doutb(w_n23294_0[1]),.din(n23294));
	jspl jspl_w_n23301_0(.douta(w_n23301_0[0]),.doutb(w_n23301_0[1]),.din(n23301));
	jspl jspl_w_n23311_0(.douta(w_n23311_0[0]),.doutb(w_n23311_0[1]),.din(n23311));
	jspl jspl_w_n23315_0(.douta(w_n23315_0[0]),.doutb(w_n23315_0[1]),.din(n23315));
	jspl jspl_w_n23326_0(.douta(w_n23326_0[0]),.doutb(w_n23326_0[1]),.din(n23326));
	jspl jspl_w_n23327_0(.douta(w_n23327_0[0]),.doutb(w_n23327_0[1]),.din(n23327));
	jspl jspl_w_n23335_0(.douta(w_n23335_0[0]),.doutb(w_n23335_0[1]),.din(n23335));
	jspl jspl_w_n23336_0(.douta(w_n23336_0[0]),.doutb(w_n23336_0[1]),.din(n23336));
	jspl jspl_w_n23339_0(.douta(w_n23339_0[0]),.doutb(w_n23339_0[1]),.din(n23339));
	jspl jspl_w_n23344_0(.douta(w_n23344_0[0]),.doutb(w_n23344_0[1]),.din(n23344));
	jspl3 jspl3_w_n23345_0(.douta(w_n23345_0[0]),.doutb(w_n23345_0[1]),.doutc(w_n23345_0[2]),.din(n23345));
	jspl3 jspl3_w_n23345_1(.douta(w_n23345_1[0]),.doutb(w_n23345_1[1]),.doutc(w_n23345_1[2]),.din(w_n23345_0[0]));
	jspl3 jspl3_w_n23345_2(.douta(w_n23345_2[0]),.doutb(w_n23345_2[1]),.doutc(w_n23345_2[2]),.din(w_n23345_0[1]));
	jspl3 jspl3_w_n23345_3(.douta(w_n23345_3[0]),.doutb(w_n23345_3[1]),.doutc(w_n23345_3[2]),.din(w_n23345_0[2]));
	jspl3 jspl3_w_n23345_4(.douta(w_n23345_4[0]),.doutb(w_n23345_4[1]),.doutc(w_n23345_4[2]),.din(w_n23345_1[0]));
	jspl3 jspl3_w_n23345_5(.douta(w_n23345_5[0]),.doutb(w_n23345_5[1]),.doutc(w_n23345_5[2]),.din(w_n23345_1[1]));
	jspl3 jspl3_w_n23345_6(.douta(w_n23345_6[0]),.doutb(w_n23345_6[1]),.doutc(w_n23345_6[2]),.din(w_n23345_1[2]));
	jspl3 jspl3_w_n23345_7(.douta(w_n23345_7[0]),.doutb(w_n23345_7[1]),.doutc(w_n23345_7[2]),.din(w_n23345_2[0]));
	jspl3 jspl3_w_n23345_8(.douta(w_n23345_8[0]),.doutb(w_n23345_8[1]),.doutc(w_n23345_8[2]),.din(w_n23345_2[1]));
	jspl3 jspl3_w_n23345_9(.douta(w_n23345_9[0]),.doutb(w_n23345_9[1]),.doutc(w_n23345_9[2]),.din(w_n23345_2[2]));
	jspl3 jspl3_w_n23345_10(.douta(w_n23345_10[0]),.doutb(w_n23345_10[1]),.doutc(w_n23345_10[2]),.din(w_n23345_3[0]));
	jspl3 jspl3_w_n23345_11(.douta(w_n23345_11[0]),.doutb(w_n23345_11[1]),.doutc(w_n23345_11[2]),.din(w_n23345_3[1]));
	jspl3 jspl3_w_n23345_12(.douta(w_n23345_12[0]),.doutb(w_n23345_12[1]),.doutc(w_n23345_12[2]),.din(w_n23345_3[2]));
	jspl3 jspl3_w_n23345_13(.douta(w_n23345_13[0]),.doutb(w_n23345_13[1]),.doutc(w_n23345_13[2]),.din(w_n23345_4[0]));
	jspl3 jspl3_w_n23345_14(.douta(w_n23345_14[0]),.doutb(w_n23345_14[1]),.doutc(w_n23345_14[2]),.din(w_n23345_4[1]));
	jspl3 jspl3_w_n23345_15(.douta(w_n23345_15[0]),.doutb(w_n23345_15[1]),.doutc(w_n23345_15[2]),.din(w_n23345_4[2]));
	jspl3 jspl3_w_n23345_16(.douta(w_n23345_16[0]),.doutb(w_n23345_16[1]),.doutc(w_n23345_16[2]),.din(w_n23345_5[0]));
	jspl3 jspl3_w_n23345_17(.douta(w_n23345_17[0]),.doutb(w_n23345_17[1]),.doutc(w_n23345_17[2]),.din(w_n23345_5[1]));
	jspl3 jspl3_w_n23345_18(.douta(w_n23345_18[0]),.doutb(w_n23345_18[1]),.doutc(w_n23345_18[2]),.din(w_n23345_5[2]));
	jspl3 jspl3_w_n23345_19(.douta(w_n23345_19[0]),.doutb(w_n23345_19[1]),.doutc(w_n23345_19[2]),.din(w_n23345_6[0]));
	jspl3 jspl3_w_n23345_20(.douta(w_n23345_20[0]),.doutb(w_n23345_20[1]),.doutc(w_n23345_20[2]),.din(w_n23345_6[1]));
	jspl3 jspl3_w_n23345_21(.douta(w_n23345_21[0]),.doutb(w_n23345_21[1]),.doutc(w_n23345_21[2]),.din(w_n23345_6[2]));
	jspl3 jspl3_w_n23345_22(.douta(w_n23345_22[0]),.doutb(w_n23345_22[1]),.doutc(w_n23345_22[2]),.din(w_n23345_7[0]));
	jspl3 jspl3_w_n23345_23(.douta(w_n23345_23[0]),.doutb(w_n23345_23[1]),.doutc(w_n23345_23[2]),.din(w_n23345_7[1]));
	jspl3 jspl3_w_n23345_24(.douta(w_n23345_24[0]),.doutb(w_n23345_24[1]),.doutc(w_n23345_24[2]),.din(w_n23345_7[2]));
	jspl3 jspl3_w_n23345_25(.douta(w_n23345_25[0]),.doutb(w_n23345_25[1]),.doutc(w_n23345_25[2]),.din(w_n23345_8[0]));
	jspl3 jspl3_w_n23345_26(.douta(w_n23345_26[0]),.doutb(w_n23345_26[1]),.doutc(w_n23345_26[2]),.din(w_n23345_8[1]));
	jspl3 jspl3_w_n23345_27(.douta(w_n23345_27[0]),.doutb(w_n23345_27[1]),.doutc(w_n23345_27[2]),.din(w_n23345_8[2]));
	jspl3 jspl3_w_n23345_28(.douta(w_n23345_28[0]),.doutb(w_n23345_28[1]),.doutc(w_n23345_28[2]),.din(w_n23345_9[0]));
	jspl3 jspl3_w_n23345_29(.douta(w_n23345_29[0]),.doutb(w_n23345_29[1]),.doutc(w_n23345_29[2]),.din(w_n23345_9[1]));
	jspl3 jspl3_w_n23345_30(.douta(w_n23345_30[0]),.doutb(w_n23345_30[1]),.doutc(w_n23345_30[2]),.din(w_n23345_9[2]));
	jspl3 jspl3_w_n23345_31(.douta(w_n23345_31[0]),.doutb(w_n23345_31[1]),.doutc(w_n23345_31[2]),.din(w_n23345_10[0]));
	jspl jspl_w_n23345_32(.douta(w_n23345_32[0]),.doutb(w_n23345_32[1]),.din(w_n23345_10[1]));
	jspl jspl_w_n23348_0(.douta(w_n23348_0[0]),.doutb(w_n23348_0[1]),.din(n23348));
	jspl3 jspl3_w_n23349_0(.douta(w_n23349_0[0]),.doutb(w_n23349_0[1]),.doutc(w_n23349_0[2]),.din(n23349));
	jspl3 jspl3_w_n23351_0(.douta(w_n23351_0[0]),.doutb(w_n23351_0[1]),.doutc(w_n23351_0[2]),.din(n23351));
	jspl jspl_w_n23351_1(.douta(w_n23351_1[0]),.doutb(w_n23351_1[1]),.din(w_n23351_0[0]));
	jspl jspl_w_n23352_0(.douta(w_n23352_0[0]),.doutb(w_n23352_0[1]),.din(n23352));
	jspl3 jspl3_w_n23353_0(.douta(w_n23353_0[0]),.doutb(w_n23353_0[1]),.doutc(w_n23353_0[2]),.din(n23353));
	jspl jspl_w_n23354_0(.douta(w_n23354_0[0]),.doutb(w_n23354_0[1]),.din(n23354));
	jspl3 jspl3_w_n23356_0(.douta(w_n23356_0[0]),.doutb(w_n23356_0[1]),.doutc(w_n23356_0[2]),.din(n23356));
	jspl jspl_w_n23357_0(.douta(w_n23357_0[0]),.doutb(w_n23357_0[1]),.din(n23357));
	jspl3 jspl3_w_n23364_0(.douta(w_n23364_0[0]),.doutb(w_n23364_0[1]),.doutc(w_n23364_0[2]),.din(n23364));
	jspl jspl_w_n23365_0(.douta(w_n23365_0[0]),.doutb(w_n23365_0[1]),.din(n23365));
	jspl jspl_w_n23368_0(.douta(w_n23368_0[0]),.doutb(w_n23368_0[1]),.din(n23368));
	jspl jspl_w_n23371_0(.douta(w_n23371_0[0]),.doutb(w_n23371_0[1]),.din(n23371));
	jspl3 jspl3_w_n23373_0(.douta(w_n23373_0[0]),.doutb(w_n23373_0[1]),.doutc(w_n23373_0[2]),.din(n23373));
	jspl jspl_w_n23374_0(.douta(w_n23374_0[0]),.doutb(w_n23374_0[1]),.din(n23374));
	jspl3 jspl3_w_n23378_0(.douta(w_n23378_0[0]),.doutb(w_n23378_0[1]),.doutc(w_n23378_0[2]),.din(n23378));
	jspl3 jspl3_w_n23380_0(.douta(w_n23380_0[0]),.doutb(w_n23380_0[1]),.doutc(w_n23380_0[2]),.din(n23380));
	jspl jspl_w_n23381_0(.douta(w_n23381_0[0]),.doutb(w_n23381_0[1]),.din(n23381));
	jspl3 jspl3_w_n23385_0(.douta(w_n23385_0[0]),.doutb(w_n23385_0[1]),.doutc(w_n23385_0[2]),.din(n23385));
	jspl3 jspl3_w_n23387_0(.douta(w_n23387_0[0]),.doutb(w_n23387_0[1]),.doutc(w_n23387_0[2]),.din(n23387));
	jspl jspl_w_n23388_0(.douta(w_n23388_0[0]),.doutb(w_n23388_0[1]),.din(n23388));
	jspl3 jspl3_w_n23392_0(.douta(w_n23392_0[0]),.doutb(w_n23392_0[1]),.doutc(w_n23392_0[2]),.din(n23392));
	jspl3 jspl3_w_n23395_0(.douta(w_n23395_0[0]),.doutb(w_n23395_0[1]),.doutc(w_n23395_0[2]),.din(n23395));
	jspl jspl_w_n23396_0(.douta(w_n23396_0[0]),.doutb(w_n23396_0[1]),.din(n23396));
	jspl3 jspl3_w_n23400_0(.douta(w_n23400_0[0]),.doutb(w_n23400_0[1]),.doutc(w_n23400_0[2]),.din(n23400));
	jspl3 jspl3_w_n23403_0(.douta(w_n23403_0[0]),.doutb(w_n23403_0[1]),.doutc(w_n23403_0[2]),.din(n23403));
	jspl jspl_w_n23404_0(.douta(w_n23404_0[0]),.doutb(w_n23404_0[1]),.din(n23404));
	jspl3 jspl3_w_n23408_0(.douta(w_n23408_0[0]),.doutb(w_n23408_0[1]),.doutc(w_n23408_0[2]),.din(n23408));
	jspl3 jspl3_w_n23411_0(.douta(w_n23411_0[0]),.doutb(w_n23411_0[1]),.doutc(w_n23411_0[2]),.din(n23411));
	jspl jspl_w_n23412_0(.douta(w_n23412_0[0]),.doutb(w_n23412_0[1]),.din(n23412));
	jspl3 jspl3_w_n23416_0(.douta(w_n23416_0[0]),.doutb(w_n23416_0[1]),.doutc(w_n23416_0[2]),.din(n23416));
	jspl3 jspl3_w_n23418_0(.douta(w_n23418_0[0]),.doutb(w_n23418_0[1]),.doutc(w_n23418_0[2]),.din(n23418));
	jspl jspl_w_n23419_0(.douta(w_n23419_0[0]),.doutb(w_n23419_0[1]),.din(n23419));
	jspl3 jspl3_w_n23423_0(.douta(w_n23423_0[0]),.doutb(w_n23423_0[1]),.doutc(w_n23423_0[2]),.din(n23423));
	jspl3 jspl3_w_n23426_0(.douta(w_n23426_0[0]),.doutb(w_n23426_0[1]),.doutc(w_n23426_0[2]),.din(n23426));
	jspl jspl_w_n23427_0(.douta(w_n23427_0[0]),.doutb(w_n23427_0[1]),.din(n23427));
	jspl3 jspl3_w_n23431_0(.douta(w_n23431_0[0]),.doutb(w_n23431_0[1]),.doutc(w_n23431_0[2]),.din(n23431));
	jspl3 jspl3_w_n23433_0(.douta(w_n23433_0[0]),.doutb(w_n23433_0[1]),.doutc(w_n23433_0[2]),.din(n23433));
	jspl jspl_w_n23434_0(.douta(w_n23434_0[0]),.doutb(w_n23434_0[1]),.din(n23434));
	jspl3 jspl3_w_n23438_0(.douta(w_n23438_0[0]),.doutb(w_n23438_0[1]),.doutc(w_n23438_0[2]),.din(n23438));
	jspl3 jspl3_w_n23441_0(.douta(w_n23441_0[0]),.doutb(w_n23441_0[1]),.doutc(w_n23441_0[2]),.din(n23441));
	jspl jspl_w_n23442_0(.douta(w_n23442_0[0]),.doutb(w_n23442_0[1]),.din(n23442));
	jspl3 jspl3_w_n23446_0(.douta(w_n23446_0[0]),.doutb(w_n23446_0[1]),.doutc(w_n23446_0[2]),.din(n23446));
	jspl3 jspl3_w_n23448_0(.douta(w_n23448_0[0]),.doutb(w_n23448_0[1]),.doutc(w_n23448_0[2]),.din(n23448));
	jspl jspl_w_n23449_0(.douta(w_n23449_0[0]),.doutb(w_n23449_0[1]),.din(n23449));
	jspl3 jspl3_w_n23453_0(.douta(w_n23453_0[0]),.doutb(w_n23453_0[1]),.doutc(w_n23453_0[2]),.din(n23453));
	jspl3 jspl3_w_n23455_0(.douta(w_n23455_0[0]),.doutb(w_n23455_0[1]),.doutc(w_n23455_0[2]),.din(n23455));
	jspl jspl_w_n23456_0(.douta(w_n23456_0[0]),.doutb(w_n23456_0[1]),.din(n23456));
	jspl3 jspl3_w_n23460_0(.douta(w_n23460_0[0]),.doutb(w_n23460_0[1]),.doutc(w_n23460_0[2]),.din(n23460));
	jspl3 jspl3_w_n23462_0(.douta(w_n23462_0[0]),.doutb(w_n23462_0[1]),.doutc(w_n23462_0[2]),.din(n23462));
	jspl jspl_w_n23463_0(.douta(w_n23463_0[0]),.doutb(w_n23463_0[1]),.din(n23463));
	jspl3 jspl3_w_n23467_0(.douta(w_n23467_0[0]),.doutb(w_n23467_0[1]),.doutc(w_n23467_0[2]),.din(n23467));
	jspl3 jspl3_w_n23470_0(.douta(w_n23470_0[0]),.doutb(w_n23470_0[1]),.doutc(w_n23470_0[2]),.din(n23470));
	jspl jspl_w_n23471_0(.douta(w_n23471_0[0]),.doutb(w_n23471_0[1]),.din(n23471));
	jspl3 jspl3_w_n23475_0(.douta(w_n23475_0[0]),.doutb(w_n23475_0[1]),.doutc(w_n23475_0[2]),.din(n23475));
	jspl3 jspl3_w_n23477_0(.douta(w_n23477_0[0]),.doutb(w_n23477_0[1]),.doutc(w_n23477_0[2]),.din(n23477));
	jspl jspl_w_n23478_0(.douta(w_n23478_0[0]),.doutb(w_n23478_0[1]),.din(n23478));
	jspl3 jspl3_w_n23482_0(.douta(w_n23482_0[0]),.doutb(w_n23482_0[1]),.doutc(w_n23482_0[2]),.din(n23482));
	jspl3 jspl3_w_n23484_0(.douta(w_n23484_0[0]),.doutb(w_n23484_0[1]),.doutc(w_n23484_0[2]),.din(n23484));
	jspl jspl_w_n23485_0(.douta(w_n23485_0[0]),.doutb(w_n23485_0[1]),.din(n23485));
	jspl3 jspl3_w_n23489_0(.douta(w_n23489_0[0]),.doutb(w_n23489_0[1]),.doutc(w_n23489_0[2]),.din(n23489));
	jspl3 jspl3_w_n23491_0(.douta(w_n23491_0[0]),.doutb(w_n23491_0[1]),.doutc(w_n23491_0[2]),.din(n23491));
	jspl jspl_w_n23492_0(.douta(w_n23492_0[0]),.doutb(w_n23492_0[1]),.din(n23492));
	jspl3 jspl3_w_n23496_0(.douta(w_n23496_0[0]),.doutb(w_n23496_0[1]),.doutc(w_n23496_0[2]),.din(n23496));
	jspl3 jspl3_w_n23499_0(.douta(w_n23499_0[0]),.doutb(w_n23499_0[1]),.doutc(w_n23499_0[2]),.din(n23499));
	jspl jspl_w_n23500_0(.douta(w_n23500_0[0]),.doutb(w_n23500_0[1]),.din(n23500));
	jspl3 jspl3_w_n23504_0(.douta(w_n23504_0[0]),.doutb(w_n23504_0[1]),.doutc(w_n23504_0[2]),.din(n23504));
	jspl3 jspl3_w_n23506_0(.douta(w_n23506_0[0]),.doutb(w_n23506_0[1]),.doutc(w_n23506_0[2]),.din(n23506));
	jspl jspl_w_n23507_0(.douta(w_n23507_0[0]),.doutb(w_n23507_0[1]),.din(n23507));
	jspl3 jspl3_w_n23511_0(.douta(w_n23511_0[0]),.doutb(w_n23511_0[1]),.doutc(w_n23511_0[2]),.din(n23511));
	jspl3 jspl3_w_n23514_0(.douta(w_n23514_0[0]),.doutb(w_n23514_0[1]),.doutc(w_n23514_0[2]),.din(n23514));
	jspl jspl_w_n23515_0(.douta(w_n23515_0[0]),.doutb(w_n23515_0[1]),.din(n23515));
	jspl3 jspl3_w_n23519_0(.douta(w_n23519_0[0]),.doutb(w_n23519_0[1]),.doutc(w_n23519_0[2]),.din(n23519));
	jspl3 jspl3_w_n23521_0(.douta(w_n23521_0[0]),.doutb(w_n23521_0[1]),.doutc(w_n23521_0[2]),.din(n23521));
	jspl jspl_w_n23522_0(.douta(w_n23522_0[0]),.doutb(w_n23522_0[1]),.din(n23522));
	jspl3 jspl3_w_n23526_0(.douta(w_n23526_0[0]),.doutb(w_n23526_0[1]),.doutc(w_n23526_0[2]),.din(n23526));
	jspl3 jspl3_w_n23529_0(.douta(w_n23529_0[0]),.doutb(w_n23529_0[1]),.doutc(w_n23529_0[2]),.din(n23529));
	jspl jspl_w_n23530_0(.douta(w_n23530_0[0]),.doutb(w_n23530_0[1]),.din(n23530));
	jspl3 jspl3_w_n23534_0(.douta(w_n23534_0[0]),.doutb(w_n23534_0[1]),.doutc(w_n23534_0[2]),.din(n23534));
	jspl3 jspl3_w_n23536_0(.douta(w_n23536_0[0]),.doutb(w_n23536_0[1]),.doutc(w_n23536_0[2]),.din(n23536));
	jspl jspl_w_n23537_0(.douta(w_n23537_0[0]),.doutb(w_n23537_0[1]),.din(n23537));
	jspl3 jspl3_w_n23541_0(.douta(w_n23541_0[0]),.doutb(w_n23541_0[1]),.doutc(w_n23541_0[2]),.din(n23541));
	jspl3 jspl3_w_n23543_0(.douta(w_n23543_0[0]),.doutb(w_n23543_0[1]),.doutc(w_n23543_0[2]),.din(n23543));
	jspl jspl_w_n23544_0(.douta(w_n23544_0[0]),.doutb(w_n23544_0[1]),.din(n23544));
	jspl3 jspl3_w_n23548_0(.douta(w_n23548_0[0]),.doutb(w_n23548_0[1]),.doutc(w_n23548_0[2]),.din(n23548));
	jspl3 jspl3_w_n23551_0(.douta(w_n23551_0[0]),.doutb(w_n23551_0[1]),.doutc(w_n23551_0[2]),.din(n23551));
	jspl jspl_w_n23552_0(.douta(w_n23552_0[0]),.doutb(w_n23552_0[1]),.din(n23552));
	jspl3 jspl3_w_n23556_0(.douta(w_n23556_0[0]),.doutb(w_n23556_0[1]),.doutc(w_n23556_0[2]),.din(n23556));
	jspl3 jspl3_w_n23559_0(.douta(w_n23559_0[0]),.doutb(w_n23559_0[1]),.doutc(w_n23559_0[2]),.din(n23559));
	jspl jspl_w_n23560_0(.douta(w_n23560_0[0]),.doutb(w_n23560_0[1]),.din(n23560));
	jspl3 jspl3_w_n23564_0(.douta(w_n23564_0[0]),.doutb(w_n23564_0[1]),.doutc(w_n23564_0[2]),.din(n23564));
	jspl3 jspl3_w_n23566_0(.douta(w_n23566_0[0]),.doutb(w_n23566_0[1]),.doutc(w_n23566_0[2]),.din(n23566));
	jspl jspl_w_n23567_0(.douta(w_n23567_0[0]),.doutb(w_n23567_0[1]),.din(n23567));
	jspl3 jspl3_w_n23571_0(.douta(w_n23571_0[0]),.doutb(w_n23571_0[1]),.doutc(w_n23571_0[2]),.din(n23571));
	jspl3 jspl3_w_n23574_0(.douta(w_n23574_0[0]),.doutb(w_n23574_0[1]),.doutc(w_n23574_0[2]),.din(n23574));
	jspl jspl_w_n23575_0(.douta(w_n23575_0[0]),.doutb(w_n23575_0[1]),.din(n23575));
	jspl3 jspl3_w_n23579_0(.douta(w_n23579_0[0]),.doutb(w_n23579_0[1]),.doutc(w_n23579_0[2]),.din(n23579));
	jspl3 jspl3_w_n23581_0(.douta(w_n23581_0[0]),.doutb(w_n23581_0[1]),.doutc(w_n23581_0[2]),.din(n23581));
	jspl jspl_w_n23582_0(.douta(w_n23582_0[0]),.doutb(w_n23582_0[1]),.din(n23582));
	jspl3 jspl3_w_n23586_0(.douta(w_n23586_0[0]),.doutb(w_n23586_0[1]),.doutc(w_n23586_0[2]),.din(n23586));
	jspl3 jspl3_w_n23589_0(.douta(w_n23589_0[0]),.doutb(w_n23589_0[1]),.doutc(w_n23589_0[2]),.din(n23589));
	jspl jspl_w_n23590_0(.douta(w_n23590_0[0]),.doutb(w_n23590_0[1]),.din(n23590));
	jspl3 jspl3_w_n23594_0(.douta(w_n23594_0[0]),.doutb(w_n23594_0[1]),.doutc(w_n23594_0[2]),.din(n23594));
	jspl3 jspl3_w_n23596_0(.douta(w_n23596_0[0]),.doutb(w_n23596_0[1]),.doutc(w_n23596_0[2]),.din(n23596));
	jspl jspl_w_n23597_0(.douta(w_n23597_0[0]),.doutb(w_n23597_0[1]),.din(n23597));
	jspl3 jspl3_w_n23601_0(.douta(w_n23601_0[0]),.doutb(w_n23601_0[1]),.doutc(w_n23601_0[2]),.din(n23601));
	jspl3 jspl3_w_n23603_0(.douta(w_n23603_0[0]),.doutb(w_n23603_0[1]),.doutc(w_n23603_0[2]),.din(n23603));
	jspl jspl_w_n23604_0(.douta(w_n23604_0[0]),.doutb(w_n23604_0[1]),.din(n23604));
	jspl3 jspl3_w_n23608_0(.douta(w_n23608_0[0]),.doutb(w_n23608_0[1]),.doutc(w_n23608_0[2]),.din(n23608));
	jspl3 jspl3_w_n23610_0(.douta(w_n23610_0[0]),.doutb(w_n23610_0[1]),.doutc(w_n23610_0[2]),.din(n23610));
	jspl jspl_w_n23611_0(.douta(w_n23611_0[0]),.doutb(w_n23611_0[1]),.din(n23611));
	jspl3 jspl3_w_n23615_0(.douta(w_n23615_0[0]),.doutb(w_n23615_0[1]),.doutc(w_n23615_0[2]),.din(n23615));
	jspl3 jspl3_w_n23618_0(.douta(w_n23618_0[0]),.doutb(w_n23618_0[1]),.doutc(w_n23618_0[2]),.din(n23618));
	jspl jspl_w_n23619_0(.douta(w_n23619_0[0]),.doutb(w_n23619_0[1]),.din(n23619));
	jspl3 jspl3_w_n23623_0(.douta(w_n23623_0[0]),.doutb(w_n23623_0[1]),.doutc(w_n23623_0[2]),.din(n23623));
	jspl3 jspl3_w_n23625_0(.douta(w_n23625_0[0]),.doutb(w_n23625_0[1]),.doutc(w_n23625_0[2]),.din(n23625));
	jspl jspl_w_n23626_0(.douta(w_n23626_0[0]),.doutb(w_n23626_0[1]),.din(n23626));
	jspl3 jspl3_w_n23630_0(.douta(w_n23630_0[0]),.doutb(w_n23630_0[1]),.doutc(w_n23630_0[2]),.din(n23630));
	jspl3 jspl3_w_n23633_0(.douta(w_n23633_0[0]),.doutb(w_n23633_0[1]),.doutc(w_n23633_0[2]),.din(n23633));
	jspl jspl_w_n23634_0(.douta(w_n23634_0[0]),.doutb(w_n23634_0[1]),.din(n23634));
	jspl3 jspl3_w_n23638_0(.douta(w_n23638_0[0]),.doutb(w_n23638_0[1]),.doutc(w_n23638_0[2]),.din(n23638));
	jspl3 jspl3_w_n23640_0(.douta(w_n23640_0[0]),.doutb(w_n23640_0[1]),.doutc(w_n23640_0[2]),.din(n23640));
	jspl jspl_w_n23641_0(.douta(w_n23641_0[0]),.doutb(w_n23641_0[1]),.din(n23641));
	jspl3 jspl3_w_n23645_0(.douta(w_n23645_0[0]),.doutb(w_n23645_0[1]),.doutc(w_n23645_0[2]),.din(n23645));
	jspl3 jspl3_w_n23648_0(.douta(w_n23648_0[0]),.doutb(w_n23648_0[1]),.doutc(w_n23648_0[2]),.din(n23648));
	jspl jspl_w_n23649_0(.douta(w_n23649_0[0]),.doutb(w_n23649_0[1]),.din(n23649));
	jspl3 jspl3_w_n23653_0(.douta(w_n23653_0[0]),.doutb(w_n23653_0[1]),.doutc(w_n23653_0[2]),.din(n23653));
	jspl3 jspl3_w_n23655_0(.douta(w_n23655_0[0]),.doutb(w_n23655_0[1]),.doutc(w_n23655_0[2]),.din(n23655));
	jspl jspl_w_n23656_0(.douta(w_n23656_0[0]),.doutb(w_n23656_0[1]),.din(n23656));
	jspl3 jspl3_w_n23660_0(.douta(w_n23660_0[0]),.doutb(w_n23660_0[1]),.doutc(w_n23660_0[2]),.din(n23660));
	jspl3 jspl3_w_n23663_0(.douta(w_n23663_0[0]),.doutb(w_n23663_0[1]),.doutc(w_n23663_0[2]),.din(n23663));
	jspl jspl_w_n23664_0(.douta(w_n23664_0[0]),.doutb(w_n23664_0[1]),.din(n23664));
	jspl3 jspl3_w_n23668_0(.douta(w_n23668_0[0]),.doutb(w_n23668_0[1]),.doutc(w_n23668_0[2]),.din(n23668));
	jspl3 jspl3_w_n23670_0(.douta(w_n23670_0[0]),.doutb(w_n23670_0[1]),.doutc(w_n23670_0[2]),.din(n23670));
	jspl jspl_w_n23671_0(.douta(w_n23671_0[0]),.doutb(w_n23671_0[1]),.din(n23671));
	jspl3 jspl3_w_n23675_0(.douta(w_n23675_0[0]),.doutb(w_n23675_0[1]),.doutc(w_n23675_0[2]),.din(n23675));
	jspl3 jspl3_w_n23677_0(.douta(w_n23677_0[0]),.doutb(w_n23677_0[1]),.doutc(w_n23677_0[2]),.din(n23677));
	jspl jspl_w_n23678_0(.douta(w_n23678_0[0]),.doutb(w_n23678_0[1]),.din(n23678));
	jspl3 jspl3_w_n23682_0(.douta(w_n23682_0[0]),.doutb(w_n23682_0[1]),.doutc(w_n23682_0[2]),.din(n23682));
	jspl3 jspl3_w_n23684_0(.douta(w_n23684_0[0]),.doutb(w_n23684_0[1]),.doutc(w_n23684_0[2]),.din(n23684));
	jspl jspl_w_n23685_0(.douta(w_n23685_0[0]),.doutb(w_n23685_0[1]),.din(n23685));
	jspl3 jspl3_w_n23689_0(.douta(w_n23689_0[0]),.doutb(w_n23689_0[1]),.doutc(w_n23689_0[2]),.din(n23689));
	jspl3 jspl3_w_n23692_0(.douta(w_n23692_0[0]),.doutb(w_n23692_0[1]),.doutc(w_n23692_0[2]),.din(n23692));
	jspl jspl_w_n23693_0(.douta(w_n23693_0[0]),.doutb(w_n23693_0[1]),.din(n23693));
	jspl3 jspl3_w_n23697_0(.douta(w_n23697_0[0]),.doutb(w_n23697_0[1]),.doutc(w_n23697_0[2]),.din(n23697));
	jspl3 jspl3_w_n23699_0(.douta(w_n23699_0[0]),.doutb(w_n23699_0[1]),.doutc(w_n23699_0[2]),.din(n23699));
	jspl jspl_w_n23700_0(.douta(w_n23700_0[0]),.doutb(w_n23700_0[1]),.din(n23700));
	jspl3 jspl3_w_n23704_0(.douta(w_n23704_0[0]),.doutb(w_n23704_0[1]),.doutc(w_n23704_0[2]),.din(n23704));
	jspl3 jspl3_w_n23706_0(.douta(w_n23706_0[0]),.doutb(w_n23706_0[1]),.doutc(w_n23706_0[2]),.din(n23706));
	jspl jspl_w_n23707_0(.douta(w_n23707_0[0]),.doutb(w_n23707_0[1]),.din(n23707));
	jspl3 jspl3_w_n23711_0(.douta(w_n23711_0[0]),.doutb(w_n23711_0[1]),.doutc(w_n23711_0[2]),.din(n23711));
	jspl3 jspl3_w_n23713_0(.douta(w_n23713_0[0]),.doutb(w_n23713_0[1]),.doutc(w_n23713_0[2]),.din(n23713));
	jspl jspl_w_n23714_0(.douta(w_n23714_0[0]),.doutb(w_n23714_0[1]),.din(n23714));
	jspl3 jspl3_w_n23718_0(.douta(w_n23718_0[0]),.doutb(w_n23718_0[1]),.doutc(w_n23718_0[2]),.din(n23718));
	jspl3 jspl3_w_n23720_0(.douta(w_n23720_0[0]),.doutb(w_n23720_0[1]),.doutc(w_n23720_0[2]),.din(n23720));
	jspl jspl_w_n23721_0(.douta(w_n23721_0[0]),.doutb(w_n23721_0[1]),.din(n23721));
	jspl3 jspl3_w_n23725_0(.douta(w_n23725_0[0]),.doutb(w_n23725_0[1]),.doutc(w_n23725_0[2]),.din(n23725));
	jspl3 jspl3_w_n23727_0(.douta(w_n23727_0[0]),.doutb(w_n23727_0[1]),.doutc(w_n23727_0[2]),.din(n23727));
	jspl jspl_w_n23728_0(.douta(w_n23728_0[0]),.doutb(w_n23728_0[1]),.din(n23728));
	jspl3 jspl3_w_n23732_0(.douta(w_n23732_0[0]),.doutb(w_n23732_0[1]),.doutc(w_n23732_0[2]),.din(n23732));
	jspl3 jspl3_w_n23735_0(.douta(w_n23735_0[0]),.doutb(w_n23735_0[1]),.doutc(w_n23735_0[2]),.din(n23735));
	jspl jspl_w_n23736_0(.douta(w_n23736_0[0]),.doutb(w_n23736_0[1]),.din(n23736));
	jspl3 jspl3_w_n23740_0(.douta(w_n23740_0[0]),.doutb(w_n23740_0[1]),.doutc(w_n23740_0[2]),.din(n23740));
	jspl3 jspl3_w_n23742_0(.douta(w_n23742_0[0]),.doutb(w_n23742_0[1]),.doutc(w_n23742_0[2]),.din(n23742));
	jspl jspl_w_n23743_0(.douta(w_n23743_0[0]),.doutb(w_n23743_0[1]),.din(n23743));
	jspl3 jspl3_w_n23747_0(.douta(w_n23747_0[0]),.doutb(w_n23747_0[1]),.doutc(w_n23747_0[2]),.din(n23747));
	jspl3 jspl3_w_n23750_0(.douta(w_n23750_0[0]),.doutb(w_n23750_0[1]),.doutc(w_n23750_0[2]),.din(n23750));
	jspl jspl_w_n23751_0(.douta(w_n23751_0[0]),.doutb(w_n23751_0[1]),.din(n23751));
	jspl3 jspl3_w_n23755_0(.douta(w_n23755_0[0]),.doutb(w_n23755_0[1]),.doutc(w_n23755_0[2]),.din(n23755));
	jspl3 jspl3_w_n23757_0(.douta(w_n23757_0[0]),.doutb(w_n23757_0[1]),.doutc(w_n23757_0[2]),.din(n23757));
	jspl jspl_w_n23758_0(.douta(w_n23758_0[0]),.doutb(w_n23758_0[1]),.din(n23758));
	jspl jspl_w_n23762_0(.douta(w_n23762_0[0]),.doutb(w_n23762_0[1]),.din(n23762));
	jspl3 jspl3_w_n23764_0(.douta(w_n23764_0[0]),.doutb(w_n23764_0[1]),.doutc(w_n23764_0[2]),.din(n23764));
	jspl jspl_w_n23765_0(.douta(w_n23765_0[0]),.doutb(w_n23765_0[1]),.din(n23765));
	jspl3 jspl3_w_n23769_0(.douta(w_n23769_0[0]),.doutb(w_n23769_0[1]),.doutc(w_n23769_0[2]),.din(n23769));
	jspl3 jspl3_w_n23772_0(.douta(w_n23772_0[0]),.doutb(w_n23772_0[1]),.doutc(w_n23772_0[2]),.din(n23772));
	jspl jspl_w_n23773_0(.douta(w_n23773_0[0]),.doutb(w_n23773_0[1]),.din(n23773));
	jspl3 jspl3_w_n23777_0(.douta(w_n23777_0[0]),.doutb(w_n23777_0[1]),.doutc(w_n23777_0[2]),.din(n23777));
	jspl3 jspl3_w_n23780_0(.douta(w_n23780_0[0]),.doutb(w_n23780_0[1]),.doutc(w_n23780_0[2]),.din(n23780));
	jspl jspl_w_n23781_0(.douta(w_n23781_0[0]),.doutb(w_n23781_0[1]),.din(n23781));
	jspl3 jspl3_w_n23785_0(.douta(w_n23785_0[0]),.doutb(w_n23785_0[1]),.doutc(w_n23785_0[2]),.din(n23785));
	jspl3 jspl3_w_n23787_0(.douta(w_n23787_0[0]),.doutb(w_n23787_0[1]),.doutc(w_n23787_0[2]),.din(n23787));
	jspl jspl_w_n23788_0(.douta(w_n23788_0[0]),.doutb(w_n23788_0[1]),.din(n23788));
	jspl3 jspl3_w_n23792_0(.douta(w_n23792_0[0]),.doutb(w_n23792_0[1]),.doutc(w_n23792_0[2]),.din(n23792));
	jspl3 jspl3_w_n23794_0(.douta(w_n23794_0[0]),.doutb(w_n23794_0[1]),.doutc(w_n23794_0[2]),.din(n23794));
	jspl jspl_w_n23794_1(.douta(w_n23794_1[0]),.doutb(w_n23794_1[1]),.din(w_n23794_0[0]));
	jspl3 jspl3_w_n23795_0(.douta(w_n23795_0[0]),.doutb(w_n23795_0[1]),.doutc(w_n23795_0[2]),.din(n23795));
	jspl jspl_w_n23796_0(.douta(w_n23796_0[0]),.doutb(w_n23796_0[1]),.din(n23796));
	jspl jspl_w_n23805_0(.douta(w_n23805_0[0]),.doutb(w_n23805_0[1]),.din(n23805));
	jspl jspl_w_n23806_0(.douta(w_n23806_0[0]),.doutb(w_n23806_0[1]),.din(n23806));
	jspl jspl_w_n23810_0(.douta(w_n23810_0[0]),.doutb(w_n23810_0[1]),.din(n23810));
	jspl jspl_w_n23811_0(.douta(w_n23811_0[0]),.doutb(w_n23811_0[1]),.din(n23811));
	jspl3 jspl3_w_n23812_0(.douta(w_n23812_0[0]),.doutb(w_n23812_0[1]),.doutc(w_n23812_0[2]),.din(n23812));
	jspl jspl_w_n23813_0(.douta(w_n23813_0[0]),.doutb(w_n23813_0[1]),.din(n23813));
	jspl jspl_w_n23818_0(.douta(w_n23818_0[0]),.doutb(w_n23818_0[1]),.din(n23818));
	jspl jspl_w_n23884_0(.douta(w_n23884_0[0]),.doutb(w_n23884_0[1]),.din(n23884));
	jspl jspl_w_n23888_0(.douta(w_n23888_0[0]),.doutb(w_n23888_0[1]),.din(n23888));
	jspl jspl_w_n24080_0(.douta(w_n24080_0[0]),.doutb(w_n24080_0[1]),.din(n24080));
	jspl jspl_w_n24097_0(.douta(w_n24097_0[0]),.doutb(w_n24097_0[1]),.din(n24097));
	jspl jspl_w_n24102_0(.douta(w_n24102_0[0]),.doutb(w_n24102_0[1]),.din(n24102));
	jspl3 jspl3_w_n24103_0(.douta(w_n24103_0[0]),.doutb(w_n24103_0[1]),.doutc(w_n24103_0[2]),.din(n24103));
	jspl3 jspl3_w_n24103_1(.douta(w_n24103_1[0]),.doutb(w_n24103_1[1]),.doutc(w_n24103_1[2]),.din(w_n24103_0[0]));
	jspl jspl_w_n24104_0(.douta(w_n24104_0[0]),.doutb(w_n24104_0[1]),.din(n24104));
	jspl jspl_w_n24105_0(.douta(w_n24105_0[0]),.doutb(w_n24105_0[1]),.din(n24105));
	jspl3 jspl3_w_n24107_0(.douta(w_n24107_0[0]),.doutb(w_n24107_0[1]),.doutc(w_n24107_0[2]),.din(n24107));
	jspl jspl_w_n24108_0(.douta(w_n24108_0[0]),.doutb(w_n24108_0[1]),.din(n24108));
	jspl jspl_w_n24112_0(.douta(w_n24112_0[0]),.doutb(w_n24112_0[1]),.din(n24112));
	jspl jspl_w_n24113_0(.douta(w_n24113_0[0]),.doutb(w_n24113_0[1]),.din(n24113));
	jspl3 jspl3_w_n24115_0(.douta(w_n24115_0[0]),.doutb(w_n24115_0[1]),.doutc(w_n24115_0[2]),.din(n24115));
	jspl jspl_w_n24116_0(.douta(w_n24116_0[0]),.doutb(w_n24116_0[1]),.din(n24116));
	jspl3 jspl3_w_n24120_0(.douta(w_n24120_0[0]),.doutb(w_n24120_0[1]),.doutc(w_n24120_0[2]),.din(n24120));
	jspl3 jspl3_w_n24122_0(.douta(w_n24122_0[0]),.doutb(w_n24122_0[1]),.doutc(w_n24122_0[2]),.din(n24122));
	jspl jspl_w_n24123_0(.douta(w_n24123_0[0]),.doutb(w_n24123_0[1]),.din(n24123));
	jspl3 jspl3_w_n24127_0(.douta(w_n24127_0[0]),.doutb(w_n24127_0[1]),.doutc(w_n24127_0[2]),.din(n24127));
	jspl3 jspl3_w_n24129_0(.douta(w_n24129_0[0]),.doutb(w_n24129_0[1]),.doutc(w_n24129_0[2]),.din(n24129));
	jspl jspl_w_n24130_0(.douta(w_n24130_0[0]),.doutb(w_n24130_0[1]),.din(n24130));
	jspl jspl_w_n24134_0(.douta(w_n24134_0[0]),.doutb(w_n24134_0[1]),.din(n24134));
	jspl jspl_w_n24135_0(.douta(w_n24135_0[0]),.doutb(w_n24135_0[1]),.din(n24135));
	jspl3 jspl3_w_n24137_0(.douta(w_n24137_0[0]),.doutb(w_n24137_0[1]),.doutc(w_n24137_0[2]),.din(n24137));
	jspl jspl_w_n24138_0(.douta(w_n24138_0[0]),.doutb(w_n24138_0[1]),.din(n24138));
	jspl jspl_w_n24142_0(.douta(w_n24142_0[0]),.doutb(w_n24142_0[1]),.din(n24142));
	jspl jspl_w_n24143_0(.douta(w_n24143_0[0]),.doutb(w_n24143_0[1]),.din(n24143));
	jspl3 jspl3_w_n24145_0(.douta(w_n24145_0[0]),.doutb(w_n24145_0[1]),.doutc(w_n24145_0[2]),.din(n24145));
	jspl jspl_w_n24146_0(.douta(w_n24146_0[0]),.doutb(w_n24146_0[1]),.din(n24146));
	jspl3 jspl3_w_n24150_0(.douta(w_n24150_0[0]),.doutb(w_n24150_0[1]),.doutc(w_n24150_0[2]),.din(n24150));
	jspl3 jspl3_w_n24152_0(.douta(w_n24152_0[0]),.doutb(w_n24152_0[1]),.doutc(w_n24152_0[2]),.din(n24152));
	jspl jspl_w_n24153_0(.douta(w_n24153_0[0]),.doutb(w_n24153_0[1]),.din(n24153));
	jspl3 jspl3_w_n24157_0(.douta(w_n24157_0[0]),.doutb(w_n24157_0[1]),.doutc(w_n24157_0[2]),.din(n24157));
	jspl3 jspl3_w_n24159_0(.douta(w_n24159_0[0]),.doutb(w_n24159_0[1]),.doutc(w_n24159_0[2]),.din(n24159));
	jspl jspl_w_n24160_0(.douta(w_n24160_0[0]),.doutb(w_n24160_0[1]),.din(n24160));
	jspl3 jspl3_w_n24164_0(.douta(w_n24164_0[0]),.doutb(w_n24164_0[1]),.doutc(w_n24164_0[2]),.din(n24164));
	jspl3 jspl3_w_n24166_0(.douta(w_n24166_0[0]),.doutb(w_n24166_0[1]),.doutc(w_n24166_0[2]),.din(n24166));
	jspl jspl_w_n24167_0(.douta(w_n24167_0[0]),.doutb(w_n24167_0[1]),.din(n24167));
	jspl jspl_w_n24171_0(.douta(w_n24171_0[0]),.doutb(w_n24171_0[1]),.din(n24171));
	jspl jspl_w_n24172_0(.douta(w_n24172_0[0]),.doutb(w_n24172_0[1]),.din(n24172));
	jspl3 jspl3_w_n24174_0(.douta(w_n24174_0[0]),.doutb(w_n24174_0[1]),.doutc(w_n24174_0[2]),.din(n24174));
	jspl jspl_w_n24175_0(.douta(w_n24175_0[0]),.doutb(w_n24175_0[1]),.din(n24175));
	jspl3 jspl3_w_n24179_0(.douta(w_n24179_0[0]),.doutb(w_n24179_0[1]),.doutc(w_n24179_0[2]),.din(n24179));
	jspl3 jspl3_w_n24181_0(.douta(w_n24181_0[0]),.doutb(w_n24181_0[1]),.doutc(w_n24181_0[2]),.din(n24181));
	jspl jspl_w_n24182_0(.douta(w_n24182_0[0]),.doutb(w_n24182_0[1]),.din(n24182));
	jspl jspl_w_n24186_0(.douta(w_n24186_0[0]),.doutb(w_n24186_0[1]),.din(n24186));
	jspl jspl_w_n24187_0(.douta(w_n24187_0[0]),.doutb(w_n24187_0[1]),.din(n24187));
	jspl3 jspl3_w_n24189_0(.douta(w_n24189_0[0]),.doutb(w_n24189_0[1]),.doutc(w_n24189_0[2]),.din(n24189));
	jspl jspl_w_n24190_0(.douta(w_n24190_0[0]),.doutb(w_n24190_0[1]),.din(n24190));
	jspl3 jspl3_w_n24194_0(.douta(w_n24194_0[0]),.doutb(w_n24194_0[1]),.doutc(w_n24194_0[2]),.din(n24194));
	jspl3 jspl3_w_n24196_0(.douta(w_n24196_0[0]),.doutb(w_n24196_0[1]),.doutc(w_n24196_0[2]),.din(n24196));
	jspl jspl_w_n24197_0(.douta(w_n24197_0[0]),.doutb(w_n24197_0[1]),.din(n24197));
	jspl jspl_w_n24201_0(.douta(w_n24201_0[0]),.doutb(w_n24201_0[1]),.din(n24201));
	jspl jspl_w_n24202_0(.douta(w_n24202_0[0]),.doutb(w_n24202_0[1]),.din(n24202));
	jspl3 jspl3_w_n24204_0(.douta(w_n24204_0[0]),.doutb(w_n24204_0[1]),.doutc(w_n24204_0[2]),.din(n24204));
	jspl jspl_w_n24205_0(.douta(w_n24205_0[0]),.doutb(w_n24205_0[1]),.din(n24205));
	jspl jspl_w_n24209_0(.douta(w_n24209_0[0]),.doutb(w_n24209_0[1]),.din(n24209));
	jspl jspl_w_n24210_0(.douta(w_n24210_0[0]),.doutb(w_n24210_0[1]),.din(n24210));
	jspl3 jspl3_w_n24212_0(.douta(w_n24212_0[0]),.doutb(w_n24212_0[1]),.doutc(w_n24212_0[2]),.din(n24212));
	jspl jspl_w_n24213_0(.douta(w_n24213_0[0]),.doutb(w_n24213_0[1]),.din(n24213));
	jspl jspl_w_n24217_0(.douta(w_n24217_0[0]),.doutb(w_n24217_0[1]),.din(n24217));
	jspl jspl_w_n24218_0(.douta(w_n24218_0[0]),.doutb(w_n24218_0[1]),.din(n24218));
	jspl3 jspl3_w_n24220_0(.douta(w_n24220_0[0]),.doutb(w_n24220_0[1]),.doutc(w_n24220_0[2]),.din(n24220));
	jspl jspl_w_n24221_0(.douta(w_n24221_0[0]),.doutb(w_n24221_0[1]),.din(n24221));
	jspl3 jspl3_w_n24225_0(.douta(w_n24225_0[0]),.doutb(w_n24225_0[1]),.doutc(w_n24225_0[2]),.din(n24225));
	jspl3 jspl3_w_n24227_0(.douta(w_n24227_0[0]),.doutb(w_n24227_0[1]),.doutc(w_n24227_0[2]),.din(n24227));
	jspl jspl_w_n24228_0(.douta(w_n24228_0[0]),.doutb(w_n24228_0[1]),.din(n24228));
	jspl jspl_w_n24232_0(.douta(w_n24232_0[0]),.doutb(w_n24232_0[1]),.din(n24232));
	jspl jspl_w_n24233_0(.douta(w_n24233_0[0]),.doutb(w_n24233_0[1]),.din(n24233));
	jspl3 jspl3_w_n24235_0(.douta(w_n24235_0[0]),.doutb(w_n24235_0[1]),.doutc(w_n24235_0[2]),.din(n24235));
	jspl jspl_w_n24236_0(.douta(w_n24236_0[0]),.doutb(w_n24236_0[1]),.din(n24236));
	jspl jspl_w_n24240_0(.douta(w_n24240_0[0]),.doutb(w_n24240_0[1]),.din(n24240));
	jspl jspl_w_n24241_0(.douta(w_n24241_0[0]),.doutb(w_n24241_0[1]),.din(n24241));
	jspl3 jspl3_w_n24243_0(.douta(w_n24243_0[0]),.doutb(w_n24243_0[1]),.doutc(w_n24243_0[2]),.din(n24243));
	jspl jspl_w_n24244_0(.douta(w_n24244_0[0]),.doutb(w_n24244_0[1]),.din(n24244));
	jspl jspl_w_n24248_0(.douta(w_n24248_0[0]),.doutb(w_n24248_0[1]),.din(n24248));
	jspl jspl_w_n24249_0(.douta(w_n24249_0[0]),.doutb(w_n24249_0[1]),.din(n24249));
	jspl3 jspl3_w_n24251_0(.douta(w_n24251_0[0]),.doutb(w_n24251_0[1]),.doutc(w_n24251_0[2]),.din(n24251));
	jspl jspl_w_n24252_0(.douta(w_n24252_0[0]),.doutb(w_n24252_0[1]),.din(n24252));
	jspl3 jspl3_w_n24256_0(.douta(w_n24256_0[0]),.doutb(w_n24256_0[1]),.doutc(w_n24256_0[2]),.din(n24256));
	jspl3 jspl3_w_n24258_0(.douta(w_n24258_0[0]),.doutb(w_n24258_0[1]),.doutc(w_n24258_0[2]),.din(n24258));
	jspl jspl_w_n24259_0(.douta(w_n24259_0[0]),.doutb(w_n24259_0[1]),.din(n24259));
	jspl jspl_w_n24263_0(.douta(w_n24263_0[0]),.doutb(w_n24263_0[1]),.din(n24263));
	jspl jspl_w_n24264_0(.douta(w_n24264_0[0]),.doutb(w_n24264_0[1]),.din(n24264));
	jspl3 jspl3_w_n24266_0(.douta(w_n24266_0[0]),.doutb(w_n24266_0[1]),.doutc(w_n24266_0[2]),.din(n24266));
	jspl jspl_w_n24267_0(.douta(w_n24267_0[0]),.doutb(w_n24267_0[1]),.din(n24267));
	jspl3 jspl3_w_n24271_0(.douta(w_n24271_0[0]),.doutb(w_n24271_0[1]),.doutc(w_n24271_0[2]),.din(n24271));
	jspl3 jspl3_w_n24273_0(.douta(w_n24273_0[0]),.doutb(w_n24273_0[1]),.doutc(w_n24273_0[2]),.din(n24273));
	jspl jspl_w_n24274_0(.douta(w_n24274_0[0]),.doutb(w_n24274_0[1]),.din(n24274));
	jspl jspl_w_n24278_0(.douta(w_n24278_0[0]),.doutb(w_n24278_0[1]),.din(n24278));
	jspl jspl_w_n24279_0(.douta(w_n24279_0[0]),.doutb(w_n24279_0[1]),.din(n24279));
	jspl3 jspl3_w_n24281_0(.douta(w_n24281_0[0]),.doutb(w_n24281_0[1]),.doutc(w_n24281_0[2]),.din(n24281));
	jspl jspl_w_n24282_0(.douta(w_n24282_0[0]),.doutb(w_n24282_0[1]),.din(n24282));
	jspl3 jspl3_w_n24286_0(.douta(w_n24286_0[0]),.doutb(w_n24286_0[1]),.doutc(w_n24286_0[2]),.din(n24286));
	jspl3 jspl3_w_n24288_0(.douta(w_n24288_0[0]),.doutb(w_n24288_0[1]),.doutc(w_n24288_0[2]),.din(n24288));
	jspl jspl_w_n24289_0(.douta(w_n24289_0[0]),.doutb(w_n24289_0[1]),.din(n24289));
	jspl jspl_w_n24293_0(.douta(w_n24293_0[0]),.doutb(w_n24293_0[1]),.din(n24293));
	jspl jspl_w_n24294_0(.douta(w_n24294_0[0]),.doutb(w_n24294_0[1]),.din(n24294));
	jspl3 jspl3_w_n24296_0(.douta(w_n24296_0[0]),.doutb(w_n24296_0[1]),.doutc(w_n24296_0[2]),.din(n24296));
	jspl jspl_w_n24297_0(.douta(w_n24297_0[0]),.doutb(w_n24297_0[1]),.din(n24297));
	jspl jspl_w_n24301_0(.douta(w_n24301_0[0]),.doutb(w_n24301_0[1]),.din(n24301));
	jspl jspl_w_n24302_0(.douta(w_n24302_0[0]),.doutb(w_n24302_0[1]),.din(n24302));
	jspl3 jspl3_w_n24304_0(.douta(w_n24304_0[0]),.doutb(w_n24304_0[1]),.doutc(w_n24304_0[2]),.din(n24304));
	jspl jspl_w_n24305_0(.douta(w_n24305_0[0]),.doutb(w_n24305_0[1]),.din(n24305));
	jspl3 jspl3_w_n24309_0(.douta(w_n24309_0[0]),.doutb(w_n24309_0[1]),.doutc(w_n24309_0[2]),.din(n24309));
	jspl3 jspl3_w_n24311_0(.douta(w_n24311_0[0]),.doutb(w_n24311_0[1]),.doutc(w_n24311_0[2]),.din(n24311));
	jspl jspl_w_n24312_0(.douta(w_n24312_0[0]),.doutb(w_n24312_0[1]),.din(n24312));
	jspl3 jspl3_w_n24316_0(.douta(w_n24316_0[0]),.doutb(w_n24316_0[1]),.doutc(w_n24316_0[2]),.din(n24316));
	jspl3 jspl3_w_n24318_0(.douta(w_n24318_0[0]),.doutb(w_n24318_0[1]),.doutc(w_n24318_0[2]),.din(n24318));
	jspl jspl_w_n24319_0(.douta(w_n24319_0[0]),.doutb(w_n24319_0[1]),.din(n24319));
	jspl jspl_w_n24323_0(.douta(w_n24323_0[0]),.doutb(w_n24323_0[1]),.din(n24323));
	jspl jspl_w_n24324_0(.douta(w_n24324_0[0]),.doutb(w_n24324_0[1]),.din(n24324));
	jspl3 jspl3_w_n24326_0(.douta(w_n24326_0[0]),.doutb(w_n24326_0[1]),.doutc(w_n24326_0[2]),.din(n24326));
	jspl jspl_w_n24327_0(.douta(w_n24327_0[0]),.doutb(w_n24327_0[1]),.din(n24327));
	jspl3 jspl3_w_n24331_0(.douta(w_n24331_0[0]),.doutb(w_n24331_0[1]),.doutc(w_n24331_0[2]),.din(n24331));
	jspl3 jspl3_w_n24333_0(.douta(w_n24333_0[0]),.doutb(w_n24333_0[1]),.doutc(w_n24333_0[2]),.din(n24333));
	jspl jspl_w_n24334_0(.douta(w_n24334_0[0]),.doutb(w_n24334_0[1]),.din(n24334));
	jspl jspl_w_n24338_0(.douta(w_n24338_0[0]),.doutb(w_n24338_0[1]),.din(n24338));
	jspl jspl_w_n24339_0(.douta(w_n24339_0[0]),.doutb(w_n24339_0[1]),.din(n24339));
	jspl3 jspl3_w_n24341_0(.douta(w_n24341_0[0]),.doutb(w_n24341_0[1]),.doutc(w_n24341_0[2]),.din(n24341));
	jspl jspl_w_n24342_0(.douta(w_n24342_0[0]),.doutb(w_n24342_0[1]),.din(n24342));
	jspl3 jspl3_w_n24346_0(.douta(w_n24346_0[0]),.doutb(w_n24346_0[1]),.doutc(w_n24346_0[2]),.din(n24346));
	jspl3 jspl3_w_n24348_0(.douta(w_n24348_0[0]),.doutb(w_n24348_0[1]),.doutc(w_n24348_0[2]),.din(n24348));
	jspl jspl_w_n24349_0(.douta(w_n24349_0[0]),.doutb(w_n24349_0[1]),.din(n24349));
	jspl jspl_w_n24353_0(.douta(w_n24353_0[0]),.doutb(w_n24353_0[1]),.din(n24353));
	jspl jspl_w_n24354_0(.douta(w_n24354_0[0]),.doutb(w_n24354_0[1]),.din(n24354));
	jspl3 jspl3_w_n24356_0(.douta(w_n24356_0[0]),.doutb(w_n24356_0[1]),.doutc(w_n24356_0[2]),.din(n24356));
	jspl jspl_w_n24357_0(.douta(w_n24357_0[0]),.doutb(w_n24357_0[1]),.din(n24357));
	jspl jspl_w_n24361_0(.douta(w_n24361_0[0]),.doutb(w_n24361_0[1]),.din(n24361));
	jspl jspl_w_n24362_0(.douta(w_n24362_0[0]),.doutb(w_n24362_0[1]),.din(n24362));
	jspl3 jspl3_w_n24364_0(.douta(w_n24364_0[0]),.doutb(w_n24364_0[1]),.doutc(w_n24364_0[2]),.din(n24364));
	jspl jspl_w_n24365_0(.douta(w_n24365_0[0]),.doutb(w_n24365_0[1]),.din(n24365));
	jspl jspl_w_n24369_0(.douta(w_n24369_0[0]),.doutb(w_n24369_0[1]),.din(n24369));
	jspl jspl_w_n24370_0(.douta(w_n24370_0[0]),.doutb(w_n24370_0[1]),.din(n24370));
	jspl3 jspl3_w_n24372_0(.douta(w_n24372_0[0]),.doutb(w_n24372_0[1]),.doutc(w_n24372_0[2]),.din(n24372));
	jspl jspl_w_n24373_0(.douta(w_n24373_0[0]),.doutb(w_n24373_0[1]),.din(n24373));
	jspl3 jspl3_w_n24377_0(.douta(w_n24377_0[0]),.doutb(w_n24377_0[1]),.doutc(w_n24377_0[2]),.din(n24377));
	jspl3 jspl3_w_n24379_0(.douta(w_n24379_0[0]),.doutb(w_n24379_0[1]),.doutc(w_n24379_0[2]),.din(n24379));
	jspl jspl_w_n24380_0(.douta(w_n24380_0[0]),.doutb(w_n24380_0[1]),.din(n24380));
	jspl jspl_w_n24384_0(.douta(w_n24384_0[0]),.doutb(w_n24384_0[1]),.din(n24384));
	jspl jspl_w_n24385_0(.douta(w_n24385_0[0]),.doutb(w_n24385_0[1]),.din(n24385));
	jspl3 jspl3_w_n24387_0(.douta(w_n24387_0[0]),.doutb(w_n24387_0[1]),.doutc(w_n24387_0[2]),.din(n24387));
	jspl jspl_w_n24388_0(.douta(w_n24388_0[0]),.doutb(w_n24388_0[1]),.din(n24388));
	jspl3 jspl3_w_n24392_0(.douta(w_n24392_0[0]),.doutb(w_n24392_0[1]),.doutc(w_n24392_0[2]),.din(n24392));
	jspl3 jspl3_w_n24394_0(.douta(w_n24394_0[0]),.doutb(w_n24394_0[1]),.doutc(w_n24394_0[2]),.din(n24394));
	jspl jspl_w_n24395_0(.douta(w_n24395_0[0]),.doutb(w_n24395_0[1]),.din(n24395));
	jspl jspl_w_n24399_0(.douta(w_n24399_0[0]),.doutb(w_n24399_0[1]),.din(n24399));
	jspl jspl_w_n24400_0(.douta(w_n24400_0[0]),.doutb(w_n24400_0[1]),.din(n24400));
	jspl3 jspl3_w_n24402_0(.douta(w_n24402_0[0]),.doutb(w_n24402_0[1]),.doutc(w_n24402_0[2]),.din(n24402));
	jspl jspl_w_n24403_0(.douta(w_n24403_0[0]),.doutb(w_n24403_0[1]),.din(n24403));
	jspl3 jspl3_w_n24407_0(.douta(w_n24407_0[0]),.doutb(w_n24407_0[1]),.doutc(w_n24407_0[2]),.din(n24407));
	jspl3 jspl3_w_n24409_0(.douta(w_n24409_0[0]),.doutb(w_n24409_0[1]),.doutc(w_n24409_0[2]),.din(n24409));
	jspl jspl_w_n24410_0(.douta(w_n24410_0[0]),.doutb(w_n24410_0[1]),.din(n24410));
	jspl jspl_w_n24414_0(.douta(w_n24414_0[0]),.doutb(w_n24414_0[1]),.din(n24414));
	jspl jspl_w_n24415_0(.douta(w_n24415_0[0]),.doutb(w_n24415_0[1]),.din(n24415));
	jspl3 jspl3_w_n24417_0(.douta(w_n24417_0[0]),.doutb(w_n24417_0[1]),.doutc(w_n24417_0[2]),.din(n24417));
	jspl jspl_w_n24418_0(.douta(w_n24418_0[0]),.doutb(w_n24418_0[1]),.din(n24418));
	jspl3 jspl3_w_n24422_0(.douta(w_n24422_0[0]),.doutb(w_n24422_0[1]),.doutc(w_n24422_0[2]),.din(n24422));
	jspl3 jspl3_w_n24424_0(.douta(w_n24424_0[0]),.doutb(w_n24424_0[1]),.doutc(w_n24424_0[2]),.din(n24424));
	jspl jspl_w_n24425_0(.douta(w_n24425_0[0]),.doutb(w_n24425_0[1]),.din(n24425));
	jspl jspl_w_n24429_0(.douta(w_n24429_0[0]),.doutb(w_n24429_0[1]),.din(n24429));
	jspl jspl_w_n24430_0(.douta(w_n24430_0[0]),.doutb(w_n24430_0[1]),.din(n24430));
	jspl3 jspl3_w_n24432_0(.douta(w_n24432_0[0]),.doutb(w_n24432_0[1]),.doutc(w_n24432_0[2]),.din(n24432));
	jspl jspl_w_n24433_0(.douta(w_n24433_0[0]),.doutb(w_n24433_0[1]),.din(n24433));
	jspl jspl_w_n24437_0(.douta(w_n24437_0[0]),.doutb(w_n24437_0[1]),.din(n24437));
	jspl jspl_w_n24438_0(.douta(w_n24438_0[0]),.doutb(w_n24438_0[1]),.din(n24438));
	jspl3 jspl3_w_n24440_0(.douta(w_n24440_0[0]),.doutb(w_n24440_0[1]),.doutc(w_n24440_0[2]),.din(n24440));
	jspl jspl_w_n24441_0(.douta(w_n24441_0[0]),.doutb(w_n24441_0[1]),.din(n24441));
	jspl jspl_w_n24445_0(.douta(w_n24445_0[0]),.doutb(w_n24445_0[1]),.din(n24445));
	jspl jspl_w_n24446_0(.douta(w_n24446_0[0]),.doutb(w_n24446_0[1]),.din(n24446));
	jspl3 jspl3_w_n24448_0(.douta(w_n24448_0[0]),.doutb(w_n24448_0[1]),.doutc(w_n24448_0[2]),.din(n24448));
	jspl jspl_w_n24449_0(.douta(w_n24449_0[0]),.doutb(w_n24449_0[1]),.din(n24449));
	jspl3 jspl3_w_n24453_0(.douta(w_n24453_0[0]),.doutb(w_n24453_0[1]),.doutc(w_n24453_0[2]),.din(n24453));
	jspl3 jspl3_w_n24455_0(.douta(w_n24455_0[0]),.doutb(w_n24455_0[1]),.doutc(w_n24455_0[2]),.din(n24455));
	jspl jspl_w_n24456_0(.douta(w_n24456_0[0]),.doutb(w_n24456_0[1]),.din(n24456));
	jspl jspl_w_n24460_0(.douta(w_n24460_0[0]),.doutb(w_n24460_0[1]),.din(n24460));
	jspl jspl_w_n24461_0(.douta(w_n24461_0[0]),.doutb(w_n24461_0[1]),.din(n24461));
	jspl3 jspl3_w_n24463_0(.douta(w_n24463_0[0]),.doutb(w_n24463_0[1]),.doutc(w_n24463_0[2]),.din(n24463));
	jspl jspl_w_n24464_0(.douta(w_n24464_0[0]),.doutb(w_n24464_0[1]),.din(n24464));
	jspl jspl_w_n24468_0(.douta(w_n24468_0[0]),.doutb(w_n24468_0[1]),.din(n24468));
	jspl jspl_w_n24469_0(.douta(w_n24469_0[0]),.doutb(w_n24469_0[1]),.din(n24469));
	jspl3 jspl3_w_n24471_0(.douta(w_n24471_0[0]),.doutb(w_n24471_0[1]),.doutc(w_n24471_0[2]),.din(n24471));
	jspl jspl_w_n24472_0(.douta(w_n24472_0[0]),.doutb(w_n24472_0[1]),.din(n24472));
	jspl jspl_w_n24476_0(.douta(w_n24476_0[0]),.doutb(w_n24476_0[1]),.din(n24476));
	jspl jspl_w_n24477_0(.douta(w_n24477_0[0]),.doutb(w_n24477_0[1]),.din(n24477));
	jspl3 jspl3_w_n24479_0(.douta(w_n24479_0[0]),.doutb(w_n24479_0[1]),.doutc(w_n24479_0[2]),.din(n24479));
	jspl jspl_w_n24480_0(.douta(w_n24480_0[0]),.doutb(w_n24480_0[1]),.din(n24480));
	jspl jspl_w_n24484_0(.douta(w_n24484_0[0]),.doutb(w_n24484_0[1]),.din(n24484));
	jspl jspl_w_n24485_0(.douta(w_n24485_0[0]),.doutb(w_n24485_0[1]),.din(n24485));
	jspl3 jspl3_w_n24487_0(.douta(w_n24487_0[0]),.doutb(w_n24487_0[1]),.doutc(w_n24487_0[2]),.din(n24487));
	jspl jspl_w_n24488_0(.douta(w_n24488_0[0]),.doutb(w_n24488_0[1]),.din(n24488));
	jspl jspl_w_n24492_0(.douta(w_n24492_0[0]),.doutb(w_n24492_0[1]),.din(n24492));
	jspl jspl_w_n24493_0(.douta(w_n24493_0[0]),.doutb(w_n24493_0[1]),.din(n24493));
	jspl3 jspl3_w_n24495_0(.douta(w_n24495_0[0]),.doutb(w_n24495_0[1]),.doutc(w_n24495_0[2]),.din(n24495));
	jspl jspl_w_n24496_0(.douta(w_n24496_0[0]),.doutb(w_n24496_0[1]),.din(n24496));
	jspl3 jspl3_w_n24500_0(.douta(w_n24500_0[0]),.doutb(w_n24500_0[1]),.doutc(w_n24500_0[2]),.din(n24500));
	jspl3 jspl3_w_n24502_0(.douta(w_n24502_0[0]),.doutb(w_n24502_0[1]),.doutc(w_n24502_0[2]),.din(n24502));
	jspl jspl_w_n24503_0(.douta(w_n24503_0[0]),.doutb(w_n24503_0[1]),.din(n24503));
	jspl jspl_w_n24507_0(.douta(w_n24507_0[0]),.doutb(w_n24507_0[1]),.din(n24507));
	jspl jspl_w_n24508_0(.douta(w_n24508_0[0]),.doutb(w_n24508_0[1]),.din(n24508));
	jspl3 jspl3_w_n24510_0(.douta(w_n24510_0[0]),.doutb(w_n24510_0[1]),.doutc(w_n24510_0[2]),.din(n24510));
	jspl jspl_w_n24511_0(.douta(w_n24511_0[0]),.doutb(w_n24511_0[1]),.din(n24511));
	jspl3 jspl3_w_n24515_0(.douta(w_n24515_0[0]),.doutb(w_n24515_0[1]),.doutc(w_n24515_0[2]),.din(n24515));
	jspl3 jspl3_w_n24517_0(.douta(w_n24517_0[0]),.doutb(w_n24517_0[1]),.doutc(w_n24517_0[2]),.din(n24517));
	jspl jspl_w_n24518_0(.douta(w_n24518_0[0]),.doutb(w_n24518_0[1]),.din(n24518));
	jspl jspl_w_n24522_0(.douta(w_n24522_0[0]),.doutb(w_n24522_0[1]),.din(n24522));
	jspl jspl_w_n24523_0(.douta(w_n24523_0[0]),.doutb(w_n24523_0[1]),.din(n24523));
	jspl3 jspl3_w_n24525_0(.douta(w_n24525_0[0]),.doutb(w_n24525_0[1]),.doutc(w_n24525_0[2]),.din(n24525));
	jspl jspl_w_n24526_0(.douta(w_n24526_0[0]),.doutb(w_n24526_0[1]),.din(n24526));
	jspl3 jspl3_w_n24530_0(.douta(w_n24530_0[0]),.doutb(w_n24530_0[1]),.doutc(w_n24530_0[2]),.din(n24530));
	jspl3 jspl3_w_n24532_0(.douta(w_n24532_0[0]),.doutb(w_n24532_0[1]),.doutc(w_n24532_0[2]),.din(n24532));
	jspl jspl_w_n24533_0(.douta(w_n24533_0[0]),.doutb(w_n24533_0[1]),.din(n24533));
	jspl3 jspl3_w_n24537_0(.douta(w_n24537_0[0]),.doutb(w_n24537_0[1]),.doutc(w_n24537_0[2]),.din(n24537));
	jspl3 jspl3_w_n24539_0(.douta(w_n24539_0[0]),.doutb(w_n24539_0[1]),.doutc(w_n24539_0[2]),.din(n24539));
	jspl jspl_w_n24540_0(.douta(w_n24540_0[0]),.doutb(w_n24540_0[1]),.din(n24540));
	jspl3 jspl3_w_n24544_0(.douta(w_n24544_0[0]),.doutb(w_n24544_0[1]),.doutc(w_n24544_0[2]),.din(n24544));
	jspl3 jspl3_w_n24546_0(.douta(w_n24546_0[0]),.doutb(w_n24546_0[1]),.doutc(w_n24546_0[2]),.din(n24546));
	jspl jspl_w_n24547_0(.douta(w_n24547_0[0]),.doutb(w_n24547_0[1]),.din(n24547));
	jspl jspl_w_n24551_0(.douta(w_n24551_0[0]),.doutb(w_n24551_0[1]),.din(n24551));
	jspl jspl_w_n24552_0(.douta(w_n24552_0[0]),.doutb(w_n24552_0[1]),.din(n24552));
	jspl3 jspl3_w_n24554_0(.douta(w_n24554_0[0]),.doutb(w_n24554_0[1]),.doutc(w_n24554_0[2]),.din(n24554));
	jspl jspl_w_n24555_0(.douta(w_n24555_0[0]),.doutb(w_n24555_0[1]),.din(n24555));
	jspl jspl_w_n24830_0(.douta(w_n24830_0[0]),.doutb(w_n24830_0[1]),.din(n24830));
	jspl jspl_w_n24831_0(.douta(w_n24831_0[0]),.doutb(w_n24831_0[1]),.din(n24831));
	jspl jspl_w_n24834_0(.douta(w_n24834_0[0]),.doutb(w_n24834_0[1]),.din(n24834));
	jspl3 jspl3_w_n24835_0(.douta(w_n24835_0[0]),.doutb(w_n24835_0[1]),.doutc(w_n24835_0[2]),.din(n24835));
	jspl jspl_w_n24836_0(.douta(w_n24836_0[0]),.doutb(w_n24836_0[1]),.din(n24836));
	jspl jspl_w_n24839_0(.douta(w_n24839_0[0]),.doutb(w_n24839_0[1]),.din(n24839));
	jspl jspl_w_n24845_0(.douta(w_n24845_0[0]),.doutb(w_n24845_0[1]),.din(n24845));
	jspl jspl_w_n24852_0(.douta(w_n24852_0[0]),.doutb(w_n24852_0[1]),.din(n24852));
	jspl3 jspl3_w_n24856_0(.douta(w_n24856_0[0]),.doutb(w_n24856_0[1]),.doutc(w_n24856_0[2]),.din(n24856));
	jspl3 jspl3_w_n24856_1(.douta(w_n24856_1[0]),.doutb(w_n24856_1[1]),.doutc(w_n24856_1[2]),.din(w_n24856_0[0]));
	jspl3 jspl3_w_n24856_2(.douta(w_n24856_2[0]),.doutb(w_n24856_2[1]),.doutc(w_n24856_2[2]),.din(w_n24856_0[1]));
	jspl3 jspl3_w_n24856_3(.douta(w_n24856_3[0]),.doutb(w_n24856_3[1]),.doutc(w_n24856_3[2]),.din(w_n24856_0[2]));
	jspl3 jspl3_w_n24856_4(.douta(w_n24856_4[0]),.doutb(w_n24856_4[1]),.doutc(w_n24856_4[2]),.din(w_n24856_1[0]));
	jspl3 jspl3_w_n24856_5(.douta(w_n24856_5[0]),.doutb(w_n24856_5[1]),.doutc(w_n24856_5[2]),.din(w_n24856_1[1]));
	jspl3 jspl3_w_n24856_6(.douta(w_n24856_6[0]),.doutb(w_n24856_6[1]),.doutc(w_n24856_6[2]),.din(w_n24856_1[2]));
	jspl3 jspl3_w_n24856_7(.douta(w_n24856_7[0]),.doutb(w_n24856_7[1]),.doutc(w_n24856_7[2]),.din(w_n24856_2[0]));
	jspl3 jspl3_w_n24856_8(.douta(w_n24856_8[0]),.doutb(w_n24856_8[1]),.doutc(w_n24856_8[2]),.din(w_n24856_2[1]));
	jspl3 jspl3_w_n24856_9(.douta(w_n24856_9[0]),.doutb(w_n24856_9[1]),.doutc(w_n24856_9[2]),.din(w_n24856_2[2]));
	jspl3 jspl3_w_n24856_10(.douta(w_n24856_10[0]),.doutb(w_n24856_10[1]),.doutc(w_n24856_10[2]),.din(w_n24856_3[0]));
	jspl3 jspl3_w_n24856_11(.douta(w_n24856_11[0]),.doutb(w_n24856_11[1]),.doutc(w_n24856_11[2]),.din(w_n24856_3[1]));
	jspl3 jspl3_w_n24856_12(.douta(w_n24856_12[0]),.doutb(w_n24856_12[1]),.doutc(w_n24856_12[2]),.din(w_n24856_3[2]));
	jspl3 jspl3_w_n24856_13(.douta(w_n24856_13[0]),.doutb(w_n24856_13[1]),.doutc(w_n24856_13[2]),.din(w_n24856_4[0]));
	jspl3 jspl3_w_n24856_14(.douta(w_n24856_14[0]),.doutb(w_n24856_14[1]),.doutc(w_n24856_14[2]),.din(w_n24856_4[1]));
	jspl3 jspl3_w_n24856_15(.douta(w_n24856_15[0]),.doutb(w_n24856_15[1]),.doutc(w_n24856_15[2]),.din(w_n24856_4[2]));
	jspl3 jspl3_w_n24856_16(.douta(w_n24856_16[0]),.doutb(w_n24856_16[1]),.doutc(w_n24856_16[2]),.din(w_n24856_5[0]));
	jspl3 jspl3_w_n24856_17(.douta(w_n24856_17[0]),.doutb(w_n24856_17[1]),.doutc(w_n24856_17[2]),.din(w_n24856_5[1]));
	jspl3 jspl3_w_n24856_18(.douta(w_n24856_18[0]),.doutb(w_n24856_18[1]),.doutc(w_n24856_18[2]),.din(w_n24856_5[2]));
	jspl3 jspl3_w_n24856_19(.douta(w_n24856_19[0]),.doutb(w_n24856_19[1]),.doutc(w_n24856_19[2]),.din(w_n24856_6[0]));
	jspl3 jspl3_w_n24856_20(.douta(w_n24856_20[0]),.doutb(w_n24856_20[1]),.doutc(w_n24856_20[2]),.din(w_n24856_6[1]));
	jspl3 jspl3_w_n24856_21(.douta(w_n24856_21[0]),.doutb(w_n24856_21[1]),.doutc(w_n24856_21[2]),.din(w_n24856_6[2]));
	jspl3 jspl3_w_n24856_22(.douta(w_n24856_22[0]),.doutb(w_n24856_22[1]),.doutc(w_n24856_22[2]),.din(w_n24856_7[0]));
	jspl3 jspl3_w_n24856_23(.douta(w_n24856_23[0]),.doutb(w_n24856_23[1]),.doutc(w_n24856_23[2]),.din(w_n24856_7[1]));
	jspl3 jspl3_w_n24856_24(.douta(w_n24856_24[0]),.doutb(w_n24856_24[1]),.doutc(w_n24856_24[2]),.din(w_n24856_7[2]));
	jspl3 jspl3_w_n24856_25(.douta(w_n24856_25[0]),.doutb(w_n24856_25[1]),.doutc(w_n24856_25[2]),.din(w_n24856_8[0]));
	jspl3 jspl3_w_n24856_26(.douta(w_n24856_26[0]),.doutb(w_n24856_26[1]),.doutc(w_n24856_26[2]),.din(w_n24856_8[1]));
	jspl3 jspl3_w_n24856_27(.douta(w_n24856_27[0]),.doutb(w_n24856_27[1]),.doutc(w_n24856_27[2]),.din(w_n24856_8[2]));
	jspl3 jspl3_w_n24856_28(.douta(w_n24856_28[0]),.doutb(w_n24856_28[1]),.doutc(w_n24856_28[2]),.din(w_n24856_9[0]));
	jspl3 jspl3_w_n24856_29(.douta(w_n24856_29[0]),.doutb(w_n24856_29[1]),.doutc(w_n24856_29[2]),.din(w_n24856_9[1]));
	jspl3 jspl3_w_n24856_30(.douta(w_n24856_30[0]),.doutb(w_n24856_30[1]),.doutc(w_n24856_30[2]),.din(w_n24856_9[2]));
	jspl jspl_w_n24859_0(.douta(w_n24859_0[0]),.doutb(w_n24859_0[1]),.din(n24859));
	jspl jspl_w_n24863_0(.douta(w_n24863_0[0]),.doutb(w_n24863_0[1]),.din(n24863));
	jspl jspl_w_n24867_0(.douta(w_n24867_0[0]),.doutb(w_n24867_0[1]),.din(n24867));
	jspl jspl_w_n24873_0(.douta(w_n24873_0[0]),.doutb(w_n24873_0[1]),.din(n24873));
	jspl jspl_w_n24877_0(.douta(w_n24877_0[0]),.doutb(w_n24877_0[1]),.din(n24877));
	jspl jspl_w_n24881_0(.douta(w_n24881_0[0]),.doutb(w_n24881_0[1]),.din(n24881));
	jspl jspl_w_n24885_0(.douta(w_n24885_0[0]),.doutb(w_n24885_0[1]),.din(n24885));
	jspl jspl_w_n24889_0(.douta(w_n24889_0[0]),.doutb(w_n24889_0[1]),.din(n24889));
	jspl jspl_w_n24893_0(.douta(w_n24893_0[0]),.doutb(w_n24893_0[1]),.din(n24893));
	jspl jspl_w_n24897_0(.douta(w_n24897_0[0]),.doutb(w_n24897_0[1]),.din(n24897));
	jspl jspl_w_n24901_0(.douta(w_n24901_0[0]),.doutb(w_n24901_0[1]),.din(n24901));
	jspl jspl_w_n24905_0(.douta(w_n24905_0[0]),.doutb(w_n24905_0[1]),.din(n24905));
	jspl jspl_w_n24909_0(.douta(w_n24909_0[0]),.doutb(w_n24909_0[1]),.din(n24909));
	jspl jspl_w_n24913_0(.douta(w_n24913_0[0]),.doutb(w_n24913_0[1]),.din(n24913));
	jspl jspl_w_n24917_0(.douta(w_n24917_0[0]),.doutb(w_n24917_0[1]),.din(n24917));
	jspl jspl_w_n24921_0(.douta(w_n24921_0[0]),.doutb(w_n24921_0[1]),.din(n24921));
	jspl jspl_w_n24925_0(.douta(w_n24925_0[0]),.doutb(w_n24925_0[1]),.din(n24925));
	jspl jspl_w_n24929_0(.douta(w_n24929_0[0]),.doutb(w_n24929_0[1]),.din(n24929));
	jspl jspl_w_n24933_0(.douta(w_n24933_0[0]),.doutb(w_n24933_0[1]),.din(n24933));
	jspl jspl_w_n24937_0(.douta(w_n24937_0[0]),.doutb(w_n24937_0[1]),.din(n24937));
	jspl jspl_w_n24941_0(.douta(w_n24941_0[0]),.doutb(w_n24941_0[1]),.din(n24941));
	jspl jspl_w_n24945_0(.douta(w_n24945_0[0]),.doutb(w_n24945_0[1]),.din(n24945));
	jspl jspl_w_n24949_0(.douta(w_n24949_0[0]),.doutb(w_n24949_0[1]),.din(n24949));
	jspl jspl_w_n24953_0(.douta(w_n24953_0[0]),.doutb(w_n24953_0[1]),.din(n24953));
	jspl jspl_w_n24958_0(.douta(w_n24958_0[0]),.doutb(w_n24958_0[1]),.din(n24958));
	jspl jspl_w_n24962_0(.douta(w_n24962_0[0]),.doutb(w_n24962_0[1]),.din(n24962));
	jspl jspl_w_n24966_0(.douta(w_n24966_0[0]),.doutb(w_n24966_0[1]),.din(n24966));
	jspl jspl_w_n24968_0(.douta(w_n24968_0[0]),.doutb(w_n24968_0[1]),.din(n24968));
	jspl jspl_w_n24971_0(.douta(w_n24971_0[0]),.doutb(w_n24971_0[1]),.din(n24971));
	jspl jspl_w_n24977_0(.douta(w_n24977_0[0]),.doutb(w_n24977_0[1]),.din(n24977));
	jspl jspl_w_n24988_0(.douta(w_n24988_0[0]),.doutb(w_n24988_0[1]),.din(n24988));
	jspl jspl_w_n24995_0(.douta(w_n24995_0[0]),.doutb(w_n24995_0[1]),.din(n24995));
	jspl jspl_w_n25014_0(.douta(w_n25014_0[0]),.doutb(w_n25014_0[1]),.din(n25014));
	jspl jspl_w_n25021_0(.douta(w_n25021_0[0]),.doutb(w_n25021_0[1]),.din(n25021));
	jspl jspl_w_n25037_0(.douta(w_n25037_0[0]),.doutb(w_n25037_0[1]),.din(n25037));
	jspl jspl_w_n25050_0(.douta(w_n25050_0[0]),.doutb(w_n25050_0[1]),.din(n25050));
	jspl jspl_w_n25057_0(.douta(w_n25057_0[0]),.doutb(w_n25057_0[1]),.din(n25057));
	jspl jspl_w_n25070_0(.douta(w_n25070_0[0]),.doutb(w_n25070_0[1]),.din(n25070));
	jspl jspl_w_n25083_0(.douta(w_n25083_0[0]),.doutb(w_n25083_0[1]),.din(n25083));
	jspl jspl_w_n25090_0(.douta(w_n25090_0[0]),.doutb(w_n25090_0[1]),.din(n25090));
	jspl jspl_w_n25097_0(.douta(w_n25097_0[0]),.doutb(w_n25097_0[1]),.din(n25097));
	jspl jspl_w_n25113_0(.douta(w_n25113_0[0]),.doutb(w_n25113_0[1]),.din(n25113));
	jspl jspl_w_n25119_0(.douta(w_n25119_0[0]),.doutb(w_n25119_0[1]),.din(n25119));
	jspl jspl_w_n25130_0(.douta(w_n25130_0[0]),.doutb(w_n25130_0[1]),.din(n25130));
	jspl jspl_w_n25137_0(.douta(w_n25137_0[0]),.doutb(w_n25137_0[1]),.din(n25137));
	jspl jspl_w_n25143_0(.douta(w_n25143_0[0]),.doutb(w_n25143_0[1]),.din(n25143));
	jspl jspl_w_n25151_0(.douta(w_n25151_0[0]),.doutb(w_n25151_0[1]),.din(n25151));
	jspl jspl_w_n25164_0(.douta(w_n25164_0[0]),.doutb(w_n25164_0[1]),.din(n25164));
	jspl jspl_w_n25171_0(.douta(w_n25171_0[0]),.doutb(w_n25171_0[1]),.din(n25171));
	jspl jspl_w_n25178_0(.douta(w_n25178_0[0]),.doutb(w_n25178_0[1]),.din(n25178));
	jspl jspl_w_n25189_0(.douta(w_n25189_0[0]),.doutb(w_n25189_0[1]),.din(n25189));
	jspl jspl_w_n25195_0(.douta(w_n25195_0[0]),.doutb(w_n25195_0[1]),.din(n25195));
	jspl jspl_w_n25208_0(.douta(w_n25208_0[0]),.doutb(w_n25208_0[1]),.din(n25208));
	jspl jspl_w_n25215_0(.douta(w_n25215_0[0]),.doutb(w_n25215_0[1]),.din(n25215));
	jspl jspl_w_n25222_0(.douta(w_n25222_0[0]),.doutb(w_n25222_0[1]),.din(n25222));
	jspl jspl_w_n25235_0(.douta(w_n25235_0[0]),.doutb(w_n25235_0[1]),.din(n25235));
	jspl jspl_w_n25246_0(.douta(w_n25246_0[0]),.doutb(w_n25246_0[1]),.din(n25246));
	jspl jspl_w_n25253_0(.douta(w_n25253_0[0]),.doutb(w_n25253_0[1]),.din(n25253));
	jspl jspl_w_n25260_0(.douta(w_n25260_0[0]),.doutb(w_n25260_0[1]),.din(n25260));
	jspl jspl_w_n25267_0(.douta(w_n25267_0[0]),.doutb(w_n25267_0[1]),.din(n25267));
	jspl jspl_w_n25273_0(.douta(w_n25273_0[0]),.doutb(w_n25273_0[1]),.din(n25273));
	jspl jspl_w_n25281_0(.douta(w_n25281_0[0]),.doutb(w_n25281_0[1]),.din(n25281));
	jspl jspl_w_n25292_0(.douta(w_n25292_0[0]),.doutb(w_n25292_0[1]),.din(n25292));
endmodule

