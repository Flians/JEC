/*

c6288:
	jxor: 446
	jspl: 940
	jspl3: 260
	jcb: 331
	jnot: 330
	jdff: 5481
	jand: 683

Summary:
	jxor: 446
	jspl: 940
	jspl3: 260
	jcb: 331
	jnot: 330
	jdff: 5481
	jand: 683
*/

module c6288(gclk, G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat, G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat, G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat, G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat, G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat, G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat, G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat, G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat, G6270gat, G6280gat, G6287gat, G6288gat);
	input gclk;
	input G1gat;
	input G18gat;
	input G35gat;
	input G52gat;
	input G69gat;
	input G86gat;
	input G103gat;
	input G120gat;
	input G137gat;
	input G154gat;
	input G171gat;
	input G188gat;
	input G205gat;
	input G222gat;
	input G239gat;
	input G256gat;
	input G273gat;
	input G290gat;
	input G307gat;
	input G324gat;
	input G341gat;
	input G358gat;
	input G375gat;
	input G392gat;
	input G409gat;
	input G426gat;
	input G443gat;
	input G460gat;
	input G477gat;
	input G494gat;
	input G511gat;
	input G528gat;
	output G545gat;
	output G1581gat;
	output G1901gat;
	output G2223gat;
	output G2548gat;
	output G2877gat;
	output G3211gat;
	output G3552gat;
	output G3895gat;
	output G4241gat;
	output G4591gat;
	output G4946gat;
	output G5308gat;
	output G5672gat;
	output G5971gat;
	output G6123gat;
	output G6150gat;
	output G6160gat;
	output G6170gat;
	output G6180gat;
	output G6190gat;
	output G6200gat;
	output G6210gat;
	output G6220gat;
	output G6230gat;
	output G6240gat;
	output G6250gat;
	output G6260gat;
	output G6270gat;
	output G6280gat;
	output G6287gat;
	output G6288gat;
	wire n65;
	wire n66;
	wire n67;
	wire n68;
	wire n69;
	wire n70;
	wire n72;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n177;
	wire n178;
	wire n179;
	wire n180;
	wire n181;
	wire n183;
	wire n184;
	wire n185;
	wire n186;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n192;
	wire n193;
	wire n194;
	wire n195;
	wire n196;
	wire n197;
	wire n198;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n204;
	wire n205;
	wire n206;
	wire n207;
	wire n208;
	wire n209;
	wire n210;
	wire n211;
	wire n212;
	wire n213;
	wire n214;
	wire n215;
	wire n216;
	wire n217;
	wire n218;
	wire n219;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n232;
	wire n233;
	wire n234;
	wire n235;
	wire n236;
	wire n237;
	wire n238;
	wire n239;
	wire n240;
	wire n241;
	wire n242;
	wire n243;
	wire n244;
	wire n245;
	wire n246;
	wire n247;
	wire n248;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n253;
	wire n254;
	wire n255;
	wire n256;
	wire n257;
	wire n258;
	wire n259;
	wire n260;
	wire n261;
	wire n262;
	wire n263;
	wire n264;
	wire n265;
	wire n266;
	wire n267;
	wire n268;
	wire n269;
	wire n270;
	wire n271;
	wire n272;
	wire n273;
	wire n274;
	wire n275;
	wire n277;
	wire n278;
	wire n279;
	wire n280;
	wire n281;
	wire n282;
	wire n283;
	wire n284;
	wire n285;
	wire n286;
	wire n287;
	wire n288;
	wire n289;
	wire n290;
	wire n291;
	wire n292;
	wire n293;
	wire n294;
	wire n295;
	wire n296;
	wire n297;
	wire n298;
	wire n299;
	wire n300;
	wire n301;
	wire n302;
	wire n303;
	wire n304;
	wire n305;
	wire n306;
	wire n307;
	wire n308;
	wire n309;
	wire n310;
	wire n311;
	wire n312;
	wire n313;
	wire n314;
	wire n315;
	wire n316;
	wire n317;
	wire n318;
	wire n319;
	wire n320;
	wire n321;
	wire n322;
	wire n323;
	wire n324;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n331;
	wire n332;
	wire n333;
	wire n335;
	wire n336;
	wire n337;
	wire n338;
	wire n339;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n344;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n349;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n354;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n359;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n448;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n555;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n608;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n653;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n662;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n672;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n710;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n743;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n757;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n770;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n778;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n790;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n805;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n815;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n827;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n838;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n851;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n868;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n875;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n888;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n899;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n915;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n927;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n966;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n983;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n997;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1011;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1020;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1029;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1047;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1054;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1061;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1068;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1075;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1083;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1091;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1099;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1107;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1115;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1123;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1131;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1139;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1156;
	wire n1157;
	wire n1158;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1164;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1170;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1176;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1183;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1191;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1198;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1206;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1212;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1219;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1226;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1233;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1241;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1250;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1259;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1266;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1273;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1280;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1288;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1296;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1304;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1312;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1320;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1336;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1344;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1387;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1453;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1598;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1616;
	wire n1617;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1623;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1640;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire n1652;
	wire n1653;
	wire n1654;
	wire n1655;
	wire n1656;
	wire n1657;
	wire n1658;
	wire n1659;
	wire n1660;
	wire n1661;
	wire n1662;
	wire n1663;
	wire n1664;
	wire n1665;
	wire n1666;
	wire n1667;
	wire n1668;
	wire n1669;
	wire n1670;
	wire n1671;
	wire n1672;
	wire n1674;
	wire n1675;
	wire n1676;
	wire n1677;
	wire n1678;
	wire n1679;
	wire n1680;
	wire n1681;
	wire n1682;
	wire n1683;
	wire n1684;
	wire n1685;
	wire n1686;
	wire n1687;
	wire n1688;
	wire n1689;
	wire n1690;
	wire n1691;
	wire n1692;
	wire n1693;
	wire n1694;
	wire n1695;
	wire n1696;
	wire n1697;
	wire n1698;
	wire n1699;
	wire n1700;
	wire n1701;
	wire n1702;
	wire n1703;
	wire n1704;
	wire n1705;
	wire n1706;
	wire n1707;
	wire n1708;
	wire n1709;
	wire n1710;
	wire n1711;
	wire n1712;
	wire n1713;
	wire n1714;
	wire n1715;
	wire n1716;
	wire n1717;
	wire n1718;
	wire n1719;
	wire n1720;
	wire n1722;
	wire n1723;
	wire n1724;
	wire n1725;
	wire n1726;
	wire n1727;
	wire n1728;
	wire n1729;
	wire n1730;
	wire n1731;
	wire n1732;
	wire n1733;
	wire n1734;
	wire n1735;
	wire n1736;
	wire n1737;
	wire n1738;
	wire n1739;
	wire n1740;
	wire n1741;
	wire n1742;
	wire n1743;
	wire n1744;
	wire n1745;
	wire n1746;
	wire n1747;
	wire n1748;
	wire n1749;
	wire n1750;
	wire n1751;
	wire n1752;
	wire n1753;
	wire n1754;
	wire n1755;
	wire n1756;
	wire n1757;
	wire n1758;
	wire n1760;
	wire n1761;
	wire n1762;
	wire n1763;
	wire n1764;
	wire n1765;
	wire n1766;
	wire n1767;
	wire n1768;
	wire n1769;
	wire n1770;
	wire n1771;
	wire n1772;
	wire n1773;
	wire n1774;
	wire n1775;
	wire n1776;
	wire n1777;
	wire n1778;
	wire n1779;
	wire n1780;
	wire n1781;
	wire n1782;
	wire n1783;
	wire n1784;
	wire n1785;
	wire n1786;
	wire n1787;
	wire n1788;
	wire n1789;
	wire n1790;
	wire n1791;
	wire n1793;
	wire n1794;
	wire n1795;
	wire n1796;
	wire n1797;
	wire n1798;
	wire n1799;
	wire n1800;
	wire n1801;
	wire n1802;
	wire n1803;
	wire n1804;
	wire n1805;
	wire n1806;
	wire n1807;
	wire n1808;
	wire n1809;
	wire n1810;
	wire n1811;
	wire n1812;
	wire n1813;
	wire n1814;
	wire n1815;
	wire n1816;
	wire n1817;
	wire n1819;
	wire n1820;
	wire n1821;
	wire n1822;
	wire n1823;
	wire n1824;
	wire n1825;
	wire n1826;
	wire n1827;
	wire n1828;
	wire n1829;
	wire n1830;
	wire n1831;
	wire n1832;
	wire n1833;
	wire n1834;
	wire n1835;
	wire n1836;
	wire n1838;
	wire n1839;
	wire n1840;
	wire n1841;
	wire n1842;
	wire n1843;
	wire n1844;
	wire n1845;
	wire n1846;
	wire n1847;
	wire n1848;
	wire n1849;
	wire n1850;
	wire n1851;
	wire [2:0] w_G1gat_0;
	wire [2:0] w_G1gat_1;
	wire [2:0] w_G1gat_2;
	wire [2:0] w_G1gat_3;
	wire [2:0] w_G1gat_4;
	wire [2:0] w_G1gat_5;
	wire [2:0] w_G1gat_6;
	wire [1:0] w_G1gat_7;
	wire [2:0] w_G18gat_0;
	wire [2:0] w_G18gat_1;
	wire [2:0] w_G18gat_2;
	wire [2:0] w_G18gat_3;
	wire [2:0] w_G18gat_4;
	wire [2:0] w_G18gat_5;
	wire [2:0] w_G18gat_6;
	wire [2:0] w_G18gat_7;
	wire [2:0] w_G35gat_0;
	wire [2:0] w_G35gat_1;
	wire [2:0] w_G35gat_2;
	wire [2:0] w_G35gat_3;
	wire [2:0] w_G35gat_4;
	wire [2:0] w_G35gat_5;
	wire [2:0] w_G35gat_6;
	wire [2:0] w_G35gat_7;
	wire [2:0] w_G52gat_0;
	wire [2:0] w_G52gat_1;
	wire [2:0] w_G52gat_2;
	wire [2:0] w_G52gat_3;
	wire [2:0] w_G52gat_4;
	wire [2:0] w_G52gat_5;
	wire [2:0] w_G52gat_6;
	wire [2:0] w_G52gat_7;
	wire [2:0] w_G69gat_0;
	wire [2:0] w_G69gat_1;
	wire [2:0] w_G69gat_2;
	wire [2:0] w_G69gat_3;
	wire [2:0] w_G69gat_4;
	wire [2:0] w_G69gat_5;
	wire [2:0] w_G69gat_6;
	wire [1:0] w_G69gat_7;
	wire [2:0] w_G86gat_0;
	wire [2:0] w_G86gat_1;
	wire [2:0] w_G86gat_2;
	wire [2:0] w_G86gat_3;
	wire [2:0] w_G86gat_4;
	wire [2:0] w_G86gat_5;
	wire [2:0] w_G86gat_6;
	wire [1:0] w_G86gat_7;
	wire [2:0] w_G103gat_0;
	wire [2:0] w_G103gat_1;
	wire [2:0] w_G103gat_2;
	wire [2:0] w_G103gat_3;
	wire [2:0] w_G103gat_4;
	wire [2:0] w_G103gat_5;
	wire [2:0] w_G103gat_6;
	wire [1:0] w_G103gat_7;
	wire [2:0] w_G120gat_0;
	wire [2:0] w_G120gat_1;
	wire [2:0] w_G120gat_2;
	wire [2:0] w_G120gat_3;
	wire [2:0] w_G120gat_4;
	wire [2:0] w_G120gat_5;
	wire [2:0] w_G120gat_6;
	wire [1:0] w_G120gat_7;
	wire [2:0] w_G137gat_0;
	wire [2:0] w_G137gat_1;
	wire [2:0] w_G137gat_2;
	wire [2:0] w_G137gat_3;
	wire [2:0] w_G137gat_4;
	wire [2:0] w_G137gat_5;
	wire [2:0] w_G137gat_6;
	wire [1:0] w_G137gat_7;
	wire [2:0] w_G154gat_0;
	wire [2:0] w_G154gat_1;
	wire [2:0] w_G154gat_2;
	wire [2:0] w_G154gat_3;
	wire [2:0] w_G154gat_4;
	wire [2:0] w_G154gat_5;
	wire [2:0] w_G154gat_6;
	wire [1:0] w_G154gat_7;
	wire [2:0] w_G171gat_0;
	wire [2:0] w_G171gat_1;
	wire [2:0] w_G171gat_2;
	wire [2:0] w_G171gat_3;
	wire [2:0] w_G171gat_4;
	wire [2:0] w_G171gat_5;
	wire [2:0] w_G171gat_6;
	wire [1:0] w_G171gat_7;
	wire [2:0] w_G188gat_0;
	wire [2:0] w_G188gat_1;
	wire [2:0] w_G188gat_2;
	wire [2:0] w_G188gat_3;
	wire [2:0] w_G188gat_4;
	wire [2:0] w_G188gat_5;
	wire [2:0] w_G188gat_6;
	wire [1:0] w_G188gat_7;
	wire [2:0] w_G205gat_0;
	wire [2:0] w_G205gat_1;
	wire [2:0] w_G205gat_2;
	wire [2:0] w_G205gat_3;
	wire [2:0] w_G205gat_4;
	wire [2:0] w_G205gat_5;
	wire [2:0] w_G205gat_6;
	wire [1:0] w_G205gat_7;
	wire [2:0] w_G222gat_0;
	wire [2:0] w_G222gat_1;
	wire [2:0] w_G222gat_2;
	wire [2:0] w_G222gat_3;
	wire [2:0] w_G222gat_4;
	wire [2:0] w_G222gat_5;
	wire [2:0] w_G222gat_6;
	wire [1:0] w_G222gat_7;
	wire [2:0] w_G239gat_0;
	wire [2:0] w_G239gat_1;
	wire [2:0] w_G239gat_2;
	wire [2:0] w_G239gat_3;
	wire [2:0] w_G239gat_4;
	wire [2:0] w_G239gat_5;
	wire [2:0] w_G239gat_6;
	wire [1:0] w_G239gat_7;
	wire [2:0] w_G256gat_0;
	wire [2:0] w_G256gat_1;
	wire [2:0] w_G256gat_2;
	wire [2:0] w_G256gat_3;
	wire [2:0] w_G256gat_4;
	wire [2:0] w_G256gat_5;
	wire [2:0] w_G256gat_6;
	wire [1:0] w_G256gat_7;
	wire [2:0] w_G273gat_0;
	wire [2:0] w_G273gat_1;
	wire [2:0] w_G273gat_2;
	wire [2:0] w_G273gat_3;
	wire [2:0] w_G273gat_4;
	wire [2:0] w_G273gat_5;
	wire [2:0] w_G273gat_6;
	wire [2:0] w_G273gat_7;
	wire [2:0] w_G290gat_0;
	wire [2:0] w_G290gat_1;
	wire [2:0] w_G290gat_2;
	wire [2:0] w_G290gat_3;
	wire [2:0] w_G290gat_4;
	wire [2:0] w_G290gat_5;
	wire [2:0] w_G290gat_6;
	wire [2:0] w_G290gat_7;
	wire [2:0] w_G307gat_0;
	wire [2:0] w_G307gat_1;
	wire [2:0] w_G307gat_2;
	wire [2:0] w_G307gat_3;
	wire [2:0] w_G307gat_4;
	wire [2:0] w_G307gat_5;
	wire [2:0] w_G307gat_6;
	wire [2:0] w_G307gat_7;
	wire [2:0] w_G324gat_0;
	wire [2:0] w_G324gat_1;
	wire [2:0] w_G324gat_2;
	wire [2:0] w_G324gat_3;
	wire [2:0] w_G324gat_4;
	wire [2:0] w_G324gat_5;
	wire [2:0] w_G324gat_6;
	wire [1:0] w_G324gat_7;
	wire [2:0] w_G341gat_0;
	wire [2:0] w_G341gat_1;
	wire [2:0] w_G341gat_2;
	wire [2:0] w_G341gat_3;
	wire [2:0] w_G341gat_4;
	wire [2:0] w_G341gat_5;
	wire [2:0] w_G341gat_6;
	wire [1:0] w_G341gat_7;
	wire [2:0] w_G358gat_0;
	wire [2:0] w_G358gat_1;
	wire [2:0] w_G358gat_2;
	wire [2:0] w_G358gat_3;
	wire [2:0] w_G358gat_4;
	wire [2:0] w_G358gat_5;
	wire [2:0] w_G358gat_6;
	wire [1:0] w_G358gat_7;
	wire [2:0] w_G375gat_0;
	wire [2:0] w_G375gat_1;
	wire [2:0] w_G375gat_2;
	wire [2:0] w_G375gat_3;
	wire [2:0] w_G375gat_4;
	wire [2:0] w_G375gat_5;
	wire [2:0] w_G375gat_6;
	wire [1:0] w_G375gat_7;
	wire [2:0] w_G392gat_0;
	wire [2:0] w_G392gat_1;
	wire [2:0] w_G392gat_2;
	wire [2:0] w_G392gat_3;
	wire [2:0] w_G392gat_4;
	wire [2:0] w_G392gat_5;
	wire [2:0] w_G392gat_6;
	wire [1:0] w_G392gat_7;
	wire [2:0] w_G409gat_0;
	wire [2:0] w_G409gat_1;
	wire [2:0] w_G409gat_2;
	wire [2:0] w_G409gat_3;
	wire [2:0] w_G409gat_4;
	wire [2:0] w_G409gat_5;
	wire [2:0] w_G409gat_6;
	wire [1:0] w_G409gat_7;
	wire [2:0] w_G426gat_0;
	wire [2:0] w_G426gat_1;
	wire [2:0] w_G426gat_2;
	wire [2:0] w_G426gat_3;
	wire [2:0] w_G426gat_4;
	wire [2:0] w_G426gat_5;
	wire [2:0] w_G426gat_6;
	wire [1:0] w_G426gat_7;
	wire [2:0] w_G443gat_0;
	wire [2:0] w_G443gat_1;
	wire [2:0] w_G443gat_2;
	wire [2:0] w_G443gat_3;
	wire [2:0] w_G443gat_4;
	wire [2:0] w_G443gat_5;
	wire [2:0] w_G443gat_6;
	wire [1:0] w_G443gat_7;
	wire [2:0] w_G460gat_0;
	wire [2:0] w_G460gat_1;
	wire [2:0] w_G460gat_2;
	wire [2:0] w_G460gat_3;
	wire [2:0] w_G460gat_4;
	wire [2:0] w_G460gat_5;
	wire [2:0] w_G460gat_6;
	wire [1:0] w_G460gat_7;
	wire [2:0] w_G477gat_0;
	wire [2:0] w_G477gat_1;
	wire [2:0] w_G477gat_2;
	wire [2:0] w_G477gat_3;
	wire [2:0] w_G477gat_4;
	wire [2:0] w_G477gat_5;
	wire [2:0] w_G477gat_6;
	wire [1:0] w_G477gat_7;
	wire [2:0] w_G494gat_0;
	wire [2:0] w_G494gat_1;
	wire [2:0] w_G494gat_2;
	wire [2:0] w_G494gat_3;
	wire [2:0] w_G494gat_4;
	wire [2:0] w_G494gat_5;
	wire [2:0] w_G494gat_6;
	wire [1:0] w_G494gat_7;
	wire [2:0] w_G511gat_0;
	wire [2:0] w_G511gat_1;
	wire [2:0] w_G511gat_2;
	wire [2:0] w_G511gat_3;
	wire [2:0] w_G511gat_4;
	wire [2:0] w_G511gat_5;
	wire [2:0] w_G511gat_6;
	wire [1:0] w_G511gat_7;
	wire [2:0] w_G528gat_0;
	wire [2:0] w_G528gat_1;
	wire [2:0] w_G528gat_2;
	wire [2:0] w_G528gat_3;
	wire [2:0] w_G528gat_4;
	wire [2:0] w_G528gat_5;
	wire [2:0] w_G528gat_6;
	wire [1:0] w_G528gat_7;
	wire w_G545gat_0;
	wire G545gat_fa_;
	wire [1:0] w_n65_0;
	wire [1:0] w_n69_0;
	wire [1:0] w_n70_0;
	wire [1:0] w_n72_0;
	wire [1:0] w_n75_0;
	wire [1:0] w_n77_0;
	wire [1:0] w_n78_0;
	wire [1:0] w_n81_0;
	wire [2:0] w_n82_0;
	wire [1:0] w_n82_1;
	wire [1:0] w_n84_0;
	wire [1:0] w_n85_0;
	wire [1:0] w_n87_0;
	wire [1:0] w_n89_0;
	wire [1:0] w_n93_0;
	wire [1:0] w_n94_0;
	wire [1:0] w_n96_0;
	wire [1:0] w_n99_0;
	wire [2:0] w_n100_0;
	wire [1:0] w_n100_1;
	wire [2:0] w_n101_0;
	wire [1:0] w_n103_0;
	wire [1:0] w_n104_0;
	wire [1:0] w_n107_0;
	wire [1:0] w_n108_0;
	wire [1:0] w_n110_0;
	wire [1:0] w_n115_0;
	wire [1:0] w_n116_0;
	wire [2:0] w_n126_0;
	wire [1:0] w_n128_0;
	wire [1:0] w_n129_0;
	wire [1:0] w_n130_0;
	wire [1:0] w_n131_0;
	wire [2:0] w_n132_0;
	wire [2:0] w_n133_0;
	wire [1:0] w_n138_0;
	wire [1:0] w_n139_0;
	wire [1:0] w_n140_0;
	wire [1:0] w_n142_0;
	wire [1:0] w_n143_0;
	wire [1:0] w_n145_0;
	wire [1:0] w_n150_0;
	wire [1:0] w_n151_0;
	wire [2:0] w_n156_0;
	wire [1:0] w_n158_0;
	wire [1:0] w_n163_0;
	wire [1:0] w_n165_0;
	wire [1:0] w_n166_0;
	wire [1:0] w_n168_0;
	wire [2:0] w_n169_0;
	wire [1:0] w_n170_0;
	wire [1:0] w_n172_0;
	wire [1:0] w_n174_0;
	wire [1:0] w_n175_0;
	wire [1:0] w_n176_0;
	wire [1:0] w_n177_0;
	wire [1:0] w_n178_0;
	wire [1:0] w_n180_0;
	wire [1:0] w_n181_0;
	wire [1:0] w_n183_0;
	wire [1:0] w_n188_0;
	wire [1:0] w_n189_0;
	wire [2:0] w_n194_0;
	wire [1:0] w_n196_0;
	wire [1:0] w_n199_0;
	wire [1:0] w_n201_0;
	wire [1:0] w_n204_0;
	wire [1:0] w_n206_0;
	wire [1:0] w_n207_0;
	wire [1:0] w_n209_0;
	wire [2:0] w_n210_0;
	wire [1:0] w_n210_1;
	wire [1:0] w_n213_0;
	wire [1:0] w_n215_0;
	wire [1:0] w_n216_0;
	wire [1:0] w_n217_0;
	wire [1:0] w_n218_0;
	wire [1:0] w_n219_0;
	wire [1:0] w_n220_0;
	wire [1:0] w_n221_0;
	wire [1:0] w_n223_0;
	wire [1:0] w_n224_0;
	wire [1:0] w_n226_0;
	wire [1:0] w_n231_0;
	wire [1:0] w_n232_0;
	wire [2:0] w_n237_0;
	wire [1:0] w_n239_0;
	wire [1:0] w_n242_0;
	wire [1:0] w_n244_0;
	wire [1:0] w_n247_0;
	wire [1:0] w_n249_0;
	wire [1:0] w_n252_0;
	wire [1:0] w_n254_0;
	wire [1:0] w_n255_0;
	wire [1:0] w_n257_0;
	wire [2:0] w_n258_0;
	wire [1:0] w_n259_0;
	wire [1:0] w_n261_0;
	wire [1:0] w_n264_0;
	wire [1:0] w_n265_0;
	wire [1:0] w_n266_0;
	wire [1:0] w_n267_0;
	wire [1:0] w_n268_0;
	wire [1:0] w_n269_0;
	wire [1:0] w_n270_0;
	wire [1:0] w_n271_0;
	wire [1:0] w_n272_0;
	wire [1:0] w_n274_0;
	wire [1:0] w_n275_0;
	wire [1:0] w_n277_0;
	wire [1:0] w_n282_0;
	wire [1:0] w_n283_0;
	wire [2:0] w_n288_0;
	wire [1:0] w_n290_0;
	wire [1:0] w_n293_0;
	wire [1:0] w_n295_0;
	wire [1:0] w_n298_0;
	wire [1:0] w_n300_0;
	wire [1:0] w_n303_0;
	wire [1:0] w_n305_0;
	wire [1:0] w_n308_0;
	wire [1:0] w_n310_0;
	wire [1:0] w_n311_0;
	wire [1:0] w_n313_0;
	wire [2:0] w_n314_0;
	wire [1:0] w_n315_0;
	wire [1:0] w_n317_0;
	wire [1:0] w_n320_0;
	wire [1:0] w_n321_0;
	wire [1:0] w_n322_0;
	wire [1:0] w_n323_0;
	wire [1:0] w_n324_0;
	wire [1:0] w_n325_0;
	wire [1:0] w_n326_0;
	wire [1:0] w_n327_0;
	wire [1:0] w_n328_0;
	wire [1:0] w_n329_0;
	wire [1:0] w_n330_0;
	wire [1:0] w_n332_0;
	wire [1:0] w_n333_0;
	wire [1:0] w_n335_0;
	wire [1:0] w_n340_0;
	wire [1:0] w_n341_0;
	wire [2:0] w_n346_0;
	wire [1:0] w_n348_0;
	wire [1:0] w_n351_0;
	wire [1:0] w_n353_0;
	wire [1:0] w_n356_0;
	wire [1:0] w_n358_0;
	wire [1:0] w_n361_0;
	wire [1:0] w_n363_0;
	wire [1:0] w_n366_0;
	wire [1:0] w_n368_0;
	wire [1:0] w_n371_0;
	wire [1:0] w_n372_0;
	wire [1:0] w_n373_0;
	wire [1:0] w_n375_0;
	wire [2:0] w_n376_0;
	wire [1:0] w_n377_0;
	wire [1:0] w_n380_0;
	wire [1:0] w_n382_0;
	wire [1:0] w_n383_0;
	wire [1:0] w_n384_0;
	wire [1:0] w_n385_0;
	wire [1:0] w_n386_0;
	wire [1:0] w_n387_0;
	wire [1:0] w_n388_0;
	wire [1:0] w_n389_0;
	wire [1:0] w_n390_0;
	wire [1:0] w_n391_0;
	wire [1:0] w_n392_0;
	wire [1:0] w_n393_0;
	wire [1:0] w_n394_0;
	wire [1:0] w_n396_0;
	wire [1:0] w_n397_0;
	wire [1:0] w_n399_0;
	wire [1:0] w_n404_0;
	wire [1:0] w_n405_0;
	wire [2:0] w_n410_0;
	wire [1:0] w_n412_0;
	wire [1:0] w_n415_0;
	wire [1:0] w_n417_0;
	wire [1:0] w_n420_0;
	wire [1:0] w_n422_0;
	wire [1:0] w_n425_0;
	wire [1:0] w_n427_0;
	wire [1:0] w_n430_0;
	wire [1:0] w_n432_0;
	wire [1:0] w_n435_0;
	wire [1:0] w_n437_0;
	wire [1:0] w_n441_0;
	wire [1:0] w_n442_0;
	wire [1:0] w_n443_0;
	wire [1:0] w_n445_0;
	wire [2:0] w_n446_0;
	wire [1:0] w_n447_0;
	wire [1:0] w_n450_0;
	wire [1:0] w_n452_0;
	wire [1:0] w_n453_0;
	wire [1:0] w_n454_0;
	wire [1:0] w_n455_0;
	wire [1:0] w_n456_0;
	wire [1:0] w_n457_0;
	wire [1:0] w_n458_0;
	wire [1:0] w_n459_0;
	wire [1:0] w_n460_0;
	wire [1:0] w_n461_0;
	wire [1:0] w_n462_0;
	wire [1:0] w_n463_0;
	wire [1:0] w_n464_0;
	wire [1:0] w_n465_0;
	wire [1:0] w_n466_0;
	wire [1:0] w_n468_0;
	wire [1:0] w_n469_0;
	wire [1:0] w_n471_0;
	wire [1:0] w_n476_0;
	wire [1:0] w_n477_0;
	wire [2:0] w_n482_0;
	wire [1:0] w_n484_0;
	wire [1:0] w_n487_0;
	wire [1:0] w_n489_0;
	wire [1:0] w_n492_0;
	wire [1:0] w_n494_0;
	wire [1:0] w_n497_0;
	wire [1:0] w_n499_0;
	wire [1:0] w_n502_0;
	wire [1:0] w_n504_0;
	wire [1:0] w_n507_0;
	wire [1:0] w_n509_0;
	wire [1:0] w_n512_0;
	wire [1:0] w_n514_0;
	wire [1:0] w_n518_0;
	wire [1:0] w_n519_0;
	wire [1:0] w_n520_0;
	wire [1:0] w_n522_0;
	wire [2:0] w_n523_0;
	wire [1:0] w_n524_0;
	wire [1:0] w_n527_0;
	wire [1:0] w_n529_0;
	wire [1:0] w_n530_0;
	wire [1:0] w_n531_0;
	wire [1:0] w_n532_0;
	wire [1:0] w_n533_0;
	wire [1:0] w_n534_0;
	wire [1:0] w_n535_0;
	wire [1:0] w_n536_0;
	wire [1:0] w_n537_0;
	wire [1:0] w_n538_0;
	wire [1:0] w_n539_0;
	wire [1:0] w_n540_0;
	wire [1:0] w_n541_0;
	wire [1:0] w_n542_0;
	wire [1:0] w_n543_0;
	wire [1:0] w_n544_0;
	wire [1:0] w_n545_0;
	wire [1:0] w_n547_0;
	wire [1:0] w_n548_0;
	wire [1:0] w_n550_0;
	wire [1:0] w_n555_0;
	wire [1:0] w_n556_0;
	wire [2:0] w_n561_0;
	wire [1:0] w_n563_0;
	wire [1:0] w_n566_0;
	wire [1:0] w_n568_0;
	wire [1:0] w_n571_0;
	wire [1:0] w_n573_0;
	wire [1:0] w_n576_0;
	wire [1:0] w_n578_0;
	wire [1:0] w_n581_0;
	wire [1:0] w_n583_0;
	wire [1:0] w_n586_0;
	wire [1:0] w_n588_0;
	wire [1:0] w_n591_0;
	wire [1:0] w_n593_0;
	wire [1:0] w_n596_0;
	wire [1:0] w_n598_0;
	wire [1:0] w_n602_0;
	wire [1:0] w_n603_0;
	wire [1:0] w_n604_0;
	wire [1:0] w_n606_0;
	wire [2:0] w_n607_0;
	wire [1:0] w_n608_0;
	wire [1:0] w_n611_0;
	wire [1:0] w_n613_0;
	wire [1:0] w_n614_0;
	wire [1:0] w_n615_0;
	wire [1:0] w_n616_0;
	wire [1:0] w_n617_0;
	wire [1:0] w_n618_0;
	wire [1:0] w_n619_0;
	wire [1:0] w_n620_0;
	wire [1:0] w_n621_0;
	wire [1:0] w_n622_0;
	wire [1:0] w_n623_0;
	wire [1:0] w_n624_0;
	wire [1:0] w_n625_0;
	wire [1:0] w_n626_0;
	wire [1:0] w_n627_0;
	wire [1:0] w_n628_0;
	wire [1:0] w_n629_0;
	wire [1:0] w_n630_0;
	wire [1:0] w_n631_0;
	wire [1:0] w_n633_0;
	wire [1:0] w_n634_0;
	wire [1:0] w_n636_0;
	wire [1:0] w_n641_0;
	wire [1:0] w_n642_0;
	wire [2:0] w_n647_0;
	wire [1:0] w_n649_0;
	wire [1:0] w_n652_0;
	wire [1:0] w_n654_0;
	wire [1:0] w_n657_0;
	wire [1:0] w_n659_0;
	wire [1:0] w_n662_0;
	wire [1:0] w_n664_0;
	wire [1:0] w_n667_0;
	wire [1:0] w_n669_0;
	wire [1:0] w_n672_0;
	wire [1:0] w_n674_0;
	wire [1:0] w_n677_0;
	wire [1:0] w_n679_0;
	wire [1:0] w_n682_0;
	wire [1:0] w_n684_0;
	wire [1:0] w_n687_0;
	wire [1:0] w_n689_0;
	wire [1:0] w_n693_0;
	wire [1:0] w_n694_0;
	wire [2:0] w_n695_0;
	wire [1:0] w_n697_0;
	wire [2:0] w_n698_0;
	wire [1:0] w_n699_0;
	wire [1:0] w_n702_0;
	wire [1:0] w_n704_0;
	wire [1:0] w_n705_0;
	wire [1:0] w_n706_0;
	wire [1:0] w_n707_0;
	wire [1:0] w_n708_0;
	wire [1:0] w_n709_0;
	wire [1:0] w_n710_0;
	wire [1:0] w_n711_0;
	wire [1:0] w_n712_0;
	wire [1:0] w_n713_0;
	wire [1:0] w_n714_0;
	wire [1:0] w_n715_0;
	wire [1:0] w_n716_0;
	wire [1:0] w_n717_0;
	wire [1:0] w_n718_0;
	wire [1:0] w_n719_0;
	wire [1:0] w_n720_0;
	wire [1:0] w_n721_0;
	wire [1:0] w_n722_0;
	wire [1:0] w_n723_0;
	wire [1:0] w_n724_0;
	wire [1:0] w_n726_0;
	wire [1:0] w_n727_0;
	wire [1:0] w_n729_0;
	wire [1:0] w_n734_0;
	wire [1:0] w_n735_0;
	wire [2:0] w_n740_0;
	wire [1:0] w_n742_0;
	wire [1:0] w_n745_0;
	wire [1:0] w_n747_0;
	wire [1:0] w_n750_0;
	wire [1:0] w_n752_0;
	wire [1:0] w_n755_0;
	wire [1:0] w_n757_0;
	wire [1:0] w_n760_0;
	wire [1:0] w_n762_0;
	wire [1:0] w_n765_0;
	wire [1:0] w_n767_0;
	wire [1:0] w_n770_0;
	wire [1:0] w_n772_0;
	wire [1:0] w_n775_0;
	wire [1:0] w_n777_0;
	wire [1:0] w_n780_0;
	wire [1:0] w_n782_0;
	wire [1:0] w_n785_0;
	wire [1:0] w_n787_0;
	wire [1:0] w_n791_0;
	wire [1:0] w_n792_0;
	wire [1:0] w_n793_0;
	wire [1:0] w_n795_0;
	wire [2:0] w_n797_0;
	wire [1:0] w_n800_0;
	wire [1:0] w_n802_0;
	wire [1:0] w_n803_0;
	wire [1:0] w_n804_0;
	wire [1:0] w_n805_0;
	wire [1:0] w_n806_0;
	wire [1:0] w_n807_0;
	wire [1:0] w_n808_0;
	wire [1:0] w_n809_0;
	wire [1:0] w_n810_0;
	wire [1:0] w_n811_0;
	wire [1:0] w_n812_0;
	wire [1:0] w_n813_0;
	wire [1:0] w_n814_0;
	wire [1:0] w_n815_0;
	wire [1:0] w_n816_0;
	wire [1:0] w_n817_0;
	wire [1:0] w_n818_0;
	wire [1:0] w_n819_0;
	wire [1:0] w_n820_0;
	wire [1:0] w_n821_0;
	wire [1:0] w_n822_0;
	wire [1:0] w_n823_0;
	wire [1:0] w_n824_0;
	wire [1:0] w_n826_0;
	wire [1:0] w_n827_0;
	wire [1:0] w_n829_0;
	wire [1:0] w_n834_0;
	wire [1:0] w_n835_0;
	wire [1:0] w_n839_0;
	wire [1:0] w_n840_0;
	wire [2:0] w_n844_0;
	wire [1:0] w_n846_0;
	wire [1:0] w_n849_0;
	wire [1:0] w_n851_0;
	wire [1:0] w_n854_0;
	wire [1:0] w_n856_0;
	wire [1:0] w_n859_0;
	wire [1:0] w_n861_0;
	wire [1:0] w_n864_0;
	wire [1:0] w_n866_0;
	wire [1:0] w_n869_0;
	wire [1:0] w_n871_0;
	wire [1:0] w_n874_0;
	wire [1:0] w_n876_0;
	wire [1:0] w_n879_0;
	wire [1:0] w_n881_0;
	wire [1:0] w_n884_0;
	wire [1:0] w_n886_0;
	wire [1:0] w_n889_0;
	wire [1:0] w_n891_0;
	wire [1:0] w_n895_0;
	wire [1:0] w_n896_0;
	wire [1:0] w_n897_0;
	wire [1:0] w_n898_0;
	wire [1:0] w_n901_0;
	wire [1:0] w_n903_0;
	wire [1:0] w_n906_0;
	wire [1:0] w_n907_0;
	wire [1:0] w_n908_0;
	wire [1:0] w_n909_0;
	wire [1:0] w_n910_0;
	wire [1:0] w_n911_0;
	wire [1:0] w_n912_0;
	wire [1:0] w_n913_0;
	wire [1:0] w_n914_0;
	wire [1:0] w_n915_0;
	wire [1:0] w_n916_0;
	wire [1:0] w_n917_0;
	wire [1:0] w_n918_0;
	wire [1:0] w_n919_0;
	wire [1:0] w_n920_0;
	wire [1:0] w_n921_0;
	wire [1:0] w_n922_0;
	wire [1:0] w_n923_0;
	wire [1:0] w_n924_0;
	wire [1:0] w_n925_0;
	wire [1:0] w_n926_0;
	wire [2:0] w_n927_0;
	wire [1:0] w_n929_0;
	wire [1:0] w_n930_0;
	wire [1:0] w_n931_0;
	wire [1:0] w_n932_0;
	wire [1:0] w_n937_0;
	wire [1:0] w_n938_0;
	wire [2:0] w_n942_0;
	wire [1:0] w_n943_0;
	wire [1:0] w_n949_0;
	wire [1:0] w_n951_0;
	wire [1:0] w_n954_0;
	wire [1:0] w_n956_0;
	wire [1:0] w_n959_0;
	wire [1:0] w_n961_0;
	wire [1:0] w_n964_0;
	wire [1:0] w_n966_0;
	wire [1:0] w_n969_0;
	wire [1:0] w_n971_0;
	wire [1:0] w_n974_0;
	wire [1:0] w_n976_0;
	wire [1:0] w_n979_0;
	wire [1:0] w_n981_0;
	wire [1:0] w_n984_0;
	wire [1:0] w_n986_0;
	wire [1:0] w_n989_0;
	wire [1:0] w_n991_0;
	wire [1:0] w_n994_0;
	wire [1:0] w_n996_0;
	wire [1:0] w_n999_0;
	wire [1:0] w_n1001_0;
	wire [1:0] w_n1005_0;
	wire [1:0] w_n1006_0;
	wire [1:0] w_n1008_0;
	wire [1:0] w_n1009_0;
	wire [1:0] w_n1010_0;
	wire [1:0] w_n1011_0;
	wire [1:0] w_n1012_0;
	wire [1:0] w_n1013_0;
	wire [1:0] w_n1014_0;
	wire [1:0] w_n1015_0;
	wire [1:0] w_n1016_0;
	wire [1:0] w_n1017_0;
	wire [1:0] w_n1018_0;
	wire [1:0] w_n1019_0;
	wire [1:0] w_n1020_0;
	wire [1:0] w_n1021_0;
	wire [1:0] w_n1022_0;
	wire [1:0] w_n1023_0;
	wire [1:0] w_n1024_0;
	wire [1:0] w_n1025_0;
	wire [1:0] w_n1026_0;
	wire [1:0] w_n1027_0;
	wire [1:0] w_n1028_0;
	wire [1:0] w_n1029_0;
	wire [1:0] w_n1030_0;
	wire [1:0] w_n1031_0;
	wire [1:0] w_n1032_0;
	wire [1:0] w_n1033_0;
	wire [1:0] w_n1034_0;
	wire [1:0] w_n1035_0;
	wire [1:0] w_n1037_0;
	wire [1:0] w_n1039_0;
	wire [1:0] w_n1043_0;
	wire [1:0] w_n1044_0;
	wire [1:0] w_n1048_0;
	wire [1:0] w_n1049_0;
	wire [1:0] w_n1052_0;
	wire [1:0] w_n1054_0;
	wire [1:0] w_n1057_0;
	wire [1:0] w_n1059_0;
	wire [1:0] w_n1062_0;
	wire [1:0] w_n1064_0;
	wire [1:0] w_n1067_0;
	wire [1:0] w_n1069_0;
	wire [1:0] w_n1072_0;
	wire [1:0] w_n1074_0;
	wire [1:0] w_n1077_0;
	wire [1:0] w_n1079_0;
	wire [1:0] w_n1082_0;
	wire [1:0] w_n1084_0;
	wire [1:0] w_n1087_0;
	wire [1:0] w_n1089_0;
	wire [1:0] w_n1092_0;
	wire [1:0] w_n1094_0;
	wire [1:0] w_n1097_0;
	wire [1:0] w_n1099_0;
	wire [1:0] w_n1102_0;
	wire [1:0] w_n1103_0;
	wire [1:0] w_n1109_0;
	wire [1:0] w_n1110_0;
	wire [1:0] w_n1114_0;
	wire [1:0] w_n1115_0;
	wire [1:0] w_n1116_0;
	wire [1:0] w_n1117_0;
	wire [1:0] w_n1118_0;
	wire [1:0] w_n1119_0;
	wire [1:0] w_n1120_0;
	wire [1:0] w_n1121_0;
	wire [1:0] w_n1122_0;
	wire [1:0] w_n1123_0;
	wire [1:0] w_n1124_0;
	wire [1:0] w_n1125_0;
	wire [1:0] w_n1126_0;
	wire [1:0] w_n1127_0;
	wire [1:0] w_n1128_0;
	wire [1:0] w_n1129_0;
	wire [1:0] w_n1130_0;
	wire [1:0] w_n1131_0;
	wire [1:0] w_n1132_0;
	wire [1:0] w_n1133_0;
	wire [1:0] w_n1134_0;
	wire [1:0] w_n1135_0;
	wire [1:0] w_n1137_0;
	wire [1:0] w_n1138_0;
	wire [1:0] w_n1139_0;
	wire [1:0] w_n1140_0;
	wire [1:0] w_n1141_0;
	wire [1:0] w_n1147_0;
	wire [1:0] w_n1151_0;
	wire [1:0] w_n1152_0;
	wire [1:0] w_n1156_0;
	wire [1:0] w_n1158_0;
	wire [1:0] w_n1161_0;
	wire [1:0] w_n1163_0;
	wire [1:0] w_n1166_0;
	wire [1:0] w_n1168_0;
	wire [1:0] w_n1171_0;
	wire [1:0] w_n1173_0;
	wire [1:0] w_n1176_0;
	wire [1:0] w_n1178_0;
	wire [1:0] w_n1181_0;
	wire [1:0] w_n1183_0;
	wire [1:0] w_n1186_0;
	wire [1:0] w_n1188_0;
	wire [1:0] w_n1191_0;
	wire [1:0] w_n1193_0;
	wire [1:0] w_n1196_0;
	wire [1:0] w_n1198_0;
	wire [1:0] w_n1201_0;
	wire [1:0] w_n1203_0;
	wire [1:0] w_n1206_0;
	wire [1:0] w_n1207_0;
	wire [1:0] w_n1208_0;
	wire [1:0] w_n1210_0;
	wire [1:0] w_n1212_0;
	wire [1:0] w_n1213_0;
	wire [1:0] w_n1214_0;
	wire [1:0] w_n1215_0;
	wire [1:0] w_n1216_0;
	wire [1:0] w_n1217_0;
	wire [1:0] w_n1218_0;
	wire [1:0] w_n1219_0;
	wire [1:0] w_n1220_0;
	wire [1:0] w_n1221_0;
	wire [1:0] w_n1222_0;
	wire [1:0] w_n1223_0;
	wire [1:0] w_n1224_0;
	wire [1:0] w_n1225_0;
	wire [1:0] w_n1226_0;
	wire [1:0] w_n1227_0;
	wire [1:0] w_n1228_0;
	wire [1:0] w_n1229_0;
	wire [1:0] w_n1230_0;
	wire [1:0] w_n1231_0;
	wire [1:0] w_n1232_0;
	wire [1:0] w_n1234_0;
	wire [1:0] w_n1236_0;
	wire [1:0] w_n1237_0;
	wire [1:0] w_n1238_0;
	wire [1:0] w_n1244_0;
	wire [1:0] w_n1247_0;
	wire [1:0] w_n1248_0;
	wire [1:0] w_n1251_0;
	wire [1:0] w_n1253_0;
	wire [1:0] w_n1256_0;
	wire [1:0] w_n1258_0;
	wire [1:0] w_n1261_0;
	wire [1:0] w_n1263_0;
	wire [1:0] w_n1266_0;
	wire [1:0] w_n1268_0;
	wire [1:0] w_n1271_0;
	wire [1:0] w_n1273_0;
	wire [1:0] w_n1276_0;
	wire [1:0] w_n1278_0;
	wire [1:0] w_n1281_0;
	wire [1:0] w_n1283_0;
	wire [1:0] w_n1286_0;
	wire [1:0] w_n1288_0;
	wire [1:0] w_n1291_0;
	wire [1:0] w_n1293_0;
	wire [1:0] w_n1296_0;
	wire [1:0] w_n1297_0;
	wire [1:0] w_n1298_0;
	wire [1:0] w_n1301_0;
	wire [1:0] w_n1303_0;
	wire [1:0] w_n1304_0;
	wire [1:0] w_n1305_0;
	wire [1:0] w_n1306_0;
	wire [1:0] w_n1307_0;
	wire [1:0] w_n1308_0;
	wire [1:0] w_n1309_0;
	wire [1:0] w_n1310_0;
	wire [1:0] w_n1311_0;
	wire [1:0] w_n1312_0;
	wire [1:0] w_n1313_0;
	wire [1:0] w_n1314_0;
	wire [1:0] w_n1315_0;
	wire [1:0] w_n1316_0;
	wire [1:0] w_n1317_0;
	wire [1:0] w_n1318_0;
	wire [1:0] w_n1319_0;
	wire [1:0] w_n1320_0;
	wire [1:0] w_n1321_0;
	wire [1:0] w_n1322_0;
	wire [1:0] w_n1324_0;
	wire [1:0] w_n1325_0;
	wire [1:0] w_n1326_0;
	wire [1:0] w_n1332_0;
	wire [1:0] w_n1337_0;
	wire [1:0] w_n1338_0;
	wire [1:0] w_n1341_0;
	wire [1:0] w_n1343_0;
	wire [1:0] w_n1346_0;
	wire [1:0] w_n1348_0;
	wire [1:0] w_n1351_0;
	wire [1:0] w_n1353_0;
	wire [1:0] w_n1356_0;
	wire [1:0] w_n1358_0;
	wire [1:0] w_n1361_0;
	wire [1:0] w_n1363_0;
	wire [1:0] w_n1366_0;
	wire [1:0] w_n1368_0;
	wire [1:0] w_n1371_0;
	wire [1:0] w_n1373_0;
	wire [1:0] w_n1376_0;
	wire [1:0] w_n1378_0;
	wire [1:0] w_n1381_0;
	wire [1:0] w_n1382_0;
	wire [1:0] w_n1383_0;
	wire [1:0] w_n1386_0;
	wire [1:0] w_n1388_0;
	wire [1:0] w_n1389_0;
	wire [1:0] w_n1390_0;
	wire [1:0] w_n1391_0;
	wire [1:0] w_n1392_0;
	wire [1:0] w_n1393_0;
	wire [1:0] w_n1394_0;
	wire [1:0] w_n1395_0;
	wire [1:0] w_n1396_0;
	wire [1:0] w_n1397_0;
	wire [1:0] w_n1398_0;
	wire [1:0] w_n1399_0;
	wire [1:0] w_n1400_0;
	wire [1:0] w_n1401_0;
	wire [1:0] w_n1402_0;
	wire [1:0] w_n1403_0;
	wire [1:0] w_n1404_0;
	wire [1:0] w_n1405_0;
	wire [1:0] w_n1407_0;
	wire [1:0] w_n1409_0;
	wire [1:0] w_n1410_0;
	wire [1:0] w_n1415_0;
	wire [1:0] w_n1420_0;
	wire [1:0] w_n1421_0;
	wire [1:0] w_n1424_0;
	wire [1:0] w_n1426_0;
	wire [1:0] w_n1429_0;
	wire [1:0] w_n1431_0;
	wire [1:0] w_n1434_0;
	wire [1:0] w_n1436_0;
	wire [1:0] w_n1439_0;
	wire [1:0] w_n1441_0;
	wire [1:0] w_n1444_0;
	wire [1:0] w_n1446_0;
	wire [1:0] w_n1449_0;
	wire [1:0] w_n1451_0;
	wire [1:0] w_n1454_0;
	wire [1:0] w_n1456_0;
	wire [1:0] w_n1459_0;
	wire [1:0] w_n1460_0;
	wire [1:0] w_n1461_0;
	wire [1:0] w_n1464_0;
	wire [1:0] w_n1466_0;
	wire [1:0] w_n1467_0;
	wire [1:0] w_n1468_0;
	wire [1:0] w_n1469_0;
	wire [1:0] w_n1470_0;
	wire [1:0] w_n1471_0;
	wire [1:0] w_n1472_0;
	wire [1:0] w_n1473_0;
	wire [1:0] w_n1474_0;
	wire [1:0] w_n1475_0;
	wire [1:0] w_n1476_0;
	wire [1:0] w_n1477_0;
	wire [1:0] w_n1478_0;
	wire [1:0] w_n1479_0;
	wire [1:0] w_n1480_0;
	wire [1:0] w_n1481_0;
	wire [1:0] w_n1483_0;
	wire [1:0] w_n1485_0;
	wire [1:0] w_n1486_0;
	wire [1:0] w_n1491_0;
	wire [1:0] w_n1496_0;
	wire [1:0] w_n1497_0;
	wire [1:0] w_n1500_0;
	wire [1:0] w_n1502_0;
	wire [1:0] w_n1505_0;
	wire [1:0] w_n1507_0;
	wire [1:0] w_n1510_0;
	wire [1:0] w_n1512_0;
	wire [1:0] w_n1515_0;
	wire [1:0] w_n1517_0;
	wire [1:0] w_n1520_0;
	wire [1:0] w_n1522_0;
	wire [1:0] w_n1525_0;
	wire [1:0] w_n1527_0;
	wire [1:0] w_n1530_0;
	wire [1:0] w_n1531_0;
	wire [1:0] w_n1532_0;
	wire [1:0] w_n1535_0;
	wire [1:0] w_n1537_0;
	wire [1:0] w_n1538_0;
	wire [1:0] w_n1539_0;
	wire [1:0] w_n1540_0;
	wire [1:0] w_n1541_0;
	wire [1:0] w_n1542_0;
	wire [1:0] w_n1543_0;
	wire [1:0] w_n1544_0;
	wire [1:0] w_n1545_0;
	wire [1:0] w_n1546_0;
	wire [1:0] w_n1547_0;
	wire [1:0] w_n1548_0;
	wire [1:0] w_n1549_0;
	wire [1:0] w_n1550_0;
	wire [1:0] w_n1552_0;
	wire [1:0] w_n1554_0;
	wire [1:0] w_n1555_0;
	wire [1:0] w_n1560_0;
	wire [1:0] w_n1565_0;
	wire [1:0] w_n1566_0;
	wire [1:0] w_n1569_0;
	wire [1:0] w_n1571_0;
	wire [1:0] w_n1574_0;
	wire [1:0] w_n1576_0;
	wire [1:0] w_n1579_0;
	wire [1:0] w_n1581_0;
	wire [1:0] w_n1584_0;
	wire [1:0] w_n1586_0;
	wire [1:0] w_n1589_0;
	wire [1:0] w_n1591_0;
	wire [1:0] w_n1594_0;
	wire [1:0] w_n1595_0;
	wire [1:0] w_n1596_0;
	wire [1:0] w_n1599_0;
	wire [1:0] w_n1601_0;
	wire [1:0] w_n1602_0;
	wire [1:0] w_n1603_0;
	wire [1:0] w_n1604_0;
	wire [1:0] w_n1605_0;
	wire [1:0] w_n1606_0;
	wire [1:0] w_n1607_0;
	wire [1:0] w_n1608_0;
	wire [1:0] w_n1609_0;
	wire [1:0] w_n1610_0;
	wire [1:0] w_n1611_0;
	wire [1:0] w_n1612_0;
	wire [1:0] w_n1614_0;
	wire [1:0] w_n1616_0;
	wire [1:0] w_n1617_0;
	wire [1:0] w_n1622_0;
	wire [1:0] w_n1627_0;
	wire [1:0] w_n1628_0;
	wire [1:0] w_n1631_0;
	wire [1:0] w_n1633_0;
	wire [1:0] w_n1636_0;
	wire [1:0] w_n1638_0;
	wire [1:0] w_n1641_0;
	wire [1:0] w_n1643_0;
	wire [1:0] w_n1646_0;
	wire [1:0] w_n1648_0;
	wire [1:0] w_n1651_0;
	wire [1:0] w_n1652_0;
	wire [1:0] w_n1653_0;
	wire [1:0] w_n1656_0;
	wire [1:0] w_n1658_0;
	wire [1:0] w_n1659_0;
	wire [1:0] w_n1660_0;
	wire [1:0] w_n1661_0;
	wire [1:0] w_n1662_0;
	wire [1:0] w_n1663_0;
	wire [1:0] w_n1664_0;
	wire [1:0] w_n1665_0;
	wire [1:0] w_n1666_0;
	wire [1:0] w_n1667_0;
	wire [1:0] w_n1669_0;
	wire [1:0] w_n1671_0;
	wire [1:0] w_n1672_0;
	wire [1:0] w_n1677_0;
	wire [1:0] w_n1682_0;
	wire [1:0] w_n1684_0;
	wire [1:0] w_n1687_0;
	wire [1:0] w_n1689_0;
	wire [1:0] w_n1692_0;
	wire [1:0] w_n1694_0;
	wire [1:0] w_n1697_0;
	wire [1:0] w_n1699_0;
	wire [1:0] w_n1702_0;
	wire [1:0] w_n1703_0;
	wire [1:0] w_n1704_0;
	wire [1:0] w_n1707_0;
	wire [1:0] w_n1709_0;
	wire [1:0] w_n1710_0;
	wire [1:0] w_n1711_0;
	wire [1:0] w_n1712_0;
	wire [1:0] w_n1713_0;
	wire [1:0] w_n1714_0;
	wire [1:0] w_n1715_0;
	wire [1:0] w_n1716_0;
	wire [1:0] w_n1717_0;
	wire [1:0] w_n1719_0;
	wire [1:0] w_n1720_0;
	wire [1:0] w_n1725_0;
	wire [1:0] w_n1728_0;
	wire [1:0] w_n1730_0;
	wire [1:0] w_n1733_0;
	wire [1:0] w_n1735_0;
	wire [1:0] w_n1738_0;
	wire [1:0] w_n1740_0;
	wire [1:0] w_n1743_0;
	wire [1:0] w_n1744_0;
	wire [1:0] w_n1745_0;
	wire [1:0] w_n1748_0;
	wire [1:0] w_n1750_0;
	wire [1:0] w_n1751_0;
	wire [1:0] w_n1752_0;
	wire [1:0] w_n1753_0;
	wire [1:0] w_n1754_0;
	wire [1:0] w_n1755_0;
	wire [1:0] w_n1756_0;
	wire [1:0] w_n1757_0;
	wire [1:0] w_n1758_0;
	wire [1:0] w_n1765_0;
	wire [1:0] w_n1768_0;
	wire [1:0] w_n1770_0;
	wire [1:0] w_n1773_0;
	wire [1:0] w_n1775_0;
	wire [1:0] w_n1778_0;
	wire [1:0] w_n1779_0;
	wire [1:0] w_n1780_0;
	wire [1:0] w_n1783_0;
	wire [1:0] w_n1785_0;
	wire [1:0] w_n1786_0;
	wire [1:0] w_n1787_0;
	wire [1:0] w_n1788_0;
	wire [1:0] w_n1789_0;
	wire [1:0] w_n1790_0;
	wire [1:0] w_n1791_0;
	wire [1:0] w_n1798_0;
	wire [1:0] w_n1801_0;
	wire [1:0] w_n1803_0;
	wire [1:0] w_n1806_0;
	wire [1:0] w_n1807_0;
	wire [1:0] w_n1808_0;
	wire [1:0] w_n1811_0;
	wire [1:0] w_n1813_0;
	wire [1:0] w_n1814_0;
	wire [1:0] w_n1815_0;
	wire [1:0] w_n1816_0;
	wire [1:0] w_n1817_0;
	wire [1:0] w_n1824_0;
	wire [1:0] w_n1827_0;
	wire [1:0] w_n1828_0;
	wire [1:0] w_n1829_0;
	wire [1:0] w_n1832_0;
	wire [1:0] w_n1834_0;
	wire [1:0] w_n1835_0;
	wire [1:0] w_n1836_0;
	wire [1:0] w_n1838_0;
	wire [1:0] w_n1841_0;
	wire [1:0] w_n1848_0;
	wire [1:0] w_n1849_0;
	wire w_dff_B_PQF7Q6RX4_1;
	wire w_dff_B_KtM7KiYd4_1;
	wire w_dff_B_ZhlSnPVz2_1;
	wire w_dff_B_n8Hb1rcW9_1;
	wire w_dff_B_tyAKh0rM9_1;
	wire w_dff_B_WsfsLaUB1_1;
	wire w_dff_B_4zMmOsTM4_1;
	wire w_dff_B_IIdfHr4V5_1;
	wire w_dff_B_dN7aLtgt7_1;
	wire w_dff_B_6OiuCooY4_1;
	wire w_dff_B_L1XRJyfl6_1;
	wire w_dff_B_ewIJIewB0_1;
	wire w_dff_B_5FevXSI36_1;
	wire w_dff_B_T589nlDk0_1;
	wire w_dff_B_ITxHWIIz4_1;
	wire w_dff_B_P9nnydua4_1;
	wire w_dff_B_UzsLI2Vz3_1;
	wire w_dff_B_PGHqKmXo0_1;
	wire w_dff_B_SWAZ2BU08_1;
	wire w_dff_B_YDVIK7HJ9_1;
	wire w_dff_B_tUTiTzBA6_1;
	wire w_dff_B_ui4FoLzg6_1;
	wire w_dff_B_ySHono3B3_1;
	wire w_dff_B_LLRp04ex6_1;
	wire w_dff_B_uMwMbtXe6_1;
	wire w_dff_B_3uSipkgl6_1;
	wire w_dff_B_v6T5OL7j9_1;
	wire w_dff_B_uknMZcEZ9_1;
	wire w_dff_B_eURwgZcN6_1;
	wire w_dff_B_E0DEu2G33_1;
	wire w_dff_B_bbbPzB4b0_1;
	wire w_dff_B_LeVcw5oU6_1;
	wire w_dff_B_vhF2fbye6_1;
	wire w_dff_B_wIIit61b4_1;
	wire w_dff_B_jyGtYMSh1_1;
	wire w_dff_B_Dfq2bJFX0_1;
	wire w_dff_B_V5S88XMb2_1;
	wire w_dff_B_1p1Cse915_1;
	wire w_dff_B_zDe0Nk612_1;
	wire w_dff_B_6DYlZ4Wv9_1;
	wire w_dff_B_iGsyV5BJ5_1;
	wire w_dff_B_2ngtrZm00_1;
	wire w_dff_B_Sw83mtes0_1;
	wire w_dff_B_Z8MvpjVb6_1;
	wire w_dff_B_r0Zve7Jg2_1;
	wire w_dff_B_hUNLCFvr1_1;
	wire w_dff_B_dhuJxHKp9_1;
	wire w_dff_B_vtWv7kPT5_1;
	wire w_dff_B_W6LWJoAP7_1;
	wire w_dff_B_5K7mlms61_1;
	wire w_dff_B_vx4ZBR9h3_1;
	wire w_dff_B_c8xqwgbt5_1;
	wire w_dff_B_feWmIk1f7_1;
	wire w_dff_B_06xoIY8R8_1;
	wire w_dff_B_o0ef297I6_1;
	wire w_dff_B_zKtuICp35_1;
	wire w_dff_B_n45O0EvX2_1;
	wire w_dff_B_4vAet7Rm0_1;
	wire w_dff_B_r0SBWScu0_1;
	wire w_dff_B_Dat5FnZs1_1;
	wire w_dff_B_vzjHGODt0_1;
	wire w_dff_B_z0CsdEBV7_1;
	wire w_dff_B_nH2cGjvr9_1;
	wire w_dff_B_G0HqAf2U0_1;
	wire w_dff_B_fB4GnBQG1_1;
	wire w_dff_B_UJBZ8oSg8_1;
	wire w_dff_B_1Mj7QbrO3_1;
	wire w_dff_B_w6z4SHnv8_1;
	wire w_dff_B_Poxu68YB1_1;
	wire w_dff_B_XUl1sJoD8_1;
	wire w_dff_B_D52GB4AA8_1;
	wire w_dff_B_vLZ0Rvma7_1;
	wire w_dff_B_DxoX74Ss2_1;
	wire w_dff_B_eGrZTmfC4_1;
	wire w_dff_B_ckDZ6xwe5_1;
	wire w_dff_B_DAPtb3rX3_1;
	wire w_dff_B_TDQN3faj4_1;
	wire w_dff_B_s6ltvAk54_1;
	wire w_dff_B_Rfj5erp36_1;
	wire w_dff_B_CrmQpBIN3_1;
	wire w_dff_B_M4qU9Zaz6_1;
	wire w_dff_B_8kJdTjWl0_1;
	wire w_dff_B_wgDUeidg0_1;
	wire w_dff_B_izKSgGRD5_1;
	wire w_dff_B_scuaBA3P9_1;
	wire w_dff_B_2MTZeLR83_1;
	wire w_dff_B_he08mcgy3_1;
	wire w_dff_B_oXdXZ9bt8_1;
	wire w_dff_B_vZmFHDus3_1;
	wire w_dff_B_9PrurzBw9_1;
	wire w_dff_B_Xsncoxn68_1;
	wire w_dff_B_uUOFw2py4_1;
	wire w_dff_B_iyDyi3uF1_1;
	wire w_dff_B_NUgGDnyd1_1;
	wire w_dff_B_ALDGzlgO8_1;
	wire w_dff_B_O8vCVjGT1_1;
	wire w_dff_B_5GsazEe12_1;
	wire w_dff_B_nh6LaOd71_1;
	wire w_dff_B_L1D3PMEI3_1;
	wire w_dff_B_t9FAN2uM4_1;
	wire w_dff_B_DFGKUIJD6_1;
	wire w_dff_B_JiFa466S7_1;
	wire w_dff_B_iI0ubWry5_1;
	wire w_dff_B_4VllvIFq9_1;
	wire w_dff_B_bIUygaES4_1;
	wire w_dff_B_e5D5TEC86_1;
	wire w_dff_B_IEq2NRb70_1;
	wire w_dff_B_N06wAm8V0_1;
	wire w_dff_B_Fg3Z1WeT2_1;
	wire w_dff_B_SLiO93it0_1;
	wire w_dff_B_uxgDp7VQ5_1;
	wire w_dff_B_iz5nuxgg5_1;
	wire w_dff_B_eCr8oSLu9_1;
	wire w_dff_B_sHMTP3JT9_1;
	wire w_dff_B_krulCJ8w6_1;
	wire w_dff_B_AavzEL6p4_1;
	wire w_dff_B_kZartvYS2_1;
	wire w_dff_B_UdHEuSoE9_1;
	wire w_dff_B_kqLUVLYO5_1;
	wire w_dff_B_VJ7UVoaq8_1;
	wire w_dff_B_nWm8VPZz1_1;
	wire w_dff_B_UTZptcMV7_1;
	wire w_dff_B_nMtdLqfT1_1;
	wire w_dff_B_XPZJBQ403_1;
	wire w_dff_B_cjVju64M6_1;
	wire w_dff_B_0Rpqzsbc9_1;
	wire w_dff_B_GjoYfDdN6_1;
	wire w_dff_B_g8md13Eg7_1;
	wire w_dff_B_Vu8awZTy1_1;
	wire w_dff_B_DllI2f9q3_1;
	wire w_dff_B_PwDdCmLD6_1;
	wire w_dff_B_0a6wVlJl0_1;
	wire w_dff_B_9jkkDO0J3_1;
	wire w_dff_B_qVpRfhja7_1;
	wire w_dff_B_unKqxwCw0_1;
	wire w_dff_B_jhY0Ph468_1;
	wire w_dff_B_a0YYHObV4_1;
	wire w_dff_B_YaDzBe1T8_1;
	wire w_dff_B_NTnK2NtP3_1;
	wire w_dff_B_WyUmnwOy7_1;
	wire w_dff_B_9MvVc6vA5_1;
	wire w_dff_B_Ix4TDhKO8_1;
	wire w_dff_B_1jI5rYFJ7_1;
	wire w_dff_B_AKd3WrEr1_1;
	wire w_dff_B_IeL3uRB35_1;
	wire w_dff_B_4wyENoWV7_1;
	wire w_dff_B_ahkEcgPM9_1;
	wire w_dff_B_t9KF2QBM8_1;
	wire w_dff_B_unEBqfAa7_1;
	wire w_dff_B_4waMXeIV3_1;
	wire w_dff_B_lGUKKiul8_1;
	wire w_dff_B_anFrpBVE5_1;
	wire w_dff_B_kVykFfvG2_1;
	wire w_dff_B_eD1xd3qJ0_1;
	wire w_dff_B_NBaIixZQ1_1;
	wire w_dff_B_ckYCSpSo5_1;
	wire w_dff_B_oGirlH2C2_1;
	wire w_dff_B_vyeF3mPc5_1;
	wire w_dff_B_mW0PzjL71_1;
	wire w_dff_B_l9DJG3cU7_1;
	wire w_dff_B_wVCT7QOs7_1;
	wire w_dff_B_FEvEN3zF4_1;
	wire w_dff_B_1YwacAhb1_1;
	wire w_dff_B_2HahP3lz4_1;
	wire w_dff_B_ALkpca9E8_1;
	wire w_dff_B_vpKDqYVp1_1;
	wire w_dff_B_1BqohqWW9_1;
	wire w_dff_B_jPJRe2Vx1_1;
	wire w_dff_B_OWW048zC0_1;
	wire w_dff_B_0nC3Wfly4_1;
	wire w_dff_B_1LKBOgen3_1;
	wire w_dff_B_aLB2d8Cb4_1;
	wire w_dff_B_nKA0yp2Q2_1;
	wire w_dff_B_cGBd3OA87_1;
	wire w_dff_B_emieqirN9_1;
	wire w_dff_B_SG3P9x418_1;
	wire w_dff_B_iHytJvjV4_1;
	wire w_dff_B_hlPpaA698_1;
	wire w_dff_B_MrbNIMoq6_1;
	wire w_dff_B_7A63QXBg4_1;
	wire w_dff_B_g4EDgwar7_1;
	wire w_dff_B_1khOGrGO3_1;
	wire w_dff_B_u7yeBYl67_1;
	wire w_dff_B_O338R50T0_1;
	wire w_dff_B_eKx4aCcY1_1;
	wire w_dff_B_pUV2rRbI9_1;
	wire w_dff_B_G6O3ndkp0_1;
	wire w_dff_B_jtLOVUAj2_1;
	wire w_dff_B_pj2vplUu7_1;
	wire w_dff_B_eX2PGYRO6_1;
	wire w_dff_B_fxTGXImx7_1;
	wire w_dff_B_wsa85A8K3_1;
	wire w_dff_B_denECjb90_1;
	wire w_dff_B_GIAdrbyx3_1;
	wire w_dff_B_gOnLd4tl9_1;
	wire w_dff_B_zQyoQ6Te9_1;
	wire w_dff_B_OFwx75Pl9_1;
	wire w_dff_B_rNN6RNev1_1;
	wire w_dff_B_I2rDsrrO3_1;
	wire w_dff_B_2AqFPdcb4_1;
	wire w_dff_B_4jyacbdo2_1;
	wire w_dff_B_j6aJq50u4_1;
	wire w_dff_B_DRoZUYa66_1;
	wire w_dff_B_x81I4trF5_1;
	wire w_dff_B_HUpk6K9F6_1;
	wire w_dff_B_aWNqCJgB3_1;
	wire w_dff_B_8IJFiap96_1;
	wire w_dff_B_t8C0qdVd1_1;
	wire w_dff_B_m85cgeEn7_1;
	wire w_dff_B_E46jhpQJ3_1;
	wire w_dff_B_6hfu1Ynt7_1;
	wire w_dff_B_OAg5oLId0_1;
	wire w_dff_B_3NDNqwgc9_1;
	wire w_dff_B_T0euW1FQ9_1;
	wire w_dff_B_TSmMUTFN5_1;
	wire w_dff_B_XOPU4qWo7_1;
	wire w_dff_B_Gxo9BsDJ1_1;
	wire w_dff_B_iiCDqQwQ1_1;
	wire w_dff_B_aoYzFfpI1_1;
	wire w_dff_B_ysdfaLGG4_1;
	wire w_dff_B_zUd21HmB0_1;
	wire w_dff_B_6PNyvwsl7_1;
	wire w_dff_B_gCuY30CU1_1;
	wire w_dff_B_UjBoxxR33_1;
	wire w_dff_B_FBqPp71W6_1;
	wire w_dff_B_MTrjtqdF6_1;
	wire w_dff_B_w9AViUWg5_1;
	wire w_dff_B_lyThDFEn0_1;
	wire w_dff_B_aiNMS3tv8_1;
	wire w_dff_B_EYClND6P2_1;
	wire w_dff_B_qpm4qKSr6_1;
	wire w_dff_B_ssHNVFP55_1;
	wire w_dff_B_fMk88tCc9_1;
	wire w_dff_B_s1iXvth84_1;
	wire w_dff_B_VmsowpXG4_1;
	wire w_dff_B_Lg2vOnfW8_1;
	wire w_dff_B_yREOMLlg4_1;
	wire w_dff_B_VBlac2Zm9_1;
	wire w_dff_B_cUcqEIWm3_1;
	wire w_dff_B_bEaYfO6w2_1;
	wire w_dff_B_XgPKrEHh5_1;
	wire w_dff_B_gsqPlIZq8_1;
	wire w_dff_B_YlZ1ifuY9_1;
	wire w_dff_B_ll7mHaFn4_1;
	wire w_dff_B_Ooq4ibow1_1;
	wire w_dff_B_r41isFue8_1;
	wire w_dff_B_9p9bTvwe7_1;
	wire w_dff_B_jwaiEsGo8_1;
	wire w_dff_B_HqmVv85Q0_1;
	wire w_dff_B_E6U2roQ78_1;
	wire w_dff_B_ZmNJV0mi8_1;
	wire w_dff_B_A8i5BUFm4_1;
	wire w_dff_B_A3nvCzqV6_1;
	wire w_dff_B_LAlxv1ln5_1;
	wire w_dff_B_jLMa77NH2_1;
	wire w_dff_B_J5pjl8qY0_0;
	wire w_dff_B_J6XJFA6V4_0;
	wire w_dff_B_Lx61Oscp4_0;
	wire w_dff_A_CEbSgHrH1_0;
	wire w_dff_A_LcoIPl2v9_0;
	wire w_dff_A_colYvOkg3_0;
	wire w_dff_A_4LDx4qi96_0;
	wire w_dff_B_XfxEq9Ce3_1;
	wire w_dff_B_yPOGelZU9_1;
	wire w_dff_B_e5lHSKNa5_2;
	wire w_dff_B_SwwazD8w1_2;
	wire w_dff_B_4uUjqRM31_2;
	wire w_dff_B_O3CQEj0Z1_2;
	wire w_dff_B_tauHEZS90_2;
	wire w_dff_B_oQ8489kV3_2;
	wire w_dff_B_WGJsjhGI8_2;
	wire w_dff_B_xwv3mdxG7_2;
	wire w_dff_B_zvLRyb8F4_2;
	wire w_dff_B_GVFpIkiz6_2;
	wire w_dff_B_SzGCV5UT3_2;
	wire w_dff_B_tjPQLyOG7_2;
	wire w_dff_B_H8b1Kziu4_2;
	wire w_dff_B_3dsv6Bni5_2;
	wire w_dff_B_tYP9EpgD4_2;
	wire w_dff_B_Gv6Quh5z0_2;
	wire w_dff_B_Qx8L1zGw4_2;
	wire w_dff_B_pW2EVA1U7_2;
	wire w_dff_B_sFI1vrC85_2;
	wire w_dff_B_9evJqlCy9_2;
	wire w_dff_B_F2CGKJ1r1_2;
	wire w_dff_B_IvaoF5hB3_2;
	wire w_dff_B_n8LDiMXb8_2;
	wire w_dff_B_ACgpmFjb1_2;
	wire w_dff_B_4HxHcM400_2;
	wire w_dff_B_lbCrCuDa2_2;
	wire w_dff_B_vsPXZqz60_2;
	wire w_dff_B_lgfc2Ygc6_2;
	wire w_dff_B_MG7DFbER2_2;
	wire w_dff_B_FXJeYFUg4_2;
	wire w_dff_B_mN9IySnE2_2;
	wire w_dff_B_ClKj2lYw6_2;
	wire w_dff_B_9NuD0v7f8_2;
	wire w_dff_B_HXCVjWyU7_2;
	wire w_dff_B_pd3gmgXl8_2;
	wire w_dff_B_nDJ2Ak723_2;
	wire w_dff_B_QWTwQzaJ9_2;
	wire w_dff_B_OkglBVIk2_2;
	wire w_dff_B_SkSwcdok2_2;
	wire w_dff_B_lEmrnIlw2_2;
	wire w_dff_B_K98NEneF9_2;
	wire w_dff_B_Kau775vn0_2;
	wire w_dff_B_ufN8n1aH5_2;
	wire w_dff_B_QjNzuNJr6_2;
	wire w_dff_B_wf5pirFW9_2;
	wire w_dff_B_no9VUopQ7_1;
	wire w_dff_B_nDhPnl7Z2_1;
	wire w_dff_B_9QfVd1cd8_1;
	wire w_dff_B_o0VQrt6u1_0;
	wire w_dff_B_bdjq8WZ84_0;
	wire w_dff_A_LHpOzrbB9_1;
	wire w_dff_A_0gs7R1tu9_1;
	wire w_dff_A_8XbjN7ht0_1;
	wire w_dff_B_KLybpQBG8_1;
	wire w_dff_B_RQidEsZv6_1;
	wire w_dff_B_J9BCiSGh4_1;
	wire w_dff_B_kL81Hs7F0_0;
	wire w_dff_B_q4rbk8rf0_0;
	wire w_dff_A_wwmBWZok5_1;
	wire w_dff_A_IKXWMXrh0_1;
	wire w_dff_A_xCr3eRnX3_1;
	wire w_dff_B_smNPmZ0o0_1;
	wire w_dff_B_mGstzwpw6_1;
	wire w_dff_B_OoUBXaLt3_1;
	wire w_dff_B_PtIjhdST2_0;
	wire w_dff_B_L95tFTN21_0;
	wire w_dff_A_KfbsAAkH5_1;
	wire w_dff_A_lGdhC9L15_1;
	wire w_dff_A_RZILa9VN8_1;
	wire w_dff_B_R2kBV6Qy2_1;
	wire w_dff_B_RHSz7nkh9_1;
	wire w_dff_B_qLp2GrJg0_1;
	wire w_dff_B_hI3AXSox5_0;
	wire w_dff_B_d0PaMaEw8_0;
	wire w_dff_A_HYyviQ8l6_1;
	wire w_dff_A_OJKRTlii0_1;
	wire w_dff_A_4zVLMqc52_1;
	wire w_dff_B_xmas2Tcw1_1;
	wire w_dff_B_fMmwneKP0_1;
	wire w_dff_B_FDF2le2Q4_1;
	wire w_dff_B_wNIJnD189_0;
	wire w_dff_A_dUeVK5hN0_1;
	wire w_dff_A_K74FCtSl7_1;
	wire w_dff_B_dlR0tHnC9_1;
	wire w_dff_B_4vwGwDhX0_1;
	wire w_dff_A_j7CybSZ25_1;
	wire w_dff_B_JRhUGIwa0_1;
	wire w_dff_B_FrfsuDlV9_1;
	wire w_dff_A_vLMIrqfW2_1;
	wire w_dff_B_cACy4Rp22_1;
	wire w_dff_B_mmxUZK7d1_1;
	wire w_dff_A_GB6k6xy42_1;
	wire w_dff_B_SMqQ1jin0_1;
	wire w_dff_B_3ViiBqlr3_1;
	wire w_dff_A_uzm3y4NF2_1;
	wire w_dff_B_51WYu2pA6_1;
	wire w_dff_B_gezxGVAF9_1;
	wire w_dff_A_NXQdRrj24_0;
	wire w_dff_B_aUjjF2ug5_1;
	wire w_dff_A_3bZjpayx8_0;
	wire w_dff_A_7yfYQd7z3_1;
	wire w_dff_B_7mxns7If6_2;
	wire w_dff_A_QGWkux4p1_1;
	wire w_dff_B_GAtqHJmd0_2;
	wire w_dff_B_BJ8Cjrj89_1;
	wire w_dff_A_M2y5S9Ic2_0;
	wire w_dff_A_A2z74COT3_0;
	wire w_dff_A_JIcAdYUM5_0;
	wire w_dff_A_JBsj4P8Y0_0;
	wire w_dff_A_mRyn88YL5_0;
	wire w_dff_A_LMH93aDI4_0;
	wire w_dff_A_4dUtf8aZ0_0;
	wire w_dff_A_HRy1BVDF9_0;
	wire w_dff_A_RA2lbvZJ3_0;
	wire w_dff_A_OuYs5i7w5_0;
	wire w_dff_A_nfBGby8k2_0;
	wire w_dff_A_CAO2L0DN0_0;
	wire w_dff_A_vVFD8ip00_0;
	wire w_dff_A_IWHs54U20_0;
	wire w_dff_A_stS7mkZF6_0;
	wire w_dff_A_LcNbG2I07_0;
	wire w_dff_A_4X7SLdyk8_0;
	wire w_dff_A_lA4eFy8G1_0;
	wire w_dff_A_Ni5oRJLR8_0;
	wire w_dff_A_VzuHRQVR7_0;
	wire w_dff_A_17Qpn3K31_0;
	wire w_dff_A_oEJZhH0h4_0;
	wire w_dff_A_NAMCyyWl9_0;
	wire w_dff_A_20oDcLU86_0;
	wire w_dff_A_b3mkxzp26_0;
	wire w_dff_A_bp1CZuUc8_0;
	wire w_dff_A_yLEvCfby4_0;
	wire w_dff_A_FKnfKZf90_0;
	wire w_dff_A_CZmSBxDb7_0;
	wire w_dff_A_TPvmPQxl1_0;
	wire w_dff_A_jiBmBqhU0_0;
	wire w_dff_A_IEtz1gEB5_0;
	wire w_dff_A_0sPTpbU60_1;
	wire w_dff_A_ckJvRe8q1_0;
	wire w_dff_A_Ni3RkCnE9_0;
	wire w_dff_A_4aLrPhyA2_0;
	wire w_dff_A_TGoF8XTR4_0;
	wire w_dff_A_SptcI34m8_0;
	wire w_dff_A_JyliSIvt9_0;
	wire w_dff_A_V9LDcEmT3_0;
	wire w_dff_A_28GU9gwZ6_0;
	wire w_dff_A_526ddzCd9_0;
	wire w_dff_A_w5edsb1a8_0;
	wire w_dff_A_YvzVBEEJ0_0;
	wire w_dff_A_C3bllVpi9_0;
	wire w_dff_A_MCFx6G085_0;
	wire w_dff_A_2c3v1nxu0_0;
	wire w_dff_A_c6Mxnvs21_0;
	wire w_dff_A_crciOiXx2_0;
	wire w_dff_A_SVvyptEf1_0;
	wire w_dff_A_nQ18yLAS9_0;
	wire w_dff_A_fvr7R8Ou9_0;
	wire w_dff_A_yM8oqcQK0_0;
	wire w_dff_A_ePW2K3FK6_0;
	wire w_dff_A_48xqbwZu3_0;
	wire w_dff_A_OxZ5SWrm2_0;
	wire w_dff_A_5tOxizFb2_0;
	wire w_dff_A_GZe99MoZ8_0;
	wire w_dff_A_hwkeze6Q3_0;
	wire w_dff_A_byWbHRO86_0;
	wire w_dff_A_5eG2FIa74_0;
	wire w_dff_A_HtM3viRm2_0;
	wire w_dff_A_1NxHfHhh4_0;
	wire w_dff_B_j1Qyn4VR3_1;
	wire w_dff_B_m8bmo6tf8_1;
	wire w_dff_B_cW4qRpP29_1;
	wire w_dff_B_hsCRbPDH6_1;
	wire w_dff_B_n8oKYvc81_1;
	wire w_dff_B_W0eCNOpV2_1;
	wire w_dff_B_WwR90PSf0_1;
	wire w_dff_B_4s2z4bQe9_1;
	wire w_dff_B_Pc03QurW3_1;
	wire w_dff_B_Q2hjMnad1_1;
	wire w_dff_B_KW99sxBe3_1;
	wire w_dff_B_KSsNT7ek7_1;
	wire w_dff_B_i4zLOusD5_1;
	wire w_dff_B_B7GCk5jB5_1;
	wire w_dff_B_5XK3Jzp21_1;
	wire w_dff_B_hk2cQKiP0_1;
	wire w_dff_B_yoX6QolF8_1;
	wire w_dff_B_gCb0fjIb4_1;
	wire w_dff_B_9Qkc2j0j4_1;
	wire w_dff_B_VAwY4NUY2_1;
	wire w_dff_B_mxfUhMI60_1;
	wire w_dff_B_jESRqfOh5_1;
	wire w_dff_B_bJiwrdoI9_1;
	wire w_dff_B_5ogWIryP1_1;
	wire w_dff_B_VyhpvSaU5_1;
	wire w_dff_B_WoRw4qqH9_1;
	wire w_dff_B_xftUq9QE4_1;
	wire w_dff_A_QRIEawwW9_0;
	wire w_dff_A_aRpb6lCj9_0;
	wire w_dff_A_h3kN2Rjy9_0;
	wire w_dff_A_aNVKrYK82_0;
	wire w_dff_A_SnlyMRNp5_0;
	wire w_dff_A_tst7LY0G2_0;
	wire w_dff_A_YoptpFe12_0;
	wire w_dff_A_r7YpmhuF6_0;
	wire w_dff_A_6CCUXlFh6_0;
	wire w_dff_A_TdwC0G0v3_0;
	wire w_dff_A_sBPdLfx06_0;
	wire w_dff_A_trkkQhNo2_0;
	wire w_dff_A_oqo6Js0f1_0;
	wire w_dff_A_4FLuXmca2_0;
	wire w_dff_A_f6sjOfPn2_0;
	wire w_dff_A_DBZipzq48_0;
	wire w_dff_A_Nd5NTdfd6_0;
	wire w_dff_A_hE6U68IY4_0;
	wire w_dff_A_0DmC97dg8_0;
	wire w_dff_A_2xMyIXmD9_0;
	wire w_dff_A_L0ZJ7ZMt8_0;
	wire w_dff_A_6eB7NOTM5_0;
	wire w_dff_A_dYDNLr6f6_0;
	wire w_dff_A_37pS510B7_0;
	wire w_dff_A_7h8LuNmB3_0;
	wire w_dff_A_5ZDX1ojs8_0;
	wire w_dff_A_t6ymttmX7_0;
	wire w_dff_A_mxYlMU4T7_0;
	wire w_dff_A_5SfzQAxg5_0;
	wire w_dff_B_Gtx6iQUT5_1;
	wire w_dff_B_wgVc6paT1_1;
	wire w_dff_B_dyBECQd94_1;
	wire w_dff_B_y7YCC6nS9_1;
	wire w_dff_B_2rtJJHXR5_1;
	wire w_dff_B_dTfkslxc8_1;
	wire w_dff_B_nRodWvVy6_1;
	wire w_dff_B_pfTDFgzc5_1;
	wire w_dff_B_xJd63XPY8_1;
	wire w_dff_B_VWS1LYYq2_1;
	wire w_dff_B_Rhx6ugLh3_1;
	wire w_dff_B_5kB4Rtwn1_1;
	wire w_dff_B_vqu4icbf5_1;
	wire w_dff_B_1ftpvpHc5_1;
	wire w_dff_B_Dpo3CHuE5_1;
	wire w_dff_B_ntEUX0s01_1;
	wire w_dff_B_LEganfDA6_1;
	wire w_dff_B_i5rTkOQc3_1;
	wire w_dff_B_1Bmrf8M43_1;
	wire w_dff_B_Hj3FjrsB0_1;
	wire w_dff_B_4Q5j9i1D5_1;
	wire w_dff_B_COvC5jYA1_1;
	wire w_dff_B_SN9eq7xb6_1;
	wire w_dff_B_yCYtyNGu2_1;
	wire w_dff_B_Y7kUWzNe8_1;
	wire w_dff_A_chNdRabH2_0;
	wire w_dff_A_t6UoPEjo7_0;
	wire w_dff_A_Xy5grSm04_0;
	wire w_dff_A_pBCy3b054_0;
	wire w_dff_A_2hueUNo63_0;
	wire w_dff_A_8YjE5BJm3_0;
	wire w_dff_A_gv21w5aP5_0;
	wire w_dff_A_kVJo1b3u0_0;
	wire w_dff_A_Olfva5oa8_0;
	wire w_dff_A_YRCqZGhF9_0;
	wire w_dff_A_USs8jSmu6_0;
	wire w_dff_A_IuOQWvfL6_0;
	wire w_dff_A_hsl7nrrv4_0;
	wire w_dff_A_BjYwVVvi0_0;
	wire w_dff_A_Swnzi0bJ0_0;
	wire w_dff_A_KXe3CEHZ1_0;
	wire w_dff_A_2BXQFruY2_0;
	wire w_dff_A_DwUuqx5f6_0;
	wire w_dff_A_7eF34zr54_0;
	wire w_dff_A_GdEAqnOh5_0;
	wire w_dff_A_LrlmMQgS7_0;
	wire w_dff_A_uvg8JFR27_0;
	wire w_dff_A_XrxlCHqV1_0;
	wire w_dff_A_lpGWMR4J8_0;
	wire w_dff_A_gx8XY1136_0;
	wire w_dff_A_DDChMjQ80_0;
	wire w_dff_A_kbhaqNm07_0;
	wire w_dff_B_0Fl91qHa7_1;
	wire w_dff_B_oQaJROwe8_1;
	wire w_dff_B_SIDBVwWf5_1;
	wire w_dff_B_B9lmbFg19_1;
	wire w_dff_B_rMR5z9EP1_1;
	wire w_dff_B_36UGUMST0_1;
	wire w_dff_B_he42QObT1_1;
	wire w_dff_B_OgHDIqo14_1;
	wire w_dff_B_zxabgURl9_1;
	wire w_dff_B_QSwSKHzD6_1;
	wire w_dff_B_TWyROOLA9_1;
	wire w_dff_B_iNmXmHwP8_1;
	wire w_dff_B_WvdwlZDU6_1;
	wire w_dff_B_r9EjzCyz0_1;
	wire w_dff_B_5UpzrQaH9_1;
	wire w_dff_B_F5M7TLqH5_1;
	wire w_dff_B_AzM9MPQw4_1;
	wire w_dff_B_XQJnSe9C6_1;
	wire w_dff_B_2D7TI53e2_1;
	wire w_dff_B_DiYja20U1_1;
	wire w_dff_B_nsyH24CG9_1;
	wire w_dff_B_u03696M12_1;
	wire w_dff_B_Bid8kzJ10_1;
	wire w_dff_A_al1351FM3_0;
	wire w_dff_A_JaPsF6wM6_0;
	wire w_dff_A_7lPUfc5j1_0;
	wire w_dff_A_GfbLkeaF8_0;
	wire w_dff_A_IARJly4G8_0;
	wire w_dff_A_S3vFVcLD6_0;
	wire w_dff_A_H2H2BRE85_0;
	wire w_dff_A_ADcGAanS1_0;
	wire w_dff_A_jQKr9a962_0;
	wire w_dff_A_jfStBTsP3_0;
	wire w_dff_A_P0llhrgA8_0;
	wire w_dff_A_QcoF8xF19_0;
	wire w_dff_A_xM9sCwMX4_0;
	wire w_dff_A_ifSAndGT2_0;
	wire w_dff_A_Z40eYaM17_0;
	wire w_dff_A_Oafz2oKT9_0;
	wire w_dff_A_CjbwsbKT4_0;
	wire w_dff_A_ysOHlpa41_0;
	wire w_dff_A_aqIJ95c39_0;
	wire w_dff_A_33K2h22O9_0;
	wire w_dff_A_mN8EVr0i4_0;
	wire w_dff_A_AR0uX3qQ2_0;
	wire w_dff_A_CxgODUZJ1_0;
	wire w_dff_A_gpPMgTpp3_0;
	wire w_dff_A_vEIwA6aA0_0;
	wire w_dff_B_ud8QjlEU3_1;
	wire w_dff_B_zmI335mi6_1;
	wire w_dff_B_bWBOJdYY1_1;
	wire w_dff_B_xr8SIehP1_1;
	wire w_dff_B_XLedBFm88_1;
	wire w_dff_B_doerRJqm9_1;
	wire w_dff_B_rLxTfpQs0_1;
	wire w_dff_B_pSRY3bP35_1;
	wire w_dff_B_eAhSCHeG3_1;
	wire w_dff_B_PQF5T7Wg5_1;
	wire w_dff_B_MtaOSoxO6_1;
	wire w_dff_B_WsdHjk4y5_1;
	wire w_dff_B_xOW5Oup12_1;
	wire w_dff_B_3l0KOHsB0_1;
	wire w_dff_B_56TIV0FV7_1;
	wire w_dff_B_R7nHuzbv0_1;
	wire w_dff_B_uNLZFaGt3_1;
	wire w_dff_B_aRHot1te5_1;
	wire w_dff_B_WnJR3tlD2_1;
	wire w_dff_B_H9cIAPfO1_1;
	wire w_dff_B_vTo9DWpq2_1;
	wire w_dff_A_swXZQXih8_0;
	wire w_dff_A_05DEkaV64_0;
	wire w_dff_A_oS9J8bpO0_0;
	wire w_dff_A_wrzDHA7Z5_0;
	wire w_dff_A_j3vvAh7y7_0;
	wire w_dff_A_ojWLVKT07_0;
	wire w_dff_A_hw03vZm11_0;
	wire w_dff_A_yvzcvKpM1_0;
	wire w_dff_A_teefEHzH5_0;
	wire w_dff_A_2KoD1YQX8_0;
	wire w_dff_A_KRqEwjQ81_0;
	wire w_dff_A_k0spBbv27_0;
	wire w_dff_A_1y2ZKeWk4_0;
	wire w_dff_A_ACy3FlvS3_0;
	wire w_dff_A_LZ60edm54_0;
	wire w_dff_A_W3yj2vlt8_0;
	wire w_dff_A_J1NUl2kS2_0;
	wire w_dff_A_dqFCisM34_0;
	wire w_dff_A_6u1ojk1k5_0;
	wire w_dff_A_U3qzrxTV4_0;
	wire w_dff_A_1xG9BDfg7_0;
	wire w_dff_A_q9OgaS2z8_0;
	wire w_dff_A_hM36iCne8_0;
	wire w_dff_B_uTZb6Z3s7_1;
	wire w_dff_B_hm1fPZAq7_1;
	wire w_dff_B_EHcLlbm60_1;
	wire w_dff_B_ODuCTbQ85_1;
	wire w_dff_B_izjg92Ap4_1;
	wire w_dff_B_L8w81y2j8_1;
	wire w_dff_B_zWcbds0U5_1;
	wire w_dff_B_5XlOMBgl2_1;
	wire w_dff_B_b5uxt2mY6_1;
	wire w_dff_B_VhGYBEJb5_1;
	wire w_dff_B_afhVULOk7_1;
	wire w_dff_B_NWYGAxDR3_1;
	wire w_dff_B_5bHmcDTs4_1;
	wire w_dff_B_RgpgXzOc0_1;
	wire w_dff_B_0SHDZ3w04_1;
	wire w_dff_B_16LtevOL6_1;
	wire w_dff_B_shtQC2Mn4_1;
	wire w_dff_B_YUNO8IgW0_1;
	wire w_dff_B_E5IsYMmE0_1;
	wire w_dff_A_TVX9hYFf4_0;
	wire w_dff_A_tJT3KFuh6_0;
	wire w_dff_A_W4EAAdrH1_0;
	wire w_dff_A_FqopWnku8_0;
	wire w_dff_A_bvsaJjqH8_0;
	wire w_dff_A_pOTCGV5m3_0;
	wire w_dff_A_aKvz969A3_0;
	wire w_dff_A_dYxmvQzE1_0;
	wire w_dff_A_py3Lhpao5_0;
	wire w_dff_A_RPAy8iYG1_0;
	wire w_dff_A_MlQGDNEl0_0;
	wire w_dff_A_8VIXhoDg6_0;
	wire w_dff_A_tTJxgcJW1_0;
	wire w_dff_A_HQMVwezQ1_0;
	wire w_dff_A_HSaA9MkR6_0;
	wire w_dff_A_iMhyR4d71_0;
	wire w_dff_A_QBgFagCF7_0;
	wire w_dff_A_6cadBoT13_0;
	wire w_dff_A_vYF5bntp6_0;
	wire w_dff_A_sOfPWkRK0_0;
	wire w_dff_A_Vez93m5r5_0;
	wire w_dff_B_m1nTTzLv5_1;
	wire w_dff_B_LcYa4VeC7_1;
	wire w_dff_B_08TmuP7q1_1;
	wire w_dff_B_2mJ8EhpL4_1;
	wire w_dff_B_3FLLYQeS5_1;
	wire w_dff_B_cA2vQFFR6_1;
	wire w_dff_B_YgSRbCQH3_1;
	wire w_dff_B_GlLYAf4y4_1;
	wire w_dff_B_nE6JvbLd3_1;
	wire w_dff_B_SP1WKq941_1;
	wire w_dff_B_etxLYvyE0_1;
	wire w_dff_B_y1UcUOWs1_1;
	wire w_dff_B_F0WfyupO0_1;
	wire w_dff_B_DNlOVOYA8_1;
	wire w_dff_B_U4FZBcFX0_1;
	wire w_dff_B_Gu4FAlXo2_1;
	wire w_dff_B_uzgOcgVR6_1;
	wire w_dff_A_2T7pXLSx7_0;
	wire w_dff_A_Pix4WXTg3_0;
	wire w_dff_A_LPLBZKPO0_0;
	wire w_dff_A_8egFxdP22_0;
	wire w_dff_A_khLpirm57_0;
	wire w_dff_A_0GYK5jNy7_0;
	wire w_dff_A_x0qTc6vE7_0;
	wire w_dff_A_DpsND7iO2_0;
	wire w_dff_A_9S7CCJsF3_0;
	wire w_dff_A_Pz0QLjXJ3_0;
	wire w_dff_A_nYuhlZqn1_0;
	wire w_dff_A_2EpMaSnq8_0;
	wire w_dff_A_673CrR0C2_0;
	wire w_dff_A_WSzD5Wpn9_0;
	wire w_dff_A_lNBjx5ke5_0;
	wire w_dff_A_CvXFFNkg9_0;
	wire w_dff_A_FdzGiTDI8_0;
	wire w_dff_A_IoO125sj7_0;
	wire w_dff_A_m3nABioh9_0;
	wire w_dff_B_bXzx77a41_1;
	wire w_dff_B_FMnajm8G4_1;
	wire w_dff_B_ccdDxJkD0_1;
	wire w_dff_B_XhRnvKZZ1_1;
	wire w_dff_B_9Rx8xwna0_1;
	wire w_dff_B_WIa8yhxu1_1;
	wire w_dff_B_hiyWUse81_1;
	wire w_dff_B_GrOBJnqH2_1;
	wire w_dff_B_u8g1M5HO3_1;
	wire w_dff_B_3KcMjNye2_1;
	wire w_dff_B_DM0c2Tpp5_1;
	wire w_dff_B_TP5Shjm96_1;
	wire w_dff_B_OB4DEuRr8_1;
	wire w_dff_B_G1KyZF0M8_1;
	wire w_dff_B_T7dveuQ82_1;
	wire w_dff_A_C95lVcqm2_0;
	wire w_dff_A_Vi6tqybi3_0;
	wire w_dff_A_J7xmdvLm9_0;
	wire w_dff_A_wcUSb0ND0_0;
	wire w_dff_A_DUiltiON6_0;
	wire w_dff_A_ZR8UbXeW8_0;
	wire w_dff_A_vdIwsETk7_0;
	wire w_dff_A_y6UBtydD0_0;
	wire w_dff_A_CgEma8ZJ4_0;
	wire w_dff_A_gl5Qt2Ot8_0;
	wire w_dff_A_7mv1w4M16_0;
	wire w_dff_A_yxy9RVM56_0;
	wire w_dff_A_cH4aSYDU7_0;
	wire w_dff_A_hKqXMD9c0_0;
	wire w_dff_A_kNtRzy8m2_0;
	wire w_dff_A_7G13RT427_0;
	wire w_dff_A_AQFbMP098_0;
	wire w_dff_B_oWFygZgG2_1;
	wire w_dff_B_akbrEpRE8_1;
	wire w_dff_B_YiAkGpZx9_1;
	wire w_dff_B_quKfcrm47_1;
	wire w_dff_B_TuJdajx77_1;
	wire w_dff_B_1WAubDVB4_1;
	wire w_dff_B_nwwEBhyz4_1;
	wire w_dff_B_zMEQz6ua2_1;
	wire w_dff_B_VDUySVi49_1;
	wire w_dff_B_UFQIP7y21_1;
	wire w_dff_B_judfDY4v3_1;
	wire w_dff_B_iS1z2tby3_1;
	wire w_dff_B_RUOdUyiF6_1;
	wire w_dff_A_oDeo4JQK6_0;
	wire w_dff_A_l3pzBfjS2_0;
	wire w_dff_A_cjgpqF0p3_0;
	wire w_dff_A_uOyZRKLN6_0;
	wire w_dff_A_xjTL6E8p5_0;
	wire w_dff_A_11UYdMps8_0;
	wire w_dff_A_Xh5PV9FL2_0;
	wire w_dff_A_3chRoaCD9_0;
	wire w_dff_A_gcf6QSsY4_0;
	wire w_dff_A_z4wlQNNV1_0;
	wire w_dff_A_5rOWLprw6_0;
	wire w_dff_A_SjSjZ8Cg4_0;
	wire w_dff_A_Ok4TBqic0_0;
	wire w_dff_A_OVDrevzS6_0;
	wire w_dff_A_mnSlSRY63_0;
	wire w_dff_B_dRsffrHs6_1;
	wire w_dff_B_hATEjAtW6_1;
	wire w_dff_B_jPMCi8ZN0_1;
	wire w_dff_B_EFirFdGd0_1;
	wire w_dff_B_FTL8EDBx4_1;
	wire w_dff_B_wnoAgGL21_1;
	wire w_dff_B_gIrIlQin4_1;
	wire w_dff_B_8VhK9wsb3_1;
	wire w_dff_B_3S00F6qj7_1;
	wire w_dff_B_E2bs8Qwu3_1;
	wire w_dff_B_FeQGZ0tg2_1;
	wire w_dff_A_LL0DfKUa1_0;
	wire w_dff_A_lOlDLeYk8_0;
	wire w_dff_A_qkiU0kGP6_0;
	wire w_dff_A_q0emCLJe2_0;
	wire w_dff_A_PlsV4TOb8_0;
	wire w_dff_A_J7J5Wt4u7_0;
	wire w_dff_A_8vUDIetG5_0;
	wire w_dff_A_cl4f1fZh7_0;
	wire w_dff_A_CP5ZuuGR5_0;
	wire w_dff_A_3dqgACn87_0;
	wire w_dff_A_G28ZyrZ98_0;
	wire w_dff_A_LcbbC6Gi6_0;
	wire w_dff_A_7HPLrMCC8_0;
	wire w_dff_B_zqWSIJpp8_1;
	wire w_dff_B_5XJ0MbIU3_1;
	wire w_dff_B_0h3XU6Cx5_1;
	wire w_dff_B_jglCie9R7_1;
	wire w_dff_B_IqNhxrqy8_1;
	wire w_dff_B_saczajSj6_1;
	wire w_dff_B_i0kVo9my7_1;
	wire w_dff_B_AjzgUDJh3_1;
	wire w_dff_B_26rhsQip6_1;
	wire w_dff_A_TenYRsws0_0;
	wire w_dff_A_1Q843crG3_0;
	wire w_dff_A_b4OC8tPc0_0;
	wire w_dff_A_6QYMP0Pm2_0;
	wire w_dff_A_AOLB0mop3_0;
	wire w_dff_A_LsVDsME93_0;
	wire w_dff_A_6rwN02mZ0_0;
	wire w_dff_A_JhvXPSSm7_0;
	wire w_dff_A_aDKKiVNS0_0;
	wire w_dff_A_wScBvGaT4_0;
	wire w_dff_A_WdwwOVyQ8_0;
	wire w_dff_B_0fv5yjhA6_1;
	wire w_dff_B_I2hCNous3_1;
	wire w_dff_B_P9ACDME41_1;
	wire w_dff_B_Jq6Qy6BN0_1;
	wire w_dff_B_nCEzdcfE5_1;
	wire w_dff_B_JC0Y6Ui80_1;
	wire w_dff_B_Wsh9ZRGM0_1;
	wire w_dff_A_lXilLWhR4_0;
	wire w_dff_B_o082cFWp4_2;
	wire w_dff_A_1MrAJqss9_0;
	wire w_dff_A_XJmi4JZf0_0;
	wire w_dff_A_TWDGeNcx3_0;
	wire w_dff_A_83xhQuQT4_0;
	wire w_dff_A_PbFVMIW76_0;
	wire w_dff_A_qbIqQljw1_0;
	wire w_dff_A_Sb20tTNi4_0;
	wire w_dff_B_97tUUQ5T3_1;
	wire w_dff_B_Ej0vGfTk0_1;
	wire w_dff_B_1my9ggDg8_1;
	wire w_dff_B_RMpO3DLV2_1;
	wire w_dff_A_QEwu1QkQ3_0;
	wire w_dff_B_jI2yWL6q9_2;
	wire w_dff_B_IDjAmrQo7_0;
	wire w_dff_A_xryOKzr28_0;
	wire w_dff_A_GTirAPbm7_0;
	wire w_dff_A_wr6o7ltw7_0;
	wire w_dff_B_Zg4WHi4m7_0;
	wire w_dff_A_PMzkp3Yy3_0;
	wire w_dff_A_iW07Qgb02_0;
	wire w_dff_B_siiwXJJ18_2;
	wire w_dff_A_JALddgvv6_1;
	wire w_dff_B_ceVyse8u0_2;
	wire w_dff_B_OsKKAQx83_2;
	wire w_dff_B_Iznw8x703_2;
	wire w_dff_B_o0OJDUGi4_2;
	wire w_dff_B_zOABYoD24_2;
	wire w_dff_B_eCn0dC6B2_2;
	wire w_dff_B_QnGobxNJ1_2;
	wire w_dff_B_pyBbdSKc3_2;
	wire w_dff_B_4dwZJS6X4_2;
	wire w_dff_B_i9d2Xck33_2;
	wire w_dff_B_v8FSVbER3_2;
	wire w_dff_B_GnhrRIJZ1_2;
	wire w_dff_B_InpRgIT89_2;
	wire w_dff_B_rlSwGTiB2_2;
	wire w_dff_B_025hKoW00_2;
	wire w_dff_B_uAvGqAgU4_2;
	wire w_dff_B_ei0xRJXx8_2;
	wire w_dff_B_jrIUrfQ32_2;
	wire w_dff_B_ptRYBJqs3_2;
	wire w_dff_B_aIr8GCuP4_2;
	wire w_dff_B_wKgyXslP4_2;
	wire w_dff_B_Xd26Q48Y8_2;
	wire w_dff_B_6hAmRQfI3_2;
	wire w_dff_B_LbHddnH23_2;
	wire w_dff_B_ifMVYr991_2;
	wire w_dff_B_rv5wyhox2_2;
	wire w_dff_B_EQrBiNvS3_2;
	wire w_dff_B_se56qiBO2_2;
	wire w_dff_B_HLMsBhxG1_2;
	wire w_dff_B_z7aPTPIf2_2;
	wire w_dff_B_wQLZOnu17_2;
	wire w_dff_B_kWfNUNAt5_2;
	wire w_dff_A_i1clNZ0m9_1;
	wire w_dff_A_um8ltIX04_2;
	wire w_dff_B_kLnAW15u8_3;
	wire w_dff_B_fPYh2NFM3_2;
	wire w_dff_B_PAx0Mzac1_2;
	wire w_dff_B_nnX5S40d4_2;
	wire w_dff_B_nKHf3q6X9_2;
	wire w_dff_B_1lRvW5IM7_2;
	wire w_dff_B_Br75LXZQ4_2;
	wire w_dff_B_foy3zvNv4_2;
	wire w_dff_B_uvZJOAsb5_2;
	wire w_dff_B_0Oqemyyk9_2;
	wire w_dff_B_gJUKotO98_2;
	wire w_dff_B_pSOEjo3U0_2;
	wire w_dff_B_gp322aiT5_2;
	wire w_dff_B_Ngf8tBR99_2;
	wire w_dff_B_HpgOyv5H4_2;
	wire w_dff_B_1vt9VwUq3_2;
	wire w_dff_B_WuLWAwiU6_2;
	wire w_dff_B_bkDjcfUG8_2;
	wire w_dff_B_DLD2mCQd1_2;
	wire w_dff_B_lZUU5Ikp7_2;
	wire w_dff_B_NNYrsWlx4_2;
	wire w_dff_B_0HmUS0n64_2;
	wire w_dff_B_4umjEWuQ9_2;
	wire w_dff_B_cgk9FrNK0_2;
	wire w_dff_B_oaxqtx8w6_2;
	wire w_dff_B_av554reE0_2;
	wire w_dff_B_bH9gXNBM5_2;
	wire w_dff_B_0x9xVjx69_2;
	wire w_dff_B_wPE0grvz8_2;
	wire w_dff_B_ik6tOIxU0_2;
	wire w_dff_B_HA4refMf4_1;
	wire w_dff_B_yZmTFvSo7_1;
	wire w_dff_B_GMRb3hFM3_1;
	wire w_dff_B_DBFYvmrq9_1;
	wire w_dff_B_LyUd0YqQ7_1;
	wire w_dff_B_mlbQyOMs1_1;
	wire w_dff_B_5eZA3ChM6_1;
	wire w_dff_B_gWK2mxjU5_1;
	wire w_dff_B_Cd67rXIQ7_1;
	wire w_dff_B_ZJLVSupR9_1;
	wire w_dff_B_g2KoK8Yr2_1;
	wire w_dff_B_6u0lKJHd8_1;
	wire w_dff_B_ZT7sgB5c1_1;
	wire w_dff_B_6EABTwI58_1;
	wire w_dff_B_xLco0Nea9_1;
	wire w_dff_B_oldjHmBk3_1;
	wire w_dff_B_r7WWhIwN8_1;
	wire w_dff_B_Enw8Q78Y7_1;
	wire w_dff_B_zQASk2fe0_1;
	wire w_dff_B_lt3OFEtz3_1;
	wire w_dff_B_P3wPA5Ou0_1;
	wire w_dff_B_uKVyaURs6_1;
	wire w_dff_B_VDgJkdLD4_1;
	wire w_dff_B_eDn57moe7_1;
	wire w_dff_B_UcabbIXb5_1;
	wire w_dff_B_GNqgMNCd9_1;
	wire w_dff_A_13aE2Vnd9_0;
	wire w_dff_A_YAHfWe8j5_0;
	wire w_dff_A_FaZnX2s07_0;
	wire w_dff_A_H2SMGDSo1_0;
	wire w_dff_A_yNDvrETi5_0;
	wire w_dff_A_pfrkrKcp0_0;
	wire w_dff_A_dziXrN4W6_0;
	wire w_dff_A_ES0o6cA46_0;
	wire w_dff_A_UXAfSEdm3_0;
	wire w_dff_A_pN94njs06_0;
	wire w_dff_A_zTvoK0eo4_0;
	wire w_dff_A_9Rvc39fk1_0;
	wire w_dff_A_dyuGMICT6_0;
	wire w_dff_A_0omNt4yn0_0;
	wire w_dff_A_0PqGSUCa3_0;
	wire w_dff_A_dzeWzO6E8_0;
	wire w_dff_A_InvzsMxT5_0;
	wire w_dff_A_e07vjjwd8_0;
	wire w_dff_A_7VtgAFAC2_0;
	wire w_dff_A_Bxd7xzdy4_0;
	wire w_dff_A_xODHA9ah0_0;
	wire w_dff_A_pRMp635i8_0;
	wire w_dff_A_yFeeqo8i6_0;
	wire w_dff_A_D1OIFUbg3_0;
	wire w_dff_A_3RniC67G8_0;
	wire w_dff_A_GQ7TLWlX5_0;
	wire w_dff_A_nn8qURut8_0;
	wire w_dff_A_ll4vw5e71_0;
	wire w_dff_A_ISoQoaIJ1_1;
	wire w_dff_A_kazzux2u8_2;
	wire w_dff_A_w9HYr66J4_0;
	wire w_dff_A_FvSOP7KV6_0;
	wire w_dff_A_43N3vsTT3_0;
	wire w_dff_A_ZYupGxZ83_0;
	wire w_dff_A_RxGa3VIE9_0;
	wire w_dff_A_2z9WHNuB5_0;
	wire w_dff_A_uezb728w2_0;
	wire w_dff_A_6NSavQqV6_0;
	wire w_dff_A_URIAhbao3_0;
	wire w_dff_A_Jd59PiaD2_0;
	wire w_dff_A_94EPOhq03_0;
	wire w_dff_A_iR2uoyDP3_0;
	wire w_dff_A_5U2JcT4S6_0;
	wire w_dff_A_wFlYTjpM2_0;
	wire w_dff_A_yAoCe94R7_0;
	wire w_dff_A_jNh70a8Q7_0;
	wire w_dff_A_JTQib3Qa8_0;
	wire w_dff_A_0CrUDDpE8_0;
	wire w_dff_A_GqDjidEL4_0;
	wire w_dff_A_VvkpVXp26_0;
	wire w_dff_A_HdapZFwp5_0;
	wire w_dff_A_uXtBycX77_0;
	wire w_dff_A_2HHX7coE5_0;
	wire w_dff_A_Y4EtgO005_0;
	wire w_dff_A_5ewLWf1x3_0;
	wire w_dff_A_aYMwcFEq6_1;
	wire w_dff_A_LtNAu88Z7_2;
	wire w_dff_A_5F9DBEBA3_0;
	wire w_dff_A_ULQI3dSY5_0;
	wire w_dff_A_mcrDvY0w8_0;
	wire w_dff_A_QeZdjYpp7_0;
	wire w_dff_A_2vJFH7uA8_0;
	wire w_dff_A_sGGiRhdj8_0;
	wire w_dff_A_mqLqVPta6_0;
	wire w_dff_A_i2KBoIBi3_0;
	wire w_dff_A_6AF8tcGX9_0;
	wire w_dff_A_r3rrGcI09_0;
	wire w_dff_A_drMLmGCL9_0;
	wire w_dff_A_1FeyGtDE7_0;
	wire w_dff_A_FCif0Lax2_0;
	wire w_dff_A_Ap4mlANs3_0;
	wire w_dff_A_4oDZ1FCG0_0;
	wire w_dff_A_YCP7jMKP2_0;
	wire w_dff_A_cksGFkhz1_0;
	wire w_dff_A_91wyghiS6_0;
	wire w_dff_A_TjezKelA1_0;
	wire w_dff_A_zeQpUz4m8_0;
	wire w_dff_A_3hgz5e1J0_0;
	wire w_dff_A_ULEY2Xh70_0;
	wire w_dff_A_feTdm7cL9_0;
	wire w_dff_A_GDWe2Ed28_1;
	wire w_dff_A_pUePyb2f4_2;
	wire w_dff_A_JZWCuGl19_0;
	wire w_dff_A_sYtQ0rJq6_0;
	wire w_dff_A_x9rTQskC1_0;
	wire w_dff_A_iy4Thptt3_0;
	wire w_dff_A_CSWz8Rh16_0;
	wire w_dff_A_NUknB0YH3_0;
	wire w_dff_A_3mMAn5rP5_0;
	wire w_dff_A_yzmVGExE3_0;
	wire w_dff_A_KZ4RsuBW9_0;
	wire w_dff_A_7MMh2dfC4_0;
	wire w_dff_A_7wMD8lrW8_0;
	wire w_dff_A_tTEfOe8G8_0;
	wire w_dff_A_G3tY7b388_0;
	wire w_dff_A_cP4hdsTT3_0;
	wire w_dff_A_3umympik8_0;
	wire w_dff_A_MHytO7VT9_0;
	wire w_dff_A_Rj0u3L2Y5_0;
	wire w_dff_A_jmfQ601j5_0;
	wire w_dff_A_ZBgEBTYf0_0;
	wire w_dff_A_YZK69PiR5_0;
	wire w_dff_A_779Ly5To1_0;
	wire w_dff_A_iwf7vElC1_1;
	wire w_dff_A_px4TwLna7_2;
	wire w_dff_A_jCGIzMeG0_0;
	wire w_dff_A_rpLt9Fpd9_0;
	wire w_dff_A_SPxXuECE0_0;
	wire w_dff_A_hxWcnJCZ1_0;
	wire w_dff_A_xlmJTAOT8_0;
	wire w_dff_A_jkvjEAHl9_0;
	wire w_dff_A_ufkRC2n31_0;
	wire w_dff_A_d0r6oMcr7_0;
	wire w_dff_A_YErHK3kd8_0;
	wire w_dff_A_5u1Lgjg41_0;
	wire w_dff_A_Fe2vuQfG0_0;
	wire w_dff_A_5Lex8d2O2_0;
	wire w_dff_A_VOALqQ4k4_0;
	wire w_dff_A_3Ld9aSWl2_0;
	wire w_dff_A_WKJmnlms2_0;
	wire w_dff_A_IYWSJVUQ9_0;
	wire w_dff_A_zbRK0Ysn1_0;
	wire w_dff_A_4QQPTkHp1_0;
	wire w_dff_A_lXR94XaA4_0;
	wire w_dff_A_vf10omxW1_1;
	wire w_dff_A_v08tLeep6_2;
	wire w_dff_A_7KpPilju2_0;
	wire w_dff_A_NIqqc0Ox9_0;
	wire w_dff_A_SL4UvMG77_0;
	wire w_dff_A_OqRlkAhm3_0;
	wire w_dff_A_R5IRv6W95_0;
	wire w_dff_A_Hz6uWMmA8_0;
	wire w_dff_A_mHD4qWy89_0;
	wire w_dff_A_qmhBJOhA2_0;
	wire w_dff_A_wQRDciC92_0;
	wire w_dff_A_MhQHdx9g9_0;
	wire w_dff_A_OMXtVIoo1_0;
	wire w_dff_A_87BUSuyJ4_0;
	wire w_dff_A_QmHmyN2l0_0;
	wire w_dff_A_tS1iXJKm9_0;
	wire w_dff_A_3JV8DRYs3_0;
	wire w_dff_A_oToKoT7i0_0;
	wire w_dff_A_bzzSIQF31_0;
	wire w_dff_A_eQlOczic5_1;
	wire w_dff_A_H17Bjt2h2_2;
	wire w_dff_A_Cqizgbsw6_0;
	wire w_dff_A_0pRyf39E5_0;
	wire w_dff_A_pqGuvdBE5_0;
	wire w_dff_A_shhzMjQP6_0;
	wire w_dff_A_uNRnbGGr9_0;
	wire w_dff_A_E78EoQLH3_0;
	wire w_dff_A_nHOhTHfi1_0;
	wire w_dff_A_F6zJR4kQ6_0;
	wire w_dff_A_O73bvBUS0_0;
	wire w_dff_A_CZPRDBnR1_0;
	wire w_dff_A_80NxXhQH0_0;
	wire w_dff_A_CoyyZRJp0_0;
	wire w_dff_A_p0w8nkSi7_0;
	wire w_dff_A_1lpFeTQs8_0;
	wire w_dff_A_Oeb4iY3b9_0;
	wire w_dff_A_dKDe0QPZ5_1;
	wire w_dff_A_DvKWN5fh7_2;
	wire w_dff_A_tDG3Qnmk9_0;
	wire w_dff_A_690nUmZT2_0;
	wire w_dff_A_6UXU6NRh0_0;
	wire w_dff_A_GKJYzaP06_0;
	wire w_dff_A_RtLgvyqS8_0;
	wire w_dff_A_wGPX2W1j9_0;
	wire w_dff_A_2zAM49FT7_0;
	wire w_dff_A_OZtLM20K6_0;
	wire w_dff_A_RDdpvEL42_0;
	wire w_dff_A_scRUgCMK7_0;
	wire w_dff_A_4rljsAHQ6_0;
	wire w_dff_A_YkYi6GKM5_0;
	wire w_dff_A_2UH2CFTH9_0;
	wire w_dff_A_3RUgPuw28_1;
	wire w_dff_A_X5hDfQDj5_2;
	wire w_dff_A_W75uVNnM6_0;
	wire w_dff_A_8ty9nFLM9_0;
	wire w_dff_A_9hHzXBpl7_0;
	wire w_dff_A_q2pGvRuu9_0;
	wire w_dff_A_v8v8RMUX2_0;
	wire w_dff_A_eazA6Cty5_0;
	wire w_dff_A_KDhbOBns9_0;
	wire w_dff_A_2nedHdpN9_0;
	wire w_dff_A_xMkIFcHq0_0;
	wire w_dff_A_gZJZmRfP0_0;
	wire w_dff_A_qj5HAMpT0_0;
	wire w_dff_A_0Nvok6OE8_1;
	wire w_dff_A_sokiXTn82_2;
	wire w_dff_A_nFyGUYEd9_0;
	wire w_dff_A_U3fbiXAi7_0;
	wire w_dff_A_AvZ2IZj87_0;
	wire w_dff_A_JTcRza669_0;
	wire w_dff_A_ojmxpyhq6_0;
	wire w_dff_A_tXUz8pSJ5_0;
	wire w_dff_A_wTMA7ou45_0;
	wire w_dff_A_s6i9fVwp6_0;
	wire w_dff_A_ZbpznAsK3_0;
	wire w_dff_A_GAQ3BWky2_1;
	wire w_dff_A_4x3nTySY4_2;
	wire w_dff_A_dgQ2v7Ka8_0;
	wire w_dff_A_obEASgJV0_0;
	wire w_dff_A_THC7F6sj7_0;
	wire w_dff_A_HKkXdrLj4_0;
	wire w_dff_A_ictpUbM78_0;
	wire w_dff_A_YbNHwdYE6_0;
	wire w_dff_A_SAPjTpMh1_0;
	wire w_dff_A_bOg8qe9P3_1;
	wire w_dff_A_bfPY2yka7_2;
	wire w_dff_B_qgd5TmgI4_3;
	wire w_dff_B_qFGeQJ162_3;
	wire w_dff_B_1uWchztE5_0;
	wire w_dff_A_mSXE5txn7_0;
	wire w_dff_A_7hvl0jIi3_0;
	wire w_dff_A_yoFFnUwE3_0;
	wire w_dff_A_dJ1rZgd00_1;
	wire w_dff_B_26h76l4t0_1;
	wire w_dff_B_cbfshor35_1;
	wire w_dff_A_b7ZXtC620_1;
	wire w_dff_A_EwX7zqbr3_2;
	wire w_dff_A_XQ7rHGXI6_2;
	wire w_dff_A_2RGpeNmG4_0;
	wire w_dff_B_j4T0AgN81_2;
	wire w_dff_B_bYJNWGcp4_2;
	wire w_dff_B_DfRfJ3bK4_2;
	wire w_dff_B_xV3L2C6S0_2;
	wire w_dff_B_mU8KX2pU1_2;
	wire w_dff_B_IK3LcRcX8_2;
	wire w_dff_B_54wJsXCZ3_2;
	wire w_dff_B_8YgzDuj16_2;
	wire w_dff_B_NEZyEFb88_2;
	wire w_dff_B_XHM7RemR6_2;
	wire w_dff_B_jd7RMWTP8_2;
	wire w_dff_B_W2ZBHAkE5_2;
	wire w_dff_B_Lm9OBGLG8_2;
	wire w_dff_B_rcAybTle5_2;
	wire w_dff_B_PRFY7O3c9_2;
	wire w_dff_B_vERN2gaO2_2;
	wire w_dff_B_PfR96urB4_2;
	wire w_dff_B_5hoGElMA3_2;
	wire w_dff_B_JI5mF0TP6_2;
	wire w_dff_B_Zt7e1kpL2_2;
	wire w_dff_B_05M2yTSO5_2;
	wire w_dff_B_zeXRbp1R3_2;
	wire w_dff_B_HuYJehbf1_2;
	wire w_dff_B_vtapNQv04_2;
	wire w_dff_B_w2uM7Xjk0_2;
	wire w_dff_B_7z2LuFvy4_2;
	wire w_dff_B_ir2jp4YY3_2;
	wire w_dff_B_LTz5XWUz2_2;
	wire w_dff_B_fINgTJaq6_2;
	wire w_dff_B_uOvMuQMc7_2;
	wire w_dff_B_871vyg922_2;
	wire w_dff_B_mE1Zy2sU9_2;
	wire w_dff_B_XkFNPjeQ5_2;
	wire w_dff_B_G2YSEwb05_2;
	wire w_dff_B_etIzj5896_2;
	wire w_dff_A_rMaboMKD7_0;
	wire w_dff_B_ZcdfPDIP9_2;
	wire w_dff_B_zEAdWz9j7_1;
	wire w_dff_B_uxGb2FZw7_2;
	wire w_dff_B_0CtX2aQn8_2;
	wire w_dff_B_gqI3gs5R0_2;
	wire w_dff_B_pOqvpxto7_2;
	wire w_dff_B_GM9vxiVN6_2;
	wire w_dff_B_TDJCfjJJ0_2;
	wire w_dff_B_MbLQsQzu0_2;
	wire w_dff_B_LdHs9k6t2_2;
	wire w_dff_B_7Z7WrGWx9_2;
	wire w_dff_B_DKYmxXIN1_2;
	wire w_dff_B_8pENd0yE5_2;
	wire w_dff_B_DV7KcakJ4_2;
	wire w_dff_B_5G5O4tAY5_2;
	wire w_dff_B_BhBgSvci0_2;
	wire w_dff_B_X2m81CUq2_2;
	wire w_dff_B_98JUuTyE8_2;
	wire w_dff_B_as2GFjCB3_2;
	wire w_dff_B_y5DIGxyD8_2;
	wire w_dff_B_pf9LINJP3_2;
	wire w_dff_B_azIu6PLv9_2;
	wire w_dff_B_ECf88KlO9_2;
	wire w_dff_B_7MgmOrwr1_2;
	wire w_dff_B_mgZhSM261_2;
	wire w_dff_B_TlewAGHq5_2;
	wire w_dff_B_2Nyxptkn9_2;
	wire w_dff_B_l3j2iUwR7_2;
	wire w_dff_B_GlrHFx7c9_2;
	wire w_dff_B_C2xiafOV4_2;
	wire w_dff_B_cCKohKyh5_2;
	wire w_dff_B_l8C2ByAj2_2;
	wire w_dff_A_qzgPrtGO7_1;
	wire w_dff_A_BJrHJgjF4_0;
	wire w_dff_A_qYJKegax7_0;
	wire w_dff_A_UiXGr92k1_0;
	wire w_dff_A_W6h5kWeR9_0;
	wire w_dff_A_tA04Wu2J0_0;
	wire w_dff_A_VvPFzFwC8_0;
	wire w_dff_A_KK9UUVl54_0;
	wire w_dff_A_EBmNu9Oy6_0;
	wire w_dff_A_kt3X1cE19_0;
	wire w_dff_A_umJctkA12_0;
	wire w_dff_A_HHGvKxhp7_0;
	wire w_dff_A_hDHH47Fi6_0;
	wire w_dff_A_4vgObg4A9_0;
	wire w_dff_A_Rpjy6oS47_0;
	wire w_dff_A_QJmZYqEV9_0;
	wire w_dff_A_fA4xHuXH3_0;
	wire w_dff_A_PLigeOWi8_0;
	wire w_dff_A_RAarvpgD9_0;
	wire w_dff_A_UgoKJSae5_0;
	wire w_dff_A_NZAsxVwn0_0;
	wire w_dff_A_9dF0jMfQ0_0;
	wire w_dff_A_bWFBy0420_0;
	wire w_dff_A_6JRJDj9P4_0;
	wire w_dff_A_vo4YJvxa3_0;
	wire w_dff_A_U6NdRyZB1_0;
	wire w_dff_A_K9vd1BE52_0;
	wire w_dff_A_X26fXPwE3_0;
	wire w_dff_A_CO6oBVJP9_0;
	wire w_dff_A_qN6gSYM48_0;
	wire w_dff_B_tdhjsvxw5_1;
	wire w_dff_B_QE2RFmPL0_2;
	wire w_dff_B_ZAk0Gr631_2;
	wire w_dff_B_uEqKH06t2_2;
	wire w_dff_B_N5zk9FHS4_2;
	wire w_dff_B_ZCwqaOg38_2;
	wire w_dff_B_A3mAc1jt2_2;
	wire w_dff_B_d7c6vFgR9_2;
	wire w_dff_B_GxW7UAtM8_2;
	wire w_dff_B_8FuUaeVB6_2;
	wire w_dff_B_3CS8Zprk9_2;
	wire w_dff_B_gtBI0k7n7_2;
	wire w_dff_B_04q9SLLh6_2;
	wire w_dff_B_IXcYr1ok6_2;
	wire w_dff_B_d3M1XEIT8_2;
	wire w_dff_B_qSNgsTXK3_2;
	wire w_dff_B_K033VI0H4_2;
	wire w_dff_B_NAH9VlkF0_2;
	wire w_dff_B_FAgdJ6M35_2;
	wire w_dff_B_F7kkwPo64_2;
	wire w_dff_B_DGOdcGys8_2;
	wire w_dff_B_qbpJxz6L6_2;
	wire w_dff_B_wvIK4g903_2;
	wire w_dff_B_jQ25XXm10_2;
	wire w_dff_B_6zgCuI5N9_2;
	wire w_dff_B_0jnZfbuD4_1;
	wire w_dff_B_d6JRT1Sj6_2;
	wire w_dff_B_F4eMiP946_2;
	wire w_dff_B_7beeHpPI5_2;
	wire w_dff_B_4RIWZMKQ9_2;
	wire w_dff_B_3VcQRmN99_2;
	wire w_dff_B_lJZefGct7_2;
	wire w_dff_B_toChjdRD8_2;
	wire w_dff_B_ORPnprfv7_2;
	wire w_dff_B_r3bPQwLu6_2;
	wire w_dff_B_DHfGuWza7_2;
	wire w_dff_B_kHAppI2U9_2;
	wire w_dff_B_W8PLt7xB4_2;
	wire w_dff_B_HNc09p799_2;
	wire w_dff_B_ZiISFO4e6_2;
	wire w_dff_B_IMh2db9w0_2;
	wire w_dff_B_nNO7I5rT4_2;
	wire w_dff_B_vAFM8nZu5_2;
	wire w_dff_B_r8pVk9yJ3_2;
	wire w_dff_B_TIh27FCV9_2;
	wire w_dff_B_9guNURWa8_2;
	wire w_dff_B_Gai22cUS9_2;
	wire w_dff_B_dD5wDP8N1_2;
	wire w_dff_B_Wmw0vaVP3_1;
	wire w_dff_B_E6csAyxh8_2;
	wire w_dff_B_PEBJSwCH4_2;
	wire w_dff_B_nJ6zdzMn2_2;
	wire w_dff_B_fGI7bQZ27_2;
	wire w_dff_B_Ul4N78Sf0_2;
	wire w_dff_B_o3rwXkbv3_2;
	wire w_dff_B_itXsQoc02_2;
	wire w_dff_B_WVbB8UgY6_2;
	wire w_dff_B_0GVjnti59_2;
	wire w_dff_B_uk17SVWN7_2;
	wire w_dff_B_s9CxG9Br1_2;
	wire w_dff_B_gHJ0ImCt1_2;
	wire w_dff_B_Ot0FYI356_2;
	wire w_dff_B_xAZXpZzQ1_2;
	wire w_dff_B_N3Gsflrv8_2;
	wire w_dff_B_ZcQzw2tB0_2;
	wire w_dff_B_um5QauEF7_2;
	wire w_dff_B_plqHSaSK6_2;
	wire w_dff_B_IYScNTsq6_2;
	wire w_dff_B_v4zCLJrf9_2;
	wire w_dff_B_mNrhr0kP7_1;
	wire w_dff_B_8uU0orkr0_2;
	wire w_dff_B_xdTh0JsV9_2;
	wire w_dff_B_ZCY2u8bj9_2;
	wire w_dff_B_uQiFdHlv7_2;
	wire w_dff_B_fGTMR4Om5_2;
	wire w_dff_B_ZolFk9wV5_2;
	wire w_dff_B_uMHjTHCD7_2;
	wire w_dff_B_lSRmAsPP8_2;
	wire w_dff_B_aSolrUlR4_2;
	wire w_dff_B_sLtem57U4_2;
	wire w_dff_B_h2M5yWJp4_2;
	wire w_dff_B_3XP1Phog8_2;
	wire w_dff_B_IPSYJc9R2_2;
	wire w_dff_B_Hn9nAkO59_2;
	wire w_dff_B_423A2rfK5_2;
	wire w_dff_B_XdpRRCVC1_2;
	wire w_dff_B_xZRDx6Bt5_2;
	wire w_dff_B_2aqVfDn05_2;
	wire w_dff_B_qGJNeFyw7_1;
	wire w_dff_B_kwKlTODZ5_2;
	wire w_dff_B_SwkXeJ1I6_2;
	wire w_dff_B_m4SnrpPw0_2;
	wire w_dff_B_AL2yACLO7_2;
	wire w_dff_B_o732N5oX6_2;
	wire w_dff_B_1rvJfPSJ5_2;
	wire w_dff_B_ikLtOuxI9_2;
	wire w_dff_B_ylp4eRFb0_2;
	wire w_dff_B_r0DdNQZO0_2;
	wire w_dff_B_x00hC7cC4_2;
	wire w_dff_B_CaJO27J65_2;
	wire w_dff_B_x11CjgDl4_2;
	wire w_dff_B_zeoYnGYG9_2;
	wire w_dff_B_bvwz06ZQ6_2;
	wire w_dff_B_XYEyF6it7_2;
	wire w_dff_B_TL6QGUTC1_2;
	wire w_dff_B_O4itNlQT3_1;
	wire w_dff_B_SR5M0VzB2_2;
	wire w_dff_B_XWv2B1TI7_2;
	wire w_dff_B_H2hSsFwG9_2;
	wire w_dff_B_UukRbFo74_2;
	wire w_dff_B_ONDBlnSX9_2;
	wire w_dff_B_J3HNgRAf3_2;
	wire w_dff_B_CzZuSfpC0_2;
	wire w_dff_B_8EGuyn8o5_2;
	wire w_dff_B_Ok4Ld4ha5_2;
	wire w_dff_B_uE7FpfDF3_2;
	wire w_dff_B_g7vvmbgS7_2;
	wire w_dff_B_6UAniggy6_2;
	wire w_dff_B_GyVhD9yX8_2;
	wire w_dff_B_P7GxG97t3_2;
	wire w_dff_B_mxWU2CBS8_1;
	wire w_dff_B_Zm67YdwU8_2;
	wire w_dff_B_g1MQVclp4_2;
	wire w_dff_B_Sv2u7VZ55_2;
	wire w_dff_B_oUyA7ZVi8_2;
	wire w_dff_B_yF7lTfJJ9_2;
	wire w_dff_B_n5xq0kya3_2;
	wire w_dff_B_lTcFdM6T7_2;
	wire w_dff_B_y9ZTsqQz0_2;
	wire w_dff_B_sHZYPjDW3_2;
	wire w_dff_B_QNXXIVyt4_2;
	wire w_dff_B_IAWsEFu13_2;
	wire w_dff_B_669JR3NH1_2;
	wire w_dff_B_Dk6URZcJ7_1;
	wire w_dff_B_3Atefzp26_2;
	wire w_dff_B_Fufmaz4c0_2;
	wire w_dff_B_6NCIYT4J2_2;
	wire w_dff_B_0UlYdXqn4_2;
	wire w_dff_B_Ppt82TVn7_2;
	wire w_dff_B_5rQPrQYp5_2;
	wire w_dff_B_NcTAceBg3_2;
	wire w_dff_B_juyQzPl45_2;
	wire w_dff_B_EknasaLQ9_2;
	wire w_dff_B_o5szB85e1_2;
	wire w_dff_B_bSS4JKmy4_1;
	wire w_dff_B_RGFVFglE4_2;
	wire w_dff_B_55E2HOtn8_2;
	wire w_dff_B_KnVzLke91_2;
	wire w_dff_B_IABejzyF6_2;
	wire w_dff_B_SxkHWhwO0_2;
	wire w_dff_B_ZFW7P50Q9_2;
	wire w_dff_B_zV0An42L0_2;
	wire w_dff_B_0YPYM2yI9_2;
	wire w_dff_B_KV0W7Hdu4_2;
	wire w_dff_B_SxyvgrUB3_1;
	wire w_dff_B_0tChY7Uu8_2;
	wire w_dff_B_oYHn7muD7_2;
	wire w_dff_B_ehy3hBab9_2;
	wire w_dff_B_ielkX7kY1_2;
	wire w_dff_B_DwabZDaX7_2;
	wire w_dff_B_d3eFCLjg4_2;
	wire w_dff_B_r8aFdsh71_2;
	wire w_dff_B_xm84fC9V6_1;
	wire w_dff_B_IADcx8xB8_1;
	wire w_dff_B_ZW6ADBYo1_1;
	wire w_dff_B_BztZO27i2_1;
	wire w_dff_B_QzidDl7h9_2;
	wire w_dff_B_QXdIKbgG8_2;
	wire w_dff_B_CZm2vIc71_2;
	wire w_dff_B_DMlKtyFT9_2;
	wire w_dff_B_VuZ7sJNf6_0;
	wire w_dff_A_MOenS5Y47_1;
	wire w_dff_A_RCAO2G978_1;
	wire w_dff_A_RUhPeT7s8_1;
	wire w_dff_A_Zns8hL4f9_2;
	wire w_dff_A_7OiKETeF1_2;
	wire w_dff_A_2DXqsfki9_0;
	wire w_dff_B_4bprLLu56_1;
	wire w_dff_B_HQ0398zs6_1;
	wire w_dff_B_rVfDrSbl7_2;
	wire w_dff_B_OUR5TpkR0_2;
	wire w_dff_B_eh1kDnH91_2;
	wire w_dff_B_0pIJejLK6_2;
	wire w_dff_B_fVgrTWcy5_2;
	wire w_dff_B_0d7leuKp4_2;
	wire w_dff_B_DZN7eg5X7_2;
	wire w_dff_B_im3r9vEP1_2;
	wire w_dff_B_shpohSec9_2;
	wire w_dff_B_z4qg006d6_2;
	wire w_dff_B_yi5zyAAe4_2;
	wire w_dff_B_OcxFxGup5_2;
	wire w_dff_B_0yLlVIZG8_2;
	wire w_dff_B_g7k0XUje4_2;
	wire w_dff_B_GV4HnXOn4_2;
	wire w_dff_B_0j2KN2Z04_2;
	wire w_dff_B_g9qiRDzU0_2;
	wire w_dff_B_WaM41Jar5_2;
	wire w_dff_B_2nsL2mIH6_2;
	wire w_dff_B_EI9rOSKt0_2;
	wire w_dff_B_IQ69olqx0_2;
	wire w_dff_B_1kY86yeo3_2;
	wire w_dff_B_OfwxjwD78_2;
	wire w_dff_B_31ez3Xxf3_2;
	wire w_dff_B_OnzbbnUu9_2;
	wire w_dff_B_d3DbEaqy9_2;
	wire w_dff_B_z20hfsCO1_2;
	wire w_dff_B_ZcSaZECM3_2;
	wire w_dff_B_95Dk3xZG3_2;
	wire w_dff_B_5QIVyAeT4_2;
	wire w_dff_B_LszWiyAZ9_2;
	wire w_dff_B_l43tMi885_2;
	wire w_dff_B_qxcq6ioB7_2;
	wire w_dff_B_UIK0X4Nc0_2;
	wire w_dff_B_dkaftnOp3_2;
	wire w_dff_B_HDeeE3zj8_2;
	wire w_dff_B_ut7Gdpue6_2;
	wire w_dff_B_8ML7WXKy8_2;
	wire w_dff_B_wVJrfpMj4_2;
	wire w_dff_B_rO9EYn8N0_2;
	wire w_dff_B_UbLV6dIC8_2;
	wire w_dff_B_SjX8Pkym2_2;
	wire w_dff_B_y31zMqjC0_2;
	wire w_dff_B_DEeYucqF6_2;
	wire w_dff_B_VICmKp3s8_2;
	wire w_dff_B_zj6j3PJl0_2;
	wire w_dff_B_lPOY5AIU6_2;
	wire w_dff_B_iulyastL8_2;
	wire w_dff_B_t9fdieQX9_2;
	wire w_dff_B_9UQMQQje6_2;
	wire w_dff_B_4HGfjpRm0_2;
	wire w_dff_B_FnRakgzV5_2;
	wire w_dff_B_TtRhlFxB1_2;
	wire w_dff_B_a8ULsxYn6_2;
	wire w_dff_B_20Hn3ifm2_2;
	wire w_dff_B_Ra7rGvSp3_2;
	wire w_dff_B_khnGhDRn9_2;
	wire w_dff_B_kwoqfqHK8_2;
	wire w_dff_B_NrlJz5gm7_2;
	wire w_dff_B_fi0giJp52_2;
	wire w_dff_B_9XSGrxv58_2;
	wire w_dff_B_oRg94UzK3_2;
	wire w_dff_B_WQnTw4us2_2;
	wire w_dff_B_0ajdEipX5_2;
	wire w_dff_B_tVRV7OsE9_2;
	wire w_dff_B_eg24WkAQ6_2;
	wire w_dff_B_0Y6pU22K5_2;
	wire w_dff_B_5BmTqeRt2_2;
	wire w_dff_B_yOVGUYnu7_1;
	wire w_dff_B_oMu2hVNG1_2;
	wire w_dff_B_jTqIiLCG7_2;
	wire w_dff_B_E9atFrem2_2;
	wire w_dff_B_kO3khuXJ1_2;
	wire w_dff_B_9Rt4fsWD2_2;
	wire w_dff_B_QPKubA1A4_2;
	wire w_dff_B_bSn9ApwM1_2;
	wire w_dff_B_lyLk7HRX3_2;
	wire w_dff_B_1QqkWXZU5_2;
	wire w_dff_B_8Gn8jUY98_2;
	wire w_dff_B_pHqETEZS1_2;
	wire w_dff_B_Aq9UJTwB0_2;
	wire w_dff_B_zHdONj456_2;
	wire w_dff_B_iHNk5Cbt5_2;
	wire w_dff_B_yhbpxAeA1_2;
	wire w_dff_B_YxOVq6wy2_2;
	wire w_dff_B_qFjfjO0G7_2;
	wire w_dff_B_uXaoQqx24_2;
	wire w_dff_B_vZC20l9v4_2;
	wire w_dff_B_paTa60LQ3_2;
	wire w_dff_B_fjui4HUZ8_2;
	wire w_dff_B_C4UnGJQX5_2;
	wire w_dff_B_wKuCAcoD5_2;
	wire w_dff_B_WxjeCSRy0_2;
	wire w_dff_B_50ZXxNf37_2;
	wire w_dff_B_yoJ1bUnw9_2;
	wire w_dff_B_BbhDxqc18_1;
	wire w_dff_B_EPVCfF0o7_2;
	wire w_dff_B_7cfyAm1b4_2;
	wire w_dff_B_RYL4EtQe0_2;
	wire w_dff_B_J7O2bJi86_2;
	wire w_dff_B_8cokMvvD1_2;
	wire w_dff_B_i6vpuMVL1_2;
	wire w_dff_B_bQlFTCX68_2;
	wire w_dff_B_mgQUN2Vv2_2;
	wire w_dff_B_U7lemMSr0_2;
	wire w_dff_B_tKcxuTBc5_2;
	wire w_dff_B_JDKuEmjY7_2;
	wire w_dff_B_lYqRj3aA4_2;
	wire w_dff_B_RSYX8dfh4_2;
	wire w_dff_B_HyYmUasu3_2;
	wire w_dff_B_GpYfbHrv9_2;
	wire w_dff_B_gCh1ZfjT8_2;
	wire w_dff_B_s7oWDwCD0_2;
	wire w_dff_B_bYBsYAXr2_2;
	wire w_dff_B_tHQkTJFO3_2;
	wire w_dff_B_Ig1ukQAh9_2;
	wire w_dff_B_f8GuRuGt0_2;
	wire w_dff_B_mtaOLY4K6_2;
	wire w_dff_B_eGaIVF2z0_2;
	wire w_dff_B_32BBUETR6_2;
	wire w_dff_B_jan9yoBt7_1;
	wire w_dff_B_QefQ0Vzc8_2;
	wire w_dff_B_EL7OHtVR9_2;
	wire w_dff_B_sPgxBzVE7_2;
	wire w_dff_B_WEC35h5t6_2;
	wire w_dff_B_P7huY2LL6_2;
	wire w_dff_B_tYv9De148_2;
	wire w_dff_B_m4lMnMzN0_2;
	wire w_dff_B_oCvDsXSc9_2;
	wire w_dff_B_OsOzXHUD2_2;
	wire w_dff_B_NWwma4Et0_2;
	wire w_dff_B_fMfR0em89_2;
	wire w_dff_B_O1raQNuD4_2;
	wire w_dff_B_43l9vTg94_2;
	wire w_dff_B_jcmNCKaf0_2;
	wire w_dff_B_ZWMPaf6m1_2;
	wire w_dff_B_nDKEzlx21_2;
	wire w_dff_B_ZeBBeoNo6_2;
	wire w_dff_B_zHdj9PRa7_2;
	wire w_dff_B_aD7xgN5p8_2;
	wire w_dff_B_ghkkU9EK4_2;
	wire w_dff_B_7XrSf3Kd8_2;
	wire w_dff_B_Ge66VRId2_2;
	wire w_dff_B_NjSLxxAi9_1;
	wire w_dff_B_0fm2pvKd1_2;
	wire w_dff_B_gOinbKHi9_2;
	wire w_dff_B_P1nDAfVW4_2;
	wire w_dff_B_jaiYtPvQ5_2;
	wire w_dff_B_ZBhRdYHg0_2;
	wire w_dff_B_sDMuL2AP2_2;
	wire w_dff_B_ZovVYjIq2_2;
	wire w_dff_B_mEMkvezv5_2;
	wire w_dff_B_wRk4F03L6_2;
	wire w_dff_B_UXcQQUlj7_2;
	wire w_dff_B_IDHaq1Xc3_2;
	wire w_dff_B_nzb8FYZJ4_2;
	wire w_dff_B_TWuDv1Zn6_2;
	wire w_dff_B_Nu0zq7kP8_2;
	wire w_dff_B_yeAU6gWp0_2;
	wire w_dff_B_3tIvfcNf7_2;
	wire w_dff_B_BjlvYQhT3_2;
	wire w_dff_B_AlUyikoN8_2;
	wire w_dff_B_bn6AZRWZ8_2;
	wire w_dff_B_jZmxLYdm6_2;
	wire w_dff_B_uqn7ykRC9_1;
	wire w_dff_B_3PRDOd840_2;
	wire w_dff_B_Nmm5tsaQ3_2;
	wire w_dff_B_66kp1h185_2;
	wire w_dff_B_2QyH3EDX1_2;
	wire w_dff_B_GYXaY3jF1_2;
	wire w_dff_B_Xbdt1keg6_2;
	wire w_dff_B_nxx84m0C9_2;
	wire w_dff_B_muiRi0J69_2;
	wire w_dff_B_MweqWHDe4_2;
	wire w_dff_B_LYJRX0Of8_2;
	wire w_dff_B_iidRc1wU2_2;
	wire w_dff_B_2SywCMjB9_2;
	wire w_dff_B_ImvNnBDr2_2;
	wire w_dff_B_mp39UK9t7_2;
	wire w_dff_B_wWR30lxS2_2;
	wire w_dff_B_75CQSFLO5_2;
	wire w_dff_B_BrbHYZtq1_2;
	wire w_dff_B_ESOkehGZ8_2;
	wire w_dff_B_DADHk8B11_1;
	wire w_dff_B_rngTF36W5_2;
	wire w_dff_B_vxPAZSQT2_2;
	wire w_dff_B_pOzWmgTj2_2;
	wire w_dff_B_2Smr4jtq5_2;
	wire w_dff_B_cRro3xIJ7_2;
	wire w_dff_B_2m9yRjZT5_2;
	wire w_dff_B_BwelrUXL4_2;
	wire w_dff_B_hE3pszSi8_2;
	wire w_dff_B_LTlBw1895_2;
	wire w_dff_B_vdoNNJG76_2;
	wire w_dff_B_XkAZ7FFS1_2;
	wire w_dff_B_dPCNRQlL7_2;
	wire w_dff_B_1rDuuBOu5_2;
	wire w_dff_B_JSPN5e8Y2_2;
	wire w_dff_B_KMEdhYIr1_2;
	wire w_dff_B_TVLIDS2Y9_2;
	wire w_dff_B_uYzApxJz9_1;
	wire w_dff_B_LR37DUxK7_2;
	wire w_dff_B_nrKd9pOE6_2;
	wire w_dff_B_EFeoN9f90_2;
	wire w_dff_B_33g02Ddm9_2;
	wire w_dff_B_f6wMn9GJ3_2;
	wire w_dff_B_6703W9K22_2;
	wire w_dff_B_iq5urRMH3_2;
	wire w_dff_B_w9PQPxu29_2;
	wire w_dff_B_Uf5WZZVs4_2;
	wire w_dff_B_V5KTX8M17_2;
	wire w_dff_B_EFP6BrTs5_2;
	wire w_dff_B_hHuZHrLA4_2;
	wire w_dff_B_jrpIEsyb2_2;
	wire w_dff_B_MGReRU7o3_2;
	wire w_dff_B_TIRuYEFC5_1;
	wire w_dff_B_ADlkfaBT0_2;
	wire w_dff_B_8riLP2J56_2;
	wire w_dff_B_qIFAkXQd9_2;
	wire w_dff_B_cxN66kwZ5_2;
	wire w_dff_B_hh2qU7rz7_2;
	wire w_dff_B_Bp5l5lz53_2;
	wire w_dff_B_TXqGHLxH2_2;
	wire w_dff_B_sN9U3zfN4_2;
	wire w_dff_B_PkOqJCLN3_2;
	wire w_dff_B_6kGhrfXn7_2;
	wire w_dff_B_wpMqGPca1_2;
	wire w_dff_B_Z8BhLEVE3_2;
	wire w_dff_B_DwjbHO0w1_1;
	wire w_dff_B_lFgjC9cs2_2;
	wire w_dff_B_FoT90ABF2_2;
	wire w_dff_B_X8NI0hMe0_2;
	wire w_dff_B_RSeWZT0v9_2;
	wire w_dff_B_hiLpQbpC1_2;
	wire w_dff_B_hTOVazCx9_2;
	wire w_dff_B_OeB7QDbi6_2;
	wire w_dff_B_z6rdy2TZ7_2;
	wire w_dff_B_ofmkEbZo1_2;
	wire w_dff_B_M5SDinXi6_2;
	wire w_dff_B_ZVn1JATL0_1;
	wire w_dff_B_CSHfwZK40_2;
	wire w_dff_B_v4tjxi2c9_2;
	wire w_dff_B_tKhnYXT06_2;
	wire w_dff_B_GTq1WUGl4_2;
	wire w_dff_B_y5b8JW3C0_2;
	wire w_dff_B_undiNxAR0_2;
	wire w_dff_B_cx3VEgZ42_2;
	wire w_dff_B_xmctGBj18_2;
	wire w_dff_B_TOOe7Jno0_2;
	wire w_dff_B_nwOQFSQ28_1;
	wire w_dff_B_t4ge3YhN4_2;
	wire w_dff_B_YoBF9TRb0_2;
	wire w_dff_B_l96uTqkB8_2;
	wire w_dff_B_Fxt6WSZz7_2;
	wire w_dff_B_nNtLFeVt4_2;
	wire w_dff_B_GK5VE46Q3_1;
	wire w_dff_B_vn3oQZHB7_0;
	wire w_dff_B_JHv1FRYm4_2;
	wire w_dff_B_GVY0OuzW2_2;
	wire w_dff_B_mHt9CsSX7_2;
	wire w_dff_B_I530oxMV5_1;
	wire w_dff_B_tNXDlT0N2_1;
	wire w_dff_A_ofpJNDQw4_0;
	wire w_dff_A_kmyc9HRq1_0;
	wire w_dff_B_TRezTEAG8_2;
	wire w_dff_B_3D2mMVj74_2;
	wire w_dff_B_cEx3tPYS7_1;
	wire w_dff_B_7UkinoS60_2;
	wire w_dff_B_6c18BDlQ0_2;
	wire w_dff_B_SdsxSNPh9_2;
	wire w_dff_B_TxGXkzvz5_2;
	wire w_dff_B_4KYFoQxi0_2;
	wire w_dff_B_lQ2G17Qz8_2;
	wire w_dff_B_9TD4OPUa6_2;
	wire w_dff_B_fNLJi2wq1_2;
	wire w_dff_B_3rR88h1H2_2;
	wire w_dff_B_DfGf5iQS9_2;
	wire w_dff_B_NE7dULgf9_2;
	wire w_dff_B_6RbOI03q7_2;
	wire w_dff_B_TIhBHJN38_2;
	wire w_dff_B_rUM1Tyhb4_2;
	wire w_dff_B_R8UWnzjE2_2;
	wire w_dff_B_04C07ge85_2;
	wire w_dff_B_5Ho9yZNc3_2;
	wire w_dff_B_vvrzDFV91_2;
	wire w_dff_B_0EluVG4F3_2;
	wire w_dff_B_3krL4CMp1_2;
	wire w_dff_B_NQtN0yqy5_2;
	wire w_dff_B_AWNRC3NM5_2;
	wire w_dff_B_g4ISwAUV5_2;
	wire w_dff_B_h22KO64B1_2;
	wire w_dff_B_XCzw0RSu3_2;
	wire w_dff_B_mfrlD0bf7_2;
	wire w_dff_B_itqNusvO0_2;
	wire w_dff_B_c6YNWpel9_2;
	wire w_dff_B_LdHS9SiW6_2;
	wire w_dff_B_BSThKHTZ2_2;
	wire w_dff_B_ce2nX3sI9_2;
	wire w_dff_B_L82pt5IS1_2;
	wire w_dff_B_rX4lAxbJ7_2;
	wire w_dff_B_n79MyZ8t5_2;
	wire w_dff_B_akaHYtU43_2;
	wire w_dff_B_NAWMwQTb3_1;
	wire w_dff_A_KykJmTCb5_1;
	wire w_dff_B_tV69P8c58_1;
	wire w_dff_B_08yCCRl85_2;
	wire w_dff_B_ega2IOAx1_2;
	wire w_dff_B_0umbl25E4_2;
	wire w_dff_B_k3nTJ9lF0_2;
	wire w_dff_B_aCZWGj4y9_2;
	wire w_dff_B_gn7HQ4dy4_2;
	wire w_dff_B_VoN6N6tk7_2;
	wire w_dff_B_F4PEiccT8_2;
	wire w_dff_B_e5iOJsHv3_2;
	wire w_dff_B_MPYbmmth5_2;
	wire w_dff_B_KSKOQreb9_2;
	wire w_dff_B_gNcDbPP20_2;
	wire w_dff_B_Q4qaNwBi7_2;
	wire w_dff_B_sWz74AKi9_2;
	wire w_dff_B_VntqsTvm2_2;
	wire w_dff_B_JaYEiOnw1_2;
	wire w_dff_B_JCp4qxlc8_2;
	wire w_dff_B_Vk6Y2Xq67_2;
	wire w_dff_B_LCS3EVqP8_2;
	wire w_dff_B_5Mp9lluc6_2;
	wire w_dff_B_twsH7dNa2_2;
	wire w_dff_B_EAR6JjCZ8_2;
	wire w_dff_B_7R9ngLxZ5_2;
	wire w_dff_B_hjvq3IXl3_2;
	wire w_dff_B_oEOBnXxC6_2;
	wire w_dff_B_zRIZoJKA2_2;
	wire w_dff_B_opiGyJHv5_2;
	wire w_dff_B_w8eQaxiw6_2;
	wire w_dff_B_TyuHfqsA3_2;
	wire w_dff_B_VjKKWoOF8_2;
	wire w_dff_B_43rU9oyq8_2;
	wire w_dff_B_isMwcS1w1_1;
	wire w_dff_B_jqSPLVzL8_2;
	wire w_dff_B_78yUqbDB2_2;
	wire w_dff_B_1kAW4RxE4_2;
	wire w_dff_B_Tf94WgGA3_2;
	wire w_dff_B_8bck2Qux5_2;
	wire w_dff_B_tnlR70Fh9_2;
	wire w_dff_B_1xSKL27U1_2;
	wire w_dff_B_1N0rZ2cL1_2;
	wire w_dff_B_U15Kks6r0_2;
	wire w_dff_B_miGCYZ6K1_2;
	wire w_dff_B_BYAOEYoV4_2;
	wire w_dff_B_VWLmRA2L7_2;
	wire w_dff_B_kBvRDchj5_2;
	wire w_dff_B_JBfInPp25_2;
	wire w_dff_B_fHX28qMm4_2;
	wire w_dff_B_3hqzMtGP8_2;
	wire w_dff_B_z7xVZdgB6_2;
	wire w_dff_B_p5BLpNmf8_2;
	wire w_dff_B_l5mYCSmb1_2;
	wire w_dff_B_oWCfsRT29_2;
	wire w_dff_B_Eag7T3Go0_2;
	wire w_dff_B_KGB44b8p5_2;
	wire w_dff_B_7FiuL1fx8_2;
	wire w_dff_B_tXmocK9L0_2;
	wire w_dff_B_LYmXnR0D6_2;
	wire w_dff_B_FUBlvQcc2_2;
	wire w_dff_B_Hh2EdLSE0_2;
	wire w_dff_B_69xcZT3g0_2;
	wire w_dff_B_Bm80gPTd6_1;
	wire w_dff_B_zM9DSR5m2_2;
	wire w_dff_B_otEsRPSG3_2;
	wire w_dff_B_1v9u5R3z3_2;
	wire w_dff_B_aZZ3vSDF5_2;
	wire w_dff_B_5ociFwIS0_2;
	wire w_dff_B_GrkhuzJ79_2;
	wire w_dff_B_2fvCIHTW9_2;
	wire w_dff_B_jSEuOTFR6_2;
	wire w_dff_B_fiqUj9wA1_2;
	wire w_dff_B_YDAYBLck8_2;
	wire w_dff_B_psnTPa0Z9_2;
	wire w_dff_B_yv0PcRP04_2;
	wire w_dff_B_bt7SzeB15_2;
	wire w_dff_B_NrTWawmi1_2;
	wire w_dff_B_0ZyU1zqh9_2;
	wire w_dff_B_AH3T2WJe9_2;
	wire w_dff_B_ZJXBQGRB7_2;
	wire w_dff_B_mMXYx8nk0_2;
	wire w_dff_B_Ih4QYTi56_2;
	wire w_dff_B_gSG37k7E7_2;
	wire w_dff_B_TyIA3mho0_2;
	wire w_dff_B_eSBkTehi6_2;
	wire w_dff_B_sjTn3Y0B7_2;
	wire w_dff_B_0ZoEKReq9_2;
	wire w_dff_B_W5g7uig16_1;
	wire w_dff_B_Iir1l9Dp0_2;
	wire w_dff_B_HFdagoan1_2;
	wire w_dff_B_cg6OqpNX8_2;
	wire w_dff_B_X8P0Gi0x9_2;
	wire w_dff_B_ILuCj0TM5_2;
	wire w_dff_B_MmafUwET9_2;
	wire w_dff_B_0DHi9rko1_2;
	wire w_dff_B_qE3pPuZD4_2;
	wire w_dff_B_HgOBbvJq6_2;
	wire w_dff_B_Xzay8MMW1_2;
	wire w_dff_B_ZadAQLYB2_2;
	wire w_dff_B_LNzFBwBl0_2;
	wire w_dff_B_jtqDpEpY8_2;
	wire w_dff_B_urQcLKTw6_2;
	wire w_dff_B_4zTlFqWa8_2;
	wire w_dff_B_makkpbhy1_2;
	wire w_dff_B_pSpKKRGM7_2;
	wire w_dff_B_TztNTQIm8_2;
	wire w_dff_B_nQIo6htB5_2;
	wire w_dff_B_iKu78UdK2_2;
	wire w_dff_B_0JwzWpsh1_2;
	wire w_dff_B_JClOxoUf1_2;
	wire w_dff_B_xYzFwxws2_1;
	wire w_dff_B_HTn8MndJ7_2;
	wire w_dff_B_GDrzHuKv3_2;
	wire w_dff_B_xfuaUkHC2_2;
	wire w_dff_B_ZgIRalUH6_2;
	wire w_dff_B_Zsz8LbIJ2_2;
	wire w_dff_B_BsRFxe4h0_2;
	wire w_dff_B_yySsxa9Q5_2;
	wire w_dff_B_AvCstIac7_2;
	wire w_dff_B_vVqxZcrC7_2;
	wire w_dff_B_4w0GsZBl6_2;
	wire w_dff_B_0DbbQjY77_2;
	wire w_dff_B_WbYEeDaZ9_2;
	wire w_dff_B_WkaWoqEY2_2;
	wire w_dff_B_EGX2etiJ9_2;
	wire w_dff_B_ogxpMXUR8_2;
	wire w_dff_B_uMQeDKnK0_2;
	wire w_dff_B_M4mJ7PxG7_2;
	wire w_dff_B_Dlr1YPDj2_2;
	wire w_dff_B_NhRtzx3h1_2;
	wire w_dff_B_G0y1hWVS6_2;
	wire w_dff_B_g5xYgFsp1_1;
	wire w_dff_B_oGO7mV1f8_2;
	wire w_dff_B_a05sQuiN5_2;
	wire w_dff_B_3Zl9v8QY2_2;
	wire w_dff_B_ktCushNk5_2;
	wire w_dff_B_92LUl3xV9_2;
	wire w_dff_B_z54okmfN2_2;
	wire w_dff_B_WmPwmEBH4_2;
	wire w_dff_B_2PPyRgBE5_2;
	wire w_dff_B_EWXT9pjb2_2;
	wire w_dff_B_Cd679bam3_2;
	wire w_dff_B_23lbCNkt2_2;
	wire w_dff_B_FLalwGIO4_2;
	wire w_dff_B_8IgrJCwc7_2;
	wire w_dff_B_EP1cTlPZ4_2;
	wire w_dff_B_Q7txkeJv4_2;
	wire w_dff_B_igt6yA2B5_2;
	wire w_dff_B_Y11jGgSH6_2;
	wire w_dff_B_VC4cduzu1_2;
	wire w_dff_B_1cPflRMl6_1;
	wire w_dff_B_lQuST4Wq9_2;
	wire w_dff_B_oD8ESpb73_2;
	wire w_dff_B_ewdMYlzB0_2;
	wire w_dff_B_QPcz9Fjk0_2;
	wire w_dff_B_88gOg1RB2_2;
	wire w_dff_B_0byU5bLA9_2;
	wire w_dff_B_lyT8jWWI9_2;
	wire w_dff_B_2LlqdzRq8_2;
	wire w_dff_B_1hXrFyqf1_2;
	wire w_dff_B_oC2zEpRx6_2;
	wire w_dff_B_AJV5VVpG4_2;
	wire w_dff_B_IauWHviK7_2;
	wire w_dff_B_6SioGfHX3_2;
	wire w_dff_B_oPqhnOSV7_2;
	wire w_dff_B_XnCFEuYz0_2;
	wire w_dff_B_RwsypYQB6_2;
	wire w_dff_B_KAUL5l4Y9_1;
	wire w_dff_B_4PnBuiIr8_2;
	wire w_dff_B_jjGp7l2O7_2;
	wire w_dff_B_gNAIgqb93_2;
	wire w_dff_B_odIHAG0E6_2;
	wire w_dff_B_SgMjPHcc9_2;
	wire w_dff_B_lPP0xdx58_2;
	wire w_dff_B_WsBLMzPU7_2;
	wire w_dff_B_PWmMLnaI0_2;
	wire w_dff_B_ekCqA8O74_2;
	wire w_dff_B_atYf08Cx5_2;
	wire w_dff_B_0N2zsqDj5_2;
	wire w_dff_B_MIiODms32_2;
	wire w_dff_B_BvjHOT067_2;
	wire w_dff_B_ioksKqhM3_2;
	wire w_dff_B_DXjHtJBZ6_1;
	wire w_dff_B_CFowmArr3_2;
	wire w_dff_B_wXFRrzH93_2;
	wire w_dff_B_pCKaer9d2_2;
	wire w_dff_B_XWvV3Zr30_2;
	wire w_dff_B_kQNePC2n0_2;
	wire w_dff_B_nUvdRr6R0_2;
	wire w_dff_B_TYFYL5hm1_2;
	wire w_dff_B_9dBaEDsj5_2;
	wire w_dff_B_XOGFjnUO3_2;
	wire w_dff_B_zWQw8quC7_2;
	wire w_dff_B_nQoFuduk2_2;
	wire w_dff_B_Gpq1DOjM2_2;
	wire w_dff_B_yDwcpi3L2_1;
	wire w_dff_B_O7eGrU9d5_2;
	wire w_dff_B_FCYgnG4M9_2;
	wire w_dff_B_HmrHlPGp3_2;
	wire w_dff_B_IJqciMO44_2;
	wire w_dff_B_F47BQwFu2_2;
	wire w_dff_B_22mCeoIk7_2;
	wire w_dff_B_va4zvVCo2_2;
	wire w_dff_B_x8aip9lM7_2;
	wire w_dff_B_rdkqiocP9_2;
	wire w_dff_B_ewWnwWek2_2;
	wire w_dff_B_Vv4HgKB73_1;
	wire w_dff_B_VYxybrD26_2;
	wire w_dff_B_5ZipRCYh4_2;
	wire w_dff_B_E1fKmDBK1_2;
	wire w_dff_B_Q8I7aWfH8_2;
	wire w_dff_B_itzwMyMP3_2;
	wire w_dff_B_7vfeekxt9_2;
	wire w_dff_B_gdRa8BAw4_2;
	wire w_dff_B_n7O6EScb1_2;
	wire w_dff_B_aRfMzHED9_1;
	wire w_dff_B_u6LFQJzG1_2;
	wire w_dff_B_pkp0MDj07_2;
	wire w_dff_B_Qo2Z6x0A8_2;
	wire w_dff_B_OLdugPB46_2;
	wire w_dff_B_3y1bZXqQ4_2;
	wire w_dff_B_TQjrYt633_2;
	wire w_dff_B_TCPyOj6B9_2;
	wire w_dff_B_lXlV1jzs3_1;
	wire w_dff_B_uPKK8ESG8_0;
	wire w_dff_B_NenG3xHE2_2;
	wire w_dff_B_hBRVaz9W2_2;
	wire w_dff_B_PZOVoV967_2;
	wire w_dff_B_iAZ0Lkdv4_1;
	wire w_dff_B_csL5jpSV9_1;
	wire w_dff_A_9f3FoyNE9_0;
	wire w_dff_A_WYSV1EYY1_0;
	wire w_dff_A_89r2owrF7_0;
	wire w_dff_A_bs6TpDgl8_1;
	wire w_dff_B_2c2Vq3eT1_2;
	wire w_dff_B_TJfsuamC7_2;
	wire w_dff_B_c0gKDITm0_1;
	wire w_dff_B_0Kt4G5Mp8_2;
	wire w_dff_B_seHp4O5c8_2;
	wire w_dff_B_xVWXescX2_2;
	wire w_dff_B_WK1KZI2k5_2;
	wire w_dff_B_NTSDQlkA8_2;
	wire w_dff_B_JeYbGqYJ3_2;
	wire w_dff_B_gII3xVBw6_2;
	wire w_dff_B_nYqfiiSP0_2;
	wire w_dff_B_KcmjyqDt9_2;
	wire w_dff_B_xPtwnFHQ8_2;
	wire w_dff_B_10X5kgUQ6_2;
	wire w_dff_B_JTzkY5tB8_2;
	wire w_dff_B_JRa8KJyg3_2;
	wire w_dff_B_2YUPKL386_2;
	wire w_dff_B_FEcWnkgH6_2;
	wire w_dff_B_E4MhIlBi4_2;
	wire w_dff_B_WxxUFk6Y8_2;
	wire w_dff_B_AzEzZdB57_2;
	wire w_dff_B_SajIirry9_2;
	wire w_dff_B_VOyzUhNY4_2;
	wire w_dff_B_E296GWDi4_2;
	wire w_dff_B_9dSD4YXs7_2;
	wire w_dff_B_2dxaVkZi9_2;
	wire w_dff_B_8zqNlNcM7_2;
	wire w_dff_B_ZGfGp6El6_2;
	wire w_dff_B_0bXkMjxX5_2;
	wire w_dff_B_Zr5J63or4_2;
	wire w_dff_B_Mn77ED753_2;
	wire w_dff_B_s20hIMS20_2;
	wire w_dff_B_0WtfogX21_2;
	wire w_dff_B_yP1yH5Mq7_2;
	wire w_dff_B_Wi9A6BGr9_2;
	wire w_dff_B_rMaPfSgc1_2;
	wire w_dff_B_NPdh8szz8_2;
	wire w_dff_B_4WINysLX4_2;
	wire w_dff_B_L9bSzvvj0_2;
	wire w_dff_B_ZuB48PZT2_1;
	wire w_dff_A_1gzZBzEp4_1;
	wire w_dff_B_PgiGbC5X8_1;
	wire w_dff_B_mxJtfWY44_2;
	wire w_dff_B_Sc34o0UJ5_2;
	wire w_dff_B_ra8v41Jb7_2;
	wire w_dff_B_9C6VkztW6_2;
	wire w_dff_B_wGCewpp48_2;
	wire w_dff_B_ZUiWFomF2_2;
	wire w_dff_B_iZjeqE6k9_2;
	wire w_dff_B_7u8kzptq9_2;
	wire w_dff_B_s4PXG8wY4_2;
	wire w_dff_B_UCp7faNg3_2;
	wire w_dff_B_Flm8jeW13_2;
	wire w_dff_B_gNCv9Isw2_2;
	wire w_dff_B_l2MS1AxN4_2;
	wire w_dff_B_wy9gGi1J2_2;
	wire w_dff_B_MIvxTpkS4_2;
	wire w_dff_B_y2qnU9p77_2;
	wire w_dff_B_ONpLwPjA6_2;
	wire w_dff_B_ixQXjcEW6_2;
	wire w_dff_B_yReINQyO8_2;
	wire w_dff_B_6gwlQc8T7_2;
	wire w_dff_B_qP3ZeTuv7_2;
	wire w_dff_B_AWwznU641_2;
	wire w_dff_B_HFhs9QCc4_2;
	wire w_dff_B_6GAkWeor2_2;
	wire w_dff_B_szGhqEO27_2;
	wire w_dff_B_VnwQJJHW4_2;
	wire w_dff_B_Yyt009D82_2;
	wire w_dff_B_u4StBFgl2_2;
	wire w_dff_B_qY5CoyaW7_2;
	wire w_dff_B_5XkrnHgD9_2;
	wire w_dff_B_IQs7OLLp0_2;
	wire w_dff_B_UP6lgHQk0_2;
	wire w_dff_B_Jm9tIshv4_1;
	wire w_dff_B_cDeRRrvT6_2;
	wire w_dff_B_beFV1w8m4_2;
	wire w_dff_B_jDNMgaUX7_2;
	wire w_dff_B_QA2I0oNs9_2;
	wire w_dff_B_3v3pc9j28_2;
	wire w_dff_B_luIh8VKD0_2;
	wire w_dff_B_WxNTYIEB8_2;
	wire w_dff_B_Qj1EpNWE3_2;
	wire w_dff_B_ZDD1f9eW5_2;
	wire w_dff_B_NlsUxI5B0_2;
	wire w_dff_B_nqMpzWkn8_2;
	wire w_dff_B_f8ji0yuA5_2;
	wire w_dff_B_8hoDUfZT0_2;
	wire w_dff_B_29rJ4ON59_2;
	wire w_dff_B_hr2CLswT9_2;
	wire w_dff_B_mYk1Dwt93_2;
	wire w_dff_B_VeL6enjW6_2;
	wire w_dff_B_ImBfs6A44_2;
	wire w_dff_B_g1M8Pnz44_2;
	wire w_dff_B_oAJ0WtWL1_2;
	wire w_dff_B_Wk6iza651_2;
	wire w_dff_B_HWLxt7d93_2;
	wire w_dff_B_6gzuIKjc0_2;
	wire w_dff_B_ruKjRQyW3_2;
	wire w_dff_B_kiwq5H8R5_2;
	wire w_dff_B_RSneklzm8_2;
	wire w_dff_B_PIQ4bFKM0_2;
	wire w_dff_B_0gddxcGe8_2;
	wire w_dff_B_NZTEQUB73_2;
	wire w_dff_B_YVApPPrf4_1;
	wire w_dff_B_u9c3TRX55_2;
	wire w_dff_B_x7z4HUUf8_2;
	wire w_dff_B_PHOpvzVV7_2;
	wire w_dff_B_BtrFSV5h5_2;
	wire w_dff_B_cMnJIbxr2_2;
	wire w_dff_B_vtyohZyJ7_2;
	wire w_dff_B_Xn3H3yZb6_2;
	wire w_dff_B_lU3I9ZbZ9_2;
	wire w_dff_B_A0LUHoC71_2;
	wire w_dff_B_YIAtZzM50_2;
	wire w_dff_B_VnqxHIum3_2;
	wire w_dff_B_oFXFmMYU7_2;
	wire w_dff_B_oh906Dl82_2;
	wire w_dff_B_hG0zkLKC8_2;
	wire w_dff_B_1Ws0COUy6_2;
	wire w_dff_B_9UBkVgE06_2;
	wire w_dff_B_e9cYIyqH7_2;
	wire w_dff_B_iJOGgfpt3_2;
	wire w_dff_B_6JW7yPFx5_2;
	wire w_dff_B_fXXlRTTR1_2;
	wire w_dff_B_1nQQUPSi4_2;
	wire w_dff_B_GGatLbCo3_2;
	wire w_dff_B_on73QUej8_2;
	wire w_dff_B_fXaeBC208_2;
	wire w_dff_B_3wbRcmS09_2;
	wire w_dff_B_ifC4YSHr9_2;
	wire w_dff_B_V46Xsi6b9_1;
	wire w_dff_B_hjCW9IC32_2;
	wire w_dff_B_sjol2ITj3_2;
	wire w_dff_B_5LxvmuZQ6_2;
	wire w_dff_B_Vtq2Wt5F8_2;
	wire w_dff_B_lJPvG3pD4_2;
	wire w_dff_B_PHTJ7ki73_2;
	wire w_dff_B_g98Uk9ux8_2;
	wire w_dff_B_pu99VB340_2;
	wire w_dff_B_kvl75geT2_2;
	wire w_dff_B_JxDq53FH1_2;
	wire w_dff_B_N4LiO5Lb4_2;
	wire w_dff_B_wTHAbH3L8_2;
	wire w_dff_B_PS2vrbAn7_2;
	wire w_dff_B_kV5qJHLH8_2;
	wire w_dff_B_IBjgHtyl9_2;
	wire w_dff_B_Yyw7O13w6_2;
	wire w_dff_B_shTCMpjF3_2;
	wire w_dff_B_nQFoaHz82_2;
	wire w_dff_B_SY5ktz1Q7_2;
	wire w_dff_B_wi7OBm364_2;
	wire w_dff_B_6qdMvcAC0_2;
	wire w_dff_B_DHkkivkZ8_2;
	wire w_dff_B_3TmBEJSr7_1;
	wire w_dff_B_A06MPEgt5_2;
	wire w_dff_B_YROz2R6i2_2;
	wire w_dff_B_tl21GLti4_2;
	wire w_dff_B_zlQkHDtW8_2;
	wire w_dff_B_xbw2aLdN8_2;
	wire w_dff_B_vR4YPr1b0_2;
	wire w_dff_B_EHT8PmzI8_2;
	wire w_dff_B_grUEZkXN1_2;
	wire w_dff_B_lf9HrfCw9_2;
	wire w_dff_B_JQ958yAm5_2;
	wire w_dff_B_PaCN99jw2_2;
	wire w_dff_B_s8jj7hbg9_2;
	wire w_dff_B_QTB9aI7J6_2;
	wire w_dff_B_M7kcno959_2;
	wire w_dff_B_a5GDJgSa4_2;
	wire w_dff_B_kVp31UCR9_2;
	wire w_dff_B_34QrVnqd4_2;
	wire w_dff_B_xZy6sAe14_2;
	wire w_dff_B_kdYGzVW45_2;
	wire w_dff_B_i3mTkYqK7_2;
	wire w_dff_B_4KcQbGzm1_1;
	wire w_dff_B_zIrAZKW33_2;
	wire w_dff_B_JPUDhBHX4_2;
	wire w_dff_B_DQ822bHd0_2;
	wire w_dff_B_GHKp6BXn5_2;
	wire w_dff_B_4wBaTMAy5_2;
	wire w_dff_B_GMCQL4WO8_2;
	wire w_dff_B_bPkKppGB2_2;
	wire w_dff_B_P3rlvkXe6_2;
	wire w_dff_B_qCujv8D04_2;
	wire w_dff_B_M3Fmb5Ys5_2;
	wire w_dff_B_XnKRtw8C6_2;
	wire w_dff_B_yHYHCaxJ8_2;
	wire w_dff_B_rNKyEzJP1_2;
	wire w_dff_B_zjjrUoGh4_2;
	wire w_dff_B_PNJ5fSUm2_2;
	wire w_dff_B_4fxM2bAj6_2;
	wire w_dff_B_OZfAXnUQ6_2;
	wire w_dff_B_tWkl39uc5_2;
	wire w_dff_B_AVYQgcJo9_1;
	wire w_dff_B_FCfwY96i0_2;
	wire w_dff_B_k2grJYnE4_2;
	wire w_dff_B_sCvb2oUk8_2;
	wire w_dff_B_z7aJZkI97_2;
	wire w_dff_B_tMEmoz6P1_2;
	wire w_dff_B_LlS9wLXh2_2;
	wire w_dff_B_slm2WGys1_2;
	wire w_dff_B_9e85SUql4_2;
	wire w_dff_B_VgODNAGO3_2;
	wire w_dff_B_MpOvCXKS5_2;
	wire w_dff_B_MkymvTnz7_2;
	wire w_dff_B_YjBIlWd48_2;
	wire w_dff_B_WURChH2z1_2;
	wire w_dff_B_nEEra4m92_2;
	wire w_dff_B_0PjRQSM98_2;
	wire w_dff_B_wrtKf0bo3_2;
	wire w_dff_B_qIP4ZgBY5_1;
	wire w_dff_B_ZVvaXVXz7_2;
	wire w_dff_B_W9ZGgO086_2;
	wire w_dff_B_Jr55POId3_2;
	wire w_dff_B_GfCCucKV8_2;
	wire w_dff_B_8GYsv1kC8_2;
	wire w_dff_B_RmaF4cQG2_2;
	wire w_dff_B_I8CXgn2L7_2;
	wire w_dff_B_XaU6V0Ck5_2;
	wire w_dff_B_3S4Kr9Iw2_2;
	wire w_dff_B_kdQc0vX30_2;
	wire w_dff_B_BbPEeNoj1_2;
	wire w_dff_B_tyw3JFfG4_2;
	wire w_dff_B_b5PoWetD6_2;
	wire w_dff_B_YeAMfOBG9_2;
	wire w_dff_B_Cn4ggaBf8_1;
	wire w_dff_B_IneA9yhg0_2;
	wire w_dff_B_sSHGSfMz1_2;
	wire w_dff_B_kFpYbUMO4_2;
	wire w_dff_B_tQsDpTIQ5_2;
	wire w_dff_B_dVGs5xcI9_2;
	wire w_dff_B_isn4nnSQ6_2;
	wire w_dff_B_1WHfJ1Hh1_2;
	wire w_dff_B_RvRI9bDG8_2;
	wire w_dff_B_Y37IMIYK6_2;
	wire w_dff_B_dfDpnIzb4_2;
	wire w_dff_B_ijB8H5kj6_2;
	wire w_dff_B_iyTxPbzz4_2;
	wire w_dff_B_Bj9aSqi12_1;
	wire w_dff_B_6jOT558k5_2;
	wire w_dff_B_a3kqAr9B3_2;
	wire w_dff_B_ZY9Ygz6Y6_2;
	wire w_dff_B_kgEVeQD81_2;
	wire w_dff_B_WWI3SvlO4_2;
	wire w_dff_B_5Nc4NQKD6_2;
	wire w_dff_B_9HaZCoiB2_2;
	wire w_dff_B_1OHFcMK08_2;
	wire w_dff_B_V6Ai4syZ5_2;
	wire w_dff_B_EA0egYHr7_2;
	wire w_dff_B_e5zG3G192_1;
	wire w_dff_B_hHF4PLv98_2;
	wire w_dff_B_vKloUbis9_2;
	wire w_dff_B_yUfKHhCJ3_2;
	wire w_dff_B_Jt8mYg262_2;
	wire w_dff_B_0rTavOea3_2;
	wire w_dff_B_J5a6kTfg1_2;
	wire w_dff_B_CyeZAuXr7_2;
	wire w_dff_B_5ER2SwBJ6_2;
	wire w_dff_B_uosZhQmA9_1;
	wire w_dff_B_fdLzkwVB3_2;
	wire w_dff_B_n7DB7ScB4_2;
	wire w_dff_B_u7KsKqec9_2;
	wire w_dff_B_b02pt5Jq6_2;
	wire w_dff_B_2xUaqW1E6_2;
	wire w_dff_B_iy6eoe9I4_2;
	wire w_dff_B_WS4OrXGn4_1;
	wire w_dff_B_y6wDHljS6_1;
	wire w_dff_B_w6gx9XeJ2_2;
	wire w_dff_B_NoHTSPrv1_2;
	wire w_dff_B_YpiywRqR1_2;
	wire w_dff_B_VKVv2ZlL7_2;
	wire w_dff_A_sffExBlQ5_1;
	wire w_dff_B_QaA4BnNI5_1;
	wire w_dff_B_nNWTPtOn8_1;
	wire w_dff_A_lTu2GWwo3_1;
	wire w_dff_A_q2YgquF76_2;
	wire w_dff_A_jkneepKI9_2;
	wire w_dff_B_kI2ENWMc5_2;
	wire w_dff_B_QXDLZGjL9_2;
	wire w_dff_B_Wc61OfOK0_1;
	wire w_dff_B_K06jwAoZ4_2;
	wire w_dff_B_jElGjNCa7_2;
	wire w_dff_B_7d8eh8lw1_2;
	wire w_dff_B_dQEkcGzT0_2;
	wire w_dff_B_sHnnsn2q7_2;
	wire w_dff_B_f2o4nSvx7_2;
	wire w_dff_B_PQGJr6EU5_2;
	wire w_dff_B_qU5riOqO4_2;
	wire w_dff_B_tyfWo8yg3_2;
	wire w_dff_B_ivJ0EobA9_2;
	wire w_dff_B_FwGifej58_2;
	wire w_dff_B_loPUOzs56_2;
	wire w_dff_B_uaAIJsIE8_2;
	wire w_dff_B_Sdx0dtdJ1_2;
	wire w_dff_B_iepCSMSW9_2;
	wire w_dff_B_fTTMvD3V9_2;
	wire w_dff_B_zdb5BAwl6_2;
	wire w_dff_B_4G62qj6k2_2;
	wire w_dff_B_Rj2vvGED0_2;
	wire w_dff_B_ngggpycu0_2;
	wire w_dff_B_Hg5LHLr43_2;
	wire w_dff_B_0299Flaz5_2;
	wire w_dff_B_o5AnkwZD8_2;
	wire w_dff_B_JPxaRGMO5_2;
	wire w_dff_B_d1YXzBx40_2;
	wire w_dff_B_qcX1VLLs6_2;
	wire w_dff_B_1zQJcAhG4_2;
	wire w_dff_B_33RengTd9_2;
	wire w_dff_B_gbkHGl7v0_2;
	wire w_dff_B_aYTb8ZT22_2;
	wire w_dff_B_iB0L1D0K5_2;
	wire w_dff_B_fvWhLSL56_2;
	wire w_dff_B_UMCpyrhA1_2;
	wire w_dff_B_DQUrikwz3_2;
	wire w_dff_B_PBkw2l3d5_2;
	wire w_dff_B_1m2STfot5_2;
	wire w_dff_B_MO3xkrHL2_2;
	wire w_dff_B_5MuID1Q30_1;
	wire w_dff_A_km6ZBDLX1_1;
	wire w_dff_B_Jch7zrMC4_1;
	wire w_dff_B_EE2ppDoD8_2;
	wire w_dff_B_LwLvKN2Y4_2;
	wire w_dff_B_3OTw13iF9_2;
	wire w_dff_B_ZclvFa4K6_2;
	wire w_dff_B_CVlt1Gry9_2;
	wire w_dff_B_69I4gQ4O2_2;
	wire w_dff_B_9nES55Xl7_2;
	wire w_dff_B_CHzIh5Jl3_2;
	wire w_dff_B_onC38s4b0_2;
	wire w_dff_B_EFiOk7zX8_2;
	wire w_dff_B_NDXDpqvm9_2;
	wire w_dff_B_VisgXv3B3_2;
	wire w_dff_B_HSC6F05V8_2;
	wire w_dff_B_D6VgF25T1_2;
	wire w_dff_B_aHyL4SUc6_2;
	wire w_dff_B_tI5ARTMl5_2;
	wire w_dff_B_5dlPVokj1_2;
	wire w_dff_B_YlMp9Zff7_2;
	wire w_dff_B_KHa3WL0A6_2;
	wire w_dff_B_hnyuUPKr5_2;
	wire w_dff_B_qWAbQCi56_2;
	wire w_dff_B_C8A15Wz96_2;
	wire w_dff_B_cpMeQEWp9_2;
	wire w_dff_B_DN7WeaL16_2;
	wire w_dff_B_9nIFu5I88_2;
	wire w_dff_B_zR0bJ7Qn3_2;
	wire w_dff_B_rsibzmaI4_2;
	wire w_dff_B_wo4XRTlx0_2;
	wire w_dff_B_xh8Ntsfk2_2;
	wire w_dff_B_W1eUP5YR8_2;
	wire w_dff_B_DKzJq4jk9_2;
	wire w_dff_B_kiAL6Qoz4_2;
	wire w_dff_B_hARVlZ0U7_2;
	wire w_dff_B_ivnOAsjy4_1;
	wire w_dff_B_LXVEP8uZ8_2;
	wire w_dff_B_4poR2CQm4_2;
	wire w_dff_B_mgOadkX03_2;
	wire w_dff_B_mgD8YAwU6_2;
	wire w_dff_B_Hdhj5BRk0_2;
	wire w_dff_B_mgW6aHdy9_2;
	wire w_dff_B_0C8RqJtJ9_2;
	wire w_dff_B_sdU84hag3_2;
	wire w_dff_B_5w8UROTJ8_2;
	wire w_dff_B_qidCpLAl7_2;
	wire w_dff_B_qwggIlGA0_2;
	wire w_dff_B_xGWCQptL5_2;
	wire w_dff_B_T0fvdXNe4_2;
	wire w_dff_B_CQLgawAo8_2;
	wire w_dff_B_HGMviyr69_2;
	wire w_dff_B_R2fiFvk72_2;
	wire w_dff_B_7a1bvLkJ6_2;
	wire w_dff_B_QMZZNcah3_2;
	wire w_dff_B_krobLoUg5_2;
	wire w_dff_B_CJxFDmu99_2;
	wire w_dff_B_Nm3JpYMv5_2;
	wire w_dff_B_rMvCm0j85_2;
	wire w_dff_B_8BFoXhsj4_2;
	wire w_dff_B_USsMmGwY4_2;
	wire w_dff_B_nIBugPL99_2;
	wire w_dff_B_wdpfAOTz2_2;
	wire w_dff_B_rBZiQDny7_2;
	wire w_dff_B_FkWhASko7_2;
	wire w_dff_B_VQgZ5SR97_2;
	wire w_dff_B_r9HkWtyQ6_2;
	wire w_dff_B_cvqoWs9e8_1;
	wire w_dff_B_FST0Ilhu0_2;
	wire w_dff_B_LsqPvrrA9_2;
	wire w_dff_B_G8WZ7BDo4_2;
	wire w_dff_B_OrqsD9Fv0_2;
	wire w_dff_B_tUHSKBNG1_2;
	wire w_dff_B_opsqlyLX3_2;
	wire w_dff_B_poDfQ2nZ2_2;
	wire w_dff_B_cOH5N3YD1_2;
	wire w_dff_B_DGMxRnhr3_2;
	wire w_dff_B_cBoDgnvL0_2;
	wire w_dff_B_nzuSHpu41_2;
	wire w_dff_B_jz5wnW713_2;
	wire w_dff_B_eTYVcJPw7_2;
	wire w_dff_B_R5c1PYkn6_2;
	wire w_dff_B_xlhFY48i7_2;
	wire w_dff_B_SJEh11Qb7_2;
	wire w_dff_B_J3K6ptWE5_2;
	wire w_dff_B_qm05tenc4_2;
	wire w_dff_B_hZB5OZ4t3_2;
	wire w_dff_B_9f49ZbKq8_2;
	wire w_dff_B_wf7cz2mD1_2;
	wire w_dff_B_zS1qtQ2l2_2;
	wire w_dff_B_OKJdbkSh3_2;
	wire w_dff_B_64zbX8iC4_2;
	wire w_dff_B_A7bc56LV9_2;
	wire w_dff_B_BeKR35A02_2;
	wire w_dff_B_xl0I0JEE5_2;
	wire w_dff_B_ELpE24bH9_1;
	wire w_dff_B_1GBAdd8W1_2;
	wire w_dff_B_QbLr8CWZ7_2;
	wire w_dff_B_JSMVuqLd7_2;
	wire w_dff_B_dMOPpgOq5_2;
	wire w_dff_B_dGfTqZLC9_2;
	wire w_dff_B_LfOXdbJe2_2;
	wire w_dff_B_S6w4rrd83_2;
	wire w_dff_B_oqevpRA25_2;
	wire w_dff_B_S6dsqgZo0_2;
	wire w_dff_B_rk6T9Vx62_2;
	wire w_dff_B_woIeXbvP3_2;
	wire w_dff_B_YXFIYIiR5_2;
	wire w_dff_B_DaPraFpZ2_2;
	wire w_dff_B_M8I1E7Xv0_2;
	wire w_dff_B_QBZIqR743_2;
	wire w_dff_B_fq7qfXWc3_2;
	wire w_dff_B_b7YJJ5Yc3_2;
	wire w_dff_B_vYV35fv94_2;
	wire w_dff_B_nzpouyKv1_2;
	wire w_dff_B_yvxZHNbN7_2;
	wire w_dff_B_2mTGSGRM8_2;
	wire w_dff_B_mg7ZoLSc5_2;
	wire w_dff_B_gIN7GL8I4_2;
	wire w_dff_B_Vk4Qj9aA2_2;
	wire w_dff_B_Usg5uhqf5_1;
	wire w_dff_B_2TfIy28O0_2;
	wire w_dff_B_OX9k87qZ1_2;
	wire w_dff_B_VpDadZwI1_2;
	wire w_dff_B_IyhPZD3n2_2;
	wire w_dff_B_1i99748o7_2;
	wire w_dff_B_Qz2hYg2v7_2;
	wire w_dff_B_4SFflszo3_2;
	wire w_dff_B_bYqvUog75_2;
	wire w_dff_B_Xcae1ElU8_2;
	wire w_dff_B_yr7H8RoG8_2;
	wire w_dff_B_dqaXI5Q01_2;
	wire w_dff_B_PoKKm8Ac3_2;
	wire w_dff_B_ehinX51G4_2;
	wire w_dff_B_BirjClnD4_2;
	wire w_dff_B_3WQ4HrMA0_2;
	wire w_dff_B_g5C6IMhb1_2;
	wire w_dff_B_y8C8BSDi7_2;
	wire w_dff_B_gtSv2GW19_2;
	wire w_dff_B_Rg2LZjCX6_2;
	wire w_dff_B_6TEB4FEv0_2;
	wire w_dff_B_KUz0OnNt7_1;
	wire w_dff_B_zYx6m8hr6_2;
	wire w_dff_B_KJ45VJJk2_2;
	wire w_dff_B_rMd0fbo21_2;
	wire w_dff_B_hTmj3hb72_2;
	wire w_dff_B_amRdSPst1_2;
	wire w_dff_B_PngaMlZc3_2;
	wire w_dff_B_m9iKnzeW7_2;
	wire w_dff_B_8wm29cfb6_2;
	wire w_dff_B_9A9bssQh9_2;
	wire w_dff_B_elLOdBSp8_2;
	wire w_dff_B_Ir5SK7Ew5_2;
	wire w_dff_B_UKXmqFIy2_2;
	wire w_dff_B_xwBRuEfy2_2;
	wire w_dff_B_BvPfyuBF3_2;
	wire w_dff_B_W5BkA0uv6_2;
	wire w_dff_B_GH7L05Zu3_2;
	wire w_dff_B_mHCpiLTu7_2;
	wire w_dff_B_BMw3Lxb49_2;
	wire w_dff_B_v6EO7e6d1_1;
	wire w_dff_B_7K2fZRS23_2;
	wire w_dff_B_6j2iQjyc0_2;
	wire w_dff_B_f2b3cNxg9_2;
	wire w_dff_B_4F8rAj4L9_2;
	wire w_dff_B_fr6qZNO09_2;
	wire w_dff_B_NHqH9jy45_2;
	wire w_dff_B_OOltNCmH7_2;
	wire w_dff_B_9sGK2Dko4_2;
	wire w_dff_B_QUELZei44_2;
	wire w_dff_B_9h4a05Wh0_2;
	wire w_dff_B_jdh6OKW50_2;
	wire w_dff_B_B8W2kcWb2_2;
	wire w_dff_B_MEA3lOOF7_2;
	wire w_dff_B_k2xht5bT4_2;
	wire w_dff_B_7TOama1m4_2;
	wire w_dff_B_531w516D6_2;
	wire w_dff_B_g8b86Sln6_1;
	wire w_dff_B_CX7Ltmiv3_2;
	wire w_dff_B_tYpSwzCP7_2;
	wire w_dff_B_kSltH5U88_2;
	wire w_dff_B_mDl3wRKA0_2;
	wire w_dff_B_wD5QUVQy1_2;
	wire w_dff_B_M3glYfEu9_2;
	wire w_dff_B_yARmHfY21_2;
	wire w_dff_B_FKyAMUxU3_2;
	wire w_dff_B_4mxO6BWl3_2;
	wire w_dff_B_OyqZG4w32_2;
	wire w_dff_B_FtxjEmG28_2;
	wire w_dff_B_s2PqJ7iJ2_2;
	wire w_dff_B_A6yDWUB58_2;
	wire w_dff_B_fyCeKIlH9_2;
	wire w_dff_B_sqlWpZ4B1_1;
	wire w_dff_B_ZtSnJRsu1_2;
	wire w_dff_B_TkVc8CnX4_2;
	wire w_dff_B_0dQqA2ul3_2;
	wire w_dff_B_U00cK3hr9_2;
	wire w_dff_B_Ar4dDLoa9_2;
	wire w_dff_B_68Tvh88u8_2;
	wire w_dff_B_mgjrZIJX6_2;
	wire w_dff_B_NSlQta5W2_2;
	wire w_dff_B_DARwgzxd6_2;
	wire w_dff_B_F2GJ0d8h3_2;
	wire w_dff_B_CPUjbOtW5_2;
	wire w_dff_B_CmZh1vkp5_2;
	wire w_dff_B_QPvjEvrN3_1;
	wire w_dff_B_yEoth6aF6_2;
	wire w_dff_B_giZl3HEc0_2;
	wire w_dff_B_OhjmHqlE3_2;
	wire w_dff_B_Ih6yjIAI0_2;
	wire w_dff_B_q63G9MCO6_2;
	wire w_dff_B_u15dV6Ig2_2;
	wire w_dff_B_d7wDfoEm9_2;
	wire w_dff_B_4bXUAm0L9_2;
	wire w_dff_B_tXKvlKa61_2;
	wire w_dff_B_lKp0G3Gz6_2;
	wire w_dff_B_dl8ogSlE8_1;
	wire w_dff_B_Brc56l3K1_2;
	wire w_dff_B_v1pP1J3C1_2;
	wire w_dff_B_J7OPjAy74_2;
	wire w_dff_B_6z5U1c8C8_2;
	wire w_dff_B_QNofcxy58_2;
	wire w_dff_B_s9SmGu9L0_2;
	wire w_dff_B_9oCeouqO9_2;
	wire w_dff_B_4f0QssU07_2;
	wire w_dff_B_jVyz4aVK1_1;
	wire w_dff_B_ZpSHMSn91_2;
	wire w_dff_B_2juTzK0k2_2;
	wire w_dff_B_jeIukxcj2_2;
	wire w_dff_B_J22aLDwg1_2;
	wire w_dff_B_TQ2jbAwY4_2;
	wire w_dff_B_2O4uTLYz9_2;
	wire w_dff_B_xZpEN1Py9_2;
	wire w_dff_B_rYc5JrPE1_1;
	wire w_dff_B_YdACboNw3_1;
	wire w_dff_B_A58hShCc8_2;
	wire w_dff_B_pAXqnY8h2_2;
	wire w_dff_B_s4uNUbwG5_2;
	wire w_dff_B_dnWkgseM9_2;
	wire w_dff_A_VcZH5Esl6_1;
	wire w_dff_B_e9Y6sfxe4_1;
	wire w_dff_B_1qBU2jhh6_1;
	wire w_dff_A_skMxtdkH5_0;
	wire w_dff_A_sg2BvyBK1_1;
	wire w_dff_A_8wznEIJ80_1;
	wire w_dff_B_DExLKsan5_2;
	wire w_dff_B_pZiXbu383_2;
	wire w_dff_B_Ha4dA8CP6_1;
	wire w_dff_B_MK926buB6_2;
	wire w_dff_B_R6zuIxg68_2;
	wire w_dff_B_xZphkrM66_2;
	wire w_dff_B_QexdX6tn6_2;
	wire w_dff_B_5OhqglfR9_2;
	wire w_dff_B_FSbp1kdf4_2;
	wire w_dff_B_dDVTMdod0_2;
	wire w_dff_B_L5UijDuh4_2;
	wire w_dff_B_ej23yrYe6_2;
	wire w_dff_B_KfLyFKoX3_2;
	wire w_dff_B_EHuwfCyy0_2;
	wire w_dff_B_TiUYpoOm2_2;
	wire w_dff_B_sbjeyHi95_2;
	wire w_dff_B_9x7PCOJT1_2;
	wire w_dff_B_WRrAVpjx7_2;
	wire w_dff_B_FpsIhPoJ8_2;
	wire w_dff_B_Eciu9rSA7_2;
	wire w_dff_B_JDcuNnem2_2;
	wire w_dff_B_GfA48xs63_2;
	wire w_dff_B_dGjPk2uv4_2;
	wire w_dff_B_8ar8sJEJ5_2;
	wire w_dff_B_Tx2FWoGG4_2;
	wire w_dff_B_BGoplHs33_2;
	wire w_dff_B_G263SDlw2_2;
	wire w_dff_B_Ftj0OEKZ3_2;
	wire w_dff_B_0m1MsdC36_2;
	wire w_dff_B_n3pEO8v07_2;
	wire w_dff_B_nJVjp2zy9_2;
	wire w_dff_B_pFTCa8SU0_2;
	wire w_dff_B_x4F5fb0j9_2;
	wire w_dff_B_GN775u902_2;
	wire w_dff_B_kbZdJDio6_2;
	wire w_dff_B_xXRxls5d9_2;
	wire w_dff_B_LFHM66KT6_2;
	wire w_dff_B_YvgYwXpD7_2;
	wire w_dff_B_BLKrYaMk7_2;
	wire w_dff_B_8MAZy0s30_2;
	wire w_dff_B_GjvakE6n3_2;
	wire w_dff_B_d35o9utC8_1;
	wire w_dff_A_lLOzs8437_1;
	wire w_dff_B_mFNHx6He1_1;
	wire w_dff_B_M6OkMOFi3_2;
	wire w_dff_B_Lk0Ern2v1_2;
	wire w_dff_B_l7GvpiWy7_2;
	wire w_dff_B_zCWGqkxA6_2;
	wire w_dff_B_wxPiLBOk4_2;
	wire w_dff_B_RUmcQ1o01_2;
	wire w_dff_B_0uzAax8D3_2;
	wire w_dff_B_DFTkswCf8_2;
	wire w_dff_B_tWpstZeL1_2;
	wire w_dff_B_lYvgkDur0_2;
	wire w_dff_B_oSR7azdG1_2;
	wire w_dff_B_cJaitoE09_2;
	wire w_dff_B_4cDCKpr24_2;
	wire w_dff_B_mzH3WjKv8_2;
	wire w_dff_B_mqHUsab91_2;
	wire w_dff_B_4Q4iHfYy6_2;
	wire w_dff_B_89uiv0Ei0_2;
	wire w_dff_B_x2PUERo15_2;
	wire w_dff_B_NyftFSa39_2;
	wire w_dff_B_ROyZ1ODi7_2;
	wire w_dff_B_27uVoUy08_2;
	wire w_dff_B_iF0Q8r5y4_2;
	wire w_dff_B_0L4tKxqg7_2;
	wire w_dff_B_FRHv0RZz6_2;
	wire w_dff_B_YiHSCAt07_2;
	wire w_dff_B_H9ZunKdY0_2;
	wire w_dff_B_8vBf2JKc0_2;
	wire w_dff_B_F8ORJLhT7_2;
	wire w_dff_B_kyjDQxZT6_2;
	wire w_dff_B_JvFmRFZb9_2;
	wire w_dff_B_yp2Jug5Y8_2;
	wire w_dff_B_YviWvkZ03_2;
	wire w_dff_B_NOISaytV5_2;
	wire w_dff_B_6w8IAF025_2;
	wire w_dff_B_PkKGRpPN5_1;
	wire w_dff_B_PliDiHTF5_2;
	wire w_dff_B_kWXhzVmt0_2;
	wire w_dff_B_1fsV6qV82_2;
	wire w_dff_B_Ma50OG3U1_2;
	wire w_dff_B_Sljro1Zy7_2;
	wire w_dff_B_RwzDse3h8_2;
	wire w_dff_B_lroheoqH4_2;
	wire w_dff_B_M4Ftwh446_2;
	wire w_dff_B_3XmlgQfQ5_2;
	wire w_dff_B_59yEYbnS4_2;
	wire w_dff_B_JFJO1CNx0_2;
	wire w_dff_B_1Go9Z96e3_2;
	wire w_dff_B_zWv3JliJ1_2;
	wire w_dff_B_Xqv6Q7457_2;
	wire w_dff_B_4bcsZa5X9_2;
	wire w_dff_B_4fgELMmN9_2;
	wire w_dff_B_SPclwaLV7_2;
	wire w_dff_B_3Jqw9cmH6_2;
	wire w_dff_B_60k9XGYn7_2;
	wire w_dff_B_eXQKReoR1_2;
	wire w_dff_B_VCaaGmXz3_2;
	wire w_dff_B_QNeD0R4d5_2;
	wire w_dff_B_wMCwo19D5_2;
	wire w_dff_B_h6mzTWY73_2;
	wire w_dff_B_MGyxqxl27_2;
	wire w_dff_B_oUFAa6B86_2;
	wire w_dff_B_fLJ3mFif7_2;
	wire w_dff_B_SUlQUeiM2_2;
	wire w_dff_B_OR7k9PM48_2;
	wire w_dff_B_rsbKbUpA0_2;
	wire w_dff_B_chs9YUMz7_2;
	wire w_dff_B_y4LofFOP8_1;
	wire w_dff_B_E9L57k8p4_2;
	wire w_dff_B_h6VIM8T74_2;
	wire w_dff_B_YXnXG3sv8_2;
	wire w_dff_B_qn7w44uf3_2;
	wire w_dff_B_p70eb7q74_2;
	wire w_dff_B_tun9RBeK1_2;
	wire w_dff_B_l7Md8jEx6_2;
	wire w_dff_B_EzdPAXDg4_2;
	wire w_dff_B_cE7u32Im9_2;
	wire w_dff_B_fcCGa3yA4_2;
	wire w_dff_B_9TCNCdbG3_2;
	wire w_dff_B_9OIgVnGx2_2;
	wire w_dff_B_JEIUrNoe7_2;
	wire w_dff_B_AQxarMdi8_2;
	wire w_dff_B_p80LeQ700_2;
	wire w_dff_B_U1qPqupJ1_2;
	wire w_dff_B_NzaRCKDZ9_2;
	wire w_dff_B_F1NjqyrD3_2;
	wire w_dff_B_lhwUwXQC5_2;
	wire w_dff_B_9tzFCHfh5_2;
	wire w_dff_B_DZAcQQot6_2;
	wire w_dff_B_1ZlTv62G8_2;
	wire w_dff_B_oVmvi1404_2;
	wire w_dff_B_FdyllLGU0_2;
	wire w_dff_B_o7DYz6aA3_2;
	wire w_dff_B_D0WC8Jrt7_2;
	wire w_dff_B_RpWXsmZk5_2;
	wire w_dff_B_aDoAwMgG7_2;
	wire w_dff_B_ppPcRfFc9_1;
	wire w_dff_B_Ts4Q0cMs5_2;
	wire w_dff_B_meOfJaf41_2;
	wire w_dff_B_5a5NhNRy2_2;
	wire w_dff_B_TMshmf287_2;
	wire w_dff_B_uvL8JNmW4_2;
	wire w_dff_B_GhrSfGCU3_2;
	wire w_dff_B_whNCTC1c4_2;
	wire w_dff_B_M4fEIXqe1_2;
	wire w_dff_B_ojp2PRcz5_2;
	wire w_dff_B_4rW8kF436_2;
	wire w_dff_B_MrBC4i2M5_2;
	wire w_dff_B_V1HKmQ0i2_2;
	wire w_dff_B_JMJMF9Th4_2;
	wire w_dff_B_63l4kO8P4_2;
	wire w_dff_B_OySR4rAB3_2;
	wire w_dff_B_jtj6jdjk9_2;
	wire w_dff_B_y9yVm9JD1_2;
	wire w_dff_B_rqqcDBgj1_2;
	wire w_dff_B_PULExbZ77_2;
	wire w_dff_B_jXIKAYn04_2;
	wire w_dff_B_GflnDjUS4_2;
	wire w_dff_B_b5PExdQZ9_2;
	wire w_dff_B_qxazGri21_2;
	wire w_dff_B_mmbLPHoG8_2;
	wire w_dff_B_kZA6OXJq2_2;
	wire w_dff_B_m3XPCPsF9_1;
	wire w_dff_B_NE20FSM95_2;
	wire w_dff_B_9KkvwDLF1_2;
	wire w_dff_B_4KqldsYg2_2;
	wire w_dff_B_ABJrZuSc0_2;
	wire w_dff_B_69rUXBt77_2;
	wire w_dff_B_QUpLqKIj1_2;
	wire w_dff_B_Hw2y83XZ8_2;
	wire w_dff_B_Q1Y3gqzV8_2;
	wire w_dff_B_R9xoNTbM5_2;
	wire w_dff_B_297dIm7T1_2;
	wire w_dff_B_G8uTXr1V5_2;
	wire w_dff_B_hRDYlOWn6_2;
	wire w_dff_B_Lblrt5vK7_2;
	wire w_dff_B_AHGs0XeU3_2;
	wire w_dff_B_SmdO51gC2_2;
	wire w_dff_B_pRq4ur5N6_2;
	wire w_dff_B_nywyIp3O3_2;
	wire w_dff_B_dzeT7FWG9_2;
	wire w_dff_B_KZ5sjCly7_2;
	wire w_dff_B_wq8TGaBw9_2;
	wire w_dff_B_jLbPvk7S3_2;
	wire w_dff_B_PT0HtWut8_2;
	wire w_dff_B_LFD6220C1_1;
	wire w_dff_B_192RJ2D25_2;
	wire w_dff_B_6tC0R6bB8_2;
	wire w_dff_B_0m1TzszK9_2;
	wire w_dff_B_CGq9dzQb2_2;
	wire w_dff_B_lK6ncWOJ1_2;
	wire w_dff_B_Jj42eF2F1_2;
	wire w_dff_B_vUeD3pRe1_2;
	wire w_dff_B_zcD1WgtR7_2;
	wire w_dff_B_ql4sEzOF1_2;
	wire w_dff_B_QwxvYzoF6_2;
	wire w_dff_B_HB8TFIOu8_2;
	wire w_dff_B_9AmG9lX73_2;
	wire w_dff_B_2FUhEZFg2_2;
	wire w_dff_B_UpF9gtnx1_2;
	wire w_dff_B_UJjaStq72_2;
	wire w_dff_B_qr3wr1s50_2;
	wire w_dff_B_FQR6UAjT8_2;
	wire w_dff_B_yGnZ6wXe5_2;
	wire w_dff_B_yxOlFviZ9_1;
	wire w_dff_B_lTUeQ3Ie8_2;
	wire w_dff_B_SiLwA4z37_2;
	wire w_dff_B_Dbxf7ptV3_2;
	wire w_dff_B_MwkCO1nP0_2;
	wire w_dff_B_ADSSVMpC1_2;
	wire w_dff_B_kmmSPiV32_2;
	wire w_dff_B_LOAHBBye1_2;
	wire w_dff_B_I3HO192n8_2;
	wire w_dff_B_cFgzPVNV1_2;
	wire w_dff_B_mw6IXts98_2;
	wire w_dff_B_8lt01LFM9_2;
	wire w_dff_B_BsrgxrED6_2;
	wire w_dff_B_X65kA0ky4_2;
	wire w_dff_B_uvbGGtbD5_2;
	wire w_dff_B_W8bDkUIY1_2;
	wire w_dff_B_jPnbXJoN6_2;
	wire w_dff_B_YeF2aOoA8_1;
	wire w_dff_B_wubA050A5_2;
	wire w_dff_B_BWComL7u2_2;
	wire w_dff_B_a1EWwCsT7_2;
	wire w_dff_B_zziIjG450_2;
	wire w_dff_B_cLeb0gH46_2;
	wire w_dff_B_al7182yJ5_2;
	wire w_dff_B_cy3n8wFt3_2;
	wire w_dff_B_qcpxDavu7_2;
	wire w_dff_B_VEfHnmUB9_2;
	wire w_dff_B_Z7UGCT8t9_2;
	wire w_dff_B_9Ao9geGd2_2;
	wire w_dff_B_SxPerF1y7_2;
	wire w_dff_B_eC0l1LTS3_2;
	wire w_dff_B_1303sco78_2;
	wire w_dff_B_RZJNQvYs6_1;
	wire w_dff_B_5wOZZdvr8_2;
	wire w_dff_B_LRAwW28o0_2;
	wire w_dff_B_nwnijX4W2_2;
	wire w_dff_B_kSxzxN4e4_2;
	wire w_dff_B_VrSglJYH0_2;
	wire w_dff_B_B5J6Viwa8_2;
	wire w_dff_B_0iOOLS0p4_2;
	wire w_dff_B_Ra50P0mj4_2;
	wire w_dff_B_otY1Qg072_2;
	wire w_dff_B_lLJRwPWq6_2;
	wire w_dff_B_ix6HIcZB0_2;
	wire w_dff_B_1cZyvX0q5_2;
	wire w_dff_B_Y9rg3qgF9_1;
	wire w_dff_B_RSKJMgTC5_2;
	wire w_dff_B_SnpKHp4H3_2;
	wire w_dff_B_r1JyNFpg6_2;
	wire w_dff_B_16yNG7l58_2;
	wire w_dff_B_HpmQSZxj5_2;
	wire w_dff_B_5FkPQTEG1_2;
	wire w_dff_B_gsQZ6bPP0_2;
	wire w_dff_B_19w1q5RB4_2;
	wire w_dff_B_fAYXX5oW1_2;
	wire w_dff_B_W8fOQmi79_2;
	wire w_dff_B_bs4LziED4_1;
	wire w_dff_B_6p1u8bTu7_2;
	wire w_dff_B_2fcZf6734_2;
	wire w_dff_B_rXYW2y8B0_2;
	wire w_dff_B_GWLpQpMt3_2;
	wire w_dff_B_ew4zP9lJ7_2;
	wire w_dff_B_49XzoXZA7_2;
	wire w_dff_B_GI6vog5R5_2;
	wire w_dff_B_pxhg50Db2_2;
	wire w_dff_B_JGGGdc0n8_1;
	wire w_dff_B_zQNwH8Bu3_2;
	wire w_dff_B_3S6wzICb9_2;
	wire w_dff_B_3Iv169k68_2;
	wire w_dff_B_7y75TMyj1_2;
	wire w_dff_B_gSJHo93y5_2;
	wire w_dff_B_q6FLbAux0_2;
	wire w_dff_B_GAwbNi6N6_2;
	wire w_dff_B_EahjSriI7_1;
	wire w_dff_B_sUcNy1gV9_1;
	wire w_dff_B_UFFyI5mw4_1;
	wire w_dff_B_hbzpAAfY3_1;
	wire w_dff_B_5JXtGLp18_0;
	wire w_dff_A_6lXKfSQ66_0;
	wire w_dff_A_vJmeg3EW2_0;
	wire w_dff_B_8PB5xVkM2_1;
	wire w_dff_B_JAaSJxCS7_1;
	wire w_dff_A_0wMb0ngO3_0;
	wire w_dff_A_TKGC6uMf4_1;
	wire w_dff_A_mzOkYWKK3_1;
	wire w_dff_A_vMC9VBYo7_1;
	wire w_dff_A_RpSN5RcD5_1;
	wire w_dff_A_2HGbCkl93_1;
	wire w_dff_A_dfd1enHt4_1;
	wire w_dff_B_WzbyGmmA2_2;
	wire w_dff_B_Q6bCvniE8_2;
	wire w_dff_B_OXtOuo0n0_1;
	wire w_dff_B_VivaAZGf5_2;
	wire w_dff_B_dxhVN85L7_2;
	wire w_dff_B_L5JB73sA2_2;
	wire w_dff_B_BaXxZ3uv4_2;
	wire w_dff_B_blhrujv86_2;
	wire w_dff_B_523Asw6t5_2;
	wire w_dff_B_XW9bV9d58_2;
	wire w_dff_B_hwGE6lXr4_2;
	wire w_dff_B_m6GYAWr86_2;
	wire w_dff_B_M8HdBnQg3_2;
	wire w_dff_B_bNLhdBen5_2;
	wire w_dff_B_jl6Qpt129_2;
	wire w_dff_B_fy9fkraS8_2;
	wire w_dff_B_vROizhuz3_2;
	wire w_dff_B_FAcelAv48_2;
	wire w_dff_B_Te6PE2su3_2;
	wire w_dff_B_4ncCPWBp1_2;
	wire w_dff_B_dtLNku6w6_2;
	wire w_dff_B_IAVikLSt5_2;
	wire w_dff_B_825JNzyU2_2;
	wire w_dff_B_D0ocor7n0_2;
	wire w_dff_B_inUuGzy63_2;
	wire w_dff_B_Kd5ISFHJ0_2;
	wire w_dff_B_0Ct8Owza1_2;
	wire w_dff_B_J01f5gZB6_2;
	wire w_dff_B_VOLourEz6_2;
	wire w_dff_B_W3bsBN664_2;
	wire w_dff_B_dv8YtCXg3_2;
	wire w_dff_B_Qm3fjjHW8_2;
	wire w_dff_B_1wvE6DfL2_2;
	wire w_dff_B_k9m4mWxG5_2;
	wire w_dff_B_kEgN8ZEG5_2;
	wire w_dff_B_bQ8ocjeg3_2;
	wire w_dff_B_jdZKA79M3_2;
	wire w_dff_B_KtU7i8xS3_2;
	wire w_dff_B_ghOwIdW76_2;
	wire w_dff_B_3zRtCl133_2;
	wire w_dff_B_UW8CfZ038_2;
	wire w_dff_B_OF2s7hnL4_2;
	wire w_dff_B_PPlTCACc9_1;
	wire w_dff_A_MJhgLnrt6_1;
	wire w_dff_B_9d5lIpiV0_1;
	wire w_dff_B_ATDfNSBi9_2;
	wire w_dff_B_LcMhr7te4_2;
	wire w_dff_B_fwAdRSxc1_2;
	wire w_dff_B_FiJ6I9Kw9_2;
	wire w_dff_B_h26dof0y6_2;
	wire w_dff_B_M13B73Rl5_2;
	wire w_dff_B_7klzmQe00_2;
	wire w_dff_B_0amQgcDR7_2;
	wire w_dff_B_0GQtr2Pz5_2;
	wire w_dff_B_Fp40F1wp5_2;
	wire w_dff_B_CQzWXpjG9_2;
	wire w_dff_B_WzPFBeTY3_2;
	wire w_dff_B_nhQxcUvz6_2;
	wire w_dff_B_buPShKzW5_2;
	wire w_dff_B_A6a9nHVX3_2;
	wire w_dff_B_UZS45at09_2;
	wire w_dff_B_tf2hMgAb3_2;
	wire w_dff_B_uVVKptxL7_2;
	wire w_dff_B_wYPlqcNd4_2;
	wire w_dff_B_BjnLBjEC6_2;
	wire w_dff_B_su1LrFrP6_2;
	wire w_dff_B_o54ktGE82_2;
	wire w_dff_B_X5jePmM40_2;
	wire w_dff_B_12YaLQ0O4_2;
	wire w_dff_B_M8pe2DeQ2_2;
	wire w_dff_B_67ubSu1H8_2;
	wire w_dff_B_RXyLOIHN0_2;
	wire w_dff_B_UKqOHD4M8_2;
	wire w_dff_B_lOJF4shG3_2;
	wire w_dff_B_61IsavOV3_2;
	wire w_dff_B_orlTxHSF1_2;
	wire w_dff_B_Aos02Svp1_2;
	wire w_dff_B_jWRVVLyV4_2;
	wire w_dff_B_cAOgaJXH0_2;
	wire w_dff_B_M9r7IJP04_2;
	wire w_dff_B_Mfh0kkv02_1;
	wire w_dff_B_23vx0GH01_2;
	wire w_dff_B_TNlgw6GN2_2;
	wire w_dff_B_WZCe2WkR3_2;
	wire w_dff_B_wkb3VJOY5_2;
	wire w_dff_B_TKPoNh7x1_2;
	wire w_dff_B_Dpjta17I5_2;
	wire w_dff_B_EooeiXEp8_2;
	wire w_dff_B_yA5dxsfP7_2;
	wire w_dff_B_BGLINkCJ1_2;
	wire w_dff_B_Itf4hP8e8_2;
	wire w_dff_B_seAxaf2Q7_2;
	wire w_dff_B_yuPoDNyZ2_2;
	wire w_dff_B_HgiqbXGI1_2;
	wire w_dff_B_2zaxelzr8_2;
	wire w_dff_B_kR7qHsBI9_2;
	wire w_dff_B_vt4oSdHW1_2;
	wire w_dff_B_jvpwUup52_2;
	wire w_dff_B_F0QEjJoF4_2;
	wire w_dff_B_qGgJHG8F2_2;
	wire w_dff_B_xnKraAcX6_2;
	wire w_dff_B_fGX8GYOV2_2;
	wire w_dff_B_dH9KQSq26_2;
	wire w_dff_B_RMtLGD6b1_2;
	wire w_dff_B_9LfUq9Ol8_2;
	wire w_dff_B_7sG1xqag1_2;
	wire w_dff_B_78oPaTnY2_2;
	wire w_dff_B_7DGOZhca9_2;
	wire w_dff_B_TDQazCe19_2;
	wire w_dff_B_ERWAJdHi6_2;
	wire w_dff_B_kC9lnoRe0_2;
	wire w_dff_B_ZIjzh16U2_2;
	wire w_dff_B_kLPA1nxm0_2;
	wire w_dff_B_t9QCbYnh7_1;
	wire w_dff_B_rFKOjRJD1_2;
	wire w_dff_B_Shkzqvwb0_2;
	wire w_dff_B_7LkwtkoP0_2;
	wire w_dff_B_kA4fFiSm0_2;
	wire w_dff_B_CWWJfgdC8_2;
	wire w_dff_B_JvBhLCxV4_2;
	wire w_dff_B_MCM2zMCV8_2;
	wire w_dff_B_OkG67PvN7_2;
	wire w_dff_B_eKw7XMBP8_2;
	wire w_dff_B_0UktzvSF0_2;
	wire w_dff_B_E0nCYUDn0_2;
	wire w_dff_B_yZNCcRCE1_2;
	wire w_dff_B_0x3WEO4a7_2;
	wire w_dff_B_HtG1hsF88_2;
	wire w_dff_B_kHof0M1V0_2;
	wire w_dff_B_dTu2bsFh9_2;
	wire w_dff_B_FBdQq1Ql5_2;
	wire w_dff_B_UotZ01n04_2;
	wire w_dff_B_kJBVrZbv9_2;
	wire w_dff_B_fiE1NPPs0_2;
	wire w_dff_B_3BSHEZxH4_2;
	wire w_dff_B_J4bdGMyz8_2;
	wire w_dff_B_iqb96eDF6_2;
	wire w_dff_B_nmskeV6s8_2;
	wire w_dff_B_ovsV0Zdr1_2;
	wire w_dff_B_4gEHlifp4_2;
	wire w_dff_B_2WrrBva48_2;
	wire w_dff_B_pZFYSmTh4_2;
	wire w_dff_B_hux4zV000_2;
	wire w_dff_B_gQxEYNeQ5_1;
	wire w_dff_B_DlDxXjjK6_2;
	wire w_dff_B_z8eyT1QK9_2;
	wire w_dff_B_6tu7Q9JE6_2;
	wire w_dff_B_6CGTOujS7_2;
	wire w_dff_B_tf71UJPL0_2;
	wire w_dff_B_vFBEuL2u5_2;
	wire w_dff_B_LYshGEXw5_2;
	wire w_dff_B_m8QAwYiR9_2;
	wire w_dff_B_0u1XMU7m9_2;
	wire w_dff_B_5OWcZrHL8_2;
	wire w_dff_B_JuhOzneL0_2;
	wire w_dff_B_LcNVsmoM5_2;
	wire w_dff_B_THtRRqyG5_2;
	wire w_dff_B_l3cwipV46_2;
	wire w_dff_B_UDJerUTc1_2;
	wire w_dff_B_9SoRBjwU6_2;
	wire w_dff_B_fBJv6lFq8_2;
	wire w_dff_B_edIW2JsD6_2;
	wire w_dff_B_Oj5RJE7y5_2;
	wire w_dff_B_cvpuUafq9_2;
	wire w_dff_B_bfJbFLVg9_2;
	wire w_dff_B_cV1fiaF85_2;
	wire w_dff_B_HyFwnOSo1_2;
	wire w_dff_B_fg2E7zCH3_2;
	wire w_dff_B_8mTW0Vt24_2;
	wire w_dff_B_OrMlmBB98_2;
	wire w_dff_B_nhgki9g39_1;
	wire w_dff_B_xIgz8OAf0_2;
	wire w_dff_B_kCjKU8d75_2;
	wire w_dff_B_CJrmh1Ng1_2;
	wire w_dff_B_6zgyirgm6_2;
	wire w_dff_B_nWS3J3vD4_2;
	wire w_dff_B_D3kcCUWA4_2;
	wire w_dff_B_XVspSW4K0_2;
	wire w_dff_B_vAV6LjBg5_2;
	wire w_dff_B_tDDOjzAo6_2;
	wire w_dff_B_YpgkdWoU9_2;
	wire w_dff_B_pg2c2Vva2_2;
	wire w_dff_B_P58eNly96_2;
	wire w_dff_B_wx3ONJIR5_2;
	wire w_dff_B_KtJuHBNA3_2;
	wire w_dff_B_Cn3U6h028_2;
	wire w_dff_B_tQZnQ0fb9_2;
	wire w_dff_B_RzYDs5yO4_2;
	wire w_dff_B_hsNE3Nwh0_2;
	wire w_dff_B_J84qplZY5_2;
	wire w_dff_B_R3Cmfkw32_2;
	wire w_dff_B_YiiwBcoV5_2;
	wire w_dff_B_qM3TMyS62_2;
	wire w_dff_B_eLwyZtca5_2;
	wire w_dff_B_J41R32b15_1;
	wire w_dff_B_SvmA60150_2;
	wire w_dff_B_HNdLjouM6_2;
	wire w_dff_B_2oalaXv76_2;
	wire w_dff_B_b7ePqXwK0_2;
	wire w_dff_B_3MM1mVp90_2;
	wire w_dff_B_KInYzAAL3_2;
	wire w_dff_B_GxmMdB2Z3_2;
	wire w_dff_B_Hfon6AiE8_2;
	wire w_dff_B_e2miI3D60_2;
	wire w_dff_B_YiRbJM8b7_2;
	wire w_dff_B_dImp38AW0_2;
	wire w_dff_B_N7fAZGqV3_2;
	wire w_dff_B_V76RIVTO0_2;
	wire w_dff_B_nntKykwv5_2;
	wire w_dff_B_SkCr0Hsw8_2;
	wire w_dff_B_N3Gz4a417_2;
	wire w_dff_B_PKsD9SUp7_2;
	wire w_dff_B_PNtD6FEn9_2;
	wire w_dff_B_PrzCxOEQ4_2;
	wire w_dff_B_JSHBTzFy4_2;
	wire w_dff_B_4RoCyyc49_1;
	wire w_dff_B_TeSDMvrh9_2;
	wire w_dff_B_aB2ruGhT5_2;
	wire w_dff_B_tHCvUFej1_2;
	wire w_dff_B_k51qxMxG3_2;
	wire w_dff_B_vwTaCo179_2;
	wire w_dff_B_dmIEIi6K7_2;
	wire w_dff_B_NfJJlwcQ6_2;
	wire w_dff_B_2ot4aw1P1_2;
	wire w_dff_B_DZ5TuKAr0_2;
	wire w_dff_B_Qr6KONTB9_2;
	wire w_dff_B_D7mpqHaZ9_2;
	wire w_dff_B_8ap9XZ2G5_2;
	wire w_dff_B_znAvAf1b6_2;
	wire w_dff_B_g7Ajp1Jz1_2;
	wire w_dff_B_2inuqmvb5_2;
	wire w_dff_B_DCbt8AsM8_2;
	wire w_dff_B_4OhSnjHB1_1;
	wire w_dff_B_BTvLNqp24_2;
	wire w_dff_B_vTRdyL2n2_2;
	wire w_dff_B_zvqJp2eF7_2;
	wire w_dff_B_cwdt00yb6_2;
	wire w_dff_B_IswTWwiX8_2;
	wire w_dff_B_jxVmJiKd6_2;
	wire w_dff_B_zh7bGbAO1_2;
	wire w_dff_B_0TuTl3f45_2;
	wire w_dff_B_d1OaOJdv0_2;
	wire w_dff_B_JPghaI0L5_2;
	wire w_dff_B_egHK3uEz1_2;
	wire w_dff_B_RZrGdPql2_2;
	wire w_dff_B_3yEfr7Fd2_2;
	wire w_dff_B_ohS8euDz2_2;
	wire w_dff_B_Z1wAO6IW1_1;
	wire w_dff_B_hYHZV2MK6_2;
	wire w_dff_B_EoSu7nZR4_2;
	wire w_dff_B_pQ7rdIDj2_2;
	wire w_dff_B_u56fcKA50_2;
	wire w_dff_B_DG8su0CU4_2;
	wire w_dff_B_YRfhCypi6_2;
	wire w_dff_B_Ir9LbLhO6_2;
	wire w_dff_B_HttjD7nw6_2;
	wire w_dff_B_DdM4YSNl6_2;
	wire w_dff_B_ojq0lhco6_2;
	wire w_dff_B_SCpfItVk0_2;
	wire w_dff_B_GRLdMi0n6_2;
	wire w_dff_B_uCF6h73s2_1;
	wire w_dff_B_GQevH8ws1_2;
	wire w_dff_B_LNr8B91J1_2;
	wire w_dff_B_sF7dip1X2_2;
	wire w_dff_B_hHMrYJ236_2;
	wire w_dff_B_TsMGOJSZ7_2;
	wire w_dff_B_ECwcD2uT7_2;
	wire w_dff_B_DyxwykNC8_2;
	wire w_dff_B_DFFMty2n4_2;
	wire w_dff_B_eRfLbmES2_2;
	wire w_dff_B_fhVItzJa8_2;
	wire w_dff_B_btSQe1sk0_1;
	wire w_dff_B_kYGGRyUY3_2;
	wire w_dff_B_ox39bHL71_2;
	wire w_dff_B_Z1Tk8c419_2;
	wire w_dff_B_WcfT0iQs9_2;
	wire w_dff_B_FmNfYIGZ8_2;
	wire w_dff_B_uwN240CB0_2;
	wire w_dff_B_JpgEOsly0_2;
	wire w_dff_B_qnHQNVmE9_2;
	wire w_dff_B_Zo9yzJzN1_1;
	wire w_dff_B_MTgunAhx5_2;
	wire w_dff_B_LxDlauum6_2;
	wire w_dff_B_OkmFtaPm9_2;
	wire w_dff_B_ZQiwqMjc1_2;
	wire w_dff_B_O92jqehP3_2;
	wire w_dff_B_4Nkw4hr37_2;
	wire w_dff_B_3rRbXLt23_2;
	wire w_dff_B_HkCdJwym8_1;
	wire w_dff_B_JjdrgagQ2_1;
	wire w_dff_B_K5lJlIMz8_1;
	wire w_dff_B_bQeuhAse3_1;
	wire w_dff_B_2vmf0QpN2_0;
	wire w_dff_A_kn0zsOHZ1_0;
	wire w_dff_A_VSjoUpi55_0;
	wire w_dff_B_q3fbxToc8_1;
	wire w_dff_B_hW2Wvec32_1;
	wire w_dff_A_LyIyUKHN6_0;
	wire w_dff_A_eDaH1P4c2_1;
	wire w_dff_A_2sY683Rr3_1;
	wire w_dff_A_A2WbjbgF7_1;
	wire w_dff_A_otQYMIni3_1;
	wire w_dff_A_BMghvNX15_1;
	wire w_dff_A_ZUEwSf3U7_1;
	wire w_dff_B_FtolqQ735_2;
	wire w_dff_B_oDu8Eos25_1;
	wire w_dff_B_wE04I4wQ7_2;
	wire w_dff_B_WPoClSER5_2;
	wire w_dff_B_9jFKQ7Qe6_2;
	wire w_dff_B_3vISEgVn9_2;
	wire w_dff_B_LMHezgEo1_2;
	wire w_dff_B_DrmD3htz3_2;
	wire w_dff_B_aRQaRnW97_2;
	wire w_dff_B_0J6AqRQK6_2;
	wire w_dff_B_oVV8g6Wz0_2;
	wire w_dff_B_b3OkEBx99_2;
	wire w_dff_B_moH1uWoa4_2;
	wire w_dff_B_KOlyZ0ow3_2;
	wire w_dff_B_l83gPR0X3_2;
	wire w_dff_B_RDXnum4J2_2;
	wire w_dff_B_wDr9hJYf0_2;
	wire w_dff_B_VMaPysuh0_2;
	wire w_dff_B_VlxA28bb9_2;
	wire w_dff_B_zUUnFJhj7_2;
	wire w_dff_B_lAzmWaIV7_2;
	wire w_dff_B_yB6oESIv2_2;
	wire w_dff_B_jwiJ97kX1_2;
	wire w_dff_B_6lEq9Y0Z3_2;
	wire w_dff_B_vqzYn8lU8_2;
	wire w_dff_B_1XG43kcY1_2;
	wire w_dff_B_gKeuf43y5_2;
	wire w_dff_B_UVIDGLvI5_2;
	wire w_dff_B_8gZXkZhv1_2;
	wire w_dff_B_mWvWq0mM1_2;
	wire w_dff_B_lfFVa1rS3_2;
	wire w_dff_B_cMm6NwEp9_2;
	wire w_dff_B_FrkmIl2f8_2;
	wire w_dff_B_A5xSx0WC3_2;
	wire w_dff_B_g4GTYxdT2_2;
	wire w_dff_B_47TwFNvY3_2;
	wire w_dff_B_hJsATW6V2_2;
	wire w_dff_B_mJNAisik9_2;
	wire w_dff_B_0SVjtCIX1_2;
	wire w_dff_B_gpdaZKjh0_2;
	wire w_dff_B_TWMzhGLa5_2;
	wire w_dff_B_fOOVUDPi4_2;
	wire w_dff_B_VtmnVXvW9_1;
	wire w_dff_A_QTN0cg9q0_1;
	wire w_dff_B_w79I0pZh7_1;
	wire w_dff_B_pUSpDTaA0_2;
	wire w_dff_B_GN3mywOV4_2;
	wire w_dff_B_Y27DkaB65_2;
	wire w_dff_B_EW2gWXP37_2;
	wire w_dff_B_OWesw7EV2_2;
	wire w_dff_B_V9dfz1PV0_2;
	wire w_dff_B_jjl6BbRA8_2;
	wire w_dff_B_TGg6UeiO9_2;
	wire w_dff_B_Zj5eYONl5_2;
	wire w_dff_B_y3aVR0YG7_2;
	wire w_dff_B_HEgBnuS27_2;
	wire w_dff_B_xXvrscyu6_2;
	wire w_dff_B_Qp1d1mau4_2;
	wire w_dff_B_lG8w9RrV6_2;
	wire w_dff_B_9QagDsVE9_2;
	wire w_dff_B_MF1CteWo4_2;
	wire w_dff_B_uNMQNpGD1_2;
	wire w_dff_B_zNvTlqqJ1_2;
	wire w_dff_B_Pu4h1Rhb2_2;
	wire w_dff_B_IE5tZrss2_2;
	wire w_dff_B_S7q4Qtl86_2;
	wire w_dff_B_GvyM50q32_2;
	wire w_dff_B_1NznSJST7_2;
	wire w_dff_B_KdSZogl33_2;
	wire w_dff_B_xeMLRUnC2_2;
	wire w_dff_B_SwXlRdzX1_2;
	wire w_dff_B_ScKyS4B77_2;
	wire w_dff_B_joK65iE04_2;
	wire w_dff_B_QiylpfWj0_2;
	wire w_dff_B_klfPiP2b1_2;
	wire w_dff_B_34A0kQTu3_2;
	wire w_dff_B_PIJFLx1L5_2;
	wire w_dff_B_prvxyJRV3_2;
	wire w_dff_B_msAlT3NN1_2;
	wire w_dff_B_cEZ81KbZ7_2;
	wire w_dff_B_e9uZd5Xu4_2;
	wire w_dff_B_uzlAELXW4_1;
	wire w_dff_B_XGLiY6PA6_2;
	wire w_dff_B_ST0ofe5k8_2;
	wire w_dff_B_8jeB2cXW2_2;
	wire w_dff_B_vdozkldW1_2;
	wire w_dff_B_hyhrJQt76_2;
	wire w_dff_B_d56VUmTU5_2;
	wire w_dff_B_uaYRbAyu2_2;
	wire w_dff_B_7Pxqdi6r0_2;
	wire w_dff_B_MRxzjgj11_2;
	wire w_dff_B_FYKSD3Pk9_2;
	wire w_dff_B_z7P477AF0_2;
	wire w_dff_B_hlM2dhGm6_2;
	wire w_dff_B_EWpUSGtz4_2;
	wire w_dff_B_t9NNhls08_2;
	wire w_dff_B_rk4pTLwE0_2;
	wire w_dff_B_7wlW9M3z8_2;
	wire w_dff_B_a7mHvGl83_2;
	wire w_dff_B_HymIFP8n3_2;
	wire w_dff_B_DW4G04bT5_2;
	wire w_dff_B_rWwPLB758_2;
	wire w_dff_B_2VQrcCgK2_2;
	wire w_dff_B_pA0W8bSL7_2;
	wire w_dff_B_y9SKUnQx5_2;
	wire w_dff_B_3HSnwsKf0_2;
	wire w_dff_B_xspFNcCs8_2;
	wire w_dff_B_uWz50CfM8_2;
	wire w_dff_B_PyGURnay0_2;
	wire w_dff_B_ZaYQw5px6_2;
	wire w_dff_B_FVaAM92D7_2;
	wire w_dff_B_I9hJsUs91_2;
	wire w_dff_B_alX2ptos8_2;
	wire w_dff_B_ecNw3eAu0_2;
	wire w_dff_B_AZwRkMcO5_2;
	wire w_dff_B_GPX5xaK20_1;
	wire w_dff_B_whCcbEjm7_2;
	wire w_dff_B_nxNef3lo2_2;
	wire w_dff_B_6tPNCA2y3_2;
	wire w_dff_B_dc0nmtWc6_2;
	wire w_dff_B_4Hn6O43Q7_2;
	wire w_dff_B_uu67OFuM1_2;
	wire w_dff_B_CVAwNBkm8_2;
	wire w_dff_B_RIA7IBCW3_2;
	wire w_dff_B_K5wy189X4_2;
	wire w_dff_B_Uy3DKsy39_2;
	wire w_dff_B_kPMyouda2_2;
	wire w_dff_B_r1ESw0DD5_2;
	wire w_dff_B_BOiVgtA71_2;
	wire w_dff_B_YE6REcEF7_2;
	wire w_dff_B_KS0eGR7P0_2;
	wire w_dff_B_3RHtpPH64_2;
	wire w_dff_B_2a2N7mhl7_2;
	wire w_dff_B_rj898B917_2;
	wire w_dff_B_weBxvRr00_2;
	wire w_dff_B_uL9aGcpt6_2;
	wire w_dff_B_YmFRj0EE0_2;
	wire w_dff_B_FbK8rl8x7_2;
	wire w_dff_B_2S5DYXY75_2;
	wire w_dff_B_BcnR6s569_2;
	wire w_dff_B_AoyNyvj77_2;
	wire w_dff_B_yGFJtCAs3_2;
	wire w_dff_B_YGfIopuj4_2;
	wire w_dff_B_2cFuOeDU0_2;
	wire w_dff_B_aRYoTqZk7_2;
	wire w_dff_B_F32ynQNJ0_2;
	wire w_dff_B_D2vrndJ97_1;
	wire w_dff_B_L17nLg5l4_2;
	wire w_dff_B_5blouBsA0_2;
	wire w_dff_B_JwvTDodC5_2;
	wire w_dff_B_If3nmpXj2_2;
	wire w_dff_B_juTBOYVR3_2;
	wire w_dff_B_Ctgey6160_2;
	wire w_dff_B_TeGskrw05_2;
	wire w_dff_B_38jb5Q205_2;
	wire w_dff_B_bV8NVUoR3_2;
	wire w_dff_B_uCV82ucR5_2;
	wire w_dff_B_gscPhUYH3_2;
	wire w_dff_B_A3GUBsnS7_2;
	wire w_dff_B_L93BWW0A6_2;
	wire w_dff_B_Q8ePGlag2_2;
	wire w_dff_B_A9V7suDM9_2;
	wire w_dff_B_6AK9eN9L2_2;
	wire w_dff_B_8UbFGlfN6_2;
	wire w_dff_B_NkJRKOzt5_2;
	wire w_dff_B_p1pj7nQ12_2;
	wire w_dff_B_WopICEiV5_2;
	wire w_dff_B_jlm51HI61_2;
	wire w_dff_B_YiQsSk0w6_2;
	wire w_dff_B_Rj7RXo2o3_2;
	wire w_dff_B_ltHDEBBi5_2;
	wire w_dff_B_w8o70wwS1_2;
	wire w_dff_B_kV5tHOnr0_2;
	wire w_dff_B_RK8XfEmu7_2;
	wire w_dff_B_xbndg6UF9_1;
	wire w_dff_B_3duHWKSw1_2;
	wire w_dff_B_hMrCfNmP0_2;
	wire w_dff_B_ued6c8hn6_2;
	wire w_dff_B_0T2T7uX31_2;
	wire w_dff_B_K473yoNF6_2;
	wire w_dff_B_eIqr0LMd6_2;
	wire w_dff_B_0MafWtwn9_2;
	wire w_dff_B_HadeiXsy8_2;
	wire w_dff_B_k6OJn5kx9_2;
	wire w_dff_B_1dDA4z7V2_2;
	wire w_dff_B_NkGUXd290_2;
	wire w_dff_B_H4ua56G17_2;
	wire w_dff_B_iNgeChwW9_2;
	wire w_dff_B_dvyf9QtG9_2;
	wire w_dff_B_tD7Grgwh6_2;
	wire w_dff_B_woIbjkXG8_2;
	wire w_dff_B_JI6S2RWY0_2;
	wire w_dff_B_1gNAIQ9X0_2;
	wire w_dff_B_fGeimlpM8_2;
	wire w_dff_B_dHQ0tyAa9_2;
	wire w_dff_B_PBiYnNvT5_2;
	wire w_dff_B_bBBRdh0W6_2;
	wire w_dff_B_fZVZwQfO1_2;
	wire w_dff_B_1zPUAOOj0_2;
	wire w_dff_B_mq9duBnh9_1;
	wire w_dff_B_qbRJKyut9_2;
	wire w_dff_B_wuosGH5V1_2;
	wire w_dff_B_c3XFSywN0_2;
	wire w_dff_B_ggIqvUyK8_2;
	wire w_dff_B_bTEMI6yI5_2;
	wire w_dff_B_A5JwVM7p1_2;
	wire w_dff_B_1IPvVJBd3_2;
	wire w_dff_B_3GYeeXMU2_2;
	wire w_dff_B_RtRMlLV93_2;
	wire w_dff_B_oVkS2rzQ3_2;
	wire w_dff_B_K4pDD6M35_2;
	wire w_dff_B_hFaZx0Bc5_2;
	wire w_dff_B_okyOLNjQ6_2;
	wire w_dff_B_Gis1WVFi2_2;
	wire w_dff_B_h9cdILAj4_2;
	wire w_dff_B_wmlXPwbF6_2;
	wire w_dff_B_aL9HpEFT0_2;
	wire w_dff_B_8lkL9us34_2;
	wire w_dff_B_9cISku7Y0_2;
	wire w_dff_B_pdMKyQz74_2;
	wire w_dff_B_4s9CXQls9_2;
	wire w_dff_B_9Uieaijd3_1;
	wire w_dff_B_Y1aFg7n48_2;
	wire w_dff_B_Q5WBLFOM6_2;
	wire w_dff_B_4CD5K0WO2_2;
	wire w_dff_B_xg1Q4P7h1_2;
	wire w_dff_B_LOaAFG0N9_2;
	wire w_dff_B_IPNKcema4_2;
	wire w_dff_B_hXwMf1Ln9_2;
	wire w_dff_B_1bsqlHYF9_2;
	wire w_dff_B_McmQJbeL0_2;
	wire w_dff_B_un1QwpFL6_2;
	wire w_dff_B_fTUIecfe6_2;
	wire w_dff_B_rUBvjqU23_2;
	wire w_dff_B_S0QUyd4z4_2;
	wire w_dff_B_cAiFs1Vr8_2;
	wire w_dff_B_UVYNXiRD1_2;
	wire w_dff_B_CYMYmG617_2;
	wire w_dff_B_uRS1Fs5X4_2;
	wire w_dff_B_q9ZmF9Nl0_2;
	wire w_dff_B_HCm4HMBu5_1;
	wire w_dff_B_q9mQfUMn5_2;
	wire w_dff_B_nfTIO8SG3_2;
	wire w_dff_B_7vMXlgty7_2;
	wire w_dff_B_zm8HHnEn6_2;
	wire w_dff_B_gcJP6ez38_2;
	wire w_dff_B_tF12xAQA2_2;
	wire w_dff_B_zzMGZgxv0_2;
	wire w_dff_B_iagYopDK9_2;
	wire w_dff_B_OfSWPD290_2;
	wire w_dff_B_3xQwQFwN0_2;
	wire w_dff_B_T1iRrGLI7_2;
	wire w_dff_B_5LjnzKQR7_2;
	wire w_dff_B_5u09NmvF9_2;
	wire w_dff_B_QM2ywPH17_2;
	wire w_dff_B_n6F9CT944_1;
	wire w_dff_B_Lq5fEtnU3_2;
	wire w_dff_B_4psRx6Yd0_2;
	wire w_dff_B_Vj1T40aS7_2;
	wire w_dff_B_2eMXGhJK5_2;
	wire w_dff_B_PvCWoQ7I2_2;
	wire w_dff_B_6PAIGnOV5_2;
	wire w_dff_B_Qs6leghL9_2;
	wire w_dff_B_aCo1Nzek7_2;
	wire w_dff_B_2KFS5uS59_2;
	wire w_dff_B_vAsbNvhD8_2;
	wire w_dff_B_JZB4b0q48_2;
	wire w_dff_B_bPAnp4Pw3_2;
	wire w_dff_B_yZPdh5aS0_1;
	wire w_dff_B_8NERdX2u5_2;
	wire w_dff_B_25ePHiwQ0_2;
	wire w_dff_B_OjrspeHH2_2;
	wire w_dff_B_PrMWFye28_2;
	wire w_dff_B_yrEi0ERg7_2;
	wire w_dff_B_hDpMZG5I2_2;
	wire w_dff_B_KrtJe9nO0_2;
	wire w_dff_B_OjXLKmvU7_2;
	wire w_dff_B_vQ5CrLRN0_2;
	wire w_dff_B_aUyLW4GW0_2;
	wire w_dff_B_9guddiw18_1;
	wire w_dff_B_eKp7kmg04_2;
	wire w_dff_B_9WnfpqXH4_2;
	wire w_dff_B_RfXqs3bx6_2;
	wire w_dff_B_FGSvVmyF6_2;
	wire w_dff_B_5VFTNBQV9_2;
	wire w_dff_B_d2WCO8lh7_2;
	wire w_dff_B_X6Lj8DZw4_2;
	wire w_dff_B_BOKcLPJE6_2;
	wire w_dff_B_3bznItpR8_1;
	wire w_dff_B_QskTUZIl3_2;
	wire w_dff_B_RYCKGT0Q5_2;
	wire w_dff_B_sJ6bMRPw3_2;
	wire w_dff_B_biN26TeG1_2;
	wire w_dff_B_wRKrBqAU8_2;
	wire w_dff_B_VWcRMS4Q8_2;
	wire w_dff_B_myQNXNk33_2;
	wire w_dff_B_Lrk1rPAU7_1;
	wire w_dff_B_kFdm4MWi7_1;
	wire w_dff_B_vvLap90t0_1;
	wire w_dff_B_SinQdaEY4_1;
	wire w_dff_B_46YEwWPG7_0;
	wire w_dff_A_7gZ8IHFB9_0;
	wire w_dff_A_KFl8vlWw0_0;
	wire w_dff_B_DXAcwMA30_1;
	wire w_dff_B_edoKP4GI5_1;
	wire w_dff_A_HhWBU4898_0;
	wire w_dff_A_lAmDUymv7_1;
	wire w_dff_A_2TJbBS0Z7_1;
	wire w_dff_A_FRrxhEYW4_1;
	wire w_dff_A_Q7cGH8RO6_1;
	wire w_dff_A_p5LVvmLl1_1;
	wire w_dff_A_RG9ph2SF1_1;
	wire w_dff_B_wybVeYra2_1;
	wire w_dff_A_u5pAxSPk8_1;
	wire w_dff_B_qjFxCdra6_1;
	wire w_dff_B_yCkoQuUi0_2;
	wire w_dff_B_1e03jPNi0_2;
	wire w_dff_B_xQoFEX040_2;
	wire w_dff_B_ra0NijEe4_2;
	wire w_dff_B_UaMnAFWO9_2;
	wire w_dff_B_qE9jf3qt6_2;
	wire w_dff_B_PUhi8Dkh0_2;
	wire w_dff_B_RF9PSkZe0_2;
	wire w_dff_B_kcai8zi98_2;
	wire w_dff_B_t9f1Af0y4_2;
	wire w_dff_B_iw2sIcTV5_2;
	wire w_dff_B_2IF9iQa65_2;
	wire w_dff_B_sjjoRjtA5_2;
	wire w_dff_B_OdVFeRCh5_2;
	wire w_dff_B_5FTypbtR2_2;
	wire w_dff_B_ch4Q0btC4_2;
	wire w_dff_B_Q97Vn3KM9_2;
	wire w_dff_B_SGvt6UJa9_2;
	wire w_dff_B_5fu915K48_2;
	wire w_dff_B_6pFmFVng7_2;
	wire w_dff_B_VwfjHoz96_2;
	wire w_dff_B_GYtKx0dE7_2;
	wire w_dff_B_KELZep1v7_2;
	wire w_dff_B_VNolA4Gw4_2;
	wire w_dff_B_OpZJGWqX4_2;
	wire w_dff_B_rAV5wLlQ9_2;
	wire w_dff_B_QVAfIkqJ5_2;
	wire w_dff_B_TYnkcW1S4_2;
	wire w_dff_B_6T2ExHXD0_2;
	wire w_dff_B_ZM7cu7DM2_2;
	wire w_dff_B_OrqWsJcW6_2;
	wire w_dff_B_A2h5ueLQ4_2;
	wire w_dff_B_Vba05DfR4_2;
	wire w_dff_B_djfyHTtY4_2;
	wire w_dff_B_CmAepxs86_2;
	wire w_dff_B_1QVlvKW01_2;
	wire w_dff_B_8tTAcvvi7_2;
	wire w_dff_B_TWgjBk507_2;
	wire w_dff_B_gMcNfZFB1_2;
	wire w_dff_B_ns7ZlvK11_2;
	wire w_dff_B_UJvMBvYk0_1;
	wire w_dff_B_EKvOAogf7_2;
	wire w_dff_B_rEQ7fuDk2_2;
	wire w_dff_B_VHdlrsMb1_2;
	wire w_dff_B_oPHqpkro3_2;
	wire w_dff_B_NDNbkwMM0_2;
	wire w_dff_B_MNBCwN6r7_2;
	wire w_dff_B_hvAPfKwF1_2;
	wire w_dff_B_3BYyu9rc2_2;
	wire w_dff_B_JPztbNPO0_2;
	wire w_dff_B_NgSs98cJ7_2;
	wire w_dff_B_kNfAVgwe7_2;
	wire w_dff_B_bGUoieEQ3_2;
	wire w_dff_B_RZa459qO5_2;
	wire w_dff_B_2FNNks7r0_2;
	wire w_dff_B_QhpERBK61_2;
	wire w_dff_B_7tr5QZs43_2;
	wire w_dff_B_wVrT1kfe4_2;
	wire w_dff_B_k7dh23Rn4_2;
	wire w_dff_B_xIQTt2et3_2;
	wire w_dff_B_rK5x8xpK2_2;
	wire w_dff_B_p2ixqy236_2;
	wire w_dff_B_MKbRpjeb4_2;
	wire w_dff_B_nL4qBlji4_2;
	wire w_dff_B_YTOHoNPs5_2;
	wire w_dff_B_L5f6J1xD0_2;
	wire w_dff_B_tBj7tZXG6_2;
	wire w_dff_B_5d7FUVW01_2;
	wire w_dff_B_FkjliwCP0_2;
	wire w_dff_B_35VTTjpI3_2;
	wire w_dff_B_XbnCMaL31_2;
	wire w_dff_B_ldc8JbMJ1_2;
	wire w_dff_B_l5SJSHRB9_2;
	wire w_dff_B_Ltf8FQDi6_2;
	wire w_dff_B_PrRunnAa2_2;
	wire w_dff_B_Bde1EA6x9_2;
	wire w_dff_B_76gp0Rog3_2;
	wire w_dff_B_iECabImR9_2;
	wire w_dff_B_nZYIJf9U5_1;
	wire w_dff_B_hAWd6X2I7_2;
	wire w_dff_B_3BXniUrU8_2;
	wire w_dff_B_1tTLeYlX7_2;
	wire w_dff_B_D4Ci9jFe0_2;
	wire w_dff_B_x38QwtGm5_2;
	wire w_dff_B_ogC7HuXu1_2;
	wire w_dff_B_ttQoC9nM3_2;
	wire w_dff_B_TMxwLvs78_2;
	wire w_dff_B_NZA6LmIg5_2;
	wire w_dff_B_v8avHYxQ2_2;
	wire w_dff_B_BqwtLHPy4_2;
	wire w_dff_B_Ls9wD5yV7_2;
	wire w_dff_B_sqKeiqba4_2;
	wire w_dff_B_uZxK1mEw5_2;
	wire w_dff_B_l02ux8P57_2;
	wire w_dff_B_VTXcpGno5_2;
	wire w_dff_B_UMHsvwog6_2;
	wire w_dff_B_uf70UhdU7_2;
	wire w_dff_B_WIREeHOA0_2;
	wire w_dff_B_Pbyvcw4L7_2;
	wire w_dff_B_TDG2Xwug7_2;
	wire w_dff_B_JPFmGs7i0_2;
	wire w_dff_B_yXhAVOAH3_2;
	wire w_dff_B_nB63w51U6_2;
	wire w_dff_B_MFAq0b0S3_2;
	wire w_dff_B_zMgc9C2y5_2;
	wire w_dff_B_gq0HB0fj5_2;
	wire w_dff_B_i1yHj2xk0_2;
	wire w_dff_B_g5n5vMzb1_2;
	wire w_dff_B_Lhsb3wVl7_2;
	wire w_dff_B_wGzqms531_2;
	wire w_dff_B_L2DbcLkm2_2;
	wire w_dff_B_MoBDJCAb9_2;
	wire w_dff_B_57WarLly3_2;
	wire w_dff_B_jYStSG8v5_1;
	wire w_dff_B_xqSHurj93_2;
	wire w_dff_B_6iikLR6j0_2;
	wire w_dff_B_nXIcOcua4_2;
	wire w_dff_B_pm0H1Snv1_2;
	wire w_dff_B_pDswfDCN9_2;
	wire w_dff_B_ygak8jyn8_2;
	wire w_dff_B_gqoH7ibT2_2;
	wire w_dff_B_TteqE1v72_2;
	wire w_dff_B_CFsi77i09_2;
	wire w_dff_B_WknhPoEQ6_2;
	wire w_dff_B_5Cuul0bY8_2;
	wire w_dff_B_TDajjuti9_2;
	wire w_dff_B_dETZ3SFf3_2;
	wire w_dff_B_fY1hOuYd8_2;
	wire w_dff_B_CFjbB4Ce4_2;
	wire w_dff_B_Nvx1jjfw8_2;
	wire w_dff_B_v4vpzgSS8_2;
	wire w_dff_B_FmWSi48O6_2;
	wire w_dff_B_uACavA1d0_2;
	wire w_dff_B_81NOX0dO1_2;
	wire w_dff_B_eVpWkW8i4_2;
	wire w_dff_B_pN7WG8NT2_2;
	wire w_dff_B_7YCPFTpR1_2;
	wire w_dff_B_ffcm9BjM2_2;
	wire w_dff_B_wrB4E1tO5_2;
	wire w_dff_B_1fi7Cs1w5_2;
	wire w_dff_B_YbbN4NXA2_2;
	wire w_dff_B_Blk3KTr49_2;
	wire w_dff_B_6fqCdItL3_2;
	wire w_dff_B_GU9LaF1R2_2;
	wire w_dff_B_NHWP0S507_2;
	wire w_dff_B_ldo93EOQ0_1;
	wire w_dff_B_NxUqrVXg7_2;
	wire w_dff_B_lasVMYWE6_2;
	wire w_dff_B_zKdzvaCg6_2;
	wire w_dff_B_MDjZycQv2_2;
	wire w_dff_B_SVJIUgvq7_2;
	wire w_dff_B_zcXRgkLW2_2;
	wire w_dff_B_rvsuLzbT2_2;
	wire w_dff_B_ajsdusPr8_2;
	wire w_dff_B_yy9Qd3dZ9_2;
	wire w_dff_B_px0OmXg14_2;
	wire w_dff_B_XR3cI6gg8_2;
	wire w_dff_B_ZDFPikBD9_2;
	wire w_dff_B_qCnLjZR68_2;
	wire w_dff_B_y3mHFv1R1_2;
	wire w_dff_B_LHox4NkO8_2;
	wire w_dff_B_sE9ohvi66_2;
	wire w_dff_B_kxkQrPRe2_2;
	wire w_dff_B_Og0ANBxg0_2;
	wire w_dff_B_9cSl21ZY9_2;
	wire w_dff_B_shtL7e940_2;
	wire w_dff_B_k2uK6uLj3_2;
	wire w_dff_B_Gg2xaO4H1_2;
	wire w_dff_B_nAWGNiAQ1_2;
	wire w_dff_B_x0g9VDz81_2;
	wire w_dff_B_GmaskMIx0_2;
	wire w_dff_B_p0mF0xOr6_2;
	wire w_dff_B_Npw3mhl04_2;
	wire w_dff_B_BGR6rjw04_2;
	wire w_dff_B_pHEnIkim6_1;
	wire w_dff_B_Vy8FtmPu6_2;
	wire w_dff_B_jQTDYqi07_2;
	wire w_dff_B_kqEpPQvl2_2;
	wire w_dff_B_XIVADeVV0_2;
	wire w_dff_B_qQgOhVCK9_2;
	wire w_dff_B_zO9pOINM7_2;
	wire w_dff_B_mZCpK91W5_2;
	wire w_dff_B_mbg4fGvC2_2;
	wire w_dff_B_Wyr8CSu17_2;
	wire w_dff_B_6lo0pbBF7_2;
	wire w_dff_B_F7dR9jbP4_2;
	wire w_dff_B_6VGobh8y4_2;
	wire w_dff_B_EPNlYuey3_2;
	wire w_dff_B_5mPfdGQY9_2;
	wire w_dff_B_ApfSoGVI9_2;
	wire w_dff_B_yi03JjiU0_2;
	wire w_dff_B_UBLS2bwR1_2;
	wire w_dff_B_3unU2PrT8_2;
	wire w_dff_B_UuLPRUt52_2;
	wire w_dff_B_chwKB6sU9_2;
	wire w_dff_B_ec3W0gK28_2;
	wire w_dff_B_g0zwmJyW6_2;
	wire w_dff_B_4YywosL63_2;
	wire w_dff_B_HexU8YbC7_2;
	wire w_dff_B_iWMEV3TI9_2;
	wire w_dff_B_HcTs0byL2_1;
	wire w_dff_B_6PVzsnq21_2;
	wire w_dff_B_psVN11xF7_2;
	wire w_dff_B_VNxKUYAG3_2;
	wire w_dff_B_8Zk1SmxN3_2;
	wire w_dff_B_RMUaedLb5_2;
	wire w_dff_B_5ekJN1di7_2;
	wire w_dff_B_Stw6vIAy9_2;
	wire w_dff_B_eyXZtImS5_2;
	wire w_dff_B_eMyVEqZ17_2;
	wire w_dff_B_HEd30MXq6_2;
	wire w_dff_B_V4XjnTm12_2;
	wire w_dff_B_VDGvfSHX1_2;
	wire w_dff_B_sH9PoYqz0_2;
	wire w_dff_B_cj7s6ouI1_2;
	wire w_dff_B_okqjrnQH7_2;
	wire w_dff_B_q0mawQe65_2;
	wire w_dff_B_EMIhYefK4_2;
	wire w_dff_B_Ezs2lTVU5_2;
	wire w_dff_B_qk7JLf7v5_2;
	wire w_dff_B_NZzFJg3M8_2;
	wire w_dff_B_D87deOIr2_2;
	wire w_dff_B_uojRNQmk5_2;
	wire w_dff_B_fGZzhjhB6_1;
	wire w_dff_B_n17ZVxRT3_2;
	wire w_dff_B_R9V95fYB0_2;
	wire w_dff_B_APApAvjJ4_2;
	wire w_dff_B_W85EUjSY1_2;
	wire w_dff_B_7EaeYfsR7_2;
	wire w_dff_B_rJfKmYiA8_2;
	wire w_dff_B_r1BfFEvS5_2;
	wire w_dff_B_qe6iiy171_2;
	wire w_dff_B_lnwLFdiM6_2;
	wire w_dff_B_tiqfHTdP7_2;
	wire w_dff_B_SaZUhaoZ5_2;
	wire w_dff_B_1QzeL0RR4_2;
	wire w_dff_B_28BcldFj2_2;
	wire w_dff_B_n20NaSMn5_2;
	wire w_dff_B_SxJkGRgQ8_2;
	wire w_dff_B_T9meeg3C1_2;
	wire w_dff_B_9GiUuddW9_2;
	wire w_dff_B_EuRzVPuY5_2;
	wire w_dff_B_s1neHrrM3_2;
	wire w_dff_B_dFsHh26v2_1;
	wire w_dff_B_oZIRDm7s4_2;
	wire w_dff_B_PgxJ4dNf9_2;
	wire w_dff_B_MByjT5W80_2;
	wire w_dff_B_3zLb4nV35_2;
	wire w_dff_B_MnFLoEPa1_2;
	wire w_dff_B_6xbD8Xho5_2;
	wire w_dff_B_paexazBJ7_2;
	wire w_dff_B_D3uaoPtH8_2;
	wire w_dff_B_v9D0bK746_2;
	wire w_dff_B_FQrQ3fBc5_2;
	wire w_dff_B_fApgYZmH1_2;
	wire w_dff_B_PdRg3K7r0_2;
	wire w_dff_B_vJ4Ybcxj4_2;
	wire w_dff_B_AIb5Liqz6_2;
	wire w_dff_B_y3BcU3Is6_2;
	wire w_dff_B_575PgbKq3_2;
	wire w_dff_B_14tFs7Lf3_1;
	wire w_dff_B_XTDYzMiw6_2;
	wire w_dff_B_u0ycFSqx9_2;
	wire w_dff_B_SyVbmMo31_2;
	wire w_dff_B_HmnsD02t1_2;
	wire w_dff_B_CrQh6mNC3_2;
	wire w_dff_B_hGdeg0wU5_2;
	wire w_dff_B_FbOgMmUl2_2;
	wire w_dff_B_q1g83Cs38_2;
	wire w_dff_B_J9m7R1mc3_2;
	wire w_dff_B_nd2iupUz6_2;
	wire w_dff_B_I7LmuTso3_2;
	wire w_dff_B_6akHVQl14_2;
	wire w_dff_B_T8q6GaV73_1;
	wire w_dff_B_ivK1VAAe2_2;
	wire w_dff_B_GLbQrpUB7_2;
	wire w_dff_B_xuHbWMUq0_2;
	wire w_dff_B_TMsJyuR51_2;
	wire w_dff_B_s0PbNZX80_2;
	wire w_dff_B_8Vj2Ag9v6_2;
	wire w_dff_B_iOK7Jftm4_2;
	wire w_dff_B_d7oiqQTm5_2;
	wire w_dff_B_tTqFB1lD5_2;
	wire w_dff_B_6PAKBTgy5_2;
	wire w_dff_B_39ySnxDb3_1;
	wire w_dff_B_OSuTQmLa3_2;
	wire w_dff_B_cWuLtvFd8_2;
	wire w_dff_B_p7ityrFI8_2;
	wire w_dff_B_RX3HDQs35_2;
	wire w_dff_B_hlA5x6yI2_2;
	wire w_dff_B_DL3pBouH4_2;
	wire w_dff_B_T1ih5VfZ8_2;
	wire w_dff_B_IYyZof909_2;
	wire w_dff_B_m2N89aZe5_1;
	wire w_dff_B_9NibFXlu7_2;
	wire w_dff_B_i5awPHmD6_2;
	wire w_dff_B_qUTHNux54_2;
	wire w_dff_B_3Qm1Dhu44_2;
	wire w_dff_B_oLzjGmyc2_2;
	wire w_dff_B_SzG0N2Y24_2;
	wire w_dff_B_wlQBLVKH0_2;
	wire w_dff_B_UipQ2Ew40_1;
	wire w_dff_B_W6KneUft4_1;
	wire w_dff_B_0mD8oNg82_1;
	wire w_dff_B_TCFaCcQC4_1;
	wire w_dff_B_Gdn853Jj8_0;
	wire w_dff_A_fWPG9oRP9_0;
	wire w_dff_A_LStzzifJ6_0;
	wire w_dff_B_VQ1qjIrd5_1;
	wire w_dff_B_VBFHxlXZ9_1;
	wire w_dff_A_jLjA2Bfy3_0;
	wire w_dff_A_UZaFVqwY3_1;
	wire w_dff_A_drno1gMW4_1;
	wire w_dff_A_cJO0RiS59_1;
	wire w_dff_A_HUDkCOMd1_1;
	wire w_dff_A_pJYFsnAs3_1;
	wire w_dff_A_G8IX5VBQ3_1;
	wire w_dff_B_qnSP67mV0_1;
	wire w_dff_A_FthOBBaS1_1;
	wire w_dff_B_6DV67CBU5_1;
	wire w_dff_B_dOGg3N0J9_2;
	wire w_dff_B_1BmlShjP1_2;
	wire w_dff_B_sBCdCDWn5_2;
	wire w_dff_B_6kVV8mKa3_2;
	wire w_dff_B_JagPo3q85_2;
	wire w_dff_B_QKmtHe0w6_2;
	wire w_dff_B_qnmEbv951_2;
	wire w_dff_B_VLBTxCBx4_2;
	wire w_dff_B_4hF8vQex5_2;
	wire w_dff_B_0wamdWPN2_2;
	wire w_dff_B_zGbEiIo27_2;
	wire w_dff_B_SJlWIMlT8_2;
	wire w_dff_B_ro1LDj600_2;
	wire w_dff_B_xn7xKFE13_2;
	wire w_dff_B_mSMf1meb0_2;
	wire w_dff_B_yLahuzfi4_2;
	wire w_dff_B_NItNMQwT1_2;
	wire w_dff_B_rNiRcqA04_2;
	wire w_dff_B_V0mWvfAB1_2;
	wire w_dff_B_e309RbpT0_2;
	wire w_dff_B_ZaQrucqD1_2;
	wire w_dff_B_Isvci4dc6_2;
	wire w_dff_B_PKbRrpm65_2;
	wire w_dff_B_fR9qGCHX3_2;
	wire w_dff_B_QmG4y5At7_2;
	wire w_dff_B_sGJlLfS49_2;
	wire w_dff_B_EUdTtewU4_2;
	wire w_dff_B_LCmBFyil5_2;
	wire w_dff_B_l3P6T8yE3_2;
	wire w_dff_B_Jp49Wk0u2_2;
	wire w_dff_B_RaOkfKwl2_2;
	wire w_dff_B_4fikkssd9_2;
	wire w_dff_B_lRKQxxSF5_2;
	wire w_dff_B_I2v5cY621_2;
	wire w_dff_B_pTGnd6c54_2;
	wire w_dff_B_TZr5F3Og9_2;
	wire w_dff_B_kR4OS3qD2_2;
	wire w_dff_B_EdX3cqby4_2;
	wire w_dff_B_MJBz7X6l3_2;
	wire w_dff_B_b5xB4cfa7_2;
	wire w_dff_B_sWLejboO0_2;
	wire w_dff_B_2il5fWCi4_1;
	wire w_dff_B_2OzbK2XA6_2;
	wire w_dff_B_EoCiPKBW8_2;
	wire w_dff_B_LwlA3ID82_2;
	wire w_dff_B_VMTBGKw68_2;
	wire w_dff_B_7hAYZ7a72_2;
	wire w_dff_B_xAbScloS1_2;
	wire w_dff_B_zgGxRnWB1_2;
	wire w_dff_B_Hf8Cv6NT2_2;
	wire w_dff_B_8mLDssmW5_2;
	wire w_dff_B_VbtoKRMe7_2;
	wire w_dff_B_vKNmCYuV2_2;
	wire w_dff_B_rJTmePHG6_2;
	wire w_dff_B_CEIZkxE79_2;
	wire w_dff_B_AHprEfiw6_2;
	wire w_dff_B_5gvjk9xL3_2;
	wire w_dff_B_1NRycjdP0_2;
	wire w_dff_B_x27BvJEP3_2;
	wire w_dff_B_ZYVl3Eh15_2;
	wire w_dff_B_1yn8CzxY3_2;
	wire w_dff_B_oyhNrCuN2_2;
	wire w_dff_B_MLqOKC2B5_2;
	wire w_dff_B_ELCuy6ku5_2;
	wire w_dff_B_t1mhuLBV3_2;
	wire w_dff_B_JsgnFewA9_2;
	wire w_dff_B_nqK2qD8L1_2;
	wire w_dff_B_9QxNETOY0_2;
	wire w_dff_B_HTZrj48d7_2;
	wire w_dff_B_8Db2viEg0_2;
	wire w_dff_B_vQSEPpxU1_2;
	wire w_dff_B_RHToYluM0_2;
	wire w_dff_B_e3zctTOZ1_2;
	wire w_dff_B_NObX8p2T4_2;
	wire w_dff_B_fnwMtLeA2_2;
	wire w_dff_B_9YwLMyqe9_2;
	wire w_dff_B_rFYf5rFh4_2;
	wire w_dff_B_cL5T4Ogy2_2;
	wire w_dff_B_3X9ysqiv8_2;
	wire w_dff_B_hmSzzKIG2_2;
	wire w_dff_B_xMcZA4CE3_1;
	wire w_dff_B_mf5Ueczm1_2;
	wire w_dff_B_GOvvzfQK0_2;
	wire w_dff_B_d4VJ3tOM3_2;
	wire w_dff_B_E3VU0BC40_2;
	wire w_dff_B_whJIcojK4_2;
	wire w_dff_B_jABkM8HR5_2;
	wire w_dff_B_nuBBTAud4_2;
	wire w_dff_B_SlEPmMjx0_2;
	wire w_dff_B_GjPHJlsT0_2;
	wire w_dff_B_kGrvL8tl5_2;
	wire w_dff_B_J9I9zmIs3_2;
	wire w_dff_B_Z8pmxG6x4_2;
	wire w_dff_B_3I2OLXAW5_2;
	wire w_dff_B_y2dODrBV9_2;
	wire w_dff_B_JycJK9A57_2;
	wire w_dff_B_skrfLLlq6_2;
	wire w_dff_B_KKwUwbUc9_2;
	wire w_dff_B_ls1dPspC9_2;
	wire w_dff_B_97ku6Fek6_2;
	wire w_dff_B_LtOycfXv9_2;
	wire w_dff_B_D7Tzzv8c7_2;
	wire w_dff_B_rQItFjMI2_2;
	wire w_dff_B_pKOH8t5A6_2;
	wire w_dff_B_BjEyFtRN9_2;
	wire w_dff_B_3KDamCFW5_2;
	wire w_dff_B_WpgIoqTT1_2;
	wire w_dff_B_98cckcgj2_2;
	wire w_dff_B_JKaAiQVz3_2;
	wire w_dff_B_OPgm1r9m1_2;
	wire w_dff_B_ptNdr2Sq4_2;
	wire w_dff_B_zABN6XwR5_2;
	wire w_dff_B_N0c5WKwz1_2;
	wire w_dff_B_eKkciStW7_2;
	wire w_dff_B_l2Pjn05G8_2;
	wire w_dff_B_OccyCEz61_2;
	wire w_dff_B_iOqyTgmz1_1;
	wire w_dff_B_YWYmBhFV4_2;
	wire w_dff_B_C5IuBdWk8_2;
	wire w_dff_B_yT3Ko8cJ6_2;
	wire w_dff_B_qp6htva55_2;
	wire w_dff_B_bvbiLwZA9_2;
	wire w_dff_B_poTebLeO3_2;
	wire w_dff_B_W7kih9lB0_2;
	wire w_dff_B_V9rExQbr4_2;
	wire w_dff_B_pRXZDnhe0_2;
	wire w_dff_B_agFrEuub0_2;
	wire w_dff_B_n9TI68tR3_2;
	wire w_dff_B_xjaRXSKH7_2;
	wire w_dff_B_9dIkEzHf6_2;
	wire w_dff_B_g1MTViux5_2;
	wire w_dff_B_d1yHmxSt4_2;
	wire w_dff_B_dreVPFfK2_2;
	wire w_dff_B_WpJs6XmR4_2;
	wire w_dff_B_aLm4x0ia2_2;
	wire w_dff_B_EZdMmF1q9_2;
	wire w_dff_B_bKkbuJZI2_2;
	wire w_dff_B_3VpGV4EA7_2;
	wire w_dff_B_qqSxGeDW7_2;
	wire w_dff_B_EqKbW2G49_2;
	wire w_dff_B_rcIcUfog5_2;
	wire w_dff_B_dCfeVtiP2_2;
	wire w_dff_B_5d7MW6cc9_2;
	wire w_dff_B_dLXWsxlb4_2;
	wire w_dff_B_Bm6amHFC5_2;
	wire w_dff_B_XaRubCkU3_2;
	wire w_dff_B_bgeYgFYi4_2;
	wire w_dff_B_fvvSlpHj4_2;
	wire w_dff_B_piK1THr49_2;
	wire w_dff_B_Nlcbd72D3_1;
	wire w_dff_B_2HPEFLM82_2;
	wire w_dff_B_vWr7eoBR6_2;
	wire w_dff_B_rg7FKUR23_2;
	wire w_dff_B_FApnZ9P93_2;
	wire w_dff_B_cUkMYVlJ3_2;
	wire w_dff_B_hDCcouWO2_2;
	wire w_dff_B_g61wtwJA1_2;
	wire w_dff_B_iicfxtvR4_2;
	wire w_dff_B_TaAUicxh6_2;
	wire w_dff_B_0qzNvZV34_2;
	wire w_dff_B_3omzJURq5_2;
	wire w_dff_B_pp4YLLXZ8_2;
	wire w_dff_B_xTuqZ6hU4_2;
	wire w_dff_B_q975WHsz1_2;
	wire w_dff_B_juriTZ5p0_2;
	wire w_dff_B_J1q0t3i26_2;
	wire w_dff_B_y6c4tBer9_2;
	wire w_dff_B_OAWuBNqb3_2;
	wire w_dff_B_VDzypX2G8_2;
	wire w_dff_B_Y4V0EiMH2_2;
	wire w_dff_B_KuJouY0T0_2;
	wire w_dff_B_YijVKpmQ0_2;
	wire w_dff_B_DomJE4z29_2;
	wire w_dff_B_1TZ6l6d11_2;
	wire w_dff_B_OnPlRJhm9_2;
	wire w_dff_B_tC22cMcN4_2;
	wire w_dff_B_5tLJTjaH8_2;
	wire w_dff_B_6DxEcXa09_2;
	wire w_dff_B_S34dDBt10_2;
	wire w_dff_B_zXMfh2tW4_1;
	wire w_dff_B_W7Dz1Qnz1_2;
	wire w_dff_B_DyLsH0OY5_2;
	wire w_dff_B_9mO2WHov3_2;
	wire w_dff_B_0bjRPH6k2_2;
	wire w_dff_B_sYUNCPeO4_2;
	wire w_dff_B_L4ykzywp6_2;
	wire w_dff_B_9VKWKBlF6_2;
	wire w_dff_B_n0VqNGXr2_2;
	wire w_dff_B_b7cB2ACx8_2;
	wire w_dff_B_mEo84peu1_2;
	wire w_dff_B_sr8ONZMh7_2;
	wire w_dff_B_hDD2sypM9_2;
	wire w_dff_B_4uzQCgt64_2;
	wire w_dff_B_Gjn9kFKJ0_2;
	wire w_dff_B_DTUizuuB1_2;
	wire w_dff_B_1rBTGPXP2_2;
	wire w_dff_B_c2ds4AcS7_2;
	wire w_dff_B_LVOKVTvM5_2;
	wire w_dff_B_7r2ABg1S5_2;
	wire w_dff_B_e1qQgB797_2;
	wire w_dff_B_GbTO9bFl8_2;
	wire w_dff_B_gEukhRpQ0_2;
	wire w_dff_B_Osy9HHTE8_2;
	wire w_dff_B_NJ0E4Suu2_2;
	wire w_dff_B_q9yyD1qM7_2;
	wire w_dff_B_Ym1N6bAQ5_2;
	wire w_dff_B_aqaLGXOT4_1;
	wire w_dff_B_oQd8Drrb6_2;
	wire w_dff_B_TgUPBvNo2_2;
	wire w_dff_B_hGutAvSs1_2;
	wire w_dff_B_dHnHjPAi6_2;
	wire w_dff_B_fdXZGFd91_2;
	wire w_dff_B_aCBknWDn7_2;
	wire w_dff_B_aRnaJa3d3_2;
	wire w_dff_B_SVsWrV5Y1_2;
	wire w_dff_B_mXgxtTEs9_2;
	wire w_dff_B_3LXiQ8wr5_2;
	wire w_dff_B_ZCPFiMjh8_2;
	wire w_dff_B_JupzjdSE7_2;
	wire w_dff_B_vwvwWmfs9_2;
	wire w_dff_B_d83LMinm0_2;
	wire w_dff_B_PT7qa8pG9_2;
	wire w_dff_B_5rfZzXRl7_2;
	wire w_dff_B_K5UsvlC36_2;
	wire w_dff_B_jN0B3Hg38_2;
	wire w_dff_B_bMWuoRQU1_2;
	wire w_dff_B_08CLUnav2_2;
	wire w_dff_B_fGMlVNJy1_2;
	wire w_dff_B_Mn7l1HXh8_2;
	wire w_dff_B_PRIeYDNt5_2;
	wire w_dff_B_kdxQH1hD6_1;
	wire w_dff_B_HCzYG60k7_2;
	wire w_dff_B_5hBk78Fa0_2;
	wire w_dff_B_D6HNnkBD1_2;
	wire w_dff_B_aUJ5hsqJ0_2;
	wire w_dff_B_eOtt4UFf4_2;
	wire w_dff_B_LHW0FfEu0_2;
	wire w_dff_B_mWpSzgvl5_2;
	wire w_dff_B_ElZNEvgM4_2;
	wire w_dff_B_SKg6nO6k2_2;
	wire w_dff_B_xaUDYiJt9_2;
	wire w_dff_B_ZLUP5LaM9_2;
	wire w_dff_B_NeEBMxcE6_2;
	wire w_dff_B_ydTr7wtZ0_2;
	wire w_dff_B_osMTjY5i1_2;
	wire w_dff_B_AffJraA94_2;
	wire w_dff_B_Z7dk3cDU5_2;
	wire w_dff_B_UubY8gNc7_2;
	wire w_dff_B_RXBU1v445_2;
	wire w_dff_B_fnGQfLsP3_2;
	wire w_dff_B_UslNWrpR7_2;
	wire w_dff_B_r7ZG6dqT3_1;
	wire w_dff_B_k6mxmWdS7_2;
	wire w_dff_B_5WVxsyCe5_2;
	wire w_dff_B_KCYjFm1k4_2;
	wire w_dff_B_6jMRu9FB5_2;
	wire w_dff_B_YS6iORA66_2;
	wire w_dff_B_P0Oa2pEG1_2;
	wire w_dff_B_oCnCQZlL4_2;
	wire w_dff_B_AMQ7jfWC0_2;
	wire w_dff_B_1RTishND9_2;
	wire w_dff_B_IwRWwSvu9_2;
	wire w_dff_B_k5bhNNs23_2;
	wire w_dff_B_A97wTBuN9_2;
	wire w_dff_B_ENSOQdib9_2;
	wire w_dff_B_WNh5RNnA5_2;
	wire w_dff_B_a5XXBoSe0_2;
	wire w_dff_B_ai4SvB5g3_2;
	wire w_dff_B_Nz2nYbTU5_2;
	wire w_dff_B_KMgHgW2O2_1;
	wire w_dff_B_QMurNLlQ7_2;
	wire w_dff_B_dzC7afe74_2;
	wire w_dff_B_B2Mgau256_2;
	wire w_dff_B_a8E0En2V6_2;
	wire w_dff_B_TzQJEmA32_2;
	wire w_dff_B_DGDETqys6_2;
	wire w_dff_B_NDSInMWX4_2;
	wire w_dff_B_h9CZyYT61_2;
	wire w_dff_B_CusKAVL52_2;
	wire w_dff_B_QxyJPTha4_2;
	wire w_dff_B_rDtdTpkI3_2;
	wire w_dff_B_yIey17ab9_2;
	wire w_dff_B_4efL7dCV5_2;
	wire w_dff_B_HU2GbyaZ7_2;
	wire w_dff_B_YI5hYO794_1;
	wire w_dff_B_4uwK1ZRk4_2;
	wire w_dff_B_z2oclxAG8_2;
	wire w_dff_B_yU3poFZb5_2;
	wire w_dff_B_5aowa2yR4_2;
	wire w_dff_B_vqkZb6233_2;
	wire w_dff_B_DwLfJLt02_2;
	wire w_dff_B_OmpSV0WB2_2;
	wire w_dff_B_AOzvZOFq4_2;
	wire w_dff_B_F4IlZSsO1_2;
	wire w_dff_B_06ARLHTF0_2;
	wire w_dff_B_0FF0RhK38_1;
	wire w_dff_B_1PVUAIIw9_2;
	wire w_dff_B_JQXRx6Ps8_2;
	wire w_dff_B_JjBpuBFH5_2;
	wire w_dff_B_hgv5c3tx9_2;
	wire w_dff_B_cRdn1g5B0_2;
	wire w_dff_B_eMgF42nM1_2;
	wire w_dff_B_DRvW5Fr76_2;
	wire w_dff_B_Zhi0614O5_2;
	wire w_dff_B_pITryFcZ5_1;
	wire w_dff_B_oXpog3fo0_2;
	wire w_dff_B_CODLarTi9_2;
	wire w_dff_B_GwxsGOQE2_2;
	wire w_dff_B_nzZv25Aw9_2;
	wire w_dff_B_Y1X9YCny9_2;
	wire w_dff_B_zeb0jvwG4_2;
	wire w_dff_B_GAMWtoFq2_2;
	wire w_dff_B_K5V2KHjU3_1;
	wire w_dff_B_wuGYaRmU8_1;
	wire w_dff_B_e5I1tcpN9_1;
	wire w_dff_B_WYYKT4UZ3_1;
	wire w_dff_B_D6eKyeyl8_0;
	wire w_dff_A_8ydGlACv3_0;
	wire w_dff_A_3m1VZbBZ2_0;
	wire w_dff_B_LyhL8Snl8_1;
	wire w_dff_B_YuHExj7R4_1;
	wire w_dff_A_48Fakt9R8_0;
	wire w_dff_A_yBVmxsN03_1;
	wire w_dff_A_1dokVTgx8_1;
	wire w_dff_A_i9qFOE6m4_1;
	wire w_dff_A_oQuvQBQq3_1;
	wire w_dff_A_EKgaLSVg7_1;
	wire w_dff_A_Kcc6bB7L1_1;
	wire w_dff_B_BIrgQ7AT7_1;
	wire w_dff_A_ssrXAKtQ0_1;
	wire w_dff_B_BXjl0G2O6_1;
	wire w_dff_B_lrFDyZ1k0_2;
	wire w_dff_B_smNHENwB4_2;
	wire w_dff_B_JHIdWpMv9_2;
	wire w_dff_B_WIShTbn59_2;
	wire w_dff_B_BgYXh6C66_2;
	wire w_dff_B_cUPdgFNU6_2;
	wire w_dff_B_VrUDwbX50_2;
	wire w_dff_B_U7BrJy915_2;
	wire w_dff_B_aF5daw8L6_2;
	wire w_dff_B_wyIyIqkM5_2;
	wire w_dff_B_3AnMBDNf9_2;
	wire w_dff_B_LBUE0QMh1_2;
	wire w_dff_B_wg6jI9769_2;
	wire w_dff_B_6ma86CHJ5_2;
	wire w_dff_B_QJhBV3h86_2;
	wire w_dff_B_RGHXScO50_2;
	wire w_dff_B_cZEYKMmO0_2;
	wire w_dff_B_DI1ZpD6Q3_2;
	wire w_dff_B_NkZ1EQx12_2;
	wire w_dff_B_aCHysf9u8_2;
	wire w_dff_B_XUzEbjbv4_2;
	wire w_dff_B_f3RHJg6j9_2;
	wire w_dff_B_UKlDCxib4_2;
	wire w_dff_B_tp7oMU3c0_2;
	wire w_dff_B_JIMLoSuW5_2;
	wire w_dff_B_x1k2WNq90_2;
	wire w_dff_B_fl0uf7fw8_2;
	wire w_dff_B_YM43M1rB6_2;
	wire w_dff_B_AZIfTLcq8_2;
	wire w_dff_B_KfcAI0Al0_2;
	wire w_dff_B_Wi7Nfyqe5_2;
	wire w_dff_B_JQGzFj0b1_2;
	wire w_dff_B_AxRDFDkS5_2;
	wire w_dff_B_qxyz7S7d4_2;
	wire w_dff_B_I5ASGsY29_2;
	wire w_dff_B_7eEp03fZ0_2;
	wire w_dff_B_gbZtysXo3_2;
	wire w_dff_B_n29bydAO2_2;
	wire w_dff_B_5048nYaS6_2;
	wire w_dff_B_0oiRhCew3_2;
	wire w_dff_B_XLEbZbGh4_2;
	wire w_dff_B_dAbLNxEq4_2;
	wire w_dff_B_PMZFNPI94_1;
	wire w_dff_B_DebyrMO77_2;
	wire w_dff_B_r8H7Kio31_2;
	wire w_dff_B_T2MKbseA9_2;
	wire w_dff_B_2iTkIsY93_2;
	wire w_dff_B_YHqQGlAz1_2;
	wire w_dff_B_pN5nbpjh8_2;
	wire w_dff_B_dYO5KS5O0_2;
	wire w_dff_B_Y8RYzSaX6_2;
	wire w_dff_B_uKw0ccgk4_2;
	wire w_dff_B_Z0Qxccvj0_2;
	wire w_dff_B_A0kbsgkX3_2;
	wire w_dff_B_qXl1i2G03_2;
	wire w_dff_B_xtNOEPbD4_2;
	wire w_dff_B_6iUx3StV5_2;
	wire w_dff_B_kumXx7DD7_2;
	wire w_dff_B_cU4ceoFc0_2;
	wire w_dff_B_shnmPZuQ9_2;
	wire w_dff_B_8xukIEZj5_2;
	wire w_dff_B_zx79VxaU5_2;
	wire w_dff_B_BJnagulE2_2;
	wire w_dff_B_RAPl8noj9_2;
	wire w_dff_B_RGUU8MWp9_2;
	wire w_dff_B_wGb0rXKg5_2;
	wire w_dff_B_VaCAp1wr0_2;
	wire w_dff_B_QG55KrUk7_2;
	wire w_dff_B_NDvpUEeQ2_2;
	wire w_dff_B_dm8KWOiU1_2;
	wire w_dff_B_p4d5zdTR9_2;
	wire w_dff_B_OBe0MAmH4_2;
	wire w_dff_B_B2EeaBhy3_2;
	wire w_dff_B_68Q8aHDQ7_2;
	wire w_dff_B_0WmD325C5_2;
	wire w_dff_B_IbqKD7kx4_2;
	wire w_dff_B_qK3gEvZR7_2;
	wire w_dff_B_MWkfWstk4_2;
	wire w_dff_B_FHrD2GwZ3_2;
	wire w_dff_B_S3idry3O1_2;
	wire w_dff_B_Onv7pv8s0_2;
	wire w_dff_B_D8AJXiMT8_2;
	wire w_dff_B_iuLwvLhL0_1;
	wire w_dff_B_hWsSLFhh0_2;
	wire w_dff_B_DnIzzPtW1_2;
	wire w_dff_B_MAOfJYIF0_2;
	wire w_dff_B_4PXKLdAN8_2;
	wire w_dff_B_LelS9Q6e1_2;
	wire w_dff_B_qlqGLVOQ4_2;
	wire w_dff_B_gk81zt5a9_2;
	wire w_dff_B_DkTaDtrc2_2;
	wire w_dff_B_BjEHUZ0o7_2;
	wire w_dff_B_i7LghEmm7_2;
	wire w_dff_B_rASNtBbA4_2;
	wire w_dff_B_OXFzaDa63_2;
	wire w_dff_B_LzKClCU40_2;
	wire w_dff_B_V4hBBEHr7_2;
	wire w_dff_B_sTsrNt3r3_2;
	wire w_dff_B_3fmE2yMf3_2;
	wire w_dff_B_HHQlUgVJ6_2;
	wire w_dff_B_St80496l2_2;
	wire w_dff_B_N4dfAHcJ7_2;
	wire w_dff_B_87HrfKX45_2;
	wire w_dff_B_JvZ0hTq43_2;
	wire w_dff_B_9JYQMTnW0_2;
	wire w_dff_B_HxcPrKRJ7_2;
	wire w_dff_B_mgRs9CGs9_2;
	wire w_dff_B_P9uCtLmh5_2;
	wire w_dff_B_cf0LEYy75_2;
	wire w_dff_B_6agVIGVX2_2;
	wire w_dff_B_Jx1P4F5i3_2;
	wire w_dff_B_k0fY72Uo3_2;
	wire w_dff_B_0i2aVSqO7_2;
	wire w_dff_B_fDFBxM5M8_2;
	wire w_dff_B_0P0nXKC87_2;
	wire w_dff_B_OcMrzMJL0_2;
	wire w_dff_B_4dq6X5jt7_2;
	wire w_dff_B_koax4oEL4_2;
	wire w_dff_B_kVKZu0VS8_2;
	wire w_dff_B_OwlYxgy72_1;
	wire w_dff_B_YMBcjPwl9_2;
	wire w_dff_B_B8rzKxcG1_2;
	wire w_dff_B_kcvzjtW91_2;
	wire w_dff_B_NGdXoPSC2_2;
	wire w_dff_B_ARNEuVDF2_2;
	wire w_dff_B_PNtMEDB15_2;
	wire w_dff_B_ac8QHhHG9_2;
	wire w_dff_B_DenZcyew2_2;
	wire w_dff_B_2cmKzP9h9_2;
	wire w_dff_B_zpyZy9Pa1_2;
	wire w_dff_B_xN4SmyIw9_2;
	wire w_dff_B_tQDyDHsC8_2;
	wire w_dff_B_DX0hPpvt7_2;
	wire w_dff_B_AI89dD9b4_2;
	wire w_dff_B_VNHZRxGO7_2;
	wire w_dff_B_z73vebUl3_2;
	wire w_dff_B_FlR1b3v91_2;
	wire w_dff_B_C8Iyb30f4_2;
	wire w_dff_B_kRxTDog36_2;
	wire w_dff_B_xG2ummhN6_2;
	wire w_dff_B_MBRnurS83_2;
	wire w_dff_B_xEkF9KEu3_2;
	wire w_dff_B_8sVaR9KL3_2;
	wire w_dff_B_JPJPO1043_2;
	wire w_dff_B_m9RY8Fbk3_2;
	wire w_dff_B_fcggUJ4O9_2;
	wire w_dff_B_yMOlkVNp5_2;
	wire w_dff_B_WWJuFx5f1_2;
	wire w_dff_B_ZbN0Ldhk4_2;
	wire w_dff_B_SCoxlTjY5_2;
	wire w_dff_B_Eb1LTRxI1_2;
	wire w_dff_B_daRlOphW0_2;
	wire w_dff_B_ZpOkK2qv5_2;
	wire w_dff_B_1zuIz7yN8_1;
	wire w_dff_B_Y9x2XN5C0_2;
	wire w_dff_B_wNIUAWUZ8_2;
	wire w_dff_B_Xu0OmIFH4_2;
	wire w_dff_B_DoZ7r9cc7_2;
	wire w_dff_B_DaC3ZOD30_2;
	wire w_dff_B_paMlMcmN3_2;
	wire w_dff_B_GaWb72g51_2;
	wire w_dff_B_TQ3OeISQ2_2;
	wire w_dff_B_uyOB9opk5_2;
	wire w_dff_B_kt6U1X2Q9_2;
	wire w_dff_B_NkYhfIoO5_2;
	wire w_dff_B_1rkvjoJp5_2;
	wire w_dff_B_2LmFrbWc1_2;
	wire w_dff_B_4n4reUpB0_2;
	wire w_dff_B_z83Qssm48_2;
	wire w_dff_B_Z9bjJAQq1_2;
	wire w_dff_B_r1vj7Apr4_2;
	wire w_dff_B_Dji2Auff5_2;
	wire w_dff_B_NvckqNtQ5_2;
	wire w_dff_B_TtPObzDc2_2;
	wire w_dff_B_615mHX7N8_2;
	wire w_dff_B_vDDfV8HK2_2;
	wire w_dff_B_UGbJX35k1_2;
	wire w_dff_B_lCaQomBp7_2;
	wire w_dff_B_WQZhWyPd8_2;
	wire w_dff_B_TyxjQAWM3_2;
	wire w_dff_B_GJlJgzFq8_2;
	wire w_dff_B_mrLY5sBn8_2;
	wire w_dff_B_mrZXleBf5_2;
	wire w_dff_B_TQ1Z6noW7_2;
	wire w_dff_B_t7lINx934_1;
	wire w_dff_B_BE4QdvDD6_2;
	wire w_dff_B_niA3mLEb2_2;
	wire w_dff_B_gshMcPLK1_2;
	wire w_dff_B_vW6fWiFr4_2;
	wire w_dff_B_phyljEV00_2;
	wire w_dff_B_WqnUaDZj3_2;
	wire w_dff_B_jViUbaNz1_2;
	wire w_dff_B_MZAUlxvx0_2;
	wire w_dff_B_V8xbDkFG8_2;
	wire w_dff_B_YEjHdRFj9_2;
	wire w_dff_B_Sx14C7uq7_2;
	wire w_dff_B_yWqDNBmV3_2;
	wire w_dff_B_kgsShTQa1_2;
	wire w_dff_B_AS5IVjcG7_2;
	wire w_dff_B_FDJxEl4k1_2;
	wire w_dff_B_ySZUNYfa5_2;
	wire w_dff_B_N1OZ2zrm9_2;
	wire w_dff_B_AYiIzIG12_2;
	wire w_dff_B_QrL7BOrv2_2;
	wire w_dff_B_9yzo2Y6g2_2;
	wire w_dff_B_UtyAaVIM3_2;
	wire w_dff_B_i1BQQSYZ2_2;
	wire w_dff_B_CdAax9ul5_2;
	wire w_dff_B_MxQTAqAG3_2;
	wire w_dff_B_9iXyJA0Q8_2;
	wire w_dff_B_SL4sG0kr9_2;
	wire w_dff_B_JTtRBhye0_2;
	wire w_dff_B_6dviGXV86_1;
	wire w_dff_B_ndH1q0i26_2;
	wire w_dff_B_PVQabe368_2;
	wire w_dff_B_UGg0x5Dn0_2;
	wire w_dff_B_CoSon9c16_2;
	wire w_dff_B_g1BDn8Lx0_2;
	wire w_dff_B_1z3AD6Fn0_2;
	wire w_dff_B_hUymP6L81_2;
	wire w_dff_B_EZTkmud71_2;
	wire w_dff_B_NktW4f2W6_2;
	wire w_dff_B_OOseTLPn8_2;
	wire w_dff_B_Eq5VuKmS1_2;
	wire w_dff_B_UNQtDASk7_2;
	wire w_dff_B_dXBavHkH6_2;
	wire w_dff_B_AnI7U8vz6_2;
	wire w_dff_B_A28RxnFs2_2;
	wire w_dff_B_tYL0F2Yq5_2;
	wire w_dff_B_VqemReL51_2;
	wire w_dff_B_FzuQiHV79_2;
	wire w_dff_B_2qdNOR3u9_2;
	wire w_dff_B_92o2sBoo8_2;
	wire w_dff_B_T9MeuH202_2;
	wire w_dff_B_kViNAkG78_2;
	wire w_dff_B_jMrDNSe89_2;
	wire w_dff_B_2McmDv8G7_2;
	wire w_dff_B_sh0dxksO2_1;
	wire w_dff_B_hC7BbIqV6_2;
	wire w_dff_B_oYRgShH11_2;
	wire w_dff_B_ZlJNZeT99_2;
	wire w_dff_B_qL4Ht7TW1_2;
	wire w_dff_B_EW52QgG49_2;
	wire w_dff_B_1LHCHdbr8_2;
	wire w_dff_B_4OjnTwQM1_2;
	wire w_dff_B_6aZBglVu5_2;
	wire w_dff_B_QUGtxAtR7_2;
	wire w_dff_B_cxL7swVY5_2;
	wire w_dff_B_OaGEaaHd2_2;
	wire w_dff_B_l6lFYMIb9_2;
	wire w_dff_B_8Lbq6cW45_2;
	wire w_dff_B_oXRt8b9B3_2;
	wire w_dff_B_sKIJYoAd3_2;
	wire w_dff_B_xL29oZzT0_2;
	wire w_dff_B_vSw9KwCM8_2;
	wire w_dff_B_nlQCxk901_2;
	wire w_dff_B_lwUCygxZ2_2;
	wire w_dff_B_iQXQbdJt5_2;
	wire w_dff_B_A0i2702a4_2;
	wire w_dff_B_INKymOYR8_1;
	wire w_dff_B_FTtdPVNL9_2;
	wire w_dff_B_SW6PhlFB7_2;
	wire w_dff_B_YgO8e70f1_2;
	wire w_dff_B_onAbcYUi9_2;
	wire w_dff_B_n3B9ZFsg5_2;
	wire w_dff_B_vp9uWi3d5_2;
	wire w_dff_B_vYbHpcV62_2;
	wire w_dff_B_4abRs4b61_2;
	wire w_dff_B_gOhZxzpu8_2;
	wire w_dff_B_N0AxYhOr4_2;
	wire w_dff_B_AzAl7yhO4_2;
	wire w_dff_B_M9jz9D8i7_2;
	wire w_dff_B_okAosbHv2_2;
	wire w_dff_B_7dBtRMgy3_2;
	wire w_dff_B_JcemjKhx5_2;
	wire w_dff_B_CRpi4ucq3_2;
	wire w_dff_B_cVNuB1795_2;
	wire w_dff_B_Lbwdgh9C9_2;
	wire w_dff_B_1n21AahF4_1;
	wire w_dff_B_wA9s5U9U5_2;
	wire w_dff_B_VIomQFwF3_2;
	wire w_dff_B_eiPr1zSx8_2;
	wire w_dff_B_6W9kCZei4_2;
	wire w_dff_B_FNUWosxc9_2;
	wire w_dff_B_OVy8mKHP4_2;
	wire w_dff_B_I23sPtR88_2;
	wire w_dff_B_UHnAMCwM8_2;
	wire w_dff_B_cItW43000_2;
	wire w_dff_B_bophiV9U5_2;
	wire w_dff_B_C0lRuRsc7_2;
	wire w_dff_B_6PEiuxw30_2;
	wire w_dff_B_63ir5bPq7_2;
	wire w_dff_B_fCsW9NnO7_2;
	wire w_dff_B_xUKLDhg11_2;
	wire w_dff_B_ztUuxrZa4_1;
	wire w_dff_B_SOjC0u682_2;
	wire w_dff_B_ZRFRRR0f1_2;
	wire w_dff_B_Lj2Y2oRF3_2;
	wire w_dff_B_fE61N04S1_2;
	wire w_dff_B_64dfNbLk6_2;
	wire w_dff_B_wlaoX3Vr8_2;
	wire w_dff_B_dfIJjtkb1_2;
	wire w_dff_B_tdHgasEH1_2;
	wire w_dff_B_FuOHYAuB3_2;
	wire w_dff_B_BrurOUzU1_2;
	wire w_dff_B_dnvH4RRW9_2;
	wire w_dff_B_bqJrps8C6_2;
	wire w_dff_B_CaNGttoo6_1;
	wire w_dff_B_AhgYcDTj0_2;
	wire w_dff_B_rWqLJzx34_2;
	wire w_dff_B_bVPYrA530_2;
	wire w_dff_B_HrkcjwoK6_2;
	wire w_dff_B_NJAO925O7_2;
	wire w_dff_B_GLmoDkf79_2;
	wire w_dff_B_eK7IfPZD4_2;
	wire w_dff_B_ixfXDMSX9_2;
	wire w_dff_B_VArijCD09_1;
	wire w_dff_B_0stsqYTI2_2;
	wire w_dff_B_LsfBhqdJ8_2;
	wire w_dff_B_IijG6F663_2;
	wire w_dff_B_gKXg3xrd9_2;
	wire w_dff_B_ytyWzPSK7_2;
	wire w_dff_B_hzNvwo292_2;
	wire w_dff_B_E2ffu9kh8_2;
	wire w_dff_B_kSwT1ifs9_1;
	wire w_dff_B_P3tf2sQs7_1;
	wire w_dff_B_VtnTitoD4_1;
	wire w_dff_B_VI7ITJyG6_1;
	wire w_dff_B_LuvGROLa3_0;
	wire w_dff_A_CUC1p7iX4_0;
	wire w_dff_A_BmmRQH6Y3_0;
	wire w_dff_B_Qoe4saXY8_1;
	wire w_dff_B_3R5BpVwG3_1;
	wire w_dff_A_rwZL9Mh59_0;
	wire w_dff_A_gPAIF4546_1;
	wire w_dff_A_MD2z5eFk2_1;
	wire w_dff_A_h7Ops2wC3_1;
	wire w_dff_A_IXjrD1I14_1;
	wire w_dff_A_Ot93eFkq0_1;
	wire w_dff_A_5nlEOUCZ1_1;
	wire w_dff_B_6dBjoyOm3_1;
	wire w_dff_B_aM5YUJHk4_1;
	wire w_dff_B_SGXXBPc45_1;
	wire w_dff_B_BcDV6mNw2_2;
	wire w_dff_B_1bGpGl5T7_2;
	wire w_dff_B_JnPmFYrf7_2;
	wire w_dff_B_ropxEmUA2_2;
	wire w_dff_B_2OdIL9367_2;
	wire w_dff_B_d6B8937O8_2;
	wire w_dff_B_vKfDsliz8_2;
	wire w_dff_B_XcEDky1r8_2;
	wire w_dff_B_D6fCJt7M3_2;
	wire w_dff_B_mQNvpyys1_2;
	wire w_dff_B_T45uRn0Q2_2;
	wire w_dff_B_rVZYlN1W7_2;
	wire w_dff_B_bKvcE4Fa9_2;
	wire w_dff_B_GC62llFU5_2;
	wire w_dff_B_6GOFvHpE6_2;
	wire w_dff_B_i5uokXZK0_2;
	wire w_dff_B_kaD8yBEQ8_2;
	wire w_dff_B_piSWNuxY6_2;
	wire w_dff_B_oFjfjcPQ5_2;
	wire w_dff_B_XIgxF0Qb7_2;
	wire w_dff_B_ZdpmQgW77_2;
	wire w_dff_B_VxsFvM9j3_2;
	wire w_dff_B_uIshidnJ9_2;
	wire w_dff_B_6EoNLDxg7_2;
	wire w_dff_B_itKKYmfu5_2;
	wire w_dff_B_26b8Wul84_2;
	wire w_dff_B_6fE9XqV78_2;
	wire w_dff_B_YvjkNsXh7_2;
	wire w_dff_B_P5Ytl9pq7_2;
	wire w_dff_B_49fqIaC37_2;
	wire w_dff_B_xwUtf7Xf2_2;
	wire w_dff_B_IA96D6sB8_2;
	wire w_dff_B_VTBg1lRU0_2;
	wire w_dff_B_JvHpUeeM8_2;
	wire w_dff_B_zCecaY1t8_2;
	wire w_dff_B_YFnOXOHD5_2;
	wire w_dff_B_H9hyc7C43_2;
	wire w_dff_B_hRj2FXJl2_2;
	wire w_dff_B_6tLBjBwn8_2;
	wire w_dff_B_SBglLqPa8_2;
	wire w_dff_B_gBHmUP9A7_2;
	wire w_dff_B_NK1gJBzJ7_2;
	wire w_dff_B_TMxCXRkN4_2;
	wire w_dff_B_4Fb7TyHm6_2;
	wire w_dff_B_4wxreOQc8_2;
	wire w_dff_B_W0A5pr7J2_2;
	wire w_dff_B_iMa9E4bR5_2;
	wire w_dff_B_pRCzIX9F5_2;
	wire w_dff_B_7Xf3GiM45_2;
	wire w_dff_B_HebX0F8X0_2;
	wire w_dff_B_nMM7Ej3k3_2;
	wire w_dff_B_HtVg4BPT0_2;
	wire w_dff_B_R35mousA7_2;
	wire w_dff_B_ZYuOm7OY3_2;
	wire w_dff_B_cioyhJK83_2;
	wire w_dff_B_elFtxs0Y6_2;
	wire w_dff_B_p9cx9ORI7_2;
	wire w_dff_B_iayFpKPe8_2;
	wire w_dff_B_d5WzPutg1_2;
	wire w_dff_B_v4QTKvHN8_2;
	wire w_dff_B_vPkN0wTH5_2;
	wire w_dff_B_xp4wdqk08_2;
	wire w_dff_B_kHzcuWf18_2;
	wire w_dff_B_jpK13zcP3_2;
	wire w_dff_B_pLF0hSJ70_2;
	wire w_dff_B_O1UkgqKR0_2;
	wire w_dff_B_lTfHWvH69_2;
	wire w_dff_B_g1daqpg70_2;
	wire w_dff_B_EBX5IZm07_2;
	wire w_dff_B_2k4ldK4S1_2;
	wire w_dff_B_hFVTBlBT9_2;
	wire w_dff_B_Qfs7R1rE8_2;
	wire w_dff_B_RCNwG5CY5_2;
	wire w_dff_B_SbH6XqLT6_2;
	wire w_dff_B_ewLWYV3L8_2;
	wire w_dff_B_sSTI7Un12_2;
	wire w_dff_B_a2c98eeB3_2;
	wire w_dff_B_XuSnMPXR4_2;
	wire w_dff_B_v3ORR4x87_2;
	wire w_dff_B_aBYn8zWe1_2;
	wire w_dff_B_RsaprTqE6_2;
	wire w_dff_B_FrYpMJtv9_2;
	wire w_dff_B_7Obk5NuS3_2;
	wire w_dff_B_xdHqNUEm5_2;
	wire w_dff_B_0P9RNZtB5_2;
	wire w_dff_B_zHkCpcXH2_2;
	wire w_dff_A_tVLqk79Y1_1;
	wire w_dff_B_zqUqH8KZ3_1;
	wire w_dff_B_RhWltqDJ3_2;
	wire w_dff_B_CnBM2kD77_2;
	wire w_dff_B_IzhKd0yn0_2;
	wire w_dff_B_XU4O6faH4_2;
	wire w_dff_B_El91niX44_2;
	wire w_dff_B_CxA3bteM8_2;
	wire w_dff_B_FdnckxMr0_2;
	wire w_dff_B_twRzAU7V4_2;
	wire w_dff_B_HEFT2mGk1_2;
	wire w_dff_B_B3WgssQZ3_2;
	wire w_dff_B_8hpJyFHe5_2;
	wire w_dff_B_34vZx5tq6_2;
	wire w_dff_B_LjR792se1_2;
	wire w_dff_B_72iKWtpb5_2;
	wire w_dff_B_rMNZlLd74_2;
	wire w_dff_B_hvEvsA8i0_2;
	wire w_dff_B_HCkalJ7L2_2;
	wire w_dff_B_Sg7lhnNc7_2;
	wire w_dff_B_dJImzno93_2;
	wire w_dff_B_vKb5FWI98_2;
	wire w_dff_B_P1kVvgXl4_2;
	wire w_dff_B_gM3Jqd4j5_2;
	wire w_dff_B_xb7wssoE8_2;
	wire w_dff_B_keaVsMcq6_2;
	wire w_dff_B_bMeNLmQj6_2;
	wire w_dff_B_ZHLi5hij9_2;
	wire w_dff_B_GekzxAFp3_2;
	wire w_dff_B_HS7poe923_2;
	wire w_dff_B_M7cw7VQS9_2;
	wire w_dff_B_IitJrHY92_2;
	wire w_dff_B_MV9rd15C1_2;
	wire w_dff_B_Xp0vBTyE8_2;
	wire w_dff_B_9c6zEnAY6_2;
	wire w_dff_B_wzbll3z81_2;
	wire w_dff_B_qBw5QAhP3_2;
	wire w_dff_B_a7HoWehd0_2;
	wire w_dff_B_ps2IY3dJ6_2;
	wire w_dff_B_mG6nYk3B3_2;
	wire w_dff_B_tztcrnI39_2;
	wire w_dff_B_ioHryxFd7_2;
	wire w_dff_B_Z7awHPYz3_2;
	wire w_dff_B_gDyZj84K6_2;
	wire w_dff_B_1Jwqxdfo2_1;
	wire w_dff_B_phKCi7S75_1;
	wire w_dff_B_tblBrehd0_2;
	wire w_dff_B_itSFHr903_2;
	wire w_dff_B_b4lFKQdd9_2;
	wire w_dff_B_EnfK4HhG4_2;
	wire w_dff_B_MBKDZO3U1_2;
	wire w_dff_B_P8wlmhnz0_2;
	wire w_dff_B_QHhqZK2W6_2;
	wire w_dff_B_ko7SEAmP5_2;
	wire w_dff_B_b9vnJDJZ6_2;
	wire w_dff_B_7xP3nVcU0_2;
	wire w_dff_B_M9E2UCpg2_2;
	wire w_dff_B_rYoCC4SL4_2;
	wire w_dff_B_0TIE7HMF9_2;
	wire w_dff_B_k06ZKsXd1_2;
	wire w_dff_B_WlkIrWxy0_2;
	wire w_dff_B_orkWzp2v5_2;
	wire w_dff_B_YvDgYskx9_2;
	wire w_dff_B_Li9pWwx11_2;
	wire w_dff_B_dpQ1y37P8_2;
	wire w_dff_B_4Kqvo8Qx4_2;
	wire w_dff_B_chCfoMZa5_2;
	wire w_dff_B_sDyJGmHR4_2;
	wire w_dff_B_iCgeaUcJ4_2;
	wire w_dff_B_3YQhtyL10_2;
	wire w_dff_B_1d5XGaJf0_2;
	wire w_dff_B_xG0VBjjW4_2;
	wire w_dff_B_8qLdaMuI1_2;
	wire w_dff_B_tNLsAqB68_2;
	wire w_dff_B_JHPb6ycA3_2;
	wire w_dff_B_hhgj1rXA4_2;
	wire w_dff_B_aJE1NL4l2_2;
	wire w_dff_B_5wSGGqLT0_2;
	wire w_dff_B_KjWQhbJj2_2;
	wire w_dff_B_Li6AQjSy2_2;
	wire w_dff_B_aDwAbSO98_2;
	wire w_dff_B_qKjbUunT4_2;
	wire w_dff_B_KgVcwmGA5_2;
	wire w_dff_B_IWPsV1KB9_2;
	wire w_dff_B_mdap9Y3v1_2;
	wire w_dff_B_ZbH0ly908_2;
	wire w_dff_B_G79aM3YV9_2;
	wire w_dff_B_6CMoaR1y9_2;
	wire w_dff_B_JcSzmsje1_2;
	wire w_dff_B_C5ETVcMd9_2;
	wire w_dff_B_WTu8ztxl0_2;
	wire w_dff_B_lOzQHJi20_2;
	wire w_dff_B_9MtAWHBZ1_2;
	wire w_dff_B_fkX8zeqN4_2;
	wire w_dff_B_5GRe2zu69_2;
	wire w_dff_B_2o673iNC0_2;
	wire w_dff_B_kSb3DJfx9_2;
	wire w_dff_B_OjADhL0S8_2;
	wire w_dff_B_vLZP8QfX8_2;
	wire w_dff_B_VJWLKmx15_2;
	wire w_dff_B_OPV2nKYI3_2;
	wire w_dff_B_QFb84w6R1_2;
	wire w_dff_B_JePpGwpI0_2;
	wire w_dff_B_1GmecIhJ0_2;
	wire w_dff_B_rzNei0n85_2;
	wire w_dff_B_juJQoHav9_2;
	wire w_dff_B_aIzD0oVX4_2;
	wire w_dff_B_cm4VAGbl5_2;
	wire w_dff_B_Cc3J9Q767_2;
	wire w_dff_B_b14ti8Um9_2;
	wire w_dff_B_DqGfZ6187_2;
	wire w_dff_B_gIpXCyK06_2;
	wire w_dff_B_XTcIuCbm7_2;
	wire w_dff_B_UtYEnfsV0_2;
	wire w_dff_B_dN1bwkGW7_2;
	wire w_dff_B_wE6vxHHD9_2;
	wire w_dff_B_tv9fE4Wm7_2;
	wire w_dff_B_r6rsoiz94_2;
	wire w_dff_B_MZF1mq131_2;
	wire w_dff_B_rBqYzJFi0_2;
	wire w_dff_B_32RysaDw5_2;
	wire w_dff_B_ELbAWnj27_2;
	wire w_dff_B_wxgzp5I84_2;
	wire w_dff_B_K1XiXgqB3_2;
	wire w_dff_B_k0NqPBpU2_2;
	wire w_dff_B_BjKCTGGi5_2;
	wire w_dff_B_ePWWhOLk3_2;
	wire w_dff_B_rylctyCW3_1;
	wire w_dff_B_h7ZEuDmb1_2;
	wire w_dff_B_XW4nAG976_2;
	wire w_dff_B_O7fUxSqP4_2;
	wire w_dff_B_cntEbQlR6_2;
	wire w_dff_B_hAMfUTEM1_2;
	wire w_dff_B_mK4vNNN49_2;
	wire w_dff_B_JrSkrzBt2_2;
	wire w_dff_B_4mXIw4G31_2;
	wire w_dff_B_s6AGkWEw1_2;
	wire w_dff_B_pmLr7PiL8_2;
	wire w_dff_B_gmcXlm5D8_2;
	wire w_dff_B_5rz6BiMc4_2;
	wire w_dff_B_q7FfvtVf9_2;
	wire w_dff_B_i1n3hgjd3_2;
	wire w_dff_B_Xuwj6L0a2_2;
	wire w_dff_B_sWDo2ve35_2;
	wire w_dff_B_KjibuJZR4_2;
	wire w_dff_B_SzcEGYeH3_2;
	wire w_dff_B_tk7FzxHW9_2;
	wire w_dff_B_GAuTDEMm7_2;
	wire w_dff_B_jngsmj9g9_2;
	wire w_dff_B_nbJs1NSe2_2;
	wire w_dff_B_1eRRJEff6_2;
	wire w_dff_B_jcR34zYb3_2;
	wire w_dff_B_RNtilsMg7_2;
	wire w_dff_B_DiD7gUH36_2;
	wire w_dff_B_rO4yVsyQ4_2;
	wire w_dff_B_yTAa6dks2_2;
	wire w_dff_B_qClnjBV82_2;
	wire w_dff_B_kczOsCVx1_2;
	wire w_dff_B_lyAVx1hT1_2;
	wire w_dff_B_kpM1PmIY4_2;
	wire w_dff_B_92dOxz244_2;
	wire w_dff_B_YdQRyXzW3_2;
	wire w_dff_B_h5K9Dn802_2;
	wire w_dff_B_z0jUJwcp6_2;
	wire w_dff_B_QHULyD6b3_2;
	wire w_dff_B_enjR0FLW7_2;
	wire w_dff_B_gbgBrA6H6_2;
	wire w_dff_B_QTjBzVB43_1;
	wire w_dff_B_i90TR0Ua5_1;
	wire w_dff_B_c4PhMsCI1_2;
	wire w_dff_B_StDVmxxv0_2;
	wire w_dff_B_3KKf0lg50_2;
	wire w_dff_B_OcTWDznu4_2;
	wire w_dff_B_MayoLo4z6_2;
	wire w_dff_B_e5Sz9ZE24_2;
	wire w_dff_B_NEolJuh88_2;
	wire w_dff_B_Eh0OcCbs4_2;
	wire w_dff_B_tK3opf0D2_2;
	wire w_dff_B_tPAK43lg2_2;
	wire w_dff_B_7Rp5K8FC7_2;
	wire w_dff_B_ONhdkeAp1_2;
	wire w_dff_B_Y9fCuxhB1_2;
	wire w_dff_B_PoFFkXua0_2;
	wire w_dff_B_9hCnEWZb8_2;
	wire w_dff_B_QbOGr7ud5_2;
	wire w_dff_B_oUIGYaME2_2;
	wire w_dff_B_cUjtq5cu9_2;
	wire w_dff_B_C092x4oO9_2;
	wire w_dff_B_QwpZgVzd6_2;
	wire w_dff_B_CrRsneMV1_2;
	wire w_dff_B_YAhGya4r9_2;
	wire w_dff_B_K7VY47iV8_2;
	wire w_dff_B_5eYdc7KG1_2;
	wire w_dff_B_3V3F6zdX0_2;
	wire w_dff_B_6iv68eh54_2;
	wire w_dff_B_XZv4HD2E6_2;
	wire w_dff_B_sRTjxp2a0_2;
	wire w_dff_B_fv8t0Bza5_2;
	wire w_dff_B_k0LAeEIJ7_2;
	wire w_dff_B_LGWN4t5i1_2;
	wire w_dff_B_51cAvMAn6_2;
	wire w_dff_B_85WyqBzm6_2;
	wire w_dff_B_pPRrrqhz7_2;
	wire w_dff_B_wOY6VAb33_2;
	wire w_dff_B_2DNCISpa2_2;
	wire w_dff_B_GmSNJfGn1_2;
	wire w_dff_B_ieUl5OA25_2;
	wire w_dff_B_Uuc2mR2h3_2;
	wire w_dff_B_LhCAu3xo2_2;
	wire w_dff_B_HMMMaqZh7_2;
	wire w_dff_B_8TgWaTU67_2;
	wire w_dff_B_zhmz6o6t0_2;
	wire w_dff_B_HJxKRaJ90_2;
	wire w_dff_B_yNmbtX614_2;
	wire w_dff_B_1r47iof57_2;
	wire w_dff_B_Q9SM2Lsz5_2;
	wire w_dff_B_olZKlNhv5_2;
	wire w_dff_B_G0wzwvvP3_2;
	wire w_dff_B_aIk4xXLa3_2;
	wire w_dff_B_FDJEGcJc0_2;
	wire w_dff_B_xo97B67i0_2;
	wire w_dff_B_xra00VK92_2;
	wire w_dff_B_7nprEDef0_2;
	wire w_dff_B_4vkip1Mz2_2;
	wire w_dff_B_HSe8mv4g1_2;
	wire w_dff_B_YrW8t61X7_2;
	wire w_dff_B_KLaxzF2E9_2;
	wire w_dff_B_9FjxJDhb4_2;
	wire w_dff_B_A17wngXb2_2;
	wire w_dff_B_rB2Act2P8_2;
	wire w_dff_B_3plsBdUM3_2;
	wire w_dff_B_902ADQ0l9_2;
	wire w_dff_B_ubUYKFxu5_2;
	wire w_dff_B_xGAa1utb7_2;
	wire w_dff_B_4sZXHQzC0_2;
	wire w_dff_B_cNkkEb6X9_2;
	wire w_dff_B_e2SNW1oG5_2;
	wire w_dff_B_rZ6eexFO1_2;
	wire w_dff_B_Tsq3goMi8_2;
	wire w_dff_B_KBcD8O4V7_2;
	wire w_dff_B_vXqmdnz53_2;
	wire w_dff_B_UX9PxSwT3_2;
	wire w_dff_B_yUI2ohxu1_2;
	wire w_dff_B_gSyS7sQ69_2;
	wire w_dff_B_Rr9uOYLY4_1;
	wire w_dff_B_okHtaBRA2_2;
	wire w_dff_B_xx9G1Dyj8_2;
	wire w_dff_B_yRag1ri84_2;
	wire w_dff_B_SIMKDxEc0_2;
	wire w_dff_B_de8eGcce1_2;
	wire w_dff_B_zNqEkX4g3_2;
	wire w_dff_B_4qnSNbtp3_2;
	wire w_dff_B_E37uSIUu7_2;
	wire w_dff_B_BU1yaWKR0_2;
	wire w_dff_B_VMAeXGvG8_2;
	wire w_dff_B_63Z5XYfG8_2;
	wire w_dff_B_ZZnGvgRo4_2;
	wire w_dff_B_f8kW5op81_2;
	wire w_dff_B_WsTIjQt01_2;
	wire w_dff_B_m4zY4HUi9_2;
	wire w_dff_B_WS1Me9cY2_2;
	wire w_dff_B_9aMRIZGK7_2;
	wire w_dff_B_gEKPAs8u9_2;
	wire w_dff_B_RWvFzPX89_2;
	wire w_dff_B_qsbvViJb7_2;
	wire w_dff_B_1hbuWucZ6_2;
	wire w_dff_B_6hZsfQ1Q4_2;
	wire w_dff_B_ztzdxNGC1_2;
	wire w_dff_B_sfmfHssI1_2;
	wire w_dff_B_W0YaUfP97_2;
	wire w_dff_B_Kx17gVau7_2;
	wire w_dff_B_A5AUQ41I8_2;
	wire w_dff_B_rjO2eZd75_2;
	wire w_dff_B_0ZIOGgvX4_2;
	wire w_dff_B_zgmLNUQJ3_2;
	wire w_dff_B_MYyxT8Ur6_2;
	wire w_dff_B_dSWEfCHf0_2;
	wire w_dff_B_hd1LKUtf0_2;
	wire w_dff_B_NPRYPLEI1_2;
	wire w_dff_B_h3LpYNfB5_2;
	wire w_dff_B_ZPhpAERb4_2;
	wire w_dff_B_SPRTuclL2_1;
	wire w_dff_B_Nayzih5N8_1;
	wire w_dff_B_stb9LMXH6_2;
	wire w_dff_B_geNNOI4z0_2;
	wire w_dff_B_JSH3k4pL4_2;
	wire w_dff_B_SQBg60se5_2;
	wire w_dff_B_Ho41pmSb0_2;
	wire w_dff_B_lZRLbIjL6_2;
	wire w_dff_B_eiNf6T714_2;
	wire w_dff_B_kNqznUS58_2;
	wire w_dff_B_gZ2N9WDJ5_2;
	wire w_dff_B_NjJntgbw3_2;
	wire w_dff_B_E0WdK6zA3_2;
	wire w_dff_B_RmcELb6R1_2;
	wire w_dff_B_HgmlUmpy4_2;
	wire w_dff_B_8zHZDOVm9_2;
	wire w_dff_B_csGE3hON3_2;
	wire w_dff_B_kQp97ZQk9_2;
	wire w_dff_B_FsmNUmCF8_2;
	wire w_dff_B_DGMFsyGd6_2;
	wire w_dff_B_fPhm7dyX2_2;
	wire w_dff_B_9guEDIXx9_2;
	wire w_dff_B_KmDdxCba2_2;
	wire w_dff_B_XNDjEVCQ2_2;
	wire w_dff_B_BCoDk1Ig3_2;
	wire w_dff_B_aPpzmYqb7_2;
	wire w_dff_B_2wQQ5OD01_2;
	wire w_dff_B_h2aLBisn5_2;
	wire w_dff_B_jQwbdlRs4_2;
	wire w_dff_B_h5EXYLZM4_2;
	wire w_dff_B_KKv14GYh4_2;
	wire w_dff_B_aLg9hG0Z2_2;
	wire w_dff_B_vmd2Q5af3_2;
	wire w_dff_B_hQc1PwNP7_2;
	wire w_dff_B_z5QIOJ2o2_2;
	wire w_dff_B_qaN1el2k1_2;
	wire w_dff_B_wUP8miuQ0_2;
	wire w_dff_B_xgifIYVK2_2;
	wire w_dff_B_YqcuE0Aq2_2;
	wire w_dff_B_at3yg0Wa3_2;
	wire w_dff_B_calvw9OX5_2;
	wire w_dff_B_FtpxofnM3_2;
	wire w_dff_B_blQ0iAMY6_2;
	wire w_dff_B_ykb41ZJk3_2;
	wire w_dff_B_HQOsVYbb9_2;
	wire w_dff_B_Zqun5X929_2;
	wire w_dff_B_8bNObTPf5_2;
	wire w_dff_B_TEvqXDKt6_2;
	wire w_dff_B_nkr8ubmc5_2;
	wire w_dff_B_Q2hQ9NlK8_2;
	wire w_dff_B_6Qqdk2Lk0_2;
	wire w_dff_B_YqCrXgWI6_2;
	wire w_dff_B_NFPIrlfV1_2;
	wire w_dff_B_RseZyUiX8_2;
	wire w_dff_B_k6nek2va8_2;
	wire w_dff_B_XgHjjRfO2_2;
	wire w_dff_B_1Z3dvCvs0_2;
	wire w_dff_B_V197taw22_2;
	wire w_dff_B_PVwL3f5e5_2;
	wire w_dff_B_poW69XPH2_2;
	wire w_dff_B_ZFnKktzJ7_2;
	wire w_dff_B_B44wpiev2_2;
	wire w_dff_B_PcvOIpH55_2;
	wire w_dff_B_LQ1euEiA0_2;
	wire w_dff_B_uX5JAVHG6_2;
	wire w_dff_B_EhALhOGY7_2;
	wire w_dff_B_IA2fbPFR6_2;
	wire w_dff_B_y9OtsbHg3_2;
	wire w_dff_B_foVNVH4X5_2;
	wire w_dff_B_bqTe6Lzj1_2;
	wire w_dff_B_c0Qs8dBf7_2;
	wire w_dff_B_IzfRDnTa7_1;
	wire w_dff_B_Zb99ZdHS8_2;
	wire w_dff_B_NgIO3hqL1_2;
	wire w_dff_B_qQrhE51o0_2;
	wire w_dff_B_9Y5WYIJl9_2;
	wire w_dff_B_OVknh3e76_2;
	wire w_dff_B_7eFjvere8_2;
	wire w_dff_B_IEnjttNr2_2;
	wire w_dff_B_Hg6inLPI1_2;
	wire w_dff_B_Cx32MKBs0_2;
	wire w_dff_B_dBCK1NDD0_2;
	wire w_dff_B_JB2dtFdm3_2;
	wire w_dff_B_WDkpkpuJ9_2;
	wire w_dff_B_lhIgNy631_2;
	wire w_dff_B_5LGLQcwG5_2;
	wire w_dff_B_0EqYBEXj0_2;
	wire w_dff_B_LxZ5clYQ8_2;
	wire w_dff_B_2JJiNf1a2_2;
	wire w_dff_B_DIhKgkga6_2;
	wire w_dff_B_6suNxC6B7_2;
	wire w_dff_B_Su5k1gae6_2;
	wire w_dff_B_PffExo7g1_2;
	wire w_dff_B_kKG2OM7H0_2;
	wire w_dff_B_O9sxoRsM0_2;
	wire w_dff_B_B6nsp8aL6_2;
	wire w_dff_B_HLwZpeXP4_2;
	wire w_dff_B_Iz2iBD161_2;
	wire w_dff_B_erGLMVOC2_2;
	wire w_dff_B_ffsAHrzV7_2;
	wire w_dff_B_YQ04Rc9S9_2;
	wire w_dff_B_Lo7HHNol8_2;
	wire w_dff_B_W0Tf1de92_2;
	wire w_dff_B_x5ZwqFSH7_2;
	wire w_dff_B_GUFsXUGN2_2;
	wire w_dff_B_PvsmpJBm4_1;
	wire w_dff_B_YErMqfjS7_1;
	wire w_dff_B_qTDl1epY8_2;
	wire w_dff_B_dDsdxMjD5_2;
	wire w_dff_B_Qzf46XOn9_2;
	wire w_dff_B_eLYoqyXj5_2;
	wire w_dff_B_XJowFD5f6_2;
	wire w_dff_B_AaeF6JTK5_2;
	wire w_dff_B_lGbbPq324_2;
	wire w_dff_B_hFDsIOkN8_2;
	wire w_dff_B_MEqaN5ff8_2;
	wire w_dff_B_aFCi0B621_2;
	wire w_dff_B_UxLDaFzC9_2;
	wire w_dff_B_knTuofbS1_2;
	wire w_dff_B_LydvIIcl3_2;
	wire w_dff_B_WdvVUIfB1_2;
	wire w_dff_B_rYtbfWX81_2;
	wire w_dff_B_nZRIjCSh5_2;
	wire w_dff_B_aE4QKcva3_2;
	wire w_dff_B_PM4EtVMa2_2;
	wire w_dff_B_20TzXt6y4_2;
	wire w_dff_B_v29Brma90_2;
	wire w_dff_B_lpNCN7Zg9_2;
	wire w_dff_B_n0dwKKlZ7_2;
	wire w_dff_B_rL8TNgld4_2;
	wire w_dff_B_fIg1iSPN4_2;
	wire w_dff_B_Ze42DfCH0_2;
	wire w_dff_B_QC5OYXZP7_2;
	wire w_dff_B_peGCjqIh5_2;
	wire w_dff_B_rNmU3GZY7_2;
	wire w_dff_B_JkyxggJK2_2;
	wire w_dff_B_mXwsCmDM5_2;
	wire w_dff_B_OUwHMjED9_2;
	wire w_dff_B_xtLV87IE7_2;
	wire w_dff_B_aJYdTGTJ0_2;
	wire w_dff_B_v1Pr301H3_2;
	wire w_dff_B_D59cdu1h4_2;
	wire w_dff_B_BMC5zDa01_2;
	wire w_dff_B_LPf4mr7G3_2;
	wire w_dff_B_K6IO6Mxv3_2;
	wire w_dff_B_ruFLtfx99_2;
	wire w_dff_B_3OtWJJV04_2;
	wire w_dff_B_beJocVUY1_2;
	wire w_dff_B_3TqRlnEJ4_2;
	wire w_dff_B_FWq85ip66_2;
	wire w_dff_B_LUNRbAaB4_2;
	wire w_dff_B_OLtQc3iX0_2;
	wire w_dff_B_vnNLjbK79_2;
	wire w_dff_B_ktNM0r6b7_2;
	wire w_dff_B_Nnb4YZRZ2_2;
	wire w_dff_B_ojFpsxO98_2;
	wire w_dff_B_IBCwZT5t5_2;
	wire w_dff_B_Pt0nCbGD5_2;
	wire w_dff_B_y7vLdVIX1_2;
	wire w_dff_B_4CbKcEhX3_2;
	wire w_dff_B_XCzWQrqQ6_2;
	wire w_dff_B_K4p38FV20_2;
	wire w_dff_B_zhm2YRNX7_2;
	wire w_dff_B_aa7M3sTb8_2;
	wire w_dff_B_R1sPw8fa1_2;
	wire w_dff_B_ZKa8ociC4_2;
	wire w_dff_B_c63vPWyR8_2;
	wire w_dff_B_xLB5aAUQ2_2;
	wire w_dff_B_QZUrIAZs9_2;
	wire w_dff_B_qSMUqC6J3_2;
	wire w_dff_B_VbSDAllf5_1;
	wire w_dff_B_hTrstGvu4_2;
	wire w_dff_B_RTlQfiI71_2;
	wire w_dff_B_gP53vt9F2_2;
	wire w_dff_B_Z5Vjm5Mo1_2;
	wire w_dff_B_vARs2y1j7_2;
	wire w_dff_B_5xtCwI856_2;
	wire w_dff_B_bR7vL1k10_2;
	wire w_dff_B_CTS5lpnv8_2;
	wire w_dff_B_StKDVNTE2_2;
	wire w_dff_B_P7lCUDBB5_2;
	wire w_dff_B_pII7MEJH8_2;
	wire w_dff_B_m5GOJuzq7_2;
	wire w_dff_B_kJtpIqHu9_2;
	wire w_dff_B_ZISNOnRE6_2;
	wire w_dff_B_OcpfefGm4_2;
	wire w_dff_B_OOQ7tIpY5_2;
	wire w_dff_B_vEivhFuV5_2;
	wire w_dff_B_66mgbrko4_2;
	wire w_dff_B_XOyCFZ7v3_2;
	wire w_dff_B_kApYDfkX9_2;
	wire w_dff_B_bakpFhan4_2;
	wire w_dff_B_HskodKWb7_2;
	wire w_dff_B_uY2M1oMY0_2;
	wire w_dff_B_BKQkdCnk2_2;
	wire w_dff_B_nv58PPcL1_2;
	wire w_dff_B_mR9KjR2E5_2;
	wire w_dff_B_QF8iOlUM9_2;
	wire w_dff_B_NEN9KgV76_2;
	wire w_dff_B_vCxmitVU2_2;
	wire w_dff_B_5vAg64vY8_2;
	wire w_dff_B_bKEYKbbV9_1;
	wire w_dff_B_3KAZd9Je8_1;
	wire w_dff_B_Vaq02DPH7_2;
	wire w_dff_B_Bnd9QY6c3_2;
	wire w_dff_B_oDdsBWCC3_2;
	wire w_dff_B_XTsRPkOW9_2;
	wire w_dff_B_QJMmha5K4_2;
	wire w_dff_B_v9qSeM8R5_2;
	wire w_dff_B_r721UY4v2_2;
	wire w_dff_B_NS5UwBBF0_2;
	wire w_dff_B_3LJWnYas0_2;
	wire w_dff_B_e273UyQ47_2;
	wire w_dff_B_sxlwXp1o0_2;
	wire w_dff_B_6ypBymCa2_2;
	wire w_dff_B_PkEeP02S0_2;
	wire w_dff_B_k5xa1wZ94_2;
	wire w_dff_B_gNcwLOgK5_2;
	wire w_dff_B_Ux6I4cQt8_2;
	wire w_dff_B_yL9mW64V9_2;
	wire w_dff_B_cpQSAWmr5_2;
	wire w_dff_B_7EwULnyV2_2;
	wire w_dff_B_41bdJH389_2;
	wire w_dff_B_J5o1CbXZ4_2;
	wire w_dff_B_mnS48AB18_2;
	wire w_dff_B_QanCfR3c3_2;
	wire w_dff_B_eef1ZK2M2_2;
	wire w_dff_B_1w2h16bM3_2;
	wire w_dff_B_nVvhYrmC6_2;
	wire w_dff_B_bsop8f2T8_2;
	wire w_dff_B_gRduZacn2_2;
	wire w_dff_B_FYGPnNpu9_2;
	wire w_dff_B_U72RIqzP6_2;
	wire w_dff_B_Ye12bHrZ4_2;
	wire w_dff_B_tdQHx3IX6_2;
	wire w_dff_B_b5n9cWZD5_2;
	wire w_dff_B_W8rA4ORs4_2;
	wire w_dff_B_RTBweTss8_2;
	wire w_dff_B_pBfnd1Mh9_2;
	wire w_dff_B_rsubGjLf5_2;
	wire w_dff_B_twt5G07e5_2;
	wire w_dff_B_AuVUz9C37_2;
	wire w_dff_B_QgPmRcTe4_2;
	wire w_dff_B_hADkqKJi8_2;
	wire w_dff_B_Iv9JaAqt2_2;
	wire w_dff_B_jJazrxyt0_2;
	wire w_dff_B_P8AMhOAB1_2;
	wire w_dff_B_nv02lWB33_2;
	wire w_dff_B_9mDozcmb5_2;
	wire w_dff_B_jrhByb670_2;
	wire w_dff_B_4XLpSYJq5_2;
	wire w_dff_B_aK6adQKb1_2;
	wire w_dff_B_xaspD9l37_2;
	wire w_dff_B_xK8wlVqX9_2;
	wire w_dff_B_IwqRa1pJ4_2;
	wire w_dff_B_RHRcBqPg9_2;
	wire w_dff_B_eRk4JWa99_2;
	wire w_dff_B_5fK0CbFV1_2;
	wire w_dff_B_Jl7bPsJO7_2;
	wire w_dff_B_ZgtcSHaY9_2;
	wire w_dff_B_8AToENM26_1;
	wire w_dff_B_hYO2MQ7m6_2;
	wire w_dff_B_wEb6SDTz8_2;
	wire w_dff_B_uJfVdAMq6_2;
	wire w_dff_B_z0AXP81o5_2;
	wire w_dff_B_54pIyioL7_2;
	wire w_dff_B_TkA8Iy4I9_2;
	wire w_dff_B_16xdJ4M99_2;
	wire w_dff_B_2lrtg4CN8_2;
	wire w_dff_B_cBxlOMyj7_2;
	wire w_dff_B_1cZNdXJN4_2;
	wire w_dff_B_HMm2gWIm2_2;
	wire w_dff_B_uROQAyYm0_2;
	wire w_dff_B_ZGHPxLHT4_2;
	wire w_dff_B_BoxmYpWt9_2;
	wire w_dff_B_s147yXgz8_2;
	wire w_dff_B_ig0Z2EHv7_2;
	wire w_dff_B_isverOzf2_2;
	wire w_dff_B_h0ACUAL07_2;
	wire w_dff_B_jxWozL602_2;
	wire w_dff_B_s3eZUIUA3_2;
	wire w_dff_B_otmrRu990_2;
	wire w_dff_B_hgAjOtlX1_2;
	wire w_dff_B_MtgfJ5PA9_2;
	wire w_dff_B_0jd2Rb4T7_2;
	wire w_dff_B_9EQoKnIl6_2;
	wire w_dff_B_WKfFzGgQ2_2;
	wire w_dff_B_ztfniFbs0_2;
	wire w_dff_B_Uqw05TLl4_1;
	wire w_dff_B_KARzh2LJ3_1;
	wire w_dff_B_SwQ8kzZG9_2;
	wire w_dff_B_qTWxOjmh9_2;
	wire w_dff_B_FArDLjPv7_2;
	wire w_dff_B_63ryLsMq7_2;
	wire w_dff_B_U8UxU3bN4_2;
	wire w_dff_B_pRJYqoAl5_2;
	wire w_dff_B_pKRAuQqg9_2;
	wire w_dff_B_n0GmbCEk2_2;
	wire w_dff_B_UmyYzFAS5_2;
	wire w_dff_B_0VikFm1P0_2;
	wire w_dff_B_U1z4qvW22_2;
	wire w_dff_B_TdHEhK7J7_2;
	wire w_dff_B_Tpj7kjtB6_2;
	wire w_dff_B_jNTNi3Tg3_2;
	wire w_dff_B_FBmyCJL18_2;
	wire w_dff_B_4SpswkaO6_2;
	wire w_dff_B_cJqfEbKN8_2;
	wire w_dff_B_yjSWSKcy7_2;
	wire w_dff_B_H6IypFwe6_2;
	wire w_dff_B_6oq6cpMR6_2;
	wire w_dff_B_H8R0rlwr1_2;
	wire w_dff_B_kh1UKGBO4_2;
	wire w_dff_B_6KOgTE5Z4_2;
	wire w_dff_B_dHTgEsif0_2;
	wire w_dff_B_PY28HlVW5_2;
	wire w_dff_B_Ntj80Knl4_2;
	wire w_dff_B_QevNkeav6_2;
	wire w_dff_B_kCvtrqo36_2;
	wire w_dff_B_wsbb7vzP7_2;
	wire w_dff_B_NwcEb03n2_2;
	wire w_dff_B_Kh6nPWOF1_2;
	wire w_dff_B_H1L0yD0s7_2;
	wire w_dff_B_FUOZRwUc9_2;
	wire w_dff_B_EG79hSRm9_2;
	wire w_dff_B_QwBL5dEG8_2;
	wire w_dff_B_r2R7smak5_2;
	wire w_dff_B_6pTO68Sw0_2;
	wire w_dff_B_T2bqYwub4_2;
	wire w_dff_B_556b7PXp0_2;
	wire w_dff_B_tYzZqhzB6_2;
	wire w_dff_B_BvMkBAov2_2;
	wire w_dff_B_OHnCXbBO7_2;
	wire w_dff_B_QJAbgZND2_2;
	wire w_dff_B_6fdHWPhQ1_2;
	wire w_dff_B_b6wd8B4S1_2;
	wire w_dff_B_bmSptCoe5_2;
	wire w_dff_B_RmDgsv8m9_2;
	wire w_dff_B_HXg69b2L5_2;
	wire w_dff_B_XzRk4iNO4_2;
	wire w_dff_B_6vXFpnbZ4_2;
	wire w_dff_B_PXxDP2ZQ2_2;
	wire w_dff_B_s0iMEh9j6_1;
	wire w_dff_B_mWOa81Rk5_2;
	wire w_dff_B_ISny6vEW4_2;
	wire w_dff_B_BvuQ1cza0_2;
	wire w_dff_B_weaMn54Z0_2;
	wire w_dff_B_rQgBqpsl1_2;
	wire w_dff_B_T6hGHSEv5_2;
	wire w_dff_B_w5wkDeUs3_2;
	wire w_dff_B_flvje6QQ0_2;
	wire w_dff_B_F6k9YprD2_2;
	wire w_dff_B_T3DxtkCa9_2;
	wire w_dff_B_yjUduDbD6_2;
	wire w_dff_B_Dk5lbwa53_2;
	wire w_dff_B_cUDNQNix4_2;
	wire w_dff_B_CaOXVu8i4_2;
	wire w_dff_B_Ssn2jGft0_2;
	wire w_dff_B_kppgszoA2_2;
	wire w_dff_B_djuiL1bi5_2;
	wire w_dff_B_RGy0bzld9_2;
	wire w_dff_B_WbMsBM4E3_2;
	wire w_dff_B_vlCMFHgH6_2;
	wire w_dff_B_NjwkrKHV4_2;
	wire w_dff_B_Ayj4Rhso9_2;
	wire w_dff_B_v7oCyk8L3_2;
	wire w_dff_B_j9F6fm7H5_2;
	wire w_dff_B_rhDUsWj34_1;
	wire w_dff_B_CsrK5ZqW4_1;
	wire w_dff_B_hXMUlXj97_2;
	wire w_dff_B_vn4HAjen4_2;
	wire w_dff_B_lLZPluQI1_2;
	wire w_dff_B_iFJeX5hP4_2;
	wire w_dff_B_2NtFqqix5_2;
	wire w_dff_B_wc4Y4toX6_2;
	wire w_dff_B_UOQsEt7c9_2;
	wire w_dff_B_Jee3Zt722_2;
	wire w_dff_B_srBTgxHS2_2;
	wire w_dff_B_4VnwhoLy7_2;
	wire w_dff_B_BPb5ynIG3_2;
	wire w_dff_B_0KARpA4n3_2;
	wire w_dff_B_FT4J4oWT7_2;
	wire w_dff_B_BY6LPpUv3_2;
	wire w_dff_B_twxpVCLP9_2;
	wire w_dff_B_xdLCfyIs9_2;
	wire w_dff_B_m9TmWIG89_2;
	wire w_dff_B_ZsXnbvxn7_2;
	wire w_dff_B_tmjAr3ij4_2;
	wire w_dff_B_xMROSzql1_2;
	wire w_dff_B_0maDXt469_2;
	wire w_dff_B_LAHOgGhx2_2;
	wire w_dff_B_rSecc6as2_2;
	wire w_dff_B_HpFlco0h5_2;
	wire w_dff_B_v9KDYvbD4_2;
	wire w_dff_B_AEgcHMBt7_2;
	wire w_dff_B_oJyGlvUs4_2;
	wire w_dff_B_oYAFx4dZ2_2;
	wire w_dff_B_pUjFk1WI7_2;
	wire w_dff_B_8zzSTvs93_2;
	wire w_dff_B_HZ1MYFKA4_2;
	wire w_dff_B_70V6dmNT8_2;
	wire w_dff_B_4YMXx4vV4_2;
	wire w_dff_B_sKToEarR1_2;
	wire w_dff_B_tsfA4iAg5_2;
	wire w_dff_B_qX6Vr7g68_2;
	wire w_dff_B_2da2878j4_2;
	wire w_dff_B_1nLpnGve6_2;
	wire w_dff_B_4t2jPIFm1_2;
	wire w_dff_B_aWmcrJ1x8_2;
	wire w_dff_B_zUJELoid4_2;
	wire w_dff_B_nslbwkcb9_2;
	wire w_dff_B_qiGqY5316_2;
	wire w_dff_B_RaaEakny6_2;
	wire w_dff_B_CT3WHjNg5_2;
	wire w_dff_B_0LPPkpTF8_1;
	wire w_dff_B_ro4fgAqA8_2;
	wire w_dff_B_HxMFnHtK6_2;
	wire w_dff_B_RU535DrL4_2;
	wire w_dff_B_VVHSkZ501_2;
	wire w_dff_B_MjfSUJft1_2;
	wire w_dff_B_zuInLHpI9_2;
	wire w_dff_B_jVXcfI5U1_2;
	wire w_dff_B_IJvuMKKD6_2;
	wire w_dff_B_KKRfMiwM5_2;
	wire w_dff_B_H35ZoJAT4_2;
	wire w_dff_B_ZHDQzUp84_2;
	wire w_dff_B_QrQq3D3c4_2;
	wire w_dff_B_6b2pPNmg5_2;
	wire w_dff_B_UfrgNYyG2_2;
	wire w_dff_B_9bSCueTo5_2;
	wire w_dff_B_45HiwsA46_2;
	wire w_dff_B_cbzno6ca3_2;
	wire w_dff_B_ijZyGR887_2;
	wire w_dff_B_KEqVdexm6_2;
	wire w_dff_B_ppiFikWv1_2;
	wire w_dff_B_kU5hk7Wz5_2;
	wire w_dff_B_4CfiHYsM2_1;
	wire w_dff_B_zYK4DSNq2_1;
	wire w_dff_B_NygoV7GR9_2;
	wire w_dff_B_PpOnQ7r68_2;
	wire w_dff_B_6OGf1WYy6_2;
	wire w_dff_B_seqL7K5u9_2;
	wire w_dff_B_vWRcOAUg8_2;
	wire w_dff_B_AZUq8oyp9_2;
	wire w_dff_B_YZTjUDOJ7_2;
	wire w_dff_B_p9zWEvwv3_2;
	wire w_dff_B_6ZL7mFoF1_2;
	wire w_dff_B_fwnuFRtw0_2;
	wire w_dff_B_vLF1sW0w2_2;
	wire w_dff_B_B6bilmLw3_2;
	wire w_dff_B_o85svmNf2_2;
	wire w_dff_B_H3ektXat2_2;
	wire w_dff_B_YJSIwh8n5_2;
	wire w_dff_B_msx7xnt23_2;
	wire w_dff_B_JBteyBSG0_2;
	wire w_dff_B_NAN3wn5C2_2;
	wire w_dff_B_9b31hflg2_2;
	wire w_dff_B_bn4XXQ5L1_2;
	wire w_dff_B_uvPZUm570_2;
	wire w_dff_B_RksPpFYX7_2;
	wire w_dff_B_JxM20JC14_2;
	wire w_dff_B_M9ak3Kws1_2;
	wire w_dff_B_ZsqlUFPP8_2;
	wire w_dff_B_MK1w0YYY3_2;
	wire w_dff_B_gioAlult0_2;
	wire w_dff_B_Gx76qa393_2;
	wire w_dff_B_kazSnlUS4_2;
	wire w_dff_B_pMtSoTl52_2;
	wire w_dff_B_0t1rKXzn2_2;
	wire w_dff_B_yEeBVL2n2_2;
	wire w_dff_B_dl3Fhrn45_2;
	wire w_dff_B_01Mgn8cX3_2;
	wire w_dff_B_LVChLgIA8_2;
	wire w_dff_B_ePEybjNl3_2;
	wire w_dff_B_SxlNqlx32_2;
	wire w_dff_B_mDRr7Giz8_2;
	wire w_dff_B_t2KKPViJ5_2;
	wire w_dff_B_85e2vVXL1_1;
	wire w_dff_B_0fauM9z03_2;
	wire w_dff_B_6jgaNYdq6_2;
	wire w_dff_B_iimuTfWp8_2;
	wire w_dff_B_0hgtJpuu2_2;
	wire w_dff_B_aqNhh1yW0_2;
	wire w_dff_B_JHAjo6kM2_2;
	wire w_dff_B_OZWJKUHE3_2;
	wire w_dff_B_Do8llFkC3_2;
	wire w_dff_B_ggfJMlwP0_2;
	wire w_dff_B_ggkfeHJt8_2;
	wire w_dff_B_E2Wox0Cw8_2;
	wire w_dff_B_FpCNkiiD7_2;
	wire w_dff_B_1GCLjYcJ5_2;
	wire w_dff_B_sSXmnpaj4_2;
	wire w_dff_B_xWS4CZJz3_2;
	wire w_dff_B_kmkDCwf04_2;
	wire w_dff_B_3HXppIed7_2;
	wire w_dff_B_L60jpsp08_2;
	wire w_dff_B_vNIMQ7pO9_1;
	wire w_dff_B_Oa0pA2St3_1;
	wire w_dff_B_VPvmGoH24_2;
	wire w_dff_B_8FBpPTDB6_2;
	wire w_dff_B_jmc6jy0Q9_2;
	wire w_dff_B_ya44IFzw8_2;
	wire w_dff_B_6rUjq6ZQ4_2;
	wire w_dff_B_rVlMZDtL8_2;
	wire w_dff_B_SVnO8GHo7_2;
	wire w_dff_B_yxSeJoTe5_2;
	wire w_dff_B_TTzUi0Sw7_2;
	wire w_dff_B_BLNBaMqb2_2;
	wire w_dff_B_qXrdNVGE2_2;
	wire w_dff_B_5f7cjCv48_2;
	wire w_dff_B_KeOJ60LY6_2;
	wire w_dff_B_XIIP9E6T4_2;
	wire w_dff_B_e44LNbve0_2;
	wire w_dff_B_pSTBK2IA9_2;
	wire w_dff_B_gUWPyqyB6_2;
	wire w_dff_B_1xTkYIv49_2;
	wire w_dff_B_EnfHMm6L9_2;
	wire w_dff_B_sFJ9tXPQ9_2;
	wire w_dff_B_vp5o16l02_2;
	wire w_dff_B_DlAJR0Oy0_2;
	wire w_dff_B_VCfUbysu6_2;
	wire w_dff_B_lrtzWRUR1_2;
	wire w_dff_B_rpekBJZO8_2;
	wire w_dff_B_VvlGChyo2_2;
	wire w_dff_B_82CmETf92_2;
	wire w_dff_B_YIzQmC5H5_2;
	wire w_dff_B_aydLwHWl5_2;
	wire w_dff_B_EmJgA1MC3_2;
	wire w_dff_B_lqajwhXR8_2;
	wire w_dff_B_GjFxFVhf7_2;
	wire w_dff_B_D4V5DroH4_2;
	wire w_dff_B_JkXbNzCC9_1;
	wire w_dff_B_hYkSZRMO2_2;
	wire w_dff_B_kk2dACGn6_2;
	wire w_dff_B_a37rvPZh4_2;
	wire w_dff_B_nlY0VBjh2_2;
	wire w_dff_B_vUYkJgk47_2;
	wire w_dff_B_lwe0PPRo7_2;
	wire w_dff_B_ojwBDWI14_2;
	wire w_dff_B_1NxNfpFi0_2;
	wire w_dff_B_u11dyIK55_2;
	wire w_dff_B_iRMJOcA28_2;
	wire w_dff_B_7NUR15Zs0_2;
	wire w_dff_B_VtKaEXlg4_2;
	wire w_dff_B_3asc5Gvr4_2;
	wire w_dff_B_IjuRj1ww2_2;
	wire w_dff_B_rKVR8sWE1_2;
	wire w_dff_B_crnr4qrw6_1;
	wire w_dff_B_moMeQzNZ4_1;
	wire w_dff_B_jArypyh02_2;
	wire w_dff_B_3EbBvGA42_2;
	wire w_dff_B_afahBYJG0_2;
	wire w_dff_B_k2p4wguJ8_2;
	wire w_dff_B_NR3jfjt91_2;
	wire w_dff_B_aPVnDS1Z4_2;
	wire w_dff_B_YXuXaoNM9_2;
	wire w_dff_B_g6RJ1NVC7_2;
	wire w_dff_B_gx6K9Wow9_2;
	wire w_dff_B_TwhgTcSW8_2;
	wire w_dff_B_4g2faHve1_2;
	wire w_dff_B_Ki1nZEhn6_2;
	wire w_dff_B_tegQGoKM7_2;
	wire w_dff_B_UgIDderV0_2;
	wire w_dff_B_NXH9GbrM0_2;
	wire w_dff_B_Twdf0ORp8_2;
	wire w_dff_B_coGlQVZF5_2;
	wire w_dff_B_4d6xiDjR5_2;
	wire w_dff_B_9w8S3GlZ9_2;
	wire w_dff_B_4pyJrmRF8_2;
	wire w_dff_B_4EOU09hD8_2;
	wire w_dff_B_POmBTAvC7_2;
	wire w_dff_B_WxnuOMZF6_2;
	wire w_dff_B_BmwIfJcz5_2;
	wire w_dff_B_cab2Nc215_2;
	wire w_dff_B_QhMgLiIT7_2;
	wire w_dff_B_JjO1MDJb9_2;
	wire w_dff_B_6OoSuzZF7_1;
	wire w_dff_B_fX8bTeqw0_2;
	wire w_dff_B_vpfPPq250_2;
	wire w_dff_B_BQqIShCe6_2;
	wire w_dff_B_lRZTpFWs1_2;
	wire w_dff_B_x1YsHaaj2_2;
	wire w_dff_B_TuaFXoE17_2;
	wire w_dff_B_pPON8ijK0_2;
	wire w_dff_B_3bezBXOB5_2;
	wire w_dff_B_6NHPVkwv5_2;
	wire w_dff_B_rBMRZ5Du1_2;
	wire w_dff_B_Sa5id6kp7_2;
	wire w_dff_B_eGtqjqZM3_2;
	wire w_dff_B_xrv1WuOu5_2;
	wire w_dff_B_Voje3uex4_2;
	wire w_dff_B_XAc0eTrz4_2;
	wire w_dff_B_KwLOO7oH1_2;
	wire w_dff_B_IdU6J5MB4_2;
	wire w_dff_B_iExQuYZR4_2;
	wire w_dff_B_3brHcHxm4_2;
	wire w_dff_B_4wJbf1jX4_2;
	wire w_dff_B_v33DHjVQ4_2;
	wire w_dff_B_RhBT1oab0_2;
	wire w_dff_B_Pc6OwOEA5_2;
	wire w_dff_B_cPFS5UMl9_2;
	wire w_dff_B_Mb4y08Yj5_2;
	wire w_dff_B_RGmyYYux5_2;
	wire w_dff_B_fQ1m8iJV7_2;
	wire w_dff_B_lfb3DuC96_2;
	wire w_dff_B_LWfmRrg24_2;
	wire w_dff_B_cbHGpwvu8_2;
	wire w_dff_B_DOCHpHWC7_2;
	wire w_dff_B_PtBSenI71_2;
	wire w_dff_B_qtCwMmqV7_2;
	wire w_dff_B_1JPldOdX0_1;
	wire w_dff_B_t2RQxvvt5_2;
	wire w_dff_B_E9dEHnKE3_2;
	wire w_dff_B_46rKKUJs4_2;
	wire w_dff_B_Q9fo6tvq9_2;
	wire w_dff_B_vmcLBHZa6_2;
	wire w_dff_B_M1cT6BMY3_2;
	wire w_dff_B_tE1xEeXB1_2;
	wire w_dff_B_ZocsiWzv7_2;
	wire w_dff_B_tmJgp1tV3_2;
	wire w_dff_A_Bpoorvzm5_0;
	wire w_dff_A_vg1N7GSx6_0;
	wire w_dff_B_BjpRqFhs3_2;
	wire w_dff_B_LsD0lV718_2;
	wire w_dff_B_VC3sdodO5_1;
	wire w_dff_B_AQKaMuAp6_1;
	wire w_dff_B_jPNVT33D5_1;
	wire w_dff_B_bUMTWNEB1_1;
	wire w_dff_B_eo89BVpV8_1;
	wire w_dff_A_MpFN9kOz1_1;
	wire w_dff_A_Dnggmsxb1_1;
	wire w_dff_A_RD7anr8l3_1;
	wire w_dff_A_OX52VQV68_1;
	wire w_dff_A_D8rU4KIX2_1;
	wire w_dff_B_unvMkBRI7_2;
	wire w_dff_B_GzSO49xg9_2;
	wire w_dff_B_3SvcwYWA5_2;
	wire w_dff_B_xoYT6RqI5_2;
	wire w_dff_B_Lo8sqDnR7_2;
	wire w_dff_B_cYi2rSmd7_2;
	wire w_dff_B_d8c3X7ZS7_2;
	wire w_dff_B_Rw9ReYqf4_2;
	wire w_dff_B_8Y9hUj1G5_2;
	wire w_dff_B_04222BGw5_1;
	wire w_dff_B_6f8sRSvr3_2;
	wire w_dff_B_jGOQpKDW6_2;
	wire w_dff_B_9LZahrSn2_2;
	wire w_dff_B_VUMRSgNd1_2;
	wire w_dff_B_UPPjNxRn4_2;
	wire w_dff_B_ImuegOsW8_2;
	wire w_dff_B_qsysMGag1_2;
	wire w_dff_B_PYu0KVco4_2;
	wire w_dff_B_fl1OZwDh9_2;
	wire w_dff_B_RUO3PTNq1_2;
	wire w_dff_A_G8AbBSSj2_0;
	wire w_dff_A_CBBvRGVn6_0;
	wire w_dff_A_be4tAm5B8_0;
	wire w_dff_A_oqTUZVoI6_1;
	wire w_dff_B_w8bbQZS44_1;
	wire w_dff_B_gOLdFHBa4_1;
	wire w_dff_B_TVSLvhh41_1;
	wire w_dff_B_NWt7fI1i0_1;
	wire w_dff_B_rAaU6uUB6_0;
	wire w_dff_A_nbVdUsEx9_0;
	wire w_dff_A_zLgoNo255_0;
	wire w_dff_A_6V0MbwZf0_1;
	wire w_dff_A_idjRVIPl0_0;
	wire w_dff_A_r6vr8Qko8_0;
	wire w_dff_B_PZUfM55S1_2;
	wire w_dff_A_BXoSWlfi3_1;
	wire w_dff_A_ztGCcWEc3_1;
	wire w_dff_A_1eNyPkSg7_1;
	wire w_dff_A_WQZtJbXd3_1;
	jand g0000(.dina(w_G273gat_7[2]),.dinb(w_G1gat_7[1]),.dout(G545gat_fa_),.clk(gclk));
	jand g0001(.dina(w_G273gat_7[1]),.dinb(w_G18gat_7[2]),.dout(n65),.clk(gclk));
	jand g0002(.dina(w_G290gat_7[2]),.dinb(w_G1gat_7[0]),.dout(n66),.clk(gclk));
	jcb g0003(.dina(n66),.dinb(w_n65_0[1]),.dout(n67));
	jand g0004(.dina(w_G290gat_7[1]),.dinb(w_G18gat_7[1]),.dout(n68),.clk(gclk));
	jand g0005(.dina(n68),.dinb(w_G545gat_0),.dout(n69),.clk(gclk));
	jnot g0006(.din(w_n69_0[1]),.dout(n70),.clk(gclk));
	jand g0007(.dina(w_n70_0[1]),.dinb(w_dff_B_KtM7KiYd4_1),.dout(G1581gat),.clk(gclk));
	jand g0008(.dina(w_G307gat_7[2]),.dinb(w_G1gat_6[2]),.dout(n72),.clk(gclk));
	jnot g0009(.din(w_n72_0[1]),.dout(n73),.clk(gclk));
	jnot g0010(.din(w_G18gat_7[0]),.dout(n74),.clk(gclk));
	jnot g0011(.din(w_G290gat_7[0]),.dout(n75),.clk(gclk));
	jcb g0012(.dina(w_n75_0[1]),.dinb(n74),.dout(n76));
	jnot g0013(.din(w_G35gat_7[2]),.dout(n77),.clk(gclk));
	jnot g0014(.din(w_G273gat_7[0]),.dout(n78),.clk(gclk));
	jcb g0015(.dina(w_n78_0[1]),.dinb(w_n77_0[1]),.dout(n79));
	jand g0016(.dina(n79),.dinb(n76),.dout(n80),.clk(gclk));
	jand g0017(.dina(w_G290gat_6[2]),.dinb(w_G35gat_7[1]),.dout(n81),.clk(gclk));
	jand g0018(.dina(w_n81_0[1]),.dinb(w_n65_0[0]),.dout(n82),.clk(gclk));
	jcb g0019(.dina(w_n82_1[1]),.dinb(n80),.dout(n83));
	jand g0020(.dina(w_dff_B_Zg4WHi4m7_0),.dinb(w_n70_0[0]),.dout(n84),.clk(gclk));
	jnot g0021(.din(w_n82_1[0]),.dout(n85),.clk(gclk));
	jand g0022(.dina(w_n85_0[1]),.dinb(w_n69_0[0]),.dout(n86),.clk(gclk));
	jcb g0023(.dina(n86),.dinb(w_n84_0[1]),.dout(n87));
	jxor g0024(.dina(w_n87_0[1]),.dinb(w_dff_B_n8Hb1rcW9_1),.dout(G1901gat),.clk(gclk));
	jand g0025(.dina(w_G324gat_7[1]),.dinb(w_G1gat_6[1]),.dout(n89),.clk(gclk));
	jnot g0026(.din(w_n89_0[1]),.dout(n90),.clk(gclk));
	jnot g0027(.din(w_n84_0[0]),.dout(n91),.clk(gclk));
	jcb g0028(.dina(w_n87_0[0]),.dinb(w_n72_0[0]),.dout(n92));
	jand g0029(.dina(w_dff_B_IDjAmrQo7_0),.dinb(n91),.dout(n93),.clk(gclk));
	jand g0030(.dina(w_G307gat_7[1]),.dinb(w_G18gat_6[2]),.dout(n94),.clk(gclk));
	jnot g0031(.din(w_n94_0[1]),.dout(n95),.clk(gclk));
	jand g0032(.dina(w_G273gat_6[2]),.dinb(w_G52gat_7[2]),.dout(n96),.clk(gclk));
	jcb g0033(.dina(w_n96_0[1]),.dinb(w_n81_0[0]),.dout(n97));
	jand g0034(.dina(w_G273gat_6[1]),.dinb(w_G35gat_7[0]),.dout(n98),.clk(gclk));
	jand g0035(.dina(w_G290gat_6[1]),.dinb(w_G52gat_7[1]),.dout(n99),.clk(gclk));
	jand g0036(.dina(w_n99_0[1]),.dinb(n98),.dout(n100),.clk(gclk));
	jnot g0037(.din(w_n100_1[1]),.dout(n101),.clk(gclk));
	jand g0038(.dina(w_n101_0[2]),.dinb(w_dff_B_cbfshor35_1),.dout(n102),.clk(gclk));
	jcb g0039(.dina(n102),.dinb(w_n82_0[2]),.dout(n103));
	jand g0040(.dina(w_n101_0[1]),.dinb(w_n82_0[1]),.dout(n104),.clk(gclk));
	jnot g0041(.din(w_n104_0[1]),.dout(n105),.clk(gclk));
	jand g0042(.dina(n105),.dinb(w_n103_0[1]),.dout(n106),.clk(gclk));
	jxor g0043(.dina(n106),.dinb(w_dff_B_RMpO3DLV2_1),.dout(n107),.clk(gclk));
	jxor g0044(.dina(w_n107_0[1]),.dinb(w_n93_0[1]),.dout(n108),.clk(gclk));
	jxor g0045(.dina(w_n108_0[1]),.dinb(w_dff_B_6OiuCooY4_1),.dout(G2223gat),.clk(gclk));
	jand g0046(.dina(w_G341gat_7[1]),.dinb(w_G1gat_6[0]),.dout(n110),.clk(gclk));
	jnot g0047(.din(w_n110_0[1]),.dout(n111),.clk(gclk));
	jnot g0048(.din(w_n107_0[0]),.dout(n112),.clk(gclk));
	jcb g0049(.dina(n112),.dinb(w_n93_0[0]),.dout(n113));
	jcb g0050(.dina(w_n108_0[0]),.dinb(w_n89_0[0]),.dout(n114));
	jand g0051(.dina(n114),.dinb(n113),.dout(n115),.clk(gclk));
	jand g0052(.dina(w_G324gat_7[0]),.dinb(w_G18gat_6[1]),.dout(n116),.clk(gclk));
	jnot g0053(.din(w_n116_0[1]),.dout(n117),.clk(gclk));
	jcb g0054(.dina(w_n75_0[0]),.dinb(w_n77_0[0]),.dout(n118));
	jnot g0055(.din(w_G52gat_7[0]),.dout(n119),.clk(gclk));
	jcb g0056(.dina(w_n78_0[0]),.dinb(n119),.dout(n120));
	jand g0057(.dina(n120),.dinb(n118),.dout(n121),.clk(gclk));
	jcb g0058(.dina(w_n100_1[0]),.dinb(n121),.dout(n122));
	jand g0059(.dina(w_dff_B_1uWchztE5_0),.dinb(w_n85_0[0]),.dout(n123),.clk(gclk));
	jcb g0060(.dina(w_n104_0[0]),.dinb(n123),.dout(n124));
	jcb g0061(.dina(n124),.dinb(w_n94_0[0]),.dout(n125));
	jand g0062(.dina(n125),.dinb(w_n103_0[0]),.dout(n126),.clk(gclk));
	jand g0063(.dina(w_G307gat_7[0]),.dinb(w_G35gat_6[2]),.dout(n127),.clk(gclk));
	jnot g0064(.din(n127),.dout(n128),.clk(gclk));
	jand g0065(.dina(w_G273gat_6[0]),.dinb(w_G69gat_7[1]),.dout(n129),.clk(gclk));
	jcb g0066(.dina(w_n129_0[1]),.dinb(w_n99_0[0]),.dout(n130));
	jand g0067(.dina(w_G290gat_6[0]),.dinb(w_G69gat_7[0]),.dout(n131),.clk(gclk));
	jand g0068(.dina(w_n131_0[1]),.dinb(w_n96_0[0]),.dout(n132),.clk(gclk));
	jnot g0069(.din(w_n132_0[2]),.dout(n133),.clk(gclk));
	jand g0070(.dina(w_n133_0[2]),.dinb(w_n130_0[1]),.dout(n134),.clk(gclk));
	jcb g0071(.dina(n134),.dinb(w_n100_0[2]),.dout(n135));
	jand g0072(.dina(w_n133_0[1]),.dinb(w_n100_0[1]),.dout(n136),.clk(gclk));
	jnot g0073(.din(n136),.dout(n137),.clk(gclk));
	jand g0074(.dina(n137),.dinb(w_dff_B_BztZO27i2_1),.dout(n138),.clk(gclk));
	jxor g0075(.dina(w_n138_0[1]),.dinb(w_n128_0[1]),.dout(n139),.clk(gclk));
	jnot g0076(.din(w_n139_0[1]),.dout(n140),.clk(gclk));
	jxor g0077(.dina(w_n140_0[1]),.dinb(w_n126_0[2]),.dout(n141),.clk(gclk));
	jxor g0078(.dina(n141),.dinb(w_dff_B_Wsh9ZRGM0_1),.dout(n142),.clk(gclk));
	jxor g0079(.dina(w_n142_0[1]),.dinb(w_n115_0[1]),.dout(n143),.clk(gclk));
	jxor g0080(.dina(w_n143_0[1]),.dinb(w_dff_B_SWAZ2BU08_1),.dout(G2548gat),.clk(gclk));
	jand g0081(.dina(w_G358gat_7[1]),.dinb(w_G1gat_5[2]),.dout(n145),.clk(gclk));
	jnot g0082(.din(w_n145_0[1]),.dout(n146),.clk(gclk));
	jnot g0083(.din(w_n142_0[0]),.dout(n147),.clk(gclk));
	jcb g0084(.dina(n147),.dinb(w_n115_0[0]),.dout(n148));
	jcb g0085(.dina(w_n143_0[0]),.dinb(w_n110_0[0]),.dout(n149));
	jand g0086(.dina(n149),.dinb(n148),.dout(n150),.clk(gclk));
	jand g0087(.dina(w_G341gat_7[0]),.dinb(w_G18gat_6[0]),.dout(n151),.clk(gclk));
	jnot g0088(.din(w_n151_0[1]),.dout(n152),.clk(gclk));
	jcb g0089(.dina(w_n140_0[0]),.dinb(w_n126_0[1]),.dout(n153));
	jxor g0090(.dina(w_n139_0[0]),.dinb(w_n126_0[0]),.dout(n154),.clk(gclk));
	jcb g0091(.dina(n154),.dinb(w_n116_0[0]),.dout(n155));
	jand g0092(.dina(n155),.dinb(n153),.dout(n156),.clk(gclk));
	jand g0093(.dina(w_G324gat_6[2]),.dinb(w_G35gat_6[1]),.dout(n157),.clk(gclk));
	jnot g0094(.din(n157),.dout(n158),.clk(gclk));
	jnot g0095(.din(w_n130_0[0]),.dout(n159),.clk(gclk));
	jcb g0096(.dina(w_n132_0[1]),.dinb(n159),.dout(n160));
	jand g0097(.dina(w_dff_B_VuZ7sJNf6_0),.dinb(w_n101_0[0]),.dout(n161),.clk(gclk));
	jand g0098(.dina(w_n138_0[0]),.dinb(w_n128_0[0]),.dout(n162),.clk(gclk));
	jcb g0099(.dina(n162),.dinb(w_dff_B_ZW6ADBYo1_1),.dout(n163));
	jand g0100(.dina(w_G307gat_6[2]),.dinb(w_G52gat_6[2]),.dout(n164),.clk(gclk));
	jnot g0101(.din(n164),.dout(n165),.clk(gclk));
	jand g0102(.dina(w_G273gat_5[2]),.dinb(w_G86gat_7[1]),.dout(n166),.clk(gclk));
	jcb g0103(.dina(w_n166_0[1]),.dinb(w_n131_0[0]),.dout(n167));
	jand g0104(.dina(w_G290gat_5[2]),.dinb(w_G86gat_7[0]),.dout(n168),.clk(gclk));
	jand g0105(.dina(w_n168_0[1]),.dinb(w_n129_0[0]),.dout(n169),.clk(gclk));
	jnot g0106(.din(w_n169_0[2]),.dout(n170),.clk(gclk));
	jand g0107(.dina(w_n170_0[1]),.dinb(w_dff_B_tNXDlT0N2_1),.dout(n171),.clk(gclk));
	jcb g0108(.dina(n171),.dinb(w_n132_0[0]),.dout(n172));
	jcb g0109(.dina(w_n169_0[1]),.dinb(w_n133_0[0]),.dout(n173));
	jand g0110(.dina(w_dff_B_vn3oQZHB7_0),.dinb(w_n172_0[1]),.dout(n174),.clk(gclk));
	jxor g0111(.dina(w_n174_0[1]),.dinb(w_n165_0[1]),.dout(n175),.clk(gclk));
	jxor g0112(.dina(w_n175_0[1]),.dinb(w_n163_0[1]),.dout(n176),.clk(gclk));
	jxor g0113(.dina(w_n176_0[1]),.dinb(w_n158_0[1]),.dout(n177),.clk(gclk));
	jnot g0114(.din(w_n177_0[1]),.dout(n178),.clk(gclk));
	jxor g0115(.dina(w_n178_0[1]),.dinb(w_n156_0[2]),.dout(n179),.clk(gclk));
	jxor g0116(.dina(n179),.dinb(w_dff_B_26rhsQip6_1),.dout(n180),.clk(gclk));
	jxor g0117(.dina(w_n180_0[1]),.dinb(w_n150_0[1]),.dout(n181),.clk(gclk));
	jxor g0118(.dina(w_n181_0[1]),.dinb(w_dff_B_E0DEu2G33_1),.dout(G2877gat),.clk(gclk));
	jand g0119(.dina(w_G375gat_7[1]),.dinb(w_G1gat_5[1]),.dout(n183),.clk(gclk));
	jnot g0120(.din(w_n183_0[1]),.dout(n184),.clk(gclk));
	jnot g0121(.din(w_n180_0[0]),.dout(n185),.clk(gclk));
	jcb g0122(.dina(n185),.dinb(w_n150_0[0]),.dout(n186));
	jcb g0123(.dina(w_n181_0[0]),.dinb(w_n145_0[0]),.dout(n187));
	jand g0124(.dina(n187),.dinb(n186),.dout(n188),.clk(gclk));
	jand g0125(.dina(w_G358gat_7[0]),.dinb(w_G18gat_5[2]),.dout(n189),.clk(gclk));
	jnot g0126(.din(w_n189_0[1]),.dout(n190),.clk(gclk));
	jcb g0127(.dina(w_n178_0[0]),.dinb(w_n156_0[1]),.dout(n191));
	jxor g0128(.dina(w_n177_0[0]),.dinb(w_n156_0[0]),.dout(n192),.clk(gclk));
	jcb g0129(.dina(n192),.dinb(w_n151_0[0]),.dout(n193));
	jand g0130(.dina(n193),.dinb(n191),.dout(n194),.clk(gclk));
	jand g0131(.dina(w_G341gat_6[2]),.dinb(w_G35gat_6[0]),.dout(n195),.clk(gclk));
	jnot g0132(.din(n195),.dout(n196),.clk(gclk));
	jand g0133(.dina(w_n175_0[0]),.dinb(w_n163_0[0]),.dout(n197),.clk(gclk));
	jand g0134(.dina(w_n176_0[0]),.dinb(w_n158_0[0]),.dout(n198),.clk(gclk));
	jcb g0135(.dina(n198),.dinb(w_dff_B_SxyvgrUB3_1),.dout(n199));
	jand g0136(.dina(w_G324gat_6[1]),.dinb(w_G52gat_6[1]),.dout(n200),.clk(gclk));
	jnot g0137(.din(n200),.dout(n201),.clk(gclk));
	jnot g0138(.din(w_n172_0[0]),.dout(n202),.clk(gclk));
	jand g0139(.dina(w_n174_0[0]),.dinb(w_n165_0[0]),.dout(n203),.clk(gclk));
	jcb g0140(.dina(n203),.dinb(w_dff_B_GK5VE46Q3_1),.dout(n204));
	jand g0141(.dina(w_G307gat_6[1]),.dinb(w_G69gat_6[2]),.dout(n205),.clk(gclk));
	jnot g0142(.din(n205),.dout(n206),.clk(gclk));
	jand g0143(.dina(w_G273gat_5[1]),.dinb(w_G103gat_7[1]),.dout(n207),.clk(gclk));
	jcb g0144(.dina(w_n207_0[1]),.dinb(w_n168_0[0]),.dout(n208));
	jand g0145(.dina(w_G290gat_5[1]),.dinb(w_G103gat_7[0]),.dout(n209),.clk(gclk));
	jand g0146(.dina(w_n209_0[1]),.dinb(w_n166_0[0]),.dout(n210),.clk(gclk));
	jnot g0147(.din(w_n210_1[1]),.dout(n211),.clk(gclk));
	jand g0148(.dina(n211),.dinb(w_dff_B_csL5jpSV9_1),.dout(n212),.clk(gclk));
	jcb g0149(.dina(n212),.dinb(w_n169_0[0]),.dout(n213));
	jcb g0150(.dina(w_n210_1[0]),.dinb(w_n170_0[0]),.dout(n214));
	jand g0151(.dina(w_dff_B_uPKK8ESG8_0),.dinb(w_n213_0[1]),.dout(n215),.clk(gclk));
	jxor g0152(.dina(w_n215_0[1]),.dinb(w_n206_0[1]),.dout(n216),.clk(gclk));
	jxor g0153(.dina(w_n216_0[1]),.dinb(w_n204_0[1]),.dout(n217),.clk(gclk));
	jxor g0154(.dina(w_n217_0[1]),.dinb(w_n201_0[1]),.dout(n218),.clk(gclk));
	jxor g0155(.dina(w_n218_0[1]),.dinb(w_n199_0[1]),.dout(n219),.clk(gclk));
	jxor g0156(.dina(w_n219_0[1]),.dinb(w_n196_0[1]),.dout(n220),.clk(gclk));
	jnot g0157(.din(w_n220_0[1]),.dout(n221),.clk(gclk));
	jxor g0158(.dina(w_n221_0[1]),.dinb(w_n194_0[2]),.dout(n222),.clk(gclk));
	jxor g0159(.dina(n222),.dinb(w_dff_B_FeQGZ0tg2_1),.dout(n223),.clk(gclk));
	jxor g0160(.dina(w_n223_0[1]),.dinb(w_n188_0[1]),.dout(n224),.clk(gclk));
	jxor g0161(.dina(w_n224_0[1]),.dinb(w_dff_B_Sw83mtes0_1),.dout(G3211gat),.clk(gclk));
	jand g0162(.dina(w_G392gat_7[1]),.dinb(w_G1gat_5[0]),.dout(n226),.clk(gclk));
	jnot g0163(.din(w_n226_0[1]),.dout(n227),.clk(gclk));
	jnot g0164(.din(w_n223_0[0]),.dout(n228),.clk(gclk));
	jcb g0165(.dina(n228),.dinb(w_n188_0[0]),.dout(n229));
	jcb g0166(.dina(w_n224_0[0]),.dinb(w_n183_0[0]),.dout(n230));
	jand g0167(.dina(n230),.dinb(n229),.dout(n231),.clk(gclk));
	jand g0168(.dina(w_G375gat_7[0]),.dinb(w_G18gat_5[1]),.dout(n232),.clk(gclk));
	jnot g0169(.din(w_n232_0[1]),.dout(n233),.clk(gclk));
	jcb g0170(.dina(w_n221_0[0]),.dinb(w_n194_0[1]),.dout(n234));
	jxor g0171(.dina(w_n220_0[0]),.dinb(w_n194_0[0]),.dout(n235),.clk(gclk));
	jcb g0172(.dina(n235),.dinb(w_n189_0[0]),.dout(n236));
	jand g0173(.dina(n236),.dinb(n234),.dout(n237),.clk(gclk));
	jand g0174(.dina(w_G358gat_6[2]),.dinb(w_G35gat_5[2]),.dout(n238),.clk(gclk));
	jnot g0175(.din(n238),.dout(n239),.clk(gclk));
	jand g0176(.dina(w_n218_0[0]),.dinb(w_n199_0[0]),.dout(n240),.clk(gclk));
	jand g0177(.dina(w_n219_0[0]),.dinb(w_n196_0[0]),.dout(n241),.clk(gclk));
	jcb g0178(.dina(n241),.dinb(w_dff_B_bSS4JKmy4_1),.dout(n242));
	jand g0179(.dina(w_G341gat_6[1]),.dinb(w_G52gat_6[0]),.dout(n243),.clk(gclk));
	jnot g0180(.din(n243),.dout(n244),.clk(gclk));
	jand g0181(.dina(w_n216_0[0]),.dinb(w_n204_0[0]),.dout(n245),.clk(gclk));
	jand g0182(.dina(w_n217_0[0]),.dinb(w_n201_0[0]),.dout(n246),.clk(gclk));
	jcb g0183(.dina(n246),.dinb(w_dff_B_nwOQFSQ28_1),.dout(n247));
	jand g0184(.dina(w_G324gat_6[0]),.dinb(w_G69gat_6[1]),.dout(n248),.clk(gclk));
	jnot g0185(.din(n248),.dout(n249),.clk(gclk));
	jnot g0186(.din(w_n213_0[0]),.dout(n250),.clk(gclk));
	jand g0187(.dina(w_n215_0[0]),.dinb(w_n206_0[0]),.dout(n251),.clk(gclk));
	jcb g0188(.dina(n251),.dinb(w_dff_B_lXlV1jzs3_1),.dout(n252));
	jand g0189(.dina(w_G307gat_6[0]),.dinb(w_G86gat_6[2]),.dout(n253),.clk(gclk));
	jnot g0190(.din(n253),.dout(n254),.clk(gclk));
	jand g0191(.dina(w_G273gat_5[0]),.dinb(w_G120gat_7[1]),.dout(n255),.clk(gclk));
	jcb g0192(.dina(w_n255_0[1]),.dinb(w_n209_0[0]),.dout(n256));
	jand g0193(.dina(w_G290gat_5[0]),.dinb(w_G120gat_7[0]),.dout(n257),.clk(gclk));
	jand g0194(.dina(w_n257_0[1]),.dinb(w_n207_0[0]),.dout(n258),.clk(gclk));
	jnot g0195(.din(w_n258_0[2]),.dout(n259),.clk(gclk));
	jand g0196(.dina(w_n259_0[1]),.dinb(w_dff_B_nNWTPtOn8_1),.dout(n260),.clk(gclk));
	jcb g0197(.dina(n260),.dinb(w_n210_0[2]),.dout(n261));
	jand g0198(.dina(w_n259_0[0]),.dinb(w_n210_0[1]),.dout(n262),.clk(gclk));
	jnot g0199(.din(n262),.dout(n263),.clk(gclk));
	jand g0200(.dina(n263),.dinb(w_n261_0[1]),.dout(n264),.clk(gclk));
	jxor g0201(.dina(w_n264_0[1]),.dinb(w_n254_0[1]),.dout(n265),.clk(gclk));
	jxor g0202(.dina(w_n265_0[1]),.dinb(w_n252_0[1]),.dout(n266),.clk(gclk));
	jxor g0203(.dina(w_n266_0[1]),.dinb(w_n249_0[1]),.dout(n267),.clk(gclk));
	jxor g0204(.dina(w_n267_0[1]),.dinb(w_n247_0[1]),.dout(n268),.clk(gclk));
	jxor g0205(.dina(w_n268_0[1]),.dinb(w_n244_0[1]),.dout(n269),.clk(gclk));
	jxor g0206(.dina(w_n269_0[1]),.dinb(w_n242_0[1]),.dout(n270),.clk(gclk));
	jxor g0207(.dina(w_n270_0[1]),.dinb(w_n239_0[1]),.dout(n271),.clk(gclk));
	jnot g0208(.din(w_n271_0[1]),.dout(n272),.clk(gclk));
	jxor g0209(.dina(w_n272_0[1]),.dinb(w_n237_0[2]),.dout(n273),.clk(gclk));
	jxor g0210(.dina(n273),.dinb(w_dff_B_RUOdUyiF6_1),.dout(n274),.clk(gclk));
	jxor g0211(.dina(w_n274_0[1]),.dinb(w_n231_0[1]),.dout(n275),.clk(gclk));
	jxor g0212(.dina(w_n275_0[1]),.dinb(w_dff_B_4vAet7Rm0_1),.dout(G3552gat),.clk(gclk));
	jand g0213(.dina(w_G409gat_7[1]),.dinb(w_G1gat_4[2]),.dout(n277),.clk(gclk));
	jnot g0214(.din(w_n277_0[1]),.dout(n278),.clk(gclk));
	jnot g0215(.din(w_n274_0[0]),.dout(n279),.clk(gclk));
	jcb g0216(.dina(n279),.dinb(w_n231_0[0]),.dout(n280));
	jcb g0217(.dina(w_n275_0[0]),.dinb(w_n226_0[0]),.dout(n281));
	jand g0218(.dina(n281),.dinb(n280),.dout(n282),.clk(gclk));
	jand g0219(.dina(w_G392gat_7[0]),.dinb(w_G18gat_5[0]),.dout(n283),.clk(gclk));
	jnot g0220(.din(w_n283_0[1]),.dout(n284),.clk(gclk));
	jcb g0221(.dina(w_n272_0[0]),.dinb(w_n237_0[1]),.dout(n285));
	jxor g0222(.dina(w_n271_0[0]),.dinb(w_n237_0[0]),.dout(n286),.clk(gclk));
	jcb g0223(.dina(n286),.dinb(w_n232_0[0]),.dout(n287));
	jand g0224(.dina(n287),.dinb(n285),.dout(n288),.clk(gclk));
	jand g0225(.dina(w_G375gat_6[2]),.dinb(w_G35gat_5[1]),.dout(n289),.clk(gclk));
	jnot g0226(.din(n289),.dout(n290),.clk(gclk));
	jand g0227(.dina(w_n269_0[0]),.dinb(w_n242_0[0]),.dout(n291),.clk(gclk));
	jand g0228(.dina(w_n270_0[0]),.dinb(w_n239_0[0]),.dout(n292),.clk(gclk));
	jcb g0229(.dina(n292),.dinb(w_dff_B_Dk6URZcJ7_1),.dout(n293));
	jand g0230(.dina(w_G358gat_6[1]),.dinb(w_G52gat_5[2]),.dout(n294),.clk(gclk));
	jnot g0231(.din(n294),.dout(n295),.clk(gclk));
	jand g0232(.dina(w_n267_0[0]),.dinb(w_n247_0[0]),.dout(n296),.clk(gclk));
	jand g0233(.dina(w_n268_0[0]),.dinb(w_n244_0[0]),.dout(n297),.clk(gclk));
	jcb g0234(.dina(n297),.dinb(w_dff_B_ZVn1JATL0_1),.dout(n298));
	jand g0235(.dina(w_G341gat_6[0]),.dinb(w_G69gat_6[0]),.dout(n299),.clk(gclk));
	jnot g0236(.din(n299),.dout(n300),.clk(gclk));
	jand g0237(.dina(w_n265_0[0]),.dinb(w_n252_0[0]),.dout(n301),.clk(gclk));
	jand g0238(.dina(w_n266_0[0]),.dinb(w_n249_0[0]),.dout(n302),.clk(gclk));
	jcb g0239(.dina(n302),.dinb(w_dff_B_aRfMzHED9_1),.dout(n303));
	jand g0240(.dina(w_G324gat_5[2]),.dinb(w_G86gat_6[1]),.dout(n304),.clk(gclk));
	jnot g0241(.din(n304),.dout(n305),.clk(gclk));
	jnot g0242(.din(w_n261_0[0]),.dout(n306),.clk(gclk));
	jand g0243(.dina(w_n264_0[0]),.dinb(w_n254_0[0]),.dout(n307),.clk(gclk));
	jcb g0244(.dina(n307),.dinb(w_dff_B_y6wDHljS6_1),.dout(n308));
	jand g0245(.dina(w_G307gat_5[2]),.dinb(w_G103gat_6[2]),.dout(n309),.clk(gclk));
	jnot g0246(.din(n309),.dout(n310),.clk(gclk));
	jand g0247(.dina(w_G273gat_4[2]),.dinb(w_G137gat_7[1]),.dout(n311),.clk(gclk));
	jcb g0248(.dina(w_n311_0[1]),.dinb(w_n257_0[0]),.dout(n312));
	jand g0249(.dina(w_G290gat_4[2]),.dinb(w_G137gat_7[0]),.dout(n313),.clk(gclk));
	jand g0250(.dina(w_n313_0[1]),.dinb(w_n255_0[0]),.dout(n314),.clk(gclk));
	jnot g0251(.din(w_n314_0[2]),.dout(n315),.clk(gclk));
	jand g0252(.dina(w_n315_0[1]),.dinb(w_dff_B_1qBU2jhh6_1),.dout(n316),.clk(gclk));
	jcb g0253(.dina(n316),.dinb(w_n258_0[1]),.dout(n317));
	jand g0254(.dina(w_n315_0[0]),.dinb(w_n258_0[0]),.dout(n318),.clk(gclk));
	jnot g0255(.din(n318),.dout(n319),.clk(gclk));
	jand g0256(.dina(n319),.dinb(w_n317_0[1]),.dout(n320),.clk(gclk));
	jxor g0257(.dina(w_n320_0[1]),.dinb(w_n310_0[1]),.dout(n321),.clk(gclk));
	jxor g0258(.dina(w_n321_0[1]),.dinb(w_n308_0[1]),.dout(n322),.clk(gclk));
	jxor g0259(.dina(w_n322_0[1]),.dinb(w_n305_0[1]),.dout(n323),.clk(gclk));
	jxor g0260(.dina(w_n323_0[1]),.dinb(w_n303_0[1]),.dout(n324),.clk(gclk));
	jxor g0261(.dina(w_n324_0[1]),.dinb(w_n300_0[1]),.dout(n325),.clk(gclk));
	jxor g0262(.dina(w_n325_0[1]),.dinb(w_n298_0[1]),.dout(n326),.clk(gclk));
	jxor g0263(.dina(w_n326_0[1]),.dinb(w_n295_0[1]),.dout(n327),.clk(gclk));
	jxor g0264(.dina(w_n327_0[1]),.dinb(w_n293_0[1]),.dout(n328),.clk(gclk));
	jxor g0265(.dina(w_n328_0[1]),.dinb(w_n290_0[1]),.dout(n329),.clk(gclk));
	jnot g0266(.din(w_n329_0[1]),.dout(n330),.clk(gclk));
	jxor g0267(.dina(w_n330_0[1]),.dinb(w_n288_0[2]),.dout(n331),.clk(gclk));
	jxor g0268(.dina(n331),.dinb(w_dff_B_T7dveuQ82_1),.dout(n332),.clk(gclk));
	jxor g0269(.dina(w_n332_0[1]),.dinb(w_n282_0[1]),.dout(n333),.clk(gclk));
	jxor g0270(.dina(w_n333_0[1]),.dinb(w_dff_B_ckDZ6xwe5_1),.dout(G3895gat),.clk(gclk));
	jand g0271(.dina(w_G426gat_7[1]),.dinb(w_G1gat_4[1]),.dout(n335),.clk(gclk));
	jnot g0272(.din(w_n335_0[1]),.dout(n336),.clk(gclk));
	jnot g0273(.din(w_n332_0[0]),.dout(n337),.clk(gclk));
	jcb g0274(.dina(n337),.dinb(w_n282_0[0]),.dout(n338));
	jcb g0275(.dina(w_n333_0[0]),.dinb(w_n277_0[0]),.dout(n339));
	jand g0276(.dina(n339),.dinb(n338),.dout(n340),.clk(gclk));
	jand g0277(.dina(w_G409gat_7[0]),.dinb(w_G18gat_4[2]),.dout(n341),.clk(gclk));
	jnot g0278(.din(w_n341_0[1]),.dout(n342),.clk(gclk));
	jcb g0279(.dina(w_n330_0[0]),.dinb(w_n288_0[1]),.dout(n343));
	jxor g0280(.dina(w_n329_0[0]),.dinb(w_n288_0[0]),.dout(n344),.clk(gclk));
	jcb g0281(.dina(n344),.dinb(w_n283_0[0]),.dout(n345));
	jand g0282(.dina(n345),.dinb(n343),.dout(n346),.clk(gclk));
	jand g0283(.dina(w_G392gat_6[2]),.dinb(w_G35gat_5[0]),.dout(n347),.clk(gclk));
	jnot g0284(.din(n347),.dout(n348),.clk(gclk));
	jand g0285(.dina(w_n327_0[0]),.dinb(w_n293_0[0]),.dout(n349),.clk(gclk));
	jand g0286(.dina(w_n328_0[0]),.dinb(w_n290_0[0]),.dout(n350),.clk(gclk));
	jcb g0287(.dina(n350),.dinb(w_dff_B_mxWU2CBS8_1),.dout(n351));
	jand g0288(.dina(w_G375gat_6[1]),.dinb(w_G52gat_5[1]),.dout(n352),.clk(gclk));
	jnot g0289(.din(n352),.dout(n353),.clk(gclk));
	jand g0290(.dina(w_n325_0[0]),.dinb(w_n298_0[0]),.dout(n354),.clk(gclk));
	jand g0291(.dina(w_n326_0[0]),.dinb(w_n295_0[0]),.dout(n355),.clk(gclk));
	jcb g0292(.dina(n355),.dinb(w_dff_B_DwjbHO0w1_1),.dout(n356));
	jand g0293(.dina(w_G358gat_6[0]),.dinb(w_G69gat_5[2]),.dout(n357),.clk(gclk));
	jnot g0294(.din(n357),.dout(n358),.clk(gclk));
	jand g0295(.dina(w_n323_0[0]),.dinb(w_n303_0[0]),.dout(n359),.clk(gclk));
	jand g0296(.dina(w_n324_0[0]),.dinb(w_n300_0[0]),.dout(n360),.clk(gclk));
	jcb g0297(.dina(n360),.dinb(w_dff_B_Vv4HgKB73_1),.dout(n361));
	jand g0298(.dina(w_G341gat_5[2]),.dinb(w_G86gat_6[0]),.dout(n362),.clk(gclk));
	jnot g0299(.din(n362),.dout(n363),.clk(gclk));
	jand g0300(.dina(w_n321_0[0]),.dinb(w_n308_0[0]),.dout(n364),.clk(gclk));
	jand g0301(.dina(w_n322_0[0]),.dinb(w_n305_0[0]),.dout(n365),.clk(gclk));
	jcb g0302(.dina(n365),.dinb(w_dff_B_uosZhQmA9_1),.dout(n366));
	jand g0303(.dina(w_G324gat_5[1]),.dinb(w_G103gat_6[1]),.dout(n367),.clk(gclk));
	jnot g0304(.din(n367),.dout(n368),.clk(gclk));
	jnot g0305(.din(w_n317_0[0]),.dout(n369),.clk(gclk));
	jand g0306(.dina(w_n320_0[0]),.dinb(w_n310_0[0]),.dout(n370),.clk(gclk));
	jcb g0307(.dina(n370),.dinb(w_dff_B_YdACboNw3_1),.dout(n371));
	jand g0308(.dina(w_G307gat_5[1]),.dinb(w_G120gat_6[2]),.dout(n372),.clk(gclk));
	jand g0309(.dina(w_G273gat_4[1]),.dinb(w_G154gat_7[1]),.dout(n373),.clk(gclk));
	jcb g0310(.dina(w_n373_0[1]),.dinb(w_n313_0[0]),.dout(n374));
	jand g0311(.dina(w_G290gat_4[1]),.dinb(w_G154gat_7[0]),.dout(n375),.clk(gclk));
	jand g0312(.dina(w_n375_0[1]),.dinb(w_n311_0[0]),.dout(n376),.clk(gclk));
	jnot g0313(.din(w_n376_0[2]),.dout(n377),.clk(gclk));
	jand g0314(.dina(w_n377_0[1]),.dinb(w_dff_B_JAaSJxCS7_1),.dout(n378),.clk(gclk));
	jcb g0315(.dina(n378),.dinb(w_n314_0[1]),.dout(n379));
	jnot g0316(.din(n379),.dout(n380),.clk(gclk));
	jand g0317(.dina(w_n377_0[0]),.dinb(w_n314_0[0]),.dout(n381),.clk(gclk));
	jcb g0318(.dina(w_dff_B_5JXtGLp18_0),.dinb(w_n380_0[1]),.dout(n382));
	jxor g0319(.dina(w_n382_0[1]),.dinb(w_n372_0[1]),.dout(n383),.clk(gclk));
	jxor g0320(.dina(w_n383_0[1]),.dinb(w_n371_0[1]),.dout(n384),.clk(gclk));
	jxor g0321(.dina(w_n384_0[1]),.dinb(w_n368_0[1]),.dout(n385),.clk(gclk));
	jxor g0322(.dina(w_n385_0[1]),.dinb(w_n366_0[1]),.dout(n386),.clk(gclk));
	jxor g0323(.dina(w_n386_0[1]),.dinb(w_n363_0[1]),.dout(n387),.clk(gclk));
	jxor g0324(.dina(w_n387_0[1]),.dinb(w_n361_0[1]),.dout(n388),.clk(gclk));
	jxor g0325(.dina(w_n388_0[1]),.dinb(w_n358_0[1]),.dout(n389),.clk(gclk));
	jxor g0326(.dina(w_n389_0[1]),.dinb(w_n356_0[1]),.dout(n390),.clk(gclk));
	jxor g0327(.dina(w_n390_0[1]),.dinb(w_n353_0[1]),.dout(n391),.clk(gclk));
	jxor g0328(.dina(w_n391_0[1]),.dinb(w_n351_0[1]),.dout(n392),.clk(gclk));
	jxor g0329(.dina(w_n392_0[1]),.dinb(w_n348_0[1]),.dout(n393),.clk(gclk));
	jnot g0330(.din(w_n393_0[1]),.dout(n394),.clk(gclk));
	jxor g0331(.dina(w_n394_0[1]),.dinb(w_n346_0[2]),.dout(n395),.clk(gclk));
	jxor g0332(.dina(n395),.dinb(w_dff_B_uzgOcgVR6_1),.dout(n396),.clk(gclk));
	jxor g0333(.dina(w_n396_0[1]),.dinb(w_n340_0[1]),.dout(n397),.clk(gclk));
	jxor g0334(.dina(w_n397_0[1]),.dinb(w_dff_B_NUgGDnyd1_1),.dout(G4241gat),.clk(gclk));
	jand g0335(.dina(w_G443gat_7[1]),.dinb(w_G1gat_4[0]),.dout(n399),.clk(gclk));
	jnot g0336(.din(w_n399_0[1]),.dout(n400),.clk(gclk));
	jnot g0337(.din(w_n396_0[0]),.dout(n401),.clk(gclk));
	jcb g0338(.dina(n401),.dinb(w_n340_0[0]),.dout(n402));
	jcb g0339(.dina(w_n397_0[0]),.dinb(w_n335_0[0]),.dout(n403));
	jand g0340(.dina(n403),.dinb(n402),.dout(n404),.clk(gclk));
	jand g0341(.dina(w_G426gat_7[0]),.dinb(w_G18gat_4[1]),.dout(n405),.clk(gclk));
	jnot g0342(.din(w_n405_0[1]),.dout(n406),.clk(gclk));
	jcb g0343(.dina(w_n394_0[0]),.dinb(w_n346_0[1]),.dout(n407));
	jxor g0344(.dina(w_n393_0[0]),.dinb(w_n346_0[0]),.dout(n408),.clk(gclk));
	jcb g0345(.dina(n408),.dinb(w_n341_0[0]),.dout(n409));
	jand g0346(.dina(n409),.dinb(n407),.dout(n410),.clk(gclk));
	jand g0347(.dina(w_G409gat_6[2]),.dinb(w_G35gat_4[2]),.dout(n411),.clk(gclk));
	jnot g0348(.din(n411),.dout(n412),.clk(gclk));
	jand g0349(.dina(w_n391_0[0]),.dinb(w_n351_0[0]),.dout(n413),.clk(gclk));
	jand g0350(.dina(w_n392_0[0]),.dinb(w_n348_0[0]),.dout(n414),.clk(gclk));
	jcb g0351(.dina(n414),.dinb(w_dff_B_O4itNlQT3_1),.dout(n415));
	jand g0352(.dina(w_G392gat_6[1]),.dinb(w_G52gat_5[0]),.dout(n416),.clk(gclk));
	jnot g0353(.din(n416),.dout(n417),.clk(gclk));
	jand g0354(.dina(w_n389_0[0]),.dinb(w_n356_0[0]),.dout(n418),.clk(gclk));
	jand g0355(.dina(w_n390_0[0]),.dinb(w_n353_0[0]),.dout(n419),.clk(gclk));
	jcb g0356(.dina(n419),.dinb(w_dff_B_TIRuYEFC5_1),.dout(n420));
	jand g0357(.dina(w_G375gat_6[0]),.dinb(w_G69gat_5[1]),.dout(n421),.clk(gclk));
	jnot g0358(.din(n421),.dout(n422),.clk(gclk));
	jand g0359(.dina(w_n387_0[0]),.dinb(w_n361_0[0]),.dout(n423),.clk(gclk));
	jand g0360(.dina(w_n388_0[0]),.dinb(w_n358_0[0]),.dout(n424),.clk(gclk));
	jcb g0361(.dina(n424),.dinb(w_dff_B_yDwcpi3L2_1),.dout(n425));
	jand g0362(.dina(w_G358gat_5[2]),.dinb(w_G86gat_5[2]),.dout(n426),.clk(gclk));
	jnot g0363(.din(n426),.dout(n427),.clk(gclk));
	jand g0364(.dina(w_n385_0[0]),.dinb(w_n366_0[0]),.dout(n428),.clk(gclk));
	jand g0365(.dina(w_n386_0[0]),.dinb(w_n363_0[0]),.dout(n429),.clk(gclk));
	jcb g0366(.dina(n429),.dinb(w_dff_B_e5zG3G192_1),.dout(n430));
	jand g0367(.dina(w_G341gat_5[1]),.dinb(w_G103gat_6[0]),.dout(n431),.clk(gclk));
	jnot g0368(.din(n431),.dout(n432),.clk(gclk));
	jand g0369(.dina(w_n383_0[0]),.dinb(w_n371_0[0]),.dout(n433),.clk(gclk));
	jand g0370(.dina(w_n384_0[0]),.dinb(w_n368_0[0]),.dout(n434),.clk(gclk));
	jcb g0371(.dina(n434),.dinb(w_dff_B_jVyz4aVK1_1),.dout(n435));
	jand g0372(.dina(w_G324gat_5[0]),.dinb(w_G120gat_6[1]),.dout(n436),.clk(gclk));
	jnot g0373(.din(n436),.dout(n437),.clk(gclk));
	jnot g0374(.din(w_n372_0[0]),.dout(n438),.clk(gclk));
	jnot g0375(.din(w_n382_0[0]),.dout(n439),.clk(gclk));
	jand g0376(.dina(n439),.dinb(w_dff_B_hbzpAAfY3_1),.dout(n440),.clk(gclk));
	jcb g0377(.dina(n440),.dinb(w_n380_0[0]),.dout(n441));
	jand g0378(.dina(w_G307gat_5[0]),.dinb(w_G137gat_6[2]),.dout(n442),.clk(gclk));
	jand g0379(.dina(w_G273gat_4[0]),.dinb(w_G171gat_7[1]),.dout(n443),.clk(gclk));
	jcb g0380(.dina(w_n443_0[1]),.dinb(w_n375_0[0]),.dout(n444));
	jand g0381(.dina(w_G290gat_4[0]),.dinb(w_G171gat_7[0]),.dout(n445),.clk(gclk));
	jand g0382(.dina(w_n445_0[1]),.dinb(w_n373_0[0]),.dout(n446),.clk(gclk));
	jnot g0383(.din(w_n446_0[2]),.dout(n447),.clk(gclk));
	jand g0384(.dina(w_n447_0[1]),.dinb(w_dff_B_hW2Wvec32_1),.dout(n448),.clk(gclk));
	jcb g0385(.dina(n448),.dinb(w_n376_0[1]),.dout(n449));
	jnot g0386(.din(n449),.dout(n450),.clk(gclk));
	jand g0387(.dina(w_n447_0[0]),.dinb(w_n376_0[0]),.dout(n451),.clk(gclk));
	jcb g0388(.dina(w_dff_B_2vmf0QpN2_0),.dinb(w_n450_0[1]),.dout(n452));
	jxor g0389(.dina(w_n452_0[1]),.dinb(w_n442_0[1]),.dout(n453),.clk(gclk));
	jxor g0390(.dina(w_n453_0[1]),.dinb(w_n441_0[1]),.dout(n454),.clk(gclk));
	jxor g0391(.dina(w_n454_0[1]),.dinb(w_n437_0[1]),.dout(n455),.clk(gclk));
	jxor g0392(.dina(w_n455_0[1]),.dinb(w_n435_0[1]),.dout(n456),.clk(gclk));
	jxor g0393(.dina(w_n456_0[1]),.dinb(w_n432_0[1]),.dout(n457),.clk(gclk));
	jxor g0394(.dina(w_n457_0[1]),.dinb(w_n430_0[1]),.dout(n458),.clk(gclk));
	jxor g0395(.dina(w_n458_0[1]),.dinb(w_n427_0[1]),.dout(n459),.clk(gclk));
	jxor g0396(.dina(w_n459_0[1]),.dinb(w_n425_0[1]),.dout(n460),.clk(gclk));
	jxor g0397(.dina(w_n460_0[1]),.dinb(w_n422_0[1]),.dout(n461),.clk(gclk));
	jxor g0398(.dina(w_n461_0[1]),.dinb(w_n420_0[1]),.dout(n462),.clk(gclk));
	jxor g0399(.dina(w_n462_0[1]),.dinb(w_n417_0[1]),.dout(n463),.clk(gclk));
	jxor g0400(.dina(w_n463_0[1]),.dinb(w_n415_0[1]),.dout(n464),.clk(gclk));
	jxor g0401(.dina(w_n464_0[1]),.dinb(w_n412_0[1]),.dout(n465),.clk(gclk));
	jnot g0402(.din(w_n465_0[1]),.dout(n466),.clk(gclk));
	jxor g0403(.dina(w_n466_0[1]),.dinb(w_n410_0[2]),.dout(n467),.clk(gclk));
	jxor g0404(.dina(n467),.dinb(w_dff_B_E5IsYMmE0_1),.dout(n468),.clk(gclk));
	jxor g0405(.dina(w_n468_0[1]),.dinb(w_n404_0[1]),.dout(n469),.clk(gclk));
	jxor g0406(.dina(w_n469_0[1]),.dinb(w_dff_B_krulCJ8w6_1),.dout(G4591gat),.clk(gclk));
	jand g0407(.dina(w_G460gat_7[1]),.dinb(w_G1gat_3[2]),.dout(n471),.clk(gclk));
	jnot g0408(.din(w_n471_0[1]),.dout(n472),.clk(gclk));
	jnot g0409(.din(w_n468_0[0]),.dout(n473),.clk(gclk));
	jcb g0410(.dina(n473),.dinb(w_n404_0[0]),.dout(n474));
	jcb g0411(.dina(w_n469_0[0]),.dinb(w_n399_0[0]),.dout(n475));
	jand g0412(.dina(n475),.dinb(n474),.dout(n476),.clk(gclk));
	jand g0413(.dina(w_G443gat_7[0]),.dinb(w_G18gat_4[0]),.dout(n477),.clk(gclk));
	jnot g0414(.din(w_n477_0[1]),.dout(n478),.clk(gclk));
	jcb g0415(.dina(w_n466_0[0]),.dinb(w_n410_0[1]),.dout(n479));
	jxor g0416(.dina(w_n465_0[0]),.dinb(w_n410_0[0]),.dout(n480),.clk(gclk));
	jcb g0417(.dina(n480),.dinb(w_n405_0[0]),.dout(n481));
	jand g0418(.dina(n481),.dinb(n479),.dout(n482),.clk(gclk));
	jand g0419(.dina(w_G426gat_6[2]),.dinb(w_G35gat_4[1]),.dout(n483),.clk(gclk));
	jnot g0420(.din(n483),.dout(n484),.clk(gclk));
	jand g0421(.dina(w_n463_0[0]),.dinb(w_n415_0[0]),.dout(n485),.clk(gclk));
	jand g0422(.dina(w_n464_0[0]),.dinb(w_n412_0[0]),.dout(n486),.clk(gclk));
	jcb g0423(.dina(n486),.dinb(w_dff_B_qGJNeFyw7_1),.dout(n487));
	jand g0424(.dina(w_G409gat_6[1]),.dinb(w_G52gat_4[2]),.dout(n488),.clk(gclk));
	jnot g0425(.din(n488),.dout(n489),.clk(gclk));
	jand g0426(.dina(w_n461_0[0]),.dinb(w_n420_0[0]),.dout(n490),.clk(gclk));
	jand g0427(.dina(w_n462_0[0]),.dinb(w_n417_0[0]),.dout(n491),.clk(gclk));
	jcb g0428(.dina(n491),.dinb(w_dff_B_uYzApxJz9_1),.dout(n492));
	jand g0429(.dina(w_G392gat_6[0]),.dinb(w_G69gat_5[0]),.dout(n493),.clk(gclk));
	jnot g0430(.din(n493),.dout(n494),.clk(gclk));
	jand g0431(.dina(w_n459_0[0]),.dinb(w_n425_0[0]),.dout(n495),.clk(gclk));
	jand g0432(.dina(w_n460_0[0]),.dinb(w_n422_0[0]),.dout(n496),.clk(gclk));
	jcb g0433(.dina(n496),.dinb(w_dff_B_DXjHtJBZ6_1),.dout(n497));
	jand g0434(.dina(w_G375gat_5[2]),.dinb(w_G86gat_5[1]),.dout(n498),.clk(gclk));
	jnot g0435(.din(n498),.dout(n499),.clk(gclk));
	jand g0436(.dina(w_n457_0[0]),.dinb(w_n430_0[0]),.dout(n500),.clk(gclk));
	jand g0437(.dina(w_n458_0[0]),.dinb(w_n427_0[0]),.dout(n501),.clk(gclk));
	jcb g0438(.dina(n501),.dinb(w_dff_B_Bj9aSqi12_1),.dout(n502));
	jand g0439(.dina(w_G358gat_5[1]),.dinb(w_G103gat_5[2]),.dout(n503),.clk(gclk));
	jnot g0440(.din(n503),.dout(n504),.clk(gclk));
	jand g0441(.dina(w_n455_0[0]),.dinb(w_n435_0[0]),.dout(n505),.clk(gclk));
	jand g0442(.dina(w_n456_0[0]),.dinb(w_n432_0[0]),.dout(n506),.clk(gclk));
	jcb g0443(.dina(n506),.dinb(w_dff_B_dl8ogSlE8_1),.dout(n507));
	jand g0444(.dina(w_G341gat_5[0]),.dinb(w_G120gat_6[0]),.dout(n508),.clk(gclk));
	jnot g0445(.din(n508),.dout(n509),.clk(gclk));
	jand g0446(.dina(w_n453_0[0]),.dinb(w_n441_0[0]),.dout(n510),.clk(gclk));
	jand g0447(.dina(w_n454_0[0]),.dinb(w_n437_0[0]),.dout(n511),.clk(gclk));
	jcb g0448(.dina(n511),.dinb(w_dff_B_JGGGdc0n8_1),.dout(n512));
	jand g0449(.dina(w_G324gat_4[2]),.dinb(w_G137gat_6[1]),.dout(n513),.clk(gclk));
	jnot g0450(.din(n513),.dout(n514),.clk(gclk));
	jnot g0451(.din(w_n442_0[0]),.dout(n515),.clk(gclk));
	jnot g0452(.din(w_n452_0[0]),.dout(n516),.clk(gclk));
	jand g0453(.dina(n516),.dinb(w_dff_B_bQeuhAse3_1),.dout(n517),.clk(gclk));
	jcb g0454(.dina(n517),.dinb(w_n450_0[0]),.dout(n518));
	jand g0455(.dina(w_G307gat_4[2]),.dinb(w_G154gat_6[2]),.dout(n519),.clk(gclk));
	jand g0456(.dina(w_G273gat_3[2]),.dinb(w_G188gat_7[1]),.dout(n520),.clk(gclk));
	jcb g0457(.dina(w_n520_0[1]),.dinb(w_n445_0[0]),.dout(n521));
	jand g0458(.dina(w_G290gat_3[2]),.dinb(w_G188gat_7[0]),.dout(n522),.clk(gclk));
	jand g0459(.dina(w_n522_0[1]),.dinb(w_n443_0[0]),.dout(n523),.clk(gclk));
	jnot g0460(.din(w_n523_0[2]),.dout(n524),.clk(gclk));
	jand g0461(.dina(w_n524_0[1]),.dinb(w_dff_B_edoKP4GI5_1),.dout(n525),.clk(gclk));
	jcb g0462(.dina(n525),.dinb(w_n446_0[1]),.dout(n526));
	jnot g0463(.din(n526),.dout(n527),.clk(gclk));
	jand g0464(.dina(w_n524_0[0]),.dinb(w_n446_0[0]),.dout(n528),.clk(gclk));
	jcb g0465(.dina(w_dff_B_46YEwWPG7_0),.dinb(w_n527_0[1]),.dout(n529));
	jxor g0466(.dina(w_n529_0[1]),.dinb(w_n519_0[1]),.dout(n530),.clk(gclk));
	jxor g0467(.dina(w_n530_0[1]),.dinb(w_n518_0[1]),.dout(n531),.clk(gclk));
	jxor g0468(.dina(w_n531_0[1]),.dinb(w_n514_0[1]),.dout(n532),.clk(gclk));
	jxor g0469(.dina(w_n532_0[1]),.dinb(w_n512_0[1]),.dout(n533),.clk(gclk));
	jxor g0470(.dina(w_n533_0[1]),.dinb(w_n509_0[1]),.dout(n534),.clk(gclk));
	jxor g0471(.dina(w_n534_0[1]),.dinb(w_n507_0[1]),.dout(n535),.clk(gclk));
	jxor g0472(.dina(w_n535_0[1]),.dinb(w_n504_0[1]),.dout(n536),.clk(gclk));
	jxor g0473(.dina(w_n536_0[1]),.dinb(w_n502_0[1]),.dout(n537),.clk(gclk));
	jxor g0474(.dina(w_n537_0[1]),.dinb(w_n499_0[1]),.dout(n538),.clk(gclk));
	jxor g0475(.dina(w_n538_0[1]),.dinb(w_n497_0[1]),.dout(n539),.clk(gclk));
	jxor g0476(.dina(w_n539_0[1]),.dinb(w_n494_0[1]),.dout(n540),.clk(gclk));
	jxor g0477(.dina(w_n540_0[1]),.dinb(w_n492_0[1]),.dout(n541),.clk(gclk));
	jxor g0478(.dina(w_n541_0[1]),.dinb(w_n489_0[1]),.dout(n542),.clk(gclk));
	jxor g0479(.dina(w_n542_0[1]),.dinb(w_n487_0[1]),.dout(n543),.clk(gclk));
	jxor g0480(.dina(w_n543_0[1]),.dinb(w_n484_0[1]),.dout(n544),.clk(gclk));
	jnot g0481(.din(w_n544_0[1]),.dout(n545),.clk(gclk));
	jxor g0482(.dina(w_n545_0[1]),.dinb(w_n482_0[2]),.dout(n546),.clk(gclk));
	jxor g0483(.dina(n546),.dinb(w_dff_B_vTo9DWpq2_1),.dout(n547),.clk(gclk));
	jxor g0484(.dina(w_n547_0[1]),.dinb(w_n476_0[1]),.dout(n548),.clk(gclk));
	jxor g0485(.dina(w_n548_0[1]),.dinb(w_dff_B_YaDzBe1T8_1),.dout(G4946gat),.clk(gclk));
	jand g0486(.dina(w_G477gat_7[1]),.dinb(w_G1gat_3[1]),.dout(n550),.clk(gclk));
	jnot g0487(.din(w_n550_0[1]),.dout(n551),.clk(gclk));
	jnot g0488(.din(w_n547_0[0]),.dout(n552),.clk(gclk));
	jcb g0489(.dina(n552),.dinb(w_n476_0[0]),.dout(n553));
	jcb g0490(.dina(w_n548_0[0]),.dinb(w_n471_0[0]),.dout(n554));
	jand g0491(.dina(n554),.dinb(n553),.dout(n555),.clk(gclk));
	jand g0492(.dina(w_G460gat_7[0]),.dinb(w_G18gat_3[2]),.dout(n556),.clk(gclk));
	jnot g0493(.din(w_n556_0[1]),.dout(n557),.clk(gclk));
	jcb g0494(.dina(w_n545_0[0]),.dinb(w_n482_0[1]),.dout(n558));
	jxor g0495(.dina(w_n544_0[0]),.dinb(w_n482_0[0]),.dout(n559),.clk(gclk));
	jcb g0496(.dina(n559),.dinb(w_n477_0[0]),.dout(n560));
	jand g0497(.dina(n560),.dinb(n558),.dout(n561),.clk(gclk));
	jand g0498(.dina(w_G443gat_6[2]),.dinb(w_G35gat_4[0]),.dout(n562),.clk(gclk));
	jnot g0499(.din(n562),.dout(n563),.clk(gclk));
	jand g0500(.dina(w_n542_0[0]),.dinb(w_n487_0[0]),.dout(n564),.clk(gclk));
	jand g0501(.dina(w_n543_0[0]),.dinb(w_n484_0[0]),.dout(n565),.clk(gclk));
	jcb g0502(.dina(n565),.dinb(w_dff_B_mNrhr0kP7_1),.dout(n566));
	jand g0503(.dina(w_G426gat_6[1]),.dinb(w_G52gat_4[1]),.dout(n567),.clk(gclk));
	jnot g0504(.din(n567),.dout(n568),.clk(gclk));
	jand g0505(.dina(w_n540_0[0]),.dinb(w_n492_0[0]),.dout(n569),.clk(gclk));
	jand g0506(.dina(w_n541_0[0]),.dinb(w_n489_0[0]),.dout(n570),.clk(gclk));
	jcb g0507(.dina(n570),.dinb(w_dff_B_DADHk8B11_1),.dout(n571));
	jand g0508(.dina(w_G409gat_6[0]),.dinb(w_G69gat_4[2]),.dout(n572),.clk(gclk));
	jnot g0509(.din(n572),.dout(n573),.clk(gclk));
	jand g0510(.dina(w_n538_0[0]),.dinb(w_n497_0[0]),.dout(n574),.clk(gclk));
	jand g0511(.dina(w_n539_0[0]),.dinb(w_n494_0[0]),.dout(n575),.clk(gclk));
	jcb g0512(.dina(n575),.dinb(w_dff_B_KAUL5l4Y9_1),.dout(n576));
	jand g0513(.dina(w_G392gat_5[2]),.dinb(w_G86gat_5[0]),.dout(n577),.clk(gclk));
	jnot g0514(.din(n577),.dout(n578),.clk(gclk));
	jand g0515(.dina(w_n536_0[0]),.dinb(w_n502_0[0]),.dout(n579),.clk(gclk));
	jand g0516(.dina(w_n537_0[0]),.dinb(w_n499_0[0]),.dout(n580),.clk(gclk));
	jcb g0517(.dina(n580),.dinb(w_dff_B_Cn4ggaBf8_1),.dout(n581));
	jand g0518(.dina(w_G375gat_5[1]),.dinb(w_G103gat_5[1]),.dout(n582),.clk(gclk));
	jnot g0519(.din(n582),.dout(n583),.clk(gclk));
	jand g0520(.dina(w_n534_0[0]),.dinb(w_n507_0[0]),.dout(n584),.clk(gclk));
	jand g0521(.dina(w_n535_0[0]),.dinb(w_n504_0[0]),.dout(n585),.clk(gclk));
	jcb g0522(.dina(n585),.dinb(w_dff_B_QPvjEvrN3_1),.dout(n586));
	jand g0523(.dina(w_G358gat_5[0]),.dinb(w_G120gat_5[2]),.dout(n587),.clk(gclk));
	jnot g0524(.din(n587),.dout(n588),.clk(gclk));
	jand g0525(.dina(w_n532_0[0]),.dinb(w_n512_0[0]),.dout(n589),.clk(gclk));
	jand g0526(.dina(w_n533_0[0]),.dinb(w_n509_0[0]),.dout(n590),.clk(gclk));
	jcb g0527(.dina(n590),.dinb(w_dff_B_bs4LziED4_1),.dout(n591));
	jand g0528(.dina(w_G341gat_4[2]),.dinb(w_G137gat_6[0]),.dout(n592),.clk(gclk));
	jnot g0529(.din(n592),.dout(n593),.clk(gclk));
	jand g0530(.dina(w_n530_0[0]),.dinb(w_n518_0[0]),.dout(n594),.clk(gclk));
	jand g0531(.dina(w_n531_0[0]),.dinb(w_n514_0[0]),.dout(n595),.clk(gclk));
	jcb g0532(.dina(n595),.dinb(w_dff_B_Zo9yzJzN1_1),.dout(n596));
	jand g0533(.dina(w_G324gat_4[1]),.dinb(w_G154gat_6[1]),.dout(n597),.clk(gclk));
	jnot g0534(.din(n597),.dout(n598),.clk(gclk));
	jnot g0535(.din(w_n519_0[0]),.dout(n599),.clk(gclk));
	jnot g0536(.din(w_n529_0[0]),.dout(n600),.clk(gclk));
	jand g0537(.dina(n600),.dinb(w_dff_B_SinQdaEY4_1),.dout(n601),.clk(gclk));
	jcb g0538(.dina(n601),.dinb(w_n527_0[0]),.dout(n602));
	jand g0539(.dina(w_G307gat_4[1]),.dinb(w_G171gat_6[2]),.dout(n603),.clk(gclk));
	jand g0540(.dina(w_G273gat_3[1]),.dinb(w_G205gat_7[1]),.dout(n604),.clk(gclk));
	jcb g0541(.dina(w_n604_0[1]),.dinb(w_n522_0[0]),.dout(n605));
	jand g0542(.dina(w_G290gat_3[1]),.dinb(w_G205gat_7[0]),.dout(n606),.clk(gclk));
	jand g0543(.dina(w_n606_0[1]),.dinb(w_n520_0[0]),.dout(n607),.clk(gclk));
	jnot g0544(.din(w_n607_0[2]),.dout(n608),.clk(gclk));
	jand g0545(.dina(w_n608_0[1]),.dinb(w_dff_B_VBFHxlXZ9_1),.dout(n609),.clk(gclk));
	jcb g0546(.dina(n609),.dinb(w_n523_0[1]),.dout(n610));
	jnot g0547(.din(n610),.dout(n611),.clk(gclk));
	jand g0548(.dina(w_n608_0[0]),.dinb(w_n523_0[0]),.dout(n612),.clk(gclk));
	jcb g0549(.dina(w_dff_B_Gdn853Jj8_0),.dinb(w_n611_0[1]),.dout(n613));
	jxor g0550(.dina(w_n613_0[1]),.dinb(w_n603_0[1]),.dout(n614),.clk(gclk));
	jxor g0551(.dina(w_n614_0[1]),.dinb(w_n602_0[1]),.dout(n615),.clk(gclk));
	jxor g0552(.dina(w_n615_0[1]),.dinb(w_n598_0[1]),.dout(n616),.clk(gclk));
	jxor g0553(.dina(w_n616_0[1]),.dinb(w_n596_0[1]),.dout(n617),.clk(gclk));
	jxor g0554(.dina(w_n617_0[1]),.dinb(w_n593_0[1]),.dout(n618),.clk(gclk));
	jxor g0555(.dina(w_n618_0[1]),.dinb(w_n591_0[1]),.dout(n619),.clk(gclk));
	jxor g0556(.dina(w_n619_0[1]),.dinb(w_n588_0[1]),.dout(n620),.clk(gclk));
	jxor g0557(.dina(w_n620_0[1]),.dinb(w_n586_0[1]),.dout(n621),.clk(gclk));
	jxor g0558(.dina(w_n621_0[1]),.dinb(w_n583_0[1]),.dout(n622),.clk(gclk));
	jxor g0559(.dina(w_n622_0[1]),.dinb(w_n581_0[1]),.dout(n623),.clk(gclk));
	jxor g0560(.dina(w_n623_0[1]),.dinb(w_n578_0[1]),.dout(n624),.clk(gclk));
	jxor g0561(.dina(w_n624_0[1]),.dinb(w_n576_0[1]),.dout(n625),.clk(gclk));
	jxor g0562(.dina(w_n625_0[1]),.dinb(w_n573_0[1]),.dout(n626),.clk(gclk));
	jxor g0563(.dina(w_n626_0[1]),.dinb(w_n571_0[1]),.dout(n627),.clk(gclk));
	jxor g0564(.dina(w_n627_0[1]),.dinb(w_n568_0[1]),.dout(n628),.clk(gclk));
	jxor g0565(.dina(w_n628_0[1]),.dinb(w_n566_0[1]),.dout(n629),.clk(gclk));
	jxor g0566(.dina(w_n629_0[1]),.dinb(w_n563_0[1]),.dout(n630),.clk(gclk));
	jnot g0567(.din(w_n630_0[1]),.dout(n631),.clk(gclk));
	jxor g0568(.dina(w_n631_0[1]),.dinb(w_n561_0[2]),.dout(n632),.clk(gclk));
	jxor g0569(.dina(n632),.dinb(w_dff_B_Bid8kzJ10_1),.dout(n633),.clk(gclk));
	jxor g0570(.dina(w_n633_0[1]),.dinb(w_n555_0[1]),.dout(n634),.clk(gclk));
	jxor g0571(.dina(w_n634_0[1]),.dinb(w_dff_B_1YwacAhb1_1),.dout(G5308gat),.clk(gclk));
	jand g0572(.dina(w_G494gat_7[1]),.dinb(w_G1gat_3[0]),.dout(n636),.clk(gclk));
	jnot g0573(.din(w_n636_0[1]),.dout(n637),.clk(gclk));
	jnot g0574(.din(w_n633_0[0]),.dout(n638),.clk(gclk));
	jcb g0575(.dina(n638),.dinb(w_n555_0[0]),.dout(n639));
	jcb g0576(.dina(w_n634_0[0]),.dinb(w_n550_0[0]),.dout(n640));
	jand g0577(.dina(n640),.dinb(n639),.dout(n641),.clk(gclk));
	jand g0578(.dina(w_G477gat_7[0]),.dinb(w_G18gat_3[1]),.dout(n642),.clk(gclk));
	jnot g0579(.din(w_n642_0[1]),.dout(n643),.clk(gclk));
	jcb g0580(.dina(w_n631_0[0]),.dinb(w_n561_0[1]),.dout(n644));
	jxor g0581(.dina(w_n630_0[0]),.dinb(w_n561_0[0]),.dout(n645),.clk(gclk));
	jcb g0582(.dina(n645),.dinb(w_n556_0[0]),.dout(n646));
	jand g0583(.dina(n646),.dinb(n644),.dout(n647),.clk(gclk));
	jand g0584(.dina(w_G460gat_6[2]),.dinb(w_G35gat_3[2]),.dout(n648),.clk(gclk));
	jnot g0585(.din(n648),.dout(n649),.clk(gclk));
	jand g0586(.dina(w_n628_0[0]),.dinb(w_n566_0[0]),.dout(n650),.clk(gclk));
	jand g0587(.dina(w_n629_0[0]),.dinb(w_n563_0[0]),.dout(n651),.clk(gclk));
	jcb g0588(.dina(n651),.dinb(w_dff_B_Wmw0vaVP3_1),.dout(n652));
	jand g0589(.dina(w_G443gat_6[1]),.dinb(w_G52gat_4[0]),.dout(n653),.clk(gclk));
	jnot g0590(.din(n653),.dout(n654),.clk(gclk));
	jand g0591(.dina(w_n626_0[0]),.dinb(w_n571_0[0]),.dout(n655),.clk(gclk));
	jand g0592(.dina(w_n627_0[0]),.dinb(w_n568_0[0]),.dout(n656),.clk(gclk));
	jcb g0593(.dina(n656),.dinb(w_dff_B_uqn7ykRC9_1),.dout(n657));
	jand g0594(.dina(w_G426gat_6[0]),.dinb(w_G69gat_4[1]),.dout(n658),.clk(gclk));
	jnot g0595(.din(n658),.dout(n659),.clk(gclk));
	jand g0596(.dina(w_n624_0[0]),.dinb(w_n576_0[0]),.dout(n660),.clk(gclk));
	jand g0597(.dina(w_n625_0[0]),.dinb(w_n573_0[0]),.dout(n661),.clk(gclk));
	jcb g0598(.dina(n661),.dinb(w_dff_B_1cPflRMl6_1),.dout(n662));
	jand g0599(.dina(w_G409gat_5[2]),.dinb(w_G86gat_4[2]),.dout(n663),.clk(gclk));
	jnot g0600(.din(n663),.dout(n664),.clk(gclk));
	jand g0601(.dina(w_n622_0[0]),.dinb(w_n581_0[0]),.dout(n665),.clk(gclk));
	jand g0602(.dina(w_n623_0[0]),.dinb(w_n578_0[0]),.dout(n666),.clk(gclk));
	jcb g0603(.dina(n666),.dinb(w_dff_B_qIP4ZgBY5_1),.dout(n667));
	jand g0604(.dina(w_G392gat_5[1]),.dinb(w_G103gat_5[0]),.dout(n668),.clk(gclk));
	jnot g0605(.din(n668),.dout(n669),.clk(gclk));
	jand g0606(.dina(w_n620_0[0]),.dinb(w_n586_0[0]),.dout(n670),.clk(gclk));
	jand g0607(.dina(w_n621_0[0]),.dinb(w_n583_0[0]),.dout(n671),.clk(gclk));
	jcb g0608(.dina(n671),.dinb(w_dff_B_sqlWpZ4B1_1),.dout(n672));
	jand g0609(.dina(w_G375gat_5[0]),.dinb(w_G120gat_5[1]),.dout(n673),.clk(gclk));
	jnot g0610(.din(n673),.dout(n674),.clk(gclk));
	jand g0611(.dina(w_n618_0[0]),.dinb(w_n591_0[0]),.dout(n675),.clk(gclk));
	jand g0612(.dina(w_n619_0[0]),.dinb(w_n588_0[0]),.dout(n676),.clk(gclk));
	jcb g0613(.dina(n676),.dinb(w_dff_B_Y9rg3qgF9_1),.dout(n677));
	jand g0614(.dina(w_G358gat_4[2]),.dinb(w_G137gat_5[2]),.dout(n678),.clk(gclk));
	jnot g0615(.din(n678),.dout(n679),.clk(gclk));
	jand g0616(.dina(w_n616_0[0]),.dinb(w_n596_0[0]),.dout(n680),.clk(gclk));
	jand g0617(.dina(w_n617_0[0]),.dinb(w_n593_0[0]),.dout(n681),.clk(gclk));
	jcb g0618(.dina(n681),.dinb(w_dff_B_btSQe1sk0_1),.dout(n682));
	jand g0619(.dina(w_G341gat_4[1]),.dinb(w_G154gat_6[0]),.dout(n683),.clk(gclk));
	jnot g0620(.din(n683),.dout(n684),.clk(gclk));
	jand g0621(.dina(w_n614_0[0]),.dinb(w_n602_0[0]),.dout(n685),.clk(gclk));
	jand g0622(.dina(w_n615_0[0]),.dinb(w_n598_0[0]),.dout(n686),.clk(gclk));
	jcb g0623(.dina(n686),.dinb(w_dff_B_3bznItpR8_1),.dout(n687));
	jand g0624(.dina(w_G324gat_4[0]),.dinb(w_G171gat_6[1]),.dout(n688),.clk(gclk));
	jnot g0625(.din(n688),.dout(n689),.clk(gclk));
	jnot g0626(.din(w_n603_0[0]),.dout(n690),.clk(gclk));
	jnot g0627(.din(w_n613_0[0]),.dout(n691),.clk(gclk));
	jand g0628(.dina(n691),.dinb(w_dff_B_TCFaCcQC4_1),.dout(n692),.clk(gclk));
	jcb g0629(.dina(n692),.dinb(w_n611_0[0]),.dout(n693));
	jand g0630(.dina(w_G307gat_4[0]),.dinb(w_G188gat_6[2]),.dout(n694),.clk(gclk));
	jand g0631(.dina(w_G273gat_3[0]),.dinb(w_G222gat_7[1]),.dout(n695),.clk(gclk));
	jcb g0632(.dina(w_n695_0[2]),.dinb(w_n606_0[0]),.dout(n696));
	jand g0633(.dina(w_G290gat_3[0]),.dinb(w_G222gat_7[0]),.dout(n697),.clk(gclk));
	jand g0634(.dina(w_n697_0[1]),.dinb(w_n604_0[0]),.dout(n698),.clk(gclk));
	jnot g0635(.din(w_n698_0[2]),.dout(n699),.clk(gclk));
	jand g0636(.dina(w_n699_0[1]),.dinb(w_dff_B_YuHExj7R4_1),.dout(n700),.clk(gclk));
	jcb g0637(.dina(n700),.dinb(w_n607_0[1]),.dout(n701));
	jnot g0638(.din(n701),.dout(n702),.clk(gclk));
	jand g0639(.dina(w_n699_0[0]),.dinb(w_n607_0[0]),.dout(n703),.clk(gclk));
	jcb g0640(.dina(w_dff_B_D6eKyeyl8_0),.dinb(w_n702_0[1]),.dout(n704));
	jxor g0641(.dina(w_n704_0[1]),.dinb(w_n694_0[1]),.dout(n705),.clk(gclk));
	jxor g0642(.dina(w_n705_0[1]),.dinb(w_n693_0[1]),.dout(n706),.clk(gclk));
	jxor g0643(.dina(w_n706_0[1]),.dinb(w_n689_0[1]),.dout(n707),.clk(gclk));
	jxor g0644(.dina(w_n707_0[1]),.dinb(w_n687_0[1]),.dout(n708),.clk(gclk));
	jxor g0645(.dina(w_n708_0[1]),.dinb(w_n684_0[1]),.dout(n709),.clk(gclk));
	jxor g0646(.dina(w_n709_0[1]),.dinb(w_n682_0[1]),.dout(n710),.clk(gclk));
	jxor g0647(.dina(w_n710_0[1]),.dinb(w_n679_0[1]),.dout(n711),.clk(gclk));
	jxor g0648(.dina(w_n711_0[1]),.dinb(w_n677_0[1]),.dout(n712),.clk(gclk));
	jxor g0649(.dina(w_n712_0[1]),.dinb(w_n674_0[1]),.dout(n713),.clk(gclk));
	jxor g0650(.dina(w_n713_0[1]),.dinb(w_n672_0[1]),.dout(n714),.clk(gclk));
	jxor g0651(.dina(w_n714_0[1]),.dinb(w_n669_0[1]),.dout(n715),.clk(gclk));
	jxor g0652(.dina(w_n715_0[1]),.dinb(w_n667_0[1]),.dout(n716),.clk(gclk));
	jxor g0653(.dina(w_n716_0[1]),.dinb(w_n664_0[1]),.dout(n717),.clk(gclk));
	jxor g0654(.dina(w_n717_0[1]),.dinb(w_n662_0[1]),.dout(n718),.clk(gclk));
	jxor g0655(.dina(w_n718_0[1]),.dinb(w_n659_0[1]),.dout(n719),.clk(gclk));
	jxor g0656(.dina(w_n719_0[1]),.dinb(w_n657_0[1]),.dout(n720),.clk(gclk));
	jxor g0657(.dina(w_n720_0[1]),.dinb(w_n654_0[1]),.dout(n721),.clk(gclk));
	jxor g0658(.dina(w_n721_0[1]),.dinb(w_n652_0[1]),.dout(n722),.clk(gclk));
	jxor g0659(.dina(w_n722_0[1]),.dinb(w_n649_0[1]),.dout(n723),.clk(gclk));
	jnot g0660(.din(w_n723_0[1]),.dout(n724),.clk(gclk));
	jxor g0661(.dina(w_n724_0[1]),.dinb(w_n647_0[2]),.dout(n725),.clk(gclk));
	jxor g0662(.dina(n725),.dinb(w_dff_B_Y7kUWzNe8_1),.dout(n726),.clk(gclk));
	jxor g0663(.dina(w_n726_0[1]),.dinb(w_n641_0[1]),.dout(n727),.clk(gclk));
	jxor g0664(.dina(w_n727_0[1]),.dinb(w_dff_B_eX2PGYRO6_1),.dout(G5672gat),.clk(gclk));
	jand g0665(.dina(w_G511gat_7[1]),.dinb(w_G1gat_2[2]),.dout(n729),.clk(gclk));
	jnot g0666(.din(w_n729_0[1]),.dout(n730),.clk(gclk));
	jnot g0667(.din(w_n726_0[0]),.dout(n731),.clk(gclk));
	jcb g0668(.dina(n731),.dinb(w_n641_0[0]),.dout(n732));
	jcb g0669(.dina(w_n727_0[0]),.dinb(w_n636_0[0]),.dout(n733));
	jand g0670(.dina(n733),.dinb(n732),.dout(n734),.clk(gclk));
	jand g0671(.dina(w_G494gat_7[0]),.dinb(w_G18gat_3[0]),.dout(n735),.clk(gclk));
	jnot g0672(.din(w_n735_0[1]),.dout(n736),.clk(gclk));
	jcb g0673(.dina(w_n724_0[0]),.dinb(w_n647_0[1]),.dout(n737));
	jxor g0674(.dina(w_n723_0[0]),.dinb(w_n647_0[0]),.dout(n738),.clk(gclk));
	jcb g0675(.dina(n738),.dinb(w_n642_0[0]),.dout(n739));
	jand g0676(.dina(n739),.dinb(n737),.dout(n740),.clk(gclk));
	jand g0677(.dina(w_G477gat_6[2]),.dinb(w_G35gat_3[1]),.dout(n741),.clk(gclk));
	jnot g0678(.din(n741),.dout(n742),.clk(gclk));
	jand g0679(.dina(w_n721_0[0]),.dinb(w_n652_0[0]),.dout(n743),.clk(gclk));
	jand g0680(.dina(w_n722_0[0]),.dinb(w_n649_0[0]),.dout(n744),.clk(gclk));
	jcb g0681(.dina(n744),.dinb(w_dff_B_0jnZfbuD4_1),.dout(n745));
	jand g0682(.dina(w_G460gat_6[1]),.dinb(w_G52gat_3[2]),.dout(n746),.clk(gclk));
	jnot g0683(.din(n746),.dout(n747),.clk(gclk));
	jand g0684(.dina(w_n719_0[0]),.dinb(w_n657_0[0]),.dout(n748),.clk(gclk));
	jand g0685(.dina(w_n720_0[0]),.dinb(w_n654_0[0]),.dout(n749),.clk(gclk));
	jcb g0686(.dina(n749),.dinb(w_dff_B_NjSLxxAi9_1),.dout(n750));
	jand g0687(.dina(w_G443gat_6[0]),.dinb(w_G69gat_4[0]),.dout(n751),.clk(gclk));
	jnot g0688(.din(n751),.dout(n752),.clk(gclk));
	jand g0689(.dina(w_n717_0[0]),.dinb(w_n662_0[0]),.dout(n753),.clk(gclk));
	jand g0690(.dina(w_n718_0[0]),.dinb(w_n659_0[0]),.dout(n754),.clk(gclk));
	jcb g0691(.dina(n754),.dinb(w_dff_B_g5xYgFsp1_1),.dout(n755));
	jand g0692(.dina(w_G426gat_5[2]),.dinb(w_G86gat_4[1]),.dout(n756),.clk(gclk));
	jnot g0693(.din(n756),.dout(n757),.clk(gclk));
	jand g0694(.dina(w_n715_0[0]),.dinb(w_n667_0[0]),.dout(n758),.clk(gclk));
	jand g0695(.dina(w_n716_0[0]),.dinb(w_n664_0[0]),.dout(n759),.clk(gclk));
	jcb g0696(.dina(n759),.dinb(w_dff_B_AVYQgcJo9_1),.dout(n760));
	jand g0697(.dina(w_G409gat_5[1]),.dinb(w_G103gat_4[2]),.dout(n761),.clk(gclk));
	jnot g0698(.din(n761),.dout(n762),.clk(gclk));
	jand g0699(.dina(w_n713_0[0]),.dinb(w_n672_0[0]),.dout(n763),.clk(gclk));
	jand g0700(.dina(w_n714_0[0]),.dinb(w_n669_0[0]),.dout(n764),.clk(gclk));
	jcb g0701(.dina(n764),.dinb(w_dff_B_g8b86Sln6_1),.dout(n765));
	jand g0702(.dina(w_G392gat_5[0]),.dinb(w_G120gat_5[0]),.dout(n766),.clk(gclk));
	jnot g0703(.din(n766),.dout(n767),.clk(gclk));
	jand g0704(.dina(w_n711_0[0]),.dinb(w_n677_0[0]),.dout(n768),.clk(gclk));
	jand g0705(.dina(w_n712_0[0]),.dinb(w_n674_0[0]),.dout(n769),.clk(gclk));
	jcb g0706(.dina(n769),.dinb(w_dff_B_RZJNQvYs6_1),.dout(n770));
	jand g0707(.dina(w_G375gat_4[2]),.dinb(w_G137gat_5[1]),.dout(n771),.clk(gclk));
	jnot g0708(.din(n771),.dout(n772),.clk(gclk));
	jand g0709(.dina(w_n709_0[0]),.dinb(w_n682_0[0]),.dout(n773),.clk(gclk));
	jand g0710(.dina(w_n710_0[0]),.dinb(w_n679_0[0]),.dout(n774),.clk(gclk));
	jcb g0711(.dina(n774),.dinb(w_dff_B_uCF6h73s2_1),.dout(n775));
	jand g0712(.dina(w_G358gat_4[1]),.dinb(w_G154gat_5[2]),.dout(n776),.clk(gclk));
	jnot g0713(.din(n776),.dout(n777),.clk(gclk));
	jand g0714(.dina(w_n707_0[0]),.dinb(w_n687_0[0]),.dout(n778),.clk(gclk));
	jand g0715(.dina(w_n708_0[0]),.dinb(w_n684_0[0]),.dout(n779),.clk(gclk));
	jcb g0716(.dina(n779),.dinb(w_dff_B_9guddiw18_1),.dout(n780));
	jand g0717(.dina(w_G341gat_4[0]),.dinb(w_G171gat_6[0]),.dout(n781),.clk(gclk));
	jnot g0718(.din(n781),.dout(n782),.clk(gclk));
	jand g0719(.dina(w_n705_0[0]),.dinb(w_n693_0[0]),.dout(n783),.clk(gclk));
	jand g0720(.dina(w_n706_0[0]),.dinb(w_n689_0[0]),.dout(n784),.clk(gclk));
	jcb g0721(.dina(n784),.dinb(w_dff_B_m2N89aZe5_1),.dout(n785));
	jand g0722(.dina(w_G324gat_3[2]),.dinb(w_G188gat_6[1]),.dout(n786),.clk(gclk));
	jnot g0723(.din(n786),.dout(n787),.clk(gclk));
	jnot g0724(.din(w_n694_0[0]),.dout(n788),.clk(gclk));
	jnot g0725(.din(w_n704_0[0]),.dout(n789),.clk(gclk));
	jand g0726(.dina(n789),.dinb(w_dff_B_WYYKT4UZ3_1),.dout(n790),.clk(gclk));
	jcb g0727(.dina(n790),.dinb(w_n702_0[0]),.dout(n791));
	jand g0728(.dina(w_G307gat_3[2]),.dinb(w_G205gat_6[2]),.dout(n792),.clk(gclk));
	jand g0729(.dina(w_G273gat_2[2]),.dinb(w_G239gat_7[1]),.dout(n793),.clk(gclk));
	jcb g0730(.dina(w_n793_0[1]),.dinb(w_n697_0[0]),.dout(n794));
	jand g0731(.dina(w_G290gat_2[2]),.dinb(w_G239gat_7[0]),.dout(n795),.clk(gclk));
	jand g0732(.dina(w_n795_0[1]),.dinb(w_n695_0[1]),.dout(n796),.clk(gclk));
	jnot g0733(.din(n796),.dout(n797),.clk(gclk));
	jand g0734(.dina(w_n797_0[2]),.dinb(w_dff_B_3R5BpVwG3_1),.dout(n798),.clk(gclk));
	jcb g0735(.dina(n798),.dinb(w_n698_0[1]),.dout(n799));
	jnot g0736(.din(n799),.dout(n800),.clk(gclk));
	jand g0737(.dina(w_n797_0[1]),.dinb(w_n698_0[0]),.dout(n801),.clk(gclk));
	jcb g0738(.dina(w_dff_B_LuvGROLa3_0),.dinb(w_n800_0[1]),.dout(n802));
	jxor g0739(.dina(w_n802_0[1]),.dinb(w_n792_0[1]),.dout(n803),.clk(gclk));
	jxor g0740(.dina(w_n803_0[1]),.dinb(w_n791_0[1]),.dout(n804),.clk(gclk));
	jxor g0741(.dina(w_n804_0[1]),.dinb(w_n787_0[1]),.dout(n805),.clk(gclk));
	jxor g0742(.dina(w_n805_0[1]),.dinb(w_n785_0[1]),.dout(n806),.clk(gclk));
	jxor g0743(.dina(w_n806_0[1]),.dinb(w_n782_0[1]),.dout(n807),.clk(gclk));
	jxor g0744(.dina(w_n807_0[1]),.dinb(w_n780_0[1]),.dout(n808),.clk(gclk));
	jxor g0745(.dina(w_n808_0[1]),.dinb(w_n777_0[1]),.dout(n809),.clk(gclk));
	jxor g0746(.dina(w_n809_0[1]),.dinb(w_n775_0[1]),.dout(n810),.clk(gclk));
	jxor g0747(.dina(w_n810_0[1]),.dinb(w_n772_0[1]),.dout(n811),.clk(gclk));
	jxor g0748(.dina(w_n811_0[1]),.dinb(w_n770_0[1]),.dout(n812),.clk(gclk));
	jxor g0749(.dina(w_n812_0[1]),.dinb(w_n767_0[1]),.dout(n813),.clk(gclk));
	jxor g0750(.dina(w_n813_0[1]),.dinb(w_n765_0[1]),.dout(n814),.clk(gclk));
	jxor g0751(.dina(w_n814_0[1]),.dinb(w_n762_0[1]),.dout(n815),.clk(gclk));
	jxor g0752(.dina(w_n815_0[1]),.dinb(w_n760_0[1]),.dout(n816),.clk(gclk));
	jxor g0753(.dina(w_n816_0[1]),.dinb(w_n757_0[1]),.dout(n817),.clk(gclk));
	jxor g0754(.dina(w_n817_0[1]),.dinb(w_n755_0[1]),.dout(n818),.clk(gclk));
	jxor g0755(.dina(w_n818_0[1]),.dinb(w_n752_0[1]),.dout(n819),.clk(gclk));
	jxor g0756(.dina(w_n819_0[1]),.dinb(w_n750_0[1]),.dout(n820),.clk(gclk));
	jxor g0757(.dina(w_n820_0[1]),.dinb(w_n747_0[1]),.dout(n821),.clk(gclk));
	jxor g0758(.dina(w_n821_0[1]),.dinb(w_n745_0[1]),.dout(n822),.clk(gclk));
	jxor g0759(.dina(w_n822_0[1]),.dinb(w_n742_0[1]),.dout(n823),.clk(gclk));
	jnot g0760(.din(w_n823_0[1]),.dout(n824),.clk(gclk));
	jxor g0761(.dina(w_n824_0[1]),.dinb(w_n740_0[2]),.dout(n825),.clk(gclk));
	jxor g0762(.dina(n825),.dinb(w_dff_B_xftUq9QE4_1),.dout(n826),.clk(gclk));
	jxor g0763(.dina(w_n826_0[1]),.dinb(w_n734_0[1]),.dout(n827),.clk(gclk));
	jxor g0764(.dina(w_n827_0[1]),.dinb(w_dff_B_aoYzFfpI1_1),.dout(G5971gat),.clk(gclk));
	jand g0765(.dina(w_G528gat_7[1]),.dinb(w_G1gat_2[1]),.dout(n829),.clk(gclk));
	jnot g0766(.din(w_n829_0[1]),.dout(n830),.clk(gclk));
	jnot g0767(.din(w_n826_0[0]),.dout(n831),.clk(gclk));
	jcb g0768(.dina(n831),.dinb(w_n734_0[0]),.dout(n832));
	jcb g0769(.dina(w_n827_0[0]),.dinb(w_n729_0[0]),.dout(n833));
	jand g0770(.dina(n833),.dinb(n832),.dout(n834),.clk(gclk));
	jand g0771(.dina(w_G511gat_7[0]),.dinb(w_G18gat_2[2]),.dout(n835),.clk(gclk));
	jcb g0772(.dina(w_n824_0[0]),.dinb(w_n740_0[1]),.dout(n836));
	jxor g0773(.dina(w_n823_0[0]),.dinb(w_n740_0[0]),.dout(n837),.clk(gclk));
	jcb g0774(.dina(n837),.dinb(w_n735_0[0]),.dout(n838));
	jand g0775(.dina(n838),.dinb(n836),.dout(n839),.clk(gclk));
	jand g0776(.dina(w_G494gat_6[2]),.dinb(w_G35gat_3[0]),.dout(n840),.clk(gclk));
	jnot g0777(.din(w_n840_0[1]),.dout(n841),.clk(gclk));
	jand g0778(.dina(w_n821_0[0]),.dinb(w_n745_0[0]),.dout(n842),.clk(gclk));
	jand g0779(.dina(w_n822_0[0]),.dinb(w_n742_0[0]),.dout(n843),.clk(gclk));
	jcb g0780(.dina(n843),.dinb(w_dff_B_tdhjsvxw5_1),.dout(n844));
	jand g0781(.dina(w_G477gat_6[1]),.dinb(w_G52gat_3[1]),.dout(n845),.clk(gclk));
	jnot g0782(.din(n845),.dout(n846),.clk(gclk));
	jand g0783(.dina(w_n819_0[0]),.dinb(w_n750_0[0]),.dout(n847),.clk(gclk));
	jand g0784(.dina(w_n820_0[0]),.dinb(w_n747_0[0]),.dout(n848),.clk(gclk));
	jcb g0785(.dina(n848),.dinb(w_dff_B_jan9yoBt7_1),.dout(n849));
	jand g0786(.dina(w_G460gat_6[0]),.dinb(w_G69gat_3[2]),.dout(n850),.clk(gclk));
	jnot g0787(.din(n850),.dout(n851),.clk(gclk));
	jand g0788(.dina(w_n817_0[0]),.dinb(w_n755_0[0]),.dout(n852),.clk(gclk));
	jand g0789(.dina(w_n818_0[0]),.dinb(w_n752_0[0]),.dout(n853),.clk(gclk));
	jcb g0790(.dina(n853),.dinb(w_dff_B_xYzFwxws2_1),.dout(n854));
	jand g0791(.dina(w_G443gat_5[2]),.dinb(w_G86gat_4[0]),.dout(n855),.clk(gclk));
	jnot g0792(.din(n855),.dout(n856),.clk(gclk));
	jand g0793(.dina(w_n815_0[0]),.dinb(w_n760_0[0]),.dout(n857),.clk(gclk));
	jand g0794(.dina(w_n816_0[0]),.dinb(w_n757_0[0]),.dout(n858),.clk(gclk));
	jcb g0795(.dina(n858),.dinb(w_dff_B_4KcQbGzm1_1),.dout(n859));
	jand g0796(.dina(w_G426gat_5[1]),.dinb(w_G103gat_4[1]),.dout(n860),.clk(gclk));
	jnot g0797(.din(n860),.dout(n861),.clk(gclk));
	jand g0798(.dina(w_n813_0[0]),.dinb(w_n765_0[0]),.dout(n862),.clk(gclk));
	jand g0799(.dina(w_n814_0[0]),.dinb(w_n762_0[0]),.dout(n863),.clk(gclk));
	jcb g0800(.dina(n863),.dinb(w_dff_B_v6EO7e6d1_1),.dout(n864));
	jand g0801(.dina(w_G409gat_5[0]),.dinb(w_G120gat_4[2]),.dout(n865),.clk(gclk));
	jnot g0802(.din(n865),.dout(n866),.clk(gclk));
	jand g0803(.dina(w_n811_0[0]),.dinb(w_n770_0[0]),.dout(n867),.clk(gclk));
	jand g0804(.dina(w_n812_0[0]),.dinb(w_n767_0[0]),.dout(n868),.clk(gclk));
	jcb g0805(.dina(n868),.dinb(w_dff_B_YeF2aOoA8_1),.dout(n869));
	jand g0806(.dina(w_G392gat_4[2]),.dinb(w_G137gat_5[0]),.dout(n870),.clk(gclk));
	jnot g0807(.din(n870),.dout(n871),.clk(gclk));
	jand g0808(.dina(w_n809_0[0]),.dinb(w_n775_0[0]),.dout(n872),.clk(gclk));
	jand g0809(.dina(w_n810_0[0]),.dinb(w_n772_0[0]),.dout(n873),.clk(gclk));
	jcb g0810(.dina(n873),.dinb(w_dff_B_Z1wAO6IW1_1),.dout(n874));
	jand g0811(.dina(w_G375gat_4[1]),.dinb(w_G154gat_5[1]),.dout(n875),.clk(gclk));
	jnot g0812(.din(n875),.dout(n876),.clk(gclk));
	jand g0813(.dina(w_n807_0[0]),.dinb(w_n780_0[0]),.dout(n877),.clk(gclk));
	jand g0814(.dina(w_n808_0[0]),.dinb(w_n777_0[0]),.dout(n878),.clk(gclk));
	jcb g0815(.dina(n878),.dinb(w_dff_B_yZPdh5aS0_1),.dout(n879));
	jand g0816(.dina(w_G358gat_4[0]),.dinb(w_G171gat_5[2]),.dout(n880),.clk(gclk));
	jnot g0817(.din(n880),.dout(n881),.clk(gclk));
	jand g0818(.dina(w_n805_0[0]),.dinb(w_n785_0[0]),.dout(n882),.clk(gclk));
	jand g0819(.dina(w_n806_0[0]),.dinb(w_n782_0[0]),.dout(n883),.clk(gclk));
	jcb g0820(.dina(n883),.dinb(w_dff_B_39ySnxDb3_1),.dout(n884));
	jand g0821(.dina(w_G341gat_3[2]),.dinb(w_G188gat_6[0]),.dout(n885),.clk(gclk));
	jnot g0822(.din(n885),.dout(n886),.clk(gclk));
	jand g0823(.dina(w_n803_0[0]),.dinb(w_n791_0[0]),.dout(n887),.clk(gclk));
	jand g0824(.dina(w_n804_0[0]),.dinb(w_n787_0[0]),.dout(n888),.clk(gclk));
	jcb g0825(.dina(n888),.dinb(w_dff_B_pITryFcZ5_1),.dout(n889));
	jand g0826(.dina(w_G324gat_3[1]),.dinb(w_G205gat_6[1]),.dout(n890),.clk(gclk));
	jnot g0827(.din(n890),.dout(n891),.clk(gclk));
	jnot g0828(.din(w_n792_0[0]),.dout(n892),.clk(gclk));
	jnot g0829(.din(w_n802_0[0]),.dout(n893),.clk(gclk));
	jand g0830(.dina(n893),.dinb(w_dff_B_VI7ITJyG6_1),.dout(n894),.clk(gclk));
	jcb g0831(.dina(n894),.dinb(w_n800_0[0]),.dout(n895));
	jand g0832(.dina(w_G307gat_3[1]),.dinb(w_G222gat_6[2]),.dout(n896),.clk(gclk));
	jnot g0833(.din(w_n795_0[0]),.dout(n897),.clk(gclk));
	jand g0834(.dina(w_G273gat_2[1]),.dinb(w_G256gat_7[1]),.dout(n898),.clk(gclk));
	jand g0835(.dina(w_n898_0[1]),.dinb(w_n897_0[1]),.dout(n899),.clk(gclk));
	jnot g0836(.din(n899),.dout(n900),.clk(gclk));
	jcb g0837(.dina(w_n898_0[0]),.dinb(w_n897_0[0]),.dout(n901));
	jand g0838(.dina(w_n901_0[1]),.dinb(w_n797_0[0]),.dout(n902),.clk(gclk));
	jand g0839(.dina(n902),.dinb(n900),.dout(n903),.clk(gclk));
	jnot g0840(.din(w_n901_0[0]),.dout(n904),.clk(gclk));
	jand g0841(.dina(n904),.dinb(w_n695_0[0]),.dout(n905),.clk(gclk));
	jcb g0842(.dina(w_dff_B_rAaU6uUB6_0),.dinb(w_n903_0[1]),.dout(n906));
	jxor g0843(.dina(w_n906_0[1]),.dinb(w_n896_0[1]),.dout(n907),.clk(gclk));
	jxor g0844(.dina(w_n907_0[1]),.dinb(w_n895_0[1]),.dout(n908),.clk(gclk));
	jxor g0845(.dina(w_n908_0[1]),.dinb(w_n891_0[1]),.dout(n909),.clk(gclk));
	jxor g0846(.dina(w_n909_0[1]),.dinb(w_n889_0[1]),.dout(n910),.clk(gclk));
	jxor g0847(.dina(w_n910_0[1]),.dinb(w_n886_0[1]),.dout(n911),.clk(gclk));
	jxor g0848(.dina(w_n911_0[1]),.dinb(w_n884_0[1]),.dout(n912),.clk(gclk));
	jxor g0849(.dina(w_n912_0[1]),.dinb(w_n881_0[1]),.dout(n913),.clk(gclk));
	jxor g0850(.dina(w_n913_0[1]),.dinb(w_n879_0[1]),.dout(n914),.clk(gclk));
	jxor g0851(.dina(w_n914_0[1]),.dinb(w_n876_0[1]),.dout(n915),.clk(gclk));
	jxor g0852(.dina(w_n915_0[1]),.dinb(w_n874_0[1]),.dout(n916),.clk(gclk));
	jxor g0853(.dina(w_n916_0[1]),.dinb(w_n871_0[1]),.dout(n917),.clk(gclk));
	jxor g0854(.dina(w_n917_0[1]),.dinb(w_n869_0[1]),.dout(n918),.clk(gclk));
	jxor g0855(.dina(w_n918_0[1]),.dinb(w_n866_0[1]),.dout(n919),.clk(gclk));
	jxor g0856(.dina(w_n919_0[1]),.dinb(w_n864_0[1]),.dout(n920),.clk(gclk));
	jxor g0857(.dina(w_n920_0[1]),.dinb(w_n861_0[1]),.dout(n921),.clk(gclk));
	jxor g0858(.dina(w_n921_0[1]),.dinb(w_n859_0[1]),.dout(n922),.clk(gclk));
	jxor g0859(.dina(w_n922_0[1]),.dinb(w_n856_0[1]),.dout(n923),.clk(gclk));
	jxor g0860(.dina(w_n923_0[1]),.dinb(w_n854_0[1]),.dout(n924),.clk(gclk));
	jxor g0861(.dina(w_n924_0[1]),.dinb(w_n851_0[1]),.dout(n925),.clk(gclk));
	jxor g0862(.dina(w_n925_0[1]),.dinb(w_n849_0[1]),.dout(n926),.clk(gclk));
	jxor g0863(.dina(w_n926_0[1]),.dinb(w_n846_0[1]),.dout(n927),.clk(gclk));
	jxor g0864(.dina(w_n927_0[2]),.dinb(w_n844_0[2]),.dout(n928),.clk(gclk));
	jxor g0865(.dina(n928),.dinb(w_dff_B_GNqgMNCd9_1),.dout(n929),.clk(gclk));
	jxor g0866(.dina(w_n929_0[1]),.dinb(w_n839_0[1]),.dout(n930),.clk(gclk));
	jxor g0867(.dina(w_n930_0[1]),.dinb(w_n835_0[1]),.dout(n931),.clk(gclk));
	jxor g0868(.dina(w_n931_0[1]),.dinb(w_n834_0[1]),.dout(n932),.clk(gclk));
	jxor g0869(.dina(w_n932_0[1]),.dinb(w_dff_B_E6U2roQ78_1),.dout(G6123gat),.clk(gclk));
	jnot g0870(.din(w_n931_0[0]),.dout(n934),.clk(gclk));
	jcb g0871(.dina(n934),.dinb(w_n834_0[0]),.dout(n935));
	jcb g0872(.dina(w_n932_0[0]),.dinb(w_n829_0[0]),.dout(n936));
	jand g0873(.dina(n936),.dinb(w_dff_B_BJ8Cjrj89_1),.dout(n937),.clk(gclk));
	jand g0874(.dina(w_G528gat_7[0]),.dinb(w_G18gat_2[1]),.dout(n938),.clk(gclk));
	jnot g0875(.din(w_n929_0[0]),.dout(n939),.clk(gclk));
	jcb g0876(.dina(n939),.dinb(w_n839_0[0]),.dout(n940));
	jcb g0877(.dina(w_n930_0[0]),.dinb(w_n835_0[0]),.dout(n941));
	jand g0878(.dina(n941),.dinb(n940),.dout(n942),.clk(gclk));
	jand g0879(.dina(w_G511gat_6[2]),.dinb(w_G35gat_2[2]),.dout(n943),.clk(gclk));
	jand g0880(.dina(w_n927_0[1]),.dinb(w_n844_0[1]),.dout(n944),.clk(gclk));
	jnot g0881(.din(n944),.dout(n945),.clk(gclk));
	jnot g0882(.din(w_n927_0[0]),.dout(n946),.clk(gclk));
	jxor g0883(.dina(n946),.dinb(w_n844_0[0]),.dout(n947),.clk(gclk));
	jcb g0884(.dina(n947),.dinb(w_n840_0[0]),.dout(n948));
	jand g0885(.dina(n948),.dinb(n945),.dout(n949),.clk(gclk));
	jand g0886(.dina(w_G494gat_6[1]),.dinb(w_G52gat_3[0]),.dout(n950),.clk(gclk));
	jnot g0887(.din(n950),.dout(n951),.clk(gclk));
	jand g0888(.dina(w_n925_0[0]),.dinb(w_n849_0[0]),.dout(n952),.clk(gclk));
	jand g0889(.dina(w_n926_0[0]),.dinb(w_n846_0[0]),.dout(n953),.clk(gclk));
	jcb g0890(.dina(n953),.dinb(w_dff_B_BbhDxqc18_1),.dout(n954));
	jand g0891(.dina(w_G477gat_6[0]),.dinb(w_G69gat_3[1]),.dout(n955),.clk(gclk));
	jnot g0892(.din(n955),.dout(n956),.clk(gclk));
	jand g0893(.dina(w_n923_0[0]),.dinb(w_n854_0[0]),.dout(n957),.clk(gclk));
	jand g0894(.dina(w_n924_0[0]),.dinb(w_n851_0[0]),.dout(n958),.clk(gclk));
	jcb g0895(.dina(n958),.dinb(w_dff_B_W5g7uig16_1),.dout(n959));
	jand g0896(.dina(w_G460gat_5[2]),.dinb(w_G86gat_3[2]),.dout(n960),.clk(gclk));
	jnot g0897(.din(n960),.dout(n961),.clk(gclk));
	jand g0898(.dina(w_n921_0[0]),.dinb(w_n859_0[0]),.dout(n962),.clk(gclk));
	jand g0899(.dina(w_n922_0[0]),.dinb(w_n856_0[0]),.dout(n963),.clk(gclk));
	jcb g0900(.dina(n963),.dinb(w_dff_B_3TmBEJSr7_1),.dout(n964));
	jand g0901(.dina(w_G443gat_5[1]),.dinb(w_G103gat_4[0]),.dout(n965),.clk(gclk));
	jnot g0902(.din(n965),.dout(n966),.clk(gclk));
	jand g0903(.dina(w_n919_0[0]),.dinb(w_n864_0[0]),.dout(n967),.clk(gclk));
	jand g0904(.dina(w_n920_0[0]),.dinb(w_n861_0[0]),.dout(n968),.clk(gclk));
	jcb g0905(.dina(n968),.dinb(w_dff_B_KUz0OnNt7_1),.dout(n969));
	jand g0906(.dina(w_G426gat_5[0]),.dinb(w_G120gat_4[1]),.dout(n970),.clk(gclk));
	jnot g0907(.din(n970),.dout(n971),.clk(gclk));
	jand g0908(.dina(w_n917_0[0]),.dinb(w_n869_0[0]),.dout(n972),.clk(gclk));
	jand g0909(.dina(w_n918_0[0]),.dinb(w_n866_0[0]),.dout(n973),.clk(gclk));
	jcb g0910(.dina(n973),.dinb(w_dff_B_yxOlFviZ9_1),.dout(n974));
	jand g0911(.dina(w_G409gat_4[2]),.dinb(w_G137gat_4[2]),.dout(n975),.clk(gclk));
	jnot g0912(.din(n975),.dout(n976),.clk(gclk));
	jand g0913(.dina(w_n915_0[0]),.dinb(w_n874_0[0]),.dout(n977),.clk(gclk));
	jand g0914(.dina(w_n916_0[0]),.dinb(w_n871_0[0]),.dout(n978),.clk(gclk));
	jcb g0915(.dina(n978),.dinb(w_dff_B_4OhSnjHB1_1),.dout(n979));
	jand g0916(.dina(w_G392gat_4[1]),.dinb(w_G154gat_5[0]),.dout(n980),.clk(gclk));
	jnot g0917(.din(n980),.dout(n981),.clk(gclk));
	jand g0918(.dina(w_n913_0[0]),.dinb(w_n879_0[0]),.dout(n982),.clk(gclk));
	jand g0919(.dina(w_n914_0[0]),.dinb(w_n876_0[0]),.dout(n983),.clk(gclk));
	jcb g0920(.dina(n983),.dinb(w_dff_B_n6F9CT944_1),.dout(n984));
	jand g0921(.dina(w_G375gat_4[0]),.dinb(w_G171gat_5[1]),.dout(n985),.clk(gclk));
	jnot g0922(.din(n985),.dout(n986),.clk(gclk));
	jand g0923(.dina(w_n911_0[0]),.dinb(w_n884_0[0]),.dout(n987),.clk(gclk));
	jand g0924(.dina(w_n912_0[0]),.dinb(w_n881_0[0]),.dout(n988),.clk(gclk));
	jcb g0925(.dina(n988),.dinb(w_dff_B_T8q6GaV73_1),.dout(n989));
	jand g0926(.dina(w_G358gat_3[2]),.dinb(w_G188gat_5[2]),.dout(n990),.clk(gclk));
	jnot g0927(.din(n990),.dout(n991),.clk(gclk));
	jand g0928(.dina(w_n909_0[0]),.dinb(w_n889_0[0]),.dout(n992),.clk(gclk));
	jand g0929(.dina(w_n910_0[0]),.dinb(w_n886_0[0]),.dout(n993),.clk(gclk));
	jcb g0930(.dina(n993),.dinb(w_dff_B_0FF0RhK38_1),.dout(n994));
	jand g0931(.dina(w_G341gat_3[1]),.dinb(w_G205gat_6[0]),.dout(n995),.clk(gclk));
	jnot g0932(.din(n995),.dout(n996),.clk(gclk));
	jand g0933(.dina(w_n907_0[0]),.dinb(w_n895_0[0]),.dout(n997),.clk(gclk));
	jand g0934(.dina(w_n908_0[0]),.dinb(w_n891_0[0]),.dout(n998),.clk(gclk));
	jcb g0935(.dina(n998),.dinb(w_dff_B_VArijCD09_1),.dout(n999));
	jand g0936(.dina(w_G324gat_3[0]),.dinb(w_G222gat_6[1]),.dout(n1000),.clk(gclk));
	jnot g0937(.din(n1000),.dout(n1001),.clk(gclk));
	jnot g0938(.din(w_n896_0[0]),.dout(n1002),.clk(gclk));
	jnot g0939(.din(w_n906_0[0]),.dout(n1003),.clk(gclk));
	jand g0940(.dina(n1003),.dinb(w_dff_B_NWt7fI1i0_1),.dout(n1004),.clk(gclk));
	jcb g0941(.dina(n1004),.dinb(w_n903_0[0]),.dout(n1005));
	jand g0942(.dina(w_G307gat_3[0]),.dinb(w_G239gat_6[2]),.dout(n1006),.clk(gclk));
	jand g0943(.dina(w_G290gat_2[1]),.dinb(w_G256gat_7[0]),.dout(n1007),.clk(gclk));
	jnot g0944(.din(n1007),.dout(n1008),.clk(gclk));
	jcb g0945(.dina(w_n1008_0[1]),.dinb(w_n793_0[0]),.dout(n1009));
	jxor g0946(.dina(w_n1009_0[1]),.dinb(w_n1006_0[1]),.dout(n1010),.clk(gclk));
	jxor g0947(.dina(w_n1010_0[1]),.dinb(w_n1005_0[1]),.dout(n1011),.clk(gclk));
	jxor g0948(.dina(w_n1011_0[1]),.dinb(w_n1001_0[1]),.dout(n1012),.clk(gclk));
	jxor g0949(.dina(w_n1012_0[1]),.dinb(w_n999_0[1]),.dout(n1013),.clk(gclk));
	jxor g0950(.dina(w_n1013_0[1]),.dinb(w_n996_0[1]),.dout(n1014),.clk(gclk));
	jxor g0951(.dina(w_n1014_0[1]),.dinb(w_n994_0[1]),.dout(n1015),.clk(gclk));
	jxor g0952(.dina(w_n1015_0[1]),.dinb(w_n991_0[1]),.dout(n1016),.clk(gclk));
	jxor g0953(.dina(w_n1016_0[1]),.dinb(w_n989_0[1]),.dout(n1017),.clk(gclk));
	jxor g0954(.dina(w_n1017_0[1]),.dinb(w_n986_0[1]),.dout(n1018),.clk(gclk));
	jxor g0955(.dina(w_n1018_0[1]),.dinb(w_n984_0[1]),.dout(n1019),.clk(gclk));
	jxor g0956(.dina(w_n1019_0[1]),.dinb(w_n981_0[1]),.dout(n1020),.clk(gclk));
	jxor g0957(.dina(w_n1020_0[1]),.dinb(w_n979_0[1]),.dout(n1021),.clk(gclk));
	jxor g0958(.dina(w_n1021_0[1]),.dinb(w_n976_0[1]),.dout(n1022),.clk(gclk));
	jxor g0959(.dina(w_n1022_0[1]),.dinb(w_n974_0[1]),.dout(n1023),.clk(gclk));
	jxor g0960(.dina(w_n1023_0[1]),.dinb(w_n971_0[1]),.dout(n1024),.clk(gclk));
	jxor g0961(.dina(w_n1024_0[1]),.dinb(w_n969_0[1]),.dout(n1025),.clk(gclk));
	jxor g0962(.dina(w_n1025_0[1]),.dinb(w_n966_0[1]),.dout(n1026),.clk(gclk));
	jxor g0963(.dina(w_n1026_0[1]),.dinb(w_n964_0[1]),.dout(n1027),.clk(gclk));
	jxor g0964(.dina(w_n1027_0[1]),.dinb(w_n961_0[1]),.dout(n1028),.clk(gclk));
	jxor g0965(.dina(w_n1028_0[1]),.dinb(w_n959_0[1]),.dout(n1029),.clk(gclk));
	jxor g0966(.dina(w_n1029_0[1]),.dinb(w_n956_0[1]),.dout(n1030),.clk(gclk));
	jxor g0967(.dina(w_n1030_0[1]),.dinb(w_n954_0[1]),.dout(n1031),.clk(gclk));
	jxor g0968(.dina(w_n1031_0[1]),.dinb(w_n951_0[1]),.dout(n1032),.clk(gclk));
	jxor g0969(.dina(w_n1032_0[1]),.dinb(w_n949_0[1]),.dout(n1033),.clk(gclk));
	jxor g0970(.dina(w_n1033_0[1]),.dinb(w_n943_0[1]),.dout(n1034),.clk(gclk));
	jnot g0971(.din(w_n1034_0[1]),.dout(n1035),.clk(gclk));
	jxor g0972(.dina(w_n1035_0[1]),.dinb(w_n942_0[2]),.dout(n1036),.clk(gclk));
	jxor g0973(.dina(n1036),.dinb(w_n938_0[1]),.dout(n1037),.clk(gclk));
	jxor g0974(.dina(w_n1037_0[1]),.dinb(w_n937_0[1]),.dout(G6150gat),.clk(gclk));
	jand g0975(.dina(w_n1037_0[0]),.dinb(w_n937_0[0]),.dout(n1039),.clk(gclk));
	jcb g0976(.dina(w_n1035_0[0]),.dinb(w_n942_0[1]),.dout(n1040));
	jxor g0977(.dina(w_n1034_0[0]),.dinb(w_n942_0[0]),.dout(n1041),.clk(gclk));
	jcb g0978(.dina(n1041),.dinb(w_n938_0[0]),.dout(n1042));
	jand g0979(.dina(n1042),.dinb(n1040),.dout(n1043),.clk(gclk));
	jand g0980(.dina(w_G528gat_6[2]),.dinb(w_G35gat_2[1]),.dout(n1044),.clk(gclk));
	jnot g0981(.din(w_n1032_0[0]),.dout(n1045),.clk(gclk));
	jcb g0982(.dina(n1045),.dinb(w_n949_0[0]),.dout(n1046));
	jcb g0983(.dina(w_n1033_0[0]),.dinb(w_n943_0[0]),.dout(n1047));
	jand g0984(.dina(n1047),.dinb(w_dff_B_zEAdWz9j7_1),.dout(n1048),.clk(gclk));
	jand g0985(.dina(w_G511gat_6[1]),.dinb(w_G52gat_2[2]),.dout(n1049),.clk(gclk));
	jand g0986(.dina(w_n1030_0[0]),.dinb(w_n954_0[0]),.dout(n1050),.clk(gclk));
	jand g0987(.dina(w_n1031_0[0]),.dinb(w_n951_0[0]),.dout(n1051),.clk(gclk));
	jcb g0988(.dina(n1051),.dinb(w_dff_B_yOVGUYnu7_1),.dout(n1052));
	jand g0989(.dina(w_G494gat_6[0]),.dinb(w_G69gat_3[0]),.dout(n1053),.clk(gclk));
	jnot g0990(.din(n1053),.dout(n1054),.clk(gclk));
	jand g0991(.dina(w_n1028_0[0]),.dinb(w_n959_0[0]),.dout(n1055),.clk(gclk));
	jand g0992(.dina(w_n1029_0[0]),.dinb(w_n956_0[0]),.dout(n1056),.clk(gclk));
	jcb g0993(.dina(n1056),.dinb(w_dff_B_Bm80gPTd6_1),.dout(n1057));
	jand g0994(.dina(w_G477gat_5[2]),.dinb(w_G86gat_3[1]),.dout(n1058),.clk(gclk));
	jnot g0995(.din(n1058),.dout(n1059),.clk(gclk));
	jand g0996(.dina(w_n1026_0[0]),.dinb(w_n964_0[0]),.dout(n1060),.clk(gclk));
	jand g0997(.dina(w_n1027_0[0]),.dinb(w_n961_0[0]),.dout(n1061),.clk(gclk));
	jcb g0998(.dina(n1061),.dinb(w_dff_B_V46Xsi6b9_1),.dout(n1062));
	jand g0999(.dina(w_G460gat_5[1]),.dinb(w_G103gat_3[2]),.dout(n1063),.clk(gclk));
	jnot g1000(.din(n1063),.dout(n1064),.clk(gclk));
	jand g1001(.dina(w_n1024_0[0]),.dinb(w_n969_0[0]),.dout(n1065),.clk(gclk));
	jand g1002(.dina(w_n1025_0[0]),.dinb(w_n966_0[0]),.dout(n1066),.clk(gclk));
	jcb g1003(.dina(n1066),.dinb(w_dff_B_Usg5uhqf5_1),.dout(n1067));
	jand g1004(.dina(w_G443gat_5[0]),.dinb(w_G120gat_4[0]),.dout(n1068),.clk(gclk));
	jnot g1005(.din(n1068),.dout(n1069),.clk(gclk));
	jand g1006(.dina(w_n1022_0[0]),.dinb(w_n974_0[0]),.dout(n1070),.clk(gclk));
	jand g1007(.dina(w_n1023_0[0]),.dinb(w_n971_0[0]),.dout(n1071),.clk(gclk));
	jcb g1008(.dina(n1071),.dinb(w_dff_B_LFD6220C1_1),.dout(n1072));
	jand g1009(.dina(w_G426gat_4[2]),.dinb(w_G137gat_4[1]),.dout(n1073),.clk(gclk));
	jnot g1010(.din(n1073),.dout(n1074),.clk(gclk));
	jand g1011(.dina(w_n1020_0[0]),.dinb(w_n979_0[0]),.dout(n1075),.clk(gclk));
	jand g1012(.dina(w_n1021_0[0]),.dinb(w_n976_0[0]),.dout(n1076),.clk(gclk));
	jcb g1013(.dina(n1076),.dinb(w_dff_B_4RoCyyc49_1),.dout(n1077));
	jand g1014(.dina(w_G409gat_4[1]),.dinb(w_G154gat_4[2]),.dout(n1078),.clk(gclk));
	jnot g1015(.din(n1078),.dout(n1079),.clk(gclk));
	jand g1016(.dina(w_n1018_0[0]),.dinb(w_n984_0[0]),.dout(n1080),.clk(gclk));
	jand g1017(.dina(w_n1019_0[0]),.dinb(w_n981_0[0]),.dout(n1081),.clk(gclk));
	jcb g1018(.dina(n1081),.dinb(w_dff_B_HCm4HMBu5_1),.dout(n1082));
	jand g1019(.dina(w_G392gat_4[0]),.dinb(w_G171gat_5[0]),.dout(n1083),.clk(gclk));
	jnot g1020(.din(n1083),.dout(n1084),.clk(gclk));
	jand g1021(.dina(w_n1016_0[0]),.dinb(w_n989_0[0]),.dout(n1085),.clk(gclk));
	jand g1022(.dina(w_n1017_0[0]),.dinb(w_n986_0[0]),.dout(n1086),.clk(gclk));
	jcb g1023(.dina(n1086),.dinb(w_dff_B_14tFs7Lf3_1),.dout(n1087));
	jand g1024(.dina(w_G375gat_3[2]),.dinb(w_G188gat_5[1]),.dout(n1088),.clk(gclk));
	jnot g1025(.din(n1088),.dout(n1089),.clk(gclk));
	jand g1026(.dina(w_n1014_0[0]),.dinb(w_n994_0[0]),.dout(n1090),.clk(gclk));
	jand g1027(.dina(w_n1015_0[0]),.dinb(w_n991_0[0]),.dout(n1091),.clk(gclk));
	jcb g1028(.dina(n1091),.dinb(w_dff_B_YI5hYO794_1),.dout(n1092));
	jand g1029(.dina(w_G358gat_3[1]),.dinb(w_G205gat_5[2]),.dout(n1093),.clk(gclk));
	jnot g1030(.din(n1093),.dout(n1094),.clk(gclk));
	jand g1031(.dina(w_n1012_0[0]),.dinb(w_n999_0[0]),.dout(n1095),.clk(gclk));
	jand g1032(.dina(w_n1013_0[0]),.dinb(w_n996_0[0]),.dout(n1096),.clk(gclk));
	jcb g1033(.dina(n1096),.dinb(w_dff_B_CaNGttoo6_1),.dout(n1097));
	jand g1034(.dina(w_G341gat_3[0]),.dinb(w_G222gat_6[0]),.dout(n1098),.clk(gclk));
	jnot g1035(.din(n1098),.dout(n1099),.clk(gclk));
	jand g1036(.dina(w_n1010_0[0]),.dinb(w_n1005_0[0]),.dout(n1100),.clk(gclk));
	jand g1037(.dina(w_n1011_0[0]),.dinb(w_n1001_0[0]),.dout(n1101),.clk(gclk));
	jcb g1038(.dina(n1101),.dinb(w_dff_B_04222BGw5_1),.dout(n1102));
	jand g1039(.dina(w_G324gat_2[2]),.dinb(w_G239gat_6[1]),.dout(n1103),.clk(gclk));
	jand g1040(.dina(w_G307gat_2[2]),.dinb(w_G256gat_6[2]),.dout(n1104),.clk(gclk));
	jnot g1041(.din(w_n1006_0[0]),.dout(n1105),.clk(gclk));
	jnot g1042(.din(w_n1009_0[0]),.dout(n1106),.clk(gclk));
	jand g1043(.dina(n1106),.dinb(w_dff_B_eo89BVpV8_1),.dout(n1107),.clk(gclk));
	jcb g1044(.dina(n1107),.dinb(w_n1008_0[0]),.dout(n1108));
	jnot g1045(.din(n1108),.dout(n1109),.clk(gclk));
	jcb g1046(.dina(w_n1109_0[1]),.dinb(w_dff_B_bUMTWNEB1_1),.dout(n1110));
	jand g1047(.dina(w_n1109_0[0]),.dinb(w_G307gat_2[1]),.dout(n1111),.clk(gclk));
	jnot g1048(.din(n1111),.dout(n1112),.clk(gclk));
	jand g1049(.dina(n1112),.dinb(w_n1110_0[1]),.dout(n1113),.clk(gclk));
	jnot g1050(.din(n1113),.dout(n1114),.clk(gclk));
	jxor g1051(.dina(w_n1114_0[1]),.dinb(w_n1103_0[1]),.dout(n1115),.clk(gclk));
	jxor g1052(.dina(w_n1115_0[1]),.dinb(w_n1102_0[1]),.dout(n1116),.clk(gclk));
	jxor g1053(.dina(w_n1116_0[1]),.dinb(w_n1099_0[1]),.dout(n1117),.clk(gclk));
	jxor g1054(.dina(w_n1117_0[1]),.dinb(w_n1097_0[1]),.dout(n1118),.clk(gclk));
	jxor g1055(.dina(w_n1118_0[1]),.dinb(w_n1094_0[1]),.dout(n1119),.clk(gclk));
	jxor g1056(.dina(w_n1119_0[1]),.dinb(w_n1092_0[1]),.dout(n1120),.clk(gclk));
	jxor g1057(.dina(w_n1120_0[1]),.dinb(w_n1089_0[1]),.dout(n1121),.clk(gclk));
	jxor g1058(.dina(w_n1121_0[1]),.dinb(w_n1087_0[1]),.dout(n1122),.clk(gclk));
	jxor g1059(.dina(w_n1122_0[1]),.dinb(w_n1084_0[1]),.dout(n1123),.clk(gclk));
	jxor g1060(.dina(w_n1123_0[1]),.dinb(w_n1082_0[1]),.dout(n1124),.clk(gclk));
	jxor g1061(.dina(w_n1124_0[1]),.dinb(w_n1079_0[1]),.dout(n1125),.clk(gclk));
	jxor g1062(.dina(w_n1125_0[1]),.dinb(w_n1077_0[1]),.dout(n1126),.clk(gclk));
	jxor g1063(.dina(w_n1126_0[1]),.dinb(w_n1074_0[1]),.dout(n1127),.clk(gclk));
	jxor g1064(.dina(w_n1127_0[1]),.dinb(w_n1072_0[1]),.dout(n1128),.clk(gclk));
	jxor g1065(.dina(w_n1128_0[1]),.dinb(w_n1069_0[1]),.dout(n1129),.clk(gclk));
	jxor g1066(.dina(w_n1129_0[1]),.dinb(w_n1067_0[1]),.dout(n1130),.clk(gclk));
	jxor g1067(.dina(w_n1130_0[1]),.dinb(w_n1064_0[1]),.dout(n1131),.clk(gclk));
	jxor g1068(.dina(w_n1131_0[1]),.dinb(w_n1062_0[1]),.dout(n1132),.clk(gclk));
	jxor g1069(.dina(w_n1132_0[1]),.dinb(w_n1059_0[1]),.dout(n1133),.clk(gclk));
	jxor g1070(.dina(w_n1133_0[1]),.dinb(w_n1057_0[1]),.dout(n1134),.clk(gclk));
	jxor g1071(.dina(w_n1134_0[1]),.dinb(w_n1054_0[1]),.dout(n1135),.clk(gclk));
	jxor g1072(.dina(w_n1135_0[1]),.dinb(w_n1052_0[1]),.dout(n1136),.clk(gclk));
	jnot g1073(.din(n1136),.dout(n1137),.clk(gclk));
	jxor g1074(.dina(w_n1137_0[1]),.dinb(w_n1049_0[1]),.dout(n1138),.clk(gclk));
	jxor g1075(.dina(w_n1138_0[1]),.dinb(w_n1048_0[1]),.dout(n1139),.clk(gclk));
	jxor g1076(.dina(w_n1139_0[1]),.dinb(w_n1044_0[1]),.dout(n1140),.clk(gclk));
	jxor g1077(.dina(w_n1140_0[1]),.dinb(w_n1043_0[1]),.dout(n1141),.clk(gclk));
	jnot g1078(.din(w_n1141_0[1]),.dout(n1142),.clk(gclk));
	jxor g1079(.dina(n1142),.dinb(w_n1039_0[1]),.dout(G6160gat),.clk(gclk));
	jnot g1080(.din(w_n1140_0[0]),.dout(n1144),.clk(gclk));
	jcb g1081(.dina(n1144),.dinb(w_n1043_0[0]),.dout(n1145));
	jcb g1082(.dina(w_n1141_0[0]),.dinb(w_n1039_0[0]),.dout(n1146));
	jand g1083(.dina(n1146),.dinb(n1145),.dout(n1147),.clk(gclk));
	jnot g1084(.din(w_n1138_0[0]),.dout(n1148),.clk(gclk));
	jcb g1085(.dina(n1148),.dinb(w_n1048_0[0]),.dout(n1149));
	jcb g1086(.dina(w_n1139_0[0]),.dinb(w_n1044_0[0]),.dout(n1150));
	jand g1087(.dina(n1150),.dinb(n1149),.dout(n1151),.clk(gclk));
	jand g1088(.dina(w_G528gat_6[1]),.dinb(w_G52gat_2[1]),.dout(n1152),.clk(gclk));
	jand g1089(.dina(w_n1135_0[0]),.dinb(w_n1052_0[0]),.dout(n1153),.clk(gclk));
	jnot g1090(.din(n1153),.dout(n1154),.clk(gclk));
	jcb g1091(.dina(w_n1137_0[0]),.dinb(w_n1049_0[0]),.dout(n1155));
	jand g1092(.dina(n1155),.dinb(n1154),.dout(n1156),.clk(gclk));
	jand g1093(.dina(w_G511gat_6[0]),.dinb(w_G69gat_2[2]),.dout(n1157),.clk(gclk));
	jnot g1094(.din(n1157),.dout(n1158),.clk(gclk));
	jand g1095(.dina(w_n1133_0[0]),.dinb(w_n1057_0[0]),.dout(n1159),.clk(gclk));
	jand g1096(.dina(w_n1134_0[0]),.dinb(w_n1054_0[0]),.dout(n1160),.clk(gclk));
	jcb g1097(.dina(n1160),.dinb(w_dff_B_isMwcS1w1_1),.dout(n1161));
	jand g1098(.dina(w_G494gat_5[2]),.dinb(w_G86gat_3[0]),.dout(n1162),.clk(gclk));
	jnot g1099(.din(n1162),.dout(n1163),.clk(gclk));
	jand g1100(.dina(w_n1131_0[0]),.dinb(w_n1062_0[0]),.dout(n1164),.clk(gclk));
	jand g1101(.dina(w_n1132_0[0]),.dinb(w_n1059_0[0]),.dout(n1165),.clk(gclk));
	jcb g1102(.dina(n1165),.dinb(w_dff_B_YVApPPrf4_1),.dout(n1166));
	jand g1103(.dina(w_G477gat_5[1]),.dinb(w_G103gat_3[1]),.dout(n1167),.clk(gclk));
	jnot g1104(.din(n1167),.dout(n1168),.clk(gclk));
	jand g1105(.dina(w_n1129_0[0]),.dinb(w_n1067_0[0]),.dout(n1169),.clk(gclk));
	jand g1106(.dina(w_n1130_0[0]),.dinb(w_n1064_0[0]),.dout(n1170),.clk(gclk));
	jcb g1107(.dina(n1170),.dinb(w_dff_B_ELpE24bH9_1),.dout(n1171));
	jand g1108(.dina(w_G460gat_5[0]),.dinb(w_G120gat_3[2]),.dout(n1172),.clk(gclk));
	jnot g1109(.din(n1172),.dout(n1173),.clk(gclk));
	jand g1110(.dina(w_n1127_0[0]),.dinb(w_n1072_0[0]),.dout(n1174),.clk(gclk));
	jand g1111(.dina(w_n1128_0[0]),.dinb(w_n1069_0[0]),.dout(n1175),.clk(gclk));
	jcb g1112(.dina(n1175),.dinb(w_dff_B_m3XPCPsF9_1),.dout(n1176));
	jand g1113(.dina(w_G443gat_4[2]),.dinb(w_G137gat_4[0]),.dout(n1177),.clk(gclk));
	jnot g1114(.din(n1177),.dout(n1178),.clk(gclk));
	jand g1115(.dina(w_n1125_0[0]),.dinb(w_n1077_0[0]),.dout(n1179),.clk(gclk));
	jand g1116(.dina(w_n1126_0[0]),.dinb(w_n1074_0[0]),.dout(n1180),.clk(gclk));
	jcb g1117(.dina(n1180),.dinb(w_dff_B_J41R32b15_1),.dout(n1181));
	jand g1118(.dina(w_G426gat_4[1]),.dinb(w_G154gat_4[1]),.dout(n1182),.clk(gclk));
	jnot g1119(.din(n1182),.dout(n1183),.clk(gclk));
	jand g1120(.dina(w_n1123_0[0]),.dinb(w_n1082_0[0]),.dout(n1184),.clk(gclk));
	jand g1121(.dina(w_n1124_0[0]),.dinb(w_n1079_0[0]),.dout(n1185),.clk(gclk));
	jcb g1122(.dina(n1185),.dinb(w_dff_B_9Uieaijd3_1),.dout(n1186));
	jand g1123(.dina(w_G409gat_4[0]),.dinb(w_G171gat_4[2]),.dout(n1187),.clk(gclk));
	jnot g1124(.din(n1187),.dout(n1188),.clk(gclk));
	jand g1125(.dina(w_n1121_0[0]),.dinb(w_n1087_0[0]),.dout(n1189),.clk(gclk));
	jand g1126(.dina(w_n1122_0[0]),.dinb(w_n1084_0[0]),.dout(n1190),.clk(gclk));
	jcb g1127(.dina(n1190),.dinb(w_dff_B_dFsHh26v2_1),.dout(n1191));
	jand g1128(.dina(w_G392gat_3[2]),.dinb(w_G188gat_5[0]),.dout(n1192),.clk(gclk));
	jnot g1129(.din(n1192),.dout(n1193),.clk(gclk));
	jand g1130(.dina(w_n1119_0[0]),.dinb(w_n1092_0[0]),.dout(n1194),.clk(gclk));
	jand g1131(.dina(w_n1120_0[0]),.dinb(w_n1089_0[0]),.dout(n1195),.clk(gclk));
	jcb g1132(.dina(n1195),.dinb(w_dff_B_KMgHgW2O2_1),.dout(n1196));
	jand g1133(.dina(w_G375gat_3[1]),.dinb(w_G205gat_5[1]),.dout(n1197),.clk(gclk));
	jnot g1134(.din(n1197),.dout(n1198),.clk(gclk));
	jand g1135(.dina(w_n1117_0[0]),.dinb(w_n1097_0[0]),.dout(n1199),.clk(gclk));
	jand g1136(.dina(w_n1118_0[0]),.dinb(w_n1094_0[0]),.dout(n1200),.clk(gclk));
	jcb g1137(.dina(n1200),.dinb(w_dff_B_ztUuxrZa4_1),.dout(n1201));
	jand g1138(.dina(w_G358gat_3[0]),.dinb(w_G222gat_5[2]),.dout(n1202),.clk(gclk));
	jnot g1139(.din(n1202),.dout(n1203),.clk(gclk));
	jand g1140(.dina(w_n1115_0[0]),.dinb(w_n1102_0[0]),.dout(n1204),.clk(gclk));
	jand g1141(.dina(w_n1116_0[0]),.dinb(w_n1099_0[0]),.dout(n1205),.clk(gclk));
	jcb g1142(.dina(n1205),.dinb(w_dff_B_1JPldOdX0_1),.dout(n1206));
	jand g1143(.dina(w_G341gat_2[2]),.dinb(w_G239gat_6[0]),.dout(n1207),.clk(gclk));
	jand g1144(.dina(w_G324gat_2[1]),.dinb(w_G256gat_6[1]),.dout(n1208),.clk(gclk));
	jcb g1145(.dina(w_n1114_0[0]),.dinb(w_n1103_0[0]),.dout(n1209));
	jand g1146(.dina(n1209),.dinb(w_n1110_0[0]),.dout(n1210),.clk(gclk));
	jxor g1147(.dina(w_n1210_0[1]),.dinb(w_n1208_0[1]),.dout(n1211),.clk(gclk));
	jnot g1148(.din(n1211),.dout(n1212),.clk(gclk));
	jxor g1149(.dina(w_n1212_0[1]),.dinb(w_n1207_0[1]),.dout(n1213),.clk(gclk));
	jxor g1150(.dina(w_n1213_0[1]),.dinb(w_n1206_0[1]),.dout(n1214),.clk(gclk));
	jxor g1151(.dina(w_n1214_0[1]),.dinb(w_n1203_0[1]),.dout(n1215),.clk(gclk));
	jxor g1152(.dina(w_n1215_0[1]),.dinb(w_n1201_0[1]),.dout(n1216),.clk(gclk));
	jxor g1153(.dina(w_n1216_0[1]),.dinb(w_n1198_0[1]),.dout(n1217),.clk(gclk));
	jxor g1154(.dina(w_n1217_0[1]),.dinb(w_n1196_0[1]),.dout(n1218),.clk(gclk));
	jxor g1155(.dina(w_n1218_0[1]),.dinb(w_n1193_0[1]),.dout(n1219),.clk(gclk));
	jxor g1156(.dina(w_n1219_0[1]),.dinb(w_n1191_0[1]),.dout(n1220),.clk(gclk));
	jxor g1157(.dina(w_n1220_0[1]),.dinb(w_n1188_0[1]),.dout(n1221),.clk(gclk));
	jxor g1158(.dina(w_n1221_0[1]),.dinb(w_n1186_0[1]),.dout(n1222),.clk(gclk));
	jxor g1159(.dina(w_n1222_0[1]),.dinb(w_n1183_0[1]),.dout(n1223),.clk(gclk));
	jxor g1160(.dina(w_n1223_0[1]),.dinb(w_n1181_0[1]),.dout(n1224),.clk(gclk));
	jxor g1161(.dina(w_n1224_0[1]),.dinb(w_n1178_0[1]),.dout(n1225),.clk(gclk));
	jxor g1162(.dina(w_n1225_0[1]),.dinb(w_n1176_0[1]),.dout(n1226),.clk(gclk));
	jxor g1163(.dina(w_n1226_0[1]),.dinb(w_n1173_0[1]),.dout(n1227),.clk(gclk));
	jxor g1164(.dina(w_n1227_0[1]),.dinb(w_n1171_0[1]),.dout(n1228),.clk(gclk));
	jxor g1165(.dina(w_n1228_0[1]),.dinb(w_n1168_0[1]),.dout(n1229),.clk(gclk));
	jxor g1166(.dina(w_n1229_0[1]),.dinb(w_n1166_0[1]),.dout(n1230),.clk(gclk));
	jxor g1167(.dina(w_n1230_0[1]),.dinb(w_n1163_0[1]),.dout(n1231),.clk(gclk));
	jxor g1168(.dina(w_n1231_0[1]),.dinb(w_n1161_0[1]),.dout(n1232),.clk(gclk));
	jxor g1169(.dina(w_n1232_0[1]),.dinb(w_n1158_0[1]),.dout(n1233),.clk(gclk));
	jnot g1170(.din(n1233),.dout(n1234),.clk(gclk));
	jxor g1171(.dina(w_n1234_0[1]),.dinb(w_n1156_0[1]),.dout(n1235),.clk(gclk));
	jnot g1172(.din(n1235),.dout(n1236),.clk(gclk));
	jxor g1173(.dina(w_n1236_0[1]),.dinb(w_n1152_0[1]),.dout(n1237),.clk(gclk));
	jxor g1174(.dina(w_n1237_0[1]),.dinb(w_n1151_0[1]),.dout(n1238),.clk(gclk));
	jnot g1175(.din(w_n1238_0[1]),.dout(n1239),.clk(gclk));
	jxor g1176(.dina(n1239),.dinb(w_n1147_0[1]),.dout(G6170gat),.clk(gclk));
	jnot g1177(.din(w_n1237_0[0]),.dout(n1241),.clk(gclk));
	jcb g1178(.dina(n1241),.dinb(w_n1151_0[0]),.dout(n1242));
	jcb g1179(.dina(w_n1238_0[0]),.dinb(w_n1147_0[0]),.dout(n1243));
	jand g1180(.dina(n1243),.dinb(n1242),.dout(n1244),.clk(gclk));
	jcb g1181(.dina(w_n1234_0[0]),.dinb(w_n1156_0[0]),.dout(n1245));
	jcb g1182(.dina(w_n1236_0[0]),.dinb(w_n1152_0[0]),.dout(n1246));
	jand g1183(.dina(n1246),.dinb(w_dff_B_HQ0398zs6_1),.dout(n1247),.clk(gclk));
	jand g1184(.dina(w_G528gat_6[0]),.dinb(w_G69gat_2[1]),.dout(n1248),.clk(gclk));
	jand g1185(.dina(w_n1231_0[0]),.dinb(w_n1161_0[0]),.dout(n1249),.clk(gclk));
	jand g1186(.dina(w_n1232_0[0]),.dinb(w_n1158_0[0]),.dout(n1250),.clk(gclk));
	jcb g1187(.dina(n1250),.dinb(w_dff_B_tV69P8c58_1),.dout(n1251));
	jand g1188(.dina(w_G511gat_5[2]),.dinb(w_G86gat_2[2]),.dout(n1252),.clk(gclk));
	jnot g1189(.din(n1252),.dout(n1253),.clk(gclk));
	jand g1190(.dina(w_n1229_0[0]),.dinb(w_n1166_0[0]),.dout(n1254),.clk(gclk));
	jand g1191(.dina(w_n1230_0[0]),.dinb(w_n1163_0[0]),.dout(n1255),.clk(gclk));
	jcb g1192(.dina(n1255),.dinb(w_dff_B_Jm9tIshv4_1),.dout(n1256));
	jand g1193(.dina(w_G494gat_5[1]),.dinb(w_G103gat_3[0]),.dout(n1257),.clk(gclk));
	jnot g1194(.din(n1257),.dout(n1258),.clk(gclk));
	jand g1195(.dina(w_n1227_0[0]),.dinb(w_n1171_0[0]),.dout(n1259),.clk(gclk));
	jand g1196(.dina(w_n1228_0[0]),.dinb(w_n1168_0[0]),.dout(n1260),.clk(gclk));
	jcb g1197(.dina(n1260),.dinb(w_dff_B_cvqoWs9e8_1),.dout(n1261));
	jand g1198(.dina(w_G477gat_5[0]),.dinb(w_G120gat_3[1]),.dout(n1262),.clk(gclk));
	jnot g1199(.din(n1262),.dout(n1263),.clk(gclk));
	jand g1200(.dina(w_n1225_0[0]),.dinb(w_n1176_0[0]),.dout(n1264),.clk(gclk));
	jand g1201(.dina(w_n1226_0[0]),.dinb(w_n1173_0[0]),.dout(n1265),.clk(gclk));
	jcb g1202(.dina(n1265),.dinb(w_dff_B_ppPcRfFc9_1),.dout(n1266));
	jand g1203(.dina(w_G460gat_4[2]),.dinb(w_G137gat_3[2]),.dout(n1267),.clk(gclk));
	jnot g1204(.din(n1267),.dout(n1268),.clk(gclk));
	jand g1205(.dina(w_n1223_0[0]),.dinb(w_n1181_0[0]),.dout(n1269),.clk(gclk));
	jand g1206(.dina(w_n1224_0[0]),.dinb(w_n1178_0[0]),.dout(n1270),.clk(gclk));
	jcb g1207(.dina(n1270),.dinb(w_dff_B_nhgki9g39_1),.dout(n1271));
	jand g1208(.dina(w_G443gat_4[1]),.dinb(w_G154gat_4[0]),.dout(n1272),.clk(gclk));
	jnot g1209(.din(n1272),.dout(n1273),.clk(gclk));
	jand g1210(.dina(w_n1221_0[0]),.dinb(w_n1186_0[0]),.dout(n1274),.clk(gclk));
	jand g1211(.dina(w_n1222_0[0]),.dinb(w_n1183_0[0]),.dout(n1275),.clk(gclk));
	jcb g1212(.dina(n1275),.dinb(w_dff_B_mq9duBnh9_1),.dout(n1276));
	jand g1213(.dina(w_G426gat_4[0]),.dinb(w_G171gat_4[1]),.dout(n1277),.clk(gclk));
	jnot g1214(.din(n1277),.dout(n1278),.clk(gclk));
	jand g1215(.dina(w_n1219_0[0]),.dinb(w_n1191_0[0]),.dout(n1279),.clk(gclk));
	jand g1216(.dina(w_n1220_0[0]),.dinb(w_n1188_0[0]),.dout(n1280),.clk(gclk));
	jcb g1217(.dina(n1280),.dinb(w_dff_B_fGZzhjhB6_1),.dout(n1281));
	jand g1218(.dina(w_G409gat_3[2]),.dinb(w_G188gat_4[2]),.dout(n1282),.clk(gclk));
	jnot g1219(.din(n1282),.dout(n1283),.clk(gclk));
	jand g1220(.dina(w_n1217_0[0]),.dinb(w_n1196_0[0]),.dout(n1284),.clk(gclk));
	jand g1221(.dina(w_n1218_0[0]),.dinb(w_n1193_0[0]),.dout(n1285),.clk(gclk));
	jcb g1222(.dina(n1285),.dinb(w_dff_B_r7ZG6dqT3_1),.dout(n1286));
	jand g1223(.dina(w_G392gat_3[1]),.dinb(w_G205gat_5[0]),.dout(n1287),.clk(gclk));
	jnot g1224(.din(n1287),.dout(n1288),.clk(gclk));
	jand g1225(.dina(w_n1215_0[0]),.dinb(w_n1201_0[0]),.dout(n1289),.clk(gclk));
	jand g1226(.dina(w_n1216_0[0]),.dinb(w_n1198_0[0]),.dout(n1290),.clk(gclk));
	jcb g1227(.dina(n1290),.dinb(w_dff_B_1n21AahF4_1),.dout(n1291));
	jand g1228(.dina(w_G375gat_3[0]),.dinb(w_G222gat_5[1]),.dout(n1292),.clk(gclk));
	jnot g1229(.din(n1292),.dout(n1293),.clk(gclk));
	jand g1230(.dina(w_n1213_0[0]),.dinb(w_n1206_0[0]),.dout(n1294),.clk(gclk));
	jand g1231(.dina(w_n1214_0[0]),.dinb(w_n1203_0[0]),.dout(n1295),.clk(gclk));
	jcb g1232(.dina(n1295),.dinb(w_dff_B_6OoSuzZF7_1),.dout(n1296));
	jand g1233(.dina(w_G358gat_2[2]),.dinb(w_G239gat_5[2]),.dout(n1297),.clk(gclk));
	jand g1234(.dina(w_G341gat_2[1]),.dinb(w_G256gat_6[0]),.dout(n1298),.clk(gclk));
	jcb g1235(.dina(w_n1210_0[0]),.dinb(w_n1208_0[0]),.dout(n1299));
	jcb g1236(.dina(w_n1212_0[0]),.dinb(w_n1207_0[0]),.dout(n1300));
	jand g1237(.dina(n1300),.dinb(w_dff_B_moMeQzNZ4_1),.dout(n1301),.clk(gclk));
	jxor g1238(.dina(w_n1301_0[1]),.dinb(w_n1298_0[1]),.dout(n1302),.clk(gclk));
	jnot g1239(.din(n1302),.dout(n1303),.clk(gclk));
	jxor g1240(.dina(w_n1303_0[1]),.dinb(w_n1297_0[1]),.dout(n1304),.clk(gclk));
	jxor g1241(.dina(w_n1304_0[1]),.dinb(w_n1296_0[1]),.dout(n1305),.clk(gclk));
	jxor g1242(.dina(w_n1305_0[1]),.dinb(w_n1293_0[1]),.dout(n1306),.clk(gclk));
	jxor g1243(.dina(w_n1306_0[1]),.dinb(w_n1291_0[1]),.dout(n1307),.clk(gclk));
	jxor g1244(.dina(w_n1307_0[1]),.dinb(w_n1288_0[1]),.dout(n1308),.clk(gclk));
	jxor g1245(.dina(w_n1308_0[1]),.dinb(w_n1286_0[1]),.dout(n1309),.clk(gclk));
	jxor g1246(.dina(w_n1309_0[1]),.dinb(w_n1283_0[1]),.dout(n1310),.clk(gclk));
	jxor g1247(.dina(w_n1310_0[1]),.dinb(w_n1281_0[1]),.dout(n1311),.clk(gclk));
	jxor g1248(.dina(w_n1311_0[1]),.dinb(w_n1278_0[1]),.dout(n1312),.clk(gclk));
	jxor g1249(.dina(w_n1312_0[1]),.dinb(w_n1276_0[1]),.dout(n1313),.clk(gclk));
	jxor g1250(.dina(w_n1313_0[1]),.dinb(w_n1273_0[1]),.dout(n1314),.clk(gclk));
	jxor g1251(.dina(w_n1314_0[1]),.dinb(w_n1271_0[1]),.dout(n1315),.clk(gclk));
	jxor g1252(.dina(w_n1315_0[1]),.dinb(w_n1268_0[1]),.dout(n1316),.clk(gclk));
	jxor g1253(.dina(w_n1316_0[1]),.dinb(w_n1266_0[1]),.dout(n1317),.clk(gclk));
	jxor g1254(.dina(w_n1317_0[1]),.dinb(w_n1263_0[1]),.dout(n1318),.clk(gclk));
	jxor g1255(.dina(w_n1318_0[1]),.dinb(w_n1261_0[1]),.dout(n1319),.clk(gclk));
	jxor g1256(.dina(w_n1319_0[1]),.dinb(w_n1258_0[1]),.dout(n1320),.clk(gclk));
	jxor g1257(.dina(w_n1320_0[1]),.dinb(w_n1256_0[1]),.dout(n1321),.clk(gclk));
	jxor g1258(.dina(w_n1321_0[1]),.dinb(w_n1253_0[1]),.dout(n1322),.clk(gclk));
	jxor g1259(.dina(w_n1322_0[1]),.dinb(w_n1251_0[1]),.dout(n1323),.clk(gclk));
	jnot g1260(.din(n1323),.dout(n1324),.clk(gclk));
	jxor g1261(.dina(w_n1324_0[1]),.dinb(w_n1248_0[1]),.dout(n1325),.clk(gclk));
	jxor g1262(.dina(w_n1325_0[1]),.dinb(w_n1247_0[1]),.dout(n1326),.clk(gclk));
	jnot g1263(.din(w_n1326_0[1]),.dout(n1327),.clk(gclk));
	jxor g1264(.dina(n1327),.dinb(w_n1244_0[1]),.dout(G6180gat),.clk(gclk));
	jnot g1265(.din(w_n1325_0[0]),.dout(n1329),.clk(gclk));
	jcb g1266(.dina(n1329),.dinb(w_n1247_0[0]),.dout(n1330));
	jcb g1267(.dina(w_n1326_0[0]),.dinb(w_n1244_0[0]),.dout(n1331));
	jand g1268(.dina(n1331),.dinb(w_dff_B_aUjjF2ug5_1),.dout(n1332),.clk(gclk));
	jnot g1269(.din(w_n1251_0[0]),.dout(n1333),.clk(gclk));
	jnot g1270(.din(w_n1322_0[0]),.dout(n1334),.clk(gclk));
	jcb g1271(.dina(n1334),.dinb(w_dff_B_NAWMwQTb3_1),.dout(n1335));
	jcb g1272(.dina(w_n1324_0[0]),.dinb(w_n1248_0[0]),.dout(n1336));
	jand g1273(.dina(n1336),.dinb(w_dff_B_cEx3tPYS7_1),.dout(n1337),.clk(gclk));
	jand g1274(.dina(w_G528gat_5[2]),.dinb(w_G86gat_2[1]),.dout(n1338),.clk(gclk));
	jand g1275(.dina(w_n1320_0[0]),.dinb(w_n1256_0[0]),.dout(n1339),.clk(gclk));
	jand g1276(.dina(w_n1321_0[0]),.dinb(w_n1253_0[0]),.dout(n1340),.clk(gclk));
	jcb g1277(.dina(n1340),.dinb(w_dff_B_PgiGbC5X8_1),.dout(n1341));
	jand g1278(.dina(w_G511gat_5[1]),.dinb(w_G103gat_2[2]),.dout(n1342),.clk(gclk));
	jnot g1279(.din(n1342),.dout(n1343),.clk(gclk));
	jand g1280(.dina(w_n1318_0[0]),.dinb(w_n1261_0[0]),.dout(n1344),.clk(gclk));
	jand g1281(.dina(w_n1319_0[0]),.dinb(w_n1258_0[0]),.dout(n1345),.clk(gclk));
	jcb g1282(.dina(n1345),.dinb(w_dff_B_ivnOAsjy4_1),.dout(n1346));
	jand g1283(.dina(w_G494gat_5[0]),.dinb(w_G120gat_3[0]),.dout(n1347),.clk(gclk));
	jnot g1284(.din(n1347),.dout(n1348),.clk(gclk));
	jand g1285(.dina(w_n1316_0[0]),.dinb(w_n1266_0[0]),.dout(n1349),.clk(gclk));
	jand g1286(.dina(w_n1317_0[0]),.dinb(w_n1263_0[0]),.dout(n1350),.clk(gclk));
	jcb g1287(.dina(n1350),.dinb(w_dff_B_y4LofFOP8_1),.dout(n1351));
	jand g1288(.dina(w_G477gat_4[2]),.dinb(w_G137gat_3[1]),.dout(n1352),.clk(gclk));
	jnot g1289(.din(n1352),.dout(n1353),.clk(gclk));
	jand g1290(.dina(w_n1314_0[0]),.dinb(w_n1271_0[0]),.dout(n1354),.clk(gclk));
	jand g1291(.dina(w_n1315_0[0]),.dinb(w_n1268_0[0]),.dout(n1355),.clk(gclk));
	jcb g1292(.dina(n1355),.dinb(w_dff_B_gQxEYNeQ5_1),.dout(n1356));
	jand g1293(.dina(w_G460gat_4[1]),.dinb(w_G154gat_3[2]),.dout(n1357),.clk(gclk));
	jnot g1294(.din(n1357),.dout(n1358),.clk(gclk));
	jand g1295(.dina(w_n1312_0[0]),.dinb(w_n1276_0[0]),.dout(n1359),.clk(gclk));
	jand g1296(.dina(w_n1313_0[0]),.dinb(w_n1273_0[0]),.dout(n1360),.clk(gclk));
	jcb g1297(.dina(n1360),.dinb(w_dff_B_xbndg6UF9_1),.dout(n1361));
	jand g1298(.dina(w_G443gat_4[0]),.dinb(w_G171gat_4[0]),.dout(n1362),.clk(gclk));
	jnot g1299(.din(n1362),.dout(n1363),.clk(gclk));
	jand g1300(.dina(w_n1310_0[0]),.dinb(w_n1281_0[0]),.dout(n1364),.clk(gclk));
	jand g1301(.dina(w_n1311_0[0]),.dinb(w_n1278_0[0]),.dout(n1365),.clk(gclk));
	jcb g1302(.dina(n1365),.dinb(w_dff_B_HcTs0byL2_1),.dout(n1366));
	jand g1303(.dina(w_G426gat_3[2]),.dinb(w_G188gat_4[1]),.dout(n1367),.clk(gclk));
	jnot g1304(.din(n1367),.dout(n1368),.clk(gclk));
	jand g1305(.dina(w_n1308_0[0]),.dinb(w_n1286_0[0]),.dout(n1369),.clk(gclk));
	jand g1306(.dina(w_n1309_0[0]),.dinb(w_n1283_0[0]),.dout(n1370),.clk(gclk));
	jcb g1307(.dina(n1370),.dinb(w_dff_B_kdxQH1hD6_1),.dout(n1371));
	jand g1308(.dina(w_G409gat_3[1]),.dinb(w_G205gat_4[2]),.dout(n1372),.clk(gclk));
	jnot g1309(.din(n1372),.dout(n1373),.clk(gclk));
	jand g1310(.dina(w_n1306_0[0]),.dinb(w_n1291_0[0]),.dout(n1374),.clk(gclk));
	jand g1311(.dina(w_n1307_0[0]),.dinb(w_n1288_0[0]),.dout(n1375),.clk(gclk));
	jcb g1312(.dina(n1375),.dinb(w_dff_B_INKymOYR8_1),.dout(n1376));
	jand g1313(.dina(w_G392gat_3[0]),.dinb(w_G222gat_5[0]),.dout(n1377),.clk(gclk));
	jnot g1314(.din(n1377),.dout(n1378),.clk(gclk));
	jand g1315(.dina(w_n1304_0[0]),.dinb(w_n1296_0[0]),.dout(n1379),.clk(gclk));
	jand g1316(.dina(w_n1305_0[0]),.dinb(w_n1293_0[0]),.dout(n1380),.clk(gclk));
	jcb g1317(.dina(n1380),.dinb(w_dff_B_JkXbNzCC9_1),.dout(n1381));
	jand g1318(.dina(w_G375gat_2[2]),.dinb(w_G239gat_5[1]),.dout(n1382),.clk(gclk));
	jand g1319(.dina(w_G358gat_2[1]),.dinb(w_G256gat_5[2]),.dout(n1383),.clk(gclk));
	jcb g1320(.dina(w_n1301_0[0]),.dinb(w_n1298_0[0]),.dout(n1384));
	jcb g1321(.dina(w_n1303_0[0]),.dinb(w_n1297_0[0]),.dout(n1385));
	jand g1322(.dina(n1385),.dinb(w_dff_B_Oa0pA2St3_1),.dout(n1386),.clk(gclk));
	jxor g1323(.dina(w_n1386_0[1]),.dinb(w_n1383_0[1]),.dout(n1387),.clk(gclk));
	jnot g1324(.din(n1387),.dout(n1388),.clk(gclk));
	jxor g1325(.dina(w_n1388_0[1]),.dinb(w_n1382_0[1]),.dout(n1389),.clk(gclk));
	jxor g1326(.dina(w_n1389_0[1]),.dinb(w_n1381_0[1]),.dout(n1390),.clk(gclk));
	jxor g1327(.dina(w_n1390_0[1]),.dinb(w_n1378_0[1]),.dout(n1391),.clk(gclk));
	jxor g1328(.dina(w_n1391_0[1]),.dinb(w_n1376_0[1]),.dout(n1392),.clk(gclk));
	jxor g1329(.dina(w_n1392_0[1]),.dinb(w_n1373_0[1]),.dout(n1393),.clk(gclk));
	jxor g1330(.dina(w_n1393_0[1]),.dinb(w_n1371_0[1]),.dout(n1394),.clk(gclk));
	jxor g1331(.dina(w_n1394_0[1]),.dinb(w_n1368_0[1]),.dout(n1395),.clk(gclk));
	jxor g1332(.dina(w_n1395_0[1]),.dinb(w_n1366_0[1]),.dout(n1396),.clk(gclk));
	jxor g1333(.dina(w_n1396_0[1]),.dinb(w_n1363_0[1]),.dout(n1397),.clk(gclk));
	jxor g1334(.dina(w_n1397_0[1]),.dinb(w_n1361_0[1]),.dout(n1398),.clk(gclk));
	jxor g1335(.dina(w_n1398_0[1]),.dinb(w_n1358_0[1]),.dout(n1399),.clk(gclk));
	jxor g1336(.dina(w_n1399_0[1]),.dinb(w_n1356_0[1]),.dout(n1400),.clk(gclk));
	jxor g1337(.dina(w_n1400_0[1]),.dinb(w_n1353_0[1]),.dout(n1401),.clk(gclk));
	jxor g1338(.dina(w_n1401_0[1]),.dinb(w_n1351_0[1]),.dout(n1402),.clk(gclk));
	jxor g1339(.dina(w_n1402_0[1]),.dinb(w_n1348_0[1]),.dout(n1403),.clk(gclk));
	jxor g1340(.dina(w_n1403_0[1]),.dinb(w_n1346_0[1]),.dout(n1404),.clk(gclk));
	jxor g1341(.dina(w_n1404_0[1]),.dinb(w_n1343_0[1]),.dout(n1405),.clk(gclk));
	jxor g1342(.dina(w_n1405_0[1]),.dinb(w_n1341_0[1]),.dout(n1406),.clk(gclk));
	jnot g1343(.din(n1406),.dout(n1407),.clk(gclk));
	jxor g1344(.dina(w_n1407_0[1]),.dinb(w_n1338_0[1]),.dout(n1408),.clk(gclk));
	jnot g1345(.din(n1408),.dout(n1409),.clk(gclk));
	jxor g1346(.dina(w_n1409_0[1]),.dinb(w_n1337_0[1]),.dout(n1410),.clk(gclk));
	jxor g1347(.dina(w_n1410_0[1]),.dinb(w_n1332_0[1]),.dout(G6190gat),.clk(gclk));
	jcb g1348(.dina(w_n1409_0[0]),.dinb(w_n1337_0[0]),.dout(n1412));
	jnot g1349(.din(w_n1410_0[0]),.dout(n1413),.clk(gclk));
	jcb g1350(.dina(n1413),.dinb(w_n1332_0[0]),.dout(n1414));
	jand g1351(.dina(n1414),.dinb(w_dff_B_gezxGVAF9_1),.dout(n1415),.clk(gclk));
	jnot g1352(.din(w_n1341_0[0]),.dout(n1416),.clk(gclk));
	jnot g1353(.din(w_n1405_0[0]),.dout(n1417),.clk(gclk));
	jcb g1354(.dina(n1417),.dinb(w_dff_B_ZuB48PZT2_1),.dout(n1418));
	jcb g1355(.dina(w_n1407_0[0]),.dinb(w_n1338_0[0]),.dout(n1419));
	jand g1356(.dina(n1419),.dinb(w_dff_B_c0gKDITm0_1),.dout(n1420),.clk(gclk));
	jand g1357(.dina(w_G528gat_5[1]),.dinb(w_G103gat_2[1]),.dout(n1421),.clk(gclk));
	jand g1358(.dina(w_n1403_0[0]),.dinb(w_n1346_0[0]),.dout(n1422),.clk(gclk));
	jand g1359(.dina(w_n1404_0[0]),.dinb(w_n1343_0[0]),.dout(n1423),.clk(gclk));
	jcb g1360(.dina(n1423),.dinb(w_dff_B_Jch7zrMC4_1),.dout(n1424));
	jand g1361(.dina(w_G511gat_5[0]),.dinb(w_G120gat_2[2]),.dout(n1425),.clk(gclk));
	jnot g1362(.din(n1425),.dout(n1426),.clk(gclk));
	jand g1363(.dina(w_n1401_0[0]),.dinb(w_n1351_0[0]),.dout(n1427),.clk(gclk));
	jand g1364(.dina(w_n1402_0[0]),.dinb(w_n1348_0[0]),.dout(n1428),.clk(gclk));
	jcb g1365(.dina(n1428),.dinb(w_dff_B_PkKGRpPN5_1),.dout(n1429));
	jand g1366(.dina(w_G494gat_4[2]),.dinb(w_G137gat_3[0]),.dout(n1430),.clk(gclk));
	jnot g1367(.din(n1430),.dout(n1431),.clk(gclk));
	jand g1368(.dina(w_n1399_0[0]),.dinb(w_n1356_0[0]),.dout(n1432),.clk(gclk));
	jand g1369(.dina(w_n1400_0[0]),.dinb(w_n1353_0[0]),.dout(n1433),.clk(gclk));
	jcb g1370(.dina(n1433),.dinb(w_dff_B_t9QCbYnh7_1),.dout(n1434));
	jand g1371(.dina(w_G477gat_4[1]),.dinb(w_G154gat_3[1]),.dout(n1435),.clk(gclk));
	jnot g1372(.din(n1435),.dout(n1436),.clk(gclk));
	jand g1373(.dina(w_n1397_0[0]),.dinb(w_n1361_0[0]),.dout(n1437),.clk(gclk));
	jand g1374(.dina(w_n1398_0[0]),.dinb(w_n1358_0[0]),.dout(n1438),.clk(gclk));
	jcb g1375(.dina(n1438),.dinb(w_dff_B_D2vrndJ97_1),.dout(n1439));
	jand g1376(.dina(w_G460gat_4[0]),.dinb(w_G171gat_3[2]),.dout(n1440),.clk(gclk));
	jnot g1377(.din(n1440),.dout(n1441),.clk(gclk));
	jand g1378(.dina(w_n1395_0[0]),.dinb(w_n1366_0[0]),.dout(n1442),.clk(gclk));
	jand g1379(.dina(w_n1396_0[0]),.dinb(w_n1363_0[0]),.dout(n1443),.clk(gclk));
	jcb g1380(.dina(n1443),.dinb(w_dff_B_pHEnIkim6_1),.dout(n1444));
	jand g1381(.dina(w_G443gat_3[2]),.dinb(w_G188gat_4[0]),.dout(n1445),.clk(gclk));
	jnot g1382(.din(n1445),.dout(n1446),.clk(gclk));
	jand g1383(.dina(w_n1393_0[0]),.dinb(w_n1371_0[0]),.dout(n1447),.clk(gclk));
	jand g1384(.dina(w_n1394_0[0]),.dinb(w_n1368_0[0]),.dout(n1448),.clk(gclk));
	jcb g1385(.dina(n1448),.dinb(w_dff_B_aqaLGXOT4_1),.dout(n1449));
	jand g1386(.dina(w_G426gat_3[1]),.dinb(w_G205gat_4[1]),.dout(n1450),.clk(gclk));
	jnot g1387(.din(n1450),.dout(n1451),.clk(gclk));
	jand g1388(.dina(w_n1391_0[0]),.dinb(w_n1376_0[0]),.dout(n1452),.clk(gclk));
	jand g1389(.dina(w_n1392_0[0]),.dinb(w_n1373_0[0]),.dout(n1453),.clk(gclk));
	jcb g1390(.dina(n1453),.dinb(w_dff_B_sh0dxksO2_1),.dout(n1454));
	jand g1391(.dina(w_G409gat_3[0]),.dinb(w_G222gat_4[2]),.dout(n1455),.clk(gclk));
	jnot g1392(.din(n1455),.dout(n1456),.clk(gclk));
	jand g1393(.dina(w_n1389_0[0]),.dinb(w_n1381_0[0]),.dout(n1457),.clk(gclk));
	jand g1394(.dina(w_n1390_0[0]),.dinb(w_n1378_0[0]),.dout(n1458),.clk(gclk));
	jcb g1395(.dina(n1458),.dinb(w_dff_B_85e2vVXL1_1),.dout(n1459));
	jand g1396(.dina(w_G392gat_2[2]),.dinb(w_G239gat_5[0]),.dout(n1460),.clk(gclk));
	jand g1397(.dina(w_G375gat_2[1]),.dinb(w_G256gat_5[1]),.dout(n1461),.clk(gclk));
	jcb g1398(.dina(w_n1386_0[0]),.dinb(w_n1383_0[0]),.dout(n1462));
	jcb g1399(.dina(w_n1388_0[0]),.dinb(w_n1382_0[0]),.dout(n1463));
	jand g1400(.dina(n1463),.dinb(w_dff_B_zYK4DSNq2_1),.dout(n1464),.clk(gclk));
	jxor g1401(.dina(w_n1464_0[1]),.dinb(w_n1461_0[1]),.dout(n1465),.clk(gclk));
	jnot g1402(.din(n1465),.dout(n1466),.clk(gclk));
	jxor g1403(.dina(w_n1466_0[1]),.dinb(w_n1460_0[1]),.dout(n1467),.clk(gclk));
	jxor g1404(.dina(w_n1467_0[1]),.dinb(w_n1459_0[1]),.dout(n1468),.clk(gclk));
	jxor g1405(.dina(w_n1468_0[1]),.dinb(w_n1456_0[1]),.dout(n1469),.clk(gclk));
	jxor g1406(.dina(w_n1469_0[1]),.dinb(w_n1454_0[1]),.dout(n1470),.clk(gclk));
	jxor g1407(.dina(w_n1470_0[1]),.dinb(w_n1451_0[1]),.dout(n1471),.clk(gclk));
	jxor g1408(.dina(w_n1471_0[1]),.dinb(w_n1449_0[1]),.dout(n1472),.clk(gclk));
	jxor g1409(.dina(w_n1472_0[1]),.dinb(w_n1446_0[1]),.dout(n1473),.clk(gclk));
	jxor g1410(.dina(w_n1473_0[1]),.dinb(w_n1444_0[1]),.dout(n1474),.clk(gclk));
	jxor g1411(.dina(w_n1474_0[1]),.dinb(w_n1441_0[1]),.dout(n1475),.clk(gclk));
	jxor g1412(.dina(w_n1475_0[1]),.dinb(w_n1439_0[1]),.dout(n1476),.clk(gclk));
	jxor g1413(.dina(w_n1476_0[1]),.dinb(w_n1436_0[1]),.dout(n1477),.clk(gclk));
	jxor g1414(.dina(w_n1477_0[1]),.dinb(w_n1434_0[1]),.dout(n1478),.clk(gclk));
	jxor g1415(.dina(w_n1478_0[1]),.dinb(w_n1431_0[1]),.dout(n1479),.clk(gclk));
	jxor g1416(.dina(w_n1479_0[1]),.dinb(w_n1429_0[1]),.dout(n1480),.clk(gclk));
	jxor g1417(.dina(w_n1480_0[1]),.dinb(w_n1426_0[1]),.dout(n1481),.clk(gclk));
	jxor g1418(.dina(w_n1481_0[1]),.dinb(w_n1424_0[1]),.dout(n1482),.clk(gclk));
	jnot g1419(.din(n1482),.dout(n1483),.clk(gclk));
	jxor g1420(.dina(w_n1483_0[1]),.dinb(w_n1421_0[1]),.dout(n1484),.clk(gclk));
	jnot g1421(.din(n1484),.dout(n1485),.clk(gclk));
	jxor g1422(.dina(w_n1485_0[1]),.dinb(w_n1420_0[1]),.dout(n1486),.clk(gclk));
	jxor g1423(.dina(w_n1486_0[1]),.dinb(w_n1415_0[1]),.dout(G6200gat),.clk(gclk));
	jcb g1424(.dina(w_n1485_0[0]),.dinb(w_n1420_0[0]),.dout(n1488));
	jnot g1425(.din(w_n1486_0[0]),.dout(n1489),.clk(gclk));
	jcb g1426(.dina(n1489),.dinb(w_n1415_0[0]),.dout(n1490));
	jand g1427(.dina(n1490),.dinb(w_dff_B_3ViiBqlr3_1),.dout(n1491),.clk(gclk));
	jnot g1428(.din(w_n1424_0[0]),.dout(n1492),.clk(gclk));
	jnot g1429(.din(w_n1481_0[0]),.dout(n1493),.clk(gclk));
	jcb g1430(.dina(n1493),.dinb(w_dff_B_5MuID1Q30_1),.dout(n1494));
	jcb g1431(.dina(w_n1483_0[0]),.dinb(w_n1421_0[0]),.dout(n1495));
	jand g1432(.dina(n1495),.dinb(w_dff_B_Wc61OfOK0_1),.dout(n1496),.clk(gclk));
	jand g1433(.dina(w_G528gat_5[0]),.dinb(w_G120gat_2[1]),.dout(n1497),.clk(gclk));
	jand g1434(.dina(w_n1479_0[0]),.dinb(w_n1429_0[0]),.dout(n1498),.clk(gclk));
	jand g1435(.dina(w_n1480_0[0]),.dinb(w_n1426_0[0]),.dout(n1499),.clk(gclk));
	jcb g1436(.dina(n1499),.dinb(w_dff_B_mFNHx6He1_1),.dout(n1500));
	jand g1437(.dina(w_G511gat_4[2]),.dinb(w_G137gat_2[2]),.dout(n1501),.clk(gclk));
	jnot g1438(.din(n1501),.dout(n1502),.clk(gclk));
	jand g1439(.dina(w_n1477_0[0]),.dinb(w_n1434_0[0]),.dout(n1503),.clk(gclk));
	jand g1440(.dina(w_n1478_0[0]),.dinb(w_n1431_0[0]),.dout(n1504),.clk(gclk));
	jcb g1441(.dina(n1504),.dinb(w_dff_B_Mfh0kkv02_1),.dout(n1505));
	jand g1442(.dina(w_G494gat_4[1]),.dinb(w_G154gat_3[0]),.dout(n1506),.clk(gclk));
	jnot g1443(.din(n1506),.dout(n1507),.clk(gclk));
	jand g1444(.dina(w_n1475_0[0]),.dinb(w_n1439_0[0]),.dout(n1508),.clk(gclk));
	jand g1445(.dina(w_n1476_0[0]),.dinb(w_n1436_0[0]),.dout(n1509),.clk(gclk));
	jcb g1446(.dina(n1509),.dinb(w_dff_B_GPX5xaK20_1),.dout(n1510));
	jand g1447(.dina(w_G477gat_4[0]),.dinb(w_G171gat_3[1]),.dout(n1511),.clk(gclk));
	jnot g1448(.din(n1511),.dout(n1512),.clk(gclk));
	jand g1449(.dina(w_n1473_0[0]),.dinb(w_n1444_0[0]),.dout(n1513),.clk(gclk));
	jand g1450(.dina(w_n1474_0[0]),.dinb(w_n1441_0[0]),.dout(n1514),.clk(gclk));
	jcb g1451(.dina(n1514),.dinb(w_dff_B_ldo93EOQ0_1),.dout(n1515));
	jand g1452(.dina(w_G460gat_3[2]),.dinb(w_G188gat_3[2]),.dout(n1516),.clk(gclk));
	jnot g1453(.din(n1516),.dout(n1517),.clk(gclk));
	jand g1454(.dina(w_n1471_0[0]),.dinb(w_n1449_0[0]),.dout(n1518),.clk(gclk));
	jand g1455(.dina(w_n1472_0[0]),.dinb(w_n1446_0[0]),.dout(n1519),.clk(gclk));
	jcb g1456(.dina(n1519),.dinb(w_dff_B_zXMfh2tW4_1),.dout(n1520));
	jand g1457(.dina(w_G443gat_3[1]),.dinb(w_G205gat_4[0]),.dout(n1521),.clk(gclk));
	jnot g1458(.din(n1521),.dout(n1522),.clk(gclk));
	jand g1459(.dina(w_n1469_0[0]),.dinb(w_n1454_0[0]),.dout(n1523),.clk(gclk));
	jand g1460(.dina(w_n1470_0[0]),.dinb(w_n1451_0[0]),.dout(n1524),.clk(gclk));
	jcb g1461(.dina(n1524),.dinb(w_dff_B_6dviGXV86_1),.dout(n1525));
	jand g1462(.dina(w_G426gat_3[0]),.dinb(w_G222gat_4[1]),.dout(n1526),.clk(gclk));
	jnot g1463(.din(n1526),.dout(n1527),.clk(gclk));
	jand g1464(.dina(w_n1467_0[0]),.dinb(w_n1459_0[0]),.dout(n1528),.clk(gclk));
	jand g1465(.dina(w_n1468_0[0]),.dinb(w_n1456_0[0]),.dout(n1529),.clk(gclk));
	jcb g1466(.dina(n1529),.dinb(w_dff_B_0LPPkpTF8_1),.dout(n1530));
	jand g1467(.dina(w_G409gat_2[2]),.dinb(w_G239gat_4[2]),.dout(n1531),.clk(gclk));
	jand g1468(.dina(w_G392gat_2[1]),.dinb(w_G256gat_5[0]),.dout(n1532),.clk(gclk));
	jcb g1469(.dina(w_n1464_0[0]),.dinb(w_n1461_0[0]),.dout(n1533));
	jcb g1470(.dina(w_n1466_0[0]),.dinb(w_n1460_0[0]),.dout(n1534));
	jand g1471(.dina(n1534),.dinb(w_dff_B_CsrK5ZqW4_1),.dout(n1535),.clk(gclk));
	jxor g1472(.dina(w_n1535_0[1]),.dinb(w_n1532_0[1]),.dout(n1536),.clk(gclk));
	jnot g1473(.din(n1536),.dout(n1537),.clk(gclk));
	jxor g1474(.dina(w_n1537_0[1]),.dinb(w_n1531_0[1]),.dout(n1538),.clk(gclk));
	jxor g1475(.dina(w_n1538_0[1]),.dinb(w_n1530_0[1]),.dout(n1539),.clk(gclk));
	jxor g1476(.dina(w_n1539_0[1]),.dinb(w_n1527_0[1]),.dout(n1540),.clk(gclk));
	jxor g1477(.dina(w_n1540_0[1]),.dinb(w_n1525_0[1]),.dout(n1541),.clk(gclk));
	jxor g1478(.dina(w_n1541_0[1]),.dinb(w_n1522_0[1]),.dout(n1542),.clk(gclk));
	jxor g1479(.dina(w_n1542_0[1]),.dinb(w_n1520_0[1]),.dout(n1543),.clk(gclk));
	jxor g1480(.dina(w_n1543_0[1]),.dinb(w_n1517_0[1]),.dout(n1544),.clk(gclk));
	jxor g1481(.dina(w_n1544_0[1]),.dinb(w_n1515_0[1]),.dout(n1545),.clk(gclk));
	jxor g1482(.dina(w_n1545_0[1]),.dinb(w_n1512_0[1]),.dout(n1546),.clk(gclk));
	jxor g1483(.dina(w_n1546_0[1]),.dinb(w_n1510_0[1]),.dout(n1547),.clk(gclk));
	jxor g1484(.dina(w_n1547_0[1]),.dinb(w_n1507_0[1]),.dout(n1548),.clk(gclk));
	jxor g1485(.dina(w_n1548_0[1]),.dinb(w_n1505_0[1]),.dout(n1549),.clk(gclk));
	jxor g1486(.dina(w_n1549_0[1]),.dinb(w_n1502_0[1]),.dout(n1550),.clk(gclk));
	jxor g1487(.dina(w_n1550_0[1]),.dinb(w_n1500_0[1]),.dout(n1551),.clk(gclk));
	jnot g1488(.din(n1551),.dout(n1552),.clk(gclk));
	jxor g1489(.dina(w_n1552_0[1]),.dinb(w_n1497_0[1]),.dout(n1553),.clk(gclk));
	jnot g1490(.din(n1553),.dout(n1554),.clk(gclk));
	jxor g1491(.dina(w_n1554_0[1]),.dinb(w_n1496_0[1]),.dout(n1555),.clk(gclk));
	jxor g1492(.dina(w_n1555_0[1]),.dinb(w_n1491_0[1]),.dout(G6210gat),.clk(gclk));
	jcb g1493(.dina(w_n1554_0[0]),.dinb(w_n1496_0[0]),.dout(n1557));
	jnot g1494(.din(w_n1555_0[0]),.dout(n1558),.clk(gclk));
	jcb g1495(.dina(n1558),.dinb(w_n1491_0[0]),.dout(n1559));
	jand g1496(.dina(n1559),.dinb(w_dff_B_mmxUZK7d1_1),.dout(n1560),.clk(gclk));
	jnot g1497(.din(w_n1500_0[0]),.dout(n1561),.clk(gclk));
	jnot g1498(.din(w_n1550_0[0]),.dout(n1562),.clk(gclk));
	jcb g1499(.dina(n1562),.dinb(w_dff_B_d35o9utC8_1),.dout(n1563));
	jcb g1500(.dina(w_n1552_0[0]),.dinb(w_n1497_0[0]),.dout(n1564));
	jand g1501(.dina(n1564),.dinb(w_dff_B_Ha4dA8CP6_1),.dout(n1565),.clk(gclk));
	jand g1502(.dina(w_G528gat_4[2]),.dinb(w_G137gat_2[1]),.dout(n1566),.clk(gclk));
	jand g1503(.dina(w_n1548_0[0]),.dinb(w_n1505_0[0]),.dout(n1567),.clk(gclk));
	jand g1504(.dina(w_n1549_0[0]),.dinb(w_n1502_0[0]),.dout(n1568),.clk(gclk));
	jcb g1505(.dina(n1568),.dinb(w_dff_B_9d5lIpiV0_1),.dout(n1569));
	jand g1506(.dina(w_G511gat_4[1]),.dinb(w_G154gat_2[2]),.dout(n1570),.clk(gclk));
	jnot g1507(.din(n1570),.dout(n1571),.clk(gclk));
	jand g1508(.dina(w_n1546_0[0]),.dinb(w_n1510_0[0]),.dout(n1572),.clk(gclk));
	jand g1509(.dina(w_n1547_0[0]),.dinb(w_n1507_0[0]),.dout(n1573),.clk(gclk));
	jcb g1510(.dina(n1573),.dinb(w_dff_B_uzlAELXW4_1),.dout(n1574));
	jand g1511(.dina(w_G494gat_4[0]),.dinb(w_G171gat_3[0]),.dout(n1575),.clk(gclk));
	jnot g1512(.din(n1575),.dout(n1576),.clk(gclk));
	jand g1513(.dina(w_n1544_0[0]),.dinb(w_n1515_0[0]),.dout(n1577),.clk(gclk));
	jand g1514(.dina(w_n1545_0[0]),.dinb(w_n1512_0[0]),.dout(n1578),.clk(gclk));
	jcb g1515(.dina(n1578),.dinb(w_dff_B_jYStSG8v5_1),.dout(n1579));
	jand g1516(.dina(w_G477gat_3[2]),.dinb(w_G188gat_3[1]),.dout(n1580),.clk(gclk));
	jnot g1517(.din(n1580),.dout(n1581),.clk(gclk));
	jand g1518(.dina(w_n1542_0[0]),.dinb(w_n1520_0[0]),.dout(n1582),.clk(gclk));
	jand g1519(.dina(w_n1543_0[0]),.dinb(w_n1517_0[0]),.dout(n1583),.clk(gclk));
	jcb g1520(.dina(n1583),.dinb(w_dff_B_Nlcbd72D3_1),.dout(n1584));
	jand g1521(.dina(w_G460gat_3[1]),.dinb(w_G205gat_3[2]),.dout(n1585),.clk(gclk));
	jnot g1522(.din(n1585),.dout(n1586),.clk(gclk));
	jand g1523(.dina(w_n1540_0[0]),.dinb(w_n1525_0[0]),.dout(n1587),.clk(gclk));
	jand g1524(.dina(w_n1541_0[0]),.dinb(w_n1522_0[0]),.dout(n1588),.clk(gclk));
	jcb g1525(.dina(n1588),.dinb(w_dff_B_t7lINx934_1),.dout(n1589));
	jand g1526(.dina(w_G443gat_3[0]),.dinb(w_G222gat_4[0]),.dout(n1590),.clk(gclk));
	jnot g1527(.din(n1590),.dout(n1591),.clk(gclk));
	jand g1528(.dina(w_n1538_0[0]),.dinb(w_n1530_0[0]),.dout(n1592),.clk(gclk));
	jand g1529(.dina(w_n1539_0[0]),.dinb(w_n1527_0[0]),.dout(n1593),.clk(gclk));
	jcb g1530(.dina(n1593),.dinb(w_dff_B_s0iMEh9j6_1),.dout(n1594));
	jand g1531(.dina(w_G426gat_2[2]),.dinb(w_G239gat_4[1]),.dout(n1595),.clk(gclk));
	jand g1532(.dina(w_G409gat_2[1]),.dinb(w_G256gat_4[2]),.dout(n1596),.clk(gclk));
	jcb g1533(.dina(w_n1535_0[0]),.dinb(w_n1532_0[0]),.dout(n1597));
	jcb g1534(.dina(w_n1537_0[0]),.dinb(w_n1531_0[0]),.dout(n1598));
	jand g1535(.dina(n1598),.dinb(w_dff_B_KARzh2LJ3_1),.dout(n1599),.clk(gclk));
	jxor g1536(.dina(w_n1599_0[1]),.dinb(w_n1596_0[1]),.dout(n1600),.clk(gclk));
	jnot g1537(.din(n1600),.dout(n1601),.clk(gclk));
	jxor g1538(.dina(w_n1601_0[1]),.dinb(w_n1595_0[1]),.dout(n1602),.clk(gclk));
	jxor g1539(.dina(w_n1602_0[1]),.dinb(w_n1594_0[1]),.dout(n1603),.clk(gclk));
	jxor g1540(.dina(w_n1603_0[1]),.dinb(w_n1591_0[1]),.dout(n1604),.clk(gclk));
	jxor g1541(.dina(w_n1604_0[1]),.dinb(w_n1589_0[1]),.dout(n1605),.clk(gclk));
	jxor g1542(.dina(w_n1605_0[1]),.dinb(w_n1586_0[1]),.dout(n1606),.clk(gclk));
	jxor g1543(.dina(w_n1606_0[1]),.dinb(w_n1584_0[1]),.dout(n1607),.clk(gclk));
	jxor g1544(.dina(w_n1607_0[1]),.dinb(w_n1581_0[1]),.dout(n1608),.clk(gclk));
	jxor g1545(.dina(w_n1608_0[1]),.dinb(w_n1579_0[1]),.dout(n1609),.clk(gclk));
	jxor g1546(.dina(w_n1609_0[1]),.dinb(w_n1576_0[1]),.dout(n1610),.clk(gclk));
	jxor g1547(.dina(w_n1610_0[1]),.dinb(w_n1574_0[1]),.dout(n1611),.clk(gclk));
	jxor g1548(.dina(w_n1611_0[1]),.dinb(w_n1571_0[1]),.dout(n1612),.clk(gclk));
	jxor g1549(.dina(w_n1612_0[1]),.dinb(w_n1569_0[1]),.dout(n1613),.clk(gclk));
	jnot g1550(.din(n1613),.dout(n1614),.clk(gclk));
	jxor g1551(.dina(w_n1614_0[1]),.dinb(w_n1566_0[1]),.dout(n1615),.clk(gclk));
	jnot g1552(.din(n1615),.dout(n1616),.clk(gclk));
	jxor g1553(.dina(w_n1616_0[1]),.dinb(w_n1565_0[1]),.dout(n1617),.clk(gclk));
	jxor g1554(.dina(w_n1617_0[1]),.dinb(w_n1560_0[1]),.dout(G6220gat),.clk(gclk));
	jcb g1555(.dina(w_n1616_0[0]),.dinb(w_n1565_0[0]),.dout(n1619));
	jnot g1556(.din(w_n1617_0[0]),.dout(n1620),.clk(gclk));
	jcb g1557(.dina(n1620),.dinb(w_n1560_0[0]),.dout(n1621));
	jand g1558(.dina(n1621),.dinb(w_dff_B_FrfsuDlV9_1),.dout(n1622),.clk(gclk));
	jnot g1559(.din(w_n1569_0[0]),.dout(n1623),.clk(gclk));
	jnot g1560(.din(w_n1612_0[0]),.dout(n1624),.clk(gclk));
	jcb g1561(.dina(n1624),.dinb(w_dff_B_PPlTCACc9_1),.dout(n1625));
	jcb g1562(.dina(w_n1614_0[0]),.dinb(w_n1566_0[0]),.dout(n1626));
	jand g1563(.dina(n1626),.dinb(w_dff_B_OXtOuo0n0_1),.dout(n1627),.clk(gclk));
	jand g1564(.dina(w_G528gat_4[1]),.dinb(w_G154gat_2[1]),.dout(n1628),.clk(gclk));
	jand g1565(.dina(w_n1610_0[0]),.dinb(w_n1574_0[0]),.dout(n1629),.clk(gclk));
	jand g1566(.dina(w_n1611_0[0]),.dinb(w_n1571_0[0]),.dout(n1630),.clk(gclk));
	jcb g1567(.dina(n1630),.dinb(w_dff_B_w79I0pZh7_1),.dout(n1631));
	jand g1568(.dina(w_G511gat_4[0]),.dinb(w_G171gat_2[2]),.dout(n1632),.clk(gclk));
	jnot g1569(.din(n1632),.dout(n1633),.clk(gclk));
	jand g1570(.dina(w_n1608_0[0]),.dinb(w_n1579_0[0]),.dout(n1634),.clk(gclk));
	jand g1571(.dina(w_n1609_0[0]),.dinb(w_n1576_0[0]),.dout(n1635),.clk(gclk));
	jcb g1572(.dina(n1635),.dinb(w_dff_B_nZYIJf9U5_1),.dout(n1636));
	jand g1573(.dina(w_G494gat_3[2]),.dinb(w_G188gat_3[0]),.dout(n1637),.clk(gclk));
	jnot g1574(.din(n1637),.dout(n1638),.clk(gclk));
	jand g1575(.dina(w_n1606_0[0]),.dinb(w_n1584_0[0]),.dout(n1639),.clk(gclk));
	jand g1576(.dina(w_n1607_0[0]),.dinb(w_n1581_0[0]),.dout(n1640),.clk(gclk));
	jcb g1577(.dina(n1640),.dinb(w_dff_B_iOqyTgmz1_1),.dout(n1641));
	jand g1578(.dina(w_G477gat_3[1]),.dinb(w_G205gat_3[1]),.dout(n1642),.clk(gclk));
	jnot g1579(.din(n1642),.dout(n1643),.clk(gclk));
	jand g1580(.dina(w_n1604_0[0]),.dinb(w_n1589_0[0]),.dout(n1644),.clk(gclk));
	jand g1581(.dina(w_n1605_0[0]),.dinb(w_n1586_0[0]),.dout(n1645),.clk(gclk));
	jcb g1582(.dina(n1645),.dinb(w_dff_B_1zuIz7yN8_1),.dout(n1646));
	jand g1583(.dina(w_G460gat_3[0]),.dinb(w_G222gat_3[2]),.dout(n1647),.clk(gclk));
	jnot g1584(.din(n1647),.dout(n1648),.clk(gclk));
	jand g1585(.dina(w_n1602_0[0]),.dinb(w_n1594_0[0]),.dout(n1649),.clk(gclk));
	jand g1586(.dina(w_n1603_0[0]),.dinb(w_n1591_0[0]),.dout(n1650),.clk(gclk));
	jcb g1587(.dina(n1650),.dinb(w_dff_B_8AToENM26_1),.dout(n1651));
	jand g1588(.dina(w_G443gat_2[2]),.dinb(w_G239gat_4[0]),.dout(n1652),.clk(gclk));
	jand g1589(.dina(w_G426gat_2[1]),.dinb(w_G256gat_4[1]),.dout(n1653),.clk(gclk));
	jcb g1590(.dina(w_n1599_0[0]),.dinb(w_n1596_0[0]),.dout(n1654));
	jcb g1591(.dina(w_n1601_0[0]),.dinb(w_n1595_0[0]),.dout(n1655));
	jand g1592(.dina(n1655),.dinb(w_dff_B_3KAZd9Je8_1),.dout(n1656),.clk(gclk));
	jxor g1593(.dina(w_n1656_0[1]),.dinb(w_n1653_0[1]),.dout(n1657),.clk(gclk));
	jnot g1594(.din(n1657),.dout(n1658),.clk(gclk));
	jxor g1595(.dina(w_n1658_0[1]),.dinb(w_n1652_0[1]),.dout(n1659),.clk(gclk));
	jxor g1596(.dina(w_n1659_0[1]),.dinb(w_n1651_0[1]),.dout(n1660),.clk(gclk));
	jxor g1597(.dina(w_n1660_0[1]),.dinb(w_n1648_0[1]),.dout(n1661),.clk(gclk));
	jxor g1598(.dina(w_n1661_0[1]),.dinb(w_n1646_0[1]),.dout(n1662),.clk(gclk));
	jxor g1599(.dina(w_n1662_0[1]),.dinb(w_n1643_0[1]),.dout(n1663),.clk(gclk));
	jxor g1600(.dina(w_n1663_0[1]),.dinb(w_n1641_0[1]),.dout(n1664),.clk(gclk));
	jxor g1601(.dina(w_n1664_0[1]),.dinb(w_n1638_0[1]),.dout(n1665),.clk(gclk));
	jxor g1602(.dina(w_n1665_0[1]),.dinb(w_n1636_0[1]),.dout(n1666),.clk(gclk));
	jxor g1603(.dina(w_n1666_0[1]),.dinb(w_n1633_0[1]),.dout(n1667),.clk(gclk));
	jxor g1604(.dina(w_n1667_0[1]),.dinb(w_n1631_0[1]),.dout(n1668),.clk(gclk));
	jnot g1605(.din(n1668),.dout(n1669),.clk(gclk));
	jxor g1606(.dina(w_n1669_0[1]),.dinb(w_n1628_0[1]),.dout(n1670),.clk(gclk));
	jnot g1607(.din(n1670),.dout(n1671),.clk(gclk));
	jxor g1608(.dina(w_n1671_0[1]),.dinb(w_n1627_0[1]),.dout(n1672),.clk(gclk));
	jxor g1609(.dina(w_n1672_0[1]),.dinb(w_n1622_0[1]),.dout(G6230gat),.clk(gclk));
	jcb g1610(.dina(w_n1671_0[0]),.dinb(w_n1627_0[0]),.dout(n1674));
	jnot g1611(.din(w_n1672_0[0]),.dout(n1675),.clk(gclk));
	jcb g1612(.dina(n1675),.dinb(w_n1622_0[0]),.dout(n1676));
	jand g1613(.dina(n1676),.dinb(w_dff_B_4vwGwDhX0_1),.dout(n1677),.clk(gclk));
	jnot g1614(.din(w_n1631_0[0]),.dout(n1678),.clk(gclk));
	jnot g1615(.din(w_n1667_0[0]),.dout(n1679),.clk(gclk));
	jcb g1616(.dina(n1679),.dinb(w_dff_B_VtmnVXvW9_1),.dout(n1680));
	jcb g1617(.dina(w_n1669_0[0]),.dinb(w_n1628_0[0]),.dout(n1681));
	jand g1618(.dina(n1681),.dinb(w_dff_B_oDu8Eos25_1),.dout(n1682),.clk(gclk));
	jand g1619(.dina(w_G528gat_4[0]),.dinb(w_G171gat_2[1]),.dout(n1683),.clk(gclk));
	jnot g1620(.din(n1683),.dout(n1684),.clk(gclk));
	jand g1621(.dina(w_n1665_0[0]),.dinb(w_n1636_0[0]),.dout(n1685),.clk(gclk));
	jand g1622(.dina(w_n1666_0[0]),.dinb(w_n1633_0[0]),.dout(n1686),.clk(gclk));
	jcb g1623(.dina(n1686),.dinb(w_dff_B_UJvMBvYk0_1),.dout(n1687));
	jand g1624(.dina(w_G511gat_3[2]),.dinb(w_G188gat_2[2]),.dout(n1688),.clk(gclk));
	jnot g1625(.din(n1688),.dout(n1689),.clk(gclk));
	jand g1626(.dina(w_n1663_0[0]),.dinb(w_n1641_0[0]),.dout(n1690),.clk(gclk));
	jand g1627(.dina(w_n1664_0[0]),.dinb(w_n1638_0[0]),.dout(n1691),.clk(gclk));
	jcb g1628(.dina(n1691),.dinb(w_dff_B_xMcZA4CE3_1),.dout(n1692));
	jand g1629(.dina(w_G494gat_3[1]),.dinb(w_G205gat_3[0]),.dout(n1693),.clk(gclk));
	jnot g1630(.din(n1693),.dout(n1694),.clk(gclk));
	jand g1631(.dina(w_n1661_0[0]),.dinb(w_n1646_0[0]),.dout(n1695),.clk(gclk));
	jand g1632(.dina(w_n1662_0[0]),.dinb(w_n1643_0[0]),.dout(n1696),.clk(gclk));
	jcb g1633(.dina(n1696),.dinb(w_dff_B_OwlYxgy72_1),.dout(n1697));
	jand g1634(.dina(w_G477gat_3[0]),.dinb(w_G222gat_3[1]),.dout(n1698),.clk(gclk));
	jnot g1635(.din(n1698),.dout(n1699),.clk(gclk));
	jand g1636(.dina(w_n1659_0[0]),.dinb(w_n1651_0[0]),.dout(n1700),.clk(gclk));
	jand g1637(.dina(w_n1660_0[0]),.dinb(w_n1648_0[0]),.dout(n1701),.clk(gclk));
	jcb g1638(.dina(n1701),.dinb(w_dff_B_VbSDAllf5_1),.dout(n1702));
	jand g1639(.dina(w_G460gat_2[2]),.dinb(w_G239gat_3[2]),.dout(n1703),.clk(gclk));
	jand g1640(.dina(w_G443gat_2[1]),.dinb(w_G256gat_4[0]),.dout(n1704),.clk(gclk));
	jcb g1641(.dina(w_n1656_0[0]),.dinb(w_n1653_0[0]),.dout(n1705));
	jcb g1642(.dina(w_n1658_0[0]),.dinb(w_n1652_0[0]),.dout(n1706));
	jand g1643(.dina(n1706),.dinb(w_dff_B_YErMqfjS7_1),.dout(n1707),.clk(gclk));
	jxor g1644(.dina(w_n1707_0[1]),.dinb(w_n1704_0[1]),.dout(n1708),.clk(gclk));
	jnot g1645(.din(n1708),.dout(n1709),.clk(gclk));
	jxor g1646(.dina(w_n1709_0[1]),.dinb(w_n1703_0[1]),.dout(n1710),.clk(gclk));
	jxor g1647(.dina(w_n1710_0[1]),.dinb(w_n1702_0[1]),.dout(n1711),.clk(gclk));
	jxor g1648(.dina(w_n1711_0[1]),.dinb(w_n1699_0[1]),.dout(n1712),.clk(gclk));
	jxor g1649(.dina(w_n1712_0[1]),.dinb(w_n1697_0[1]),.dout(n1713),.clk(gclk));
	jxor g1650(.dina(w_n1713_0[1]),.dinb(w_n1694_0[1]),.dout(n1714),.clk(gclk));
	jxor g1651(.dina(w_n1714_0[1]),.dinb(w_n1692_0[1]),.dout(n1715),.clk(gclk));
	jxor g1652(.dina(w_n1715_0[1]),.dinb(w_n1689_0[1]),.dout(n1716),.clk(gclk));
	jxor g1653(.dina(w_n1716_0[1]),.dinb(w_n1687_0[1]),.dout(n1717),.clk(gclk));
	jxor g1654(.dina(w_n1717_0[1]),.dinb(w_n1684_0[1]),.dout(n1718),.clk(gclk));
	jnot g1655(.din(n1718),.dout(n1719),.clk(gclk));
	jxor g1656(.dina(w_n1719_0[1]),.dinb(w_n1682_0[1]),.dout(n1720),.clk(gclk));
	jxor g1657(.dina(w_n1720_0[1]),.dinb(w_n1677_0[1]),.dout(G6240gat),.clk(gclk));
	jcb g1658(.dina(w_n1719_0[0]),.dinb(w_n1682_0[0]),.dout(n1722));
	jnot g1659(.din(w_n1720_0[0]),.dout(n1723),.clk(gclk));
	jcb g1660(.dina(w_dff_B_wNIJnD189_0),.dinb(w_n1677_0[0]),.dout(n1724));
	jand g1661(.dina(n1724),.dinb(w_dff_B_FDF2le2Q4_1),.dout(n1725),.clk(gclk));
	jand g1662(.dina(w_n1716_0[0]),.dinb(w_n1687_0[0]),.dout(n1726),.clk(gclk));
	jand g1663(.dina(w_n1717_0[0]),.dinb(w_n1684_0[0]),.dout(n1727),.clk(gclk));
	jcb g1664(.dina(n1727),.dinb(w_dff_B_qjFxCdra6_1),.dout(n1728));
	jand g1665(.dina(w_G528gat_3[2]),.dinb(w_G188gat_2[1]),.dout(n1729),.clk(gclk));
	jnot g1666(.din(n1729),.dout(n1730),.clk(gclk));
	jand g1667(.dina(w_n1714_0[0]),.dinb(w_n1692_0[0]),.dout(n1731),.clk(gclk));
	jand g1668(.dina(w_n1715_0[0]),.dinb(w_n1689_0[0]),.dout(n1732),.clk(gclk));
	jcb g1669(.dina(n1732),.dinb(w_dff_B_2il5fWCi4_1),.dout(n1733));
	jand g1670(.dina(w_G511gat_3[1]),.dinb(w_G205gat_2[2]),.dout(n1734),.clk(gclk));
	jnot g1671(.din(n1734),.dout(n1735),.clk(gclk));
	jand g1672(.dina(w_n1712_0[0]),.dinb(w_n1697_0[0]),.dout(n1736),.clk(gclk));
	jand g1673(.dina(w_n1713_0[0]),.dinb(w_n1694_0[0]),.dout(n1737),.clk(gclk));
	jcb g1674(.dina(n1737),.dinb(w_dff_B_iuLwvLhL0_1),.dout(n1738));
	jand g1675(.dina(w_G494gat_3[0]),.dinb(w_G222gat_3[0]),.dout(n1739),.clk(gclk));
	jnot g1676(.din(n1739),.dout(n1740),.clk(gclk));
	jand g1677(.dina(w_n1710_0[0]),.dinb(w_n1702_0[0]),.dout(n1741),.clk(gclk));
	jand g1678(.dina(w_n1711_0[0]),.dinb(w_n1699_0[0]),.dout(n1742),.clk(gclk));
	jcb g1679(.dina(n1742),.dinb(w_dff_B_IzfRDnTa7_1),.dout(n1743));
	jand g1680(.dina(w_G477gat_2[2]),.dinb(w_G239gat_3[1]),.dout(n1744),.clk(gclk));
	jand g1681(.dina(w_G460gat_2[1]),.dinb(w_G256gat_3[2]),.dout(n1745),.clk(gclk));
	jcb g1682(.dina(w_n1707_0[0]),.dinb(w_n1704_0[0]),.dout(n1746));
	jcb g1683(.dina(w_n1709_0[0]),.dinb(w_n1703_0[0]),.dout(n1747));
	jand g1684(.dina(n1747),.dinb(w_dff_B_Nayzih5N8_1),.dout(n1748),.clk(gclk));
	jxor g1685(.dina(w_n1748_0[1]),.dinb(w_n1745_0[1]),.dout(n1749),.clk(gclk));
	jnot g1686(.din(n1749),.dout(n1750),.clk(gclk));
	jxor g1687(.dina(w_n1750_0[1]),.dinb(w_n1744_0[1]),.dout(n1751),.clk(gclk));
	jxor g1688(.dina(w_n1751_0[1]),.dinb(w_n1743_0[1]),.dout(n1752),.clk(gclk));
	jxor g1689(.dina(w_n1752_0[1]),.dinb(w_n1740_0[1]),.dout(n1753),.clk(gclk));
	jxor g1690(.dina(w_n1753_0[1]),.dinb(w_n1738_0[1]),.dout(n1754),.clk(gclk));
	jxor g1691(.dina(w_n1754_0[1]),.dinb(w_n1735_0[1]),.dout(n1755),.clk(gclk));
	jxor g1692(.dina(w_n1755_0[1]),.dinb(w_n1733_0[1]),.dout(n1756),.clk(gclk));
	jxor g1693(.dina(w_n1756_0[1]),.dinb(w_n1730_0[1]),.dout(n1757),.clk(gclk));
	jxor g1694(.dina(w_n1757_0[1]),.dinb(w_n1728_0[1]),.dout(n1758),.clk(gclk));
	jxor g1695(.dina(w_n1758_0[1]),.dinb(w_n1725_0[1]),.dout(G6250gat),.clk(gclk));
	jnot g1696(.din(w_n1728_0[0]),.dout(n1760),.clk(gclk));
	jnot g1697(.din(w_n1757_0[0]),.dout(n1761),.clk(gclk));
	jcb g1698(.dina(n1761),.dinb(w_dff_B_wybVeYra2_1),.dout(n1762));
	jnot g1699(.din(w_n1758_0[0]),.dout(n1763),.clk(gclk));
	jcb g1700(.dina(w_dff_B_d0PaMaEw8_0),.dinb(w_n1725_0[0]),.dout(n1764));
	jand g1701(.dina(n1764),.dinb(w_dff_B_qLp2GrJg0_1),.dout(n1765),.clk(gclk));
	jand g1702(.dina(w_n1755_0[0]),.dinb(w_n1733_0[0]),.dout(n1766),.clk(gclk));
	jand g1703(.dina(w_n1756_0[0]),.dinb(w_n1730_0[0]),.dout(n1767),.clk(gclk));
	jcb g1704(.dina(n1767),.dinb(w_dff_B_6DV67CBU5_1),.dout(n1768));
	jand g1705(.dina(w_G528gat_3[1]),.dinb(w_G205gat_2[1]),.dout(n1769),.clk(gclk));
	jnot g1706(.din(n1769),.dout(n1770),.clk(gclk));
	jand g1707(.dina(w_n1753_0[0]),.dinb(w_n1738_0[0]),.dout(n1771),.clk(gclk));
	jand g1708(.dina(w_n1754_0[0]),.dinb(w_n1735_0[0]),.dout(n1772),.clk(gclk));
	jcb g1709(.dina(n1772),.dinb(w_dff_B_PMZFNPI94_1),.dout(n1773));
	jand g1710(.dina(w_G511gat_3[0]),.dinb(w_G222gat_2[2]),.dout(n1774),.clk(gclk));
	jnot g1711(.din(n1774),.dout(n1775),.clk(gclk));
	jand g1712(.dina(w_n1751_0[0]),.dinb(w_n1743_0[0]),.dout(n1776),.clk(gclk));
	jand g1713(.dina(w_n1752_0[0]),.dinb(w_n1740_0[0]),.dout(n1777),.clk(gclk));
	jcb g1714(.dina(n1777),.dinb(w_dff_B_Rr9uOYLY4_1),.dout(n1778));
	jand g1715(.dina(w_G494gat_2[2]),.dinb(w_G239gat_3[0]),.dout(n1779),.clk(gclk));
	jand g1716(.dina(w_G477gat_2[1]),.dinb(w_G256gat_3[1]),.dout(n1780),.clk(gclk));
	jcb g1717(.dina(w_n1748_0[0]),.dinb(w_n1745_0[0]),.dout(n1781));
	jcb g1718(.dina(w_n1750_0[0]),.dinb(w_n1744_0[0]),.dout(n1782));
	jand g1719(.dina(n1782),.dinb(w_dff_B_i90TR0Ua5_1),.dout(n1783),.clk(gclk));
	jxor g1720(.dina(w_n1783_0[1]),.dinb(w_n1780_0[1]),.dout(n1784),.clk(gclk));
	jnot g1721(.din(n1784),.dout(n1785),.clk(gclk));
	jxor g1722(.dina(w_n1785_0[1]),.dinb(w_n1779_0[1]),.dout(n1786),.clk(gclk));
	jxor g1723(.dina(w_n1786_0[1]),.dinb(w_n1778_0[1]),.dout(n1787),.clk(gclk));
	jxor g1724(.dina(w_n1787_0[1]),.dinb(w_n1775_0[1]),.dout(n1788),.clk(gclk));
	jxor g1725(.dina(w_n1788_0[1]),.dinb(w_n1773_0[1]),.dout(n1789),.clk(gclk));
	jxor g1726(.dina(w_n1789_0[1]),.dinb(w_n1770_0[1]),.dout(n1790),.clk(gclk));
	jxor g1727(.dina(w_n1790_0[1]),.dinb(w_n1768_0[1]),.dout(n1791),.clk(gclk));
	jxor g1728(.dina(w_n1791_0[1]),.dinb(w_n1765_0[1]),.dout(G6260gat),.clk(gclk));
	jnot g1729(.din(w_n1768_0[0]),.dout(n1793),.clk(gclk));
	jnot g1730(.din(w_n1790_0[0]),.dout(n1794),.clk(gclk));
	jcb g1731(.dina(n1794),.dinb(w_dff_B_qnSP67mV0_1),.dout(n1795));
	jnot g1732(.din(w_n1791_0[0]),.dout(n1796),.clk(gclk));
	jcb g1733(.dina(w_dff_B_L95tFTN21_0),.dinb(w_n1765_0[0]),.dout(n1797));
	jand g1734(.dina(n1797),.dinb(w_dff_B_OoUBXaLt3_1),.dout(n1798),.clk(gclk));
	jand g1735(.dina(w_n1788_0[0]),.dinb(w_n1773_0[0]),.dout(n1799),.clk(gclk));
	jand g1736(.dina(w_n1789_0[0]),.dinb(w_n1770_0[0]),.dout(n1800),.clk(gclk));
	jcb g1737(.dina(n1800),.dinb(w_dff_B_BXjl0G2O6_1),.dout(n1801));
	jand g1738(.dina(w_G528gat_3[0]),.dinb(w_G222gat_2[1]),.dout(n1802),.clk(gclk));
	jnot g1739(.din(n1802),.dout(n1803),.clk(gclk));
	jand g1740(.dina(w_n1786_0[0]),.dinb(w_n1778_0[0]),.dout(n1804),.clk(gclk));
	jand g1741(.dina(w_n1787_0[0]),.dinb(w_n1775_0[0]),.dout(n1805),.clk(gclk));
	jcb g1742(.dina(n1805),.dinb(w_dff_B_rylctyCW3_1),.dout(n1806));
	jand g1743(.dina(w_G511gat_2[2]),.dinb(w_G239gat_2[2]),.dout(n1807),.clk(gclk));
	jand g1744(.dina(w_G494gat_2[1]),.dinb(w_G256gat_3[0]),.dout(n1808),.clk(gclk));
	jcb g1745(.dina(w_n1783_0[0]),.dinb(w_n1780_0[0]),.dout(n1809));
	jcb g1746(.dina(w_n1785_0[0]),.dinb(w_n1779_0[0]),.dout(n1810));
	jand g1747(.dina(n1810),.dinb(w_dff_B_phKCi7S75_1),.dout(n1811),.clk(gclk));
	jxor g1748(.dina(w_n1811_0[1]),.dinb(w_n1808_0[1]),.dout(n1812),.clk(gclk));
	jnot g1749(.din(n1812),.dout(n1813),.clk(gclk));
	jxor g1750(.dina(w_n1813_0[1]),.dinb(w_n1807_0[1]),.dout(n1814),.clk(gclk));
	jxor g1751(.dina(w_n1814_0[1]),.dinb(w_n1806_0[1]),.dout(n1815),.clk(gclk));
	jxor g1752(.dina(w_n1815_0[1]),.dinb(w_n1803_0[1]),.dout(n1816),.clk(gclk));
	jxor g1753(.dina(w_n1816_0[1]),.dinb(w_n1801_0[1]),.dout(n1817),.clk(gclk));
	jxor g1754(.dina(w_n1817_0[1]),.dinb(w_n1798_0[1]),.dout(G6270gat),.clk(gclk));
	jnot g1755(.din(w_n1801_0[0]),.dout(n1819),.clk(gclk));
	jnot g1756(.din(w_n1816_0[0]),.dout(n1820),.clk(gclk));
	jcb g1757(.dina(n1820),.dinb(w_dff_B_BIrgQ7AT7_1),.dout(n1821));
	jnot g1758(.din(w_n1817_0[0]),.dout(n1822),.clk(gclk));
	jcb g1759(.dina(w_dff_B_q4rbk8rf0_0),.dinb(w_n1798_0[0]),.dout(n1823));
	jand g1760(.dina(n1823),.dinb(w_dff_B_J9BCiSGh4_1),.dout(n1824),.clk(gclk));
	jand g1761(.dina(w_n1814_0[0]),.dinb(w_n1806_0[0]),.dout(n1825),.clk(gclk));
	jand g1762(.dina(w_n1815_0[0]),.dinb(w_n1803_0[0]),.dout(n1826),.clk(gclk));
	jcb g1763(.dina(n1826),.dinb(w_dff_B_zqUqH8KZ3_1),.dout(n1827));
	jand g1764(.dina(w_G528gat_2[2]),.dinb(w_G239gat_2[1]),.dout(n1828),.clk(gclk));
	jand g1765(.dina(w_G511gat_2[1]),.dinb(w_G256gat_2[2]),.dout(n1829),.clk(gclk));
	jcb g1766(.dina(w_n1811_0[0]),.dinb(w_n1808_0[0]),.dout(n1830));
	jcb g1767(.dina(w_n1813_0[0]),.dinb(w_n1807_0[0]),.dout(n1831));
	jand g1768(.dina(n1831),.dinb(w_dff_B_SGXXBPc45_1),.dout(n1832),.clk(gclk));
	jxor g1769(.dina(w_n1832_0[1]),.dinb(w_n1829_0[1]),.dout(n1833),.clk(gclk));
	jnot g1770(.din(n1833),.dout(n1834),.clk(gclk));
	jxor g1771(.dina(w_n1834_0[1]),.dinb(w_n1828_0[1]),.dout(n1835),.clk(gclk));
	jxor g1772(.dina(w_n1835_0[1]),.dinb(w_n1827_0[1]),.dout(n1836),.clk(gclk));
	jxor g1773(.dina(w_n1836_0[1]),.dinb(w_n1824_0[1]),.dout(G6280gat),.clk(gclk));
	jand g1774(.dina(w_G528gat_2[1]),.dinb(w_G256gat_2[1]),.dout(n1838),.clk(gclk));
	jcb g1775(.dina(w_n1832_0[0]),.dinb(w_n1829_0[0]),.dout(n1839));
	jcb g1776(.dina(w_n1834_0[0]),.dinb(w_n1828_0[0]),.dout(n1840));
	jand g1777(.dina(n1840),.dinb(w_dff_B_yPOGelZU9_1),.dout(n1841),.clk(gclk));
	jcb g1778(.dina(w_n1841_0[1]),.dinb(w_n1838_0[1]),.dout(n1842));
	jnot g1779(.din(w_n1827_0[0]),.dout(n1843),.clk(gclk));
	jnot g1780(.din(w_n1835_0[0]),.dout(n1844),.clk(gclk));
	jcb g1781(.dina(n1844),.dinb(w_dff_B_6dBjoyOm3_1),.dout(n1845));
	jnot g1782(.din(w_n1836_0[0]),.dout(n1846),.clk(gclk));
	jcb g1783(.dina(w_dff_B_bdjq8WZ84_0),.dinb(w_n1824_0[0]),.dout(n1847));
	jand g1784(.dina(n1847),.dinb(w_dff_B_9QfVd1cd8_1),.dout(n1848),.clk(gclk));
	jxor g1785(.dina(w_n1841_0[0]),.dinb(w_n1838_0[0]),.dout(n1849),.clk(gclk));
	jnot g1786(.din(w_n1849_0[1]),.dout(n1850),.clk(gclk));
	jcb g1787(.dina(w_dff_B_Lx61Oscp4_0),.dinb(w_n1848_0[1]),.dout(n1851));
	jand g1788(.dina(n1851),.dinb(w_dff_B_jLMa77NH2_1),.dout(G6287gat),.clk(gclk));
	jxor g1789(.dina(w_n1849_0[0]),.dinb(w_n1848_0[0]),.dout(G6288gat),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_G1gat_0[0]),.doutb(w_G1gat_0[1]),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G1gat_1(.douta(w_G1gat_1[0]),.doutb(w_G1gat_1[1]),.doutc(w_G1gat_1[2]),.din(w_G1gat_0[0]));
	jspl3 jspl3_w_G1gat_2(.douta(w_G1gat_2[0]),.doutb(w_G1gat_2[1]),.doutc(w_G1gat_2[2]),.din(w_G1gat_0[1]));
	jspl3 jspl3_w_G1gat_3(.douta(w_G1gat_3[0]),.doutb(w_G1gat_3[1]),.doutc(w_G1gat_3[2]),.din(w_G1gat_0[2]));
	jspl3 jspl3_w_G1gat_4(.douta(w_G1gat_4[0]),.doutb(w_G1gat_4[1]),.doutc(w_G1gat_4[2]),.din(w_G1gat_1[0]));
	jspl3 jspl3_w_G1gat_5(.douta(w_G1gat_5[0]),.doutb(w_G1gat_5[1]),.doutc(w_G1gat_5[2]),.din(w_G1gat_1[1]));
	jspl3 jspl3_w_G1gat_6(.douta(w_G1gat_6[0]),.doutb(w_G1gat_6[1]),.doutc(w_G1gat_6[2]),.din(w_G1gat_1[2]));
	jspl jspl_w_G1gat_7(.douta(w_G1gat_7[0]),.doutb(w_G1gat_7[1]),.din(w_G1gat_2[0]));
	jspl3 jspl3_w_G18gat_0(.douta(w_G18gat_0[0]),.doutb(w_G18gat_0[1]),.doutc(w_G18gat_0[2]),.din(G18gat));
	jspl3 jspl3_w_G18gat_1(.douta(w_G18gat_1[0]),.doutb(w_G18gat_1[1]),.doutc(w_G18gat_1[2]),.din(w_G18gat_0[0]));
	jspl3 jspl3_w_G18gat_2(.douta(w_G18gat_2[0]),.doutb(w_G18gat_2[1]),.doutc(w_G18gat_2[2]),.din(w_G18gat_0[1]));
	jspl3 jspl3_w_G18gat_3(.douta(w_G18gat_3[0]),.doutb(w_G18gat_3[1]),.doutc(w_G18gat_3[2]),.din(w_G18gat_0[2]));
	jspl3 jspl3_w_G18gat_4(.douta(w_G18gat_4[0]),.doutb(w_G18gat_4[1]),.doutc(w_G18gat_4[2]),.din(w_G18gat_1[0]));
	jspl3 jspl3_w_G18gat_5(.douta(w_G18gat_5[0]),.doutb(w_G18gat_5[1]),.doutc(w_G18gat_5[2]),.din(w_G18gat_1[1]));
	jspl3 jspl3_w_G18gat_6(.douta(w_G18gat_6[0]),.doutb(w_G18gat_6[1]),.doutc(w_G18gat_6[2]),.din(w_G18gat_1[2]));
	jspl3 jspl3_w_G18gat_7(.douta(w_G18gat_7[0]),.doutb(w_G18gat_7[1]),.doutc(w_G18gat_7[2]),.din(w_G18gat_2[0]));
	jspl3 jspl3_w_G35gat_0(.douta(w_G35gat_0[0]),.doutb(w_G35gat_0[1]),.doutc(w_G35gat_0[2]),.din(G35gat));
	jspl3 jspl3_w_G35gat_1(.douta(w_G35gat_1[0]),.doutb(w_G35gat_1[1]),.doutc(w_G35gat_1[2]),.din(w_G35gat_0[0]));
	jspl3 jspl3_w_G35gat_2(.douta(w_G35gat_2[0]),.doutb(w_G35gat_2[1]),.doutc(w_G35gat_2[2]),.din(w_G35gat_0[1]));
	jspl3 jspl3_w_G35gat_3(.douta(w_G35gat_3[0]),.doutb(w_G35gat_3[1]),.doutc(w_G35gat_3[2]),.din(w_G35gat_0[2]));
	jspl3 jspl3_w_G35gat_4(.douta(w_G35gat_4[0]),.doutb(w_G35gat_4[1]),.doutc(w_G35gat_4[2]),.din(w_G35gat_1[0]));
	jspl3 jspl3_w_G35gat_5(.douta(w_G35gat_5[0]),.doutb(w_G35gat_5[1]),.doutc(w_G35gat_5[2]),.din(w_G35gat_1[1]));
	jspl3 jspl3_w_G35gat_6(.douta(w_G35gat_6[0]),.doutb(w_G35gat_6[1]),.doutc(w_G35gat_6[2]),.din(w_G35gat_1[2]));
	jspl3 jspl3_w_G35gat_7(.douta(w_G35gat_7[0]),.doutb(w_G35gat_7[1]),.doutc(w_G35gat_7[2]),.din(w_G35gat_2[0]));
	jspl3 jspl3_w_G52gat_0(.douta(w_G52gat_0[0]),.doutb(w_G52gat_0[1]),.doutc(w_G52gat_0[2]),.din(G52gat));
	jspl3 jspl3_w_G52gat_1(.douta(w_G52gat_1[0]),.doutb(w_G52gat_1[1]),.doutc(w_G52gat_1[2]),.din(w_G52gat_0[0]));
	jspl3 jspl3_w_G52gat_2(.douta(w_G52gat_2[0]),.doutb(w_G52gat_2[1]),.doutc(w_G52gat_2[2]),.din(w_G52gat_0[1]));
	jspl3 jspl3_w_G52gat_3(.douta(w_G52gat_3[0]),.doutb(w_G52gat_3[1]),.doutc(w_G52gat_3[2]),.din(w_G52gat_0[2]));
	jspl3 jspl3_w_G52gat_4(.douta(w_G52gat_4[0]),.doutb(w_G52gat_4[1]),.doutc(w_G52gat_4[2]),.din(w_G52gat_1[0]));
	jspl3 jspl3_w_G52gat_5(.douta(w_G52gat_5[0]),.doutb(w_G52gat_5[1]),.doutc(w_G52gat_5[2]),.din(w_G52gat_1[1]));
	jspl3 jspl3_w_G52gat_6(.douta(w_G52gat_6[0]),.doutb(w_G52gat_6[1]),.doutc(w_G52gat_6[2]),.din(w_G52gat_1[2]));
	jspl3 jspl3_w_G52gat_7(.douta(w_G52gat_7[0]),.doutb(w_G52gat_7[1]),.doutc(w_G52gat_7[2]),.din(w_G52gat_2[0]));
	jspl3 jspl3_w_G69gat_0(.douta(w_G69gat_0[0]),.doutb(w_G69gat_0[1]),.doutc(w_G69gat_0[2]),.din(G69gat));
	jspl3 jspl3_w_G69gat_1(.douta(w_G69gat_1[0]),.doutb(w_G69gat_1[1]),.doutc(w_G69gat_1[2]),.din(w_G69gat_0[0]));
	jspl3 jspl3_w_G69gat_2(.douta(w_G69gat_2[0]),.doutb(w_G69gat_2[1]),.doutc(w_G69gat_2[2]),.din(w_G69gat_0[1]));
	jspl3 jspl3_w_G69gat_3(.douta(w_G69gat_3[0]),.doutb(w_G69gat_3[1]),.doutc(w_G69gat_3[2]),.din(w_G69gat_0[2]));
	jspl3 jspl3_w_G69gat_4(.douta(w_G69gat_4[0]),.doutb(w_G69gat_4[1]),.doutc(w_G69gat_4[2]),.din(w_G69gat_1[0]));
	jspl3 jspl3_w_G69gat_5(.douta(w_G69gat_5[0]),.doutb(w_G69gat_5[1]),.doutc(w_G69gat_5[2]),.din(w_G69gat_1[1]));
	jspl3 jspl3_w_G69gat_6(.douta(w_G69gat_6[0]),.doutb(w_G69gat_6[1]),.doutc(w_G69gat_6[2]),.din(w_G69gat_1[2]));
	jspl jspl_w_G69gat_7(.douta(w_G69gat_7[0]),.doutb(w_G69gat_7[1]),.din(w_G69gat_2[0]));
	jspl3 jspl3_w_G86gat_0(.douta(w_G86gat_0[0]),.doutb(w_G86gat_0[1]),.doutc(w_G86gat_0[2]),.din(G86gat));
	jspl3 jspl3_w_G86gat_1(.douta(w_G86gat_1[0]),.doutb(w_G86gat_1[1]),.doutc(w_G86gat_1[2]),.din(w_G86gat_0[0]));
	jspl3 jspl3_w_G86gat_2(.douta(w_G86gat_2[0]),.doutb(w_G86gat_2[1]),.doutc(w_G86gat_2[2]),.din(w_G86gat_0[1]));
	jspl3 jspl3_w_G86gat_3(.douta(w_G86gat_3[0]),.doutb(w_G86gat_3[1]),.doutc(w_G86gat_3[2]),.din(w_G86gat_0[2]));
	jspl3 jspl3_w_G86gat_4(.douta(w_G86gat_4[0]),.doutb(w_G86gat_4[1]),.doutc(w_G86gat_4[2]),.din(w_G86gat_1[0]));
	jspl3 jspl3_w_G86gat_5(.douta(w_G86gat_5[0]),.doutb(w_G86gat_5[1]),.doutc(w_G86gat_5[2]),.din(w_G86gat_1[1]));
	jspl3 jspl3_w_G86gat_6(.douta(w_G86gat_6[0]),.doutb(w_G86gat_6[1]),.doutc(w_G86gat_6[2]),.din(w_G86gat_1[2]));
	jspl jspl_w_G86gat_7(.douta(w_G86gat_7[0]),.doutb(w_G86gat_7[1]),.din(w_G86gat_2[0]));
	jspl3 jspl3_w_G103gat_0(.douta(w_G103gat_0[0]),.doutb(w_G103gat_0[1]),.doutc(w_G103gat_0[2]),.din(G103gat));
	jspl3 jspl3_w_G103gat_1(.douta(w_G103gat_1[0]),.doutb(w_G103gat_1[1]),.doutc(w_G103gat_1[2]),.din(w_G103gat_0[0]));
	jspl3 jspl3_w_G103gat_2(.douta(w_G103gat_2[0]),.doutb(w_G103gat_2[1]),.doutc(w_G103gat_2[2]),.din(w_G103gat_0[1]));
	jspl3 jspl3_w_G103gat_3(.douta(w_G103gat_3[0]),.doutb(w_G103gat_3[1]),.doutc(w_G103gat_3[2]),.din(w_G103gat_0[2]));
	jspl3 jspl3_w_G103gat_4(.douta(w_G103gat_4[0]),.doutb(w_G103gat_4[1]),.doutc(w_G103gat_4[2]),.din(w_G103gat_1[0]));
	jspl3 jspl3_w_G103gat_5(.douta(w_G103gat_5[0]),.doutb(w_G103gat_5[1]),.doutc(w_G103gat_5[2]),.din(w_G103gat_1[1]));
	jspl3 jspl3_w_G103gat_6(.douta(w_G103gat_6[0]),.doutb(w_G103gat_6[1]),.doutc(w_G103gat_6[2]),.din(w_G103gat_1[2]));
	jspl jspl_w_G103gat_7(.douta(w_G103gat_7[0]),.doutb(w_G103gat_7[1]),.din(w_G103gat_2[0]));
	jspl3 jspl3_w_G120gat_0(.douta(w_G120gat_0[0]),.doutb(w_G120gat_0[1]),.doutc(w_G120gat_0[2]),.din(G120gat));
	jspl3 jspl3_w_G120gat_1(.douta(w_G120gat_1[0]),.doutb(w_G120gat_1[1]),.doutc(w_G120gat_1[2]),.din(w_G120gat_0[0]));
	jspl3 jspl3_w_G120gat_2(.douta(w_G120gat_2[0]),.doutb(w_G120gat_2[1]),.doutc(w_G120gat_2[2]),.din(w_G120gat_0[1]));
	jspl3 jspl3_w_G120gat_3(.douta(w_G120gat_3[0]),.doutb(w_G120gat_3[1]),.doutc(w_G120gat_3[2]),.din(w_G120gat_0[2]));
	jspl3 jspl3_w_G120gat_4(.douta(w_G120gat_4[0]),.doutb(w_G120gat_4[1]),.doutc(w_G120gat_4[2]),.din(w_G120gat_1[0]));
	jspl3 jspl3_w_G120gat_5(.douta(w_G120gat_5[0]),.doutb(w_G120gat_5[1]),.doutc(w_G120gat_5[2]),.din(w_G120gat_1[1]));
	jspl3 jspl3_w_G120gat_6(.douta(w_G120gat_6[0]),.doutb(w_G120gat_6[1]),.doutc(w_G120gat_6[2]),.din(w_G120gat_1[2]));
	jspl jspl_w_G120gat_7(.douta(w_G120gat_7[0]),.doutb(w_G120gat_7[1]),.din(w_G120gat_2[0]));
	jspl3 jspl3_w_G137gat_0(.douta(w_G137gat_0[0]),.doutb(w_G137gat_0[1]),.doutc(w_G137gat_0[2]),.din(G137gat));
	jspl3 jspl3_w_G137gat_1(.douta(w_G137gat_1[0]),.doutb(w_G137gat_1[1]),.doutc(w_G137gat_1[2]),.din(w_G137gat_0[0]));
	jspl3 jspl3_w_G137gat_2(.douta(w_G137gat_2[0]),.doutb(w_G137gat_2[1]),.doutc(w_G137gat_2[2]),.din(w_G137gat_0[1]));
	jspl3 jspl3_w_G137gat_3(.douta(w_G137gat_3[0]),.doutb(w_G137gat_3[1]),.doutc(w_G137gat_3[2]),.din(w_G137gat_0[2]));
	jspl3 jspl3_w_G137gat_4(.douta(w_G137gat_4[0]),.doutb(w_G137gat_4[1]),.doutc(w_G137gat_4[2]),.din(w_G137gat_1[0]));
	jspl3 jspl3_w_G137gat_5(.douta(w_G137gat_5[0]),.doutb(w_G137gat_5[1]),.doutc(w_G137gat_5[2]),.din(w_G137gat_1[1]));
	jspl3 jspl3_w_G137gat_6(.douta(w_G137gat_6[0]),.doutb(w_G137gat_6[1]),.doutc(w_G137gat_6[2]),.din(w_G137gat_1[2]));
	jspl jspl_w_G137gat_7(.douta(w_G137gat_7[0]),.doutb(w_G137gat_7[1]),.din(w_G137gat_2[0]));
	jspl3 jspl3_w_G154gat_0(.douta(w_G154gat_0[0]),.doutb(w_G154gat_0[1]),.doutc(w_G154gat_0[2]),.din(G154gat));
	jspl3 jspl3_w_G154gat_1(.douta(w_G154gat_1[0]),.doutb(w_G154gat_1[1]),.doutc(w_G154gat_1[2]),.din(w_G154gat_0[0]));
	jspl3 jspl3_w_G154gat_2(.douta(w_G154gat_2[0]),.doutb(w_G154gat_2[1]),.doutc(w_G154gat_2[2]),.din(w_G154gat_0[1]));
	jspl3 jspl3_w_G154gat_3(.douta(w_G154gat_3[0]),.doutb(w_G154gat_3[1]),.doutc(w_G154gat_3[2]),.din(w_G154gat_0[2]));
	jspl3 jspl3_w_G154gat_4(.douta(w_G154gat_4[0]),.doutb(w_G154gat_4[1]),.doutc(w_G154gat_4[2]),.din(w_G154gat_1[0]));
	jspl3 jspl3_w_G154gat_5(.douta(w_G154gat_5[0]),.doutb(w_G154gat_5[1]),.doutc(w_G154gat_5[2]),.din(w_G154gat_1[1]));
	jspl3 jspl3_w_G154gat_6(.douta(w_G154gat_6[0]),.doutb(w_G154gat_6[1]),.doutc(w_G154gat_6[2]),.din(w_G154gat_1[2]));
	jspl jspl_w_G154gat_7(.douta(w_G154gat_7[0]),.doutb(w_G154gat_7[1]),.din(w_G154gat_2[0]));
	jspl3 jspl3_w_G171gat_0(.douta(w_G171gat_0[0]),.doutb(w_G171gat_0[1]),.doutc(w_G171gat_0[2]),.din(G171gat));
	jspl3 jspl3_w_G171gat_1(.douta(w_G171gat_1[0]),.doutb(w_G171gat_1[1]),.doutc(w_G171gat_1[2]),.din(w_G171gat_0[0]));
	jspl3 jspl3_w_G171gat_2(.douta(w_G171gat_2[0]),.doutb(w_G171gat_2[1]),.doutc(w_G171gat_2[2]),.din(w_G171gat_0[1]));
	jspl3 jspl3_w_G171gat_3(.douta(w_G171gat_3[0]),.doutb(w_G171gat_3[1]),.doutc(w_G171gat_3[2]),.din(w_G171gat_0[2]));
	jspl3 jspl3_w_G171gat_4(.douta(w_G171gat_4[0]),.doutb(w_G171gat_4[1]),.doutc(w_G171gat_4[2]),.din(w_G171gat_1[0]));
	jspl3 jspl3_w_G171gat_5(.douta(w_G171gat_5[0]),.doutb(w_G171gat_5[1]),.doutc(w_G171gat_5[2]),.din(w_G171gat_1[1]));
	jspl3 jspl3_w_G171gat_6(.douta(w_G171gat_6[0]),.doutb(w_G171gat_6[1]),.doutc(w_G171gat_6[2]),.din(w_G171gat_1[2]));
	jspl jspl_w_G171gat_7(.douta(w_G171gat_7[0]),.doutb(w_G171gat_7[1]),.din(w_G171gat_2[0]));
	jspl3 jspl3_w_G188gat_0(.douta(w_G188gat_0[0]),.doutb(w_G188gat_0[1]),.doutc(w_G188gat_0[2]),.din(G188gat));
	jspl3 jspl3_w_G188gat_1(.douta(w_G188gat_1[0]),.doutb(w_G188gat_1[1]),.doutc(w_G188gat_1[2]),.din(w_G188gat_0[0]));
	jspl3 jspl3_w_G188gat_2(.douta(w_G188gat_2[0]),.doutb(w_G188gat_2[1]),.doutc(w_G188gat_2[2]),.din(w_G188gat_0[1]));
	jspl3 jspl3_w_G188gat_3(.douta(w_G188gat_3[0]),.doutb(w_G188gat_3[1]),.doutc(w_G188gat_3[2]),.din(w_G188gat_0[2]));
	jspl3 jspl3_w_G188gat_4(.douta(w_G188gat_4[0]),.doutb(w_G188gat_4[1]),.doutc(w_G188gat_4[2]),.din(w_G188gat_1[0]));
	jspl3 jspl3_w_G188gat_5(.douta(w_G188gat_5[0]),.doutb(w_G188gat_5[1]),.doutc(w_G188gat_5[2]),.din(w_G188gat_1[1]));
	jspl3 jspl3_w_G188gat_6(.douta(w_G188gat_6[0]),.doutb(w_G188gat_6[1]),.doutc(w_G188gat_6[2]),.din(w_G188gat_1[2]));
	jspl jspl_w_G188gat_7(.douta(w_G188gat_7[0]),.doutb(w_G188gat_7[1]),.din(w_G188gat_2[0]));
	jspl3 jspl3_w_G205gat_0(.douta(w_G205gat_0[0]),.doutb(w_G205gat_0[1]),.doutc(w_G205gat_0[2]),.din(G205gat));
	jspl3 jspl3_w_G205gat_1(.douta(w_G205gat_1[0]),.doutb(w_G205gat_1[1]),.doutc(w_G205gat_1[2]),.din(w_G205gat_0[0]));
	jspl3 jspl3_w_G205gat_2(.douta(w_G205gat_2[0]),.doutb(w_G205gat_2[1]),.doutc(w_G205gat_2[2]),.din(w_G205gat_0[1]));
	jspl3 jspl3_w_G205gat_3(.douta(w_G205gat_3[0]),.doutb(w_G205gat_3[1]),.doutc(w_G205gat_3[2]),.din(w_G205gat_0[2]));
	jspl3 jspl3_w_G205gat_4(.douta(w_G205gat_4[0]),.doutb(w_G205gat_4[1]),.doutc(w_G205gat_4[2]),.din(w_G205gat_1[0]));
	jspl3 jspl3_w_G205gat_5(.douta(w_G205gat_5[0]),.doutb(w_G205gat_5[1]),.doutc(w_G205gat_5[2]),.din(w_G205gat_1[1]));
	jspl3 jspl3_w_G205gat_6(.douta(w_G205gat_6[0]),.doutb(w_G205gat_6[1]),.doutc(w_G205gat_6[2]),.din(w_G205gat_1[2]));
	jspl jspl_w_G205gat_7(.douta(w_G205gat_7[0]),.doutb(w_G205gat_7[1]),.din(w_G205gat_2[0]));
	jspl3 jspl3_w_G222gat_0(.douta(w_G222gat_0[0]),.doutb(w_G222gat_0[1]),.doutc(w_G222gat_0[2]),.din(G222gat));
	jspl3 jspl3_w_G222gat_1(.douta(w_G222gat_1[0]),.doutb(w_G222gat_1[1]),.doutc(w_G222gat_1[2]),.din(w_G222gat_0[0]));
	jspl3 jspl3_w_G222gat_2(.douta(w_G222gat_2[0]),.doutb(w_G222gat_2[1]),.doutc(w_G222gat_2[2]),.din(w_G222gat_0[1]));
	jspl3 jspl3_w_G222gat_3(.douta(w_G222gat_3[0]),.doutb(w_G222gat_3[1]),.doutc(w_G222gat_3[2]),.din(w_G222gat_0[2]));
	jspl3 jspl3_w_G222gat_4(.douta(w_G222gat_4[0]),.doutb(w_G222gat_4[1]),.doutc(w_G222gat_4[2]),.din(w_G222gat_1[0]));
	jspl3 jspl3_w_G222gat_5(.douta(w_G222gat_5[0]),.doutb(w_G222gat_5[1]),.doutc(w_G222gat_5[2]),.din(w_G222gat_1[1]));
	jspl3 jspl3_w_G222gat_6(.douta(w_G222gat_6[0]),.doutb(w_G222gat_6[1]),.doutc(w_G222gat_6[2]),.din(w_G222gat_1[2]));
	jspl jspl_w_G222gat_7(.douta(w_G222gat_7[0]),.doutb(w_G222gat_7[1]),.din(w_G222gat_2[0]));
	jspl3 jspl3_w_G239gat_0(.douta(w_G239gat_0[0]),.doutb(w_G239gat_0[1]),.doutc(w_G239gat_0[2]),.din(G239gat));
	jspl3 jspl3_w_G239gat_1(.douta(w_G239gat_1[0]),.doutb(w_G239gat_1[1]),.doutc(w_G239gat_1[2]),.din(w_G239gat_0[0]));
	jspl3 jspl3_w_G239gat_2(.douta(w_G239gat_2[0]),.doutb(w_G239gat_2[1]),.doutc(w_G239gat_2[2]),.din(w_G239gat_0[1]));
	jspl3 jspl3_w_G239gat_3(.douta(w_G239gat_3[0]),.doutb(w_G239gat_3[1]),.doutc(w_G239gat_3[2]),.din(w_G239gat_0[2]));
	jspl3 jspl3_w_G239gat_4(.douta(w_G239gat_4[0]),.doutb(w_G239gat_4[1]),.doutc(w_G239gat_4[2]),.din(w_G239gat_1[0]));
	jspl3 jspl3_w_G239gat_5(.douta(w_G239gat_5[0]),.doutb(w_G239gat_5[1]),.doutc(w_G239gat_5[2]),.din(w_G239gat_1[1]));
	jspl3 jspl3_w_G239gat_6(.douta(w_G239gat_6[0]),.doutb(w_G239gat_6[1]),.doutc(w_G239gat_6[2]),.din(w_G239gat_1[2]));
	jspl jspl_w_G239gat_7(.douta(w_G239gat_7[0]),.doutb(w_G239gat_7[1]),.din(w_G239gat_2[0]));
	jspl3 jspl3_w_G256gat_0(.douta(w_G256gat_0[0]),.doutb(w_G256gat_0[1]),.doutc(w_G256gat_0[2]),.din(G256gat));
	jspl3 jspl3_w_G256gat_1(.douta(w_G256gat_1[0]),.doutb(w_G256gat_1[1]),.doutc(w_G256gat_1[2]),.din(w_G256gat_0[0]));
	jspl3 jspl3_w_G256gat_2(.douta(w_G256gat_2[0]),.doutb(w_G256gat_2[1]),.doutc(w_G256gat_2[2]),.din(w_G256gat_0[1]));
	jspl3 jspl3_w_G256gat_3(.douta(w_G256gat_3[0]),.doutb(w_G256gat_3[1]),.doutc(w_G256gat_3[2]),.din(w_G256gat_0[2]));
	jspl3 jspl3_w_G256gat_4(.douta(w_G256gat_4[0]),.doutb(w_G256gat_4[1]),.doutc(w_G256gat_4[2]),.din(w_G256gat_1[0]));
	jspl3 jspl3_w_G256gat_5(.douta(w_G256gat_5[0]),.doutb(w_G256gat_5[1]),.doutc(w_G256gat_5[2]),.din(w_G256gat_1[1]));
	jspl3 jspl3_w_G256gat_6(.douta(w_G256gat_6[0]),.doutb(w_G256gat_6[1]),.doutc(w_G256gat_6[2]),.din(w_G256gat_1[2]));
	jspl jspl_w_G256gat_7(.douta(w_G256gat_7[0]),.doutb(w_G256gat_7[1]),.din(w_G256gat_2[0]));
	jspl3 jspl3_w_G273gat_0(.douta(w_G273gat_0[0]),.doutb(w_G273gat_0[1]),.doutc(w_G273gat_0[2]),.din(G273gat));
	jspl3 jspl3_w_G273gat_1(.douta(w_G273gat_1[0]),.doutb(w_G273gat_1[1]),.doutc(w_G273gat_1[2]),.din(w_G273gat_0[0]));
	jspl3 jspl3_w_G273gat_2(.douta(w_G273gat_2[0]),.doutb(w_G273gat_2[1]),.doutc(w_G273gat_2[2]),.din(w_G273gat_0[1]));
	jspl3 jspl3_w_G273gat_3(.douta(w_G273gat_3[0]),.doutb(w_G273gat_3[1]),.doutc(w_G273gat_3[2]),.din(w_G273gat_0[2]));
	jspl3 jspl3_w_G273gat_4(.douta(w_G273gat_4[0]),.doutb(w_G273gat_4[1]),.doutc(w_G273gat_4[2]),.din(w_G273gat_1[0]));
	jspl3 jspl3_w_G273gat_5(.douta(w_G273gat_5[0]),.doutb(w_G273gat_5[1]),.doutc(w_G273gat_5[2]),.din(w_G273gat_1[1]));
	jspl3 jspl3_w_G273gat_6(.douta(w_G273gat_6[0]),.doutb(w_G273gat_6[1]),.doutc(w_G273gat_6[2]),.din(w_G273gat_1[2]));
	jspl3 jspl3_w_G273gat_7(.douta(w_G273gat_7[0]),.doutb(w_G273gat_7[1]),.doutc(w_G273gat_7[2]),.din(w_G273gat_2[0]));
	jspl3 jspl3_w_G290gat_0(.douta(w_G290gat_0[0]),.doutb(w_G290gat_0[1]),.doutc(w_G290gat_0[2]),.din(G290gat));
	jspl3 jspl3_w_G290gat_1(.douta(w_G290gat_1[0]),.doutb(w_G290gat_1[1]),.doutc(w_G290gat_1[2]),.din(w_G290gat_0[0]));
	jspl3 jspl3_w_G290gat_2(.douta(w_G290gat_2[0]),.doutb(w_G290gat_2[1]),.doutc(w_G290gat_2[2]),.din(w_G290gat_0[1]));
	jspl3 jspl3_w_G290gat_3(.douta(w_G290gat_3[0]),.doutb(w_G290gat_3[1]),.doutc(w_G290gat_3[2]),.din(w_G290gat_0[2]));
	jspl3 jspl3_w_G290gat_4(.douta(w_G290gat_4[0]),.doutb(w_G290gat_4[1]),.doutc(w_G290gat_4[2]),.din(w_G290gat_1[0]));
	jspl3 jspl3_w_G290gat_5(.douta(w_G290gat_5[0]),.doutb(w_G290gat_5[1]),.doutc(w_G290gat_5[2]),.din(w_G290gat_1[1]));
	jspl3 jspl3_w_G290gat_6(.douta(w_G290gat_6[0]),.doutb(w_G290gat_6[1]),.doutc(w_G290gat_6[2]),.din(w_G290gat_1[2]));
	jspl3 jspl3_w_G290gat_7(.douta(w_G290gat_7[0]),.doutb(w_G290gat_7[1]),.doutc(w_G290gat_7[2]),.din(w_G290gat_2[0]));
	jspl3 jspl3_w_G307gat_0(.douta(w_G307gat_0[0]),.doutb(w_G307gat_0[1]),.doutc(w_G307gat_0[2]),.din(G307gat));
	jspl3 jspl3_w_G307gat_1(.douta(w_G307gat_1[0]),.doutb(w_G307gat_1[1]),.doutc(w_G307gat_1[2]),.din(w_G307gat_0[0]));
	jspl3 jspl3_w_G307gat_2(.douta(w_G307gat_2[0]),.doutb(w_dff_A_D8rU4KIX2_1),.doutc(w_G307gat_2[2]),.din(w_G307gat_0[1]));
	jspl3 jspl3_w_G307gat_3(.douta(w_G307gat_3[0]),.doutb(w_G307gat_3[1]),.doutc(w_G307gat_3[2]),.din(w_G307gat_0[2]));
	jspl3 jspl3_w_G307gat_4(.douta(w_G307gat_4[0]),.doutb(w_G307gat_4[1]),.doutc(w_G307gat_4[2]),.din(w_G307gat_1[0]));
	jspl3 jspl3_w_G307gat_5(.douta(w_G307gat_5[0]),.doutb(w_G307gat_5[1]),.doutc(w_G307gat_5[2]),.din(w_G307gat_1[1]));
	jspl3 jspl3_w_G307gat_6(.douta(w_G307gat_6[0]),.doutb(w_G307gat_6[1]),.doutc(w_G307gat_6[2]),.din(w_G307gat_1[2]));
	jspl3 jspl3_w_G307gat_7(.douta(w_G307gat_7[0]),.doutb(w_G307gat_7[1]),.doutc(w_G307gat_7[2]),.din(w_G307gat_2[0]));
	jspl3 jspl3_w_G324gat_0(.douta(w_G324gat_0[0]),.doutb(w_G324gat_0[1]),.doutc(w_G324gat_0[2]),.din(G324gat));
	jspl3 jspl3_w_G324gat_1(.douta(w_G324gat_1[0]),.doutb(w_G324gat_1[1]),.doutc(w_G324gat_1[2]),.din(w_G324gat_0[0]));
	jspl3 jspl3_w_G324gat_2(.douta(w_G324gat_2[0]),.doutb(w_G324gat_2[1]),.doutc(w_G324gat_2[2]),.din(w_G324gat_0[1]));
	jspl3 jspl3_w_G324gat_3(.douta(w_G324gat_3[0]),.doutb(w_G324gat_3[1]),.doutc(w_G324gat_3[2]),.din(w_G324gat_0[2]));
	jspl3 jspl3_w_G324gat_4(.douta(w_G324gat_4[0]),.doutb(w_G324gat_4[1]),.doutc(w_G324gat_4[2]),.din(w_G324gat_1[0]));
	jspl3 jspl3_w_G324gat_5(.douta(w_G324gat_5[0]),.doutb(w_G324gat_5[1]),.doutc(w_G324gat_5[2]),.din(w_G324gat_1[1]));
	jspl3 jspl3_w_G324gat_6(.douta(w_G324gat_6[0]),.doutb(w_G324gat_6[1]),.doutc(w_G324gat_6[2]),.din(w_G324gat_1[2]));
	jspl jspl_w_G324gat_7(.douta(w_G324gat_7[0]),.doutb(w_G324gat_7[1]),.din(w_G324gat_2[0]));
	jspl3 jspl3_w_G341gat_0(.douta(w_G341gat_0[0]),.doutb(w_G341gat_0[1]),.doutc(w_G341gat_0[2]),.din(G341gat));
	jspl3 jspl3_w_G341gat_1(.douta(w_G341gat_1[0]),.doutb(w_G341gat_1[1]),.doutc(w_G341gat_1[2]),.din(w_G341gat_0[0]));
	jspl3 jspl3_w_G341gat_2(.douta(w_G341gat_2[0]),.doutb(w_G341gat_2[1]),.doutc(w_G341gat_2[2]),.din(w_G341gat_0[1]));
	jspl3 jspl3_w_G341gat_3(.douta(w_G341gat_3[0]),.doutb(w_G341gat_3[1]),.doutc(w_G341gat_3[2]),.din(w_G341gat_0[2]));
	jspl3 jspl3_w_G341gat_4(.douta(w_G341gat_4[0]),.doutb(w_G341gat_4[1]),.doutc(w_G341gat_4[2]),.din(w_G341gat_1[0]));
	jspl3 jspl3_w_G341gat_5(.douta(w_G341gat_5[0]),.doutb(w_G341gat_5[1]),.doutc(w_G341gat_5[2]),.din(w_G341gat_1[1]));
	jspl3 jspl3_w_G341gat_6(.douta(w_G341gat_6[0]),.doutb(w_G341gat_6[1]),.doutc(w_G341gat_6[2]),.din(w_G341gat_1[2]));
	jspl jspl_w_G341gat_7(.douta(w_G341gat_7[0]),.doutb(w_G341gat_7[1]),.din(w_G341gat_2[0]));
	jspl3 jspl3_w_G358gat_0(.douta(w_G358gat_0[0]),.doutb(w_G358gat_0[1]),.doutc(w_G358gat_0[2]),.din(G358gat));
	jspl3 jspl3_w_G358gat_1(.douta(w_G358gat_1[0]),.doutb(w_G358gat_1[1]),.doutc(w_G358gat_1[2]),.din(w_G358gat_0[0]));
	jspl3 jspl3_w_G358gat_2(.douta(w_G358gat_2[0]),.doutb(w_G358gat_2[1]),.doutc(w_G358gat_2[2]),.din(w_G358gat_0[1]));
	jspl3 jspl3_w_G358gat_3(.douta(w_G358gat_3[0]),.doutb(w_G358gat_3[1]),.doutc(w_G358gat_3[2]),.din(w_G358gat_0[2]));
	jspl3 jspl3_w_G358gat_4(.douta(w_G358gat_4[0]),.doutb(w_G358gat_4[1]),.doutc(w_G358gat_4[2]),.din(w_G358gat_1[0]));
	jspl3 jspl3_w_G358gat_5(.douta(w_G358gat_5[0]),.doutb(w_G358gat_5[1]),.doutc(w_G358gat_5[2]),.din(w_G358gat_1[1]));
	jspl3 jspl3_w_G358gat_6(.douta(w_G358gat_6[0]),.doutb(w_G358gat_6[1]),.doutc(w_G358gat_6[2]),.din(w_G358gat_1[2]));
	jspl jspl_w_G358gat_7(.douta(w_G358gat_7[0]),.doutb(w_G358gat_7[1]),.din(w_G358gat_2[0]));
	jspl3 jspl3_w_G375gat_0(.douta(w_G375gat_0[0]),.doutb(w_G375gat_0[1]),.doutc(w_G375gat_0[2]),.din(G375gat));
	jspl3 jspl3_w_G375gat_1(.douta(w_G375gat_1[0]),.doutb(w_G375gat_1[1]),.doutc(w_G375gat_1[2]),.din(w_G375gat_0[0]));
	jspl3 jspl3_w_G375gat_2(.douta(w_G375gat_2[0]),.doutb(w_G375gat_2[1]),.doutc(w_G375gat_2[2]),.din(w_G375gat_0[1]));
	jspl3 jspl3_w_G375gat_3(.douta(w_G375gat_3[0]),.doutb(w_G375gat_3[1]),.doutc(w_G375gat_3[2]),.din(w_G375gat_0[2]));
	jspl3 jspl3_w_G375gat_4(.douta(w_G375gat_4[0]),.doutb(w_G375gat_4[1]),.doutc(w_G375gat_4[2]),.din(w_G375gat_1[0]));
	jspl3 jspl3_w_G375gat_5(.douta(w_G375gat_5[0]),.doutb(w_G375gat_5[1]),.doutc(w_G375gat_5[2]),.din(w_G375gat_1[1]));
	jspl3 jspl3_w_G375gat_6(.douta(w_G375gat_6[0]),.doutb(w_G375gat_6[1]),.doutc(w_G375gat_6[2]),.din(w_G375gat_1[2]));
	jspl jspl_w_G375gat_7(.douta(w_G375gat_7[0]),.doutb(w_G375gat_7[1]),.din(w_G375gat_2[0]));
	jspl3 jspl3_w_G392gat_0(.douta(w_G392gat_0[0]),.doutb(w_G392gat_0[1]),.doutc(w_G392gat_0[2]),.din(G392gat));
	jspl3 jspl3_w_G392gat_1(.douta(w_G392gat_1[0]),.doutb(w_G392gat_1[1]),.doutc(w_G392gat_1[2]),.din(w_G392gat_0[0]));
	jspl3 jspl3_w_G392gat_2(.douta(w_G392gat_2[0]),.doutb(w_G392gat_2[1]),.doutc(w_G392gat_2[2]),.din(w_G392gat_0[1]));
	jspl3 jspl3_w_G392gat_3(.douta(w_G392gat_3[0]),.doutb(w_G392gat_3[1]),.doutc(w_G392gat_3[2]),.din(w_G392gat_0[2]));
	jspl3 jspl3_w_G392gat_4(.douta(w_G392gat_4[0]),.doutb(w_G392gat_4[1]),.doutc(w_G392gat_4[2]),.din(w_G392gat_1[0]));
	jspl3 jspl3_w_G392gat_5(.douta(w_G392gat_5[0]),.doutb(w_G392gat_5[1]),.doutc(w_G392gat_5[2]),.din(w_G392gat_1[1]));
	jspl3 jspl3_w_G392gat_6(.douta(w_G392gat_6[0]),.doutb(w_G392gat_6[1]),.doutc(w_G392gat_6[2]),.din(w_G392gat_1[2]));
	jspl jspl_w_G392gat_7(.douta(w_G392gat_7[0]),.doutb(w_G392gat_7[1]),.din(w_G392gat_2[0]));
	jspl3 jspl3_w_G409gat_0(.douta(w_G409gat_0[0]),.doutb(w_G409gat_0[1]),.doutc(w_G409gat_0[2]),.din(G409gat));
	jspl3 jspl3_w_G409gat_1(.douta(w_G409gat_1[0]),.doutb(w_G409gat_1[1]),.doutc(w_G409gat_1[2]),.din(w_G409gat_0[0]));
	jspl3 jspl3_w_G409gat_2(.douta(w_G409gat_2[0]),.doutb(w_G409gat_2[1]),.doutc(w_G409gat_2[2]),.din(w_G409gat_0[1]));
	jspl3 jspl3_w_G409gat_3(.douta(w_G409gat_3[0]),.doutb(w_G409gat_3[1]),.doutc(w_G409gat_3[2]),.din(w_G409gat_0[2]));
	jspl3 jspl3_w_G409gat_4(.douta(w_G409gat_4[0]),.doutb(w_G409gat_4[1]),.doutc(w_G409gat_4[2]),.din(w_G409gat_1[0]));
	jspl3 jspl3_w_G409gat_5(.douta(w_G409gat_5[0]),.doutb(w_G409gat_5[1]),.doutc(w_G409gat_5[2]),.din(w_G409gat_1[1]));
	jspl3 jspl3_w_G409gat_6(.douta(w_G409gat_6[0]),.doutb(w_G409gat_6[1]),.doutc(w_G409gat_6[2]),.din(w_G409gat_1[2]));
	jspl jspl_w_G409gat_7(.douta(w_G409gat_7[0]),.doutb(w_G409gat_7[1]),.din(w_G409gat_2[0]));
	jspl3 jspl3_w_G426gat_0(.douta(w_G426gat_0[0]),.doutb(w_G426gat_0[1]),.doutc(w_G426gat_0[2]),.din(G426gat));
	jspl3 jspl3_w_G426gat_1(.douta(w_G426gat_1[0]),.doutb(w_G426gat_1[1]),.doutc(w_G426gat_1[2]),.din(w_G426gat_0[0]));
	jspl3 jspl3_w_G426gat_2(.douta(w_G426gat_2[0]),.doutb(w_G426gat_2[1]),.doutc(w_G426gat_2[2]),.din(w_G426gat_0[1]));
	jspl3 jspl3_w_G426gat_3(.douta(w_G426gat_3[0]),.doutb(w_G426gat_3[1]),.doutc(w_G426gat_3[2]),.din(w_G426gat_0[2]));
	jspl3 jspl3_w_G426gat_4(.douta(w_G426gat_4[0]),.doutb(w_G426gat_4[1]),.doutc(w_G426gat_4[2]),.din(w_G426gat_1[0]));
	jspl3 jspl3_w_G426gat_5(.douta(w_G426gat_5[0]),.doutb(w_G426gat_5[1]),.doutc(w_G426gat_5[2]),.din(w_G426gat_1[1]));
	jspl3 jspl3_w_G426gat_6(.douta(w_G426gat_6[0]),.doutb(w_G426gat_6[1]),.doutc(w_G426gat_6[2]),.din(w_G426gat_1[2]));
	jspl jspl_w_G426gat_7(.douta(w_G426gat_7[0]),.doutb(w_G426gat_7[1]),.din(w_G426gat_2[0]));
	jspl3 jspl3_w_G443gat_0(.douta(w_G443gat_0[0]),.doutb(w_G443gat_0[1]),.doutc(w_G443gat_0[2]),.din(G443gat));
	jspl3 jspl3_w_G443gat_1(.douta(w_G443gat_1[0]),.doutb(w_G443gat_1[1]),.doutc(w_G443gat_1[2]),.din(w_G443gat_0[0]));
	jspl3 jspl3_w_G443gat_2(.douta(w_G443gat_2[0]),.doutb(w_G443gat_2[1]),.doutc(w_G443gat_2[2]),.din(w_G443gat_0[1]));
	jspl3 jspl3_w_G443gat_3(.douta(w_G443gat_3[0]),.doutb(w_G443gat_3[1]),.doutc(w_G443gat_3[2]),.din(w_G443gat_0[2]));
	jspl3 jspl3_w_G443gat_4(.douta(w_G443gat_4[0]),.doutb(w_G443gat_4[1]),.doutc(w_G443gat_4[2]),.din(w_G443gat_1[0]));
	jspl3 jspl3_w_G443gat_5(.douta(w_G443gat_5[0]),.doutb(w_G443gat_5[1]),.doutc(w_G443gat_5[2]),.din(w_G443gat_1[1]));
	jspl3 jspl3_w_G443gat_6(.douta(w_G443gat_6[0]),.doutb(w_G443gat_6[1]),.doutc(w_G443gat_6[2]),.din(w_G443gat_1[2]));
	jspl jspl_w_G443gat_7(.douta(w_G443gat_7[0]),.doutb(w_G443gat_7[1]),.din(w_G443gat_2[0]));
	jspl3 jspl3_w_G460gat_0(.douta(w_G460gat_0[0]),.doutb(w_G460gat_0[1]),.doutc(w_G460gat_0[2]),.din(G460gat));
	jspl3 jspl3_w_G460gat_1(.douta(w_G460gat_1[0]),.doutb(w_G460gat_1[1]),.doutc(w_G460gat_1[2]),.din(w_G460gat_0[0]));
	jspl3 jspl3_w_G460gat_2(.douta(w_G460gat_2[0]),.doutb(w_G460gat_2[1]),.doutc(w_G460gat_2[2]),.din(w_G460gat_0[1]));
	jspl3 jspl3_w_G460gat_3(.douta(w_G460gat_3[0]),.doutb(w_G460gat_3[1]),.doutc(w_G460gat_3[2]),.din(w_G460gat_0[2]));
	jspl3 jspl3_w_G460gat_4(.douta(w_G460gat_4[0]),.doutb(w_G460gat_4[1]),.doutc(w_G460gat_4[2]),.din(w_G460gat_1[0]));
	jspl3 jspl3_w_G460gat_5(.douta(w_G460gat_5[0]),.doutb(w_G460gat_5[1]),.doutc(w_G460gat_5[2]),.din(w_G460gat_1[1]));
	jspl3 jspl3_w_G460gat_6(.douta(w_G460gat_6[0]),.doutb(w_G460gat_6[1]),.doutc(w_G460gat_6[2]),.din(w_G460gat_1[2]));
	jspl jspl_w_G460gat_7(.douta(w_G460gat_7[0]),.doutb(w_G460gat_7[1]),.din(w_G460gat_2[0]));
	jspl3 jspl3_w_G477gat_0(.douta(w_G477gat_0[0]),.doutb(w_G477gat_0[1]),.doutc(w_G477gat_0[2]),.din(G477gat));
	jspl3 jspl3_w_G477gat_1(.douta(w_G477gat_1[0]),.doutb(w_G477gat_1[1]),.doutc(w_G477gat_1[2]),.din(w_G477gat_0[0]));
	jspl3 jspl3_w_G477gat_2(.douta(w_G477gat_2[0]),.doutb(w_G477gat_2[1]),.doutc(w_G477gat_2[2]),.din(w_G477gat_0[1]));
	jspl3 jspl3_w_G477gat_3(.douta(w_G477gat_3[0]),.doutb(w_G477gat_3[1]),.doutc(w_G477gat_3[2]),.din(w_G477gat_0[2]));
	jspl3 jspl3_w_G477gat_4(.douta(w_G477gat_4[0]),.doutb(w_G477gat_4[1]),.doutc(w_G477gat_4[2]),.din(w_G477gat_1[0]));
	jspl3 jspl3_w_G477gat_5(.douta(w_G477gat_5[0]),.doutb(w_G477gat_5[1]),.doutc(w_G477gat_5[2]),.din(w_G477gat_1[1]));
	jspl3 jspl3_w_G477gat_6(.douta(w_G477gat_6[0]),.doutb(w_G477gat_6[1]),.doutc(w_G477gat_6[2]),.din(w_G477gat_1[2]));
	jspl jspl_w_G477gat_7(.douta(w_G477gat_7[0]),.doutb(w_G477gat_7[1]),.din(w_G477gat_2[0]));
	jspl3 jspl3_w_G494gat_0(.douta(w_G494gat_0[0]),.doutb(w_G494gat_0[1]),.doutc(w_G494gat_0[2]),.din(G494gat));
	jspl3 jspl3_w_G494gat_1(.douta(w_G494gat_1[0]),.doutb(w_G494gat_1[1]),.doutc(w_G494gat_1[2]),.din(w_G494gat_0[0]));
	jspl3 jspl3_w_G494gat_2(.douta(w_G494gat_2[0]),.doutb(w_G494gat_2[1]),.doutc(w_G494gat_2[2]),.din(w_G494gat_0[1]));
	jspl3 jspl3_w_G494gat_3(.douta(w_G494gat_3[0]),.doutb(w_G494gat_3[1]),.doutc(w_G494gat_3[2]),.din(w_G494gat_0[2]));
	jspl3 jspl3_w_G494gat_4(.douta(w_G494gat_4[0]),.doutb(w_G494gat_4[1]),.doutc(w_G494gat_4[2]),.din(w_G494gat_1[0]));
	jspl3 jspl3_w_G494gat_5(.douta(w_G494gat_5[0]),.doutb(w_G494gat_5[1]),.doutc(w_G494gat_5[2]),.din(w_G494gat_1[1]));
	jspl3 jspl3_w_G494gat_6(.douta(w_G494gat_6[0]),.doutb(w_G494gat_6[1]),.doutc(w_G494gat_6[2]),.din(w_G494gat_1[2]));
	jspl jspl_w_G494gat_7(.douta(w_G494gat_7[0]),.doutb(w_G494gat_7[1]),.din(w_G494gat_2[0]));
	jspl3 jspl3_w_G511gat_0(.douta(w_G511gat_0[0]),.doutb(w_G511gat_0[1]),.doutc(w_G511gat_0[2]),.din(G511gat));
	jspl3 jspl3_w_G511gat_1(.douta(w_G511gat_1[0]),.doutb(w_G511gat_1[1]),.doutc(w_G511gat_1[2]),.din(w_G511gat_0[0]));
	jspl3 jspl3_w_G511gat_2(.douta(w_G511gat_2[0]),.doutb(w_G511gat_2[1]),.doutc(w_G511gat_2[2]),.din(w_G511gat_0[1]));
	jspl3 jspl3_w_G511gat_3(.douta(w_G511gat_3[0]),.doutb(w_G511gat_3[1]),.doutc(w_G511gat_3[2]),.din(w_G511gat_0[2]));
	jspl3 jspl3_w_G511gat_4(.douta(w_G511gat_4[0]),.doutb(w_G511gat_4[1]),.doutc(w_G511gat_4[2]),.din(w_G511gat_1[0]));
	jspl3 jspl3_w_G511gat_5(.douta(w_G511gat_5[0]),.doutb(w_G511gat_5[1]),.doutc(w_G511gat_5[2]),.din(w_G511gat_1[1]));
	jspl3 jspl3_w_G511gat_6(.douta(w_G511gat_6[0]),.doutb(w_G511gat_6[1]),.doutc(w_G511gat_6[2]),.din(w_G511gat_1[2]));
	jspl jspl_w_G511gat_7(.douta(w_G511gat_7[0]),.doutb(w_G511gat_7[1]),.din(w_G511gat_2[0]));
	jspl3 jspl3_w_G528gat_0(.douta(w_G528gat_0[0]),.doutb(w_G528gat_0[1]),.doutc(w_G528gat_0[2]),.din(G528gat));
	jspl3 jspl3_w_G528gat_1(.douta(w_G528gat_1[0]),.doutb(w_G528gat_1[1]),.doutc(w_G528gat_1[2]),.din(w_G528gat_0[0]));
	jspl3 jspl3_w_G528gat_2(.douta(w_G528gat_2[0]),.doutb(w_G528gat_2[1]),.doutc(w_G528gat_2[2]),.din(w_G528gat_0[1]));
	jspl3 jspl3_w_G528gat_3(.douta(w_G528gat_3[0]),.doutb(w_G528gat_3[1]),.doutc(w_G528gat_3[2]),.din(w_G528gat_0[2]));
	jspl3 jspl3_w_G528gat_4(.douta(w_G528gat_4[0]),.doutb(w_G528gat_4[1]),.doutc(w_G528gat_4[2]),.din(w_G528gat_1[0]));
	jspl3 jspl3_w_G528gat_5(.douta(w_G528gat_5[0]),.doutb(w_G528gat_5[1]),.doutc(w_G528gat_5[2]),.din(w_G528gat_1[1]));
	jspl3 jspl3_w_G528gat_6(.douta(w_G528gat_6[0]),.doutb(w_G528gat_6[1]),.doutc(w_G528gat_6[2]),.din(w_G528gat_1[2]));
	jspl jspl_w_G528gat_7(.douta(w_G528gat_7[0]),.doutb(w_G528gat_7[1]),.din(w_G528gat_2[0]));
	jspl jspl_w_G545gat_0(.douta(w_G545gat_0),.doutb(G545gat),.din(G545gat_fa_));
	jspl jspl_w_n65_0(.douta(w_n65_0[0]),.doutb(w_n65_0[1]),.din(n65));
	jspl jspl_w_n69_0(.douta(w_dff_A_PMzkp3Yy3_0),.doutb(w_n69_0[1]),.din(n69));
	jspl jspl_w_n70_0(.douta(w_n70_0[0]),.doutb(w_n70_0[1]),.din(n70));
	jspl jspl_w_n72_0(.douta(w_dff_A_wr6o7ltw7_0),.doutb(w_n72_0[1]),.din(n72));
	jspl jspl_w_n75_0(.douta(w_n75_0[0]),.doutb(w_n75_0[1]),.din(n75));
	jspl jspl_w_n77_0(.douta(w_n77_0[0]),.doutb(w_n77_0[1]),.din(n77));
	jspl jspl_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.din(n78));
	jspl jspl_w_n81_0(.douta(w_n81_0[0]),.doutb(w_n81_0[1]),.din(n81));
	jspl3 jspl3_w_n82_0(.douta(w_n82_0[0]),.doutb(w_dff_A_b7ZXtC620_1),.doutc(w_dff_A_XQ7rHGXI6_2),.din(n82));
	jspl jspl_w_n82_1(.douta(w_n82_1[0]),.doutb(w_n82_1[1]),.din(w_n82_0[0]));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl jspl_w_n85_0(.douta(w_n85_0[0]),.doutb(w_n85_0[1]),.din(n85));
	jspl jspl_w_n87_0(.douta(w_n87_0[0]),.doutb(w_n87_0[1]),.din(n87));
	jspl jspl_w_n89_0(.douta(w_dff_A_Sb20tTNi4_0),.doutb(w_n89_0[1]),.din(n89));
	jspl jspl_w_n93_0(.douta(w_dff_A_QEwu1QkQ3_0),.doutb(w_n93_0[1]),.din(w_dff_B_jI2yWL6q9_2));
	jspl jspl_w_n94_0(.douta(w_dff_A_yoFFnUwE3_0),.doutb(w_n94_0[1]),.din(n94));
	jspl jspl_w_n96_0(.douta(w_n96_0[0]),.doutb(w_n96_0[1]),.din(n96));
	jspl jspl_w_n99_0(.douta(w_n99_0[0]),.doutb(w_n99_0[1]),.din(n99));
	jspl3 jspl3_w_n100_0(.douta(w_n100_0[0]),.doutb(w_dff_A_RUhPeT7s8_1),.doutc(w_dff_A_7OiKETeF1_2),.din(n100));
	jspl jspl_w_n100_1(.douta(w_n100_1[0]),.doutb(w_n100_1[1]),.din(w_n100_0[0]));
	jspl3 jspl3_w_n101_0(.douta(w_n101_0[0]),.doutb(w_n101_0[1]),.doutc(w_n101_0[2]),.din(n101));
	jspl jspl_w_n103_0(.douta(w_n103_0[0]),.doutb(w_dff_A_dJ1rZgd00_1),.din(n103));
	jspl jspl_w_n104_0(.douta(w_n104_0[0]),.doutb(w_n104_0[1]),.din(n104));
	jspl jspl_w_n107_0(.douta(w_n107_0[0]),.doutb(w_n107_0[1]),.din(n107));
	jspl jspl_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n110_0(.douta(w_dff_A_WdwwOVyQ8_0),.doutb(w_n110_0[1]),.din(n110));
	jspl jspl_w_n115_0(.douta(w_dff_A_lXilLWhR4_0),.doutb(w_n115_0[1]),.din(w_dff_B_o082cFWp4_2));
	jspl jspl_w_n116_0(.douta(w_dff_A_SAPjTpMh1_0),.doutb(w_n116_0[1]),.din(n116));
	jspl3 jspl3_w_n126_0(.douta(w_n126_0[0]),.doutb(w_dff_A_bOg8qe9P3_1),.doutc(w_dff_A_bfPY2yka7_2),.din(w_dff_B_qFGeQJ162_3));
	jspl jspl_w_n128_0(.douta(w_n128_0[0]),.doutb(w_n128_0[1]),.din(w_dff_B_DMlKtyFT9_2));
	jspl jspl_w_n129_0(.douta(w_n129_0[0]),.doutb(w_n129_0[1]),.din(n129));
	jspl jspl_w_n130_0(.douta(w_n130_0[0]),.doutb(w_dff_A_RCAO2G978_1),.din(n130));
	jspl jspl_w_n131_0(.douta(w_n131_0[0]),.doutb(w_n131_0[1]),.din(n131));
	jspl3 jspl3_w_n132_0(.douta(w_dff_A_kmyc9HRq1_0),.doutb(w_n132_0[1]),.doutc(w_n132_0[2]),.din(n132));
	jspl3 jspl3_w_n133_0(.douta(w_n133_0[0]),.doutb(w_n133_0[1]),.doutc(w_n133_0[2]),.din(n133));
	jspl jspl_w_n138_0(.douta(w_n138_0[0]),.doutb(w_n138_0[1]),.din(n138));
	jspl jspl_w_n139_0(.douta(w_n139_0[0]),.doutb(w_n139_0[1]),.din(n139));
	jspl jspl_w_n140_0(.douta(w_n140_0[0]),.doutb(w_n140_0[1]),.din(n140));
	jspl jspl_w_n142_0(.douta(w_n142_0[0]),.doutb(w_n142_0[1]),.din(n142));
	jspl jspl_w_n143_0(.douta(w_n143_0[0]),.doutb(w_n143_0[1]),.din(n143));
	jspl jspl_w_n145_0(.douta(w_dff_A_7HPLrMCC8_0),.doutb(w_n145_0[1]),.din(n145));
	jspl jspl_w_n150_0(.douta(w_dff_A_TenYRsws0_0),.doutb(w_n150_0[1]),.din(n150));
	jspl jspl_w_n151_0(.douta(w_dff_A_ZbpznAsK3_0),.doutb(w_n151_0[1]),.din(n151));
	jspl3 jspl3_w_n156_0(.douta(w_n156_0[0]),.doutb(w_dff_A_GAQ3BWky2_1),.doutc(w_dff_A_4x3nTySY4_2),.din(n156));
	jspl jspl_w_n158_0(.douta(w_n158_0[0]),.doutb(w_n158_0[1]),.din(w_dff_B_d3eFCLjg4_2));
	jspl jspl_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.din(n163));
	jspl jspl_w_n165_0(.douta(w_n165_0[0]),.doutb(w_n165_0[1]),.din(w_dff_B_mHt9CsSX7_2));
	jspl jspl_w_n166_0(.douta(w_n166_0[0]),.doutb(w_n166_0[1]),.din(n166));
	jspl jspl_w_n168_0(.douta(w_n168_0[0]),.doutb(w_n168_0[1]),.din(n168));
	jspl3 jspl3_w_n169_0(.douta(w_dff_A_89r2owrF7_0),.doutb(w_dff_A_bs6TpDgl8_1),.doutc(w_n169_0[2]),.din(n169));
	jspl jspl_w_n170_0(.douta(w_n170_0[0]),.doutb(w_n170_0[1]),.din(n170));
	jspl jspl_w_n172_0(.douta(w_n172_0[0]),.doutb(w_n172_0[1]),.din(n172));
	jspl jspl_w_n174_0(.douta(w_n174_0[0]),.doutb(w_n174_0[1]),.din(n174));
	jspl jspl_w_n175_0(.douta(w_n175_0[0]),.doutb(w_n175_0[1]),.din(w_dff_B_r8aFdsh71_2));
	jspl jspl_w_n176_0(.douta(w_n176_0[0]),.doutb(w_n176_0[1]),.din(n176));
	jspl jspl_w_n177_0(.douta(w_n177_0[0]),.doutb(w_n177_0[1]),.din(n177));
	jspl jspl_w_n178_0(.douta(w_n178_0[0]),.doutb(w_n178_0[1]),.din(n178));
	jspl jspl_w_n180_0(.douta(w_n180_0[0]),.doutb(w_n180_0[1]),.din(n180));
	jspl jspl_w_n181_0(.douta(w_n181_0[0]),.doutb(w_n181_0[1]),.din(n181));
	jspl jspl_w_n183_0(.douta(w_dff_A_mnSlSRY63_0),.doutb(w_n183_0[1]),.din(n183));
	jspl jspl_w_n188_0(.douta(w_dff_A_LL0DfKUa1_0),.doutb(w_n188_0[1]),.din(n188));
	jspl jspl_w_n189_0(.douta(w_dff_A_qj5HAMpT0_0),.doutb(w_n189_0[1]),.din(n189));
	jspl3 jspl3_w_n194_0(.douta(w_n194_0[0]),.doutb(w_dff_A_0Nvok6OE8_1),.doutc(w_dff_A_sokiXTn82_2),.din(n194));
	jspl jspl_w_n196_0(.douta(w_n196_0[0]),.doutb(w_n196_0[1]),.din(w_dff_B_0YPYM2yI9_2));
	jspl jspl_w_n199_0(.douta(w_n199_0[0]),.doutb(w_n199_0[1]),.din(n199));
	jspl jspl_w_n201_0(.douta(w_n201_0[0]),.doutb(w_n201_0[1]),.din(w_dff_B_nNtLFeVt4_2));
	jspl jspl_w_n204_0(.douta(w_n204_0[0]),.doutb(w_n204_0[1]),.din(n204));
	jspl jspl_w_n206_0(.douta(w_n206_0[0]),.doutb(w_n206_0[1]),.din(w_dff_B_PZOVoV967_2));
	jspl jspl_w_n207_0(.douta(w_n207_0[0]),.doutb(w_n207_0[1]),.din(n207));
	jspl jspl_w_n209_0(.douta(w_n209_0[0]),.doutb(w_n209_0[1]),.din(n209));
	jspl3 jspl3_w_n210_0(.douta(w_n210_0[0]),.doutb(w_dff_A_lTu2GWwo3_1),.doutc(w_dff_A_jkneepKI9_2),.din(n210));
	jspl jspl_w_n210_1(.douta(w_dff_A_9f3FoyNE9_0),.doutb(w_n210_1[1]),.din(w_n210_0[0]));
	jspl jspl_w_n213_0(.douta(w_n213_0[0]),.doutb(w_n213_0[1]),.din(n213));
	jspl jspl_w_n215_0(.douta(w_n215_0[0]),.doutb(w_n215_0[1]),.din(n215));
	jspl jspl_w_n216_0(.douta(w_n216_0[0]),.doutb(w_n216_0[1]),.din(n216));
	jspl jspl_w_n217_0(.douta(w_n217_0[0]),.doutb(w_n217_0[1]),.din(n217));
	jspl jspl_w_n218_0(.douta(w_n218_0[0]),.doutb(w_n218_0[1]),.din(w_dff_B_KV0W7Hdu4_2));
	jspl jspl_w_n219_0(.douta(w_n219_0[0]),.doutb(w_n219_0[1]),.din(n219));
	jspl jspl_w_n220_0(.douta(w_n220_0[0]),.doutb(w_n220_0[1]),.din(n220));
	jspl jspl_w_n221_0(.douta(w_n221_0[0]),.doutb(w_n221_0[1]),.din(n221));
	jspl jspl_w_n223_0(.douta(w_n223_0[0]),.doutb(w_n223_0[1]),.din(n223));
	jspl jspl_w_n224_0(.douta(w_n224_0[0]),.doutb(w_n224_0[1]),.din(n224));
	jspl jspl_w_n226_0(.douta(w_dff_A_AQFbMP098_0),.doutb(w_n226_0[1]),.din(n226));
	jspl jspl_w_n231_0(.douta(w_dff_A_oDeo4JQK6_0),.doutb(w_n231_0[1]),.din(n231));
	jspl jspl_w_n232_0(.douta(w_dff_A_2UH2CFTH9_0),.doutb(w_n232_0[1]),.din(n232));
	jspl3 jspl3_w_n237_0(.douta(w_n237_0[0]),.doutb(w_dff_A_3RUgPuw28_1),.doutc(w_dff_A_X5hDfQDj5_2),.din(n237));
	jspl jspl_w_n239_0(.douta(w_n239_0[0]),.doutb(w_n239_0[1]),.din(w_dff_B_o5szB85e1_2));
	jspl jspl_w_n242_0(.douta(w_n242_0[0]),.doutb(w_n242_0[1]),.din(n242));
	jspl jspl_w_n244_0(.douta(w_n244_0[0]),.doutb(w_n244_0[1]),.din(w_dff_B_xmctGBj18_2));
	jspl jspl_w_n247_0(.douta(w_n247_0[0]),.doutb(w_n247_0[1]),.din(w_dff_B_TOOe7Jno0_2));
	jspl jspl_w_n249_0(.douta(w_n249_0[0]),.doutb(w_n249_0[1]),.din(w_dff_B_TQjrYt633_2));
	jspl jspl_w_n252_0(.douta(w_n252_0[0]),.doutb(w_n252_0[1]),.din(w_dff_B_TCPyOj6B9_2));
	jspl jspl_w_n254_0(.douta(w_n254_0[0]),.doutb(w_n254_0[1]),.din(w_dff_B_VKVv2ZlL7_2));
	jspl jspl_w_n255_0(.douta(w_n255_0[0]),.doutb(w_n255_0[1]),.din(n255));
	jspl jspl_w_n257_0(.douta(w_n257_0[0]),.doutb(w_n257_0[1]),.din(n257));
	jspl3 jspl3_w_n258_0(.douta(w_dff_A_skMxtdkH5_0),.doutb(w_dff_A_8wznEIJ80_1),.doutc(w_n258_0[2]),.din(n258));
	jspl jspl_w_n259_0(.douta(w_n259_0[0]),.doutb(w_n259_0[1]),.din(n259));
	jspl jspl_w_n261_0(.douta(w_n261_0[0]),.doutb(w_dff_A_sffExBlQ5_1),.din(n261));
	jspl jspl_w_n264_0(.douta(w_n264_0[0]),.doutb(w_n264_0[1]),.din(n264));
	jspl jspl_w_n265_0(.douta(w_n265_0[0]),.doutb(w_n265_0[1]),.din(n265));
	jspl jspl_w_n266_0(.douta(w_n266_0[0]),.doutb(w_n266_0[1]),.din(n266));
	jspl jspl_w_n267_0(.douta(w_n267_0[0]),.doutb(w_n267_0[1]),.din(n267));
	jspl jspl_w_n268_0(.douta(w_n268_0[0]),.doutb(w_n268_0[1]),.din(n268));
	jspl jspl_w_n269_0(.douta(w_n269_0[0]),.doutb(w_n269_0[1]),.din(n269));
	jspl jspl_w_n270_0(.douta(w_n270_0[0]),.doutb(w_n270_0[1]),.din(n270));
	jspl jspl_w_n271_0(.douta(w_n271_0[0]),.doutb(w_n271_0[1]),.din(n271));
	jspl jspl_w_n272_0(.douta(w_n272_0[0]),.doutb(w_n272_0[1]),.din(n272));
	jspl jspl_w_n274_0(.douta(w_n274_0[0]),.doutb(w_n274_0[1]),.din(n274));
	jspl jspl_w_n275_0(.douta(w_n275_0[0]),.doutb(w_n275_0[1]),.din(n275));
	jspl jspl_w_n277_0(.douta(w_dff_A_m3nABioh9_0),.doutb(w_n277_0[1]),.din(n277));
	jspl jspl_w_n282_0(.douta(w_dff_A_C95lVcqm2_0),.doutb(w_n282_0[1]),.din(n282));
	jspl jspl_w_n283_0(.douta(w_dff_A_Oeb4iY3b9_0),.doutb(w_n283_0[1]),.din(n283));
	jspl3 jspl3_w_n288_0(.douta(w_n288_0[0]),.doutb(w_dff_A_dKDe0QPZ5_1),.doutc(w_dff_A_DvKWN5fh7_2),.din(n288));
	jspl jspl_w_n290_0(.douta(w_n290_0[0]),.doutb(w_n290_0[1]),.din(w_dff_B_669JR3NH1_2));
	jspl jspl_w_n293_0(.douta(w_n293_0[0]),.doutb(w_n293_0[1]),.din(n293));
	jspl jspl_w_n295_0(.douta(w_n295_0[0]),.doutb(w_n295_0[1]),.din(w_dff_B_M5SDinXi6_2));
	jspl jspl_w_n298_0(.douta(w_n298_0[0]),.doutb(w_n298_0[1]),.din(n298));
	jspl jspl_w_n300_0(.douta(w_n300_0[0]),.doutb(w_n300_0[1]),.din(w_dff_B_n7O6EScb1_2));
	jspl jspl_w_n303_0(.douta(w_n303_0[0]),.doutb(w_n303_0[1]),.din(n303));
	jspl jspl_w_n305_0(.douta(w_n305_0[0]),.doutb(w_n305_0[1]),.din(w_dff_B_iy6eoe9I4_2));
	jspl jspl_w_n308_0(.douta(w_n308_0[0]),.doutb(w_n308_0[1]),.din(n308));
	jspl jspl_w_n310_0(.douta(w_n310_0[0]),.doutb(w_n310_0[1]),.din(w_dff_B_dnWkgseM9_2));
	jspl jspl_w_n311_0(.douta(w_n311_0[0]),.doutb(w_n311_0[1]),.din(n311));
	jspl jspl_w_n313_0(.douta(w_n313_0[0]),.doutb(w_n313_0[1]),.din(n313));
	jspl3 jspl3_w_n314_0(.douta(w_dff_A_0wMb0ngO3_0),.doutb(w_dff_A_mzOkYWKK3_1),.doutc(w_n314_0[2]),.din(n314));
	jspl jspl_w_n315_0(.douta(w_n315_0[0]),.doutb(w_n315_0[1]),.din(n315));
	jspl jspl_w_n317_0(.douta(w_n317_0[0]),.doutb(w_dff_A_VcZH5Esl6_1),.din(n317));
	jspl jspl_w_n320_0(.douta(w_n320_0[0]),.doutb(w_n320_0[1]),.din(n320));
	jspl jspl_w_n321_0(.douta(w_n321_0[0]),.doutb(w_n321_0[1]),.din(n321));
	jspl jspl_w_n322_0(.douta(w_n322_0[0]),.doutb(w_n322_0[1]),.din(n322));
	jspl jspl_w_n323_0(.douta(w_n323_0[0]),.doutb(w_n323_0[1]),.din(n323));
	jspl jspl_w_n324_0(.douta(w_n324_0[0]),.doutb(w_n324_0[1]),.din(n324));
	jspl jspl_w_n325_0(.douta(w_n325_0[0]),.doutb(w_n325_0[1]),.din(n325));
	jspl jspl_w_n326_0(.douta(w_n326_0[0]),.doutb(w_n326_0[1]),.din(n326));
	jspl jspl_w_n327_0(.douta(w_n327_0[0]),.doutb(w_n327_0[1]),.din(n327));
	jspl jspl_w_n328_0(.douta(w_n328_0[0]),.doutb(w_n328_0[1]),.din(n328));
	jspl jspl_w_n329_0(.douta(w_n329_0[0]),.doutb(w_n329_0[1]),.din(n329));
	jspl jspl_w_n330_0(.douta(w_n330_0[0]),.doutb(w_n330_0[1]),.din(n330));
	jspl jspl_w_n332_0(.douta(w_n332_0[0]),.doutb(w_n332_0[1]),.din(n332));
	jspl jspl_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.din(n333));
	jspl jspl_w_n335_0(.douta(w_dff_A_Vez93m5r5_0),.doutb(w_n335_0[1]),.din(n335));
	jspl jspl_w_n340_0(.douta(w_dff_A_2T7pXLSx7_0),.doutb(w_n340_0[1]),.din(n340));
	jspl jspl_w_n341_0(.douta(w_dff_A_bzzSIQF31_0),.doutb(w_n341_0[1]),.din(n341));
	jspl3 jspl3_w_n346_0(.douta(w_n346_0[0]),.doutb(w_dff_A_eQlOczic5_1),.doutc(w_dff_A_H17Bjt2h2_2),.din(n346));
	jspl jspl_w_n348_0(.douta(w_n348_0[0]),.doutb(w_n348_0[1]),.din(w_dff_B_P7GxG97t3_2));
	jspl jspl_w_n351_0(.douta(w_n351_0[0]),.doutb(w_n351_0[1]),.din(n351));
	jspl jspl_w_n353_0(.douta(w_n353_0[0]),.doutb(w_n353_0[1]),.din(w_dff_B_Z8BhLEVE3_2));
	jspl jspl_w_n356_0(.douta(w_n356_0[0]),.doutb(w_n356_0[1]),.din(n356));
	jspl jspl_w_n358_0(.douta(w_n358_0[0]),.doutb(w_n358_0[1]),.din(w_dff_B_ewWnwWek2_2));
	jspl jspl_w_n361_0(.douta(w_n361_0[0]),.doutb(w_n361_0[1]),.din(n361));
	jspl jspl_w_n363_0(.douta(w_n363_0[0]),.doutb(w_n363_0[1]),.din(w_dff_B_5ER2SwBJ6_2));
	jspl jspl_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.din(n366));
	jspl jspl_w_n368_0(.douta(w_n368_0[0]),.doutb(w_n368_0[1]),.din(w_dff_B_2O4uTLYz9_2));
	jspl jspl_w_n371_0(.douta(w_n371_0[0]),.doutb(w_n371_0[1]),.din(n371));
	jspl jspl_w_n372_0(.douta(w_n372_0[0]),.doutb(w_dff_A_dfd1enHt4_1),.din(n372));
	jspl jspl_w_n373_0(.douta(w_n373_0[0]),.doutb(w_n373_0[1]),.din(n373));
	jspl jspl_w_n375_0(.douta(w_n375_0[0]),.doutb(w_n375_0[1]),.din(n375));
	jspl3 jspl3_w_n376_0(.douta(w_dff_A_LyIyUKHN6_0),.doutb(w_dff_A_2sY683Rr3_1),.doutc(w_n376_0[2]),.din(n376));
	jspl jspl_w_n377_0(.douta(w_n377_0[0]),.doutb(w_n377_0[1]),.din(n377));
	jspl jspl_w_n380_0(.douta(w_dff_A_vJmeg3EW2_0),.doutb(w_n380_0[1]),.din(n380));
	jspl jspl_w_n382_0(.douta(w_n382_0[0]),.doutb(w_n382_0[1]),.din(n382));
	jspl jspl_w_n383_0(.douta(w_n383_0[0]),.doutb(w_n383_0[1]),.din(w_dff_B_xZpEN1Py9_2));
	jspl jspl_w_n384_0(.douta(w_n384_0[0]),.doutb(w_n384_0[1]),.din(n384));
	jspl jspl_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.din(n385));
	jspl jspl_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.din(n386));
	jspl jspl_w_n387_0(.douta(w_n387_0[0]),.doutb(w_n387_0[1]),.din(n387));
	jspl jspl_w_n388_0(.douta(w_n388_0[0]),.doutb(w_n388_0[1]),.din(n388));
	jspl jspl_w_n389_0(.douta(w_n389_0[0]),.doutb(w_n389_0[1]),.din(n389));
	jspl jspl_w_n390_0(.douta(w_n390_0[0]),.doutb(w_n390_0[1]),.din(n390));
	jspl jspl_w_n391_0(.douta(w_n391_0[0]),.doutb(w_n391_0[1]),.din(n391));
	jspl jspl_w_n392_0(.douta(w_n392_0[0]),.doutb(w_n392_0[1]),.din(n392));
	jspl jspl_w_n393_0(.douta(w_n393_0[0]),.doutb(w_n393_0[1]),.din(n393));
	jspl jspl_w_n394_0(.douta(w_n394_0[0]),.doutb(w_n394_0[1]),.din(n394));
	jspl jspl_w_n396_0(.douta(w_n396_0[0]),.doutb(w_n396_0[1]),.din(n396));
	jspl jspl_w_n397_0(.douta(w_n397_0[0]),.doutb(w_n397_0[1]),.din(n397));
	jspl jspl_w_n399_0(.douta(w_dff_A_hM36iCne8_0),.doutb(w_n399_0[1]),.din(n399));
	jspl jspl_w_n404_0(.douta(w_dff_A_TVX9hYFf4_0),.doutb(w_n404_0[1]),.din(n404));
	jspl jspl_w_n405_0(.douta(w_dff_A_lXR94XaA4_0),.doutb(w_n405_0[1]),.din(n405));
	jspl3 jspl3_w_n410_0(.douta(w_n410_0[0]),.doutb(w_dff_A_vf10omxW1_1),.doutc(w_dff_A_v08tLeep6_2),.din(n410));
	jspl jspl_w_n412_0(.douta(w_n412_0[0]),.doutb(w_n412_0[1]),.din(w_dff_B_TL6QGUTC1_2));
	jspl jspl_w_n415_0(.douta(w_n415_0[0]),.doutb(w_n415_0[1]),.din(n415));
	jspl jspl_w_n417_0(.douta(w_n417_0[0]),.doutb(w_n417_0[1]),.din(w_dff_B_MGReRU7o3_2));
	jspl jspl_w_n420_0(.douta(w_n420_0[0]),.doutb(w_n420_0[1]),.din(n420));
	jspl jspl_w_n422_0(.douta(w_n422_0[0]),.doutb(w_n422_0[1]),.din(w_dff_B_Gpq1DOjM2_2));
	jspl jspl_w_n425_0(.douta(w_n425_0[0]),.doutb(w_n425_0[1]),.din(n425));
	jspl jspl_w_n427_0(.douta(w_n427_0[0]),.doutb(w_n427_0[1]),.din(w_dff_B_EA0egYHr7_2));
	jspl jspl_w_n430_0(.douta(w_n430_0[0]),.doutb(w_n430_0[1]),.din(n430));
	jspl jspl_w_n432_0(.douta(w_n432_0[0]),.doutb(w_n432_0[1]),.din(w_dff_B_4f0QssU07_2));
	jspl jspl_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.din(n435));
	jspl jspl_w_n437_0(.douta(w_n437_0[0]),.doutb(w_n437_0[1]),.din(w_dff_B_q6FLbAux0_2));
	jspl jspl_w_n441_0(.douta(w_n441_0[0]),.doutb(w_n441_0[1]),.din(n441));
	jspl jspl_w_n442_0(.douta(w_n442_0[0]),.doutb(w_dff_A_ZUEwSf3U7_1),.din(n442));
	jspl jspl_w_n443_0(.douta(w_n443_0[0]),.doutb(w_n443_0[1]),.din(n443));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl3 jspl3_w_n446_0(.douta(w_dff_A_HhWBU4898_0),.doutb(w_dff_A_2TJbBS0Z7_1),.doutc(w_n446_0[2]),.din(n446));
	jspl jspl_w_n447_0(.douta(w_n447_0[0]),.doutb(w_n447_0[1]),.din(n447));
	jspl jspl_w_n450_0(.douta(w_dff_A_VSjoUpi55_0),.doutb(w_n450_0[1]),.din(n450));
	jspl jspl_w_n452_0(.douta(w_n452_0[0]),.doutb(w_n452_0[1]),.din(n452));
	jspl jspl_w_n453_0(.douta(w_n453_0[0]),.doutb(w_n453_0[1]),.din(w_dff_B_GAwbNi6N6_2));
	jspl jspl_w_n454_0(.douta(w_n454_0[0]),.doutb(w_n454_0[1]),.din(n454));
	jspl jspl_w_n455_0(.douta(w_n455_0[0]),.doutb(w_n455_0[1]),.din(n455));
	jspl jspl_w_n456_0(.douta(w_n456_0[0]),.doutb(w_n456_0[1]),.din(n456));
	jspl jspl_w_n457_0(.douta(w_n457_0[0]),.doutb(w_n457_0[1]),.din(n457));
	jspl jspl_w_n458_0(.douta(w_n458_0[0]),.doutb(w_n458_0[1]),.din(n458));
	jspl jspl_w_n459_0(.douta(w_n459_0[0]),.doutb(w_n459_0[1]),.din(n459));
	jspl jspl_w_n460_0(.douta(w_n460_0[0]),.doutb(w_n460_0[1]),.din(n460));
	jspl jspl_w_n461_0(.douta(w_n461_0[0]),.doutb(w_n461_0[1]),.din(n461));
	jspl jspl_w_n462_0(.douta(w_n462_0[0]),.doutb(w_n462_0[1]),.din(n462));
	jspl jspl_w_n463_0(.douta(w_n463_0[0]),.doutb(w_n463_0[1]),.din(n463));
	jspl jspl_w_n464_0(.douta(w_n464_0[0]),.doutb(w_n464_0[1]),.din(n464));
	jspl jspl_w_n465_0(.douta(w_n465_0[0]),.doutb(w_n465_0[1]),.din(n465));
	jspl jspl_w_n466_0(.douta(w_n466_0[0]),.doutb(w_n466_0[1]),.din(n466));
	jspl jspl_w_n468_0(.douta(w_n468_0[0]),.doutb(w_n468_0[1]),.din(n468));
	jspl jspl_w_n469_0(.douta(w_n469_0[0]),.doutb(w_n469_0[1]),.din(n469));
	jspl jspl_w_n471_0(.douta(w_dff_A_vEIwA6aA0_0),.doutb(w_n471_0[1]),.din(n471));
	jspl jspl_w_n476_0(.douta(w_dff_A_swXZQXih8_0),.doutb(w_n476_0[1]),.din(n476));
	jspl jspl_w_n477_0(.douta(w_dff_A_779Ly5To1_0),.doutb(w_n477_0[1]),.din(n477));
	jspl3 jspl3_w_n482_0(.douta(w_n482_0[0]),.doutb(w_dff_A_iwf7vElC1_1),.doutc(w_dff_A_px4TwLna7_2),.din(n482));
	jspl jspl_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.din(w_dff_B_2aqVfDn05_2));
	jspl jspl_w_n487_0(.douta(w_n487_0[0]),.doutb(w_n487_0[1]),.din(n487));
	jspl jspl_w_n489_0(.douta(w_n489_0[0]),.doutb(w_n489_0[1]),.din(w_dff_B_TVLIDS2Y9_2));
	jspl jspl_w_n492_0(.douta(w_n492_0[0]),.doutb(w_n492_0[1]),.din(n492));
	jspl jspl_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.din(w_dff_B_ioksKqhM3_2));
	jspl jspl_w_n497_0(.douta(w_n497_0[0]),.doutb(w_n497_0[1]),.din(n497));
	jspl jspl_w_n499_0(.douta(w_n499_0[0]),.doutb(w_n499_0[1]),.din(w_dff_B_iyTxPbzz4_2));
	jspl jspl_w_n502_0(.douta(w_n502_0[0]),.doutb(w_n502_0[1]),.din(n502));
	jspl jspl_w_n504_0(.douta(w_n504_0[0]),.doutb(w_n504_0[1]),.din(w_dff_B_lKp0G3Gz6_2));
	jspl jspl_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.din(n507));
	jspl jspl_w_n509_0(.douta(w_n509_0[0]),.doutb(w_n509_0[1]),.din(w_dff_B_pxhg50Db2_2));
	jspl jspl_w_n512_0(.douta(w_n512_0[0]),.doutb(w_n512_0[1]),.din(n512));
	jspl jspl_w_n514_0(.douta(w_n514_0[0]),.doutb(w_n514_0[1]),.din(w_dff_B_4Nkw4hr37_2));
	jspl jspl_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.din(n518));
	jspl jspl_w_n519_0(.douta(w_n519_0[0]),.doutb(w_dff_A_RG9ph2SF1_1),.din(n519));
	jspl jspl_w_n520_0(.douta(w_n520_0[0]),.doutb(w_n520_0[1]),.din(n520));
	jspl jspl_w_n522_0(.douta(w_n522_0[0]),.doutb(w_n522_0[1]),.din(n522));
	jspl3 jspl3_w_n523_0(.douta(w_dff_A_jLjA2Bfy3_0),.doutb(w_dff_A_drno1gMW4_1),.doutc(w_n523_0[2]),.din(n523));
	jspl jspl_w_n524_0(.douta(w_n524_0[0]),.doutb(w_n524_0[1]),.din(n524));
	jspl jspl_w_n527_0(.douta(w_dff_A_KFl8vlWw0_0),.doutb(w_n527_0[1]),.din(n527));
	jspl jspl_w_n529_0(.douta(w_n529_0[0]),.doutb(w_n529_0[1]),.din(n529));
	jspl jspl_w_n530_0(.douta(w_n530_0[0]),.doutb(w_n530_0[1]),.din(w_dff_B_3rRbXLt23_2));
	jspl jspl_w_n531_0(.douta(w_n531_0[0]),.doutb(w_n531_0[1]),.din(n531));
	jspl jspl_w_n532_0(.douta(w_n532_0[0]),.doutb(w_n532_0[1]),.din(n532));
	jspl jspl_w_n533_0(.douta(w_n533_0[0]),.doutb(w_n533_0[1]),.din(n533));
	jspl jspl_w_n534_0(.douta(w_n534_0[0]),.doutb(w_n534_0[1]),.din(n534));
	jspl jspl_w_n535_0(.douta(w_n535_0[0]),.doutb(w_n535_0[1]),.din(n535));
	jspl jspl_w_n536_0(.douta(w_n536_0[0]),.doutb(w_n536_0[1]),.din(n536));
	jspl jspl_w_n537_0(.douta(w_n537_0[0]),.doutb(w_n537_0[1]),.din(n537));
	jspl jspl_w_n538_0(.douta(w_n538_0[0]),.doutb(w_n538_0[1]),.din(n538));
	jspl jspl_w_n539_0(.douta(w_n539_0[0]),.doutb(w_n539_0[1]),.din(n539));
	jspl jspl_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.din(n540));
	jspl jspl_w_n541_0(.douta(w_n541_0[0]),.doutb(w_n541_0[1]),.din(n541));
	jspl jspl_w_n542_0(.douta(w_n542_0[0]),.doutb(w_n542_0[1]),.din(n542));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_n543_0[1]),.din(n543));
	jspl jspl_w_n544_0(.douta(w_n544_0[0]),.doutb(w_n544_0[1]),.din(n544));
	jspl jspl_w_n545_0(.douta(w_n545_0[0]),.doutb(w_n545_0[1]),.din(n545));
	jspl jspl_w_n547_0(.douta(w_n547_0[0]),.doutb(w_n547_0[1]),.din(n547));
	jspl jspl_w_n548_0(.douta(w_n548_0[0]),.doutb(w_n548_0[1]),.din(n548));
	jspl jspl_w_n550_0(.douta(w_dff_A_kbhaqNm07_0),.doutb(w_n550_0[1]),.din(n550));
	jspl jspl_w_n555_0(.douta(w_dff_A_al1351FM3_0),.doutb(w_n555_0[1]),.din(n555));
	jspl jspl_w_n556_0(.douta(w_dff_A_feTdm7cL9_0),.doutb(w_n556_0[1]),.din(n556));
	jspl3 jspl3_w_n561_0(.douta(w_n561_0[0]),.doutb(w_dff_A_GDWe2Ed28_1),.doutc(w_dff_A_pUePyb2f4_2),.din(n561));
	jspl jspl_w_n563_0(.douta(w_n563_0[0]),.doutb(w_n563_0[1]),.din(w_dff_B_v4zCLJrf9_2));
	jspl jspl_w_n566_0(.douta(w_n566_0[0]),.doutb(w_n566_0[1]),.din(n566));
	jspl jspl_w_n568_0(.douta(w_n568_0[0]),.doutb(w_n568_0[1]),.din(w_dff_B_ESOkehGZ8_2));
	jspl jspl_w_n571_0(.douta(w_n571_0[0]),.doutb(w_n571_0[1]),.din(n571));
	jspl jspl_w_n573_0(.douta(w_n573_0[0]),.doutb(w_n573_0[1]),.din(w_dff_B_RwsypYQB6_2));
	jspl jspl_w_n576_0(.douta(w_n576_0[0]),.doutb(w_n576_0[1]),.din(n576));
	jspl jspl_w_n578_0(.douta(w_n578_0[0]),.doutb(w_n578_0[1]),.din(w_dff_B_YeAMfOBG9_2));
	jspl jspl_w_n581_0(.douta(w_n581_0[0]),.doutb(w_n581_0[1]),.din(n581));
	jspl jspl_w_n583_0(.douta(w_n583_0[0]),.doutb(w_n583_0[1]),.din(w_dff_B_CmZh1vkp5_2));
	jspl jspl_w_n586_0(.douta(w_n586_0[0]),.doutb(w_n586_0[1]),.din(n586));
	jspl jspl_w_n588_0(.douta(w_n588_0[0]),.doutb(w_n588_0[1]),.din(w_dff_B_W8fOQmi79_2));
	jspl jspl_w_n591_0(.douta(w_n591_0[0]),.doutb(w_n591_0[1]),.din(n591));
	jspl jspl_w_n593_0(.douta(w_n593_0[0]),.doutb(w_n593_0[1]),.din(w_dff_B_qnHQNVmE9_2));
	jspl jspl_w_n596_0(.douta(w_n596_0[0]),.doutb(w_n596_0[1]),.din(n596));
	jspl jspl_w_n598_0(.douta(w_n598_0[0]),.doutb(w_n598_0[1]),.din(w_dff_B_VWcRMS4Q8_2));
	jspl jspl_w_n602_0(.douta(w_n602_0[0]),.doutb(w_n602_0[1]),.din(n602));
	jspl jspl_w_n603_0(.douta(w_n603_0[0]),.doutb(w_dff_A_G8IX5VBQ3_1),.din(n603));
	jspl jspl_w_n604_0(.douta(w_n604_0[0]),.doutb(w_n604_0[1]),.din(n604));
	jspl jspl_w_n606_0(.douta(w_n606_0[0]),.doutb(w_n606_0[1]),.din(n606));
	jspl3 jspl3_w_n607_0(.douta(w_dff_A_48Fakt9R8_0),.doutb(w_dff_A_1dokVTgx8_1),.doutc(w_n607_0[2]),.din(n607));
	jspl jspl_w_n608_0(.douta(w_n608_0[0]),.doutb(w_n608_0[1]),.din(n608));
	jspl jspl_w_n611_0(.douta(w_dff_A_LStzzifJ6_0),.doutb(w_n611_0[1]),.din(n611));
	jspl jspl_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.din(n613));
	jspl jspl_w_n614_0(.douta(w_n614_0[0]),.doutb(w_n614_0[1]),.din(w_dff_B_myQNXNk33_2));
	jspl jspl_w_n615_0(.douta(w_n615_0[0]),.doutb(w_n615_0[1]),.din(n615));
	jspl jspl_w_n616_0(.douta(w_n616_0[0]),.doutb(w_n616_0[1]),.din(n616));
	jspl jspl_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.din(n617));
	jspl jspl_w_n618_0(.douta(w_n618_0[0]),.doutb(w_n618_0[1]),.din(n618));
	jspl jspl_w_n619_0(.douta(w_n619_0[0]),.doutb(w_n619_0[1]),.din(n619));
	jspl jspl_w_n620_0(.douta(w_n620_0[0]),.doutb(w_n620_0[1]),.din(n620));
	jspl jspl_w_n621_0(.douta(w_n621_0[0]),.doutb(w_n621_0[1]),.din(n621));
	jspl jspl_w_n622_0(.douta(w_n622_0[0]),.doutb(w_n622_0[1]),.din(n622));
	jspl jspl_w_n623_0(.douta(w_n623_0[0]),.doutb(w_n623_0[1]),.din(n623));
	jspl jspl_w_n624_0(.douta(w_n624_0[0]),.doutb(w_n624_0[1]),.din(n624));
	jspl jspl_w_n625_0(.douta(w_n625_0[0]),.doutb(w_n625_0[1]),.din(n625));
	jspl jspl_w_n626_0(.douta(w_n626_0[0]),.doutb(w_n626_0[1]),.din(n626));
	jspl jspl_w_n627_0(.douta(w_n627_0[0]),.doutb(w_n627_0[1]),.din(n627));
	jspl jspl_w_n628_0(.douta(w_n628_0[0]),.doutb(w_n628_0[1]),.din(n628));
	jspl jspl_w_n629_0(.douta(w_n629_0[0]),.doutb(w_n629_0[1]),.din(n629));
	jspl jspl_w_n630_0(.douta(w_n630_0[0]),.doutb(w_n630_0[1]),.din(n630));
	jspl jspl_w_n631_0(.douta(w_n631_0[0]),.doutb(w_n631_0[1]),.din(n631));
	jspl jspl_w_n633_0(.douta(w_n633_0[0]),.doutb(w_n633_0[1]),.din(n633));
	jspl jspl_w_n634_0(.douta(w_n634_0[0]),.doutb(w_n634_0[1]),.din(n634));
	jspl jspl_w_n636_0(.douta(w_dff_A_5SfzQAxg5_0),.doutb(w_n636_0[1]),.din(n636));
	jspl jspl_w_n641_0(.douta(w_dff_A_chNdRabH2_0),.doutb(w_n641_0[1]),.din(n641));
	jspl jspl_w_n642_0(.douta(w_dff_A_5ewLWf1x3_0),.doutb(w_n642_0[1]),.din(n642));
	jspl3 jspl3_w_n647_0(.douta(w_n647_0[0]),.doutb(w_dff_A_aYMwcFEq6_1),.doutc(w_dff_A_LtNAu88Z7_2),.din(n647));
	jspl jspl_w_n649_0(.douta(w_n649_0[0]),.doutb(w_n649_0[1]),.din(w_dff_B_dD5wDP8N1_2));
	jspl jspl_w_n652_0(.douta(w_n652_0[0]),.doutb(w_n652_0[1]),.din(n652));
	jspl jspl_w_n654_0(.douta(w_n654_0[0]),.doutb(w_n654_0[1]),.din(w_dff_B_jZmxLYdm6_2));
	jspl jspl_w_n657_0(.douta(w_n657_0[0]),.doutb(w_n657_0[1]),.din(n657));
	jspl jspl_w_n659_0(.douta(w_n659_0[0]),.doutb(w_n659_0[1]),.din(w_dff_B_VC4cduzu1_2));
	jspl jspl_w_n662_0(.douta(w_n662_0[0]),.doutb(w_n662_0[1]),.din(n662));
	jspl jspl_w_n664_0(.douta(w_n664_0[0]),.doutb(w_n664_0[1]),.din(w_dff_B_wrtKf0bo3_2));
	jspl jspl_w_n667_0(.douta(w_n667_0[0]),.doutb(w_n667_0[1]),.din(n667));
	jspl jspl_w_n669_0(.douta(w_n669_0[0]),.doutb(w_n669_0[1]),.din(w_dff_B_fyCeKIlH9_2));
	jspl jspl_w_n672_0(.douta(w_n672_0[0]),.doutb(w_n672_0[1]),.din(n672));
	jspl jspl_w_n674_0(.douta(w_n674_0[0]),.doutb(w_n674_0[1]),.din(w_dff_B_1cZyvX0q5_2));
	jspl jspl_w_n677_0(.douta(w_n677_0[0]),.doutb(w_n677_0[1]),.din(n677));
	jspl jspl_w_n679_0(.douta(w_n679_0[0]),.doutb(w_n679_0[1]),.din(w_dff_B_fhVItzJa8_2));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.din(n682));
	jspl jspl_w_n684_0(.douta(w_n684_0[0]),.doutb(w_n684_0[1]),.din(w_dff_B_BOKcLPJE6_2));
	jspl jspl_w_n687_0(.douta(w_n687_0[0]),.doutb(w_n687_0[1]),.din(n687));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(w_dff_B_SzG0N2Y24_2));
	jspl jspl_w_n693_0(.douta(w_n693_0[0]),.doutb(w_n693_0[1]),.din(n693));
	jspl jspl_w_n694_0(.douta(w_n694_0[0]),.doutb(w_dff_A_Kcc6bB7L1_1),.din(n694));
	jspl3 jspl3_w_n695_0(.douta(w_dff_A_r6vr8Qko8_0),.doutb(w_n695_0[1]),.doutc(w_n695_0[2]),.din(n695));
	jspl jspl_w_n697_0(.douta(w_n697_0[0]),.doutb(w_n697_0[1]),.din(n697));
	jspl3 jspl3_w_n698_0(.douta(w_dff_A_rwZL9Mh59_0),.doutb(w_dff_A_MD2z5eFk2_1),.doutc(w_n698_0[2]),.din(n698));
	jspl jspl_w_n699_0(.douta(w_n699_0[0]),.doutb(w_n699_0[1]),.din(n699));
	jspl jspl_w_n702_0(.douta(w_dff_A_3m1VZbBZ2_0),.doutb(w_n702_0[1]),.din(n702));
	jspl jspl_w_n704_0(.douta(w_n704_0[0]),.doutb(w_n704_0[1]),.din(n704));
	jspl jspl_w_n705_0(.douta(w_n705_0[0]),.doutb(w_n705_0[1]),.din(w_dff_B_wlQBLVKH0_2));
	jspl jspl_w_n706_0(.douta(w_n706_0[0]),.doutb(w_n706_0[1]),.din(n706));
	jspl jspl_w_n707_0(.douta(w_n707_0[0]),.doutb(w_n707_0[1]),.din(n707));
	jspl jspl_w_n708_0(.douta(w_n708_0[0]),.doutb(w_n708_0[1]),.din(n708));
	jspl jspl_w_n709_0(.douta(w_n709_0[0]),.doutb(w_n709_0[1]),.din(n709));
	jspl jspl_w_n710_0(.douta(w_n710_0[0]),.doutb(w_n710_0[1]),.din(n710));
	jspl jspl_w_n711_0(.douta(w_n711_0[0]),.doutb(w_n711_0[1]),.din(n711));
	jspl jspl_w_n712_0(.douta(w_n712_0[0]),.doutb(w_n712_0[1]),.din(n712));
	jspl jspl_w_n713_0(.douta(w_n713_0[0]),.doutb(w_n713_0[1]),.din(n713));
	jspl jspl_w_n714_0(.douta(w_n714_0[0]),.doutb(w_n714_0[1]),.din(n714));
	jspl jspl_w_n715_0(.douta(w_n715_0[0]),.doutb(w_n715_0[1]),.din(n715));
	jspl jspl_w_n716_0(.douta(w_n716_0[0]),.doutb(w_n716_0[1]),.din(n716));
	jspl jspl_w_n717_0(.douta(w_n717_0[0]),.doutb(w_n717_0[1]),.din(n717));
	jspl jspl_w_n718_0(.douta(w_n718_0[0]),.doutb(w_n718_0[1]),.din(n718));
	jspl jspl_w_n719_0(.douta(w_n719_0[0]),.doutb(w_n719_0[1]),.din(n719));
	jspl jspl_w_n720_0(.douta(w_n720_0[0]),.doutb(w_n720_0[1]),.din(n720));
	jspl jspl_w_n721_0(.douta(w_n721_0[0]),.doutb(w_n721_0[1]),.din(n721));
	jspl jspl_w_n722_0(.douta(w_n722_0[0]),.doutb(w_n722_0[1]),.din(n722));
	jspl jspl_w_n723_0(.douta(w_n723_0[0]),.doutb(w_n723_0[1]),.din(n723));
	jspl jspl_w_n724_0(.douta(w_n724_0[0]),.doutb(w_n724_0[1]),.din(n724));
	jspl jspl_w_n726_0(.douta(w_n726_0[0]),.doutb(w_n726_0[1]),.din(n726));
	jspl jspl_w_n727_0(.douta(w_n727_0[0]),.doutb(w_n727_0[1]),.din(n727));
	jspl jspl_w_n729_0(.douta(w_dff_A_1NxHfHhh4_0),.doutb(w_n729_0[1]),.din(n729));
	jspl jspl_w_n734_0(.douta(w_dff_A_QRIEawwW9_0),.doutb(w_n734_0[1]),.din(n734));
	jspl jspl_w_n735_0(.douta(w_dff_A_ll4vw5e71_0),.doutb(w_n735_0[1]),.din(n735));
	jspl3 jspl3_w_n740_0(.douta(w_n740_0[0]),.doutb(w_dff_A_ISoQoaIJ1_1),.doutc(w_dff_A_kazzux2u8_2),.din(n740));
	jspl jspl_w_n742_0(.douta(w_n742_0[0]),.doutb(w_n742_0[1]),.din(w_dff_B_6zgCuI5N9_2));
	jspl jspl_w_n745_0(.douta(w_n745_0[0]),.doutb(w_n745_0[1]),.din(n745));
	jspl jspl_w_n747_0(.douta(w_n747_0[0]),.doutb(w_n747_0[1]),.din(w_dff_B_Ge66VRId2_2));
	jspl jspl_w_n750_0(.douta(w_n750_0[0]),.doutb(w_n750_0[1]),.din(n750));
	jspl jspl_w_n752_0(.douta(w_n752_0[0]),.doutb(w_n752_0[1]),.din(w_dff_B_G0y1hWVS6_2));
	jspl jspl_w_n755_0(.douta(w_n755_0[0]),.doutb(w_n755_0[1]),.din(n755));
	jspl jspl_w_n757_0(.douta(w_n757_0[0]),.doutb(w_n757_0[1]),.din(w_dff_B_tWkl39uc5_2));
	jspl jspl_w_n760_0(.douta(w_n760_0[0]),.doutb(w_n760_0[1]),.din(n760));
	jspl jspl_w_n762_0(.douta(w_n762_0[0]),.doutb(w_n762_0[1]),.din(w_dff_B_531w516D6_2));
	jspl jspl_w_n765_0(.douta(w_n765_0[0]),.doutb(w_n765_0[1]),.din(n765));
	jspl jspl_w_n767_0(.douta(w_n767_0[0]),.doutb(w_n767_0[1]),.din(w_dff_B_1303sco78_2));
	jspl jspl_w_n770_0(.douta(w_n770_0[0]),.doutb(w_n770_0[1]),.din(n770));
	jspl jspl_w_n772_0(.douta(w_n772_0[0]),.doutb(w_n772_0[1]),.din(w_dff_B_GRLdMi0n6_2));
	jspl jspl_w_n775_0(.douta(w_n775_0[0]),.doutb(w_n775_0[1]),.din(n775));
	jspl jspl_w_n777_0(.douta(w_n777_0[0]),.doutb(w_n777_0[1]),.din(w_dff_B_aUyLW4GW0_2));
	jspl jspl_w_n780_0(.douta(w_n780_0[0]),.doutb(w_n780_0[1]),.din(n780));
	jspl jspl_w_n782_0(.douta(w_n782_0[0]),.doutb(w_n782_0[1]),.din(w_dff_B_IYyZof909_2));
	jspl jspl_w_n785_0(.douta(w_n785_0[0]),.doutb(w_n785_0[1]),.din(n785));
	jspl jspl_w_n787_0(.douta(w_n787_0[0]),.doutb(w_n787_0[1]),.din(w_dff_B_zeb0jvwG4_2));
	jspl jspl_w_n791_0(.douta(w_n791_0[0]),.doutb(w_n791_0[1]),.din(n791));
	jspl jspl_w_n792_0(.douta(w_n792_0[0]),.doutb(w_dff_A_5nlEOUCZ1_1),.din(n792));
	jspl jspl_w_n793_0(.douta(w_dff_A_be4tAm5B8_0),.doutb(w_n793_0[1]),.din(n793));
	jspl jspl_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.din(n795));
	jspl3 jspl3_w_n797_0(.douta(w_n797_0[0]),.doutb(w_n797_0[1]),.doutc(w_n797_0[2]),.din(n797));
	jspl jspl_w_n800_0(.douta(w_dff_A_BmmRQH6Y3_0),.doutb(w_n800_0[1]),.din(n800));
	jspl jspl_w_n802_0(.douta(w_n802_0[0]),.doutb(w_n802_0[1]),.din(n802));
	jspl jspl_w_n803_0(.douta(w_n803_0[0]),.doutb(w_n803_0[1]),.din(w_dff_B_GAMWtoFq2_2));
	jspl jspl_w_n804_0(.douta(w_n804_0[0]),.doutb(w_n804_0[1]),.din(n804));
	jspl jspl_w_n805_0(.douta(w_n805_0[0]),.doutb(w_n805_0[1]),.din(n805));
	jspl jspl_w_n806_0(.douta(w_n806_0[0]),.doutb(w_n806_0[1]),.din(n806));
	jspl jspl_w_n807_0(.douta(w_n807_0[0]),.doutb(w_n807_0[1]),.din(n807));
	jspl jspl_w_n808_0(.douta(w_n808_0[0]),.doutb(w_n808_0[1]),.din(n808));
	jspl jspl_w_n809_0(.douta(w_n809_0[0]),.doutb(w_n809_0[1]),.din(n809));
	jspl jspl_w_n810_0(.douta(w_n810_0[0]),.doutb(w_n810_0[1]),.din(n810));
	jspl jspl_w_n811_0(.douta(w_n811_0[0]),.doutb(w_n811_0[1]),.din(n811));
	jspl jspl_w_n812_0(.douta(w_n812_0[0]),.doutb(w_n812_0[1]),.din(n812));
	jspl jspl_w_n813_0(.douta(w_n813_0[0]),.doutb(w_n813_0[1]),.din(n813));
	jspl jspl_w_n814_0(.douta(w_n814_0[0]),.doutb(w_n814_0[1]),.din(n814));
	jspl jspl_w_n815_0(.douta(w_n815_0[0]),.doutb(w_n815_0[1]),.din(n815));
	jspl jspl_w_n816_0(.douta(w_n816_0[0]),.doutb(w_n816_0[1]),.din(n816));
	jspl jspl_w_n817_0(.douta(w_n817_0[0]),.doutb(w_n817_0[1]),.din(n817));
	jspl jspl_w_n818_0(.douta(w_n818_0[0]),.doutb(w_n818_0[1]),.din(n818));
	jspl jspl_w_n819_0(.douta(w_n819_0[0]),.doutb(w_n819_0[1]),.din(n819));
	jspl jspl_w_n820_0(.douta(w_n820_0[0]),.doutb(w_n820_0[1]),.din(n820));
	jspl jspl_w_n821_0(.douta(w_n821_0[0]),.doutb(w_n821_0[1]),.din(n821));
	jspl jspl_w_n822_0(.douta(w_n822_0[0]),.doutb(w_n822_0[1]),.din(n822));
	jspl jspl_w_n823_0(.douta(w_n823_0[0]),.doutb(w_n823_0[1]),.din(n823));
	jspl jspl_w_n824_0(.douta(w_n824_0[0]),.doutb(w_n824_0[1]),.din(n824));
	jspl jspl_w_n826_0(.douta(w_n826_0[0]),.doutb(w_n826_0[1]),.din(n826));
	jspl jspl_w_n827_0(.douta(w_n827_0[0]),.doutb(w_n827_0[1]),.din(n827));
	jspl jspl_w_n829_0(.douta(w_dff_A_IEtz1gEB5_0),.doutb(w_n829_0[1]),.din(n829));
	jspl jspl_w_n834_0(.douta(w_n834_0[0]),.doutb(w_n834_0[1]),.din(n834));
	jspl jspl_w_n835_0(.douta(w_n835_0[0]),.doutb(w_n835_0[1]),.din(w_dff_B_ik6tOIxU0_2));
	jspl jspl_w_n839_0(.douta(w_dff_A_13aE2Vnd9_0),.doutb(w_n839_0[1]),.din(n839));
	jspl jspl_w_n840_0(.douta(w_dff_A_CO6oBVJP9_0),.doutb(w_n840_0[1]),.din(n840));
	jspl3 jspl3_w_n844_0(.douta(w_dff_A_qN6gSYM48_0),.doutb(w_n844_0[1]),.doutc(w_n844_0[2]),.din(n844));
	jspl jspl_w_n846_0(.douta(w_n846_0[0]),.doutb(w_n846_0[1]),.din(w_dff_B_32BBUETR6_2));
	jspl jspl_w_n849_0(.douta(w_n849_0[0]),.doutb(w_n849_0[1]),.din(n849));
	jspl jspl_w_n851_0(.douta(w_n851_0[0]),.doutb(w_n851_0[1]),.din(w_dff_B_JClOxoUf1_2));
	jspl jspl_w_n854_0(.douta(w_n854_0[0]),.doutb(w_n854_0[1]),.din(n854));
	jspl jspl_w_n856_0(.douta(w_n856_0[0]),.doutb(w_n856_0[1]),.din(w_dff_B_i3mTkYqK7_2));
	jspl jspl_w_n859_0(.douta(w_n859_0[0]),.doutb(w_n859_0[1]),.din(n859));
	jspl jspl_w_n861_0(.douta(w_n861_0[0]),.doutb(w_n861_0[1]),.din(w_dff_B_BMw3Lxb49_2));
	jspl jspl_w_n864_0(.douta(w_n864_0[0]),.doutb(w_n864_0[1]),.din(n864));
	jspl jspl_w_n866_0(.douta(w_n866_0[0]),.doutb(w_n866_0[1]),.din(w_dff_B_jPnbXJoN6_2));
	jspl jspl_w_n869_0(.douta(w_n869_0[0]),.doutb(w_n869_0[1]),.din(n869));
	jspl jspl_w_n871_0(.douta(w_n871_0[0]),.doutb(w_n871_0[1]),.din(w_dff_B_ohS8euDz2_2));
	jspl jspl_w_n874_0(.douta(w_n874_0[0]),.doutb(w_n874_0[1]),.din(n874));
	jspl jspl_w_n876_0(.douta(w_n876_0[0]),.doutb(w_n876_0[1]),.din(w_dff_B_bPAnp4Pw3_2));
	jspl jspl_w_n879_0(.douta(w_n879_0[0]),.doutb(w_n879_0[1]),.din(n879));
	jspl jspl_w_n881_0(.douta(w_n881_0[0]),.doutb(w_n881_0[1]),.din(w_dff_B_6PAKBTgy5_2));
	jspl jspl_w_n884_0(.douta(w_n884_0[0]),.doutb(w_n884_0[1]),.din(n884));
	jspl jspl_w_n886_0(.douta(w_n886_0[0]),.doutb(w_n886_0[1]),.din(w_dff_B_Zhi0614O5_2));
	jspl jspl_w_n889_0(.douta(w_n889_0[0]),.doutb(w_n889_0[1]),.din(n889));
	jspl jspl_w_n891_0(.douta(w_n891_0[0]),.doutb(w_n891_0[1]),.din(w_dff_B_hzNvwo292_2));
	jspl jspl_w_n895_0(.douta(w_n895_0[0]),.doutb(w_n895_0[1]),.din(n895));
	jspl jspl_w_n896_0(.douta(w_n896_0[0]),.doutb(w_dff_A_WQZtJbXd3_1),.din(n896));
	jspl jspl_w_n897_0(.douta(w_n897_0[0]),.doutb(w_n897_0[1]),.din(n897));
	jspl jspl_w_n898_0(.douta(w_n898_0[0]),.doutb(w_n898_0[1]),.din(w_dff_B_PZUfM55S1_2));
	jspl jspl_w_n901_0(.douta(w_n901_0[0]),.doutb(w_dff_A_6V0MbwZf0_1),.din(n901));
	jspl jspl_w_n903_0(.douta(w_dff_A_zLgoNo255_0),.doutb(w_n903_0[1]),.din(n903));
	jspl jspl_w_n906_0(.douta(w_n906_0[0]),.doutb(w_n906_0[1]),.din(n906));
	jspl jspl_w_n907_0(.douta(w_n907_0[0]),.doutb(w_n907_0[1]),.din(w_dff_B_E2ffu9kh8_2));
	jspl jspl_w_n908_0(.douta(w_n908_0[0]),.doutb(w_n908_0[1]),.din(n908));
	jspl jspl_w_n909_0(.douta(w_n909_0[0]),.doutb(w_n909_0[1]),.din(n909));
	jspl jspl_w_n910_0(.douta(w_n910_0[0]),.doutb(w_n910_0[1]),.din(n910));
	jspl jspl_w_n911_0(.douta(w_n911_0[0]),.doutb(w_n911_0[1]),.din(n911));
	jspl jspl_w_n912_0(.douta(w_n912_0[0]),.doutb(w_n912_0[1]),.din(n912));
	jspl jspl_w_n913_0(.douta(w_n913_0[0]),.doutb(w_n913_0[1]),.din(n913));
	jspl jspl_w_n914_0(.douta(w_n914_0[0]),.doutb(w_n914_0[1]),.din(n914));
	jspl jspl_w_n915_0(.douta(w_n915_0[0]),.doutb(w_n915_0[1]),.din(n915));
	jspl jspl_w_n916_0(.douta(w_n916_0[0]),.doutb(w_n916_0[1]),.din(n916));
	jspl jspl_w_n917_0(.douta(w_n917_0[0]),.doutb(w_n917_0[1]),.din(n917));
	jspl jspl_w_n918_0(.douta(w_n918_0[0]),.doutb(w_n918_0[1]),.din(n918));
	jspl jspl_w_n919_0(.douta(w_n919_0[0]),.doutb(w_n919_0[1]),.din(n919));
	jspl jspl_w_n920_0(.douta(w_n920_0[0]),.doutb(w_n920_0[1]),.din(n920));
	jspl jspl_w_n921_0(.douta(w_n921_0[0]),.doutb(w_n921_0[1]),.din(n921));
	jspl jspl_w_n922_0(.douta(w_n922_0[0]),.doutb(w_n922_0[1]),.din(n922));
	jspl jspl_w_n923_0(.douta(w_n923_0[0]),.doutb(w_n923_0[1]),.din(n923));
	jspl jspl_w_n924_0(.douta(w_n924_0[0]),.doutb(w_n924_0[1]),.din(n924));
	jspl jspl_w_n925_0(.douta(w_n925_0[0]),.doutb(w_n925_0[1]),.din(n925));
	jspl jspl_w_n926_0(.douta(w_n926_0[0]),.doutb(w_n926_0[1]),.din(n926));
	jspl3 jspl3_w_n927_0(.douta(w_n927_0[0]),.doutb(w_n927_0[1]),.doutc(w_n927_0[2]),.din(n927));
	jspl jspl_w_n929_0(.douta(w_n929_0[0]),.doutb(w_n929_0[1]),.din(n929));
	jspl jspl_w_n930_0(.douta(w_n930_0[0]),.doutb(w_n930_0[1]),.din(n930));
	jspl jspl_w_n931_0(.douta(w_n931_0[0]),.doutb(w_dff_A_0sPTpbU60_1),.din(n931));
	jspl jspl_w_n932_0(.douta(w_n932_0[0]),.doutb(w_n932_0[1]),.din(n932));
	jspl jspl_w_n937_0(.douta(w_n937_0[0]),.doutb(w_n937_0[1]),.din(w_dff_B_GAtqHJmd0_2));
	jspl jspl_w_n938_0(.douta(w_n938_0[0]),.doutb(w_dff_A_JALddgvv6_1),.din(w_dff_B_kWfNUNAt5_2));
	jspl3 jspl3_w_n942_0(.douta(w_n942_0[0]),.doutb(w_dff_A_i1clNZ0m9_1),.doutc(w_dff_A_um8ltIX04_2),.din(w_dff_B_kLnAW15u8_3));
	jspl jspl_w_n943_0(.douta(w_n943_0[0]),.doutb(w_n943_0[1]),.din(w_dff_B_l8C2ByAj2_2));
	jspl jspl_w_n949_0(.douta(w_n949_0[0]),.doutb(w_n949_0[1]),.din(n949));
	jspl jspl_w_n951_0(.douta(w_n951_0[0]),.doutb(w_n951_0[1]),.din(w_dff_B_yoJ1bUnw9_2));
	jspl jspl_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.din(n954));
	jspl jspl_w_n956_0(.douta(w_n956_0[0]),.doutb(w_n956_0[1]),.din(w_dff_B_0ZoEKReq9_2));
	jspl jspl_w_n959_0(.douta(w_n959_0[0]),.doutb(w_n959_0[1]),.din(n959));
	jspl jspl_w_n961_0(.douta(w_n961_0[0]),.doutb(w_n961_0[1]),.din(w_dff_B_DHkkivkZ8_2));
	jspl jspl_w_n964_0(.douta(w_n964_0[0]),.doutb(w_n964_0[1]),.din(n964));
	jspl jspl_w_n966_0(.douta(w_n966_0[0]),.doutb(w_n966_0[1]),.din(w_dff_B_6TEB4FEv0_2));
	jspl jspl_w_n969_0(.douta(w_n969_0[0]),.doutb(w_n969_0[1]),.din(n969));
	jspl jspl_w_n971_0(.douta(w_n971_0[0]),.doutb(w_n971_0[1]),.din(w_dff_B_yGnZ6wXe5_2));
	jspl jspl_w_n974_0(.douta(w_n974_0[0]),.doutb(w_n974_0[1]),.din(n974));
	jspl jspl_w_n976_0(.douta(w_n976_0[0]),.doutb(w_n976_0[1]),.din(w_dff_B_DCbt8AsM8_2));
	jspl jspl_w_n979_0(.douta(w_n979_0[0]),.doutb(w_n979_0[1]),.din(n979));
	jspl jspl_w_n981_0(.douta(w_n981_0[0]),.doutb(w_n981_0[1]),.din(w_dff_B_QM2ywPH17_2));
	jspl jspl_w_n984_0(.douta(w_n984_0[0]),.doutb(w_n984_0[1]),.din(n984));
	jspl jspl_w_n986_0(.douta(w_n986_0[0]),.doutb(w_n986_0[1]),.din(w_dff_B_6akHVQl14_2));
	jspl jspl_w_n989_0(.douta(w_n989_0[0]),.doutb(w_n989_0[1]),.din(n989));
	jspl jspl_w_n991_0(.douta(w_n991_0[0]),.doutb(w_n991_0[1]),.din(w_dff_B_06ARLHTF0_2));
	jspl jspl_w_n994_0(.douta(w_n994_0[0]),.doutb(w_n994_0[1]),.din(n994));
	jspl jspl_w_n996_0(.douta(w_n996_0[0]),.doutb(w_n996_0[1]),.din(w_dff_B_ixfXDMSX9_2));
	jspl jspl_w_n999_0(.douta(w_n999_0[0]),.doutb(w_n999_0[1]),.din(n999));
	jspl jspl_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.din(w_dff_B_ImuegOsW8_2));
	jspl jspl_w_n1005_0(.douta(w_n1005_0[0]),.doutb(w_n1005_0[1]),.din(n1005));
	jspl jspl_w_n1006_0(.douta(w_n1006_0[0]),.doutb(w_dff_A_oqTUZVoI6_1),.din(n1006));
	jspl jspl_w_n1008_0(.douta(w_dff_A_CBBvRGVn6_0),.doutb(w_n1008_0[1]),.din(n1008));
	jspl jspl_w_n1009_0(.douta(w_n1009_0[0]),.doutb(w_n1009_0[1]),.din(n1009));
	jspl jspl_w_n1010_0(.douta(w_n1010_0[0]),.doutb(w_n1010_0[1]),.din(w_dff_B_RUO3PTNq1_2));
	jspl jspl_w_n1011_0(.douta(w_n1011_0[0]),.doutb(w_n1011_0[1]),.din(n1011));
	jspl jspl_w_n1012_0(.douta(w_n1012_0[0]),.doutb(w_n1012_0[1]),.din(n1012));
	jspl jspl_w_n1013_0(.douta(w_n1013_0[0]),.doutb(w_n1013_0[1]),.din(n1013));
	jspl jspl_w_n1014_0(.douta(w_n1014_0[0]),.doutb(w_n1014_0[1]),.din(n1014));
	jspl jspl_w_n1015_0(.douta(w_n1015_0[0]),.doutb(w_n1015_0[1]),.din(n1015));
	jspl jspl_w_n1016_0(.douta(w_n1016_0[0]),.doutb(w_n1016_0[1]),.din(n1016));
	jspl jspl_w_n1017_0(.douta(w_n1017_0[0]),.doutb(w_n1017_0[1]),.din(n1017));
	jspl jspl_w_n1018_0(.douta(w_n1018_0[0]),.doutb(w_n1018_0[1]),.din(n1018));
	jspl jspl_w_n1019_0(.douta(w_n1019_0[0]),.doutb(w_n1019_0[1]),.din(n1019));
	jspl jspl_w_n1020_0(.douta(w_n1020_0[0]),.doutb(w_n1020_0[1]),.din(n1020));
	jspl jspl_w_n1021_0(.douta(w_n1021_0[0]),.doutb(w_n1021_0[1]),.din(n1021));
	jspl jspl_w_n1022_0(.douta(w_n1022_0[0]),.doutb(w_n1022_0[1]),.din(n1022));
	jspl jspl_w_n1023_0(.douta(w_n1023_0[0]),.doutb(w_n1023_0[1]),.din(n1023));
	jspl jspl_w_n1024_0(.douta(w_n1024_0[0]),.doutb(w_n1024_0[1]),.din(n1024));
	jspl jspl_w_n1025_0(.douta(w_n1025_0[0]),.doutb(w_n1025_0[1]),.din(n1025));
	jspl jspl_w_n1026_0(.douta(w_n1026_0[0]),.doutb(w_n1026_0[1]),.din(n1026));
	jspl jspl_w_n1027_0(.douta(w_n1027_0[0]),.doutb(w_n1027_0[1]),.din(n1027));
	jspl jspl_w_n1028_0(.douta(w_n1028_0[0]),.doutb(w_n1028_0[1]),.din(n1028));
	jspl jspl_w_n1029_0(.douta(w_n1029_0[0]),.doutb(w_n1029_0[1]),.din(n1029));
	jspl jspl_w_n1030_0(.douta(w_n1030_0[0]),.doutb(w_n1030_0[1]),.din(n1030));
	jspl jspl_w_n1031_0(.douta(w_n1031_0[0]),.doutb(w_n1031_0[1]),.din(n1031));
	jspl jspl_w_n1032_0(.douta(w_n1032_0[0]),.doutb(w_dff_A_qzgPrtGO7_1),.din(n1032));
	jspl jspl_w_n1033_0(.douta(w_n1033_0[0]),.doutb(w_n1033_0[1]),.din(n1033));
	jspl jspl_w_n1034_0(.douta(w_n1034_0[0]),.doutb(w_n1034_0[1]),.din(n1034));
	jspl jspl_w_n1035_0(.douta(w_n1035_0[0]),.doutb(w_n1035_0[1]),.din(n1035));
	jspl jspl_w_n1037_0(.douta(w_n1037_0[0]),.doutb(w_n1037_0[1]),.din(n1037));
	jspl jspl_w_n1039_0(.douta(w_n1039_0[0]),.doutb(w_dff_A_QGWkux4p1_1),.din(n1039));
	jspl jspl_w_n1043_0(.douta(w_dff_A_iW07Qgb02_0),.doutb(w_n1043_0[1]),.din(w_dff_B_siiwXJJ18_2));
	jspl jspl_w_n1044_0(.douta(w_n1044_0[0]),.doutb(w_n1044_0[1]),.din(w_dff_B_etIzj5896_2));
	jspl jspl_w_n1048_0(.douta(w_dff_A_rMaboMKD7_0),.doutb(w_n1048_0[1]),.din(w_dff_B_ZcdfPDIP9_2));
	jspl jspl_w_n1049_0(.douta(w_n1049_0[0]),.doutb(w_n1049_0[1]),.din(w_dff_B_0Y6pU22K5_2));
	jspl jspl_w_n1052_0(.douta(w_n1052_0[0]),.doutb(w_n1052_0[1]),.din(w_dff_B_5BmTqeRt2_2));
	jspl jspl_w_n1054_0(.douta(w_n1054_0[0]),.doutb(w_n1054_0[1]),.din(w_dff_B_Hh2EdLSE0_2));
	jspl jspl_w_n1057_0(.douta(w_n1057_0[0]),.doutb(w_n1057_0[1]),.din(w_dff_B_69xcZT3g0_2));
	jspl jspl_w_n1059_0(.douta(w_n1059_0[0]),.doutb(w_n1059_0[1]),.din(w_dff_B_3wbRcmS09_2));
	jspl jspl_w_n1062_0(.douta(w_n1062_0[0]),.doutb(w_n1062_0[1]),.din(w_dff_B_ifC4YSHr9_2));
	jspl jspl_w_n1064_0(.douta(w_n1064_0[0]),.doutb(w_n1064_0[1]),.din(w_dff_B_gIN7GL8I4_2));
	jspl jspl_w_n1067_0(.douta(w_n1067_0[0]),.doutb(w_n1067_0[1]),.din(w_dff_B_Vk4Qj9aA2_2));
	jspl jspl_w_n1069_0(.douta(w_n1069_0[0]),.doutb(w_n1069_0[1]),.din(w_dff_B_jLbPvk7S3_2));
	jspl jspl_w_n1072_0(.douta(w_n1072_0[0]),.doutb(w_n1072_0[1]),.din(w_dff_B_PT0HtWut8_2));
	jspl jspl_w_n1074_0(.douta(w_n1074_0[0]),.doutb(w_n1074_0[1]),.din(w_dff_B_PrzCxOEQ4_2));
	jspl jspl_w_n1077_0(.douta(w_n1077_0[0]),.doutb(w_n1077_0[1]),.din(w_dff_B_JSHBTzFy4_2));
	jspl jspl_w_n1079_0(.douta(w_n1079_0[0]),.doutb(w_n1079_0[1]),.din(w_dff_B_uRS1Fs5X4_2));
	jspl jspl_w_n1082_0(.douta(w_n1082_0[0]),.doutb(w_n1082_0[1]),.din(w_dff_B_q9ZmF9Nl0_2));
	jspl jspl_w_n1084_0(.douta(w_n1084_0[0]),.doutb(w_n1084_0[1]),.din(w_dff_B_y3BcU3Is6_2));
	jspl jspl_w_n1087_0(.douta(w_n1087_0[0]),.doutb(w_n1087_0[1]),.din(w_dff_B_575PgbKq3_2));
	jspl jspl_w_n1089_0(.douta(w_n1089_0[0]),.doutb(w_n1089_0[1]),.din(w_dff_B_4efL7dCV5_2));
	jspl jspl_w_n1092_0(.douta(w_n1092_0[0]),.doutb(w_n1092_0[1]),.din(w_dff_B_HU2GbyaZ7_2));
	jspl jspl_w_n1094_0(.douta(w_n1094_0[0]),.doutb(w_n1094_0[1]),.din(w_dff_B_dnvH4RRW9_2));
	jspl jspl_w_n1097_0(.douta(w_n1097_0[0]),.doutb(w_n1097_0[1]),.din(w_dff_B_bqJrps8C6_2));
	jspl jspl_w_n1099_0(.douta(w_n1099_0[0]),.doutb(w_n1099_0[1]),.din(w_dff_B_tmJgp1tV3_2));
	jspl jspl_w_n1102_0(.douta(w_n1102_0[0]),.doutb(w_n1102_0[1]),.din(w_dff_B_8Y9hUj1G5_2));
	jspl jspl_w_n1103_0(.douta(w_n1103_0[0]),.doutb(w_n1103_0[1]),.din(w_dff_B_Rw9ReYqf4_2));
	jspl jspl_w_n1109_0(.douta(w_n1109_0[0]),.doutb(w_n1109_0[1]),.din(n1109));
	jspl jspl_w_n1110_0(.douta(w_dff_A_vg1N7GSx6_0),.doutb(w_n1110_0[1]),.din(w_dff_B_LsD0lV718_2));
	jspl jspl_w_n1114_0(.douta(w_n1114_0[0]),.doutb(w_n1114_0[1]),.din(n1114));
	jspl jspl_w_n1115_0(.douta(w_n1115_0[0]),.doutb(w_n1115_0[1]),.din(n1115));
	jspl jspl_w_n1116_0(.douta(w_n1116_0[0]),.doutb(w_n1116_0[1]),.din(n1116));
	jspl jspl_w_n1117_0(.douta(w_n1117_0[0]),.doutb(w_n1117_0[1]),.din(n1117));
	jspl jspl_w_n1118_0(.douta(w_n1118_0[0]),.doutb(w_n1118_0[1]),.din(n1118));
	jspl jspl_w_n1119_0(.douta(w_n1119_0[0]),.doutb(w_n1119_0[1]),.din(n1119));
	jspl jspl_w_n1120_0(.douta(w_n1120_0[0]),.doutb(w_n1120_0[1]),.din(n1120));
	jspl jspl_w_n1121_0(.douta(w_n1121_0[0]),.doutb(w_n1121_0[1]),.din(n1121));
	jspl jspl_w_n1122_0(.douta(w_n1122_0[0]),.doutb(w_n1122_0[1]),.din(n1122));
	jspl jspl_w_n1123_0(.douta(w_n1123_0[0]),.doutb(w_n1123_0[1]),.din(n1123));
	jspl jspl_w_n1124_0(.douta(w_n1124_0[0]),.doutb(w_n1124_0[1]),.din(n1124));
	jspl jspl_w_n1125_0(.douta(w_n1125_0[0]),.doutb(w_n1125_0[1]),.din(n1125));
	jspl jspl_w_n1126_0(.douta(w_n1126_0[0]),.doutb(w_n1126_0[1]),.din(n1126));
	jspl jspl_w_n1127_0(.douta(w_n1127_0[0]),.doutb(w_n1127_0[1]),.din(n1127));
	jspl jspl_w_n1128_0(.douta(w_n1128_0[0]),.doutb(w_n1128_0[1]),.din(n1128));
	jspl jspl_w_n1129_0(.douta(w_n1129_0[0]),.doutb(w_n1129_0[1]),.din(n1129));
	jspl jspl_w_n1130_0(.douta(w_n1130_0[0]),.doutb(w_n1130_0[1]),.din(n1130));
	jspl jspl_w_n1131_0(.douta(w_n1131_0[0]),.doutb(w_n1131_0[1]),.din(n1131));
	jspl jspl_w_n1132_0(.douta(w_n1132_0[0]),.doutb(w_n1132_0[1]),.din(n1132));
	jspl jspl_w_n1133_0(.douta(w_n1133_0[0]),.doutb(w_n1133_0[1]),.din(n1133));
	jspl jspl_w_n1134_0(.douta(w_n1134_0[0]),.doutb(w_n1134_0[1]),.din(n1134));
	jspl jspl_w_n1135_0(.douta(w_n1135_0[0]),.doutb(w_n1135_0[1]),.din(n1135));
	jspl jspl_w_n1137_0(.douta(w_n1137_0[0]),.doutb(w_n1137_0[1]),.din(n1137));
	jspl jspl_w_n1138_0(.douta(w_n1138_0[0]),.doutb(w_n1138_0[1]),.din(n1138));
	jspl jspl_w_n1139_0(.douta(w_n1139_0[0]),.doutb(w_n1139_0[1]),.din(n1139));
	jspl jspl_w_n1140_0(.douta(w_n1140_0[0]),.doutb(w_n1140_0[1]),.din(n1140));
	jspl jspl_w_n1141_0(.douta(w_n1141_0[0]),.doutb(w_n1141_0[1]),.din(n1141));
	jspl jspl_w_n1147_0(.douta(w_n1147_0[0]),.doutb(w_dff_A_7yfYQd7z3_1),.din(w_dff_B_7mxns7If6_2));
	jspl jspl_w_n1151_0(.douta(w_dff_A_2RGpeNmG4_0),.doutb(w_n1151_0[1]),.din(w_dff_B_bYJNWGcp4_2));
	jspl jspl_w_n1152_0(.douta(w_n1152_0[0]),.doutb(w_n1152_0[1]),.din(w_dff_B_dkaftnOp3_2));
	jspl jspl_w_n1156_0(.douta(w_n1156_0[0]),.doutb(w_n1156_0[1]),.din(w_dff_B_HDeeE3zj8_2));
	jspl jspl_w_n1158_0(.douta(w_n1158_0[0]),.doutb(w_n1158_0[1]),.din(w_dff_B_VjKKWoOF8_2));
	jspl jspl_w_n1161_0(.douta(w_n1161_0[0]),.doutb(w_n1161_0[1]),.din(w_dff_B_43rU9oyq8_2));
	jspl jspl_w_n1163_0(.douta(w_n1163_0[0]),.doutb(w_n1163_0[1]),.din(w_dff_B_0gddxcGe8_2));
	jspl jspl_w_n1166_0(.douta(w_n1166_0[0]),.doutb(w_n1166_0[1]),.din(w_dff_B_NZTEQUB73_2));
	jspl jspl_w_n1168_0(.douta(w_n1168_0[0]),.doutb(w_n1168_0[1]),.din(w_dff_B_BeKR35A02_2));
	jspl jspl_w_n1171_0(.douta(w_n1171_0[0]),.doutb(w_n1171_0[1]),.din(w_dff_B_xl0I0JEE5_2));
	jspl jspl_w_n1173_0(.douta(w_n1173_0[0]),.doutb(w_n1173_0[1]),.din(w_dff_B_mmbLPHoG8_2));
	jspl jspl_w_n1176_0(.douta(w_n1176_0[0]),.doutb(w_n1176_0[1]),.din(w_dff_B_kZA6OXJq2_2));
	jspl jspl_w_n1178_0(.douta(w_n1178_0[0]),.doutb(w_n1178_0[1]),.din(w_dff_B_qM3TMyS62_2));
	jspl jspl_w_n1181_0(.douta(w_n1181_0[0]),.doutb(w_n1181_0[1]),.din(w_dff_B_eLwyZtca5_2));
	jspl jspl_w_n1183_0(.douta(w_n1183_0[0]),.doutb(w_n1183_0[1]),.din(w_dff_B_pdMKyQz74_2));
	jspl jspl_w_n1186_0(.douta(w_n1186_0[0]),.doutb(w_n1186_0[1]),.din(w_dff_B_4s9CXQls9_2));
	jspl jspl_w_n1188_0(.douta(w_n1188_0[0]),.doutb(w_n1188_0[1]),.din(w_dff_B_EuRzVPuY5_2));
	jspl jspl_w_n1191_0(.douta(w_n1191_0[0]),.doutb(w_n1191_0[1]),.din(w_dff_B_s1neHrrM3_2));
	jspl jspl_w_n1193_0(.douta(w_n1193_0[0]),.doutb(w_n1193_0[1]),.din(w_dff_B_ai4SvB5g3_2));
	jspl jspl_w_n1196_0(.douta(w_n1196_0[0]),.doutb(w_n1196_0[1]),.din(w_dff_B_Nz2nYbTU5_2));
	jspl jspl_w_n1198_0(.douta(w_n1198_0[0]),.doutb(w_n1198_0[1]),.din(w_dff_B_fCsW9NnO7_2));
	jspl jspl_w_n1201_0(.douta(w_n1201_0[0]),.doutb(w_n1201_0[1]),.din(w_dff_B_xUKLDhg11_2));
	jspl jspl_w_n1203_0(.douta(w_n1203_0[0]),.doutb(w_n1203_0[1]),.din(w_dff_B_eGtqjqZM3_2));
	jspl jspl_w_n1206_0(.douta(w_n1206_0[0]),.doutb(w_n1206_0[1]),.din(w_dff_B_qtCwMmqV7_2));
	jspl jspl_w_n1207_0(.douta(w_n1207_0[0]),.doutb(w_n1207_0[1]),.din(w_dff_B_PtBSenI71_2));
	jspl jspl_w_n1208_0(.douta(w_n1208_0[0]),.doutb(w_n1208_0[1]),.din(w_dff_B_v33DHjVQ4_2));
	jspl jspl_w_n1210_0(.douta(w_n1210_0[0]),.doutb(w_n1210_0[1]),.din(n1210));
	jspl jspl_w_n1212_0(.douta(w_n1212_0[0]),.doutb(w_n1212_0[1]),.din(n1212));
	jspl jspl_w_n1213_0(.douta(w_n1213_0[0]),.doutb(w_n1213_0[1]),.din(n1213));
	jspl jspl_w_n1214_0(.douta(w_n1214_0[0]),.doutb(w_n1214_0[1]),.din(n1214));
	jspl jspl_w_n1215_0(.douta(w_n1215_0[0]),.doutb(w_n1215_0[1]),.din(n1215));
	jspl jspl_w_n1216_0(.douta(w_n1216_0[0]),.doutb(w_n1216_0[1]),.din(n1216));
	jspl jspl_w_n1217_0(.douta(w_n1217_0[0]),.doutb(w_n1217_0[1]),.din(n1217));
	jspl jspl_w_n1218_0(.douta(w_n1218_0[0]),.doutb(w_n1218_0[1]),.din(n1218));
	jspl jspl_w_n1219_0(.douta(w_n1219_0[0]),.doutb(w_n1219_0[1]),.din(n1219));
	jspl jspl_w_n1220_0(.douta(w_n1220_0[0]),.doutb(w_n1220_0[1]),.din(n1220));
	jspl jspl_w_n1221_0(.douta(w_n1221_0[0]),.doutb(w_n1221_0[1]),.din(n1221));
	jspl jspl_w_n1222_0(.douta(w_n1222_0[0]),.doutb(w_n1222_0[1]),.din(n1222));
	jspl jspl_w_n1223_0(.douta(w_n1223_0[0]),.doutb(w_n1223_0[1]),.din(n1223));
	jspl jspl_w_n1224_0(.douta(w_n1224_0[0]),.doutb(w_n1224_0[1]),.din(n1224));
	jspl jspl_w_n1225_0(.douta(w_n1225_0[0]),.doutb(w_n1225_0[1]),.din(n1225));
	jspl jspl_w_n1226_0(.douta(w_n1226_0[0]),.doutb(w_n1226_0[1]),.din(n1226));
	jspl jspl_w_n1227_0(.douta(w_n1227_0[0]),.doutb(w_n1227_0[1]),.din(n1227));
	jspl jspl_w_n1228_0(.douta(w_n1228_0[0]),.doutb(w_n1228_0[1]),.din(n1228));
	jspl jspl_w_n1229_0(.douta(w_n1229_0[0]),.doutb(w_n1229_0[1]),.din(n1229));
	jspl jspl_w_n1230_0(.douta(w_n1230_0[0]),.doutb(w_n1230_0[1]),.din(n1230));
	jspl jspl_w_n1231_0(.douta(w_n1231_0[0]),.doutb(w_n1231_0[1]),.din(n1231));
	jspl jspl_w_n1232_0(.douta(w_n1232_0[0]),.doutb(w_n1232_0[1]),.din(n1232));
	jspl jspl_w_n1234_0(.douta(w_n1234_0[0]),.doutb(w_n1234_0[1]),.din(n1234));
	jspl jspl_w_n1236_0(.douta(w_n1236_0[0]),.doutb(w_n1236_0[1]),.din(n1236));
	jspl jspl_w_n1237_0(.douta(w_n1237_0[0]),.doutb(w_n1237_0[1]),.din(n1237));
	jspl jspl_w_n1238_0(.douta(w_n1238_0[0]),.doutb(w_n1238_0[1]),.din(n1238));
	jspl jspl_w_n1244_0(.douta(w_n1244_0[0]),.doutb(w_n1244_0[1]),.din(n1244));
	jspl jspl_w_n1247_0(.douta(w_dff_A_2DXqsfki9_0),.doutb(w_n1247_0[1]),.din(n1247));
	jspl jspl_w_n1248_0(.douta(w_n1248_0[0]),.doutb(w_n1248_0[1]),.din(w_dff_B_akaHYtU43_2));
	jspl jspl_w_n1251_0(.douta(w_n1251_0[0]),.doutb(w_dff_A_KykJmTCb5_1),.din(n1251));
	jspl jspl_w_n1253_0(.douta(w_n1253_0[0]),.doutb(w_n1253_0[1]),.din(w_dff_B_IQs7OLLp0_2));
	jspl jspl_w_n1256_0(.douta(w_n1256_0[0]),.doutb(w_n1256_0[1]),.din(w_dff_B_UP6lgHQk0_2));
	jspl jspl_w_n1258_0(.douta(w_n1258_0[0]),.doutb(w_n1258_0[1]),.din(w_dff_B_VQgZ5SR97_2));
	jspl jspl_w_n1261_0(.douta(w_n1261_0[0]),.doutb(w_n1261_0[1]),.din(w_dff_B_r9HkWtyQ6_2));
	jspl jspl_w_n1263_0(.douta(w_n1263_0[0]),.doutb(w_n1263_0[1]),.din(w_dff_B_RpWXsmZk5_2));
	jspl jspl_w_n1266_0(.douta(w_n1266_0[0]),.doutb(w_n1266_0[1]),.din(w_dff_B_aDoAwMgG7_2));
	jspl jspl_w_n1268_0(.douta(w_n1268_0[0]),.doutb(w_n1268_0[1]),.din(w_dff_B_8mTW0Vt24_2));
	jspl jspl_w_n1271_0(.douta(w_n1271_0[0]),.doutb(w_n1271_0[1]),.din(w_dff_B_OrMlmBB98_2));
	jspl jspl_w_n1273_0(.douta(w_n1273_0[0]),.doutb(w_n1273_0[1]),.din(w_dff_B_fZVZwQfO1_2));
	jspl jspl_w_n1276_0(.douta(w_n1276_0[0]),.doutb(w_n1276_0[1]),.din(w_dff_B_1zPUAOOj0_2));
	jspl jspl_w_n1278_0(.douta(w_n1278_0[0]),.doutb(w_n1278_0[1]),.din(w_dff_B_D87deOIr2_2));
	jspl jspl_w_n1281_0(.douta(w_n1281_0[0]),.doutb(w_n1281_0[1]),.din(w_dff_B_uojRNQmk5_2));
	jspl jspl_w_n1283_0(.douta(w_n1283_0[0]),.doutb(w_n1283_0[1]),.din(w_dff_B_fnGQfLsP3_2));
	jspl jspl_w_n1286_0(.douta(w_n1286_0[0]),.doutb(w_n1286_0[1]),.din(w_dff_B_UslNWrpR7_2));
	jspl jspl_w_n1288_0(.douta(w_n1288_0[0]),.doutb(w_n1288_0[1]),.din(w_dff_B_cVNuB1795_2));
	jspl jspl_w_n1291_0(.douta(w_n1291_0[0]),.doutb(w_n1291_0[1]),.din(w_dff_B_Lbwdgh9C9_2));
	jspl jspl_w_n1293_0(.douta(w_n1293_0[0]),.doutb(w_n1293_0[1]),.din(w_dff_B_rKVR8sWE1_2));
	jspl jspl_w_n1296_0(.douta(w_n1296_0[0]),.doutb(w_n1296_0[1]),.din(w_dff_B_JjO1MDJb9_2));
	jspl jspl_w_n1297_0(.douta(w_n1297_0[0]),.doutb(w_n1297_0[1]),.din(w_dff_B_QhMgLiIT7_2));
	jspl jspl_w_n1298_0(.douta(w_n1298_0[0]),.doutb(w_n1298_0[1]),.din(w_dff_B_Ki1nZEhn6_2));
	jspl jspl_w_n1301_0(.douta(w_n1301_0[0]),.doutb(w_n1301_0[1]),.din(n1301));
	jspl jspl_w_n1303_0(.douta(w_n1303_0[0]),.doutb(w_n1303_0[1]),.din(n1303));
	jspl jspl_w_n1304_0(.douta(w_n1304_0[0]),.doutb(w_n1304_0[1]),.din(n1304));
	jspl jspl_w_n1305_0(.douta(w_n1305_0[0]),.doutb(w_n1305_0[1]),.din(n1305));
	jspl jspl_w_n1306_0(.douta(w_n1306_0[0]),.doutb(w_n1306_0[1]),.din(n1306));
	jspl jspl_w_n1307_0(.douta(w_n1307_0[0]),.doutb(w_n1307_0[1]),.din(n1307));
	jspl jspl_w_n1308_0(.douta(w_n1308_0[0]),.doutb(w_n1308_0[1]),.din(n1308));
	jspl jspl_w_n1309_0(.douta(w_n1309_0[0]),.doutb(w_n1309_0[1]),.din(n1309));
	jspl jspl_w_n1310_0(.douta(w_n1310_0[0]),.doutb(w_n1310_0[1]),.din(n1310));
	jspl jspl_w_n1311_0(.douta(w_n1311_0[0]),.doutb(w_n1311_0[1]),.din(n1311));
	jspl jspl_w_n1312_0(.douta(w_n1312_0[0]),.doutb(w_n1312_0[1]),.din(n1312));
	jspl jspl_w_n1313_0(.douta(w_n1313_0[0]),.doutb(w_n1313_0[1]),.din(n1313));
	jspl jspl_w_n1314_0(.douta(w_n1314_0[0]),.doutb(w_n1314_0[1]),.din(n1314));
	jspl jspl_w_n1315_0(.douta(w_n1315_0[0]),.doutb(w_n1315_0[1]),.din(n1315));
	jspl jspl_w_n1316_0(.douta(w_n1316_0[0]),.doutb(w_n1316_0[1]),.din(n1316));
	jspl jspl_w_n1317_0(.douta(w_n1317_0[0]),.doutb(w_n1317_0[1]),.din(n1317));
	jspl jspl_w_n1318_0(.douta(w_n1318_0[0]),.doutb(w_n1318_0[1]),.din(n1318));
	jspl jspl_w_n1319_0(.douta(w_n1319_0[0]),.doutb(w_n1319_0[1]),.din(n1319));
	jspl jspl_w_n1320_0(.douta(w_n1320_0[0]),.doutb(w_n1320_0[1]),.din(n1320));
	jspl jspl_w_n1321_0(.douta(w_n1321_0[0]),.doutb(w_n1321_0[1]),.din(n1321));
	jspl jspl_w_n1322_0(.douta(w_n1322_0[0]),.doutb(w_n1322_0[1]),.din(n1322));
	jspl jspl_w_n1324_0(.douta(w_n1324_0[0]),.doutb(w_n1324_0[1]),.din(n1324));
	jspl jspl_w_n1325_0(.douta(w_n1325_0[0]),.doutb(w_n1325_0[1]),.din(n1325));
	jspl jspl_w_n1326_0(.douta(w_dff_A_3bZjpayx8_0),.doutb(w_n1326_0[1]),.din(n1326));
	jspl jspl_w_n1332_0(.douta(w_dff_A_NXQdRrj24_0),.doutb(w_n1332_0[1]),.din(n1332));
	jspl jspl_w_n1337_0(.douta(w_n1337_0[0]),.doutb(w_n1337_0[1]),.din(w_dff_B_3D2mMVj74_2));
	jspl jspl_w_n1338_0(.douta(w_n1338_0[0]),.doutb(w_n1338_0[1]),.din(w_dff_B_L9bSzvvj0_2));
	jspl jspl_w_n1341_0(.douta(w_n1341_0[0]),.doutb(w_dff_A_1gzZBzEp4_1),.din(n1341));
	jspl jspl_w_n1343_0(.douta(w_n1343_0[0]),.doutb(w_n1343_0[1]),.din(w_dff_B_kiAL6Qoz4_2));
	jspl jspl_w_n1346_0(.douta(w_n1346_0[0]),.doutb(w_n1346_0[1]),.din(w_dff_B_hARVlZ0U7_2));
	jspl jspl_w_n1348_0(.douta(w_n1348_0[0]),.doutb(w_n1348_0[1]),.din(w_dff_B_rsbKbUpA0_2));
	jspl jspl_w_n1351_0(.douta(w_n1351_0[0]),.doutb(w_n1351_0[1]),.din(w_dff_B_chs9YUMz7_2));
	jspl jspl_w_n1353_0(.douta(w_n1353_0[0]),.doutb(w_n1353_0[1]),.din(w_dff_B_pZFYSmTh4_2));
	jspl jspl_w_n1356_0(.douta(w_n1356_0[0]),.doutb(w_n1356_0[1]),.din(w_dff_B_hux4zV000_2));
	jspl jspl_w_n1358_0(.douta(w_n1358_0[0]),.doutb(w_n1358_0[1]),.din(w_dff_B_kV5tHOnr0_2));
	jspl jspl_w_n1361_0(.douta(w_n1361_0[0]),.doutb(w_n1361_0[1]),.din(w_dff_B_RK8XfEmu7_2));
	jspl jspl_w_n1363_0(.douta(w_n1363_0[0]),.doutb(w_n1363_0[1]),.din(w_dff_B_HexU8YbC7_2));
	jspl jspl_w_n1366_0(.douta(w_n1366_0[0]),.doutb(w_n1366_0[1]),.din(w_dff_B_iWMEV3TI9_2));
	jspl jspl_w_n1368_0(.douta(w_n1368_0[0]),.doutb(w_n1368_0[1]),.din(w_dff_B_Mn7l1HXh8_2));
	jspl jspl_w_n1371_0(.douta(w_n1371_0[0]),.doutb(w_n1371_0[1]),.din(w_dff_B_PRIeYDNt5_2));
	jspl jspl_w_n1373_0(.douta(w_n1373_0[0]),.doutb(w_n1373_0[1]),.din(w_dff_B_iQXQbdJt5_2));
	jspl jspl_w_n1376_0(.douta(w_n1376_0[0]),.doutb(w_n1376_0[1]),.din(w_dff_B_A0i2702a4_2));
	jspl jspl_w_n1378_0(.douta(w_n1378_0[0]),.doutb(w_n1378_0[1]),.din(w_dff_B_L60jpsp08_2));
	jspl jspl_w_n1381_0(.douta(w_n1381_0[0]),.doutb(w_n1381_0[1]),.din(w_dff_B_D4V5DroH4_2));
	jspl jspl_w_n1382_0(.douta(w_n1382_0[0]),.doutb(w_n1382_0[1]),.din(w_dff_B_GjFxFVhf7_2));
	jspl jspl_w_n1383_0(.douta(w_n1383_0[0]),.doutb(w_n1383_0[1]),.din(w_dff_B_e44LNbve0_2));
	jspl jspl_w_n1386_0(.douta(w_n1386_0[0]),.doutb(w_n1386_0[1]),.din(n1386));
	jspl jspl_w_n1388_0(.douta(w_n1388_0[0]),.doutb(w_n1388_0[1]),.din(n1388));
	jspl jspl_w_n1389_0(.douta(w_n1389_0[0]),.doutb(w_n1389_0[1]),.din(n1389));
	jspl jspl_w_n1390_0(.douta(w_n1390_0[0]),.doutb(w_n1390_0[1]),.din(n1390));
	jspl jspl_w_n1391_0(.douta(w_n1391_0[0]),.doutb(w_n1391_0[1]),.din(n1391));
	jspl jspl_w_n1392_0(.douta(w_n1392_0[0]),.doutb(w_n1392_0[1]),.din(n1392));
	jspl jspl_w_n1393_0(.douta(w_n1393_0[0]),.doutb(w_n1393_0[1]),.din(n1393));
	jspl jspl_w_n1394_0(.douta(w_n1394_0[0]),.doutb(w_n1394_0[1]),.din(n1394));
	jspl jspl_w_n1395_0(.douta(w_n1395_0[0]),.doutb(w_n1395_0[1]),.din(n1395));
	jspl jspl_w_n1396_0(.douta(w_n1396_0[0]),.doutb(w_n1396_0[1]),.din(n1396));
	jspl jspl_w_n1397_0(.douta(w_n1397_0[0]),.doutb(w_n1397_0[1]),.din(n1397));
	jspl jspl_w_n1398_0(.douta(w_n1398_0[0]),.doutb(w_n1398_0[1]),.din(n1398));
	jspl jspl_w_n1399_0(.douta(w_n1399_0[0]),.doutb(w_n1399_0[1]),.din(n1399));
	jspl jspl_w_n1400_0(.douta(w_n1400_0[0]),.doutb(w_n1400_0[1]),.din(n1400));
	jspl jspl_w_n1401_0(.douta(w_n1401_0[0]),.doutb(w_n1401_0[1]),.din(n1401));
	jspl jspl_w_n1402_0(.douta(w_n1402_0[0]),.doutb(w_n1402_0[1]),.din(n1402));
	jspl jspl_w_n1403_0(.douta(w_n1403_0[0]),.doutb(w_n1403_0[1]),.din(n1403));
	jspl jspl_w_n1404_0(.douta(w_n1404_0[0]),.doutb(w_n1404_0[1]),.din(n1404));
	jspl jspl_w_n1405_0(.douta(w_n1405_0[0]),.doutb(w_n1405_0[1]),.din(n1405));
	jspl jspl_w_n1407_0(.douta(w_n1407_0[0]),.doutb(w_n1407_0[1]),.din(n1407));
	jspl jspl_w_n1409_0(.douta(w_n1409_0[0]),.doutb(w_n1409_0[1]),.din(n1409));
	jspl jspl_w_n1410_0(.douta(w_n1410_0[0]),.doutb(w_n1410_0[1]),.din(n1410));
	jspl jspl_w_n1415_0(.douta(w_n1415_0[0]),.doutb(w_n1415_0[1]),.din(n1415));
	jspl jspl_w_n1420_0(.douta(w_n1420_0[0]),.doutb(w_n1420_0[1]),.din(w_dff_B_TJfsuamC7_2));
	jspl jspl_w_n1421_0(.douta(w_n1421_0[0]),.doutb(w_n1421_0[1]),.din(w_dff_B_MO3xkrHL2_2));
	jspl jspl_w_n1424_0(.douta(w_n1424_0[0]),.doutb(w_dff_A_km6ZBDLX1_1),.din(n1424));
	jspl jspl_w_n1426_0(.douta(w_n1426_0[0]),.doutb(w_n1426_0[1]),.din(w_dff_B_NOISaytV5_2));
	jspl jspl_w_n1429_0(.douta(w_n1429_0[0]),.doutb(w_n1429_0[1]),.din(w_dff_B_6w8IAF025_2));
	jspl jspl_w_n1431_0(.douta(w_n1431_0[0]),.doutb(w_n1431_0[1]),.din(w_dff_B_ZIjzh16U2_2));
	jspl jspl_w_n1434_0(.douta(w_n1434_0[0]),.doutb(w_n1434_0[1]),.din(w_dff_B_kLPA1nxm0_2));
	jspl jspl_w_n1436_0(.douta(w_n1436_0[0]),.doutb(w_n1436_0[1]),.din(w_dff_B_aRYoTqZk7_2));
	jspl jspl_w_n1439_0(.douta(w_n1439_0[0]),.doutb(w_n1439_0[1]),.din(w_dff_B_F32ynQNJ0_2));
	jspl jspl_w_n1441_0(.douta(w_n1441_0[0]),.doutb(w_n1441_0[1]),.din(w_dff_B_Npw3mhl04_2));
	jspl jspl_w_n1444_0(.douta(w_n1444_0[0]),.doutb(w_n1444_0[1]),.din(w_dff_B_BGR6rjw04_2));
	jspl jspl_w_n1446_0(.douta(w_n1446_0[0]),.doutb(w_n1446_0[1]),.din(w_dff_B_q9yyD1qM7_2));
	jspl jspl_w_n1449_0(.douta(w_n1449_0[0]),.doutb(w_n1449_0[1]),.din(w_dff_B_Ym1N6bAQ5_2));
	jspl jspl_w_n1451_0(.douta(w_n1451_0[0]),.doutb(w_n1451_0[1]),.din(w_dff_B_jMrDNSe89_2));
	jspl jspl_w_n1454_0(.douta(w_n1454_0[0]),.doutb(w_n1454_0[1]),.din(w_dff_B_2McmDv8G7_2));
	jspl jspl_w_n1456_0(.douta(w_n1456_0[0]),.doutb(w_n1456_0[1]),.din(w_dff_B_kU5hk7Wz5_2));
	jspl jspl_w_n1459_0(.douta(w_n1459_0[0]),.doutb(w_n1459_0[1]),.din(w_dff_B_t2KKPViJ5_2));
	jspl jspl_w_n1460_0(.douta(w_n1460_0[0]),.doutb(w_n1460_0[1]),.din(w_dff_B_mDRr7Giz8_2));
	jspl jspl_w_n1461_0(.douta(w_n1461_0[0]),.doutb(w_n1461_0[1]),.din(w_dff_B_NAN3wn5C2_2));
	jspl jspl_w_n1464_0(.douta(w_n1464_0[0]),.doutb(w_n1464_0[1]),.din(n1464));
	jspl jspl_w_n1466_0(.douta(w_n1466_0[0]),.doutb(w_n1466_0[1]),.din(n1466));
	jspl jspl_w_n1467_0(.douta(w_n1467_0[0]),.doutb(w_n1467_0[1]),.din(n1467));
	jspl jspl_w_n1468_0(.douta(w_n1468_0[0]),.doutb(w_n1468_0[1]),.din(n1468));
	jspl jspl_w_n1469_0(.douta(w_n1469_0[0]),.doutb(w_n1469_0[1]),.din(n1469));
	jspl jspl_w_n1470_0(.douta(w_n1470_0[0]),.doutb(w_n1470_0[1]),.din(n1470));
	jspl jspl_w_n1471_0(.douta(w_n1471_0[0]),.doutb(w_n1471_0[1]),.din(n1471));
	jspl jspl_w_n1472_0(.douta(w_n1472_0[0]),.doutb(w_n1472_0[1]),.din(n1472));
	jspl jspl_w_n1473_0(.douta(w_n1473_0[0]),.doutb(w_n1473_0[1]),.din(n1473));
	jspl jspl_w_n1474_0(.douta(w_n1474_0[0]),.doutb(w_n1474_0[1]),.din(n1474));
	jspl jspl_w_n1475_0(.douta(w_n1475_0[0]),.doutb(w_n1475_0[1]),.din(n1475));
	jspl jspl_w_n1476_0(.douta(w_n1476_0[0]),.doutb(w_n1476_0[1]),.din(n1476));
	jspl jspl_w_n1477_0(.douta(w_n1477_0[0]),.doutb(w_n1477_0[1]),.din(n1477));
	jspl jspl_w_n1478_0(.douta(w_n1478_0[0]),.doutb(w_n1478_0[1]),.din(n1478));
	jspl jspl_w_n1479_0(.douta(w_n1479_0[0]),.doutb(w_n1479_0[1]),.din(n1479));
	jspl jspl_w_n1480_0(.douta(w_n1480_0[0]),.doutb(w_n1480_0[1]),.din(n1480));
	jspl jspl_w_n1481_0(.douta(w_n1481_0[0]),.doutb(w_n1481_0[1]),.din(n1481));
	jspl jspl_w_n1483_0(.douta(w_n1483_0[0]),.doutb(w_n1483_0[1]),.din(n1483));
	jspl jspl_w_n1485_0(.douta(w_n1485_0[0]),.doutb(w_n1485_0[1]),.din(n1485));
	jspl jspl_w_n1486_0(.douta(w_n1486_0[0]),.doutb(w_dff_A_uzm3y4NF2_1),.din(n1486));
	jspl jspl_w_n1491_0(.douta(w_n1491_0[0]),.doutb(w_n1491_0[1]),.din(n1491));
	jspl jspl_w_n1496_0(.douta(w_n1496_0[0]),.doutb(w_n1496_0[1]),.din(w_dff_B_QXDLZGjL9_2));
	jspl jspl_w_n1497_0(.douta(w_n1497_0[0]),.doutb(w_n1497_0[1]),.din(w_dff_B_GjvakE6n3_2));
	jspl jspl_w_n1500_0(.douta(w_n1500_0[0]),.doutb(w_dff_A_lLOzs8437_1),.din(n1500));
	jspl jspl_w_n1502_0(.douta(w_n1502_0[0]),.doutb(w_n1502_0[1]),.din(w_dff_B_cAOgaJXH0_2));
	jspl jspl_w_n1505_0(.douta(w_n1505_0[0]),.doutb(w_n1505_0[1]),.din(w_dff_B_M9r7IJP04_2));
	jspl jspl_w_n1507_0(.douta(w_n1507_0[0]),.doutb(w_n1507_0[1]),.din(w_dff_B_ecNw3eAu0_2));
	jspl jspl_w_n1510_0(.douta(w_n1510_0[0]),.doutb(w_n1510_0[1]),.din(w_dff_B_AZwRkMcO5_2));
	jspl jspl_w_n1512_0(.douta(w_n1512_0[0]),.doutb(w_n1512_0[1]),.din(w_dff_B_GU9LaF1R2_2));
	jspl jspl_w_n1515_0(.douta(w_n1515_0[0]),.doutb(w_n1515_0[1]),.din(w_dff_B_NHWP0S507_2));
	jspl jspl_w_n1517_0(.douta(w_n1517_0[0]),.doutb(w_n1517_0[1]),.din(w_dff_B_6DxEcXa09_2));
	jspl jspl_w_n1520_0(.douta(w_n1520_0[0]),.doutb(w_n1520_0[1]),.din(w_dff_B_S34dDBt10_2));
	jspl jspl_w_n1522_0(.douta(w_n1522_0[0]),.doutb(w_n1522_0[1]),.din(w_dff_B_SL4sG0kr9_2));
	jspl jspl_w_n1525_0(.douta(w_n1525_0[0]),.doutb(w_n1525_0[1]),.din(w_dff_B_JTtRBhye0_2));
	jspl jspl_w_n1527_0(.douta(w_n1527_0[0]),.doutb(w_n1527_0[1]),.din(w_dff_B_j9F6fm7H5_2));
	jspl jspl_w_n1530_0(.douta(w_n1530_0[0]),.doutb(w_n1530_0[1]),.din(w_dff_B_CT3WHjNg5_2));
	jspl jspl_w_n1531_0(.douta(w_n1531_0[0]),.doutb(w_n1531_0[1]),.din(w_dff_B_RaaEakny6_2));
	jspl jspl_w_n1532_0(.douta(w_n1532_0[0]),.doutb(w_n1532_0[1]),.din(w_dff_B_0maDXt469_2));
	jspl jspl_w_n1535_0(.douta(w_n1535_0[0]),.doutb(w_n1535_0[1]),.din(n1535));
	jspl jspl_w_n1537_0(.douta(w_n1537_0[0]),.doutb(w_n1537_0[1]),.din(n1537));
	jspl jspl_w_n1538_0(.douta(w_n1538_0[0]),.doutb(w_n1538_0[1]),.din(n1538));
	jspl jspl_w_n1539_0(.douta(w_n1539_0[0]),.doutb(w_n1539_0[1]),.din(n1539));
	jspl jspl_w_n1540_0(.douta(w_n1540_0[0]),.doutb(w_n1540_0[1]),.din(n1540));
	jspl jspl_w_n1541_0(.douta(w_n1541_0[0]),.doutb(w_n1541_0[1]),.din(n1541));
	jspl jspl_w_n1542_0(.douta(w_n1542_0[0]),.doutb(w_n1542_0[1]),.din(n1542));
	jspl jspl_w_n1543_0(.douta(w_n1543_0[0]),.doutb(w_n1543_0[1]),.din(n1543));
	jspl jspl_w_n1544_0(.douta(w_n1544_0[0]),.doutb(w_n1544_0[1]),.din(n1544));
	jspl jspl_w_n1545_0(.douta(w_n1545_0[0]),.doutb(w_n1545_0[1]),.din(n1545));
	jspl jspl_w_n1546_0(.douta(w_n1546_0[0]),.doutb(w_n1546_0[1]),.din(n1546));
	jspl jspl_w_n1547_0(.douta(w_n1547_0[0]),.doutb(w_n1547_0[1]),.din(n1547));
	jspl jspl_w_n1548_0(.douta(w_n1548_0[0]),.doutb(w_n1548_0[1]),.din(n1548));
	jspl jspl_w_n1549_0(.douta(w_n1549_0[0]),.doutb(w_n1549_0[1]),.din(n1549));
	jspl jspl_w_n1550_0(.douta(w_n1550_0[0]),.doutb(w_n1550_0[1]),.din(n1550));
	jspl jspl_w_n1552_0(.douta(w_n1552_0[0]),.doutb(w_n1552_0[1]),.din(n1552));
	jspl jspl_w_n1554_0(.douta(w_n1554_0[0]),.doutb(w_n1554_0[1]),.din(n1554));
	jspl jspl_w_n1555_0(.douta(w_n1555_0[0]),.doutb(w_dff_A_GB6k6xy42_1),.din(n1555));
	jspl jspl_w_n1560_0(.douta(w_n1560_0[0]),.doutb(w_n1560_0[1]),.din(n1560));
	jspl jspl_w_n1565_0(.douta(w_n1565_0[0]),.doutb(w_n1565_0[1]),.din(w_dff_B_pZiXbu383_2));
	jspl jspl_w_n1566_0(.douta(w_n1566_0[0]),.doutb(w_n1566_0[1]),.din(w_dff_B_OF2s7hnL4_2));
	jspl jspl_w_n1569_0(.douta(w_n1569_0[0]),.doutb(w_dff_A_MJhgLnrt6_1),.din(n1569));
	jspl jspl_w_n1571_0(.douta(w_n1571_0[0]),.doutb(w_n1571_0[1]),.din(w_dff_B_cEZ81KbZ7_2));
	jspl jspl_w_n1574_0(.douta(w_n1574_0[0]),.doutb(w_n1574_0[1]),.din(w_dff_B_e9uZd5Xu4_2));
	jspl jspl_w_n1576_0(.douta(w_n1576_0[0]),.doutb(w_n1576_0[1]),.din(w_dff_B_MoBDJCAb9_2));
	jspl jspl_w_n1579_0(.douta(w_n1579_0[0]),.doutb(w_n1579_0[1]),.din(w_dff_B_57WarLly3_2));
	jspl jspl_w_n1581_0(.douta(w_n1581_0[0]),.doutb(w_n1581_0[1]),.din(w_dff_B_fvvSlpHj4_2));
	jspl jspl_w_n1584_0(.douta(w_n1584_0[0]),.doutb(w_n1584_0[1]),.din(w_dff_B_piK1THr49_2));
	jspl jspl_w_n1586_0(.douta(w_n1586_0[0]),.doutb(w_n1586_0[1]),.din(w_dff_B_mrZXleBf5_2));
	jspl jspl_w_n1589_0(.douta(w_n1589_0[0]),.doutb(w_n1589_0[1]),.din(w_dff_B_TQ1Z6noW7_2));
	jspl jspl_w_n1591_0(.douta(w_n1591_0[0]),.doutb(w_n1591_0[1]),.din(w_dff_B_ztfniFbs0_2));
	jspl jspl_w_n1594_0(.douta(w_n1594_0[0]),.doutb(w_n1594_0[1]),.din(w_dff_B_PXxDP2ZQ2_2));
	jspl jspl_w_n1595_0(.douta(w_n1595_0[0]),.doutb(w_n1595_0[1]),.din(w_dff_B_6vXFpnbZ4_2));
	jspl jspl_w_n1596_0(.douta(w_n1596_0[0]),.doutb(w_n1596_0[1]),.din(w_dff_B_dHTgEsif0_2));
	jspl jspl_w_n1599_0(.douta(w_n1599_0[0]),.doutb(w_n1599_0[1]),.din(n1599));
	jspl jspl_w_n1601_0(.douta(w_n1601_0[0]),.doutb(w_n1601_0[1]),.din(n1601));
	jspl jspl_w_n1602_0(.douta(w_n1602_0[0]),.doutb(w_n1602_0[1]),.din(n1602));
	jspl jspl_w_n1603_0(.douta(w_n1603_0[0]),.doutb(w_n1603_0[1]),.din(n1603));
	jspl jspl_w_n1604_0(.douta(w_n1604_0[0]),.doutb(w_n1604_0[1]),.din(n1604));
	jspl jspl_w_n1605_0(.douta(w_n1605_0[0]),.doutb(w_n1605_0[1]),.din(n1605));
	jspl jspl_w_n1606_0(.douta(w_n1606_0[0]),.doutb(w_n1606_0[1]),.din(n1606));
	jspl jspl_w_n1607_0(.douta(w_n1607_0[0]),.doutb(w_n1607_0[1]),.din(n1607));
	jspl jspl_w_n1608_0(.douta(w_n1608_0[0]),.doutb(w_n1608_0[1]),.din(n1608));
	jspl jspl_w_n1609_0(.douta(w_n1609_0[0]),.doutb(w_n1609_0[1]),.din(n1609));
	jspl jspl_w_n1610_0(.douta(w_n1610_0[0]),.doutb(w_n1610_0[1]),.din(n1610));
	jspl jspl_w_n1611_0(.douta(w_n1611_0[0]),.doutb(w_n1611_0[1]),.din(n1611));
	jspl jspl_w_n1612_0(.douta(w_n1612_0[0]),.doutb(w_n1612_0[1]),.din(n1612));
	jspl jspl_w_n1614_0(.douta(w_n1614_0[0]),.doutb(w_n1614_0[1]),.din(n1614));
	jspl jspl_w_n1616_0(.douta(w_n1616_0[0]),.doutb(w_n1616_0[1]),.din(n1616));
	jspl jspl_w_n1617_0(.douta(w_n1617_0[0]),.doutb(w_dff_A_vLMIrqfW2_1),.din(n1617));
	jspl jspl_w_n1622_0(.douta(w_n1622_0[0]),.doutb(w_n1622_0[1]),.din(n1622));
	jspl jspl_w_n1627_0(.douta(w_n1627_0[0]),.doutb(w_n1627_0[1]),.din(w_dff_B_Q6bCvniE8_2));
	jspl jspl_w_n1628_0(.douta(w_n1628_0[0]),.doutb(w_n1628_0[1]),.din(w_dff_B_fOOVUDPi4_2));
	jspl jspl_w_n1631_0(.douta(w_n1631_0[0]),.doutb(w_dff_A_QTN0cg9q0_1),.din(n1631));
	jspl jspl_w_n1633_0(.douta(w_n1633_0[0]),.doutb(w_n1633_0[1]),.din(w_dff_B_76gp0Rog3_2));
	jspl jspl_w_n1636_0(.douta(w_n1636_0[0]),.doutb(w_n1636_0[1]),.din(w_dff_B_iECabImR9_2));
	jspl jspl_w_n1638_0(.douta(w_n1638_0[0]),.doutb(w_n1638_0[1]),.din(w_dff_B_l2Pjn05G8_2));
	jspl jspl_w_n1641_0(.douta(w_n1641_0[0]),.doutb(w_n1641_0[1]),.din(w_dff_B_OccyCEz61_2));
	jspl jspl_w_n1643_0(.douta(w_n1643_0[0]),.doutb(w_n1643_0[1]),.din(w_dff_B_daRlOphW0_2));
	jspl jspl_w_n1646_0(.douta(w_n1646_0[0]),.doutb(w_n1646_0[1]),.din(w_dff_B_ZpOkK2qv5_2));
	jspl jspl_w_n1648_0(.douta(w_n1648_0[0]),.doutb(w_n1648_0[1]),.din(w_dff_B_5vAg64vY8_2));
	jspl jspl_w_n1651_0(.douta(w_n1651_0[0]),.doutb(w_n1651_0[1]),.din(w_dff_B_ZgtcSHaY9_2));
	jspl jspl_w_n1652_0(.douta(w_n1652_0[0]),.doutb(w_n1652_0[1]),.din(w_dff_B_Jl7bPsJO7_2));
	jspl jspl_w_n1653_0(.douta(w_n1653_0[0]),.doutb(w_n1653_0[1]),.din(w_dff_B_bsop8f2T8_2));
	jspl jspl_w_n1656_0(.douta(w_n1656_0[0]),.doutb(w_n1656_0[1]),.din(n1656));
	jspl jspl_w_n1658_0(.douta(w_n1658_0[0]),.doutb(w_n1658_0[1]),.din(n1658));
	jspl jspl_w_n1659_0(.douta(w_n1659_0[0]),.doutb(w_n1659_0[1]),.din(n1659));
	jspl jspl_w_n1660_0(.douta(w_n1660_0[0]),.doutb(w_n1660_0[1]),.din(n1660));
	jspl jspl_w_n1661_0(.douta(w_n1661_0[0]),.doutb(w_n1661_0[1]),.din(n1661));
	jspl jspl_w_n1662_0(.douta(w_n1662_0[0]),.doutb(w_n1662_0[1]),.din(n1662));
	jspl jspl_w_n1663_0(.douta(w_n1663_0[0]),.doutb(w_n1663_0[1]),.din(n1663));
	jspl jspl_w_n1664_0(.douta(w_n1664_0[0]),.doutb(w_n1664_0[1]),.din(n1664));
	jspl jspl_w_n1665_0(.douta(w_n1665_0[0]),.doutb(w_n1665_0[1]),.din(n1665));
	jspl jspl_w_n1666_0(.douta(w_n1666_0[0]),.doutb(w_n1666_0[1]),.din(n1666));
	jspl jspl_w_n1667_0(.douta(w_n1667_0[0]),.doutb(w_n1667_0[1]),.din(n1667));
	jspl jspl_w_n1669_0(.douta(w_n1669_0[0]),.doutb(w_n1669_0[1]),.din(n1669));
	jspl jspl_w_n1671_0(.douta(w_n1671_0[0]),.doutb(w_n1671_0[1]),.din(n1671));
	jspl jspl_w_n1672_0(.douta(w_n1672_0[0]),.doutb(w_dff_A_j7CybSZ25_1),.din(n1672));
	jspl jspl_w_n1677_0(.douta(w_n1677_0[0]),.doutb(w_n1677_0[1]),.din(n1677));
	jspl jspl_w_n1682_0(.douta(w_n1682_0[0]),.doutb(w_n1682_0[1]),.din(w_dff_B_FtolqQ735_2));
	jspl jspl_w_n1684_0(.douta(w_n1684_0[0]),.doutb(w_n1684_0[1]),.din(w_dff_B_gMcNfZFB1_2));
	jspl jspl_w_n1687_0(.douta(w_n1687_0[0]),.doutb(w_n1687_0[1]),.din(w_dff_B_ns7ZlvK11_2));
	jspl jspl_w_n1689_0(.douta(w_n1689_0[0]),.doutb(w_n1689_0[1]),.din(w_dff_B_3X9ysqiv8_2));
	jspl jspl_w_n1692_0(.douta(w_n1692_0[0]),.doutb(w_n1692_0[1]),.din(w_dff_B_hmSzzKIG2_2));
	jspl jspl_w_n1694_0(.douta(w_n1694_0[0]),.doutb(w_n1694_0[1]),.din(w_dff_B_koax4oEL4_2));
	jspl jspl_w_n1697_0(.douta(w_n1697_0[0]),.doutb(w_n1697_0[1]),.din(w_dff_B_kVKZu0VS8_2));
	jspl jspl_w_n1699_0(.douta(w_n1699_0[0]),.doutb(w_n1699_0[1]),.din(w_dff_B_GUFsXUGN2_2));
	jspl jspl_w_n1702_0(.douta(w_n1702_0[0]),.doutb(w_n1702_0[1]),.din(w_dff_B_qSMUqC6J3_2));
	jspl jspl_w_n1703_0(.douta(w_n1703_0[0]),.doutb(w_n1703_0[1]),.din(w_dff_B_QZUrIAZs9_2));
	jspl jspl_w_n1704_0(.douta(w_n1704_0[0]),.doutb(w_n1704_0[1]),.din(w_dff_B_mXwsCmDM5_2));
	jspl jspl_w_n1707_0(.douta(w_n1707_0[0]),.doutb(w_n1707_0[1]),.din(n1707));
	jspl jspl_w_n1709_0(.douta(w_n1709_0[0]),.doutb(w_n1709_0[1]),.din(n1709));
	jspl jspl_w_n1710_0(.douta(w_n1710_0[0]),.doutb(w_n1710_0[1]),.din(n1710));
	jspl jspl_w_n1711_0(.douta(w_n1711_0[0]),.doutb(w_n1711_0[1]),.din(n1711));
	jspl jspl_w_n1712_0(.douta(w_n1712_0[0]),.doutb(w_n1712_0[1]),.din(n1712));
	jspl jspl_w_n1713_0(.douta(w_n1713_0[0]),.doutb(w_n1713_0[1]),.din(n1713));
	jspl jspl_w_n1714_0(.douta(w_n1714_0[0]),.doutb(w_n1714_0[1]),.din(n1714));
	jspl jspl_w_n1715_0(.douta(w_n1715_0[0]),.doutb(w_n1715_0[1]),.din(n1715));
	jspl jspl_w_n1716_0(.douta(w_n1716_0[0]),.doutb(w_n1716_0[1]),.din(n1716));
	jspl jspl_w_n1717_0(.douta(w_n1717_0[0]),.doutb(w_n1717_0[1]),.din(n1717));
	jspl jspl_w_n1719_0(.douta(w_n1719_0[0]),.doutb(w_n1719_0[1]),.din(n1719));
	jspl jspl_w_n1720_0(.douta(w_n1720_0[0]),.doutb(w_dff_A_K74FCtSl7_1),.din(n1720));
	jspl jspl_w_n1725_0(.douta(w_n1725_0[0]),.doutb(w_n1725_0[1]),.din(n1725));
	jspl jspl_w_n1728_0(.douta(w_n1728_0[0]),.doutb(w_dff_A_u5pAxSPk8_1),.din(n1728));
	jspl jspl_w_n1730_0(.douta(w_n1730_0[0]),.doutb(w_n1730_0[1]),.din(w_dff_B_b5xB4cfa7_2));
	jspl jspl_w_n1733_0(.douta(w_n1733_0[0]),.doutb(w_n1733_0[1]),.din(w_dff_B_sWLejboO0_2));
	jspl jspl_w_n1735_0(.douta(w_n1735_0[0]),.doutb(w_n1735_0[1]),.din(w_dff_B_Onv7pv8s0_2));
	jspl jspl_w_n1738_0(.douta(w_n1738_0[0]),.doutb(w_n1738_0[1]),.din(w_dff_B_D8AJXiMT8_2));
	jspl jspl_w_n1740_0(.douta(w_n1740_0[0]),.doutb(w_n1740_0[1]),.din(w_dff_B_ZPhpAERb4_2));
	jspl jspl_w_n1743_0(.douta(w_n1743_0[0]),.doutb(w_n1743_0[1]),.din(w_dff_B_c0Qs8dBf7_2));
	jspl jspl_w_n1744_0(.douta(w_n1744_0[0]),.doutb(w_n1744_0[1]),.din(w_dff_B_bqTe6Lzj1_2));
	jspl jspl_w_n1745_0(.douta(w_n1745_0[0]),.doutb(w_n1745_0[1]),.din(w_dff_B_z5QIOJ2o2_2));
	jspl jspl_w_n1748_0(.douta(w_n1748_0[0]),.doutb(w_n1748_0[1]),.din(n1748));
	jspl jspl_w_n1750_0(.douta(w_n1750_0[0]),.doutb(w_n1750_0[1]),.din(n1750));
	jspl jspl_w_n1751_0(.douta(w_n1751_0[0]),.doutb(w_n1751_0[1]),.din(n1751));
	jspl jspl_w_n1752_0(.douta(w_n1752_0[0]),.doutb(w_n1752_0[1]),.din(n1752));
	jspl jspl_w_n1753_0(.douta(w_n1753_0[0]),.doutb(w_n1753_0[1]),.din(n1753));
	jspl jspl_w_n1754_0(.douta(w_n1754_0[0]),.doutb(w_n1754_0[1]),.din(n1754));
	jspl jspl_w_n1755_0(.douta(w_n1755_0[0]),.doutb(w_n1755_0[1]),.din(n1755));
	jspl jspl_w_n1756_0(.douta(w_n1756_0[0]),.doutb(w_n1756_0[1]),.din(n1756));
	jspl jspl_w_n1757_0(.douta(w_n1757_0[0]),.doutb(w_n1757_0[1]),.din(n1757));
	jspl jspl_w_n1758_0(.douta(w_n1758_0[0]),.doutb(w_dff_A_4zVLMqc52_1),.din(n1758));
	jspl jspl_w_n1765_0(.douta(w_n1765_0[0]),.doutb(w_n1765_0[1]),.din(n1765));
	jspl jspl_w_n1768_0(.douta(w_n1768_0[0]),.doutb(w_dff_A_FthOBBaS1_1),.din(n1768));
	jspl jspl_w_n1770_0(.douta(w_n1770_0[0]),.doutb(w_n1770_0[1]),.din(w_dff_B_XLEbZbGh4_2));
	jspl jspl_w_n1773_0(.douta(w_n1773_0[0]),.doutb(w_n1773_0[1]),.din(w_dff_B_dAbLNxEq4_2));
	jspl jspl_w_n1775_0(.douta(w_n1775_0[0]),.doutb(w_n1775_0[1]),.din(w_dff_B_gbgBrA6H6_2));
	jspl jspl_w_n1778_0(.douta(w_n1778_0[0]),.doutb(w_n1778_0[1]),.din(w_dff_B_gSyS7sQ69_2));
	jspl jspl_w_n1779_0(.douta(w_n1779_0[0]),.doutb(w_n1779_0[1]),.din(w_dff_B_yUI2ohxu1_2));
	jspl jspl_w_n1780_0(.douta(w_n1780_0[0]),.doutb(w_n1780_0[1]),.din(w_dff_B_2DNCISpa2_2));
	jspl jspl_w_n1783_0(.douta(w_n1783_0[0]),.doutb(w_n1783_0[1]),.din(n1783));
	jspl jspl_w_n1785_0(.douta(w_n1785_0[0]),.doutb(w_n1785_0[1]),.din(n1785));
	jspl jspl_w_n1786_0(.douta(w_n1786_0[0]),.doutb(w_n1786_0[1]),.din(n1786));
	jspl jspl_w_n1787_0(.douta(w_n1787_0[0]),.doutb(w_n1787_0[1]),.din(n1787));
	jspl jspl_w_n1788_0(.douta(w_n1788_0[0]),.doutb(w_n1788_0[1]),.din(n1788));
	jspl jspl_w_n1789_0(.douta(w_n1789_0[0]),.doutb(w_n1789_0[1]),.din(n1789));
	jspl jspl_w_n1790_0(.douta(w_n1790_0[0]),.doutb(w_n1790_0[1]),.din(n1790));
	jspl jspl_w_n1791_0(.douta(w_n1791_0[0]),.doutb(w_dff_A_RZILa9VN8_1),.din(n1791));
	jspl jspl_w_n1798_0(.douta(w_n1798_0[0]),.doutb(w_n1798_0[1]),.din(n1798));
	jspl jspl_w_n1801_0(.douta(w_n1801_0[0]),.doutb(w_dff_A_ssrXAKtQ0_1),.din(n1801));
	jspl jspl_w_n1803_0(.douta(w_n1803_0[0]),.doutb(w_n1803_0[1]),.din(w_dff_B_gDyZj84K6_2));
	jspl jspl_w_n1806_0(.douta(w_n1806_0[0]),.doutb(w_n1806_0[1]),.din(w_dff_B_ePWWhOLk3_2));
	jspl jspl_w_n1807_0(.douta(w_n1807_0[0]),.doutb(w_n1807_0[1]),.din(w_dff_B_BjKCTGGi5_2));
	jspl jspl_w_n1808_0(.douta(w_n1808_0[0]),.doutb(w_n1808_0[1]),.din(w_dff_B_mdap9Y3v1_2));
	jspl jspl_w_n1811_0(.douta(w_n1811_0[0]),.doutb(w_n1811_0[1]),.din(n1811));
	jspl jspl_w_n1813_0(.douta(w_n1813_0[0]),.doutb(w_n1813_0[1]),.din(n1813));
	jspl jspl_w_n1814_0(.douta(w_n1814_0[0]),.doutb(w_n1814_0[1]),.din(n1814));
	jspl jspl_w_n1815_0(.douta(w_n1815_0[0]),.doutb(w_n1815_0[1]),.din(n1815));
	jspl jspl_w_n1816_0(.douta(w_n1816_0[0]),.doutb(w_n1816_0[1]),.din(n1816));
	jspl jspl_w_n1817_0(.douta(w_n1817_0[0]),.doutb(w_dff_A_xCr3eRnX3_1),.din(n1817));
	jspl jspl_w_n1824_0(.douta(w_n1824_0[0]),.doutb(w_n1824_0[1]),.din(n1824));
	jspl jspl_w_n1827_0(.douta(w_n1827_0[0]),.doutb(w_dff_A_tVLqk79Y1_1),.din(n1827));
	jspl jspl_w_n1828_0(.douta(w_n1828_0[0]),.doutb(w_n1828_0[1]),.din(w_dff_B_zHkCpcXH2_2));
	jspl jspl_w_n1829_0(.douta(w_n1829_0[0]),.doutb(w_n1829_0[1]),.din(w_dff_B_NK1gJBzJ7_2));
	jspl jspl_w_n1832_0(.douta(w_n1832_0[0]),.doutb(w_n1832_0[1]),.din(n1832));
	jspl jspl_w_n1834_0(.douta(w_n1834_0[0]),.doutb(w_n1834_0[1]),.din(n1834));
	jspl jspl_w_n1835_0(.douta(w_n1835_0[0]),.doutb(w_n1835_0[1]),.din(n1835));
	jspl jspl_w_n1836_0(.douta(w_n1836_0[0]),.doutb(w_dff_A_8XbjN7ht0_1),.din(n1836));
	jspl jspl_w_n1838_0(.douta(w_n1838_0[0]),.doutb(w_n1838_0[1]),.din(w_dff_B_wf5pirFW9_2));
	jspl jspl_w_n1841_0(.douta(w_n1841_0[0]),.doutb(w_n1841_0[1]),.din(n1841));
	jspl jspl_w_n1848_0(.douta(w_n1848_0[0]),.doutb(w_n1848_0[1]),.din(n1848));
	jspl jspl_w_n1849_0(.douta(w_dff_A_4LDx4qi96_0),.doutb(w_n1849_0[1]),.din(n1849));
	jdff dff_B_PQF7Q6RX4_1(.din(n67),.dout(w_dff_B_PQF7Q6RX4_1),.clk(gclk));
	jdff dff_B_KtM7KiYd4_1(.din(w_dff_B_PQF7Q6RX4_1),.dout(w_dff_B_KtM7KiYd4_1),.clk(gclk));
	jdff dff_B_ZhlSnPVz2_1(.din(n73),.dout(w_dff_B_ZhlSnPVz2_1),.clk(gclk));
	jdff dff_B_n8Hb1rcW9_1(.din(w_dff_B_ZhlSnPVz2_1),.dout(w_dff_B_n8Hb1rcW9_1),.clk(gclk));
	jdff dff_B_tyAKh0rM9_1(.din(n90),.dout(w_dff_B_tyAKh0rM9_1),.clk(gclk));
	jdff dff_B_WsfsLaUB1_1(.din(w_dff_B_tyAKh0rM9_1),.dout(w_dff_B_WsfsLaUB1_1),.clk(gclk));
	jdff dff_B_4zMmOsTM4_1(.din(w_dff_B_WsfsLaUB1_1),.dout(w_dff_B_4zMmOsTM4_1),.clk(gclk));
	jdff dff_B_IIdfHr4V5_1(.din(w_dff_B_4zMmOsTM4_1),.dout(w_dff_B_IIdfHr4V5_1),.clk(gclk));
	jdff dff_B_dN7aLtgt7_1(.din(w_dff_B_IIdfHr4V5_1),.dout(w_dff_B_dN7aLtgt7_1),.clk(gclk));
	jdff dff_B_6OiuCooY4_1(.din(w_dff_B_dN7aLtgt7_1),.dout(w_dff_B_6OiuCooY4_1),.clk(gclk));
	jdff dff_B_L1XRJyfl6_1(.din(n111),.dout(w_dff_B_L1XRJyfl6_1),.clk(gclk));
	jdff dff_B_ewIJIewB0_1(.din(w_dff_B_L1XRJyfl6_1),.dout(w_dff_B_ewIJIewB0_1),.clk(gclk));
	jdff dff_B_5FevXSI36_1(.din(w_dff_B_ewIJIewB0_1),.dout(w_dff_B_5FevXSI36_1),.clk(gclk));
	jdff dff_B_T589nlDk0_1(.din(w_dff_B_5FevXSI36_1),.dout(w_dff_B_T589nlDk0_1),.clk(gclk));
	jdff dff_B_ITxHWIIz4_1(.din(w_dff_B_T589nlDk0_1),.dout(w_dff_B_ITxHWIIz4_1),.clk(gclk));
	jdff dff_B_P9nnydua4_1(.din(w_dff_B_ITxHWIIz4_1),.dout(w_dff_B_P9nnydua4_1),.clk(gclk));
	jdff dff_B_UzsLI2Vz3_1(.din(w_dff_B_P9nnydua4_1),.dout(w_dff_B_UzsLI2Vz3_1),.clk(gclk));
	jdff dff_B_PGHqKmXo0_1(.din(w_dff_B_UzsLI2Vz3_1),.dout(w_dff_B_PGHqKmXo0_1),.clk(gclk));
	jdff dff_B_SWAZ2BU08_1(.din(w_dff_B_PGHqKmXo0_1),.dout(w_dff_B_SWAZ2BU08_1),.clk(gclk));
	jdff dff_B_YDVIK7HJ9_1(.din(n146),.dout(w_dff_B_YDVIK7HJ9_1),.clk(gclk));
	jdff dff_B_tUTiTzBA6_1(.din(w_dff_B_YDVIK7HJ9_1),.dout(w_dff_B_tUTiTzBA6_1),.clk(gclk));
	jdff dff_B_ui4FoLzg6_1(.din(w_dff_B_tUTiTzBA6_1),.dout(w_dff_B_ui4FoLzg6_1),.clk(gclk));
	jdff dff_B_ySHono3B3_1(.din(w_dff_B_ui4FoLzg6_1),.dout(w_dff_B_ySHono3B3_1),.clk(gclk));
	jdff dff_B_LLRp04ex6_1(.din(w_dff_B_ySHono3B3_1),.dout(w_dff_B_LLRp04ex6_1),.clk(gclk));
	jdff dff_B_uMwMbtXe6_1(.din(w_dff_B_LLRp04ex6_1),.dout(w_dff_B_uMwMbtXe6_1),.clk(gclk));
	jdff dff_B_3uSipkgl6_1(.din(w_dff_B_uMwMbtXe6_1),.dout(w_dff_B_3uSipkgl6_1),.clk(gclk));
	jdff dff_B_v6T5OL7j9_1(.din(w_dff_B_3uSipkgl6_1),.dout(w_dff_B_v6T5OL7j9_1),.clk(gclk));
	jdff dff_B_uknMZcEZ9_1(.din(w_dff_B_v6T5OL7j9_1),.dout(w_dff_B_uknMZcEZ9_1),.clk(gclk));
	jdff dff_B_eURwgZcN6_1(.din(w_dff_B_uknMZcEZ9_1),.dout(w_dff_B_eURwgZcN6_1),.clk(gclk));
	jdff dff_B_E0DEu2G33_1(.din(w_dff_B_eURwgZcN6_1),.dout(w_dff_B_E0DEu2G33_1),.clk(gclk));
	jdff dff_B_bbbPzB4b0_1(.din(n184),.dout(w_dff_B_bbbPzB4b0_1),.clk(gclk));
	jdff dff_B_LeVcw5oU6_1(.din(w_dff_B_bbbPzB4b0_1),.dout(w_dff_B_LeVcw5oU6_1),.clk(gclk));
	jdff dff_B_vhF2fbye6_1(.din(w_dff_B_LeVcw5oU6_1),.dout(w_dff_B_vhF2fbye6_1),.clk(gclk));
	jdff dff_B_wIIit61b4_1(.din(w_dff_B_vhF2fbye6_1),.dout(w_dff_B_wIIit61b4_1),.clk(gclk));
	jdff dff_B_jyGtYMSh1_1(.din(w_dff_B_wIIit61b4_1),.dout(w_dff_B_jyGtYMSh1_1),.clk(gclk));
	jdff dff_B_Dfq2bJFX0_1(.din(w_dff_B_jyGtYMSh1_1),.dout(w_dff_B_Dfq2bJFX0_1),.clk(gclk));
	jdff dff_B_V5S88XMb2_1(.din(w_dff_B_Dfq2bJFX0_1),.dout(w_dff_B_V5S88XMb2_1),.clk(gclk));
	jdff dff_B_1p1Cse915_1(.din(w_dff_B_V5S88XMb2_1),.dout(w_dff_B_1p1Cse915_1),.clk(gclk));
	jdff dff_B_zDe0Nk612_1(.din(w_dff_B_1p1Cse915_1),.dout(w_dff_B_zDe0Nk612_1),.clk(gclk));
	jdff dff_B_6DYlZ4Wv9_1(.din(w_dff_B_zDe0Nk612_1),.dout(w_dff_B_6DYlZ4Wv9_1),.clk(gclk));
	jdff dff_B_iGsyV5BJ5_1(.din(w_dff_B_6DYlZ4Wv9_1),.dout(w_dff_B_iGsyV5BJ5_1),.clk(gclk));
	jdff dff_B_2ngtrZm00_1(.din(w_dff_B_iGsyV5BJ5_1),.dout(w_dff_B_2ngtrZm00_1),.clk(gclk));
	jdff dff_B_Sw83mtes0_1(.din(w_dff_B_2ngtrZm00_1),.dout(w_dff_B_Sw83mtes0_1),.clk(gclk));
	jdff dff_B_Z8MvpjVb6_1(.din(n227),.dout(w_dff_B_Z8MvpjVb6_1),.clk(gclk));
	jdff dff_B_r0Zve7Jg2_1(.din(w_dff_B_Z8MvpjVb6_1),.dout(w_dff_B_r0Zve7Jg2_1),.clk(gclk));
	jdff dff_B_hUNLCFvr1_1(.din(w_dff_B_r0Zve7Jg2_1),.dout(w_dff_B_hUNLCFvr1_1),.clk(gclk));
	jdff dff_B_dhuJxHKp9_1(.din(w_dff_B_hUNLCFvr1_1),.dout(w_dff_B_dhuJxHKp9_1),.clk(gclk));
	jdff dff_B_vtWv7kPT5_1(.din(w_dff_B_dhuJxHKp9_1),.dout(w_dff_B_vtWv7kPT5_1),.clk(gclk));
	jdff dff_B_W6LWJoAP7_1(.din(w_dff_B_vtWv7kPT5_1),.dout(w_dff_B_W6LWJoAP7_1),.clk(gclk));
	jdff dff_B_5K7mlms61_1(.din(w_dff_B_W6LWJoAP7_1),.dout(w_dff_B_5K7mlms61_1),.clk(gclk));
	jdff dff_B_vx4ZBR9h3_1(.din(w_dff_B_5K7mlms61_1),.dout(w_dff_B_vx4ZBR9h3_1),.clk(gclk));
	jdff dff_B_c8xqwgbt5_1(.din(w_dff_B_vx4ZBR9h3_1),.dout(w_dff_B_c8xqwgbt5_1),.clk(gclk));
	jdff dff_B_feWmIk1f7_1(.din(w_dff_B_c8xqwgbt5_1),.dout(w_dff_B_feWmIk1f7_1),.clk(gclk));
	jdff dff_B_06xoIY8R8_1(.din(w_dff_B_feWmIk1f7_1),.dout(w_dff_B_06xoIY8R8_1),.clk(gclk));
	jdff dff_B_o0ef297I6_1(.din(w_dff_B_06xoIY8R8_1),.dout(w_dff_B_o0ef297I6_1),.clk(gclk));
	jdff dff_B_zKtuICp35_1(.din(w_dff_B_o0ef297I6_1),.dout(w_dff_B_zKtuICp35_1),.clk(gclk));
	jdff dff_B_n45O0EvX2_1(.din(w_dff_B_zKtuICp35_1),.dout(w_dff_B_n45O0EvX2_1),.clk(gclk));
	jdff dff_B_4vAet7Rm0_1(.din(w_dff_B_n45O0EvX2_1),.dout(w_dff_B_4vAet7Rm0_1),.clk(gclk));
	jdff dff_B_r0SBWScu0_1(.din(n278),.dout(w_dff_B_r0SBWScu0_1),.clk(gclk));
	jdff dff_B_Dat5FnZs1_1(.din(w_dff_B_r0SBWScu0_1),.dout(w_dff_B_Dat5FnZs1_1),.clk(gclk));
	jdff dff_B_vzjHGODt0_1(.din(w_dff_B_Dat5FnZs1_1),.dout(w_dff_B_vzjHGODt0_1),.clk(gclk));
	jdff dff_B_z0CsdEBV7_1(.din(w_dff_B_vzjHGODt0_1),.dout(w_dff_B_z0CsdEBV7_1),.clk(gclk));
	jdff dff_B_nH2cGjvr9_1(.din(w_dff_B_z0CsdEBV7_1),.dout(w_dff_B_nH2cGjvr9_1),.clk(gclk));
	jdff dff_B_G0HqAf2U0_1(.din(w_dff_B_nH2cGjvr9_1),.dout(w_dff_B_G0HqAf2U0_1),.clk(gclk));
	jdff dff_B_fB4GnBQG1_1(.din(w_dff_B_G0HqAf2U0_1),.dout(w_dff_B_fB4GnBQG1_1),.clk(gclk));
	jdff dff_B_UJBZ8oSg8_1(.din(w_dff_B_fB4GnBQG1_1),.dout(w_dff_B_UJBZ8oSg8_1),.clk(gclk));
	jdff dff_B_1Mj7QbrO3_1(.din(w_dff_B_UJBZ8oSg8_1),.dout(w_dff_B_1Mj7QbrO3_1),.clk(gclk));
	jdff dff_B_w6z4SHnv8_1(.din(w_dff_B_1Mj7QbrO3_1),.dout(w_dff_B_w6z4SHnv8_1),.clk(gclk));
	jdff dff_B_Poxu68YB1_1(.din(w_dff_B_w6z4SHnv8_1),.dout(w_dff_B_Poxu68YB1_1),.clk(gclk));
	jdff dff_B_XUl1sJoD8_1(.din(w_dff_B_Poxu68YB1_1),.dout(w_dff_B_XUl1sJoD8_1),.clk(gclk));
	jdff dff_B_D52GB4AA8_1(.din(w_dff_B_XUl1sJoD8_1),.dout(w_dff_B_D52GB4AA8_1),.clk(gclk));
	jdff dff_B_vLZ0Rvma7_1(.din(w_dff_B_D52GB4AA8_1),.dout(w_dff_B_vLZ0Rvma7_1),.clk(gclk));
	jdff dff_B_DxoX74Ss2_1(.din(w_dff_B_vLZ0Rvma7_1),.dout(w_dff_B_DxoX74Ss2_1),.clk(gclk));
	jdff dff_B_eGrZTmfC4_1(.din(w_dff_B_DxoX74Ss2_1),.dout(w_dff_B_eGrZTmfC4_1),.clk(gclk));
	jdff dff_B_ckDZ6xwe5_1(.din(w_dff_B_eGrZTmfC4_1),.dout(w_dff_B_ckDZ6xwe5_1),.clk(gclk));
	jdff dff_B_DAPtb3rX3_1(.din(n336),.dout(w_dff_B_DAPtb3rX3_1),.clk(gclk));
	jdff dff_B_TDQN3faj4_1(.din(w_dff_B_DAPtb3rX3_1),.dout(w_dff_B_TDQN3faj4_1),.clk(gclk));
	jdff dff_B_s6ltvAk54_1(.din(w_dff_B_TDQN3faj4_1),.dout(w_dff_B_s6ltvAk54_1),.clk(gclk));
	jdff dff_B_Rfj5erp36_1(.din(w_dff_B_s6ltvAk54_1),.dout(w_dff_B_Rfj5erp36_1),.clk(gclk));
	jdff dff_B_CrmQpBIN3_1(.din(w_dff_B_Rfj5erp36_1),.dout(w_dff_B_CrmQpBIN3_1),.clk(gclk));
	jdff dff_B_M4qU9Zaz6_1(.din(w_dff_B_CrmQpBIN3_1),.dout(w_dff_B_M4qU9Zaz6_1),.clk(gclk));
	jdff dff_B_8kJdTjWl0_1(.din(w_dff_B_M4qU9Zaz6_1),.dout(w_dff_B_8kJdTjWl0_1),.clk(gclk));
	jdff dff_B_wgDUeidg0_1(.din(w_dff_B_8kJdTjWl0_1),.dout(w_dff_B_wgDUeidg0_1),.clk(gclk));
	jdff dff_B_izKSgGRD5_1(.din(w_dff_B_wgDUeidg0_1),.dout(w_dff_B_izKSgGRD5_1),.clk(gclk));
	jdff dff_B_scuaBA3P9_1(.din(w_dff_B_izKSgGRD5_1),.dout(w_dff_B_scuaBA3P9_1),.clk(gclk));
	jdff dff_B_2MTZeLR83_1(.din(w_dff_B_scuaBA3P9_1),.dout(w_dff_B_2MTZeLR83_1),.clk(gclk));
	jdff dff_B_he08mcgy3_1(.din(w_dff_B_2MTZeLR83_1),.dout(w_dff_B_he08mcgy3_1),.clk(gclk));
	jdff dff_B_oXdXZ9bt8_1(.din(w_dff_B_he08mcgy3_1),.dout(w_dff_B_oXdXZ9bt8_1),.clk(gclk));
	jdff dff_B_vZmFHDus3_1(.din(w_dff_B_oXdXZ9bt8_1),.dout(w_dff_B_vZmFHDus3_1),.clk(gclk));
	jdff dff_B_9PrurzBw9_1(.din(w_dff_B_vZmFHDus3_1),.dout(w_dff_B_9PrurzBw9_1),.clk(gclk));
	jdff dff_B_Xsncoxn68_1(.din(w_dff_B_9PrurzBw9_1),.dout(w_dff_B_Xsncoxn68_1),.clk(gclk));
	jdff dff_B_uUOFw2py4_1(.din(w_dff_B_Xsncoxn68_1),.dout(w_dff_B_uUOFw2py4_1),.clk(gclk));
	jdff dff_B_iyDyi3uF1_1(.din(w_dff_B_uUOFw2py4_1),.dout(w_dff_B_iyDyi3uF1_1),.clk(gclk));
	jdff dff_B_NUgGDnyd1_1(.din(w_dff_B_iyDyi3uF1_1),.dout(w_dff_B_NUgGDnyd1_1),.clk(gclk));
	jdff dff_B_ALDGzlgO8_1(.din(n400),.dout(w_dff_B_ALDGzlgO8_1),.clk(gclk));
	jdff dff_B_O8vCVjGT1_1(.din(w_dff_B_ALDGzlgO8_1),.dout(w_dff_B_O8vCVjGT1_1),.clk(gclk));
	jdff dff_B_5GsazEe12_1(.din(w_dff_B_O8vCVjGT1_1),.dout(w_dff_B_5GsazEe12_1),.clk(gclk));
	jdff dff_B_nh6LaOd71_1(.din(w_dff_B_5GsazEe12_1),.dout(w_dff_B_nh6LaOd71_1),.clk(gclk));
	jdff dff_B_L1D3PMEI3_1(.din(w_dff_B_nh6LaOd71_1),.dout(w_dff_B_L1D3PMEI3_1),.clk(gclk));
	jdff dff_B_t9FAN2uM4_1(.din(w_dff_B_L1D3PMEI3_1),.dout(w_dff_B_t9FAN2uM4_1),.clk(gclk));
	jdff dff_B_DFGKUIJD6_1(.din(w_dff_B_t9FAN2uM4_1),.dout(w_dff_B_DFGKUIJD6_1),.clk(gclk));
	jdff dff_B_JiFa466S7_1(.din(w_dff_B_DFGKUIJD6_1),.dout(w_dff_B_JiFa466S7_1),.clk(gclk));
	jdff dff_B_iI0ubWry5_1(.din(w_dff_B_JiFa466S7_1),.dout(w_dff_B_iI0ubWry5_1),.clk(gclk));
	jdff dff_B_4VllvIFq9_1(.din(w_dff_B_iI0ubWry5_1),.dout(w_dff_B_4VllvIFq9_1),.clk(gclk));
	jdff dff_B_bIUygaES4_1(.din(w_dff_B_4VllvIFq9_1),.dout(w_dff_B_bIUygaES4_1),.clk(gclk));
	jdff dff_B_e5D5TEC86_1(.din(w_dff_B_bIUygaES4_1),.dout(w_dff_B_e5D5TEC86_1),.clk(gclk));
	jdff dff_B_IEq2NRb70_1(.din(w_dff_B_e5D5TEC86_1),.dout(w_dff_B_IEq2NRb70_1),.clk(gclk));
	jdff dff_B_N06wAm8V0_1(.din(w_dff_B_IEq2NRb70_1),.dout(w_dff_B_N06wAm8V0_1),.clk(gclk));
	jdff dff_B_Fg3Z1WeT2_1(.din(w_dff_B_N06wAm8V0_1),.dout(w_dff_B_Fg3Z1WeT2_1),.clk(gclk));
	jdff dff_B_SLiO93it0_1(.din(w_dff_B_Fg3Z1WeT2_1),.dout(w_dff_B_SLiO93it0_1),.clk(gclk));
	jdff dff_B_uxgDp7VQ5_1(.din(w_dff_B_SLiO93it0_1),.dout(w_dff_B_uxgDp7VQ5_1),.clk(gclk));
	jdff dff_B_iz5nuxgg5_1(.din(w_dff_B_uxgDp7VQ5_1),.dout(w_dff_B_iz5nuxgg5_1),.clk(gclk));
	jdff dff_B_eCr8oSLu9_1(.din(w_dff_B_iz5nuxgg5_1),.dout(w_dff_B_eCr8oSLu9_1),.clk(gclk));
	jdff dff_B_sHMTP3JT9_1(.din(w_dff_B_eCr8oSLu9_1),.dout(w_dff_B_sHMTP3JT9_1),.clk(gclk));
	jdff dff_B_krulCJ8w6_1(.din(w_dff_B_sHMTP3JT9_1),.dout(w_dff_B_krulCJ8w6_1),.clk(gclk));
	jdff dff_B_AavzEL6p4_1(.din(n472),.dout(w_dff_B_AavzEL6p4_1),.clk(gclk));
	jdff dff_B_kZartvYS2_1(.din(w_dff_B_AavzEL6p4_1),.dout(w_dff_B_kZartvYS2_1),.clk(gclk));
	jdff dff_B_UdHEuSoE9_1(.din(w_dff_B_kZartvYS2_1),.dout(w_dff_B_UdHEuSoE9_1),.clk(gclk));
	jdff dff_B_kqLUVLYO5_1(.din(w_dff_B_UdHEuSoE9_1),.dout(w_dff_B_kqLUVLYO5_1),.clk(gclk));
	jdff dff_B_VJ7UVoaq8_1(.din(w_dff_B_kqLUVLYO5_1),.dout(w_dff_B_VJ7UVoaq8_1),.clk(gclk));
	jdff dff_B_nWm8VPZz1_1(.din(w_dff_B_VJ7UVoaq8_1),.dout(w_dff_B_nWm8VPZz1_1),.clk(gclk));
	jdff dff_B_UTZptcMV7_1(.din(w_dff_B_nWm8VPZz1_1),.dout(w_dff_B_UTZptcMV7_1),.clk(gclk));
	jdff dff_B_nMtdLqfT1_1(.din(w_dff_B_UTZptcMV7_1),.dout(w_dff_B_nMtdLqfT1_1),.clk(gclk));
	jdff dff_B_XPZJBQ403_1(.din(w_dff_B_nMtdLqfT1_1),.dout(w_dff_B_XPZJBQ403_1),.clk(gclk));
	jdff dff_B_cjVju64M6_1(.din(w_dff_B_XPZJBQ403_1),.dout(w_dff_B_cjVju64M6_1),.clk(gclk));
	jdff dff_B_0Rpqzsbc9_1(.din(w_dff_B_cjVju64M6_1),.dout(w_dff_B_0Rpqzsbc9_1),.clk(gclk));
	jdff dff_B_GjoYfDdN6_1(.din(w_dff_B_0Rpqzsbc9_1),.dout(w_dff_B_GjoYfDdN6_1),.clk(gclk));
	jdff dff_B_g8md13Eg7_1(.din(w_dff_B_GjoYfDdN6_1),.dout(w_dff_B_g8md13Eg7_1),.clk(gclk));
	jdff dff_B_Vu8awZTy1_1(.din(w_dff_B_g8md13Eg7_1),.dout(w_dff_B_Vu8awZTy1_1),.clk(gclk));
	jdff dff_B_DllI2f9q3_1(.din(w_dff_B_Vu8awZTy1_1),.dout(w_dff_B_DllI2f9q3_1),.clk(gclk));
	jdff dff_B_PwDdCmLD6_1(.din(w_dff_B_DllI2f9q3_1),.dout(w_dff_B_PwDdCmLD6_1),.clk(gclk));
	jdff dff_B_0a6wVlJl0_1(.din(w_dff_B_PwDdCmLD6_1),.dout(w_dff_B_0a6wVlJl0_1),.clk(gclk));
	jdff dff_B_9jkkDO0J3_1(.din(w_dff_B_0a6wVlJl0_1),.dout(w_dff_B_9jkkDO0J3_1),.clk(gclk));
	jdff dff_B_qVpRfhja7_1(.din(w_dff_B_9jkkDO0J3_1),.dout(w_dff_B_qVpRfhja7_1),.clk(gclk));
	jdff dff_B_unKqxwCw0_1(.din(w_dff_B_qVpRfhja7_1),.dout(w_dff_B_unKqxwCw0_1),.clk(gclk));
	jdff dff_B_jhY0Ph468_1(.din(w_dff_B_unKqxwCw0_1),.dout(w_dff_B_jhY0Ph468_1),.clk(gclk));
	jdff dff_B_a0YYHObV4_1(.din(w_dff_B_jhY0Ph468_1),.dout(w_dff_B_a0YYHObV4_1),.clk(gclk));
	jdff dff_B_YaDzBe1T8_1(.din(w_dff_B_a0YYHObV4_1),.dout(w_dff_B_YaDzBe1T8_1),.clk(gclk));
	jdff dff_B_NTnK2NtP3_1(.din(n551),.dout(w_dff_B_NTnK2NtP3_1),.clk(gclk));
	jdff dff_B_WyUmnwOy7_1(.din(w_dff_B_NTnK2NtP3_1),.dout(w_dff_B_WyUmnwOy7_1),.clk(gclk));
	jdff dff_B_9MvVc6vA5_1(.din(w_dff_B_WyUmnwOy7_1),.dout(w_dff_B_9MvVc6vA5_1),.clk(gclk));
	jdff dff_B_Ix4TDhKO8_1(.din(w_dff_B_9MvVc6vA5_1),.dout(w_dff_B_Ix4TDhKO8_1),.clk(gclk));
	jdff dff_B_1jI5rYFJ7_1(.din(w_dff_B_Ix4TDhKO8_1),.dout(w_dff_B_1jI5rYFJ7_1),.clk(gclk));
	jdff dff_B_AKd3WrEr1_1(.din(w_dff_B_1jI5rYFJ7_1),.dout(w_dff_B_AKd3WrEr1_1),.clk(gclk));
	jdff dff_B_IeL3uRB35_1(.din(w_dff_B_AKd3WrEr1_1),.dout(w_dff_B_IeL3uRB35_1),.clk(gclk));
	jdff dff_B_4wyENoWV7_1(.din(w_dff_B_IeL3uRB35_1),.dout(w_dff_B_4wyENoWV7_1),.clk(gclk));
	jdff dff_B_ahkEcgPM9_1(.din(w_dff_B_4wyENoWV7_1),.dout(w_dff_B_ahkEcgPM9_1),.clk(gclk));
	jdff dff_B_t9KF2QBM8_1(.din(w_dff_B_ahkEcgPM9_1),.dout(w_dff_B_t9KF2QBM8_1),.clk(gclk));
	jdff dff_B_unEBqfAa7_1(.din(w_dff_B_t9KF2QBM8_1),.dout(w_dff_B_unEBqfAa7_1),.clk(gclk));
	jdff dff_B_4waMXeIV3_1(.din(w_dff_B_unEBqfAa7_1),.dout(w_dff_B_4waMXeIV3_1),.clk(gclk));
	jdff dff_B_lGUKKiul8_1(.din(w_dff_B_4waMXeIV3_1),.dout(w_dff_B_lGUKKiul8_1),.clk(gclk));
	jdff dff_B_anFrpBVE5_1(.din(w_dff_B_lGUKKiul8_1),.dout(w_dff_B_anFrpBVE5_1),.clk(gclk));
	jdff dff_B_kVykFfvG2_1(.din(w_dff_B_anFrpBVE5_1),.dout(w_dff_B_kVykFfvG2_1),.clk(gclk));
	jdff dff_B_eD1xd3qJ0_1(.din(w_dff_B_kVykFfvG2_1),.dout(w_dff_B_eD1xd3qJ0_1),.clk(gclk));
	jdff dff_B_NBaIixZQ1_1(.din(w_dff_B_eD1xd3qJ0_1),.dout(w_dff_B_NBaIixZQ1_1),.clk(gclk));
	jdff dff_B_ckYCSpSo5_1(.din(w_dff_B_NBaIixZQ1_1),.dout(w_dff_B_ckYCSpSo5_1),.clk(gclk));
	jdff dff_B_oGirlH2C2_1(.din(w_dff_B_ckYCSpSo5_1),.dout(w_dff_B_oGirlH2C2_1),.clk(gclk));
	jdff dff_B_vyeF3mPc5_1(.din(w_dff_B_oGirlH2C2_1),.dout(w_dff_B_vyeF3mPc5_1),.clk(gclk));
	jdff dff_B_mW0PzjL71_1(.din(w_dff_B_vyeF3mPc5_1),.dout(w_dff_B_mW0PzjL71_1),.clk(gclk));
	jdff dff_B_l9DJG3cU7_1(.din(w_dff_B_mW0PzjL71_1),.dout(w_dff_B_l9DJG3cU7_1),.clk(gclk));
	jdff dff_B_wVCT7QOs7_1(.din(w_dff_B_l9DJG3cU7_1),.dout(w_dff_B_wVCT7QOs7_1),.clk(gclk));
	jdff dff_B_FEvEN3zF4_1(.din(w_dff_B_wVCT7QOs7_1),.dout(w_dff_B_FEvEN3zF4_1),.clk(gclk));
	jdff dff_B_1YwacAhb1_1(.din(w_dff_B_FEvEN3zF4_1),.dout(w_dff_B_1YwacAhb1_1),.clk(gclk));
	jdff dff_B_2HahP3lz4_1(.din(n637),.dout(w_dff_B_2HahP3lz4_1),.clk(gclk));
	jdff dff_B_ALkpca9E8_1(.din(w_dff_B_2HahP3lz4_1),.dout(w_dff_B_ALkpca9E8_1),.clk(gclk));
	jdff dff_B_vpKDqYVp1_1(.din(w_dff_B_ALkpca9E8_1),.dout(w_dff_B_vpKDqYVp1_1),.clk(gclk));
	jdff dff_B_1BqohqWW9_1(.din(w_dff_B_vpKDqYVp1_1),.dout(w_dff_B_1BqohqWW9_1),.clk(gclk));
	jdff dff_B_jPJRe2Vx1_1(.din(w_dff_B_1BqohqWW9_1),.dout(w_dff_B_jPJRe2Vx1_1),.clk(gclk));
	jdff dff_B_OWW048zC0_1(.din(w_dff_B_jPJRe2Vx1_1),.dout(w_dff_B_OWW048zC0_1),.clk(gclk));
	jdff dff_B_0nC3Wfly4_1(.din(w_dff_B_OWW048zC0_1),.dout(w_dff_B_0nC3Wfly4_1),.clk(gclk));
	jdff dff_B_1LKBOgen3_1(.din(w_dff_B_0nC3Wfly4_1),.dout(w_dff_B_1LKBOgen3_1),.clk(gclk));
	jdff dff_B_aLB2d8Cb4_1(.din(w_dff_B_1LKBOgen3_1),.dout(w_dff_B_aLB2d8Cb4_1),.clk(gclk));
	jdff dff_B_nKA0yp2Q2_1(.din(w_dff_B_aLB2d8Cb4_1),.dout(w_dff_B_nKA0yp2Q2_1),.clk(gclk));
	jdff dff_B_cGBd3OA87_1(.din(w_dff_B_nKA0yp2Q2_1),.dout(w_dff_B_cGBd3OA87_1),.clk(gclk));
	jdff dff_B_emieqirN9_1(.din(w_dff_B_cGBd3OA87_1),.dout(w_dff_B_emieqirN9_1),.clk(gclk));
	jdff dff_B_SG3P9x418_1(.din(w_dff_B_emieqirN9_1),.dout(w_dff_B_SG3P9x418_1),.clk(gclk));
	jdff dff_B_iHytJvjV4_1(.din(w_dff_B_SG3P9x418_1),.dout(w_dff_B_iHytJvjV4_1),.clk(gclk));
	jdff dff_B_hlPpaA698_1(.din(w_dff_B_iHytJvjV4_1),.dout(w_dff_B_hlPpaA698_1),.clk(gclk));
	jdff dff_B_MrbNIMoq6_1(.din(w_dff_B_hlPpaA698_1),.dout(w_dff_B_MrbNIMoq6_1),.clk(gclk));
	jdff dff_B_7A63QXBg4_1(.din(w_dff_B_MrbNIMoq6_1),.dout(w_dff_B_7A63QXBg4_1),.clk(gclk));
	jdff dff_B_g4EDgwar7_1(.din(w_dff_B_7A63QXBg4_1),.dout(w_dff_B_g4EDgwar7_1),.clk(gclk));
	jdff dff_B_1khOGrGO3_1(.din(w_dff_B_g4EDgwar7_1),.dout(w_dff_B_1khOGrGO3_1),.clk(gclk));
	jdff dff_B_u7yeBYl67_1(.din(w_dff_B_1khOGrGO3_1),.dout(w_dff_B_u7yeBYl67_1),.clk(gclk));
	jdff dff_B_O338R50T0_1(.din(w_dff_B_u7yeBYl67_1),.dout(w_dff_B_O338R50T0_1),.clk(gclk));
	jdff dff_B_eKx4aCcY1_1(.din(w_dff_B_O338R50T0_1),.dout(w_dff_B_eKx4aCcY1_1),.clk(gclk));
	jdff dff_B_pUV2rRbI9_1(.din(w_dff_B_eKx4aCcY1_1),.dout(w_dff_B_pUV2rRbI9_1),.clk(gclk));
	jdff dff_B_G6O3ndkp0_1(.din(w_dff_B_pUV2rRbI9_1),.dout(w_dff_B_G6O3ndkp0_1),.clk(gclk));
	jdff dff_B_jtLOVUAj2_1(.din(w_dff_B_G6O3ndkp0_1),.dout(w_dff_B_jtLOVUAj2_1),.clk(gclk));
	jdff dff_B_pj2vplUu7_1(.din(w_dff_B_jtLOVUAj2_1),.dout(w_dff_B_pj2vplUu7_1),.clk(gclk));
	jdff dff_B_eX2PGYRO6_1(.din(w_dff_B_pj2vplUu7_1),.dout(w_dff_B_eX2PGYRO6_1),.clk(gclk));
	jdff dff_B_fxTGXImx7_1(.din(n730),.dout(w_dff_B_fxTGXImx7_1),.clk(gclk));
	jdff dff_B_wsa85A8K3_1(.din(w_dff_B_fxTGXImx7_1),.dout(w_dff_B_wsa85A8K3_1),.clk(gclk));
	jdff dff_B_denECjb90_1(.din(w_dff_B_wsa85A8K3_1),.dout(w_dff_B_denECjb90_1),.clk(gclk));
	jdff dff_B_GIAdrbyx3_1(.din(w_dff_B_denECjb90_1),.dout(w_dff_B_GIAdrbyx3_1),.clk(gclk));
	jdff dff_B_gOnLd4tl9_1(.din(w_dff_B_GIAdrbyx3_1),.dout(w_dff_B_gOnLd4tl9_1),.clk(gclk));
	jdff dff_B_zQyoQ6Te9_1(.din(w_dff_B_gOnLd4tl9_1),.dout(w_dff_B_zQyoQ6Te9_1),.clk(gclk));
	jdff dff_B_OFwx75Pl9_1(.din(w_dff_B_zQyoQ6Te9_1),.dout(w_dff_B_OFwx75Pl9_1),.clk(gclk));
	jdff dff_B_rNN6RNev1_1(.din(w_dff_B_OFwx75Pl9_1),.dout(w_dff_B_rNN6RNev1_1),.clk(gclk));
	jdff dff_B_I2rDsrrO3_1(.din(w_dff_B_rNN6RNev1_1),.dout(w_dff_B_I2rDsrrO3_1),.clk(gclk));
	jdff dff_B_2AqFPdcb4_1(.din(w_dff_B_I2rDsrrO3_1),.dout(w_dff_B_2AqFPdcb4_1),.clk(gclk));
	jdff dff_B_4jyacbdo2_1(.din(w_dff_B_2AqFPdcb4_1),.dout(w_dff_B_4jyacbdo2_1),.clk(gclk));
	jdff dff_B_j6aJq50u4_1(.din(w_dff_B_4jyacbdo2_1),.dout(w_dff_B_j6aJq50u4_1),.clk(gclk));
	jdff dff_B_DRoZUYa66_1(.din(w_dff_B_j6aJq50u4_1),.dout(w_dff_B_DRoZUYa66_1),.clk(gclk));
	jdff dff_B_x81I4trF5_1(.din(w_dff_B_DRoZUYa66_1),.dout(w_dff_B_x81I4trF5_1),.clk(gclk));
	jdff dff_B_HUpk6K9F6_1(.din(w_dff_B_x81I4trF5_1),.dout(w_dff_B_HUpk6K9F6_1),.clk(gclk));
	jdff dff_B_aWNqCJgB3_1(.din(w_dff_B_HUpk6K9F6_1),.dout(w_dff_B_aWNqCJgB3_1),.clk(gclk));
	jdff dff_B_8IJFiap96_1(.din(w_dff_B_aWNqCJgB3_1),.dout(w_dff_B_8IJFiap96_1),.clk(gclk));
	jdff dff_B_t8C0qdVd1_1(.din(w_dff_B_8IJFiap96_1),.dout(w_dff_B_t8C0qdVd1_1),.clk(gclk));
	jdff dff_B_m85cgeEn7_1(.din(w_dff_B_t8C0qdVd1_1),.dout(w_dff_B_m85cgeEn7_1),.clk(gclk));
	jdff dff_B_E46jhpQJ3_1(.din(w_dff_B_m85cgeEn7_1),.dout(w_dff_B_E46jhpQJ3_1),.clk(gclk));
	jdff dff_B_6hfu1Ynt7_1(.din(w_dff_B_E46jhpQJ3_1),.dout(w_dff_B_6hfu1Ynt7_1),.clk(gclk));
	jdff dff_B_OAg5oLId0_1(.din(w_dff_B_6hfu1Ynt7_1),.dout(w_dff_B_OAg5oLId0_1),.clk(gclk));
	jdff dff_B_3NDNqwgc9_1(.din(w_dff_B_OAg5oLId0_1),.dout(w_dff_B_3NDNqwgc9_1),.clk(gclk));
	jdff dff_B_T0euW1FQ9_1(.din(w_dff_B_3NDNqwgc9_1),.dout(w_dff_B_T0euW1FQ9_1),.clk(gclk));
	jdff dff_B_TSmMUTFN5_1(.din(w_dff_B_T0euW1FQ9_1),.dout(w_dff_B_TSmMUTFN5_1),.clk(gclk));
	jdff dff_B_XOPU4qWo7_1(.din(w_dff_B_TSmMUTFN5_1),.dout(w_dff_B_XOPU4qWo7_1),.clk(gclk));
	jdff dff_B_Gxo9BsDJ1_1(.din(w_dff_B_XOPU4qWo7_1),.dout(w_dff_B_Gxo9BsDJ1_1),.clk(gclk));
	jdff dff_B_iiCDqQwQ1_1(.din(w_dff_B_Gxo9BsDJ1_1),.dout(w_dff_B_iiCDqQwQ1_1),.clk(gclk));
	jdff dff_B_aoYzFfpI1_1(.din(w_dff_B_iiCDqQwQ1_1),.dout(w_dff_B_aoYzFfpI1_1),.clk(gclk));
	jdff dff_B_ysdfaLGG4_1(.din(n830),.dout(w_dff_B_ysdfaLGG4_1),.clk(gclk));
	jdff dff_B_zUd21HmB0_1(.din(w_dff_B_ysdfaLGG4_1),.dout(w_dff_B_zUd21HmB0_1),.clk(gclk));
	jdff dff_B_6PNyvwsl7_1(.din(w_dff_B_zUd21HmB0_1),.dout(w_dff_B_6PNyvwsl7_1),.clk(gclk));
	jdff dff_B_gCuY30CU1_1(.din(w_dff_B_6PNyvwsl7_1),.dout(w_dff_B_gCuY30CU1_1),.clk(gclk));
	jdff dff_B_UjBoxxR33_1(.din(w_dff_B_gCuY30CU1_1),.dout(w_dff_B_UjBoxxR33_1),.clk(gclk));
	jdff dff_B_FBqPp71W6_1(.din(w_dff_B_UjBoxxR33_1),.dout(w_dff_B_FBqPp71W6_1),.clk(gclk));
	jdff dff_B_MTrjtqdF6_1(.din(w_dff_B_FBqPp71W6_1),.dout(w_dff_B_MTrjtqdF6_1),.clk(gclk));
	jdff dff_B_w9AViUWg5_1(.din(w_dff_B_MTrjtqdF6_1),.dout(w_dff_B_w9AViUWg5_1),.clk(gclk));
	jdff dff_B_lyThDFEn0_1(.din(w_dff_B_w9AViUWg5_1),.dout(w_dff_B_lyThDFEn0_1),.clk(gclk));
	jdff dff_B_aiNMS3tv8_1(.din(w_dff_B_lyThDFEn0_1),.dout(w_dff_B_aiNMS3tv8_1),.clk(gclk));
	jdff dff_B_EYClND6P2_1(.din(w_dff_B_aiNMS3tv8_1),.dout(w_dff_B_EYClND6P2_1),.clk(gclk));
	jdff dff_B_qpm4qKSr6_1(.din(w_dff_B_EYClND6P2_1),.dout(w_dff_B_qpm4qKSr6_1),.clk(gclk));
	jdff dff_B_ssHNVFP55_1(.din(w_dff_B_qpm4qKSr6_1),.dout(w_dff_B_ssHNVFP55_1),.clk(gclk));
	jdff dff_B_fMk88tCc9_1(.din(w_dff_B_ssHNVFP55_1),.dout(w_dff_B_fMk88tCc9_1),.clk(gclk));
	jdff dff_B_s1iXvth84_1(.din(w_dff_B_fMk88tCc9_1),.dout(w_dff_B_s1iXvth84_1),.clk(gclk));
	jdff dff_B_VmsowpXG4_1(.din(w_dff_B_s1iXvth84_1),.dout(w_dff_B_VmsowpXG4_1),.clk(gclk));
	jdff dff_B_Lg2vOnfW8_1(.din(w_dff_B_VmsowpXG4_1),.dout(w_dff_B_Lg2vOnfW8_1),.clk(gclk));
	jdff dff_B_yREOMLlg4_1(.din(w_dff_B_Lg2vOnfW8_1),.dout(w_dff_B_yREOMLlg4_1),.clk(gclk));
	jdff dff_B_VBlac2Zm9_1(.din(w_dff_B_yREOMLlg4_1),.dout(w_dff_B_VBlac2Zm9_1),.clk(gclk));
	jdff dff_B_cUcqEIWm3_1(.din(w_dff_B_VBlac2Zm9_1),.dout(w_dff_B_cUcqEIWm3_1),.clk(gclk));
	jdff dff_B_bEaYfO6w2_1(.din(w_dff_B_cUcqEIWm3_1),.dout(w_dff_B_bEaYfO6w2_1),.clk(gclk));
	jdff dff_B_XgPKrEHh5_1(.din(w_dff_B_bEaYfO6w2_1),.dout(w_dff_B_XgPKrEHh5_1),.clk(gclk));
	jdff dff_B_gsqPlIZq8_1(.din(w_dff_B_XgPKrEHh5_1),.dout(w_dff_B_gsqPlIZq8_1),.clk(gclk));
	jdff dff_B_YlZ1ifuY9_1(.din(w_dff_B_gsqPlIZq8_1),.dout(w_dff_B_YlZ1ifuY9_1),.clk(gclk));
	jdff dff_B_ll7mHaFn4_1(.din(w_dff_B_YlZ1ifuY9_1),.dout(w_dff_B_ll7mHaFn4_1),.clk(gclk));
	jdff dff_B_Ooq4ibow1_1(.din(w_dff_B_ll7mHaFn4_1),.dout(w_dff_B_Ooq4ibow1_1),.clk(gclk));
	jdff dff_B_r41isFue8_1(.din(w_dff_B_Ooq4ibow1_1),.dout(w_dff_B_r41isFue8_1),.clk(gclk));
	jdff dff_B_9p9bTvwe7_1(.din(w_dff_B_r41isFue8_1),.dout(w_dff_B_9p9bTvwe7_1),.clk(gclk));
	jdff dff_B_jwaiEsGo8_1(.din(w_dff_B_9p9bTvwe7_1),.dout(w_dff_B_jwaiEsGo8_1),.clk(gclk));
	jdff dff_B_HqmVv85Q0_1(.din(w_dff_B_jwaiEsGo8_1),.dout(w_dff_B_HqmVv85Q0_1),.clk(gclk));
	jdff dff_B_E6U2roQ78_1(.din(w_dff_B_HqmVv85Q0_1),.dout(w_dff_B_E6U2roQ78_1),.clk(gclk));
	jdff dff_B_ZmNJV0mi8_1(.din(n1842),.dout(w_dff_B_ZmNJV0mi8_1),.clk(gclk));
	jdff dff_B_A8i5BUFm4_1(.din(w_dff_B_ZmNJV0mi8_1),.dout(w_dff_B_A8i5BUFm4_1),.clk(gclk));
	jdff dff_B_A3nvCzqV6_1(.din(w_dff_B_A8i5BUFm4_1),.dout(w_dff_B_A3nvCzqV6_1),.clk(gclk));
	jdff dff_B_LAlxv1ln5_1(.din(w_dff_B_A3nvCzqV6_1),.dout(w_dff_B_LAlxv1ln5_1),.clk(gclk));
	jdff dff_B_jLMa77NH2_1(.din(w_dff_B_LAlxv1ln5_1),.dout(w_dff_B_jLMa77NH2_1),.clk(gclk));
	jdff dff_B_J5pjl8qY0_0(.din(n1850),.dout(w_dff_B_J5pjl8qY0_0),.clk(gclk));
	jdff dff_B_J6XJFA6V4_0(.din(w_dff_B_J5pjl8qY0_0),.dout(w_dff_B_J6XJFA6V4_0),.clk(gclk));
	jdff dff_B_Lx61Oscp4_0(.din(w_dff_B_J6XJFA6V4_0),.dout(w_dff_B_Lx61Oscp4_0),.clk(gclk));
	jdff dff_A_CEbSgHrH1_0(.dout(w_n1849_0[0]),.din(w_dff_A_CEbSgHrH1_0),.clk(gclk));
	jdff dff_A_LcoIPl2v9_0(.dout(w_dff_A_CEbSgHrH1_0),.din(w_dff_A_LcoIPl2v9_0),.clk(gclk));
	jdff dff_A_colYvOkg3_0(.dout(w_dff_A_LcoIPl2v9_0),.din(w_dff_A_colYvOkg3_0),.clk(gclk));
	jdff dff_A_4LDx4qi96_0(.dout(w_dff_A_colYvOkg3_0),.din(w_dff_A_4LDx4qi96_0),.clk(gclk));
	jdff dff_B_XfxEq9Ce3_1(.din(n1839),.dout(w_dff_B_XfxEq9Ce3_1),.clk(gclk));
	jdff dff_B_yPOGelZU9_1(.din(w_dff_B_XfxEq9Ce3_1),.dout(w_dff_B_yPOGelZU9_1),.clk(gclk));
	jdff dff_B_e5lHSKNa5_2(.din(n1838),.dout(w_dff_B_e5lHSKNa5_2),.clk(gclk));
	jdff dff_B_SwwazD8w1_2(.din(w_dff_B_e5lHSKNa5_2),.dout(w_dff_B_SwwazD8w1_2),.clk(gclk));
	jdff dff_B_4uUjqRM31_2(.din(w_dff_B_SwwazD8w1_2),.dout(w_dff_B_4uUjqRM31_2),.clk(gclk));
	jdff dff_B_O3CQEj0Z1_2(.din(w_dff_B_4uUjqRM31_2),.dout(w_dff_B_O3CQEj0Z1_2),.clk(gclk));
	jdff dff_B_tauHEZS90_2(.din(w_dff_B_O3CQEj0Z1_2),.dout(w_dff_B_tauHEZS90_2),.clk(gclk));
	jdff dff_B_oQ8489kV3_2(.din(w_dff_B_tauHEZS90_2),.dout(w_dff_B_oQ8489kV3_2),.clk(gclk));
	jdff dff_B_WGJsjhGI8_2(.din(w_dff_B_oQ8489kV3_2),.dout(w_dff_B_WGJsjhGI8_2),.clk(gclk));
	jdff dff_B_xwv3mdxG7_2(.din(w_dff_B_WGJsjhGI8_2),.dout(w_dff_B_xwv3mdxG7_2),.clk(gclk));
	jdff dff_B_zvLRyb8F4_2(.din(w_dff_B_xwv3mdxG7_2),.dout(w_dff_B_zvLRyb8F4_2),.clk(gclk));
	jdff dff_B_GVFpIkiz6_2(.din(w_dff_B_zvLRyb8F4_2),.dout(w_dff_B_GVFpIkiz6_2),.clk(gclk));
	jdff dff_B_SzGCV5UT3_2(.din(w_dff_B_GVFpIkiz6_2),.dout(w_dff_B_SzGCV5UT3_2),.clk(gclk));
	jdff dff_B_tjPQLyOG7_2(.din(w_dff_B_SzGCV5UT3_2),.dout(w_dff_B_tjPQLyOG7_2),.clk(gclk));
	jdff dff_B_H8b1Kziu4_2(.din(w_dff_B_tjPQLyOG7_2),.dout(w_dff_B_H8b1Kziu4_2),.clk(gclk));
	jdff dff_B_3dsv6Bni5_2(.din(w_dff_B_H8b1Kziu4_2),.dout(w_dff_B_3dsv6Bni5_2),.clk(gclk));
	jdff dff_B_tYP9EpgD4_2(.din(w_dff_B_3dsv6Bni5_2),.dout(w_dff_B_tYP9EpgD4_2),.clk(gclk));
	jdff dff_B_Gv6Quh5z0_2(.din(w_dff_B_tYP9EpgD4_2),.dout(w_dff_B_Gv6Quh5z0_2),.clk(gclk));
	jdff dff_B_Qx8L1zGw4_2(.din(w_dff_B_Gv6Quh5z0_2),.dout(w_dff_B_Qx8L1zGw4_2),.clk(gclk));
	jdff dff_B_pW2EVA1U7_2(.din(w_dff_B_Qx8L1zGw4_2),.dout(w_dff_B_pW2EVA1U7_2),.clk(gclk));
	jdff dff_B_sFI1vrC85_2(.din(w_dff_B_pW2EVA1U7_2),.dout(w_dff_B_sFI1vrC85_2),.clk(gclk));
	jdff dff_B_9evJqlCy9_2(.din(w_dff_B_sFI1vrC85_2),.dout(w_dff_B_9evJqlCy9_2),.clk(gclk));
	jdff dff_B_F2CGKJ1r1_2(.din(w_dff_B_9evJqlCy9_2),.dout(w_dff_B_F2CGKJ1r1_2),.clk(gclk));
	jdff dff_B_IvaoF5hB3_2(.din(w_dff_B_F2CGKJ1r1_2),.dout(w_dff_B_IvaoF5hB3_2),.clk(gclk));
	jdff dff_B_n8LDiMXb8_2(.din(w_dff_B_IvaoF5hB3_2),.dout(w_dff_B_n8LDiMXb8_2),.clk(gclk));
	jdff dff_B_ACgpmFjb1_2(.din(w_dff_B_n8LDiMXb8_2),.dout(w_dff_B_ACgpmFjb1_2),.clk(gclk));
	jdff dff_B_4HxHcM400_2(.din(w_dff_B_ACgpmFjb1_2),.dout(w_dff_B_4HxHcM400_2),.clk(gclk));
	jdff dff_B_lbCrCuDa2_2(.din(w_dff_B_4HxHcM400_2),.dout(w_dff_B_lbCrCuDa2_2),.clk(gclk));
	jdff dff_B_vsPXZqz60_2(.din(w_dff_B_lbCrCuDa2_2),.dout(w_dff_B_vsPXZqz60_2),.clk(gclk));
	jdff dff_B_lgfc2Ygc6_2(.din(w_dff_B_vsPXZqz60_2),.dout(w_dff_B_lgfc2Ygc6_2),.clk(gclk));
	jdff dff_B_MG7DFbER2_2(.din(w_dff_B_lgfc2Ygc6_2),.dout(w_dff_B_MG7DFbER2_2),.clk(gclk));
	jdff dff_B_FXJeYFUg4_2(.din(w_dff_B_MG7DFbER2_2),.dout(w_dff_B_FXJeYFUg4_2),.clk(gclk));
	jdff dff_B_mN9IySnE2_2(.din(w_dff_B_FXJeYFUg4_2),.dout(w_dff_B_mN9IySnE2_2),.clk(gclk));
	jdff dff_B_ClKj2lYw6_2(.din(w_dff_B_mN9IySnE2_2),.dout(w_dff_B_ClKj2lYw6_2),.clk(gclk));
	jdff dff_B_9NuD0v7f8_2(.din(w_dff_B_ClKj2lYw6_2),.dout(w_dff_B_9NuD0v7f8_2),.clk(gclk));
	jdff dff_B_HXCVjWyU7_2(.din(w_dff_B_9NuD0v7f8_2),.dout(w_dff_B_HXCVjWyU7_2),.clk(gclk));
	jdff dff_B_pd3gmgXl8_2(.din(w_dff_B_HXCVjWyU7_2),.dout(w_dff_B_pd3gmgXl8_2),.clk(gclk));
	jdff dff_B_nDJ2Ak723_2(.din(w_dff_B_pd3gmgXl8_2),.dout(w_dff_B_nDJ2Ak723_2),.clk(gclk));
	jdff dff_B_QWTwQzaJ9_2(.din(w_dff_B_nDJ2Ak723_2),.dout(w_dff_B_QWTwQzaJ9_2),.clk(gclk));
	jdff dff_B_OkglBVIk2_2(.din(w_dff_B_QWTwQzaJ9_2),.dout(w_dff_B_OkglBVIk2_2),.clk(gclk));
	jdff dff_B_SkSwcdok2_2(.din(w_dff_B_OkglBVIk2_2),.dout(w_dff_B_SkSwcdok2_2),.clk(gclk));
	jdff dff_B_lEmrnIlw2_2(.din(w_dff_B_SkSwcdok2_2),.dout(w_dff_B_lEmrnIlw2_2),.clk(gclk));
	jdff dff_B_K98NEneF9_2(.din(w_dff_B_lEmrnIlw2_2),.dout(w_dff_B_K98NEneF9_2),.clk(gclk));
	jdff dff_B_Kau775vn0_2(.din(w_dff_B_K98NEneF9_2),.dout(w_dff_B_Kau775vn0_2),.clk(gclk));
	jdff dff_B_ufN8n1aH5_2(.din(w_dff_B_Kau775vn0_2),.dout(w_dff_B_ufN8n1aH5_2),.clk(gclk));
	jdff dff_B_QjNzuNJr6_2(.din(w_dff_B_ufN8n1aH5_2),.dout(w_dff_B_QjNzuNJr6_2),.clk(gclk));
	jdff dff_B_wf5pirFW9_2(.din(w_dff_B_QjNzuNJr6_2),.dout(w_dff_B_wf5pirFW9_2),.clk(gclk));
	jdff dff_B_no9VUopQ7_1(.din(n1845),.dout(w_dff_B_no9VUopQ7_1),.clk(gclk));
	jdff dff_B_nDhPnl7Z2_1(.din(w_dff_B_no9VUopQ7_1),.dout(w_dff_B_nDhPnl7Z2_1),.clk(gclk));
	jdff dff_B_9QfVd1cd8_1(.din(w_dff_B_nDhPnl7Z2_1),.dout(w_dff_B_9QfVd1cd8_1),.clk(gclk));
	jdff dff_B_o0VQrt6u1_0(.din(n1846),.dout(w_dff_B_o0VQrt6u1_0),.clk(gclk));
	jdff dff_B_bdjq8WZ84_0(.din(w_dff_B_o0VQrt6u1_0),.dout(w_dff_B_bdjq8WZ84_0),.clk(gclk));
	jdff dff_A_LHpOzrbB9_1(.dout(w_n1836_0[1]),.din(w_dff_A_LHpOzrbB9_1),.clk(gclk));
	jdff dff_A_0gs7R1tu9_1(.dout(w_dff_A_LHpOzrbB9_1),.din(w_dff_A_0gs7R1tu9_1),.clk(gclk));
	jdff dff_A_8XbjN7ht0_1(.dout(w_dff_A_0gs7R1tu9_1),.din(w_dff_A_8XbjN7ht0_1),.clk(gclk));
	jdff dff_B_KLybpQBG8_1(.din(n1821),.dout(w_dff_B_KLybpQBG8_1),.clk(gclk));
	jdff dff_B_RQidEsZv6_1(.din(w_dff_B_KLybpQBG8_1),.dout(w_dff_B_RQidEsZv6_1),.clk(gclk));
	jdff dff_B_J9BCiSGh4_1(.din(w_dff_B_RQidEsZv6_1),.dout(w_dff_B_J9BCiSGh4_1),.clk(gclk));
	jdff dff_B_kL81Hs7F0_0(.din(n1822),.dout(w_dff_B_kL81Hs7F0_0),.clk(gclk));
	jdff dff_B_q4rbk8rf0_0(.din(w_dff_B_kL81Hs7F0_0),.dout(w_dff_B_q4rbk8rf0_0),.clk(gclk));
	jdff dff_A_wwmBWZok5_1(.dout(w_n1817_0[1]),.din(w_dff_A_wwmBWZok5_1),.clk(gclk));
	jdff dff_A_IKXWMXrh0_1(.dout(w_dff_A_wwmBWZok5_1),.din(w_dff_A_IKXWMXrh0_1),.clk(gclk));
	jdff dff_A_xCr3eRnX3_1(.dout(w_dff_A_IKXWMXrh0_1),.din(w_dff_A_xCr3eRnX3_1),.clk(gclk));
	jdff dff_B_smNPmZ0o0_1(.din(n1795),.dout(w_dff_B_smNPmZ0o0_1),.clk(gclk));
	jdff dff_B_mGstzwpw6_1(.din(w_dff_B_smNPmZ0o0_1),.dout(w_dff_B_mGstzwpw6_1),.clk(gclk));
	jdff dff_B_OoUBXaLt3_1(.din(w_dff_B_mGstzwpw6_1),.dout(w_dff_B_OoUBXaLt3_1),.clk(gclk));
	jdff dff_B_PtIjhdST2_0(.din(n1796),.dout(w_dff_B_PtIjhdST2_0),.clk(gclk));
	jdff dff_B_L95tFTN21_0(.din(w_dff_B_PtIjhdST2_0),.dout(w_dff_B_L95tFTN21_0),.clk(gclk));
	jdff dff_A_KfbsAAkH5_1(.dout(w_n1791_0[1]),.din(w_dff_A_KfbsAAkH5_1),.clk(gclk));
	jdff dff_A_lGdhC9L15_1(.dout(w_dff_A_KfbsAAkH5_1),.din(w_dff_A_lGdhC9L15_1),.clk(gclk));
	jdff dff_A_RZILa9VN8_1(.dout(w_dff_A_lGdhC9L15_1),.din(w_dff_A_RZILa9VN8_1),.clk(gclk));
	jdff dff_B_R2kBV6Qy2_1(.din(n1762),.dout(w_dff_B_R2kBV6Qy2_1),.clk(gclk));
	jdff dff_B_RHSz7nkh9_1(.din(w_dff_B_R2kBV6Qy2_1),.dout(w_dff_B_RHSz7nkh9_1),.clk(gclk));
	jdff dff_B_qLp2GrJg0_1(.din(w_dff_B_RHSz7nkh9_1),.dout(w_dff_B_qLp2GrJg0_1),.clk(gclk));
	jdff dff_B_hI3AXSox5_0(.din(n1763),.dout(w_dff_B_hI3AXSox5_0),.clk(gclk));
	jdff dff_B_d0PaMaEw8_0(.din(w_dff_B_hI3AXSox5_0),.dout(w_dff_B_d0PaMaEw8_0),.clk(gclk));
	jdff dff_A_HYyviQ8l6_1(.dout(w_n1758_0[1]),.din(w_dff_A_HYyviQ8l6_1),.clk(gclk));
	jdff dff_A_OJKRTlii0_1(.dout(w_dff_A_HYyviQ8l6_1),.din(w_dff_A_OJKRTlii0_1),.clk(gclk));
	jdff dff_A_4zVLMqc52_1(.dout(w_dff_A_OJKRTlii0_1),.din(w_dff_A_4zVLMqc52_1),.clk(gclk));
	jdff dff_B_xmas2Tcw1_1(.din(n1722),.dout(w_dff_B_xmas2Tcw1_1),.clk(gclk));
	jdff dff_B_fMmwneKP0_1(.din(w_dff_B_xmas2Tcw1_1),.dout(w_dff_B_fMmwneKP0_1),.clk(gclk));
	jdff dff_B_FDF2le2Q4_1(.din(w_dff_B_fMmwneKP0_1),.dout(w_dff_B_FDF2le2Q4_1),.clk(gclk));
	jdff dff_B_wNIJnD189_0(.din(n1723),.dout(w_dff_B_wNIJnD189_0),.clk(gclk));
	jdff dff_A_dUeVK5hN0_1(.dout(w_n1720_0[1]),.din(w_dff_A_dUeVK5hN0_1),.clk(gclk));
	jdff dff_A_K74FCtSl7_1(.dout(w_dff_A_dUeVK5hN0_1),.din(w_dff_A_K74FCtSl7_1),.clk(gclk));
	jdff dff_B_dlR0tHnC9_1(.din(n1674),.dout(w_dff_B_dlR0tHnC9_1),.clk(gclk));
	jdff dff_B_4vwGwDhX0_1(.din(w_dff_B_dlR0tHnC9_1),.dout(w_dff_B_4vwGwDhX0_1),.clk(gclk));
	jdff dff_A_j7CybSZ25_1(.dout(w_n1672_0[1]),.din(w_dff_A_j7CybSZ25_1),.clk(gclk));
	jdff dff_B_JRhUGIwa0_1(.din(n1619),.dout(w_dff_B_JRhUGIwa0_1),.clk(gclk));
	jdff dff_B_FrfsuDlV9_1(.din(w_dff_B_JRhUGIwa0_1),.dout(w_dff_B_FrfsuDlV9_1),.clk(gclk));
	jdff dff_A_vLMIrqfW2_1(.dout(w_n1617_0[1]),.din(w_dff_A_vLMIrqfW2_1),.clk(gclk));
	jdff dff_B_cACy4Rp22_1(.din(n1557),.dout(w_dff_B_cACy4Rp22_1),.clk(gclk));
	jdff dff_B_mmxUZK7d1_1(.din(w_dff_B_cACy4Rp22_1),.dout(w_dff_B_mmxUZK7d1_1),.clk(gclk));
	jdff dff_A_GB6k6xy42_1(.dout(w_n1555_0[1]),.din(w_dff_A_GB6k6xy42_1),.clk(gclk));
	jdff dff_B_SMqQ1jin0_1(.din(n1488),.dout(w_dff_B_SMqQ1jin0_1),.clk(gclk));
	jdff dff_B_3ViiBqlr3_1(.din(w_dff_B_SMqQ1jin0_1),.dout(w_dff_B_3ViiBqlr3_1),.clk(gclk));
	jdff dff_A_uzm3y4NF2_1(.dout(w_n1486_0[1]),.din(w_dff_A_uzm3y4NF2_1),.clk(gclk));
	jdff dff_B_51WYu2pA6_1(.din(n1412),.dout(w_dff_B_51WYu2pA6_1),.clk(gclk));
	jdff dff_B_gezxGVAF9_1(.din(w_dff_B_51WYu2pA6_1),.dout(w_dff_B_gezxGVAF9_1),.clk(gclk));
	jdff dff_A_NXQdRrj24_0(.dout(w_n1332_0[0]),.din(w_dff_A_NXQdRrj24_0),.clk(gclk));
	jdff dff_B_aUjjF2ug5_1(.din(n1330),.dout(w_dff_B_aUjjF2ug5_1),.clk(gclk));
	jdff dff_A_3bZjpayx8_0(.dout(w_n1326_0[0]),.din(w_dff_A_3bZjpayx8_0),.clk(gclk));
	jdff dff_A_7yfYQd7z3_1(.dout(w_n1147_0[1]),.din(w_dff_A_7yfYQd7z3_1),.clk(gclk));
	jdff dff_B_7mxns7If6_2(.din(n1147),.dout(w_dff_B_7mxns7If6_2),.clk(gclk));
	jdff dff_A_QGWkux4p1_1(.dout(w_n1039_0[1]),.din(w_dff_A_QGWkux4p1_1),.clk(gclk));
	jdff dff_B_GAtqHJmd0_2(.din(n937),.dout(w_dff_B_GAtqHJmd0_2),.clk(gclk));
	jdff dff_B_BJ8Cjrj89_1(.din(n935),.dout(w_dff_B_BJ8Cjrj89_1),.clk(gclk));
	jdff dff_A_M2y5S9Ic2_0(.dout(w_n829_0[0]),.din(w_dff_A_M2y5S9Ic2_0),.clk(gclk));
	jdff dff_A_A2z74COT3_0(.dout(w_dff_A_M2y5S9Ic2_0),.din(w_dff_A_A2z74COT3_0),.clk(gclk));
	jdff dff_A_JIcAdYUM5_0(.dout(w_dff_A_A2z74COT3_0),.din(w_dff_A_JIcAdYUM5_0),.clk(gclk));
	jdff dff_A_JBsj4P8Y0_0(.dout(w_dff_A_JIcAdYUM5_0),.din(w_dff_A_JBsj4P8Y0_0),.clk(gclk));
	jdff dff_A_mRyn88YL5_0(.dout(w_dff_A_JBsj4P8Y0_0),.din(w_dff_A_mRyn88YL5_0),.clk(gclk));
	jdff dff_A_LMH93aDI4_0(.dout(w_dff_A_mRyn88YL5_0),.din(w_dff_A_LMH93aDI4_0),.clk(gclk));
	jdff dff_A_4dUtf8aZ0_0(.dout(w_dff_A_LMH93aDI4_0),.din(w_dff_A_4dUtf8aZ0_0),.clk(gclk));
	jdff dff_A_HRy1BVDF9_0(.dout(w_dff_A_4dUtf8aZ0_0),.din(w_dff_A_HRy1BVDF9_0),.clk(gclk));
	jdff dff_A_RA2lbvZJ3_0(.dout(w_dff_A_HRy1BVDF9_0),.din(w_dff_A_RA2lbvZJ3_0),.clk(gclk));
	jdff dff_A_OuYs5i7w5_0(.dout(w_dff_A_RA2lbvZJ3_0),.din(w_dff_A_OuYs5i7w5_0),.clk(gclk));
	jdff dff_A_nfBGby8k2_0(.dout(w_dff_A_OuYs5i7w5_0),.din(w_dff_A_nfBGby8k2_0),.clk(gclk));
	jdff dff_A_CAO2L0DN0_0(.dout(w_dff_A_nfBGby8k2_0),.din(w_dff_A_CAO2L0DN0_0),.clk(gclk));
	jdff dff_A_vVFD8ip00_0(.dout(w_dff_A_CAO2L0DN0_0),.din(w_dff_A_vVFD8ip00_0),.clk(gclk));
	jdff dff_A_IWHs54U20_0(.dout(w_dff_A_vVFD8ip00_0),.din(w_dff_A_IWHs54U20_0),.clk(gclk));
	jdff dff_A_stS7mkZF6_0(.dout(w_dff_A_IWHs54U20_0),.din(w_dff_A_stS7mkZF6_0),.clk(gclk));
	jdff dff_A_LcNbG2I07_0(.dout(w_dff_A_stS7mkZF6_0),.din(w_dff_A_LcNbG2I07_0),.clk(gclk));
	jdff dff_A_4X7SLdyk8_0(.dout(w_dff_A_LcNbG2I07_0),.din(w_dff_A_4X7SLdyk8_0),.clk(gclk));
	jdff dff_A_lA4eFy8G1_0(.dout(w_dff_A_4X7SLdyk8_0),.din(w_dff_A_lA4eFy8G1_0),.clk(gclk));
	jdff dff_A_Ni5oRJLR8_0(.dout(w_dff_A_lA4eFy8G1_0),.din(w_dff_A_Ni5oRJLR8_0),.clk(gclk));
	jdff dff_A_VzuHRQVR7_0(.dout(w_dff_A_Ni5oRJLR8_0),.din(w_dff_A_VzuHRQVR7_0),.clk(gclk));
	jdff dff_A_17Qpn3K31_0(.dout(w_dff_A_VzuHRQVR7_0),.din(w_dff_A_17Qpn3K31_0),.clk(gclk));
	jdff dff_A_oEJZhH0h4_0(.dout(w_dff_A_17Qpn3K31_0),.din(w_dff_A_oEJZhH0h4_0),.clk(gclk));
	jdff dff_A_NAMCyyWl9_0(.dout(w_dff_A_oEJZhH0h4_0),.din(w_dff_A_NAMCyyWl9_0),.clk(gclk));
	jdff dff_A_20oDcLU86_0(.dout(w_dff_A_NAMCyyWl9_0),.din(w_dff_A_20oDcLU86_0),.clk(gclk));
	jdff dff_A_b3mkxzp26_0(.dout(w_dff_A_20oDcLU86_0),.din(w_dff_A_b3mkxzp26_0),.clk(gclk));
	jdff dff_A_bp1CZuUc8_0(.dout(w_dff_A_b3mkxzp26_0),.din(w_dff_A_bp1CZuUc8_0),.clk(gclk));
	jdff dff_A_yLEvCfby4_0(.dout(w_dff_A_bp1CZuUc8_0),.din(w_dff_A_yLEvCfby4_0),.clk(gclk));
	jdff dff_A_FKnfKZf90_0(.dout(w_dff_A_yLEvCfby4_0),.din(w_dff_A_FKnfKZf90_0),.clk(gclk));
	jdff dff_A_CZmSBxDb7_0(.dout(w_dff_A_FKnfKZf90_0),.din(w_dff_A_CZmSBxDb7_0),.clk(gclk));
	jdff dff_A_TPvmPQxl1_0(.dout(w_dff_A_CZmSBxDb7_0),.din(w_dff_A_TPvmPQxl1_0),.clk(gclk));
	jdff dff_A_jiBmBqhU0_0(.dout(w_dff_A_TPvmPQxl1_0),.din(w_dff_A_jiBmBqhU0_0),.clk(gclk));
	jdff dff_A_IEtz1gEB5_0(.dout(w_dff_A_jiBmBqhU0_0),.din(w_dff_A_IEtz1gEB5_0),.clk(gclk));
	jdff dff_A_0sPTpbU60_1(.dout(w_n931_0[1]),.din(w_dff_A_0sPTpbU60_1),.clk(gclk));
	jdff dff_A_ckJvRe8q1_0(.dout(w_n729_0[0]),.din(w_dff_A_ckJvRe8q1_0),.clk(gclk));
	jdff dff_A_Ni3RkCnE9_0(.dout(w_dff_A_ckJvRe8q1_0),.din(w_dff_A_Ni3RkCnE9_0),.clk(gclk));
	jdff dff_A_4aLrPhyA2_0(.dout(w_dff_A_Ni3RkCnE9_0),.din(w_dff_A_4aLrPhyA2_0),.clk(gclk));
	jdff dff_A_TGoF8XTR4_0(.dout(w_dff_A_4aLrPhyA2_0),.din(w_dff_A_TGoF8XTR4_0),.clk(gclk));
	jdff dff_A_SptcI34m8_0(.dout(w_dff_A_TGoF8XTR4_0),.din(w_dff_A_SptcI34m8_0),.clk(gclk));
	jdff dff_A_JyliSIvt9_0(.dout(w_dff_A_SptcI34m8_0),.din(w_dff_A_JyliSIvt9_0),.clk(gclk));
	jdff dff_A_V9LDcEmT3_0(.dout(w_dff_A_JyliSIvt9_0),.din(w_dff_A_V9LDcEmT3_0),.clk(gclk));
	jdff dff_A_28GU9gwZ6_0(.dout(w_dff_A_V9LDcEmT3_0),.din(w_dff_A_28GU9gwZ6_0),.clk(gclk));
	jdff dff_A_526ddzCd9_0(.dout(w_dff_A_28GU9gwZ6_0),.din(w_dff_A_526ddzCd9_0),.clk(gclk));
	jdff dff_A_w5edsb1a8_0(.dout(w_dff_A_526ddzCd9_0),.din(w_dff_A_w5edsb1a8_0),.clk(gclk));
	jdff dff_A_YvzVBEEJ0_0(.dout(w_dff_A_w5edsb1a8_0),.din(w_dff_A_YvzVBEEJ0_0),.clk(gclk));
	jdff dff_A_C3bllVpi9_0(.dout(w_dff_A_YvzVBEEJ0_0),.din(w_dff_A_C3bllVpi9_0),.clk(gclk));
	jdff dff_A_MCFx6G085_0(.dout(w_dff_A_C3bllVpi9_0),.din(w_dff_A_MCFx6G085_0),.clk(gclk));
	jdff dff_A_2c3v1nxu0_0(.dout(w_dff_A_MCFx6G085_0),.din(w_dff_A_2c3v1nxu0_0),.clk(gclk));
	jdff dff_A_c6Mxnvs21_0(.dout(w_dff_A_2c3v1nxu0_0),.din(w_dff_A_c6Mxnvs21_0),.clk(gclk));
	jdff dff_A_crciOiXx2_0(.dout(w_dff_A_c6Mxnvs21_0),.din(w_dff_A_crciOiXx2_0),.clk(gclk));
	jdff dff_A_SVvyptEf1_0(.dout(w_dff_A_crciOiXx2_0),.din(w_dff_A_SVvyptEf1_0),.clk(gclk));
	jdff dff_A_nQ18yLAS9_0(.dout(w_dff_A_SVvyptEf1_0),.din(w_dff_A_nQ18yLAS9_0),.clk(gclk));
	jdff dff_A_fvr7R8Ou9_0(.dout(w_dff_A_nQ18yLAS9_0),.din(w_dff_A_fvr7R8Ou9_0),.clk(gclk));
	jdff dff_A_yM8oqcQK0_0(.dout(w_dff_A_fvr7R8Ou9_0),.din(w_dff_A_yM8oqcQK0_0),.clk(gclk));
	jdff dff_A_ePW2K3FK6_0(.dout(w_dff_A_yM8oqcQK0_0),.din(w_dff_A_ePW2K3FK6_0),.clk(gclk));
	jdff dff_A_48xqbwZu3_0(.dout(w_dff_A_ePW2K3FK6_0),.din(w_dff_A_48xqbwZu3_0),.clk(gclk));
	jdff dff_A_OxZ5SWrm2_0(.dout(w_dff_A_48xqbwZu3_0),.din(w_dff_A_OxZ5SWrm2_0),.clk(gclk));
	jdff dff_A_5tOxizFb2_0(.dout(w_dff_A_OxZ5SWrm2_0),.din(w_dff_A_5tOxizFb2_0),.clk(gclk));
	jdff dff_A_GZe99MoZ8_0(.dout(w_dff_A_5tOxizFb2_0),.din(w_dff_A_GZe99MoZ8_0),.clk(gclk));
	jdff dff_A_hwkeze6Q3_0(.dout(w_dff_A_GZe99MoZ8_0),.din(w_dff_A_hwkeze6Q3_0),.clk(gclk));
	jdff dff_A_byWbHRO86_0(.dout(w_dff_A_hwkeze6Q3_0),.din(w_dff_A_byWbHRO86_0),.clk(gclk));
	jdff dff_A_5eG2FIa74_0(.dout(w_dff_A_byWbHRO86_0),.din(w_dff_A_5eG2FIa74_0),.clk(gclk));
	jdff dff_A_HtM3viRm2_0(.dout(w_dff_A_5eG2FIa74_0),.din(w_dff_A_HtM3viRm2_0),.clk(gclk));
	jdff dff_A_1NxHfHhh4_0(.dout(w_dff_A_HtM3viRm2_0),.din(w_dff_A_1NxHfHhh4_0),.clk(gclk));
	jdff dff_B_j1Qyn4VR3_1(.din(n736),.dout(w_dff_B_j1Qyn4VR3_1),.clk(gclk));
	jdff dff_B_m8bmo6tf8_1(.din(w_dff_B_j1Qyn4VR3_1),.dout(w_dff_B_m8bmo6tf8_1),.clk(gclk));
	jdff dff_B_cW4qRpP29_1(.din(w_dff_B_m8bmo6tf8_1),.dout(w_dff_B_cW4qRpP29_1),.clk(gclk));
	jdff dff_B_hsCRbPDH6_1(.din(w_dff_B_cW4qRpP29_1),.dout(w_dff_B_hsCRbPDH6_1),.clk(gclk));
	jdff dff_B_n8oKYvc81_1(.din(w_dff_B_hsCRbPDH6_1),.dout(w_dff_B_n8oKYvc81_1),.clk(gclk));
	jdff dff_B_W0eCNOpV2_1(.din(w_dff_B_n8oKYvc81_1),.dout(w_dff_B_W0eCNOpV2_1),.clk(gclk));
	jdff dff_B_WwR90PSf0_1(.din(w_dff_B_W0eCNOpV2_1),.dout(w_dff_B_WwR90PSf0_1),.clk(gclk));
	jdff dff_B_4s2z4bQe9_1(.din(w_dff_B_WwR90PSf0_1),.dout(w_dff_B_4s2z4bQe9_1),.clk(gclk));
	jdff dff_B_Pc03QurW3_1(.din(w_dff_B_4s2z4bQe9_1),.dout(w_dff_B_Pc03QurW3_1),.clk(gclk));
	jdff dff_B_Q2hjMnad1_1(.din(w_dff_B_Pc03QurW3_1),.dout(w_dff_B_Q2hjMnad1_1),.clk(gclk));
	jdff dff_B_KW99sxBe3_1(.din(w_dff_B_Q2hjMnad1_1),.dout(w_dff_B_KW99sxBe3_1),.clk(gclk));
	jdff dff_B_KSsNT7ek7_1(.din(w_dff_B_KW99sxBe3_1),.dout(w_dff_B_KSsNT7ek7_1),.clk(gclk));
	jdff dff_B_i4zLOusD5_1(.din(w_dff_B_KSsNT7ek7_1),.dout(w_dff_B_i4zLOusD5_1),.clk(gclk));
	jdff dff_B_B7GCk5jB5_1(.din(w_dff_B_i4zLOusD5_1),.dout(w_dff_B_B7GCk5jB5_1),.clk(gclk));
	jdff dff_B_5XK3Jzp21_1(.din(w_dff_B_B7GCk5jB5_1),.dout(w_dff_B_5XK3Jzp21_1),.clk(gclk));
	jdff dff_B_hk2cQKiP0_1(.din(w_dff_B_5XK3Jzp21_1),.dout(w_dff_B_hk2cQKiP0_1),.clk(gclk));
	jdff dff_B_yoX6QolF8_1(.din(w_dff_B_hk2cQKiP0_1),.dout(w_dff_B_yoX6QolF8_1),.clk(gclk));
	jdff dff_B_gCb0fjIb4_1(.din(w_dff_B_yoX6QolF8_1),.dout(w_dff_B_gCb0fjIb4_1),.clk(gclk));
	jdff dff_B_9Qkc2j0j4_1(.din(w_dff_B_gCb0fjIb4_1),.dout(w_dff_B_9Qkc2j0j4_1),.clk(gclk));
	jdff dff_B_VAwY4NUY2_1(.din(w_dff_B_9Qkc2j0j4_1),.dout(w_dff_B_VAwY4NUY2_1),.clk(gclk));
	jdff dff_B_mxfUhMI60_1(.din(w_dff_B_VAwY4NUY2_1),.dout(w_dff_B_mxfUhMI60_1),.clk(gclk));
	jdff dff_B_jESRqfOh5_1(.din(w_dff_B_mxfUhMI60_1),.dout(w_dff_B_jESRqfOh5_1),.clk(gclk));
	jdff dff_B_bJiwrdoI9_1(.din(w_dff_B_jESRqfOh5_1),.dout(w_dff_B_bJiwrdoI9_1),.clk(gclk));
	jdff dff_B_5ogWIryP1_1(.din(w_dff_B_bJiwrdoI9_1),.dout(w_dff_B_5ogWIryP1_1),.clk(gclk));
	jdff dff_B_VyhpvSaU5_1(.din(w_dff_B_5ogWIryP1_1),.dout(w_dff_B_VyhpvSaU5_1),.clk(gclk));
	jdff dff_B_WoRw4qqH9_1(.din(w_dff_B_VyhpvSaU5_1),.dout(w_dff_B_WoRw4qqH9_1),.clk(gclk));
	jdff dff_B_xftUq9QE4_1(.din(w_dff_B_WoRw4qqH9_1),.dout(w_dff_B_xftUq9QE4_1),.clk(gclk));
	jdff dff_A_QRIEawwW9_0(.dout(w_n734_0[0]),.din(w_dff_A_QRIEawwW9_0),.clk(gclk));
	jdff dff_A_aRpb6lCj9_0(.dout(w_n636_0[0]),.din(w_dff_A_aRpb6lCj9_0),.clk(gclk));
	jdff dff_A_h3kN2Rjy9_0(.dout(w_dff_A_aRpb6lCj9_0),.din(w_dff_A_h3kN2Rjy9_0),.clk(gclk));
	jdff dff_A_aNVKrYK82_0(.dout(w_dff_A_h3kN2Rjy9_0),.din(w_dff_A_aNVKrYK82_0),.clk(gclk));
	jdff dff_A_SnlyMRNp5_0(.dout(w_dff_A_aNVKrYK82_0),.din(w_dff_A_SnlyMRNp5_0),.clk(gclk));
	jdff dff_A_tst7LY0G2_0(.dout(w_dff_A_SnlyMRNp5_0),.din(w_dff_A_tst7LY0G2_0),.clk(gclk));
	jdff dff_A_YoptpFe12_0(.dout(w_dff_A_tst7LY0G2_0),.din(w_dff_A_YoptpFe12_0),.clk(gclk));
	jdff dff_A_r7YpmhuF6_0(.dout(w_dff_A_YoptpFe12_0),.din(w_dff_A_r7YpmhuF6_0),.clk(gclk));
	jdff dff_A_6CCUXlFh6_0(.dout(w_dff_A_r7YpmhuF6_0),.din(w_dff_A_6CCUXlFh6_0),.clk(gclk));
	jdff dff_A_TdwC0G0v3_0(.dout(w_dff_A_6CCUXlFh6_0),.din(w_dff_A_TdwC0G0v3_0),.clk(gclk));
	jdff dff_A_sBPdLfx06_0(.dout(w_dff_A_TdwC0G0v3_0),.din(w_dff_A_sBPdLfx06_0),.clk(gclk));
	jdff dff_A_trkkQhNo2_0(.dout(w_dff_A_sBPdLfx06_0),.din(w_dff_A_trkkQhNo2_0),.clk(gclk));
	jdff dff_A_oqo6Js0f1_0(.dout(w_dff_A_trkkQhNo2_0),.din(w_dff_A_oqo6Js0f1_0),.clk(gclk));
	jdff dff_A_4FLuXmca2_0(.dout(w_dff_A_oqo6Js0f1_0),.din(w_dff_A_4FLuXmca2_0),.clk(gclk));
	jdff dff_A_f6sjOfPn2_0(.dout(w_dff_A_4FLuXmca2_0),.din(w_dff_A_f6sjOfPn2_0),.clk(gclk));
	jdff dff_A_DBZipzq48_0(.dout(w_dff_A_f6sjOfPn2_0),.din(w_dff_A_DBZipzq48_0),.clk(gclk));
	jdff dff_A_Nd5NTdfd6_0(.dout(w_dff_A_DBZipzq48_0),.din(w_dff_A_Nd5NTdfd6_0),.clk(gclk));
	jdff dff_A_hE6U68IY4_0(.dout(w_dff_A_Nd5NTdfd6_0),.din(w_dff_A_hE6U68IY4_0),.clk(gclk));
	jdff dff_A_0DmC97dg8_0(.dout(w_dff_A_hE6U68IY4_0),.din(w_dff_A_0DmC97dg8_0),.clk(gclk));
	jdff dff_A_2xMyIXmD9_0(.dout(w_dff_A_0DmC97dg8_0),.din(w_dff_A_2xMyIXmD9_0),.clk(gclk));
	jdff dff_A_L0ZJ7ZMt8_0(.dout(w_dff_A_2xMyIXmD9_0),.din(w_dff_A_L0ZJ7ZMt8_0),.clk(gclk));
	jdff dff_A_6eB7NOTM5_0(.dout(w_dff_A_L0ZJ7ZMt8_0),.din(w_dff_A_6eB7NOTM5_0),.clk(gclk));
	jdff dff_A_dYDNLr6f6_0(.dout(w_dff_A_6eB7NOTM5_0),.din(w_dff_A_dYDNLr6f6_0),.clk(gclk));
	jdff dff_A_37pS510B7_0(.dout(w_dff_A_dYDNLr6f6_0),.din(w_dff_A_37pS510B7_0),.clk(gclk));
	jdff dff_A_7h8LuNmB3_0(.dout(w_dff_A_37pS510B7_0),.din(w_dff_A_7h8LuNmB3_0),.clk(gclk));
	jdff dff_A_5ZDX1ojs8_0(.dout(w_dff_A_7h8LuNmB3_0),.din(w_dff_A_5ZDX1ojs8_0),.clk(gclk));
	jdff dff_A_t6ymttmX7_0(.dout(w_dff_A_5ZDX1ojs8_0),.din(w_dff_A_t6ymttmX7_0),.clk(gclk));
	jdff dff_A_mxYlMU4T7_0(.dout(w_dff_A_t6ymttmX7_0),.din(w_dff_A_mxYlMU4T7_0),.clk(gclk));
	jdff dff_A_5SfzQAxg5_0(.dout(w_dff_A_mxYlMU4T7_0),.din(w_dff_A_5SfzQAxg5_0),.clk(gclk));
	jdff dff_B_Gtx6iQUT5_1(.din(n643),.dout(w_dff_B_Gtx6iQUT5_1),.clk(gclk));
	jdff dff_B_wgVc6paT1_1(.din(w_dff_B_Gtx6iQUT5_1),.dout(w_dff_B_wgVc6paT1_1),.clk(gclk));
	jdff dff_B_dyBECQd94_1(.din(w_dff_B_wgVc6paT1_1),.dout(w_dff_B_dyBECQd94_1),.clk(gclk));
	jdff dff_B_y7YCC6nS9_1(.din(w_dff_B_dyBECQd94_1),.dout(w_dff_B_y7YCC6nS9_1),.clk(gclk));
	jdff dff_B_2rtJJHXR5_1(.din(w_dff_B_y7YCC6nS9_1),.dout(w_dff_B_2rtJJHXR5_1),.clk(gclk));
	jdff dff_B_dTfkslxc8_1(.din(w_dff_B_2rtJJHXR5_1),.dout(w_dff_B_dTfkslxc8_1),.clk(gclk));
	jdff dff_B_nRodWvVy6_1(.din(w_dff_B_dTfkslxc8_1),.dout(w_dff_B_nRodWvVy6_1),.clk(gclk));
	jdff dff_B_pfTDFgzc5_1(.din(w_dff_B_nRodWvVy6_1),.dout(w_dff_B_pfTDFgzc5_1),.clk(gclk));
	jdff dff_B_xJd63XPY8_1(.din(w_dff_B_pfTDFgzc5_1),.dout(w_dff_B_xJd63XPY8_1),.clk(gclk));
	jdff dff_B_VWS1LYYq2_1(.din(w_dff_B_xJd63XPY8_1),.dout(w_dff_B_VWS1LYYq2_1),.clk(gclk));
	jdff dff_B_Rhx6ugLh3_1(.din(w_dff_B_VWS1LYYq2_1),.dout(w_dff_B_Rhx6ugLh3_1),.clk(gclk));
	jdff dff_B_5kB4Rtwn1_1(.din(w_dff_B_Rhx6ugLh3_1),.dout(w_dff_B_5kB4Rtwn1_1),.clk(gclk));
	jdff dff_B_vqu4icbf5_1(.din(w_dff_B_5kB4Rtwn1_1),.dout(w_dff_B_vqu4icbf5_1),.clk(gclk));
	jdff dff_B_1ftpvpHc5_1(.din(w_dff_B_vqu4icbf5_1),.dout(w_dff_B_1ftpvpHc5_1),.clk(gclk));
	jdff dff_B_Dpo3CHuE5_1(.din(w_dff_B_1ftpvpHc5_1),.dout(w_dff_B_Dpo3CHuE5_1),.clk(gclk));
	jdff dff_B_ntEUX0s01_1(.din(w_dff_B_Dpo3CHuE5_1),.dout(w_dff_B_ntEUX0s01_1),.clk(gclk));
	jdff dff_B_LEganfDA6_1(.din(w_dff_B_ntEUX0s01_1),.dout(w_dff_B_LEganfDA6_1),.clk(gclk));
	jdff dff_B_i5rTkOQc3_1(.din(w_dff_B_LEganfDA6_1),.dout(w_dff_B_i5rTkOQc3_1),.clk(gclk));
	jdff dff_B_1Bmrf8M43_1(.din(w_dff_B_i5rTkOQc3_1),.dout(w_dff_B_1Bmrf8M43_1),.clk(gclk));
	jdff dff_B_Hj3FjrsB0_1(.din(w_dff_B_1Bmrf8M43_1),.dout(w_dff_B_Hj3FjrsB0_1),.clk(gclk));
	jdff dff_B_4Q5j9i1D5_1(.din(w_dff_B_Hj3FjrsB0_1),.dout(w_dff_B_4Q5j9i1D5_1),.clk(gclk));
	jdff dff_B_COvC5jYA1_1(.din(w_dff_B_4Q5j9i1D5_1),.dout(w_dff_B_COvC5jYA1_1),.clk(gclk));
	jdff dff_B_SN9eq7xb6_1(.din(w_dff_B_COvC5jYA1_1),.dout(w_dff_B_SN9eq7xb6_1),.clk(gclk));
	jdff dff_B_yCYtyNGu2_1(.din(w_dff_B_SN9eq7xb6_1),.dout(w_dff_B_yCYtyNGu2_1),.clk(gclk));
	jdff dff_B_Y7kUWzNe8_1(.din(w_dff_B_yCYtyNGu2_1),.dout(w_dff_B_Y7kUWzNe8_1),.clk(gclk));
	jdff dff_A_chNdRabH2_0(.dout(w_n641_0[0]),.din(w_dff_A_chNdRabH2_0),.clk(gclk));
	jdff dff_A_t6UoPEjo7_0(.dout(w_n550_0[0]),.din(w_dff_A_t6UoPEjo7_0),.clk(gclk));
	jdff dff_A_Xy5grSm04_0(.dout(w_dff_A_t6UoPEjo7_0),.din(w_dff_A_Xy5grSm04_0),.clk(gclk));
	jdff dff_A_pBCy3b054_0(.dout(w_dff_A_Xy5grSm04_0),.din(w_dff_A_pBCy3b054_0),.clk(gclk));
	jdff dff_A_2hueUNo63_0(.dout(w_dff_A_pBCy3b054_0),.din(w_dff_A_2hueUNo63_0),.clk(gclk));
	jdff dff_A_8YjE5BJm3_0(.dout(w_dff_A_2hueUNo63_0),.din(w_dff_A_8YjE5BJm3_0),.clk(gclk));
	jdff dff_A_gv21w5aP5_0(.dout(w_dff_A_8YjE5BJm3_0),.din(w_dff_A_gv21w5aP5_0),.clk(gclk));
	jdff dff_A_kVJo1b3u0_0(.dout(w_dff_A_gv21w5aP5_0),.din(w_dff_A_kVJo1b3u0_0),.clk(gclk));
	jdff dff_A_Olfva5oa8_0(.dout(w_dff_A_kVJo1b3u0_0),.din(w_dff_A_Olfva5oa8_0),.clk(gclk));
	jdff dff_A_YRCqZGhF9_0(.dout(w_dff_A_Olfva5oa8_0),.din(w_dff_A_YRCqZGhF9_0),.clk(gclk));
	jdff dff_A_USs8jSmu6_0(.dout(w_dff_A_YRCqZGhF9_0),.din(w_dff_A_USs8jSmu6_0),.clk(gclk));
	jdff dff_A_IuOQWvfL6_0(.dout(w_dff_A_USs8jSmu6_0),.din(w_dff_A_IuOQWvfL6_0),.clk(gclk));
	jdff dff_A_hsl7nrrv4_0(.dout(w_dff_A_IuOQWvfL6_0),.din(w_dff_A_hsl7nrrv4_0),.clk(gclk));
	jdff dff_A_BjYwVVvi0_0(.dout(w_dff_A_hsl7nrrv4_0),.din(w_dff_A_BjYwVVvi0_0),.clk(gclk));
	jdff dff_A_Swnzi0bJ0_0(.dout(w_dff_A_BjYwVVvi0_0),.din(w_dff_A_Swnzi0bJ0_0),.clk(gclk));
	jdff dff_A_KXe3CEHZ1_0(.dout(w_dff_A_Swnzi0bJ0_0),.din(w_dff_A_KXe3CEHZ1_0),.clk(gclk));
	jdff dff_A_2BXQFruY2_0(.dout(w_dff_A_KXe3CEHZ1_0),.din(w_dff_A_2BXQFruY2_0),.clk(gclk));
	jdff dff_A_DwUuqx5f6_0(.dout(w_dff_A_2BXQFruY2_0),.din(w_dff_A_DwUuqx5f6_0),.clk(gclk));
	jdff dff_A_7eF34zr54_0(.dout(w_dff_A_DwUuqx5f6_0),.din(w_dff_A_7eF34zr54_0),.clk(gclk));
	jdff dff_A_GdEAqnOh5_0(.dout(w_dff_A_7eF34zr54_0),.din(w_dff_A_GdEAqnOh5_0),.clk(gclk));
	jdff dff_A_LrlmMQgS7_0(.dout(w_dff_A_GdEAqnOh5_0),.din(w_dff_A_LrlmMQgS7_0),.clk(gclk));
	jdff dff_A_uvg8JFR27_0(.dout(w_dff_A_LrlmMQgS7_0),.din(w_dff_A_uvg8JFR27_0),.clk(gclk));
	jdff dff_A_XrxlCHqV1_0(.dout(w_dff_A_uvg8JFR27_0),.din(w_dff_A_XrxlCHqV1_0),.clk(gclk));
	jdff dff_A_lpGWMR4J8_0(.dout(w_dff_A_XrxlCHqV1_0),.din(w_dff_A_lpGWMR4J8_0),.clk(gclk));
	jdff dff_A_gx8XY1136_0(.dout(w_dff_A_lpGWMR4J8_0),.din(w_dff_A_gx8XY1136_0),.clk(gclk));
	jdff dff_A_DDChMjQ80_0(.dout(w_dff_A_gx8XY1136_0),.din(w_dff_A_DDChMjQ80_0),.clk(gclk));
	jdff dff_A_kbhaqNm07_0(.dout(w_dff_A_DDChMjQ80_0),.din(w_dff_A_kbhaqNm07_0),.clk(gclk));
	jdff dff_B_0Fl91qHa7_1(.din(n557),.dout(w_dff_B_0Fl91qHa7_1),.clk(gclk));
	jdff dff_B_oQaJROwe8_1(.din(w_dff_B_0Fl91qHa7_1),.dout(w_dff_B_oQaJROwe8_1),.clk(gclk));
	jdff dff_B_SIDBVwWf5_1(.din(w_dff_B_oQaJROwe8_1),.dout(w_dff_B_SIDBVwWf5_1),.clk(gclk));
	jdff dff_B_B9lmbFg19_1(.din(w_dff_B_SIDBVwWf5_1),.dout(w_dff_B_B9lmbFg19_1),.clk(gclk));
	jdff dff_B_rMR5z9EP1_1(.din(w_dff_B_B9lmbFg19_1),.dout(w_dff_B_rMR5z9EP1_1),.clk(gclk));
	jdff dff_B_36UGUMST0_1(.din(w_dff_B_rMR5z9EP1_1),.dout(w_dff_B_36UGUMST0_1),.clk(gclk));
	jdff dff_B_he42QObT1_1(.din(w_dff_B_36UGUMST0_1),.dout(w_dff_B_he42QObT1_1),.clk(gclk));
	jdff dff_B_OgHDIqo14_1(.din(w_dff_B_he42QObT1_1),.dout(w_dff_B_OgHDIqo14_1),.clk(gclk));
	jdff dff_B_zxabgURl9_1(.din(w_dff_B_OgHDIqo14_1),.dout(w_dff_B_zxabgURl9_1),.clk(gclk));
	jdff dff_B_QSwSKHzD6_1(.din(w_dff_B_zxabgURl9_1),.dout(w_dff_B_QSwSKHzD6_1),.clk(gclk));
	jdff dff_B_TWyROOLA9_1(.din(w_dff_B_QSwSKHzD6_1),.dout(w_dff_B_TWyROOLA9_1),.clk(gclk));
	jdff dff_B_iNmXmHwP8_1(.din(w_dff_B_TWyROOLA9_1),.dout(w_dff_B_iNmXmHwP8_1),.clk(gclk));
	jdff dff_B_WvdwlZDU6_1(.din(w_dff_B_iNmXmHwP8_1),.dout(w_dff_B_WvdwlZDU6_1),.clk(gclk));
	jdff dff_B_r9EjzCyz0_1(.din(w_dff_B_WvdwlZDU6_1),.dout(w_dff_B_r9EjzCyz0_1),.clk(gclk));
	jdff dff_B_5UpzrQaH9_1(.din(w_dff_B_r9EjzCyz0_1),.dout(w_dff_B_5UpzrQaH9_1),.clk(gclk));
	jdff dff_B_F5M7TLqH5_1(.din(w_dff_B_5UpzrQaH9_1),.dout(w_dff_B_F5M7TLqH5_1),.clk(gclk));
	jdff dff_B_AzM9MPQw4_1(.din(w_dff_B_F5M7TLqH5_1),.dout(w_dff_B_AzM9MPQw4_1),.clk(gclk));
	jdff dff_B_XQJnSe9C6_1(.din(w_dff_B_AzM9MPQw4_1),.dout(w_dff_B_XQJnSe9C6_1),.clk(gclk));
	jdff dff_B_2D7TI53e2_1(.din(w_dff_B_XQJnSe9C6_1),.dout(w_dff_B_2D7TI53e2_1),.clk(gclk));
	jdff dff_B_DiYja20U1_1(.din(w_dff_B_2D7TI53e2_1),.dout(w_dff_B_DiYja20U1_1),.clk(gclk));
	jdff dff_B_nsyH24CG9_1(.din(w_dff_B_DiYja20U1_1),.dout(w_dff_B_nsyH24CG9_1),.clk(gclk));
	jdff dff_B_u03696M12_1(.din(w_dff_B_nsyH24CG9_1),.dout(w_dff_B_u03696M12_1),.clk(gclk));
	jdff dff_B_Bid8kzJ10_1(.din(w_dff_B_u03696M12_1),.dout(w_dff_B_Bid8kzJ10_1),.clk(gclk));
	jdff dff_A_al1351FM3_0(.dout(w_n555_0[0]),.din(w_dff_A_al1351FM3_0),.clk(gclk));
	jdff dff_A_JaPsF6wM6_0(.dout(w_n471_0[0]),.din(w_dff_A_JaPsF6wM6_0),.clk(gclk));
	jdff dff_A_7lPUfc5j1_0(.dout(w_dff_A_JaPsF6wM6_0),.din(w_dff_A_7lPUfc5j1_0),.clk(gclk));
	jdff dff_A_GfbLkeaF8_0(.dout(w_dff_A_7lPUfc5j1_0),.din(w_dff_A_GfbLkeaF8_0),.clk(gclk));
	jdff dff_A_IARJly4G8_0(.dout(w_dff_A_GfbLkeaF8_0),.din(w_dff_A_IARJly4G8_0),.clk(gclk));
	jdff dff_A_S3vFVcLD6_0(.dout(w_dff_A_IARJly4G8_0),.din(w_dff_A_S3vFVcLD6_0),.clk(gclk));
	jdff dff_A_H2H2BRE85_0(.dout(w_dff_A_S3vFVcLD6_0),.din(w_dff_A_H2H2BRE85_0),.clk(gclk));
	jdff dff_A_ADcGAanS1_0(.dout(w_dff_A_H2H2BRE85_0),.din(w_dff_A_ADcGAanS1_0),.clk(gclk));
	jdff dff_A_jQKr9a962_0(.dout(w_dff_A_ADcGAanS1_0),.din(w_dff_A_jQKr9a962_0),.clk(gclk));
	jdff dff_A_jfStBTsP3_0(.dout(w_dff_A_jQKr9a962_0),.din(w_dff_A_jfStBTsP3_0),.clk(gclk));
	jdff dff_A_P0llhrgA8_0(.dout(w_dff_A_jfStBTsP3_0),.din(w_dff_A_P0llhrgA8_0),.clk(gclk));
	jdff dff_A_QcoF8xF19_0(.dout(w_dff_A_P0llhrgA8_0),.din(w_dff_A_QcoF8xF19_0),.clk(gclk));
	jdff dff_A_xM9sCwMX4_0(.dout(w_dff_A_QcoF8xF19_0),.din(w_dff_A_xM9sCwMX4_0),.clk(gclk));
	jdff dff_A_ifSAndGT2_0(.dout(w_dff_A_xM9sCwMX4_0),.din(w_dff_A_ifSAndGT2_0),.clk(gclk));
	jdff dff_A_Z40eYaM17_0(.dout(w_dff_A_ifSAndGT2_0),.din(w_dff_A_Z40eYaM17_0),.clk(gclk));
	jdff dff_A_Oafz2oKT9_0(.dout(w_dff_A_Z40eYaM17_0),.din(w_dff_A_Oafz2oKT9_0),.clk(gclk));
	jdff dff_A_CjbwsbKT4_0(.dout(w_dff_A_Oafz2oKT9_0),.din(w_dff_A_CjbwsbKT4_0),.clk(gclk));
	jdff dff_A_ysOHlpa41_0(.dout(w_dff_A_CjbwsbKT4_0),.din(w_dff_A_ysOHlpa41_0),.clk(gclk));
	jdff dff_A_aqIJ95c39_0(.dout(w_dff_A_ysOHlpa41_0),.din(w_dff_A_aqIJ95c39_0),.clk(gclk));
	jdff dff_A_33K2h22O9_0(.dout(w_dff_A_aqIJ95c39_0),.din(w_dff_A_33K2h22O9_0),.clk(gclk));
	jdff dff_A_mN8EVr0i4_0(.dout(w_dff_A_33K2h22O9_0),.din(w_dff_A_mN8EVr0i4_0),.clk(gclk));
	jdff dff_A_AR0uX3qQ2_0(.dout(w_dff_A_mN8EVr0i4_0),.din(w_dff_A_AR0uX3qQ2_0),.clk(gclk));
	jdff dff_A_CxgODUZJ1_0(.dout(w_dff_A_AR0uX3qQ2_0),.din(w_dff_A_CxgODUZJ1_0),.clk(gclk));
	jdff dff_A_gpPMgTpp3_0(.dout(w_dff_A_CxgODUZJ1_0),.din(w_dff_A_gpPMgTpp3_0),.clk(gclk));
	jdff dff_A_vEIwA6aA0_0(.dout(w_dff_A_gpPMgTpp3_0),.din(w_dff_A_vEIwA6aA0_0),.clk(gclk));
	jdff dff_B_ud8QjlEU3_1(.din(n478),.dout(w_dff_B_ud8QjlEU3_1),.clk(gclk));
	jdff dff_B_zmI335mi6_1(.din(w_dff_B_ud8QjlEU3_1),.dout(w_dff_B_zmI335mi6_1),.clk(gclk));
	jdff dff_B_bWBOJdYY1_1(.din(w_dff_B_zmI335mi6_1),.dout(w_dff_B_bWBOJdYY1_1),.clk(gclk));
	jdff dff_B_xr8SIehP1_1(.din(w_dff_B_bWBOJdYY1_1),.dout(w_dff_B_xr8SIehP1_1),.clk(gclk));
	jdff dff_B_XLedBFm88_1(.din(w_dff_B_xr8SIehP1_1),.dout(w_dff_B_XLedBFm88_1),.clk(gclk));
	jdff dff_B_doerRJqm9_1(.din(w_dff_B_XLedBFm88_1),.dout(w_dff_B_doerRJqm9_1),.clk(gclk));
	jdff dff_B_rLxTfpQs0_1(.din(w_dff_B_doerRJqm9_1),.dout(w_dff_B_rLxTfpQs0_1),.clk(gclk));
	jdff dff_B_pSRY3bP35_1(.din(w_dff_B_rLxTfpQs0_1),.dout(w_dff_B_pSRY3bP35_1),.clk(gclk));
	jdff dff_B_eAhSCHeG3_1(.din(w_dff_B_pSRY3bP35_1),.dout(w_dff_B_eAhSCHeG3_1),.clk(gclk));
	jdff dff_B_PQF5T7Wg5_1(.din(w_dff_B_eAhSCHeG3_1),.dout(w_dff_B_PQF5T7Wg5_1),.clk(gclk));
	jdff dff_B_MtaOSoxO6_1(.din(w_dff_B_PQF5T7Wg5_1),.dout(w_dff_B_MtaOSoxO6_1),.clk(gclk));
	jdff dff_B_WsdHjk4y5_1(.din(w_dff_B_MtaOSoxO6_1),.dout(w_dff_B_WsdHjk4y5_1),.clk(gclk));
	jdff dff_B_xOW5Oup12_1(.din(w_dff_B_WsdHjk4y5_1),.dout(w_dff_B_xOW5Oup12_1),.clk(gclk));
	jdff dff_B_3l0KOHsB0_1(.din(w_dff_B_xOW5Oup12_1),.dout(w_dff_B_3l0KOHsB0_1),.clk(gclk));
	jdff dff_B_56TIV0FV7_1(.din(w_dff_B_3l0KOHsB0_1),.dout(w_dff_B_56TIV0FV7_1),.clk(gclk));
	jdff dff_B_R7nHuzbv0_1(.din(w_dff_B_56TIV0FV7_1),.dout(w_dff_B_R7nHuzbv0_1),.clk(gclk));
	jdff dff_B_uNLZFaGt3_1(.din(w_dff_B_R7nHuzbv0_1),.dout(w_dff_B_uNLZFaGt3_1),.clk(gclk));
	jdff dff_B_aRHot1te5_1(.din(w_dff_B_uNLZFaGt3_1),.dout(w_dff_B_aRHot1te5_1),.clk(gclk));
	jdff dff_B_WnJR3tlD2_1(.din(w_dff_B_aRHot1te5_1),.dout(w_dff_B_WnJR3tlD2_1),.clk(gclk));
	jdff dff_B_H9cIAPfO1_1(.din(w_dff_B_WnJR3tlD2_1),.dout(w_dff_B_H9cIAPfO1_1),.clk(gclk));
	jdff dff_B_vTo9DWpq2_1(.din(w_dff_B_H9cIAPfO1_1),.dout(w_dff_B_vTo9DWpq2_1),.clk(gclk));
	jdff dff_A_swXZQXih8_0(.dout(w_n476_0[0]),.din(w_dff_A_swXZQXih8_0),.clk(gclk));
	jdff dff_A_05DEkaV64_0(.dout(w_n399_0[0]),.din(w_dff_A_05DEkaV64_0),.clk(gclk));
	jdff dff_A_oS9J8bpO0_0(.dout(w_dff_A_05DEkaV64_0),.din(w_dff_A_oS9J8bpO0_0),.clk(gclk));
	jdff dff_A_wrzDHA7Z5_0(.dout(w_dff_A_oS9J8bpO0_0),.din(w_dff_A_wrzDHA7Z5_0),.clk(gclk));
	jdff dff_A_j3vvAh7y7_0(.dout(w_dff_A_wrzDHA7Z5_0),.din(w_dff_A_j3vvAh7y7_0),.clk(gclk));
	jdff dff_A_ojWLVKT07_0(.dout(w_dff_A_j3vvAh7y7_0),.din(w_dff_A_ojWLVKT07_0),.clk(gclk));
	jdff dff_A_hw03vZm11_0(.dout(w_dff_A_ojWLVKT07_0),.din(w_dff_A_hw03vZm11_0),.clk(gclk));
	jdff dff_A_yvzcvKpM1_0(.dout(w_dff_A_hw03vZm11_0),.din(w_dff_A_yvzcvKpM1_0),.clk(gclk));
	jdff dff_A_teefEHzH5_0(.dout(w_dff_A_yvzcvKpM1_0),.din(w_dff_A_teefEHzH5_0),.clk(gclk));
	jdff dff_A_2KoD1YQX8_0(.dout(w_dff_A_teefEHzH5_0),.din(w_dff_A_2KoD1YQX8_0),.clk(gclk));
	jdff dff_A_KRqEwjQ81_0(.dout(w_dff_A_2KoD1YQX8_0),.din(w_dff_A_KRqEwjQ81_0),.clk(gclk));
	jdff dff_A_k0spBbv27_0(.dout(w_dff_A_KRqEwjQ81_0),.din(w_dff_A_k0spBbv27_0),.clk(gclk));
	jdff dff_A_1y2ZKeWk4_0(.dout(w_dff_A_k0spBbv27_0),.din(w_dff_A_1y2ZKeWk4_0),.clk(gclk));
	jdff dff_A_ACy3FlvS3_0(.dout(w_dff_A_1y2ZKeWk4_0),.din(w_dff_A_ACy3FlvS3_0),.clk(gclk));
	jdff dff_A_LZ60edm54_0(.dout(w_dff_A_ACy3FlvS3_0),.din(w_dff_A_LZ60edm54_0),.clk(gclk));
	jdff dff_A_W3yj2vlt8_0(.dout(w_dff_A_LZ60edm54_0),.din(w_dff_A_W3yj2vlt8_0),.clk(gclk));
	jdff dff_A_J1NUl2kS2_0(.dout(w_dff_A_W3yj2vlt8_0),.din(w_dff_A_J1NUl2kS2_0),.clk(gclk));
	jdff dff_A_dqFCisM34_0(.dout(w_dff_A_J1NUl2kS2_0),.din(w_dff_A_dqFCisM34_0),.clk(gclk));
	jdff dff_A_6u1ojk1k5_0(.dout(w_dff_A_dqFCisM34_0),.din(w_dff_A_6u1ojk1k5_0),.clk(gclk));
	jdff dff_A_U3qzrxTV4_0(.dout(w_dff_A_6u1ojk1k5_0),.din(w_dff_A_U3qzrxTV4_0),.clk(gclk));
	jdff dff_A_1xG9BDfg7_0(.dout(w_dff_A_U3qzrxTV4_0),.din(w_dff_A_1xG9BDfg7_0),.clk(gclk));
	jdff dff_A_q9OgaS2z8_0(.dout(w_dff_A_1xG9BDfg7_0),.din(w_dff_A_q9OgaS2z8_0),.clk(gclk));
	jdff dff_A_hM36iCne8_0(.dout(w_dff_A_q9OgaS2z8_0),.din(w_dff_A_hM36iCne8_0),.clk(gclk));
	jdff dff_B_uTZb6Z3s7_1(.din(n406),.dout(w_dff_B_uTZb6Z3s7_1),.clk(gclk));
	jdff dff_B_hm1fPZAq7_1(.din(w_dff_B_uTZb6Z3s7_1),.dout(w_dff_B_hm1fPZAq7_1),.clk(gclk));
	jdff dff_B_EHcLlbm60_1(.din(w_dff_B_hm1fPZAq7_1),.dout(w_dff_B_EHcLlbm60_1),.clk(gclk));
	jdff dff_B_ODuCTbQ85_1(.din(w_dff_B_EHcLlbm60_1),.dout(w_dff_B_ODuCTbQ85_1),.clk(gclk));
	jdff dff_B_izjg92Ap4_1(.din(w_dff_B_ODuCTbQ85_1),.dout(w_dff_B_izjg92Ap4_1),.clk(gclk));
	jdff dff_B_L8w81y2j8_1(.din(w_dff_B_izjg92Ap4_1),.dout(w_dff_B_L8w81y2j8_1),.clk(gclk));
	jdff dff_B_zWcbds0U5_1(.din(w_dff_B_L8w81y2j8_1),.dout(w_dff_B_zWcbds0U5_1),.clk(gclk));
	jdff dff_B_5XlOMBgl2_1(.din(w_dff_B_zWcbds0U5_1),.dout(w_dff_B_5XlOMBgl2_1),.clk(gclk));
	jdff dff_B_b5uxt2mY6_1(.din(w_dff_B_5XlOMBgl2_1),.dout(w_dff_B_b5uxt2mY6_1),.clk(gclk));
	jdff dff_B_VhGYBEJb5_1(.din(w_dff_B_b5uxt2mY6_1),.dout(w_dff_B_VhGYBEJb5_1),.clk(gclk));
	jdff dff_B_afhVULOk7_1(.din(w_dff_B_VhGYBEJb5_1),.dout(w_dff_B_afhVULOk7_1),.clk(gclk));
	jdff dff_B_NWYGAxDR3_1(.din(w_dff_B_afhVULOk7_1),.dout(w_dff_B_NWYGAxDR3_1),.clk(gclk));
	jdff dff_B_5bHmcDTs4_1(.din(w_dff_B_NWYGAxDR3_1),.dout(w_dff_B_5bHmcDTs4_1),.clk(gclk));
	jdff dff_B_RgpgXzOc0_1(.din(w_dff_B_5bHmcDTs4_1),.dout(w_dff_B_RgpgXzOc0_1),.clk(gclk));
	jdff dff_B_0SHDZ3w04_1(.din(w_dff_B_RgpgXzOc0_1),.dout(w_dff_B_0SHDZ3w04_1),.clk(gclk));
	jdff dff_B_16LtevOL6_1(.din(w_dff_B_0SHDZ3w04_1),.dout(w_dff_B_16LtevOL6_1),.clk(gclk));
	jdff dff_B_shtQC2Mn4_1(.din(w_dff_B_16LtevOL6_1),.dout(w_dff_B_shtQC2Mn4_1),.clk(gclk));
	jdff dff_B_YUNO8IgW0_1(.din(w_dff_B_shtQC2Mn4_1),.dout(w_dff_B_YUNO8IgW0_1),.clk(gclk));
	jdff dff_B_E5IsYMmE0_1(.din(w_dff_B_YUNO8IgW0_1),.dout(w_dff_B_E5IsYMmE0_1),.clk(gclk));
	jdff dff_A_TVX9hYFf4_0(.dout(w_n404_0[0]),.din(w_dff_A_TVX9hYFf4_0),.clk(gclk));
	jdff dff_A_tJT3KFuh6_0(.dout(w_n335_0[0]),.din(w_dff_A_tJT3KFuh6_0),.clk(gclk));
	jdff dff_A_W4EAAdrH1_0(.dout(w_dff_A_tJT3KFuh6_0),.din(w_dff_A_W4EAAdrH1_0),.clk(gclk));
	jdff dff_A_FqopWnku8_0(.dout(w_dff_A_W4EAAdrH1_0),.din(w_dff_A_FqopWnku8_0),.clk(gclk));
	jdff dff_A_bvsaJjqH8_0(.dout(w_dff_A_FqopWnku8_0),.din(w_dff_A_bvsaJjqH8_0),.clk(gclk));
	jdff dff_A_pOTCGV5m3_0(.dout(w_dff_A_bvsaJjqH8_0),.din(w_dff_A_pOTCGV5m3_0),.clk(gclk));
	jdff dff_A_aKvz969A3_0(.dout(w_dff_A_pOTCGV5m3_0),.din(w_dff_A_aKvz969A3_0),.clk(gclk));
	jdff dff_A_dYxmvQzE1_0(.dout(w_dff_A_aKvz969A3_0),.din(w_dff_A_dYxmvQzE1_0),.clk(gclk));
	jdff dff_A_py3Lhpao5_0(.dout(w_dff_A_dYxmvQzE1_0),.din(w_dff_A_py3Lhpao5_0),.clk(gclk));
	jdff dff_A_RPAy8iYG1_0(.dout(w_dff_A_py3Lhpao5_0),.din(w_dff_A_RPAy8iYG1_0),.clk(gclk));
	jdff dff_A_MlQGDNEl0_0(.dout(w_dff_A_RPAy8iYG1_0),.din(w_dff_A_MlQGDNEl0_0),.clk(gclk));
	jdff dff_A_8VIXhoDg6_0(.dout(w_dff_A_MlQGDNEl0_0),.din(w_dff_A_8VIXhoDg6_0),.clk(gclk));
	jdff dff_A_tTJxgcJW1_0(.dout(w_dff_A_8VIXhoDg6_0),.din(w_dff_A_tTJxgcJW1_0),.clk(gclk));
	jdff dff_A_HQMVwezQ1_0(.dout(w_dff_A_tTJxgcJW1_0),.din(w_dff_A_HQMVwezQ1_0),.clk(gclk));
	jdff dff_A_HSaA9MkR6_0(.dout(w_dff_A_HQMVwezQ1_0),.din(w_dff_A_HSaA9MkR6_0),.clk(gclk));
	jdff dff_A_iMhyR4d71_0(.dout(w_dff_A_HSaA9MkR6_0),.din(w_dff_A_iMhyR4d71_0),.clk(gclk));
	jdff dff_A_QBgFagCF7_0(.dout(w_dff_A_iMhyR4d71_0),.din(w_dff_A_QBgFagCF7_0),.clk(gclk));
	jdff dff_A_6cadBoT13_0(.dout(w_dff_A_QBgFagCF7_0),.din(w_dff_A_6cadBoT13_0),.clk(gclk));
	jdff dff_A_vYF5bntp6_0(.dout(w_dff_A_6cadBoT13_0),.din(w_dff_A_vYF5bntp6_0),.clk(gclk));
	jdff dff_A_sOfPWkRK0_0(.dout(w_dff_A_vYF5bntp6_0),.din(w_dff_A_sOfPWkRK0_0),.clk(gclk));
	jdff dff_A_Vez93m5r5_0(.dout(w_dff_A_sOfPWkRK0_0),.din(w_dff_A_Vez93m5r5_0),.clk(gclk));
	jdff dff_B_m1nTTzLv5_1(.din(n342),.dout(w_dff_B_m1nTTzLv5_1),.clk(gclk));
	jdff dff_B_LcYa4VeC7_1(.din(w_dff_B_m1nTTzLv5_1),.dout(w_dff_B_LcYa4VeC7_1),.clk(gclk));
	jdff dff_B_08TmuP7q1_1(.din(w_dff_B_LcYa4VeC7_1),.dout(w_dff_B_08TmuP7q1_1),.clk(gclk));
	jdff dff_B_2mJ8EhpL4_1(.din(w_dff_B_08TmuP7q1_1),.dout(w_dff_B_2mJ8EhpL4_1),.clk(gclk));
	jdff dff_B_3FLLYQeS5_1(.din(w_dff_B_2mJ8EhpL4_1),.dout(w_dff_B_3FLLYQeS5_1),.clk(gclk));
	jdff dff_B_cA2vQFFR6_1(.din(w_dff_B_3FLLYQeS5_1),.dout(w_dff_B_cA2vQFFR6_1),.clk(gclk));
	jdff dff_B_YgSRbCQH3_1(.din(w_dff_B_cA2vQFFR6_1),.dout(w_dff_B_YgSRbCQH3_1),.clk(gclk));
	jdff dff_B_GlLYAf4y4_1(.din(w_dff_B_YgSRbCQH3_1),.dout(w_dff_B_GlLYAf4y4_1),.clk(gclk));
	jdff dff_B_nE6JvbLd3_1(.din(w_dff_B_GlLYAf4y4_1),.dout(w_dff_B_nE6JvbLd3_1),.clk(gclk));
	jdff dff_B_SP1WKq941_1(.din(w_dff_B_nE6JvbLd3_1),.dout(w_dff_B_SP1WKq941_1),.clk(gclk));
	jdff dff_B_etxLYvyE0_1(.din(w_dff_B_SP1WKq941_1),.dout(w_dff_B_etxLYvyE0_1),.clk(gclk));
	jdff dff_B_y1UcUOWs1_1(.din(w_dff_B_etxLYvyE0_1),.dout(w_dff_B_y1UcUOWs1_1),.clk(gclk));
	jdff dff_B_F0WfyupO0_1(.din(w_dff_B_y1UcUOWs1_1),.dout(w_dff_B_F0WfyupO0_1),.clk(gclk));
	jdff dff_B_DNlOVOYA8_1(.din(w_dff_B_F0WfyupO0_1),.dout(w_dff_B_DNlOVOYA8_1),.clk(gclk));
	jdff dff_B_U4FZBcFX0_1(.din(w_dff_B_DNlOVOYA8_1),.dout(w_dff_B_U4FZBcFX0_1),.clk(gclk));
	jdff dff_B_Gu4FAlXo2_1(.din(w_dff_B_U4FZBcFX0_1),.dout(w_dff_B_Gu4FAlXo2_1),.clk(gclk));
	jdff dff_B_uzgOcgVR6_1(.din(w_dff_B_Gu4FAlXo2_1),.dout(w_dff_B_uzgOcgVR6_1),.clk(gclk));
	jdff dff_A_2T7pXLSx7_0(.dout(w_n340_0[0]),.din(w_dff_A_2T7pXLSx7_0),.clk(gclk));
	jdff dff_A_Pix4WXTg3_0(.dout(w_n277_0[0]),.din(w_dff_A_Pix4WXTg3_0),.clk(gclk));
	jdff dff_A_LPLBZKPO0_0(.dout(w_dff_A_Pix4WXTg3_0),.din(w_dff_A_LPLBZKPO0_0),.clk(gclk));
	jdff dff_A_8egFxdP22_0(.dout(w_dff_A_LPLBZKPO0_0),.din(w_dff_A_8egFxdP22_0),.clk(gclk));
	jdff dff_A_khLpirm57_0(.dout(w_dff_A_8egFxdP22_0),.din(w_dff_A_khLpirm57_0),.clk(gclk));
	jdff dff_A_0GYK5jNy7_0(.dout(w_dff_A_khLpirm57_0),.din(w_dff_A_0GYK5jNy7_0),.clk(gclk));
	jdff dff_A_x0qTc6vE7_0(.dout(w_dff_A_0GYK5jNy7_0),.din(w_dff_A_x0qTc6vE7_0),.clk(gclk));
	jdff dff_A_DpsND7iO2_0(.dout(w_dff_A_x0qTc6vE7_0),.din(w_dff_A_DpsND7iO2_0),.clk(gclk));
	jdff dff_A_9S7CCJsF3_0(.dout(w_dff_A_DpsND7iO2_0),.din(w_dff_A_9S7CCJsF3_0),.clk(gclk));
	jdff dff_A_Pz0QLjXJ3_0(.dout(w_dff_A_9S7CCJsF3_0),.din(w_dff_A_Pz0QLjXJ3_0),.clk(gclk));
	jdff dff_A_nYuhlZqn1_0(.dout(w_dff_A_Pz0QLjXJ3_0),.din(w_dff_A_nYuhlZqn1_0),.clk(gclk));
	jdff dff_A_2EpMaSnq8_0(.dout(w_dff_A_nYuhlZqn1_0),.din(w_dff_A_2EpMaSnq8_0),.clk(gclk));
	jdff dff_A_673CrR0C2_0(.dout(w_dff_A_2EpMaSnq8_0),.din(w_dff_A_673CrR0C2_0),.clk(gclk));
	jdff dff_A_WSzD5Wpn9_0(.dout(w_dff_A_673CrR0C2_0),.din(w_dff_A_WSzD5Wpn9_0),.clk(gclk));
	jdff dff_A_lNBjx5ke5_0(.dout(w_dff_A_WSzD5Wpn9_0),.din(w_dff_A_lNBjx5ke5_0),.clk(gclk));
	jdff dff_A_CvXFFNkg9_0(.dout(w_dff_A_lNBjx5ke5_0),.din(w_dff_A_CvXFFNkg9_0),.clk(gclk));
	jdff dff_A_FdzGiTDI8_0(.dout(w_dff_A_CvXFFNkg9_0),.din(w_dff_A_FdzGiTDI8_0),.clk(gclk));
	jdff dff_A_IoO125sj7_0(.dout(w_dff_A_FdzGiTDI8_0),.din(w_dff_A_IoO125sj7_0),.clk(gclk));
	jdff dff_A_m3nABioh9_0(.dout(w_dff_A_IoO125sj7_0),.din(w_dff_A_m3nABioh9_0),.clk(gclk));
	jdff dff_B_bXzx77a41_1(.din(n284),.dout(w_dff_B_bXzx77a41_1),.clk(gclk));
	jdff dff_B_FMnajm8G4_1(.din(w_dff_B_bXzx77a41_1),.dout(w_dff_B_FMnajm8G4_1),.clk(gclk));
	jdff dff_B_ccdDxJkD0_1(.din(w_dff_B_FMnajm8G4_1),.dout(w_dff_B_ccdDxJkD0_1),.clk(gclk));
	jdff dff_B_XhRnvKZZ1_1(.din(w_dff_B_ccdDxJkD0_1),.dout(w_dff_B_XhRnvKZZ1_1),.clk(gclk));
	jdff dff_B_9Rx8xwna0_1(.din(w_dff_B_XhRnvKZZ1_1),.dout(w_dff_B_9Rx8xwna0_1),.clk(gclk));
	jdff dff_B_WIa8yhxu1_1(.din(w_dff_B_9Rx8xwna0_1),.dout(w_dff_B_WIa8yhxu1_1),.clk(gclk));
	jdff dff_B_hiyWUse81_1(.din(w_dff_B_WIa8yhxu1_1),.dout(w_dff_B_hiyWUse81_1),.clk(gclk));
	jdff dff_B_GrOBJnqH2_1(.din(w_dff_B_hiyWUse81_1),.dout(w_dff_B_GrOBJnqH2_1),.clk(gclk));
	jdff dff_B_u8g1M5HO3_1(.din(w_dff_B_GrOBJnqH2_1),.dout(w_dff_B_u8g1M5HO3_1),.clk(gclk));
	jdff dff_B_3KcMjNye2_1(.din(w_dff_B_u8g1M5HO3_1),.dout(w_dff_B_3KcMjNye2_1),.clk(gclk));
	jdff dff_B_DM0c2Tpp5_1(.din(w_dff_B_3KcMjNye2_1),.dout(w_dff_B_DM0c2Tpp5_1),.clk(gclk));
	jdff dff_B_TP5Shjm96_1(.din(w_dff_B_DM0c2Tpp5_1),.dout(w_dff_B_TP5Shjm96_1),.clk(gclk));
	jdff dff_B_OB4DEuRr8_1(.din(w_dff_B_TP5Shjm96_1),.dout(w_dff_B_OB4DEuRr8_1),.clk(gclk));
	jdff dff_B_G1KyZF0M8_1(.din(w_dff_B_OB4DEuRr8_1),.dout(w_dff_B_G1KyZF0M8_1),.clk(gclk));
	jdff dff_B_T7dveuQ82_1(.din(w_dff_B_G1KyZF0M8_1),.dout(w_dff_B_T7dveuQ82_1),.clk(gclk));
	jdff dff_A_C95lVcqm2_0(.dout(w_n282_0[0]),.din(w_dff_A_C95lVcqm2_0),.clk(gclk));
	jdff dff_A_Vi6tqybi3_0(.dout(w_n226_0[0]),.din(w_dff_A_Vi6tqybi3_0),.clk(gclk));
	jdff dff_A_J7xmdvLm9_0(.dout(w_dff_A_Vi6tqybi3_0),.din(w_dff_A_J7xmdvLm9_0),.clk(gclk));
	jdff dff_A_wcUSb0ND0_0(.dout(w_dff_A_J7xmdvLm9_0),.din(w_dff_A_wcUSb0ND0_0),.clk(gclk));
	jdff dff_A_DUiltiON6_0(.dout(w_dff_A_wcUSb0ND0_0),.din(w_dff_A_DUiltiON6_0),.clk(gclk));
	jdff dff_A_ZR8UbXeW8_0(.dout(w_dff_A_DUiltiON6_0),.din(w_dff_A_ZR8UbXeW8_0),.clk(gclk));
	jdff dff_A_vdIwsETk7_0(.dout(w_dff_A_ZR8UbXeW8_0),.din(w_dff_A_vdIwsETk7_0),.clk(gclk));
	jdff dff_A_y6UBtydD0_0(.dout(w_dff_A_vdIwsETk7_0),.din(w_dff_A_y6UBtydD0_0),.clk(gclk));
	jdff dff_A_CgEma8ZJ4_0(.dout(w_dff_A_y6UBtydD0_0),.din(w_dff_A_CgEma8ZJ4_0),.clk(gclk));
	jdff dff_A_gl5Qt2Ot8_0(.dout(w_dff_A_CgEma8ZJ4_0),.din(w_dff_A_gl5Qt2Ot8_0),.clk(gclk));
	jdff dff_A_7mv1w4M16_0(.dout(w_dff_A_gl5Qt2Ot8_0),.din(w_dff_A_7mv1w4M16_0),.clk(gclk));
	jdff dff_A_yxy9RVM56_0(.dout(w_dff_A_7mv1w4M16_0),.din(w_dff_A_yxy9RVM56_0),.clk(gclk));
	jdff dff_A_cH4aSYDU7_0(.dout(w_dff_A_yxy9RVM56_0),.din(w_dff_A_cH4aSYDU7_0),.clk(gclk));
	jdff dff_A_hKqXMD9c0_0(.dout(w_dff_A_cH4aSYDU7_0),.din(w_dff_A_hKqXMD9c0_0),.clk(gclk));
	jdff dff_A_kNtRzy8m2_0(.dout(w_dff_A_hKqXMD9c0_0),.din(w_dff_A_kNtRzy8m2_0),.clk(gclk));
	jdff dff_A_7G13RT427_0(.dout(w_dff_A_kNtRzy8m2_0),.din(w_dff_A_7G13RT427_0),.clk(gclk));
	jdff dff_A_AQFbMP098_0(.dout(w_dff_A_7G13RT427_0),.din(w_dff_A_AQFbMP098_0),.clk(gclk));
	jdff dff_B_oWFygZgG2_1(.din(n233),.dout(w_dff_B_oWFygZgG2_1),.clk(gclk));
	jdff dff_B_akbrEpRE8_1(.din(w_dff_B_oWFygZgG2_1),.dout(w_dff_B_akbrEpRE8_1),.clk(gclk));
	jdff dff_B_YiAkGpZx9_1(.din(w_dff_B_akbrEpRE8_1),.dout(w_dff_B_YiAkGpZx9_1),.clk(gclk));
	jdff dff_B_quKfcrm47_1(.din(w_dff_B_YiAkGpZx9_1),.dout(w_dff_B_quKfcrm47_1),.clk(gclk));
	jdff dff_B_TuJdajx77_1(.din(w_dff_B_quKfcrm47_1),.dout(w_dff_B_TuJdajx77_1),.clk(gclk));
	jdff dff_B_1WAubDVB4_1(.din(w_dff_B_TuJdajx77_1),.dout(w_dff_B_1WAubDVB4_1),.clk(gclk));
	jdff dff_B_nwwEBhyz4_1(.din(w_dff_B_1WAubDVB4_1),.dout(w_dff_B_nwwEBhyz4_1),.clk(gclk));
	jdff dff_B_zMEQz6ua2_1(.din(w_dff_B_nwwEBhyz4_1),.dout(w_dff_B_zMEQz6ua2_1),.clk(gclk));
	jdff dff_B_VDUySVi49_1(.din(w_dff_B_zMEQz6ua2_1),.dout(w_dff_B_VDUySVi49_1),.clk(gclk));
	jdff dff_B_UFQIP7y21_1(.din(w_dff_B_VDUySVi49_1),.dout(w_dff_B_UFQIP7y21_1),.clk(gclk));
	jdff dff_B_judfDY4v3_1(.din(w_dff_B_UFQIP7y21_1),.dout(w_dff_B_judfDY4v3_1),.clk(gclk));
	jdff dff_B_iS1z2tby3_1(.din(w_dff_B_judfDY4v3_1),.dout(w_dff_B_iS1z2tby3_1),.clk(gclk));
	jdff dff_B_RUOdUyiF6_1(.din(w_dff_B_iS1z2tby3_1),.dout(w_dff_B_RUOdUyiF6_1),.clk(gclk));
	jdff dff_A_oDeo4JQK6_0(.dout(w_n231_0[0]),.din(w_dff_A_oDeo4JQK6_0),.clk(gclk));
	jdff dff_A_l3pzBfjS2_0(.dout(w_n183_0[0]),.din(w_dff_A_l3pzBfjS2_0),.clk(gclk));
	jdff dff_A_cjgpqF0p3_0(.dout(w_dff_A_l3pzBfjS2_0),.din(w_dff_A_cjgpqF0p3_0),.clk(gclk));
	jdff dff_A_uOyZRKLN6_0(.dout(w_dff_A_cjgpqF0p3_0),.din(w_dff_A_uOyZRKLN6_0),.clk(gclk));
	jdff dff_A_xjTL6E8p5_0(.dout(w_dff_A_uOyZRKLN6_0),.din(w_dff_A_xjTL6E8p5_0),.clk(gclk));
	jdff dff_A_11UYdMps8_0(.dout(w_dff_A_xjTL6E8p5_0),.din(w_dff_A_11UYdMps8_0),.clk(gclk));
	jdff dff_A_Xh5PV9FL2_0(.dout(w_dff_A_11UYdMps8_0),.din(w_dff_A_Xh5PV9FL2_0),.clk(gclk));
	jdff dff_A_3chRoaCD9_0(.dout(w_dff_A_Xh5PV9FL2_0),.din(w_dff_A_3chRoaCD9_0),.clk(gclk));
	jdff dff_A_gcf6QSsY4_0(.dout(w_dff_A_3chRoaCD9_0),.din(w_dff_A_gcf6QSsY4_0),.clk(gclk));
	jdff dff_A_z4wlQNNV1_0(.dout(w_dff_A_gcf6QSsY4_0),.din(w_dff_A_z4wlQNNV1_0),.clk(gclk));
	jdff dff_A_5rOWLprw6_0(.dout(w_dff_A_z4wlQNNV1_0),.din(w_dff_A_5rOWLprw6_0),.clk(gclk));
	jdff dff_A_SjSjZ8Cg4_0(.dout(w_dff_A_5rOWLprw6_0),.din(w_dff_A_SjSjZ8Cg4_0),.clk(gclk));
	jdff dff_A_Ok4TBqic0_0(.dout(w_dff_A_SjSjZ8Cg4_0),.din(w_dff_A_Ok4TBqic0_0),.clk(gclk));
	jdff dff_A_OVDrevzS6_0(.dout(w_dff_A_Ok4TBqic0_0),.din(w_dff_A_OVDrevzS6_0),.clk(gclk));
	jdff dff_A_mnSlSRY63_0(.dout(w_dff_A_OVDrevzS6_0),.din(w_dff_A_mnSlSRY63_0),.clk(gclk));
	jdff dff_B_dRsffrHs6_1(.din(n190),.dout(w_dff_B_dRsffrHs6_1),.clk(gclk));
	jdff dff_B_hATEjAtW6_1(.din(w_dff_B_dRsffrHs6_1),.dout(w_dff_B_hATEjAtW6_1),.clk(gclk));
	jdff dff_B_jPMCi8ZN0_1(.din(w_dff_B_hATEjAtW6_1),.dout(w_dff_B_jPMCi8ZN0_1),.clk(gclk));
	jdff dff_B_EFirFdGd0_1(.din(w_dff_B_jPMCi8ZN0_1),.dout(w_dff_B_EFirFdGd0_1),.clk(gclk));
	jdff dff_B_FTL8EDBx4_1(.din(w_dff_B_EFirFdGd0_1),.dout(w_dff_B_FTL8EDBx4_1),.clk(gclk));
	jdff dff_B_wnoAgGL21_1(.din(w_dff_B_FTL8EDBx4_1),.dout(w_dff_B_wnoAgGL21_1),.clk(gclk));
	jdff dff_B_gIrIlQin4_1(.din(w_dff_B_wnoAgGL21_1),.dout(w_dff_B_gIrIlQin4_1),.clk(gclk));
	jdff dff_B_8VhK9wsb3_1(.din(w_dff_B_gIrIlQin4_1),.dout(w_dff_B_8VhK9wsb3_1),.clk(gclk));
	jdff dff_B_3S00F6qj7_1(.din(w_dff_B_8VhK9wsb3_1),.dout(w_dff_B_3S00F6qj7_1),.clk(gclk));
	jdff dff_B_E2bs8Qwu3_1(.din(w_dff_B_3S00F6qj7_1),.dout(w_dff_B_E2bs8Qwu3_1),.clk(gclk));
	jdff dff_B_FeQGZ0tg2_1(.din(w_dff_B_E2bs8Qwu3_1),.dout(w_dff_B_FeQGZ0tg2_1),.clk(gclk));
	jdff dff_A_LL0DfKUa1_0(.dout(w_n188_0[0]),.din(w_dff_A_LL0DfKUa1_0),.clk(gclk));
	jdff dff_A_lOlDLeYk8_0(.dout(w_n145_0[0]),.din(w_dff_A_lOlDLeYk8_0),.clk(gclk));
	jdff dff_A_qkiU0kGP6_0(.dout(w_dff_A_lOlDLeYk8_0),.din(w_dff_A_qkiU0kGP6_0),.clk(gclk));
	jdff dff_A_q0emCLJe2_0(.dout(w_dff_A_qkiU0kGP6_0),.din(w_dff_A_q0emCLJe2_0),.clk(gclk));
	jdff dff_A_PlsV4TOb8_0(.dout(w_dff_A_q0emCLJe2_0),.din(w_dff_A_PlsV4TOb8_0),.clk(gclk));
	jdff dff_A_J7J5Wt4u7_0(.dout(w_dff_A_PlsV4TOb8_0),.din(w_dff_A_J7J5Wt4u7_0),.clk(gclk));
	jdff dff_A_8vUDIetG5_0(.dout(w_dff_A_J7J5Wt4u7_0),.din(w_dff_A_8vUDIetG5_0),.clk(gclk));
	jdff dff_A_cl4f1fZh7_0(.dout(w_dff_A_8vUDIetG5_0),.din(w_dff_A_cl4f1fZh7_0),.clk(gclk));
	jdff dff_A_CP5ZuuGR5_0(.dout(w_dff_A_cl4f1fZh7_0),.din(w_dff_A_CP5ZuuGR5_0),.clk(gclk));
	jdff dff_A_3dqgACn87_0(.dout(w_dff_A_CP5ZuuGR5_0),.din(w_dff_A_3dqgACn87_0),.clk(gclk));
	jdff dff_A_G28ZyrZ98_0(.dout(w_dff_A_3dqgACn87_0),.din(w_dff_A_G28ZyrZ98_0),.clk(gclk));
	jdff dff_A_LcbbC6Gi6_0(.dout(w_dff_A_G28ZyrZ98_0),.din(w_dff_A_LcbbC6Gi6_0),.clk(gclk));
	jdff dff_A_7HPLrMCC8_0(.dout(w_dff_A_LcbbC6Gi6_0),.din(w_dff_A_7HPLrMCC8_0),.clk(gclk));
	jdff dff_B_zqWSIJpp8_1(.din(n152),.dout(w_dff_B_zqWSIJpp8_1),.clk(gclk));
	jdff dff_B_5XJ0MbIU3_1(.din(w_dff_B_zqWSIJpp8_1),.dout(w_dff_B_5XJ0MbIU3_1),.clk(gclk));
	jdff dff_B_0h3XU6Cx5_1(.din(w_dff_B_5XJ0MbIU3_1),.dout(w_dff_B_0h3XU6Cx5_1),.clk(gclk));
	jdff dff_B_jglCie9R7_1(.din(w_dff_B_0h3XU6Cx5_1),.dout(w_dff_B_jglCie9R7_1),.clk(gclk));
	jdff dff_B_IqNhxrqy8_1(.din(w_dff_B_jglCie9R7_1),.dout(w_dff_B_IqNhxrqy8_1),.clk(gclk));
	jdff dff_B_saczajSj6_1(.din(w_dff_B_IqNhxrqy8_1),.dout(w_dff_B_saczajSj6_1),.clk(gclk));
	jdff dff_B_i0kVo9my7_1(.din(w_dff_B_saczajSj6_1),.dout(w_dff_B_i0kVo9my7_1),.clk(gclk));
	jdff dff_B_AjzgUDJh3_1(.din(w_dff_B_i0kVo9my7_1),.dout(w_dff_B_AjzgUDJh3_1),.clk(gclk));
	jdff dff_B_26rhsQip6_1(.din(w_dff_B_AjzgUDJh3_1),.dout(w_dff_B_26rhsQip6_1),.clk(gclk));
	jdff dff_A_TenYRsws0_0(.dout(w_n150_0[0]),.din(w_dff_A_TenYRsws0_0),.clk(gclk));
	jdff dff_A_1Q843crG3_0(.dout(w_n110_0[0]),.din(w_dff_A_1Q843crG3_0),.clk(gclk));
	jdff dff_A_b4OC8tPc0_0(.dout(w_dff_A_1Q843crG3_0),.din(w_dff_A_b4OC8tPc0_0),.clk(gclk));
	jdff dff_A_6QYMP0Pm2_0(.dout(w_dff_A_b4OC8tPc0_0),.din(w_dff_A_6QYMP0Pm2_0),.clk(gclk));
	jdff dff_A_AOLB0mop3_0(.dout(w_dff_A_6QYMP0Pm2_0),.din(w_dff_A_AOLB0mop3_0),.clk(gclk));
	jdff dff_A_LsVDsME93_0(.dout(w_dff_A_AOLB0mop3_0),.din(w_dff_A_LsVDsME93_0),.clk(gclk));
	jdff dff_A_6rwN02mZ0_0(.dout(w_dff_A_LsVDsME93_0),.din(w_dff_A_6rwN02mZ0_0),.clk(gclk));
	jdff dff_A_JhvXPSSm7_0(.dout(w_dff_A_6rwN02mZ0_0),.din(w_dff_A_JhvXPSSm7_0),.clk(gclk));
	jdff dff_A_aDKKiVNS0_0(.dout(w_dff_A_JhvXPSSm7_0),.din(w_dff_A_aDKKiVNS0_0),.clk(gclk));
	jdff dff_A_wScBvGaT4_0(.dout(w_dff_A_aDKKiVNS0_0),.din(w_dff_A_wScBvGaT4_0),.clk(gclk));
	jdff dff_A_WdwwOVyQ8_0(.dout(w_dff_A_wScBvGaT4_0),.din(w_dff_A_WdwwOVyQ8_0),.clk(gclk));
	jdff dff_B_0fv5yjhA6_1(.din(n117),.dout(w_dff_B_0fv5yjhA6_1),.clk(gclk));
	jdff dff_B_I2hCNous3_1(.din(w_dff_B_0fv5yjhA6_1),.dout(w_dff_B_I2hCNous3_1),.clk(gclk));
	jdff dff_B_P9ACDME41_1(.din(w_dff_B_I2hCNous3_1),.dout(w_dff_B_P9ACDME41_1),.clk(gclk));
	jdff dff_B_Jq6Qy6BN0_1(.din(w_dff_B_P9ACDME41_1),.dout(w_dff_B_Jq6Qy6BN0_1),.clk(gclk));
	jdff dff_B_nCEzdcfE5_1(.din(w_dff_B_Jq6Qy6BN0_1),.dout(w_dff_B_nCEzdcfE5_1),.clk(gclk));
	jdff dff_B_JC0Y6Ui80_1(.din(w_dff_B_nCEzdcfE5_1),.dout(w_dff_B_JC0Y6Ui80_1),.clk(gclk));
	jdff dff_B_Wsh9ZRGM0_1(.din(w_dff_B_JC0Y6Ui80_1),.dout(w_dff_B_Wsh9ZRGM0_1),.clk(gclk));
	jdff dff_A_lXilLWhR4_0(.dout(w_n115_0[0]),.din(w_dff_A_lXilLWhR4_0),.clk(gclk));
	jdff dff_B_o082cFWp4_2(.din(n115),.dout(w_dff_B_o082cFWp4_2),.clk(gclk));
	jdff dff_A_1MrAJqss9_0(.dout(w_n89_0[0]),.din(w_dff_A_1MrAJqss9_0),.clk(gclk));
	jdff dff_A_XJmi4JZf0_0(.dout(w_dff_A_1MrAJqss9_0),.din(w_dff_A_XJmi4JZf0_0),.clk(gclk));
	jdff dff_A_TWDGeNcx3_0(.dout(w_dff_A_XJmi4JZf0_0),.din(w_dff_A_TWDGeNcx3_0),.clk(gclk));
	jdff dff_A_83xhQuQT4_0(.dout(w_dff_A_TWDGeNcx3_0),.din(w_dff_A_83xhQuQT4_0),.clk(gclk));
	jdff dff_A_PbFVMIW76_0(.dout(w_dff_A_83xhQuQT4_0),.din(w_dff_A_PbFVMIW76_0),.clk(gclk));
	jdff dff_A_qbIqQljw1_0(.dout(w_dff_A_PbFVMIW76_0),.din(w_dff_A_qbIqQljw1_0),.clk(gclk));
	jdff dff_A_Sb20tTNi4_0(.dout(w_dff_A_qbIqQljw1_0),.din(w_dff_A_Sb20tTNi4_0),.clk(gclk));
	jdff dff_B_97tUUQ5T3_1(.din(n95),.dout(w_dff_B_97tUUQ5T3_1),.clk(gclk));
	jdff dff_B_Ej0vGfTk0_1(.din(w_dff_B_97tUUQ5T3_1),.dout(w_dff_B_Ej0vGfTk0_1),.clk(gclk));
	jdff dff_B_1my9ggDg8_1(.din(w_dff_B_Ej0vGfTk0_1),.dout(w_dff_B_1my9ggDg8_1),.clk(gclk));
	jdff dff_B_RMpO3DLV2_1(.din(w_dff_B_1my9ggDg8_1),.dout(w_dff_B_RMpO3DLV2_1),.clk(gclk));
	jdff dff_A_QEwu1QkQ3_0(.dout(w_n93_0[0]),.din(w_dff_A_QEwu1QkQ3_0),.clk(gclk));
	jdff dff_B_jI2yWL6q9_2(.din(n93),.dout(w_dff_B_jI2yWL6q9_2),.clk(gclk));
	jdff dff_B_IDjAmrQo7_0(.din(n92),.dout(w_dff_B_IDjAmrQo7_0),.clk(gclk));
	jdff dff_A_xryOKzr28_0(.dout(w_n72_0[0]),.din(w_dff_A_xryOKzr28_0),.clk(gclk));
	jdff dff_A_GTirAPbm7_0(.dout(w_dff_A_xryOKzr28_0),.din(w_dff_A_GTirAPbm7_0),.clk(gclk));
	jdff dff_A_wr6o7ltw7_0(.dout(w_dff_A_GTirAPbm7_0),.din(w_dff_A_wr6o7ltw7_0),.clk(gclk));
	jdff dff_B_Zg4WHi4m7_0(.din(n83),.dout(w_dff_B_Zg4WHi4m7_0),.clk(gclk));
	jdff dff_A_PMzkp3Yy3_0(.dout(w_n69_0[0]),.din(w_dff_A_PMzkp3Yy3_0),.clk(gclk));
	jdff dff_A_iW07Qgb02_0(.dout(w_n1043_0[0]),.din(w_dff_A_iW07Qgb02_0),.clk(gclk));
	jdff dff_B_siiwXJJ18_2(.din(n1043),.dout(w_dff_B_siiwXJJ18_2),.clk(gclk));
	jdff dff_A_JALddgvv6_1(.dout(w_n938_0[1]),.din(w_dff_A_JALddgvv6_1),.clk(gclk));
	jdff dff_B_ceVyse8u0_2(.din(n938),.dout(w_dff_B_ceVyse8u0_2),.clk(gclk));
	jdff dff_B_OsKKAQx83_2(.din(w_dff_B_ceVyse8u0_2),.dout(w_dff_B_OsKKAQx83_2),.clk(gclk));
	jdff dff_B_Iznw8x703_2(.din(w_dff_B_OsKKAQx83_2),.dout(w_dff_B_Iznw8x703_2),.clk(gclk));
	jdff dff_B_o0OJDUGi4_2(.din(w_dff_B_Iznw8x703_2),.dout(w_dff_B_o0OJDUGi4_2),.clk(gclk));
	jdff dff_B_zOABYoD24_2(.din(w_dff_B_o0OJDUGi4_2),.dout(w_dff_B_zOABYoD24_2),.clk(gclk));
	jdff dff_B_eCn0dC6B2_2(.din(w_dff_B_zOABYoD24_2),.dout(w_dff_B_eCn0dC6B2_2),.clk(gclk));
	jdff dff_B_QnGobxNJ1_2(.din(w_dff_B_eCn0dC6B2_2),.dout(w_dff_B_QnGobxNJ1_2),.clk(gclk));
	jdff dff_B_pyBbdSKc3_2(.din(w_dff_B_QnGobxNJ1_2),.dout(w_dff_B_pyBbdSKc3_2),.clk(gclk));
	jdff dff_B_4dwZJS6X4_2(.din(w_dff_B_pyBbdSKc3_2),.dout(w_dff_B_4dwZJS6X4_2),.clk(gclk));
	jdff dff_B_i9d2Xck33_2(.din(w_dff_B_4dwZJS6X4_2),.dout(w_dff_B_i9d2Xck33_2),.clk(gclk));
	jdff dff_B_v8FSVbER3_2(.din(w_dff_B_i9d2Xck33_2),.dout(w_dff_B_v8FSVbER3_2),.clk(gclk));
	jdff dff_B_GnhrRIJZ1_2(.din(w_dff_B_v8FSVbER3_2),.dout(w_dff_B_GnhrRIJZ1_2),.clk(gclk));
	jdff dff_B_InpRgIT89_2(.din(w_dff_B_GnhrRIJZ1_2),.dout(w_dff_B_InpRgIT89_2),.clk(gclk));
	jdff dff_B_rlSwGTiB2_2(.din(w_dff_B_InpRgIT89_2),.dout(w_dff_B_rlSwGTiB2_2),.clk(gclk));
	jdff dff_B_025hKoW00_2(.din(w_dff_B_rlSwGTiB2_2),.dout(w_dff_B_025hKoW00_2),.clk(gclk));
	jdff dff_B_uAvGqAgU4_2(.din(w_dff_B_025hKoW00_2),.dout(w_dff_B_uAvGqAgU4_2),.clk(gclk));
	jdff dff_B_ei0xRJXx8_2(.din(w_dff_B_uAvGqAgU4_2),.dout(w_dff_B_ei0xRJXx8_2),.clk(gclk));
	jdff dff_B_jrIUrfQ32_2(.din(w_dff_B_ei0xRJXx8_2),.dout(w_dff_B_jrIUrfQ32_2),.clk(gclk));
	jdff dff_B_ptRYBJqs3_2(.din(w_dff_B_jrIUrfQ32_2),.dout(w_dff_B_ptRYBJqs3_2),.clk(gclk));
	jdff dff_B_aIr8GCuP4_2(.din(w_dff_B_ptRYBJqs3_2),.dout(w_dff_B_aIr8GCuP4_2),.clk(gclk));
	jdff dff_B_wKgyXslP4_2(.din(w_dff_B_aIr8GCuP4_2),.dout(w_dff_B_wKgyXslP4_2),.clk(gclk));
	jdff dff_B_Xd26Q48Y8_2(.din(w_dff_B_wKgyXslP4_2),.dout(w_dff_B_Xd26Q48Y8_2),.clk(gclk));
	jdff dff_B_6hAmRQfI3_2(.din(w_dff_B_Xd26Q48Y8_2),.dout(w_dff_B_6hAmRQfI3_2),.clk(gclk));
	jdff dff_B_LbHddnH23_2(.din(w_dff_B_6hAmRQfI3_2),.dout(w_dff_B_LbHddnH23_2),.clk(gclk));
	jdff dff_B_ifMVYr991_2(.din(w_dff_B_LbHddnH23_2),.dout(w_dff_B_ifMVYr991_2),.clk(gclk));
	jdff dff_B_rv5wyhox2_2(.din(w_dff_B_ifMVYr991_2),.dout(w_dff_B_rv5wyhox2_2),.clk(gclk));
	jdff dff_B_EQrBiNvS3_2(.din(w_dff_B_rv5wyhox2_2),.dout(w_dff_B_EQrBiNvS3_2),.clk(gclk));
	jdff dff_B_se56qiBO2_2(.din(w_dff_B_EQrBiNvS3_2),.dout(w_dff_B_se56qiBO2_2),.clk(gclk));
	jdff dff_B_HLMsBhxG1_2(.din(w_dff_B_se56qiBO2_2),.dout(w_dff_B_HLMsBhxG1_2),.clk(gclk));
	jdff dff_B_z7aPTPIf2_2(.din(w_dff_B_HLMsBhxG1_2),.dout(w_dff_B_z7aPTPIf2_2),.clk(gclk));
	jdff dff_B_wQLZOnu17_2(.din(w_dff_B_z7aPTPIf2_2),.dout(w_dff_B_wQLZOnu17_2),.clk(gclk));
	jdff dff_B_kWfNUNAt5_2(.din(w_dff_B_wQLZOnu17_2),.dout(w_dff_B_kWfNUNAt5_2),.clk(gclk));
	jdff dff_A_i1clNZ0m9_1(.dout(w_n942_0[1]),.din(w_dff_A_i1clNZ0m9_1),.clk(gclk));
	jdff dff_A_um8ltIX04_2(.dout(w_n942_0[2]),.din(w_dff_A_um8ltIX04_2),.clk(gclk));
	jdff dff_B_kLnAW15u8_3(.din(n942),.dout(w_dff_B_kLnAW15u8_3),.clk(gclk));
	jdff dff_B_fPYh2NFM3_2(.din(n835),.dout(w_dff_B_fPYh2NFM3_2),.clk(gclk));
	jdff dff_B_PAx0Mzac1_2(.din(w_dff_B_fPYh2NFM3_2),.dout(w_dff_B_PAx0Mzac1_2),.clk(gclk));
	jdff dff_B_nnX5S40d4_2(.din(w_dff_B_PAx0Mzac1_2),.dout(w_dff_B_nnX5S40d4_2),.clk(gclk));
	jdff dff_B_nKHf3q6X9_2(.din(w_dff_B_nnX5S40d4_2),.dout(w_dff_B_nKHf3q6X9_2),.clk(gclk));
	jdff dff_B_1lRvW5IM7_2(.din(w_dff_B_nKHf3q6X9_2),.dout(w_dff_B_1lRvW5IM7_2),.clk(gclk));
	jdff dff_B_Br75LXZQ4_2(.din(w_dff_B_1lRvW5IM7_2),.dout(w_dff_B_Br75LXZQ4_2),.clk(gclk));
	jdff dff_B_foy3zvNv4_2(.din(w_dff_B_Br75LXZQ4_2),.dout(w_dff_B_foy3zvNv4_2),.clk(gclk));
	jdff dff_B_uvZJOAsb5_2(.din(w_dff_B_foy3zvNv4_2),.dout(w_dff_B_uvZJOAsb5_2),.clk(gclk));
	jdff dff_B_0Oqemyyk9_2(.din(w_dff_B_uvZJOAsb5_2),.dout(w_dff_B_0Oqemyyk9_2),.clk(gclk));
	jdff dff_B_gJUKotO98_2(.din(w_dff_B_0Oqemyyk9_2),.dout(w_dff_B_gJUKotO98_2),.clk(gclk));
	jdff dff_B_pSOEjo3U0_2(.din(w_dff_B_gJUKotO98_2),.dout(w_dff_B_pSOEjo3U0_2),.clk(gclk));
	jdff dff_B_gp322aiT5_2(.din(w_dff_B_pSOEjo3U0_2),.dout(w_dff_B_gp322aiT5_2),.clk(gclk));
	jdff dff_B_Ngf8tBR99_2(.din(w_dff_B_gp322aiT5_2),.dout(w_dff_B_Ngf8tBR99_2),.clk(gclk));
	jdff dff_B_HpgOyv5H4_2(.din(w_dff_B_Ngf8tBR99_2),.dout(w_dff_B_HpgOyv5H4_2),.clk(gclk));
	jdff dff_B_1vt9VwUq3_2(.din(w_dff_B_HpgOyv5H4_2),.dout(w_dff_B_1vt9VwUq3_2),.clk(gclk));
	jdff dff_B_WuLWAwiU6_2(.din(w_dff_B_1vt9VwUq3_2),.dout(w_dff_B_WuLWAwiU6_2),.clk(gclk));
	jdff dff_B_bkDjcfUG8_2(.din(w_dff_B_WuLWAwiU6_2),.dout(w_dff_B_bkDjcfUG8_2),.clk(gclk));
	jdff dff_B_DLD2mCQd1_2(.din(w_dff_B_bkDjcfUG8_2),.dout(w_dff_B_DLD2mCQd1_2),.clk(gclk));
	jdff dff_B_lZUU5Ikp7_2(.din(w_dff_B_DLD2mCQd1_2),.dout(w_dff_B_lZUU5Ikp7_2),.clk(gclk));
	jdff dff_B_NNYrsWlx4_2(.din(w_dff_B_lZUU5Ikp7_2),.dout(w_dff_B_NNYrsWlx4_2),.clk(gclk));
	jdff dff_B_0HmUS0n64_2(.din(w_dff_B_NNYrsWlx4_2),.dout(w_dff_B_0HmUS0n64_2),.clk(gclk));
	jdff dff_B_4umjEWuQ9_2(.din(w_dff_B_0HmUS0n64_2),.dout(w_dff_B_4umjEWuQ9_2),.clk(gclk));
	jdff dff_B_cgk9FrNK0_2(.din(w_dff_B_4umjEWuQ9_2),.dout(w_dff_B_cgk9FrNK0_2),.clk(gclk));
	jdff dff_B_oaxqtx8w6_2(.din(w_dff_B_cgk9FrNK0_2),.dout(w_dff_B_oaxqtx8w6_2),.clk(gclk));
	jdff dff_B_av554reE0_2(.din(w_dff_B_oaxqtx8w6_2),.dout(w_dff_B_av554reE0_2),.clk(gclk));
	jdff dff_B_bH9gXNBM5_2(.din(w_dff_B_av554reE0_2),.dout(w_dff_B_bH9gXNBM5_2),.clk(gclk));
	jdff dff_B_0x9xVjx69_2(.din(w_dff_B_bH9gXNBM5_2),.dout(w_dff_B_0x9xVjx69_2),.clk(gclk));
	jdff dff_B_wPE0grvz8_2(.din(w_dff_B_0x9xVjx69_2),.dout(w_dff_B_wPE0grvz8_2),.clk(gclk));
	jdff dff_B_ik6tOIxU0_2(.din(w_dff_B_wPE0grvz8_2),.dout(w_dff_B_ik6tOIxU0_2),.clk(gclk));
	jdff dff_B_HA4refMf4_1(.din(n841),.dout(w_dff_B_HA4refMf4_1),.clk(gclk));
	jdff dff_B_yZmTFvSo7_1(.din(w_dff_B_HA4refMf4_1),.dout(w_dff_B_yZmTFvSo7_1),.clk(gclk));
	jdff dff_B_GMRb3hFM3_1(.din(w_dff_B_yZmTFvSo7_1),.dout(w_dff_B_GMRb3hFM3_1),.clk(gclk));
	jdff dff_B_DBFYvmrq9_1(.din(w_dff_B_GMRb3hFM3_1),.dout(w_dff_B_DBFYvmrq9_1),.clk(gclk));
	jdff dff_B_LyUd0YqQ7_1(.din(w_dff_B_DBFYvmrq9_1),.dout(w_dff_B_LyUd0YqQ7_1),.clk(gclk));
	jdff dff_B_mlbQyOMs1_1(.din(w_dff_B_LyUd0YqQ7_1),.dout(w_dff_B_mlbQyOMs1_1),.clk(gclk));
	jdff dff_B_5eZA3ChM6_1(.din(w_dff_B_mlbQyOMs1_1),.dout(w_dff_B_5eZA3ChM6_1),.clk(gclk));
	jdff dff_B_gWK2mxjU5_1(.din(w_dff_B_5eZA3ChM6_1),.dout(w_dff_B_gWK2mxjU5_1),.clk(gclk));
	jdff dff_B_Cd67rXIQ7_1(.din(w_dff_B_gWK2mxjU5_1),.dout(w_dff_B_Cd67rXIQ7_1),.clk(gclk));
	jdff dff_B_ZJLVSupR9_1(.din(w_dff_B_Cd67rXIQ7_1),.dout(w_dff_B_ZJLVSupR9_1),.clk(gclk));
	jdff dff_B_g2KoK8Yr2_1(.din(w_dff_B_ZJLVSupR9_1),.dout(w_dff_B_g2KoK8Yr2_1),.clk(gclk));
	jdff dff_B_6u0lKJHd8_1(.din(w_dff_B_g2KoK8Yr2_1),.dout(w_dff_B_6u0lKJHd8_1),.clk(gclk));
	jdff dff_B_ZT7sgB5c1_1(.din(w_dff_B_6u0lKJHd8_1),.dout(w_dff_B_ZT7sgB5c1_1),.clk(gclk));
	jdff dff_B_6EABTwI58_1(.din(w_dff_B_ZT7sgB5c1_1),.dout(w_dff_B_6EABTwI58_1),.clk(gclk));
	jdff dff_B_xLco0Nea9_1(.din(w_dff_B_6EABTwI58_1),.dout(w_dff_B_xLco0Nea9_1),.clk(gclk));
	jdff dff_B_oldjHmBk3_1(.din(w_dff_B_xLco0Nea9_1),.dout(w_dff_B_oldjHmBk3_1),.clk(gclk));
	jdff dff_B_r7WWhIwN8_1(.din(w_dff_B_oldjHmBk3_1),.dout(w_dff_B_r7WWhIwN8_1),.clk(gclk));
	jdff dff_B_Enw8Q78Y7_1(.din(w_dff_B_r7WWhIwN8_1),.dout(w_dff_B_Enw8Q78Y7_1),.clk(gclk));
	jdff dff_B_zQASk2fe0_1(.din(w_dff_B_Enw8Q78Y7_1),.dout(w_dff_B_zQASk2fe0_1),.clk(gclk));
	jdff dff_B_lt3OFEtz3_1(.din(w_dff_B_zQASk2fe0_1),.dout(w_dff_B_lt3OFEtz3_1),.clk(gclk));
	jdff dff_B_P3wPA5Ou0_1(.din(w_dff_B_lt3OFEtz3_1),.dout(w_dff_B_P3wPA5Ou0_1),.clk(gclk));
	jdff dff_B_uKVyaURs6_1(.din(w_dff_B_P3wPA5Ou0_1),.dout(w_dff_B_uKVyaURs6_1),.clk(gclk));
	jdff dff_B_VDgJkdLD4_1(.din(w_dff_B_uKVyaURs6_1),.dout(w_dff_B_VDgJkdLD4_1),.clk(gclk));
	jdff dff_B_eDn57moe7_1(.din(w_dff_B_VDgJkdLD4_1),.dout(w_dff_B_eDn57moe7_1),.clk(gclk));
	jdff dff_B_UcabbIXb5_1(.din(w_dff_B_eDn57moe7_1),.dout(w_dff_B_UcabbIXb5_1),.clk(gclk));
	jdff dff_B_GNqgMNCd9_1(.din(w_dff_B_UcabbIXb5_1),.dout(w_dff_B_GNqgMNCd9_1),.clk(gclk));
	jdff dff_A_13aE2Vnd9_0(.dout(w_n839_0[0]),.din(w_dff_A_13aE2Vnd9_0),.clk(gclk));
	jdff dff_A_YAHfWe8j5_0(.dout(w_n735_0[0]),.din(w_dff_A_YAHfWe8j5_0),.clk(gclk));
	jdff dff_A_FaZnX2s07_0(.dout(w_dff_A_YAHfWe8j5_0),.din(w_dff_A_FaZnX2s07_0),.clk(gclk));
	jdff dff_A_H2SMGDSo1_0(.dout(w_dff_A_FaZnX2s07_0),.din(w_dff_A_H2SMGDSo1_0),.clk(gclk));
	jdff dff_A_yNDvrETi5_0(.dout(w_dff_A_H2SMGDSo1_0),.din(w_dff_A_yNDvrETi5_0),.clk(gclk));
	jdff dff_A_pfrkrKcp0_0(.dout(w_dff_A_yNDvrETi5_0),.din(w_dff_A_pfrkrKcp0_0),.clk(gclk));
	jdff dff_A_dziXrN4W6_0(.dout(w_dff_A_pfrkrKcp0_0),.din(w_dff_A_dziXrN4W6_0),.clk(gclk));
	jdff dff_A_ES0o6cA46_0(.dout(w_dff_A_dziXrN4W6_0),.din(w_dff_A_ES0o6cA46_0),.clk(gclk));
	jdff dff_A_UXAfSEdm3_0(.dout(w_dff_A_ES0o6cA46_0),.din(w_dff_A_UXAfSEdm3_0),.clk(gclk));
	jdff dff_A_pN94njs06_0(.dout(w_dff_A_UXAfSEdm3_0),.din(w_dff_A_pN94njs06_0),.clk(gclk));
	jdff dff_A_zTvoK0eo4_0(.dout(w_dff_A_pN94njs06_0),.din(w_dff_A_zTvoK0eo4_0),.clk(gclk));
	jdff dff_A_9Rvc39fk1_0(.dout(w_dff_A_zTvoK0eo4_0),.din(w_dff_A_9Rvc39fk1_0),.clk(gclk));
	jdff dff_A_dyuGMICT6_0(.dout(w_dff_A_9Rvc39fk1_0),.din(w_dff_A_dyuGMICT6_0),.clk(gclk));
	jdff dff_A_0omNt4yn0_0(.dout(w_dff_A_dyuGMICT6_0),.din(w_dff_A_0omNt4yn0_0),.clk(gclk));
	jdff dff_A_0PqGSUCa3_0(.dout(w_dff_A_0omNt4yn0_0),.din(w_dff_A_0PqGSUCa3_0),.clk(gclk));
	jdff dff_A_dzeWzO6E8_0(.dout(w_dff_A_0PqGSUCa3_0),.din(w_dff_A_dzeWzO6E8_0),.clk(gclk));
	jdff dff_A_InvzsMxT5_0(.dout(w_dff_A_dzeWzO6E8_0),.din(w_dff_A_InvzsMxT5_0),.clk(gclk));
	jdff dff_A_e07vjjwd8_0(.dout(w_dff_A_InvzsMxT5_0),.din(w_dff_A_e07vjjwd8_0),.clk(gclk));
	jdff dff_A_7VtgAFAC2_0(.dout(w_dff_A_e07vjjwd8_0),.din(w_dff_A_7VtgAFAC2_0),.clk(gclk));
	jdff dff_A_Bxd7xzdy4_0(.dout(w_dff_A_7VtgAFAC2_0),.din(w_dff_A_Bxd7xzdy4_0),.clk(gclk));
	jdff dff_A_xODHA9ah0_0(.dout(w_dff_A_Bxd7xzdy4_0),.din(w_dff_A_xODHA9ah0_0),.clk(gclk));
	jdff dff_A_pRMp635i8_0(.dout(w_dff_A_xODHA9ah0_0),.din(w_dff_A_pRMp635i8_0),.clk(gclk));
	jdff dff_A_yFeeqo8i6_0(.dout(w_dff_A_pRMp635i8_0),.din(w_dff_A_yFeeqo8i6_0),.clk(gclk));
	jdff dff_A_D1OIFUbg3_0(.dout(w_dff_A_yFeeqo8i6_0),.din(w_dff_A_D1OIFUbg3_0),.clk(gclk));
	jdff dff_A_3RniC67G8_0(.dout(w_dff_A_D1OIFUbg3_0),.din(w_dff_A_3RniC67G8_0),.clk(gclk));
	jdff dff_A_GQ7TLWlX5_0(.dout(w_dff_A_3RniC67G8_0),.din(w_dff_A_GQ7TLWlX5_0),.clk(gclk));
	jdff dff_A_nn8qURut8_0(.dout(w_dff_A_GQ7TLWlX5_0),.din(w_dff_A_nn8qURut8_0),.clk(gclk));
	jdff dff_A_ll4vw5e71_0(.dout(w_dff_A_nn8qURut8_0),.din(w_dff_A_ll4vw5e71_0),.clk(gclk));
	jdff dff_A_ISoQoaIJ1_1(.dout(w_n740_0[1]),.din(w_dff_A_ISoQoaIJ1_1),.clk(gclk));
	jdff dff_A_kazzux2u8_2(.dout(w_n740_0[2]),.din(w_dff_A_kazzux2u8_2),.clk(gclk));
	jdff dff_A_w9HYr66J4_0(.dout(w_n642_0[0]),.din(w_dff_A_w9HYr66J4_0),.clk(gclk));
	jdff dff_A_FvSOP7KV6_0(.dout(w_dff_A_w9HYr66J4_0),.din(w_dff_A_FvSOP7KV6_0),.clk(gclk));
	jdff dff_A_43N3vsTT3_0(.dout(w_dff_A_FvSOP7KV6_0),.din(w_dff_A_43N3vsTT3_0),.clk(gclk));
	jdff dff_A_ZYupGxZ83_0(.dout(w_dff_A_43N3vsTT3_0),.din(w_dff_A_ZYupGxZ83_0),.clk(gclk));
	jdff dff_A_RxGa3VIE9_0(.dout(w_dff_A_ZYupGxZ83_0),.din(w_dff_A_RxGa3VIE9_0),.clk(gclk));
	jdff dff_A_2z9WHNuB5_0(.dout(w_dff_A_RxGa3VIE9_0),.din(w_dff_A_2z9WHNuB5_0),.clk(gclk));
	jdff dff_A_uezb728w2_0(.dout(w_dff_A_2z9WHNuB5_0),.din(w_dff_A_uezb728w2_0),.clk(gclk));
	jdff dff_A_6NSavQqV6_0(.dout(w_dff_A_uezb728w2_0),.din(w_dff_A_6NSavQqV6_0),.clk(gclk));
	jdff dff_A_URIAhbao3_0(.dout(w_dff_A_6NSavQqV6_0),.din(w_dff_A_URIAhbao3_0),.clk(gclk));
	jdff dff_A_Jd59PiaD2_0(.dout(w_dff_A_URIAhbao3_0),.din(w_dff_A_Jd59PiaD2_0),.clk(gclk));
	jdff dff_A_94EPOhq03_0(.dout(w_dff_A_Jd59PiaD2_0),.din(w_dff_A_94EPOhq03_0),.clk(gclk));
	jdff dff_A_iR2uoyDP3_0(.dout(w_dff_A_94EPOhq03_0),.din(w_dff_A_iR2uoyDP3_0),.clk(gclk));
	jdff dff_A_5U2JcT4S6_0(.dout(w_dff_A_iR2uoyDP3_0),.din(w_dff_A_5U2JcT4S6_0),.clk(gclk));
	jdff dff_A_wFlYTjpM2_0(.dout(w_dff_A_5U2JcT4S6_0),.din(w_dff_A_wFlYTjpM2_0),.clk(gclk));
	jdff dff_A_yAoCe94R7_0(.dout(w_dff_A_wFlYTjpM2_0),.din(w_dff_A_yAoCe94R7_0),.clk(gclk));
	jdff dff_A_jNh70a8Q7_0(.dout(w_dff_A_yAoCe94R7_0),.din(w_dff_A_jNh70a8Q7_0),.clk(gclk));
	jdff dff_A_JTQib3Qa8_0(.dout(w_dff_A_jNh70a8Q7_0),.din(w_dff_A_JTQib3Qa8_0),.clk(gclk));
	jdff dff_A_0CrUDDpE8_0(.dout(w_dff_A_JTQib3Qa8_0),.din(w_dff_A_0CrUDDpE8_0),.clk(gclk));
	jdff dff_A_GqDjidEL4_0(.dout(w_dff_A_0CrUDDpE8_0),.din(w_dff_A_GqDjidEL4_0),.clk(gclk));
	jdff dff_A_VvkpVXp26_0(.dout(w_dff_A_GqDjidEL4_0),.din(w_dff_A_VvkpVXp26_0),.clk(gclk));
	jdff dff_A_HdapZFwp5_0(.dout(w_dff_A_VvkpVXp26_0),.din(w_dff_A_HdapZFwp5_0),.clk(gclk));
	jdff dff_A_uXtBycX77_0(.dout(w_dff_A_HdapZFwp5_0),.din(w_dff_A_uXtBycX77_0),.clk(gclk));
	jdff dff_A_2HHX7coE5_0(.dout(w_dff_A_uXtBycX77_0),.din(w_dff_A_2HHX7coE5_0),.clk(gclk));
	jdff dff_A_Y4EtgO005_0(.dout(w_dff_A_2HHX7coE5_0),.din(w_dff_A_Y4EtgO005_0),.clk(gclk));
	jdff dff_A_5ewLWf1x3_0(.dout(w_dff_A_Y4EtgO005_0),.din(w_dff_A_5ewLWf1x3_0),.clk(gclk));
	jdff dff_A_aYMwcFEq6_1(.dout(w_n647_0[1]),.din(w_dff_A_aYMwcFEq6_1),.clk(gclk));
	jdff dff_A_LtNAu88Z7_2(.dout(w_n647_0[2]),.din(w_dff_A_LtNAu88Z7_2),.clk(gclk));
	jdff dff_A_5F9DBEBA3_0(.dout(w_n556_0[0]),.din(w_dff_A_5F9DBEBA3_0),.clk(gclk));
	jdff dff_A_ULQI3dSY5_0(.dout(w_dff_A_5F9DBEBA3_0),.din(w_dff_A_ULQI3dSY5_0),.clk(gclk));
	jdff dff_A_mcrDvY0w8_0(.dout(w_dff_A_ULQI3dSY5_0),.din(w_dff_A_mcrDvY0w8_0),.clk(gclk));
	jdff dff_A_QeZdjYpp7_0(.dout(w_dff_A_mcrDvY0w8_0),.din(w_dff_A_QeZdjYpp7_0),.clk(gclk));
	jdff dff_A_2vJFH7uA8_0(.dout(w_dff_A_QeZdjYpp7_0),.din(w_dff_A_2vJFH7uA8_0),.clk(gclk));
	jdff dff_A_sGGiRhdj8_0(.dout(w_dff_A_2vJFH7uA8_0),.din(w_dff_A_sGGiRhdj8_0),.clk(gclk));
	jdff dff_A_mqLqVPta6_0(.dout(w_dff_A_sGGiRhdj8_0),.din(w_dff_A_mqLqVPta6_0),.clk(gclk));
	jdff dff_A_i2KBoIBi3_0(.dout(w_dff_A_mqLqVPta6_0),.din(w_dff_A_i2KBoIBi3_0),.clk(gclk));
	jdff dff_A_6AF8tcGX9_0(.dout(w_dff_A_i2KBoIBi3_0),.din(w_dff_A_6AF8tcGX9_0),.clk(gclk));
	jdff dff_A_r3rrGcI09_0(.dout(w_dff_A_6AF8tcGX9_0),.din(w_dff_A_r3rrGcI09_0),.clk(gclk));
	jdff dff_A_drMLmGCL9_0(.dout(w_dff_A_r3rrGcI09_0),.din(w_dff_A_drMLmGCL9_0),.clk(gclk));
	jdff dff_A_1FeyGtDE7_0(.dout(w_dff_A_drMLmGCL9_0),.din(w_dff_A_1FeyGtDE7_0),.clk(gclk));
	jdff dff_A_FCif0Lax2_0(.dout(w_dff_A_1FeyGtDE7_0),.din(w_dff_A_FCif0Lax2_0),.clk(gclk));
	jdff dff_A_Ap4mlANs3_0(.dout(w_dff_A_FCif0Lax2_0),.din(w_dff_A_Ap4mlANs3_0),.clk(gclk));
	jdff dff_A_4oDZ1FCG0_0(.dout(w_dff_A_Ap4mlANs3_0),.din(w_dff_A_4oDZ1FCG0_0),.clk(gclk));
	jdff dff_A_YCP7jMKP2_0(.dout(w_dff_A_4oDZ1FCG0_0),.din(w_dff_A_YCP7jMKP2_0),.clk(gclk));
	jdff dff_A_cksGFkhz1_0(.dout(w_dff_A_YCP7jMKP2_0),.din(w_dff_A_cksGFkhz1_0),.clk(gclk));
	jdff dff_A_91wyghiS6_0(.dout(w_dff_A_cksGFkhz1_0),.din(w_dff_A_91wyghiS6_0),.clk(gclk));
	jdff dff_A_TjezKelA1_0(.dout(w_dff_A_91wyghiS6_0),.din(w_dff_A_TjezKelA1_0),.clk(gclk));
	jdff dff_A_zeQpUz4m8_0(.dout(w_dff_A_TjezKelA1_0),.din(w_dff_A_zeQpUz4m8_0),.clk(gclk));
	jdff dff_A_3hgz5e1J0_0(.dout(w_dff_A_zeQpUz4m8_0),.din(w_dff_A_3hgz5e1J0_0),.clk(gclk));
	jdff dff_A_ULEY2Xh70_0(.dout(w_dff_A_3hgz5e1J0_0),.din(w_dff_A_ULEY2Xh70_0),.clk(gclk));
	jdff dff_A_feTdm7cL9_0(.dout(w_dff_A_ULEY2Xh70_0),.din(w_dff_A_feTdm7cL9_0),.clk(gclk));
	jdff dff_A_GDWe2Ed28_1(.dout(w_n561_0[1]),.din(w_dff_A_GDWe2Ed28_1),.clk(gclk));
	jdff dff_A_pUePyb2f4_2(.dout(w_n561_0[2]),.din(w_dff_A_pUePyb2f4_2),.clk(gclk));
	jdff dff_A_JZWCuGl19_0(.dout(w_n477_0[0]),.din(w_dff_A_JZWCuGl19_0),.clk(gclk));
	jdff dff_A_sYtQ0rJq6_0(.dout(w_dff_A_JZWCuGl19_0),.din(w_dff_A_sYtQ0rJq6_0),.clk(gclk));
	jdff dff_A_x9rTQskC1_0(.dout(w_dff_A_sYtQ0rJq6_0),.din(w_dff_A_x9rTQskC1_0),.clk(gclk));
	jdff dff_A_iy4Thptt3_0(.dout(w_dff_A_x9rTQskC1_0),.din(w_dff_A_iy4Thptt3_0),.clk(gclk));
	jdff dff_A_CSWz8Rh16_0(.dout(w_dff_A_iy4Thptt3_0),.din(w_dff_A_CSWz8Rh16_0),.clk(gclk));
	jdff dff_A_NUknB0YH3_0(.dout(w_dff_A_CSWz8Rh16_0),.din(w_dff_A_NUknB0YH3_0),.clk(gclk));
	jdff dff_A_3mMAn5rP5_0(.dout(w_dff_A_NUknB0YH3_0),.din(w_dff_A_3mMAn5rP5_0),.clk(gclk));
	jdff dff_A_yzmVGExE3_0(.dout(w_dff_A_3mMAn5rP5_0),.din(w_dff_A_yzmVGExE3_0),.clk(gclk));
	jdff dff_A_KZ4RsuBW9_0(.dout(w_dff_A_yzmVGExE3_0),.din(w_dff_A_KZ4RsuBW9_0),.clk(gclk));
	jdff dff_A_7MMh2dfC4_0(.dout(w_dff_A_KZ4RsuBW9_0),.din(w_dff_A_7MMh2dfC4_0),.clk(gclk));
	jdff dff_A_7wMD8lrW8_0(.dout(w_dff_A_7MMh2dfC4_0),.din(w_dff_A_7wMD8lrW8_0),.clk(gclk));
	jdff dff_A_tTEfOe8G8_0(.dout(w_dff_A_7wMD8lrW8_0),.din(w_dff_A_tTEfOe8G8_0),.clk(gclk));
	jdff dff_A_G3tY7b388_0(.dout(w_dff_A_tTEfOe8G8_0),.din(w_dff_A_G3tY7b388_0),.clk(gclk));
	jdff dff_A_cP4hdsTT3_0(.dout(w_dff_A_G3tY7b388_0),.din(w_dff_A_cP4hdsTT3_0),.clk(gclk));
	jdff dff_A_3umympik8_0(.dout(w_dff_A_cP4hdsTT3_0),.din(w_dff_A_3umympik8_0),.clk(gclk));
	jdff dff_A_MHytO7VT9_0(.dout(w_dff_A_3umympik8_0),.din(w_dff_A_MHytO7VT9_0),.clk(gclk));
	jdff dff_A_Rj0u3L2Y5_0(.dout(w_dff_A_MHytO7VT9_0),.din(w_dff_A_Rj0u3L2Y5_0),.clk(gclk));
	jdff dff_A_jmfQ601j5_0(.dout(w_dff_A_Rj0u3L2Y5_0),.din(w_dff_A_jmfQ601j5_0),.clk(gclk));
	jdff dff_A_ZBgEBTYf0_0(.dout(w_dff_A_jmfQ601j5_0),.din(w_dff_A_ZBgEBTYf0_0),.clk(gclk));
	jdff dff_A_YZK69PiR5_0(.dout(w_dff_A_ZBgEBTYf0_0),.din(w_dff_A_YZK69PiR5_0),.clk(gclk));
	jdff dff_A_779Ly5To1_0(.dout(w_dff_A_YZK69PiR5_0),.din(w_dff_A_779Ly5To1_0),.clk(gclk));
	jdff dff_A_iwf7vElC1_1(.dout(w_n482_0[1]),.din(w_dff_A_iwf7vElC1_1),.clk(gclk));
	jdff dff_A_px4TwLna7_2(.dout(w_n482_0[2]),.din(w_dff_A_px4TwLna7_2),.clk(gclk));
	jdff dff_A_jCGIzMeG0_0(.dout(w_n405_0[0]),.din(w_dff_A_jCGIzMeG0_0),.clk(gclk));
	jdff dff_A_rpLt9Fpd9_0(.dout(w_dff_A_jCGIzMeG0_0),.din(w_dff_A_rpLt9Fpd9_0),.clk(gclk));
	jdff dff_A_SPxXuECE0_0(.dout(w_dff_A_rpLt9Fpd9_0),.din(w_dff_A_SPxXuECE0_0),.clk(gclk));
	jdff dff_A_hxWcnJCZ1_0(.dout(w_dff_A_SPxXuECE0_0),.din(w_dff_A_hxWcnJCZ1_0),.clk(gclk));
	jdff dff_A_xlmJTAOT8_0(.dout(w_dff_A_hxWcnJCZ1_0),.din(w_dff_A_xlmJTAOT8_0),.clk(gclk));
	jdff dff_A_jkvjEAHl9_0(.dout(w_dff_A_xlmJTAOT8_0),.din(w_dff_A_jkvjEAHl9_0),.clk(gclk));
	jdff dff_A_ufkRC2n31_0(.dout(w_dff_A_jkvjEAHl9_0),.din(w_dff_A_ufkRC2n31_0),.clk(gclk));
	jdff dff_A_d0r6oMcr7_0(.dout(w_dff_A_ufkRC2n31_0),.din(w_dff_A_d0r6oMcr7_0),.clk(gclk));
	jdff dff_A_YErHK3kd8_0(.dout(w_dff_A_d0r6oMcr7_0),.din(w_dff_A_YErHK3kd8_0),.clk(gclk));
	jdff dff_A_5u1Lgjg41_0(.dout(w_dff_A_YErHK3kd8_0),.din(w_dff_A_5u1Lgjg41_0),.clk(gclk));
	jdff dff_A_Fe2vuQfG0_0(.dout(w_dff_A_5u1Lgjg41_0),.din(w_dff_A_Fe2vuQfG0_0),.clk(gclk));
	jdff dff_A_5Lex8d2O2_0(.dout(w_dff_A_Fe2vuQfG0_0),.din(w_dff_A_5Lex8d2O2_0),.clk(gclk));
	jdff dff_A_VOALqQ4k4_0(.dout(w_dff_A_5Lex8d2O2_0),.din(w_dff_A_VOALqQ4k4_0),.clk(gclk));
	jdff dff_A_3Ld9aSWl2_0(.dout(w_dff_A_VOALqQ4k4_0),.din(w_dff_A_3Ld9aSWl2_0),.clk(gclk));
	jdff dff_A_WKJmnlms2_0(.dout(w_dff_A_3Ld9aSWl2_0),.din(w_dff_A_WKJmnlms2_0),.clk(gclk));
	jdff dff_A_IYWSJVUQ9_0(.dout(w_dff_A_WKJmnlms2_0),.din(w_dff_A_IYWSJVUQ9_0),.clk(gclk));
	jdff dff_A_zbRK0Ysn1_0(.dout(w_dff_A_IYWSJVUQ9_0),.din(w_dff_A_zbRK0Ysn1_0),.clk(gclk));
	jdff dff_A_4QQPTkHp1_0(.dout(w_dff_A_zbRK0Ysn1_0),.din(w_dff_A_4QQPTkHp1_0),.clk(gclk));
	jdff dff_A_lXR94XaA4_0(.dout(w_dff_A_4QQPTkHp1_0),.din(w_dff_A_lXR94XaA4_0),.clk(gclk));
	jdff dff_A_vf10omxW1_1(.dout(w_n410_0[1]),.din(w_dff_A_vf10omxW1_1),.clk(gclk));
	jdff dff_A_v08tLeep6_2(.dout(w_n410_0[2]),.din(w_dff_A_v08tLeep6_2),.clk(gclk));
	jdff dff_A_7KpPilju2_0(.dout(w_n341_0[0]),.din(w_dff_A_7KpPilju2_0),.clk(gclk));
	jdff dff_A_NIqqc0Ox9_0(.dout(w_dff_A_7KpPilju2_0),.din(w_dff_A_NIqqc0Ox9_0),.clk(gclk));
	jdff dff_A_SL4UvMG77_0(.dout(w_dff_A_NIqqc0Ox9_0),.din(w_dff_A_SL4UvMG77_0),.clk(gclk));
	jdff dff_A_OqRlkAhm3_0(.dout(w_dff_A_SL4UvMG77_0),.din(w_dff_A_OqRlkAhm3_0),.clk(gclk));
	jdff dff_A_R5IRv6W95_0(.dout(w_dff_A_OqRlkAhm3_0),.din(w_dff_A_R5IRv6W95_0),.clk(gclk));
	jdff dff_A_Hz6uWMmA8_0(.dout(w_dff_A_R5IRv6W95_0),.din(w_dff_A_Hz6uWMmA8_0),.clk(gclk));
	jdff dff_A_mHD4qWy89_0(.dout(w_dff_A_Hz6uWMmA8_0),.din(w_dff_A_mHD4qWy89_0),.clk(gclk));
	jdff dff_A_qmhBJOhA2_0(.dout(w_dff_A_mHD4qWy89_0),.din(w_dff_A_qmhBJOhA2_0),.clk(gclk));
	jdff dff_A_wQRDciC92_0(.dout(w_dff_A_qmhBJOhA2_0),.din(w_dff_A_wQRDciC92_0),.clk(gclk));
	jdff dff_A_MhQHdx9g9_0(.dout(w_dff_A_wQRDciC92_0),.din(w_dff_A_MhQHdx9g9_0),.clk(gclk));
	jdff dff_A_OMXtVIoo1_0(.dout(w_dff_A_MhQHdx9g9_0),.din(w_dff_A_OMXtVIoo1_0),.clk(gclk));
	jdff dff_A_87BUSuyJ4_0(.dout(w_dff_A_OMXtVIoo1_0),.din(w_dff_A_87BUSuyJ4_0),.clk(gclk));
	jdff dff_A_QmHmyN2l0_0(.dout(w_dff_A_87BUSuyJ4_0),.din(w_dff_A_QmHmyN2l0_0),.clk(gclk));
	jdff dff_A_tS1iXJKm9_0(.dout(w_dff_A_QmHmyN2l0_0),.din(w_dff_A_tS1iXJKm9_0),.clk(gclk));
	jdff dff_A_3JV8DRYs3_0(.dout(w_dff_A_tS1iXJKm9_0),.din(w_dff_A_3JV8DRYs3_0),.clk(gclk));
	jdff dff_A_oToKoT7i0_0(.dout(w_dff_A_3JV8DRYs3_0),.din(w_dff_A_oToKoT7i0_0),.clk(gclk));
	jdff dff_A_bzzSIQF31_0(.dout(w_dff_A_oToKoT7i0_0),.din(w_dff_A_bzzSIQF31_0),.clk(gclk));
	jdff dff_A_eQlOczic5_1(.dout(w_n346_0[1]),.din(w_dff_A_eQlOczic5_1),.clk(gclk));
	jdff dff_A_H17Bjt2h2_2(.dout(w_n346_0[2]),.din(w_dff_A_H17Bjt2h2_2),.clk(gclk));
	jdff dff_A_Cqizgbsw6_0(.dout(w_n283_0[0]),.din(w_dff_A_Cqizgbsw6_0),.clk(gclk));
	jdff dff_A_0pRyf39E5_0(.dout(w_dff_A_Cqizgbsw6_0),.din(w_dff_A_0pRyf39E5_0),.clk(gclk));
	jdff dff_A_pqGuvdBE5_0(.dout(w_dff_A_0pRyf39E5_0),.din(w_dff_A_pqGuvdBE5_0),.clk(gclk));
	jdff dff_A_shhzMjQP6_0(.dout(w_dff_A_pqGuvdBE5_0),.din(w_dff_A_shhzMjQP6_0),.clk(gclk));
	jdff dff_A_uNRnbGGr9_0(.dout(w_dff_A_shhzMjQP6_0),.din(w_dff_A_uNRnbGGr9_0),.clk(gclk));
	jdff dff_A_E78EoQLH3_0(.dout(w_dff_A_uNRnbGGr9_0),.din(w_dff_A_E78EoQLH3_0),.clk(gclk));
	jdff dff_A_nHOhTHfi1_0(.dout(w_dff_A_E78EoQLH3_0),.din(w_dff_A_nHOhTHfi1_0),.clk(gclk));
	jdff dff_A_F6zJR4kQ6_0(.dout(w_dff_A_nHOhTHfi1_0),.din(w_dff_A_F6zJR4kQ6_0),.clk(gclk));
	jdff dff_A_O73bvBUS0_0(.dout(w_dff_A_F6zJR4kQ6_0),.din(w_dff_A_O73bvBUS0_0),.clk(gclk));
	jdff dff_A_CZPRDBnR1_0(.dout(w_dff_A_O73bvBUS0_0),.din(w_dff_A_CZPRDBnR1_0),.clk(gclk));
	jdff dff_A_80NxXhQH0_0(.dout(w_dff_A_CZPRDBnR1_0),.din(w_dff_A_80NxXhQH0_0),.clk(gclk));
	jdff dff_A_CoyyZRJp0_0(.dout(w_dff_A_80NxXhQH0_0),.din(w_dff_A_CoyyZRJp0_0),.clk(gclk));
	jdff dff_A_p0w8nkSi7_0(.dout(w_dff_A_CoyyZRJp0_0),.din(w_dff_A_p0w8nkSi7_0),.clk(gclk));
	jdff dff_A_1lpFeTQs8_0(.dout(w_dff_A_p0w8nkSi7_0),.din(w_dff_A_1lpFeTQs8_0),.clk(gclk));
	jdff dff_A_Oeb4iY3b9_0(.dout(w_dff_A_1lpFeTQs8_0),.din(w_dff_A_Oeb4iY3b9_0),.clk(gclk));
	jdff dff_A_dKDe0QPZ5_1(.dout(w_n288_0[1]),.din(w_dff_A_dKDe0QPZ5_1),.clk(gclk));
	jdff dff_A_DvKWN5fh7_2(.dout(w_n288_0[2]),.din(w_dff_A_DvKWN5fh7_2),.clk(gclk));
	jdff dff_A_tDG3Qnmk9_0(.dout(w_n232_0[0]),.din(w_dff_A_tDG3Qnmk9_0),.clk(gclk));
	jdff dff_A_690nUmZT2_0(.dout(w_dff_A_tDG3Qnmk9_0),.din(w_dff_A_690nUmZT2_0),.clk(gclk));
	jdff dff_A_6UXU6NRh0_0(.dout(w_dff_A_690nUmZT2_0),.din(w_dff_A_6UXU6NRh0_0),.clk(gclk));
	jdff dff_A_GKJYzaP06_0(.dout(w_dff_A_6UXU6NRh0_0),.din(w_dff_A_GKJYzaP06_0),.clk(gclk));
	jdff dff_A_RtLgvyqS8_0(.dout(w_dff_A_GKJYzaP06_0),.din(w_dff_A_RtLgvyqS8_0),.clk(gclk));
	jdff dff_A_wGPX2W1j9_0(.dout(w_dff_A_RtLgvyqS8_0),.din(w_dff_A_wGPX2W1j9_0),.clk(gclk));
	jdff dff_A_2zAM49FT7_0(.dout(w_dff_A_wGPX2W1j9_0),.din(w_dff_A_2zAM49FT7_0),.clk(gclk));
	jdff dff_A_OZtLM20K6_0(.dout(w_dff_A_2zAM49FT7_0),.din(w_dff_A_OZtLM20K6_0),.clk(gclk));
	jdff dff_A_RDdpvEL42_0(.dout(w_dff_A_OZtLM20K6_0),.din(w_dff_A_RDdpvEL42_0),.clk(gclk));
	jdff dff_A_scRUgCMK7_0(.dout(w_dff_A_RDdpvEL42_0),.din(w_dff_A_scRUgCMK7_0),.clk(gclk));
	jdff dff_A_4rljsAHQ6_0(.dout(w_dff_A_scRUgCMK7_0),.din(w_dff_A_4rljsAHQ6_0),.clk(gclk));
	jdff dff_A_YkYi6GKM5_0(.dout(w_dff_A_4rljsAHQ6_0),.din(w_dff_A_YkYi6GKM5_0),.clk(gclk));
	jdff dff_A_2UH2CFTH9_0(.dout(w_dff_A_YkYi6GKM5_0),.din(w_dff_A_2UH2CFTH9_0),.clk(gclk));
	jdff dff_A_3RUgPuw28_1(.dout(w_n237_0[1]),.din(w_dff_A_3RUgPuw28_1),.clk(gclk));
	jdff dff_A_X5hDfQDj5_2(.dout(w_n237_0[2]),.din(w_dff_A_X5hDfQDj5_2),.clk(gclk));
	jdff dff_A_W75uVNnM6_0(.dout(w_n189_0[0]),.din(w_dff_A_W75uVNnM6_0),.clk(gclk));
	jdff dff_A_8ty9nFLM9_0(.dout(w_dff_A_W75uVNnM6_0),.din(w_dff_A_8ty9nFLM9_0),.clk(gclk));
	jdff dff_A_9hHzXBpl7_0(.dout(w_dff_A_8ty9nFLM9_0),.din(w_dff_A_9hHzXBpl7_0),.clk(gclk));
	jdff dff_A_q2pGvRuu9_0(.dout(w_dff_A_9hHzXBpl7_0),.din(w_dff_A_q2pGvRuu9_0),.clk(gclk));
	jdff dff_A_v8v8RMUX2_0(.dout(w_dff_A_q2pGvRuu9_0),.din(w_dff_A_v8v8RMUX2_0),.clk(gclk));
	jdff dff_A_eazA6Cty5_0(.dout(w_dff_A_v8v8RMUX2_0),.din(w_dff_A_eazA6Cty5_0),.clk(gclk));
	jdff dff_A_KDhbOBns9_0(.dout(w_dff_A_eazA6Cty5_0),.din(w_dff_A_KDhbOBns9_0),.clk(gclk));
	jdff dff_A_2nedHdpN9_0(.dout(w_dff_A_KDhbOBns9_0),.din(w_dff_A_2nedHdpN9_0),.clk(gclk));
	jdff dff_A_xMkIFcHq0_0(.dout(w_dff_A_2nedHdpN9_0),.din(w_dff_A_xMkIFcHq0_0),.clk(gclk));
	jdff dff_A_gZJZmRfP0_0(.dout(w_dff_A_xMkIFcHq0_0),.din(w_dff_A_gZJZmRfP0_0),.clk(gclk));
	jdff dff_A_qj5HAMpT0_0(.dout(w_dff_A_gZJZmRfP0_0),.din(w_dff_A_qj5HAMpT0_0),.clk(gclk));
	jdff dff_A_0Nvok6OE8_1(.dout(w_n194_0[1]),.din(w_dff_A_0Nvok6OE8_1),.clk(gclk));
	jdff dff_A_sokiXTn82_2(.dout(w_n194_0[2]),.din(w_dff_A_sokiXTn82_2),.clk(gclk));
	jdff dff_A_nFyGUYEd9_0(.dout(w_n151_0[0]),.din(w_dff_A_nFyGUYEd9_0),.clk(gclk));
	jdff dff_A_U3fbiXAi7_0(.dout(w_dff_A_nFyGUYEd9_0),.din(w_dff_A_U3fbiXAi7_0),.clk(gclk));
	jdff dff_A_AvZ2IZj87_0(.dout(w_dff_A_U3fbiXAi7_0),.din(w_dff_A_AvZ2IZj87_0),.clk(gclk));
	jdff dff_A_JTcRza669_0(.dout(w_dff_A_AvZ2IZj87_0),.din(w_dff_A_JTcRza669_0),.clk(gclk));
	jdff dff_A_ojmxpyhq6_0(.dout(w_dff_A_JTcRza669_0),.din(w_dff_A_ojmxpyhq6_0),.clk(gclk));
	jdff dff_A_tXUz8pSJ5_0(.dout(w_dff_A_ojmxpyhq6_0),.din(w_dff_A_tXUz8pSJ5_0),.clk(gclk));
	jdff dff_A_wTMA7ou45_0(.dout(w_dff_A_tXUz8pSJ5_0),.din(w_dff_A_wTMA7ou45_0),.clk(gclk));
	jdff dff_A_s6i9fVwp6_0(.dout(w_dff_A_wTMA7ou45_0),.din(w_dff_A_s6i9fVwp6_0),.clk(gclk));
	jdff dff_A_ZbpznAsK3_0(.dout(w_dff_A_s6i9fVwp6_0),.din(w_dff_A_ZbpznAsK3_0),.clk(gclk));
	jdff dff_A_GAQ3BWky2_1(.dout(w_n156_0[1]),.din(w_dff_A_GAQ3BWky2_1),.clk(gclk));
	jdff dff_A_4x3nTySY4_2(.dout(w_n156_0[2]),.din(w_dff_A_4x3nTySY4_2),.clk(gclk));
	jdff dff_A_dgQ2v7Ka8_0(.dout(w_n116_0[0]),.din(w_dff_A_dgQ2v7Ka8_0),.clk(gclk));
	jdff dff_A_obEASgJV0_0(.dout(w_dff_A_dgQ2v7Ka8_0),.din(w_dff_A_obEASgJV0_0),.clk(gclk));
	jdff dff_A_THC7F6sj7_0(.dout(w_dff_A_obEASgJV0_0),.din(w_dff_A_THC7F6sj7_0),.clk(gclk));
	jdff dff_A_HKkXdrLj4_0(.dout(w_dff_A_THC7F6sj7_0),.din(w_dff_A_HKkXdrLj4_0),.clk(gclk));
	jdff dff_A_ictpUbM78_0(.dout(w_dff_A_HKkXdrLj4_0),.din(w_dff_A_ictpUbM78_0),.clk(gclk));
	jdff dff_A_YbNHwdYE6_0(.dout(w_dff_A_ictpUbM78_0),.din(w_dff_A_YbNHwdYE6_0),.clk(gclk));
	jdff dff_A_SAPjTpMh1_0(.dout(w_dff_A_YbNHwdYE6_0),.din(w_dff_A_SAPjTpMh1_0),.clk(gclk));
	jdff dff_A_bOg8qe9P3_1(.dout(w_n126_0[1]),.din(w_dff_A_bOg8qe9P3_1),.clk(gclk));
	jdff dff_A_bfPY2yka7_2(.dout(w_n126_0[2]),.din(w_dff_A_bfPY2yka7_2),.clk(gclk));
	jdff dff_B_qgd5TmgI4_3(.din(n126),.dout(w_dff_B_qgd5TmgI4_3),.clk(gclk));
	jdff dff_B_qFGeQJ162_3(.din(w_dff_B_qgd5TmgI4_3),.dout(w_dff_B_qFGeQJ162_3),.clk(gclk));
	jdff dff_B_1uWchztE5_0(.din(n122),.dout(w_dff_B_1uWchztE5_0),.clk(gclk));
	jdff dff_A_mSXE5txn7_0(.dout(w_n94_0[0]),.din(w_dff_A_mSXE5txn7_0),.clk(gclk));
	jdff dff_A_7hvl0jIi3_0(.dout(w_dff_A_mSXE5txn7_0),.din(w_dff_A_7hvl0jIi3_0),.clk(gclk));
	jdff dff_A_yoFFnUwE3_0(.dout(w_dff_A_7hvl0jIi3_0),.din(w_dff_A_yoFFnUwE3_0),.clk(gclk));
	jdff dff_A_dJ1rZgd00_1(.dout(w_n103_0[1]),.din(w_dff_A_dJ1rZgd00_1),.clk(gclk));
	jdff dff_B_26h76l4t0_1(.din(n97),.dout(w_dff_B_26h76l4t0_1),.clk(gclk));
	jdff dff_B_cbfshor35_1(.din(w_dff_B_26h76l4t0_1),.dout(w_dff_B_cbfshor35_1),.clk(gclk));
	jdff dff_A_b7ZXtC620_1(.dout(w_n82_0[1]),.din(w_dff_A_b7ZXtC620_1),.clk(gclk));
	jdff dff_A_EwX7zqbr3_2(.dout(w_n82_0[2]),.din(w_dff_A_EwX7zqbr3_2),.clk(gclk));
	jdff dff_A_XQ7rHGXI6_2(.dout(w_dff_A_EwX7zqbr3_2),.din(w_dff_A_XQ7rHGXI6_2),.clk(gclk));
	jdff dff_A_2RGpeNmG4_0(.dout(w_n1151_0[0]),.din(w_dff_A_2RGpeNmG4_0),.clk(gclk));
	jdff dff_B_j4T0AgN81_2(.din(n1151),.dout(w_dff_B_j4T0AgN81_2),.clk(gclk));
	jdff dff_B_bYJNWGcp4_2(.din(w_dff_B_j4T0AgN81_2),.dout(w_dff_B_bYJNWGcp4_2),.clk(gclk));
	jdff dff_B_DfRfJ3bK4_2(.din(n1044),.dout(w_dff_B_DfRfJ3bK4_2),.clk(gclk));
	jdff dff_B_xV3L2C6S0_2(.din(w_dff_B_DfRfJ3bK4_2),.dout(w_dff_B_xV3L2C6S0_2),.clk(gclk));
	jdff dff_B_mU8KX2pU1_2(.din(w_dff_B_xV3L2C6S0_2),.dout(w_dff_B_mU8KX2pU1_2),.clk(gclk));
	jdff dff_B_IK3LcRcX8_2(.din(w_dff_B_mU8KX2pU1_2),.dout(w_dff_B_IK3LcRcX8_2),.clk(gclk));
	jdff dff_B_54wJsXCZ3_2(.din(w_dff_B_IK3LcRcX8_2),.dout(w_dff_B_54wJsXCZ3_2),.clk(gclk));
	jdff dff_B_8YgzDuj16_2(.din(w_dff_B_54wJsXCZ3_2),.dout(w_dff_B_8YgzDuj16_2),.clk(gclk));
	jdff dff_B_NEZyEFb88_2(.din(w_dff_B_8YgzDuj16_2),.dout(w_dff_B_NEZyEFb88_2),.clk(gclk));
	jdff dff_B_XHM7RemR6_2(.din(w_dff_B_NEZyEFb88_2),.dout(w_dff_B_XHM7RemR6_2),.clk(gclk));
	jdff dff_B_jd7RMWTP8_2(.din(w_dff_B_XHM7RemR6_2),.dout(w_dff_B_jd7RMWTP8_2),.clk(gclk));
	jdff dff_B_W2ZBHAkE5_2(.din(w_dff_B_jd7RMWTP8_2),.dout(w_dff_B_W2ZBHAkE5_2),.clk(gclk));
	jdff dff_B_Lm9OBGLG8_2(.din(w_dff_B_W2ZBHAkE5_2),.dout(w_dff_B_Lm9OBGLG8_2),.clk(gclk));
	jdff dff_B_rcAybTle5_2(.din(w_dff_B_Lm9OBGLG8_2),.dout(w_dff_B_rcAybTle5_2),.clk(gclk));
	jdff dff_B_PRFY7O3c9_2(.din(w_dff_B_rcAybTle5_2),.dout(w_dff_B_PRFY7O3c9_2),.clk(gclk));
	jdff dff_B_vERN2gaO2_2(.din(w_dff_B_PRFY7O3c9_2),.dout(w_dff_B_vERN2gaO2_2),.clk(gclk));
	jdff dff_B_PfR96urB4_2(.din(w_dff_B_vERN2gaO2_2),.dout(w_dff_B_PfR96urB4_2),.clk(gclk));
	jdff dff_B_5hoGElMA3_2(.din(w_dff_B_PfR96urB4_2),.dout(w_dff_B_5hoGElMA3_2),.clk(gclk));
	jdff dff_B_JI5mF0TP6_2(.din(w_dff_B_5hoGElMA3_2),.dout(w_dff_B_JI5mF0TP6_2),.clk(gclk));
	jdff dff_B_Zt7e1kpL2_2(.din(w_dff_B_JI5mF0TP6_2),.dout(w_dff_B_Zt7e1kpL2_2),.clk(gclk));
	jdff dff_B_05M2yTSO5_2(.din(w_dff_B_Zt7e1kpL2_2),.dout(w_dff_B_05M2yTSO5_2),.clk(gclk));
	jdff dff_B_zeXRbp1R3_2(.din(w_dff_B_05M2yTSO5_2),.dout(w_dff_B_zeXRbp1R3_2),.clk(gclk));
	jdff dff_B_HuYJehbf1_2(.din(w_dff_B_zeXRbp1R3_2),.dout(w_dff_B_HuYJehbf1_2),.clk(gclk));
	jdff dff_B_vtapNQv04_2(.din(w_dff_B_HuYJehbf1_2),.dout(w_dff_B_vtapNQv04_2),.clk(gclk));
	jdff dff_B_w2uM7Xjk0_2(.din(w_dff_B_vtapNQv04_2),.dout(w_dff_B_w2uM7Xjk0_2),.clk(gclk));
	jdff dff_B_7z2LuFvy4_2(.din(w_dff_B_w2uM7Xjk0_2),.dout(w_dff_B_7z2LuFvy4_2),.clk(gclk));
	jdff dff_B_ir2jp4YY3_2(.din(w_dff_B_7z2LuFvy4_2),.dout(w_dff_B_ir2jp4YY3_2),.clk(gclk));
	jdff dff_B_LTz5XWUz2_2(.din(w_dff_B_ir2jp4YY3_2),.dout(w_dff_B_LTz5XWUz2_2),.clk(gclk));
	jdff dff_B_fINgTJaq6_2(.din(w_dff_B_LTz5XWUz2_2),.dout(w_dff_B_fINgTJaq6_2),.clk(gclk));
	jdff dff_B_uOvMuQMc7_2(.din(w_dff_B_fINgTJaq6_2),.dout(w_dff_B_uOvMuQMc7_2),.clk(gclk));
	jdff dff_B_871vyg922_2(.din(w_dff_B_uOvMuQMc7_2),.dout(w_dff_B_871vyg922_2),.clk(gclk));
	jdff dff_B_mE1Zy2sU9_2(.din(w_dff_B_871vyg922_2),.dout(w_dff_B_mE1Zy2sU9_2),.clk(gclk));
	jdff dff_B_XkFNPjeQ5_2(.din(w_dff_B_mE1Zy2sU9_2),.dout(w_dff_B_XkFNPjeQ5_2),.clk(gclk));
	jdff dff_B_G2YSEwb05_2(.din(w_dff_B_XkFNPjeQ5_2),.dout(w_dff_B_G2YSEwb05_2),.clk(gclk));
	jdff dff_B_etIzj5896_2(.din(w_dff_B_G2YSEwb05_2),.dout(w_dff_B_etIzj5896_2),.clk(gclk));
	jdff dff_A_rMaboMKD7_0(.dout(w_n1048_0[0]),.din(w_dff_A_rMaboMKD7_0),.clk(gclk));
	jdff dff_B_ZcdfPDIP9_2(.din(n1048),.dout(w_dff_B_ZcdfPDIP9_2),.clk(gclk));
	jdff dff_B_zEAdWz9j7_1(.din(n1046),.dout(w_dff_B_zEAdWz9j7_1),.clk(gclk));
	jdff dff_B_uxGb2FZw7_2(.din(n943),.dout(w_dff_B_uxGb2FZw7_2),.clk(gclk));
	jdff dff_B_0CtX2aQn8_2(.din(w_dff_B_uxGb2FZw7_2),.dout(w_dff_B_0CtX2aQn8_2),.clk(gclk));
	jdff dff_B_gqI3gs5R0_2(.din(w_dff_B_0CtX2aQn8_2),.dout(w_dff_B_gqI3gs5R0_2),.clk(gclk));
	jdff dff_B_pOqvpxto7_2(.din(w_dff_B_gqI3gs5R0_2),.dout(w_dff_B_pOqvpxto7_2),.clk(gclk));
	jdff dff_B_GM9vxiVN6_2(.din(w_dff_B_pOqvpxto7_2),.dout(w_dff_B_GM9vxiVN6_2),.clk(gclk));
	jdff dff_B_TDJCfjJJ0_2(.din(w_dff_B_GM9vxiVN6_2),.dout(w_dff_B_TDJCfjJJ0_2),.clk(gclk));
	jdff dff_B_MbLQsQzu0_2(.din(w_dff_B_TDJCfjJJ0_2),.dout(w_dff_B_MbLQsQzu0_2),.clk(gclk));
	jdff dff_B_LdHs9k6t2_2(.din(w_dff_B_MbLQsQzu0_2),.dout(w_dff_B_LdHs9k6t2_2),.clk(gclk));
	jdff dff_B_7Z7WrGWx9_2(.din(w_dff_B_LdHs9k6t2_2),.dout(w_dff_B_7Z7WrGWx9_2),.clk(gclk));
	jdff dff_B_DKYmxXIN1_2(.din(w_dff_B_7Z7WrGWx9_2),.dout(w_dff_B_DKYmxXIN1_2),.clk(gclk));
	jdff dff_B_8pENd0yE5_2(.din(w_dff_B_DKYmxXIN1_2),.dout(w_dff_B_8pENd0yE5_2),.clk(gclk));
	jdff dff_B_DV7KcakJ4_2(.din(w_dff_B_8pENd0yE5_2),.dout(w_dff_B_DV7KcakJ4_2),.clk(gclk));
	jdff dff_B_5G5O4tAY5_2(.din(w_dff_B_DV7KcakJ4_2),.dout(w_dff_B_5G5O4tAY5_2),.clk(gclk));
	jdff dff_B_BhBgSvci0_2(.din(w_dff_B_5G5O4tAY5_2),.dout(w_dff_B_BhBgSvci0_2),.clk(gclk));
	jdff dff_B_X2m81CUq2_2(.din(w_dff_B_BhBgSvci0_2),.dout(w_dff_B_X2m81CUq2_2),.clk(gclk));
	jdff dff_B_98JUuTyE8_2(.din(w_dff_B_X2m81CUq2_2),.dout(w_dff_B_98JUuTyE8_2),.clk(gclk));
	jdff dff_B_as2GFjCB3_2(.din(w_dff_B_98JUuTyE8_2),.dout(w_dff_B_as2GFjCB3_2),.clk(gclk));
	jdff dff_B_y5DIGxyD8_2(.din(w_dff_B_as2GFjCB3_2),.dout(w_dff_B_y5DIGxyD8_2),.clk(gclk));
	jdff dff_B_pf9LINJP3_2(.din(w_dff_B_y5DIGxyD8_2),.dout(w_dff_B_pf9LINJP3_2),.clk(gclk));
	jdff dff_B_azIu6PLv9_2(.din(w_dff_B_pf9LINJP3_2),.dout(w_dff_B_azIu6PLv9_2),.clk(gclk));
	jdff dff_B_ECf88KlO9_2(.din(w_dff_B_azIu6PLv9_2),.dout(w_dff_B_ECf88KlO9_2),.clk(gclk));
	jdff dff_B_7MgmOrwr1_2(.din(w_dff_B_ECf88KlO9_2),.dout(w_dff_B_7MgmOrwr1_2),.clk(gclk));
	jdff dff_B_mgZhSM261_2(.din(w_dff_B_7MgmOrwr1_2),.dout(w_dff_B_mgZhSM261_2),.clk(gclk));
	jdff dff_B_TlewAGHq5_2(.din(w_dff_B_mgZhSM261_2),.dout(w_dff_B_TlewAGHq5_2),.clk(gclk));
	jdff dff_B_2Nyxptkn9_2(.din(w_dff_B_TlewAGHq5_2),.dout(w_dff_B_2Nyxptkn9_2),.clk(gclk));
	jdff dff_B_l3j2iUwR7_2(.din(w_dff_B_2Nyxptkn9_2),.dout(w_dff_B_l3j2iUwR7_2),.clk(gclk));
	jdff dff_B_GlrHFx7c9_2(.din(w_dff_B_l3j2iUwR7_2),.dout(w_dff_B_GlrHFx7c9_2),.clk(gclk));
	jdff dff_B_C2xiafOV4_2(.din(w_dff_B_GlrHFx7c9_2),.dout(w_dff_B_C2xiafOV4_2),.clk(gclk));
	jdff dff_B_cCKohKyh5_2(.din(w_dff_B_C2xiafOV4_2),.dout(w_dff_B_cCKohKyh5_2),.clk(gclk));
	jdff dff_B_l8C2ByAj2_2(.din(w_dff_B_cCKohKyh5_2),.dout(w_dff_B_l8C2ByAj2_2),.clk(gclk));
	jdff dff_A_qzgPrtGO7_1(.dout(w_n1032_0[1]),.din(w_dff_A_qzgPrtGO7_1),.clk(gclk));
	jdff dff_A_BJrHJgjF4_0(.dout(w_n840_0[0]),.din(w_dff_A_BJrHJgjF4_0),.clk(gclk));
	jdff dff_A_qYJKegax7_0(.dout(w_dff_A_BJrHJgjF4_0),.din(w_dff_A_qYJKegax7_0),.clk(gclk));
	jdff dff_A_UiXGr92k1_0(.dout(w_dff_A_qYJKegax7_0),.din(w_dff_A_UiXGr92k1_0),.clk(gclk));
	jdff dff_A_W6h5kWeR9_0(.dout(w_dff_A_UiXGr92k1_0),.din(w_dff_A_W6h5kWeR9_0),.clk(gclk));
	jdff dff_A_tA04Wu2J0_0(.dout(w_dff_A_W6h5kWeR9_0),.din(w_dff_A_tA04Wu2J0_0),.clk(gclk));
	jdff dff_A_VvPFzFwC8_0(.dout(w_dff_A_tA04Wu2J0_0),.din(w_dff_A_VvPFzFwC8_0),.clk(gclk));
	jdff dff_A_KK9UUVl54_0(.dout(w_dff_A_VvPFzFwC8_0),.din(w_dff_A_KK9UUVl54_0),.clk(gclk));
	jdff dff_A_EBmNu9Oy6_0(.dout(w_dff_A_KK9UUVl54_0),.din(w_dff_A_EBmNu9Oy6_0),.clk(gclk));
	jdff dff_A_kt3X1cE19_0(.dout(w_dff_A_EBmNu9Oy6_0),.din(w_dff_A_kt3X1cE19_0),.clk(gclk));
	jdff dff_A_umJctkA12_0(.dout(w_dff_A_kt3X1cE19_0),.din(w_dff_A_umJctkA12_0),.clk(gclk));
	jdff dff_A_HHGvKxhp7_0(.dout(w_dff_A_umJctkA12_0),.din(w_dff_A_HHGvKxhp7_0),.clk(gclk));
	jdff dff_A_hDHH47Fi6_0(.dout(w_dff_A_HHGvKxhp7_0),.din(w_dff_A_hDHH47Fi6_0),.clk(gclk));
	jdff dff_A_4vgObg4A9_0(.dout(w_dff_A_hDHH47Fi6_0),.din(w_dff_A_4vgObg4A9_0),.clk(gclk));
	jdff dff_A_Rpjy6oS47_0(.dout(w_dff_A_4vgObg4A9_0),.din(w_dff_A_Rpjy6oS47_0),.clk(gclk));
	jdff dff_A_QJmZYqEV9_0(.dout(w_dff_A_Rpjy6oS47_0),.din(w_dff_A_QJmZYqEV9_0),.clk(gclk));
	jdff dff_A_fA4xHuXH3_0(.dout(w_dff_A_QJmZYqEV9_0),.din(w_dff_A_fA4xHuXH3_0),.clk(gclk));
	jdff dff_A_PLigeOWi8_0(.dout(w_dff_A_fA4xHuXH3_0),.din(w_dff_A_PLigeOWi8_0),.clk(gclk));
	jdff dff_A_RAarvpgD9_0(.dout(w_dff_A_PLigeOWi8_0),.din(w_dff_A_RAarvpgD9_0),.clk(gclk));
	jdff dff_A_UgoKJSae5_0(.dout(w_dff_A_RAarvpgD9_0),.din(w_dff_A_UgoKJSae5_0),.clk(gclk));
	jdff dff_A_NZAsxVwn0_0(.dout(w_dff_A_UgoKJSae5_0),.din(w_dff_A_NZAsxVwn0_0),.clk(gclk));
	jdff dff_A_9dF0jMfQ0_0(.dout(w_dff_A_NZAsxVwn0_0),.din(w_dff_A_9dF0jMfQ0_0),.clk(gclk));
	jdff dff_A_bWFBy0420_0(.dout(w_dff_A_9dF0jMfQ0_0),.din(w_dff_A_bWFBy0420_0),.clk(gclk));
	jdff dff_A_6JRJDj9P4_0(.dout(w_dff_A_bWFBy0420_0),.din(w_dff_A_6JRJDj9P4_0),.clk(gclk));
	jdff dff_A_vo4YJvxa3_0(.dout(w_dff_A_6JRJDj9P4_0),.din(w_dff_A_vo4YJvxa3_0),.clk(gclk));
	jdff dff_A_U6NdRyZB1_0(.dout(w_dff_A_vo4YJvxa3_0),.din(w_dff_A_U6NdRyZB1_0),.clk(gclk));
	jdff dff_A_K9vd1BE52_0(.dout(w_dff_A_U6NdRyZB1_0),.din(w_dff_A_K9vd1BE52_0),.clk(gclk));
	jdff dff_A_X26fXPwE3_0(.dout(w_dff_A_K9vd1BE52_0),.din(w_dff_A_X26fXPwE3_0),.clk(gclk));
	jdff dff_A_CO6oBVJP9_0(.dout(w_dff_A_X26fXPwE3_0),.din(w_dff_A_CO6oBVJP9_0),.clk(gclk));
	jdff dff_A_qN6gSYM48_0(.dout(w_n844_0[0]),.din(w_dff_A_qN6gSYM48_0),.clk(gclk));
	jdff dff_B_tdhjsvxw5_1(.din(n842),.dout(w_dff_B_tdhjsvxw5_1),.clk(gclk));
	jdff dff_B_QE2RFmPL0_2(.din(n742),.dout(w_dff_B_QE2RFmPL0_2),.clk(gclk));
	jdff dff_B_ZAk0Gr631_2(.din(w_dff_B_QE2RFmPL0_2),.dout(w_dff_B_ZAk0Gr631_2),.clk(gclk));
	jdff dff_B_uEqKH06t2_2(.din(w_dff_B_ZAk0Gr631_2),.dout(w_dff_B_uEqKH06t2_2),.clk(gclk));
	jdff dff_B_N5zk9FHS4_2(.din(w_dff_B_uEqKH06t2_2),.dout(w_dff_B_N5zk9FHS4_2),.clk(gclk));
	jdff dff_B_ZCwqaOg38_2(.din(w_dff_B_N5zk9FHS4_2),.dout(w_dff_B_ZCwqaOg38_2),.clk(gclk));
	jdff dff_B_A3mAc1jt2_2(.din(w_dff_B_ZCwqaOg38_2),.dout(w_dff_B_A3mAc1jt2_2),.clk(gclk));
	jdff dff_B_d7c6vFgR9_2(.din(w_dff_B_A3mAc1jt2_2),.dout(w_dff_B_d7c6vFgR9_2),.clk(gclk));
	jdff dff_B_GxW7UAtM8_2(.din(w_dff_B_d7c6vFgR9_2),.dout(w_dff_B_GxW7UAtM8_2),.clk(gclk));
	jdff dff_B_8FuUaeVB6_2(.din(w_dff_B_GxW7UAtM8_2),.dout(w_dff_B_8FuUaeVB6_2),.clk(gclk));
	jdff dff_B_3CS8Zprk9_2(.din(w_dff_B_8FuUaeVB6_2),.dout(w_dff_B_3CS8Zprk9_2),.clk(gclk));
	jdff dff_B_gtBI0k7n7_2(.din(w_dff_B_3CS8Zprk9_2),.dout(w_dff_B_gtBI0k7n7_2),.clk(gclk));
	jdff dff_B_04q9SLLh6_2(.din(w_dff_B_gtBI0k7n7_2),.dout(w_dff_B_04q9SLLh6_2),.clk(gclk));
	jdff dff_B_IXcYr1ok6_2(.din(w_dff_B_04q9SLLh6_2),.dout(w_dff_B_IXcYr1ok6_2),.clk(gclk));
	jdff dff_B_d3M1XEIT8_2(.din(w_dff_B_IXcYr1ok6_2),.dout(w_dff_B_d3M1XEIT8_2),.clk(gclk));
	jdff dff_B_qSNgsTXK3_2(.din(w_dff_B_d3M1XEIT8_2),.dout(w_dff_B_qSNgsTXK3_2),.clk(gclk));
	jdff dff_B_K033VI0H4_2(.din(w_dff_B_qSNgsTXK3_2),.dout(w_dff_B_K033VI0H4_2),.clk(gclk));
	jdff dff_B_NAH9VlkF0_2(.din(w_dff_B_K033VI0H4_2),.dout(w_dff_B_NAH9VlkF0_2),.clk(gclk));
	jdff dff_B_FAgdJ6M35_2(.din(w_dff_B_NAH9VlkF0_2),.dout(w_dff_B_FAgdJ6M35_2),.clk(gclk));
	jdff dff_B_F7kkwPo64_2(.din(w_dff_B_FAgdJ6M35_2),.dout(w_dff_B_F7kkwPo64_2),.clk(gclk));
	jdff dff_B_DGOdcGys8_2(.din(w_dff_B_F7kkwPo64_2),.dout(w_dff_B_DGOdcGys8_2),.clk(gclk));
	jdff dff_B_qbpJxz6L6_2(.din(w_dff_B_DGOdcGys8_2),.dout(w_dff_B_qbpJxz6L6_2),.clk(gclk));
	jdff dff_B_wvIK4g903_2(.din(w_dff_B_qbpJxz6L6_2),.dout(w_dff_B_wvIK4g903_2),.clk(gclk));
	jdff dff_B_jQ25XXm10_2(.din(w_dff_B_wvIK4g903_2),.dout(w_dff_B_jQ25XXm10_2),.clk(gclk));
	jdff dff_B_6zgCuI5N9_2(.din(w_dff_B_jQ25XXm10_2),.dout(w_dff_B_6zgCuI5N9_2),.clk(gclk));
	jdff dff_B_0jnZfbuD4_1(.din(n743),.dout(w_dff_B_0jnZfbuD4_1),.clk(gclk));
	jdff dff_B_d6JRT1Sj6_2(.din(n649),.dout(w_dff_B_d6JRT1Sj6_2),.clk(gclk));
	jdff dff_B_F4eMiP946_2(.din(w_dff_B_d6JRT1Sj6_2),.dout(w_dff_B_F4eMiP946_2),.clk(gclk));
	jdff dff_B_7beeHpPI5_2(.din(w_dff_B_F4eMiP946_2),.dout(w_dff_B_7beeHpPI5_2),.clk(gclk));
	jdff dff_B_4RIWZMKQ9_2(.din(w_dff_B_7beeHpPI5_2),.dout(w_dff_B_4RIWZMKQ9_2),.clk(gclk));
	jdff dff_B_3VcQRmN99_2(.din(w_dff_B_4RIWZMKQ9_2),.dout(w_dff_B_3VcQRmN99_2),.clk(gclk));
	jdff dff_B_lJZefGct7_2(.din(w_dff_B_3VcQRmN99_2),.dout(w_dff_B_lJZefGct7_2),.clk(gclk));
	jdff dff_B_toChjdRD8_2(.din(w_dff_B_lJZefGct7_2),.dout(w_dff_B_toChjdRD8_2),.clk(gclk));
	jdff dff_B_ORPnprfv7_2(.din(w_dff_B_toChjdRD8_2),.dout(w_dff_B_ORPnprfv7_2),.clk(gclk));
	jdff dff_B_r3bPQwLu6_2(.din(w_dff_B_ORPnprfv7_2),.dout(w_dff_B_r3bPQwLu6_2),.clk(gclk));
	jdff dff_B_DHfGuWza7_2(.din(w_dff_B_r3bPQwLu6_2),.dout(w_dff_B_DHfGuWza7_2),.clk(gclk));
	jdff dff_B_kHAppI2U9_2(.din(w_dff_B_DHfGuWza7_2),.dout(w_dff_B_kHAppI2U9_2),.clk(gclk));
	jdff dff_B_W8PLt7xB4_2(.din(w_dff_B_kHAppI2U9_2),.dout(w_dff_B_W8PLt7xB4_2),.clk(gclk));
	jdff dff_B_HNc09p799_2(.din(w_dff_B_W8PLt7xB4_2),.dout(w_dff_B_HNc09p799_2),.clk(gclk));
	jdff dff_B_ZiISFO4e6_2(.din(w_dff_B_HNc09p799_2),.dout(w_dff_B_ZiISFO4e6_2),.clk(gclk));
	jdff dff_B_IMh2db9w0_2(.din(w_dff_B_ZiISFO4e6_2),.dout(w_dff_B_IMh2db9w0_2),.clk(gclk));
	jdff dff_B_nNO7I5rT4_2(.din(w_dff_B_IMh2db9w0_2),.dout(w_dff_B_nNO7I5rT4_2),.clk(gclk));
	jdff dff_B_vAFM8nZu5_2(.din(w_dff_B_nNO7I5rT4_2),.dout(w_dff_B_vAFM8nZu5_2),.clk(gclk));
	jdff dff_B_r8pVk9yJ3_2(.din(w_dff_B_vAFM8nZu5_2),.dout(w_dff_B_r8pVk9yJ3_2),.clk(gclk));
	jdff dff_B_TIh27FCV9_2(.din(w_dff_B_r8pVk9yJ3_2),.dout(w_dff_B_TIh27FCV9_2),.clk(gclk));
	jdff dff_B_9guNURWa8_2(.din(w_dff_B_TIh27FCV9_2),.dout(w_dff_B_9guNURWa8_2),.clk(gclk));
	jdff dff_B_Gai22cUS9_2(.din(w_dff_B_9guNURWa8_2),.dout(w_dff_B_Gai22cUS9_2),.clk(gclk));
	jdff dff_B_dD5wDP8N1_2(.din(w_dff_B_Gai22cUS9_2),.dout(w_dff_B_dD5wDP8N1_2),.clk(gclk));
	jdff dff_B_Wmw0vaVP3_1(.din(n650),.dout(w_dff_B_Wmw0vaVP3_1),.clk(gclk));
	jdff dff_B_E6csAyxh8_2(.din(n563),.dout(w_dff_B_E6csAyxh8_2),.clk(gclk));
	jdff dff_B_PEBJSwCH4_2(.din(w_dff_B_E6csAyxh8_2),.dout(w_dff_B_PEBJSwCH4_2),.clk(gclk));
	jdff dff_B_nJ6zdzMn2_2(.din(w_dff_B_PEBJSwCH4_2),.dout(w_dff_B_nJ6zdzMn2_2),.clk(gclk));
	jdff dff_B_fGI7bQZ27_2(.din(w_dff_B_nJ6zdzMn2_2),.dout(w_dff_B_fGI7bQZ27_2),.clk(gclk));
	jdff dff_B_Ul4N78Sf0_2(.din(w_dff_B_fGI7bQZ27_2),.dout(w_dff_B_Ul4N78Sf0_2),.clk(gclk));
	jdff dff_B_o3rwXkbv3_2(.din(w_dff_B_Ul4N78Sf0_2),.dout(w_dff_B_o3rwXkbv3_2),.clk(gclk));
	jdff dff_B_itXsQoc02_2(.din(w_dff_B_o3rwXkbv3_2),.dout(w_dff_B_itXsQoc02_2),.clk(gclk));
	jdff dff_B_WVbB8UgY6_2(.din(w_dff_B_itXsQoc02_2),.dout(w_dff_B_WVbB8UgY6_2),.clk(gclk));
	jdff dff_B_0GVjnti59_2(.din(w_dff_B_WVbB8UgY6_2),.dout(w_dff_B_0GVjnti59_2),.clk(gclk));
	jdff dff_B_uk17SVWN7_2(.din(w_dff_B_0GVjnti59_2),.dout(w_dff_B_uk17SVWN7_2),.clk(gclk));
	jdff dff_B_s9CxG9Br1_2(.din(w_dff_B_uk17SVWN7_2),.dout(w_dff_B_s9CxG9Br1_2),.clk(gclk));
	jdff dff_B_gHJ0ImCt1_2(.din(w_dff_B_s9CxG9Br1_2),.dout(w_dff_B_gHJ0ImCt1_2),.clk(gclk));
	jdff dff_B_Ot0FYI356_2(.din(w_dff_B_gHJ0ImCt1_2),.dout(w_dff_B_Ot0FYI356_2),.clk(gclk));
	jdff dff_B_xAZXpZzQ1_2(.din(w_dff_B_Ot0FYI356_2),.dout(w_dff_B_xAZXpZzQ1_2),.clk(gclk));
	jdff dff_B_N3Gsflrv8_2(.din(w_dff_B_xAZXpZzQ1_2),.dout(w_dff_B_N3Gsflrv8_2),.clk(gclk));
	jdff dff_B_ZcQzw2tB0_2(.din(w_dff_B_N3Gsflrv8_2),.dout(w_dff_B_ZcQzw2tB0_2),.clk(gclk));
	jdff dff_B_um5QauEF7_2(.din(w_dff_B_ZcQzw2tB0_2),.dout(w_dff_B_um5QauEF7_2),.clk(gclk));
	jdff dff_B_plqHSaSK6_2(.din(w_dff_B_um5QauEF7_2),.dout(w_dff_B_plqHSaSK6_2),.clk(gclk));
	jdff dff_B_IYScNTsq6_2(.din(w_dff_B_plqHSaSK6_2),.dout(w_dff_B_IYScNTsq6_2),.clk(gclk));
	jdff dff_B_v4zCLJrf9_2(.din(w_dff_B_IYScNTsq6_2),.dout(w_dff_B_v4zCLJrf9_2),.clk(gclk));
	jdff dff_B_mNrhr0kP7_1(.din(n564),.dout(w_dff_B_mNrhr0kP7_1),.clk(gclk));
	jdff dff_B_8uU0orkr0_2(.din(n484),.dout(w_dff_B_8uU0orkr0_2),.clk(gclk));
	jdff dff_B_xdTh0JsV9_2(.din(w_dff_B_8uU0orkr0_2),.dout(w_dff_B_xdTh0JsV9_2),.clk(gclk));
	jdff dff_B_ZCY2u8bj9_2(.din(w_dff_B_xdTh0JsV9_2),.dout(w_dff_B_ZCY2u8bj9_2),.clk(gclk));
	jdff dff_B_uQiFdHlv7_2(.din(w_dff_B_ZCY2u8bj9_2),.dout(w_dff_B_uQiFdHlv7_2),.clk(gclk));
	jdff dff_B_fGTMR4Om5_2(.din(w_dff_B_uQiFdHlv7_2),.dout(w_dff_B_fGTMR4Om5_2),.clk(gclk));
	jdff dff_B_ZolFk9wV5_2(.din(w_dff_B_fGTMR4Om5_2),.dout(w_dff_B_ZolFk9wV5_2),.clk(gclk));
	jdff dff_B_uMHjTHCD7_2(.din(w_dff_B_ZolFk9wV5_2),.dout(w_dff_B_uMHjTHCD7_2),.clk(gclk));
	jdff dff_B_lSRmAsPP8_2(.din(w_dff_B_uMHjTHCD7_2),.dout(w_dff_B_lSRmAsPP8_2),.clk(gclk));
	jdff dff_B_aSolrUlR4_2(.din(w_dff_B_lSRmAsPP8_2),.dout(w_dff_B_aSolrUlR4_2),.clk(gclk));
	jdff dff_B_sLtem57U4_2(.din(w_dff_B_aSolrUlR4_2),.dout(w_dff_B_sLtem57U4_2),.clk(gclk));
	jdff dff_B_h2M5yWJp4_2(.din(w_dff_B_sLtem57U4_2),.dout(w_dff_B_h2M5yWJp4_2),.clk(gclk));
	jdff dff_B_3XP1Phog8_2(.din(w_dff_B_h2M5yWJp4_2),.dout(w_dff_B_3XP1Phog8_2),.clk(gclk));
	jdff dff_B_IPSYJc9R2_2(.din(w_dff_B_3XP1Phog8_2),.dout(w_dff_B_IPSYJc9R2_2),.clk(gclk));
	jdff dff_B_Hn9nAkO59_2(.din(w_dff_B_IPSYJc9R2_2),.dout(w_dff_B_Hn9nAkO59_2),.clk(gclk));
	jdff dff_B_423A2rfK5_2(.din(w_dff_B_Hn9nAkO59_2),.dout(w_dff_B_423A2rfK5_2),.clk(gclk));
	jdff dff_B_XdpRRCVC1_2(.din(w_dff_B_423A2rfK5_2),.dout(w_dff_B_XdpRRCVC1_2),.clk(gclk));
	jdff dff_B_xZRDx6Bt5_2(.din(w_dff_B_XdpRRCVC1_2),.dout(w_dff_B_xZRDx6Bt5_2),.clk(gclk));
	jdff dff_B_2aqVfDn05_2(.din(w_dff_B_xZRDx6Bt5_2),.dout(w_dff_B_2aqVfDn05_2),.clk(gclk));
	jdff dff_B_qGJNeFyw7_1(.din(n485),.dout(w_dff_B_qGJNeFyw7_1),.clk(gclk));
	jdff dff_B_kwKlTODZ5_2(.din(n412),.dout(w_dff_B_kwKlTODZ5_2),.clk(gclk));
	jdff dff_B_SwkXeJ1I6_2(.din(w_dff_B_kwKlTODZ5_2),.dout(w_dff_B_SwkXeJ1I6_2),.clk(gclk));
	jdff dff_B_m4SnrpPw0_2(.din(w_dff_B_SwkXeJ1I6_2),.dout(w_dff_B_m4SnrpPw0_2),.clk(gclk));
	jdff dff_B_AL2yACLO7_2(.din(w_dff_B_m4SnrpPw0_2),.dout(w_dff_B_AL2yACLO7_2),.clk(gclk));
	jdff dff_B_o732N5oX6_2(.din(w_dff_B_AL2yACLO7_2),.dout(w_dff_B_o732N5oX6_2),.clk(gclk));
	jdff dff_B_1rvJfPSJ5_2(.din(w_dff_B_o732N5oX6_2),.dout(w_dff_B_1rvJfPSJ5_2),.clk(gclk));
	jdff dff_B_ikLtOuxI9_2(.din(w_dff_B_1rvJfPSJ5_2),.dout(w_dff_B_ikLtOuxI9_2),.clk(gclk));
	jdff dff_B_ylp4eRFb0_2(.din(w_dff_B_ikLtOuxI9_2),.dout(w_dff_B_ylp4eRFb0_2),.clk(gclk));
	jdff dff_B_r0DdNQZO0_2(.din(w_dff_B_ylp4eRFb0_2),.dout(w_dff_B_r0DdNQZO0_2),.clk(gclk));
	jdff dff_B_x00hC7cC4_2(.din(w_dff_B_r0DdNQZO0_2),.dout(w_dff_B_x00hC7cC4_2),.clk(gclk));
	jdff dff_B_CaJO27J65_2(.din(w_dff_B_x00hC7cC4_2),.dout(w_dff_B_CaJO27J65_2),.clk(gclk));
	jdff dff_B_x11CjgDl4_2(.din(w_dff_B_CaJO27J65_2),.dout(w_dff_B_x11CjgDl4_2),.clk(gclk));
	jdff dff_B_zeoYnGYG9_2(.din(w_dff_B_x11CjgDl4_2),.dout(w_dff_B_zeoYnGYG9_2),.clk(gclk));
	jdff dff_B_bvwz06ZQ6_2(.din(w_dff_B_zeoYnGYG9_2),.dout(w_dff_B_bvwz06ZQ6_2),.clk(gclk));
	jdff dff_B_XYEyF6it7_2(.din(w_dff_B_bvwz06ZQ6_2),.dout(w_dff_B_XYEyF6it7_2),.clk(gclk));
	jdff dff_B_TL6QGUTC1_2(.din(w_dff_B_XYEyF6it7_2),.dout(w_dff_B_TL6QGUTC1_2),.clk(gclk));
	jdff dff_B_O4itNlQT3_1(.din(n413),.dout(w_dff_B_O4itNlQT3_1),.clk(gclk));
	jdff dff_B_SR5M0VzB2_2(.din(n348),.dout(w_dff_B_SR5M0VzB2_2),.clk(gclk));
	jdff dff_B_XWv2B1TI7_2(.din(w_dff_B_SR5M0VzB2_2),.dout(w_dff_B_XWv2B1TI7_2),.clk(gclk));
	jdff dff_B_H2hSsFwG9_2(.din(w_dff_B_XWv2B1TI7_2),.dout(w_dff_B_H2hSsFwG9_2),.clk(gclk));
	jdff dff_B_UukRbFo74_2(.din(w_dff_B_H2hSsFwG9_2),.dout(w_dff_B_UukRbFo74_2),.clk(gclk));
	jdff dff_B_ONDBlnSX9_2(.din(w_dff_B_UukRbFo74_2),.dout(w_dff_B_ONDBlnSX9_2),.clk(gclk));
	jdff dff_B_J3HNgRAf3_2(.din(w_dff_B_ONDBlnSX9_2),.dout(w_dff_B_J3HNgRAf3_2),.clk(gclk));
	jdff dff_B_CzZuSfpC0_2(.din(w_dff_B_J3HNgRAf3_2),.dout(w_dff_B_CzZuSfpC0_2),.clk(gclk));
	jdff dff_B_8EGuyn8o5_2(.din(w_dff_B_CzZuSfpC0_2),.dout(w_dff_B_8EGuyn8o5_2),.clk(gclk));
	jdff dff_B_Ok4Ld4ha5_2(.din(w_dff_B_8EGuyn8o5_2),.dout(w_dff_B_Ok4Ld4ha5_2),.clk(gclk));
	jdff dff_B_uE7FpfDF3_2(.din(w_dff_B_Ok4Ld4ha5_2),.dout(w_dff_B_uE7FpfDF3_2),.clk(gclk));
	jdff dff_B_g7vvmbgS7_2(.din(w_dff_B_uE7FpfDF3_2),.dout(w_dff_B_g7vvmbgS7_2),.clk(gclk));
	jdff dff_B_6UAniggy6_2(.din(w_dff_B_g7vvmbgS7_2),.dout(w_dff_B_6UAniggy6_2),.clk(gclk));
	jdff dff_B_GyVhD9yX8_2(.din(w_dff_B_6UAniggy6_2),.dout(w_dff_B_GyVhD9yX8_2),.clk(gclk));
	jdff dff_B_P7GxG97t3_2(.din(w_dff_B_GyVhD9yX8_2),.dout(w_dff_B_P7GxG97t3_2),.clk(gclk));
	jdff dff_B_mxWU2CBS8_1(.din(n349),.dout(w_dff_B_mxWU2CBS8_1),.clk(gclk));
	jdff dff_B_Zm67YdwU8_2(.din(n290),.dout(w_dff_B_Zm67YdwU8_2),.clk(gclk));
	jdff dff_B_g1MQVclp4_2(.din(w_dff_B_Zm67YdwU8_2),.dout(w_dff_B_g1MQVclp4_2),.clk(gclk));
	jdff dff_B_Sv2u7VZ55_2(.din(w_dff_B_g1MQVclp4_2),.dout(w_dff_B_Sv2u7VZ55_2),.clk(gclk));
	jdff dff_B_oUyA7ZVi8_2(.din(w_dff_B_Sv2u7VZ55_2),.dout(w_dff_B_oUyA7ZVi8_2),.clk(gclk));
	jdff dff_B_yF7lTfJJ9_2(.din(w_dff_B_oUyA7ZVi8_2),.dout(w_dff_B_yF7lTfJJ9_2),.clk(gclk));
	jdff dff_B_n5xq0kya3_2(.din(w_dff_B_yF7lTfJJ9_2),.dout(w_dff_B_n5xq0kya3_2),.clk(gclk));
	jdff dff_B_lTcFdM6T7_2(.din(w_dff_B_n5xq0kya3_2),.dout(w_dff_B_lTcFdM6T7_2),.clk(gclk));
	jdff dff_B_y9ZTsqQz0_2(.din(w_dff_B_lTcFdM6T7_2),.dout(w_dff_B_y9ZTsqQz0_2),.clk(gclk));
	jdff dff_B_sHZYPjDW3_2(.din(w_dff_B_y9ZTsqQz0_2),.dout(w_dff_B_sHZYPjDW3_2),.clk(gclk));
	jdff dff_B_QNXXIVyt4_2(.din(w_dff_B_sHZYPjDW3_2),.dout(w_dff_B_QNXXIVyt4_2),.clk(gclk));
	jdff dff_B_IAWsEFu13_2(.din(w_dff_B_QNXXIVyt4_2),.dout(w_dff_B_IAWsEFu13_2),.clk(gclk));
	jdff dff_B_669JR3NH1_2(.din(w_dff_B_IAWsEFu13_2),.dout(w_dff_B_669JR3NH1_2),.clk(gclk));
	jdff dff_B_Dk6URZcJ7_1(.din(n291),.dout(w_dff_B_Dk6URZcJ7_1),.clk(gclk));
	jdff dff_B_3Atefzp26_2(.din(n239),.dout(w_dff_B_3Atefzp26_2),.clk(gclk));
	jdff dff_B_Fufmaz4c0_2(.din(w_dff_B_3Atefzp26_2),.dout(w_dff_B_Fufmaz4c0_2),.clk(gclk));
	jdff dff_B_6NCIYT4J2_2(.din(w_dff_B_Fufmaz4c0_2),.dout(w_dff_B_6NCIYT4J2_2),.clk(gclk));
	jdff dff_B_0UlYdXqn4_2(.din(w_dff_B_6NCIYT4J2_2),.dout(w_dff_B_0UlYdXqn4_2),.clk(gclk));
	jdff dff_B_Ppt82TVn7_2(.din(w_dff_B_0UlYdXqn4_2),.dout(w_dff_B_Ppt82TVn7_2),.clk(gclk));
	jdff dff_B_5rQPrQYp5_2(.din(w_dff_B_Ppt82TVn7_2),.dout(w_dff_B_5rQPrQYp5_2),.clk(gclk));
	jdff dff_B_NcTAceBg3_2(.din(w_dff_B_5rQPrQYp5_2),.dout(w_dff_B_NcTAceBg3_2),.clk(gclk));
	jdff dff_B_juyQzPl45_2(.din(w_dff_B_NcTAceBg3_2),.dout(w_dff_B_juyQzPl45_2),.clk(gclk));
	jdff dff_B_EknasaLQ9_2(.din(w_dff_B_juyQzPl45_2),.dout(w_dff_B_EknasaLQ9_2),.clk(gclk));
	jdff dff_B_o5szB85e1_2(.din(w_dff_B_EknasaLQ9_2),.dout(w_dff_B_o5szB85e1_2),.clk(gclk));
	jdff dff_B_bSS4JKmy4_1(.din(n240),.dout(w_dff_B_bSS4JKmy4_1),.clk(gclk));
	jdff dff_B_RGFVFglE4_2(.din(n196),.dout(w_dff_B_RGFVFglE4_2),.clk(gclk));
	jdff dff_B_55E2HOtn8_2(.din(w_dff_B_RGFVFglE4_2),.dout(w_dff_B_55E2HOtn8_2),.clk(gclk));
	jdff dff_B_KnVzLke91_2(.din(w_dff_B_55E2HOtn8_2),.dout(w_dff_B_KnVzLke91_2),.clk(gclk));
	jdff dff_B_IABejzyF6_2(.din(w_dff_B_KnVzLke91_2),.dout(w_dff_B_IABejzyF6_2),.clk(gclk));
	jdff dff_B_SxkHWhwO0_2(.din(w_dff_B_IABejzyF6_2),.dout(w_dff_B_SxkHWhwO0_2),.clk(gclk));
	jdff dff_B_ZFW7P50Q9_2(.din(w_dff_B_SxkHWhwO0_2),.dout(w_dff_B_ZFW7P50Q9_2),.clk(gclk));
	jdff dff_B_zV0An42L0_2(.din(w_dff_B_ZFW7P50Q9_2),.dout(w_dff_B_zV0An42L0_2),.clk(gclk));
	jdff dff_B_0YPYM2yI9_2(.din(w_dff_B_zV0An42L0_2),.dout(w_dff_B_0YPYM2yI9_2),.clk(gclk));
	jdff dff_B_KV0W7Hdu4_2(.din(n218),.dout(w_dff_B_KV0W7Hdu4_2),.clk(gclk));
	jdff dff_B_SxyvgrUB3_1(.din(n197),.dout(w_dff_B_SxyvgrUB3_1),.clk(gclk));
	jdff dff_B_0tChY7Uu8_2(.din(n158),.dout(w_dff_B_0tChY7Uu8_2),.clk(gclk));
	jdff dff_B_oYHn7muD7_2(.din(w_dff_B_0tChY7Uu8_2),.dout(w_dff_B_oYHn7muD7_2),.clk(gclk));
	jdff dff_B_ehy3hBab9_2(.din(w_dff_B_oYHn7muD7_2),.dout(w_dff_B_ehy3hBab9_2),.clk(gclk));
	jdff dff_B_ielkX7kY1_2(.din(w_dff_B_ehy3hBab9_2),.dout(w_dff_B_ielkX7kY1_2),.clk(gclk));
	jdff dff_B_DwabZDaX7_2(.din(w_dff_B_ielkX7kY1_2),.dout(w_dff_B_DwabZDaX7_2),.clk(gclk));
	jdff dff_B_d3eFCLjg4_2(.din(w_dff_B_DwabZDaX7_2),.dout(w_dff_B_d3eFCLjg4_2),.clk(gclk));
	jdff dff_B_r8aFdsh71_2(.din(n175),.dout(w_dff_B_r8aFdsh71_2),.clk(gclk));
	jdff dff_B_xm84fC9V6_1(.din(n161),.dout(w_dff_B_xm84fC9V6_1),.clk(gclk));
	jdff dff_B_IADcx8xB8_1(.din(w_dff_B_xm84fC9V6_1),.dout(w_dff_B_IADcx8xB8_1),.clk(gclk));
	jdff dff_B_ZW6ADBYo1_1(.din(w_dff_B_IADcx8xB8_1),.dout(w_dff_B_ZW6ADBYo1_1),.clk(gclk));
	jdff dff_B_BztZO27i2_1(.din(n135),.dout(w_dff_B_BztZO27i2_1),.clk(gclk));
	jdff dff_B_QzidDl7h9_2(.din(n128),.dout(w_dff_B_QzidDl7h9_2),.clk(gclk));
	jdff dff_B_QXdIKbgG8_2(.din(w_dff_B_QzidDl7h9_2),.dout(w_dff_B_QXdIKbgG8_2),.clk(gclk));
	jdff dff_B_CZm2vIc71_2(.din(w_dff_B_QXdIKbgG8_2),.dout(w_dff_B_CZm2vIc71_2),.clk(gclk));
	jdff dff_B_DMlKtyFT9_2(.din(w_dff_B_CZm2vIc71_2),.dout(w_dff_B_DMlKtyFT9_2),.clk(gclk));
	jdff dff_B_VuZ7sJNf6_0(.din(n160),.dout(w_dff_B_VuZ7sJNf6_0),.clk(gclk));
	jdff dff_A_MOenS5Y47_1(.dout(w_n130_0[1]),.din(w_dff_A_MOenS5Y47_1),.clk(gclk));
	jdff dff_A_RCAO2G978_1(.dout(w_dff_A_MOenS5Y47_1),.din(w_dff_A_RCAO2G978_1),.clk(gclk));
	jdff dff_A_RUhPeT7s8_1(.dout(w_n100_0[1]),.din(w_dff_A_RUhPeT7s8_1),.clk(gclk));
	jdff dff_A_Zns8hL4f9_2(.dout(w_n100_0[2]),.din(w_dff_A_Zns8hL4f9_2),.clk(gclk));
	jdff dff_A_7OiKETeF1_2(.dout(w_dff_A_Zns8hL4f9_2),.din(w_dff_A_7OiKETeF1_2),.clk(gclk));
	jdff dff_A_2DXqsfki9_0(.dout(w_n1247_0[0]),.din(w_dff_A_2DXqsfki9_0),.clk(gclk));
	jdff dff_B_4bprLLu56_1(.din(n1245),.dout(w_dff_B_4bprLLu56_1),.clk(gclk));
	jdff dff_B_HQ0398zs6_1(.din(w_dff_B_4bprLLu56_1),.dout(w_dff_B_HQ0398zs6_1),.clk(gclk));
	jdff dff_B_rVfDrSbl7_2(.din(n1152),.dout(w_dff_B_rVfDrSbl7_2),.clk(gclk));
	jdff dff_B_OUR5TpkR0_2(.din(w_dff_B_rVfDrSbl7_2),.dout(w_dff_B_OUR5TpkR0_2),.clk(gclk));
	jdff dff_B_eh1kDnH91_2(.din(w_dff_B_OUR5TpkR0_2),.dout(w_dff_B_eh1kDnH91_2),.clk(gclk));
	jdff dff_B_0pIJejLK6_2(.din(w_dff_B_eh1kDnH91_2),.dout(w_dff_B_0pIJejLK6_2),.clk(gclk));
	jdff dff_B_fVgrTWcy5_2(.din(w_dff_B_0pIJejLK6_2),.dout(w_dff_B_fVgrTWcy5_2),.clk(gclk));
	jdff dff_B_0d7leuKp4_2(.din(w_dff_B_fVgrTWcy5_2),.dout(w_dff_B_0d7leuKp4_2),.clk(gclk));
	jdff dff_B_DZN7eg5X7_2(.din(w_dff_B_0d7leuKp4_2),.dout(w_dff_B_DZN7eg5X7_2),.clk(gclk));
	jdff dff_B_im3r9vEP1_2(.din(w_dff_B_DZN7eg5X7_2),.dout(w_dff_B_im3r9vEP1_2),.clk(gclk));
	jdff dff_B_shpohSec9_2(.din(w_dff_B_im3r9vEP1_2),.dout(w_dff_B_shpohSec9_2),.clk(gclk));
	jdff dff_B_z4qg006d6_2(.din(w_dff_B_shpohSec9_2),.dout(w_dff_B_z4qg006d6_2),.clk(gclk));
	jdff dff_B_yi5zyAAe4_2(.din(w_dff_B_z4qg006d6_2),.dout(w_dff_B_yi5zyAAe4_2),.clk(gclk));
	jdff dff_B_OcxFxGup5_2(.din(w_dff_B_yi5zyAAe4_2),.dout(w_dff_B_OcxFxGup5_2),.clk(gclk));
	jdff dff_B_0yLlVIZG8_2(.din(w_dff_B_OcxFxGup5_2),.dout(w_dff_B_0yLlVIZG8_2),.clk(gclk));
	jdff dff_B_g7k0XUje4_2(.din(w_dff_B_0yLlVIZG8_2),.dout(w_dff_B_g7k0XUje4_2),.clk(gclk));
	jdff dff_B_GV4HnXOn4_2(.din(w_dff_B_g7k0XUje4_2),.dout(w_dff_B_GV4HnXOn4_2),.clk(gclk));
	jdff dff_B_0j2KN2Z04_2(.din(w_dff_B_GV4HnXOn4_2),.dout(w_dff_B_0j2KN2Z04_2),.clk(gclk));
	jdff dff_B_g9qiRDzU0_2(.din(w_dff_B_0j2KN2Z04_2),.dout(w_dff_B_g9qiRDzU0_2),.clk(gclk));
	jdff dff_B_WaM41Jar5_2(.din(w_dff_B_g9qiRDzU0_2),.dout(w_dff_B_WaM41Jar5_2),.clk(gclk));
	jdff dff_B_2nsL2mIH6_2(.din(w_dff_B_WaM41Jar5_2),.dout(w_dff_B_2nsL2mIH6_2),.clk(gclk));
	jdff dff_B_EI9rOSKt0_2(.din(w_dff_B_2nsL2mIH6_2),.dout(w_dff_B_EI9rOSKt0_2),.clk(gclk));
	jdff dff_B_IQ69olqx0_2(.din(w_dff_B_EI9rOSKt0_2),.dout(w_dff_B_IQ69olqx0_2),.clk(gclk));
	jdff dff_B_1kY86yeo3_2(.din(w_dff_B_IQ69olqx0_2),.dout(w_dff_B_1kY86yeo3_2),.clk(gclk));
	jdff dff_B_OfwxjwD78_2(.din(w_dff_B_1kY86yeo3_2),.dout(w_dff_B_OfwxjwD78_2),.clk(gclk));
	jdff dff_B_31ez3Xxf3_2(.din(w_dff_B_OfwxjwD78_2),.dout(w_dff_B_31ez3Xxf3_2),.clk(gclk));
	jdff dff_B_OnzbbnUu9_2(.din(w_dff_B_31ez3Xxf3_2),.dout(w_dff_B_OnzbbnUu9_2),.clk(gclk));
	jdff dff_B_d3DbEaqy9_2(.din(w_dff_B_OnzbbnUu9_2),.dout(w_dff_B_d3DbEaqy9_2),.clk(gclk));
	jdff dff_B_z20hfsCO1_2(.din(w_dff_B_d3DbEaqy9_2),.dout(w_dff_B_z20hfsCO1_2),.clk(gclk));
	jdff dff_B_ZcSaZECM3_2(.din(w_dff_B_z20hfsCO1_2),.dout(w_dff_B_ZcSaZECM3_2),.clk(gclk));
	jdff dff_B_95Dk3xZG3_2(.din(w_dff_B_ZcSaZECM3_2),.dout(w_dff_B_95Dk3xZG3_2),.clk(gclk));
	jdff dff_B_5QIVyAeT4_2(.din(w_dff_B_95Dk3xZG3_2),.dout(w_dff_B_5QIVyAeT4_2),.clk(gclk));
	jdff dff_B_LszWiyAZ9_2(.din(w_dff_B_5QIVyAeT4_2),.dout(w_dff_B_LszWiyAZ9_2),.clk(gclk));
	jdff dff_B_l43tMi885_2(.din(w_dff_B_LszWiyAZ9_2),.dout(w_dff_B_l43tMi885_2),.clk(gclk));
	jdff dff_B_qxcq6ioB7_2(.din(w_dff_B_l43tMi885_2),.dout(w_dff_B_qxcq6ioB7_2),.clk(gclk));
	jdff dff_B_UIK0X4Nc0_2(.din(w_dff_B_qxcq6ioB7_2),.dout(w_dff_B_UIK0X4Nc0_2),.clk(gclk));
	jdff dff_B_dkaftnOp3_2(.din(w_dff_B_UIK0X4Nc0_2),.dout(w_dff_B_dkaftnOp3_2),.clk(gclk));
	jdff dff_B_HDeeE3zj8_2(.din(n1156),.dout(w_dff_B_HDeeE3zj8_2),.clk(gclk));
	jdff dff_B_ut7Gdpue6_2(.din(n1049),.dout(w_dff_B_ut7Gdpue6_2),.clk(gclk));
	jdff dff_B_8ML7WXKy8_2(.din(w_dff_B_ut7Gdpue6_2),.dout(w_dff_B_8ML7WXKy8_2),.clk(gclk));
	jdff dff_B_wVJrfpMj4_2(.din(w_dff_B_8ML7WXKy8_2),.dout(w_dff_B_wVJrfpMj4_2),.clk(gclk));
	jdff dff_B_rO9EYn8N0_2(.din(w_dff_B_wVJrfpMj4_2),.dout(w_dff_B_rO9EYn8N0_2),.clk(gclk));
	jdff dff_B_UbLV6dIC8_2(.din(w_dff_B_rO9EYn8N0_2),.dout(w_dff_B_UbLV6dIC8_2),.clk(gclk));
	jdff dff_B_SjX8Pkym2_2(.din(w_dff_B_UbLV6dIC8_2),.dout(w_dff_B_SjX8Pkym2_2),.clk(gclk));
	jdff dff_B_y31zMqjC0_2(.din(w_dff_B_SjX8Pkym2_2),.dout(w_dff_B_y31zMqjC0_2),.clk(gclk));
	jdff dff_B_DEeYucqF6_2(.din(w_dff_B_y31zMqjC0_2),.dout(w_dff_B_DEeYucqF6_2),.clk(gclk));
	jdff dff_B_VICmKp3s8_2(.din(w_dff_B_DEeYucqF6_2),.dout(w_dff_B_VICmKp3s8_2),.clk(gclk));
	jdff dff_B_zj6j3PJl0_2(.din(w_dff_B_VICmKp3s8_2),.dout(w_dff_B_zj6j3PJl0_2),.clk(gclk));
	jdff dff_B_lPOY5AIU6_2(.din(w_dff_B_zj6j3PJl0_2),.dout(w_dff_B_lPOY5AIU6_2),.clk(gclk));
	jdff dff_B_iulyastL8_2(.din(w_dff_B_lPOY5AIU6_2),.dout(w_dff_B_iulyastL8_2),.clk(gclk));
	jdff dff_B_t9fdieQX9_2(.din(w_dff_B_iulyastL8_2),.dout(w_dff_B_t9fdieQX9_2),.clk(gclk));
	jdff dff_B_9UQMQQje6_2(.din(w_dff_B_t9fdieQX9_2),.dout(w_dff_B_9UQMQQje6_2),.clk(gclk));
	jdff dff_B_4HGfjpRm0_2(.din(w_dff_B_9UQMQQje6_2),.dout(w_dff_B_4HGfjpRm0_2),.clk(gclk));
	jdff dff_B_FnRakgzV5_2(.din(w_dff_B_4HGfjpRm0_2),.dout(w_dff_B_FnRakgzV5_2),.clk(gclk));
	jdff dff_B_TtRhlFxB1_2(.din(w_dff_B_FnRakgzV5_2),.dout(w_dff_B_TtRhlFxB1_2),.clk(gclk));
	jdff dff_B_a8ULsxYn6_2(.din(w_dff_B_TtRhlFxB1_2),.dout(w_dff_B_a8ULsxYn6_2),.clk(gclk));
	jdff dff_B_20Hn3ifm2_2(.din(w_dff_B_a8ULsxYn6_2),.dout(w_dff_B_20Hn3ifm2_2),.clk(gclk));
	jdff dff_B_Ra7rGvSp3_2(.din(w_dff_B_20Hn3ifm2_2),.dout(w_dff_B_Ra7rGvSp3_2),.clk(gclk));
	jdff dff_B_khnGhDRn9_2(.din(w_dff_B_Ra7rGvSp3_2),.dout(w_dff_B_khnGhDRn9_2),.clk(gclk));
	jdff dff_B_kwoqfqHK8_2(.din(w_dff_B_khnGhDRn9_2),.dout(w_dff_B_kwoqfqHK8_2),.clk(gclk));
	jdff dff_B_NrlJz5gm7_2(.din(w_dff_B_kwoqfqHK8_2),.dout(w_dff_B_NrlJz5gm7_2),.clk(gclk));
	jdff dff_B_fi0giJp52_2(.din(w_dff_B_NrlJz5gm7_2),.dout(w_dff_B_fi0giJp52_2),.clk(gclk));
	jdff dff_B_9XSGrxv58_2(.din(w_dff_B_fi0giJp52_2),.dout(w_dff_B_9XSGrxv58_2),.clk(gclk));
	jdff dff_B_oRg94UzK3_2(.din(w_dff_B_9XSGrxv58_2),.dout(w_dff_B_oRg94UzK3_2),.clk(gclk));
	jdff dff_B_WQnTw4us2_2(.din(w_dff_B_oRg94UzK3_2),.dout(w_dff_B_WQnTw4us2_2),.clk(gclk));
	jdff dff_B_0ajdEipX5_2(.din(w_dff_B_WQnTw4us2_2),.dout(w_dff_B_0ajdEipX5_2),.clk(gclk));
	jdff dff_B_tVRV7OsE9_2(.din(w_dff_B_0ajdEipX5_2),.dout(w_dff_B_tVRV7OsE9_2),.clk(gclk));
	jdff dff_B_eg24WkAQ6_2(.din(w_dff_B_tVRV7OsE9_2),.dout(w_dff_B_eg24WkAQ6_2),.clk(gclk));
	jdff dff_B_0Y6pU22K5_2(.din(w_dff_B_eg24WkAQ6_2),.dout(w_dff_B_0Y6pU22K5_2),.clk(gclk));
	jdff dff_B_5BmTqeRt2_2(.din(n1052),.dout(w_dff_B_5BmTqeRt2_2),.clk(gclk));
	jdff dff_B_yOVGUYnu7_1(.din(n1050),.dout(w_dff_B_yOVGUYnu7_1),.clk(gclk));
	jdff dff_B_oMu2hVNG1_2(.din(n951),.dout(w_dff_B_oMu2hVNG1_2),.clk(gclk));
	jdff dff_B_jTqIiLCG7_2(.din(w_dff_B_oMu2hVNG1_2),.dout(w_dff_B_jTqIiLCG7_2),.clk(gclk));
	jdff dff_B_E9atFrem2_2(.din(w_dff_B_jTqIiLCG7_2),.dout(w_dff_B_E9atFrem2_2),.clk(gclk));
	jdff dff_B_kO3khuXJ1_2(.din(w_dff_B_E9atFrem2_2),.dout(w_dff_B_kO3khuXJ1_2),.clk(gclk));
	jdff dff_B_9Rt4fsWD2_2(.din(w_dff_B_kO3khuXJ1_2),.dout(w_dff_B_9Rt4fsWD2_2),.clk(gclk));
	jdff dff_B_QPKubA1A4_2(.din(w_dff_B_9Rt4fsWD2_2),.dout(w_dff_B_QPKubA1A4_2),.clk(gclk));
	jdff dff_B_bSn9ApwM1_2(.din(w_dff_B_QPKubA1A4_2),.dout(w_dff_B_bSn9ApwM1_2),.clk(gclk));
	jdff dff_B_lyLk7HRX3_2(.din(w_dff_B_bSn9ApwM1_2),.dout(w_dff_B_lyLk7HRX3_2),.clk(gclk));
	jdff dff_B_1QqkWXZU5_2(.din(w_dff_B_lyLk7HRX3_2),.dout(w_dff_B_1QqkWXZU5_2),.clk(gclk));
	jdff dff_B_8Gn8jUY98_2(.din(w_dff_B_1QqkWXZU5_2),.dout(w_dff_B_8Gn8jUY98_2),.clk(gclk));
	jdff dff_B_pHqETEZS1_2(.din(w_dff_B_8Gn8jUY98_2),.dout(w_dff_B_pHqETEZS1_2),.clk(gclk));
	jdff dff_B_Aq9UJTwB0_2(.din(w_dff_B_pHqETEZS1_2),.dout(w_dff_B_Aq9UJTwB0_2),.clk(gclk));
	jdff dff_B_zHdONj456_2(.din(w_dff_B_Aq9UJTwB0_2),.dout(w_dff_B_zHdONj456_2),.clk(gclk));
	jdff dff_B_iHNk5Cbt5_2(.din(w_dff_B_zHdONj456_2),.dout(w_dff_B_iHNk5Cbt5_2),.clk(gclk));
	jdff dff_B_yhbpxAeA1_2(.din(w_dff_B_iHNk5Cbt5_2),.dout(w_dff_B_yhbpxAeA1_2),.clk(gclk));
	jdff dff_B_YxOVq6wy2_2(.din(w_dff_B_yhbpxAeA1_2),.dout(w_dff_B_YxOVq6wy2_2),.clk(gclk));
	jdff dff_B_qFjfjO0G7_2(.din(w_dff_B_YxOVq6wy2_2),.dout(w_dff_B_qFjfjO0G7_2),.clk(gclk));
	jdff dff_B_uXaoQqx24_2(.din(w_dff_B_qFjfjO0G7_2),.dout(w_dff_B_uXaoQqx24_2),.clk(gclk));
	jdff dff_B_vZC20l9v4_2(.din(w_dff_B_uXaoQqx24_2),.dout(w_dff_B_vZC20l9v4_2),.clk(gclk));
	jdff dff_B_paTa60LQ3_2(.din(w_dff_B_vZC20l9v4_2),.dout(w_dff_B_paTa60LQ3_2),.clk(gclk));
	jdff dff_B_fjui4HUZ8_2(.din(w_dff_B_paTa60LQ3_2),.dout(w_dff_B_fjui4HUZ8_2),.clk(gclk));
	jdff dff_B_C4UnGJQX5_2(.din(w_dff_B_fjui4HUZ8_2),.dout(w_dff_B_C4UnGJQX5_2),.clk(gclk));
	jdff dff_B_wKuCAcoD5_2(.din(w_dff_B_C4UnGJQX5_2),.dout(w_dff_B_wKuCAcoD5_2),.clk(gclk));
	jdff dff_B_WxjeCSRy0_2(.din(w_dff_B_wKuCAcoD5_2),.dout(w_dff_B_WxjeCSRy0_2),.clk(gclk));
	jdff dff_B_50ZXxNf37_2(.din(w_dff_B_WxjeCSRy0_2),.dout(w_dff_B_50ZXxNf37_2),.clk(gclk));
	jdff dff_B_yoJ1bUnw9_2(.din(w_dff_B_50ZXxNf37_2),.dout(w_dff_B_yoJ1bUnw9_2),.clk(gclk));
	jdff dff_B_BbhDxqc18_1(.din(n952),.dout(w_dff_B_BbhDxqc18_1),.clk(gclk));
	jdff dff_B_EPVCfF0o7_2(.din(n846),.dout(w_dff_B_EPVCfF0o7_2),.clk(gclk));
	jdff dff_B_7cfyAm1b4_2(.din(w_dff_B_EPVCfF0o7_2),.dout(w_dff_B_7cfyAm1b4_2),.clk(gclk));
	jdff dff_B_RYL4EtQe0_2(.din(w_dff_B_7cfyAm1b4_2),.dout(w_dff_B_RYL4EtQe0_2),.clk(gclk));
	jdff dff_B_J7O2bJi86_2(.din(w_dff_B_RYL4EtQe0_2),.dout(w_dff_B_J7O2bJi86_2),.clk(gclk));
	jdff dff_B_8cokMvvD1_2(.din(w_dff_B_J7O2bJi86_2),.dout(w_dff_B_8cokMvvD1_2),.clk(gclk));
	jdff dff_B_i6vpuMVL1_2(.din(w_dff_B_8cokMvvD1_2),.dout(w_dff_B_i6vpuMVL1_2),.clk(gclk));
	jdff dff_B_bQlFTCX68_2(.din(w_dff_B_i6vpuMVL1_2),.dout(w_dff_B_bQlFTCX68_2),.clk(gclk));
	jdff dff_B_mgQUN2Vv2_2(.din(w_dff_B_bQlFTCX68_2),.dout(w_dff_B_mgQUN2Vv2_2),.clk(gclk));
	jdff dff_B_U7lemMSr0_2(.din(w_dff_B_mgQUN2Vv2_2),.dout(w_dff_B_U7lemMSr0_2),.clk(gclk));
	jdff dff_B_tKcxuTBc5_2(.din(w_dff_B_U7lemMSr0_2),.dout(w_dff_B_tKcxuTBc5_2),.clk(gclk));
	jdff dff_B_JDKuEmjY7_2(.din(w_dff_B_tKcxuTBc5_2),.dout(w_dff_B_JDKuEmjY7_2),.clk(gclk));
	jdff dff_B_lYqRj3aA4_2(.din(w_dff_B_JDKuEmjY7_2),.dout(w_dff_B_lYqRj3aA4_2),.clk(gclk));
	jdff dff_B_RSYX8dfh4_2(.din(w_dff_B_lYqRj3aA4_2),.dout(w_dff_B_RSYX8dfh4_2),.clk(gclk));
	jdff dff_B_HyYmUasu3_2(.din(w_dff_B_RSYX8dfh4_2),.dout(w_dff_B_HyYmUasu3_2),.clk(gclk));
	jdff dff_B_GpYfbHrv9_2(.din(w_dff_B_HyYmUasu3_2),.dout(w_dff_B_GpYfbHrv9_2),.clk(gclk));
	jdff dff_B_gCh1ZfjT8_2(.din(w_dff_B_GpYfbHrv9_2),.dout(w_dff_B_gCh1ZfjT8_2),.clk(gclk));
	jdff dff_B_s7oWDwCD0_2(.din(w_dff_B_gCh1ZfjT8_2),.dout(w_dff_B_s7oWDwCD0_2),.clk(gclk));
	jdff dff_B_bYBsYAXr2_2(.din(w_dff_B_s7oWDwCD0_2),.dout(w_dff_B_bYBsYAXr2_2),.clk(gclk));
	jdff dff_B_tHQkTJFO3_2(.din(w_dff_B_bYBsYAXr2_2),.dout(w_dff_B_tHQkTJFO3_2),.clk(gclk));
	jdff dff_B_Ig1ukQAh9_2(.din(w_dff_B_tHQkTJFO3_2),.dout(w_dff_B_Ig1ukQAh9_2),.clk(gclk));
	jdff dff_B_f8GuRuGt0_2(.din(w_dff_B_Ig1ukQAh9_2),.dout(w_dff_B_f8GuRuGt0_2),.clk(gclk));
	jdff dff_B_mtaOLY4K6_2(.din(w_dff_B_f8GuRuGt0_2),.dout(w_dff_B_mtaOLY4K6_2),.clk(gclk));
	jdff dff_B_eGaIVF2z0_2(.din(w_dff_B_mtaOLY4K6_2),.dout(w_dff_B_eGaIVF2z0_2),.clk(gclk));
	jdff dff_B_32BBUETR6_2(.din(w_dff_B_eGaIVF2z0_2),.dout(w_dff_B_32BBUETR6_2),.clk(gclk));
	jdff dff_B_jan9yoBt7_1(.din(n847),.dout(w_dff_B_jan9yoBt7_1),.clk(gclk));
	jdff dff_B_QefQ0Vzc8_2(.din(n747),.dout(w_dff_B_QefQ0Vzc8_2),.clk(gclk));
	jdff dff_B_EL7OHtVR9_2(.din(w_dff_B_QefQ0Vzc8_2),.dout(w_dff_B_EL7OHtVR9_2),.clk(gclk));
	jdff dff_B_sPgxBzVE7_2(.din(w_dff_B_EL7OHtVR9_2),.dout(w_dff_B_sPgxBzVE7_2),.clk(gclk));
	jdff dff_B_WEC35h5t6_2(.din(w_dff_B_sPgxBzVE7_2),.dout(w_dff_B_WEC35h5t6_2),.clk(gclk));
	jdff dff_B_P7huY2LL6_2(.din(w_dff_B_WEC35h5t6_2),.dout(w_dff_B_P7huY2LL6_2),.clk(gclk));
	jdff dff_B_tYv9De148_2(.din(w_dff_B_P7huY2LL6_2),.dout(w_dff_B_tYv9De148_2),.clk(gclk));
	jdff dff_B_m4lMnMzN0_2(.din(w_dff_B_tYv9De148_2),.dout(w_dff_B_m4lMnMzN0_2),.clk(gclk));
	jdff dff_B_oCvDsXSc9_2(.din(w_dff_B_m4lMnMzN0_2),.dout(w_dff_B_oCvDsXSc9_2),.clk(gclk));
	jdff dff_B_OsOzXHUD2_2(.din(w_dff_B_oCvDsXSc9_2),.dout(w_dff_B_OsOzXHUD2_2),.clk(gclk));
	jdff dff_B_NWwma4Et0_2(.din(w_dff_B_OsOzXHUD2_2),.dout(w_dff_B_NWwma4Et0_2),.clk(gclk));
	jdff dff_B_fMfR0em89_2(.din(w_dff_B_NWwma4Et0_2),.dout(w_dff_B_fMfR0em89_2),.clk(gclk));
	jdff dff_B_O1raQNuD4_2(.din(w_dff_B_fMfR0em89_2),.dout(w_dff_B_O1raQNuD4_2),.clk(gclk));
	jdff dff_B_43l9vTg94_2(.din(w_dff_B_O1raQNuD4_2),.dout(w_dff_B_43l9vTg94_2),.clk(gclk));
	jdff dff_B_jcmNCKaf0_2(.din(w_dff_B_43l9vTg94_2),.dout(w_dff_B_jcmNCKaf0_2),.clk(gclk));
	jdff dff_B_ZWMPaf6m1_2(.din(w_dff_B_jcmNCKaf0_2),.dout(w_dff_B_ZWMPaf6m1_2),.clk(gclk));
	jdff dff_B_nDKEzlx21_2(.din(w_dff_B_ZWMPaf6m1_2),.dout(w_dff_B_nDKEzlx21_2),.clk(gclk));
	jdff dff_B_ZeBBeoNo6_2(.din(w_dff_B_nDKEzlx21_2),.dout(w_dff_B_ZeBBeoNo6_2),.clk(gclk));
	jdff dff_B_zHdj9PRa7_2(.din(w_dff_B_ZeBBeoNo6_2),.dout(w_dff_B_zHdj9PRa7_2),.clk(gclk));
	jdff dff_B_aD7xgN5p8_2(.din(w_dff_B_zHdj9PRa7_2),.dout(w_dff_B_aD7xgN5p8_2),.clk(gclk));
	jdff dff_B_ghkkU9EK4_2(.din(w_dff_B_aD7xgN5p8_2),.dout(w_dff_B_ghkkU9EK4_2),.clk(gclk));
	jdff dff_B_7XrSf3Kd8_2(.din(w_dff_B_ghkkU9EK4_2),.dout(w_dff_B_7XrSf3Kd8_2),.clk(gclk));
	jdff dff_B_Ge66VRId2_2(.din(w_dff_B_7XrSf3Kd8_2),.dout(w_dff_B_Ge66VRId2_2),.clk(gclk));
	jdff dff_B_NjSLxxAi9_1(.din(n748),.dout(w_dff_B_NjSLxxAi9_1),.clk(gclk));
	jdff dff_B_0fm2pvKd1_2(.din(n654),.dout(w_dff_B_0fm2pvKd1_2),.clk(gclk));
	jdff dff_B_gOinbKHi9_2(.din(w_dff_B_0fm2pvKd1_2),.dout(w_dff_B_gOinbKHi9_2),.clk(gclk));
	jdff dff_B_P1nDAfVW4_2(.din(w_dff_B_gOinbKHi9_2),.dout(w_dff_B_P1nDAfVW4_2),.clk(gclk));
	jdff dff_B_jaiYtPvQ5_2(.din(w_dff_B_P1nDAfVW4_2),.dout(w_dff_B_jaiYtPvQ5_2),.clk(gclk));
	jdff dff_B_ZBhRdYHg0_2(.din(w_dff_B_jaiYtPvQ5_2),.dout(w_dff_B_ZBhRdYHg0_2),.clk(gclk));
	jdff dff_B_sDMuL2AP2_2(.din(w_dff_B_ZBhRdYHg0_2),.dout(w_dff_B_sDMuL2AP2_2),.clk(gclk));
	jdff dff_B_ZovVYjIq2_2(.din(w_dff_B_sDMuL2AP2_2),.dout(w_dff_B_ZovVYjIq2_2),.clk(gclk));
	jdff dff_B_mEMkvezv5_2(.din(w_dff_B_ZovVYjIq2_2),.dout(w_dff_B_mEMkvezv5_2),.clk(gclk));
	jdff dff_B_wRk4F03L6_2(.din(w_dff_B_mEMkvezv5_2),.dout(w_dff_B_wRk4F03L6_2),.clk(gclk));
	jdff dff_B_UXcQQUlj7_2(.din(w_dff_B_wRk4F03L6_2),.dout(w_dff_B_UXcQQUlj7_2),.clk(gclk));
	jdff dff_B_IDHaq1Xc3_2(.din(w_dff_B_UXcQQUlj7_2),.dout(w_dff_B_IDHaq1Xc3_2),.clk(gclk));
	jdff dff_B_nzb8FYZJ4_2(.din(w_dff_B_IDHaq1Xc3_2),.dout(w_dff_B_nzb8FYZJ4_2),.clk(gclk));
	jdff dff_B_TWuDv1Zn6_2(.din(w_dff_B_nzb8FYZJ4_2),.dout(w_dff_B_TWuDv1Zn6_2),.clk(gclk));
	jdff dff_B_Nu0zq7kP8_2(.din(w_dff_B_TWuDv1Zn6_2),.dout(w_dff_B_Nu0zq7kP8_2),.clk(gclk));
	jdff dff_B_yeAU6gWp0_2(.din(w_dff_B_Nu0zq7kP8_2),.dout(w_dff_B_yeAU6gWp0_2),.clk(gclk));
	jdff dff_B_3tIvfcNf7_2(.din(w_dff_B_yeAU6gWp0_2),.dout(w_dff_B_3tIvfcNf7_2),.clk(gclk));
	jdff dff_B_BjlvYQhT3_2(.din(w_dff_B_3tIvfcNf7_2),.dout(w_dff_B_BjlvYQhT3_2),.clk(gclk));
	jdff dff_B_AlUyikoN8_2(.din(w_dff_B_BjlvYQhT3_2),.dout(w_dff_B_AlUyikoN8_2),.clk(gclk));
	jdff dff_B_bn6AZRWZ8_2(.din(w_dff_B_AlUyikoN8_2),.dout(w_dff_B_bn6AZRWZ8_2),.clk(gclk));
	jdff dff_B_jZmxLYdm6_2(.din(w_dff_B_bn6AZRWZ8_2),.dout(w_dff_B_jZmxLYdm6_2),.clk(gclk));
	jdff dff_B_uqn7ykRC9_1(.din(n655),.dout(w_dff_B_uqn7ykRC9_1),.clk(gclk));
	jdff dff_B_3PRDOd840_2(.din(n568),.dout(w_dff_B_3PRDOd840_2),.clk(gclk));
	jdff dff_B_Nmm5tsaQ3_2(.din(w_dff_B_3PRDOd840_2),.dout(w_dff_B_Nmm5tsaQ3_2),.clk(gclk));
	jdff dff_B_66kp1h185_2(.din(w_dff_B_Nmm5tsaQ3_2),.dout(w_dff_B_66kp1h185_2),.clk(gclk));
	jdff dff_B_2QyH3EDX1_2(.din(w_dff_B_66kp1h185_2),.dout(w_dff_B_2QyH3EDX1_2),.clk(gclk));
	jdff dff_B_GYXaY3jF1_2(.din(w_dff_B_2QyH3EDX1_2),.dout(w_dff_B_GYXaY3jF1_2),.clk(gclk));
	jdff dff_B_Xbdt1keg6_2(.din(w_dff_B_GYXaY3jF1_2),.dout(w_dff_B_Xbdt1keg6_2),.clk(gclk));
	jdff dff_B_nxx84m0C9_2(.din(w_dff_B_Xbdt1keg6_2),.dout(w_dff_B_nxx84m0C9_2),.clk(gclk));
	jdff dff_B_muiRi0J69_2(.din(w_dff_B_nxx84m0C9_2),.dout(w_dff_B_muiRi0J69_2),.clk(gclk));
	jdff dff_B_MweqWHDe4_2(.din(w_dff_B_muiRi0J69_2),.dout(w_dff_B_MweqWHDe4_2),.clk(gclk));
	jdff dff_B_LYJRX0Of8_2(.din(w_dff_B_MweqWHDe4_2),.dout(w_dff_B_LYJRX0Of8_2),.clk(gclk));
	jdff dff_B_iidRc1wU2_2(.din(w_dff_B_LYJRX0Of8_2),.dout(w_dff_B_iidRc1wU2_2),.clk(gclk));
	jdff dff_B_2SywCMjB9_2(.din(w_dff_B_iidRc1wU2_2),.dout(w_dff_B_2SywCMjB9_2),.clk(gclk));
	jdff dff_B_ImvNnBDr2_2(.din(w_dff_B_2SywCMjB9_2),.dout(w_dff_B_ImvNnBDr2_2),.clk(gclk));
	jdff dff_B_mp39UK9t7_2(.din(w_dff_B_ImvNnBDr2_2),.dout(w_dff_B_mp39UK9t7_2),.clk(gclk));
	jdff dff_B_wWR30lxS2_2(.din(w_dff_B_mp39UK9t7_2),.dout(w_dff_B_wWR30lxS2_2),.clk(gclk));
	jdff dff_B_75CQSFLO5_2(.din(w_dff_B_wWR30lxS2_2),.dout(w_dff_B_75CQSFLO5_2),.clk(gclk));
	jdff dff_B_BrbHYZtq1_2(.din(w_dff_B_75CQSFLO5_2),.dout(w_dff_B_BrbHYZtq1_2),.clk(gclk));
	jdff dff_B_ESOkehGZ8_2(.din(w_dff_B_BrbHYZtq1_2),.dout(w_dff_B_ESOkehGZ8_2),.clk(gclk));
	jdff dff_B_DADHk8B11_1(.din(n569),.dout(w_dff_B_DADHk8B11_1),.clk(gclk));
	jdff dff_B_rngTF36W5_2(.din(n489),.dout(w_dff_B_rngTF36W5_2),.clk(gclk));
	jdff dff_B_vxPAZSQT2_2(.din(w_dff_B_rngTF36W5_2),.dout(w_dff_B_vxPAZSQT2_2),.clk(gclk));
	jdff dff_B_pOzWmgTj2_2(.din(w_dff_B_vxPAZSQT2_2),.dout(w_dff_B_pOzWmgTj2_2),.clk(gclk));
	jdff dff_B_2Smr4jtq5_2(.din(w_dff_B_pOzWmgTj2_2),.dout(w_dff_B_2Smr4jtq5_2),.clk(gclk));
	jdff dff_B_cRro3xIJ7_2(.din(w_dff_B_2Smr4jtq5_2),.dout(w_dff_B_cRro3xIJ7_2),.clk(gclk));
	jdff dff_B_2m9yRjZT5_2(.din(w_dff_B_cRro3xIJ7_2),.dout(w_dff_B_2m9yRjZT5_2),.clk(gclk));
	jdff dff_B_BwelrUXL4_2(.din(w_dff_B_2m9yRjZT5_2),.dout(w_dff_B_BwelrUXL4_2),.clk(gclk));
	jdff dff_B_hE3pszSi8_2(.din(w_dff_B_BwelrUXL4_2),.dout(w_dff_B_hE3pszSi8_2),.clk(gclk));
	jdff dff_B_LTlBw1895_2(.din(w_dff_B_hE3pszSi8_2),.dout(w_dff_B_LTlBw1895_2),.clk(gclk));
	jdff dff_B_vdoNNJG76_2(.din(w_dff_B_LTlBw1895_2),.dout(w_dff_B_vdoNNJG76_2),.clk(gclk));
	jdff dff_B_XkAZ7FFS1_2(.din(w_dff_B_vdoNNJG76_2),.dout(w_dff_B_XkAZ7FFS1_2),.clk(gclk));
	jdff dff_B_dPCNRQlL7_2(.din(w_dff_B_XkAZ7FFS1_2),.dout(w_dff_B_dPCNRQlL7_2),.clk(gclk));
	jdff dff_B_1rDuuBOu5_2(.din(w_dff_B_dPCNRQlL7_2),.dout(w_dff_B_1rDuuBOu5_2),.clk(gclk));
	jdff dff_B_JSPN5e8Y2_2(.din(w_dff_B_1rDuuBOu5_2),.dout(w_dff_B_JSPN5e8Y2_2),.clk(gclk));
	jdff dff_B_KMEdhYIr1_2(.din(w_dff_B_JSPN5e8Y2_2),.dout(w_dff_B_KMEdhYIr1_2),.clk(gclk));
	jdff dff_B_TVLIDS2Y9_2(.din(w_dff_B_KMEdhYIr1_2),.dout(w_dff_B_TVLIDS2Y9_2),.clk(gclk));
	jdff dff_B_uYzApxJz9_1(.din(n490),.dout(w_dff_B_uYzApxJz9_1),.clk(gclk));
	jdff dff_B_LR37DUxK7_2(.din(n417),.dout(w_dff_B_LR37DUxK7_2),.clk(gclk));
	jdff dff_B_nrKd9pOE6_2(.din(w_dff_B_LR37DUxK7_2),.dout(w_dff_B_nrKd9pOE6_2),.clk(gclk));
	jdff dff_B_EFeoN9f90_2(.din(w_dff_B_nrKd9pOE6_2),.dout(w_dff_B_EFeoN9f90_2),.clk(gclk));
	jdff dff_B_33g02Ddm9_2(.din(w_dff_B_EFeoN9f90_2),.dout(w_dff_B_33g02Ddm9_2),.clk(gclk));
	jdff dff_B_f6wMn9GJ3_2(.din(w_dff_B_33g02Ddm9_2),.dout(w_dff_B_f6wMn9GJ3_2),.clk(gclk));
	jdff dff_B_6703W9K22_2(.din(w_dff_B_f6wMn9GJ3_2),.dout(w_dff_B_6703W9K22_2),.clk(gclk));
	jdff dff_B_iq5urRMH3_2(.din(w_dff_B_6703W9K22_2),.dout(w_dff_B_iq5urRMH3_2),.clk(gclk));
	jdff dff_B_w9PQPxu29_2(.din(w_dff_B_iq5urRMH3_2),.dout(w_dff_B_w9PQPxu29_2),.clk(gclk));
	jdff dff_B_Uf5WZZVs4_2(.din(w_dff_B_w9PQPxu29_2),.dout(w_dff_B_Uf5WZZVs4_2),.clk(gclk));
	jdff dff_B_V5KTX8M17_2(.din(w_dff_B_Uf5WZZVs4_2),.dout(w_dff_B_V5KTX8M17_2),.clk(gclk));
	jdff dff_B_EFP6BrTs5_2(.din(w_dff_B_V5KTX8M17_2),.dout(w_dff_B_EFP6BrTs5_2),.clk(gclk));
	jdff dff_B_hHuZHrLA4_2(.din(w_dff_B_EFP6BrTs5_2),.dout(w_dff_B_hHuZHrLA4_2),.clk(gclk));
	jdff dff_B_jrpIEsyb2_2(.din(w_dff_B_hHuZHrLA4_2),.dout(w_dff_B_jrpIEsyb2_2),.clk(gclk));
	jdff dff_B_MGReRU7o3_2(.din(w_dff_B_jrpIEsyb2_2),.dout(w_dff_B_MGReRU7o3_2),.clk(gclk));
	jdff dff_B_TIRuYEFC5_1(.din(n418),.dout(w_dff_B_TIRuYEFC5_1),.clk(gclk));
	jdff dff_B_ADlkfaBT0_2(.din(n353),.dout(w_dff_B_ADlkfaBT0_2),.clk(gclk));
	jdff dff_B_8riLP2J56_2(.din(w_dff_B_ADlkfaBT0_2),.dout(w_dff_B_8riLP2J56_2),.clk(gclk));
	jdff dff_B_qIFAkXQd9_2(.din(w_dff_B_8riLP2J56_2),.dout(w_dff_B_qIFAkXQd9_2),.clk(gclk));
	jdff dff_B_cxN66kwZ5_2(.din(w_dff_B_qIFAkXQd9_2),.dout(w_dff_B_cxN66kwZ5_2),.clk(gclk));
	jdff dff_B_hh2qU7rz7_2(.din(w_dff_B_cxN66kwZ5_2),.dout(w_dff_B_hh2qU7rz7_2),.clk(gclk));
	jdff dff_B_Bp5l5lz53_2(.din(w_dff_B_hh2qU7rz7_2),.dout(w_dff_B_Bp5l5lz53_2),.clk(gclk));
	jdff dff_B_TXqGHLxH2_2(.din(w_dff_B_Bp5l5lz53_2),.dout(w_dff_B_TXqGHLxH2_2),.clk(gclk));
	jdff dff_B_sN9U3zfN4_2(.din(w_dff_B_TXqGHLxH2_2),.dout(w_dff_B_sN9U3zfN4_2),.clk(gclk));
	jdff dff_B_PkOqJCLN3_2(.din(w_dff_B_sN9U3zfN4_2),.dout(w_dff_B_PkOqJCLN3_2),.clk(gclk));
	jdff dff_B_6kGhrfXn7_2(.din(w_dff_B_PkOqJCLN3_2),.dout(w_dff_B_6kGhrfXn7_2),.clk(gclk));
	jdff dff_B_wpMqGPca1_2(.din(w_dff_B_6kGhrfXn7_2),.dout(w_dff_B_wpMqGPca1_2),.clk(gclk));
	jdff dff_B_Z8BhLEVE3_2(.din(w_dff_B_wpMqGPca1_2),.dout(w_dff_B_Z8BhLEVE3_2),.clk(gclk));
	jdff dff_B_DwjbHO0w1_1(.din(n354),.dout(w_dff_B_DwjbHO0w1_1),.clk(gclk));
	jdff dff_B_lFgjC9cs2_2(.din(n295),.dout(w_dff_B_lFgjC9cs2_2),.clk(gclk));
	jdff dff_B_FoT90ABF2_2(.din(w_dff_B_lFgjC9cs2_2),.dout(w_dff_B_FoT90ABF2_2),.clk(gclk));
	jdff dff_B_X8NI0hMe0_2(.din(w_dff_B_FoT90ABF2_2),.dout(w_dff_B_X8NI0hMe0_2),.clk(gclk));
	jdff dff_B_RSeWZT0v9_2(.din(w_dff_B_X8NI0hMe0_2),.dout(w_dff_B_RSeWZT0v9_2),.clk(gclk));
	jdff dff_B_hiLpQbpC1_2(.din(w_dff_B_RSeWZT0v9_2),.dout(w_dff_B_hiLpQbpC1_2),.clk(gclk));
	jdff dff_B_hTOVazCx9_2(.din(w_dff_B_hiLpQbpC1_2),.dout(w_dff_B_hTOVazCx9_2),.clk(gclk));
	jdff dff_B_OeB7QDbi6_2(.din(w_dff_B_hTOVazCx9_2),.dout(w_dff_B_OeB7QDbi6_2),.clk(gclk));
	jdff dff_B_z6rdy2TZ7_2(.din(w_dff_B_OeB7QDbi6_2),.dout(w_dff_B_z6rdy2TZ7_2),.clk(gclk));
	jdff dff_B_ofmkEbZo1_2(.din(w_dff_B_z6rdy2TZ7_2),.dout(w_dff_B_ofmkEbZo1_2),.clk(gclk));
	jdff dff_B_M5SDinXi6_2(.din(w_dff_B_ofmkEbZo1_2),.dout(w_dff_B_M5SDinXi6_2),.clk(gclk));
	jdff dff_B_ZVn1JATL0_1(.din(n296),.dout(w_dff_B_ZVn1JATL0_1),.clk(gclk));
	jdff dff_B_CSHfwZK40_2(.din(n244),.dout(w_dff_B_CSHfwZK40_2),.clk(gclk));
	jdff dff_B_v4tjxi2c9_2(.din(w_dff_B_CSHfwZK40_2),.dout(w_dff_B_v4tjxi2c9_2),.clk(gclk));
	jdff dff_B_tKhnYXT06_2(.din(w_dff_B_v4tjxi2c9_2),.dout(w_dff_B_tKhnYXT06_2),.clk(gclk));
	jdff dff_B_GTq1WUGl4_2(.din(w_dff_B_tKhnYXT06_2),.dout(w_dff_B_GTq1WUGl4_2),.clk(gclk));
	jdff dff_B_y5b8JW3C0_2(.din(w_dff_B_GTq1WUGl4_2),.dout(w_dff_B_y5b8JW3C0_2),.clk(gclk));
	jdff dff_B_undiNxAR0_2(.din(w_dff_B_y5b8JW3C0_2),.dout(w_dff_B_undiNxAR0_2),.clk(gclk));
	jdff dff_B_cx3VEgZ42_2(.din(w_dff_B_undiNxAR0_2),.dout(w_dff_B_cx3VEgZ42_2),.clk(gclk));
	jdff dff_B_xmctGBj18_2(.din(w_dff_B_cx3VEgZ42_2),.dout(w_dff_B_xmctGBj18_2),.clk(gclk));
	jdff dff_B_TOOe7Jno0_2(.din(n247),.dout(w_dff_B_TOOe7Jno0_2),.clk(gclk));
	jdff dff_B_nwOQFSQ28_1(.din(n245),.dout(w_dff_B_nwOQFSQ28_1),.clk(gclk));
	jdff dff_B_t4ge3YhN4_2(.din(n201),.dout(w_dff_B_t4ge3YhN4_2),.clk(gclk));
	jdff dff_B_YoBF9TRb0_2(.din(w_dff_B_t4ge3YhN4_2),.dout(w_dff_B_YoBF9TRb0_2),.clk(gclk));
	jdff dff_B_l96uTqkB8_2(.din(w_dff_B_YoBF9TRb0_2),.dout(w_dff_B_l96uTqkB8_2),.clk(gclk));
	jdff dff_B_Fxt6WSZz7_2(.din(w_dff_B_l96uTqkB8_2),.dout(w_dff_B_Fxt6WSZz7_2),.clk(gclk));
	jdff dff_B_nNtLFeVt4_2(.din(w_dff_B_Fxt6WSZz7_2),.dout(w_dff_B_nNtLFeVt4_2),.clk(gclk));
	jdff dff_B_GK5VE46Q3_1(.din(n202),.dout(w_dff_B_GK5VE46Q3_1),.clk(gclk));
	jdff dff_B_vn3oQZHB7_0(.din(n173),.dout(w_dff_B_vn3oQZHB7_0),.clk(gclk));
	jdff dff_B_JHv1FRYm4_2(.din(n165),.dout(w_dff_B_JHv1FRYm4_2),.clk(gclk));
	jdff dff_B_GVY0OuzW2_2(.din(w_dff_B_JHv1FRYm4_2),.dout(w_dff_B_GVY0OuzW2_2),.clk(gclk));
	jdff dff_B_mHt9CsSX7_2(.din(w_dff_B_GVY0OuzW2_2),.dout(w_dff_B_mHt9CsSX7_2),.clk(gclk));
	jdff dff_B_I530oxMV5_1(.din(n167),.dout(w_dff_B_I530oxMV5_1),.clk(gclk));
	jdff dff_B_tNXDlT0N2_1(.din(w_dff_B_I530oxMV5_1),.dout(w_dff_B_tNXDlT0N2_1),.clk(gclk));
	jdff dff_A_ofpJNDQw4_0(.dout(w_n132_0[0]),.din(w_dff_A_ofpJNDQw4_0),.clk(gclk));
	jdff dff_A_kmyc9HRq1_0(.dout(w_dff_A_ofpJNDQw4_0),.din(w_dff_A_kmyc9HRq1_0),.clk(gclk));
	jdff dff_B_TRezTEAG8_2(.din(n1337),.dout(w_dff_B_TRezTEAG8_2),.clk(gclk));
	jdff dff_B_3D2mMVj74_2(.din(w_dff_B_TRezTEAG8_2),.dout(w_dff_B_3D2mMVj74_2),.clk(gclk));
	jdff dff_B_cEx3tPYS7_1(.din(n1335),.dout(w_dff_B_cEx3tPYS7_1),.clk(gclk));
	jdff dff_B_7UkinoS60_2(.din(n1248),.dout(w_dff_B_7UkinoS60_2),.clk(gclk));
	jdff dff_B_6c18BDlQ0_2(.din(w_dff_B_7UkinoS60_2),.dout(w_dff_B_6c18BDlQ0_2),.clk(gclk));
	jdff dff_B_SdsxSNPh9_2(.din(w_dff_B_6c18BDlQ0_2),.dout(w_dff_B_SdsxSNPh9_2),.clk(gclk));
	jdff dff_B_TxGXkzvz5_2(.din(w_dff_B_SdsxSNPh9_2),.dout(w_dff_B_TxGXkzvz5_2),.clk(gclk));
	jdff dff_B_4KYFoQxi0_2(.din(w_dff_B_TxGXkzvz5_2),.dout(w_dff_B_4KYFoQxi0_2),.clk(gclk));
	jdff dff_B_lQ2G17Qz8_2(.din(w_dff_B_4KYFoQxi0_2),.dout(w_dff_B_lQ2G17Qz8_2),.clk(gclk));
	jdff dff_B_9TD4OPUa6_2(.din(w_dff_B_lQ2G17Qz8_2),.dout(w_dff_B_9TD4OPUa6_2),.clk(gclk));
	jdff dff_B_fNLJi2wq1_2(.din(w_dff_B_9TD4OPUa6_2),.dout(w_dff_B_fNLJi2wq1_2),.clk(gclk));
	jdff dff_B_3rR88h1H2_2(.din(w_dff_B_fNLJi2wq1_2),.dout(w_dff_B_3rR88h1H2_2),.clk(gclk));
	jdff dff_B_DfGf5iQS9_2(.din(w_dff_B_3rR88h1H2_2),.dout(w_dff_B_DfGf5iQS9_2),.clk(gclk));
	jdff dff_B_NE7dULgf9_2(.din(w_dff_B_DfGf5iQS9_2),.dout(w_dff_B_NE7dULgf9_2),.clk(gclk));
	jdff dff_B_6RbOI03q7_2(.din(w_dff_B_NE7dULgf9_2),.dout(w_dff_B_6RbOI03q7_2),.clk(gclk));
	jdff dff_B_TIhBHJN38_2(.din(w_dff_B_6RbOI03q7_2),.dout(w_dff_B_TIhBHJN38_2),.clk(gclk));
	jdff dff_B_rUM1Tyhb4_2(.din(w_dff_B_TIhBHJN38_2),.dout(w_dff_B_rUM1Tyhb4_2),.clk(gclk));
	jdff dff_B_R8UWnzjE2_2(.din(w_dff_B_rUM1Tyhb4_2),.dout(w_dff_B_R8UWnzjE2_2),.clk(gclk));
	jdff dff_B_04C07ge85_2(.din(w_dff_B_R8UWnzjE2_2),.dout(w_dff_B_04C07ge85_2),.clk(gclk));
	jdff dff_B_5Ho9yZNc3_2(.din(w_dff_B_04C07ge85_2),.dout(w_dff_B_5Ho9yZNc3_2),.clk(gclk));
	jdff dff_B_vvrzDFV91_2(.din(w_dff_B_5Ho9yZNc3_2),.dout(w_dff_B_vvrzDFV91_2),.clk(gclk));
	jdff dff_B_0EluVG4F3_2(.din(w_dff_B_vvrzDFV91_2),.dout(w_dff_B_0EluVG4F3_2),.clk(gclk));
	jdff dff_B_3krL4CMp1_2(.din(w_dff_B_0EluVG4F3_2),.dout(w_dff_B_3krL4CMp1_2),.clk(gclk));
	jdff dff_B_NQtN0yqy5_2(.din(w_dff_B_3krL4CMp1_2),.dout(w_dff_B_NQtN0yqy5_2),.clk(gclk));
	jdff dff_B_AWNRC3NM5_2(.din(w_dff_B_NQtN0yqy5_2),.dout(w_dff_B_AWNRC3NM5_2),.clk(gclk));
	jdff dff_B_g4ISwAUV5_2(.din(w_dff_B_AWNRC3NM5_2),.dout(w_dff_B_g4ISwAUV5_2),.clk(gclk));
	jdff dff_B_h22KO64B1_2(.din(w_dff_B_g4ISwAUV5_2),.dout(w_dff_B_h22KO64B1_2),.clk(gclk));
	jdff dff_B_XCzw0RSu3_2(.din(w_dff_B_h22KO64B1_2),.dout(w_dff_B_XCzw0RSu3_2),.clk(gclk));
	jdff dff_B_mfrlD0bf7_2(.din(w_dff_B_XCzw0RSu3_2),.dout(w_dff_B_mfrlD0bf7_2),.clk(gclk));
	jdff dff_B_itqNusvO0_2(.din(w_dff_B_mfrlD0bf7_2),.dout(w_dff_B_itqNusvO0_2),.clk(gclk));
	jdff dff_B_c6YNWpel9_2(.din(w_dff_B_itqNusvO0_2),.dout(w_dff_B_c6YNWpel9_2),.clk(gclk));
	jdff dff_B_LdHS9SiW6_2(.din(w_dff_B_c6YNWpel9_2),.dout(w_dff_B_LdHS9SiW6_2),.clk(gclk));
	jdff dff_B_BSThKHTZ2_2(.din(w_dff_B_LdHS9SiW6_2),.dout(w_dff_B_BSThKHTZ2_2),.clk(gclk));
	jdff dff_B_ce2nX3sI9_2(.din(w_dff_B_BSThKHTZ2_2),.dout(w_dff_B_ce2nX3sI9_2),.clk(gclk));
	jdff dff_B_L82pt5IS1_2(.din(w_dff_B_ce2nX3sI9_2),.dout(w_dff_B_L82pt5IS1_2),.clk(gclk));
	jdff dff_B_rX4lAxbJ7_2(.din(w_dff_B_L82pt5IS1_2),.dout(w_dff_B_rX4lAxbJ7_2),.clk(gclk));
	jdff dff_B_n79MyZ8t5_2(.din(w_dff_B_rX4lAxbJ7_2),.dout(w_dff_B_n79MyZ8t5_2),.clk(gclk));
	jdff dff_B_akaHYtU43_2(.din(w_dff_B_n79MyZ8t5_2),.dout(w_dff_B_akaHYtU43_2),.clk(gclk));
	jdff dff_B_NAWMwQTb3_1(.din(n1333),.dout(w_dff_B_NAWMwQTb3_1),.clk(gclk));
	jdff dff_A_KykJmTCb5_1(.dout(w_n1251_0[1]),.din(w_dff_A_KykJmTCb5_1),.clk(gclk));
	jdff dff_B_tV69P8c58_1(.din(n1249),.dout(w_dff_B_tV69P8c58_1),.clk(gclk));
	jdff dff_B_08yCCRl85_2(.din(n1158),.dout(w_dff_B_08yCCRl85_2),.clk(gclk));
	jdff dff_B_ega2IOAx1_2(.din(w_dff_B_08yCCRl85_2),.dout(w_dff_B_ega2IOAx1_2),.clk(gclk));
	jdff dff_B_0umbl25E4_2(.din(w_dff_B_ega2IOAx1_2),.dout(w_dff_B_0umbl25E4_2),.clk(gclk));
	jdff dff_B_k3nTJ9lF0_2(.din(w_dff_B_0umbl25E4_2),.dout(w_dff_B_k3nTJ9lF0_2),.clk(gclk));
	jdff dff_B_aCZWGj4y9_2(.din(w_dff_B_k3nTJ9lF0_2),.dout(w_dff_B_aCZWGj4y9_2),.clk(gclk));
	jdff dff_B_gn7HQ4dy4_2(.din(w_dff_B_aCZWGj4y9_2),.dout(w_dff_B_gn7HQ4dy4_2),.clk(gclk));
	jdff dff_B_VoN6N6tk7_2(.din(w_dff_B_gn7HQ4dy4_2),.dout(w_dff_B_VoN6N6tk7_2),.clk(gclk));
	jdff dff_B_F4PEiccT8_2(.din(w_dff_B_VoN6N6tk7_2),.dout(w_dff_B_F4PEiccT8_2),.clk(gclk));
	jdff dff_B_e5iOJsHv3_2(.din(w_dff_B_F4PEiccT8_2),.dout(w_dff_B_e5iOJsHv3_2),.clk(gclk));
	jdff dff_B_MPYbmmth5_2(.din(w_dff_B_e5iOJsHv3_2),.dout(w_dff_B_MPYbmmth5_2),.clk(gclk));
	jdff dff_B_KSKOQreb9_2(.din(w_dff_B_MPYbmmth5_2),.dout(w_dff_B_KSKOQreb9_2),.clk(gclk));
	jdff dff_B_gNcDbPP20_2(.din(w_dff_B_KSKOQreb9_2),.dout(w_dff_B_gNcDbPP20_2),.clk(gclk));
	jdff dff_B_Q4qaNwBi7_2(.din(w_dff_B_gNcDbPP20_2),.dout(w_dff_B_Q4qaNwBi7_2),.clk(gclk));
	jdff dff_B_sWz74AKi9_2(.din(w_dff_B_Q4qaNwBi7_2),.dout(w_dff_B_sWz74AKi9_2),.clk(gclk));
	jdff dff_B_VntqsTvm2_2(.din(w_dff_B_sWz74AKi9_2),.dout(w_dff_B_VntqsTvm2_2),.clk(gclk));
	jdff dff_B_JaYEiOnw1_2(.din(w_dff_B_VntqsTvm2_2),.dout(w_dff_B_JaYEiOnw1_2),.clk(gclk));
	jdff dff_B_JCp4qxlc8_2(.din(w_dff_B_JaYEiOnw1_2),.dout(w_dff_B_JCp4qxlc8_2),.clk(gclk));
	jdff dff_B_Vk6Y2Xq67_2(.din(w_dff_B_JCp4qxlc8_2),.dout(w_dff_B_Vk6Y2Xq67_2),.clk(gclk));
	jdff dff_B_LCS3EVqP8_2(.din(w_dff_B_Vk6Y2Xq67_2),.dout(w_dff_B_LCS3EVqP8_2),.clk(gclk));
	jdff dff_B_5Mp9lluc6_2(.din(w_dff_B_LCS3EVqP8_2),.dout(w_dff_B_5Mp9lluc6_2),.clk(gclk));
	jdff dff_B_twsH7dNa2_2(.din(w_dff_B_5Mp9lluc6_2),.dout(w_dff_B_twsH7dNa2_2),.clk(gclk));
	jdff dff_B_EAR6JjCZ8_2(.din(w_dff_B_twsH7dNa2_2),.dout(w_dff_B_EAR6JjCZ8_2),.clk(gclk));
	jdff dff_B_7R9ngLxZ5_2(.din(w_dff_B_EAR6JjCZ8_2),.dout(w_dff_B_7R9ngLxZ5_2),.clk(gclk));
	jdff dff_B_hjvq3IXl3_2(.din(w_dff_B_7R9ngLxZ5_2),.dout(w_dff_B_hjvq3IXl3_2),.clk(gclk));
	jdff dff_B_oEOBnXxC6_2(.din(w_dff_B_hjvq3IXl3_2),.dout(w_dff_B_oEOBnXxC6_2),.clk(gclk));
	jdff dff_B_zRIZoJKA2_2(.din(w_dff_B_oEOBnXxC6_2),.dout(w_dff_B_zRIZoJKA2_2),.clk(gclk));
	jdff dff_B_opiGyJHv5_2(.din(w_dff_B_zRIZoJKA2_2),.dout(w_dff_B_opiGyJHv5_2),.clk(gclk));
	jdff dff_B_w8eQaxiw6_2(.din(w_dff_B_opiGyJHv5_2),.dout(w_dff_B_w8eQaxiw6_2),.clk(gclk));
	jdff dff_B_TyuHfqsA3_2(.din(w_dff_B_w8eQaxiw6_2),.dout(w_dff_B_TyuHfqsA3_2),.clk(gclk));
	jdff dff_B_VjKKWoOF8_2(.din(w_dff_B_TyuHfqsA3_2),.dout(w_dff_B_VjKKWoOF8_2),.clk(gclk));
	jdff dff_B_43rU9oyq8_2(.din(n1161),.dout(w_dff_B_43rU9oyq8_2),.clk(gclk));
	jdff dff_B_isMwcS1w1_1(.din(n1159),.dout(w_dff_B_isMwcS1w1_1),.clk(gclk));
	jdff dff_B_jqSPLVzL8_2(.din(n1054),.dout(w_dff_B_jqSPLVzL8_2),.clk(gclk));
	jdff dff_B_78yUqbDB2_2(.din(w_dff_B_jqSPLVzL8_2),.dout(w_dff_B_78yUqbDB2_2),.clk(gclk));
	jdff dff_B_1kAW4RxE4_2(.din(w_dff_B_78yUqbDB2_2),.dout(w_dff_B_1kAW4RxE4_2),.clk(gclk));
	jdff dff_B_Tf94WgGA3_2(.din(w_dff_B_1kAW4RxE4_2),.dout(w_dff_B_Tf94WgGA3_2),.clk(gclk));
	jdff dff_B_8bck2Qux5_2(.din(w_dff_B_Tf94WgGA3_2),.dout(w_dff_B_8bck2Qux5_2),.clk(gclk));
	jdff dff_B_tnlR70Fh9_2(.din(w_dff_B_8bck2Qux5_2),.dout(w_dff_B_tnlR70Fh9_2),.clk(gclk));
	jdff dff_B_1xSKL27U1_2(.din(w_dff_B_tnlR70Fh9_2),.dout(w_dff_B_1xSKL27U1_2),.clk(gclk));
	jdff dff_B_1N0rZ2cL1_2(.din(w_dff_B_1xSKL27U1_2),.dout(w_dff_B_1N0rZ2cL1_2),.clk(gclk));
	jdff dff_B_U15Kks6r0_2(.din(w_dff_B_1N0rZ2cL1_2),.dout(w_dff_B_U15Kks6r0_2),.clk(gclk));
	jdff dff_B_miGCYZ6K1_2(.din(w_dff_B_U15Kks6r0_2),.dout(w_dff_B_miGCYZ6K1_2),.clk(gclk));
	jdff dff_B_BYAOEYoV4_2(.din(w_dff_B_miGCYZ6K1_2),.dout(w_dff_B_BYAOEYoV4_2),.clk(gclk));
	jdff dff_B_VWLmRA2L7_2(.din(w_dff_B_BYAOEYoV4_2),.dout(w_dff_B_VWLmRA2L7_2),.clk(gclk));
	jdff dff_B_kBvRDchj5_2(.din(w_dff_B_VWLmRA2L7_2),.dout(w_dff_B_kBvRDchj5_2),.clk(gclk));
	jdff dff_B_JBfInPp25_2(.din(w_dff_B_kBvRDchj5_2),.dout(w_dff_B_JBfInPp25_2),.clk(gclk));
	jdff dff_B_fHX28qMm4_2(.din(w_dff_B_JBfInPp25_2),.dout(w_dff_B_fHX28qMm4_2),.clk(gclk));
	jdff dff_B_3hqzMtGP8_2(.din(w_dff_B_fHX28qMm4_2),.dout(w_dff_B_3hqzMtGP8_2),.clk(gclk));
	jdff dff_B_z7xVZdgB6_2(.din(w_dff_B_3hqzMtGP8_2),.dout(w_dff_B_z7xVZdgB6_2),.clk(gclk));
	jdff dff_B_p5BLpNmf8_2(.din(w_dff_B_z7xVZdgB6_2),.dout(w_dff_B_p5BLpNmf8_2),.clk(gclk));
	jdff dff_B_l5mYCSmb1_2(.din(w_dff_B_p5BLpNmf8_2),.dout(w_dff_B_l5mYCSmb1_2),.clk(gclk));
	jdff dff_B_oWCfsRT29_2(.din(w_dff_B_l5mYCSmb1_2),.dout(w_dff_B_oWCfsRT29_2),.clk(gclk));
	jdff dff_B_Eag7T3Go0_2(.din(w_dff_B_oWCfsRT29_2),.dout(w_dff_B_Eag7T3Go0_2),.clk(gclk));
	jdff dff_B_KGB44b8p5_2(.din(w_dff_B_Eag7T3Go0_2),.dout(w_dff_B_KGB44b8p5_2),.clk(gclk));
	jdff dff_B_7FiuL1fx8_2(.din(w_dff_B_KGB44b8p5_2),.dout(w_dff_B_7FiuL1fx8_2),.clk(gclk));
	jdff dff_B_tXmocK9L0_2(.din(w_dff_B_7FiuL1fx8_2),.dout(w_dff_B_tXmocK9L0_2),.clk(gclk));
	jdff dff_B_LYmXnR0D6_2(.din(w_dff_B_tXmocK9L0_2),.dout(w_dff_B_LYmXnR0D6_2),.clk(gclk));
	jdff dff_B_FUBlvQcc2_2(.din(w_dff_B_LYmXnR0D6_2),.dout(w_dff_B_FUBlvQcc2_2),.clk(gclk));
	jdff dff_B_Hh2EdLSE0_2(.din(w_dff_B_FUBlvQcc2_2),.dout(w_dff_B_Hh2EdLSE0_2),.clk(gclk));
	jdff dff_B_69xcZT3g0_2(.din(n1057),.dout(w_dff_B_69xcZT3g0_2),.clk(gclk));
	jdff dff_B_Bm80gPTd6_1(.din(n1055),.dout(w_dff_B_Bm80gPTd6_1),.clk(gclk));
	jdff dff_B_zM9DSR5m2_2(.din(n956),.dout(w_dff_B_zM9DSR5m2_2),.clk(gclk));
	jdff dff_B_otEsRPSG3_2(.din(w_dff_B_zM9DSR5m2_2),.dout(w_dff_B_otEsRPSG3_2),.clk(gclk));
	jdff dff_B_1v9u5R3z3_2(.din(w_dff_B_otEsRPSG3_2),.dout(w_dff_B_1v9u5R3z3_2),.clk(gclk));
	jdff dff_B_aZZ3vSDF5_2(.din(w_dff_B_1v9u5R3z3_2),.dout(w_dff_B_aZZ3vSDF5_2),.clk(gclk));
	jdff dff_B_5ociFwIS0_2(.din(w_dff_B_aZZ3vSDF5_2),.dout(w_dff_B_5ociFwIS0_2),.clk(gclk));
	jdff dff_B_GrkhuzJ79_2(.din(w_dff_B_5ociFwIS0_2),.dout(w_dff_B_GrkhuzJ79_2),.clk(gclk));
	jdff dff_B_2fvCIHTW9_2(.din(w_dff_B_GrkhuzJ79_2),.dout(w_dff_B_2fvCIHTW9_2),.clk(gclk));
	jdff dff_B_jSEuOTFR6_2(.din(w_dff_B_2fvCIHTW9_2),.dout(w_dff_B_jSEuOTFR6_2),.clk(gclk));
	jdff dff_B_fiqUj9wA1_2(.din(w_dff_B_jSEuOTFR6_2),.dout(w_dff_B_fiqUj9wA1_2),.clk(gclk));
	jdff dff_B_YDAYBLck8_2(.din(w_dff_B_fiqUj9wA1_2),.dout(w_dff_B_YDAYBLck8_2),.clk(gclk));
	jdff dff_B_psnTPa0Z9_2(.din(w_dff_B_YDAYBLck8_2),.dout(w_dff_B_psnTPa0Z9_2),.clk(gclk));
	jdff dff_B_yv0PcRP04_2(.din(w_dff_B_psnTPa0Z9_2),.dout(w_dff_B_yv0PcRP04_2),.clk(gclk));
	jdff dff_B_bt7SzeB15_2(.din(w_dff_B_yv0PcRP04_2),.dout(w_dff_B_bt7SzeB15_2),.clk(gclk));
	jdff dff_B_NrTWawmi1_2(.din(w_dff_B_bt7SzeB15_2),.dout(w_dff_B_NrTWawmi1_2),.clk(gclk));
	jdff dff_B_0ZyU1zqh9_2(.din(w_dff_B_NrTWawmi1_2),.dout(w_dff_B_0ZyU1zqh9_2),.clk(gclk));
	jdff dff_B_AH3T2WJe9_2(.din(w_dff_B_0ZyU1zqh9_2),.dout(w_dff_B_AH3T2WJe9_2),.clk(gclk));
	jdff dff_B_ZJXBQGRB7_2(.din(w_dff_B_AH3T2WJe9_2),.dout(w_dff_B_ZJXBQGRB7_2),.clk(gclk));
	jdff dff_B_mMXYx8nk0_2(.din(w_dff_B_ZJXBQGRB7_2),.dout(w_dff_B_mMXYx8nk0_2),.clk(gclk));
	jdff dff_B_Ih4QYTi56_2(.din(w_dff_B_mMXYx8nk0_2),.dout(w_dff_B_Ih4QYTi56_2),.clk(gclk));
	jdff dff_B_gSG37k7E7_2(.din(w_dff_B_Ih4QYTi56_2),.dout(w_dff_B_gSG37k7E7_2),.clk(gclk));
	jdff dff_B_TyIA3mho0_2(.din(w_dff_B_gSG37k7E7_2),.dout(w_dff_B_TyIA3mho0_2),.clk(gclk));
	jdff dff_B_eSBkTehi6_2(.din(w_dff_B_TyIA3mho0_2),.dout(w_dff_B_eSBkTehi6_2),.clk(gclk));
	jdff dff_B_sjTn3Y0B7_2(.din(w_dff_B_eSBkTehi6_2),.dout(w_dff_B_sjTn3Y0B7_2),.clk(gclk));
	jdff dff_B_0ZoEKReq9_2(.din(w_dff_B_sjTn3Y0B7_2),.dout(w_dff_B_0ZoEKReq9_2),.clk(gclk));
	jdff dff_B_W5g7uig16_1(.din(n957),.dout(w_dff_B_W5g7uig16_1),.clk(gclk));
	jdff dff_B_Iir1l9Dp0_2(.din(n851),.dout(w_dff_B_Iir1l9Dp0_2),.clk(gclk));
	jdff dff_B_HFdagoan1_2(.din(w_dff_B_Iir1l9Dp0_2),.dout(w_dff_B_HFdagoan1_2),.clk(gclk));
	jdff dff_B_cg6OqpNX8_2(.din(w_dff_B_HFdagoan1_2),.dout(w_dff_B_cg6OqpNX8_2),.clk(gclk));
	jdff dff_B_X8P0Gi0x9_2(.din(w_dff_B_cg6OqpNX8_2),.dout(w_dff_B_X8P0Gi0x9_2),.clk(gclk));
	jdff dff_B_ILuCj0TM5_2(.din(w_dff_B_X8P0Gi0x9_2),.dout(w_dff_B_ILuCj0TM5_2),.clk(gclk));
	jdff dff_B_MmafUwET9_2(.din(w_dff_B_ILuCj0TM5_2),.dout(w_dff_B_MmafUwET9_2),.clk(gclk));
	jdff dff_B_0DHi9rko1_2(.din(w_dff_B_MmafUwET9_2),.dout(w_dff_B_0DHi9rko1_2),.clk(gclk));
	jdff dff_B_qE3pPuZD4_2(.din(w_dff_B_0DHi9rko1_2),.dout(w_dff_B_qE3pPuZD4_2),.clk(gclk));
	jdff dff_B_HgOBbvJq6_2(.din(w_dff_B_qE3pPuZD4_2),.dout(w_dff_B_HgOBbvJq6_2),.clk(gclk));
	jdff dff_B_Xzay8MMW1_2(.din(w_dff_B_HgOBbvJq6_2),.dout(w_dff_B_Xzay8MMW1_2),.clk(gclk));
	jdff dff_B_ZadAQLYB2_2(.din(w_dff_B_Xzay8MMW1_2),.dout(w_dff_B_ZadAQLYB2_2),.clk(gclk));
	jdff dff_B_LNzFBwBl0_2(.din(w_dff_B_ZadAQLYB2_2),.dout(w_dff_B_LNzFBwBl0_2),.clk(gclk));
	jdff dff_B_jtqDpEpY8_2(.din(w_dff_B_LNzFBwBl0_2),.dout(w_dff_B_jtqDpEpY8_2),.clk(gclk));
	jdff dff_B_urQcLKTw6_2(.din(w_dff_B_jtqDpEpY8_2),.dout(w_dff_B_urQcLKTw6_2),.clk(gclk));
	jdff dff_B_4zTlFqWa8_2(.din(w_dff_B_urQcLKTw6_2),.dout(w_dff_B_4zTlFqWa8_2),.clk(gclk));
	jdff dff_B_makkpbhy1_2(.din(w_dff_B_4zTlFqWa8_2),.dout(w_dff_B_makkpbhy1_2),.clk(gclk));
	jdff dff_B_pSpKKRGM7_2(.din(w_dff_B_makkpbhy1_2),.dout(w_dff_B_pSpKKRGM7_2),.clk(gclk));
	jdff dff_B_TztNTQIm8_2(.din(w_dff_B_pSpKKRGM7_2),.dout(w_dff_B_TztNTQIm8_2),.clk(gclk));
	jdff dff_B_nQIo6htB5_2(.din(w_dff_B_TztNTQIm8_2),.dout(w_dff_B_nQIo6htB5_2),.clk(gclk));
	jdff dff_B_iKu78UdK2_2(.din(w_dff_B_nQIo6htB5_2),.dout(w_dff_B_iKu78UdK2_2),.clk(gclk));
	jdff dff_B_0JwzWpsh1_2(.din(w_dff_B_iKu78UdK2_2),.dout(w_dff_B_0JwzWpsh1_2),.clk(gclk));
	jdff dff_B_JClOxoUf1_2(.din(w_dff_B_0JwzWpsh1_2),.dout(w_dff_B_JClOxoUf1_2),.clk(gclk));
	jdff dff_B_xYzFwxws2_1(.din(n852),.dout(w_dff_B_xYzFwxws2_1),.clk(gclk));
	jdff dff_B_HTn8MndJ7_2(.din(n752),.dout(w_dff_B_HTn8MndJ7_2),.clk(gclk));
	jdff dff_B_GDrzHuKv3_2(.din(w_dff_B_HTn8MndJ7_2),.dout(w_dff_B_GDrzHuKv3_2),.clk(gclk));
	jdff dff_B_xfuaUkHC2_2(.din(w_dff_B_GDrzHuKv3_2),.dout(w_dff_B_xfuaUkHC2_2),.clk(gclk));
	jdff dff_B_ZgIRalUH6_2(.din(w_dff_B_xfuaUkHC2_2),.dout(w_dff_B_ZgIRalUH6_2),.clk(gclk));
	jdff dff_B_Zsz8LbIJ2_2(.din(w_dff_B_ZgIRalUH6_2),.dout(w_dff_B_Zsz8LbIJ2_2),.clk(gclk));
	jdff dff_B_BsRFxe4h0_2(.din(w_dff_B_Zsz8LbIJ2_2),.dout(w_dff_B_BsRFxe4h0_2),.clk(gclk));
	jdff dff_B_yySsxa9Q5_2(.din(w_dff_B_BsRFxe4h0_2),.dout(w_dff_B_yySsxa9Q5_2),.clk(gclk));
	jdff dff_B_AvCstIac7_2(.din(w_dff_B_yySsxa9Q5_2),.dout(w_dff_B_AvCstIac7_2),.clk(gclk));
	jdff dff_B_vVqxZcrC7_2(.din(w_dff_B_AvCstIac7_2),.dout(w_dff_B_vVqxZcrC7_2),.clk(gclk));
	jdff dff_B_4w0GsZBl6_2(.din(w_dff_B_vVqxZcrC7_2),.dout(w_dff_B_4w0GsZBl6_2),.clk(gclk));
	jdff dff_B_0DbbQjY77_2(.din(w_dff_B_4w0GsZBl6_2),.dout(w_dff_B_0DbbQjY77_2),.clk(gclk));
	jdff dff_B_WbYEeDaZ9_2(.din(w_dff_B_0DbbQjY77_2),.dout(w_dff_B_WbYEeDaZ9_2),.clk(gclk));
	jdff dff_B_WkaWoqEY2_2(.din(w_dff_B_WbYEeDaZ9_2),.dout(w_dff_B_WkaWoqEY2_2),.clk(gclk));
	jdff dff_B_EGX2etiJ9_2(.din(w_dff_B_WkaWoqEY2_2),.dout(w_dff_B_EGX2etiJ9_2),.clk(gclk));
	jdff dff_B_ogxpMXUR8_2(.din(w_dff_B_EGX2etiJ9_2),.dout(w_dff_B_ogxpMXUR8_2),.clk(gclk));
	jdff dff_B_uMQeDKnK0_2(.din(w_dff_B_ogxpMXUR8_2),.dout(w_dff_B_uMQeDKnK0_2),.clk(gclk));
	jdff dff_B_M4mJ7PxG7_2(.din(w_dff_B_uMQeDKnK0_2),.dout(w_dff_B_M4mJ7PxG7_2),.clk(gclk));
	jdff dff_B_Dlr1YPDj2_2(.din(w_dff_B_M4mJ7PxG7_2),.dout(w_dff_B_Dlr1YPDj2_2),.clk(gclk));
	jdff dff_B_NhRtzx3h1_2(.din(w_dff_B_Dlr1YPDj2_2),.dout(w_dff_B_NhRtzx3h1_2),.clk(gclk));
	jdff dff_B_G0y1hWVS6_2(.din(w_dff_B_NhRtzx3h1_2),.dout(w_dff_B_G0y1hWVS6_2),.clk(gclk));
	jdff dff_B_g5xYgFsp1_1(.din(n753),.dout(w_dff_B_g5xYgFsp1_1),.clk(gclk));
	jdff dff_B_oGO7mV1f8_2(.din(n659),.dout(w_dff_B_oGO7mV1f8_2),.clk(gclk));
	jdff dff_B_a05sQuiN5_2(.din(w_dff_B_oGO7mV1f8_2),.dout(w_dff_B_a05sQuiN5_2),.clk(gclk));
	jdff dff_B_3Zl9v8QY2_2(.din(w_dff_B_a05sQuiN5_2),.dout(w_dff_B_3Zl9v8QY2_2),.clk(gclk));
	jdff dff_B_ktCushNk5_2(.din(w_dff_B_3Zl9v8QY2_2),.dout(w_dff_B_ktCushNk5_2),.clk(gclk));
	jdff dff_B_92LUl3xV9_2(.din(w_dff_B_ktCushNk5_2),.dout(w_dff_B_92LUl3xV9_2),.clk(gclk));
	jdff dff_B_z54okmfN2_2(.din(w_dff_B_92LUl3xV9_2),.dout(w_dff_B_z54okmfN2_2),.clk(gclk));
	jdff dff_B_WmPwmEBH4_2(.din(w_dff_B_z54okmfN2_2),.dout(w_dff_B_WmPwmEBH4_2),.clk(gclk));
	jdff dff_B_2PPyRgBE5_2(.din(w_dff_B_WmPwmEBH4_2),.dout(w_dff_B_2PPyRgBE5_2),.clk(gclk));
	jdff dff_B_EWXT9pjb2_2(.din(w_dff_B_2PPyRgBE5_2),.dout(w_dff_B_EWXT9pjb2_2),.clk(gclk));
	jdff dff_B_Cd679bam3_2(.din(w_dff_B_EWXT9pjb2_2),.dout(w_dff_B_Cd679bam3_2),.clk(gclk));
	jdff dff_B_23lbCNkt2_2(.din(w_dff_B_Cd679bam3_2),.dout(w_dff_B_23lbCNkt2_2),.clk(gclk));
	jdff dff_B_FLalwGIO4_2(.din(w_dff_B_23lbCNkt2_2),.dout(w_dff_B_FLalwGIO4_2),.clk(gclk));
	jdff dff_B_8IgrJCwc7_2(.din(w_dff_B_FLalwGIO4_2),.dout(w_dff_B_8IgrJCwc7_2),.clk(gclk));
	jdff dff_B_EP1cTlPZ4_2(.din(w_dff_B_8IgrJCwc7_2),.dout(w_dff_B_EP1cTlPZ4_2),.clk(gclk));
	jdff dff_B_Q7txkeJv4_2(.din(w_dff_B_EP1cTlPZ4_2),.dout(w_dff_B_Q7txkeJv4_2),.clk(gclk));
	jdff dff_B_igt6yA2B5_2(.din(w_dff_B_Q7txkeJv4_2),.dout(w_dff_B_igt6yA2B5_2),.clk(gclk));
	jdff dff_B_Y11jGgSH6_2(.din(w_dff_B_igt6yA2B5_2),.dout(w_dff_B_Y11jGgSH6_2),.clk(gclk));
	jdff dff_B_VC4cduzu1_2(.din(w_dff_B_Y11jGgSH6_2),.dout(w_dff_B_VC4cduzu1_2),.clk(gclk));
	jdff dff_B_1cPflRMl6_1(.din(n660),.dout(w_dff_B_1cPflRMl6_1),.clk(gclk));
	jdff dff_B_lQuST4Wq9_2(.din(n573),.dout(w_dff_B_lQuST4Wq9_2),.clk(gclk));
	jdff dff_B_oD8ESpb73_2(.din(w_dff_B_lQuST4Wq9_2),.dout(w_dff_B_oD8ESpb73_2),.clk(gclk));
	jdff dff_B_ewdMYlzB0_2(.din(w_dff_B_oD8ESpb73_2),.dout(w_dff_B_ewdMYlzB0_2),.clk(gclk));
	jdff dff_B_QPcz9Fjk0_2(.din(w_dff_B_ewdMYlzB0_2),.dout(w_dff_B_QPcz9Fjk0_2),.clk(gclk));
	jdff dff_B_88gOg1RB2_2(.din(w_dff_B_QPcz9Fjk0_2),.dout(w_dff_B_88gOg1RB2_2),.clk(gclk));
	jdff dff_B_0byU5bLA9_2(.din(w_dff_B_88gOg1RB2_2),.dout(w_dff_B_0byU5bLA9_2),.clk(gclk));
	jdff dff_B_lyT8jWWI9_2(.din(w_dff_B_0byU5bLA9_2),.dout(w_dff_B_lyT8jWWI9_2),.clk(gclk));
	jdff dff_B_2LlqdzRq8_2(.din(w_dff_B_lyT8jWWI9_2),.dout(w_dff_B_2LlqdzRq8_2),.clk(gclk));
	jdff dff_B_1hXrFyqf1_2(.din(w_dff_B_2LlqdzRq8_2),.dout(w_dff_B_1hXrFyqf1_2),.clk(gclk));
	jdff dff_B_oC2zEpRx6_2(.din(w_dff_B_1hXrFyqf1_2),.dout(w_dff_B_oC2zEpRx6_2),.clk(gclk));
	jdff dff_B_AJV5VVpG4_2(.din(w_dff_B_oC2zEpRx6_2),.dout(w_dff_B_AJV5VVpG4_2),.clk(gclk));
	jdff dff_B_IauWHviK7_2(.din(w_dff_B_AJV5VVpG4_2),.dout(w_dff_B_IauWHviK7_2),.clk(gclk));
	jdff dff_B_6SioGfHX3_2(.din(w_dff_B_IauWHviK7_2),.dout(w_dff_B_6SioGfHX3_2),.clk(gclk));
	jdff dff_B_oPqhnOSV7_2(.din(w_dff_B_6SioGfHX3_2),.dout(w_dff_B_oPqhnOSV7_2),.clk(gclk));
	jdff dff_B_XnCFEuYz0_2(.din(w_dff_B_oPqhnOSV7_2),.dout(w_dff_B_XnCFEuYz0_2),.clk(gclk));
	jdff dff_B_RwsypYQB6_2(.din(w_dff_B_XnCFEuYz0_2),.dout(w_dff_B_RwsypYQB6_2),.clk(gclk));
	jdff dff_B_KAUL5l4Y9_1(.din(n574),.dout(w_dff_B_KAUL5l4Y9_1),.clk(gclk));
	jdff dff_B_4PnBuiIr8_2(.din(n494),.dout(w_dff_B_4PnBuiIr8_2),.clk(gclk));
	jdff dff_B_jjGp7l2O7_2(.din(w_dff_B_4PnBuiIr8_2),.dout(w_dff_B_jjGp7l2O7_2),.clk(gclk));
	jdff dff_B_gNAIgqb93_2(.din(w_dff_B_jjGp7l2O7_2),.dout(w_dff_B_gNAIgqb93_2),.clk(gclk));
	jdff dff_B_odIHAG0E6_2(.din(w_dff_B_gNAIgqb93_2),.dout(w_dff_B_odIHAG0E6_2),.clk(gclk));
	jdff dff_B_SgMjPHcc9_2(.din(w_dff_B_odIHAG0E6_2),.dout(w_dff_B_SgMjPHcc9_2),.clk(gclk));
	jdff dff_B_lPP0xdx58_2(.din(w_dff_B_SgMjPHcc9_2),.dout(w_dff_B_lPP0xdx58_2),.clk(gclk));
	jdff dff_B_WsBLMzPU7_2(.din(w_dff_B_lPP0xdx58_2),.dout(w_dff_B_WsBLMzPU7_2),.clk(gclk));
	jdff dff_B_PWmMLnaI0_2(.din(w_dff_B_WsBLMzPU7_2),.dout(w_dff_B_PWmMLnaI0_2),.clk(gclk));
	jdff dff_B_ekCqA8O74_2(.din(w_dff_B_PWmMLnaI0_2),.dout(w_dff_B_ekCqA8O74_2),.clk(gclk));
	jdff dff_B_atYf08Cx5_2(.din(w_dff_B_ekCqA8O74_2),.dout(w_dff_B_atYf08Cx5_2),.clk(gclk));
	jdff dff_B_0N2zsqDj5_2(.din(w_dff_B_atYf08Cx5_2),.dout(w_dff_B_0N2zsqDj5_2),.clk(gclk));
	jdff dff_B_MIiODms32_2(.din(w_dff_B_0N2zsqDj5_2),.dout(w_dff_B_MIiODms32_2),.clk(gclk));
	jdff dff_B_BvjHOT067_2(.din(w_dff_B_MIiODms32_2),.dout(w_dff_B_BvjHOT067_2),.clk(gclk));
	jdff dff_B_ioksKqhM3_2(.din(w_dff_B_BvjHOT067_2),.dout(w_dff_B_ioksKqhM3_2),.clk(gclk));
	jdff dff_B_DXjHtJBZ6_1(.din(n495),.dout(w_dff_B_DXjHtJBZ6_1),.clk(gclk));
	jdff dff_B_CFowmArr3_2(.din(n422),.dout(w_dff_B_CFowmArr3_2),.clk(gclk));
	jdff dff_B_wXFRrzH93_2(.din(w_dff_B_CFowmArr3_2),.dout(w_dff_B_wXFRrzH93_2),.clk(gclk));
	jdff dff_B_pCKaer9d2_2(.din(w_dff_B_wXFRrzH93_2),.dout(w_dff_B_pCKaer9d2_2),.clk(gclk));
	jdff dff_B_XWvV3Zr30_2(.din(w_dff_B_pCKaer9d2_2),.dout(w_dff_B_XWvV3Zr30_2),.clk(gclk));
	jdff dff_B_kQNePC2n0_2(.din(w_dff_B_XWvV3Zr30_2),.dout(w_dff_B_kQNePC2n0_2),.clk(gclk));
	jdff dff_B_nUvdRr6R0_2(.din(w_dff_B_kQNePC2n0_2),.dout(w_dff_B_nUvdRr6R0_2),.clk(gclk));
	jdff dff_B_TYFYL5hm1_2(.din(w_dff_B_nUvdRr6R0_2),.dout(w_dff_B_TYFYL5hm1_2),.clk(gclk));
	jdff dff_B_9dBaEDsj5_2(.din(w_dff_B_TYFYL5hm1_2),.dout(w_dff_B_9dBaEDsj5_2),.clk(gclk));
	jdff dff_B_XOGFjnUO3_2(.din(w_dff_B_9dBaEDsj5_2),.dout(w_dff_B_XOGFjnUO3_2),.clk(gclk));
	jdff dff_B_zWQw8quC7_2(.din(w_dff_B_XOGFjnUO3_2),.dout(w_dff_B_zWQw8quC7_2),.clk(gclk));
	jdff dff_B_nQoFuduk2_2(.din(w_dff_B_zWQw8quC7_2),.dout(w_dff_B_nQoFuduk2_2),.clk(gclk));
	jdff dff_B_Gpq1DOjM2_2(.din(w_dff_B_nQoFuduk2_2),.dout(w_dff_B_Gpq1DOjM2_2),.clk(gclk));
	jdff dff_B_yDwcpi3L2_1(.din(n423),.dout(w_dff_B_yDwcpi3L2_1),.clk(gclk));
	jdff dff_B_O7eGrU9d5_2(.din(n358),.dout(w_dff_B_O7eGrU9d5_2),.clk(gclk));
	jdff dff_B_FCYgnG4M9_2(.din(w_dff_B_O7eGrU9d5_2),.dout(w_dff_B_FCYgnG4M9_2),.clk(gclk));
	jdff dff_B_HmrHlPGp3_2(.din(w_dff_B_FCYgnG4M9_2),.dout(w_dff_B_HmrHlPGp3_2),.clk(gclk));
	jdff dff_B_IJqciMO44_2(.din(w_dff_B_HmrHlPGp3_2),.dout(w_dff_B_IJqciMO44_2),.clk(gclk));
	jdff dff_B_F47BQwFu2_2(.din(w_dff_B_IJqciMO44_2),.dout(w_dff_B_F47BQwFu2_2),.clk(gclk));
	jdff dff_B_22mCeoIk7_2(.din(w_dff_B_F47BQwFu2_2),.dout(w_dff_B_22mCeoIk7_2),.clk(gclk));
	jdff dff_B_va4zvVCo2_2(.din(w_dff_B_22mCeoIk7_2),.dout(w_dff_B_va4zvVCo2_2),.clk(gclk));
	jdff dff_B_x8aip9lM7_2(.din(w_dff_B_va4zvVCo2_2),.dout(w_dff_B_x8aip9lM7_2),.clk(gclk));
	jdff dff_B_rdkqiocP9_2(.din(w_dff_B_x8aip9lM7_2),.dout(w_dff_B_rdkqiocP9_2),.clk(gclk));
	jdff dff_B_ewWnwWek2_2(.din(w_dff_B_rdkqiocP9_2),.dout(w_dff_B_ewWnwWek2_2),.clk(gclk));
	jdff dff_B_Vv4HgKB73_1(.din(n359),.dout(w_dff_B_Vv4HgKB73_1),.clk(gclk));
	jdff dff_B_VYxybrD26_2(.din(n300),.dout(w_dff_B_VYxybrD26_2),.clk(gclk));
	jdff dff_B_5ZipRCYh4_2(.din(w_dff_B_VYxybrD26_2),.dout(w_dff_B_5ZipRCYh4_2),.clk(gclk));
	jdff dff_B_E1fKmDBK1_2(.din(w_dff_B_5ZipRCYh4_2),.dout(w_dff_B_E1fKmDBK1_2),.clk(gclk));
	jdff dff_B_Q8I7aWfH8_2(.din(w_dff_B_E1fKmDBK1_2),.dout(w_dff_B_Q8I7aWfH8_2),.clk(gclk));
	jdff dff_B_itzwMyMP3_2(.din(w_dff_B_Q8I7aWfH8_2),.dout(w_dff_B_itzwMyMP3_2),.clk(gclk));
	jdff dff_B_7vfeekxt9_2(.din(w_dff_B_itzwMyMP3_2),.dout(w_dff_B_7vfeekxt9_2),.clk(gclk));
	jdff dff_B_gdRa8BAw4_2(.din(w_dff_B_7vfeekxt9_2),.dout(w_dff_B_gdRa8BAw4_2),.clk(gclk));
	jdff dff_B_n7O6EScb1_2(.din(w_dff_B_gdRa8BAw4_2),.dout(w_dff_B_n7O6EScb1_2),.clk(gclk));
	jdff dff_B_aRfMzHED9_1(.din(n301),.dout(w_dff_B_aRfMzHED9_1),.clk(gclk));
	jdff dff_B_u6LFQJzG1_2(.din(n249),.dout(w_dff_B_u6LFQJzG1_2),.clk(gclk));
	jdff dff_B_pkp0MDj07_2(.din(w_dff_B_u6LFQJzG1_2),.dout(w_dff_B_pkp0MDj07_2),.clk(gclk));
	jdff dff_B_Qo2Z6x0A8_2(.din(w_dff_B_pkp0MDj07_2),.dout(w_dff_B_Qo2Z6x0A8_2),.clk(gclk));
	jdff dff_B_OLdugPB46_2(.din(w_dff_B_Qo2Z6x0A8_2),.dout(w_dff_B_OLdugPB46_2),.clk(gclk));
	jdff dff_B_3y1bZXqQ4_2(.din(w_dff_B_OLdugPB46_2),.dout(w_dff_B_3y1bZXqQ4_2),.clk(gclk));
	jdff dff_B_TQjrYt633_2(.din(w_dff_B_3y1bZXqQ4_2),.dout(w_dff_B_TQjrYt633_2),.clk(gclk));
	jdff dff_B_TCPyOj6B9_2(.din(n252),.dout(w_dff_B_TCPyOj6B9_2),.clk(gclk));
	jdff dff_B_lXlV1jzs3_1(.din(n250),.dout(w_dff_B_lXlV1jzs3_1),.clk(gclk));
	jdff dff_B_uPKK8ESG8_0(.din(n214),.dout(w_dff_B_uPKK8ESG8_0),.clk(gclk));
	jdff dff_B_NenG3xHE2_2(.din(n206),.dout(w_dff_B_NenG3xHE2_2),.clk(gclk));
	jdff dff_B_hBRVaz9W2_2(.din(w_dff_B_NenG3xHE2_2),.dout(w_dff_B_hBRVaz9W2_2),.clk(gclk));
	jdff dff_B_PZOVoV967_2(.din(w_dff_B_hBRVaz9W2_2),.dout(w_dff_B_PZOVoV967_2),.clk(gclk));
	jdff dff_B_iAZ0Lkdv4_1(.din(n208),.dout(w_dff_B_iAZ0Lkdv4_1),.clk(gclk));
	jdff dff_B_csL5jpSV9_1(.din(w_dff_B_iAZ0Lkdv4_1),.dout(w_dff_B_csL5jpSV9_1),.clk(gclk));
	jdff dff_A_9f3FoyNE9_0(.dout(w_n210_1[0]),.din(w_dff_A_9f3FoyNE9_0),.clk(gclk));
	jdff dff_A_WYSV1EYY1_0(.dout(w_n169_0[0]),.din(w_dff_A_WYSV1EYY1_0),.clk(gclk));
	jdff dff_A_89r2owrF7_0(.dout(w_dff_A_WYSV1EYY1_0),.din(w_dff_A_89r2owrF7_0),.clk(gclk));
	jdff dff_A_bs6TpDgl8_1(.dout(w_n169_0[1]),.din(w_dff_A_bs6TpDgl8_1),.clk(gclk));
	jdff dff_B_2c2Vq3eT1_2(.din(n1420),.dout(w_dff_B_2c2Vq3eT1_2),.clk(gclk));
	jdff dff_B_TJfsuamC7_2(.din(w_dff_B_2c2Vq3eT1_2),.dout(w_dff_B_TJfsuamC7_2),.clk(gclk));
	jdff dff_B_c0gKDITm0_1(.din(n1418),.dout(w_dff_B_c0gKDITm0_1),.clk(gclk));
	jdff dff_B_0Kt4G5Mp8_2(.din(n1338),.dout(w_dff_B_0Kt4G5Mp8_2),.clk(gclk));
	jdff dff_B_seHp4O5c8_2(.din(w_dff_B_0Kt4G5Mp8_2),.dout(w_dff_B_seHp4O5c8_2),.clk(gclk));
	jdff dff_B_xVWXescX2_2(.din(w_dff_B_seHp4O5c8_2),.dout(w_dff_B_xVWXescX2_2),.clk(gclk));
	jdff dff_B_WK1KZI2k5_2(.din(w_dff_B_xVWXescX2_2),.dout(w_dff_B_WK1KZI2k5_2),.clk(gclk));
	jdff dff_B_NTSDQlkA8_2(.din(w_dff_B_WK1KZI2k5_2),.dout(w_dff_B_NTSDQlkA8_2),.clk(gclk));
	jdff dff_B_JeYbGqYJ3_2(.din(w_dff_B_NTSDQlkA8_2),.dout(w_dff_B_JeYbGqYJ3_2),.clk(gclk));
	jdff dff_B_gII3xVBw6_2(.din(w_dff_B_JeYbGqYJ3_2),.dout(w_dff_B_gII3xVBw6_2),.clk(gclk));
	jdff dff_B_nYqfiiSP0_2(.din(w_dff_B_gII3xVBw6_2),.dout(w_dff_B_nYqfiiSP0_2),.clk(gclk));
	jdff dff_B_KcmjyqDt9_2(.din(w_dff_B_nYqfiiSP0_2),.dout(w_dff_B_KcmjyqDt9_2),.clk(gclk));
	jdff dff_B_xPtwnFHQ8_2(.din(w_dff_B_KcmjyqDt9_2),.dout(w_dff_B_xPtwnFHQ8_2),.clk(gclk));
	jdff dff_B_10X5kgUQ6_2(.din(w_dff_B_xPtwnFHQ8_2),.dout(w_dff_B_10X5kgUQ6_2),.clk(gclk));
	jdff dff_B_JTzkY5tB8_2(.din(w_dff_B_10X5kgUQ6_2),.dout(w_dff_B_JTzkY5tB8_2),.clk(gclk));
	jdff dff_B_JRa8KJyg3_2(.din(w_dff_B_JTzkY5tB8_2),.dout(w_dff_B_JRa8KJyg3_2),.clk(gclk));
	jdff dff_B_2YUPKL386_2(.din(w_dff_B_JRa8KJyg3_2),.dout(w_dff_B_2YUPKL386_2),.clk(gclk));
	jdff dff_B_FEcWnkgH6_2(.din(w_dff_B_2YUPKL386_2),.dout(w_dff_B_FEcWnkgH6_2),.clk(gclk));
	jdff dff_B_E4MhIlBi4_2(.din(w_dff_B_FEcWnkgH6_2),.dout(w_dff_B_E4MhIlBi4_2),.clk(gclk));
	jdff dff_B_WxxUFk6Y8_2(.din(w_dff_B_E4MhIlBi4_2),.dout(w_dff_B_WxxUFk6Y8_2),.clk(gclk));
	jdff dff_B_AzEzZdB57_2(.din(w_dff_B_WxxUFk6Y8_2),.dout(w_dff_B_AzEzZdB57_2),.clk(gclk));
	jdff dff_B_SajIirry9_2(.din(w_dff_B_AzEzZdB57_2),.dout(w_dff_B_SajIirry9_2),.clk(gclk));
	jdff dff_B_VOyzUhNY4_2(.din(w_dff_B_SajIirry9_2),.dout(w_dff_B_VOyzUhNY4_2),.clk(gclk));
	jdff dff_B_E296GWDi4_2(.din(w_dff_B_VOyzUhNY4_2),.dout(w_dff_B_E296GWDi4_2),.clk(gclk));
	jdff dff_B_9dSD4YXs7_2(.din(w_dff_B_E296GWDi4_2),.dout(w_dff_B_9dSD4YXs7_2),.clk(gclk));
	jdff dff_B_2dxaVkZi9_2(.din(w_dff_B_9dSD4YXs7_2),.dout(w_dff_B_2dxaVkZi9_2),.clk(gclk));
	jdff dff_B_8zqNlNcM7_2(.din(w_dff_B_2dxaVkZi9_2),.dout(w_dff_B_8zqNlNcM7_2),.clk(gclk));
	jdff dff_B_ZGfGp6El6_2(.din(w_dff_B_8zqNlNcM7_2),.dout(w_dff_B_ZGfGp6El6_2),.clk(gclk));
	jdff dff_B_0bXkMjxX5_2(.din(w_dff_B_ZGfGp6El6_2),.dout(w_dff_B_0bXkMjxX5_2),.clk(gclk));
	jdff dff_B_Zr5J63or4_2(.din(w_dff_B_0bXkMjxX5_2),.dout(w_dff_B_Zr5J63or4_2),.clk(gclk));
	jdff dff_B_Mn77ED753_2(.din(w_dff_B_Zr5J63or4_2),.dout(w_dff_B_Mn77ED753_2),.clk(gclk));
	jdff dff_B_s20hIMS20_2(.din(w_dff_B_Mn77ED753_2),.dout(w_dff_B_s20hIMS20_2),.clk(gclk));
	jdff dff_B_0WtfogX21_2(.din(w_dff_B_s20hIMS20_2),.dout(w_dff_B_0WtfogX21_2),.clk(gclk));
	jdff dff_B_yP1yH5Mq7_2(.din(w_dff_B_0WtfogX21_2),.dout(w_dff_B_yP1yH5Mq7_2),.clk(gclk));
	jdff dff_B_Wi9A6BGr9_2(.din(w_dff_B_yP1yH5Mq7_2),.dout(w_dff_B_Wi9A6BGr9_2),.clk(gclk));
	jdff dff_B_rMaPfSgc1_2(.din(w_dff_B_Wi9A6BGr9_2),.dout(w_dff_B_rMaPfSgc1_2),.clk(gclk));
	jdff dff_B_NPdh8szz8_2(.din(w_dff_B_rMaPfSgc1_2),.dout(w_dff_B_NPdh8szz8_2),.clk(gclk));
	jdff dff_B_4WINysLX4_2(.din(w_dff_B_NPdh8szz8_2),.dout(w_dff_B_4WINysLX4_2),.clk(gclk));
	jdff dff_B_L9bSzvvj0_2(.din(w_dff_B_4WINysLX4_2),.dout(w_dff_B_L9bSzvvj0_2),.clk(gclk));
	jdff dff_B_ZuB48PZT2_1(.din(n1416),.dout(w_dff_B_ZuB48PZT2_1),.clk(gclk));
	jdff dff_A_1gzZBzEp4_1(.dout(w_n1341_0[1]),.din(w_dff_A_1gzZBzEp4_1),.clk(gclk));
	jdff dff_B_PgiGbC5X8_1(.din(n1339),.dout(w_dff_B_PgiGbC5X8_1),.clk(gclk));
	jdff dff_B_mxJtfWY44_2(.din(n1253),.dout(w_dff_B_mxJtfWY44_2),.clk(gclk));
	jdff dff_B_Sc34o0UJ5_2(.din(w_dff_B_mxJtfWY44_2),.dout(w_dff_B_Sc34o0UJ5_2),.clk(gclk));
	jdff dff_B_ra8v41Jb7_2(.din(w_dff_B_Sc34o0UJ5_2),.dout(w_dff_B_ra8v41Jb7_2),.clk(gclk));
	jdff dff_B_9C6VkztW6_2(.din(w_dff_B_ra8v41Jb7_2),.dout(w_dff_B_9C6VkztW6_2),.clk(gclk));
	jdff dff_B_wGCewpp48_2(.din(w_dff_B_9C6VkztW6_2),.dout(w_dff_B_wGCewpp48_2),.clk(gclk));
	jdff dff_B_ZUiWFomF2_2(.din(w_dff_B_wGCewpp48_2),.dout(w_dff_B_ZUiWFomF2_2),.clk(gclk));
	jdff dff_B_iZjeqE6k9_2(.din(w_dff_B_ZUiWFomF2_2),.dout(w_dff_B_iZjeqE6k9_2),.clk(gclk));
	jdff dff_B_7u8kzptq9_2(.din(w_dff_B_iZjeqE6k9_2),.dout(w_dff_B_7u8kzptq9_2),.clk(gclk));
	jdff dff_B_s4PXG8wY4_2(.din(w_dff_B_7u8kzptq9_2),.dout(w_dff_B_s4PXG8wY4_2),.clk(gclk));
	jdff dff_B_UCp7faNg3_2(.din(w_dff_B_s4PXG8wY4_2),.dout(w_dff_B_UCp7faNg3_2),.clk(gclk));
	jdff dff_B_Flm8jeW13_2(.din(w_dff_B_UCp7faNg3_2),.dout(w_dff_B_Flm8jeW13_2),.clk(gclk));
	jdff dff_B_gNCv9Isw2_2(.din(w_dff_B_Flm8jeW13_2),.dout(w_dff_B_gNCv9Isw2_2),.clk(gclk));
	jdff dff_B_l2MS1AxN4_2(.din(w_dff_B_gNCv9Isw2_2),.dout(w_dff_B_l2MS1AxN4_2),.clk(gclk));
	jdff dff_B_wy9gGi1J2_2(.din(w_dff_B_l2MS1AxN4_2),.dout(w_dff_B_wy9gGi1J2_2),.clk(gclk));
	jdff dff_B_MIvxTpkS4_2(.din(w_dff_B_wy9gGi1J2_2),.dout(w_dff_B_MIvxTpkS4_2),.clk(gclk));
	jdff dff_B_y2qnU9p77_2(.din(w_dff_B_MIvxTpkS4_2),.dout(w_dff_B_y2qnU9p77_2),.clk(gclk));
	jdff dff_B_ONpLwPjA6_2(.din(w_dff_B_y2qnU9p77_2),.dout(w_dff_B_ONpLwPjA6_2),.clk(gclk));
	jdff dff_B_ixQXjcEW6_2(.din(w_dff_B_ONpLwPjA6_2),.dout(w_dff_B_ixQXjcEW6_2),.clk(gclk));
	jdff dff_B_yReINQyO8_2(.din(w_dff_B_ixQXjcEW6_2),.dout(w_dff_B_yReINQyO8_2),.clk(gclk));
	jdff dff_B_6gwlQc8T7_2(.din(w_dff_B_yReINQyO8_2),.dout(w_dff_B_6gwlQc8T7_2),.clk(gclk));
	jdff dff_B_qP3ZeTuv7_2(.din(w_dff_B_6gwlQc8T7_2),.dout(w_dff_B_qP3ZeTuv7_2),.clk(gclk));
	jdff dff_B_AWwznU641_2(.din(w_dff_B_qP3ZeTuv7_2),.dout(w_dff_B_AWwznU641_2),.clk(gclk));
	jdff dff_B_HFhs9QCc4_2(.din(w_dff_B_AWwznU641_2),.dout(w_dff_B_HFhs9QCc4_2),.clk(gclk));
	jdff dff_B_6GAkWeor2_2(.din(w_dff_B_HFhs9QCc4_2),.dout(w_dff_B_6GAkWeor2_2),.clk(gclk));
	jdff dff_B_szGhqEO27_2(.din(w_dff_B_6GAkWeor2_2),.dout(w_dff_B_szGhqEO27_2),.clk(gclk));
	jdff dff_B_VnwQJJHW4_2(.din(w_dff_B_szGhqEO27_2),.dout(w_dff_B_VnwQJJHW4_2),.clk(gclk));
	jdff dff_B_Yyt009D82_2(.din(w_dff_B_VnwQJJHW4_2),.dout(w_dff_B_Yyt009D82_2),.clk(gclk));
	jdff dff_B_u4StBFgl2_2(.din(w_dff_B_Yyt009D82_2),.dout(w_dff_B_u4StBFgl2_2),.clk(gclk));
	jdff dff_B_qY5CoyaW7_2(.din(w_dff_B_u4StBFgl2_2),.dout(w_dff_B_qY5CoyaW7_2),.clk(gclk));
	jdff dff_B_5XkrnHgD9_2(.din(w_dff_B_qY5CoyaW7_2),.dout(w_dff_B_5XkrnHgD9_2),.clk(gclk));
	jdff dff_B_IQs7OLLp0_2(.din(w_dff_B_5XkrnHgD9_2),.dout(w_dff_B_IQs7OLLp0_2),.clk(gclk));
	jdff dff_B_UP6lgHQk0_2(.din(n1256),.dout(w_dff_B_UP6lgHQk0_2),.clk(gclk));
	jdff dff_B_Jm9tIshv4_1(.din(n1254),.dout(w_dff_B_Jm9tIshv4_1),.clk(gclk));
	jdff dff_B_cDeRRrvT6_2(.din(n1163),.dout(w_dff_B_cDeRRrvT6_2),.clk(gclk));
	jdff dff_B_beFV1w8m4_2(.din(w_dff_B_cDeRRrvT6_2),.dout(w_dff_B_beFV1w8m4_2),.clk(gclk));
	jdff dff_B_jDNMgaUX7_2(.din(w_dff_B_beFV1w8m4_2),.dout(w_dff_B_jDNMgaUX7_2),.clk(gclk));
	jdff dff_B_QA2I0oNs9_2(.din(w_dff_B_jDNMgaUX7_2),.dout(w_dff_B_QA2I0oNs9_2),.clk(gclk));
	jdff dff_B_3v3pc9j28_2(.din(w_dff_B_QA2I0oNs9_2),.dout(w_dff_B_3v3pc9j28_2),.clk(gclk));
	jdff dff_B_luIh8VKD0_2(.din(w_dff_B_3v3pc9j28_2),.dout(w_dff_B_luIh8VKD0_2),.clk(gclk));
	jdff dff_B_WxNTYIEB8_2(.din(w_dff_B_luIh8VKD0_2),.dout(w_dff_B_WxNTYIEB8_2),.clk(gclk));
	jdff dff_B_Qj1EpNWE3_2(.din(w_dff_B_WxNTYIEB8_2),.dout(w_dff_B_Qj1EpNWE3_2),.clk(gclk));
	jdff dff_B_ZDD1f9eW5_2(.din(w_dff_B_Qj1EpNWE3_2),.dout(w_dff_B_ZDD1f9eW5_2),.clk(gclk));
	jdff dff_B_NlsUxI5B0_2(.din(w_dff_B_ZDD1f9eW5_2),.dout(w_dff_B_NlsUxI5B0_2),.clk(gclk));
	jdff dff_B_nqMpzWkn8_2(.din(w_dff_B_NlsUxI5B0_2),.dout(w_dff_B_nqMpzWkn8_2),.clk(gclk));
	jdff dff_B_f8ji0yuA5_2(.din(w_dff_B_nqMpzWkn8_2),.dout(w_dff_B_f8ji0yuA5_2),.clk(gclk));
	jdff dff_B_8hoDUfZT0_2(.din(w_dff_B_f8ji0yuA5_2),.dout(w_dff_B_8hoDUfZT0_2),.clk(gclk));
	jdff dff_B_29rJ4ON59_2(.din(w_dff_B_8hoDUfZT0_2),.dout(w_dff_B_29rJ4ON59_2),.clk(gclk));
	jdff dff_B_hr2CLswT9_2(.din(w_dff_B_29rJ4ON59_2),.dout(w_dff_B_hr2CLswT9_2),.clk(gclk));
	jdff dff_B_mYk1Dwt93_2(.din(w_dff_B_hr2CLswT9_2),.dout(w_dff_B_mYk1Dwt93_2),.clk(gclk));
	jdff dff_B_VeL6enjW6_2(.din(w_dff_B_mYk1Dwt93_2),.dout(w_dff_B_VeL6enjW6_2),.clk(gclk));
	jdff dff_B_ImBfs6A44_2(.din(w_dff_B_VeL6enjW6_2),.dout(w_dff_B_ImBfs6A44_2),.clk(gclk));
	jdff dff_B_g1M8Pnz44_2(.din(w_dff_B_ImBfs6A44_2),.dout(w_dff_B_g1M8Pnz44_2),.clk(gclk));
	jdff dff_B_oAJ0WtWL1_2(.din(w_dff_B_g1M8Pnz44_2),.dout(w_dff_B_oAJ0WtWL1_2),.clk(gclk));
	jdff dff_B_Wk6iza651_2(.din(w_dff_B_oAJ0WtWL1_2),.dout(w_dff_B_Wk6iza651_2),.clk(gclk));
	jdff dff_B_HWLxt7d93_2(.din(w_dff_B_Wk6iza651_2),.dout(w_dff_B_HWLxt7d93_2),.clk(gclk));
	jdff dff_B_6gzuIKjc0_2(.din(w_dff_B_HWLxt7d93_2),.dout(w_dff_B_6gzuIKjc0_2),.clk(gclk));
	jdff dff_B_ruKjRQyW3_2(.din(w_dff_B_6gzuIKjc0_2),.dout(w_dff_B_ruKjRQyW3_2),.clk(gclk));
	jdff dff_B_kiwq5H8R5_2(.din(w_dff_B_ruKjRQyW3_2),.dout(w_dff_B_kiwq5H8R5_2),.clk(gclk));
	jdff dff_B_RSneklzm8_2(.din(w_dff_B_kiwq5H8R5_2),.dout(w_dff_B_RSneklzm8_2),.clk(gclk));
	jdff dff_B_PIQ4bFKM0_2(.din(w_dff_B_RSneklzm8_2),.dout(w_dff_B_PIQ4bFKM0_2),.clk(gclk));
	jdff dff_B_0gddxcGe8_2(.din(w_dff_B_PIQ4bFKM0_2),.dout(w_dff_B_0gddxcGe8_2),.clk(gclk));
	jdff dff_B_NZTEQUB73_2(.din(n1166),.dout(w_dff_B_NZTEQUB73_2),.clk(gclk));
	jdff dff_B_YVApPPrf4_1(.din(n1164),.dout(w_dff_B_YVApPPrf4_1),.clk(gclk));
	jdff dff_B_u9c3TRX55_2(.din(n1059),.dout(w_dff_B_u9c3TRX55_2),.clk(gclk));
	jdff dff_B_x7z4HUUf8_2(.din(w_dff_B_u9c3TRX55_2),.dout(w_dff_B_x7z4HUUf8_2),.clk(gclk));
	jdff dff_B_PHOpvzVV7_2(.din(w_dff_B_x7z4HUUf8_2),.dout(w_dff_B_PHOpvzVV7_2),.clk(gclk));
	jdff dff_B_BtrFSV5h5_2(.din(w_dff_B_PHOpvzVV7_2),.dout(w_dff_B_BtrFSV5h5_2),.clk(gclk));
	jdff dff_B_cMnJIbxr2_2(.din(w_dff_B_BtrFSV5h5_2),.dout(w_dff_B_cMnJIbxr2_2),.clk(gclk));
	jdff dff_B_vtyohZyJ7_2(.din(w_dff_B_cMnJIbxr2_2),.dout(w_dff_B_vtyohZyJ7_2),.clk(gclk));
	jdff dff_B_Xn3H3yZb6_2(.din(w_dff_B_vtyohZyJ7_2),.dout(w_dff_B_Xn3H3yZb6_2),.clk(gclk));
	jdff dff_B_lU3I9ZbZ9_2(.din(w_dff_B_Xn3H3yZb6_2),.dout(w_dff_B_lU3I9ZbZ9_2),.clk(gclk));
	jdff dff_B_A0LUHoC71_2(.din(w_dff_B_lU3I9ZbZ9_2),.dout(w_dff_B_A0LUHoC71_2),.clk(gclk));
	jdff dff_B_YIAtZzM50_2(.din(w_dff_B_A0LUHoC71_2),.dout(w_dff_B_YIAtZzM50_2),.clk(gclk));
	jdff dff_B_VnqxHIum3_2(.din(w_dff_B_YIAtZzM50_2),.dout(w_dff_B_VnqxHIum3_2),.clk(gclk));
	jdff dff_B_oFXFmMYU7_2(.din(w_dff_B_VnqxHIum3_2),.dout(w_dff_B_oFXFmMYU7_2),.clk(gclk));
	jdff dff_B_oh906Dl82_2(.din(w_dff_B_oFXFmMYU7_2),.dout(w_dff_B_oh906Dl82_2),.clk(gclk));
	jdff dff_B_hG0zkLKC8_2(.din(w_dff_B_oh906Dl82_2),.dout(w_dff_B_hG0zkLKC8_2),.clk(gclk));
	jdff dff_B_1Ws0COUy6_2(.din(w_dff_B_hG0zkLKC8_2),.dout(w_dff_B_1Ws0COUy6_2),.clk(gclk));
	jdff dff_B_9UBkVgE06_2(.din(w_dff_B_1Ws0COUy6_2),.dout(w_dff_B_9UBkVgE06_2),.clk(gclk));
	jdff dff_B_e9cYIyqH7_2(.din(w_dff_B_9UBkVgE06_2),.dout(w_dff_B_e9cYIyqH7_2),.clk(gclk));
	jdff dff_B_iJOGgfpt3_2(.din(w_dff_B_e9cYIyqH7_2),.dout(w_dff_B_iJOGgfpt3_2),.clk(gclk));
	jdff dff_B_6JW7yPFx5_2(.din(w_dff_B_iJOGgfpt3_2),.dout(w_dff_B_6JW7yPFx5_2),.clk(gclk));
	jdff dff_B_fXXlRTTR1_2(.din(w_dff_B_6JW7yPFx5_2),.dout(w_dff_B_fXXlRTTR1_2),.clk(gclk));
	jdff dff_B_1nQQUPSi4_2(.din(w_dff_B_fXXlRTTR1_2),.dout(w_dff_B_1nQQUPSi4_2),.clk(gclk));
	jdff dff_B_GGatLbCo3_2(.din(w_dff_B_1nQQUPSi4_2),.dout(w_dff_B_GGatLbCo3_2),.clk(gclk));
	jdff dff_B_on73QUej8_2(.din(w_dff_B_GGatLbCo3_2),.dout(w_dff_B_on73QUej8_2),.clk(gclk));
	jdff dff_B_fXaeBC208_2(.din(w_dff_B_on73QUej8_2),.dout(w_dff_B_fXaeBC208_2),.clk(gclk));
	jdff dff_B_3wbRcmS09_2(.din(w_dff_B_fXaeBC208_2),.dout(w_dff_B_3wbRcmS09_2),.clk(gclk));
	jdff dff_B_ifC4YSHr9_2(.din(n1062),.dout(w_dff_B_ifC4YSHr9_2),.clk(gclk));
	jdff dff_B_V46Xsi6b9_1(.din(n1060),.dout(w_dff_B_V46Xsi6b9_1),.clk(gclk));
	jdff dff_B_hjCW9IC32_2(.din(n961),.dout(w_dff_B_hjCW9IC32_2),.clk(gclk));
	jdff dff_B_sjol2ITj3_2(.din(w_dff_B_hjCW9IC32_2),.dout(w_dff_B_sjol2ITj3_2),.clk(gclk));
	jdff dff_B_5LxvmuZQ6_2(.din(w_dff_B_sjol2ITj3_2),.dout(w_dff_B_5LxvmuZQ6_2),.clk(gclk));
	jdff dff_B_Vtq2Wt5F8_2(.din(w_dff_B_5LxvmuZQ6_2),.dout(w_dff_B_Vtq2Wt5F8_2),.clk(gclk));
	jdff dff_B_lJPvG3pD4_2(.din(w_dff_B_Vtq2Wt5F8_2),.dout(w_dff_B_lJPvG3pD4_2),.clk(gclk));
	jdff dff_B_PHTJ7ki73_2(.din(w_dff_B_lJPvG3pD4_2),.dout(w_dff_B_PHTJ7ki73_2),.clk(gclk));
	jdff dff_B_g98Uk9ux8_2(.din(w_dff_B_PHTJ7ki73_2),.dout(w_dff_B_g98Uk9ux8_2),.clk(gclk));
	jdff dff_B_pu99VB340_2(.din(w_dff_B_g98Uk9ux8_2),.dout(w_dff_B_pu99VB340_2),.clk(gclk));
	jdff dff_B_kvl75geT2_2(.din(w_dff_B_pu99VB340_2),.dout(w_dff_B_kvl75geT2_2),.clk(gclk));
	jdff dff_B_JxDq53FH1_2(.din(w_dff_B_kvl75geT2_2),.dout(w_dff_B_JxDq53FH1_2),.clk(gclk));
	jdff dff_B_N4LiO5Lb4_2(.din(w_dff_B_JxDq53FH1_2),.dout(w_dff_B_N4LiO5Lb4_2),.clk(gclk));
	jdff dff_B_wTHAbH3L8_2(.din(w_dff_B_N4LiO5Lb4_2),.dout(w_dff_B_wTHAbH3L8_2),.clk(gclk));
	jdff dff_B_PS2vrbAn7_2(.din(w_dff_B_wTHAbH3L8_2),.dout(w_dff_B_PS2vrbAn7_2),.clk(gclk));
	jdff dff_B_kV5qJHLH8_2(.din(w_dff_B_PS2vrbAn7_2),.dout(w_dff_B_kV5qJHLH8_2),.clk(gclk));
	jdff dff_B_IBjgHtyl9_2(.din(w_dff_B_kV5qJHLH8_2),.dout(w_dff_B_IBjgHtyl9_2),.clk(gclk));
	jdff dff_B_Yyw7O13w6_2(.din(w_dff_B_IBjgHtyl9_2),.dout(w_dff_B_Yyw7O13w6_2),.clk(gclk));
	jdff dff_B_shTCMpjF3_2(.din(w_dff_B_Yyw7O13w6_2),.dout(w_dff_B_shTCMpjF3_2),.clk(gclk));
	jdff dff_B_nQFoaHz82_2(.din(w_dff_B_shTCMpjF3_2),.dout(w_dff_B_nQFoaHz82_2),.clk(gclk));
	jdff dff_B_SY5ktz1Q7_2(.din(w_dff_B_nQFoaHz82_2),.dout(w_dff_B_SY5ktz1Q7_2),.clk(gclk));
	jdff dff_B_wi7OBm364_2(.din(w_dff_B_SY5ktz1Q7_2),.dout(w_dff_B_wi7OBm364_2),.clk(gclk));
	jdff dff_B_6qdMvcAC0_2(.din(w_dff_B_wi7OBm364_2),.dout(w_dff_B_6qdMvcAC0_2),.clk(gclk));
	jdff dff_B_DHkkivkZ8_2(.din(w_dff_B_6qdMvcAC0_2),.dout(w_dff_B_DHkkivkZ8_2),.clk(gclk));
	jdff dff_B_3TmBEJSr7_1(.din(n962),.dout(w_dff_B_3TmBEJSr7_1),.clk(gclk));
	jdff dff_B_A06MPEgt5_2(.din(n856),.dout(w_dff_B_A06MPEgt5_2),.clk(gclk));
	jdff dff_B_YROz2R6i2_2(.din(w_dff_B_A06MPEgt5_2),.dout(w_dff_B_YROz2R6i2_2),.clk(gclk));
	jdff dff_B_tl21GLti4_2(.din(w_dff_B_YROz2R6i2_2),.dout(w_dff_B_tl21GLti4_2),.clk(gclk));
	jdff dff_B_zlQkHDtW8_2(.din(w_dff_B_tl21GLti4_2),.dout(w_dff_B_zlQkHDtW8_2),.clk(gclk));
	jdff dff_B_xbw2aLdN8_2(.din(w_dff_B_zlQkHDtW8_2),.dout(w_dff_B_xbw2aLdN8_2),.clk(gclk));
	jdff dff_B_vR4YPr1b0_2(.din(w_dff_B_xbw2aLdN8_2),.dout(w_dff_B_vR4YPr1b0_2),.clk(gclk));
	jdff dff_B_EHT8PmzI8_2(.din(w_dff_B_vR4YPr1b0_2),.dout(w_dff_B_EHT8PmzI8_2),.clk(gclk));
	jdff dff_B_grUEZkXN1_2(.din(w_dff_B_EHT8PmzI8_2),.dout(w_dff_B_grUEZkXN1_2),.clk(gclk));
	jdff dff_B_lf9HrfCw9_2(.din(w_dff_B_grUEZkXN1_2),.dout(w_dff_B_lf9HrfCw9_2),.clk(gclk));
	jdff dff_B_JQ958yAm5_2(.din(w_dff_B_lf9HrfCw9_2),.dout(w_dff_B_JQ958yAm5_2),.clk(gclk));
	jdff dff_B_PaCN99jw2_2(.din(w_dff_B_JQ958yAm5_2),.dout(w_dff_B_PaCN99jw2_2),.clk(gclk));
	jdff dff_B_s8jj7hbg9_2(.din(w_dff_B_PaCN99jw2_2),.dout(w_dff_B_s8jj7hbg9_2),.clk(gclk));
	jdff dff_B_QTB9aI7J6_2(.din(w_dff_B_s8jj7hbg9_2),.dout(w_dff_B_QTB9aI7J6_2),.clk(gclk));
	jdff dff_B_M7kcno959_2(.din(w_dff_B_QTB9aI7J6_2),.dout(w_dff_B_M7kcno959_2),.clk(gclk));
	jdff dff_B_a5GDJgSa4_2(.din(w_dff_B_M7kcno959_2),.dout(w_dff_B_a5GDJgSa4_2),.clk(gclk));
	jdff dff_B_kVp31UCR9_2(.din(w_dff_B_a5GDJgSa4_2),.dout(w_dff_B_kVp31UCR9_2),.clk(gclk));
	jdff dff_B_34QrVnqd4_2(.din(w_dff_B_kVp31UCR9_2),.dout(w_dff_B_34QrVnqd4_2),.clk(gclk));
	jdff dff_B_xZy6sAe14_2(.din(w_dff_B_34QrVnqd4_2),.dout(w_dff_B_xZy6sAe14_2),.clk(gclk));
	jdff dff_B_kdYGzVW45_2(.din(w_dff_B_xZy6sAe14_2),.dout(w_dff_B_kdYGzVW45_2),.clk(gclk));
	jdff dff_B_i3mTkYqK7_2(.din(w_dff_B_kdYGzVW45_2),.dout(w_dff_B_i3mTkYqK7_2),.clk(gclk));
	jdff dff_B_4KcQbGzm1_1(.din(n857),.dout(w_dff_B_4KcQbGzm1_1),.clk(gclk));
	jdff dff_B_zIrAZKW33_2(.din(n757),.dout(w_dff_B_zIrAZKW33_2),.clk(gclk));
	jdff dff_B_JPUDhBHX4_2(.din(w_dff_B_zIrAZKW33_2),.dout(w_dff_B_JPUDhBHX4_2),.clk(gclk));
	jdff dff_B_DQ822bHd0_2(.din(w_dff_B_JPUDhBHX4_2),.dout(w_dff_B_DQ822bHd0_2),.clk(gclk));
	jdff dff_B_GHKp6BXn5_2(.din(w_dff_B_DQ822bHd0_2),.dout(w_dff_B_GHKp6BXn5_2),.clk(gclk));
	jdff dff_B_4wBaTMAy5_2(.din(w_dff_B_GHKp6BXn5_2),.dout(w_dff_B_4wBaTMAy5_2),.clk(gclk));
	jdff dff_B_GMCQL4WO8_2(.din(w_dff_B_4wBaTMAy5_2),.dout(w_dff_B_GMCQL4WO8_2),.clk(gclk));
	jdff dff_B_bPkKppGB2_2(.din(w_dff_B_GMCQL4WO8_2),.dout(w_dff_B_bPkKppGB2_2),.clk(gclk));
	jdff dff_B_P3rlvkXe6_2(.din(w_dff_B_bPkKppGB2_2),.dout(w_dff_B_P3rlvkXe6_2),.clk(gclk));
	jdff dff_B_qCujv8D04_2(.din(w_dff_B_P3rlvkXe6_2),.dout(w_dff_B_qCujv8D04_2),.clk(gclk));
	jdff dff_B_M3Fmb5Ys5_2(.din(w_dff_B_qCujv8D04_2),.dout(w_dff_B_M3Fmb5Ys5_2),.clk(gclk));
	jdff dff_B_XnKRtw8C6_2(.din(w_dff_B_M3Fmb5Ys5_2),.dout(w_dff_B_XnKRtw8C6_2),.clk(gclk));
	jdff dff_B_yHYHCaxJ8_2(.din(w_dff_B_XnKRtw8C6_2),.dout(w_dff_B_yHYHCaxJ8_2),.clk(gclk));
	jdff dff_B_rNKyEzJP1_2(.din(w_dff_B_yHYHCaxJ8_2),.dout(w_dff_B_rNKyEzJP1_2),.clk(gclk));
	jdff dff_B_zjjrUoGh4_2(.din(w_dff_B_rNKyEzJP1_2),.dout(w_dff_B_zjjrUoGh4_2),.clk(gclk));
	jdff dff_B_PNJ5fSUm2_2(.din(w_dff_B_zjjrUoGh4_2),.dout(w_dff_B_PNJ5fSUm2_2),.clk(gclk));
	jdff dff_B_4fxM2bAj6_2(.din(w_dff_B_PNJ5fSUm2_2),.dout(w_dff_B_4fxM2bAj6_2),.clk(gclk));
	jdff dff_B_OZfAXnUQ6_2(.din(w_dff_B_4fxM2bAj6_2),.dout(w_dff_B_OZfAXnUQ6_2),.clk(gclk));
	jdff dff_B_tWkl39uc5_2(.din(w_dff_B_OZfAXnUQ6_2),.dout(w_dff_B_tWkl39uc5_2),.clk(gclk));
	jdff dff_B_AVYQgcJo9_1(.din(n758),.dout(w_dff_B_AVYQgcJo9_1),.clk(gclk));
	jdff dff_B_FCfwY96i0_2(.din(n664),.dout(w_dff_B_FCfwY96i0_2),.clk(gclk));
	jdff dff_B_k2grJYnE4_2(.din(w_dff_B_FCfwY96i0_2),.dout(w_dff_B_k2grJYnE4_2),.clk(gclk));
	jdff dff_B_sCvb2oUk8_2(.din(w_dff_B_k2grJYnE4_2),.dout(w_dff_B_sCvb2oUk8_2),.clk(gclk));
	jdff dff_B_z7aJZkI97_2(.din(w_dff_B_sCvb2oUk8_2),.dout(w_dff_B_z7aJZkI97_2),.clk(gclk));
	jdff dff_B_tMEmoz6P1_2(.din(w_dff_B_z7aJZkI97_2),.dout(w_dff_B_tMEmoz6P1_2),.clk(gclk));
	jdff dff_B_LlS9wLXh2_2(.din(w_dff_B_tMEmoz6P1_2),.dout(w_dff_B_LlS9wLXh2_2),.clk(gclk));
	jdff dff_B_slm2WGys1_2(.din(w_dff_B_LlS9wLXh2_2),.dout(w_dff_B_slm2WGys1_2),.clk(gclk));
	jdff dff_B_9e85SUql4_2(.din(w_dff_B_slm2WGys1_2),.dout(w_dff_B_9e85SUql4_2),.clk(gclk));
	jdff dff_B_VgODNAGO3_2(.din(w_dff_B_9e85SUql4_2),.dout(w_dff_B_VgODNAGO3_2),.clk(gclk));
	jdff dff_B_MpOvCXKS5_2(.din(w_dff_B_VgODNAGO3_2),.dout(w_dff_B_MpOvCXKS5_2),.clk(gclk));
	jdff dff_B_MkymvTnz7_2(.din(w_dff_B_MpOvCXKS5_2),.dout(w_dff_B_MkymvTnz7_2),.clk(gclk));
	jdff dff_B_YjBIlWd48_2(.din(w_dff_B_MkymvTnz7_2),.dout(w_dff_B_YjBIlWd48_2),.clk(gclk));
	jdff dff_B_WURChH2z1_2(.din(w_dff_B_YjBIlWd48_2),.dout(w_dff_B_WURChH2z1_2),.clk(gclk));
	jdff dff_B_nEEra4m92_2(.din(w_dff_B_WURChH2z1_2),.dout(w_dff_B_nEEra4m92_2),.clk(gclk));
	jdff dff_B_0PjRQSM98_2(.din(w_dff_B_nEEra4m92_2),.dout(w_dff_B_0PjRQSM98_2),.clk(gclk));
	jdff dff_B_wrtKf0bo3_2(.din(w_dff_B_0PjRQSM98_2),.dout(w_dff_B_wrtKf0bo3_2),.clk(gclk));
	jdff dff_B_qIP4ZgBY5_1(.din(n665),.dout(w_dff_B_qIP4ZgBY5_1),.clk(gclk));
	jdff dff_B_ZVvaXVXz7_2(.din(n578),.dout(w_dff_B_ZVvaXVXz7_2),.clk(gclk));
	jdff dff_B_W9ZGgO086_2(.din(w_dff_B_ZVvaXVXz7_2),.dout(w_dff_B_W9ZGgO086_2),.clk(gclk));
	jdff dff_B_Jr55POId3_2(.din(w_dff_B_W9ZGgO086_2),.dout(w_dff_B_Jr55POId3_2),.clk(gclk));
	jdff dff_B_GfCCucKV8_2(.din(w_dff_B_Jr55POId3_2),.dout(w_dff_B_GfCCucKV8_2),.clk(gclk));
	jdff dff_B_8GYsv1kC8_2(.din(w_dff_B_GfCCucKV8_2),.dout(w_dff_B_8GYsv1kC8_2),.clk(gclk));
	jdff dff_B_RmaF4cQG2_2(.din(w_dff_B_8GYsv1kC8_2),.dout(w_dff_B_RmaF4cQG2_2),.clk(gclk));
	jdff dff_B_I8CXgn2L7_2(.din(w_dff_B_RmaF4cQG2_2),.dout(w_dff_B_I8CXgn2L7_2),.clk(gclk));
	jdff dff_B_XaU6V0Ck5_2(.din(w_dff_B_I8CXgn2L7_2),.dout(w_dff_B_XaU6V0Ck5_2),.clk(gclk));
	jdff dff_B_3S4Kr9Iw2_2(.din(w_dff_B_XaU6V0Ck5_2),.dout(w_dff_B_3S4Kr9Iw2_2),.clk(gclk));
	jdff dff_B_kdQc0vX30_2(.din(w_dff_B_3S4Kr9Iw2_2),.dout(w_dff_B_kdQc0vX30_2),.clk(gclk));
	jdff dff_B_BbPEeNoj1_2(.din(w_dff_B_kdQc0vX30_2),.dout(w_dff_B_BbPEeNoj1_2),.clk(gclk));
	jdff dff_B_tyw3JFfG4_2(.din(w_dff_B_BbPEeNoj1_2),.dout(w_dff_B_tyw3JFfG4_2),.clk(gclk));
	jdff dff_B_b5PoWetD6_2(.din(w_dff_B_tyw3JFfG4_2),.dout(w_dff_B_b5PoWetD6_2),.clk(gclk));
	jdff dff_B_YeAMfOBG9_2(.din(w_dff_B_b5PoWetD6_2),.dout(w_dff_B_YeAMfOBG9_2),.clk(gclk));
	jdff dff_B_Cn4ggaBf8_1(.din(n579),.dout(w_dff_B_Cn4ggaBf8_1),.clk(gclk));
	jdff dff_B_IneA9yhg0_2(.din(n499),.dout(w_dff_B_IneA9yhg0_2),.clk(gclk));
	jdff dff_B_sSHGSfMz1_2(.din(w_dff_B_IneA9yhg0_2),.dout(w_dff_B_sSHGSfMz1_2),.clk(gclk));
	jdff dff_B_kFpYbUMO4_2(.din(w_dff_B_sSHGSfMz1_2),.dout(w_dff_B_kFpYbUMO4_2),.clk(gclk));
	jdff dff_B_tQsDpTIQ5_2(.din(w_dff_B_kFpYbUMO4_2),.dout(w_dff_B_tQsDpTIQ5_2),.clk(gclk));
	jdff dff_B_dVGs5xcI9_2(.din(w_dff_B_tQsDpTIQ5_2),.dout(w_dff_B_dVGs5xcI9_2),.clk(gclk));
	jdff dff_B_isn4nnSQ6_2(.din(w_dff_B_dVGs5xcI9_2),.dout(w_dff_B_isn4nnSQ6_2),.clk(gclk));
	jdff dff_B_1WHfJ1Hh1_2(.din(w_dff_B_isn4nnSQ6_2),.dout(w_dff_B_1WHfJ1Hh1_2),.clk(gclk));
	jdff dff_B_RvRI9bDG8_2(.din(w_dff_B_1WHfJ1Hh1_2),.dout(w_dff_B_RvRI9bDG8_2),.clk(gclk));
	jdff dff_B_Y37IMIYK6_2(.din(w_dff_B_RvRI9bDG8_2),.dout(w_dff_B_Y37IMIYK6_2),.clk(gclk));
	jdff dff_B_dfDpnIzb4_2(.din(w_dff_B_Y37IMIYK6_2),.dout(w_dff_B_dfDpnIzb4_2),.clk(gclk));
	jdff dff_B_ijB8H5kj6_2(.din(w_dff_B_dfDpnIzb4_2),.dout(w_dff_B_ijB8H5kj6_2),.clk(gclk));
	jdff dff_B_iyTxPbzz4_2(.din(w_dff_B_ijB8H5kj6_2),.dout(w_dff_B_iyTxPbzz4_2),.clk(gclk));
	jdff dff_B_Bj9aSqi12_1(.din(n500),.dout(w_dff_B_Bj9aSqi12_1),.clk(gclk));
	jdff dff_B_6jOT558k5_2(.din(n427),.dout(w_dff_B_6jOT558k5_2),.clk(gclk));
	jdff dff_B_a3kqAr9B3_2(.din(w_dff_B_6jOT558k5_2),.dout(w_dff_B_a3kqAr9B3_2),.clk(gclk));
	jdff dff_B_ZY9Ygz6Y6_2(.din(w_dff_B_a3kqAr9B3_2),.dout(w_dff_B_ZY9Ygz6Y6_2),.clk(gclk));
	jdff dff_B_kgEVeQD81_2(.din(w_dff_B_ZY9Ygz6Y6_2),.dout(w_dff_B_kgEVeQD81_2),.clk(gclk));
	jdff dff_B_WWI3SvlO4_2(.din(w_dff_B_kgEVeQD81_2),.dout(w_dff_B_WWI3SvlO4_2),.clk(gclk));
	jdff dff_B_5Nc4NQKD6_2(.din(w_dff_B_WWI3SvlO4_2),.dout(w_dff_B_5Nc4NQKD6_2),.clk(gclk));
	jdff dff_B_9HaZCoiB2_2(.din(w_dff_B_5Nc4NQKD6_2),.dout(w_dff_B_9HaZCoiB2_2),.clk(gclk));
	jdff dff_B_1OHFcMK08_2(.din(w_dff_B_9HaZCoiB2_2),.dout(w_dff_B_1OHFcMK08_2),.clk(gclk));
	jdff dff_B_V6Ai4syZ5_2(.din(w_dff_B_1OHFcMK08_2),.dout(w_dff_B_V6Ai4syZ5_2),.clk(gclk));
	jdff dff_B_EA0egYHr7_2(.din(w_dff_B_V6Ai4syZ5_2),.dout(w_dff_B_EA0egYHr7_2),.clk(gclk));
	jdff dff_B_e5zG3G192_1(.din(n428),.dout(w_dff_B_e5zG3G192_1),.clk(gclk));
	jdff dff_B_hHF4PLv98_2(.din(n363),.dout(w_dff_B_hHF4PLv98_2),.clk(gclk));
	jdff dff_B_vKloUbis9_2(.din(w_dff_B_hHF4PLv98_2),.dout(w_dff_B_vKloUbis9_2),.clk(gclk));
	jdff dff_B_yUfKHhCJ3_2(.din(w_dff_B_vKloUbis9_2),.dout(w_dff_B_yUfKHhCJ3_2),.clk(gclk));
	jdff dff_B_Jt8mYg262_2(.din(w_dff_B_yUfKHhCJ3_2),.dout(w_dff_B_Jt8mYg262_2),.clk(gclk));
	jdff dff_B_0rTavOea3_2(.din(w_dff_B_Jt8mYg262_2),.dout(w_dff_B_0rTavOea3_2),.clk(gclk));
	jdff dff_B_J5a6kTfg1_2(.din(w_dff_B_0rTavOea3_2),.dout(w_dff_B_J5a6kTfg1_2),.clk(gclk));
	jdff dff_B_CyeZAuXr7_2(.din(w_dff_B_J5a6kTfg1_2),.dout(w_dff_B_CyeZAuXr7_2),.clk(gclk));
	jdff dff_B_5ER2SwBJ6_2(.din(w_dff_B_CyeZAuXr7_2),.dout(w_dff_B_5ER2SwBJ6_2),.clk(gclk));
	jdff dff_B_uosZhQmA9_1(.din(n364),.dout(w_dff_B_uosZhQmA9_1),.clk(gclk));
	jdff dff_B_fdLzkwVB3_2(.din(n305),.dout(w_dff_B_fdLzkwVB3_2),.clk(gclk));
	jdff dff_B_n7DB7ScB4_2(.din(w_dff_B_fdLzkwVB3_2),.dout(w_dff_B_n7DB7ScB4_2),.clk(gclk));
	jdff dff_B_u7KsKqec9_2(.din(w_dff_B_n7DB7ScB4_2),.dout(w_dff_B_u7KsKqec9_2),.clk(gclk));
	jdff dff_B_b02pt5Jq6_2(.din(w_dff_B_u7KsKqec9_2),.dout(w_dff_B_b02pt5Jq6_2),.clk(gclk));
	jdff dff_B_2xUaqW1E6_2(.din(w_dff_B_b02pt5Jq6_2),.dout(w_dff_B_2xUaqW1E6_2),.clk(gclk));
	jdff dff_B_iy6eoe9I4_2(.din(w_dff_B_2xUaqW1E6_2),.dout(w_dff_B_iy6eoe9I4_2),.clk(gclk));
	jdff dff_B_WS4OrXGn4_1(.din(n306),.dout(w_dff_B_WS4OrXGn4_1),.clk(gclk));
	jdff dff_B_y6wDHljS6_1(.din(w_dff_B_WS4OrXGn4_1),.dout(w_dff_B_y6wDHljS6_1),.clk(gclk));
	jdff dff_B_w6gx9XeJ2_2(.din(n254),.dout(w_dff_B_w6gx9XeJ2_2),.clk(gclk));
	jdff dff_B_NoHTSPrv1_2(.din(w_dff_B_w6gx9XeJ2_2),.dout(w_dff_B_NoHTSPrv1_2),.clk(gclk));
	jdff dff_B_YpiywRqR1_2(.din(w_dff_B_NoHTSPrv1_2),.dout(w_dff_B_YpiywRqR1_2),.clk(gclk));
	jdff dff_B_VKVv2ZlL7_2(.din(w_dff_B_YpiywRqR1_2),.dout(w_dff_B_VKVv2ZlL7_2),.clk(gclk));
	jdff dff_A_sffExBlQ5_1(.dout(w_n261_0[1]),.din(w_dff_A_sffExBlQ5_1),.clk(gclk));
	jdff dff_B_QaA4BnNI5_1(.din(n256),.dout(w_dff_B_QaA4BnNI5_1),.clk(gclk));
	jdff dff_B_nNWTPtOn8_1(.din(w_dff_B_QaA4BnNI5_1),.dout(w_dff_B_nNWTPtOn8_1),.clk(gclk));
	jdff dff_A_lTu2GWwo3_1(.dout(w_n210_0[1]),.din(w_dff_A_lTu2GWwo3_1),.clk(gclk));
	jdff dff_A_q2YgquF76_2(.dout(w_n210_0[2]),.din(w_dff_A_q2YgquF76_2),.clk(gclk));
	jdff dff_A_jkneepKI9_2(.dout(w_dff_A_q2YgquF76_2),.din(w_dff_A_jkneepKI9_2),.clk(gclk));
	jdff dff_B_kI2ENWMc5_2(.din(n1496),.dout(w_dff_B_kI2ENWMc5_2),.clk(gclk));
	jdff dff_B_QXDLZGjL9_2(.din(w_dff_B_kI2ENWMc5_2),.dout(w_dff_B_QXDLZGjL9_2),.clk(gclk));
	jdff dff_B_Wc61OfOK0_1(.din(n1494),.dout(w_dff_B_Wc61OfOK0_1),.clk(gclk));
	jdff dff_B_K06jwAoZ4_2(.din(n1421),.dout(w_dff_B_K06jwAoZ4_2),.clk(gclk));
	jdff dff_B_jElGjNCa7_2(.din(w_dff_B_K06jwAoZ4_2),.dout(w_dff_B_jElGjNCa7_2),.clk(gclk));
	jdff dff_B_7d8eh8lw1_2(.din(w_dff_B_jElGjNCa7_2),.dout(w_dff_B_7d8eh8lw1_2),.clk(gclk));
	jdff dff_B_dQEkcGzT0_2(.din(w_dff_B_7d8eh8lw1_2),.dout(w_dff_B_dQEkcGzT0_2),.clk(gclk));
	jdff dff_B_sHnnsn2q7_2(.din(w_dff_B_dQEkcGzT0_2),.dout(w_dff_B_sHnnsn2q7_2),.clk(gclk));
	jdff dff_B_f2o4nSvx7_2(.din(w_dff_B_sHnnsn2q7_2),.dout(w_dff_B_f2o4nSvx7_2),.clk(gclk));
	jdff dff_B_PQGJr6EU5_2(.din(w_dff_B_f2o4nSvx7_2),.dout(w_dff_B_PQGJr6EU5_2),.clk(gclk));
	jdff dff_B_qU5riOqO4_2(.din(w_dff_B_PQGJr6EU5_2),.dout(w_dff_B_qU5riOqO4_2),.clk(gclk));
	jdff dff_B_tyfWo8yg3_2(.din(w_dff_B_qU5riOqO4_2),.dout(w_dff_B_tyfWo8yg3_2),.clk(gclk));
	jdff dff_B_ivJ0EobA9_2(.din(w_dff_B_tyfWo8yg3_2),.dout(w_dff_B_ivJ0EobA9_2),.clk(gclk));
	jdff dff_B_FwGifej58_2(.din(w_dff_B_ivJ0EobA9_2),.dout(w_dff_B_FwGifej58_2),.clk(gclk));
	jdff dff_B_loPUOzs56_2(.din(w_dff_B_FwGifej58_2),.dout(w_dff_B_loPUOzs56_2),.clk(gclk));
	jdff dff_B_uaAIJsIE8_2(.din(w_dff_B_loPUOzs56_2),.dout(w_dff_B_uaAIJsIE8_2),.clk(gclk));
	jdff dff_B_Sdx0dtdJ1_2(.din(w_dff_B_uaAIJsIE8_2),.dout(w_dff_B_Sdx0dtdJ1_2),.clk(gclk));
	jdff dff_B_iepCSMSW9_2(.din(w_dff_B_Sdx0dtdJ1_2),.dout(w_dff_B_iepCSMSW9_2),.clk(gclk));
	jdff dff_B_fTTMvD3V9_2(.din(w_dff_B_iepCSMSW9_2),.dout(w_dff_B_fTTMvD3V9_2),.clk(gclk));
	jdff dff_B_zdb5BAwl6_2(.din(w_dff_B_fTTMvD3V9_2),.dout(w_dff_B_zdb5BAwl6_2),.clk(gclk));
	jdff dff_B_4G62qj6k2_2(.din(w_dff_B_zdb5BAwl6_2),.dout(w_dff_B_4G62qj6k2_2),.clk(gclk));
	jdff dff_B_Rj2vvGED0_2(.din(w_dff_B_4G62qj6k2_2),.dout(w_dff_B_Rj2vvGED0_2),.clk(gclk));
	jdff dff_B_ngggpycu0_2(.din(w_dff_B_Rj2vvGED0_2),.dout(w_dff_B_ngggpycu0_2),.clk(gclk));
	jdff dff_B_Hg5LHLr43_2(.din(w_dff_B_ngggpycu0_2),.dout(w_dff_B_Hg5LHLr43_2),.clk(gclk));
	jdff dff_B_0299Flaz5_2(.din(w_dff_B_Hg5LHLr43_2),.dout(w_dff_B_0299Flaz5_2),.clk(gclk));
	jdff dff_B_o5AnkwZD8_2(.din(w_dff_B_0299Flaz5_2),.dout(w_dff_B_o5AnkwZD8_2),.clk(gclk));
	jdff dff_B_JPxaRGMO5_2(.din(w_dff_B_o5AnkwZD8_2),.dout(w_dff_B_JPxaRGMO5_2),.clk(gclk));
	jdff dff_B_d1YXzBx40_2(.din(w_dff_B_JPxaRGMO5_2),.dout(w_dff_B_d1YXzBx40_2),.clk(gclk));
	jdff dff_B_qcX1VLLs6_2(.din(w_dff_B_d1YXzBx40_2),.dout(w_dff_B_qcX1VLLs6_2),.clk(gclk));
	jdff dff_B_1zQJcAhG4_2(.din(w_dff_B_qcX1VLLs6_2),.dout(w_dff_B_1zQJcAhG4_2),.clk(gclk));
	jdff dff_B_33RengTd9_2(.din(w_dff_B_1zQJcAhG4_2),.dout(w_dff_B_33RengTd9_2),.clk(gclk));
	jdff dff_B_gbkHGl7v0_2(.din(w_dff_B_33RengTd9_2),.dout(w_dff_B_gbkHGl7v0_2),.clk(gclk));
	jdff dff_B_aYTb8ZT22_2(.din(w_dff_B_gbkHGl7v0_2),.dout(w_dff_B_aYTb8ZT22_2),.clk(gclk));
	jdff dff_B_iB0L1D0K5_2(.din(w_dff_B_aYTb8ZT22_2),.dout(w_dff_B_iB0L1D0K5_2),.clk(gclk));
	jdff dff_B_fvWhLSL56_2(.din(w_dff_B_iB0L1D0K5_2),.dout(w_dff_B_fvWhLSL56_2),.clk(gclk));
	jdff dff_B_UMCpyrhA1_2(.din(w_dff_B_fvWhLSL56_2),.dout(w_dff_B_UMCpyrhA1_2),.clk(gclk));
	jdff dff_B_DQUrikwz3_2(.din(w_dff_B_UMCpyrhA1_2),.dout(w_dff_B_DQUrikwz3_2),.clk(gclk));
	jdff dff_B_PBkw2l3d5_2(.din(w_dff_B_DQUrikwz3_2),.dout(w_dff_B_PBkw2l3d5_2),.clk(gclk));
	jdff dff_B_1m2STfot5_2(.din(w_dff_B_PBkw2l3d5_2),.dout(w_dff_B_1m2STfot5_2),.clk(gclk));
	jdff dff_B_MO3xkrHL2_2(.din(w_dff_B_1m2STfot5_2),.dout(w_dff_B_MO3xkrHL2_2),.clk(gclk));
	jdff dff_B_5MuID1Q30_1(.din(n1492),.dout(w_dff_B_5MuID1Q30_1),.clk(gclk));
	jdff dff_A_km6ZBDLX1_1(.dout(w_n1424_0[1]),.din(w_dff_A_km6ZBDLX1_1),.clk(gclk));
	jdff dff_B_Jch7zrMC4_1(.din(n1422),.dout(w_dff_B_Jch7zrMC4_1),.clk(gclk));
	jdff dff_B_EE2ppDoD8_2(.din(n1343),.dout(w_dff_B_EE2ppDoD8_2),.clk(gclk));
	jdff dff_B_LwLvKN2Y4_2(.din(w_dff_B_EE2ppDoD8_2),.dout(w_dff_B_LwLvKN2Y4_2),.clk(gclk));
	jdff dff_B_3OTw13iF9_2(.din(w_dff_B_LwLvKN2Y4_2),.dout(w_dff_B_3OTw13iF9_2),.clk(gclk));
	jdff dff_B_ZclvFa4K6_2(.din(w_dff_B_3OTw13iF9_2),.dout(w_dff_B_ZclvFa4K6_2),.clk(gclk));
	jdff dff_B_CVlt1Gry9_2(.din(w_dff_B_ZclvFa4K6_2),.dout(w_dff_B_CVlt1Gry9_2),.clk(gclk));
	jdff dff_B_69I4gQ4O2_2(.din(w_dff_B_CVlt1Gry9_2),.dout(w_dff_B_69I4gQ4O2_2),.clk(gclk));
	jdff dff_B_9nES55Xl7_2(.din(w_dff_B_69I4gQ4O2_2),.dout(w_dff_B_9nES55Xl7_2),.clk(gclk));
	jdff dff_B_CHzIh5Jl3_2(.din(w_dff_B_9nES55Xl7_2),.dout(w_dff_B_CHzIh5Jl3_2),.clk(gclk));
	jdff dff_B_onC38s4b0_2(.din(w_dff_B_CHzIh5Jl3_2),.dout(w_dff_B_onC38s4b0_2),.clk(gclk));
	jdff dff_B_EFiOk7zX8_2(.din(w_dff_B_onC38s4b0_2),.dout(w_dff_B_EFiOk7zX8_2),.clk(gclk));
	jdff dff_B_NDXDpqvm9_2(.din(w_dff_B_EFiOk7zX8_2),.dout(w_dff_B_NDXDpqvm9_2),.clk(gclk));
	jdff dff_B_VisgXv3B3_2(.din(w_dff_B_NDXDpqvm9_2),.dout(w_dff_B_VisgXv3B3_2),.clk(gclk));
	jdff dff_B_HSC6F05V8_2(.din(w_dff_B_VisgXv3B3_2),.dout(w_dff_B_HSC6F05V8_2),.clk(gclk));
	jdff dff_B_D6VgF25T1_2(.din(w_dff_B_HSC6F05V8_2),.dout(w_dff_B_D6VgF25T1_2),.clk(gclk));
	jdff dff_B_aHyL4SUc6_2(.din(w_dff_B_D6VgF25T1_2),.dout(w_dff_B_aHyL4SUc6_2),.clk(gclk));
	jdff dff_B_tI5ARTMl5_2(.din(w_dff_B_aHyL4SUc6_2),.dout(w_dff_B_tI5ARTMl5_2),.clk(gclk));
	jdff dff_B_5dlPVokj1_2(.din(w_dff_B_tI5ARTMl5_2),.dout(w_dff_B_5dlPVokj1_2),.clk(gclk));
	jdff dff_B_YlMp9Zff7_2(.din(w_dff_B_5dlPVokj1_2),.dout(w_dff_B_YlMp9Zff7_2),.clk(gclk));
	jdff dff_B_KHa3WL0A6_2(.din(w_dff_B_YlMp9Zff7_2),.dout(w_dff_B_KHa3WL0A6_2),.clk(gclk));
	jdff dff_B_hnyuUPKr5_2(.din(w_dff_B_KHa3WL0A6_2),.dout(w_dff_B_hnyuUPKr5_2),.clk(gclk));
	jdff dff_B_qWAbQCi56_2(.din(w_dff_B_hnyuUPKr5_2),.dout(w_dff_B_qWAbQCi56_2),.clk(gclk));
	jdff dff_B_C8A15Wz96_2(.din(w_dff_B_qWAbQCi56_2),.dout(w_dff_B_C8A15Wz96_2),.clk(gclk));
	jdff dff_B_cpMeQEWp9_2(.din(w_dff_B_C8A15Wz96_2),.dout(w_dff_B_cpMeQEWp9_2),.clk(gclk));
	jdff dff_B_DN7WeaL16_2(.din(w_dff_B_cpMeQEWp9_2),.dout(w_dff_B_DN7WeaL16_2),.clk(gclk));
	jdff dff_B_9nIFu5I88_2(.din(w_dff_B_DN7WeaL16_2),.dout(w_dff_B_9nIFu5I88_2),.clk(gclk));
	jdff dff_B_zR0bJ7Qn3_2(.din(w_dff_B_9nIFu5I88_2),.dout(w_dff_B_zR0bJ7Qn3_2),.clk(gclk));
	jdff dff_B_rsibzmaI4_2(.din(w_dff_B_zR0bJ7Qn3_2),.dout(w_dff_B_rsibzmaI4_2),.clk(gclk));
	jdff dff_B_wo4XRTlx0_2(.din(w_dff_B_rsibzmaI4_2),.dout(w_dff_B_wo4XRTlx0_2),.clk(gclk));
	jdff dff_B_xh8Ntsfk2_2(.din(w_dff_B_wo4XRTlx0_2),.dout(w_dff_B_xh8Ntsfk2_2),.clk(gclk));
	jdff dff_B_W1eUP5YR8_2(.din(w_dff_B_xh8Ntsfk2_2),.dout(w_dff_B_W1eUP5YR8_2),.clk(gclk));
	jdff dff_B_DKzJq4jk9_2(.din(w_dff_B_W1eUP5YR8_2),.dout(w_dff_B_DKzJq4jk9_2),.clk(gclk));
	jdff dff_B_kiAL6Qoz4_2(.din(w_dff_B_DKzJq4jk9_2),.dout(w_dff_B_kiAL6Qoz4_2),.clk(gclk));
	jdff dff_B_hARVlZ0U7_2(.din(n1346),.dout(w_dff_B_hARVlZ0U7_2),.clk(gclk));
	jdff dff_B_ivnOAsjy4_1(.din(n1344),.dout(w_dff_B_ivnOAsjy4_1),.clk(gclk));
	jdff dff_B_LXVEP8uZ8_2(.din(n1258),.dout(w_dff_B_LXVEP8uZ8_2),.clk(gclk));
	jdff dff_B_4poR2CQm4_2(.din(w_dff_B_LXVEP8uZ8_2),.dout(w_dff_B_4poR2CQm4_2),.clk(gclk));
	jdff dff_B_mgOadkX03_2(.din(w_dff_B_4poR2CQm4_2),.dout(w_dff_B_mgOadkX03_2),.clk(gclk));
	jdff dff_B_mgD8YAwU6_2(.din(w_dff_B_mgOadkX03_2),.dout(w_dff_B_mgD8YAwU6_2),.clk(gclk));
	jdff dff_B_Hdhj5BRk0_2(.din(w_dff_B_mgD8YAwU6_2),.dout(w_dff_B_Hdhj5BRk0_2),.clk(gclk));
	jdff dff_B_mgW6aHdy9_2(.din(w_dff_B_Hdhj5BRk0_2),.dout(w_dff_B_mgW6aHdy9_2),.clk(gclk));
	jdff dff_B_0C8RqJtJ9_2(.din(w_dff_B_mgW6aHdy9_2),.dout(w_dff_B_0C8RqJtJ9_2),.clk(gclk));
	jdff dff_B_sdU84hag3_2(.din(w_dff_B_0C8RqJtJ9_2),.dout(w_dff_B_sdU84hag3_2),.clk(gclk));
	jdff dff_B_5w8UROTJ8_2(.din(w_dff_B_sdU84hag3_2),.dout(w_dff_B_5w8UROTJ8_2),.clk(gclk));
	jdff dff_B_qidCpLAl7_2(.din(w_dff_B_5w8UROTJ8_2),.dout(w_dff_B_qidCpLAl7_2),.clk(gclk));
	jdff dff_B_qwggIlGA0_2(.din(w_dff_B_qidCpLAl7_2),.dout(w_dff_B_qwggIlGA0_2),.clk(gclk));
	jdff dff_B_xGWCQptL5_2(.din(w_dff_B_qwggIlGA0_2),.dout(w_dff_B_xGWCQptL5_2),.clk(gclk));
	jdff dff_B_T0fvdXNe4_2(.din(w_dff_B_xGWCQptL5_2),.dout(w_dff_B_T0fvdXNe4_2),.clk(gclk));
	jdff dff_B_CQLgawAo8_2(.din(w_dff_B_T0fvdXNe4_2),.dout(w_dff_B_CQLgawAo8_2),.clk(gclk));
	jdff dff_B_HGMviyr69_2(.din(w_dff_B_CQLgawAo8_2),.dout(w_dff_B_HGMviyr69_2),.clk(gclk));
	jdff dff_B_R2fiFvk72_2(.din(w_dff_B_HGMviyr69_2),.dout(w_dff_B_R2fiFvk72_2),.clk(gclk));
	jdff dff_B_7a1bvLkJ6_2(.din(w_dff_B_R2fiFvk72_2),.dout(w_dff_B_7a1bvLkJ6_2),.clk(gclk));
	jdff dff_B_QMZZNcah3_2(.din(w_dff_B_7a1bvLkJ6_2),.dout(w_dff_B_QMZZNcah3_2),.clk(gclk));
	jdff dff_B_krobLoUg5_2(.din(w_dff_B_QMZZNcah3_2),.dout(w_dff_B_krobLoUg5_2),.clk(gclk));
	jdff dff_B_CJxFDmu99_2(.din(w_dff_B_krobLoUg5_2),.dout(w_dff_B_CJxFDmu99_2),.clk(gclk));
	jdff dff_B_Nm3JpYMv5_2(.din(w_dff_B_CJxFDmu99_2),.dout(w_dff_B_Nm3JpYMv5_2),.clk(gclk));
	jdff dff_B_rMvCm0j85_2(.din(w_dff_B_Nm3JpYMv5_2),.dout(w_dff_B_rMvCm0j85_2),.clk(gclk));
	jdff dff_B_8BFoXhsj4_2(.din(w_dff_B_rMvCm0j85_2),.dout(w_dff_B_8BFoXhsj4_2),.clk(gclk));
	jdff dff_B_USsMmGwY4_2(.din(w_dff_B_8BFoXhsj4_2),.dout(w_dff_B_USsMmGwY4_2),.clk(gclk));
	jdff dff_B_nIBugPL99_2(.din(w_dff_B_USsMmGwY4_2),.dout(w_dff_B_nIBugPL99_2),.clk(gclk));
	jdff dff_B_wdpfAOTz2_2(.din(w_dff_B_nIBugPL99_2),.dout(w_dff_B_wdpfAOTz2_2),.clk(gclk));
	jdff dff_B_rBZiQDny7_2(.din(w_dff_B_wdpfAOTz2_2),.dout(w_dff_B_rBZiQDny7_2),.clk(gclk));
	jdff dff_B_FkWhASko7_2(.din(w_dff_B_rBZiQDny7_2),.dout(w_dff_B_FkWhASko7_2),.clk(gclk));
	jdff dff_B_VQgZ5SR97_2(.din(w_dff_B_FkWhASko7_2),.dout(w_dff_B_VQgZ5SR97_2),.clk(gclk));
	jdff dff_B_r9HkWtyQ6_2(.din(n1261),.dout(w_dff_B_r9HkWtyQ6_2),.clk(gclk));
	jdff dff_B_cvqoWs9e8_1(.din(n1259),.dout(w_dff_B_cvqoWs9e8_1),.clk(gclk));
	jdff dff_B_FST0Ilhu0_2(.din(n1168),.dout(w_dff_B_FST0Ilhu0_2),.clk(gclk));
	jdff dff_B_LsqPvrrA9_2(.din(w_dff_B_FST0Ilhu0_2),.dout(w_dff_B_LsqPvrrA9_2),.clk(gclk));
	jdff dff_B_G8WZ7BDo4_2(.din(w_dff_B_LsqPvrrA9_2),.dout(w_dff_B_G8WZ7BDo4_2),.clk(gclk));
	jdff dff_B_OrqsD9Fv0_2(.din(w_dff_B_G8WZ7BDo4_2),.dout(w_dff_B_OrqsD9Fv0_2),.clk(gclk));
	jdff dff_B_tUHSKBNG1_2(.din(w_dff_B_OrqsD9Fv0_2),.dout(w_dff_B_tUHSKBNG1_2),.clk(gclk));
	jdff dff_B_opsqlyLX3_2(.din(w_dff_B_tUHSKBNG1_2),.dout(w_dff_B_opsqlyLX3_2),.clk(gclk));
	jdff dff_B_poDfQ2nZ2_2(.din(w_dff_B_opsqlyLX3_2),.dout(w_dff_B_poDfQ2nZ2_2),.clk(gclk));
	jdff dff_B_cOH5N3YD1_2(.din(w_dff_B_poDfQ2nZ2_2),.dout(w_dff_B_cOH5N3YD1_2),.clk(gclk));
	jdff dff_B_DGMxRnhr3_2(.din(w_dff_B_cOH5N3YD1_2),.dout(w_dff_B_DGMxRnhr3_2),.clk(gclk));
	jdff dff_B_cBoDgnvL0_2(.din(w_dff_B_DGMxRnhr3_2),.dout(w_dff_B_cBoDgnvL0_2),.clk(gclk));
	jdff dff_B_nzuSHpu41_2(.din(w_dff_B_cBoDgnvL0_2),.dout(w_dff_B_nzuSHpu41_2),.clk(gclk));
	jdff dff_B_jz5wnW713_2(.din(w_dff_B_nzuSHpu41_2),.dout(w_dff_B_jz5wnW713_2),.clk(gclk));
	jdff dff_B_eTYVcJPw7_2(.din(w_dff_B_jz5wnW713_2),.dout(w_dff_B_eTYVcJPw7_2),.clk(gclk));
	jdff dff_B_R5c1PYkn6_2(.din(w_dff_B_eTYVcJPw7_2),.dout(w_dff_B_R5c1PYkn6_2),.clk(gclk));
	jdff dff_B_xlhFY48i7_2(.din(w_dff_B_R5c1PYkn6_2),.dout(w_dff_B_xlhFY48i7_2),.clk(gclk));
	jdff dff_B_SJEh11Qb7_2(.din(w_dff_B_xlhFY48i7_2),.dout(w_dff_B_SJEh11Qb7_2),.clk(gclk));
	jdff dff_B_J3K6ptWE5_2(.din(w_dff_B_SJEh11Qb7_2),.dout(w_dff_B_J3K6ptWE5_2),.clk(gclk));
	jdff dff_B_qm05tenc4_2(.din(w_dff_B_J3K6ptWE5_2),.dout(w_dff_B_qm05tenc4_2),.clk(gclk));
	jdff dff_B_hZB5OZ4t3_2(.din(w_dff_B_qm05tenc4_2),.dout(w_dff_B_hZB5OZ4t3_2),.clk(gclk));
	jdff dff_B_9f49ZbKq8_2(.din(w_dff_B_hZB5OZ4t3_2),.dout(w_dff_B_9f49ZbKq8_2),.clk(gclk));
	jdff dff_B_wf7cz2mD1_2(.din(w_dff_B_9f49ZbKq8_2),.dout(w_dff_B_wf7cz2mD1_2),.clk(gclk));
	jdff dff_B_zS1qtQ2l2_2(.din(w_dff_B_wf7cz2mD1_2),.dout(w_dff_B_zS1qtQ2l2_2),.clk(gclk));
	jdff dff_B_OKJdbkSh3_2(.din(w_dff_B_zS1qtQ2l2_2),.dout(w_dff_B_OKJdbkSh3_2),.clk(gclk));
	jdff dff_B_64zbX8iC4_2(.din(w_dff_B_OKJdbkSh3_2),.dout(w_dff_B_64zbX8iC4_2),.clk(gclk));
	jdff dff_B_A7bc56LV9_2(.din(w_dff_B_64zbX8iC4_2),.dout(w_dff_B_A7bc56LV9_2),.clk(gclk));
	jdff dff_B_BeKR35A02_2(.din(w_dff_B_A7bc56LV9_2),.dout(w_dff_B_BeKR35A02_2),.clk(gclk));
	jdff dff_B_xl0I0JEE5_2(.din(n1171),.dout(w_dff_B_xl0I0JEE5_2),.clk(gclk));
	jdff dff_B_ELpE24bH9_1(.din(n1169),.dout(w_dff_B_ELpE24bH9_1),.clk(gclk));
	jdff dff_B_1GBAdd8W1_2(.din(n1064),.dout(w_dff_B_1GBAdd8W1_2),.clk(gclk));
	jdff dff_B_QbLr8CWZ7_2(.din(w_dff_B_1GBAdd8W1_2),.dout(w_dff_B_QbLr8CWZ7_2),.clk(gclk));
	jdff dff_B_JSMVuqLd7_2(.din(w_dff_B_QbLr8CWZ7_2),.dout(w_dff_B_JSMVuqLd7_2),.clk(gclk));
	jdff dff_B_dMOPpgOq5_2(.din(w_dff_B_JSMVuqLd7_2),.dout(w_dff_B_dMOPpgOq5_2),.clk(gclk));
	jdff dff_B_dGfTqZLC9_2(.din(w_dff_B_dMOPpgOq5_2),.dout(w_dff_B_dGfTqZLC9_2),.clk(gclk));
	jdff dff_B_LfOXdbJe2_2(.din(w_dff_B_dGfTqZLC9_2),.dout(w_dff_B_LfOXdbJe2_2),.clk(gclk));
	jdff dff_B_S6w4rrd83_2(.din(w_dff_B_LfOXdbJe2_2),.dout(w_dff_B_S6w4rrd83_2),.clk(gclk));
	jdff dff_B_oqevpRA25_2(.din(w_dff_B_S6w4rrd83_2),.dout(w_dff_B_oqevpRA25_2),.clk(gclk));
	jdff dff_B_S6dsqgZo0_2(.din(w_dff_B_oqevpRA25_2),.dout(w_dff_B_S6dsqgZo0_2),.clk(gclk));
	jdff dff_B_rk6T9Vx62_2(.din(w_dff_B_S6dsqgZo0_2),.dout(w_dff_B_rk6T9Vx62_2),.clk(gclk));
	jdff dff_B_woIeXbvP3_2(.din(w_dff_B_rk6T9Vx62_2),.dout(w_dff_B_woIeXbvP3_2),.clk(gclk));
	jdff dff_B_YXFIYIiR5_2(.din(w_dff_B_woIeXbvP3_2),.dout(w_dff_B_YXFIYIiR5_2),.clk(gclk));
	jdff dff_B_DaPraFpZ2_2(.din(w_dff_B_YXFIYIiR5_2),.dout(w_dff_B_DaPraFpZ2_2),.clk(gclk));
	jdff dff_B_M8I1E7Xv0_2(.din(w_dff_B_DaPraFpZ2_2),.dout(w_dff_B_M8I1E7Xv0_2),.clk(gclk));
	jdff dff_B_QBZIqR743_2(.din(w_dff_B_M8I1E7Xv0_2),.dout(w_dff_B_QBZIqR743_2),.clk(gclk));
	jdff dff_B_fq7qfXWc3_2(.din(w_dff_B_QBZIqR743_2),.dout(w_dff_B_fq7qfXWc3_2),.clk(gclk));
	jdff dff_B_b7YJJ5Yc3_2(.din(w_dff_B_fq7qfXWc3_2),.dout(w_dff_B_b7YJJ5Yc3_2),.clk(gclk));
	jdff dff_B_vYV35fv94_2(.din(w_dff_B_b7YJJ5Yc3_2),.dout(w_dff_B_vYV35fv94_2),.clk(gclk));
	jdff dff_B_nzpouyKv1_2(.din(w_dff_B_vYV35fv94_2),.dout(w_dff_B_nzpouyKv1_2),.clk(gclk));
	jdff dff_B_yvxZHNbN7_2(.din(w_dff_B_nzpouyKv1_2),.dout(w_dff_B_yvxZHNbN7_2),.clk(gclk));
	jdff dff_B_2mTGSGRM8_2(.din(w_dff_B_yvxZHNbN7_2),.dout(w_dff_B_2mTGSGRM8_2),.clk(gclk));
	jdff dff_B_mg7ZoLSc5_2(.din(w_dff_B_2mTGSGRM8_2),.dout(w_dff_B_mg7ZoLSc5_2),.clk(gclk));
	jdff dff_B_gIN7GL8I4_2(.din(w_dff_B_mg7ZoLSc5_2),.dout(w_dff_B_gIN7GL8I4_2),.clk(gclk));
	jdff dff_B_Vk4Qj9aA2_2(.din(n1067),.dout(w_dff_B_Vk4Qj9aA2_2),.clk(gclk));
	jdff dff_B_Usg5uhqf5_1(.din(n1065),.dout(w_dff_B_Usg5uhqf5_1),.clk(gclk));
	jdff dff_B_2TfIy28O0_2(.din(n966),.dout(w_dff_B_2TfIy28O0_2),.clk(gclk));
	jdff dff_B_OX9k87qZ1_2(.din(w_dff_B_2TfIy28O0_2),.dout(w_dff_B_OX9k87qZ1_2),.clk(gclk));
	jdff dff_B_VpDadZwI1_2(.din(w_dff_B_OX9k87qZ1_2),.dout(w_dff_B_VpDadZwI1_2),.clk(gclk));
	jdff dff_B_IyhPZD3n2_2(.din(w_dff_B_VpDadZwI1_2),.dout(w_dff_B_IyhPZD3n2_2),.clk(gclk));
	jdff dff_B_1i99748o7_2(.din(w_dff_B_IyhPZD3n2_2),.dout(w_dff_B_1i99748o7_2),.clk(gclk));
	jdff dff_B_Qz2hYg2v7_2(.din(w_dff_B_1i99748o7_2),.dout(w_dff_B_Qz2hYg2v7_2),.clk(gclk));
	jdff dff_B_4SFflszo3_2(.din(w_dff_B_Qz2hYg2v7_2),.dout(w_dff_B_4SFflszo3_2),.clk(gclk));
	jdff dff_B_bYqvUog75_2(.din(w_dff_B_4SFflszo3_2),.dout(w_dff_B_bYqvUog75_2),.clk(gclk));
	jdff dff_B_Xcae1ElU8_2(.din(w_dff_B_bYqvUog75_2),.dout(w_dff_B_Xcae1ElU8_2),.clk(gclk));
	jdff dff_B_yr7H8RoG8_2(.din(w_dff_B_Xcae1ElU8_2),.dout(w_dff_B_yr7H8RoG8_2),.clk(gclk));
	jdff dff_B_dqaXI5Q01_2(.din(w_dff_B_yr7H8RoG8_2),.dout(w_dff_B_dqaXI5Q01_2),.clk(gclk));
	jdff dff_B_PoKKm8Ac3_2(.din(w_dff_B_dqaXI5Q01_2),.dout(w_dff_B_PoKKm8Ac3_2),.clk(gclk));
	jdff dff_B_ehinX51G4_2(.din(w_dff_B_PoKKm8Ac3_2),.dout(w_dff_B_ehinX51G4_2),.clk(gclk));
	jdff dff_B_BirjClnD4_2(.din(w_dff_B_ehinX51G4_2),.dout(w_dff_B_BirjClnD4_2),.clk(gclk));
	jdff dff_B_3WQ4HrMA0_2(.din(w_dff_B_BirjClnD4_2),.dout(w_dff_B_3WQ4HrMA0_2),.clk(gclk));
	jdff dff_B_g5C6IMhb1_2(.din(w_dff_B_3WQ4HrMA0_2),.dout(w_dff_B_g5C6IMhb1_2),.clk(gclk));
	jdff dff_B_y8C8BSDi7_2(.din(w_dff_B_g5C6IMhb1_2),.dout(w_dff_B_y8C8BSDi7_2),.clk(gclk));
	jdff dff_B_gtSv2GW19_2(.din(w_dff_B_y8C8BSDi7_2),.dout(w_dff_B_gtSv2GW19_2),.clk(gclk));
	jdff dff_B_Rg2LZjCX6_2(.din(w_dff_B_gtSv2GW19_2),.dout(w_dff_B_Rg2LZjCX6_2),.clk(gclk));
	jdff dff_B_6TEB4FEv0_2(.din(w_dff_B_Rg2LZjCX6_2),.dout(w_dff_B_6TEB4FEv0_2),.clk(gclk));
	jdff dff_B_KUz0OnNt7_1(.din(n967),.dout(w_dff_B_KUz0OnNt7_1),.clk(gclk));
	jdff dff_B_zYx6m8hr6_2(.din(n861),.dout(w_dff_B_zYx6m8hr6_2),.clk(gclk));
	jdff dff_B_KJ45VJJk2_2(.din(w_dff_B_zYx6m8hr6_2),.dout(w_dff_B_KJ45VJJk2_2),.clk(gclk));
	jdff dff_B_rMd0fbo21_2(.din(w_dff_B_KJ45VJJk2_2),.dout(w_dff_B_rMd0fbo21_2),.clk(gclk));
	jdff dff_B_hTmj3hb72_2(.din(w_dff_B_rMd0fbo21_2),.dout(w_dff_B_hTmj3hb72_2),.clk(gclk));
	jdff dff_B_amRdSPst1_2(.din(w_dff_B_hTmj3hb72_2),.dout(w_dff_B_amRdSPst1_2),.clk(gclk));
	jdff dff_B_PngaMlZc3_2(.din(w_dff_B_amRdSPst1_2),.dout(w_dff_B_PngaMlZc3_2),.clk(gclk));
	jdff dff_B_m9iKnzeW7_2(.din(w_dff_B_PngaMlZc3_2),.dout(w_dff_B_m9iKnzeW7_2),.clk(gclk));
	jdff dff_B_8wm29cfb6_2(.din(w_dff_B_m9iKnzeW7_2),.dout(w_dff_B_8wm29cfb6_2),.clk(gclk));
	jdff dff_B_9A9bssQh9_2(.din(w_dff_B_8wm29cfb6_2),.dout(w_dff_B_9A9bssQh9_2),.clk(gclk));
	jdff dff_B_elLOdBSp8_2(.din(w_dff_B_9A9bssQh9_2),.dout(w_dff_B_elLOdBSp8_2),.clk(gclk));
	jdff dff_B_Ir5SK7Ew5_2(.din(w_dff_B_elLOdBSp8_2),.dout(w_dff_B_Ir5SK7Ew5_2),.clk(gclk));
	jdff dff_B_UKXmqFIy2_2(.din(w_dff_B_Ir5SK7Ew5_2),.dout(w_dff_B_UKXmqFIy2_2),.clk(gclk));
	jdff dff_B_xwBRuEfy2_2(.din(w_dff_B_UKXmqFIy2_2),.dout(w_dff_B_xwBRuEfy2_2),.clk(gclk));
	jdff dff_B_BvPfyuBF3_2(.din(w_dff_B_xwBRuEfy2_2),.dout(w_dff_B_BvPfyuBF3_2),.clk(gclk));
	jdff dff_B_W5BkA0uv6_2(.din(w_dff_B_BvPfyuBF3_2),.dout(w_dff_B_W5BkA0uv6_2),.clk(gclk));
	jdff dff_B_GH7L05Zu3_2(.din(w_dff_B_W5BkA0uv6_2),.dout(w_dff_B_GH7L05Zu3_2),.clk(gclk));
	jdff dff_B_mHCpiLTu7_2(.din(w_dff_B_GH7L05Zu3_2),.dout(w_dff_B_mHCpiLTu7_2),.clk(gclk));
	jdff dff_B_BMw3Lxb49_2(.din(w_dff_B_mHCpiLTu7_2),.dout(w_dff_B_BMw3Lxb49_2),.clk(gclk));
	jdff dff_B_v6EO7e6d1_1(.din(n862),.dout(w_dff_B_v6EO7e6d1_1),.clk(gclk));
	jdff dff_B_7K2fZRS23_2(.din(n762),.dout(w_dff_B_7K2fZRS23_2),.clk(gclk));
	jdff dff_B_6j2iQjyc0_2(.din(w_dff_B_7K2fZRS23_2),.dout(w_dff_B_6j2iQjyc0_2),.clk(gclk));
	jdff dff_B_f2b3cNxg9_2(.din(w_dff_B_6j2iQjyc0_2),.dout(w_dff_B_f2b3cNxg9_2),.clk(gclk));
	jdff dff_B_4F8rAj4L9_2(.din(w_dff_B_f2b3cNxg9_2),.dout(w_dff_B_4F8rAj4L9_2),.clk(gclk));
	jdff dff_B_fr6qZNO09_2(.din(w_dff_B_4F8rAj4L9_2),.dout(w_dff_B_fr6qZNO09_2),.clk(gclk));
	jdff dff_B_NHqH9jy45_2(.din(w_dff_B_fr6qZNO09_2),.dout(w_dff_B_NHqH9jy45_2),.clk(gclk));
	jdff dff_B_OOltNCmH7_2(.din(w_dff_B_NHqH9jy45_2),.dout(w_dff_B_OOltNCmH7_2),.clk(gclk));
	jdff dff_B_9sGK2Dko4_2(.din(w_dff_B_OOltNCmH7_2),.dout(w_dff_B_9sGK2Dko4_2),.clk(gclk));
	jdff dff_B_QUELZei44_2(.din(w_dff_B_9sGK2Dko4_2),.dout(w_dff_B_QUELZei44_2),.clk(gclk));
	jdff dff_B_9h4a05Wh0_2(.din(w_dff_B_QUELZei44_2),.dout(w_dff_B_9h4a05Wh0_2),.clk(gclk));
	jdff dff_B_jdh6OKW50_2(.din(w_dff_B_9h4a05Wh0_2),.dout(w_dff_B_jdh6OKW50_2),.clk(gclk));
	jdff dff_B_B8W2kcWb2_2(.din(w_dff_B_jdh6OKW50_2),.dout(w_dff_B_B8W2kcWb2_2),.clk(gclk));
	jdff dff_B_MEA3lOOF7_2(.din(w_dff_B_B8W2kcWb2_2),.dout(w_dff_B_MEA3lOOF7_2),.clk(gclk));
	jdff dff_B_k2xht5bT4_2(.din(w_dff_B_MEA3lOOF7_2),.dout(w_dff_B_k2xht5bT4_2),.clk(gclk));
	jdff dff_B_7TOama1m4_2(.din(w_dff_B_k2xht5bT4_2),.dout(w_dff_B_7TOama1m4_2),.clk(gclk));
	jdff dff_B_531w516D6_2(.din(w_dff_B_7TOama1m4_2),.dout(w_dff_B_531w516D6_2),.clk(gclk));
	jdff dff_B_g8b86Sln6_1(.din(n763),.dout(w_dff_B_g8b86Sln6_1),.clk(gclk));
	jdff dff_B_CX7Ltmiv3_2(.din(n669),.dout(w_dff_B_CX7Ltmiv3_2),.clk(gclk));
	jdff dff_B_tYpSwzCP7_2(.din(w_dff_B_CX7Ltmiv3_2),.dout(w_dff_B_tYpSwzCP7_2),.clk(gclk));
	jdff dff_B_kSltH5U88_2(.din(w_dff_B_tYpSwzCP7_2),.dout(w_dff_B_kSltH5U88_2),.clk(gclk));
	jdff dff_B_mDl3wRKA0_2(.din(w_dff_B_kSltH5U88_2),.dout(w_dff_B_mDl3wRKA0_2),.clk(gclk));
	jdff dff_B_wD5QUVQy1_2(.din(w_dff_B_mDl3wRKA0_2),.dout(w_dff_B_wD5QUVQy1_2),.clk(gclk));
	jdff dff_B_M3glYfEu9_2(.din(w_dff_B_wD5QUVQy1_2),.dout(w_dff_B_M3glYfEu9_2),.clk(gclk));
	jdff dff_B_yARmHfY21_2(.din(w_dff_B_M3glYfEu9_2),.dout(w_dff_B_yARmHfY21_2),.clk(gclk));
	jdff dff_B_FKyAMUxU3_2(.din(w_dff_B_yARmHfY21_2),.dout(w_dff_B_FKyAMUxU3_2),.clk(gclk));
	jdff dff_B_4mxO6BWl3_2(.din(w_dff_B_FKyAMUxU3_2),.dout(w_dff_B_4mxO6BWl3_2),.clk(gclk));
	jdff dff_B_OyqZG4w32_2(.din(w_dff_B_4mxO6BWl3_2),.dout(w_dff_B_OyqZG4w32_2),.clk(gclk));
	jdff dff_B_FtxjEmG28_2(.din(w_dff_B_OyqZG4w32_2),.dout(w_dff_B_FtxjEmG28_2),.clk(gclk));
	jdff dff_B_s2PqJ7iJ2_2(.din(w_dff_B_FtxjEmG28_2),.dout(w_dff_B_s2PqJ7iJ2_2),.clk(gclk));
	jdff dff_B_A6yDWUB58_2(.din(w_dff_B_s2PqJ7iJ2_2),.dout(w_dff_B_A6yDWUB58_2),.clk(gclk));
	jdff dff_B_fyCeKIlH9_2(.din(w_dff_B_A6yDWUB58_2),.dout(w_dff_B_fyCeKIlH9_2),.clk(gclk));
	jdff dff_B_sqlWpZ4B1_1(.din(n670),.dout(w_dff_B_sqlWpZ4B1_1),.clk(gclk));
	jdff dff_B_ZtSnJRsu1_2(.din(n583),.dout(w_dff_B_ZtSnJRsu1_2),.clk(gclk));
	jdff dff_B_TkVc8CnX4_2(.din(w_dff_B_ZtSnJRsu1_2),.dout(w_dff_B_TkVc8CnX4_2),.clk(gclk));
	jdff dff_B_0dQqA2ul3_2(.din(w_dff_B_TkVc8CnX4_2),.dout(w_dff_B_0dQqA2ul3_2),.clk(gclk));
	jdff dff_B_U00cK3hr9_2(.din(w_dff_B_0dQqA2ul3_2),.dout(w_dff_B_U00cK3hr9_2),.clk(gclk));
	jdff dff_B_Ar4dDLoa9_2(.din(w_dff_B_U00cK3hr9_2),.dout(w_dff_B_Ar4dDLoa9_2),.clk(gclk));
	jdff dff_B_68Tvh88u8_2(.din(w_dff_B_Ar4dDLoa9_2),.dout(w_dff_B_68Tvh88u8_2),.clk(gclk));
	jdff dff_B_mgjrZIJX6_2(.din(w_dff_B_68Tvh88u8_2),.dout(w_dff_B_mgjrZIJX6_2),.clk(gclk));
	jdff dff_B_NSlQta5W2_2(.din(w_dff_B_mgjrZIJX6_2),.dout(w_dff_B_NSlQta5W2_2),.clk(gclk));
	jdff dff_B_DARwgzxd6_2(.din(w_dff_B_NSlQta5W2_2),.dout(w_dff_B_DARwgzxd6_2),.clk(gclk));
	jdff dff_B_F2GJ0d8h3_2(.din(w_dff_B_DARwgzxd6_2),.dout(w_dff_B_F2GJ0d8h3_2),.clk(gclk));
	jdff dff_B_CPUjbOtW5_2(.din(w_dff_B_F2GJ0d8h3_2),.dout(w_dff_B_CPUjbOtW5_2),.clk(gclk));
	jdff dff_B_CmZh1vkp5_2(.din(w_dff_B_CPUjbOtW5_2),.dout(w_dff_B_CmZh1vkp5_2),.clk(gclk));
	jdff dff_B_QPvjEvrN3_1(.din(n584),.dout(w_dff_B_QPvjEvrN3_1),.clk(gclk));
	jdff dff_B_yEoth6aF6_2(.din(n504),.dout(w_dff_B_yEoth6aF6_2),.clk(gclk));
	jdff dff_B_giZl3HEc0_2(.din(w_dff_B_yEoth6aF6_2),.dout(w_dff_B_giZl3HEc0_2),.clk(gclk));
	jdff dff_B_OhjmHqlE3_2(.din(w_dff_B_giZl3HEc0_2),.dout(w_dff_B_OhjmHqlE3_2),.clk(gclk));
	jdff dff_B_Ih6yjIAI0_2(.din(w_dff_B_OhjmHqlE3_2),.dout(w_dff_B_Ih6yjIAI0_2),.clk(gclk));
	jdff dff_B_q63G9MCO6_2(.din(w_dff_B_Ih6yjIAI0_2),.dout(w_dff_B_q63G9MCO6_2),.clk(gclk));
	jdff dff_B_u15dV6Ig2_2(.din(w_dff_B_q63G9MCO6_2),.dout(w_dff_B_u15dV6Ig2_2),.clk(gclk));
	jdff dff_B_d7wDfoEm9_2(.din(w_dff_B_u15dV6Ig2_2),.dout(w_dff_B_d7wDfoEm9_2),.clk(gclk));
	jdff dff_B_4bXUAm0L9_2(.din(w_dff_B_d7wDfoEm9_2),.dout(w_dff_B_4bXUAm0L9_2),.clk(gclk));
	jdff dff_B_tXKvlKa61_2(.din(w_dff_B_4bXUAm0L9_2),.dout(w_dff_B_tXKvlKa61_2),.clk(gclk));
	jdff dff_B_lKp0G3Gz6_2(.din(w_dff_B_tXKvlKa61_2),.dout(w_dff_B_lKp0G3Gz6_2),.clk(gclk));
	jdff dff_B_dl8ogSlE8_1(.din(n505),.dout(w_dff_B_dl8ogSlE8_1),.clk(gclk));
	jdff dff_B_Brc56l3K1_2(.din(n432),.dout(w_dff_B_Brc56l3K1_2),.clk(gclk));
	jdff dff_B_v1pP1J3C1_2(.din(w_dff_B_Brc56l3K1_2),.dout(w_dff_B_v1pP1J3C1_2),.clk(gclk));
	jdff dff_B_J7OPjAy74_2(.din(w_dff_B_v1pP1J3C1_2),.dout(w_dff_B_J7OPjAy74_2),.clk(gclk));
	jdff dff_B_6z5U1c8C8_2(.din(w_dff_B_J7OPjAy74_2),.dout(w_dff_B_6z5U1c8C8_2),.clk(gclk));
	jdff dff_B_QNofcxy58_2(.din(w_dff_B_6z5U1c8C8_2),.dout(w_dff_B_QNofcxy58_2),.clk(gclk));
	jdff dff_B_s9SmGu9L0_2(.din(w_dff_B_QNofcxy58_2),.dout(w_dff_B_s9SmGu9L0_2),.clk(gclk));
	jdff dff_B_9oCeouqO9_2(.din(w_dff_B_s9SmGu9L0_2),.dout(w_dff_B_9oCeouqO9_2),.clk(gclk));
	jdff dff_B_4f0QssU07_2(.din(w_dff_B_9oCeouqO9_2),.dout(w_dff_B_4f0QssU07_2),.clk(gclk));
	jdff dff_B_jVyz4aVK1_1(.din(n433),.dout(w_dff_B_jVyz4aVK1_1),.clk(gclk));
	jdff dff_B_ZpSHMSn91_2(.din(n368),.dout(w_dff_B_ZpSHMSn91_2),.clk(gclk));
	jdff dff_B_2juTzK0k2_2(.din(w_dff_B_ZpSHMSn91_2),.dout(w_dff_B_2juTzK0k2_2),.clk(gclk));
	jdff dff_B_jeIukxcj2_2(.din(w_dff_B_2juTzK0k2_2),.dout(w_dff_B_jeIukxcj2_2),.clk(gclk));
	jdff dff_B_J22aLDwg1_2(.din(w_dff_B_jeIukxcj2_2),.dout(w_dff_B_J22aLDwg1_2),.clk(gclk));
	jdff dff_B_TQ2jbAwY4_2(.din(w_dff_B_J22aLDwg1_2),.dout(w_dff_B_TQ2jbAwY4_2),.clk(gclk));
	jdff dff_B_2O4uTLYz9_2(.din(w_dff_B_TQ2jbAwY4_2),.dout(w_dff_B_2O4uTLYz9_2),.clk(gclk));
	jdff dff_B_xZpEN1Py9_2(.din(n383),.dout(w_dff_B_xZpEN1Py9_2),.clk(gclk));
	jdff dff_B_rYc5JrPE1_1(.din(n369),.dout(w_dff_B_rYc5JrPE1_1),.clk(gclk));
	jdff dff_B_YdACboNw3_1(.din(w_dff_B_rYc5JrPE1_1),.dout(w_dff_B_YdACboNw3_1),.clk(gclk));
	jdff dff_B_A58hShCc8_2(.din(n310),.dout(w_dff_B_A58hShCc8_2),.clk(gclk));
	jdff dff_B_pAXqnY8h2_2(.din(w_dff_B_A58hShCc8_2),.dout(w_dff_B_pAXqnY8h2_2),.clk(gclk));
	jdff dff_B_s4uNUbwG5_2(.din(w_dff_B_pAXqnY8h2_2),.dout(w_dff_B_s4uNUbwG5_2),.clk(gclk));
	jdff dff_B_dnWkgseM9_2(.din(w_dff_B_s4uNUbwG5_2),.dout(w_dff_B_dnWkgseM9_2),.clk(gclk));
	jdff dff_A_VcZH5Esl6_1(.dout(w_n317_0[1]),.din(w_dff_A_VcZH5Esl6_1),.clk(gclk));
	jdff dff_B_e9Y6sfxe4_1(.din(n312),.dout(w_dff_B_e9Y6sfxe4_1),.clk(gclk));
	jdff dff_B_1qBU2jhh6_1(.din(w_dff_B_e9Y6sfxe4_1),.dout(w_dff_B_1qBU2jhh6_1),.clk(gclk));
	jdff dff_A_skMxtdkH5_0(.dout(w_n258_0[0]),.din(w_dff_A_skMxtdkH5_0),.clk(gclk));
	jdff dff_A_sg2BvyBK1_1(.dout(w_n258_0[1]),.din(w_dff_A_sg2BvyBK1_1),.clk(gclk));
	jdff dff_A_8wznEIJ80_1(.dout(w_dff_A_sg2BvyBK1_1),.din(w_dff_A_8wznEIJ80_1),.clk(gclk));
	jdff dff_B_DExLKsan5_2(.din(n1565),.dout(w_dff_B_DExLKsan5_2),.clk(gclk));
	jdff dff_B_pZiXbu383_2(.din(w_dff_B_DExLKsan5_2),.dout(w_dff_B_pZiXbu383_2),.clk(gclk));
	jdff dff_B_Ha4dA8CP6_1(.din(n1563),.dout(w_dff_B_Ha4dA8CP6_1),.clk(gclk));
	jdff dff_B_MK926buB6_2(.din(n1497),.dout(w_dff_B_MK926buB6_2),.clk(gclk));
	jdff dff_B_R6zuIxg68_2(.din(w_dff_B_MK926buB6_2),.dout(w_dff_B_R6zuIxg68_2),.clk(gclk));
	jdff dff_B_xZphkrM66_2(.din(w_dff_B_R6zuIxg68_2),.dout(w_dff_B_xZphkrM66_2),.clk(gclk));
	jdff dff_B_QexdX6tn6_2(.din(w_dff_B_xZphkrM66_2),.dout(w_dff_B_QexdX6tn6_2),.clk(gclk));
	jdff dff_B_5OhqglfR9_2(.din(w_dff_B_QexdX6tn6_2),.dout(w_dff_B_5OhqglfR9_2),.clk(gclk));
	jdff dff_B_FSbp1kdf4_2(.din(w_dff_B_5OhqglfR9_2),.dout(w_dff_B_FSbp1kdf4_2),.clk(gclk));
	jdff dff_B_dDVTMdod0_2(.din(w_dff_B_FSbp1kdf4_2),.dout(w_dff_B_dDVTMdod0_2),.clk(gclk));
	jdff dff_B_L5UijDuh4_2(.din(w_dff_B_dDVTMdod0_2),.dout(w_dff_B_L5UijDuh4_2),.clk(gclk));
	jdff dff_B_ej23yrYe6_2(.din(w_dff_B_L5UijDuh4_2),.dout(w_dff_B_ej23yrYe6_2),.clk(gclk));
	jdff dff_B_KfLyFKoX3_2(.din(w_dff_B_ej23yrYe6_2),.dout(w_dff_B_KfLyFKoX3_2),.clk(gclk));
	jdff dff_B_EHuwfCyy0_2(.din(w_dff_B_KfLyFKoX3_2),.dout(w_dff_B_EHuwfCyy0_2),.clk(gclk));
	jdff dff_B_TiUYpoOm2_2(.din(w_dff_B_EHuwfCyy0_2),.dout(w_dff_B_TiUYpoOm2_2),.clk(gclk));
	jdff dff_B_sbjeyHi95_2(.din(w_dff_B_TiUYpoOm2_2),.dout(w_dff_B_sbjeyHi95_2),.clk(gclk));
	jdff dff_B_9x7PCOJT1_2(.din(w_dff_B_sbjeyHi95_2),.dout(w_dff_B_9x7PCOJT1_2),.clk(gclk));
	jdff dff_B_WRrAVpjx7_2(.din(w_dff_B_9x7PCOJT1_2),.dout(w_dff_B_WRrAVpjx7_2),.clk(gclk));
	jdff dff_B_FpsIhPoJ8_2(.din(w_dff_B_WRrAVpjx7_2),.dout(w_dff_B_FpsIhPoJ8_2),.clk(gclk));
	jdff dff_B_Eciu9rSA7_2(.din(w_dff_B_FpsIhPoJ8_2),.dout(w_dff_B_Eciu9rSA7_2),.clk(gclk));
	jdff dff_B_JDcuNnem2_2(.din(w_dff_B_Eciu9rSA7_2),.dout(w_dff_B_JDcuNnem2_2),.clk(gclk));
	jdff dff_B_GfA48xs63_2(.din(w_dff_B_JDcuNnem2_2),.dout(w_dff_B_GfA48xs63_2),.clk(gclk));
	jdff dff_B_dGjPk2uv4_2(.din(w_dff_B_GfA48xs63_2),.dout(w_dff_B_dGjPk2uv4_2),.clk(gclk));
	jdff dff_B_8ar8sJEJ5_2(.din(w_dff_B_dGjPk2uv4_2),.dout(w_dff_B_8ar8sJEJ5_2),.clk(gclk));
	jdff dff_B_Tx2FWoGG4_2(.din(w_dff_B_8ar8sJEJ5_2),.dout(w_dff_B_Tx2FWoGG4_2),.clk(gclk));
	jdff dff_B_BGoplHs33_2(.din(w_dff_B_Tx2FWoGG4_2),.dout(w_dff_B_BGoplHs33_2),.clk(gclk));
	jdff dff_B_G263SDlw2_2(.din(w_dff_B_BGoplHs33_2),.dout(w_dff_B_G263SDlw2_2),.clk(gclk));
	jdff dff_B_Ftj0OEKZ3_2(.din(w_dff_B_G263SDlw2_2),.dout(w_dff_B_Ftj0OEKZ3_2),.clk(gclk));
	jdff dff_B_0m1MsdC36_2(.din(w_dff_B_Ftj0OEKZ3_2),.dout(w_dff_B_0m1MsdC36_2),.clk(gclk));
	jdff dff_B_n3pEO8v07_2(.din(w_dff_B_0m1MsdC36_2),.dout(w_dff_B_n3pEO8v07_2),.clk(gclk));
	jdff dff_B_nJVjp2zy9_2(.din(w_dff_B_n3pEO8v07_2),.dout(w_dff_B_nJVjp2zy9_2),.clk(gclk));
	jdff dff_B_pFTCa8SU0_2(.din(w_dff_B_nJVjp2zy9_2),.dout(w_dff_B_pFTCa8SU0_2),.clk(gclk));
	jdff dff_B_x4F5fb0j9_2(.din(w_dff_B_pFTCa8SU0_2),.dout(w_dff_B_x4F5fb0j9_2),.clk(gclk));
	jdff dff_B_GN775u902_2(.din(w_dff_B_x4F5fb0j9_2),.dout(w_dff_B_GN775u902_2),.clk(gclk));
	jdff dff_B_kbZdJDio6_2(.din(w_dff_B_GN775u902_2),.dout(w_dff_B_kbZdJDio6_2),.clk(gclk));
	jdff dff_B_xXRxls5d9_2(.din(w_dff_B_kbZdJDio6_2),.dout(w_dff_B_xXRxls5d9_2),.clk(gclk));
	jdff dff_B_LFHM66KT6_2(.din(w_dff_B_xXRxls5d9_2),.dout(w_dff_B_LFHM66KT6_2),.clk(gclk));
	jdff dff_B_YvgYwXpD7_2(.din(w_dff_B_LFHM66KT6_2),.dout(w_dff_B_YvgYwXpD7_2),.clk(gclk));
	jdff dff_B_BLKrYaMk7_2(.din(w_dff_B_YvgYwXpD7_2),.dout(w_dff_B_BLKrYaMk7_2),.clk(gclk));
	jdff dff_B_8MAZy0s30_2(.din(w_dff_B_BLKrYaMk7_2),.dout(w_dff_B_8MAZy0s30_2),.clk(gclk));
	jdff dff_B_GjvakE6n3_2(.din(w_dff_B_8MAZy0s30_2),.dout(w_dff_B_GjvakE6n3_2),.clk(gclk));
	jdff dff_B_d35o9utC8_1(.din(n1561),.dout(w_dff_B_d35o9utC8_1),.clk(gclk));
	jdff dff_A_lLOzs8437_1(.dout(w_n1500_0[1]),.din(w_dff_A_lLOzs8437_1),.clk(gclk));
	jdff dff_B_mFNHx6He1_1(.din(n1498),.dout(w_dff_B_mFNHx6He1_1),.clk(gclk));
	jdff dff_B_M6OkMOFi3_2(.din(n1426),.dout(w_dff_B_M6OkMOFi3_2),.clk(gclk));
	jdff dff_B_Lk0Ern2v1_2(.din(w_dff_B_M6OkMOFi3_2),.dout(w_dff_B_Lk0Ern2v1_2),.clk(gclk));
	jdff dff_B_l7GvpiWy7_2(.din(w_dff_B_Lk0Ern2v1_2),.dout(w_dff_B_l7GvpiWy7_2),.clk(gclk));
	jdff dff_B_zCWGqkxA6_2(.din(w_dff_B_l7GvpiWy7_2),.dout(w_dff_B_zCWGqkxA6_2),.clk(gclk));
	jdff dff_B_wxPiLBOk4_2(.din(w_dff_B_zCWGqkxA6_2),.dout(w_dff_B_wxPiLBOk4_2),.clk(gclk));
	jdff dff_B_RUmcQ1o01_2(.din(w_dff_B_wxPiLBOk4_2),.dout(w_dff_B_RUmcQ1o01_2),.clk(gclk));
	jdff dff_B_0uzAax8D3_2(.din(w_dff_B_RUmcQ1o01_2),.dout(w_dff_B_0uzAax8D3_2),.clk(gclk));
	jdff dff_B_DFTkswCf8_2(.din(w_dff_B_0uzAax8D3_2),.dout(w_dff_B_DFTkswCf8_2),.clk(gclk));
	jdff dff_B_tWpstZeL1_2(.din(w_dff_B_DFTkswCf8_2),.dout(w_dff_B_tWpstZeL1_2),.clk(gclk));
	jdff dff_B_lYvgkDur0_2(.din(w_dff_B_tWpstZeL1_2),.dout(w_dff_B_lYvgkDur0_2),.clk(gclk));
	jdff dff_B_oSR7azdG1_2(.din(w_dff_B_lYvgkDur0_2),.dout(w_dff_B_oSR7azdG1_2),.clk(gclk));
	jdff dff_B_cJaitoE09_2(.din(w_dff_B_oSR7azdG1_2),.dout(w_dff_B_cJaitoE09_2),.clk(gclk));
	jdff dff_B_4cDCKpr24_2(.din(w_dff_B_cJaitoE09_2),.dout(w_dff_B_4cDCKpr24_2),.clk(gclk));
	jdff dff_B_mzH3WjKv8_2(.din(w_dff_B_4cDCKpr24_2),.dout(w_dff_B_mzH3WjKv8_2),.clk(gclk));
	jdff dff_B_mqHUsab91_2(.din(w_dff_B_mzH3WjKv8_2),.dout(w_dff_B_mqHUsab91_2),.clk(gclk));
	jdff dff_B_4Q4iHfYy6_2(.din(w_dff_B_mqHUsab91_2),.dout(w_dff_B_4Q4iHfYy6_2),.clk(gclk));
	jdff dff_B_89uiv0Ei0_2(.din(w_dff_B_4Q4iHfYy6_2),.dout(w_dff_B_89uiv0Ei0_2),.clk(gclk));
	jdff dff_B_x2PUERo15_2(.din(w_dff_B_89uiv0Ei0_2),.dout(w_dff_B_x2PUERo15_2),.clk(gclk));
	jdff dff_B_NyftFSa39_2(.din(w_dff_B_x2PUERo15_2),.dout(w_dff_B_NyftFSa39_2),.clk(gclk));
	jdff dff_B_ROyZ1ODi7_2(.din(w_dff_B_NyftFSa39_2),.dout(w_dff_B_ROyZ1ODi7_2),.clk(gclk));
	jdff dff_B_27uVoUy08_2(.din(w_dff_B_ROyZ1ODi7_2),.dout(w_dff_B_27uVoUy08_2),.clk(gclk));
	jdff dff_B_iF0Q8r5y4_2(.din(w_dff_B_27uVoUy08_2),.dout(w_dff_B_iF0Q8r5y4_2),.clk(gclk));
	jdff dff_B_0L4tKxqg7_2(.din(w_dff_B_iF0Q8r5y4_2),.dout(w_dff_B_0L4tKxqg7_2),.clk(gclk));
	jdff dff_B_FRHv0RZz6_2(.din(w_dff_B_0L4tKxqg7_2),.dout(w_dff_B_FRHv0RZz6_2),.clk(gclk));
	jdff dff_B_YiHSCAt07_2(.din(w_dff_B_FRHv0RZz6_2),.dout(w_dff_B_YiHSCAt07_2),.clk(gclk));
	jdff dff_B_H9ZunKdY0_2(.din(w_dff_B_YiHSCAt07_2),.dout(w_dff_B_H9ZunKdY0_2),.clk(gclk));
	jdff dff_B_8vBf2JKc0_2(.din(w_dff_B_H9ZunKdY0_2),.dout(w_dff_B_8vBf2JKc0_2),.clk(gclk));
	jdff dff_B_F8ORJLhT7_2(.din(w_dff_B_8vBf2JKc0_2),.dout(w_dff_B_F8ORJLhT7_2),.clk(gclk));
	jdff dff_B_kyjDQxZT6_2(.din(w_dff_B_F8ORJLhT7_2),.dout(w_dff_B_kyjDQxZT6_2),.clk(gclk));
	jdff dff_B_JvFmRFZb9_2(.din(w_dff_B_kyjDQxZT6_2),.dout(w_dff_B_JvFmRFZb9_2),.clk(gclk));
	jdff dff_B_yp2Jug5Y8_2(.din(w_dff_B_JvFmRFZb9_2),.dout(w_dff_B_yp2Jug5Y8_2),.clk(gclk));
	jdff dff_B_YviWvkZ03_2(.din(w_dff_B_yp2Jug5Y8_2),.dout(w_dff_B_YviWvkZ03_2),.clk(gclk));
	jdff dff_B_NOISaytV5_2(.din(w_dff_B_YviWvkZ03_2),.dout(w_dff_B_NOISaytV5_2),.clk(gclk));
	jdff dff_B_6w8IAF025_2(.din(n1429),.dout(w_dff_B_6w8IAF025_2),.clk(gclk));
	jdff dff_B_PkKGRpPN5_1(.din(n1427),.dout(w_dff_B_PkKGRpPN5_1),.clk(gclk));
	jdff dff_B_PliDiHTF5_2(.din(n1348),.dout(w_dff_B_PliDiHTF5_2),.clk(gclk));
	jdff dff_B_kWXhzVmt0_2(.din(w_dff_B_PliDiHTF5_2),.dout(w_dff_B_kWXhzVmt0_2),.clk(gclk));
	jdff dff_B_1fsV6qV82_2(.din(w_dff_B_kWXhzVmt0_2),.dout(w_dff_B_1fsV6qV82_2),.clk(gclk));
	jdff dff_B_Ma50OG3U1_2(.din(w_dff_B_1fsV6qV82_2),.dout(w_dff_B_Ma50OG3U1_2),.clk(gclk));
	jdff dff_B_Sljro1Zy7_2(.din(w_dff_B_Ma50OG3U1_2),.dout(w_dff_B_Sljro1Zy7_2),.clk(gclk));
	jdff dff_B_RwzDse3h8_2(.din(w_dff_B_Sljro1Zy7_2),.dout(w_dff_B_RwzDse3h8_2),.clk(gclk));
	jdff dff_B_lroheoqH4_2(.din(w_dff_B_RwzDse3h8_2),.dout(w_dff_B_lroheoqH4_2),.clk(gclk));
	jdff dff_B_M4Ftwh446_2(.din(w_dff_B_lroheoqH4_2),.dout(w_dff_B_M4Ftwh446_2),.clk(gclk));
	jdff dff_B_3XmlgQfQ5_2(.din(w_dff_B_M4Ftwh446_2),.dout(w_dff_B_3XmlgQfQ5_2),.clk(gclk));
	jdff dff_B_59yEYbnS4_2(.din(w_dff_B_3XmlgQfQ5_2),.dout(w_dff_B_59yEYbnS4_2),.clk(gclk));
	jdff dff_B_JFJO1CNx0_2(.din(w_dff_B_59yEYbnS4_2),.dout(w_dff_B_JFJO1CNx0_2),.clk(gclk));
	jdff dff_B_1Go9Z96e3_2(.din(w_dff_B_JFJO1CNx0_2),.dout(w_dff_B_1Go9Z96e3_2),.clk(gclk));
	jdff dff_B_zWv3JliJ1_2(.din(w_dff_B_1Go9Z96e3_2),.dout(w_dff_B_zWv3JliJ1_2),.clk(gclk));
	jdff dff_B_Xqv6Q7457_2(.din(w_dff_B_zWv3JliJ1_2),.dout(w_dff_B_Xqv6Q7457_2),.clk(gclk));
	jdff dff_B_4bcsZa5X9_2(.din(w_dff_B_Xqv6Q7457_2),.dout(w_dff_B_4bcsZa5X9_2),.clk(gclk));
	jdff dff_B_4fgELMmN9_2(.din(w_dff_B_4bcsZa5X9_2),.dout(w_dff_B_4fgELMmN9_2),.clk(gclk));
	jdff dff_B_SPclwaLV7_2(.din(w_dff_B_4fgELMmN9_2),.dout(w_dff_B_SPclwaLV7_2),.clk(gclk));
	jdff dff_B_3Jqw9cmH6_2(.din(w_dff_B_SPclwaLV7_2),.dout(w_dff_B_3Jqw9cmH6_2),.clk(gclk));
	jdff dff_B_60k9XGYn7_2(.din(w_dff_B_3Jqw9cmH6_2),.dout(w_dff_B_60k9XGYn7_2),.clk(gclk));
	jdff dff_B_eXQKReoR1_2(.din(w_dff_B_60k9XGYn7_2),.dout(w_dff_B_eXQKReoR1_2),.clk(gclk));
	jdff dff_B_VCaaGmXz3_2(.din(w_dff_B_eXQKReoR1_2),.dout(w_dff_B_VCaaGmXz3_2),.clk(gclk));
	jdff dff_B_QNeD0R4d5_2(.din(w_dff_B_VCaaGmXz3_2),.dout(w_dff_B_QNeD0R4d5_2),.clk(gclk));
	jdff dff_B_wMCwo19D5_2(.din(w_dff_B_QNeD0R4d5_2),.dout(w_dff_B_wMCwo19D5_2),.clk(gclk));
	jdff dff_B_h6mzTWY73_2(.din(w_dff_B_wMCwo19D5_2),.dout(w_dff_B_h6mzTWY73_2),.clk(gclk));
	jdff dff_B_MGyxqxl27_2(.din(w_dff_B_h6mzTWY73_2),.dout(w_dff_B_MGyxqxl27_2),.clk(gclk));
	jdff dff_B_oUFAa6B86_2(.din(w_dff_B_MGyxqxl27_2),.dout(w_dff_B_oUFAa6B86_2),.clk(gclk));
	jdff dff_B_fLJ3mFif7_2(.din(w_dff_B_oUFAa6B86_2),.dout(w_dff_B_fLJ3mFif7_2),.clk(gclk));
	jdff dff_B_SUlQUeiM2_2(.din(w_dff_B_fLJ3mFif7_2),.dout(w_dff_B_SUlQUeiM2_2),.clk(gclk));
	jdff dff_B_OR7k9PM48_2(.din(w_dff_B_SUlQUeiM2_2),.dout(w_dff_B_OR7k9PM48_2),.clk(gclk));
	jdff dff_B_rsbKbUpA0_2(.din(w_dff_B_OR7k9PM48_2),.dout(w_dff_B_rsbKbUpA0_2),.clk(gclk));
	jdff dff_B_chs9YUMz7_2(.din(n1351),.dout(w_dff_B_chs9YUMz7_2),.clk(gclk));
	jdff dff_B_y4LofFOP8_1(.din(n1349),.dout(w_dff_B_y4LofFOP8_1),.clk(gclk));
	jdff dff_B_E9L57k8p4_2(.din(n1263),.dout(w_dff_B_E9L57k8p4_2),.clk(gclk));
	jdff dff_B_h6VIM8T74_2(.din(w_dff_B_E9L57k8p4_2),.dout(w_dff_B_h6VIM8T74_2),.clk(gclk));
	jdff dff_B_YXnXG3sv8_2(.din(w_dff_B_h6VIM8T74_2),.dout(w_dff_B_YXnXG3sv8_2),.clk(gclk));
	jdff dff_B_qn7w44uf3_2(.din(w_dff_B_YXnXG3sv8_2),.dout(w_dff_B_qn7w44uf3_2),.clk(gclk));
	jdff dff_B_p70eb7q74_2(.din(w_dff_B_qn7w44uf3_2),.dout(w_dff_B_p70eb7q74_2),.clk(gclk));
	jdff dff_B_tun9RBeK1_2(.din(w_dff_B_p70eb7q74_2),.dout(w_dff_B_tun9RBeK1_2),.clk(gclk));
	jdff dff_B_l7Md8jEx6_2(.din(w_dff_B_tun9RBeK1_2),.dout(w_dff_B_l7Md8jEx6_2),.clk(gclk));
	jdff dff_B_EzdPAXDg4_2(.din(w_dff_B_l7Md8jEx6_2),.dout(w_dff_B_EzdPAXDg4_2),.clk(gclk));
	jdff dff_B_cE7u32Im9_2(.din(w_dff_B_EzdPAXDg4_2),.dout(w_dff_B_cE7u32Im9_2),.clk(gclk));
	jdff dff_B_fcCGa3yA4_2(.din(w_dff_B_cE7u32Im9_2),.dout(w_dff_B_fcCGa3yA4_2),.clk(gclk));
	jdff dff_B_9TCNCdbG3_2(.din(w_dff_B_fcCGa3yA4_2),.dout(w_dff_B_9TCNCdbG3_2),.clk(gclk));
	jdff dff_B_9OIgVnGx2_2(.din(w_dff_B_9TCNCdbG3_2),.dout(w_dff_B_9OIgVnGx2_2),.clk(gclk));
	jdff dff_B_JEIUrNoe7_2(.din(w_dff_B_9OIgVnGx2_2),.dout(w_dff_B_JEIUrNoe7_2),.clk(gclk));
	jdff dff_B_AQxarMdi8_2(.din(w_dff_B_JEIUrNoe7_2),.dout(w_dff_B_AQxarMdi8_2),.clk(gclk));
	jdff dff_B_p80LeQ700_2(.din(w_dff_B_AQxarMdi8_2),.dout(w_dff_B_p80LeQ700_2),.clk(gclk));
	jdff dff_B_U1qPqupJ1_2(.din(w_dff_B_p80LeQ700_2),.dout(w_dff_B_U1qPqupJ1_2),.clk(gclk));
	jdff dff_B_NzaRCKDZ9_2(.din(w_dff_B_U1qPqupJ1_2),.dout(w_dff_B_NzaRCKDZ9_2),.clk(gclk));
	jdff dff_B_F1NjqyrD3_2(.din(w_dff_B_NzaRCKDZ9_2),.dout(w_dff_B_F1NjqyrD3_2),.clk(gclk));
	jdff dff_B_lhwUwXQC5_2(.din(w_dff_B_F1NjqyrD3_2),.dout(w_dff_B_lhwUwXQC5_2),.clk(gclk));
	jdff dff_B_9tzFCHfh5_2(.din(w_dff_B_lhwUwXQC5_2),.dout(w_dff_B_9tzFCHfh5_2),.clk(gclk));
	jdff dff_B_DZAcQQot6_2(.din(w_dff_B_9tzFCHfh5_2),.dout(w_dff_B_DZAcQQot6_2),.clk(gclk));
	jdff dff_B_1ZlTv62G8_2(.din(w_dff_B_DZAcQQot6_2),.dout(w_dff_B_1ZlTv62G8_2),.clk(gclk));
	jdff dff_B_oVmvi1404_2(.din(w_dff_B_1ZlTv62G8_2),.dout(w_dff_B_oVmvi1404_2),.clk(gclk));
	jdff dff_B_FdyllLGU0_2(.din(w_dff_B_oVmvi1404_2),.dout(w_dff_B_FdyllLGU0_2),.clk(gclk));
	jdff dff_B_o7DYz6aA3_2(.din(w_dff_B_FdyllLGU0_2),.dout(w_dff_B_o7DYz6aA3_2),.clk(gclk));
	jdff dff_B_D0WC8Jrt7_2(.din(w_dff_B_o7DYz6aA3_2),.dout(w_dff_B_D0WC8Jrt7_2),.clk(gclk));
	jdff dff_B_RpWXsmZk5_2(.din(w_dff_B_D0WC8Jrt7_2),.dout(w_dff_B_RpWXsmZk5_2),.clk(gclk));
	jdff dff_B_aDoAwMgG7_2(.din(n1266),.dout(w_dff_B_aDoAwMgG7_2),.clk(gclk));
	jdff dff_B_ppPcRfFc9_1(.din(n1264),.dout(w_dff_B_ppPcRfFc9_1),.clk(gclk));
	jdff dff_B_Ts4Q0cMs5_2(.din(n1173),.dout(w_dff_B_Ts4Q0cMs5_2),.clk(gclk));
	jdff dff_B_meOfJaf41_2(.din(w_dff_B_Ts4Q0cMs5_2),.dout(w_dff_B_meOfJaf41_2),.clk(gclk));
	jdff dff_B_5a5NhNRy2_2(.din(w_dff_B_meOfJaf41_2),.dout(w_dff_B_5a5NhNRy2_2),.clk(gclk));
	jdff dff_B_TMshmf287_2(.din(w_dff_B_5a5NhNRy2_2),.dout(w_dff_B_TMshmf287_2),.clk(gclk));
	jdff dff_B_uvL8JNmW4_2(.din(w_dff_B_TMshmf287_2),.dout(w_dff_B_uvL8JNmW4_2),.clk(gclk));
	jdff dff_B_GhrSfGCU3_2(.din(w_dff_B_uvL8JNmW4_2),.dout(w_dff_B_GhrSfGCU3_2),.clk(gclk));
	jdff dff_B_whNCTC1c4_2(.din(w_dff_B_GhrSfGCU3_2),.dout(w_dff_B_whNCTC1c4_2),.clk(gclk));
	jdff dff_B_M4fEIXqe1_2(.din(w_dff_B_whNCTC1c4_2),.dout(w_dff_B_M4fEIXqe1_2),.clk(gclk));
	jdff dff_B_ojp2PRcz5_2(.din(w_dff_B_M4fEIXqe1_2),.dout(w_dff_B_ojp2PRcz5_2),.clk(gclk));
	jdff dff_B_4rW8kF436_2(.din(w_dff_B_ojp2PRcz5_2),.dout(w_dff_B_4rW8kF436_2),.clk(gclk));
	jdff dff_B_MrBC4i2M5_2(.din(w_dff_B_4rW8kF436_2),.dout(w_dff_B_MrBC4i2M5_2),.clk(gclk));
	jdff dff_B_V1HKmQ0i2_2(.din(w_dff_B_MrBC4i2M5_2),.dout(w_dff_B_V1HKmQ0i2_2),.clk(gclk));
	jdff dff_B_JMJMF9Th4_2(.din(w_dff_B_V1HKmQ0i2_2),.dout(w_dff_B_JMJMF9Th4_2),.clk(gclk));
	jdff dff_B_63l4kO8P4_2(.din(w_dff_B_JMJMF9Th4_2),.dout(w_dff_B_63l4kO8P4_2),.clk(gclk));
	jdff dff_B_OySR4rAB3_2(.din(w_dff_B_63l4kO8P4_2),.dout(w_dff_B_OySR4rAB3_2),.clk(gclk));
	jdff dff_B_jtj6jdjk9_2(.din(w_dff_B_OySR4rAB3_2),.dout(w_dff_B_jtj6jdjk9_2),.clk(gclk));
	jdff dff_B_y9yVm9JD1_2(.din(w_dff_B_jtj6jdjk9_2),.dout(w_dff_B_y9yVm9JD1_2),.clk(gclk));
	jdff dff_B_rqqcDBgj1_2(.din(w_dff_B_y9yVm9JD1_2),.dout(w_dff_B_rqqcDBgj1_2),.clk(gclk));
	jdff dff_B_PULExbZ77_2(.din(w_dff_B_rqqcDBgj1_2),.dout(w_dff_B_PULExbZ77_2),.clk(gclk));
	jdff dff_B_jXIKAYn04_2(.din(w_dff_B_PULExbZ77_2),.dout(w_dff_B_jXIKAYn04_2),.clk(gclk));
	jdff dff_B_GflnDjUS4_2(.din(w_dff_B_jXIKAYn04_2),.dout(w_dff_B_GflnDjUS4_2),.clk(gclk));
	jdff dff_B_b5PExdQZ9_2(.din(w_dff_B_GflnDjUS4_2),.dout(w_dff_B_b5PExdQZ9_2),.clk(gclk));
	jdff dff_B_qxazGri21_2(.din(w_dff_B_b5PExdQZ9_2),.dout(w_dff_B_qxazGri21_2),.clk(gclk));
	jdff dff_B_mmbLPHoG8_2(.din(w_dff_B_qxazGri21_2),.dout(w_dff_B_mmbLPHoG8_2),.clk(gclk));
	jdff dff_B_kZA6OXJq2_2(.din(n1176),.dout(w_dff_B_kZA6OXJq2_2),.clk(gclk));
	jdff dff_B_m3XPCPsF9_1(.din(n1174),.dout(w_dff_B_m3XPCPsF9_1),.clk(gclk));
	jdff dff_B_NE20FSM95_2(.din(n1069),.dout(w_dff_B_NE20FSM95_2),.clk(gclk));
	jdff dff_B_9KkvwDLF1_2(.din(w_dff_B_NE20FSM95_2),.dout(w_dff_B_9KkvwDLF1_2),.clk(gclk));
	jdff dff_B_4KqldsYg2_2(.din(w_dff_B_9KkvwDLF1_2),.dout(w_dff_B_4KqldsYg2_2),.clk(gclk));
	jdff dff_B_ABJrZuSc0_2(.din(w_dff_B_4KqldsYg2_2),.dout(w_dff_B_ABJrZuSc0_2),.clk(gclk));
	jdff dff_B_69rUXBt77_2(.din(w_dff_B_ABJrZuSc0_2),.dout(w_dff_B_69rUXBt77_2),.clk(gclk));
	jdff dff_B_QUpLqKIj1_2(.din(w_dff_B_69rUXBt77_2),.dout(w_dff_B_QUpLqKIj1_2),.clk(gclk));
	jdff dff_B_Hw2y83XZ8_2(.din(w_dff_B_QUpLqKIj1_2),.dout(w_dff_B_Hw2y83XZ8_2),.clk(gclk));
	jdff dff_B_Q1Y3gqzV8_2(.din(w_dff_B_Hw2y83XZ8_2),.dout(w_dff_B_Q1Y3gqzV8_2),.clk(gclk));
	jdff dff_B_R9xoNTbM5_2(.din(w_dff_B_Q1Y3gqzV8_2),.dout(w_dff_B_R9xoNTbM5_2),.clk(gclk));
	jdff dff_B_297dIm7T1_2(.din(w_dff_B_R9xoNTbM5_2),.dout(w_dff_B_297dIm7T1_2),.clk(gclk));
	jdff dff_B_G8uTXr1V5_2(.din(w_dff_B_297dIm7T1_2),.dout(w_dff_B_G8uTXr1V5_2),.clk(gclk));
	jdff dff_B_hRDYlOWn6_2(.din(w_dff_B_G8uTXr1V5_2),.dout(w_dff_B_hRDYlOWn6_2),.clk(gclk));
	jdff dff_B_Lblrt5vK7_2(.din(w_dff_B_hRDYlOWn6_2),.dout(w_dff_B_Lblrt5vK7_2),.clk(gclk));
	jdff dff_B_AHGs0XeU3_2(.din(w_dff_B_Lblrt5vK7_2),.dout(w_dff_B_AHGs0XeU3_2),.clk(gclk));
	jdff dff_B_SmdO51gC2_2(.din(w_dff_B_AHGs0XeU3_2),.dout(w_dff_B_SmdO51gC2_2),.clk(gclk));
	jdff dff_B_pRq4ur5N6_2(.din(w_dff_B_SmdO51gC2_2),.dout(w_dff_B_pRq4ur5N6_2),.clk(gclk));
	jdff dff_B_nywyIp3O3_2(.din(w_dff_B_pRq4ur5N6_2),.dout(w_dff_B_nywyIp3O3_2),.clk(gclk));
	jdff dff_B_dzeT7FWG9_2(.din(w_dff_B_nywyIp3O3_2),.dout(w_dff_B_dzeT7FWG9_2),.clk(gclk));
	jdff dff_B_KZ5sjCly7_2(.din(w_dff_B_dzeT7FWG9_2),.dout(w_dff_B_KZ5sjCly7_2),.clk(gclk));
	jdff dff_B_wq8TGaBw9_2(.din(w_dff_B_KZ5sjCly7_2),.dout(w_dff_B_wq8TGaBw9_2),.clk(gclk));
	jdff dff_B_jLbPvk7S3_2(.din(w_dff_B_wq8TGaBw9_2),.dout(w_dff_B_jLbPvk7S3_2),.clk(gclk));
	jdff dff_B_PT0HtWut8_2(.din(n1072),.dout(w_dff_B_PT0HtWut8_2),.clk(gclk));
	jdff dff_B_LFD6220C1_1(.din(n1070),.dout(w_dff_B_LFD6220C1_1),.clk(gclk));
	jdff dff_B_192RJ2D25_2(.din(n971),.dout(w_dff_B_192RJ2D25_2),.clk(gclk));
	jdff dff_B_6tC0R6bB8_2(.din(w_dff_B_192RJ2D25_2),.dout(w_dff_B_6tC0R6bB8_2),.clk(gclk));
	jdff dff_B_0m1TzszK9_2(.din(w_dff_B_6tC0R6bB8_2),.dout(w_dff_B_0m1TzszK9_2),.clk(gclk));
	jdff dff_B_CGq9dzQb2_2(.din(w_dff_B_0m1TzszK9_2),.dout(w_dff_B_CGq9dzQb2_2),.clk(gclk));
	jdff dff_B_lK6ncWOJ1_2(.din(w_dff_B_CGq9dzQb2_2),.dout(w_dff_B_lK6ncWOJ1_2),.clk(gclk));
	jdff dff_B_Jj42eF2F1_2(.din(w_dff_B_lK6ncWOJ1_2),.dout(w_dff_B_Jj42eF2F1_2),.clk(gclk));
	jdff dff_B_vUeD3pRe1_2(.din(w_dff_B_Jj42eF2F1_2),.dout(w_dff_B_vUeD3pRe1_2),.clk(gclk));
	jdff dff_B_zcD1WgtR7_2(.din(w_dff_B_vUeD3pRe1_2),.dout(w_dff_B_zcD1WgtR7_2),.clk(gclk));
	jdff dff_B_ql4sEzOF1_2(.din(w_dff_B_zcD1WgtR7_2),.dout(w_dff_B_ql4sEzOF1_2),.clk(gclk));
	jdff dff_B_QwxvYzoF6_2(.din(w_dff_B_ql4sEzOF1_2),.dout(w_dff_B_QwxvYzoF6_2),.clk(gclk));
	jdff dff_B_HB8TFIOu8_2(.din(w_dff_B_QwxvYzoF6_2),.dout(w_dff_B_HB8TFIOu8_2),.clk(gclk));
	jdff dff_B_9AmG9lX73_2(.din(w_dff_B_HB8TFIOu8_2),.dout(w_dff_B_9AmG9lX73_2),.clk(gclk));
	jdff dff_B_2FUhEZFg2_2(.din(w_dff_B_9AmG9lX73_2),.dout(w_dff_B_2FUhEZFg2_2),.clk(gclk));
	jdff dff_B_UpF9gtnx1_2(.din(w_dff_B_2FUhEZFg2_2),.dout(w_dff_B_UpF9gtnx1_2),.clk(gclk));
	jdff dff_B_UJjaStq72_2(.din(w_dff_B_UpF9gtnx1_2),.dout(w_dff_B_UJjaStq72_2),.clk(gclk));
	jdff dff_B_qr3wr1s50_2(.din(w_dff_B_UJjaStq72_2),.dout(w_dff_B_qr3wr1s50_2),.clk(gclk));
	jdff dff_B_FQR6UAjT8_2(.din(w_dff_B_qr3wr1s50_2),.dout(w_dff_B_FQR6UAjT8_2),.clk(gclk));
	jdff dff_B_yGnZ6wXe5_2(.din(w_dff_B_FQR6UAjT8_2),.dout(w_dff_B_yGnZ6wXe5_2),.clk(gclk));
	jdff dff_B_yxOlFviZ9_1(.din(n972),.dout(w_dff_B_yxOlFviZ9_1),.clk(gclk));
	jdff dff_B_lTUeQ3Ie8_2(.din(n866),.dout(w_dff_B_lTUeQ3Ie8_2),.clk(gclk));
	jdff dff_B_SiLwA4z37_2(.din(w_dff_B_lTUeQ3Ie8_2),.dout(w_dff_B_SiLwA4z37_2),.clk(gclk));
	jdff dff_B_Dbxf7ptV3_2(.din(w_dff_B_SiLwA4z37_2),.dout(w_dff_B_Dbxf7ptV3_2),.clk(gclk));
	jdff dff_B_MwkCO1nP0_2(.din(w_dff_B_Dbxf7ptV3_2),.dout(w_dff_B_MwkCO1nP0_2),.clk(gclk));
	jdff dff_B_ADSSVMpC1_2(.din(w_dff_B_MwkCO1nP0_2),.dout(w_dff_B_ADSSVMpC1_2),.clk(gclk));
	jdff dff_B_kmmSPiV32_2(.din(w_dff_B_ADSSVMpC1_2),.dout(w_dff_B_kmmSPiV32_2),.clk(gclk));
	jdff dff_B_LOAHBBye1_2(.din(w_dff_B_kmmSPiV32_2),.dout(w_dff_B_LOAHBBye1_2),.clk(gclk));
	jdff dff_B_I3HO192n8_2(.din(w_dff_B_LOAHBBye1_2),.dout(w_dff_B_I3HO192n8_2),.clk(gclk));
	jdff dff_B_cFgzPVNV1_2(.din(w_dff_B_I3HO192n8_2),.dout(w_dff_B_cFgzPVNV1_2),.clk(gclk));
	jdff dff_B_mw6IXts98_2(.din(w_dff_B_cFgzPVNV1_2),.dout(w_dff_B_mw6IXts98_2),.clk(gclk));
	jdff dff_B_8lt01LFM9_2(.din(w_dff_B_mw6IXts98_2),.dout(w_dff_B_8lt01LFM9_2),.clk(gclk));
	jdff dff_B_BsrgxrED6_2(.din(w_dff_B_8lt01LFM9_2),.dout(w_dff_B_BsrgxrED6_2),.clk(gclk));
	jdff dff_B_X65kA0ky4_2(.din(w_dff_B_BsrgxrED6_2),.dout(w_dff_B_X65kA0ky4_2),.clk(gclk));
	jdff dff_B_uvbGGtbD5_2(.din(w_dff_B_X65kA0ky4_2),.dout(w_dff_B_uvbGGtbD5_2),.clk(gclk));
	jdff dff_B_W8bDkUIY1_2(.din(w_dff_B_uvbGGtbD5_2),.dout(w_dff_B_W8bDkUIY1_2),.clk(gclk));
	jdff dff_B_jPnbXJoN6_2(.din(w_dff_B_W8bDkUIY1_2),.dout(w_dff_B_jPnbXJoN6_2),.clk(gclk));
	jdff dff_B_YeF2aOoA8_1(.din(n867),.dout(w_dff_B_YeF2aOoA8_1),.clk(gclk));
	jdff dff_B_wubA050A5_2(.din(n767),.dout(w_dff_B_wubA050A5_2),.clk(gclk));
	jdff dff_B_BWComL7u2_2(.din(w_dff_B_wubA050A5_2),.dout(w_dff_B_BWComL7u2_2),.clk(gclk));
	jdff dff_B_a1EWwCsT7_2(.din(w_dff_B_BWComL7u2_2),.dout(w_dff_B_a1EWwCsT7_2),.clk(gclk));
	jdff dff_B_zziIjG450_2(.din(w_dff_B_a1EWwCsT7_2),.dout(w_dff_B_zziIjG450_2),.clk(gclk));
	jdff dff_B_cLeb0gH46_2(.din(w_dff_B_zziIjG450_2),.dout(w_dff_B_cLeb0gH46_2),.clk(gclk));
	jdff dff_B_al7182yJ5_2(.din(w_dff_B_cLeb0gH46_2),.dout(w_dff_B_al7182yJ5_2),.clk(gclk));
	jdff dff_B_cy3n8wFt3_2(.din(w_dff_B_al7182yJ5_2),.dout(w_dff_B_cy3n8wFt3_2),.clk(gclk));
	jdff dff_B_qcpxDavu7_2(.din(w_dff_B_cy3n8wFt3_2),.dout(w_dff_B_qcpxDavu7_2),.clk(gclk));
	jdff dff_B_VEfHnmUB9_2(.din(w_dff_B_qcpxDavu7_2),.dout(w_dff_B_VEfHnmUB9_2),.clk(gclk));
	jdff dff_B_Z7UGCT8t9_2(.din(w_dff_B_VEfHnmUB9_2),.dout(w_dff_B_Z7UGCT8t9_2),.clk(gclk));
	jdff dff_B_9Ao9geGd2_2(.din(w_dff_B_Z7UGCT8t9_2),.dout(w_dff_B_9Ao9geGd2_2),.clk(gclk));
	jdff dff_B_SxPerF1y7_2(.din(w_dff_B_9Ao9geGd2_2),.dout(w_dff_B_SxPerF1y7_2),.clk(gclk));
	jdff dff_B_eC0l1LTS3_2(.din(w_dff_B_SxPerF1y7_2),.dout(w_dff_B_eC0l1LTS3_2),.clk(gclk));
	jdff dff_B_1303sco78_2(.din(w_dff_B_eC0l1LTS3_2),.dout(w_dff_B_1303sco78_2),.clk(gclk));
	jdff dff_B_RZJNQvYs6_1(.din(n768),.dout(w_dff_B_RZJNQvYs6_1),.clk(gclk));
	jdff dff_B_5wOZZdvr8_2(.din(n674),.dout(w_dff_B_5wOZZdvr8_2),.clk(gclk));
	jdff dff_B_LRAwW28o0_2(.din(w_dff_B_5wOZZdvr8_2),.dout(w_dff_B_LRAwW28o0_2),.clk(gclk));
	jdff dff_B_nwnijX4W2_2(.din(w_dff_B_LRAwW28o0_2),.dout(w_dff_B_nwnijX4W2_2),.clk(gclk));
	jdff dff_B_kSxzxN4e4_2(.din(w_dff_B_nwnijX4W2_2),.dout(w_dff_B_kSxzxN4e4_2),.clk(gclk));
	jdff dff_B_VrSglJYH0_2(.din(w_dff_B_kSxzxN4e4_2),.dout(w_dff_B_VrSglJYH0_2),.clk(gclk));
	jdff dff_B_B5J6Viwa8_2(.din(w_dff_B_VrSglJYH0_2),.dout(w_dff_B_B5J6Viwa8_2),.clk(gclk));
	jdff dff_B_0iOOLS0p4_2(.din(w_dff_B_B5J6Viwa8_2),.dout(w_dff_B_0iOOLS0p4_2),.clk(gclk));
	jdff dff_B_Ra50P0mj4_2(.din(w_dff_B_0iOOLS0p4_2),.dout(w_dff_B_Ra50P0mj4_2),.clk(gclk));
	jdff dff_B_otY1Qg072_2(.din(w_dff_B_Ra50P0mj4_2),.dout(w_dff_B_otY1Qg072_2),.clk(gclk));
	jdff dff_B_lLJRwPWq6_2(.din(w_dff_B_otY1Qg072_2),.dout(w_dff_B_lLJRwPWq6_2),.clk(gclk));
	jdff dff_B_ix6HIcZB0_2(.din(w_dff_B_lLJRwPWq6_2),.dout(w_dff_B_ix6HIcZB0_2),.clk(gclk));
	jdff dff_B_1cZyvX0q5_2(.din(w_dff_B_ix6HIcZB0_2),.dout(w_dff_B_1cZyvX0q5_2),.clk(gclk));
	jdff dff_B_Y9rg3qgF9_1(.din(n675),.dout(w_dff_B_Y9rg3qgF9_1),.clk(gclk));
	jdff dff_B_RSKJMgTC5_2(.din(n588),.dout(w_dff_B_RSKJMgTC5_2),.clk(gclk));
	jdff dff_B_SnpKHp4H3_2(.din(w_dff_B_RSKJMgTC5_2),.dout(w_dff_B_SnpKHp4H3_2),.clk(gclk));
	jdff dff_B_r1JyNFpg6_2(.din(w_dff_B_SnpKHp4H3_2),.dout(w_dff_B_r1JyNFpg6_2),.clk(gclk));
	jdff dff_B_16yNG7l58_2(.din(w_dff_B_r1JyNFpg6_2),.dout(w_dff_B_16yNG7l58_2),.clk(gclk));
	jdff dff_B_HpmQSZxj5_2(.din(w_dff_B_16yNG7l58_2),.dout(w_dff_B_HpmQSZxj5_2),.clk(gclk));
	jdff dff_B_5FkPQTEG1_2(.din(w_dff_B_HpmQSZxj5_2),.dout(w_dff_B_5FkPQTEG1_2),.clk(gclk));
	jdff dff_B_gsQZ6bPP0_2(.din(w_dff_B_5FkPQTEG1_2),.dout(w_dff_B_gsQZ6bPP0_2),.clk(gclk));
	jdff dff_B_19w1q5RB4_2(.din(w_dff_B_gsQZ6bPP0_2),.dout(w_dff_B_19w1q5RB4_2),.clk(gclk));
	jdff dff_B_fAYXX5oW1_2(.din(w_dff_B_19w1q5RB4_2),.dout(w_dff_B_fAYXX5oW1_2),.clk(gclk));
	jdff dff_B_W8fOQmi79_2(.din(w_dff_B_fAYXX5oW1_2),.dout(w_dff_B_W8fOQmi79_2),.clk(gclk));
	jdff dff_B_bs4LziED4_1(.din(n589),.dout(w_dff_B_bs4LziED4_1),.clk(gclk));
	jdff dff_B_6p1u8bTu7_2(.din(n509),.dout(w_dff_B_6p1u8bTu7_2),.clk(gclk));
	jdff dff_B_2fcZf6734_2(.din(w_dff_B_6p1u8bTu7_2),.dout(w_dff_B_2fcZf6734_2),.clk(gclk));
	jdff dff_B_rXYW2y8B0_2(.din(w_dff_B_2fcZf6734_2),.dout(w_dff_B_rXYW2y8B0_2),.clk(gclk));
	jdff dff_B_GWLpQpMt3_2(.din(w_dff_B_rXYW2y8B0_2),.dout(w_dff_B_GWLpQpMt3_2),.clk(gclk));
	jdff dff_B_ew4zP9lJ7_2(.din(w_dff_B_GWLpQpMt3_2),.dout(w_dff_B_ew4zP9lJ7_2),.clk(gclk));
	jdff dff_B_49XzoXZA7_2(.din(w_dff_B_ew4zP9lJ7_2),.dout(w_dff_B_49XzoXZA7_2),.clk(gclk));
	jdff dff_B_GI6vog5R5_2(.din(w_dff_B_49XzoXZA7_2),.dout(w_dff_B_GI6vog5R5_2),.clk(gclk));
	jdff dff_B_pxhg50Db2_2(.din(w_dff_B_GI6vog5R5_2),.dout(w_dff_B_pxhg50Db2_2),.clk(gclk));
	jdff dff_B_JGGGdc0n8_1(.din(n510),.dout(w_dff_B_JGGGdc0n8_1),.clk(gclk));
	jdff dff_B_zQNwH8Bu3_2(.din(n437),.dout(w_dff_B_zQNwH8Bu3_2),.clk(gclk));
	jdff dff_B_3S6wzICb9_2(.din(w_dff_B_zQNwH8Bu3_2),.dout(w_dff_B_3S6wzICb9_2),.clk(gclk));
	jdff dff_B_3Iv169k68_2(.din(w_dff_B_3S6wzICb9_2),.dout(w_dff_B_3Iv169k68_2),.clk(gclk));
	jdff dff_B_7y75TMyj1_2(.din(w_dff_B_3Iv169k68_2),.dout(w_dff_B_7y75TMyj1_2),.clk(gclk));
	jdff dff_B_gSJHo93y5_2(.din(w_dff_B_7y75TMyj1_2),.dout(w_dff_B_gSJHo93y5_2),.clk(gclk));
	jdff dff_B_q6FLbAux0_2(.din(w_dff_B_gSJHo93y5_2),.dout(w_dff_B_q6FLbAux0_2),.clk(gclk));
	jdff dff_B_GAwbNi6N6_2(.din(n453),.dout(w_dff_B_GAwbNi6N6_2),.clk(gclk));
	jdff dff_B_EahjSriI7_1(.din(n438),.dout(w_dff_B_EahjSriI7_1),.clk(gclk));
	jdff dff_B_sUcNy1gV9_1(.din(w_dff_B_EahjSriI7_1),.dout(w_dff_B_sUcNy1gV9_1),.clk(gclk));
	jdff dff_B_UFFyI5mw4_1(.din(w_dff_B_sUcNy1gV9_1),.dout(w_dff_B_UFFyI5mw4_1),.clk(gclk));
	jdff dff_B_hbzpAAfY3_1(.din(w_dff_B_UFFyI5mw4_1),.dout(w_dff_B_hbzpAAfY3_1),.clk(gclk));
	jdff dff_B_5JXtGLp18_0(.din(n381),.dout(w_dff_B_5JXtGLp18_0),.clk(gclk));
	jdff dff_A_6lXKfSQ66_0(.dout(w_n380_0[0]),.din(w_dff_A_6lXKfSQ66_0),.clk(gclk));
	jdff dff_A_vJmeg3EW2_0(.dout(w_dff_A_6lXKfSQ66_0),.din(w_dff_A_vJmeg3EW2_0),.clk(gclk));
	jdff dff_B_8PB5xVkM2_1(.din(n374),.dout(w_dff_B_8PB5xVkM2_1),.clk(gclk));
	jdff dff_B_JAaSJxCS7_1(.din(w_dff_B_8PB5xVkM2_1),.dout(w_dff_B_JAaSJxCS7_1),.clk(gclk));
	jdff dff_A_0wMb0ngO3_0(.dout(w_n314_0[0]),.din(w_dff_A_0wMb0ngO3_0),.clk(gclk));
	jdff dff_A_TKGC6uMf4_1(.dout(w_n314_0[1]),.din(w_dff_A_TKGC6uMf4_1),.clk(gclk));
	jdff dff_A_mzOkYWKK3_1(.dout(w_dff_A_TKGC6uMf4_1),.din(w_dff_A_mzOkYWKK3_1),.clk(gclk));
	jdff dff_A_vMC9VBYo7_1(.dout(w_n372_0[1]),.din(w_dff_A_vMC9VBYo7_1),.clk(gclk));
	jdff dff_A_RpSN5RcD5_1(.dout(w_dff_A_vMC9VBYo7_1),.din(w_dff_A_RpSN5RcD5_1),.clk(gclk));
	jdff dff_A_2HGbCkl93_1(.dout(w_dff_A_RpSN5RcD5_1),.din(w_dff_A_2HGbCkl93_1),.clk(gclk));
	jdff dff_A_dfd1enHt4_1(.dout(w_dff_A_2HGbCkl93_1),.din(w_dff_A_dfd1enHt4_1),.clk(gclk));
	jdff dff_B_WzbyGmmA2_2(.din(n1627),.dout(w_dff_B_WzbyGmmA2_2),.clk(gclk));
	jdff dff_B_Q6bCvniE8_2(.din(w_dff_B_WzbyGmmA2_2),.dout(w_dff_B_Q6bCvniE8_2),.clk(gclk));
	jdff dff_B_OXtOuo0n0_1(.din(n1625),.dout(w_dff_B_OXtOuo0n0_1),.clk(gclk));
	jdff dff_B_VivaAZGf5_2(.din(n1566),.dout(w_dff_B_VivaAZGf5_2),.clk(gclk));
	jdff dff_B_dxhVN85L7_2(.din(w_dff_B_VivaAZGf5_2),.dout(w_dff_B_dxhVN85L7_2),.clk(gclk));
	jdff dff_B_L5JB73sA2_2(.din(w_dff_B_dxhVN85L7_2),.dout(w_dff_B_L5JB73sA2_2),.clk(gclk));
	jdff dff_B_BaXxZ3uv4_2(.din(w_dff_B_L5JB73sA2_2),.dout(w_dff_B_BaXxZ3uv4_2),.clk(gclk));
	jdff dff_B_blhrujv86_2(.din(w_dff_B_BaXxZ3uv4_2),.dout(w_dff_B_blhrujv86_2),.clk(gclk));
	jdff dff_B_523Asw6t5_2(.din(w_dff_B_blhrujv86_2),.dout(w_dff_B_523Asw6t5_2),.clk(gclk));
	jdff dff_B_XW9bV9d58_2(.din(w_dff_B_523Asw6t5_2),.dout(w_dff_B_XW9bV9d58_2),.clk(gclk));
	jdff dff_B_hwGE6lXr4_2(.din(w_dff_B_XW9bV9d58_2),.dout(w_dff_B_hwGE6lXr4_2),.clk(gclk));
	jdff dff_B_m6GYAWr86_2(.din(w_dff_B_hwGE6lXr4_2),.dout(w_dff_B_m6GYAWr86_2),.clk(gclk));
	jdff dff_B_M8HdBnQg3_2(.din(w_dff_B_m6GYAWr86_2),.dout(w_dff_B_M8HdBnQg3_2),.clk(gclk));
	jdff dff_B_bNLhdBen5_2(.din(w_dff_B_M8HdBnQg3_2),.dout(w_dff_B_bNLhdBen5_2),.clk(gclk));
	jdff dff_B_jl6Qpt129_2(.din(w_dff_B_bNLhdBen5_2),.dout(w_dff_B_jl6Qpt129_2),.clk(gclk));
	jdff dff_B_fy9fkraS8_2(.din(w_dff_B_jl6Qpt129_2),.dout(w_dff_B_fy9fkraS8_2),.clk(gclk));
	jdff dff_B_vROizhuz3_2(.din(w_dff_B_fy9fkraS8_2),.dout(w_dff_B_vROizhuz3_2),.clk(gclk));
	jdff dff_B_FAcelAv48_2(.din(w_dff_B_vROizhuz3_2),.dout(w_dff_B_FAcelAv48_2),.clk(gclk));
	jdff dff_B_Te6PE2su3_2(.din(w_dff_B_FAcelAv48_2),.dout(w_dff_B_Te6PE2su3_2),.clk(gclk));
	jdff dff_B_4ncCPWBp1_2(.din(w_dff_B_Te6PE2su3_2),.dout(w_dff_B_4ncCPWBp1_2),.clk(gclk));
	jdff dff_B_dtLNku6w6_2(.din(w_dff_B_4ncCPWBp1_2),.dout(w_dff_B_dtLNku6w6_2),.clk(gclk));
	jdff dff_B_IAVikLSt5_2(.din(w_dff_B_dtLNku6w6_2),.dout(w_dff_B_IAVikLSt5_2),.clk(gclk));
	jdff dff_B_825JNzyU2_2(.din(w_dff_B_IAVikLSt5_2),.dout(w_dff_B_825JNzyU2_2),.clk(gclk));
	jdff dff_B_D0ocor7n0_2(.din(w_dff_B_825JNzyU2_2),.dout(w_dff_B_D0ocor7n0_2),.clk(gclk));
	jdff dff_B_inUuGzy63_2(.din(w_dff_B_D0ocor7n0_2),.dout(w_dff_B_inUuGzy63_2),.clk(gclk));
	jdff dff_B_Kd5ISFHJ0_2(.din(w_dff_B_inUuGzy63_2),.dout(w_dff_B_Kd5ISFHJ0_2),.clk(gclk));
	jdff dff_B_0Ct8Owza1_2(.din(w_dff_B_Kd5ISFHJ0_2),.dout(w_dff_B_0Ct8Owza1_2),.clk(gclk));
	jdff dff_B_J01f5gZB6_2(.din(w_dff_B_0Ct8Owza1_2),.dout(w_dff_B_J01f5gZB6_2),.clk(gclk));
	jdff dff_B_VOLourEz6_2(.din(w_dff_B_J01f5gZB6_2),.dout(w_dff_B_VOLourEz6_2),.clk(gclk));
	jdff dff_B_W3bsBN664_2(.din(w_dff_B_VOLourEz6_2),.dout(w_dff_B_W3bsBN664_2),.clk(gclk));
	jdff dff_B_dv8YtCXg3_2(.din(w_dff_B_W3bsBN664_2),.dout(w_dff_B_dv8YtCXg3_2),.clk(gclk));
	jdff dff_B_Qm3fjjHW8_2(.din(w_dff_B_dv8YtCXg3_2),.dout(w_dff_B_Qm3fjjHW8_2),.clk(gclk));
	jdff dff_B_1wvE6DfL2_2(.din(w_dff_B_Qm3fjjHW8_2),.dout(w_dff_B_1wvE6DfL2_2),.clk(gclk));
	jdff dff_B_k9m4mWxG5_2(.din(w_dff_B_1wvE6DfL2_2),.dout(w_dff_B_k9m4mWxG5_2),.clk(gclk));
	jdff dff_B_kEgN8ZEG5_2(.din(w_dff_B_k9m4mWxG5_2),.dout(w_dff_B_kEgN8ZEG5_2),.clk(gclk));
	jdff dff_B_bQ8ocjeg3_2(.din(w_dff_B_kEgN8ZEG5_2),.dout(w_dff_B_bQ8ocjeg3_2),.clk(gclk));
	jdff dff_B_jdZKA79M3_2(.din(w_dff_B_bQ8ocjeg3_2),.dout(w_dff_B_jdZKA79M3_2),.clk(gclk));
	jdff dff_B_KtU7i8xS3_2(.din(w_dff_B_jdZKA79M3_2),.dout(w_dff_B_KtU7i8xS3_2),.clk(gclk));
	jdff dff_B_ghOwIdW76_2(.din(w_dff_B_KtU7i8xS3_2),.dout(w_dff_B_ghOwIdW76_2),.clk(gclk));
	jdff dff_B_3zRtCl133_2(.din(w_dff_B_ghOwIdW76_2),.dout(w_dff_B_3zRtCl133_2),.clk(gclk));
	jdff dff_B_UW8CfZ038_2(.din(w_dff_B_3zRtCl133_2),.dout(w_dff_B_UW8CfZ038_2),.clk(gclk));
	jdff dff_B_OF2s7hnL4_2(.din(w_dff_B_UW8CfZ038_2),.dout(w_dff_B_OF2s7hnL4_2),.clk(gclk));
	jdff dff_B_PPlTCACc9_1(.din(n1623),.dout(w_dff_B_PPlTCACc9_1),.clk(gclk));
	jdff dff_A_MJhgLnrt6_1(.dout(w_n1569_0[1]),.din(w_dff_A_MJhgLnrt6_1),.clk(gclk));
	jdff dff_B_9d5lIpiV0_1(.din(n1567),.dout(w_dff_B_9d5lIpiV0_1),.clk(gclk));
	jdff dff_B_ATDfNSBi9_2(.din(n1502),.dout(w_dff_B_ATDfNSBi9_2),.clk(gclk));
	jdff dff_B_LcMhr7te4_2(.din(w_dff_B_ATDfNSBi9_2),.dout(w_dff_B_LcMhr7te4_2),.clk(gclk));
	jdff dff_B_fwAdRSxc1_2(.din(w_dff_B_LcMhr7te4_2),.dout(w_dff_B_fwAdRSxc1_2),.clk(gclk));
	jdff dff_B_FiJ6I9Kw9_2(.din(w_dff_B_fwAdRSxc1_2),.dout(w_dff_B_FiJ6I9Kw9_2),.clk(gclk));
	jdff dff_B_h26dof0y6_2(.din(w_dff_B_FiJ6I9Kw9_2),.dout(w_dff_B_h26dof0y6_2),.clk(gclk));
	jdff dff_B_M13B73Rl5_2(.din(w_dff_B_h26dof0y6_2),.dout(w_dff_B_M13B73Rl5_2),.clk(gclk));
	jdff dff_B_7klzmQe00_2(.din(w_dff_B_M13B73Rl5_2),.dout(w_dff_B_7klzmQe00_2),.clk(gclk));
	jdff dff_B_0amQgcDR7_2(.din(w_dff_B_7klzmQe00_2),.dout(w_dff_B_0amQgcDR7_2),.clk(gclk));
	jdff dff_B_0GQtr2Pz5_2(.din(w_dff_B_0amQgcDR7_2),.dout(w_dff_B_0GQtr2Pz5_2),.clk(gclk));
	jdff dff_B_Fp40F1wp5_2(.din(w_dff_B_0GQtr2Pz5_2),.dout(w_dff_B_Fp40F1wp5_2),.clk(gclk));
	jdff dff_B_CQzWXpjG9_2(.din(w_dff_B_Fp40F1wp5_2),.dout(w_dff_B_CQzWXpjG9_2),.clk(gclk));
	jdff dff_B_WzPFBeTY3_2(.din(w_dff_B_CQzWXpjG9_2),.dout(w_dff_B_WzPFBeTY3_2),.clk(gclk));
	jdff dff_B_nhQxcUvz6_2(.din(w_dff_B_WzPFBeTY3_2),.dout(w_dff_B_nhQxcUvz6_2),.clk(gclk));
	jdff dff_B_buPShKzW5_2(.din(w_dff_B_nhQxcUvz6_2),.dout(w_dff_B_buPShKzW5_2),.clk(gclk));
	jdff dff_B_A6a9nHVX3_2(.din(w_dff_B_buPShKzW5_2),.dout(w_dff_B_A6a9nHVX3_2),.clk(gclk));
	jdff dff_B_UZS45at09_2(.din(w_dff_B_A6a9nHVX3_2),.dout(w_dff_B_UZS45at09_2),.clk(gclk));
	jdff dff_B_tf2hMgAb3_2(.din(w_dff_B_UZS45at09_2),.dout(w_dff_B_tf2hMgAb3_2),.clk(gclk));
	jdff dff_B_uVVKptxL7_2(.din(w_dff_B_tf2hMgAb3_2),.dout(w_dff_B_uVVKptxL7_2),.clk(gclk));
	jdff dff_B_wYPlqcNd4_2(.din(w_dff_B_uVVKptxL7_2),.dout(w_dff_B_wYPlqcNd4_2),.clk(gclk));
	jdff dff_B_BjnLBjEC6_2(.din(w_dff_B_wYPlqcNd4_2),.dout(w_dff_B_BjnLBjEC6_2),.clk(gclk));
	jdff dff_B_su1LrFrP6_2(.din(w_dff_B_BjnLBjEC6_2),.dout(w_dff_B_su1LrFrP6_2),.clk(gclk));
	jdff dff_B_o54ktGE82_2(.din(w_dff_B_su1LrFrP6_2),.dout(w_dff_B_o54ktGE82_2),.clk(gclk));
	jdff dff_B_X5jePmM40_2(.din(w_dff_B_o54ktGE82_2),.dout(w_dff_B_X5jePmM40_2),.clk(gclk));
	jdff dff_B_12YaLQ0O4_2(.din(w_dff_B_X5jePmM40_2),.dout(w_dff_B_12YaLQ0O4_2),.clk(gclk));
	jdff dff_B_M8pe2DeQ2_2(.din(w_dff_B_12YaLQ0O4_2),.dout(w_dff_B_M8pe2DeQ2_2),.clk(gclk));
	jdff dff_B_67ubSu1H8_2(.din(w_dff_B_M8pe2DeQ2_2),.dout(w_dff_B_67ubSu1H8_2),.clk(gclk));
	jdff dff_B_RXyLOIHN0_2(.din(w_dff_B_67ubSu1H8_2),.dout(w_dff_B_RXyLOIHN0_2),.clk(gclk));
	jdff dff_B_UKqOHD4M8_2(.din(w_dff_B_RXyLOIHN0_2),.dout(w_dff_B_UKqOHD4M8_2),.clk(gclk));
	jdff dff_B_lOJF4shG3_2(.din(w_dff_B_UKqOHD4M8_2),.dout(w_dff_B_lOJF4shG3_2),.clk(gclk));
	jdff dff_B_61IsavOV3_2(.din(w_dff_B_lOJF4shG3_2),.dout(w_dff_B_61IsavOV3_2),.clk(gclk));
	jdff dff_B_orlTxHSF1_2(.din(w_dff_B_61IsavOV3_2),.dout(w_dff_B_orlTxHSF1_2),.clk(gclk));
	jdff dff_B_Aos02Svp1_2(.din(w_dff_B_orlTxHSF1_2),.dout(w_dff_B_Aos02Svp1_2),.clk(gclk));
	jdff dff_B_jWRVVLyV4_2(.din(w_dff_B_Aos02Svp1_2),.dout(w_dff_B_jWRVVLyV4_2),.clk(gclk));
	jdff dff_B_cAOgaJXH0_2(.din(w_dff_B_jWRVVLyV4_2),.dout(w_dff_B_cAOgaJXH0_2),.clk(gclk));
	jdff dff_B_M9r7IJP04_2(.din(n1505),.dout(w_dff_B_M9r7IJP04_2),.clk(gclk));
	jdff dff_B_Mfh0kkv02_1(.din(n1503),.dout(w_dff_B_Mfh0kkv02_1),.clk(gclk));
	jdff dff_B_23vx0GH01_2(.din(n1431),.dout(w_dff_B_23vx0GH01_2),.clk(gclk));
	jdff dff_B_TNlgw6GN2_2(.din(w_dff_B_23vx0GH01_2),.dout(w_dff_B_TNlgw6GN2_2),.clk(gclk));
	jdff dff_B_WZCe2WkR3_2(.din(w_dff_B_TNlgw6GN2_2),.dout(w_dff_B_WZCe2WkR3_2),.clk(gclk));
	jdff dff_B_wkb3VJOY5_2(.din(w_dff_B_WZCe2WkR3_2),.dout(w_dff_B_wkb3VJOY5_2),.clk(gclk));
	jdff dff_B_TKPoNh7x1_2(.din(w_dff_B_wkb3VJOY5_2),.dout(w_dff_B_TKPoNh7x1_2),.clk(gclk));
	jdff dff_B_Dpjta17I5_2(.din(w_dff_B_TKPoNh7x1_2),.dout(w_dff_B_Dpjta17I5_2),.clk(gclk));
	jdff dff_B_EooeiXEp8_2(.din(w_dff_B_Dpjta17I5_2),.dout(w_dff_B_EooeiXEp8_2),.clk(gclk));
	jdff dff_B_yA5dxsfP7_2(.din(w_dff_B_EooeiXEp8_2),.dout(w_dff_B_yA5dxsfP7_2),.clk(gclk));
	jdff dff_B_BGLINkCJ1_2(.din(w_dff_B_yA5dxsfP7_2),.dout(w_dff_B_BGLINkCJ1_2),.clk(gclk));
	jdff dff_B_Itf4hP8e8_2(.din(w_dff_B_BGLINkCJ1_2),.dout(w_dff_B_Itf4hP8e8_2),.clk(gclk));
	jdff dff_B_seAxaf2Q7_2(.din(w_dff_B_Itf4hP8e8_2),.dout(w_dff_B_seAxaf2Q7_2),.clk(gclk));
	jdff dff_B_yuPoDNyZ2_2(.din(w_dff_B_seAxaf2Q7_2),.dout(w_dff_B_yuPoDNyZ2_2),.clk(gclk));
	jdff dff_B_HgiqbXGI1_2(.din(w_dff_B_yuPoDNyZ2_2),.dout(w_dff_B_HgiqbXGI1_2),.clk(gclk));
	jdff dff_B_2zaxelzr8_2(.din(w_dff_B_HgiqbXGI1_2),.dout(w_dff_B_2zaxelzr8_2),.clk(gclk));
	jdff dff_B_kR7qHsBI9_2(.din(w_dff_B_2zaxelzr8_2),.dout(w_dff_B_kR7qHsBI9_2),.clk(gclk));
	jdff dff_B_vt4oSdHW1_2(.din(w_dff_B_kR7qHsBI9_2),.dout(w_dff_B_vt4oSdHW1_2),.clk(gclk));
	jdff dff_B_jvpwUup52_2(.din(w_dff_B_vt4oSdHW1_2),.dout(w_dff_B_jvpwUup52_2),.clk(gclk));
	jdff dff_B_F0QEjJoF4_2(.din(w_dff_B_jvpwUup52_2),.dout(w_dff_B_F0QEjJoF4_2),.clk(gclk));
	jdff dff_B_qGgJHG8F2_2(.din(w_dff_B_F0QEjJoF4_2),.dout(w_dff_B_qGgJHG8F2_2),.clk(gclk));
	jdff dff_B_xnKraAcX6_2(.din(w_dff_B_qGgJHG8F2_2),.dout(w_dff_B_xnKraAcX6_2),.clk(gclk));
	jdff dff_B_fGX8GYOV2_2(.din(w_dff_B_xnKraAcX6_2),.dout(w_dff_B_fGX8GYOV2_2),.clk(gclk));
	jdff dff_B_dH9KQSq26_2(.din(w_dff_B_fGX8GYOV2_2),.dout(w_dff_B_dH9KQSq26_2),.clk(gclk));
	jdff dff_B_RMtLGD6b1_2(.din(w_dff_B_dH9KQSq26_2),.dout(w_dff_B_RMtLGD6b1_2),.clk(gclk));
	jdff dff_B_9LfUq9Ol8_2(.din(w_dff_B_RMtLGD6b1_2),.dout(w_dff_B_9LfUq9Ol8_2),.clk(gclk));
	jdff dff_B_7sG1xqag1_2(.din(w_dff_B_9LfUq9Ol8_2),.dout(w_dff_B_7sG1xqag1_2),.clk(gclk));
	jdff dff_B_78oPaTnY2_2(.din(w_dff_B_7sG1xqag1_2),.dout(w_dff_B_78oPaTnY2_2),.clk(gclk));
	jdff dff_B_7DGOZhca9_2(.din(w_dff_B_78oPaTnY2_2),.dout(w_dff_B_7DGOZhca9_2),.clk(gclk));
	jdff dff_B_TDQazCe19_2(.din(w_dff_B_7DGOZhca9_2),.dout(w_dff_B_TDQazCe19_2),.clk(gclk));
	jdff dff_B_ERWAJdHi6_2(.din(w_dff_B_TDQazCe19_2),.dout(w_dff_B_ERWAJdHi6_2),.clk(gclk));
	jdff dff_B_kC9lnoRe0_2(.din(w_dff_B_ERWAJdHi6_2),.dout(w_dff_B_kC9lnoRe0_2),.clk(gclk));
	jdff dff_B_ZIjzh16U2_2(.din(w_dff_B_kC9lnoRe0_2),.dout(w_dff_B_ZIjzh16U2_2),.clk(gclk));
	jdff dff_B_kLPA1nxm0_2(.din(n1434),.dout(w_dff_B_kLPA1nxm0_2),.clk(gclk));
	jdff dff_B_t9QCbYnh7_1(.din(n1432),.dout(w_dff_B_t9QCbYnh7_1),.clk(gclk));
	jdff dff_B_rFKOjRJD1_2(.din(n1353),.dout(w_dff_B_rFKOjRJD1_2),.clk(gclk));
	jdff dff_B_Shkzqvwb0_2(.din(w_dff_B_rFKOjRJD1_2),.dout(w_dff_B_Shkzqvwb0_2),.clk(gclk));
	jdff dff_B_7LkwtkoP0_2(.din(w_dff_B_Shkzqvwb0_2),.dout(w_dff_B_7LkwtkoP0_2),.clk(gclk));
	jdff dff_B_kA4fFiSm0_2(.din(w_dff_B_7LkwtkoP0_2),.dout(w_dff_B_kA4fFiSm0_2),.clk(gclk));
	jdff dff_B_CWWJfgdC8_2(.din(w_dff_B_kA4fFiSm0_2),.dout(w_dff_B_CWWJfgdC8_2),.clk(gclk));
	jdff dff_B_JvBhLCxV4_2(.din(w_dff_B_CWWJfgdC8_2),.dout(w_dff_B_JvBhLCxV4_2),.clk(gclk));
	jdff dff_B_MCM2zMCV8_2(.din(w_dff_B_JvBhLCxV4_2),.dout(w_dff_B_MCM2zMCV8_2),.clk(gclk));
	jdff dff_B_OkG67PvN7_2(.din(w_dff_B_MCM2zMCV8_2),.dout(w_dff_B_OkG67PvN7_2),.clk(gclk));
	jdff dff_B_eKw7XMBP8_2(.din(w_dff_B_OkG67PvN7_2),.dout(w_dff_B_eKw7XMBP8_2),.clk(gclk));
	jdff dff_B_0UktzvSF0_2(.din(w_dff_B_eKw7XMBP8_2),.dout(w_dff_B_0UktzvSF0_2),.clk(gclk));
	jdff dff_B_E0nCYUDn0_2(.din(w_dff_B_0UktzvSF0_2),.dout(w_dff_B_E0nCYUDn0_2),.clk(gclk));
	jdff dff_B_yZNCcRCE1_2(.din(w_dff_B_E0nCYUDn0_2),.dout(w_dff_B_yZNCcRCE1_2),.clk(gclk));
	jdff dff_B_0x3WEO4a7_2(.din(w_dff_B_yZNCcRCE1_2),.dout(w_dff_B_0x3WEO4a7_2),.clk(gclk));
	jdff dff_B_HtG1hsF88_2(.din(w_dff_B_0x3WEO4a7_2),.dout(w_dff_B_HtG1hsF88_2),.clk(gclk));
	jdff dff_B_kHof0M1V0_2(.din(w_dff_B_HtG1hsF88_2),.dout(w_dff_B_kHof0M1V0_2),.clk(gclk));
	jdff dff_B_dTu2bsFh9_2(.din(w_dff_B_kHof0M1V0_2),.dout(w_dff_B_dTu2bsFh9_2),.clk(gclk));
	jdff dff_B_FBdQq1Ql5_2(.din(w_dff_B_dTu2bsFh9_2),.dout(w_dff_B_FBdQq1Ql5_2),.clk(gclk));
	jdff dff_B_UotZ01n04_2(.din(w_dff_B_FBdQq1Ql5_2),.dout(w_dff_B_UotZ01n04_2),.clk(gclk));
	jdff dff_B_kJBVrZbv9_2(.din(w_dff_B_UotZ01n04_2),.dout(w_dff_B_kJBVrZbv9_2),.clk(gclk));
	jdff dff_B_fiE1NPPs0_2(.din(w_dff_B_kJBVrZbv9_2),.dout(w_dff_B_fiE1NPPs0_2),.clk(gclk));
	jdff dff_B_3BSHEZxH4_2(.din(w_dff_B_fiE1NPPs0_2),.dout(w_dff_B_3BSHEZxH4_2),.clk(gclk));
	jdff dff_B_J4bdGMyz8_2(.din(w_dff_B_3BSHEZxH4_2),.dout(w_dff_B_J4bdGMyz8_2),.clk(gclk));
	jdff dff_B_iqb96eDF6_2(.din(w_dff_B_J4bdGMyz8_2),.dout(w_dff_B_iqb96eDF6_2),.clk(gclk));
	jdff dff_B_nmskeV6s8_2(.din(w_dff_B_iqb96eDF6_2),.dout(w_dff_B_nmskeV6s8_2),.clk(gclk));
	jdff dff_B_ovsV0Zdr1_2(.din(w_dff_B_nmskeV6s8_2),.dout(w_dff_B_ovsV0Zdr1_2),.clk(gclk));
	jdff dff_B_4gEHlifp4_2(.din(w_dff_B_ovsV0Zdr1_2),.dout(w_dff_B_4gEHlifp4_2),.clk(gclk));
	jdff dff_B_2WrrBva48_2(.din(w_dff_B_4gEHlifp4_2),.dout(w_dff_B_2WrrBva48_2),.clk(gclk));
	jdff dff_B_pZFYSmTh4_2(.din(w_dff_B_2WrrBva48_2),.dout(w_dff_B_pZFYSmTh4_2),.clk(gclk));
	jdff dff_B_hux4zV000_2(.din(n1356),.dout(w_dff_B_hux4zV000_2),.clk(gclk));
	jdff dff_B_gQxEYNeQ5_1(.din(n1354),.dout(w_dff_B_gQxEYNeQ5_1),.clk(gclk));
	jdff dff_B_DlDxXjjK6_2(.din(n1268),.dout(w_dff_B_DlDxXjjK6_2),.clk(gclk));
	jdff dff_B_z8eyT1QK9_2(.din(w_dff_B_DlDxXjjK6_2),.dout(w_dff_B_z8eyT1QK9_2),.clk(gclk));
	jdff dff_B_6tu7Q9JE6_2(.din(w_dff_B_z8eyT1QK9_2),.dout(w_dff_B_6tu7Q9JE6_2),.clk(gclk));
	jdff dff_B_6CGTOujS7_2(.din(w_dff_B_6tu7Q9JE6_2),.dout(w_dff_B_6CGTOujS7_2),.clk(gclk));
	jdff dff_B_tf71UJPL0_2(.din(w_dff_B_6CGTOujS7_2),.dout(w_dff_B_tf71UJPL0_2),.clk(gclk));
	jdff dff_B_vFBEuL2u5_2(.din(w_dff_B_tf71UJPL0_2),.dout(w_dff_B_vFBEuL2u5_2),.clk(gclk));
	jdff dff_B_LYshGEXw5_2(.din(w_dff_B_vFBEuL2u5_2),.dout(w_dff_B_LYshGEXw5_2),.clk(gclk));
	jdff dff_B_m8QAwYiR9_2(.din(w_dff_B_LYshGEXw5_2),.dout(w_dff_B_m8QAwYiR9_2),.clk(gclk));
	jdff dff_B_0u1XMU7m9_2(.din(w_dff_B_m8QAwYiR9_2),.dout(w_dff_B_0u1XMU7m9_2),.clk(gclk));
	jdff dff_B_5OWcZrHL8_2(.din(w_dff_B_0u1XMU7m9_2),.dout(w_dff_B_5OWcZrHL8_2),.clk(gclk));
	jdff dff_B_JuhOzneL0_2(.din(w_dff_B_5OWcZrHL8_2),.dout(w_dff_B_JuhOzneL0_2),.clk(gclk));
	jdff dff_B_LcNVsmoM5_2(.din(w_dff_B_JuhOzneL0_2),.dout(w_dff_B_LcNVsmoM5_2),.clk(gclk));
	jdff dff_B_THtRRqyG5_2(.din(w_dff_B_LcNVsmoM5_2),.dout(w_dff_B_THtRRqyG5_2),.clk(gclk));
	jdff dff_B_l3cwipV46_2(.din(w_dff_B_THtRRqyG5_2),.dout(w_dff_B_l3cwipV46_2),.clk(gclk));
	jdff dff_B_UDJerUTc1_2(.din(w_dff_B_l3cwipV46_2),.dout(w_dff_B_UDJerUTc1_2),.clk(gclk));
	jdff dff_B_9SoRBjwU6_2(.din(w_dff_B_UDJerUTc1_2),.dout(w_dff_B_9SoRBjwU6_2),.clk(gclk));
	jdff dff_B_fBJv6lFq8_2(.din(w_dff_B_9SoRBjwU6_2),.dout(w_dff_B_fBJv6lFq8_2),.clk(gclk));
	jdff dff_B_edIW2JsD6_2(.din(w_dff_B_fBJv6lFq8_2),.dout(w_dff_B_edIW2JsD6_2),.clk(gclk));
	jdff dff_B_Oj5RJE7y5_2(.din(w_dff_B_edIW2JsD6_2),.dout(w_dff_B_Oj5RJE7y5_2),.clk(gclk));
	jdff dff_B_cvpuUafq9_2(.din(w_dff_B_Oj5RJE7y5_2),.dout(w_dff_B_cvpuUafq9_2),.clk(gclk));
	jdff dff_B_bfJbFLVg9_2(.din(w_dff_B_cvpuUafq9_2),.dout(w_dff_B_bfJbFLVg9_2),.clk(gclk));
	jdff dff_B_cV1fiaF85_2(.din(w_dff_B_bfJbFLVg9_2),.dout(w_dff_B_cV1fiaF85_2),.clk(gclk));
	jdff dff_B_HyFwnOSo1_2(.din(w_dff_B_cV1fiaF85_2),.dout(w_dff_B_HyFwnOSo1_2),.clk(gclk));
	jdff dff_B_fg2E7zCH3_2(.din(w_dff_B_HyFwnOSo1_2),.dout(w_dff_B_fg2E7zCH3_2),.clk(gclk));
	jdff dff_B_8mTW0Vt24_2(.din(w_dff_B_fg2E7zCH3_2),.dout(w_dff_B_8mTW0Vt24_2),.clk(gclk));
	jdff dff_B_OrMlmBB98_2(.din(n1271),.dout(w_dff_B_OrMlmBB98_2),.clk(gclk));
	jdff dff_B_nhgki9g39_1(.din(n1269),.dout(w_dff_B_nhgki9g39_1),.clk(gclk));
	jdff dff_B_xIgz8OAf0_2(.din(n1178),.dout(w_dff_B_xIgz8OAf0_2),.clk(gclk));
	jdff dff_B_kCjKU8d75_2(.din(w_dff_B_xIgz8OAf0_2),.dout(w_dff_B_kCjKU8d75_2),.clk(gclk));
	jdff dff_B_CJrmh1Ng1_2(.din(w_dff_B_kCjKU8d75_2),.dout(w_dff_B_CJrmh1Ng1_2),.clk(gclk));
	jdff dff_B_6zgyirgm6_2(.din(w_dff_B_CJrmh1Ng1_2),.dout(w_dff_B_6zgyirgm6_2),.clk(gclk));
	jdff dff_B_nWS3J3vD4_2(.din(w_dff_B_6zgyirgm6_2),.dout(w_dff_B_nWS3J3vD4_2),.clk(gclk));
	jdff dff_B_D3kcCUWA4_2(.din(w_dff_B_nWS3J3vD4_2),.dout(w_dff_B_D3kcCUWA4_2),.clk(gclk));
	jdff dff_B_XVspSW4K0_2(.din(w_dff_B_D3kcCUWA4_2),.dout(w_dff_B_XVspSW4K0_2),.clk(gclk));
	jdff dff_B_vAV6LjBg5_2(.din(w_dff_B_XVspSW4K0_2),.dout(w_dff_B_vAV6LjBg5_2),.clk(gclk));
	jdff dff_B_tDDOjzAo6_2(.din(w_dff_B_vAV6LjBg5_2),.dout(w_dff_B_tDDOjzAo6_2),.clk(gclk));
	jdff dff_B_YpgkdWoU9_2(.din(w_dff_B_tDDOjzAo6_2),.dout(w_dff_B_YpgkdWoU9_2),.clk(gclk));
	jdff dff_B_pg2c2Vva2_2(.din(w_dff_B_YpgkdWoU9_2),.dout(w_dff_B_pg2c2Vva2_2),.clk(gclk));
	jdff dff_B_P58eNly96_2(.din(w_dff_B_pg2c2Vva2_2),.dout(w_dff_B_P58eNly96_2),.clk(gclk));
	jdff dff_B_wx3ONJIR5_2(.din(w_dff_B_P58eNly96_2),.dout(w_dff_B_wx3ONJIR5_2),.clk(gclk));
	jdff dff_B_KtJuHBNA3_2(.din(w_dff_B_wx3ONJIR5_2),.dout(w_dff_B_KtJuHBNA3_2),.clk(gclk));
	jdff dff_B_Cn3U6h028_2(.din(w_dff_B_KtJuHBNA3_2),.dout(w_dff_B_Cn3U6h028_2),.clk(gclk));
	jdff dff_B_tQZnQ0fb9_2(.din(w_dff_B_Cn3U6h028_2),.dout(w_dff_B_tQZnQ0fb9_2),.clk(gclk));
	jdff dff_B_RzYDs5yO4_2(.din(w_dff_B_tQZnQ0fb9_2),.dout(w_dff_B_RzYDs5yO4_2),.clk(gclk));
	jdff dff_B_hsNE3Nwh0_2(.din(w_dff_B_RzYDs5yO4_2),.dout(w_dff_B_hsNE3Nwh0_2),.clk(gclk));
	jdff dff_B_J84qplZY5_2(.din(w_dff_B_hsNE3Nwh0_2),.dout(w_dff_B_J84qplZY5_2),.clk(gclk));
	jdff dff_B_R3Cmfkw32_2(.din(w_dff_B_J84qplZY5_2),.dout(w_dff_B_R3Cmfkw32_2),.clk(gclk));
	jdff dff_B_YiiwBcoV5_2(.din(w_dff_B_R3Cmfkw32_2),.dout(w_dff_B_YiiwBcoV5_2),.clk(gclk));
	jdff dff_B_qM3TMyS62_2(.din(w_dff_B_YiiwBcoV5_2),.dout(w_dff_B_qM3TMyS62_2),.clk(gclk));
	jdff dff_B_eLwyZtca5_2(.din(n1181),.dout(w_dff_B_eLwyZtca5_2),.clk(gclk));
	jdff dff_B_J41R32b15_1(.din(n1179),.dout(w_dff_B_J41R32b15_1),.clk(gclk));
	jdff dff_B_SvmA60150_2(.din(n1074),.dout(w_dff_B_SvmA60150_2),.clk(gclk));
	jdff dff_B_HNdLjouM6_2(.din(w_dff_B_SvmA60150_2),.dout(w_dff_B_HNdLjouM6_2),.clk(gclk));
	jdff dff_B_2oalaXv76_2(.din(w_dff_B_HNdLjouM6_2),.dout(w_dff_B_2oalaXv76_2),.clk(gclk));
	jdff dff_B_b7ePqXwK0_2(.din(w_dff_B_2oalaXv76_2),.dout(w_dff_B_b7ePqXwK0_2),.clk(gclk));
	jdff dff_B_3MM1mVp90_2(.din(w_dff_B_b7ePqXwK0_2),.dout(w_dff_B_3MM1mVp90_2),.clk(gclk));
	jdff dff_B_KInYzAAL3_2(.din(w_dff_B_3MM1mVp90_2),.dout(w_dff_B_KInYzAAL3_2),.clk(gclk));
	jdff dff_B_GxmMdB2Z3_2(.din(w_dff_B_KInYzAAL3_2),.dout(w_dff_B_GxmMdB2Z3_2),.clk(gclk));
	jdff dff_B_Hfon6AiE8_2(.din(w_dff_B_GxmMdB2Z3_2),.dout(w_dff_B_Hfon6AiE8_2),.clk(gclk));
	jdff dff_B_e2miI3D60_2(.din(w_dff_B_Hfon6AiE8_2),.dout(w_dff_B_e2miI3D60_2),.clk(gclk));
	jdff dff_B_YiRbJM8b7_2(.din(w_dff_B_e2miI3D60_2),.dout(w_dff_B_YiRbJM8b7_2),.clk(gclk));
	jdff dff_B_dImp38AW0_2(.din(w_dff_B_YiRbJM8b7_2),.dout(w_dff_B_dImp38AW0_2),.clk(gclk));
	jdff dff_B_N7fAZGqV3_2(.din(w_dff_B_dImp38AW0_2),.dout(w_dff_B_N7fAZGqV3_2),.clk(gclk));
	jdff dff_B_V76RIVTO0_2(.din(w_dff_B_N7fAZGqV3_2),.dout(w_dff_B_V76RIVTO0_2),.clk(gclk));
	jdff dff_B_nntKykwv5_2(.din(w_dff_B_V76RIVTO0_2),.dout(w_dff_B_nntKykwv5_2),.clk(gclk));
	jdff dff_B_SkCr0Hsw8_2(.din(w_dff_B_nntKykwv5_2),.dout(w_dff_B_SkCr0Hsw8_2),.clk(gclk));
	jdff dff_B_N3Gz4a417_2(.din(w_dff_B_SkCr0Hsw8_2),.dout(w_dff_B_N3Gz4a417_2),.clk(gclk));
	jdff dff_B_PKsD9SUp7_2(.din(w_dff_B_N3Gz4a417_2),.dout(w_dff_B_PKsD9SUp7_2),.clk(gclk));
	jdff dff_B_PNtD6FEn9_2(.din(w_dff_B_PKsD9SUp7_2),.dout(w_dff_B_PNtD6FEn9_2),.clk(gclk));
	jdff dff_B_PrzCxOEQ4_2(.din(w_dff_B_PNtD6FEn9_2),.dout(w_dff_B_PrzCxOEQ4_2),.clk(gclk));
	jdff dff_B_JSHBTzFy4_2(.din(n1077),.dout(w_dff_B_JSHBTzFy4_2),.clk(gclk));
	jdff dff_B_4RoCyyc49_1(.din(n1075),.dout(w_dff_B_4RoCyyc49_1),.clk(gclk));
	jdff dff_B_TeSDMvrh9_2(.din(n976),.dout(w_dff_B_TeSDMvrh9_2),.clk(gclk));
	jdff dff_B_aB2ruGhT5_2(.din(w_dff_B_TeSDMvrh9_2),.dout(w_dff_B_aB2ruGhT5_2),.clk(gclk));
	jdff dff_B_tHCvUFej1_2(.din(w_dff_B_aB2ruGhT5_2),.dout(w_dff_B_tHCvUFej1_2),.clk(gclk));
	jdff dff_B_k51qxMxG3_2(.din(w_dff_B_tHCvUFej1_2),.dout(w_dff_B_k51qxMxG3_2),.clk(gclk));
	jdff dff_B_vwTaCo179_2(.din(w_dff_B_k51qxMxG3_2),.dout(w_dff_B_vwTaCo179_2),.clk(gclk));
	jdff dff_B_dmIEIi6K7_2(.din(w_dff_B_vwTaCo179_2),.dout(w_dff_B_dmIEIi6K7_2),.clk(gclk));
	jdff dff_B_NfJJlwcQ6_2(.din(w_dff_B_dmIEIi6K7_2),.dout(w_dff_B_NfJJlwcQ6_2),.clk(gclk));
	jdff dff_B_2ot4aw1P1_2(.din(w_dff_B_NfJJlwcQ6_2),.dout(w_dff_B_2ot4aw1P1_2),.clk(gclk));
	jdff dff_B_DZ5TuKAr0_2(.din(w_dff_B_2ot4aw1P1_2),.dout(w_dff_B_DZ5TuKAr0_2),.clk(gclk));
	jdff dff_B_Qr6KONTB9_2(.din(w_dff_B_DZ5TuKAr0_2),.dout(w_dff_B_Qr6KONTB9_2),.clk(gclk));
	jdff dff_B_D7mpqHaZ9_2(.din(w_dff_B_Qr6KONTB9_2),.dout(w_dff_B_D7mpqHaZ9_2),.clk(gclk));
	jdff dff_B_8ap9XZ2G5_2(.din(w_dff_B_D7mpqHaZ9_2),.dout(w_dff_B_8ap9XZ2G5_2),.clk(gclk));
	jdff dff_B_znAvAf1b6_2(.din(w_dff_B_8ap9XZ2G5_2),.dout(w_dff_B_znAvAf1b6_2),.clk(gclk));
	jdff dff_B_g7Ajp1Jz1_2(.din(w_dff_B_znAvAf1b6_2),.dout(w_dff_B_g7Ajp1Jz1_2),.clk(gclk));
	jdff dff_B_2inuqmvb5_2(.din(w_dff_B_g7Ajp1Jz1_2),.dout(w_dff_B_2inuqmvb5_2),.clk(gclk));
	jdff dff_B_DCbt8AsM8_2(.din(w_dff_B_2inuqmvb5_2),.dout(w_dff_B_DCbt8AsM8_2),.clk(gclk));
	jdff dff_B_4OhSnjHB1_1(.din(n977),.dout(w_dff_B_4OhSnjHB1_1),.clk(gclk));
	jdff dff_B_BTvLNqp24_2(.din(n871),.dout(w_dff_B_BTvLNqp24_2),.clk(gclk));
	jdff dff_B_vTRdyL2n2_2(.din(w_dff_B_BTvLNqp24_2),.dout(w_dff_B_vTRdyL2n2_2),.clk(gclk));
	jdff dff_B_zvqJp2eF7_2(.din(w_dff_B_vTRdyL2n2_2),.dout(w_dff_B_zvqJp2eF7_2),.clk(gclk));
	jdff dff_B_cwdt00yb6_2(.din(w_dff_B_zvqJp2eF7_2),.dout(w_dff_B_cwdt00yb6_2),.clk(gclk));
	jdff dff_B_IswTWwiX8_2(.din(w_dff_B_cwdt00yb6_2),.dout(w_dff_B_IswTWwiX8_2),.clk(gclk));
	jdff dff_B_jxVmJiKd6_2(.din(w_dff_B_IswTWwiX8_2),.dout(w_dff_B_jxVmJiKd6_2),.clk(gclk));
	jdff dff_B_zh7bGbAO1_2(.din(w_dff_B_jxVmJiKd6_2),.dout(w_dff_B_zh7bGbAO1_2),.clk(gclk));
	jdff dff_B_0TuTl3f45_2(.din(w_dff_B_zh7bGbAO1_2),.dout(w_dff_B_0TuTl3f45_2),.clk(gclk));
	jdff dff_B_d1OaOJdv0_2(.din(w_dff_B_0TuTl3f45_2),.dout(w_dff_B_d1OaOJdv0_2),.clk(gclk));
	jdff dff_B_JPghaI0L5_2(.din(w_dff_B_d1OaOJdv0_2),.dout(w_dff_B_JPghaI0L5_2),.clk(gclk));
	jdff dff_B_egHK3uEz1_2(.din(w_dff_B_JPghaI0L5_2),.dout(w_dff_B_egHK3uEz1_2),.clk(gclk));
	jdff dff_B_RZrGdPql2_2(.din(w_dff_B_egHK3uEz1_2),.dout(w_dff_B_RZrGdPql2_2),.clk(gclk));
	jdff dff_B_3yEfr7Fd2_2(.din(w_dff_B_RZrGdPql2_2),.dout(w_dff_B_3yEfr7Fd2_2),.clk(gclk));
	jdff dff_B_ohS8euDz2_2(.din(w_dff_B_3yEfr7Fd2_2),.dout(w_dff_B_ohS8euDz2_2),.clk(gclk));
	jdff dff_B_Z1wAO6IW1_1(.din(n872),.dout(w_dff_B_Z1wAO6IW1_1),.clk(gclk));
	jdff dff_B_hYHZV2MK6_2(.din(n772),.dout(w_dff_B_hYHZV2MK6_2),.clk(gclk));
	jdff dff_B_EoSu7nZR4_2(.din(w_dff_B_hYHZV2MK6_2),.dout(w_dff_B_EoSu7nZR4_2),.clk(gclk));
	jdff dff_B_pQ7rdIDj2_2(.din(w_dff_B_EoSu7nZR4_2),.dout(w_dff_B_pQ7rdIDj2_2),.clk(gclk));
	jdff dff_B_u56fcKA50_2(.din(w_dff_B_pQ7rdIDj2_2),.dout(w_dff_B_u56fcKA50_2),.clk(gclk));
	jdff dff_B_DG8su0CU4_2(.din(w_dff_B_u56fcKA50_2),.dout(w_dff_B_DG8su0CU4_2),.clk(gclk));
	jdff dff_B_YRfhCypi6_2(.din(w_dff_B_DG8su0CU4_2),.dout(w_dff_B_YRfhCypi6_2),.clk(gclk));
	jdff dff_B_Ir9LbLhO6_2(.din(w_dff_B_YRfhCypi6_2),.dout(w_dff_B_Ir9LbLhO6_2),.clk(gclk));
	jdff dff_B_HttjD7nw6_2(.din(w_dff_B_Ir9LbLhO6_2),.dout(w_dff_B_HttjD7nw6_2),.clk(gclk));
	jdff dff_B_DdM4YSNl6_2(.din(w_dff_B_HttjD7nw6_2),.dout(w_dff_B_DdM4YSNl6_2),.clk(gclk));
	jdff dff_B_ojq0lhco6_2(.din(w_dff_B_DdM4YSNl6_2),.dout(w_dff_B_ojq0lhco6_2),.clk(gclk));
	jdff dff_B_SCpfItVk0_2(.din(w_dff_B_ojq0lhco6_2),.dout(w_dff_B_SCpfItVk0_2),.clk(gclk));
	jdff dff_B_GRLdMi0n6_2(.din(w_dff_B_SCpfItVk0_2),.dout(w_dff_B_GRLdMi0n6_2),.clk(gclk));
	jdff dff_B_uCF6h73s2_1(.din(n773),.dout(w_dff_B_uCF6h73s2_1),.clk(gclk));
	jdff dff_B_GQevH8ws1_2(.din(n679),.dout(w_dff_B_GQevH8ws1_2),.clk(gclk));
	jdff dff_B_LNr8B91J1_2(.din(w_dff_B_GQevH8ws1_2),.dout(w_dff_B_LNr8B91J1_2),.clk(gclk));
	jdff dff_B_sF7dip1X2_2(.din(w_dff_B_LNr8B91J1_2),.dout(w_dff_B_sF7dip1X2_2),.clk(gclk));
	jdff dff_B_hHMrYJ236_2(.din(w_dff_B_sF7dip1X2_2),.dout(w_dff_B_hHMrYJ236_2),.clk(gclk));
	jdff dff_B_TsMGOJSZ7_2(.din(w_dff_B_hHMrYJ236_2),.dout(w_dff_B_TsMGOJSZ7_2),.clk(gclk));
	jdff dff_B_ECwcD2uT7_2(.din(w_dff_B_TsMGOJSZ7_2),.dout(w_dff_B_ECwcD2uT7_2),.clk(gclk));
	jdff dff_B_DyxwykNC8_2(.din(w_dff_B_ECwcD2uT7_2),.dout(w_dff_B_DyxwykNC8_2),.clk(gclk));
	jdff dff_B_DFFMty2n4_2(.din(w_dff_B_DyxwykNC8_2),.dout(w_dff_B_DFFMty2n4_2),.clk(gclk));
	jdff dff_B_eRfLbmES2_2(.din(w_dff_B_DFFMty2n4_2),.dout(w_dff_B_eRfLbmES2_2),.clk(gclk));
	jdff dff_B_fhVItzJa8_2(.din(w_dff_B_eRfLbmES2_2),.dout(w_dff_B_fhVItzJa8_2),.clk(gclk));
	jdff dff_B_btSQe1sk0_1(.din(n680),.dout(w_dff_B_btSQe1sk0_1),.clk(gclk));
	jdff dff_B_kYGGRyUY3_2(.din(n593),.dout(w_dff_B_kYGGRyUY3_2),.clk(gclk));
	jdff dff_B_ox39bHL71_2(.din(w_dff_B_kYGGRyUY3_2),.dout(w_dff_B_ox39bHL71_2),.clk(gclk));
	jdff dff_B_Z1Tk8c419_2(.din(w_dff_B_ox39bHL71_2),.dout(w_dff_B_Z1Tk8c419_2),.clk(gclk));
	jdff dff_B_WcfT0iQs9_2(.din(w_dff_B_Z1Tk8c419_2),.dout(w_dff_B_WcfT0iQs9_2),.clk(gclk));
	jdff dff_B_FmNfYIGZ8_2(.din(w_dff_B_WcfT0iQs9_2),.dout(w_dff_B_FmNfYIGZ8_2),.clk(gclk));
	jdff dff_B_uwN240CB0_2(.din(w_dff_B_FmNfYIGZ8_2),.dout(w_dff_B_uwN240CB0_2),.clk(gclk));
	jdff dff_B_JpgEOsly0_2(.din(w_dff_B_uwN240CB0_2),.dout(w_dff_B_JpgEOsly0_2),.clk(gclk));
	jdff dff_B_qnHQNVmE9_2(.din(w_dff_B_JpgEOsly0_2),.dout(w_dff_B_qnHQNVmE9_2),.clk(gclk));
	jdff dff_B_Zo9yzJzN1_1(.din(n594),.dout(w_dff_B_Zo9yzJzN1_1),.clk(gclk));
	jdff dff_B_MTgunAhx5_2(.din(n514),.dout(w_dff_B_MTgunAhx5_2),.clk(gclk));
	jdff dff_B_LxDlauum6_2(.din(w_dff_B_MTgunAhx5_2),.dout(w_dff_B_LxDlauum6_2),.clk(gclk));
	jdff dff_B_OkmFtaPm9_2(.din(w_dff_B_LxDlauum6_2),.dout(w_dff_B_OkmFtaPm9_2),.clk(gclk));
	jdff dff_B_ZQiwqMjc1_2(.din(w_dff_B_OkmFtaPm9_2),.dout(w_dff_B_ZQiwqMjc1_2),.clk(gclk));
	jdff dff_B_O92jqehP3_2(.din(w_dff_B_ZQiwqMjc1_2),.dout(w_dff_B_O92jqehP3_2),.clk(gclk));
	jdff dff_B_4Nkw4hr37_2(.din(w_dff_B_O92jqehP3_2),.dout(w_dff_B_4Nkw4hr37_2),.clk(gclk));
	jdff dff_B_3rRbXLt23_2(.din(n530),.dout(w_dff_B_3rRbXLt23_2),.clk(gclk));
	jdff dff_B_HkCdJwym8_1(.din(n515),.dout(w_dff_B_HkCdJwym8_1),.clk(gclk));
	jdff dff_B_JjdrgagQ2_1(.din(w_dff_B_HkCdJwym8_1),.dout(w_dff_B_JjdrgagQ2_1),.clk(gclk));
	jdff dff_B_K5lJlIMz8_1(.din(w_dff_B_JjdrgagQ2_1),.dout(w_dff_B_K5lJlIMz8_1),.clk(gclk));
	jdff dff_B_bQeuhAse3_1(.din(w_dff_B_K5lJlIMz8_1),.dout(w_dff_B_bQeuhAse3_1),.clk(gclk));
	jdff dff_B_2vmf0QpN2_0(.din(n451),.dout(w_dff_B_2vmf0QpN2_0),.clk(gclk));
	jdff dff_A_kn0zsOHZ1_0(.dout(w_n450_0[0]),.din(w_dff_A_kn0zsOHZ1_0),.clk(gclk));
	jdff dff_A_VSjoUpi55_0(.dout(w_dff_A_kn0zsOHZ1_0),.din(w_dff_A_VSjoUpi55_0),.clk(gclk));
	jdff dff_B_q3fbxToc8_1(.din(n444),.dout(w_dff_B_q3fbxToc8_1),.clk(gclk));
	jdff dff_B_hW2Wvec32_1(.din(w_dff_B_q3fbxToc8_1),.dout(w_dff_B_hW2Wvec32_1),.clk(gclk));
	jdff dff_A_LyIyUKHN6_0(.dout(w_n376_0[0]),.din(w_dff_A_LyIyUKHN6_0),.clk(gclk));
	jdff dff_A_eDaH1P4c2_1(.dout(w_n376_0[1]),.din(w_dff_A_eDaH1P4c2_1),.clk(gclk));
	jdff dff_A_2sY683Rr3_1(.dout(w_dff_A_eDaH1P4c2_1),.din(w_dff_A_2sY683Rr3_1),.clk(gclk));
	jdff dff_A_A2WbjbgF7_1(.dout(w_n442_0[1]),.din(w_dff_A_A2WbjbgF7_1),.clk(gclk));
	jdff dff_A_otQYMIni3_1(.dout(w_dff_A_A2WbjbgF7_1),.din(w_dff_A_otQYMIni3_1),.clk(gclk));
	jdff dff_A_BMghvNX15_1(.dout(w_dff_A_otQYMIni3_1),.din(w_dff_A_BMghvNX15_1),.clk(gclk));
	jdff dff_A_ZUEwSf3U7_1(.dout(w_dff_A_BMghvNX15_1),.din(w_dff_A_ZUEwSf3U7_1),.clk(gclk));
	jdff dff_B_FtolqQ735_2(.din(n1682),.dout(w_dff_B_FtolqQ735_2),.clk(gclk));
	jdff dff_B_oDu8Eos25_1(.din(n1680),.dout(w_dff_B_oDu8Eos25_1),.clk(gclk));
	jdff dff_B_wE04I4wQ7_2(.din(n1628),.dout(w_dff_B_wE04I4wQ7_2),.clk(gclk));
	jdff dff_B_WPoClSER5_2(.din(w_dff_B_wE04I4wQ7_2),.dout(w_dff_B_WPoClSER5_2),.clk(gclk));
	jdff dff_B_9jFKQ7Qe6_2(.din(w_dff_B_WPoClSER5_2),.dout(w_dff_B_9jFKQ7Qe6_2),.clk(gclk));
	jdff dff_B_3vISEgVn9_2(.din(w_dff_B_9jFKQ7Qe6_2),.dout(w_dff_B_3vISEgVn9_2),.clk(gclk));
	jdff dff_B_LMHezgEo1_2(.din(w_dff_B_3vISEgVn9_2),.dout(w_dff_B_LMHezgEo1_2),.clk(gclk));
	jdff dff_B_DrmD3htz3_2(.din(w_dff_B_LMHezgEo1_2),.dout(w_dff_B_DrmD3htz3_2),.clk(gclk));
	jdff dff_B_aRQaRnW97_2(.din(w_dff_B_DrmD3htz3_2),.dout(w_dff_B_aRQaRnW97_2),.clk(gclk));
	jdff dff_B_0J6AqRQK6_2(.din(w_dff_B_aRQaRnW97_2),.dout(w_dff_B_0J6AqRQK6_2),.clk(gclk));
	jdff dff_B_oVV8g6Wz0_2(.din(w_dff_B_0J6AqRQK6_2),.dout(w_dff_B_oVV8g6Wz0_2),.clk(gclk));
	jdff dff_B_b3OkEBx99_2(.din(w_dff_B_oVV8g6Wz0_2),.dout(w_dff_B_b3OkEBx99_2),.clk(gclk));
	jdff dff_B_moH1uWoa4_2(.din(w_dff_B_b3OkEBx99_2),.dout(w_dff_B_moH1uWoa4_2),.clk(gclk));
	jdff dff_B_KOlyZ0ow3_2(.din(w_dff_B_moH1uWoa4_2),.dout(w_dff_B_KOlyZ0ow3_2),.clk(gclk));
	jdff dff_B_l83gPR0X3_2(.din(w_dff_B_KOlyZ0ow3_2),.dout(w_dff_B_l83gPR0X3_2),.clk(gclk));
	jdff dff_B_RDXnum4J2_2(.din(w_dff_B_l83gPR0X3_2),.dout(w_dff_B_RDXnum4J2_2),.clk(gclk));
	jdff dff_B_wDr9hJYf0_2(.din(w_dff_B_RDXnum4J2_2),.dout(w_dff_B_wDr9hJYf0_2),.clk(gclk));
	jdff dff_B_VMaPysuh0_2(.din(w_dff_B_wDr9hJYf0_2),.dout(w_dff_B_VMaPysuh0_2),.clk(gclk));
	jdff dff_B_VlxA28bb9_2(.din(w_dff_B_VMaPysuh0_2),.dout(w_dff_B_VlxA28bb9_2),.clk(gclk));
	jdff dff_B_zUUnFJhj7_2(.din(w_dff_B_VlxA28bb9_2),.dout(w_dff_B_zUUnFJhj7_2),.clk(gclk));
	jdff dff_B_lAzmWaIV7_2(.din(w_dff_B_zUUnFJhj7_2),.dout(w_dff_B_lAzmWaIV7_2),.clk(gclk));
	jdff dff_B_yB6oESIv2_2(.din(w_dff_B_lAzmWaIV7_2),.dout(w_dff_B_yB6oESIv2_2),.clk(gclk));
	jdff dff_B_jwiJ97kX1_2(.din(w_dff_B_yB6oESIv2_2),.dout(w_dff_B_jwiJ97kX1_2),.clk(gclk));
	jdff dff_B_6lEq9Y0Z3_2(.din(w_dff_B_jwiJ97kX1_2),.dout(w_dff_B_6lEq9Y0Z3_2),.clk(gclk));
	jdff dff_B_vqzYn8lU8_2(.din(w_dff_B_6lEq9Y0Z3_2),.dout(w_dff_B_vqzYn8lU8_2),.clk(gclk));
	jdff dff_B_1XG43kcY1_2(.din(w_dff_B_vqzYn8lU8_2),.dout(w_dff_B_1XG43kcY1_2),.clk(gclk));
	jdff dff_B_gKeuf43y5_2(.din(w_dff_B_1XG43kcY1_2),.dout(w_dff_B_gKeuf43y5_2),.clk(gclk));
	jdff dff_B_UVIDGLvI5_2(.din(w_dff_B_gKeuf43y5_2),.dout(w_dff_B_UVIDGLvI5_2),.clk(gclk));
	jdff dff_B_8gZXkZhv1_2(.din(w_dff_B_UVIDGLvI5_2),.dout(w_dff_B_8gZXkZhv1_2),.clk(gclk));
	jdff dff_B_mWvWq0mM1_2(.din(w_dff_B_8gZXkZhv1_2),.dout(w_dff_B_mWvWq0mM1_2),.clk(gclk));
	jdff dff_B_lfFVa1rS3_2(.din(w_dff_B_mWvWq0mM1_2),.dout(w_dff_B_lfFVa1rS3_2),.clk(gclk));
	jdff dff_B_cMm6NwEp9_2(.din(w_dff_B_lfFVa1rS3_2),.dout(w_dff_B_cMm6NwEp9_2),.clk(gclk));
	jdff dff_B_FrkmIl2f8_2(.din(w_dff_B_cMm6NwEp9_2),.dout(w_dff_B_FrkmIl2f8_2),.clk(gclk));
	jdff dff_B_A5xSx0WC3_2(.din(w_dff_B_FrkmIl2f8_2),.dout(w_dff_B_A5xSx0WC3_2),.clk(gclk));
	jdff dff_B_g4GTYxdT2_2(.din(w_dff_B_A5xSx0WC3_2),.dout(w_dff_B_g4GTYxdT2_2),.clk(gclk));
	jdff dff_B_47TwFNvY3_2(.din(w_dff_B_g4GTYxdT2_2),.dout(w_dff_B_47TwFNvY3_2),.clk(gclk));
	jdff dff_B_hJsATW6V2_2(.din(w_dff_B_47TwFNvY3_2),.dout(w_dff_B_hJsATW6V2_2),.clk(gclk));
	jdff dff_B_mJNAisik9_2(.din(w_dff_B_hJsATW6V2_2),.dout(w_dff_B_mJNAisik9_2),.clk(gclk));
	jdff dff_B_0SVjtCIX1_2(.din(w_dff_B_mJNAisik9_2),.dout(w_dff_B_0SVjtCIX1_2),.clk(gclk));
	jdff dff_B_gpdaZKjh0_2(.din(w_dff_B_0SVjtCIX1_2),.dout(w_dff_B_gpdaZKjh0_2),.clk(gclk));
	jdff dff_B_TWMzhGLa5_2(.din(w_dff_B_gpdaZKjh0_2),.dout(w_dff_B_TWMzhGLa5_2),.clk(gclk));
	jdff dff_B_fOOVUDPi4_2(.din(w_dff_B_TWMzhGLa5_2),.dout(w_dff_B_fOOVUDPi4_2),.clk(gclk));
	jdff dff_B_VtmnVXvW9_1(.din(n1678),.dout(w_dff_B_VtmnVXvW9_1),.clk(gclk));
	jdff dff_A_QTN0cg9q0_1(.dout(w_n1631_0[1]),.din(w_dff_A_QTN0cg9q0_1),.clk(gclk));
	jdff dff_B_w79I0pZh7_1(.din(n1629),.dout(w_dff_B_w79I0pZh7_1),.clk(gclk));
	jdff dff_B_pUSpDTaA0_2(.din(n1571),.dout(w_dff_B_pUSpDTaA0_2),.clk(gclk));
	jdff dff_B_GN3mywOV4_2(.din(w_dff_B_pUSpDTaA0_2),.dout(w_dff_B_GN3mywOV4_2),.clk(gclk));
	jdff dff_B_Y27DkaB65_2(.din(w_dff_B_GN3mywOV4_2),.dout(w_dff_B_Y27DkaB65_2),.clk(gclk));
	jdff dff_B_EW2gWXP37_2(.din(w_dff_B_Y27DkaB65_2),.dout(w_dff_B_EW2gWXP37_2),.clk(gclk));
	jdff dff_B_OWesw7EV2_2(.din(w_dff_B_EW2gWXP37_2),.dout(w_dff_B_OWesw7EV2_2),.clk(gclk));
	jdff dff_B_V9dfz1PV0_2(.din(w_dff_B_OWesw7EV2_2),.dout(w_dff_B_V9dfz1PV0_2),.clk(gclk));
	jdff dff_B_jjl6BbRA8_2(.din(w_dff_B_V9dfz1PV0_2),.dout(w_dff_B_jjl6BbRA8_2),.clk(gclk));
	jdff dff_B_TGg6UeiO9_2(.din(w_dff_B_jjl6BbRA8_2),.dout(w_dff_B_TGg6UeiO9_2),.clk(gclk));
	jdff dff_B_Zj5eYONl5_2(.din(w_dff_B_TGg6UeiO9_2),.dout(w_dff_B_Zj5eYONl5_2),.clk(gclk));
	jdff dff_B_y3aVR0YG7_2(.din(w_dff_B_Zj5eYONl5_2),.dout(w_dff_B_y3aVR0YG7_2),.clk(gclk));
	jdff dff_B_HEgBnuS27_2(.din(w_dff_B_y3aVR0YG7_2),.dout(w_dff_B_HEgBnuS27_2),.clk(gclk));
	jdff dff_B_xXvrscyu6_2(.din(w_dff_B_HEgBnuS27_2),.dout(w_dff_B_xXvrscyu6_2),.clk(gclk));
	jdff dff_B_Qp1d1mau4_2(.din(w_dff_B_xXvrscyu6_2),.dout(w_dff_B_Qp1d1mau4_2),.clk(gclk));
	jdff dff_B_lG8w9RrV6_2(.din(w_dff_B_Qp1d1mau4_2),.dout(w_dff_B_lG8w9RrV6_2),.clk(gclk));
	jdff dff_B_9QagDsVE9_2(.din(w_dff_B_lG8w9RrV6_2),.dout(w_dff_B_9QagDsVE9_2),.clk(gclk));
	jdff dff_B_MF1CteWo4_2(.din(w_dff_B_9QagDsVE9_2),.dout(w_dff_B_MF1CteWo4_2),.clk(gclk));
	jdff dff_B_uNMQNpGD1_2(.din(w_dff_B_MF1CteWo4_2),.dout(w_dff_B_uNMQNpGD1_2),.clk(gclk));
	jdff dff_B_zNvTlqqJ1_2(.din(w_dff_B_uNMQNpGD1_2),.dout(w_dff_B_zNvTlqqJ1_2),.clk(gclk));
	jdff dff_B_Pu4h1Rhb2_2(.din(w_dff_B_zNvTlqqJ1_2),.dout(w_dff_B_Pu4h1Rhb2_2),.clk(gclk));
	jdff dff_B_IE5tZrss2_2(.din(w_dff_B_Pu4h1Rhb2_2),.dout(w_dff_B_IE5tZrss2_2),.clk(gclk));
	jdff dff_B_S7q4Qtl86_2(.din(w_dff_B_IE5tZrss2_2),.dout(w_dff_B_S7q4Qtl86_2),.clk(gclk));
	jdff dff_B_GvyM50q32_2(.din(w_dff_B_S7q4Qtl86_2),.dout(w_dff_B_GvyM50q32_2),.clk(gclk));
	jdff dff_B_1NznSJST7_2(.din(w_dff_B_GvyM50q32_2),.dout(w_dff_B_1NznSJST7_2),.clk(gclk));
	jdff dff_B_KdSZogl33_2(.din(w_dff_B_1NznSJST7_2),.dout(w_dff_B_KdSZogl33_2),.clk(gclk));
	jdff dff_B_xeMLRUnC2_2(.din(w_dff_B_KdSZogl33_2),.dout(w_dff_B_xeMLRUnC2_2),.clk(gclk));
	jdff dff_B_SwXlRdzX1_2(.din(w_dff_B_xeMLRUnC2_2),.dout(w_dff_B_SwXlRdzX1_2),.clk(gclk));
	jdff dff_B_ScKyS4B77_2(.din(w_dff_B_SwXlRdzX1_2),.dout(w_dff_B_ScKyS4B77_2),.clk(gclk));
	jdff dff_B_joK65iE04_2(.din(w_dff_B_ScKyS4B77_2),.dout(w_dff_B_joK65iE04_2),.clk(gclk));
	jdff dff_B_QiylpfWj0_2(.din(w_dff_B_joK65iE04_2),.dout(w_dff_B_QiylpfWj0_2),.clk(gclk));
	jdff dff_B_klfPiP2b1_2(.din(w_dff_B_QiylpfWj0_2),.dout(w_dff_B_klfPiP2b1_2),.clk(gclk));
	jdff dff_B_34A0kQTu3_2(.din(w_dff_B_klfPiP2b1_2),.dout(w_dff_B_34A0kQTu3_2),.clk(gclk));
	jdff dff_B_PIJFLx1L5_2(.din(w_dff_B_34A0kQTu3_2),.dout(w_dff_B_PIJFLx1L5_2),.clk(gclk));
	jdff dff_B_prvxyJRV3_2(.din(w_dff_B_PIJFLx1L5_2),.dout(w_dff_B_prvxyJRV3_2),.clk(gclk));
	jdff dff_B_msAlT3NN1_2(.din(w_dff_B_prvxyJRV3_2),.dout(w_dff_B_msAlT3NN1_2),.clk(gclk));
	jdff dff_B_cEZ81KbZ7_2(.din(w_dff_B_msAlT3NN1_2),.dout(w_dff_B_cEZ81KbZ7_2),.clk(gclk));
	jdff dff_B_e9uZd5Xu4_2(.din(n1574),.dout(w_dff_B_e9uZd5Xu4_2),.clk(gclk));
	jdff dff_B_uzlAELXW4_1(.din(n1572),.dout(w_dff_B_uzlAELXW4_1),.clk(gclk));
	jdff dff_B_XGLiY6PA6_2(.din(n1507),.dout(w_dff_B_XGLiY6PA6_2),.clk(gclk));
	jdff dff_B_ST0ofe5k8_2(.din(w_dff_B_XGLiY6PA6_2),.dout(w_dff_B_ST0ofe5k8_2),.clk(gclk));
	jdff dff_B_8jeB2cXW2_2(.din(w_dff_B_ST0ofe5k8_2),.dout(w_dff_B_8jeB2cXW2_2),.clk(gclk));
	jdff dff_B_vdozkldW1_2(.din(w_dff_B_8jeB2cXW2_2),.dout(w_dff_B_vdozkldW1_2),.clk(gclk));
	jdff dff_B_hyhrJQt76_2(.din(w_dff_B_vdozkldW1_2),.dout(w_dff_B_hyhrJQt76_2),.clk(gclk));
	jdff dff_B_d56VUmTU5_2(.din(w_dff_B_hyhrJQt76_2),.dout(w_dff_B_d56VUmTU5_2),.clk(gclk));
	jdff dff_B_uaYRbAyu2_2(.din(w_dff_B_d56VUmTU5_2),.dout(w_dff_B_uaYRbAyu2_2),.clk(gclk));
	jdff dff_B_7Pxqdi6r0_2(.din(w_dff_B_uaYRbAyu2_2),.dout(w_dff_B_7Pxqdi6r0_2),.clk(gclk));
	jdff dff_B_MRxzjgj11_2(.din(w_dff_B_7Pxqdi6r0_2),.dout(w_dff_B_MRxzjgj11_2),.clk(gclk));
	jdff dff_B_FYKSD3Pk9_2(.din(w_dff_B_MRxzjgj11_2),.dout(w_dff_B_FYKSD3Pk9_2),.clk(gclk));
	jdff dff_B_z7P477AF0_2(.din(w_dff_B_FYKSD3Pk9_2),.dout(w_dff_B_z7P477AF0_2),.clk(gclk));
	jdff dff_B_hlM2dhGm6_2(.din(w_dff_B_z7P477AF0_2),.dout(w_dff_B_hlM2dhGm6_2),.clk(gclk));
	jdff dff_B_EWpUSGtz4_2(.din(w_dff_B_hlM2dhGm6_2),.dout(w_dff_B_EWpUSGtz4_2),.clk(gclk));
	jdff dff_B_t9NNhls08_2(.din(w_dff_B_EWpUSGtz4_2),.dout(w_dff_B_t9NNhls08_2),.clk(gclk));
	jdff dff_B_rk4pTLwE0_2(.din(w_dff_B_t9NNhls08_2),.dout(w_dff_B_rk4pTLwE0_2),.clk(gclk));
	jdff dff_B_7wlW9M3z8_2(.din(w_dff_B_rk4pTLwE0_2),.dout(w_dff_B_7wlW9M3z8_2),.clk(gclk));
	jdff dff_B_a7mHvGl83_2(.din(w_dff_B_7wlW9M3z8_2),.dout(w_dff_B_a7mHvGl83_2),.clk(gclk));
	jdff dff_B_HymIFP8n3_2(.din(w_dff_B_a7mHvGl83_2),.dout(w_dff_B_HymIFP8n3_2),.clk(gclk));
	jdff dff_B_DW4G04bT5_2(.din(w_dff_B_HymIFP8n3_2),.dout(w_dff_B_DW4G04bT5_2),.clk(gclk));
	jdff dff_B_rWwPLB758_2(.din(w_dff_B_DW4G04bT5_2),.dout(w_dff_B_rWwPLB758_2),.clk(gclk));
	jdff dff_B_2VQrcCgK2_2(.din(w_dff_B_rWwPLB758_2),.dout(w_dff_B_2VQrcCgK2_2),.clk(gclk));
	jdff dff_B_pA0W8bSL7_2(.din(w_dff_B_2VQrcCgK2_2),.dout(w_dff_B_pA0W8bSL7_2),.clk(gclk));
	jdff dff_B_y9SKUnQx5_2(.din(w_dff_B_pA0W8bSL7_2),.dout(w_dff_B_y9SKUnQx5_2),.clk(gclk));
	jdff dff_B_3HSnwsKf0_2(.din(w_dff_B_y9SKUnQx5_2),.dout(w_dff_B_3HSnwsKf0_2),.clk(gclk));
	jdff dff_B_xspFNcCs8_2(.din(w_dff_B_3HSnwsKf0_2),.dout(w_dff_B_xspFNcCs8_2),.clk(gclk));
	jdff dff_B_uWz50CfM8_2(.din(w_dff_B_xspFNcCs8_2),.dout(w_dff_B_uWz50CfM8_2),.clk(gclk));
	jdff dff_B_PyGURnay0_2(.din(w_dff_B_uWz50CfM8_2),.dout(w_dff_B_PyGURnay0_2),.clk(gclk));
	jdff dff_B_ZaYQw5px6_2(.din(w_dff_B_PyGURnay0_2),.dout(w_dff_B_ZaYQw5px6_2),.clk(gclk));
	jdff dff_B_FVaAM92D7_2(.din(w_dff_B_ZaYQw5px6_2),.dout(w_dff_B_FVaAM92D7_2),.clk(gclk));
	jdff dff_B_I9hJsUs91_2(.din(w_dff_B_FVaAM92D7_2),.dout(w_dff_B_I9hJsUs91_2),.clk(gclk));
	jdff dff_B_alX2ptos8_2(.din(w_dff_B_I9hJsUs91_2),.dout(w_dff_B_alX2ptos8_2),.clk(gclk));
	jdff dff_B_ecNw3eAu0_2(.din(w_dff_B_alX2ptos8_2),.dout(w_dff_B_ecNw3eAu0_2),.clk(gclk));
	jdff dff_B_AZwRkMcO5_2(.din(n1510),.dout(w_dff_B_AZwRkMcO5_2),.clk(gclk));
	jdff dff_B_GPX5xaK20_1(.din(n1508),.dout(w_dff_B_GPX5xaK20_1),.clk(gclk));
	jdff dff_B_whCcbEjm7_2(.din(n1436),.dout(w_dff_B_whCcbEjm7_2),.clk(gclk));
	jdff dff_B_nxNef3lo2_2(.din(w_dff_B_whCcbEjm7_2),.dout(w_dff_B_nxNef3lo2_2),.clk(gclk));
	jdff dff_B_6tPNCA2y3_2(.din(w_dff_B_nxNef3lo2_2),.dout(w_dff_B_6tPNCA2y3_2),.clk(gclk));
	jdff dff_B_dc0nmtWc6_2(.din(w_dff_B_6tPNCA2y3_2),.dout(w_dff_B_dc0nmtWc6_2),.clk(gclk));
	jdff dff_B_4Hn6O43Q7_2(.din(w_dff_B_dc0nmtWc6_2),.dout(w_dff_B_4Hn6O43Q7_2),.clk(gclk));
	jdff dff_B_uu67OFuM1_2(.din(w_dff_B_4Hn6O43Q7_2),.dout(w_dff_B_uu67OFuM1_2),.clk(gclk));
	jdff dff_B_CVAwNBkm8_2(.din(w_dff_B_uu67OFuM1_2),.dout(w_dff_B_CVAwNBkm8_2),.clk(gclk));
	jdff dff_B_RIA7IBCW3_2(.din(w_dff_B_CVAwNBkm8_2),.dout(w_dff_B_RIA7IBCW3_2),.clk(gclk));
	jdff dff_B_K5wy189X4_2(.din(w_dff_B_RIA7IBCW3_2),.dout(w_dff_B_K5wy189X4_2),.clk(gclk));
	jdff dff_B_Uy3DKsy39_2(.din(w_dff_B_K5wy189X4_2),.dout(w_dff_B_Uy3DKsy39_2),.clk(gclk));
	jdff dff_B_kPMyouda2_2(.din(w_dff_B_Uy3DKsy39_2),.dout(w_dff_B_kPMyouda2_2),.clk(gclk));
	jdff dff_B_r1ESw0DD5_2(.din(w_dff_B_kPMyouda2_2),.dout(w_dff_B_r1ESw0DD5_2),.clk(gclk));
	jdff dff_B_BOiVgtA71_2(.din(w_dff_B_r1ESw0DD5_2),.dout(w_dff_B_BOiVgtA71_2),.clk(gclk));
	jdff dff_B_YE6REcEF7_2(.din(w_dff_B_BOiVgtA71_2),.dout(w_dff_B_YE6REcEF7_2),.clk(gclk));
	jdff dff_B_KS0eGR7P0_2(.din(w_dff_B_YE6REcEF7_2),.dout(w_dff_B_KS0eGR7P0_2),.clk(gclk));
	jdff dff_B_3RHtpPH64_2(.din(w_dff_B_KS0eGR7P0_2),.dout(w_dff_B_3RHtpPH64_2),.clk(gclk));
	jdff dff_B_2a2N7mhl7_2(.din(w_dff_B_3RHtpPH64_2),.dout(w_dff_B_2a2N7mhl7_2),.clk(gclk));
	jdff dff_B_rj898B917_2(.din(w_dff_B_2a2N7mhl7_2),.dout(w_dff_B_rj898B917_2),.clk(gclk));
	jdff dff_B_weBxvRr00_2(.din(w_dff_B_rj898B917_2),.dout(w_dff_B_weBxvRr00_2),.clk(gclk));
	jdff dff_B_uL9aGcpt6_2(.din(w_dff_B_weBxvRr00_2),.dout(w_dff_B_uL9aGcpt6_2),.clk(gclk));
	jdff dff_B_YmFRj0EE0_2(.din(w_dff_B_uL9aGcpt6_2),.dout(w_dff_B_YmFRj0EE0_2),.clk(gclk));
	jdff dff_B_FbK8rl8x7_2(.din(w_dff_B_YmFRj0EE0_2),.dout(w_dff_B_FbK8rl8x7_2),.clk(gclk));
	jdff dff_B_2S5DYXY75_2(.din(w_dff_B_FbK8rl8x7_2),.dout(w_dff_B_2S5DYXY75_2),.clk(gclk));
	jdff dff_B_BcnR6s569_2(.din(w_dff_B_2S5DYXY75_2),.dout(w_dff_B_BcnR6s569_2),.clk(gclk));
	jdff dff_B_AoyNyvj77_2(.din(w_dff_B_BcnR6s569_2),.dout(w_dff_B_AoyNyvj77_2),.clk(gclk));
	jdff dff_B_yGFJtCAs3_2(.din(w_dff_B_AoyNyvj77_2),.dout(w_dff_B_yGFJtCAs3_2),.clk(gclk));
	jdff dff_B_YGfIopuj4_2(.din(w_dff_B_yGFJtCAs3_2),.dout(w_dff_B_YGfIopuj4_2),.clk(gclk));
	jdff dff_B_2cFuOeDU0_2(.din(w_dff_B_YGfIopuj4_2),.dout(w_dff_B_2cFuOeDU0_2),.clk(gclk));
	jdff dff_B_aRYoTqZk7_2(.din(w_dff_B_2cFuOeDU0_2),.dout(w_dff_B_aRYoTqZk7_2),.clk(gclk));
	jdff dff_B_F32ynQNJ0_2(.din(n1439),.dout(w_dff_B_F32ynQNJ0_2),.clk(gclk));
	jdff dff_B_D2vrndJ97_1(.din(n1437),.dout(w_dff_B_D2vrndJ97_1),.clk(gclk));
	jdff dff_B_L17nLg5l4_2(.din(n1358),.dout(w_dff_B_L17nLg5l4_2),.clk(gclk));
	jdff dff_B_5blouBsA0_2(.din(w_dff_B_L17nLg5l4_2),.dout(w_dff_B_5blouBsA0_2),.clk(gclk));
	jdff dff_B_JwvTDodC5_2(.din(w_dff_B_5blouBsA0_2),.dout(w_dff_B_JwvTDodC5_2),.clk(gclk));
	jdff dff_B_If3nmpXj2_2(.din(w_dff_B_JwvTDodC5_2),.dout(w_dff_B_If3nmpXj2_2),.clk(gclk));
	jdff dff_B_juTBOYVR3_2(.din(w_dff_B_If3nmpXj2_2),.dout(w_dff_B_juTBOYVR3_2),.clk(gclk));
	jdff dff_B_Ctgey6160_2(.din(w_dff_B_juTBOYVR3_2),.dout(w_dff_B_Ctgey6160_2),.clk(gclk));
	jdff dff_B_TeGskrw05_2(.din(w_dff_B_Ctgey6160_2),.dout(w_dff_B_TeGskrw05_2),.clk(gclk));
	jdff dff_B_38jb5Q205_2(.din(w_dff_B_TeGskrw05_2),.dout(w_dff_B_38jb5Q205_2),.clk(gclk));
	jdff dff_B_bV8NVUoR3_2(.din(w_dff_B_38jb5Q205_2),.dout(w_dff_B_bV8NVUoR3_2),.clk(gclk));
	jdff dff_B_uCV82ucR5_2(.din(w_dff_B_bV8NVUoR3_2),.dout(w_dff_B_uCV82ucR5_2),.clk(gclk));
	jdff dff_B_gscPhUYH3_2(.din(w_dff_B_uCV82ucR5_2),.dout(w_dff_B_gscPhUYH3_2),.clk(gclk));
	jdff dff_B_A3GUBsnS7_2(.din(w_dff_B_gscPhUYH3_2),.dout(w_dff_B_A3GUBsnS7_2),.clk(gclk));
	jdff dff_B_L93BWW0A6_2(.din(w_dff_B_A3GUBsnS7_2),.dout(w_dff_B_L93BWW0A6_2),.clk(gclk));
	jdff dff_B_Q8ePGlag2_2(.din(w_dff_B_L93BWW0A6_2),.dout(w_dff_B_Q8ePGlag2_2),.clk(gclk));
	jdff dff_B_A9V7suDM9_2(.din(w_dff_B_Q8ePGlag2_2),.dout(w_dff_B_A9V7suDM9_2),.clk(gclk));
	jdff dff_B_6AK9eN9L2_2(.din(w_dff_B_A9V7suDM9_2),.dout(w_dff_B_6AK9eN9L2_2),.clk(gclk));
	jdff dff_B_8UbFGlfN6_2(.din(w_dff_B_6AK9eN9L2_2),.dout(w_dff_B_8UbFGlfN6_2),.clk(gclk));
	jdff dff_B_NkJRKOzt5_2(.din(w_dff_B_8UbFGlfN6_2),.dout(w_dff_B_NkJRKOzt5_2),.clk(gclk));
	jdff dff_B_p1pj7nQ12_2(.din(w_dff_B_NkJRKOzt5_2),.dout(w_dff_B_p1pj7nQ12_2),.clk(gclk));
	jdff dff_B_WopICEiV5_2(.din(w_dff_B_p1pj7nQ12_2),.dout(w_dff_B_WopICEiV5_2),.clk(gclk));
	jdff dff_B_jlm51HI61_2(.din(w_dff_B_WopICEiV5_2),.dout(w_dff_B_jlm51HI61_2),.clk(gclk));
	jdff dff_B_YiQsSk0w6_2(.din(w_dff_B_jlm51HI61_2),.dout(w_dff_B_YiQsSk0w6_2),.clk(gclk));
	jdff dff_B_Rj7RXo2o3_2(.din(w_dff_B_YiQsSk0w6_2),.dout(w_dff_B_Rj7RXo2o3_2),.clk(gclk));
	jdff dff_B_ltHDEBBi5_2(.din(w_dff_B_Rj7RXo2o3_2),.dout(w_dff_B_ltHDEBBi5_2),.clk(gclk));
	jdff dff_B_w8o70wwS1_2(.din(w_dff_B_ltHDEBBi5_2),.dout(w_dff_B_w8o70wwS1_2),.clk(gclk));
	jdff dff_B_kV5tHOnr0_2(.din(w_dff_B_w8o70wwS1_2),.dout(w_dff_B_kV5tHOnr0_2),.clk(gclk));
	jdff dff_B_RK8XfEmu7_2(.din(n1361),.dout(w_dff_B_RK8XfEmu7_2),.clk(gclk));
	jdff dff_B_xbndg6UF9_1(.din(n1359),.dout(w_dff_B_xbndg6UF9_1),.clk(gclk));
	jdff dff_B_3duHWKSw1_2(.din(n1273),.dout(w_dff_B_3duHWKSw1_2),.clk(gclk));
	jdff dff_B_hMrCfNmP0_2(.din(w_dff_B_3duHWKSw1_2),.dout(w_dff_B_hMrCfNmP0_2),.clk(gclk));
	jdff dff_B_ued6c8hn6_2(.din(w_dff_B_hMrCfNmP0_2),.dout(w_dff_B_ued6c8hn6_2),.clk(gclk));
	jdff dff_B_0T2T7uX31_2(.din(w_dff_B_ued6c8hn6_2),.dout(w_dff_B_0T2T7uX31_2),.clk(gclk));
	jdff dff_B_K473yoNF6_2(.din(w_dff_B_0T2T7uX31_2),.dout(w_dff_B_K473yoNF6_2),.clk(gclk));
	jdff dff_B_eIqr0LMd6_2(.din(w_dff_B_K473yoNF6_2),.dout(w_dff_B_eIqr0LMd6_2),.clk(gclk));
	jdff dff_B_0MafWtwn9_2(.din(w_dff_B_eIqr0LMd6_2),.dout(w_dff_B_0MafWtwn9_2),.clk(gclk));
	jdff dff_B_HadeiXsy8_2(.din(w_dff_B_0MafWtwn9_2),.dout(w_dff_B_HadeiXsy8_2),.clk(gclk));
	jdff dff_B_k6OJn5kx9_2(.din(w_dff_B_HadeiXsy8_2),.dout(w_dff_B_k6OJn5kx9_2),.clk(gclk));
	jdff dff_B_1dDA4z7V2_2(.din(w_dff_B_k6OJn5kx9_2),.dout(w_dff_B_1dDA4z7V2_2),.clk(gclk));
	jdff dff_B_NkGUXd290_2(.din(w_dff_B_1dDA4z7V2_2),.dout(w_dff_B_NkGUXd290_2),.clk(gclk));
	jdff dff_B_H4ua56G17_2(.din(w_dff_B_NkGUXd290_2),.dout(w_dff_B_H4ua56G17_2),.clk(gclk));
	jdff dff_B_iNgeChwW9_2(.din(w_dff_B_H4ua56G17_2),.dout(w_dff_B_iNgeChwW9_2),.clk(gclk));
	jdff dff_B_dvyf9QtG9_2(.din(w_dff_B_iNgeChwW9_2),.dout(w_dff_B_dvyf9QtG9_2),.clk(gclk));
	jdff dff_B_tD7Grgwh6_2(.din(w_dff_B_dvyf9QtG9_2),.dout(w_dff_B_tD7Grgwh6_2),.clk(gclk));
	jdff dff_B_woIbjkXG8_2(.din(w_dff_B_tD7Grgwh6_2),.dout(w_dff_B_woIbjkXG8_2),.clk(gclk));
	jdff dff_B_JI6S2RWY0_2(.din(w_dff_B_woIbjkXG8_2),.dout(w_dff_B_JI6S2RWY0_2),.clk(gclk));
	jdff dff_B_1gNAIQ9X0_2(.din(w_dff_B_JI6S2RWY0_2),.dout(w_dff_B_1gNAIQ9X0_2),.clk(gclk));
	jdff dff_B_fGeimlpM8_2(.din(w_dff_B_1gNAIQ9X0_2),.dout(w_dff_B_fGeimlpM8_2),.clk(gclk));
	jdff dff_B_dHQ0tyAa9_2(.din(w_dff_B_fGeimlpM8_2),.dout(w_dff_B_dHQ0tyAa9_2),.clk(gclk));
	jdff dff_B_PBiYnNvT5_2(.din(w_dff_B_dHQ0tyAa9_2),.dout(w_dff_B_PBiYnNvT5_2),.clk(gclk));
	jdff dff_B_bBBRdh0W6_2(.din(w_dff_B_PBiYnNvT5_2),.dout(w_dff_B_bBBRdh0W6_2),.clk(gclk));
	jdff dff_B_fZVZwQfO1_2(.din(w_dff_B_bBBRdh0W6_2),.dout(w_dff_B_fZVZwQfO1_2),.clk(gclk));
	jdff dff_B_1zPUAOOj0_2(.din(n1276),.dout(w_dff_B_1zPUAOOj0_2),.clk(gclk));
	jdff dff_B_mq9duBnh9_1(.din(n1274),.dout(w_dff_B_mq9duBnh9_1),.clk(gclk));
	jdff dff_B_qbRJKyut9_2(.din(n1183),.dout(w_dff_B_qbRJKyut9_2),.clk(gclk));
	jdff dff_B_wuosGH5V1_2(.din(w_dff_B_qbRJKyut9_2),.dout(w_dff_B_wuosGH5V1_2),.clk(gclk));
	jdff dff_B_c3XFSywN0_2(.din(w_dff_B_wuosGH5V1_2),.dout(w_dff_B_c3XFSywN0_2),.clk(gclk));
	jdff dff_B_ggIqvUyK8_2(.din(w_dff_B_c3XFSywN0_2),.dout(w_dff_B_ggIqvUyK8_2),.clk(gclk));
	jdff dff_B_bTEMI6yI5_2(.din(w_dff_B_ggIqvUyK8_2),.dout(w_dff_B_bTEMI6yI5_2),.clk(gclk));
	jdff dff_B_A5JwVM7p1_2(.din(w_dff_B_bTEMI6yI5_2),.dout(w_dff_B_A5JwVM7p1_2),.clk(gclk));
	jdff dff_B_1IPvVJBd3_2(.din(w_dff_B_A5JwVM7p1_2),.dout(w_dff_B_1IPvVJBd3_2),.clk(gclk));
	jdff dff_B_3GYeeXMU2_2(.din(w_dff_B_1IPvVJBd3_2),.dout(w_dff_B_3GYeeXMU2_2),.clk(gclk));
	jdff dff_B_RtRMlLV93_2(.din(w_dff_B_3GYeeXMU2_2),.dout(w_dff_B_RtRMlLV93_2),.clk(gclk));
	jdff dff_B_oVkS2rzQ3_2(.din(w_dff_B_RtRMlLV93_2),.dout(w_dff_B_oVkS2rzQ3_2),.clk(gclk));
	jdff dff_B_K4pDD6M35_2(.din(w_dff_B_oVkS2rzQ3_2),.dout(w_dff_B_K4pDD6M35_2),.clk(gclk));
	jdff dff_B_hFaZx0Bc5_2(.din(w_dff_B_K4pDD6M35_2),.dout(w_dff_B_hFaZx0Bc5_2),.clk(gclk));
	jdff dff_B_okyOLNjQ6_2(.din(w_dff_B_hFaZx0Bc5_2),.dout(w_dff_B_okyOLNjQ6_2),.clk(gclk));
	jdff dff_B_Gis1WVFi2_2(.din(w_dff_B_okyOLNjQ6_2),.dout(w_dff_B_Gis1WVFi2_2),.clk(gclk));
	jdff dff_B_h9cdILAj4_2(.din(w_dff_B_Gis1WVFi2_2),.dout(w_dff_B_h9cdILAj4_2),.clk(gclk));
	jdff dff_B_wmlXPwbF6_2(.din(w_dff_B_h9cdILAj4_2),.dout(w_dff_B_wmlXPwbF6_2),.clk(gclk));
	jdff dff_B_aL9HpEFT0_2(.din(w_dff_B_wmlXPwbF6_2),.dout(w_dff_B_aL9HpEFT0_2),.clk(gclk));
	jdff dff_B_8lkL9us34_2(.din(w_dff_B_aL9HpEFT0_2),.dout(w_dff_B_8lkL9us34_2),.clk(gclk));
	jdff dff_B_9cISku7Y0_2(.din(w_dff_B_8lkL9us34_2),.dout(w_dff_B_9cISku7Y0_2),.clk(gclk));
	jdff dff_B_pdMKyQz74_2(.din(w_dff_B_9cISku7Y0_2),.dout(w_dff_B_pdMKyQz74_2),.clk(gclk));
	jdff dff_B_4s9CXQls9_2(.din(n1186),.dout(w_dff_B_4s9CXQls9_2),.clk(gclk));
	jdff dff_B_9Uieaijd3_1(.din(n1184),.dout(w_dff_B_9Uieaijd3_1),.clk(gclk));
	jdff dff_B_Y1aFg7n48_2(.din(n1079),.dout(w_dff_B_Y1aFg7n48_2),.clk(gclk));
	jdff dff_B_Q5WBLFOM6_2(.din(w_dff_B_Y1aFg7n48_2),.dout(w_dff_B_Q5WBLFOM6_2),.clk(gclk));
	jdff dff_B_4CD5K0WO2_2(.din(w_dff_B_Q5WBLFOM6_2),.dout(w_dff_B_4CD5K0WO2_2),.clk(gclk));
	jdff dff_B_xg1Q4P7h1_2(.din(w_dff_B_4CD5K0WO2_2),.dout(w_dff_B_xg1Q4P7h1_2),.clk(gclk));
	jdff dff_B_LOaAFG0N9_2(.din(w_dff_B_xg1Q4P7h1_2),.dout(w_dff_B_LOaAFG0N9_2),.clk(gclk));
	jdff dff_B_IPNKcema4_2(.din(w_dff_B_LOaAFG0N9_2),.dout(w_dff_B_IPNKcema4_2),.clk(gclk));
	jdff dff_B_hXwMf1Ln9_2(.din(w_dff_B_IPNKcema4_2),.dout(w_dff_B_hXwMf1Ln9_2),.clk(gclk));
	jdff dff_B_1bsqlHYF9_2(.din(w_dff_B_hXwMf1Ln9_2),.dout(w_dff_B_1bsqlHYF9_2),.clk(gclk));
	jdff dff_B_McmQJbeL0_2(.din(w_dff_B_1bsqlHYF9_2),.dout(w_dff_B_McmQJbeL0_2),.clk(gclk));
	jdff dff_B_un1QwpFL6_2(.din(w_dff_B_McmQJbeL0_2),.dout(w_dff_B_un1QwpFL6_2),.clk(gclk));
	jdff dff_B_fTUIecfe6_2(.din(w_dff_B_un1QwpFL6_2),.dout(w_dff_B_fTUIecfe6_2),.clk(gclk));
	jdff dff_B_rUBvjqU23_2(.din(w_dff_B_fTUIecfe6_2),.dout(w_dff_B_rUBvjqU23_2),.clk(gclk));
	jdff dff_B_S0QUyd4z4_2(.din(w_dff_B_rUBvjqU23_2),.dout(w_dff_B_S0QUyd4z4_2),.clk(gclk));
	jdff dff_B_cAiFs1Vr8_2(.din(w_dff_B_S0QUyd4z4_2),.dout(w_dff_B_cAiFs1Vr8_2),.clk(gclk));
	jdff dff_B_UVYNXiRD1_2(.din(w_dff_B_cAiFs1Vr8_2),.dout(w_dff_B_UVYNXiRD1_2),.clk(gclk));
	jdff dff_B_CYMYmG617_2(.din(w_dff_B_UVYNXiRD1_2),.dout(w_dff_B_CYMYmG617_2),.clk(gclk));
	jdff dff_B_uRS1Fs5X4_2(.din(w_dff_B_CYMYmG617_2),.dout(w_dff_B_uRS1Fs5X4_2),.clk(gclk));
	jdff dff_B_q9ZmF9Nl0_2(.din(n1082),.dout(w_dff_B_q9ZmF9Nl0_2),.clk(gclk));
	jdff dff_B_HCm4HMBu5_1(.din(n1080),.dout(w_dff_B_HCm4HMBu5_1),.clk(gclk));
	jdff dff_B_q9mQfUMn5_2(.din(n981),.dout(w_dff_B_q9mQfUMn5_2),.clk(gclk));
	jdff dff_B_nfTIO8SG3_2(.din(w_dff_B_q9mQfUMn5_2),.dout(w_dff_B_nfTIO8SG3_2),.clk(gclk));
	jdff dff_B_7vMXlgty7_2(.din(w_dff_B_nfTIO8SG3_2),.dout(w_dff_B_7vMXlgty7_2),.clk(gclk));
	jdff dff_B_zm8HHnEn6_2(.din(w_dff_B_7vMXlgty7_2),.dout(w_dff_B_zm8HHnEn6_2),.clk(gclk));
	jdff dff_B_gcJP6ez38_2(.din(w_dff_B_zm8HHnEn6_2),.dout(w_dff_B_gcJP6ez38_2),.clk(gclk));
	jdff dff_B_tF12xAQA2_2(.din(w_dff_B_gcJP6ez38_2),.dout(w_dff_B_tF12xAQA2_2),.clk(gclk));
	jdff dff_B_zzMGZgxv0_2(.din(w_dff_B_tF12xAQA2_2),.dout(w_dff_B_zzMGZgxv0_2),.clk(gclk));
	jdff dff_B_iagYopDK9_2(.din(w_dff_B_zzMGZgxv0_2),.dout(w_dff_B_iagYopDK9_2),.clk(gclk));
	jdff dff_B_OfSWPD290_2(.din(w_dff_B_iagYopDK9_2),.dout(w_dff_B_OfSWPD290_2),.clk(gclk));
	jdff dff_B_3xQwQFwN0_2(.din(w_dff_B_OfSWPD290_2),.dout(w_dff_B_3xQwQFwN0_2),.clk(gclk));
	jdff dff_B_T1iRrGLI7_2(.din(w_dff_B_3xQwQFwN0_2),.dout(w_dff_B_T1iRrGLI7_2),.clk(gclk));
	jdff dff_B_5LjnzKQR7_2(.din(w_dff_B_T1iRrGLI7_2),.dout(w_dff_B_5LjnzKQR7_2),.clk(gclk));
	jdff dff_B_5u09NmvF9_2(.din(w_dff_B_5LjnzKQR7_2),.dout(w_dff_B_5u09NmvF9_2),.clk(gclk));
	jdff dff_B_QM2ywPH17_2(.din(w_dff_B_5u09NmvF9_2),.dout(w_dff_B_QM2ywPH17_2),.clk(gclk));
	jdff dff_B_n6F9CT944_1(.din(n982),.dout(w_dff_B_n6F9CT944_1),.clk(gclk));
	jdff dff_B_Lq5fEtnU3_2(.din(n876),.dout(w_dff_B_Lq5fEtnU3_2),.clk(gclk));
	jdff dff_B_4psRx6Yd0_2(.din(w_dff_B_Lq5fEtnU3_2),.dout(w_dff_B_4psRx6Yd0_2),.clk(gclk));
	jdff dff_B_Vj1T40aS7_2(.din(w_dff_B_4psRx6Yd0_2),.dout(w_dff_B_Vj1T40aS7_2),.clk(gclk));
	jdff dff_B_2eMXGhJK5_2(.din(w_dff_B_Vj1T40aS7_2),.dout(w_dff_B_2eMXGhJK5_2),.clk(gclk));
	jdff dff_B_PvCWoQ7I2_2(.din(w_dff_B_2eMXGhJK5_2),.dout(w_dff_B_PvCWoQ7I2_2),.clk(gclk));
	jdff dff_B_6PAIGnOV5_2(.din(w_dff_B_PvCWoQ7I2_2),.dout(w_dff_B_6PAIGnOV5_2),.clk(gclk));
	jdff dff_B_Qs6leghL9_2(.din(w_dff_B_6PAIGnOV5_2),.dout(w_dff_B_Qs6leghL9_2),.clk(gclk));
	jdff dff_B_aCo1Nzek7_2(.din(w_dff_B_Qs6leghL9_2),.dout(w_dff_B_aCo1Nzek7_2),.clk(gclk));
	jdff dff_B_2KFS5uS59_2(.din(w_dff_B_aCo1Nzek7_2),.dout(w_dff_B_2KFS5uS59_2),.clk(gclk));
	jdff dff_B_vAsbNvhD8_2(.din(w_dff_B_2KFS5uS59_2),.dout(w_dff_B_vAsbNvhD8_2),.clk(gclk));
	jdff dff_B_JZB4b0q48_2(.din(w_dff_B_vAsbNvhD8_2),.dout(w_dff_B_JZB4b0q48_2),.clk(gclk));
	jdff dff_B_bPAnp4Pw3_2(.din(w_dff_B_JZB4b0q48_2),.dout(w_dff_B_bPAnp4Pw3_2),.clk(gclk));
	jdff dff_B_yZPdh5aS0_1(.din(n877),.dout(w_dff_B_yZPdh5aS0_1),.clk(gclk));
	jdff dff_B_8NERdX2u5_2(.din(n777),.dout(w_dff_B_8NERdX2u5_2),.clk(gclk));
	jdff dff_B_25ePHiwQ0_2(.din(w_dff_B_8NERdX2u5_2),.dout(w_dff_B_25ePHiwQ0_2),.clk(gclk));
	jdff dff_B_OjrspeHH2_2(.din(w_dff_B_25ePHiwQ0_2),.dout(w_dff_B_OjrspeHH2_2),.clk(gclk));
	jdff dff_B_PrMWFye28_2(.din(w_dff_B_OjrspeHH2_2),.dout(w_dff_B_PrMWFye28_2),.clk(gclk));
	jdff dff_B_yrEi0ERg7_2(.din(w_dff_B_PrMWFye28_2),.dout(w_dff_B_yrEi0ERg7_2),.clk(gclk));
	jdff dff_B_hDpMZG5I2_2(.din(w_dff_B_yrEi0ERg7_2),.dout(w_dff_B_hDpMZG5I2_2),.clk(gclk));
	jdff dff_B_KrtJe9nO0_2(.din(w_dff_B_hDpMZG5I2_2),.dout(w_dff_B_KrtJe9nO0_2),.clk(gclk));
	jdff dff_B_OjXLKmvU7_2(.din(w_dff_B_KrtJe9nO0_2),.dout(w_dff_B_OjXLKmvU7_2),.clk(gclk));
	jdff dff_B_vQ5CrLRN0_2(.din(w_dff_B_OjXLKmvU7_2),.dout(w_dff_B_vQ5CrLRN0_2),.clk(gclk));
	jdff dff_B_aUyLW4GW0_2(.din(w_dff_B_vQ5CrLRN0_2),.dout(w_dff_B_aUyLW4GW0_2),.clk(gclk));
	jdff dff_B_9guddiw18_1(.din(n778),.dout(w_dff_B_9guddiw18_1),.clk(gclk));
	jdff dff_B_eKp7kmg04_2(.din(n684),.dout(w_dff_B_eKp7kmg04_2),.clk(gclk));
	jdff dff_B_9WnfpqXH4_2(.din(w_dff_B_eKp7kmg04_2),.dout(w_dff_B_9WnfpqXH4_2),.clk(gclk));
	jdff dff_B_RfXqs3bx6_2(.din(w_dff_B_9WnfpqXH4_2),.dout(w_dff_B_RfXqs3bx6_2),.clk(gclk));
	jdff dff_B_FGSvVmyF6_2(.din(w_dff_B_RfXqs3bx6_2),.dout(w_dff_B_FGSvVmyF6_2),.clk(gclk));
	jdff dff_B_5VFTNBQV9_2(.din(w_dff_B_FGSvVmyF6_2),.dout(w_dff_B_5VFTNBQV9_2),.clk(gclk));
	jdff dff_B_d2WCO8lh7_2(.din(w_dff_B_5VFTNBQV9_2),.dout(w_dff_B_d2WCO8lh7_2),.clk(gclk));
	jdff dff_B_X6Lj8DZw4_2(.din(w_dff_B_d2WCO8lh7_2),.dout(w_dff_B_X6Lj8DZw4_2),.clk(gclk));
	jdff dff_B_BOKcLPJE6_2(.din(w_dff_B_X6Lj8DZw4_2),.dout(w_dff_B_BOKcLPJE6_2),.clk(gclk));
	jdff dff_B_3bznItpR8_1(.din(n685),.dout(w_dff_B_3bznItpR8_1),.clk(gclk));
	jdff dff_B_QskTUZIl3_2(.din(n598),.dout(w_dff_B_QskTUZIl3_2),.clk(gclk));
	jdff dff_B_RYCKGT0Q5_2(.din(w_dff_B_QskTUZIl3_2),.dout(w_dff_B_RYCKGT0Q5_2),.clk(gclk));
	jdff dff_B_sJ6bMRPw3_2(.din(w_dff_B_RYCKGT0Q5_2),.dout(w_dff_B_sJ6bMRPw3_2),.clk(gclk));
	jdff dff_B_biN26TeG1_2(.din(w_dff_B_sJ6bMRPw3_2),.dout(w_dff_B_biN26TeG1_2),.clk(gclk));
	jdff dff_B_wRKrBqAU8_2(.din(w_dff_B_biN26TeG1_2),.dout(w_dff_B_wRKrBqAU8_2),.clk(gclk));
	jdff dff_B_VWcRMS4Q8_2(.din(w_dff_B_wRKrBqAU8_2),.dout(w_dff_B_VWcRMS4Q8_2),.clk(gclk));
	jdff dff_B_myQNXNk33_2(.din(n614),.dout(w_dff_B_myQNXNk33_2),.clk(gclk));
	jdff dff_B_Lrk1rPAU7_1(.din(n599),.dout(w_dff_B_Lrk1rPAU7_1),.clk(gclk));
	jdff dff_B_kFdm4MWi7_1(.din(w_dff_B_Lrk1rPAU7_1),.dout(w_dff_B_kFdm4MWi7_1),.clk(gclk));
	jdff dff_B_vvLap90t0_1(.din(w_dff_B_kFdm4MWi7_1),.dout(w_dff_B_vvLap90t0_1),.clk(gclk));
	jdff dff_B_SinQdaEY4_1(.din(w_dff_B_vvLap90t0_1),.dout(w_dff_B_SinQdaEY4_1),.clk(gclk));
	jdff dff_B_46YEwWPG7_0(.din(n528),.dout(w_dff_B_46YEwWPG7_0),.clk(gclk));
	jdff dff_A_7gZ8IHFB9_0(.dout(w_n527_0[0]),.din(w_dff_A_7gZ8IHFB9_0),.clk(gclk));
	jdff dff_A_KFl8vlWw0_0(.dout(w_dff_A_7gZ8IHFB9_0),.din(w_dff_A_KFl8vlWw0_0),.clk(gclk));
	jdff dff_B_DXAcwMA30_1(.din(n521),.dout(w_dff_B_DXAcwMA30_1),.clk(gclk));
	jdff dff_B_edoKP4GI5_1(.din(w_dff_B_DXAcwMA30_1),.dout(w_dff_B_edoKP4GI5_1),.clk(gclk));
	jdff dff_A_HhWBU4898_0(.dout(w_n446_0[0]),.din(w_dff_A_HhWBU4898_0),.clk(gclk));
	jdff dff_A_lAmDUymv7_1(.dout(w_n446_0[1]),.din(w_dff_A_lAmDUymv7_1),.clk(gclk));
	jdff dff_A_2TJbBS0Z7_1(.dout(w_dff_A_lAmDUymv7_1),.din(w_dff_A_2TJbBS0Z7_1),.clk(gclk));
	jdff dff_A_FRrxhEYW4_1(.dout(w_n519_0[1]),.din(w_dff_A_FRrxhEYW4_1),.clk(gclk));
	jdff dff_A_Q7cGH8RO6_1(.dout(w_dff_A_FRrxhEYW4_1),.din(w_dff_A_Q7cGH8RO6_1),.clk(gclk));
	jdff dff_A_p5LVvmLl1_1(.dout(w_dff_A_Q7cGH8RO6_1),.din(w_dff_A_p5LVvmLl1_1),.clk(gclk));
	jdff dff_A_RG9ph2SF1_1(.dout(w_dff_A_p5LVvmLl1_1),.din(w_dff_A_RG9ph2SF1_1),.clk(gclk));
	jdff dff_B_wybVeYra2_1(.din(n1760),.dout(w_dff_B_wybVeYra2_1),.clk(gclk));
	jdff dff_A_u5pAxSPk8_1(.dout(w_n1728_0[1]),.din(w_dff_A_u5pAxSPk8_1),.clk(gclk));
	jdff dff_B_qjFxCdra6_1(.din(n1726),.dout(w_dff_B_qjFxCdra6_1),.clk(gclk));
	jdff dff_B_yCkoQuUi0_2(.din(n1684),.dout(w_dff_B_yCkoQuUi0_2),.clk(gclk));
	jdff dff_B_1e03jPNi0_2(.din(w_dff_B_yCkoQuUi0_2),.dout(w_dff_B_1e03jPNi0_2),.clk(gclk));
	jdff dff_B_xQoFEX040_2(.din(w_dff_B_1e03jPNi0_2),.dout(w_dff_B_xQoFEX040_2),.clk(gclk));
	jdff dff_B_ra0NijEe4_2(.din(w_dff_B_xQoFEX040_2),.dout(w_dff_B_ra0NijEe4_2),.clk(gclk));
	jdff dff_B_UaMnAFWO9_2(.din(w_dff_B_ra0NijEe4_2),.dout(w_dff_B_UaMnAFWO9_2),.clk(gclk));
	jdff dff_B_qE9jf3qt6_2(.din(w_dff_B_UaMnAFWO9_2),.dout(w_dff_B_qE9jf3qt6_2),.clk(gclk));
	jdff dff_B_PUhi8Dkh0_2(.din(w_dff_B_qE9jf3qt6_2),.dout(w_dff_B_PUhi8Dkh0_2),.clk(gclk));
	jdff dff_B_RF9PSkZe0_2(.din(w_dff_B_PUhi8Dkh0_2),.dout(w_dff_B_RF9PSkZe0_2),.clk(gclk));
	jdff dff_B_kcai8zi98_2(.din(w_dff_B_RF9PSkZe0_2),.dout(w_dff_B_kcai8zi98_2),.clk(gclk));
	jdff dff_B_t9f1Af0y4_2(.din(w_dff_B_kcai8zi98_2),.dout(w_dff_B_t9f1Af0y4_2),.clk(gclk));
	jdff dff_B_iw2sIcTV5_2(.din(w_dff_B_t9f1Af0y4_2),.dout(w_dff_B_iw2sIcTV5_2),.clk(gclk));
	jdff dff_B_2IF9iQa65_2(.din(w_dff_B_iw2sIcTV5_2),.dout(w_dff_B_2IF9iQa65_2),.clk(gclk));
	jdff dff_B_sjjoRjtA5_2(.din(w_dff_B_2IF9iQa65_2),.dout(w_dff_B_sjjoRjtA5_2),.clk(gclk));
	jdff dff_B_OdVFeRCh5_2(.din(w_dff_B_sjjoRjtA5_2),.dout(w_dff_B_OdVFeRCh5_2),.clk(gclk));
	jdff dff_B_5FTypbtR2_2(.din(w_dff_B_OdVFeRCh5_2),.dout(w_dff_B_5FTypbtR2_2),.clk(gclk));
	jdff dff_B_ch4Q0btC4_2(.din(w_dff_B_5FTypbtR2_2),.dout(w_dff_B_ch4Q0btC4_2),.clk(gclk));
	jdff dff_B_Q97Vn3KM9_2(.din(w_dff_B_ch4Q0btC4_2),.dout(w_dff_B_Q97Vn3KM9_2),.clk(gclk));
	jdff dff_B_SGvt6UJa9_2(.din(w_dff_B_Q97Vn3KM9_2),.dout(w_dff_B_SGvt6UJa9_2),.clk(gclk));
	jdff dff_B_5fu915K48_2(.din(w_dff_B_SGvt6UJa9_2),.dout(w_dff_B_5fu915K48_2),.clk(gclk));
	jdff dff_B_6pFmFVng7_2(.din(w_dff_B_5fu915K48_2),.dout(w_dff_B_6pFmFVng7_2),.clk(gclk));
	jdff dff_B_VwfjHoz96_2(.din(w_dff_B_6pFmFVng7_2),.dout(w_dff_B_VwfjHoz96_2),.clk(gclk));
	jdff dff_B_GYtKx0dE7_2(.din(w_dff_B_VwfjHoz96_2),.dout(w_dff_B_GYtKx0dE7_2),.clk(gclk));
	jdff dff_B_KELZep1v7_2(.din(w_dff_B_GYtKx0dE7_2),.dout(w_dff_B_KELZep1v7_2),.clk(gclk));
	jdff dff_B_VNolA4Gw4_2(.din(w_dff_B_KELZep1v7_2),.dout(w_dff_B_VNolA4Gw4_2),.clk(gclk));
	jdff dff_B_OpZJGWqX4_2(.din(w_dff_B_VNolA4Gw4_2),.dout(w_dff_B_OpZJGWqX4_2),.clk(gclk));
	jdff dff_B_rAV5wLlQ9_2(.din(w_dff_B_OpZJGWqX4_2),.dout(w_dff_B_rAV5wLlQ9_2),.clk(gclk));
	jdff dff_B_QVAfIkqJ5_2(.din(w_dff_B_rAV5wLlQ9_2),.dout(w_dff_B_QVAfIkqJ5_2),.clk(gclk));
	jdff dff_B_TYnkcW1S4_2(.din(w_dff_B_QVAfIkqJ5_2),.dout(w_dff_B_TYnkcW1S4_2),.clk(gclk));
	jdff dff_B_6T2ExHXD0_2(.din(w_dff_B_TYnkcW1S4_2),.dout(w_dff_B_6T2ExHXD0_2),.clk(gclk));
	jdff dff_B_ZM7cu7DM2_2(.din(w_dff_B_6T2ExHXD0_2),.dout(w_dff_B_ZM7cu7DM2_2),.clk(gclk));
	jdff dff_B_OrqWsJcW6_2(.din(w_dff_B_ZM7cu7DM2_2),.dout(w_dff_B_OrqWsJcW6_2),.clk(gclk));
	jdff dff_B_A2h5ueLQ4_2(.din(w_dff_B_OrqWsJcW6_2),.dout(w_dff_B_A2h5ueLQ4_2),.clk(gclk));
	jdff dff_B_Vba05DfR4_2(.din(w_dff_B_A2h5ueLQ4_2),.dout(w_dff_B_Vba05DfR4_2),.clk(gclk));
	jdff dff_B_djfyHTtY4_2(.din(w_dff_B_Vba05DfR4_2),.dout(w_dff_B_djfyHTtY4_2),.clk(gclk));
	jdff dff_B_CmAepxs86_2(.din(w_dff_B_djfyHTtY4_2),.dout(w_dff_B_CmAepxs86_2),.clk(gclk));
	jdff dff_B_1QVlvKW01_2(.din(w_dff_B_CmAepxs86_2),.dout(w_dff_B_1QVlvKW01_2),.clk(gclk));
	jdff dff_B_8tTAcvvi7_2(.din(w_dff_B_1QVlvKW01_2),.dout(w_dff_B_8tTAcvvi7_2),.clk(gclk));
	jdff dff_B_TWgjBk507_2(.din(w_dff_B_8tTAcvvi7_2),.dout(w_dff_B_TWgjBk507_2),.clk(gclk));
	jdff dff_B_gMcNfZFB1_2(.din(w_dff_B_TWgjBk507_2),.dout(w_dff_B_gMcNfZFB1_2),.clk(gclk));
	jdff dff_B_ns7ZlvK11_2(.din(n1687),.dout(w_dff_B_ns7ZlvK11_2),.clk(gclk));
	jdff dff_B_UJvMBvYk0_1(.din(n1685),.dout(w_dff_B_UJvMBvYk0_1),.clk(gclk));
	jdff dff_B_EKvOAogf7_2(.din(n1633),.dout(w_dff_B_EKvOAogf7_2),.clk(gclk));
	jdff dff_B_rEQ7fuDk2_2(.din(w_dff_B_EKvOAogf7_2),.dout(w_dff_B_rEQ7fuDk2_2),.clk(gclk));
	jdff dff_B_VHdlrsMb1_2(.din(w_dff_B_rEQ7fuDk2_2),.dout(w_dff_B_VHdlrsMb1_2),.clk(gclk));
	jdff dff_B_oPHqpkro3_2(.din(w_dff_B_VHdlrsMb1_2),.dout(w_dff_B_oPHqpkro3_2),.clk(gclk));
	jdff dff_B_NDNbkwMM0_2(.din(w_dff_B_oPHqpkro3_2),.dout(w_dff_B_NDNbkwMM0_2),.clk(gclk));
	jdff dff_B_MNBCwN6r7_2(.din(w_dff_B_NDNbkwMM0_2),.dout(w_dff_B_MNBCwN6r7_2),.clk(gclk));
	jdff dff_B_hvAPfKwF1_2(.din(w_dff_B_MNBCwN6r7_2),.dout(w_dff_B_hvAPfKwF1_2),.clk(gclk));
	jdff dff_B_3BYyu9rc2_2(.din(w_dff_B_hvAPfKwF1_2),.dout(w_dff_B_3BYyu9rc2_2),.clk(gclk));
	jdff dff_B_JPztbNPO0_2(.din(w_dff_B_3BYyu9rc2_2),.dout(w_dff_B_JPztbNPO0_2),.clk(gclk));
	jdff dff_B_NgSs98cJ7_2(.din(w_dff_B_JPztbNPO0_2),.dout(w_dff_B_NgSs98cJ7_2),.clk(gclk));
	jdff dff_B_kNfAVgwe7_2(.din(w_dff_B_NgSs98cJ7_2),.dout(w_dff_B_kNfAVgwe7_2),.clk(gclk));
	jdff dff_B_bGUoieEQ3_2(.din(w_dff_B_kNfAVgwe7_2),.dout(w_dff_B_bGUoieEQ3_2),.clk(gclk));
	jdff dff_B_RZa459qO5_2(.din(w_dff_B_bGUoieEQ3_2),.dout(w_dff_B_RZa459qO5_2),.clk(gclk));
	jdff dff_B_2FNNks7r0_2(.din(w_dff_B_RZa459qO5_2),.dout(w_dff_B_2FNNks7r0_2),.clk(gclk));
	jdff dff_B_QhpERBK61_2(.din(w_dff_B_2FNNks7r0_2),.dout(w_dff_B_QhpERBK61_2),.clk(gclk));
	jdff dff_B_7tr5QZs43_2(.din(w_dff_B_QhpERBK61_2),.dout(w_dff_B_7tr5QZs43_2),.clk(gclk));
	jdff dff_B_wVrT1kfe4_2(.din(w_dff_B_7tr5QZs43_2),.dout(w_dff_B_wVrT1kfe4_2),.clk(gclk));
	jdff dff_B_k7dh23Rn4_2(.din(w_dff_B_wVrT1kfe4_2),.dout(w_dff_B_k7dh23Rn4_2),.clk(gclk));
	jdff dff_B_xIQTt2et3_2(.din(w_dff_B_k7dh23Rn4_2),.dout(w_dff_B_xIQTt2et3_2),.clk(gclk));
	jdff dff_B_rK5x8xpK2_2(.din(w_dff_B_xIQTt2et3_2),.dout(w_dff_B_rK5x8xpK2_2),.clk(gclk));
	jdff dff_B_p2ixqy236_2(.din(w_dff_B_rK5x8xpK2_2),.dout(w_dff_B_p2ixqy236_2),.clk(gclk));
	jdff dff_B_MKbRpjeb4_2(.din(w_dff_B_p2ixqy236_2),.dout(w_dff_B_MKbRpjeb4_2),.clk(gclk));
	jdff dff_B_nL4qBlji4_2(.din(w_dff_B_MKbRpjeb4_2),.dout(w_dff_B_nL4qBlji4_2),.clk(gclk));
	jdff dff_B_YTOHoNPs5_2(.din(w_dff_B_nL4qBlji4_2),.dout(w_dff_B_YTOHoNPs5_2),.clk(gclk));
	jdff dff_B_L5f6J1xD0_2(.din(w_dff_B_YTOHoNPs5_2),.dout(w_dff_B_L5f6J1xD0_2),.clk(gclk));
	jdff dff_B_tBj7tZXG6_2(.din(w_dff_B_L5f6J1xD0_2),.dout(w_dff_B_tBj7tZXG6_2),.clk(gclk));
	jdff dff_B_5d7FUVW01_2(.din(w_dff_B_tBj7tZXG6_2),.dout(w_dff_B_5d7FUVW01_2),.clk(gclk));
	jdff dff_B_FkjliwCP0_2(.din(w_dff_B_5d7FUVW01_2),.dout(w_dff_B_FkjliwCP0_2),.clk(gclk));
	jdff dff_B_35VTTjpI3_2(.din(w_dff_B_FkjliwCP0_2),.dout(w_dff_B_35VTTjpI3_2),.clk(gclk));
	jdff dff_B_XbnCMaL31_2(.din(w_dff_B_35VTTjpI3_2),.dout(w_dff_B_XbnCMaL31_2),.clk(gclk));
	jdff dff_B_ldc8JbMJ1_2(.din(w_dff_B_XbnCMaL31_2),.dout(w_dff_B_ldc8JbMJ1_2),.clk(gclk));
	jdff dff_B_l5SJSHRB9_2(.din(w_dff_B_ldc8JbMJ1_2),.dout(w_dff_B_l5SJSHRB9_2),.clk(gclk));
	jdff dff_B_Ltf8FQDi6_2(.din(w_dff_B_l5SJSHRB9_2),.dout(w_dff_B_Ltf8FQDi6_2),.clk(gclk));
	jdff dff_B_PrRunnAa2_2(.din(w_dff_B_Ltf8FQDi6_2),.dout(w_dff_B_PrRunnAa2_2),.clk(gclk));
	jdff dff_B_Bde1EA6x9_2(.din(w_dff_B_PrRunnAa2_2),.dout(w_dff_B_Bde1EA6x9_2),.clk(gclk));
	jdff dff_B_76gp0Rog3_2(.din(w_dff_B_Bde1EA6x9_2),.dout(w_dff_B_76gp0Rog3_2),.clk(gclk));
	jdff dff_B_iECabImR9_2(.din(n1636),.dout(w_dff_B_iECabImR9_2),.clk(gclk));
	jdff dff_B_nZYIJf9U5_1(.din(n1634),.dout(w_dff_B_nZYIJf9U5_1),.clk(gclk));
	jdff dff_B_hAWd6X2I7_2(.din(n1576),.dout(w_dff_B_hAWd6X2I7_2),.clk(gclk));
	jdff dff_B_3BXniUrU8_2(.din(w_dff_B_hAWd6X2I7_2),.dout(w_dff_B_3BXniUrU8_2),.clk(gclk));
	jdff dff_B_1tTLeYlX7_2(.din(w_dff_B_3BXniUrU8_2),.dout(w_dff_B_1tTLeYlX7_2),.clk(gclk));
	jdff dff_B_D4Ci9jFe0_2(.din(w_dff_B_1tTLeYlX7_2),.dout(w_dff_B_D4Ci9jFe0_2),.clk(gclk));
	jdff dff_B_x38QwtGm5_2(.din(w_dff_B_D4Ci9jFe0_2),.dout(w_dff_B_x38QwtGm5_2),.clk(gclk));
	jdff dff_B_ogC7HuXu1_2(.din(w_dff_B_x38QwtGm5_2),.dout(w_dff_B_ogC7HuXu1_2),.clk(gclk));
	jdff dff_B_ttQoC9nM3_2(.din(w_dff_B_ogC7HuXu1_2),.dout(w_dff_B_ttQoC9nM3_2),.clk(gclk));
	jdff dff_B_TMxwLvs78_2(.din(w_dff_B_ttQoC9nM3_2),.dout(w_dff_B_TMxwLvs78_2),.clk(gclk));
	jdff dff_B_NZA6LmIg5_2(.din(w_dff_B_TMxwLvs78_2),.dout(w_dff_B_NZA6LmIg5_2),.clk(gclk));
	jdff dff_B_v8avHYxQ2_2(.din(w_dff_B_NZA6LmIg5_2),.dout(w_dff_B_v8avHYxQ2_2),.clk(gclk));
	jdff dff_B_BqwtLHPy4_2(.din(w_dff_B_v8avHYxQ2_2),.dout(w_dff_B_BqwtLHPy4_2),.clk(gclk));
	jdff dff_B_Ls9wD5yV7_2(.din(w_dff_B_BqwtLHPy4_2),.dout(w_dff_B_Ls9wD5yV7_2),.clk(gclk));
	jdff dff_B_sqKeiqba4_2(.din(w_dff_B_Ls9wD5yV7_2),.dout(w_dff_B_sqKeiqba4_2),.clk(gclk));
	jdff dff_B_uZxK1mEw5_2(.din(w_dff_B_sqKeiqba4_2),.dout(w_dff_B_uZxK1mEw5_2),.clk(gclk));
	jdff dff_B_l02ux8P57_2(.din(w_dff_B_uZxK1mEw5_2),.dout(w_dff_B_l02ux8P57_2),.clk(gclk));
	jdff dff_B_VTXcpGno5_2(.din(w_dff_B_l02ux8P57_2),.dout(w_dff_B_VTXcpGno5_2),.clk(gclk));
	jdff dff_B_UMHsvwog6_2(.din(w_dff_B_VTXcpGno5_2),.dout(w_dff_B_UMHsvwog6_2),.clk(gclk));
	jdff dff_B_uf70UhdU7_2(.din(w_dff_B_UMHsvwog6_2),.dout(w_dff_B_uf70UhdU7_2),.clk(gclk));
	jdff dff_B_WIREeHOA0_2(.din(w_dff_B_uf70UhdU7_2),.dout(w_dff_B_WIREeHOA0_2),.clk(gclk));
	jdff dff_B_Pbyvcw4L7_2(.din(w_dff_B_WIREeHOA0_2),.dout(w_dff_B_Pbyvcw4L7_2),.clk(gclk));
	jdff dff_B_TDG2Xwug7_2(.din(w_dff_B_Pbyvcw4L7_2),.dout(w_dff_B_TDG2Xwug7_2),.clk(gclk));
	jdff dff_B_JPFmGs7i0_2(.din(w_dff_B_TDG2Xwug7_2),.dout(w_dff_B_JPFmGs7i0_2),.clk(gclk));
	jdff dff_B_yXhAVOAH3_2(.din(w_dff_B_JPFmGs7i0_2),.dout(w_dff_B_yXhAVOAH3_2),.clk(gclk));
	jdff dff_B_nB63w51U6_2(.din(w_dff_B_yXhAVOAH3_2),.dout(w_dff_B_nB63w51U6_2),.clk(gclk));
	jdff dff_B_MFAq0b0S3_2(.din(w_dff_B_nB63w51U6_2),.dout(w_dff_B_MFAq0b0S3_2),.clk(gclk));
	jdff dff_B_zMgc9C2y5_2(.din(w_dff_B_MFAq0b0S3_2),.dout(w_dff_B_zMgc9C2y5_2),.clk(gclk));
	jdff dff_B_gq0HB0fj5_2(.din(w_dff_B_zMgc9C2y5_2),.dout(w_dff_B_gq0HB0fj5_2),.clk(gclk));
	jdff dff_B_i1yHj2xk0_2(.din(w_dff_B_gq0HB0fj5_2),.dout(w_dff_B_i1yHj2xk0_2),.clk(gclk));
	jdff dff_B_g5n5vMzb1_2(.din(w_dff_B_i1yHj2xk0_2),.dout(w_dff_B_g5n5vMzb1_2),.clk(gclk));
	jdff dff_B_Lhsb3wVl7_2(.din(w_dff_B_g5n5vMzb1_2),.dout(w_dff_B_Lhsb3wVl7_2),.clk(gclk));
	jdff dff_B_wGzqms531_2(.din(w_dff_B_Lhsb3wVl7_2),.dout(w_dff_B_wGzqms531_2),.clk(gclk));
	jdff dff_B_L2DbcLkm2_2(.din(w_dff_B_wGzqms531_2),.dout(w_dff_B_L2DbcLkm2_2),.clk(gclk));
	jdff dff_B_MoBDJCAb9_2(.din(w_dff_B_L2DbcLkm2_2),.dout(w_dff_B_MoBDJCAb9_2),.clk(gclk));
	jdff dff_B_57WarLly3_2(.din(n1579),.dout(w_dff_B_57WarLly3_2),.clk(gclk));
	jdff dff_B_jYStSG8v5_1(.din(n1577),.dout(w_dff_B_jYStSG8v5_1),.clk(gclk));
	jdff dff_B_xqSHurj93_2(.din(n1512),.dout(w_dff_B_xqSHurj93_2),.clk(gclk));
	jdff dff_B_6iikLR6j0_2(.din(w_dff_B_xqSHurj93_2),.dout(w_dff_B_6iikLR6j0_2),.clk(gclk));
	jdff dff_B_nXIcOcua4_2(.din(w_dff_B_6iikLR6j0_2),.dout(w_dff_B_nXIcOcua4_2),.clk(gclk));
	jdff dff_B_pm0H1Snv1_2(.din(w_dff_B_nXIcOcua4_2),.dout(w_dff_B_pm0H1Snv1_2),.clk(gclk));
	jdff dff_B_pDswfDCN9_2(.din(w_dff_B_pm0H1Snv1_2),.dout(w_dff_B_pDswfDCN9_2),.clk(gclk));
	jdff dff_B_ygak8jyn8_2(.din(w_dff_B_pDswfDCN9_2),.dout(w_dff_B_ygak8jyn8_2),.clk(gclk));
	jdff dff_B_gqoH7ibT2_2(.din(w_dff_B_ygak8jyn8_2),.dout(w_dff_B_gqoH7ibT2_2),.clk(gclk));
	jdff dff_B_TteqE1v72_2(.din(w_dff_B_gqoH7ibT2_2),.dout(w_dff_B_TteqE1v72_2),.clk(gclk));
	jdff dff_B_CFsi77i09_2(.din(w_dff_B_TteqE1v72_2),.dout(w_dff_B_CFsi77i09_2),.clk(gclk));
	jdff dff_B_WknhPoEQ6_2(.din(w_dff_B_CFsi77i09_2),.dout(w_dff_B_WknhPoEQ6_2),.clk(gclk));
	jdff dff_B_5Cuul0bY8_2(.din(w_dff_B_WknhPoEQ6_2),.dout(w_dff_B_5Cuul0bY8_2),.clk(gclk));
	jdff dff_B_TDajjuti9_2(.din(w_dff_B_5Cuul0bY8_2),.dout(w_dff_B_TDajjuti9_2),.clk(gclk));
	jdff dff_B_dETZ3SFf3_2(.din(w_dff_B_TDajjuti9_2),.dout(w_dff_B_dETZ3SFf3_2),.clk(gclk));
	jdff dff_B_fY1hOuYd8_2(.din(w_dff_B_dETZ3SFf3_2),.dout(w_dff_B_fY1hOuYd8_2),.clk(gclk));
	jdff dff_B_CFjbB4Ce4_2(.din(w_dff_B_fY1hOuYd8_2),.dout(w_dff_B_CFjbB4Ce4_2),.clk(gclk));
	jdff dff_B_Nvx1jjfw8_2(.din(w_dff_B_CFjbB4Ce4_2),.dout(w_dff_B_Nvx1jjfw8_2),.clk(gclk));
	jdff dff_B_v4vpzgSS8_2(.din(w_dff_B_Nvx1jjfw8_2),.dout(w_dff_B_v4vpzgSS8_2),.clk(gclk));
	jdff dff_B_FmWSi48O6_2(.din(w_dff_B_v4vpzgSS8_2),.dout(w_dff_B_FmWSi48O6_2),.clk(gclk));
	jdff dff_B_uACavA1d0_2(.din(w_dff_B_FmWSi48O6_2),.dout(w_dff_B_uACavA1d0_2),.clk(gclk));
	jdff dff_B_81NOX0dO1_2(.din(w_dff_B_uACavA1d0_2),.dout(w_dff_B_81NOX0dO1_2),.clk(gclk));
	jdff dff_B_eVpWkW8i4_2(.din(w_dff_B_81NOX0dO1_2),.dout(w_dff_B_eVpWkW8i4_2),.clk(gclk));
	jdff dff_B_pN7WG8NT2_2(.din(w_dff_B_eVpWkW8i4_2),.dout(w_dff_B_pN7WG8NT2_2),.clk(gclk));
	jdff dff_B_7YCPFTpR1_2(.din(w_dff_B_pN7WG8NT2_2),.dout(w_dff_B_7YCPFTpR1_2),.clk(gclk));
	jdff dff_B_ffcm9BjM2_2(.din(w_dff_B_7YCPFTpR1_2),.dout(w_dff_B_ffcm9BjM2_2),.clk(gclk));
	jdff dff_B_wrB4E1tO5_2(.din(w_dff_B_ffcm9BjM2_2),.dout(w_dff_B_wrB4E1tO5_2),.clk(gclk));
	jdff dff_B_1fi7Cs1w5_2(.din(w_dff_B_wrB4E1tO5_2),.dout(w_dff_B_1fi7Cs1w5_2),.clk(gclk));
	jdff dff_B_YbbN4NXA2_2(.din(w_dff_B_1fi7Cs1w5_2),.dout(w_dff_B_YbbN4NXA2_2),.clk(gclk));
	jdff dff_B_Blk3KTr49_2(.din(w_dff_B_YbbN4NXA2_2),.dout(w_dff_B_Blk3KTr49_2),.clk(gclk));
	jdff dff_B_6fqCdItL3_2(.din(w_dff_B_Blk3KTr49_2),.dout(w_dff_B_6fqCdItL3_2),.clk(gclk));
	jdff dff_B_GU9LaF1R2_2(.din(w_dff_B_6fqCdItL3_2),.dout(w_dff_B_GU9LaF1R2_2),.clk(gclk));
	jdff dff_B_NHWP0S507_2(.din(n1515),.dout(w_dff_B_NHWP0S507_2),.clk(gclk));
	jdff dff_B_ldo93EOQ0_1(.din(n1513),.dout(w_dff_B_ldo93EOQ0_1),.clk(gclk));
	jdff dff_B_NxUqrVXg7_2(.din(n1441),.dout(w_dff_B_NxUqrVXg7_2),.clk(gclk));
	jdff dff_B_lasVMYWE6_2(.din(w_dff_B_NxUqrVXg7_2),.dout(w_dff_B_lasVMYWE6_2),.clk(gclk));
	jdff dff_B_zKdzvaCg6_2(.din(w_dff_B_lasVMYWE6_2),.dout(w_dff_B_zKdzvaCg6_2),.clk(gclk));
	jdff dff_B_MDjZycQv2_2(.din(w_dff_B_zKdzvaCg6_2),.dout(w_dff_B_MDjZycQv2_2),.clk(gclk));
	jdff dff_B_SVJIUgvq7_2(.din(w_dff_B_MDjZycQv2_2),.dout(w_dff_B_SVJIUgvq7_2),.clk(gclk));
	jdff dff_B_zcXRgkLW2_2(.din(w_dff_B_SVJIUgvq7_2),.dout(w_dff_B_zcXRgkLW2_2),.clk(gclk));
	jdff dff_B_rvsuLzbT2_2(.din(w_dff_B_zcXRgkLW2_2),.dout(w_dff_B_rvsuLzbT2_2),.clk(gclk));
	jdff dff_B_ajsdusPr8_2(.din(w_dff_B_rvsuLzbT2_2),.dout(w_dff_B_ajsdusPr8_2),.clk(gclk));
	jdff dff_B_yy9Qd3dZ9_2(.din(w_dff_B_ajsdusPr8_2),.dout(w_dff_B_yy9Qd3dZ9_2),.clk(gclk));
	jdff dff_B_px0OmXg14_2(.din(w_dff_B_yy9Qd3dZ9_2),.dout(w_dff_B_px0OmXg14_2),.clk(gclk));
	jdff dff_B_XR3cI6gg8_2(.din(w_dff_B_px0OmXg14_2),.dout(w_dff_B_XR3cI6gg8_2),.clk(gclk));
	jdff dff_B_ZDFPikBD9_2(.din(w_dff_B_XR3cI6gg8_2),.dout(w_dff_B_ZDFPikBD9_2),.clk(gclk));
	jdff dff_B_qCnLjZR68_2(.din(w_dff_B_ZDFPikBD9_2),.dout(w_dff_B_qCnLjZR68_2),.clk(gclk));
	jdff dff_B_y3mHFv1R1_2(.din(w_dff_B_qCnLjZR68_2),.dout(w_dff_B_y3mHFv1R1_2),.clk(gclk));
	jdff dff_B_LHox4NkO8_2(.din(w_dff_B_y3mHFv1R1_2),.dout(w_dff_B_LHox4NkO8_2),.clk(gclk));
	jdff dff_B_sE9ohvi66_2(.din(w_dff_B_LHox4NkO8_2),.dout(w_dff_B_sE9ohvi66_2),.clk(gclk));
	jdff dff_B_kxkQrPRe2_2(.din(w_dff_B_sE9ohvi66_2),.dout(w_dff_B_kxkQrPRe2_2),.clk(gclk));
	jdff dff_B_Og0ANBxg0_2(.din(w_dff_B_kxkQrPRe2_2),.dout(w_dff_B_Og0ANBxg0_2),.clk(gclk));
	jdff dff_B_9cSl21ZY9_2(.din(w_dff_B_Og0ANBxg0_2),.dout(w_dff_B_9cSl21ZY9_2),.clk(gclk));
	jdff dff_B_shtL7e940_2(.din(w_dff_B_9cSl21ZY9_2),.dout(w_dff_B_shtL7e940_2),.clk(gclk));
	jdff dff_B_k2uK6uLj3_2(.din(w_dff_B_shtL7e940_2),.dout(w_dff_B_k2uK6uLj3_2),.clk(gclk));
	jdff dff_B_Gg2xaO4H1_2(.din(w_dff_B_k2uK6uLj3_2),.dout(w_dff_B_Gg2xaO4H1_2),.clk(gclk));
	jdff dff_B_nAWGNiAQ1_2(.din(w_dff_B_Gg2xaO4H1_2),.dout(w_dff_B_nAWGNiAQ1_2),.clk(gclk));
	jdff dff_B_x0g9VDz81_2(.din(w_dff_B_nAWGNiAQ1_2),.dout(w_dff_B_x0g9VDz81_2),.clk(gclk));
	jdff dff_B_GmaskMIx0_2(.din(w_dff_B_x0g9VDz81_2),.dout(w_dff_B_GmaskMIx0_2),.clk(gclk));
	jdff dff_B_p0mF0xOr6_2(.din(w_dff_B_GmaskMIx0_2),.dout(w_dff_B_p0mF0xOr6_2),.clk(gclk));
	jdff dff_B_Npw3mhl04_2(.din(w_dff_B_p0mF0xOr6_2),.dout(w_dff_B_Npw3mhl04_2),.clk(gclk));
	jdff dff_B_BGR6rjw04_2(.din(n1444),.dout(w_dff_B_BGR6rjw04_2),.clk(gclk));
	jdff dff_B_pHEnIkim6_1(.din(n1442),.dout(w_dff_B_pHEnIkim6_1),.clk(gclk));
	jdff dff_B_Vy8FtmPu6_2(.din(n1363),.dout(w_dff_B_Vy8FtmPu6_2),.clk(gclk));
	jdff dff_B_jQTDYqi07_2(.din(w_dff_B_Vy8FtmPu6_2),.dout(w_dff_B_jQTDYqi07_2),.clk(gclk));
	jdff dff_B_kqEpPQvl2_2(.din(w_dff_B_jQTDYqi07_2),.dout(w_dff_B_kqEpPQvl2_2),.clk(gclk));
	jdff dff_B_XIVADeVV0_2(.din(w_dff_B_kqEpPQvl2_2),.dout(w_dff_B_XIVADeVV0_2),.clk(gclk));
	jdff dff_B_qQgOhVCK9_2(.din(w_dff_B_XIVADeVV0_2),.dout(w_dff_B_qQgOhVCK9_2),.clk(gclk));
	jdff dff_B_zO9pOINM7_2(.din(w_dff_B_qQgOhVCK9_2),.dout(w_dff_B_zO9pOINM7_2),.clk(gclk));
	jdff dff_B_mZCpK91W5_2(.din(w_dff_B_zO9pOINM7_2),.dout(w_dff_B_mZCpK91W5_2),.clk(gclk));
	jdff dff_B_mbg4fGvC2_2(.din(w_dff_B_mZCpK91W5_2),.dout(w_dff_B_mbg4fGvC2_2),.clk(gclk));
	jdff dff_B_Wyr8CSu17_2(.din(w_dff_B_mbg4fGvC2_2),.dout(w_dff_B_Wyr8CSu17_2),.clk(gclk));
	jdff dff_B_6lo0pbBF7_2(.din(w_dff_B_Wyr8CSu17_2),.dout(w_dff_B_6lo0pbBF7_2),.clk(gclk));
	jdff dff_B_F7dR9jbP4_2(.din(w_dff_B_6lo0pbBF7_2),.dout(w_dff_B_F7dR9jbP4_2),.clk(gclk));
	jdff dff_B_6VGobh8y4_2(.din(w_dff_B_F7dR9jbP4_2),.dout(w_dff_B_6VGobh8y4_2),.clk(gclk));
	jdff dff_B_EPNlYuey3_2(.din(w_dff_B_6VGobh8y4_2),.dout(w_dff_B_EPNlYuey3_2),.clk(gclk));
	jdff dff_B_5mPfdGQY9_2(.din(w_dff_B_EPNlYuey3_2),.dout(w_dff_B_5mPfdGQY9_2),.clk(gclk));
	jdff dff_B_ApfSoGVI9_2(.din(w_dff_B_5mPfdGQY9_2),.dout(w_dff_B_ApfSoGVI9_2),.clk(gclk));
	jdff dff_B_yi03JjiU0_2(.din(w_dff_B_ApfSoGVI9_2),.dout(w_dff_B_yi03JjiU0_2),.clk(gclk));
	jdff dff_B_UBLS2bwR1_2(.din(w_dff_B_yi03JjiU0_2),.dout(w_dff_B_UBLS2bwR1_2),.clk(gclk));
	jdff dff_B_3unU2PrT8_2(.din(w_dff_B_UBLS2bwR1_2),.dout(w_dff_B_3unU2PrT8_2),.clk(gclk));
	jdff dff_B_UuLPRUt52_2(.din(w_dff_B_3unU2PrT8_2),.dout(w_dff_B_UuLPRUt52_2),.clk(gclk));
	jdff dff_B_chwKB6sU9_2(.din(w_dff_B_UuLPRUt52_2),.dout(w_dff_B_chwKB6sU9_2),.clk(gclk));
	jdff dff_B_ec3W0gK28_2(.din(w_dff_B_chwKB6sU9_2),.dout(w_dff_B_ec3W0gK28_2),.clk(gclk));
	jdff dff_B_g0zwmJyW6_2(.din(w_dff_B_ec3W0gK28_2),.dout(w_dff_B_g0zwmJyW6_2),.clk(gclk));
	jdff dff_B_4YywosL63_2(.din(w_dff_B_g0zwmJyW6_2),.dout(w_dff_B_4YywosL63_2),.clk(gclk));
	jdff dff_B_HexU8YbC7_2(.din(w_dff_B_4YywosL63_2),.dout(w_dff_B_HexU8YbC7_2),.clk(gclk));
	jdff dff_B_iWMEV3TI9_2(.din(n1366),.dout(w_dff_B_iWMEV3TI9_2),.clk(gclk));
	jdff dff_B_HcTs0byL2_1(.din(n1364),.dout(w_dff_B_HcTs0byL2_1),.clk(gclk));
	jdff dff_B_6PVzsnq21_2(.din(n1278),.dout(w_dff_B_6PVzsnq21_2),.clk(gclk));
	jdff dff_B_psVN11xF7_2(.din(w_dff_B_6PVzsnq21_2),.dout(w_dff_B_psVN11xF7_2),.clk(gclk));
	jdff dff_B_VNxKUYAG3_2(.din(w_dff_B_psVN11xF7_2),.dout(w_dff_B_VNxKUYAG3_2),.clk(gclk));
	jdff dff_B_8Zk1SmxN3_2(.din(w_dff_B_VNxKUYAG3_2),.dout(w_dff_B_8Zk1SmxN3_2),.clk(gclk));
	jdff dff_B_RMUaedLb5_2(.din(w_dff_B_8Zk1SmxN3_2),.dout(w_dff_B_RMUaedLb5_2),.clk(gclk));
	jdff dff_B_5ekJN1di7_2(.din(w_dff_B_RMUaedLb5_2),.dout(w_dff_B_5ekJN1di7_2),.clk(gclk));
	jdff dff_B_Stw6vIAy9_2(.din(w_dff_B_5ekJN1di7_2),.dout(w_dff_B_Stw6vIAy9_2),.clk(gclk));
	jdff dff_B_eyXZtImS5_2(.din(w_dff_B_Stw6vIAy9_2),.dout(w_dff_B_eyXZtImS5_2),.clk(gclk));
	jdff dff_B_eMyVEqZ17_2(.din(w_dff_B_eyXZtImS5_2),.dout(w_dff_B_eMyVEqZ17_2),.clk(gclk));
	jdff dff_B_HEd30MXq6_2(.din(w_dff_B_eMyVEqZ17_2),.dout(w_dff_B_HEd30MXq6_2),.clk(gclk));
	jdff dff_B_V4XjnTm12_2(.din(w_dff_B_HEd30MXq6_2),.dout(w_dff_B_V4XjnTm12_2),.clk(gclk));
	jdff dff_B_VDGvfSHX1_2(.din(w_dff_B_V4XjnTm12_2),.dout(w_dff_B_VDGvfSHX1_2),.clk(gclk));
	jdff dff_B_sH9PoYqz0_2(.din(w_dff_B_VDGvfSHX1_2),.dout(w_dff_B_sH9PoYqz0_2),.clk(gclk));
	jdff dff_B_cj7s6ouI1_2(.din(w_dff_B_sH9PoYqz0_2),.dout(w_dff_B_cj7s6ouI1_2),.clk(gclk));
	jdff dff_B_okqjrnQH7_2(.din(w_dff_B_cj7s6ouI1_2),.dout(w_dff_B_okqjrnQH7_2),.clk(gclk));
	jdff dff_B_q0mawQe65_2(.din(w_dff_B_okqjrnQH7_2),.dout(w_dff_B_q0mawQe65_2),.clk(gclk));
	jdff dff_B_EMIhYefK4_2(.din(w_dff_B_q0mawQe65_2),.dout(w_dff_B_EMIhYefK4_2),.clk(gclk));
	jdff dff_B_Ezs2lTVU5_2(.din(w_dff_B_EMIhYefK4_2),.dout(w_dff_B_Ezs2lTVU5_2),.clk(gclk));
	jdff dff_B_qk7JLf7v5_2(.din(w_dff_B_Ezs2lTVU5_2),.dout(w_dff_B_qk7JLf7v5_2),.clk(gclk));
	jdff dff_B_NZzFJg3M8_2(.din(w_dff_B_qk7JLf7v5_2),.dout(w_dff_B_NZzFJg3M8_2),.clk(gclk));
	jdff dff_B_D87deOIr2_2(.din(w_dff_B_NZzFJg3M8_2),.dout(w_dff_B_D87deOIr2_2),.clk(gclk));
	jdff dff_B_uojRNQmk5_2(.din(n1281),.dout(w_dff_B_uojRNQmk5_2),.clk(gclk));
	jdff dff_B_fGZzhjhB6_1(.din(n1279),.dout(w_dff_B_fGZzhjhB6_1),.clk(gclk));
	jdff dff_B_n17ZVxRT3_2(.din(n1188),.dout(w_dff_B_n17ZVxRT3_2),.clk(gclk));
	jdff dff_B_R9V95fYB0_2(.din(w_dff_B_n17ZVxRT3_2),.dout(w_dff_B_R9V95fYB0_2),.clk(gclk));
	jdff dff_B_APApAvjJ4_2(.din(w_dff_B_R9V95fYB0_2),.dout(w_dff_B_APApAvjJ4_2),.clk(gclk));
	jdff dff_B_W85EUjSY1_2(.din(w_dff_B_APApAvjJ4_2),.dout(w_dff_B_W85EUjSY1_2),.clk(gclk));
	jdff dff_B_7EaeYfsR7_2(.din(w_dff_B_W85EUjSY1_2),.dout(w_dff_B_7EaeYfsR7_2),.clk(gclk));
	jdff dff_B_rJfKmYiA8_2(.din(w_dff_B_7EaeYfsR7_2),.dout(w_dff_B_rJfKmYiA8_2),.clk(gclk));
	jdff dff_B_r1BfFEvS5_2(.din(w_dff_B_rJfKmYiA8_2),.dout(w_dff_B_r1BfFEvS5_2),.clk(gclk));
	jdff dff_B_qe6iiy171_2(.din(w_dff_B_r1BfFEvS5_2),.dout(w_dff_B_qe6iiy171_2),.clk(gclk));
	jdff dff_B_lnwLFdiM6_2(.din(w_dff_B_qe6iiy171_2),.dout(w_dff_B_lnwLFdiM6_2),.clk(gclk));
	jdff dff_B_tiqfHTdP7_2(.din(w_dff_B_lnwLFdiM6_2),.dout(w_dff_B_tiqfHTdP7_2),.clk(gclk));
	jdff dff_B_SaZUhaoZ5_2(.din(w_dff_B_tiqfHTdP7_2),.dout(w_dff_B_SaZUhaoZ5_2),.clk(gclk));
	jdff dff_B_1QzeL0RR4_2(.din(w_dff_B_SaZUhaoZ5_2),.dout(w_dff_B_1QzeL0RR4_2),.clk(gclk));
	jdff dff_B_28BcldFj2_2(.din(w_dff_B_1QzeL0RR4_2),.dout(w_dff_B_28BcldFj2_2),.clk(gclk));
	jdff dff_B_n20NaSMn5_2(.din(w_dff_B_28BcldFj2_2),.dout(w_dff_B_n20NaSMn5_2),.clk(gclk));
	jdff dff_B_SxJkGRgQ8_2(.din(w_dff_B_n20NaSMn5_2),.dout(w_dff_B_SxJkGRgQ8_2),.clk(gclk));
	jdff dff_B_T9meeg3C1_2(.din(w_dff_B_SxJkGRgQ8_2),.dout(w_dff_B_T9meeg3C1_2),.clk(gclk));
	jdff dff_B_9GiUuddW9_2(.din(w_dff_B_T9meeg3C1_2),.dout(w_dff_B_9GiUuddW9_2),.clk(gclk));
	jdff dff_B_EuRzVPuY5_2(.din(w_dff_B_9GiUuddW9_2),.dout(w_dff_B_EuRzVPuY5_2),.clk(gclk));
	jdff dff_B_s1neHrrM3_2(.din(n1191),.dout(w_dff_B_s1neHrrM3_2),.clk(gclk));
	jdff dff_B_dFsHh26v2_1(.din(n1189),.dout(w_dff_B_dFsHh26v2_1),.clk(gclk));
	jdff dff_B_oZIRDm7s4_2(.din(n1084),.dout(w_dff_B_oZIRDm7s4_2),.clk(gclk));
	jdff dff_B_PgxJ4dNf9_2(.din(w_dff_B_oZIRDm7s4_2),.dout(w_dff_B_PgxJ4dNf9_2),.clk(gclk));
	jdff dff_B_MByjT5W80_2(.din(w_dff_B_PgxJ4dNf9_2),.dout(w_dff_B_MByjT5W80_2),.clk(gclk));
	jdff dff_B_3zLb4nV35_2(.din(w_dff_B_MByjT5W80_2),.dout(w_dff_B_3zLb4nV35_2),.clk(gclk));
	jdff dff_B_MnFLoEPa1_2(.din(w_dff_B_3zLb4nV35_2),.dout(w_dff_B_MnFLoEPa1_2),.clk(gclk));
	jdff dff_B_6xbD8Xho5_2(.din(w_dff_B_MnFLoEPa1_2),.dout(w_dff_B_6xbD8Xho5_2),.clk(gclk));
	jdff dff_B_paexazBJ7_2(.din(w_dff_B_6xbD8Xho5_2),.dout(w_dff_B_paexazBJ7_2),.clk(gclk));
	jdff dff_B_D3uaoPtH8_2(.din(w_dff_B_paexazBJ7_2),.dout(w_dff_B_D3uaoPtH8_2),.clk(gclk));
	jdff dff_B_v9D0bK746_2(.din(w_dff_B_D3uaoPtH8_2),.dout(w_dff_B_v9D0bK746_2),.clk(gclk));
	jdff dff_B_FQrQ3fBc5_2(.din(w_dff_B_v9D0bK746_2),.dout(w_dff_B_FQrQ3fBc5_2),.clk(gclk));
	jdff dff_B_fApgYZmH1_2(.din(w_dff_B_FQrQ3fBc5_2),.dout(w_dff_B_fApgYZmH1_2),.clk(gclk));
	jdff dff_B_PdRg3K7r0_2(.din(w_dff_B_fApgYZmH1_2),.dout(w_dff_B_PdRg3K7r0_2),.clk(gclk));
	jdff dff_B_vJ4Ybcxj4_2(.din(w_dff_B_PdRg3K7r0_2),.dout(w_dff_B_vJ4Ybcxj4_2),.clk(gclk));
	jdff dff_B_AIb5Liqz6_2(.din(w_dff_B_vJ4Ybcxj4_2),.dout(w_dff_B_AIb5Liqz6_2),.clk(gclk));
	jdff dff_B_y3BcU3Is6_2(.din(w_dff_B_AIb5Liqz6_2),.dout(w_dff_B_y3BcU3Is6_2),.clk(gclk));
	jdff dff_B_575PgbKq3_2(.din(n1087),.dout(w_dff_B_575PgbKq3_2),.clk(gclk));
	jdff dff_B_14tFs7Lf3_1(.din(n1085),.dout(w_dff_B_14tFs7Lf3_1),.clk(gclk));
	jdff dff_B_XTDYzMiw6_2(.din(n986),.dout(w_dff_B_XTDYzMiw6_2),.clk(gclk));
	jdff dff_B_u0ycFSqx9_2(.din(w_dff_B_XTDYzMiw6_2),.dout(w_dff_B_u0ycFSqx9_2),.clk(gclk));
	jdff dff_B_SyVbmMo31_2(.din(w_dff_B_u0ycFSqx9_2),.dout(w_dff_B_SyVbmMo31_2),.clk(gclk));
	jdff dff_B_HmnsD02t1_2(.din(w_dff_B_SyVbmMo31_2),.dout(w_dff_B_HmnsD02t1_2),.clk(gclk));
	jdff dff_B_CrQh6mNC3_2(.din(w_dff_B_HmnsD02t1_2),.dout(w_dff_B_CrQh6mNC3_2),.clk(gclk));
	jdff dff_B_hGdeg0wU5_2(.din(w_dff_B_CrQh6mNC3_2),.dout(w_dff_B_hGdeg0wU5_2),.clk(gclk));
	jdff dff_B_FbOgMmUl2_2(.din(w_dff_B_hGdeg0wU5_2),.dout(w_dff_B_FbOgMmUl2_2),.clk(gclk));
	jdff dff_B_q1g83Cs38_2(.din(w_dff_B_FbOgMmUl2_2),.dout(w_dff_B_q1g83Cs38_2),.clk(gclk));
	jdff dff_B_J9m7R1mc3_2(.din(w_dff_B_q1g83Cs38_2),.dout(w_dff_B_J9m7R1mc3_2),.clk(gclk));
	jdff dff_B_nd2iupUz6_2(.din(w_dff_B_J9m7R1mc3_2),.dout(w_dff_B_nd2iupUz6_2),.clk(gclk));
	jdff dff_B_I7LmuTso3_2(.din(w_dff_B_nd2iupUz6_2),.dout(w_dff_B_I7LmuTso3_2),.clk(gclk));
	jdff dff_B_6akHVQl14_2(.din(w_dff_B_I7LmuTso3_2),.dout(w_dff_B_6akHVQl14_2),.clk(gclk));
	jdff dff_B_T8q6GaV73_1(.din(n987),.dout(w_dff_B_T8q6GaV73_1),.clk(gclk));
	jdff dff_B_ivK1VAAe2_2(.din(n881),.dout(w_dff_B_ivK1VAAe2_2),.clk(gclk));
	jdff dff_B_GLbQrpUB7_2(.din(w_dff_B_ivK1VAAe2_2),.dout(w_dff_B_GLbQrpUB7_2),.clk(gclk));
	jdff dff_B_xuHbWMUq0_2(.din(w_dff_B_GLbQrpUB7_2),.dout(w_dff_B_xuHbWMUq0_2),.clk(gclk));
	jdff dff_B_TMsJyuR51_2(.din(w_dff_B_xuHbWMUq0_2),.dout(w_dff_B_TMsJyuR51_2),.clk(gclk));
	jdff dff_B_s0PbNZX80_2(.din(w_dff_B_TMsJyuR51_2),.dout(w_dff_B_s0PbNZX80_2),.clk(gclk));
	jdff dff_B_8Vj2Ag9v6_2(.din(w_dff_B_s0PbNZX80_2),.dout(w_dff_B_8Vj2Ag9v6_2),.clk(gclk));
	jdff dff_B_iOK7Jftm4_2(.din(w_dff_B_8Vj2Ag9v6_2),.dout(w_dff_B_iOK7Jftm4_2),.clk(gclk));
	jdff dff_B_d7oiqQTm5_2(.din(w_dff_B_iOK7Jftm4_2),.dout(w_dff_B_d7oiqQTm5_2),.clk(gclk));
	jdff dff_B_tTqFB1lD5_2(.din(w_dff_B_d7oiqQTm5_2),.dout(w_dff_B_tTqFB1lD5_2),.clk(gclk));
	jdff dff_B_6PAKBTgy5_2(.din(w_dff_B_tTqFB1lD5_2),.dout(w_dff_B_6PAKBTgy5_2),.clk(gclk));
	jdff dff_B_39ySnxDb3_1(.din(n882),.dout(w_dff_B_39ySnxDb3_1),.clk(gclk));
	jdff dff_B_OSuTQmLa3_2(.din(n782),.dout(w_dff_B_OSuTQmLa3_2),.clk(gclk));
	jdff dff_B_cWuLtvFd8_2(.din(w_dff_B_OSuTQmLa3_2),.dout(w_dff_B_cWuLtvFd8_2),.clk(gclk));
	jdff dff_B_p7ityrFI8_2(.din(w_dff_B_cWuLtvFd8_2),.dout(w_dff_B_p7ityrFI8_2),.clk(gclk));
	jdff dff_B_RX3HDQs35_2(.din(w_dff_B_p7ityrFI8_2),.dout(w_dff_B_RX3HDQs35_2),.clk(gclk));
	jdff dff_B_hlA5x6yI2_2(.din(w_dff_B_RX3HDQs35_2),.dout(w_dff_B_hlA5x6yI2_2),.clk(gclk));
	jdff dff_B_DL3pBouH4_2(.din(w_dff_B_hlA5x6yI2_2),.dout(w_dff_B_DL3pBouH4_2),.clk(gclk));
	jdff dff_B_T1ih5VfZ8_2(.din(w_dff_B_DL3pBouH4_2),.dout(w_dff_B_T1ih5VfZ8_2),.clk(gclk));
	jdff dff_B_IYyZof909_2(.din(w_dff_B_T1ih5VfZ8_2),.dout(w_dff_B_IYyZof909_2),.clk(gclk));
	jdff dff_B_m2N89aZe5_1(.din(n783),.dout(w_dff_B_m2N89aZe5_1),.clk(gclk));
	jdff dff_B_9NibFXlu7_2(.din(n689),.dout(w_dff_B_9NibFXlu7_2),.clk(gclk));
	jdff dff_B_i5awPHmD6_2(.din(w_dff_B_9NibFXlu7_2),.dout(w_dff_B_i5awPHmD6_2),.clk(gclk));
	jdff dff_B_qUTHNux54_2(.din(w_dff_B_i5awPHmD6_2),.dout(w_dff_B_qUTHNux54_2),.clk(gclk));
	jdff dff_B_3Qm1Dhu44_2(.din(w_dff_B_qUTHNux54_2),.dout(w_dff_B_3Qm1Dhu44_2),.clk(gclk));
	jdff dff_B_oLzjGmyc2_2(.din(w_dff_B_3Qm1Dhu44_2),.dout(w_dff_B_oLzjGmyc2_2),.clk(gclk));
	jdff dff_B_SzG0N2Y24_2(.din(w_dff_B_oLzjGmyc2_2),.dout(w_dff_B_SzG0N2Y24_2),.clk(gclk));
	jdff dff_B_wlQBLVKH0_2(.din(n705),.dout(w_dff_B_wlQBLVKH0_2),.clk(gclk));
	jdff dff_B_UipQ2Ew40_1(.din(n690),.dout(w_dff_B_UipQ2Ew40_1),.clk(gclk));
	jdff dff_B_W6KneUft4_1(.din(w_dff_B_UipQ2Ew40_1),.dout(w_dff_B_W6KneUft4_1),.clk(gclk));
	jdff dff_B_0mD8oNg82_1(.din(w_dff_B_W6KneUft4_1),.dout(w_dff_B_0mD8oNg82_1),.clk(gclk));
	jdff dff_B_TCFaCcQC4_1(.din(w_dff_B_0mD8oNg82_1),.dout(w_dff_B_TCFaCcQC4_1),.clk(gclk));
	jdff dff_B_Gdn853Jj8_0(.din(n612),.dout(w_dff_B_Gdn853Jj8_0),.clk(gclk));
	jdff dff_A_fWPG9oRP9_0(.dout(w_n611_0[0]),.din(w_dff_A_fWPG9oRP9_0),.clk(gclk));
	jdff dff_A_LStzzifJ6_0(.dout(w_dff_A_fWPG9oRP9_0),.din(w_dff_A_LStzzifJ6_0),.clk(gclk));
	jdff dff_B_VQ1qjIrd5_1(.din(n605),.dout(w_dff_B_VQ1qjIrd5_1),.clk(gclk));
	jdff dff_B_VBFHxlXZ9_1(.din(w_dff_B_VQ1qjIrd5_1),.dout(w_dff_B_VBFHxlXZ9_1),.clk(gclk));
	jdff dff_A_jLjA2Bfy3_0(.dout(w_n523_0[0]),.din(w_dff_A_jLjA2Bfy3_0),.clk(gclk));
	jdff dff_A_UZaFVqwY3_1(.dout(w_n523_0[1]),.din(w_dff_A_UZaFVqwY3_1),.clk(gclk));
	jdff dff_A_drno1gMW4_1(.dout(w_dff_A_UZaFVqwY3_1),.din(w_dff_A_drno1gMW4_1),.clk(gclk));
	jdff dff_A_cJO0RiS59_1(.dout(w_n603_0[1]),.din(w_dff_A_cJO0RiS59_1),.clk(gclk));
	jdff dff_A_HUDkCOMd1_1(.dout(w_dff_A_cJO0RiS59_1),.din(w_dff_A_HUDkCOMd1_1),.clk(gclk));
	jdff dff_A_pJYFsnAs3_1(.dout(w_dff_A_HUDkCOMd1_1),.din(w_dff_A_pJYFsnAs3_1),.clk(gclk));
	jdff dff_A_G8IX5VBQ3_1(.dout(w_dff_A_pJYFsnAs3_1),.din(w_dff_A_G8IX5VBQ3_1),.clk(gclk));
	jdff dff_B_qnSP67mV0_1(.din(n1793),.dout(w_dff_B_qnSP67mV0_1),.clk(gclk));
	jdff dff_A_FthOBBaS1_1(.dout(w_n1768_0[1]),.din(w_dff_A_FthOBBaS1_1),.clk(gclk));
	jdff dff_B_6DV67CBU5_1(.din(n1766),.dout(w_dff_B_6DV67CBU5_1),.clk(gclk));
	jdff dff_B_dOGg3N0J9_2(.din(n1730),.dout(w_dff_B_dOGg3N0J9_2),.clk(gclk));
	jdff dff_B_1BmlShjP1_2(.din(w_dff_B_dOGg3N0J9_2),.dout(w_dff_B_1BmlShjP1_2),.clk(gclk));
	jdff dff_B_sBCdCDWn5_2(.din(w_dff_B_1BmlShjP1_2),.dout(w_dff_B_sBCdCDWn5_2),.clk(gclk));
	jdff dff_B_6kVV8mKa3_2(.din(w_dff_B_sBCdCDWn5_2),.dout(w_dff_B_6kVV8mKa3_2),.clk(gclk));
	jdff dff_B_JagPo3q85_2(.din(w_dff_B_6kVV8mKa3_2),.dout(w_dff_B_JagPo3q85_2),.clk(gclk));
	jdff dff_B_QKmtHe0w6_2(.din(w_dff_B_JagPo3q85_2),.dout(w_dff_B_QKmtHe0w6_2),.clk(gclk));
	jdff dff_B_qnmEbv951_2(.din(w_dff_B_QKmtHe0w6_2),.dout(w_dff_B_qnmEbv951_2),.clk(gclk));
	jdff dff_B_VLBTxCBx4_2(.din(w_dff_B_qnmEbv951_2),.dout(w_dff_B_VLBTxCBx4_2),.clk(gclk));
	jdff dff_B_4hF8vQex5_2(.din(w_dff_B_VLBTxCBx4_2),.dout(w_dff_B_4hF8vQex5_2),.clk(gclk));
	jdff dff_B_0wamdWPN2_2(.din(w_dff_B_4hF8vQex5_2),.dout(w_dff_B_0wamdWPN2_2),.clk(gclk));
	jdff dff_B_zGbEiIo27_2(.din(w_dff_B_0wamdWPN2_2),.dout(w_dff_B_zGbEiIo27_2),.clk(gclk));
	jdff dff_B_SJlWIMlT8_2(.din(w_dff_B_zGbEiIo27_2),.dout(w_dff_B_SJlWIMlT8_2),.clk(gclk));
	jdff dff_B_ro1LDj600_2(.din(w_dff_B_SJlWIMlT8_2),.dout(w_dff_B_ro1LDj600_2),.clk(gclk));
	jdff dff_B_xn7xKFE13_2(.din(w_dff_B_ro1LDj600_2),.dout(w_dff_B_xn7xKFE13_2),.clk(gclk));
	jdff dff_B_mSMf1meb0_2(.din(w_dff_B_xn7xKFE13_2),.dout(w_dff_B_mSMf1meb0_2),.clk(gclk));
	jdff dff_B_yLahuzfi4_2(.din(w_dff_B_mSMf1meb0_2),.dout(w_dff_B_yLahuzfi4_2),.clk(gclk));
	jdff dff_B_NItNMQwT1_2(.din(w_dff_B_yLahuzfi4_2),.dout(w_dff_B_NItNMQwT1_2),.clk(gclk));
	jdff dff_B_rNiRcqA04_2(.din(w_dff_B_NItNMQwT1_2),.dout(w_dff_B_rNiRcqA04_2),.clk(gclk));
	jdff dff_B_V0mWvfAB1_2(.din(w_dff_B_rNiRcqA04_2),.dout(w_dff_B_V0mWvfAB1_2),.clk(gclk));
	jdff dff_B_e309RbpT0_2(.din(w_dff_B_V0mWvfAB1_2),.dout(w_dff_B_e309RbpT0_2),.clk(gclk));
	jdff dff_B_ZaQrucqD1_2(.din(w_dff_B_e309RbpT0_2),.dout(w_dff_B_ZaQrucqD1_2),.clk(gclk));
	jdff dff_B_Isvci4dc6_2(.din(w_dff_B_ZaQrucqD1_2),.dout(w_dff_B_Isvci4dc6_2),.clk(gclk));
	jdff dff_B_PKbRrpm65_2(.din(w_dff_B_Isvci4dc6_2),.dout(w_dff_B_PKbRrpm65_2),.clk(gclk));
	jdff dff_B_fR9qGCHX3_2(.din(w_dff_B_PKbRrpm65_2),.dout(w_dff_B_fR9qGCHX3_2),.clk(gclk));
	jdff dff_B_QmG4y5At7_2(.din(w_dff_B_fR9qGCHX3_2),.dout(w_dff_B_QmG4y5At7_2),.clk(gclk));
	jdff dff_B_sGJlLfS49_2(.din(w_dff_B_QmG4y5At7_2),.dout(w_dff_B_sGJlLfS49_2),.clk(gclk));
	jdff dff_B_EUdTtewU4_2(.din(w_dff_B_sGJlLfS49_2),.dout(w_dff_B_EUdTtewU4_2),.clk(gclk));
	jdff dff_B_LCmBFyil5_2(.din(w_dff_B_EUdTtewU4_2),.dout(w_dff_B_LCmBFyil5_2),.clk(gclk));
	jdff dff_B_l3P6T8yE3_2(.din(w_dff_B_LCmBFyil5_2),.dout(w_dff_B_l3P6T8yE3_2),.clk(gclk));
	jdff dff_B_Jp49Wk0u2_2(.din(w_dff_B_l3P6T8yE3_2),.dout(w_dff_B_Jp49Wk0u2_2),.clk(gclk));
	jdff dff_B_RaOkfKwl2_2(.din(w_dff_B_Jp49Wk0u2_2),.dout(w_dff_B_RaOkfKwl2_2),.clk(gclk));
	jdff dff_B_4fikkssd9_2(.din(w_dff_B_RaOkfKwl2_2),.dout(w_dff_B_4fikkssd9_2),.clk(gclk));
	jdff dff_B_lRKQxxSF5_2(.din(w_dff_B_4fikkssd9_2),.dout(w_dff_B_lRKQxxSF5_2),.clk(gclk));
	jdff dff_B_I2v5cY621_2(.din(w_dff_B_lRKQxxSF5_2),.dout(w_dff_B_I2v5cY621_2),.clk(gclk));
	jdff dff_B_pTGnd6c54_2(.din(w_dff_B_I2v5cY621_2),.dout(w_dff_B_pTGnd6c54_2),.clk(gclk));
	jdff dff_B_TZr5F3Og9_2(.din(w_dff_B_pTGnd6c54_2),.dout(w_dff_B_TZr5F3Og9_2),.clk(gclk));
	jdff dff_B_kR4OS3qD2_2(.din(w_dff_B_TZr5F3Og9_2),.dout(w_dff_B_kR4OS3qD2_2),.clk(gclk));
	jdff dff_B_EdX3cqby4_2(.din(w_dff_B_kR4OS3qD2_2),.dout(w_dff_B_EdX3cqby4_2),.clk(gclk));
	jdff dff_B_MJBz7X6l3_2(.din(w_dff_B_EdX3cqby4_2),.dout(w_dff_B_MJBz7X6l3_2),.clk(gclk));
	jdff dff_B_b5xB4cfa7_2(.din(w_dff_B_MJBz7X6l3_2),.dout(w_dff_B_b5xB4cfa7_2),.clk(gclk));
	jdff dff_B_sWLejboO0_2(.din(n1733),.dout(w_dff_B_sWLejboO0_2),.clk(gclk));
	jdff dff_B_2il5fWCi4_1(.din(n1731),.dout(w_dff_B_2il5fWCi4_1),.clk(gclk));
	jdff dff_B_2OzbK2XA6_2(.din(n1689),.dout(w_dff_B_2OzbK2XA6_2),.clk(gclk));
	jdff dff_B_EoCiPKBW8_2(.din(w_dff_B_2OzbK2XA6_2),.dout(w_dff_B_EoCiPKBW8_2),.clk(gclk));
	jdff dff_B_LwlA3ID82_2(.din(w_dff_B_EoCiPKBW8_2),.dout(w_dff_B_LwlA3ID82_2),.clk(gclk));
	jdff dff_B_VMTBGKw68_2(.din(w_dff_B_LwlA3ID82_2),.dout(w_dff_B_VMTBGKw68_2),.clk(gclk));
	jdff dff_B_7hAYZ7a72_2(.din(w_dff_B_VMTBGKw68_2),.dout(w_dff_B_7hAYZ7a72_2),.clk(gclk));
	jdff dff_B_xAbScloS1_2(.din(w_dff_B_7hAYZ7a72_2),.dout(w_dff_B_xAbScloS1_2),.clk(gclk));
	jdff dff_B_zgGxRnWB1_2(.din(w_dff_B_xAbScloS1_2),.dout(w_dff_B_zgGxRnWB1_2),.clk(gclk));
	jdff dff_B_Hf8Cv6NT2_2(.din(w_dff_B_zgGxRnWB1_2),.dout(w_dff_B_Hf8Cv6NT2_2),.clk(gclk));
	jdff dff_B_8mLDssmW5_2(.din(w_dff_B_Hf8Cv6NT2_2),.dout(w_dff_B_8mLDssmW5_2),.clk(gclk));
	jdff dff_B_VbtoKRMe7_2(.din(w_dff_B_8mLDssmW5_2),.dout(w_dff_B_VbtoKRMe7_2),.clk(gclk));
	jdff dff_B_vKNmCYuV2_2(.din(w_dff_B_VbtoKRMe7_2),.dout(w_dff_B_vKNmCYuV2_2),.clk(gclk));
	jdff dff_B_rJTmePHG6_2(.din(w_dff_B_vKNmCYuV2_2),.dout(w_dff_B_rJTmePHG6_2),.clk(gclk));
	jdff dff_B_CEIZkxE79_2(.din(w_dff_B_rJTmePHG6_2),.dout(w_dff_B_CEIZkxE79_2),.clk(gclk));
	jdff dff_B_AHprEfiw6_2(.din(w_dff_B_CEIZkxE79_2),.dout(w_dff_B_AHprEfiw6_2),.clk(gclk));
	jdff dff_B_5gvjk9xL3_2(.din(w_dff_B_AHprEfiw6_2),.dout(w_dff_B_5gvjk9xL3_2),.clk(gclk));
	jdff dff_B_1NRycjdP0_2(.din(w_dff_B_5gvjk9xL3_2),.dout(w_dff_B_1NRycjdP0_2),.clk(gclk));
	jdff dff_B_x27BvJEP3_2(.din(w_dff_B_1NRycjdP0_2),.dout(w_dff_B_x27BvJEP3_2),.clk(gclk));
	jdff dff_B_ZYVl3Eh15_2(.din(w_dff_B_x27BvJEP3_2),.dout(w_dff_B_ZYVl3Eh15_2),.clk(gclk));
	jdff dff_B_1yn8CzxY3_2(.din(w_dff_B_ZYVl3Eh15_2),.dout(w_dff_B_1yn8CzxY3_2),.clk(gclk));
	jdff dff_B_oyhNrCuN2_2(.din(w_dff_B_1yn8CzxY3_2),.dout(w_dff_B_oyhNrCuN2_2),.clk(gclk));
	jdff dff_B_MLqOKC2B5_2(.din(w_dff_B_oyhNrCuN2_2),.dout(w_dff_B_MLqOKC2B5_2),.clk(gclk));
	jdff dff_B_ELCuy6ku5_2(.din(w_dff_B_MLqOKC2B5_2),.dout(w_dff_B_ELCuy6ku5_2),.clk(gclk));
	jdff dff_B_t1mhuLBV3_2(.din(w_dff_B_ELCuy6ku5_2),.dout(w_dff_B_t1mhuLBV3_2),.clk(gclk));
	jdff dff_B_JsgnFewA9_2(.din(w_dff_B_t1mhuLBV3_2),.dout(w_dff_B_JsgnFewA9_2),.clk(gclk));
	jdff dff_B_nqK2qD8L1_2(.din(w_dff_B_JsgnFewA9_2),.dout(w_dff_B_nqK2qD8L1_2),.clk(gclk));
	jdff dff_B_9QxNETOY0_2(.din(w_dff_B_nqK2qD8L1_2),.dout(w_dff_B_9QxNETOY0_2),.clk(gclk));
	jdff dff_B_HTZrj48d7_2(.din(w_dff_B_9QxNETOY0_2),.dout(w_dff_B_HTZrj48d7_2),.clk(gclk));
	jdff dff_B_8Db2viEg0_2(.din(w_dff_B_HTZrj48d7_2),.dout(w_dff_B_8Db2viEg0_2),.clk(gclk));
	jdff dff_B_vQSEPpxU1_2(.din(w_dff_B_8Db2viEg0_2),.dout(w_dff_B_vQSEPpxU1_2),.clk(gclk));
	jdff dff_B_RHToYluM0_2(.din(w_dff_B_vQSEPpxU1_2),.dout(w_dff_B_RHToYluM0_2),.clk(gclk));
	jdff dff_B_e3zctTOZ1_2(.din(w_dff_B_RHToYluM0_2),.dout(w_dff_B_e3zctTOZ1_2),.clk(gclk));
	jdff dff_B_NObX8p2T4_2(.din(w_dff_B_e3zctTOZ1_2),.dout(w_dff_B_NObX8p2T4_2),.clk(gclk));
	jdff dff_B_fnwMtLeA2_2(.din(w_dff_B_NObX8p2T4_2),.dout(w_dff_B_fnwMtLeA2_2),.clk(gclk));
	jdff dff_B_9YwLMyqe9_2(.din(w_dff_B_fnwMtLeA2_2),.dout(w_dff_B_9YwLMyqe9_2),.clk(gclk));
	jdff dff_B_rFYf5rFh4_2(.din(w_dff_B_9YwLMyqe9_2),.dout(w_dff_B_rFYf5rFh4_2),.clk(gclk));
	jdff dff_B_cL5T4Ogy2_2(.din(w_dff_B_rFYf5rFh4_2),.dout(w_dff_B_cL5T4Ogy2_2),.clk(gclk));
	jdff dff_B_3X9ysqiv8_2(.din(w_dff_B_cL5T4Ogy2_2),.dout(w_dff_B_3X9ysqiv8_2),.clk(gclk));
	jdff dff_B_hmSzzKIG2_2(.din(n1692),.dout(w_dff_B_hmSzzKIG2_2),.clk(gclk));
	jdff dff_B_xMcZA4CE3_1(.din(n1690),.dout(w_dff_B_xMcZA4CE3_1),.clk(gclk));
	jdff dff_B_mf5Ueczm1_2(.din(n1638),.dout(w_dff_B_mf5Ueczm1_2),.clk(gclk));
	jdff dff_B_GOvvzfQK0_2(.din(w_dff_B_mf5Ueczm1_2),.dout(w_dff_B_GOvvzfQK0_2),.clk(gclk));
	jdff dff_B_d4VJ3tOM3_2(.din(w_dff_B_GOvvzfQK0_2),.dout(w_dff_B_d4VJ3tOM3_2),.clk(gclk));
	jdff dff_B_E3VU0BC40_2(.din(w_dff_B_d4VJ3tOM3_2),.dout(w_dff_B_E3VU0BC40_2),.clk(gclk));
	jdff dff_B_whJIcojK4_2(.din(w_dff_B_E3VU0BC40_2),.dout(w_dff_B_whJIcojK4_2),.clk(gclk));
	jdff dff_B_jABkM8HR5_2(.din(w_dff_B_whJIcojK4_2),.dout(w_dff_B_jABkM8HR5_2),.clk(gclk));
	jdff dff_B_nuBBTAud4_2(.din(w_dff_B_jABkM8HR5_2),.dout(w_dff_B_nuBBTAud4_2),.clk(gclk));
	jdff dff_B_SlEPmMjx0_2(.din(w_dff_B_nuBBTAud4_2),.dout(w_dff_B_SlEPmMjx0_2),.clk(gclk));
	jdff dff_B_GjPHJlsT0_2(.din(w_dff_B_SlEPmMjx0_2),.dout(w_dff_B_GjPHJlsT0_2),.clk(gclk));
	jdff dff_B_kGrvL8tl5_2(.din(w_dff_B_GjPHJlsT0_2),.dout(w_dff_B_kGrvL8tl5_2),.clk(gclk));
	jdff dff_B_J9I9zmIs3_2(.din(w_dff_B_kGrvL8tl5_2),.dout(w_dff_B_J9I9zmIs3_2),.clk(gclk));
	jdff dff_B_Z8pmxG6x4_2(.din(w_dff_B_J9I9zmIs3_2),.dout(w_dff_B_Z8pmxG6x4_2),.clk(gclk));
	jdff dff_B_3I2OLXAW5_2(.din(w_dff_B_Z8pmxG6x4_2),.dout(w_dff_B_3I2OLXAW5_2),.clk(gclk));
	jdff dff_B_y2dODrBV9_2(.din(w_dff_B_3I2OLXAW5_2),.dout(w_dff_B_y2dODrBV9_2),.clk(gclk));
	jdff dff_B_JycJK9A57_2(.din(w_dff_B_y2dODrBV9_2),.dout(w_dff_B_JycJK9A57_2),.clk(gclk));
	jdff dff_B_skrfLLlq6_2(.din(w_dff_B_JycJK9A57_2),.dout(w_dff_B_skrfLLlq6_2),.clk(gclk));
	jdff dff_B_KKwUwbUc9_2(.din(w_dff_B_skrfLLlq6_2),.dout(w_dff_B_KKwUwbUc9_2),.clk(gclk));
	jdff dff_B_ls1dPspC9_2(.din(w_dff_B_KKwUwbUc9_2),.dout(w_dff_B_ls1dPspC9_2),.clk(gclk));
	jdff dff_B_97ku6Fek6_2(.din(w_dff_B_ls1dPspC9_2),.dout(w_dff_B_97ku6Fek6_2),.clk(gclk));
	jdff dff_B_LtOycfXv9_2(.din(w_dff_B_97ku6Fek6_2),.dout(w_dff_B_LtOycfXv9_2),.clk(gclk));
	jdff dff_B_D7Tzzv8c7_2(.din(w_dff_B_LtOycfXv9_2),.dout(w_dff_B_D7Tzzv8c7_2),.clk(gclk));
	jdff dff_B_rQItFjMI2_2(.din(w_dff_B_D7Tzzv8c7_2),.dout(w_dff_B_rQItFjMI2_2),.clk(gclk));
	jdff dff_B_pKOH8t5A6_2(.din(w_dff_B_rQItFjMI2_2),.dout(w_dff_B_pKOH8t5A6_2),.clk(gclk));
	jdff dff_B_BjEyFtRN9_2(.din(w_dff_B_pKOH8t5A6_2),.dout(w_dff_B_BjEyFtRN9_2),.clk(gclk));
	jdff dff_B_3KDamCFW5_2(.din(w_dff_B_BjEyFtRN9_2),.dout(w_dff_B_3KDamCFW5_2),.clk(gclk));
	jdff dff_B_WpgIoqTT1_2(.din(w_dff_B_3KDamCFW5_2),.dout(w_dff_B_WpgIoqTT1_2),.clk(gclk));
	jdff dff_B_98cckcgj2_2(.din(w_dff_B_WpgIoqTT1_2),.dout(w_dff_B_98cckcgj2_2),.clk(gclk));
	jdff dff_B_JKaAiQVz3_2(.din(w_dff_B_98cckcgj2_2),.dout(w_dff_B_JKaAiQVz3_2),.clk(gclk));
	jdff dff_B_OPgm1r9m1_2(.din(w_dff_B_JKaAiQVz3_2),.dout(w_dff_B_OPgm1r9m1_2),.clk(gclk));
	jdff dff_B_ptNdr2Sq4_2(.din(w_dff_B_OPgm1r9m1_2),.dout(w_dff_B_ptNdr2Sq4_2),.clk(gclk));
	jdff dff_B_zABN6XwR5_2(.din(w_dff_B_ptNdr2Sq4_2),.dout(w_dff_B_zABN6XwR5_2),.clk(gclk));
	jdff dff_B_N0c5WKwz1_2(.din(w_dff_B_zABN6XwR5_2),.dout(w_dff_B_N0c5WKwz1_2),.clk(gclk));
	jdff dff_B_eKkciStW7_2(.din(w_dff_B_N0c5WKwz1_2),.dout(w_dff_B_eKkciStW7_2),.clk(gclk));
	jdff dff_B_l2Pjn05G8_2(.din(w_dff_B_eKkciStW7_2),.dout(w_dff_B_l2Pjn05G8_2),.clk(gclk));
	jdff dff_B_OccyCEz61_2(.din(n1641),.dout(w_dff_B_OccyCEz61_2),.clk(gclk));
	jdff dff_B_iOqyTgmz1_1(.din(n1639),.dout(w_dff_B_iOqyTgmz1_1),.clk(gclk));
	jdff dff_B_YWYmBhFV4_2(.din(n1581),.dout(w_dff_B_YWYmBhFV4_2),.clk(gclk));
	jdff dff_B_C5IuBdWk8_2(.din(w_dff_B_YWYmBhFV4_2),.dout(w_dff_B_C5IuBdWk8_2),.clk(gclk));
	jdff dff_B_yT3Ko8cJ6_2(.din(w_dff_B_C5IuBdWk8_2),.dout(w_dff_B_yT3Ko8cJ6_2),.clk(gclk));
	jdff dff_B_qp6htva55_2(.din(w_dff_B_yT3Ko8cJ6_2),.dout(w_dff_B_qp6htva55_2),.clk(gclk));
	jdff dff_B_bvbiLwZA9_2(.din(w_dff_B_qp6htva55_2),.dout(w_dff_B_bvbiLwZA9_2),.clk(gclk));
	jdff dff_B_poTebLeO3_2(.din(w_dff_B_bvbiLwZA9_2),.dout(w_dff_B_poTebLeO3_2),.clk(gclk));
	jdff dff_B_W7kih9lB0_2(.din(w_dff_B_poTebLeO3_2),.dout(w_dff_B_W7kih9lB0_2),.clk(gclk));
	jdff dff_B_V9rExQbr4_2(.din(w_dff_B_W7kih9lB0_2),.dout(w_dff_B_V9rExQbr4_2),.clk(gclk));
	jdff dff_B_pRXZDnhe0_2(.din(w_dff_B_V9rExQbr4_2),.dout(w_dff_B_pRXZDnhe0_2),.clk(gclk));
	jdff dff_B_agFrEuub0_2(.din(w_dff_B_pRXZDnhe0_2),.dout(w_dff_B_agFrEuub0_2),.clk(gclk));
	jdff dff_B_n9TI68tR3_2(.din(w_dff_B_agFrEuub0_2),.dout(w_dff_B_n9TI68tR3_2),.clk(gclk));
	jdff dff_B_xjaRXSKH7_2(.din(w_dff_B_n9TI68tR3_2),.dout(w_dff_B_xjaRXSKH7_2),.clk(gclk));
	jdff dff_B_9dIkEzHf6_2(.din(w_dff_B_xjaRXSKH7_2),.dout(w_dff_B_9dIkEzHf6_2),.clk(gclk));
	jdff dff_B_g1MTViux5_2(.din(w_dff_B_9dIkEzHf6_2),.dout(w_dff_B_g1MTViux5_2),.clk(gclk));
	jdff dff_B_d1yHmxSt4_2(.din(w_dff_B_g1MTViux5_2),.dout(w_dff_B_d1yHmxSt4_2),.clk(gclk));
	jdff dff_B_dreVPFfK2_2(.din(w_dff_B_d1yHmxSt4_2),.dout(w_dff_B_dreVPFfK2_2),.clk(gclk));
	jdff dff_B_WpJs6XmR4_2(.din(w_dff_B_dreVPFfK2_2),.dout(w_dff_B_WpJs6XmR4_2),.clk(gclk));
	jdff dff_B_aLm4x0ia2_2(.din(w_dff_B_WpJs6XmR4_2),.dout(w_dff_B_aLm4x0ia2_2),.clk(gclk));
	jdff dff_B_EZdMmF1q9_2(.din(w_dff_B_aLm4x0ia2_2),.dout(w_dff_B_EZdMmF1q9_2),.clk(gclk));
	jdff dff_B_bKkbuJZI2_2(.din(w_dff_B_EZdMmF1q9_2),.dout(w_dff_B_bKkbuJZI2_2),.clk(gclk));
	jdff dff_B_3VpGV4EA7_2(.din(w_dff_B_bKkbuJZI2_2),.dout(w_dff_B_3VpGV4EA7_2),.clk(gclk));
	jdff dff_B_qqSxGeDW7_2(.din(w_dff_B_3VpGV4EA7_2),.dout(w_dff_B_qqSxGeDW7_2),.clk(gclk));
	jdff dff_B_EqKbW2G49_2(.din(w_dff_B_qqSxGeDW7_2),.dout(w_dff_B_EqKbW2G49_2),.clk(gclk));
	jdff dff_B_rcIcUfog5_2(.din(w_dff_B_EqKbW2G49_2),.dout(w_dff_B_rcIcUfog5_2),.clk(gclk));
	jdff dff_B_dCfeVtiP2_2(.din(w_dff_B_rcIcUfog5_2),.dout(w_dff_B_dCfeVtiP2_2),.clk(gclk));
	jdff dff_B_5d7MW6cc9_2(.din(w_dff_B_dCfeVtiP2_2),.dout(w_dff_B_5d7MW6cc9_2),.clk(gclk));
	jdff dff_B_dLXWsxlb4_2(.din(w_dff_B_5d7MW6cc9_2),.dout(w_dff_B_dLXWsxlb4_2),.clk(gclk));
	jdff dff_B_Bm6amHFC5_2(.din(w_dff_B_dLXWsxlb4_2),.dout(w_dff_B_Bm6amHFC5_2),.clk(gclk));
	jdff dff_B_XaRubCkU3_2(.din(w_dff_B_Bm6amHFC5_2),.dout(w_dff_B_XaRubCkU3_2),.clk(gclk));
	jdff dff_B_bgeYgFYi4_2(.din(w_dff_B_XaRubCkU3_2),.dout(w_dff_B_bgeYgFYi4_2),.clk(gclk));
	jdff dff_B_fvvSlpHj4_2(.din(w_dff_B_bgeYgFYi4_2),.dout(w_dff_B_fvvSlpHj4_2),.clk(gclk));
	jdff dff_B_piK1THr49_2(.din(n1584),.dout(w_dff_B_piK1THr49_2),.clk(gclk));
	jdff dff_B_Nlcbd72D3_1(.din(n1582),.dout(w_dff_B_Nlcbd72D3_1),.clk(gclk));
	jdff dff_B_2HPEFLM82_2(.din(n1517),.dout(w_dff_B_2HPEFLM82_2),.clk(gclk));
	jdff dff_B_vWr7eoBR6_2(.din(w_dff_B_2HPEFLM82_2),.dout(w_dff_B_vWr7eoBR6_2),.clk(gclk));
	jdff dff_B_rg7FKUR23_2(.din(w_dff_B_vWr7eoBR6_2),.dout(w_dff_B_rg7FKUR23_2),.clk(gclk));
	jdff dff_B_FApnZ9P93_2(.din(w_dff_B_rg7FKUR23_2),.dout(w_dff_B_FApnZ9P93_2),.clk(gclk));
	jdff dff_B_cUkMYVlJ3_2(.din(w_dff_B_FApnZ9P93_2),.dout(w_dff_B_cUkMYVlJ3_2),.clk(gclk));
	jdff dff_B_hDCcouWO2_2(.din(w_dff_B_cUkMYVlJ3_2),.dout(w_dff_B_hDCcouWO2_2),.clk(gclk));
	jdff dff_B_g61wtwJA1_2(.din(w_dff_B_hDCcouWO2_2),.dout(w_dff_B_g61wtwJA1_2),.clk(gclk));
	jdff dff_B_iicfxtvR4_2(.din(w_dff_B_g61wtwJA1_2),.dout(w_dff_B_iicfxtvR4_2),.clk(gclk));
	jdff dff_B_TaAUicxh6_2(.din(w_dff_B_iicfxtvR4_2),.dout(w_dff_B_TaAUicxh6_2),.clk(gclk));
	jdff dff_B_0qzNvZV34_2(.din(w_dff_B_TaAUicxh6_2),.dout(w_dff_B_0qzNvZV34_2),.clk(gclk));
	jdff dff_B_3omzJURq5_2(.din(w_dff_B_0qzNvZV34_2),.dout(w_dff_B_3omzJURq5_2),.clk(gclk));
	jdff dff_B_pp4YLLXZ8_2(.din(w_dff_B_3omzJURq5_2),.dout(w_dff_B_pp4YLLXZ8_2),.clk(gclk));
	jdff dff_B_xTuqZ6hU4_2(.din(w_dff_B_pp4YLLXZ8_2),.dout(w_dff_B_xTuqZ6hU4_2),.clk(gclk));
	jdff dff_B_q975WHsz1_2(.din(w_dff_B_xTuqZ6hU4_2),.dout(w_dff_B_q975WHsz1_2),.clk(gclk));
	jdff dff_B_juriTZ5p0_2(.din(w_dff_B_q975WHsz1_2),.dout(w_dff_B_juriTZ5p0_2),.clk(gclk));
	jdff dff_B_J1q0t3i26_2(.din(w_dff_B_juriTZ5p0_2),.dout(w_dff_B_J1q0t3i26_2),.clk(gclk));
	jdff dff_B_y6c4tBer9_2(.din(w_dff_B_J1q0t3i26_2),.dout(w_dff_B_y6c4tBer9_2),.clk(gclk));
	jdff dff_B_OAWuBNqb3_2(.din(w_dff_B_y6c4tBer9_2),.dout(w_dff_B_OAWuBNqb3_2),.clk(gclk));
	jdff dff_B_VDzypX2G8_2(.din(w_dff_B_OAWuBNqb3_2),.dout(w_dff_B_VDzypX2G8_2),.clk(gclk));
	jdff dff_B_Y4V0EiMH2_2(.din(w_dff_B_VDzypX2G8_2),.dout(w_dff_B_Y4V0EiMH2_2),.clk(gclk));
	jdff dff_B_KuJouY0T0_2(.din(w_dff_B_Y4V0EiMH2_2),.dout(w_dff_B_KuJouY0T0_2),.clk(gclk));
	jdff dff_B_YijVKpmQ0_2(.din(w_dff_B_KuJouY0T0_2),.dout(w_dff_B_YijVKpmQ0_2),.clk(gclk));
	jdff dff_B_DomJE4z29_2(.din(w_dff_B_YijVKpmQ0_2),.dout(w_dff_B_DomJE4z29_2),.clk(gclk));
	jdff dff_B_1TZ6l6d11_2(.din(w_dff_B_DomJE4z29_2),.dout(w_dff_B_1TZ6l6d11_2),.clk(gclk));
	jdff dff_B_OnPlRJhm9_2(.din(w_dff_B_1TZ6l6d11_2),.dout(w_dff_B_OnPlRJhm9_2),.clk(gclk));
	jdff dff_B_tC22cMcN4_2(.din(w_dff_B_OnPlRJhm9_2),.dout(w_dff_B_tC22cMcN4_2),.clk(gclk));
	jdff dff_B_5tLJTjaH8_2(.din(w_dff_B_tC22cMcN4_2),.dout(w_dff_B_5tLJTjaH8_2),.clk(gclk));
	jdff dff_B_6DxEcXa09_2(.din(w_dff_B_5tLJTjaH8_2),.dout(w_dff_B_6DxEcXa09_2),.clk(gclk));
	jdff dff_B_S34dDBt10_2(.din(n1520),.dout(w_dff_B_S34dDBt10_2),.clk(gclk));
	jdff dff_B_zXMfh2tW4_1(.din(n1518),.dout(w_dff_B_zXMfh2tW4_1),.clk(gclk));
	jdff dff_B_W7Dz1Qnz1_2(.din(n1446),.dout(w_dff_B_W7Dz1Qnz1_2),.clk(gclk));
	jdff dff_B_DyLsH0OY5_2(.din(w_dff_B_W7Dz1Qnz1_2),.dout(w_dff_B_DyLsH0OY5_2),.clk(gclk));
	jdff dff_B_9mO2WHov3_2(.din(w_dff_B_DyLsH0OY5_2),.dout(w_dff_B_9mO2WHov3_2),.clk(gclk));
	jdff dff_B_0bjRPH6k2_2(.din(w_dff_B_9mO2WHov3_2),.dout(w_dff_B_0bjRPH6k2_2),.clk(gclk));
	jdff dff_B_sYUNCPeO4_2(.din(w_dff_B_0bjRPH6k2_2),.dout(w_dff_B_sYUNCPeO4_2),.clk(gclk));
	jdff dff_B_L4ykzywp6_2(.din(w_dff_B_sYUNCPeO4_2),.dout(w_dff_B_L4ykzywp6_2),.clk(gclk));
	jdff dff_B_9VKWKBlF6_2(.din(w_dff_B_L4ykzywp6_2),.dout(w_dff_B_9VKWKBlF6_2),.clk(gclk));
	jdff dff_B_n0VqNGXr2_2(.din(w_dff_B_9VKWKBlF6_2),.dout(w_dff_B_n0VqNGXr2_2),.clk(gclk));
	jdff dff_B_b7cB2ACx8_2(.din(w_dff_B_n0VqNGXr2_2),.dout(w_dff_B_b7cB2ACx8_2),.clk(gclk));
	jdff dff_B_mEo84peu1_2(.din(w_dff_B_b7cB2ACx8_2),.dout(w_dff_B_mEo84peu1_2),.clk(gclk));
	jdff dff_B_sr8ONZMh7_2(.din(w_dff_B_mEo84peu1_2),.dout(w_dff_B_sr8ONZMh7_2),.clk(gclk));
	jdff dff_B_hDD2sypM9_2(.din(w_dff_B_sr8ONZMh7_2),.dout(w_dff_B_hDD2sypM9_2),.clk(gclk));
	jdff dff_B_4uzQCgt64_2(.din(w_dff_B_hDD2sypM9_2),.dout(w_dff_B_4uzQCgt64_2),.clk(gclk));
	jdff dff_B_Gjn9kFKJ0_2(.din(w_dff_B_4uzQCgt64_2),.dout(w_dff_B_Gjn9kFKJ0_2),.clk(gclk));
	jdff dff_B_DTUizuuB1_2(.din(w_dff_B_Gjn9kFKJ0_2),.dout(w_dff_B_DTUizuuB1_2),.clk(gclk));
	jdff dff_B_1rBTGPXP2_2(.din(w_dff_B_DTUizuuB1_2),.dout(w_dff_B_1rBTGPXP2_2),.clk(gclk));
	jdff dff_B_c2ds4AcS7_2(.din(w_dff_B_1rBTGPXP2_2),.dout(w_dff_B_c2ds4AcS7_2),.clk(gclk));
	jdff dff_B_LVOKVTvM5_2(.din(w_dff_B_c2ds4AcS7_2),.dout(w_dff_B_LVOKVTvM5_2),.clk(gclk));
	jdff dff_B_7r2ABg1S5_2(.din(w_dff_B_LVOKVTvM5_2),.dout(w_dff_B_7r2ABg1S5_2),.clk(gclk));
	jdff dff_B_e1qQgB797_2(.din(w_dff_B_7r2ABg1S5_2),.dout(w_dff_B_e1qQgB797_2),.clk(gclk));
	jdff dff_B_GbTO9bFl8_2(.din(w_dff_B_e1qQgB797_2),.dout(w_dff_B_GbTO9bFl8_2),.clk(gclk));
	jdff dff_B_gEukhRpQ0_2(.din(w_dff_B_GbTO9bFl8_2),.dout(w_dff_B_gEukhRpQ0_2),.clk(gclk));
	jdff dff_B_Osy9HHTE8_2(.din(w_dff_B_gEukhRpQ0_2),.dout(w_dff_B_Osy9HHTE8_2),.clk(gclk));
	jdff dff_B_NJ0E4Suu2_2(.din(w_dff_B_Osy9HHTE8_2),.dout(w_dff_B_NJ0E4Suu2_2),.clk(gclk));
	jdff dff_B_q9yyD1qM7_2(.din(w_dff_B_NJ0E4Suu2_2),.dout(w_dff_B_q9yyD1qM7_2),.clk(gclk));
	jdff dff_B_Ym1N6bAQ5_2(.din(n1449),.dout(w_dff_B_Ym1N6bAQ5_2),.clk(gclk));
	jdff dff_B_aqaLGXOT4_1(.din(n1447),.dout(w_dff_B_aqaLGXOT4_1),.clk(gclk));
	jdff dff_B_oQd8Drrb6_2(.din(n1368),.dout(w_dff_B_oQd8Drrb6_2),.clk(gclk));
	jdff dff_B_TgUPBvNo2_2(.din(w_dff_B_oQd8Drrb6_2),.dout(w_dff_B_TgUPBvNo2_2),.clk(gclk));
	jdff dff_B_hGutAvSs1_2(.din(w_dff_B_TgUPBvNo2_2),.dout(w_dff_B_hGutAvSs1_2),.clk(gclk));
	jdff dff_B_dHnHjPAi6_2(.din(w_dff_B_hGutAvSs1_2),.dout(w_dff_B_dHnHjPAi6_2),.clk(gclk));
	jdff dff_B_fdXZGFd91_2(.din(w_dff_B_dHnHjPAi6_2),.dout(w_dff_B_fdXZGFd91_2),.clk(gclk));
	jdff dff_B_aCBknWDn7_2(.din(w_dff_B_fdXZGFd91_2),.dout(w_dff_B_aCBknWDn7_2),.clk(gclk));
	jdff dff_B_aRnaJa3d3_2(.din(w_dff_B_aCBknWDn7_2),.dout(w_dff_B_aRnaJa3d3_2),.clk(gclk));
	jdff dff_B_SVsWrV5Y1_2(.din(w_dff_B_aRnaJa3d3_2),.dout(w_dff_B_SVsWrV5Y1_2),.clk(gclk));
	jdff dff_B_mXgxtTEs9_2(.din(w_dff_B_SVsWrV5Y1_2),.dout(w_dff_B_mXgxtTEs9_2),.clk(gclk));
	jdff dff_B_3LXiQ8wr5_2(.din(w_dff_B_mXgxtTEs9_2),.dout(w_dff_B_3LXiQ8wr5_2),.clk(gclk));
	jdff dff_B_ZCPFiMjh8_2(.din(w_dff_B_3LXiQ8wr5_2),.dout(w_dff_B_ZCPFiMjh8_2),.clk(gclk));
	jdff dff_B_JupzjdSE7_2(.din(w_dff_B_ZCPFiMjh8_2),.dout(w_dff_B_JupzjdSE7_2),.clk(gclk));
	jdff dff_B_vwvwWmfs9_2(.din(w_dff_B_JupzjdSE7_2),.dout(w_dff_B_vwvwWmfs9_2),.clk(gclk));
	jdff dff_B_d83LMinm0_2(.din(w_dff_B_vwvwWmfs9_2),.dout(w_dff_B_d83LMinm0_2),.clk(gclk));
	jdff dff_B_PT7qa8pG9_2(.din(w_dff_B_d83LMinm0_2),.dout(w_dff_B_PT7qa8pG9_2),.clk(gclk));
	jdff dff_B_5rfZzXRl7_2(.din(w_dff_B_PT7qa8pG9_2),.dout(w_dff_B_5rfZzXRl7_2),.clk(gclk));
	jdff dff_B_K5UsvlC36_2(.din(w_dff_B_5rfZzXRl7_2),.dout(w_dff_B_K5UsvlC36_2),.clk(gclk));
	jdff dff_B_jN0B3Hg38_2(.din(w_dff_B_K5UsvlC36_2),.dout(w_dff_B_jN0B3Hg38_2),.clk(gclk));
	jdff dff_B_bMWuoRQU1_2(.din(w_dff_B_jN0B3Hg38_2),.dout(w_dff_B_bMWuoRQU1_2),.clk(gclk));
	jdff dff_B_08CLUnav2_2(.din(w_dff_B_bMWuoRQU1_2),.dout(w_dff_B_08CLUnav2_2),.clk(gclk));
	jdff dff_B_fGMlVNJy1_2(.din(w_dff_B_08CLUnav2_2),.dout(w_dff_B_fGMlVNJy1_2),.clk(gclk));
	jdff dff_B_Mn7l1HXh8_2(.din(w_dff_B_fGMlVNJy1_2),.dout(w_dff_B_Mn7l1HXh8_2),.clk(gclk));
	jdff dff_B_PRIeYDNt5_2(.din(n1371),.dout(w_dff_B_PRIeYDNt5_2),.clk(gclk));
	jdff dff_B_kdxQH1hD6_1(.din(n1369),.dout(w_dff_B_kdxQH1hD6_1),.clk(gclk));
	jdff dff_B_HCzYG60k7_2(.din(n1283),.dout(w_dff_B_HCzYG60k7_2),.clk(gclk));
	jdff dff_B_5hBk78Fa0_2(.din(w_dff_B_HCzYG60k7_2),.dout(w_dff_B_5hBk78Fa0_2),.clk(gclk));
	jdff dff_B_D6HNnkBD1_2(.din(w_dff_B_5hBk78Fa0_2),.dout(w_dff_B_D6HNnkBD1_2),.clk(gclk));
	jdff dff_B_aUJ5hsqJ0_2(.din(w_dff_B_D6HNnkBD1_2),.dout(w_dff_B_aUJ5hsqJ0_2),.clk(gclk));
	jdff dff_B_eOtt4UFf4_2(.din(w_dff_B_aUJ5hsqJ0_2),.dout(w_dff_B_eOtt4UFf4_2),.clk(gclk));
	jdff dff_B_LHW0FfEu0_2(.din(w_dff_B_eOtt4UFf4_2),.dout(w_dff_B_LHW0FfEu0_2),.clk(gclk));
	jdff dff_B_mWpSzgvl5_2(.din(w_dff_B_LHW0FfEu0_2),.dout(w_dff_B_mWpSzgvl5_2),.clk(gclk));
	jdff dff_B_ElZNEvgM4_2(.din(w_dff_B_mWpSzgvl5_2),.dout(w_dff_B_ElZNEvgM4_2),.clk(gclk));
	jdff dff_B_SKg6nO6k2_2(.din(w_dff_B_ElZNEvgM4_2),.dout(w_dff_B_SKg6nO6k2_2),.clk(gclk));
	jdff dff_B_xaUDYiJt9_2(.din(w_dff_B_SKg6nO6k2_2),.dout(w_dff_B_xaUDYiJt9_2),.clk(gclk));
	jdff dff_B_ZLUP5LaM9_2(.din(w_dff_B_xaUDYiJt9_2),.dout(w_dff_B_ZLUP5LaM9_2),.clk(gclk));
	jdff dff_B_NeEBMxcE6_2(.din(w_dff_B_ZLUP5LaM9_2),.dout(w_dff_B_NeEBMxcE6_2),.clk(gclk));
	jdff dff_B_ydTr7wtZ0_2(.din(w_dff_B_NeEBMxcE6_2),.dout(w_dff_B_ydTr7wtZ0_2),.clk(gclk));
	jdff dff_B_osMTjY5i1_2(.din(w_dff_B_ydTr7wtZ0_2),.dout(w_dff_B_osMTjY5i1_2),.clk(gclk));
	jdff dff_B_AffJraA94_2(.din(w_dff_B_osMTjY5i1_2),.dout(w_dff_B_AffJraA94_2),.clk(gclk));
	jdff dff_B_Z7dk3cDU5_2(.din(w_dff_B_AffJraA94_2),.dout(w_dff_B_Z7dk3cDU5_2),.clk(gclk));
	jdff dff_B_UubY8gNc7_2(.din(w_dff_B_Z7dk3cDU5_2),.dout(w_dff_B_UubY8gNc7_2),.clk(gclk));
	jdff dff_B_RXBU1v445_2(.din(w_dff_B_UubY8gNc7_2),.dout(w_dff_B_RXBU1v445_2),.clk(gclk));
	jdff dff_B_fnGQfLsP3_2(.din(w_dff_B_RXBU1v445_2),.dout(w_dff_B_fnGQfLsP3_2),.clk(gclk));
	jdff dff_B_UslNWrpR7_2(.din(n1286),.dout(w_dff_B_UslNWrpR7_2),.clk(gclk));
	jdff dff_B_r7ZG6dqT3_1(.din(n1284),.dout(w_dff_B_r7ZG6dqT3_1),.clk(gclk));
	jdff dff_B_k6mxmWdS7_2(.din(n1193),.dout(w_dff_B_k6mxmWdS7_2),.clk(gclk));
	jdff dff_B_5WVxsyCe5_2(.din(w_dff_B_k6mxmWdS7_2),.dout(w_dff_B_5WVxsyCe5_2),.clk(gclk));
	jdff dff_B_KCYjFm1k4_2(.din(w_dff_B_5WVxsyCe5_2),.dout(w_dff_B_KCYjFm1k4_2),.clk(gclk));
	jdff dff_B_6jMRu9FB5_2(.din(w_dff_B_KCYjFm1k4_2),.dout(w_dff_B_6jMRu9FB5_2),.clk(gclk));
	jdff dff_B_YS6iORA66_2(.din(w_dff_B_6jMRu9FB5_2),.dout(w_dff_B_YS6iORA66_2),.clk(gclk));
	jdff dff_B_P0Oa2pEG1_2(.din(w_dff_B_YS6iORA66_2),.dout(w_dff_B_P0Oa2pEG1_2),.clk(gclk));
	jdff dff_B_oCnCQZlL4_2(.din(w_dff_B_P0Oa2pEG1_2),.dout(w_dff_B_oCnCQZlL4_2),.clk(gclk));
	jdff dff_B_AMQ7jfWC0_2(.din(w_dff_B_oCnCQZlL4_2),.dout(w_dff_B_AMQ7jfWC0_2),.clk(gclk));
	jdff dff_B_1RTishND9_2(.din(w_dff_B_AMQ7jfWC0_2),.dout(w_dff_B_1RTishND9_2),.clk(gclk));
	jdff dff_B_IwRWwSvu9_2(.din(w_dff_B_1RTishND9_2),.dout(w_dff_B_IwRWwSvu9_2),.clk(gclk));
	jdff dff_B_k5bhNNs23_2(.din(w_dff_B_IwRWwSvu9_2),.dout(w_dff_B_k5bhNNs23_2),.clk(gclk));
	jdff dff_B_A97wTBuN9_2(.din(w_dff_B_k5bhNNs23_2),.dout(w_dff_B_A97wTBuN9_2),.clk(gclk));
	jdff dff_B_ENSOQdib9_2(.din(w_dff_B_A97wTBuN9_2),.dout(w_dff_B_ENSOQdib9_2),.clk(gclk));
	jdff dff_B_WNh5RNnA5_2(.din(w_dff_B_ENSOQdib9_2),.dout(w_dff_B_WNh5RNnA5_2),.clk(gclk));
	jdff dff_B_a5XXBoSe0_2(.din(w_dff_B_WNh5RNnA5_2),.dout(w_dff_B_a5XXBoSe0_2),.clk(gclk));
	jdff dff_B_ai4SvB5g3_2(.din(w_dff_B_a5XXBoSe0_2),.dout(w_dff_B_ai4SvB5g3_2),.clk(gclk));
	jdff dff_B_Nz2nYbTU5_2(.din(n1196),.dout(w_dff_B_Nz2nYbTU5_2),.clk(gclk));
	jdff dff_B_KMgHgW2O2_1(.din(n1194),.dout(w_dff_B_KMgHgW2O2_1),.clk(gclk));
	jdff dff_B_QMurNLlQ7_2(.din(n1089),.dout(w_dff_B_QMurNLlQ7_2),.clk(gclk));
	jdff dff_B_dzC7afe74_2(.din(w_dff_B_QMurNLlQ7_2),.dout(w_dff_B_dzC7afe74_2),.clk(gclk));
	jdff dff_B_B2Mgau256_2(.din(w_dff_B_dzC7afe74_2),.dout(w_dff_B_B2Mgau256_2),.clk(gclk));
	jdff dff_B_a8E0En2V6_2(.din(w_dff_B_B2Mgau256_2),.dout(w_dff_B_a8E0En2V6_2),.clk(gclk));
	jdff dff_B_TzQJEmA32_2(.din(w_dff_B_a8E0En2V6_2),.dout(w_dff_B_TzQJEmA32_2),.clk(gclk));
	jdff dff_B_DGDETqys6_2(.din(w_dff_B_TzQJEmA32_2),.dout(w_dff_B_DGDETqys6_2),.clk(gclk));
	jdff dff_B_NDSInMWX4_2(.din(w_dff_B_DGDETqys6_2),.dout(w_dff_B_NDSInMWX4_2),.clk(gclk));
	jdff dff_B_h9CZyYT61_2(.din(w_dff_B_NDSInMWX4_2),.dout(w_dff_B_h9CZyYT61_2),.clk(gclk));
	jdff dff_B_CusKAVL52_2(.din(w_dff_B_h9CZyYT61_2),.dout(w_dff_B_CusKAVL52_2),.clk(gclk));
	jdff dff_B_QxyJPTha4_2(.din(w_dff_B_CusKAVL52_2),.dout(w_dff_B_QxyJPTha4_2),.clk(gclk));
	jdff dff_B_rDtdTpkI3_2(.din(w_dff_B_QxyJPTha4_2),.dout(w_dff_B_rDtdTpkI3_2),.clk(gclk));
	jdff dff_B_yIey17ab9_2(.din(w_dff_B_rDtdTpkI3_2),.dout(w_dff_B_yIey17ab9_2),.clk(gclk));
	jdff dff_B_4efL7dCV5_2(.din(w_dff_B_yIey17ab9_2),.dout(w_dff_B_4efL7dCV5_2),.clk(gclk));
	jdff dff_B_HU2GbyaZ7_2(.din(n1092),.dout(w_dff_B_HU2GbyaZ7_2),.clk(gclk));
	jdff dff_B_YI5hYO794_1(.din(n1090),.dout(w_dff_B_YI5hYO794_1),.clk(gclk));
	jdff dff_B_4uwK1ZRk4_2(.din(n991),.dout(w_dff_B_4uwK1ZRk4_2),.clk(gclk));
	jdff dff_B_z2oclxAG8_2(.din(w_dff_B_4uwK1ZRk4_2),.dout(w_dff_B_z2oclxAG8_2),.clk(gclk));
	jdff dff_B_yU3poFZb5_2(.din(w_dff_B_z2oclxAG8_2),.dout(w_dff_B_yU3poFZb5_2),.clk(gclk));
	jdff dff_B_5aowa2yR4_2(.din(w_dff_B_yU3poFZb5_2),.dout(w_dff_B_5aowa2yR4_2),.clk(gclk));
	jdff dff_B_vqkZb6233_2(.din(w_dff_B_5aowa2yR4_2),.dout(w_dff_B_vqkZb6233_2),.clk(gclk));
	jdff dff_B_DwLfJLt02_2(.din(w_dff_B_vqkZb6233_2),.dout(w_dff_B_DwLfJLt02_2),.clk(gclk));
	jdff dff_B_OmpSV0WB2_2(.din(w_dff_B_DwLfJLt02_2),.dout(w_dff_B_OmpSV0WB2_2),.clk(gclk));
	jdff dff_B_AOzvZOFq4_2(.din(w_dff_B_OmpSV0WB2_2),.dout(w_dff_B_AOzvZOFq4_2),.clk(gclk));
	jdff dff_B_F4IlZSsO1_2(.din(w_dff_B_AOzvZOFq4_2),.dout(w_dff_B_F4IlZSsO1_2),.clk(gclk));
	jdff dff_B_06ARLHTF0_2(.din(w_dff_B_F4IlZSsO1_2),.dout(w_dff_B_06ARLHTF0_2),.clk(gclk));
	jdff dff_B_0FF0RhK38_1(.din(n992),.dout(w_dff_B_0FF0RhK38_1),.clk(gclk));
	jdff dff_B_1PVUAIIw9_2(.din(n886),.dout(w_dff_B_1PVUAIIw9_2),.clk(gclk));
	jdff dff_B_JQXRx6Ps8_2(.din(w_dff_B_1PVUAIIw9_2),.dout(w_dff_B_JQXRx6Ps8_2),.clk(gclk));
	jdff dff_B_JjBpuBFH5_2(.din(w_dff_B_JQXRx6Ps8_2),.dout(w_dff_B_JjBpuBFH5_2),.clk(gclk));
	jdff dff_B_hgv5c3tx9_2(.din(w_dff_B_JjBpuBFH5_2),.dout(w_dff_B_hgv5c3tx9_2),.clk(gclk));
	jdff dff_B_cRdn1g5B0_2(.din(w_dff_B_hgv5c3tx9_2),.dout(w_dff_B_cRdn1g5B0_2),.clk(gclk));
	jdff dff_B_eMgF42nM1_2(.din(w_dff_B_cRdn1g5B0_2),.dout(w_dff_B_eMgF42nM1_2),.clk(gclk));
	jdff dff_B_DRvW5Fr76_2(.din(w_dff_B_eMgF42nM1_2),.dout(w_dff_B_DRvW5Fr76_2),.clk(gclk));
	jdff dff_B_Zhi0614O5_2(.din(w_dff_B_DRvW5Fr76_2),.dout(w_dff_B_Zhi0614O5_2),.clk(gclk));
	jdff dff_B_pITryFcZ5_1(.din(n887),.dout(w_dff_B_pITryFcZ5_1),.clk(gclk));
	jdff dff_B_oXpog3fo0_2(.din(n787),.dout(w_dff_B_oXpog3fo0_2),.clk(gclk));
	jdff dff_B_CODLarTi9_2(.din(w_dff_B_oXpog3fo0_2),.dout(w_dff_B_CODLarTi9_2),.clk(gclk));
	jdff dff_B_GwxsGOQE2_2(.din(w_dff_B_CODLarTi9_2),.dout(w_dff_B_GwxsGOQE2_2),.clk(gclk));
	jdff dff_B_nzZv25Aw9_2(.din(w_dff_B_GwxsGOQE2_2),.dout(w_dff_B_nzZv25Aw9_2),.clk(gclk));
	jdff dff_B_Y1X9YCny9_2(.din(w_dff_B_nzZv25Aw9_2),.dout(w_dff_B_Y1X9YCny9_2),.clk(gclk));
	jdff dff_B_zeb0jvwG4_2(.din(w_dff_B_Y1X9YCny9_2),.dout(w_dff_B_zeb0jvwG4_2),.clk(gclk));
	jdff dff_B_GAMWtoFq2_2(.din(n803),.dout(w_dff_B_GAMWtoFq2_2),.clk(gclk));
	jdff dff_B_K5V2KHjU3_1(.din(n788),.dout(w_dff_B_K5V2KHjU3_1),.clk(gclk));
	jdff dff_B_wuGYaRmU8_1(.din(w_dff_B_K5V2KHjU3_1),.dout(w_dff_B_wuGYaRmU8_1),.clk(gclk));
	jdff dff_B_e5I1tcpN9_1(.din(w_dff_B_wuGYaRmU8_1),.dout(w_dff_B_e5I1tcpN9_1),.clk(gclk));
	jdff dff_B_WYYKT4UZ3_1(.din(w_dff_B_e5I1tcpN9_1),.dout(w_dff_B_WYYKT4UZ3_1),.clk(gclk));
	jdff dff_B_D6eKyeyl8_0(.din(n703),.dout(w_dff_B_D6eKyeyl8_0),.clk(gclk));
	jdff dff_A_8ydGlACv3_0(.dout(w_n702_0[0]),.din(w_dff_A_8ydGlACv3_0),.clk(gclk));
	jdff dff_A_3m1VZbBZ2_0(.dout(w_dff_A_8ydGlACv3_0),.din(w_dff_A_3m1VZbBZ2_0),.clk(gclk));
	jdff dff_B_LyhL8Snl8_1(.din(n696),.dout(w_dff_B_LyhL8Snl8_1),.clk(gclk));
	jdff dff_B_YuHExj7R4_1(.din(w_dff_B_LyhL8Snl8_1),.dout(w_dff_B_YuHExj7R4_1),.clk(gclk));
	jdff dff_A_48Fakt9R8_0(.dout(w_n607_0[0]),.din(w_dff_A_48Fakt9R8_0),.clk(gclk));
	jdff dff_A_yBVmxsN03_1(.dout(w_n607_0[1]),.din(w_dff_A_yBVmxsN03_1),.clk(gclk));
	jdff dff_A_1dokVTgx8_1(.dout(w_dff_A_yBVmxsN03_1),.din(w_dff_A_1dokVTgx8_1),.clk(gclk));
	jdff dff_A_i9qFOE6m4_1(.dout(w_n694_0[1]),.din(w_dff_A_i9qFOE6m4_1),.clk(gclk));
	jdff dff_A_oQuvQBQq3_1(.dout(w_dff_A_i9qFOE6m4_1),.din(w_dff_A_oQuvQBQq3_1),.clk(gclk));
	jdff dff_A_EKgaLSVg7_1(.dout(w_dff_A_oQuvQBQq3_1),.din(w_dff_A_EKgaLSVg7_1),.clk(gclk));
	jdff dff_A_Kcc6bB7L1_1(.dout(w_dff_A_EKgaLSVg7_1),.din(w_dff_A_Kcc6bB7L1_1),.clk(gclk));
	jdff dff_B_BIrgQ7AT7_1(.din(n1819),.dout(w_dff_B_BIrgQ7AT7_1),.clk(gclk));
	jdff dff_A_ssrXAKtQ0_1(.dout(w_n1801_0[1]),.din(w_dff_A_ssrXAKtQ0_1),.clk(gclk));
	jdff dff_B_BXjl0G2O6_1(.din(n1799),.dout(w_dff_B_BXjl0G2O6_1),.clk(gclk));
	jdff dff_B_lrFDyZ1k0_2(.din(n1770),.dout(w_dff_B_lrFDyZ1k0_2),.clk(gclk));
	jdff dff_B_smNHENwB4_2(.din(w_dff_B_lrFDyZ1k0_2),.dout(w_dff_B_smNHENwB4_2),.clk(gclk));
	jdff dff_B_JHIdWpMv9_2(.din(w_dff_B_smNHENwB4_2),.dout(w_dff_B_JHIdWpMv9_2),.clk(gclk));
	jdff dff_B_WIShTbn59_2(.din(w_dff_B_JHIdWpMv9_2),.dout(w_dff_B_WIShTbn59_2),.clk(gclk));
	jdff dff_B_BgYXh6C66_2(.din(w_dff_B_WIShTbn59_2),.dout(w_dff_B_BgYXh6C66_2),.clk(gclk));
	jdff dff_B_cUPdgFNU6_2(.din(w_dff_B_BgYXh6C66_2),.dout(w_dff_B_cUPdgFNU6_2),.clk(gclk));
	jdff dff_B_VrUDwbX50_2(.din(w_dff_B_cUPdgFNU6_2),.dout(w_dff_B_VrUDwbX50_2),.clk(gclk));
	jdff dff_B_U7BrJy915_2(.din(w_dff_B_VrUDwbX50_2),.dout(w_dff_B_U7BrJy915_2),.clk(gclk));
	jdff dff_B_aF5daw8L6_2(.din(w_dff_B_U7BrJy915_2),.dout(w_dff_B_aF5daw8L6_2),.clk(gclk));
	jdff dff_B_wyIyIqkM5_2(.din(w_dff_B_aF5daw8L6_2),.dout(w_dff_B_wyIyIqkM5_2),.clk(gclk));
	jdff dff_B_3AnMBDNf9_2(.din(w_dff_B_wyIyIqkM5_2),.dout(w_dff_B_3AnMBDNf9_2),.clk(gclk));
	jdff dff_B_LBUE0QMh1_2(.din(w_dff_B_3AnMBDNf9_2),.dout(w_dff_B_LBUE0QMh1_2),.clk(gclk));
	jdff dff_B_wg6jI9769_2(.din(w_dff_B_LBUE0QMh1_2),.dout(w_dff_B_wg6jI9769_2),.clk(gclk));
	jdff dff_B_6ma86CHJ5_2(.din(w_dff_B_wg6jI9769_2),.dout(w_dff_B_6ma86CHJ5_2),.clk(gclk));
	jdff dff_B_QJhBV3h86_2(.din(w_dff_B_6ma86CHJ5_2),.dout(w_dff_B_QJhBV3h86_2),.clk(gclk));
	jdff dff_B_RGHXScO50_2(.din(w_dff_B_QJhBV3h86_2),.dout(w_dff_B_RGHXScO50_2),.clk(gclk));
	jdff dff_B_cZEYKMmO0_2(.din(w_dff_B_RGHXScO50_2),.dout(w_dff_B_cZEYKMmO0_2),.clk(gclk));
	jdff dff_B_DI1ZpD6Q3_2(.din(w_dff_B_cZEYKMmO0_2),.dout(w_dff_B_DI1ZpD6Q3_2),.clk(gclk));
	jdff dff_B_NkZ1EQx12_2(.din(w_dff_B_DI1ZpD6Q3_2),.dout(w_dff_B_NkZ1EQx12_2),.clk(gclk));
	jdff dff_B_aCHysf9u8_2(.din(w_dff_B_NkZ1EQx12_2),.dout(w_dff_B_aCHysf9u8_2),.clk(gclk));
	jdff dff_B_XUzEbjbv4_2(.din(w_dff_B_aCHysf9u8_2),.dout(w_dff_B_XUzEbjbv4_2),.clk(gclk));
	jdff dff_B_f3RHJg6j9_2(.din(w_dff_B_XUzEbjbv4_2),.dout(w_dff_B_f3RHJg6j9_2),.clk(gclk));
	jdff dff_B_UKlDCxib4_2(.din(w_dff_B_f3RHJg6j9_2),.dout(w_dff_B_UKlDCxib4_2),.clk(gclk));
	jdff dff_B_tp7oMU3c0_2(.din(w_dff_B_UKlDCxib4_2),.dout(w_dff_B_tp7oMU3c0_2),.clk(gclk));
	jdff dff_B_JIMLoSuW5_2(.din(w_dff_B_tp7oMU3c0_2),.dout(w_dff_B_JIMLoSuW5_2),.clk(gclk));
	jdff dff_B_x1k2WNq90_2(.din(w_dff_B_JIMLoSuW5_2),.dout(w_dff_B_x1k2WNq90_2),.clk(gclk));
	jdff dff_B_fl0uf7fw8_2(.din(w_dff_B_x1k2WNq90_2),.dout(w_dff_B_fl0uf7fw8_2),.clk(gclk));
	jdff dff_B_YM43M1rB6_2(.din(w_dff_B_fl0uf7fw8_2),.dout(w_dff_B_YM43M1rB6_2),.clk(gclk));
	jdff dff_B_AZIfTLcq8_2(.din(w_dff_B_YM43M1rB6_2),.dout(w_dff_B_AZIfTLcq8_2),.clk(gclk));
	jdff dff_B_KfcAI0Al0_2(.din(w_dff_B_AZIfTLcq8_2),.dout(w_dff_B_KfcAI0Al0_2),.clk(gclk));
	jdff dff_B_Wi7Nfyqe5_2(.din(w_dff_B_KfcAI0Al0_2),.dout(w_dff_B_Wi7Nfyqe5_2),.clk(gclk));
	jdff dff_B_JQGzFj0b1_2(.din(w_dff_B_Wi7Nfyqe5_2),.dout(w_dff_B_JQGzFj0b1_2),.clk(gclk));
	jdff dff_B_AxRDFDkS5_2(.din(w_dff_B_JQGzFj0b1_2),.dout(w_dff_B_AxRDFDkS5_2),.clk(gclk));
	jdff dff_B_qxyz7S7d4_2(.din(w_dff_B_AxRDFDkS5_2),.dout(w_dff_B_qxyz7S7d4_2),.clk(gclk));
	jdff dff_B_I5ASGsY29_2(.din(w_dff_B_qxyz7S7d4_2),.dout(w_dff_B_I5ASGsY29_2),.clk(gclk));
	jdff dff_B_7eEp03fZ0_2(.din(w_dff_B_I5ASGsY29_2),.dout(w_dff_B_7eEp03fZ0_2),.clk(gclk));
	jdff dff_B_gbZtysXo3_2(.din(w_dff_B_7eEp03fZ0_2),.dout(w_dff_B_gbZtysXo3_2),.clk(gclk));
	jdff dff_B_n29bydAO2_2(.din(w_dff_B_gbZtysXo3_2),.dout(w_dff_B_n29bydAO2_2),.clk(gclk));
	jdff dff_B_5048nYaS6_2(.din(w_dff_B_n29bydAO2_2),.dout(w_dff_B_5048nYaS6_2),.clk(gclk));
	jdff dff_B_0oiRhCew3_2(.din(w_dff_B_5048nYaS6_2),.dout(w_dff_B_0oiRhCew3_2),.clk(gclk));
	jdff dff_B_XLEbZbGh4_2(.din(w_dff_B_0oiRhCew3_2),.dout(w_dff_B_XLEbZbGh4_2),.clk(gclk));
	jdff dff_B_dAbLNxEq4_2(.din(n1773),.dout(w_dff_B_dAbLNxEq4_2),.clk(gclk));
	jdff dff_B_PMZFNPI94_1(.din(n1771),.dout(w_dff_B_PMZFNPI94_1),.clk(gclk));
	jdff dff_B_DebyrMO77_2(.din(n1735),.dout(w_dff_B_DebyrMO77_2),.clk(gclk));
	jdff dff_B_r8H7Kio31_2(.din(w_dff_B_DebyrMO77_2),.dout(w_dff_B_r8H7Kio31_2),.clk(gclk));
	jdff dff_B_T2MKbseA9_2(.din(w_dff_B_r8H7Kio31_2),.dout(w_dff_B_T2MKbseA9_2),.clk(gclk));
	jdff dff_B_2iTkIsY93_2(.din(w_dff_B_T2MKbseA9_2),.dout(w_dff_B_2iTkIsY93_2),.clk(gclk));
	jdff dff_B_YHqQGlAz1_2(.din(w_dff_B_2iTkIsY93_2),.dout(w_dff_B_YHqQGlAz1_2),.clk(gclk));
	jdff dff_B_pN5nbpjh8_2(.din(w_dff_B_YHqQGlAz1_2),.dout(w_dff_B_pN5nbpjh8_2),.clk(gclk));
	jdff dff_B_dYO5KS5O0_2(.din(w_dff_B_pN5nbpjh8_2),.dout(w_dff_B_dYO5KS5O0_2),.clk(gclk));
	jdff dff_B_Y8RYzSaX6_2(.din(w_dff_B_dYO5KS5O0_2),.dout(w_dff_B_Y8RYzSaX6_2),.clk(gclk));
	jdff dff_B_uKw0ccgk4_2(.din(w_dff_B_Y8RYzSaX6_2),.dout(w_dff_B_uKw0ccgk4_2),.clk(gclk));
	jdff dff_B_Z0Qxccvj0_2(.din(w_dff_B_uKw0ccgk4_2),.dout(w_dff_B_Z0Qxccvj0_2),.clk(gclk));
	jdff dff_B_A0kbsgkX3_2(.din(w_dff_B_Z0Qxccvj0_2),.dout(w_dff_B_A0kbsgkX3_2),.clk(gclk));
	jdff dff_B_qXl1i2G03_2(.din(w_dff_B_A0kbsgkX3_2),.dout(w_dff_B_qXl1i2G03_2),.clk(gclk));
	jdff dff_B_xtNOEPbD4_2(.din(w_dff_B_qXl1i2G03_2),.dout(w_dff_B_xtNOEPbD4_2),.clk(gclk));
	jdff dff_B_6iUx3StV5_2(.din(w_dff_B_xtNOEPbD4_2),.dout(w_dff_B_6iUx3StV5_2),.clk(gclk));
	jdff dff_B_kumXx7DD7_2(.din(w_dff_B_6iUx3StV5_2),.dout(w_dff_B_kumXx7DD7_2),.clk(gclk));
	jdff dff_B_cU4ceoFc0_2(.din(w_dff_B_kumXx7DD7_2),.dout(w_dff_B_cU4ceoFc0_2),.clk(gclk));
	jdff dff_B_shnmPZuQ9_2(.din(w_dff_B_cU4ceoFc0_2),.dout(w_dff_B_shnmPZuQ9_2),.clk(gclk));
	jdff dff_B_8xukIEZj5_2(.din(w_dff_B_shnmPZuQ9_2),.dout(w_dff_B_8xukIEZj5_2),.clk(gclk));
	jdff dff_B_zx79VxaU5_2(.din(w_dff_B_8xukIEZj5_2),.dout(w_dff_B_zx79VxaU5_2),.clk(gclk));
	jdff dff_B_BJnagulE2_2(.din(w_dff_B_zx79VxaU5_2),.dout(w_dff_B_BJnagulE2_2),.clk(gclk));
	jdff dff_B_RAPl8noj9_2(.din(w_dff_B_BJnagulE2_2),.dout(w_dff_B_RAPl8noj9_2),.clk(gclk));
	jdff dff_B_RGUU8MWp9_2(.din(w_dff_B_RAPl8noj9_2),.dout(w_dff_B_RGUU8MWp9_2),.clk(gclk));
	jdff dff_B_wGb0rXKg5_2(.din(w_dff_B_RGUU8MWp9_2),.dout(w_dff_B_wGb0rXKg5_2),.clk(gclk));
	jdff dff_B_VaCAp1wr0_2(.din(w_dff_B_wGb0rXKg5_2),.dout(w_dff_B_VaCAp1wr0_2),.clk(gclk));
	jdff dff_B_QG55KrUk7_2(.din(w_dff_B_VaCAp1wr0_2),.dout(w_dff_B_QG55KrUk7_2),.clk(gclk));
	jdff dff_B_NDvpUEeQ2_2(.din(w_dff_B_QG55KrUk7_2),.dout(w_dff_B_NDvpUEeQ2_2),.clk(gclk));
	jdff dff_B_dm8KWOiU1_2(.din(w_dff_B_NDvpUEeQ2_2),.dout(w_dff_B_dm8KWOiU1_2),.clk(gclk));
	jdff dff_B_p4d5zdTR9_2(.din(w_dff_B_dm8KWOiU1_2),.dout(w_dff_B_p4d5zdTR9_2),.clk(gclk));
	jdff dff_B_OBe0MAmH4_2(.din(w_dff_B_p4d5zdTR9_2),.dout(w_dff_B_OBe0MAmH4_2),.clk(gclk));
	jdff dff_B_B2EeaBhy3_2(.din(w_dff_B_OBe0MAmH4_2),.dout(w_dff_B_B2EeaBhy3_2),.clk(gclk));
	jdff dff_B_68Q8aHDQ7_2(.din(w_dff_B_B2EeaBhy3_2),.dout(w_dff_B_68Q8aHDQ7_2),.clk(gclk));
	jdff dff_B_0WmD325C5_2(.din(w_dff_B_68Q8aHDQ7_2),.dout(w_dff_B_0WmD325C5_2),.clk(gclk));
	jdff dff_B_IbqKD7kx4_2(.din(w_dff_B_0WmD325C5_2),.dout(w_dff_B_IbqKD7kx4_2),.clk(gclk));
	jdff dff_B_qK3gEvZR7_2(.din(w_dff_B_IbqKD7kx4_2),.dout(w_dff_B_qK3gEvZR7_2),.clk(gclk));
	jdff dff_B_MWkfWstk4_2(.din(w_dff_B_qK3gEvZR7_2),.dout(w_dff_B_MWkfWstk4_2),.clk(gclk));
	jdff dff_B_FHrD2GwZ3_2(.din(w_dff_B_MWkfWstk4_2),.dout(w_dff_B_FHrD2GwZ3_2),.clk(gclk));
	jdff dff_B_S3idry3O1_2(.din(w_dff_B_FHrD2GwZ3_2),.dout(w_dff_B_S3idry3O1_2),.clk(gclk));
	jdff dff_B_Onv7pv8s0_2(.din(w_dff_B_S3idry3O1_2),.dout(w_dff_B_Onv7pv8s0_2),.clk(gclk));
	jdff dff_B_D8AJXiMT8_2(.din(n1738),.dout(w_dff_B_D8AJXiMT8_2),.clk(gclk));
	jdff dff_B_iuLwvLhL0_1(.din(n1736),.dout(w_dff_B_iuLwvLhL0_1),.clk(gclk));
	jdff dff_B_hWsSLFhh0_2(.din(n1694),.dout(w_dff_B_hWsSLFhh0_2),.clk(gclk));
	jdff dff_B_DnIzzPtW1_2(.din(w_dff_B_hWsSLFhh0_2),.dout(w_dff_B_DnIzzPtW1_2),.clk(gclk));
	jdff dff_B_MAOfJYIF0_2(.din(w_dff_B_DnIzzPtW1_2),.dout(w_dff_B_MAOfJYIF0_2),.clk(gclk));
	jdff dff_B_4PXKLdAN8_2(.din(w_dff_B_MAOfJYIF0_2),.dout(w_dff_B_4PXKLdAN8_2),.clk(gclk));
	jdff dff_B_LelS9Q6e1_2(.din(w_dff_B_4PXKLdAN8_2),.dout(w_dff_B_LelS9Q6e1_2),.clk(gclk));
	jdff dff_B_qlqGLVOQ4_2(.din(w_dff_B_LelS9Q6e1_2),.dout(w_dff_B_qlqGLVOQ4_2),.clk(gclk));
	jdff dff_B_gk81zt5a9_2(.din(w_dff_B_qlqGLVOQ4_2),.dout(w_dff_B_gk81zt5a9_2),.clk(gclk));
	jdff dff_B_DkTaDtrc2_2(.din(w_dff_B_gk81zt5a9_2),.dout(w_dff_B_DkTaDtrc2_2),.clk(gclk));
	jdff dff_B_BjEHUZ0o7_2(.din(w_dff_B_DkTaDtrc2_2),.dout(w_dff_B_BjEHUZ0o7_2),.clk(gclk));
	jdff dff_B_i7LghEmm7_2(.din(w_dff_B_BjEHUZ0o7_2),.dout(w_dff_B_i7LghEmm7_2),.clk(gclk));
	jdff dff_B_rASNtBbA4_2(.din(w_dff_B_i7LghEmm7_2),.dout(w_dff_B_rASNtBbA4_2),.clk(gclk));
	jdff dff_B_OXFzaDa63_2(.din(w_dff_B_rASNtBbA4_2),.dout(w_dff_B_OXFzaDa63_2),.clk(gclk));
	jdff dff_B_LzKClCU40_2(.din(w_dff_B_OXFzaDa63_2),.dout(w_dff_B_LzKClCU40_2),.clk(gclk));
	jdff dff_B_V4hBBEHr7_2(.din(w_dff_B_LzKClCU40_2),.dout(w_dff_B_V4hBBEHr7_2),.clk(gclk));
	jdff dff_B_sTsrNt3r3_2(.din(w_dff_B_V4hBBEHr7_2),.dout(w_dff_B_sTsrNt3r3_2),.clk(gclk));
	jdff dff_B_3fmE2yMf3_2(.din(w_dff_B_sTsrNt3r3_2),.dout(w_dff_B_3fmE2yMf3_2),.clk(gclk));
	jdff dff_B_HHQlUgVJ6_2(.din(w_dff_B_3fmE2yMf3_2),.dout(w_dff_B_HHQlUgVJ6_2),.clk(gclk));
	jdff dff_B_St80496l2_2(.din(w_dff_B_HHQlUgVJ6_2),.dout(w_dff_B_St80496l2_2),.clk(gclk));
	jdff dff_B_N4dfAHcJ7_2(.din(w_dff_B_St80496l2_2),.dout(w_dff_B_N4dfAHcJ7_2),.clk(gclk));
	jdff dff_B_87HrfKX45_2(.din(w_dff_B_N4dfAHcJ7_2),.dout(w_dff_B_87HrfKX45_2),.clk(gclk));
	jdff dff_B_JvZ0hTq43_2(.din(w_dff_B_87HrfKX45_2),.dout(w_dff_B_JvZ0hTq43_2),.clk(gclk));
	jdff dff_B_9JYQMTnW0_2(.din(w_dff_B_JvZ0hTq43_2),.dout(w_dff_B_9JYQMTnW0_2),.clk(gclk));
	jdff dff_B_HxcPrKRJ7_2(.din(w_dff_B_9JYQMTnW0_2),.dout(w_dff_B_HxcPrKRJ7_2),.clk(gclk));
	jdff dff_B_mgRs9CGs9_2(.din(w_dff_B_HxcPrKRJ7_2),.dout(w_dff_B_mgRs9CGs9_2),.clk(gclk));
	jdff dff_B_P9uCtLmh5_2(.din(w_dff_B_mgRs9CGs9_2),.dout(w_dff_B_P9uCtLmh5_2),.clk(gclk));
	jdff dff_B_cf0LEYy75_2(.din(w_dff_B_P9uCtLmh5_2),.dout(w_dff_B_cf0LEYy75_2),.clk(gclk));
	jdff dff_B_6agVIGVX2_2(.din(w_dff_B_cf0LEYy75_2),.dout(w_dff_B_6agVIGVX2_2),.clk(gclk));
	jdff dff_B_Jx1P4F5i3_2(.din(w_dff_B_6agVIGVX2_2),.dout(w_dff_B_Jx1P4F5i3_2),.clk(gclk));
	jdff dff_B_k0fY72Uo3_2(.din(w_dff_B_Jx1P4F5i3_2),.dout(w_dff_B_k0fY72Uo3_2),.clk(gclk));
	jdff dff_B_0i2aVSqO7_2(.din(w_dff_B_k0fY72Uo3_2),.dout(w_dff_B_0i2aVSqO7_2),.clk(gclk));
	jdff dff_B_fDFBxM5M8_2(.din(w_dff_B_0i2aVSqO7_2),.dout(w_dff_B_fDFBxM5M8_2),.clk(gclk));
	jdff dff_B_0P0nXKC87_2(.din(w_dff_B_fDFBxM5M8_2),.dout(w_dff_B_0P0nXKC87_2),.clk(gclk));
	jdff dff_B_OcMrzMJL0_2(.din(w_dff_B_0P0nXKC87_2),.dout(w_dff_B_OcMrzMJL0_2),.clk(gclk));
	jdff dff_B_4dq6X5jt7_2(.din(w_dff_B_OcMrzMJL0_2),.dout(w_dff_B_4dq6X5jt7_2),.clk(gclk));
	jdff dff_B_koax4oEL4_2(.din(w_dff_B_4dq6X5jt7_2),.dout(w_dff_B_koax4oEL4_2),.clk(gclk));
	jdff dff_B_kVKZu0VS8_2(.din(n1697),.dout(w_dff_B_kVKZu0VS8_2),.clk(gclk));
	jdff dff_B_OwlYxgy72_1(.din(n1695),.dout(w_dff_B_OwlYxgy72_1),.clk(gclk));
	jdff dff_B_YMBcjPwl9_2(.din(n1643),.dout(w_dff_B_YMBcjPwl9_2),.clk(gclk));
	jdff dff_B_B8rzKxcG1_2(.din(w_dff_B_YMBcjPwl9_2),.dout(w_dff_B_B8rzKxcG1_2),.clk(gclk));
	jdff dff_B_kcvzjtW91_2(.din(w_dff_B_B8rzKxcG1_2),.dout(w_dff_B_kcvzjtW91_2),.clk(gclk));
	jdff dff_B_NGdXoPSC2_2(.din(w_dff_B_kcvzjtW91_2),.dout(w_dff_B_NGdXoPSC2_2),.clk(gclk));
	jdff dff_B_ARNEuVDF2_2(.din(w_dff_B_NGdXoPSC2_2),.dout(w_dff_B_ARNEuVDF2_2),.clk(gclk));
	jdff dff_B_PNtMEDB15_2(.din(w_dff_B_ARNEuVDF2_2),.dout(w_dff_B_PNtMEDB15_2),.clk(gclk));
	jdff dff_B_ac8QHhHG9_2(.din(w_dff_B_PNtMEDB15_2),.dout(w_dff_B_ac8QHhHG9_2),.clk(gclk));
	jdff dff_B_DenZcyew2_2(.din(w_dff_B_ac8QHhHG9_2),.dout(w_dff_B_DenZcyew2_2),.clk(gclk));
	jdff dff_B_2cmKzP9h9_2(.din(w_dff_B_DenZcyew2_2),.dout(w_dff_B_2cmKzP9h9_2),.clk(gclk));
	jdff dff_B_zpyZy9Pa1_2(.din(w_dff_B_2cmKzP9h9_2),.dout(w_dff_B_zpyZy9Pa1_2),.clk(gclk));
	jdff dff_B_xN4SmyIw9_2(.din(w_dff_B_zpyZy9Pa1_2),.dout(w_dff_B_xN4SmyIw9_2),.clk(gclk));
	jdff dff_B_tQDyDHsC8_2(.din(w_dff_B_xN4SmyIw9_2),.dout(w_dff_B_tQDyDHsC8_2),.clk(gclk));
	jdff dff_B_DX0hPpvt7_2(.din(w_dff_B_tQDyDHsC8_2),.dout(w_dff_B_DX0hPpvt7_2),.clk(gclk));
	jdff dff_B_AI89dD9b4_2(.din(w_dff_B_DX0hPpvt7_2),.dout(w_dff_B_AI89dD9b4_2),.clk(gclk));
	jdff dff_B_VNHZRxGO7_2(.din(w_dff_B_AI89dD9b4_2),.dout(w_dff_B_VNHZRxGO7_2),.clk(gclk));
	jdff dff_B_z73vebUl3_2(.din(w_dff_B_VNHZRxGO7_2),.dout(w_dff_B_z73vebUl3_2),.clk(gclk));
	jdff dff_B_FlR1b3v91_2(.din(w_dff_B_z73vebUl3_2),.dout(w_dff_B_FlR1b3v91_2),.clk(gclk));
	jdff dff_B_C8Iyb30f4_2(.din(w_dff_B_FlR1b3v91_2),.dout(w_dff_B_C8Iyb30f4_2),.clk(gclk));
	jdff dff_B_kRxTDog36_2(.din(w_dff_B_C8Iyb30f4_2),.dout(w_dff_B_kRxTDog36_2),.clk(gclk));
	jdff dff_B_xG2ummhN6_2(.din(w_dff_B_kRxTDog36_2),.dout(w_dff_B_xG2ummhN6_2),.clk(gclk));
	jdff dff_B_MBRnurS83_2(.din(w_dff_B_xG2ummhN6_2),.dout(w_dff_B_MBRnurS83_2),.clk(gclk));
	jdff dff_B_xEkF9KEu3_2(.din(w_dff_B_MBRnurS83_2),.dout(w_dff_B_xEkF9KEu3_2),.clk(gclk));
	jdff dff_B_8sVaR9KL3_2(.din(w_dff_B_xEkF9KEu3_2),.dout(w_dff_B_8sVaR9KL3_2),.clk(gclk));
	jdff dff_B_JPJPO1043_2(.din(w_dff_B_8sVaR9KL3_2),.dout(w_dff_B_JPJPO1043_2),.clk(gclk));
	jdff dff_B_m9RY8Fbk3_2(.din(w_dff_B_JPJPO1043_2),.dout(w_dff_B_m9RY8Fbk3_2),.clk(gclk));
	jdff dff_B_fcggUJ4O9_2(.din(w_dff_B_m9RY8Fbk3_2),.dout(w_dff_B_fcggUJ4O9_2),.clk(gclk));
	jdff dff_B_yMOlkVNp5_2(.din(w_dff_B_fcggUJ4O9_2),.dout(w_dff_B_yMOlkVNp5_2),.clk(gclk));
	jdff dff_B_WWJuFx5f1_2(.din(w_dff_B_yMOlkVNp5_2),.dout(w_dff_B_WWJuFx5f1_2),.clk(gclk));
	jdff dff_B_ZbN0Ldhk4_2(.din(w_dff_B_WWJuFx5f1_2),.dout(w_dff_B_ZbN0Ldhk4_2),.clk(gclk));
	jdff dff_B_SCoxlTjY5_2(.din(w_dff_B_ZbN0Ldhk4_2),.dout(w_dff_B_SCoxlTjY5_2),.clk(gclk));
	jdff dff_B_Eb1LTRxI1_2(.din(w_dff_B_SCoxlTjY5_2),.dout(w_dff_B_Eb1LTRxI1_2),.clk(gclk));
	jdff dff_B_daRlOphW0_2(.din(w_dff_B_Eb1LTRxI1_2),.dout(w_dff_B_daRlOphW0_2),.clk(gclk));
	jdff dff_B_ZpOkK2qv5_2(.din(n1646),.dout(w_dff_B_ZpOkK2qv5_2),.clk(gclk));
	jdff dff_B_1zuIz7yN8_1(.din(n1644),.dout(w_dff_B_1zuIz7yN8_1),.clk(gclk));
	jdff dff_B_Y9x2XN5C0_2(.din(n1586),.dout(w_dff_B_Y9x2XN5C0_2),.clk(gclk));
	jdff dff_B_wNIUAWUZ8_2(.din(w_dff_B_Y9x2XN5C0_2),.dout(w_dff_B_wNIUAWUZ8_2),.clk(gclk));
	jdff dff_B_Xu0OmIFH4_2(.din(w_dff_B_wNIUAWUZ8_2),.dout(w_dff_B_Xu0OmIFH4_2),.clk(gclk));
	jdff dff_B_DoZ7r9cc7_2(.din(w_dff_B_Xu0OmIFH4_2),.dout(w_dff_B_DoZ7r9cc7_2),.clk(gclk));
	jdff dff_B_DaC3ZOD30_2(.din(w_dff_B_DoZ7r9cc7_2),.dout(w_dff_B_DaC3ZOD30_2),.clk(gclk));
	jdff dff_B_paMlMcmN3_2(.din(w_dff_B_DaC3ZOD30_2),.dout(w_dff_B_paMlMcmN3_2),.clk(gclk));
	jdff dff_B_GaWb72g51_2(.din(w_dff_B_paMlMcmN3_2),.dout(w_dff_B_GaWb72g51_2),.clk(gclk));
	jdff dff_B_TQ3OeISQ2_2(.din(w_dff_B_GaWb72g51_2),.dout(w_dff_B_TQ3OeISQ2_2),.clk(gclk));
	jdff dff_B_uyOB9opk5_2(.din(w_dff_B_TQ3OeISQ2_2),.dout(w_dff_B_uyOB9opk5_2),.clk(gclk));
	jdff dff_B_kt6U1X2Q9_2(.din(w_dff_B_uyOB9opk5_2),.dout(w_dff_B_kt6U1X2Q9_2),.clk(gclk));
	jdff dff_B_NkYhfIoO5_2(.din(w_dff_B_kt6U1X2Q9_2),.dout(w_dff_B_NkYhfIoO5_2),.clk(gclk));
	jdff dff_B_1rkvjoJp5_2(.din(w_dff_B_NkYhfIoO5_2),.dout(w_dff_B_1rkvjoJp5_2),.clk(gclk));
	jdff dff_B_2LmFrbWc1_2(.din(w_dff_B_1rkvjoJp5_2),.dout(w_dff_B_2LmFrbWc1_2),.clk(gclk));
	jdff dff_B_4n4reUpB0_2(.din(w_dff_B_2LmFrbWc1_2),.dout(w_dff_B_4n4reUpB0_2),.clk(gclk));
	jdff dff_B_z83Qssm48_2(.din(w_dff_B_4n4reUpB0_2),.dout(w_dff_B_z83Qssm48_2),.clk(gclk));
	jdff dff_B_Z9bjJAQq1_2(.din(w_dff_B_z83Qssm48_2),.dout(w_dff_B_Z9bjJAQq1_2),.clk(gclk));
	jdff dff_B_r1vj7Apr4_2(.din(w_dff_B_Z9bjJAQq1_2),.dout(w_dff_B_r1vj7Apr4_2),.clk(gclk));
	jdff dff_B_Dji2Auff5_2(.din(w_dff_B_r1vj7Apr4_2),.dout(w_dff_B_Dji2Auff5_2),.clk(gclk));
	jdff dff_B_NvckqNtQ5_2(.din(w_dff_B_Dji2Auff5_2),.dout(w_dff_B_NvckqNtQ5_2),.clk(gclk));
	jdff dff_B_TtPObzDc2_2(.din(w_dff_B_NvckqNtQ5_2),.dout(w_dff_B_TtPObzDc2_2),.clk(gclk));
	jdff dff_B_615mHX7N8_2(.din(w_dff_B_TtPObzDc2_2),.dout(w_dff_B_615mHX7N8_2),.clk(gclk));
	jdff dff_B_vDDfV8HK2_2(.din(w_dff_B_615mHX7N8_2),.dout(w_dff_B_vDDfV8HK2_2),.clk(gclk));
	jdff dff_B_UGbJX35k1_2(.din(w_dff_B_vDDfV8HK2_2),.dout(w_dff_B_UGbJX35k1_2),.clk(gclk));
	jdff dff_B_lCaQomBp7_2(.din(w_dff_B_UGbJX35k1_2),.dout(w_dff_B_lCaQomBp7_2),.clk(gclk));
	jdff dff_B_WQZhWyPd8_2(.din(w_dff_B_lCaQomBp7_2),.dout(w_dff_B_WQZhWyPd8_2),.clk(gclk));
	jdff dff_B_TyxjQAWM3_2(.din(w_dff_B_WQZhWyPd8_2),.dout(w_dff_B_TyxjQAWM3_2),.clk(gclk));
	jdff dff_B_GJlJgzFq8_2(.din(w_dff_B_TyxjQAWM3_2),.dout(w_dff_B_GJlJgzFq8_2),.clk(gclk));
	jdff dff_B_mrLY5sBn8_2(.din(w_dff_B_GJlJgzFq8_2),.dout(w_dff_B_mrLY5sBn8_2),.clk(gclk));
	jdff dff_B_mrZXleBf5_2(.din(w_dff_B_mrLY5sBn8_2),.dout(w_dff_B_mrZXleBf5_2),.clk(gclk));
	jdff dff_B_TQ1Z6noW7_2(.din(n1589),.dout(w_dff_B_TQ1Z6noW7_2),.clk(gclk));
	jdff dff_B_t7lINx934_1(.din(n1587),.dout(w_dff_B_t7lINx934_1),.clk(gclk));
	jdff dff_B_BE4QdvDD6_2(.din(n1522),.dout(w_dff_B_BE4QdvDD6_2),.clk(gclk));
	jdff dff_B_niA3mLEb2_2(.din(w_dff_B_BE4QdvDD6_2),.dout(w_dff_B_niA3mLEb2_2),.clk(gclk));
	jdff dff_B_gshMcPLK1_2(.din(w_dff_B_niA3mLEb2_2),.dout(w_dff_B_gshMcPLK1_2),.clk(gclk));
	jdff dff_B_vW6fWiFr4_2(.din(w_dff_B_gshMcPLK1_2),.dout(w_dff_B_vW6fWiFr4_2),.clk(gclk));
	jdff dff_B_phyljEV00_2(.din(w_dff_B_vW6fWiFr4_2),.dout(w_dff_B_phyljEV00_2),.clk(gclk));
	jdff dff_B_WqnUaDZj3_2(.din(w_dff_B_phyljEV00_2),.dout(w_dff_B_WqnUaDZj3_2),.clk(gclk));
	jdff dff_B_jViUbaNz1_2(.din(w_dff_B_WqnUaDZj3_2),.dout(w_dff_B_jViUbaNz1_2),.clk(gclk));
	jdff dff_B_MZAUlxvx0_2(.din(w_dff_B_jViUbaNz1_2),.dout(w_dff_B_MZAUlxvx0_2),.clk(gclk));
	jdff dff_B_V8xbDkFG8_2(.din(w_dff_B_MZAUlxvx0_2),.dout(w_dff_B_V8xbDkFG8_2),.clk(gclk));
	jdff dff_B_YEjHdRFj9_2(.din(w_dff_B_V8xbDkFG8_2),.dout(w_dff_B_YEjHdRFj9_2),.clk(gclk));
	jdff dff_B_Sx14C7uq7_2(.din(w_dff_B_YEjHdRFj9_2),.dout(w_dff_B_Sx14C7uq7_2),.clk(gclk));
	jdff dff_B_yWqDNBmV3_2(.din(w_dff_B_Sx14C7uq7_2),.dout(w_dff_B_yWqDNBmV3_2),.clk(gclk));
	jdff dff_B_kgsShTQa1_2(.din(w_dff_B_yWqDNBmV3_2),.dout(w_dff_B_kgsShTQa1_2),.clk(gclk));
	jdff dff_B_AS5IVjcG7_2(.din(w_dff_B_kgsShTQa1_2),.dout(w_dff_B_AS5IVjcG7_2),.clk(gclk));
	jdff dff_B_FDJxEl4k1_2(.din(w_dff_B_AS5IVjcG7_2),.dout(w_dff_B_FDJxEl4k1_2),.clk(gclk));
	jdff dff_B_ySZUNYfa5_2(.din(w_dff_B_FDJxEl4k1_2),.dout(w_dff_B_ySZUNYfa5_2),.clk(gclk));
	jdff dff_B_N1OZ2zrm9_2(.din(w_dff_B_ySZUNYfa5_2),.dout(w_dff_B_N1OZ2zrm9_2),.clk(gclk));
	jdff dff_B_AYiIzIG12_2(.din(w_dff_B_N1OZ2zrm9_2),.dout(w_dff_B_AYiIzIG12_2),.clk(gclk));
	jdff dff_B_QrL7BOrv2_2(.din(w_dff_B_AYiIzIG12_2),.dout(w_dff_B_QrL7BOrv2_2),.clk(gclk));
	jdff dff_B_9yzo2Y6g2_2(.din(w_dff_B_QrL7BOrv2_2),.dout(w_dff_B_9yzo2Y6g2_2),.clk(gclk));
	jdff dff_B_UtyAaVIM3_2(.din(w_dff_B_9yzo2Y6g2_2),.dout(w_dff_B_UtyAaVIM3_2),.clk(gclk));
	jdff dff_B_i1BQQSYZ2_2(.din(w_dff_B_UtyAaVIM3_2),.dout(w_dff_B_i1BQQSYZ2_2),.clk(gclk));
	jdff dff_B_CdAax9ul5_2(.din(w_dff_B_i1BQQSYZ2_2),.dout(w_dff_B_CdAax9ul5_2),.clk(gclk));
	jdff dff_B_MxQTAqAG3_2(.din(w_dff_B_CdAax9ul5_2),.dout(w_dff_B_MxQTAqAG3_2),.clk(gclk));
	jdff dff_B_9iXyJA0Q8_2(.din(w_dff_B_MxQTAqAG3_2),.dout(w_dff_B_9iXyJA0Q8_2),.clk(gclk));
	jdff dff_B_SL4sG0kr9_2(.din(w_dff_B_9iXyJA0Q8_2),.dout(w_dff_B_SL4sG0kr9_2),.clk(gclk));
	jdff dff_B_JTtRBhye0_2(.din(n1525),.dout(w_dff_B_JTtRBhye0_2),.clk(gclk));
	jdff dff_B_6dviGXV86_1(.din(n1523),.dout(w_dff_B_6dviGXV86_1),.clk(gclk));
	jdff dff_B_ndH1q0i26_2(.din(n1451),.dout(w_dff_B_ndH1q0i26_2),.clk(gclk));
	jdff dff_B_PVQabe368_2(.din(w_dff_B_ndH1q0i26_2),.dout(w_dff_B_PVQabe368_2),.clk(gclk));
	jdff dff_B_UGg0x5Dn0_2(.din(w_dff_B_PVQabe368_2),.dout(w_dff_B_UGg0x5Dn0_2),.clk(gclk));
	jdff dff_B_CoSon9c16_2(.din(w_dff_B_UGg0x5Dn0_2),.dout(w_dff_B_CoSon9c16_2),.clk(gclk));
	jdff dff_B_g1BDn8Lx0_2(.din(w_dff_B_CoSon9c16_2),.dout(w_dff_B_g1BDn8Lx0_2),.clk(gclk));
	jdff dff_B_1z3AD6Fn0_2(.din(w_dff_B_g1BDn8Lx0_2),.dout(w_dff_B_1z3AD6Fn0_2),.clk(gclk));
	jdff dff_B_hUymP6L81_2(.din(w_dff_B_1z3AD6Fn0_2),.dout(w_dff_B_hUymP6L81_2),.clk(gclk));
	jdff dff_B_EZTkmud71_2(.din(w_dff_B_hUymP6L81_2),.dout(w_dff_B_EZTkmud71_2),.clk(gclk));
	jdff dff_B_NktW4f2W6_2(.din(w_dff_B_EZTkmud71_2),.dout(w_dff_B_NktW4f2W6_2),.clk(gclk));
	jdff dff_B_OOseTLPn8_2(.din(w_dff_B_NktW4f2W6_2),.dout(w_dff_B_OOseTLPn8_2),.clk(gclk));
	jdff dff_B_Eq5VuKmS1_2(.din(w_dff_B_OOseTLPn8_2),.dout(w_dff_B_Eq5VuKmS1_2),.clk(gclk));
	jdff dff_B_UNQtDASk7_2(.din(w_dff_B_Eq5VuKmS1_2),.dout(w_dff_B_UNQtDASk7_2),.clk(gclk));
	jdff dff_B_dXBavHkH6_2(.din(w_dff_B_UNQtDASk7_2),.dout(w_dff_B_dXBavHkH6_2),.clk(gclk));
	jdff dff_B_AnI7U8vz6_2(.din(w_dff_B_dXBavHkH6_2),.dout(w_dff_B_AnI7U8vz6_2),.clk(gclk));
	jdff dff_B_A28RxnFs2_2(.din(w_dff_B_AnI7U8vz6_2),.dout(w_dff_B_A28RxnFs2_2),.clk(gclk));
	jdff dff_B_tYL0F2Yq5_2(.din(w_dff_B_A28RxnFs2_2),.dout(w_dff_B_tYL0F2Yq5_2),.clk(gclk));
	jdff dff_B_VqemReL51_2(.din(w_dff_B_tYL0F2Yq5_2),.dout(w_dff_B_VqemReL51_2),.clk(gclk));
	jdff dff_B_FzuQiHV79_2(.din(w_dff_B_VqemReL51_2),.dout(w_dff_B_FzuQiHV79_2),.clk(gclk));
	jdff dff_B_2qdNOR3u9_2(.din(w_dff_B_FzuQiHV79_2),.dout(w_dff_B_2qdNOR3u9_2),.clk(gclk));
	jdff dff_B_92o2sBoo8_2(.din(w_dff_B_2qdNOR3u9_2),.dout(w_dff_B_92o2sBoo8_2),.clk(gclk));
	jdff dff_B_T9MeuH202_2(.din(w_dff_B_92o2sBoo8_2),.dout(w_dff_B_T9MeuH202_2),.clk(gclk));
	jdff dff_B_kViNAkG78_2(.din(w_dff_B_T9MeuH202_2),.dout(w_dff_B_kViNAkG78_2),.clk(gclk));
	jdff dff_B_jMrDNSe89_2(.din(w_dff_B_kViNAkG78_2),.dout(w_dff_B_jMrDNSe89_2),.clk(gclk));
	jdff dff_B_2McmDv8G7_2(.din(n1454),.dout(w_dff_B_2McmDv8G7_2),.clk(gclk));
	jdff dff_B_sh0dxksO2_1(.din(n1452),.dout(w_dff_B_sh0dxksO2_1),.clk(gclk));
	jdff dff_B_hC7BbIqV6_2(.din(n1373),.dout(w_dff_B_hC7BbIqV6_2),.clk(gclk));
	jdff dff_B_oYRgShH11_2(.din(w_dff_B_hC7BbIqV6_2),.dout(w_dff_B_oYRgShH11_2),.clk(gclk));
	jdff dff_B_ZlJNZeT99_2(.din(w_dff_B_oYRgShH11_2),.dout(w_dff_B_ZlJNZeT99_2),.clk(gclk));
	jdff dff_B_qL4Ht7TW1_2(.din(w_dff_B_ZlJNZeT99_2),.dout(w_dff_B_qL4Ht7TW1_2),.clk(gclk));
	jdff dff_B_EW52QgG49_2(.din(w_dff_B_qL4Ht7TW1_2),.dout(w_dff_B_EW52QgG49_2),.clk(gclk));
	jdff dff_B_1LHCHdbr8_2(.din(w_dff_B_EW52QgG49_2),.dout(w_dff_B_1LHCHdbr8_2),.clk(gclk));
	jdff dff_B_4OjnTwQM1_2(.din(w_dff_B_1LHCHdbr8_2),.dout(w_dff_B_4OjnTwQM1_2),.clk(gclk));
	jdff dff_B_6aZBglVu5_2(.din(w_dff_B_4OjnTwQM1_2),.dout(w_dff_B_6aZBglVu5_2),.clk(gclk));
	jdff dff_B_QUGtxAtR7_2(.din(w_dff_B_6aZBglVu5_2),.dout(w_dff_B_QUGtxAtR7_2),.clk(gclk));
	jdff dff_B_cxL7swVY5_2(.din(w_dff_B_QUGtxAtR7_2),.dout(w_dff_B_cxL7swVY5_2),.clk(gclk));
	jdff dff_B_OaGEaaHd2_2(.din(w_dff_B_cxL7swVY5_2),.dout(w_dff_B_OaGEaaHd2_2),.clk(gclk));
	jdff dff_B_l6lFYMIb9_2(.din(w_dff_B_OaGEaaHd2_2),.dout(w_dff_B_l6lFYMIb9_2),.clk(gclk));
	jdff dff_B_8Lbq6cW45_2(.din(w_dff_B_l6lFYMIb9_2),.dout(w_dff_B_8Lbq6cW45_2),.clk(gclk));
	jdff dff_B_oXRt8b9B3_2(.din(w_dff_B_8Lbq6cW45_2),.dout(w_dff_B_oXRt8b9B3_2),.clk(gclk));
	jdff dff_B_sKIJYoAd3_2(.din(w_dff_B_oXRt8b9B3_2),.dout(w_dff_B_sKIJYoAd3_2),.clk(gclk));
	jdff dff_B_xL29oZzT0_2(.din(w_dff_B_sKIJYoAd3_2),.dout(w_dff_B_xL29oZzT0_2),.clk(gclk));
	jdff dff_B_vSw9KwCM8_2(.din(w_dff_B_xL29oZzT0_2),.dout(w_dff_B_vSw9KwCM8_2),.clk(gclk));
	jdff dff_B_nlQCxk901_2(.din(w_dff_B_vSw9KwCM8_2),.dout(w_dff_B_nlQCxk901_2),.clk(gclk));
	jdff dff_B_lwUCygxZ2_2(.din(w_dff_B_nlQCxk901_2),.dout(w_dff_B_lwUCygxZ2_2),.clk(gclk));
	jdff dff_B_iQXQbdJt5_2(.din(w_dff_B_lwUCygxZ2_2),.dout(w_dff_B_iQXQbdJt5_2),.clk(gclk));
	jdff dff_B_A0i2702a4_2(.din(n1376),.dout(w_dff_B_A0i2702a4_2),.clk(gclk));
	jdff dff_B_INKymOYR8_1(.din(n1374),.dout(w_dff_B_INKymOYR8_1),.clk(gclk));
	jdff dff_B_FTtdPVNL9_2(.din(n1288),.dout(w_dff_B_FTtdPVNL9_2),.clk(gclk));
	jdff dff_B_SW6PhlFB7_2(.din(w_dff_B_FTtdPVNL9_2),.dout(w_dff_B_SW6PhlFB7_2),.clk(gclk));
	jdff dff_B_YgO8e70f1_2(.din(w_dff_B_SW6PhlFB7_2),.dout(w_dff_B_YgO8e70f1_2),.clk(gclk));
	jdff dff_B_onAbcYUi9_2(.din(w_dff_B_YgO8e70f1_2),.dout(w_dff_B_onAbcYUi9_2),.clk(gclk));
	jdff dff_B_n3B9ZFsg5_2(.din(w_dff_B_onAbcYUi9_2),.dout(w_dff_B_n3B9ZFsg5_2),.clk(gclk));
	jdff dff_B_vp9uWi3d5_2(.din(w_dff_B_n3B9ZFsg5_2),.dout(w_dff_B_vp9uWi3d5_2),.clk(gclk));
	jdff dff_B_vYbHpcV62_2(.din(w_dff_B_vp9uWi3d5_2),.dout(w_dff_B_vYbHpcV62_2),.clk(gclk));
	jdff dff_B_4abRs4b61_2(.din(w_dff_B_vYbHpcV62_2),.dout(w_dff_B_4abRs4b61_2),.clk(gclk));
	jdff dff_B_gOhZxzpu8_2(.din(w_dff_B_4abRs4b61_2),.dout(w_dff_B_gOhZxzpu8_2),.clk(gclk));
	jdff dff_B_N0AxYhOr4_2(.din(w_dff_B_gOhZxzpu8_2),.dout(w_dff_B_N0AxYhOr4_2),.clk(gclk));
	jdff dff_B_AzAl7yhO4_2(.din(w_dff_B_N0AxYhOr4_2),.dout(w_dff_B_AzAl7yhO4_2),.clk(gclk));
	jdff dff_B_M9jz9D8i7_2(.din(w_dff_B_AzAl7yhO4_2),.dout(w_dff_B_M9jz9D8i7_2),.clk(gclk));
	jdff dff_B_okAosbHv2_2(.din(w_dff_B_M9jz9D8i7_2),.dout(w_dff_B_okAosbHv2_2),.clk(gclk));
	jdff dff_B_7dBtRMgy3_2(.din(w_dff_B_okAosbHv2_2),.dout(w_dff_B_7dBtRMgy3_2),.clk(gclk));
	jdff dff_B_JcemjKhx5_2(.din(w_dff_B_7dBtRMgy3_2),.dout(w_dff_B_JcemjKhx5_2),.clk(gclk));
	jdff dff_B_CRpi4ucq3_2(.din(w_dff_B_JcemjKhx5_2),.dout(w_dff_B_CRpi4ucq3_2),.clk(gclk));
	jdff dff_B_cVNuB1795_2(.din(w_dff_B_CRpi4ucq3_2),.dout(w_dff_B_cVNuB1795_2),.clk(gclk));
	jdff dff_B_Lbwdgh9C9_2(.din(n1291),.dout(w_dff_B_Lbwdgh9C9_2),.clk(gclk));
	jdff dff_B_1n21AahF4_1(.din(n1289),.dout(w_dff_B_1n21AahF4_1),.clk(gclk));
	jdff dff_B_wA9s5U9U5_2(.din(n1198),.dout(w_dff_B_wA9s5U9U5_2),.clk(gclk));
	jdff dff_B_VIomQFwF3_2(.din(w_dff_B_wA9s5U9U5_2),.dout(w_dff_B_VIomQFwF3_2),.clk(gclk));
	jdff dff_B_eiPr1zSx8_2(.din(w_dff_B_VIomQFwF3_2),.dout(w_dff_B_eiPr1zSx8_2),.clk(gclk));
	jdff dff_B_6W9kCZei4_2(.din(w_dff_B_eiPr1zSx8_2),.dout(w_dff_B_6W9kCZei4_2),.clk(gclk));
	jdff dff_B_FNUWosxc9_2(.din(w_dff_B_6W9kCZei4_2),.dout(w_dff_B_FNUWosxc9_2),.clk(gclk));
	jdff dff_B_OVy8mKHP4_2(.din(w_dff_B_FNUWosxc9_2),.dout(w_dff_B_OVy8mKHP4_2),.clk(gclk));
	jdff dff_B_I23sPtR88_2(.din(w_dff_B_OVy8mKHP4_2),.dout(w_dff_B_I23sPtR88_2),.clk(gclk));
	jdff dff_B_UHnAMCwM8_2(.din(w_dff_B_I23sPtR88_2),.dout(w_dff_B_UHnAMCwM8_2),.clk(gclk));
	jdff dff_B_cItW43000_2(.din(w_dff_B_UHnAMCwM8_2),.dout(w_dff_B_cItW43000_2),.clk(gclk));
	jdff dff_B_bophiV9U5_2(.din(w_dff_B_cItW43000_2),.dout(w_dff_B_bophiV9U5_2),.clk(gclk));
	jdff dff_B_C0lRuRsc7_2(.din(w_dff_B_bophiV9U5_2),.dout(w_dff_B_C0lRuRsc7_2),.clk(gclk));
	jdff dff_B_6PEiuxw30_2(.din(w_dff_B_C0lRuRsc7_2),.dout(w_dff_B_6PEiuxw30_2),.clk(gclk));
	jdff dff_B_63ir5bPq7_2(.din(w_dff_B_6PEiuxw30_2),.dout(w_dff_B_63ir5bPq7_2),.clk(gclk));
	jdff dff_B_fCsW9NnO7_2(.din(w_dff_B_63ir5bPq7_2),.dout(w_dff_B_fCsW9NnO7_2),.clk(gclk));
	jdff dff_B_xUKLDhg11_2(.din(n1201),.dout(w_dff_B_xUKLDhg11_2),.clk(gclk));
	jdff dff_B_ztUuxrZa4_1(.din(n1199),.dout(w_dff_B_ztUuxrZa4_1),.clk(gclk));
	jdff dff_B_SOjC0u682_2(.din(n1094),.dout(w_dff_B_SOjC0u682_2),.clk(gclk));
	jdff dff_B_ZRFRRR0f1_2(.din(w_dff_B_SOjC0u682_2),.dout(w_dff_B_ZRFRRR0f1_2),.clk(gclk));
	jdff dff_B_Lj2Y2oRF3_2(.din(w_dff_B_ZRFRRR0f1_2),.dout(w_dff_B_Lj2Y2oRF3_2),.clk(gclk));
	jdff dff_B_fE61N04S1_2(.din(w_dff_B_Lj2Y2oRF3_2),.dout(w_dff_B_fE61N04S1_2),.clk(gclk));
	jdff dff_B_64dfNbLk6_2(.din(w_dff_B_fE61N04S1_2),.dout(w_dff_B_64dfNbLk6_2),.clk(gclk));
	jdff dff_B_wlaoX3Vr8_2(.din(w_dff_B_64dfNbLk6_2),.dout(w_dff_B_wlaoX3Vr8_2),.clk(gclk));
	jdff dff_B_dfIJjtkb1_2(.din(w_dff_B_wlaoX3Vr8_2),.dout(w_dff_B_dfIJjtkb1_2),.clk(gclk));
	jdff dff_B_tdHgasEH1_2(.din(w_dff_B_dfIJjtkb1_2),.dout(w_dff_B_tdHgasEH1_2),.clk(gclk));
	jdff dff_B_FuOHYAuB3_2(.din(w_dff_B_tdHgasEH1_2),.dout(w_dff_B_FuOHYAuB3_2),.clk(gclk));
	jdff dff_B_BrurOUzU1_2(.din(w_dff_B_FuOHYAuB3_2),.dout(w_dff_B_BrurOUzU1_2),.clk(gclk));
	jdff dff_B_dnvH4RRW9_2(.din(w_dff_B_BrurOUzU1_2),.dout(w_dff_B_dnvH4RRW9_2),.clk(gclk));
	jdff dff_B_bqJrps8C6_2(.din(n1097),.dout(w_dff_B_bqJrps8C6_2),.clk(gclk));
	jdff dff_B_CaNGttoo6_1(.din(n1095),.dout(w_dff_B_CaNGttoo6_1),.clk(gclk));
	jdff dff_B_AhgYcDTj0_2(.din(n996),.dout(w_dff_B_AhgYcDTj0_2),.clk(gclk));
	jdff dff_B_rWqLJzx34_2(.din(w_dff_B_AhgYcDTj0_2),.dout(w_dff_B_rWqLJzx34_2),.clk(gclk));
	jdff dff_B_bVPYrA530_2(.din(w_dff_B_rWqLJzx34_2),.dout(w_dff_B_bVPYrA530_2),.clk(gclk));
	jdff dff_B_HrkcjwoK6_2(.din(w_dff_B_bVPYrA530_2),.dout(w_dff_B_HrkcjwoK6_2),.clk(gclk));
	jdff dff_B_NJAO925O7_2(.din(w_dff_B_HrkcjwoK6_2),.dout(w_dff_B_NJAO925O7_2),.clk(gclk));
	jdff dff_B_GLmoDkf79_2(.din(w_dff_B_NJAO925O7_2),.dout(w_dff_B_GLmoDkf79_2),.clk(gclk));
	jdff dff_B_eK7IfPZD4_2(.din(w_dff_B_GLmoDkf79_2),.dout(w_dff_B_eK7IfPZD4_2),.clk(gclk));
	jdff dff_B_ixfXDMSX9_2(.din(w_dff_B_eK7IfPZD4_2),.dout(w_dff_B_ixfXDMSX9_2),.clk(gclk));
	jdff dff_B_VArijCD09_1(.din(n997),.dout(w_dff_B_VArijCD09_1),.clk(gclk));
	jdff dff_B_0stsqYTI2_2(.din(n891),.dout(w_dff_B_0stsqYTI2_2),.clk(gclk));
	jdff dff_B_LsfBhqdJ8_2(.din(w_dff_B_0stsqYTI2_2),.dout(w_dff_B_LsfBhqdJ8_2),.clk(gclk));
	jdff dff_B_IijG6F663_2(.din(w_dff_B_LsfBhqdJ8_2),.dout(w_dff_B_IijG6F663_2),.clk(gclk));
	jdff dff_B_gKXg3xrd9_2(.din(w_dff_B_IijG6F663_2),.dout(w_dff_B_gKXg3xrd9_2),.clk(gclk));
	jdff dff_B_ytyWzPSK7_2(.din(w_dff_B_gKXg3xrd9_2),.dout(w_dff_B_ytyWzPSK7_2),.clk(gclk));
	jdff dff_B_hzNvwo292_2(.din(w_dff_B_ytyWzPSK7_2),.dout(w_dff_B_hzNvwo292_2),.clk(gclk));
	jdff dff_B_E2ffu9kh8_2(.din(n907),.dout(w_dff_B_E2ffu9kh8_2),.clk(gclk));
	jdff dff_B_kSwT1ifs9_1(.din(n892),.dout(w_dff_B_kSwT1ifs9_1),.clk(gclk));
	jdff dff_B_P3tf2sQs7_1(.din(w_dff_B_kSwT1ifs9_1),.dout(w_dff_B_P3tf2sQs7_1),.clk(gclk));
	jdff dff_B_VtnTitoD4_1(.din(w_dff_B_P3tf2sQs7_1),.dout(w_dff_B_VtnTitoD4_1),.clk(gclk));
	jdff dff_B_VI7ITJyG6_1(.din(w_dff_B_VtnTitoD4_1),.dout(w_dff_B_VI7ITJyG6_1),.clk(gclk));
	jdff dff_B_LuvGROLa3_0(.din(n801),.dout(w_dff_B_LuvGROLa3_0),.clk(gclk));
	jdff dff_A_CUC1p7iX4_0(.dout(w_n800_0[0]),.din(w_dff_A_CUC1p7iX4_0),.clk(gclk));
	jdff dff_A_BmmRQH6Y3_0(.dout(w_dff_A_CUC1p7iX4_0),.din(w_dff_A_BmmRQH6Y3_0),.clk(gclk));
	jdff dff_B_Qoe4saXY8_1(.din(n794),.dout(w_dff_B_Qoe4saXY8_1),.clk(gclk));
	jdff dff_B_3R5BpVwG3_1(.din(w_dff_B_Qoe4saXY8_1),.dout(w_dff_B_3R5BpVwG3_1),.clk(gclk));
	jdff dff_A_rwZL9Mh59_0(.dout(w_n698_0[0]),.din(w_dff_A_rwZL9Mh59_0),.clk(gclk));
	jdff dff_A_gPAIF4546_1(.dout(w_n698_0[1]),.din(w_dff_A_gPAIF4546_1),.clk(gclk));
	jdff dff_A_MD2z5eFk2_1(.dout(w_dff_A_gPAIF4546_1),.din(w_dff_A_MD2z5eFk2_1),.clk(gclk));
	jdff dff_A_h7Ops2wC3_1(.dout(w_n792_0[1]),.din(w_dff_A_h7Ops2wC3_1),.clk(gclk));
	jdff dff_A_IXjrD1I14_1(.dout(w_dff_A_h7Ops2wC3_1),.din(w_dff_A_IXjrD1I14_1),.clk(gclk));
	jdff dff_A_Ot93eFkq0_1(.dout(w_dff_A_IXjrD1I14_1),.din(w_dff_A_Ot93eFkq0_1),.clk(gclk));
	jdff dff_A_5nlEOUCZ1_1(.dout(w_dff_A_Ot93eFkq0_1),.din(w_dff_A_5nlEOUCZ1_1),.clk(gclk));
	jdff dff_B_6dBjoyOm3_1(.din(n1843),.dout(w_dff_B_6dBjoyOm3_1),.clk(gclk));
	jdff dff_B_aM5YUJHk4_1(.din(n1830),.dout(w_dff_B_aM5YUJHk4_1),.clk(gclk));
	jdff dff_B_SGXXBPc45_1(.din(w_dff_B_aM5YUJHk4_1),.dout(w_dff_B_SGXXBPc45_1),.clk(gclk));
	jdff dff_B_BcDV6mNw2_2(.din(n1829),.dout(w_dff_B_BcDV6mNw2_2),.clk(gclk));
	jdff dff_B_1bGpGl5T7_2(.din(w_dff_B_BcDV6mNw2_2),.dout(w_dff_B_1bGpGl5T7_2),.clk(gclk));
	jdff dff_B_JnPmFYrf7_2(.din(w_dff_B_1bGpGl5T7_2),.dout(w_dff_B_JnPmFYrf7_2),.clk(gclk));
	jdff dff_B_ropxEmUA2_2(.din(w_dff_B_JnPmFYrf7_2),.dout(w_dff_B_ropxEmUA2_2),.clk(gclk));
	jdff dff_B_2OdIL9367_2(.din(w_dff_B_ropxEmUA2_2),.dout(w_dff_B_2OdIL9367_2),.clk(gclk));
	jdff dff_B_d6B8937O8_2(.din(w_dff_B_2OdIL9367_2),.dout(w_dff_B_d6B8937O8_2),.clk(gclk));
	jdff dff_B_vKfDsliz8_2(.din(w_dff_B_d6B8937O8_2),.dout(w_dff_B_vKfDsliz8_2),.clk(gclk));
	jdff dff_B_XcEDky1r8_2(.din(w_dff_B_vKfDsliz8_2),.dout(w_dff_B_XcEDky1r8_2),.clk(gclk));
	jdff dff_B_D6fCJt7M3_2(.din(w_dff_B_XcEDky1r8_2),.dout(w_dff_B_D6fCJt7M3_2),.clk(gclk));
	jdff dff_B_mQNvpyys1_2(.din(w_dff_B_D6fCJt7M3_2),.dout(w_dff_B_mQNvpyys1_2),.clk(gclk));
	jdff dff_B_T45uRn0Q2_2(.din(w_dff_B_mQNvpyys1_2),.dout(w_dff_B_T45uRn0Q2_2),.clk(gclk));
	jdff dff_B_rVZYlN1W7_2(.din(w_dff_B_T45uRn0Q2_2),.dout(w_dff_B_rVZYlN1W7_2),.clk(gclk));
	jdff dff_B_bKvcE4Fa9_2(.din(w_dff_B_rVZYlN1W7_2),.dout(w_dff_B_bKvcE4Fa9_2),.clk(gclk));
	jdff dff_B_GC62llFU5_2(.din(w_dff_B_bKvcE4Fa9_2),.dout(w_dff_B_GC62llFU5_2),.clk(gclk));
	jdff dff_B_6GOFvHpE6_2(.din(w_dff_B_GC62llFU5_2),.dout(w_dff_B_6GOFvHpE6_2),.clk(gclk));
	jdff dff_B_i5uokXZK0_2(.din(w_dff_B_6GOFvHpE6_2),.dout(w_dff_B_i5uokXZK0_2),.clk(gclk));
	jdff dff_B_kaD8yBEQ8_2(.din(w_dff_B_i5uokXZK0_2),.dout(w_dff_B_kaD8yBEQ8_2),.clk(gclk));
	jdff dff_B_piSWNuxY6_2(.din(w_dff_B_kaD8yBEQ8_2),.dout(w_dff_B_piSWNuxY6_2),.clk(gclk));
	jdff dff_B_oFjfjcPQ5_2(.din(w_dff_B_piSWNuxY6_2),.dout(w_dff_B_oFjfjcPQ5_2),.clk(gclk));
	jdff dff_B_XIgxF0Qb7_2(.din(w_dff_B_oFjfjcPQ5_2),.dout(w_dff_B_XIgxF0Qb7_2),.clk(gclk));
	jdff dff_B_ZdpmQgW77_2(.din(w_dff_B_XIgxF0Qb7_2),.dout(w_dff_B_ZdpmQgW77_2),.clk(gclk));
	jdff dff_B_VxsFvM9j3_2(.din(w_dff_B_ZdpmQgW77_2),.dout(w_dff_B_VxsFvM9j3_2),.clk(gclk));
	jdff dff_B_uIshidnJ9_2(.din(w_dff_B_VxsFvM9j3_2),.dout(w_dff_B_uIshidnJ9_2),.clk(gclk));
	jdff dff_B_6EoNLDxg7_2(.din(w_dff_B_uIshidnJ9_2),.dout(w_dff_B_6EoNLDxg7_2),.clk(gclk));
	jdff dff_B_itKKYmfu5_2(.din(w_dff_B_6EoNLDxg7_2),.dout(w_dff_B_itKKYmfu5_2),.clk(gclk));
	jdff dff_B_26b8Wul84_2(.din(w_dff_B_itKKYmfu5_2),.dout(w_dff_B_26b8Wul84_2),.clk(gclk));
	jdff dff_B_6fE9XqV78_2(.din(w_dff_B_26b8Wul84_2),.dout(w_dff_B_6fE9XqV78_2),.clk(gclk));
	jdff dff_B_YvjkNsXh7_2(.din(w_dff_B_6fE9XqV78_2),.dout(w_dff_B_YvjkNsXh7_2),.clk(gclk));
	jdff dff_B_P5Ytl9pq7_2(.din(w_dff_B_YvjkNsXh7_2),.dout(w_dff_B_P5Ytl9pq7_2),.clk(gclk));
	jdff dff_B_49fqIaC37_2(.din(w_dff_B_P5Ytl9pq7_2),.dout(w_dff_B_49fqIaC37_2),.clk(gclk));
	jdff dff_B_xwUtf7Xf2_2(.din(w_dff_B_49fqIaC37_2),.dout(w_dff_B_xwUtf7Xf2_2),.clk(gclk));
	jdff dff_B_IA96D6sB8_2(.din(w_dff_B_xwUtf7Xf2_2),.dout(w_dff_B_IA96D6sB8_2),.clk(gclk));
	jdff dff_B_VTBg1lRU0_2(.din(w_dff_B_IA96D6sB8_2),.dout(w_dff_B_VTBg1lRU0_2),.clk(gclk));
	jdff dff_B_JvHpUeeM8_2(.din(w_dff_B_VTBg1lRU0_2),.dout(w_dff_B_JvHpUeeM8_2),.clk(gclk));
	jdff dff_B_zCecaY1t8_2(.din(w_dff_B_JvHpUeeM8_2),.dout(w_dff_B_zCecaY1t8_2),.clk(gclk));
	jdff dff_B_YFnOXOHD5_2(.din(w_dff_B_zCecaY1t8_2),.dout(w_dff_B_YFnOXOHD5_2),.clk(gclk));
	jdff dff_B_H9hyc7C43_2(.din(w_dff_B_YFnOXOHD5_2),.dout(w_dff_B_H9hyc7C43_2),.clk(gclk));
	jdff dff_B_hRj2FXJl2_2(.din(w_dff_B_H9hyc7C43_2),.dout(w_dff_B_hRj2FXJl2_2),.clk(gclk));
	jdff dff_B_6tLBjBwn8_2(.din(w_dff_B_hRj2FXJl2_2),.dout(w_dff_B_6tLBjBwn8_2),.clk(gclk));
	jdff dff_B_SBglLqPa8_2(.din(w_dff_B_6tLBjBwn8_2),.dout(w_dff_B_SBglLqPa8_2),.clk(gclk));
	jdff dff_B_gBHmUP9A7_2(.din(w_dff_B_SBglLqPa8_2),.dout(w_dff_B_gBHmUP9A7_2),.clk(gclk));
	jdff dff_B_NK1gJBzJ7_2(.din(w_dff_B_gBHmUP9A7_2),.dout(w_dff_B_NK1gJBzJ7_2),.clk(gclk));
	jdff dff_B_TMxCXRkN4_2(.din(n1828),.dout(w_dff_B_TMxCXRkN4_2),.clk(gclk));
	jdff dff_B_4Fb7TyHm6_2(.din(w_dff_B_TMxCXRkN4_2),.dout(w_dff_B_4Fb7TyHm6_2),.clk(gclk));
	jdff dff_B_4wxreOQc8_2(.din(w_dff_B_4Fb7TyHm6_2),.dout(w_dff_B_4wxreOQc8_2),.clk(gclk));
	jdff dff_B_W0A5pr7J2_2(.din(w_dff_B_4wxreOQc8_2),.dout(w_dff_B_W0A5pr7J2_2),.clk(gclk));
	jdff dff_B_iMa9E4bR5_2(.din(w_dff_B_W0A5pr7J2_2),.dout(w_dff_B_iMa9E4bR5_2),.clk(gclk));
	jdff dff_B_pRCzIX9F5_2(.din(w_dff_B_iMa9E4bR5_2),.dout(w_dff_B_pRCzIX9F5_2),.clk(gclk));
	jdff dff_B_7Xf3GiM45_2(.din(w_dff_B_pRCzIX9F5_2),.dout(w_dff_B_7Xf3GiM45_2),.clk(gclk));
	jdff dff_B_HebX0F8X0_2(.din(w_dff_B_7Xf3GiM45_2),.dout(w_dff_B_HebX0F8X0_2),.clk(gclk));
	jdff dff_B_nMM7Ej3k3_2(.din(w_dff_B_HebX0F8X0_2),.dout(w_dff_B_nMM7Ej3k3_2),.clk(gclk));
	jdff dff_B_HtVg4BPT0_2(.din(w_dff_B_nMM7Ej3k3_2),.dout(w_dff_B_HtVg4BPT0_2),.clk(gclk));
	jdff dff_B_R35mousA7_2(.din(w_dff_B_HtVg4BPT0_2),.dout(w_dff_B_R35mousA7_2),.clk(gclk));
	jdff dff_B_ZYuOm7OY3_2(.din(w_dff_B_R35mousA7_2),.dout(w_dff_B_ZYuOm7OY3_2),.clk(gclk));
	jdff dff_B_cioyhJK83_2(.din(w_dff_B_ZYuOm7OY3_2),.dout(w_dff_B_cioyhJK83_2),.clk(gclk));
	jdff dff_B_elFtxs0Y6_2(.din(w_dff_B_cioyhJK83_2),.dout(w_dff_B_elFtxs0Y6_2),.clk(gclk));
	jdff dff_B_p9cx9ORI7_2(.din(w_dff_B_elFtxs0Y6_2),.dout(w_dff_B_p9cx9ORI7_2),.clk(gclk));
	jdff dff_B_iayFpKPe8_2(.din(w_dff_B_p9cx9ORI7_2),.dout(w_dff_B_iayFpKPe8_2),.clk(gclk));
	jdff dff_B_d5WzPutg1_2(.din(w_dff_B_iayFpKPe8_2),.dout(w_dff_B_d5WzPutg1_2),.clk(gclk));
	jdff dff_B_v4QTKvHN8_2(.din(w_dff_B_d5WzPutg1_2),.dout(w_dff_B_v4QTKvHN8_2),.clk(gclk));
	jdff dff_B_vPkN0wTH5_2(.din(w_dff_B_v4QTKvHN8_2),.dout(w_dff_B_vPkN0wTH5_2),.clk(gclk));
	jdff dff_B_xp4wdqk08_2(.din(w_dff_B_vPkN0wTH5_2),.dout(w_dff_B_xp4wdqk08_2),.clk(gclk));
	jdff dff_B_kHzcuWf18_2(.din(w_dff_B_xp4wdqk08_2),.dout(w_dff_B_kHzcuWf18_2),.clk(gclk));
	jdff dff_B_jpK13zcP3_2(.din(w_dff_B_kHzcuWf18_2),.dout(w_dff_B_jpK13zcP3_2),.clk(gclk));
	jdff dff_B_pLF0hSJ70_2(.din(w_dff_B_jpK13zcP3_2),.dout(w_dff_B_pLF0hSJ70_2),.clk(gclk));
	jdff dff_B_O1UkgqKR0_2(.din(w_dff_B_pLF0hSJ70_2),.dout(w_dff_B_O1UkgqKR0_2),.clk(gclk));
	jdff dff_B_lTfHWvH69_2(.din(w_dff_B_O1UkgqKR0_2),.dout(w_dff_B_lTfHWvH69_2),.clk(gclk));
	jdff dff_B_g1daqpg70_2(.din(w_dff_B_lTfHWvH69_2),.dout(w_dff_B_g1daqpg70_2),.clk(gclk));
	jdff dff_B_EBX5IZm07_2(.din(w_dff_B_g1daqpg70_2),.dout(w_dff_B_EBX5IZm07_2),.clk(gclk));
	jdff dff_B_2k4ldK4S1_2(.din(w_dff_B_EBX5IZm07_2),.dout(w_dff_B_2k4ldK4S1_2),.clk(gclk));
	jdff dff_B_hFVTBlBT9_2(.din(w_dff_B_2k4ldK4S1_2),.dout(w_dff_B_hFVTBlBT9_2),.clk(gclk));
	jdff dff_B_Qfs7R1rE8_2(.din(w_dff_B_hFVTBlBT9_2),.dout(w_dff_B_Qfs7R1rE8_2),.clk(gclk));
	jdff dff_B_RCNwG5CY5_2(.din(w_dff_B_Qfs7R1rE8_2),.dout(w_dff_B_RCNwG5CY5_2),.clk(gclk));
	jdff dff_B_SbH6XqLT6_2(.din(w_dff_B_RCNwG5CY5_2),.dout(w_dff_B_SbH6XqLT6_2),.clk(gclk));
	jdff dff_B_ewLWYV3L8_2(.din(w_dff_B_SbH6XqLT6_2),.dout(w_dff_B_ewLWYV3L8_2),.clk(gclk));
	jdff dff_B_sSTI7Un12_2(.din(w_dff_B_ewLWYV3L8_2),.dout(w_dff_B_sSTI7Un12_2),.clk(gclk));
	jdff dff_B_a2c98eeB3_2(.din(w_dff_B_sSTI7Un12_2),.dout(w_dff_B_a2c98eeB3_2),.clk(gclk));
	jdff dff_B_XuSnMPXR4_2(.din(w_dff_B_a2c98eeB3_2),.dout(w_dff_B_XuSnMPXR4_2),.clk(gclk));
	jdff dff_B_v3ORR4x87_2(.din(w_dff_B_XuSnMPXR4_2),.dout(w_dff_B_v3ORR4x87_2),.clk(gclk));
	jdff dff_B_aBYn8zWe1_2(.din(w_dff_B_v3ORR4x87_2),.dout(w_dff_B_aBYn8zWe1_2),.clk(gclk));
	jdff dff_B_RsaprTqE6_2(.din(w_dff_B_aBYn8zWe1_2),.dout(w_dff_B_RsaprTqE6_2),.clk(gclk));
	jdff dff_B_FrYpMJtv9_2(.din(w_dff_B_RsaprTqE6_2),.dout(w_dff_B_FrYpMJtv9_2),.clk(gclk));
	jdff dff_B_7Obk5NuS3_2(.din(w_dff_B_FrYpMJtv9_2),.dout(w_dff_B_7Obk5NuS3_2),.clk(gclk));
	jdff dff_B_xdHqNUEm5_2(.din(w_dff_B_7Obk5NuS3_2),.dout(w_dff_B_xdHqNUEm5_2),.clk(gclk));
	jdff dff_B_0P9RNZtB5_2(.din(w_dff_B_xdHqNUEm5_2),.dout(w_dff_B_0P9RNZtB5_2),.clk(gclk));
	jdff dff_B_zHkCpcXH2_2(.din(w_dff_B_0P9RNZtB5_2),.dout(w_dff_B_zHkCpcXH2_2),.clk(gclk));
	jdff dff_A_tVLqk79Y1_1(.dout(w_n1827_0[1]),.din(w_dff_A_tVLqk79Y1_1),.clk(gclk));
	jdff dff_B_zqUqH8KZ3_1(.din(n1825),.dout(w_dff_B_zqUqH8KZ3_1),.clk(gclk));
	jdff dff_B_RhWltqDJ3_2(.din(n1803),.dout(w_dff_B_RhWltqDJ3_2),.clk(gclk));
	jdff dff_B_CnBM2kD77_2(.din(w_dff_B_RhWltqDJ3_2),.dout(w_dff_B_CnBM2kD77_2),.clk(gclk));
	jdff dff_B_IzhKd0yn0_2(.din(w_dff_B_CnBM2kD77_2),.dout(w_dff_B_IzhKd0yn0_2),.clk(gclk));
	jdff dff_B_XU4O6faH4_2(.din(w_dff_B_IzhKd0yn0_2),.dout(w_dff_B_XU4O6faH4_2),.clk(gclk));
	jdff dff_B_El91niX44_2(.din(w_dff_B_XU4O6faH4_2),.dout(w_dff_B_El91niX44_2),.clk(gclk));
	jdff dff_B_CxA3bteM8_2(.din(w_dff_B_El91niX44_2),.dout(w_dff_B_CxA3bteM8_2),.clk(gclk));
	jdff dff_B_FdnckxMr0_2(.din(w_dff_B_CxA3bteM8_2),.dout(w_dff_B_FdnckxMr0_2),.clk(gclk));
	jdff dff_B_twRzAU7V4_2(.din(w_dff_B_FdnckxMr0_2),.dout(w_dff_B_twRzAU7V4_2),.clk(gclk));
	jdff dff_B_HEFT2mGk1_2(.din(w_dff_B_twRzAU7V4_2),.dout(w_dff_B_HEFT2mGk1_2),.clk(gclk));
	jdff dff_B_B3WgssQZ3_2(.din(w_dff_B_HEFT2mGk1_2),.dout(w_dff_B_B3WgssQZ3_2),.clk(gclk));
	jdff dff_B_8hpJyFHe5_2(.din(w_dff_B_B3WgssQZ3_2),.dout(w_dff_B_8hpJyFHe5_2),.clk(gclk));
	jdff dff_B_34vZx5tq6_2(.din(w_dff_B_8hpJyFHe5_2),.dout(w_dff_B_34vZx5tq6_2),.clk(gclk));
	jdff dff_B_LjR792se1_2(.din(w_dff_B_34vZx5tq6_2),.dout(w_dff_B_LjR792se1_2),.clk(gclk));
	jdff dff_B_72iKWtpb5_2(.din(w_dff_B_LjR792se1_2),.dout(w_dff_B_72iKWtpb5_2),.clk(gclk));
	jdff dff_B_rMNZlLd74_2(.din(w_dff_B_72iKWtpb5_2),.dout(w_dff_B_rMNZlLd74_2),.clk(gclk));
	jdff dff_B_hvEvsA8i0_2(.din(w_dff_B_rMNZlLd74_2),.dout(w_dff_B_hvEvsA8i0_2),.clk(gclk));
	jdff dff_B_HCkalJ7L2_2(.din(w_dff_B_hvEvsA8i0_2),.dout(w_dff_B_HCkalJ7L2_2),.clk(gclk));
	jdff dff_B_Sg7lhnNc7_2(.din(w_dff_B_HCkalJ7L2_2),.dout(w_dff_B_Sg7lhnNc7_2),.clk(gclk));
	jdff dff_B_dJImzno93_2(.din(w_dff_B_Sg7lhnNc7_2),.dout(w_dff_B_dJImzno93_2),.clk(gclk));
	jdff dff_B_vKb5FWI98_2(.din(w_dff_B_dJImzno93_2),.dout(w_dff_B_vKb5FWI98_2),.clk(gclk));
	jdff dff_B_P1kVvgXl4_2(.din(w_dff_B_vKb5FWI98_2),.dout(w_dff_B_P1kVvgXl4_2),.clk(gclk));
	jdff dff_B_gM3Jqd4j5_2(.din(w_dff_B_P1kVvgXl4_2),.dout(w_dff_B_gM3Jqd4j5_2),.clk(gclk));
	jdff dff_B_xb7wssoE8_2(.din(w_dff_B_gM3Jqd4j5_2),.dout(w_dff_B_xb7wssoE8_2),.clk(gclk));
	jdff dff_B_keaVsMcq6_2(.din(w_dff_B_xb7wssoE8_2),.dout(w_dff_B_keaVsMcq6_2),.clk(gclk));
	jdff dff_B_bMeNLmQj6_2(.din(w_dff_B_keaVsMcq6_2),.dout(w_dff_B_bMeNLmQj6_2),.clk(gclk));
	jdff dff_B_ZHLi5hij9_2(.din(w_dff_B_bMeNLmQj6_2),.dout(w_dff_B_ZHLi5hij9_2),.clk(gclk));
	jdff dff_B_GekzxAFp3_2(.din(w_dff_B_ZHLi5hij9_2),.dout(w_dff_B_GekzxAFp3_2),.clk(gclk));
	jdff dff_B_HS7poe923_2(.din(w_dff_B_GekzxAFp3_2),.dout(w_dff_B_HS7poe923_2),.clk(gclk));
	jdff dff_B_M7cw7VQS9_2(.din(w_dff_B_HS7poe923_2),.dout(w_dff_B_M7cw7VQS9_2),.clk(gclk));
	jdff dff_B_IitJrHY92_2(.din(w_dff_B_M7cw7VQS9_2),.dout(w_dff_B_IitJrHY92_2),.clk(gclk));
	jdff dff_B_MV9rd15C1_2(.din(w_dff_B_IitJrHY92_2),.dout(w_dff_B_MV9rd15C1_2),.clk(gclk));
	jdff dff_B_Xp0vBTyE8_2(.din(w_dff_B_MV9rd15C1_2),.dout(w_dff_B_Xp0vBTyE8_2),.clk(gclk));
	jdff dff_B_9c6zEnAY6_2(.din(w_dff_B_Xp0vBTyE8_2),.dout(w_dff_B_9c6zEnAY6_2),.clk(gclk));
	jdff dff_B_wzbll3z81_2(.din(w_dff_B_9c6zEnAY6_2),.dout(w_dff_B_wzbll3z81_2),.clk(gclk));
	jdff dff_B_qBw5QAhP3_2(.din(w_dff_B_wzbll3z81_2),.dout(w_dff_B_qBw5QAhP3_2),.clk(gclk));
	jdff dff_B_a7HoWehd0_2(.din(w_dff_B_qBw5QAhP3_2),.dout(w_dff_B_a7HoWehd0_2),.clk(gclk));
	jdff dff_B_ps2IY3dJ6_2(.din(w_dff_B_a7HoWehd0_2),.dout(w_dff_B_ps2IY3dJ6_2),.clk(gclk));
	jdff dff_B_mG6nYk3B3_2(.din(w_dff_B_ps2IY3dJ6_2),.dout(w_dff_B_mG6nYk3B3_2),.clk(gclk));
	jdff dff_B_tztcrnI39_2(.din(w_dff_B_mG6nYk3B3_2),.dout(w_dff_B_tztcrnI39_2),.clk(gclk));
	jdff dff_B_ioHryxFd7_2(.din(w_dff_B_tztcrnI39_2),.dout(w_dff_B_ioHryxFd7_2),.clk(gclk));
	jdff dff_B_Z7awHPYz3_2(.din(w_dff_B_ioHryxFd7_2),.dout(w_dff_B_Z7awHPYz3_2),.clk(gclk));
	jdff dff_B_gDyZj84K6_2(.din(w_dff_B_Z7awHPYz3_2),.dout(w_dff_B_gDyZj84K6_2),.clk(gclk));
	jdff dff_B_1Jwqxdfo2_1(.din(n1809),.dout(w_dff_B_1Jwqxdfo2_1),.clk(gclk));
	jdff dff_B_phKCi7S75_1(.din(w_dff_B_1Jwqxdfo2_1),.dout(w_dff_B_phKCi7S75_1),.clk(gclk));
	jdff dff_B_tblBrehd0_2(.din(n1808),.dout(w_dff_B_tblBrehd0_2),.clk(gclk));
	jdff dff_B_itSFHr903_2(.din(w_dff_B_tblBrehd0_2),.dout(w_dff_B_itSFHr903_2),.clk(gclk));
	jdff dff_B_b4lFKQdd9_2(.din(w_dff_B_itSFHr903_2),.dout(w_dff_B_b4lFKQdd9_2),.clk(gclk));
	jdff dff_B_EnfK4HhG4_2(.din(w_dff_B_b4lFKQdd9_2),.dout(w_dff_B_EnfK4HhG4_2),.clk(gclk));
	jdff dff_B_MBKDZO3U1_2(.din(w_dff_B_EnfK4HhG4_2),.dout(w_dff_B_MBKDZO3U1_2),.clk(gclk));
	jdff dff_B_P8wlmhnz0_2(.din(w_dff_B_MBKDZO3U1_2),.dout(w_dff_B_P8wlmhnz0_2),.clk(gclk));
	jdff dff_B_QHhqZK2W6_2(.din(w_dff_B_P8wlmhnz0_2),.dout(w_dff_B_QHhqZK2W6_2),.clk(gclk));
	jdff dff_B_ko7SEAmP5_2(.din(w_dff_B_QHhqZK2W6_2),.dout(w_dff_B_ko7SEAmP5_2),.clk(gclk));
	jdff dff_B_b9vnJDJZ6_2(.din(w_dff_B_ko7SEAmP5_2),.dout(w_dff_B_b9vnJDJZ6_2),.clk(gclk));
	jdff dff_B_7xP3nVcU0_2(.din(w_dff_B_b9vnJDJZ6_2),.dout(w_dff_B_7xP3nVcU0_2),.clk(gclk));
	jdff dff_B_M9E2UCpg2_2(.din(w_dff_B_7xP3nVcU0_2),.dout(w_dff_B_M9E2UCpg2_2),.clk(gclk));
	jdff dff_B_rYoCC4SL4_2(.din(w_dff_B_M9E2UCpg2_2),.dout(w_dff_B_rYoCC4SL4_2),.clk(gclk));
	jdff dff_B_0TIE7HMF9_2(.din(w_dff_B_rYoCC4SL4_2),.dout(w_dff_B_0TIE7HMF9_2),.clk(gclk));
	jdff dff_B_k06ZKsXd1_2(.din(w_dff_B_0TIE7HMF9_2),.dout(w_dff_B_k06ZKsXd1_2),.clk(gclk));
	jdff dff_B_WlkIrWxy0_2(.din(w_dff_B_k06ZKsXd1_2),.dout(w_dff_B_WlkIrWxy0_2),.clk(gclk));
	jdff dff_B_orkWzp2v5_2(.din(w_dff_B_WlkIrWxy0_2),.dout(w_dff_B_orkWzp2v5_2),.clk(gclk));
	jdff dff_B_YvDgYskx9_2(.din(w_dff_B_orkWzp2v5_2),.dout(w_dff_B_YvDgYskx9_2),.clk(gclk));
	jdff dff_B_Li9pWwx11_2(.din(w_dff_B_YvDgYskx9_2),.dout(w_dff_B_Li9pWwx11_2),.clk(gclk));
	jdff dff_B_dpQ1y37P8_2(.din(w_dff_B_Li9pWwx11_2),.dout(w_dff_B_dpQ1y37P8_2),.clk(gclk));
	jdff dff_B_4Kqvo8Qx4_2(.din(w_dff_B_dpQ1y37P8_2),.dout(w_dff_B_4Kqvo8Qx4_2),.clk(gclk));
	jdff dff_B_chCfoMZa5_2(.din(w_dff_B_4Kqvo8Qx4_2),.dout(w_dff_B_chCfoMZa5_2),.clk(gclk));
	jdff dff_B_sDyJGmHR4_2(.din(w_dff_B_chCfoMZa5_2),.dout(w_dff_B_sDyJGmHR4_2),.clk(gclk));
	jdff dff_B_iCgeaUcJ4_2(.din(w_dff_B_sDyJGmHR4_2),.dout(w_dff_B_iCgeaUcJ4_2),.clk(gclk));
	jdff dff_B_3YQhtyL10_2(.din(w_dff_B_iCgeaUcJ4_2),.dout(w_dff_B_3YQhtyL10_2),.clk(gclk));
	jdff dff_B_1d5XGaJf0_2(.din(w_dff_B_3YQhtyL10_2),.dout(w_dff_B_1d5XGaJf0_2),.clk(gclk));
	jdff dff_B_xG0VBjjW4_2(.din(w_dff_B_1d5XGaJf0_2),.dout(w_dff_B_xG0VBjjW4_2),.clk(gclk));
	jdff dff_B_8qLdaMuI1_2(.din(w_dff_B_xG0VBjjW4_2),.dout(w_dff_B_8qLdaMuI1_2),.clk(gclk));
	jdff dff_B_tNLsAqB68_2(.din(w_dff_B_8qLdaMuI1_2),.dout(w_dff_B_tNLsAqB68_2),.clk(gclk));
	jdff dff_B_JHPb6ycA3_2(.din(w_dff_B_tNLsAqB68_2),.dout(w_dff_B_JHPb6ycA3_2),.clk(gclk));
	jdff dff_B_hhgj1rXA4_2(.din(w_dff_B_JHPb6ycA3_2),.dout(w_dff_B_hhgj1rXA4_2),.clk(gclk));
	jdff dff_B_aJE1NL4l2_2(.din(w_dff_B_hhgj1rXA4_2),.dout(w_dff_B_aJE1NL4l2_2),.clk(gclk));
	jdff dff_B_5wSGGqLT0_2(.din(w_dff_B_aJE1NL4l2_2),.dout(w_dff_B_5wSGGqLT0_2),.clk(gclk));
	jdff dff_B_KjWQhbJj2_2(.din(w_dff_B_5wSGGqLT0_2),.dout(w_dff_B_KjWQhbJj2_2),.clk(gclk));
	jdff dff_B_Li6AQjSy2_2(.din(w_dff_B_KjWQhbJj2_2),.dout(w_dff_B_Li6AQjSy2_2),.clk(gclk));
	jdff dff_B_aDwAbSO98_2(.din(w_dff_B_Li6AQjSy2_2),.dout(w_dff_B_aDwAbSO98_2),.clk(gclk));
	jdff dff_B_qKjbUunT4_2(.din(w_dff_B_aDwAbSO98_2),.dout(w_dff_B_qKjbUunT4_2),.clk(gclk));
	jdff dff_B_KgVcwmGA5_2(.din(w_dff_B_qKjbUunT4_2),.dout(w_dff_B_KgVcwmGA5_2),.clk(gclk));
	jdff dff_B_IWPsV1KB9_2(.din(w_dff_B_KgVcwmGA5_2),.dout(w_dff_B_IWPsV1KB9_2),.clk(gclk));
	jdff dff_B_mdap9Y3v1_2(.din(w_dff_B_IWPsV1KB9_2),.dout(w_dff_B_mdap9Y3v1_2),.clk(gclk));
	jdff dff_B_ZbH0ly908_2(.din(n1807),.dout(w_dff_B_ZbH0ly908_2),.clk(gclk));
	jdff dff_B_G79aM3YV9_2(.din(w_dff_B_ZbH0ly908_2),.dout(w_dff_B_G79aM3YV9_2),.clk(gclk));
	jdff dff_B_6CMoaR1y9_2(.din(w_dff_B_G79aM3YV9_2),.dout(w_dff_B_6CMoaR1y9_2),.clk(gclk));
	jdff dff_B_JcSzmsje1_2(.din(w_dff_B_6CMoaR1y9_2),.dout(w_dff_B_JcSzmsje1_2),.clk(gclk));
	jdff dff_B_C5ETVcMd9_2(.din(w_dff_B_JcSzmsje1_2),.dout(w_dff_B_C5ETVcMd9_2),.clk(gclk));
	jdff dff_B_WTu8ztxl0_2(.din(w_dff_B_C5ETVcMd9_2),.dout(w_dff_B_WTu8ztxl0_2),.clk(gclk));
	jdff dff_B_lOzQHJi20_2(.din(w_dff_B_WTu8ztxl0_2),.dout(w_dff_B_lOzQHJi20_2),.clk(gclk));
	jdff dff_B_9MtAWHBZ1_2(.din(w_dff_B_lOzQHJi20_2),.dout(w_dff_B_9MtAWHBZ1_2),.clk(gclk));
	jdff dff_B_fkX8zeqN4_2(.din(w_dff_B_9MtAWHBZ1_2),.dout(w_dff_B_fkX8zeqN4_2),.clk(gclk));
	jdff dff_B_5GRe2zu69_2(.din(w_dff_B_fkX8zeqN4_2),.dout(w_dff_B_5GRe2zu69_2),.clk(gclk));
	jdff dff_B_2o673iNC0_2(.din(w_dff_B_5GRe2zu69_2),.dout(w_dff_B_2o673iNC0_2),.clk(gclk));
	jdff dff_B_kSb3DJfx9_2(.din(w_dff_B_2o673iNC0_2),.dout(w_dff_B_kSb3DJfx9_2),.clk(gclk));
	jdff dff_B_OjADhL0S8_2(.din(w_dff_B_kSb3DJfx9_2),.dout(w_dff_B_OjADhL0S8_2),.clk(gclk));
	jdff dff_B_vLZP8QfX8_2(.din(w_dff_B_OjADhL0S8_2),.dout(w_dff_B_vLZP8QfX8_2),.clk(gclk));
	jdff dff_B_VJWLKmx15_2(.din(w_dff_B_vLZP8QfX8_2),.dout(w_dff_B_VJWLKmx15_2),.clk(gclk));
	jdff dff_B_OPV2nKYI3_2(.din(w_dff_B_VJWLKmx15_2),.dout(w_dff_B_OPV2nKYI3_2),.clk(gclk));
	jdff dff_B_QFb84w6R1_2(.din(w_dff_B_OPV2nKYI3_2),.dout(w_dff_B_QFb84w6R1_2),.clk(gclk));
	jdff dff_B_JePpGwpI0_2(.din(w_dff_B_QFb84w6R1_2),.dout(w_dff_B_JePpGwpI0_2),.clk(gclk));
	jdff dff_B_1GmecIhJ0_2(.din(w_dff_B_JePpGwpI0_2),.dout(w_dff_B_1GmecIhJ0_2),.clk(gclk));
	jdff dff_B_rzNei0n85_2(.din(w_dff_B_1GmecIhJ0_2),.dout(w_dff_B_rzNei0n85_2),.clk(gclk));
	jdff dff_B_juJQoHav9_2(.din(w_dff_B_rzNei0n85_2),.dout(w_dff_B_juJQoHav9_2),.clk(gclk));
	jdff dff_B_aIzD0oVX4_2(.din(w_dff_B_juJQoHav9_2),.dout(w_dff_B_aIzD0oVX4_2),.clk(gclk));
	jdff dff_B_cm4VAGbl5_2(.din(w_dff_B_aIzD0oVX4_2),.dout(w_dff_B_cm4VAGbl5_2),.clk(gclk));
	jdff dff_B_Cc3J9Q767_2(.din(w_dff_B_cm4VAGbl5_2),.dout(w_dff_B_Cc3J9Q767_2),.clk(gclk));
	jdff dff_B_b14ti8Um9_2(.din(w_dff_B_Cc3J9Q767_2),.dout(w_dff_B_b14ti8Um9_2),.clk(gclk));
	jdff dff_B_DqGfZ6187_2(.din(w_dff_B_b14ti8Um9_2),.dout(w_dff_B_DqGfZ6187_2),.clk(gclk));
	jdff dff_B_gIpXCyK06_2(.din(w_dff_B_DqGfZ6187_2),.dout(w_dff_B_gIpXCyK06_2),.clk(gclk));
	jdff dff_B_XTcIuCbm7_2(.din(w_dff_B_gIpXCyK06_2),.dout(w_dff_B_XTcIuCbm7_2),.clk(gclk));
	jdff dff_B_UtYEnfsV0_2(.din(w_dff_B_XTcIuCbm7_2),.dout(w_dff_B_UtYEnfsV0_2),.clk(gclk));
	jdff dff_B_dN1bwkGW7_2(.din(w_dff_B_UtYEnfsV0_2),.dout(w_dff_B_dN1bwkGW7_2),.clk(gclk));
	jdff dff_B_wE6vxHHD9_2(.din(w_dff_B_dN1bwkGW7_2),.dout(w_dff_B_wE6vxHHD9_2),.clk(gclk));
	jdff dff_B_tv9fE4Wm7_2(.din(w_dff_B_wE6vxHHD9_2),.dout(w_dff_B_tv9fE4Wm7_2),.clk(gclk));
	jdff dff_B_r6rsoiz94_2(.din(w_dff_B_tv9fE4Wm7_2),.dout(w_dff_B_r6rsoiz94_2),.clk(gclk));
	jdff dff_B_MZF1mq131_2(.din(w_dff_B_r6rsoiz94_2),.dout(w_dff_B_MZF1mq131_2),.clk(gclk));
	jdff dff_B_rBqYzJFi0_2(.din(w_dff_B_MZF1mq131_2),.dout(w_dff_B_rBqYzJFi0_2),.clk(gclk));
	jdff dff_B_32RysaDw5_2(.din(w_dff_B_rBqYzJFi0_2),.dout(w_dff_B_32RysaDw5_2),.clk(gclk));
	jdff dff_B_ELbAWnj27_2(.din(w_dff_B_32RysaDw5_2),.dout(w_dff_B_ELbAWnj27_2),.clk(gclk));
	jdff dff_B_wxgzp5I84_2(.din(w_dff_B_ELbAWnj27_2),.dout(w_dff_B_wxgzp5I84_2),.clk(gclk));
	jdff dff_B_K1XiXgqB3_2(.din(w_dff_B_wxgzp5I84_2),.dout(w_dff_B_K1XiXgqB3_2),.clk(gclk));
	jdff dff_B_k0NqPBpU2_2(.din(w_dff_B_K1XiXgqB3_2),.dout(w_dff_B_k0NqPBpU2_2),.clk(gclk));
	jdff dff_B_BjKCTGGi5_2(.din(w_dff_B_k0NqPBpU2_2),.dout(w_dff_B_BjKCTGGi5_2),.clk(gclk));
	jdff dff_B_ePWWhOLk3_2(.din(n1806),.dout(w_dff_B_ePWWhOLk3_2),.clk(gclk));
	jdff dff_B_rylctyCW3_1(.din(n1804),.dout(w_dff_B_rylctyCW3_1),.clk(gclk));
	jdff dff_B_h7ZEuDmb1_2(.din(n1775),.dout(w_dff_B_h7ZEuDmb1_2),.clk(gclk));
	jdff dff_B_XW4nAG976_2(.din(w_dff_B_h7ZEuDmb1_2),.dout(w_dff_B_XW4nAG976_2),.clk(gclk));
	jdff dff_B_O7fUxSqP4_2(.din(w_dff_B_XW4nAG976_2),.dout(w_dff_B_O7fUxSqP4_2),.clk(gclk));
	jdff dff_B_cntEbQlR6_2(.din(w_dff_B_O7fUxSqP4_2),.dout(w_dff_B_cntEbQlR6_2),.clk(gclk));
	jdff dff_B_hAMfUTEM1_2(.din(w_dff_B_cntEbQlR6_2),.dout(w_dff_B_hAMfUTEM1_2),.clk(gclk));
	jdff dff_B_mK4vNNN49_2(.din(w_dff_B_hAMfUTEM1_2),.dout(w_dff_B_mK4vNNN49_2),.clk(gclk));
	jdff dff_B_JrSkrzBt2_2(.din(w_dff_B_mK4vNNN49_2),.dout(w_dff_B_JrSkrzBt2_2),.clk(gclk));
	jdff dff_B_4mXIw4G31_2(.din(w_dff_B_JrSkrzBt2_2),.dout(w_dff_B_4mXIw4G31_2),.clk(gclk));
	jdff dff_B_s6AGkWEw1_2(.din(w_dff_B_4mXIw4G31_2),.dout(w_dff_B_s6AGkWEw1_2),.clk(gclk));
	jdff dff_B_pmLr7PiL8_2(.din(w_dff_B_s6AGkWEw1_2),.dout(w_dff_B_pmLr7PiL8_2),.clk(gclk));
	jdff dff_B_gmcXlm5D8_2(.din(w_dff_B_pmLr7PiL8_2),.dout(w_dff_B_gmcXlm5D8_2),.clk(gclk));
	jdff dff_B_5rz6BiMc4_2(.din(w_dff_B_gmcXlm5D8_2),.dout(w_dff_B_5rz6BiMc4_2),.clk(gclk));
	jdff dff_B_q7FfvtVf9_2(.din(w_dff_B_5rz6BiMc4_2),.dout(w_dff_B_q7FfvtVf9_2),.clk(gclk));
	jdff dff_B_i1n3hgjd3_2(.din(w_dff_B_q7FfvtVf9_2),.dout(w_dff_B_i1n3hgjd3_2),.clk(gclk));
	jdff dff_B_Xuwj6L0a2_2(.din(w_dff_B_i1n3hgjd3_2),.dout(w_dff_B_Xuwj6L0a2_2),.clk(gclk));
	jdff dff_B_sWDo2ve35_2(.din(w_dff_B_Xuwj6L0a2_2),.dout(w_dff_B_sWDo2ve35_2),.clk(gclk));
	jdff dff_B_KjibuJZR4_2(.din(w_dff_B_sWDo2ve35_2),.dout(w_dff_B_KjibuJZR4_2),.clk(gclk));
	jdff dff_B_SzcEGYeH3_2(.din(w_dff_B_KjibuJZR4_2),.dout(w_dff_B_SzcEGYeH3_2),.clk(gclk));
	jdff dff_B_tk7FzxHW9_2(.din(w_dff_B_SzcEGYeH3_2),.dout(w_dff_B_tk7FzxHW9_2),.clk(gclk));
	jdff dff_B_GAuTDEMm7_2(.din(w_dff_B_tk7FzxHW9_2),.dout(w_dff_B_GAuTDEMm7_2),.clk(gclk));
	jdff dff_B_jngsmj9g9_2(.din(w_dff_B_GAuTDEMm7_2),.dout(w_dff_B_jngsmj9g9_2),.clk(gclk));
	jdff dff_B_nbJs1NSe2_2(.din(w_dff_B_jngsmj9g9_2),.dout(w_dff_B_nbJs1NSe2_2),.clk(gclk));
	jdff dff_B_1eRRJEff6_2(.din(w_dff_B_nbJs1NSe2_2),.dout(w_dff_B_1eRRJEff6_2),.clk(gclk));
	jdff dff_B_jcR34zYb3_2(.din(w_dff_B_1eRRJEff6_2),.dout(w_dff_B_jcR34zYb3_2),.clk(gclk));
	jdff dff_B_RNtilsMg7_2(.din(w_dff_B_jcR34zYb3_2),.dout(w_dff_B_RNtilsMg7_2),.clk(gclk));
	jdff dff_B_DiD7gUH36_2(.din(w_dff_B_RNtilsMg7_2),.dout(w_dff_B_DiD7gUH36_2),.clk(gclk));
	jdff dff_B_rO4yVsyQ4_2(.din(w_dff_B_DiD7gUH36_2),.dout(w_dff_B_rO4yVsyQ4_2),.clk(gclk));
	jdff dff_B_yTAa6dks2_2(.din(w_dff_B_rO4yVsyQ4_2),.dout(w_dff_B_yTAa6dks2_2),.clk(gclk));
	jdff dff_B_qClnjBV82_2(.din(w_dff_B_yTAa6dks2_2),.dout(w_dff_B_qClnjBV82_2),.clk(gclk));
	jdff dff_B_kczOsCVx1_2(.din(w_dff_B_qClnjBV82_2),.dout(w_dff_B_kczOsCVx1_2),.clk(gclk));
	jdff dff_B_lyAVx1hT1_2(.din(w_dff_B_kczOsCVx1_2),.dout(w_dff_B_lyAVx1hT1_2),.clk(gclk));
	jdff dff_B_kpM1PmIY4_2(.din(w_dff_B_lyAVx1hT1_2),.dout(w_dff_B_kpM1PmIY4_2),.clk(gclk));
	jdff dff_B_92dOxz244_2(.din(w_dff_B_kpM1PmIY4_2),.dout(w_dff_B_92dOxz244_2),.clk(gclk));
	jdff dff_B_YdQRyXzW3_2(.din(w_dff_B_92dOxz244_2),.dout(w_dff_B_YdQRyXzW3_2),.clk(gclk));
	jdff dff_B_h5K9Dn802_2(.din(w_dff_B_YdQRyXzW3_2),.dout(w_dff_B_h5K9Dn802_2),.clk(gclk));
	jdff dff_B_z0jUJwcp6_2(.din(w_dff_B_h5K9Dn802_2),.dout(w_dff_B_z0jUJwcp6_2),.clk(gclk));
	jdff dff_B_QHULyD6b3_2(.din(w_dff_B_z0jUJwcp6_2),.dout(w_dff_B_QHULyD6b3_2),.clk(gclk));
	jdff dff_B_enjR0FLW7_2(.din(w_dff_B_QHULyD6b3_2),.dout(w_dff_B_enjR0FLW7_2),.clk(gclk));
	jdff dff_B_gbgBrA6H6_2(.din(w_dff_B_enjR0FLW7_2),.dout(w_dff_B_gbgBrA6H6_2),.clk(gclk));
	jdff dff_B_QTjBzVB43_1(.din(n1781),.dout(w_dff_B_QTjBzVB43_1),.clk(gclk));
	jdff dff_B_i90TR0Ua5_1(.din(w_dff_B_QTjBzVB43_1),.dout(w_dff_B_i90TR0Ua5_1),.clk(gclk));
	jdff dff_B_c4PhMsCI1_2(.din(n1780),.dout(w_dff_B_c4PhMsCI1_2),.clk(gclk));
	jdff dff_B_StDVmxxv0_2(.din(w_dff_B_c4PhMsCI1_2),.dout(w_dff_B_StDVmxxv0_2),.clk(gclk));
	jdff dff_B_3KKf0lg50_2(.din(w_dff_B_StDVmxxv0_2),.dout(w_dff_B_3KKf0lg50_2),.clk(gclk));
	jdff dff_B_OcTWDznu4_2(.din(w_dff_B_3KKf0lg50_2),.dout(w_dff_B_OcTWDznu4_2),.clk(gclk));
	jdff dff_B_MayoLo4z6_2(.din(w_dff_B_OcTWDznu4_2),.dout(w_dff_B_MayoLo4z6_2),.clk(gclk));
	jdff dff_B_e5Sz9ZE24_2(.din(w_dff_B_MayoLo4z6_2),.dout(w_dff_B_e5Sz9ZE24_2),.clk(gclk));
	jdff dff_B_NEolJuh88_2(.din(w_dff_B_e5Sz9ZE24_2),.dout(w_dff_B_NEolJuh88_2),.clk(gclk));
	jdff dff_B_Eh0OcCbs4_2(.din(w_dff_B_NEolJuh88_2),.dout(w_dff_B_Eh0OcCbs4_2),.clk(gclk));
	jdff dff_B_tK3opf0D2_2(.din(w_dff_B_Eh0OcCbs4_2),.dout(w_dff_B_tK3opf0D2_2),.clk(gclk));
	jdff dff_B_tPAK43lg2_2(.din(w_dff_B_tK3opf0D2_2),.dout(w_dff_B_tPAK43lg2_2),.clk(gclk));
	jdff dff_B_7Rp5K8FC7_2(.din(w_dff_B_tPAK43lg2_2),.dout(w_dff_B_7Rp5K8FC7_2),.clk(gclk));
	jdff dff_B_ONhdkeAp1_2(.din(w_dff_B_7Rp5K8FC7_2),.dout(w_dff_B_ONhdkeAp1_2),.clk(gclk));
	jdff dff_B_Y9fCuxhB1_2(.din(w_dff_B_ONhdkeAp1_2),.dout(w_dff_B_Y9fCuxhB1_2),.clk(gclk));
	jdff dff_B_PoFFkXua0_2(.din(w_dff_B_Y9fCuxhB1_2),.dout(w_dff_B_PoFFkXua0_2),.clk(gclk));
	jdff dff_B_9hCnEWZb8_2(.din(w_dff_B_PoFFkXua0_2),.dout(w_dff_B_9hCnEWZb8_2),.clk(gclk));
	jdff dff_B_QbOGr7ud5_2(.din(w_dff_B_9hCnEWZb8_2),.dout(w_dff_B_QbOGr7ud5_2),.clk(gclk));
	jdff dff_B_oUIGYaME2_2(.din(w_dff_B_QbOGr7ud5_2),.dout(w_dff_B_oUIGYaME2_2),.clk(gclk));
	jdff dff_B_cUjtq5cu9_2(.din(w_dff_B_oUIGYaME2_2),.dout(w_dff_B_cUjtq5cu9_2),.clk(gclk));
	jdff dff_B_C092x4oO9_2(.din(w_dff_B_cUjtq5cu9_2),.dout(w_dff_B_C092x4oO9_2),.clk(gclk));
	jdff dff_B_QwpZgVzd6_2(.din(w_dff_B_C092x4oO9_2),.dout(w_dff_B_QwpZgVzd6_2),.clk(gclk));
	jdff dff_B_CrRsneMV1_2(.din(w_dff_B_QwpZgVzd6_2),.dout(w_dff_B_CrRsneMV1_2),.clk(gclk));
	jdff dff_B_YAhGya4r9_2(.din(w_dff_B_CrRsneMV1_2),.dout(w_dff_B_YAhGya4r9_2),.clk(gclk));
	jdff dff_B_K7VY47iV8_2(.din(w_dff_B_YAhGya4r9_2),.dout(w_dff_B_K7VY47iV8_2),.clk(gclk));
	jdff dff_B_5eYdc7KG1_2(.din(w_dff_B_K7VY47iV8_2),.dout(w_dff_B_5eYdc7KG1_2),.clk(gclk));
	jdff dff_B_3V3F6zdX0_2(.din(w_dff_B_5eYdc7KG1_2),.dout(w_dff_B_3V3F6zdX0_2),.clk(gclk));
	jdff dff_B_6iv68eh54_2(.din(w_dff_B_3V3F6zdX0_2),.dout(w_dff_B_6iv68eh54_2),.clk(gclk));
	jdff dff_B_XZv4HD2E6_2(.din(w_dff_B_6iv68eh54_2),.dout(w_dff_B_XZv4HD2E6_2),.clk(gclk));
	jdff dff_B_sRTjxp2a0_2(.din(w_dff_B_XZv4HD2E6_2),.dout(w_dff_B_sRTjxp2a0_2),.clk(gclk));
	jdff dff_B_fv8t0Bza5_2(.din(w_dff_B_sRTjxp2a0_2),.dout(w_dff_B_fv8t0Bza5_2),.clk(gclk));
	jdff dff_B_k0LAeEIJ7_2(.din(w_dff_B_fv8t0Bza5_2),.dout(w_dff_B_k0LAeEIJ7_2),.clk(gclk));
	jdff dff_B_LGWN4t5i1_2(.din(w_dff_B_k0LAeEIJ7_2),.dout(w_dff_B_LGWN4t5i1_2),.clk(gclk));
	jdff dff_B_51cAvMAn6_2(.din(w_dff_B_LGWN4t5i1_2),.dout(w_dff_B_51cAvMAn6_2),.clk(gclk));
	jdff dff_B_85WyqBzm6_2(.din(w_dff_B_51cAvMAn6_2),.dout(w_dff_B_85WyqBzm6_2),.clk(gclk));
	jdff dff_B_pPRrrqhz7_2(.din(w_dff_B_85WyqBzm6_2),.dout(w_dff_B_pPRrrqhz7_2),.clk(gclk));
	jdff dff_B_wOY6VAb33_2(.din(w_dff_B_pPRrrqhz7_2),.dout(w_dff_B_wOY6VAb33_2),.clk(gclk));
	jdff dff_B_2DNCISpa2_2(.din(w_dff_B_wOY6VAb33_2),.dout(w_dff_B_2DNCISpa2_2),.clk(gclk));
	jdff dff_B_GmSNJfGn1_2(.din(n1779),.dout(w_dff_B_GmSNJfGn1_2),.clk(gclk));
	jdff dff_B_ieUl5OA25_2(.din(w_dff_B_GmSNJfGn1_2),.dout(w_dff_B_ieUl5OA25_2),.clk(gclk));
	jdff dff_B_Uuc2mR2h3_2(.din(w_dff_B_ieUl5OA25_2),.dout(w_dff_B_Uuc2mR2h3_2),.clk(gclk));
	jdff dff_B_LhCAu3xo2_2(.din(w_dff_B_Uuc2mR2h3_2),.dout(w_dff_B_LhCAu3xo2_2),.clk(gclk));
	jdff dff_B_HMMMaqZh7_2(.din(w_dff_B_LhCAu3xo2_2),.dout(w_dff_B_HMMMaqZh7_2),.clk(gclk));
	jdff dff_B_8TgWaTU67_2(.din(w_dff_B_HMMMaqZh7_2),.dout(w_dff_B_8TgWaTU67_2),.clk(gclk));
	jdff dff_B_zhmz6o6t0_2(.din(w_dff_B_8TgWaTU67_2),.dout(w_dff_B_zhmz6o6t0_2),.clk(gclk));
	jdff dff_B_HJxKRaJ90_2(.din(w_dff_B_zhmz6o6t0_2),.dout(w_dff_B_HJxKRaJ90_2),.clk(gclk));
	jdff dff_B_yNmbtX614_2(.din(w_dff_B_HJxKRaJ90_2),.dout(w_dff_B_yNmbtX614_2),.clk(gclk));
	jdff dff_B_1r47iof57_2(.din(w_dff_B_yNmbtX614_2),.dout(w_dff_B_1r47iof57_2),.clk(gclk));
	jdff dff_B_Q9SM2Lsz5_2(.din(w_dff_B_1r47iof57_2),.dout(w_dff_B_Q9SM2Lsz5_2),.clk(gclk));
	jdff dff_B_olZKlNhv5_2(.din(w_dff_B_Q9SM2Lsz5_2),.dout(w_dff_B_olZKlNhv5_2),.clk(gclk));
	jdff dff_B_G0wzwvvP3_2(.din(w_dff_B_olZKlNhv5_2),.dout(w_dff_B_G0wzwvvP3_2),.clk(gclk));
	jdff dff_B_aIk4xXLa3_2(.din(w_dff_B_G0wzwvvP3_2),.dout(w_dff_B_aIk4xXLa3_2),.clk(gclk));
	jdff dff_B_FDJEGcJc0_2(.din(w_dff_B_aIk4xXLa3_2),.dout(w_dff_B_FDJEGcJc0_2),.clk(gclk));
	jdff dff_B_xo97B67i0_2(.din(w_dff_B_FDJEGcJc0_2),.dout(w_dff_B_xo97B67i0_2),.clk(gclk));
	jdff dff_B_xra00VK92_2(.din(w_dff_B_xo97B67i0_2),.dout(w_dff_B_xra00VK92_2),.clk(gclk));
	jdff dff_B_7nprEDef0_2(.din(w_dff_B_xra00VK92_2),.dout(w_dff_B_7nprEDef0_2),.clk(gclk));
	jdff dff_B_4vkip1Mz2_2(.din(w_dff_B_7nprEDef0_2),.dout(w_dff_B_4vkip1Mz2_2),.clk(gclk));
	jdff dff_B_HSe8mv4g1_2(.din(w_dff_B_4vkip1Mz2_2),.dout(w_dff_B_HSe8mv4g1_2),.clk(gclk));
	jdff dff_B_YrW8t61X7_2(.din(w_dff_B_HSe8mv4g1_2),.dout(w_dff_B_YrW8t61X7_2),.clk(gclk));
	jdff dff_B_KLaxzF2E9_2(.din(w_dff_B_YrW8t61X7_2),.dout(w_dff_B_KLaxzF2E9_2),.clk(gclk));
	jdff dff_B_9FjxJDhb4_2(.din(w_dff_B_KLaxzF2E9_2),.dout(w_dff_B_9FjxJDhb4_2),.clk(gclk));
	jdff dff_B_A17wngXb2_2(.din(w_dff_B_9FjxJDhb4_2),.dout(w_dff_B_A17wngXb2_2),.clk(gclk));
	jdff dff_B_rB2Act2P8_2(.din(w_dff_B_A17wngXb2_2),.dout(w_dff_B_rB2Act2P8_2),.clk(gclk));
	jdff dff_B_3plsBdUM3_2(.din(w_dff_B_rB2Act2P8_2),.dout(w_dff_B_3plsBdUM3_2),.clk(gclk));
	jdff dff_B_902ADQ0l9_2(.din(w_dff_B_3plsBdUM3_2),.dout(w_dff_B_902ADQ0l9_2),.clk(gclk));
	jdff dff_B_ubUYKFxu5_2(.din(w_dff_B_902ADQ0l9_2),.dout(w_dff_B_ubUYKFxu5_2),.clk(gclk));
	jdff dff_B_xGAa1utb7_2(.din(w_dff_B_ubUYKFxu5_2),.dout(w_dff_B_xGAa1utb7_2),.clk(gclk));
	jdff dff_B_4sZXHQzC0_2(.din(w_dff_B_xGAa1utb7_2),.dout(w_dff_B_4sZXHQzC0_2),.clk(gclk));
	jdff dff_B_cNkkEb6X9_2(.din(w_dff_B_4sZXHQzC0_2),.dout(w_dff_B_cNkkEb6X9_2),.clk(gclk));
	jdff dff_B_e2SNW1oG5_2(.din(w_dff_B_cNkkEb6X9_2),.dout(w_dff_B_e2SNW1oG5_2),.clk(gclk));
	jdff dff_B_rZ6eexFO1_2(.din(w_dff_B_e2SNW1oG5_2),.dout(w_dff_B_rZ6eexFO1_2),.clk(gclk));
	jdff dff_B_Tsq3goMi8_2(.din(w_dff_B_rZ6eexFO1_2),.dout(w_dff_B_Tsq3goMi8_2),.clk(gclk));
	jdff dff_B_KBcD8O4V7_2(.din(w_dff_B_Tsq3goMi8_2),.dout(w_dff_B_KBcD8O4V7_2),.clk(gclk));
	jdff dff_B_vXqmdnz53_2(.din(w_dff_B_KBcD8O4V7_2),.dout(w_dff_B_vXqmdnz53_2),.clk(gclk));
	jdff dff_B_UX9PxSwT3_2(.din(w_dff_B_vXqmdnz53_2),.dout(w_dff_B_UX9PxSwT3_2),.clk(gclk));
	jdff dff_B_yUI2ohxu1_2(.din(w_dff_B_UX9PxSwT3_2),.dout(w_dff_B_yUI2ohxu1_2),.clk(gclk));
	jdff dff_B_gSyS7sQ69_2(.din(n1778),.dout(w_dff_B_gSyS7sQ69_2),.clk(gclk));
	jdff dff_B_Rr9uOYLY4_1(.din(n1776),.dout(w_dff_B_Rr9uOYLY4_1),.clk(gclk));
	jdff dff_B_okHtaBRA2_2(.din(n1740),.dout(w_dff_B_okHtaBRA2_2),.clk(gclk));
	jdff dff_B_xx9G1Dyj8_2(.din(w_dff_B_okHtaBRA2_2),.dout(w_dff_B_xx9G1Dyj8_2),.clk(gclk));
	jdff dff_B_yRag1ri84_2(.din(w_dff_B_xx9G1Dyj8_2),.dout(w_dff_B_yRag1ri84_2),.clk(gclk));
	jdff dff_B_SIMKDxEc0_2(.din(w_dff_B_yRag1ri84_2),.dout(w_dff_B_SIMKDxEc0_2),.clk(gclk));
	jdff dff_B_de8eGcce1_2(.din(w_dff_B_SIMKDxEc0_2),.dout(w_dff_B_de8eGcce1_2),.clk(gclk));
	jdff dff_B_zNqEkX4g3_2(.din(w_dff_B_de8eGcce1_2),.dout(w_dff_B_zNqEkX4g3_2),.clk(gclk));
	jdff dff_B_4qnSNbtp3_2(.din(w_dff_B_zNqEkX4g3_2),.dout(w_dff_B_4qnSNbtp3_2),.clk(gclk));
	jdff dff_B_E37uSIUu7_2(.din(w_dff_B_4qnSNbtp3_2),.dout(w_dff_B_E37uSIUu7_2),.clk(gclk));
	jdff dff_B_BU1yaWKR0_2(.din(w_dff_B_E37uSIUu7_2),.dout(w_dff_B_BU1yaWKR0_2),.clk(gclk));
	jdff dff_B_VMAeXGvG8_2(.din(w_dff_B_BU1yaWKR0_2),.dout(w_dff_B_VMAeXGvG8_2),.clk(gclk));
	jdff dff_B_63Z5XYfG8_2(.din(w_dff_B_VMAeXGvG8_2),.dout(w_dff_B_63Z5XYfG8_2),.clk(gclk));
	jdff dff_B_ZZnGvgRo4_2(.din(w_dff_B_63Z5XYfG8_2),.dout(w_dff_B_ZZnGvgRo4_2),.clk(gclk));
	jdff dff_B_f8kW5op81_2(.din(w_dff_B_ZZnGvgRo4_2),.dout(w_dff_B_f8kW5op81_2),.clk(gclk));
	jdff dff_B_WsTIjQt01_2(.din(w_dff_B_f8kW5op81_2),.dout(w_dff_B_WsTIjQt01_2),.clk(gclk));
	jdff dff_B_m4zY4HUi9_2(.din(w_dff_B_WsTIjQt01_2),.dout(w_dff_B_m4zY4HUi9_2),.clk(gclk));
	jdff dff_B_WS1Me9cY2_2(.din(w_dff_B_m4zY4HUi9_2),.dout(w_dff_B_WS1Me9cY2_2),.clk(gclk));
	jdff dff_B_9aMRIZGK7_2(.din(w_dff_B_WS1Me9cY2_2),.dout(w_dff_B_9aMRIZGK7_2),.clk(gclk));
	jdff dff_B_gEKPAs8u9_2(.din(w_dff_B_9aMRIZGK7_2),.dout(w_dff_B_gEKPAs8u9_2),.clk(gclk));
	jdff dff_B_RWvFzPX89_2(.din(w_dff_B_gEKPAs8u9_2),.dout(w_dff_B_RWvFzPX89_2),.clk(gclk));
	jdff dff_B_qsbvViJb7_2(.din(w_dff_B_RWvFzPX89_2),.dout(w_dff_B_qsbvViJb7_2),.clk(gclk));
	jdff dff_B_1hbuWucZ6_2(.din(w_dff_B_qsbvViJb7_2),.dout(w_dff_B_1hbuWucZ6_2),.clk(gclk));
	jdff dff_B_6hZsfQ1Q4_2(.din(w_dff_B_1hbuWucZ6_2),.dout(w_dff_B_6hZsfQ1Q4_2),.clk(gclk));
	jdff dff_B_ztzdxNGC1_2(.din(w_dff_B_6hZsfQ1Q4_2),.dout(w_dff_B_ztzdxNGC1_2),.clk(gclk));
	jdff dff_B_sfmfHssI1_2(.din(w_dff_B_ztzdxNGC1_2),.dout(w_dff_B_sfmfHssI1_2),.clk(gclk));
	jdff dff_B_W0YaUfP97_2(.din(w_dff_B_sfmfHssI1_2),.dout(w_dff_B_W0YaUfP97_2),.clk(gclk));
	jdff dff_B_Kx17gVau7_2(.din(w_dff_B_W0YaUfP97_2),.dout(w_dff_B_Kx17gVau7_2),.clk(gclk));
	jdff dff_B_A5AUQ41I8_2(.din(w_dff_B_Kx17gVau7_2),.dout(w_dff_B_A5AUQ41I8_2),.clk(gclk));
	jdff dff_B_rjO2eZd75_2(.din(w_dff_B_A5AUQ41I8_2),.dout(w_dff_B_rjO2eZd75_2),.clk(gclk));
	jdff dff_B_0ZIOGgvX4_2(.din(w_dff_B_rjO2eZd75_2),.dout(w_dff_B_0ZIOGgvX4_2),.clk(gclk));
	jdff dff_B_zgmLNUQJ3_2(.din(w_dff_B_0ZIOGgvX4_2),.dout(w_dff_B_zgmLNUQJ3_2),.clk(gclk));
	jdff dff_B_MYyxT8Ur6_2(.din(w_dff_B_zgmLNUQJ3_2),.dout(w_dff_B_MYyxT8Ur6_2),.clk(gclk));
	jdff dff_B_dSWEfCHf0_2(.din(w_dff_B_MYyxT8Ur6_2),.dout(w_dff_B_dSWEfCHf0_2),.clk(gclk));
	jdff dff_B_hd1LKUtf0_2(.din(w_dff_B_dSWEfCHf0_2),.dout(w_dff_B_hd1LKUtf0_2),.clk(gclk));
	jdff dff_B_NPRYPLEI1_2(.din(w_dff_B_hd1LKUtf0_2),.dout(w_dff_B_NPRYPLEI1_2),.clk(gclk));
	jdff dff_B_h3LpYNfB5_2(.din(w_dff_B_NPRYPLEI1_2),.dout(w_dff_B_h3LpYNfB5_2),.clk(gclk));
	jdff dff_B_ZPhpAERb4_2(.din(w_dff_B_h3LpYNfB5_2),.dout(w_dff_B_ZPhpAERb4_2),.clk(gclk));
	jdff dff_B_SPRTuclL2_1(.din(n1746),.dout(w_dff_B_SPRTuclL2_1),.clk(gclk));
	jdff dff_B_Nayzih5N8_1(.din(w_dff_B_SPRTuclL2_1),.dout(w_dff_B_Nayzih5N8_1),.clk(gclk));
	jdff dff_B_stb9LMXH6_2(.din(n1745),.dout(w_dff_B_stb9LMXH6_2),.clk(gclk));
	jdff dff_B_geNNOI4z0_2(.din(w_dff_B_stb9LMXH6_2),.dout(w_dff_B_geNNOI4z0_2),.clk(gclk));
	jdff dff_B_JSH3k4pL4_2(.din(w_dff_B_geNNOI4z0_2),.dout(w_dff_B_JSH3k4pL4_2),.clk(gclk));
	jdff dff_B_SQBg60se5_2(.din(w_dff_B_JSH3k4pL4_2),.dout(w_dff_B_SQBg60se5_2),.clk(gclk));
	jdff dff_B_Ho41pmSb0_2(.din(w_dff_B_SQBg60se5_2),.dout(w_dff_B_Ho41pmSb0_2),.clk(gclk));
	jdff dff_B_lZRLbIjL6_2(.din(w_dff_B_Ho41pmSb0_2),.dout(w_dff_B_lZRLbIjL6_2),.clk(gclk));
	jdff dff_B_eiNf6T714_2(.din(w_dff_B_lZRLbIjL6_2),.dout(w_dff_B_eiNf6T714_2),.clk(gclk));
	jdff dff_B_kNqznUS58_2(.din(w_dff_B_eiNf6T714_2),.dout(w_dff_B_kNqznUS58_2),.clk(gclk));
	jdff dff_B_gZ2N9WDJ5_2(.din(w_dff_B_kNqznUS58_2),.dout(w_dff_B_gZ2N9WDJ5_2),.clk(gclk));
	jdff dff_B_NjJntgbw3_2(.din(w_dff_B_gZ2N9WDJ5_2),.dout(w_dff_B_NjJntgbw3_2),.clk(gclk));
	jdff dff_B_E0WdK6zA3_2(.din(w_dff_B_NjJntgbw3_2),.dout(w_dff_B_E0WdK6zA3_2),.clk(gclk));
	jdff dff_B_RmcELb6R1_2(.din(w_dff_B_E0WdK6zA3_2),.dout(w_dff_B_RmcELb6R1_2),.clk(gclk));
	jdff dff_B_HgmlUmpy4_2(.din(w_dff_B_RmcELb6R1_2),.dout(w_dff_B_HgmlUmpy4_2),.clk(gclk));
	jdff dff_B_8zHZDOVm9_2(.din(w_dff_B_HgmlUmpy4_2),.dout(w_dff_B_8zHZDOVm9_2),.clk(gclk));
	jdff dff_B_csGE3hON3_2(.din(w_dff_B_8zHZDOVm9_2),.dout(w_dff_B_csGE3hON3_2),.clk(gclk));
	jdff dff_B_kQp97ZQk9_2(.din(w_dff_B_csGE3hON3_2),.dout(w_dff_B_kQp97ZQk9_2),.clk(gclk));
	jdff dff_B_FsmNUmCF8_2(.din(w_dff_B_kQp97ZQk9_2),.dout(w_dff_B_FsmNUmCF8_2),.clk(gclk));
	jdff dff_B_DGMFsyGd6_2(.din(w_dff_B_FsmNUmCF8_2),.dout(w_dff_B_DGMFsyGd6_2),.clk(gclk));
	jdff dff_B_fPhm7dyX2_2(.din(w_dff_B_DGMFsyGd6_2),.dout(w_dff_B_fPhm7dyX2_2),.clk(gclk));
	jdff dff_B_9guEDIXx9_2(.din(w_dff_B_fPhm7dyX2_2),.dout(w_dff_B_9guEDIXx9_2),.clk(gclk));
	jdff dff_B_KmDdxCba2_2(.din(w_dff_B_9guEDIXx9_2),.dout(w_dff_B_KmDdxCba2_2),.clk(gclk));
	jdff dff_B_XNDjEVCQ2_2(.din(w_dff_B_KmDdxCba2_2),.dout(w_dff_B_XNDjEVCQ2_2),.clk(gclk));
	jdff dff_B_BCoDk1Ig3_2(.din(w_dff_B_XNDjEVCQ2_2),.dout(w_dff_B_BCoDk1Ig3_2),.clk(gclk));
	jdff dff_B_aPpzmYqb7_2(.din(w_dff_B_BCoDk1Ig3_2),.dout(w_dff_B_aPpzmYqb7_2),.clk(gclk));
	jdff dff_B_2wQQ5OD01_2(.din(w_dff_B_aPpzmYqb7_2),.dout(w_dff_B_2wQQ5OD01_2),.clk(gclk));
	jdff dff_B_h2aLBisn5_2(.din(w_dff_B_2wQQ5OD01_2),.dout(w_dff_B_h2aLBisn5_2),.clk(gclk));
	jdff dff_B_jQwbdlRs4_2(.din(w_dff_B_h2aLBisn5_2),.dout(w_dff_B_jQwbdlRs4_2),.clk(gclk));
	jdff dff_B_h5EXYLZM4_2(.din(w_dff_B_jQwbdlRs4_2),.dout(w_dff_B_h5EXYLZM4_2),.clk(gclk));
	jdff dff_B_KKv14GYh4_2(.din(w_dff_B_h5EXYLZM4_2),.dout(w_dff_B_KKv14GYh4_2),.clk(gclk));
	jdff dff_B_aLg9hG0Z2_2(.din(w_dff_B_KKv14GYh4_2),.dout(w_dff_B_aLg9hG0Z2_2),.clk(gclk));
	jdff dff_B_vmd2Q5af3_2(.din(w_dff_B_aLg9hG0Z2_2),.dout(w_dff_B_vmd2Q5af3_2),.clk(gclk));
	jdff dff_B_hQc1PwNP7_2(.din(w_dff_B_vmd2Q5af3_2),.dout(w_dff_B_hQc1PwNP7_2),.clk(gclk));
	jdff dff_B_z5QIOJ2o2_2(.din(w_dff_B_hQc1PwNP7_2),.dout(w_dff_B_z5QIOJ2o2_2),.clk(gclk));
	jdff dff_B_qaN1el2k1_2(.din(n1744),.dout(w_dff_B_qaN1el2k1_2),.clk(gclk));
	jdff dff_B_wUP8miuQ0_2(.din(w_dff_B_qaN1el2k1_2),.dout(w_dff_B_wUP8miuQ0_2),.clk(gclk));
	jdff dff_B_xgifIYVK2_2(.din(w_dff_B_wUP8miuQ0_2),.dout(w_dff_B_xgifIYVK2_2),.clk(gclk));
	jdff dff_B_YqcuE0Aq2_2(.din(w_dff_B_xgifIYVK2_2),.dout(w_dff_B_YqcuE0Aq2_2),.clk(gclk));
	jdff dff_B_at3yg0Wa3_2(.din(w_dff_B_YqcuE0Aq2_2),.dout(w_dff_B_at3yg0Wa3_2),.clk(gclk));
	jdff dff_B_calvw9OX5_2(.din(w_dff_B_at3yg0Wa3_2),.dout(w_dff_B_calvw9OX5_2),.clk(gclk));
	jdff dff_B_FtpxofnM3_2(.din(w_dff_B_calvw9OX5_2),.dout(w_dff_B_FtpxofnM3_2),.clk(gclk));
	jdff dff_B_blQ0iAMY6_2(.din(w_dff_B_FtpxofnM3_2),.dout(w_dff_B_blQ0iAMY6_2),.clk(gclk));
	jdff dff_B_ykb41ZJk3_2(.din(w_dff_B_blQ0iAMY6_2),.dout(w_dff_B_ykb41ZJk3_2),.clk(gclk));
	jdff dff_B_HQOsVYbb9_2(.din(w_dff_B_ykb41ZJk3_2),.dout(w_dff_B_HQOsVYbb9_2),.clk(gclk));
	jdff dff_B_Zqun5X929_2(.din(w_dff_B_HQOsVYbb9_2),.dout(w_dff_B_Zqun5X929_2),.clk(gclk));
	jdff dff_B_8bNObTPf5_2(.din(w_dff_B_Zqun5X929_2),.dout(w_dff_B_8bNObTPf5_2),.clk(gclk));
	jdff dff_B_TEvqXDKt6_2(.din(w_dff_B_8bNObTPf5_2),.dout(w_dff_B_TEvqXDKt6_2),.clk(gclk));
	jdff dff_B_nkr8ubmc5_2(.din(w_dff_B_TEvqXDKt6_2),.dout(w_dff_B_nkr8ubmc5_2),.clk(gclk));
	jdff dff_B_Q2hQ9NlK8_2(.din(w_dff_B_nkr8ubmc5_2),.dout(w_dff_B_Q2hQ9NlK8_2),.clk(gclk));
	jdff dff_B_6Qqdk2Lk0_2(.din(w_dff_B_Q2hQ9NlK8_2),.dout(w_dff_B_6Qqdk2Lk0_2),.clk(gclk));
	jdff dff_B_YqCrXgWI6_2(.din(w_dff_B_6Qqdk2Lk0_2),.dout(w_dff_B_YqCrXgWI6_2),.clk(gclk));
	jdff dff_B_NFPIrlfV1_2(.din(w_dff_B_YqCrXgWI6_2),.dout(w_dff_B_NFPIrlfV1_2),.clk(gclk));
	jdff dff_B_RseZyUiX8_2(.din(w_dff_B_NFPIrlfV1_2),.dout(w_dff_B_RseZyUiX8_2),.clk(gclk));
	jdff dff_B_k6nek2va8_2(.din(w_dff_B_RseZyUiX8_2),.dout(w_dff_B_k6nek2va8_2),.clk(gclk));
	jdff dff_B_XgHjjRfO2_2(.din(w_dff_B_k6nek2va8_2),.dout(w_dff_B_XgHjjRfO2_2),.clk(gclk));
	jdff dff_B_1Z3dvCvs0_2(.din(w_dff_B_XgHjjRfO2_2),.dout(w_dff_B_1Z3dvCvs0_2),.clk(gclk));
	jdff dff_B_V197taw22_2(.din(w_dff_B_1Z3dvCvs0_2),.dout(w_dff_B_V197taw22_2),.clk(gclk));
	jdff dff_B_PVwL3f5e5_2(.din(w_dff_B_V197taw22_2),.dout(w_dff_B_PVwL3f5e5_2),.clk(gclk));
	jdff dff_B_poW69XPH2_2(.din(w_dff_B_PVwL3f5e5_2),.dout(w_dff_B_poW69XPH2_2),.clk(gclk));
	jdff dff_B_ZFnKktzJ7_2(.din(w_dff_B_poW69XPH2_2),.dout(w_dff_B_ZFnKktzJ7_2),.clk(gclk));
	jdff dff_B_B44wpiev2_2(.din(w_dff_B_ZFnKktzJ7_2),.dout(w_dff_B_B44wpiev2_2),.clk(gclk));
	jdff dff_B_PcvOIpH55_2(.din(w_dff_B_B44wpiev2_2),.dout(w_dff_B_PcvOIpH55_2),.clk(gclk));
	jdff dff_B_LQ1euEiA0_2(.din(w_dff_B_PcvOIpH55_2),.dout(w_dff_B_LQ1euEiA0_2),.clk(gclk));
	jdff dff_B_uX5JAVHG6_2(.din(w_dff_B_LQ1euEiA0_2),.dout(w_dff_B_uX5JAVHG6_2),.clk(gclk));
	jdff dff_B_EhALhOGY7_2(.din(w_dff_B_uX5JAVHG6_2),.dout(w_dff_B_EhALhOGY7_2),.clk(gclk));
	jdff dff_B_IA2fbPFR6_2(.din(w_dff_B_EhALhOGY7_2),.dout(w_dff_B_IA2fbPFR6_2),.clk(gclk));
	jdff dff_B_y9OtsbHg3_2(.din(w_dff_B_IA2fbPFR6_2),.dout(w_dff_B_y9OtsbHg3_2),.clk(gclk));
	jdff dff_B_foVNVH4X5_2(.din(w_dff_B_y9OtsbHg3_2),.dout(w_dff_B_foVNVH4X5_2),.clk(gclk));
	jdff dff_B_bqTe6Lzj1_2(.din(w_dff_B_foVNVH4X5_2),.dout(w_dff_B_bqTe6Lzj1_2),.clk(gclk));
	jdff dff_B_c0Qs8dBf7_2(.din(n1743),.dout(w_dff_B_c0Qs8dBf7_2),.clk(gclk));
	jdff dff_B_IzfRDnTa7_1(.din(n1741),.dout(w_dff_B_IzfRDnTa7_1),.clk(gclk));
	jdff dff_B_Zb99ZdHS8_2(.din(n1699),.dout(w_dff_B_Zb99ZdHS8_2),.clk(gclk));
	jdff dff_B_NgIO3hqL1_2(.din(w_dff_B_Zb99ZdHS8_2),.dout(w_dff_B_NgIO3hqL1_2),.clk(gclk));
	jdff dff_B_qQrhE51o0_2(.din(w_dff_B_NgIO3hqL1_2),.dout(w_dff_B_qQrhE51o0_2),.clk(gclk));
	jdff dff_B_9Y5WYIJl9_2(.din(w_dff_B_qQrhE51o0_2),.dout(w_dff_B_9Y5WYIJl9_2),.clk(gclk));
	jdff dff_B_OVknh3e76_2(.din(w_dff_B_9Y5WYIJl9_2),.dout(w_dff_B_OVknh3e76_2),.clk(gclk));
	jdff dff_B_7eFjvere8_2(.din(w_dff_B_OVknh3e76_2),.dout(w_dff_B_7eFjvere8_2),.clk(gclk));
	jdff dff_B_IEnjttNr2_2(.din(w_dff_B_7eFjvere8_2),.dout(w_dff_B_IEnjttNr2_2),.clk(gclk));
	jdff dff_B_Hg6inLPI1_2(.din(w_dff_B_IEnjttNr2_2),.dout(w_dff_B_Hg6inLPI1_2),.clk(gclk));
	jdff dff_B_Cx32MKBs0_2(.din(w_dff_B_Hg6inLPI1_2),.dout(w_dff_B_Cx32MKBs0_2),.clk(gclk));
	jdff dff_B_dBCK1NDD0_2(.din(w_dff_B_Cx32MKBs0_2),.dout(w_dff_B_dBCK1NDD0_2),.clk(gclk));
	jdff dff_B_JB2dtFdm3_2(.din(w_dff_B_dBCK1NDD0_2),.dout(w_dff_B_JB2dtFdm3_2),.clk(gclk));
	jdff dff_B_WDkpkpuJ9_2(.din(w_dff_B_JB2dtFdm3_2),.dout(w_dff_B_WDkpkpuJ9_2),.clk(gclk));
	jdff dff_B_lhIgNy631_2(.din(w_dff_B_WDkpkpuJ9_2),.dout(w_dff_B_lhIgNy631_2),.clk(gclk));
	jdff dff_B_5LGLQcwG5_2(.din(w_dff_B_lhIgNy631_2),.dout(w_dff_B_5LGLQcwG5_2),.clk(gclk));
	jdff dff_B_0EqYBEXj0_2(.din(w_dff_B_5LGLQcwG5_2),.dout(w_dff_B_0EqYBEXj0_2),.clk(gclk));
	jdff dff_B_LxZ5clYQ8_2(.din(w_dff_B_0EqYBEXj0_2),.dout(w_dff_B_LxZ5clYQ8_2),.clk(gclk));
	jdff dff_B_2JJiNf1a2_2(.din(w_dff_B_LxZ5clYQ8_2),.dout(w_dff_B_2JJiNf1a2_2),.clk(gclk));
	jdff dff_B_DIhKgkga6_2(.din(w_dff_B_2JJiNf1a2_2),.dout(w_dff_B_DIhKgkga6_2),.clk(gclk));
	jdff dff_B_6suNxC6B7_2(.din(w_dff_B_DIhKgkga6_2),.dout(w_dff_B_6suNxC6B7_2),.clk(gclk));
	jdff dff_B_Su5k1gae6_2(.din(w_dff_B_6suNxC6B7_2),.dout(w_dff_B_Su5k1gae6_2),.clk(gclk));
	jdff dff_B_PffExo7g1_2(.din(w_dff_B_Su5k1gae6_2),.dout(w_dff_B_PffExo7g1_2),.clk(gclk));
	jdff dff_B_kKG2OM7H0_2(.din(w_dff_B_PffExo7g1_2),.dout(w_dff_B_kKG2OM7H0_2),.clk(gclk));
	jdff dff_B_O9sxoRsM0_2(.din(w_dff_B_kKG2OM7H0_2),.dout(w_dff_B_O9sxoRsM0_2),.clk(gclk));
	jdff dff_B_B6nsp8aL6_2(.din(w_dff_B_O9sxoRsM0_2),.dout(w_dff_B_B6nsp8aL6_2),.clk(gclk));
	jdff dff_B_HLwZpeXP4_2(.din(w_dff_B_B6nsp8aL6_2),.dout(w_dff_B_HLwZpeXP4_2),.clk(gclk));
	jdff dff_B_Iz2iBD161_2(.din(w_dff_B_HLwZpeXP4_2),.dout(w_dff_B_Iz2iBD161_2),.clk(gclk));
	jdff dff_B_erGLMVOC2_2(.din(w_dff_B_Iz2iBD161_2),.dout(w_dff_B_erGLMVOC2_2),.clk(gclk));
	jdff dff_B_ffsAHrzV7_2(.din(w_dff_B_erGLMVOC2_2),.dout(w_dff_B_ffsAHrzV7_2),.clk(gclk));
	jdff dff_B_YQ04Rc9S9_2(.din(w_dff_B_ffsAHrzV7_2),.dout(w_dff_B_YQ04Rc9S9_2),.clk(gclk));
	jdff dff_B_Lo7HHNol8_2(.din(w_dff_B_YQ04Rc9S9_2),.dout(w_dff_B_Lo7HHNol8_2),.clk(gclk));
	jdff dff_B_W0Tf1de92_2(.din(w_dff_B_Lo7HHNol8_2),.dout(w_dff_B_W0Tf1de92_2),.clk(gclk));
	jdff dff_B_x5ZwqFSH7_2(.din(w_dff_B_W0Tf1de92_2),.dout(w_dff_B_x5ZwqFSH7_2),.clk(gclk));
	jdff dff_B_GUFsXUGN2_2(.din(w_dff_B_x5ZwqFSH7_2),.dout(w_dff_B_GUFsXUGN2_2),.clk(gclk));
	jdff dff_B_PvsmpJBm4_1(.din(n1705),.dout(w_dff_B_PvsmpJBm4_1),.clk(gclk));
	jdff dff_B_YErMqfjS7_1(.din(w_dff_B_PvsmpJBm4_1),.dout(w_dff_B_YErMqfjS7_1),.clk(gclk));
	jdff dff_B_qTDl1epY8_2(.din(n1704),.dout(w_dff_B_qTDl1epY8_2),.clk(gclk));
	jdff dff_B_dDsdxMjD5_2(.din(w_dff_B_qTDl1epY8_2),.dout(w_dff_B_dDsdxMjD5_2),.clk(gclk));
	jdff dff_B_Qzf46XOn9_2(.din(w_dff_B_dDsdxMjD5_2),.dout(w_dff_B_Qzf46XOn9_2),.clk(gclk));
	jdff dff_B_eLYoqyXj5_2(.din(w_dff_B_Qzf46XOn9_2),.dout(w_dff_B_eLYoqyXj5_2),.clk(gclk));
	jdff dff_B_XJowFD5f6_2(.din(w_dff_B_eLYoqyXj5_2),.dout(w_dff_B_XJowFD5f6_2),.clk(gclk));
	jdff dff_B_AaeF6JTK5_2(.din(w_dff_B_XJowFD5f6_2),.dout(w_dff_B_AaeF6JTK5_2),.clk(gclk));
	jdff dff_B_lGbbPq324_2(.din(w_dff_B_AaeF6JTK5_2),.dout(w_dff_B_lGbbPq324_2),.clk(gclk));
	jdff dff_B_hFDsIOkN8_2(.din(w_dff_B_lGbbPq324_2),.dout(w_dff_B_hFDsIOkN8_2),.clk(gclk));
	jdff dff_B_MEqaN5ff8_2(.din(w_dff_B_hFDsIOkN8_2),.dout(w_dff_B_MEqaN5ff8_2),.clk(gclk));
	jdff dff_B_aFCi0B621_2(.din(w_dff_B_MEqaN5ff8_2),.dout(w_dff_B_aFCi0B621_2),.clk(gclk));
	jdff dff_B_UxLDaFzC9_2(.din(w_dff_B_aFCi0B621_2),.dout(w_dff_B_UxLDaFzC9_2),.clk(gclk));
	jdff dff_B_knTuofbS1_2(.din(w_dff_B_UxLDaFzC9_2),.dout(w_dff_B_knTuofbS1_2),.clk(gclk));
	jdff dff_B_LydvIIcl3_2(.din(w_dff_B_knTuofbS1_2),.dout(w_dff_B_LydvIIcl3_2),.clk(gclk));
	jdff dff_B_WdvVUIfB1_2(.din(w_dff_B_LydvIIcl3_2),.dout(w_dff_B_WdvVUIfB1_2),.clk(gclk));
	jdff dff_B_rYtbfWX81_2(.din(w_dff_B_WdvVUIfB1_2),.dout(w_dff_B_rYtbfWX81_2),.clk(gclk));
	jdff dff_B_nZRIjCSh5_2(.din(w_dff_B_rYtbfWX81_2),.dout(w_dff_B_nZRIjCSh5_2),.clk(gclk));
	jdff dff_B_aE4QKcva3_2(.din(w_dff_B_nZRIjCSh5_2),.dout(w_dff_B_aE4QKcva3_2),.clk(gclk));
	jdff dff_B_PM4EtVMa2_2(.din(w_dff_B_aE4QKcva3_2),.dout(w_dff_B_PM4EtVMa2_2),.clk(gclk));
	jdff dff_B_20TzXt6y4_2(.din(w_dff_B_PM4EtVMa2_2),.dout(w_dff_B_20TzXt6y4_2),.clk(gclk));
	jdff dff_B_v29Brma90_2(.din(w_dff_B_20TzXt6y4_2),.dout(w_dff_B_v29Brma90_2),.clk(gclk));
	jdff dff_B_lpNCN7Zg9_2(.din(w_dff_B_v29Brma90_2),.dout(w_dff_B_lpNCN7Zg9_2),.clk(gclk));
	jdff dff_B_n0dwKKlZ7_2(.din(w_dff_B_lpNCN7Zg9_2),.dout(w_dff_B_n0dwKKlZ7_2),.clk(gclk));
	jdff dff_B_rL8TNgld4_2(.din(w_dff_B_n0dwKKlZ7_2),.dout(w_dff_B_rL8TNgld4_2),.clk(gclk));
	jdff dff_B_fIg1iSPN4_2(.din(w_dff_B_rL8TNgld4_2),.dout(w_dff_B_fIg1iSPN4_2),.clk(gclk));
	jdff dff_B_Ze42DfCH0_2(.din(w_dff_B_fIg1iSPN4_2),.dout(w_dff_B_Ze42DfCH0_2),.clk(gclk));
	jdff dff_B_QC5OYXZP7_2(.din(w_dff_B_Ze42DfCH0_2),.dout(w_dff_B_QC5OYXZP7_2),.clk(gclk));
	jdff dff_B_peGCjqIh5_2(.din(w_dff_B_QC5OYXZP7_2),.dout(w_dff_B_peGCjqIh5_2),.clk(gclk));
	jdff dff_B_rNmU3GZY7_2(.din(w_dff_B_peGCjqIh5_2),.dout(w_dff_B_rNmU3GZY7_2),.clk(gclk));
	jdff dff_B_JkyxggJK2_2(.din(w_dff_B_rNmU3GZY7_2),.dout(w_dff_B_JkyxggJK2_2),.clk(gclk));
	jdff dff_B_mXwsCmDM5_2(.din(w_dff_B_JkyxggJK2_2),.dout(w_dff_B_mXwsCmDM5_2),.clk(gclk));
	jdff dff_B_OUwHMjED9_2(.din(n1703),.dout(w_dff_B_OUwHMjED9_2),.clk(gclk));
	jdff dff_B_xtLV87IE7_2(.din(w_dff_B_OUwHMjED9_2),.dout(w_dff_B_xtLV87IE7_2),.clk(gclk));
	jdff dff_B_aJYdTGTJ0_2(.din(w_dff_B_xtLV87IE7_2),.dout(w_dff_B_aJYdTGTJ0_2),.clk(gclk));
	jdff dff_B_v1Pr301H3_2(.din(w_dff_B_aJYdTGTJ0_2),.dout(w_dff_B_v1Pr301H3_2),.clk(gclk));
	jdff dff_B_D59cdu1h4_2(.din(w_dff_B_v1Pr301H3_2),.dout(w_dff_B_D59cdu1h4_2),.clk(gclk));
	jdff dff_B_BMC5zDa01_2(.din(w_dff_B_D59cdu1h4_2),.dout(w_dff_B_BMC5zDa01_2),.clk(gclk));
	jdff dff_B_LPf4mr7G3_2(.din(w_dff_B_BMC5zDa01_2),.dout(w_dff_B_LPf4mr7G3_2),.clk(gclk));
	jdff dff_B_K6IO6Mxv3_2(.din(w_dff_B_LPf4mr7G3_2),.dout(w_dff_B_K6IO6Mxv3_2),.clk(gclk));
	jdff dff_B_ruFLtfx99_2(.din(w_dff_B_K6IO6Mxv3_2),.dout(w_dff_B_ruFLtfx99_2),.clk(gclk));
	jdff dff_B_3OtWJJV04_2(.din(w_dff_B_ruFLtfx99_2),.dout(w_dff_B_3OtWJJV04_2),.clk(gclk));
	jdff dff_B_beJocVUY1_2(.din(w_dff_B_3OtWJJV04_2),.dout(w_dff_B_beJocVUY1_2),.clk(gclk));
	jdff dff_B_3TqRlnEJ4_2(.din(w_dff_B_beJocVUY1_2),.dout(w_dff_B_3TqRlnEJ4_2),.clk(gclk));
	jdff dff_B_FWq85ip66_2(.din(w_dff_B_3TqRlnEJ4_2),.dout(w_dff_B_FWq85ip66_2),.clk(gclk));
	jdff dff_B_LUNRbAaB4_2(.din(w_dff_B_FWq85ip66_2),.dout(w_dff_B_LUNRbAaB4_2),.clk(gclk));
	jdff dff_B_OLtQc3iX0_2(.din(w_dff_B_LUNRbAaB4_2),.dout(w_dff_B_OLtQc3iX0_2),.clk(gclk));
	jdff dff_B_vnNLjbK79_2(.din(w_dff_B_OLtQc3iX0_2),.dout(w_dff_B_vnNLjbK79_2),.clk(gclk));
	jdff dff_B_ktNM0r6b7_2(.din(w_dff_B_vnNLjbK79_2),.dout(w_dff_B_ktNM0r6b7_2),.clk(gclk));
	jdff dff_B_Nnb4YZRZ2_2(.din(w_dff_B_ktNM0r6b7_2),.dout(w_dff_B_Nnb4YZRZ2_2),.clk(gclk));
	jdff dff_B_ojFpsxO98_2(.din(w_dff_B_Nnb4YZRZ2_2),.dout(w_dff_B_ojFpsxO98_2),.clk(gclk));
	jdff dff_B_IBCwZT5t5_2(.din(w_dff_B_ojFpsxO98_2),.dout(w_dff_B_IBCwZT5t5_2),.clk(gclk));
	jdff dff_B_Pt0nCbGD5_2(.din(w_dff_B_IBCwZT5t5_2),.dout(w_dff_B_Pt0nCbGD5_2),.clk(gclk));
	jdff dff_B_y7vLdVIX1_2(.din(w_dff_B_Pt0nCbGD5_2),.dout(w_dff_B_y7vLdVIX1_2),.clk(gclk));
	jdff dff_B_4CbKcEhX3_2(.din(w_dff_B_y7vLdVIX1_2),.dout(w_dff_B_4CbKcEhX3_2),.clk(gclk));
	jdff dff_B_XCzWQrqQ6_2(.din(w_dff_B_4CbKcEhX3_2),.dout(w_dff_B_XCzWQrqQ6_2),.clk(gclk));
	jdff dff_B_K4p38FV20_2(.din(w_dff_B_XCzWQrqQ6_2),.dout(w_dff_B_K4p38FV20_2),.clk(gclk));
	jdff dff_B_zhm2YRNX7_2(.din(w_dff_B_K4p38FV20_2),.dout(w_dff_B_zhm2YRNX7_2),.clk(gclk));
	jdff dff_B_aa7M3sTb8_2(.din(w_dff_B_zhm2YRNX7_2),.dout(w_dff_B_aa7M3sTb8_2),.clk(gclk));
	jdff dff_B_R1sPw8fa1_2(.din(w_dff_B_aa7M3sTb8_2),.dout(w_dff_B_R1sPw8fa1_2),.clk(gclk));
	jdff dff_B_ZKa8ociC4_2(.din(w_dff_B_R1sPw8fa1_2),.dout(w_dff_B_ZKa8ociC4_2),.clk(gclk));
	jdff dff_B_c63vPWyR8_2(.din(w_dff_B_ZKa8ociC4_2),.dout(w_dff_B_c63vPWyR8_2),.clk(gclk));
	jdff dff_B_xLB5aAUQ2_2(.din(w_dff_B_c63vPWyR8_2),.dout(w_dff_B_xLB5aAUQ2_2),.clk(gclk));
	jdff dff_B_QZUrIAZs9_2(.din(w_dff_B_xLB5aAUQ2_2),.dout(w_dff_B_QZUrIAZs9_2),.clk(gclk));
	jdff dff_B_qSMUqC6J3_2(.din(n1702),.dout(w_dff_B_qSMUqC6J3_2),.clk(gclk));
	jdff dff_B_VbSDAllf5_1(.din(n1700),.dout(w_dff_B_VbSDAllf5_1),.clk(gclk));
	jdff dff_B_hTrstGvu4_2(.din(n1648),.dout(w_dff_B_hTrstGvu4_2),.clk(gclk));
	jdff dff_B_RTlQfiI71_2(.din(w_dff_B_hTrstGvu4_2),.dout(w_dff_B_RTlQfiI71_2),.clk(gclk));
	jdff dff_B_gP53vt9F2_2(.din(w_dff_B_RTlQfiI71_2),.dout(w_dff_B_gP53vt9F2_2),.clk(gclk));
	jdff dff_B_Z5Vjm5Mo1_2(.din(w_dff_B_gP53vt9F2_2),.dout(w_dff_B_Z5Vjm5Mo1_2),.clk(gclk));
	jdff dff_B_vARs2y1j7_2(.din(w_dff_B_Z5Vjm5Mo1_2),.dout(w_dff_B_vARs2y1j7_2),.clk(gclk));
	jdff dff_B_5xtCwI856_2(.din(w_dff_B_vARs2y1j7_2),.dout(w_dff_B_5xtCwI856_2),.clk(gclk));
	jdff dff_B_bR7vL1k10_2(.din(w_dff_B_5xtCwI856_2),.dout(w_dff_B_bR7vL1k10_2),.clk(gclk));
	jdff dff_B_CTS5lpnv8_2(.din(w_dff_B_bR7vL1k10_2),.dout(w_dff_B_CTS5lpnv8_2),.clk(gclk));
	jdff dff_B_StKDVNTE2_2(.din(w_dff_B_CTS5lpnv8_2),.dout(w_dff_B_StKDVNTE2_2),.clk(gclk));
	jdff dff_B_P7lCUDBB5_2(.din(w_dff_B_StKDVNTE2_2),.dout(w_dff_B_P7lCUDBB5_2),.clk(gclk));
	jdff dff_B_pII7MEJH8_2(.din(w_dff_B_P7lCUDBB5_2),.dout(w_dff_B_pII7MEJH8_2),.clk(gclk));
	jdff dff_B_m5GOJuzq7_2(.din(w_dff_B_pII7MEJH8_2),.dout(w_dff_B_m5GOJuzq7_2),.clk(gclk));
	jdff dff_B_kJtpIqHu9_2(.din(w_dff_B_m5GOJuzq7_2),.dout(w_dff_B_kJtpIqHu9_2),.clk(gclk));
	jdff dff_B_ZISNOnRE6_2(.din(w_dff_B_kJtpIqHu9_2),.dout(w_dff_B_ZISNOnRE6_2),.clk(gclk));
	jdff dff_B_OcpfefGm4_2(.din(w_dff_B_ZISNOnRE6_2),.dout(w_dff_B_OcpfefGm4_2),.clk(gclk));
	jdff dff_B_OOQ7tIpY5_2(.din(w_dff_B_OcpfefGm4_2),.dout(w_dff_B_OOQ7tIpY5_2),.clk(gclk));
	jdff dff_B_vEivhFuV5_2(.din(w_dff_B_OOQ7tIpY5_2),.dout(w_dff_B_vEivhFuV5_2),.clk(gclk));
	jdff dff_B_66mgbrko4_2(.din(w_dff_B_vEivhFuV5_2),.dout(w_dff_B_66mgbrko4_2),.clk(gclk));
	jdff dff_B_XOyCFZ7v3_2(.din(w_dff_B_66mgbrko4_2),.dout(w_dff_B_XOyCFZ7v3_2),.clk(gclk));
	jdff dff_B_kApYDfkX9_2(.din(w_dff_B_XOyCFZ7v3_2),.dout(w_dff_B_kApYDfkX9_2),.clk(gclk));
	jdff dff_B_bakpFhan4_2(.din(w_dff_B_kApYDfkX9_2),.dout(w_dff_B_bakpFhan4_2),.clk(gclk));
	jdff dff_B_HskodKWb7_2(.din(w_dff_B_bakpFhan4_2),.dout(w_dff_B_HskodKWb7_2),.clk(gclk));
	jdff dff_B_uY2M1oMY0_2(.din(w_dff_B_HskodKWb7_2),.dout(w_dff_B_uY2M1oMY0_2),.clk(gclk));
	jdff dff_B_BKQkdCnk2_2(.din(w_dff_B_uY2M1oMY0_2),.dout(w_dff_B_BKQkdCnk2_2),.clk(gclk));
	jdff dff_B_nv58PPcL1_2(.din(w_dff_B_BKQkdCnk2_2),.dout(w_dff_B_nv58PPcL1_2),.clk(gclk));
	jdff dff_B_mR9KjR2E5_2(.din(w_dff_B_nv58PPcL1_2),.dout(w_dff_B_mR9KjR2E5_2),.clk(gclk));
	jdff dff_B_QF8iOlUM9_2(.din(w_dff_B_mR9KjR2E5_2),.dout(w_dff_B_QF8iOlUM9_2),.clk(gclk));
	jdff dff_B_NEN9KgV76_2(.din(w_dff_B_QF8iOlUM9_2),.dout(w_dff_B_NEN9KgV76_2),.clk(gclk));
	jdff dff_B_vCxmitVU2_2(.din(w_dff_B_NEN9KgV76_2),.dout(w_dff_B_vCxmitVU2_2),.clk(gclk));
	jdff dff_B_5vAg64vY8_2(.din(w_dff_B_vCxmitVU2_2),.dout(w_dff_B_5vAg64vY8_2),.clk(gclk));
	jdff dff_B_bKEYKbbV9_1(.din(n1654),.dout(w_dff_B_bKEYKbbV9_1),.clk(gclk));
	jdff dff_B_3KAZd9Je8_1(.din(w_dff_B_bKEYKbbV9_1),.dout(w_dff_B_3KAZd9Je8_1),.clk(gclk));
	jdff dff_B_Vaq02DPH7_2(.din(n1653),.dout(w_dff_B_Vaq02DPH7_2),.clk(gclk));
	jdff dff_B_Bnd9QY6c3_2(.din(w_dff_B_Vaq02DPH7_2),.dout(w_dff_B_Bnd9QY6c3_2),.clk(gclk));
	jdff dff_B_oDdsBWCC3_2(.din(w_dff_B_Bnd9QY6c3_2),.dout(w_dff_B_oDdsBWCC3_2),.clk(gclk));
	jdff dff_B_XTsRPkOW9_2(.din(w_dff_B_oDdsBWCC3_2),.dout(w_dff_B_XTsRPkOW9_2),.clk(gclk));
	jdff dff_B_QJMmha5K4_2(.din(w_dff_B_XTsRPkOW9_2),.dout(w_dff_B_QJMmha5K4_2),.clk(gclk));
	jdff dff_B_v9qSeM8R5_2(.din(w_dff_B_QJMmha5K4_2),.dout(w_dff_B_v9qSeM8R5_2),.clk(gclk));
	jdff dff_B_r721UY4v2_2(.din(w_dff_B_v9qSeM8R5_2),.dout(w_dff_B_r721UY4v2_2),.clk(gclk));
	jdff dff_B_NS5UwBBF0_2(.din(w_dff_B_r721UY4v2_2),.dout(w_dff_B_NS5UwBBF0_2),.clk(gclk));
	jdff dff_B_3LJWnYas0_2(.din(w_dff_B_NS5UwBBF0_2),.dout(w_dff_B_3LJWnYas0_2),.clk(gclk));
	jdff dff_B_e273UyQ47_2(.din(w_dff_B_3LJWnYas0_2),.dout(w_dff_B_e273UyQ47_2),.clk(gclk));
	jdff dff_B_sxlwXp1o0_2(.din(w_dff_B_e273UyQ47_2),.dout(w_dff_B_sxlwXp1o0_2),.clk(gclk));
	jdff dff_B_6ypBymCa2_2(.din(w_dff_B_sxlwXp1o0_2),.dout(w_dff_B_6ypBymCa2_2),.clk(gclk));
	jdff dff_B_PkEeP02S0_2(.din(w_dff_B_6ypBymCa2_2),.dout(w_dff_B_PkEeP02S0_2),.clk(gclk));
	jdff dff_B_k5xa1wZ94_2(.din(w_dff_B_PkEeP02S0_2),.dout(w_dff_B_k5xa1wZ94_2),.clk(gclk));
	jdff dff_B_gNcwLOgK5_2(.din(w_dff_B_k5xa1wZ94_2),.dout(w_dff_B_gNcwLOgK5_2),.clk(gclk));
	jdff dff_B_Ux6I4cQt8_2(.din(w_dff_B_gNcwLOgK5_2),.dout(w_dff_B_Ux6I4cQt8_2),.clk(gclk));
	jdff dff_B_yL9mW64V9_2(.din(w_dff_B_Ux6I4cQt8_2),.dout(w_dff_B_yL9mW64V9_2),.clk(gclk));
	jdff dff_B_cpQSAWmr5_2(.din(w_dff_B_yL9mW64V9_2),.dout(w_dff_B_cpQSAWmr5_2),.clk(gclk));
	jdff dff_B_7EwULnyV2_2(.din(w_dff_B_cpQSAWmr5_2),.dout(w_dff_B_7EwULnyV2_2),.clk(gclk));
	jdff dff_B_41bdJH389_2(.din(w_dff_B_7EwULnyV2_2),.dout(w_dff_B_41bdJH389_2),.clk(gclk));
	jdff dff_B_J5o1CbXZ4_2(.din(w_dff_B_41bdJH389_2),.dout(w_dff_B_J5o1CbXZ4_2),.clk(gclk));
	jdff dff_B_mnS48AB18_2(.din(w_dff_B_J5o1CbXZ4_2),.dout(w_dff_B_mnS48AB18_2),.clk(gclk));
	jdff dff_B_QanCfR3c3_2(.din(w_dff_B_mnS48AB18_2),.dout(w_dff_B_QanCfR3c3_2),.clk(gclk));
	jdff dff_B_eef1ZK2M2_2(.din(w_dff_B_QanCfR3c3_2),.dout(w_dff_B_eef1ZK2M2_2),.clk(gclk));
	jdff dff_B_1w2h16bM3_2(.din(w_dff_B_eef1ZK2M2_2),.dout(w_dff_B_1w2h16bM3_2),.clk(gclk));
	jdff dff_B_nVvhYrmC6_2(.din(w_dff_B_1w2h16bM3_2),.dout(w_dff_B_nVvhYrmC6_2),.clk(gclk));
	jdff dff_B_bsop8f2T8_2(.din(w_dff_B_nVvhYrmC6_2),.dout(w_dff_B_bsop8f2T8_2),.clk(gclk));
	jdff dff_B_gRduZacn2_2(.din(n1652),.dout(w_dff_B_gRduZacn2_2),.clk(gclk));
	jdff dff_B_FYGPnNpu9_2(.din(w_dff_B_gRduZacn2_2),.dout(w_dff_B_FYGPnNpu9_2),.clk(gclk));
	jdff dff_B_U72RIqzP6_2(.din(w_dff_B_FYGPnNpu9_2),.dout(w_dff_B_U72RIqzP6_2),.clk(gclk));
	jdff dff_B_Ye12bHrZ4_2(.din(w_dff_B_U72RIqzP6_2),.dout(w_dff_B_Ye12bHrZ4_2),.clk(gclk));
	jdff dff_B_tdQHx3IX6_2(.din(w_dff_B_Ye12bHrZ4_2),.dout(w_dff_B_tdQHx3IX6_2),.clk(gclk));
	jdff dff_B_b5n9cWZD5_2(.din(w_dff_B_tdQHx3IX6_2),.dout(w_dff_B_b5n9cWZD5_2),.clk(gclk));
	jdff dff_B_W8rA4ORs4_2(.din(w_dff_B_b5n9cWZD5_2),.dout(w_dff_B_W8rA4ORs4_2),.clk(gclk));
	jdff dff_B_RTBweTss8_2(.din(w_dff_B_W8rA4ORs4_2),.dout(w_dff_B_RTBweTss8_2),.clk(gclk));
	jdff dff_B_pBfnd1Mh9_2(.din(w_dff_B_RTBweTss8_2),.dout(w_dff_B_pBfnd1Mh9_2),.clk(gclk));
	jdff dff_B_rsubGjLf5_2(.din(w_dff_B_pBfnd1Mh9_2),.dout(w_dff_B_rsubGjLf5_2),.clk(gclk));
	jdff dff_B_twt5G07e5_2(.din(w_dff_B_rsubGjLf5_2),.dout(w_dff_B_twt5G07e5_2),.clk(gclk));
	jdff dff_B_AuVUz9C37_2(.din(w_dff_B_twt5G07e5_2),.dout(w_dff_B_AuVUz9C37_2),.clk(gclk));
	jdff dff_B_QgPmRcTe4_2(.din(w_dff_B_AuVUz9C37_2),.dout(w_dff_B_QgPmRcTe4_2),.clk(gclk));
	jdff dff_B_hADkqKJi8_2(.din(w_dff_B_QgPmRcTe4_2),.dout(w_dff_B_hADkqKJi8_2),.clk(gclk));
	jdff dff_B_Iv9JaAqt2_2(.din(w_dff_B_hADkqKJi8_2),.dout(w_dff_B_Iv9JaAqt2_2),.clk(gclk));
	jdff dff_B_jJazrxyt0_2(.din(w_dff_B_Iv9JaAqt2_2),.dout(w_dff_B_jJazrxyt0_2),.clk(gclk));
	jdff dff_B_P8AMhOAB1_2(.din(w_dff_B_jJazrxyt0_2),.dout(w_dff_B_P8AMhOAB1_2),.clk(gclk));
	jdff dff_B_nv02lWB33_2(.din(w_dff_B_P8AMhOAB1_2),.dout(w_dff_B_nv02lWB33_2),.clk(gclk));
	jdff dff_B_9mDozcmb5_2(.din(w_dff_B_nv02lWB33_2),.dout(w_dff_B_9mDozcmb5_2),.clk(gclk));
	jdff dff_B_jrhByb670_2(.din(w_dff_B_9mDozcmb5_2),.dout(w_dff_B_jrhByb670_2),.clk(gclk));
	jdff dff_B_4XLpSYJq5_2(.din(w_dff_B_jrhByb670_2),.dout(w_dff_B_4XLpSYJq5_2),.clk(gclk));
	jdff dff_B_aK6adQKb1_2(.din(w_dff_B_4XLpSYJq5_2),.dout(w_dff_B_aK6adQKb1_2),.clk(gclk));
	jdff dff_B_xaspD9l37_2(.din(w_dff_B_aK6adQKb1_2),.dout(w_dff_B_xaspD9l37_2),.clk(gclk));
	jdff dff_B_xK8wlVqX9_2(.din(w_dff_B_xaspD9l37_2),.dout(w_dff_B_xK8wlVqX9_2),.clk(gclk));
	jdff dff_B_IwqRa1pJ4_2(.din(w_dff_B_xK8wlVqX9_2),.dout(w_dff_B_IwqRa1pJ4_2),.clk(gclk));
	jdff dff_B_RHRcBqPg9_2(.din(w_dff_B_IwqRa1pJ4_2),.dout(w_dff_B_RHRcBqPg9_2),.clk(gclk));
	jdff dff_B_eRk4JWa99_2(.din(w_dff_B_RHRcBqPg9_2),.dout(w_dff_B_eRk4JWa99_2),.clk(gclk));
	jdff dff_B_5fK0CbFV1_2(.din(w_dff_B_eRk4JWa99_2),.dout(w_dff_B_5fK0CbFV1_2),.clk(gclk));
	jdff dff_B_Jl7bPsJO7_2(.din(w_dff_B_5fK0CbFV1_2),.dout(w_dff_B_Jl7bPsJO7_2),.clk(gclk));
	jdff dff_B_ZgtcSHaY9_2(.din(n1651),.dout(w_dff_B_ZgtcSHaY9_2),.clk(gclk));
	jdff dff_B_8AToENM26_1(.din(n1649),.dout(w_dff_B_8AToENM26_1),.clk(gclk));
	jdff dff_B_hYO2MQ7m6_2(.din(n1591),.dout(w_dff_B_hYO2MQ7m6_2),.clk(gclk));
	jdff dff_B_wEb6SDTz8_2(.din(w_dff_B_hYO2MQ7m6_2),.dout(w_dff_B_wEb6SDTz8_2),.clk(gclk));
	jdff dff_B_uJfVdAMq6_2(.din(w_dff_B_wEb6SDTz8_2),.dout(w_dff_B_uJfVdAMq6_2),.clk(gclk));
	jdff dff_B_z0AXP81o5_2(.din(w_dff_B_uJfVdAMq6_2),.dout(w_dff_B_z0AXP81o5_2),.clk(gclk));
	jdff dff_B_54pIyioL7_2(.din(w_dff_B_z0AXP81o5_2),.dout(w_dff_B_54pIyioL7_2),.clk(gclk));
	jdff dff_B_TkA8Iy4I9_2(.din(w_dff_B_54pIyioL7_2),.dout(w_dff_B_TkA8Iy4I9_2),.clk(gclk));
	jdff dff_B_16xdJ4M99_2(.din(w_dff_B_TkA8Iy4I9_2),.dout(w_dff_B_16xdJ4M99_2),.clk(gclk));
	jdff dff_B_2lrtg4CN8_2(.din(w_dff_B_16xdJ4M99_2),.dout(w_dff_B_2lrtg4CN8_2),.clk(gclk));
	jdff dff_B_cBxlOMyj7_2(.din(w_dff_B_2lrtg4CN8_2),.dout(w_dff_B_cBxlOMyj7_2),.clk(gclk));
	jdff dff_B_1cZNdXJN4_2(.din(w_dff_B_cBxlOMyj7_2),.dout(w_dff_B_1cZNdXJN4_2),.clk(gclk));
	jdff dff_B_HMm2gWIm2_2(.din(w_dff_B_1cZNdXJN4_2),.dout(w_dff_B_HMm2gWIm2_2),.clk(gclk));
	jdff dff_B_uROQAyYm0_2(.din(w_dff_B_HMm2gWIm2_2),.dout(w_dff_B_uROQAyYm0_2),.clk(gclk));
	jdff dff_B_ZGHPxLHT4_2(.din(w_dff_B_uROQAyYm0_2),.dout(w_dff_B_ZGHPxLHT4_2),.clk(gclk));
	jdff dff_B_BoxmYpWt9_2(.din(w_dff_B_ZGHPxLHT4_2),.dout(w_dff_B_BoxmYpWt9_2),.clk(gclk));
	jdff dff_B_s147yXgz8_2(.din(w_dff_B_BoxmYpWt9_2),.dout(w_dff_B_s147yXgz8_2),.clk(gclk));
	jdff dff_B_ig0Z2EHv7_2(.din(w_dff_B_s147yXgz8_2),.dout(w_dff_B_ig0Z2EHv7_2),.clk(gclk));
	jdff dff_B_isverOzf2_2(.din(w_dff_B_ig0Z2EHv7_2),.dout(w_dff_B_isverOzf2_2),.clk(gclk));
	jdff dff_B_h0ACUAL07_2(.din(w_dff_B_isverOzf2_2),.dout(w_dff_B_h0ACUAL07_2),.clk(gclk));
	jdff dff_B_jxWozL602_2(.din(w_dff_B_h0ACUAL07_2),.dout(w_dff_B_jxWozL602_2),.clk(gclk));
	jdff dff_B_s3eZUIUA3_2(.din(w_dff_B_jxWozL602_2),.dout(w_dff_B_s3eZUIUA3_2),.clk(gclk));
	jdff dff_B_otmrRu990_2(.din(w_dff_B_s3eZUIUA3_2),.dout(w_dff_B_otmrRu990_2),.clk(gclk));
	jdff dff_B_hgAjOtlX1_2(.din(w_dff_B_otmrRu990_2),.dout(w_dff_B_hgAjOtlX1_2),.clk(gclk));
	jdff dff_B_MtgfJ5PA9_2(.din(w_dff_B_hgAjOtlX1_2),.dout(w_dff_B_MtgfJ5PA9_2),.clk(gclk));
	jdff dff_B_0jd2Rb4T7_2(.din(w_dff_B_MtgfJ5PA9_2),.dout(w_dff_B_0jd2Rb4T7_2),.clk(gclk));
	jdff dff_B_9EQoKnIl6_2(.din(w_dff_B_0jd2Rb4T7_2),.dout(w_dff_B_9EQoKnIl6_2),.clk(gclk));
	jdff dff_B_WKfFzGgQ2_2(.din(w_dff_B_9EQoKnIl6_2),.dout(w_dff_B_WKfFzGgQ2_2),.clk(gclk));
	jdff dff_B_ztfniFbs0_2(.din(w_dff_B_WKfFzGgQ2_2),.dout(w_dff_B_ztfniFbs0_2),.clk(gclk));
	jdff dff_B_Uqw05TLl4_1(.din(n1597),.dout(w_dff_B_Uqw05TLl4_1),.clk(gclk));
	jdff dff_B_KARzh2LJ3_1(.din(w_dff_B_Uqw05TLl4_1),.dout(w_dff_B_KARzh2LJ3_1),.clk(gclk));
	jdff dff_B_SwQ8kzZG9_2(.din(n1596),.dout(w_dff_B_SwQ8kzZG9_2),.clk(gclk));
	jdff dff_B_qTWxOjmh9_2(.din(w_dff_B_SwQ8kzZG9_2),.dout(w_dff_B_qTWxOjmh9_2),.clk(gclk));
	jdff dff_B_FArDLjPv7_2(.din(w_dff_B_qTWxOjmh9_2),.dout(w_dff_B_FArDLjPv7_2),.clk(gclk));
	jdff dff_B_63ryLsMq7_2(.din(w_dff_B_FArDLjPv7_2),.dout(w_dff_B_63ryLsMq7_2),.clk(gclk));
	jdff dff_B_U8UxU3bN4_2(.din(w_dff_B_63ryLsMq7_2),.dout(w_dff_B_U8UxU3bN4_2),.clk(gclk));
	jdff dff_B_pRJYqoAl5_2(.din(w_dff_B_U8UxU3bN4_2),.dout(w_dff_B_pRJYqoAl5_2),.clk(gclk));
	jdff dff_B_pKRAuQqg9_2(.din(w_dff_B_pRJYqoAl5_2),.dout(w_dff_B_pKRAuQqg9_2),.clk(gclk));
	jdff dff_B_n0GmbCEk2_2(.din(w_dff_B_pKRAuQqg9_2),.dout(w_dff_B_n0GmbCEk2_2),.clk(gclk));
	jdff dff_B_UmyYzFAS5_2(.din(w_dff_B_n0GmbCEk2_2),.dout(w_dff_B_UmyYzFAS5_2),.clk(gclk));
	jdff dff_B_0VikFm1P0_2(.din(w_dff_B_UmyYzFAS5_2),.dout(w_dff_B_0VikFm1P0_2),.clk(gclk));
	jdff dff_B_U1z4qvW22_2(.din(w_dff_B_0VikFm1P0_2),.dout(w_dff_B_U1z4qvW22_2),.clk(gclk));
	jdff dff_B_TdHEhK7J7_2(.din(w_dff_B_U1z4qvW22_2),.dout(w_dff_B_TdHEhK7J7_2),.clk(gclk));
	jdff dff_B_Tpj7kjtB6_2(.din(w_dff_B_TdHEhK7J7_2),.dout(w_dff_B_Tpj7kjtB6_2),.clk(gclk));
	jdff dff_B_jNTNi3Tg3_2(.din(w_dff_B_Tpj7kjtB6_2),.dout(w_dff_B_jNTNi3Tg3_2),.clk(gclk));
	jdff dff_B_FBmyCJL18_2(.din(w_dff_B_jNTNi3Tg3_2),.dout(w_dff_B_FBmyCJL18_2),.clk(gclk));
	jdff dff_B_4SpswkaO6_2(.din(w_dff_B_FBmyCJL18_2),.dout(w_dff_B_4SpswkaO6_2),.clk(gclk));
	jdff dff_B_cJqfEbKN8_2(.din(w_dff_B_4SpswkaO6_2),.dout(w_dff_B_cJqfEbKN8_2),.clk(gclk));
	jdff dff_B_yjSWSKcy7_2(.din(w_dff_B_cJqfEbKN8_2),.dout(w_dff_B_yjSWSKcy7_2),.clk(gclk));
	jdff dff_B_H6IypFwe6_2(.din(w_dff_B_yjSWSKcy7_2),.dout(w_dff_B_H6IypFwe6_2),.clk(gclk));
	jdff dff_B_6oq6cpMR6_2(.din(w_dff_B_H6IypFwe6_2),.dout(w_dff_B_6oq6cpMR6_2),.clk(gclk));
	jdff dff_B_H8R0rlwr1_2(.din(w_dff_B_6oq6cpMR6_2),.dout(w_dff_B_H8R0rlwr1_2),.clk(gclk));
	jdff dff_B_kh1UKGBO4_2(.din(w_dff_B_H8R0rlwr1_2),.dout(w_dff_B_kh1UKGBO4_2),.clk(gclk));
	jdff dff_B_6KOgTE5Z4_2(.din(w_dff_B_kh1UKGBO4_2),.dout(w_dff_B_6KOgTE5Z4_2),.clk(gclk));
	jdff dff_B_dHTgEsif0_2(.din(w_dff_B_6KOgTE5Z4_2),.dout(w_dff_B_dHTgEsif0_2),.clk(gclk));
	jdff dff_B_PY28HlVW5_2(.din(n1595),.dout(w_dff_B_PY28HlVW5_2),.clk(gclk));
	jdff dff_B_Ntj80Knl4_2(.din(w_dff_B_PY28HlVW5_2),.dout(w_dff_B_Ntj80Knl4_2),.clk(gclk));
	jdff dff_B_QevNkeav6_2(.din(w_dff_B_Ntj80Knl4_2),.dout(w_dff_B_QevNkeav6_2),.clk(gclk));
	jdff dff_B_kCvtrqo36_2(.din(w_dff_B_QevNkeav6_2),.dout(w_dff_B_kCvtrqo36_2),.clk(gclk));
	jdff dff_B_wsbb7vzP7_2(.din(w_dff_B_kCvtrqo36_2),.dout(w_dff_B_wsbb7vzP7_2),.clk(gclk));
	jdff dff_B_NwcEb03n2_2(.din(w_dff_B_wsbb7vzP7_2),.dout(w_dff_B_NwcEb03n2_2),.clk(gclk));
	jdff dff_B_Kh6nPWOF1_2(.din(w_dff_B_NwcEb03n2_2),.dout(w_dff_B_Kh6nPWOF1_2),.clk(gclk));
	jdff dff_B_H1L0yD0s7_2(.din(w_dff_B_Kh6nPWOF1_2),.dout(w_dff_B_H1L0yD0s7_2),.clk(gclk));
	jdff dff_B_FUOZRwUc9_2(.din(w_dff_B_H1L0yD0s7_2),.dout(w_dff_B_FUOZRwUc9_2),.clk(gclk));
	jdff dff_B_EG79hSRm9_2(.din(w_dff_B_FUOZRwUc9_2),.dout(w_dff_B_EG79hSRm9_2),.clk(gclk));
	jdff dff_B_QwBL5dEG8_2(.din(w_dff_B_EG79hSRm9_2),.dout(w_dff_B_QwBL5dEG8_2),.clk(gclk));
	jdff dff_B_r2R7smak5_2(.din(w_dff_B_QwBL5dEG8_2),.dout(w_dff_B_r2R7smak5_2),.clk(gclk));
	jdff dff_B_6pTO68Sw0_2(.din(w_dff_B_r2R7smak5_2),.dout(w_dff_B_6pTO68Sw0_2),.clk(gclk));
	jdff dff_B_T2bqYwub4_2(.din(w_dff_B_6pTO68Sw0_2),.dout(w_dff_B_T2bqYwub4_2),.clk(gclk));
	jdff dff_B_556b7PXp0_2(.din(w_dff_B_T2bqYwub4_2),.dout(w_dff_B_556b7PXp0_2),.clk(gclk));
	jdff dff_B_tYzZqhzB6_2(.din(w_dff_B_556b7PXp0_2),.dout(w_dff_B_tYzZqhzB6_2),.clk(gclk));
	jdff dff_B_BvMkBAov2_2(.din(w_dff_B_tYzZqhzB6_2),.dout(w_dff_B_BvMkBAov2_2),.clk(gclk));
	jdff dff_B_OHnCXbBO7_2(.din(w_dff_B_BvMkBAov2_2),.dout(w_dff_B_OHnCXbBO7_2),.clk(gclk));
	jdff dff_B_QJAbgZND2_2(.din(w_dff_B_OHnCXbBO7_2),.dout(w_dff_B_QJAbgZND2_2),.clk(gclk));
	jdff dff_B_6fdHWPhQ1_2(.din(w_dff_B_QJAbgZND2_2),.dout(w_dff_B_6fdHWPhQ1_2),.clk(gclk));
	jdff dff_B_b6wd8B4S1_2(.din(w_dff_B_6fdHWPhQ1_2),.dout(w_dff_B_b6wd8B4S1_2),.clk(gclk));
	jdff dff_B_bmSptCoe5_2(.din(w_dff_B_b6wd8B4S1_2),.dout(w_dff_B_bmSptCoe5_2),.clk(gclk));
	jdff dff_B_RmDgsv8m9_2(.din(w_dff_B_bmSptCoe5_2),.dout(w_dff_B_RmDgsv8m9_2),.clk(gclk));
	jdff dff_B_HXg69b2L5_2(.din(w_dff_B_RmDgsv8m9_2),.dout(w_dff_B_HXg69b2L5_2),.clk(gclk));
	jdff dff_B_XzRk4iNO4_2(.din(w_dff_B_HXg69b2L5_2),.dout(w_dff_B_XzRk4iNO4_2),.clk(gclk));
	jdff dff_B_6vXFpnbZ4_2(.din(w_dff_B_XzRk4iNO4_2),.dout(w_dff_B_6vXFpnbZ4_2),.clk(gclk));
	jdff dff_B_PXxDP2ZQ2_2(.din(n1594),.dout(w_dff_B_PXxDP2ZQ2_2),.clk(gclk));
	jdff dff_B_s0iMEh9j6_1(.din(n1592),.dout(w_dff_B_s0iMEh9j6_1),.clk(gclk));
	jdff dff_B_mWOa81Rk5_2(.din(n1527),.dout(w_dff_B_mWOa81Rk5_2),.clk(gclk));
	jdff dff_B_ISny6vEW4_2(.din(w_dff_B_mWOa81Rk5_2),.dout(w_dff_B_ISny6vEW4_2),.clk(gclk));
	jdff dff_B_BvuQ1cza0_2(.din(w_dff_B_ISny6vEW4_2),.dout(w_dff_B_BvuQ1cza0_2),.clk(gclk));
	jdff dff_B_weaMn54Z0_2(.din(w_dff_B_BvuQ1cza0_2),.dout(w_dff_B_weaMn54Z0_2),.clk(gclk));
	jdff dff_B_rQgBqpsl1_2(.din(w_dff_B_weaMn54Z0_2),.dout(w_dff_B_rQgBqpsl1_2),.clk(gclk));
	jdff dff_B_T6hGHSEv5_2(.din(w_dff_B_rQgBqpsl1_2),.dout(w_dff_B_T6hGHSEv5_2),.clk(gclk));
	jdff dff_B_w5wkDeUs3_2(.din(w_dff_B_T6hGHSEv5_2),.dout(w_dff_B_w5wkDeUs3_2),.clk(gclk));
	jdff dff_B_flvje6QQ0_2(.din(w_dff_B_w5wkDeUs3_2),.dout(w_dff_B_flvje6QQ0_2),.clk(gclk));
	jdff dff_B_F6k9YprD2_2(.din(w_dff_B_flvje6QQ0_2),.dout(w_dff_B_F6k9YprD2_2),.clk(gclk));
	jdff dff_B_T3DxtkCa9_2(.din(w_dff_B_F6k9YprD2_2),.dout(w_dff_B_T3DxtkCa9_2),.clk(gclk));
	jdff dff_B_yjUduDbD6_2(.din(w_dff_B_T3DxtkCa9_2),.dout(w_dff_B_yjUduDbD6_2),.clk(gclk));
	jdff dff_B_Dk5lbwa53_2(.din(w_dff_B_yjUduDbD6_2),.dout(w_dff_B_Dk5lbwa53_2),.clk(gclk));
	jdff dff_B_cUDNQNix4_2(.din(w_dff_B_Dk5lbwa53_2),.dout(w_dff_B_cUDNQNix4_2),.clk(gclk));
	jdff dff_B_CaOXVu8i4_2(.din(w_dff_B_cUDNQNix4_2),.dout(w_dff_B_CaOXVu8i4_2),.clk(gclk));
	jdff dff_B_Ssn2jGft0_2(.din(w_dff_B_CaOXVu8i4_2),.dout(w_dff_B_Ssn2jGft0_2),.clk(gclk));
	jdff dff_B_kppgszoA2_2(.din(w_dff_B_Ssn2jGft0_2),.dout(w_dff_B_kppgszoA2_2),.clk(gclk));
	jdff dff_B_djuiL1bi5_2(.din(w_dff_B_kppgszoA2_2),.dout(w_dff_B_djuiL1bi5_2),.clk(gclk));
	jdff dff_B_RGy0bzld9_2(.din(w_dff_B_djuiL1bi5_2),.dout(w_dff_B_RGy0bzld9_2),.clk(gclk));
	jdff dff_B_WbMsBM4E3_2(.din(w_dff_B_RGy0bzld9_2),.dout(w_dff_B_WbMsBM4E3_2),.clk(gclk));
	jdff dff_B_vlCMFHgH6_2(.din(w_dff_B_WbMsBM4E3_2),.dout(w_dff_B_vlCMFHgH6_2),.clk(gclk));
	jdff dff_B_NjwkrKHV4_2(.din(w_dff_B_vlCMFHgH6_2),.dout(w_dff_B_NjwkrKHV4_2),.clk(gclk));
	jdff dff_B_Ayj4Rhso9_2(.din(w_dff_B_NjwkrKHV4_2),.dout(w_dff_B_Ayj4Rhso9_2),.clk(gclk));
	jdff dff_B_v7oCyk8L3_2(.din(w_dff_B_Ayj4Rhso9_2),.dout(w_dff_B_v7oCyk8L3_2),.clk(gclk));
	jdff dff_B_j9F6fm7H5_2(.din(w_dff_B_v7oCyk8L3_2),.dout(w_dff_B_j9F6fm7H5_2),.clk(gclk));
	jdff dff_B_rhDUsWj34_1(.din(n1533),.dout(w_dff_B_rhDUsWj34_1),.clk(gclk));
	jdff dff_B_CsrK5ZqW4_1(.din(w_dff_B_rhDUsWj34_1),.dout(w_dff_B_CsrK5ZqW4_1),.clk(gclk));
	jdff dff_B_hXMUlXj97_2(.din(n1532),.dout(w_dff_B_hXMUlXj97_2),.clk(gclk));
	jdff dff_B_vn4HAjen4_2(.din(w_dff_B_hXMUlXj97_2),.dout(w_dff_B_vn4HAjen4_2),.clk(gclk));
	jdff dff_B_lLZPluQI1_2(.din(w_dff_B_vn4HAjen4_2),.dout(w_dff_B_lLZPluQI1_2),.clk(gclk));
	jdff dff_B_iFJeX5hP4_2(.din(w_dff_B_lLZPluQI1_2),.dout(w_dff_B_iFJeX5hP4_2),.clk(gclk));
	jdff dff_B_2NtFqqix5_2(.din(w_dff_B_iFJeX5hP4_2),.dout(w_dff_B_2NtFqqix5_2),.clk(gclk));
	jdff dff_B_wc4Y4toX6_2(.din(w_dff_B_2NtFqqix5_2),.dout(w_dff_B_wc4Y4toX6_2),.clk(gclk));
	jdff dff_B_UOQsEt7c9_2(.din(w_dff_B_wc4Y4toX6_2),.dout(w_dff_B_UOQsEt7c9_2),.clk(gclk));
	jdff dff_B_Jee3Zt722_2(.din(w_dff_B_UOQsEt7c9_2),.dout(w_dff_B_Jee3Zt722_2),.clk(gclk));
	jdff dff_B_srBTgxHS2_2(.din(w_dff_B_Jee3Zt722_2),.dout(w_dff_B_srBTgxHS2_2),.clk(gclk));
	jdff dff_B_4VnwhoLy7_2(.din(w_dff_B_srBTgxHS2_2),.dout(w_dff_B_4VnwhoLy7_2),.clk(gclk));
	jdff dff_B_BPb5ynIG3_2(.din(w_dff_B_4VnwhoLy7_2),.dout(w_dff_B_BPb5ynIG3_2),.clk(gclk));
	jdff dff_B_0KARpA4n3_2(.din(w_dff_B_BPb5ynIG3_2),.dout(w_dff_B_0KARpA4n3_2),.clk(gclk));
	jdff dff_B_FT4J4oWT7_2(.din(w_dff_B_0KARpA4n3_2),.dout(w_dff_B_FT4J4oWT7_2),.clk(gclk));
	jdff dff_B_BY6LPpUv3_2(.din(w_dff_B_FT4J4oWT7_2),.dout(w_dff_B_BY6LPpUv3_2),.clk(gclk));
	jdff dff_B_twxpVCLP9_2(.din(w_dff_B_BY6LPpUv3_2),.dout(w_dff_B_twxpVCLP9_2),.clk(gclk));
	jdff dff_B_xdLCfyIs9_2(.din(w_dff_B_twxpVCLP9_2),.dout(w_dff_B_xdLCfyIs9_2),.clk(gclk));
	jdff dff_B_m9TmWIG89_2(.din(w_dff_B_xdLCfyIs9_2),.dout(w_dff_B_m9TmWIG89_2),.clk(gclk));
	jdff dff_B_ZsXnbvxn7_2(.din(w_dff_B_m9TmWIG89_2),.dout(w_dff_B_ZsXnbvxn7_2),.clk(gclk));
	jdff dff_B_tmjAr3ij4_2(.din(w_dff_B_ZsXnbvxn7_2),.dout(w_dff_B_tmjAr3ij4_2),.clk(gclk));
	jdff dff_B_xMROSzql1_2(.din(w_dff_B_tmjAr3ij4_2),.dout(w_dff_B_xMROSzql1_2),.clk(gclk));
	jdff dff_B_0maDXt469_2(.din(w_dff_B_xMROSzql1_2),.dout(w_dff_B_0maDXt469_2),.clk(gclk));
	jdff dff_B_LAHOgGhx2_2(.din(n1531),.dout(w_dff_B_LAHOgGhx2_2),.clk(gclk));
	jdff dff_B_rSecc6as2_2(.din(w_dff_B_LAHOgGhx2_2),.dout(w_dff_B_rSecc6as2_2),.clk(gclk));
	jdff dff_B_HpFlco0h5_2(.din(w_dff_B_rSecc6as2_2),.dout(w_dff_B_HpFlco0h5_2),.clk(gclk));
	jdff dff_B_v9KDYvbD4_2(.din(w_dff_B_HpFlco0h5_2),.dout(w_dff_B_v9KDYvbD4_2),.clk(gclk));
	jdff dff_B_AEgcHMBt7_2(.din(w_dff_B_v9KDYvbD4_2),.dout(w_dff_B_AEgcHMBt7_2),.clk(gclk));
	jdff dff_B_oJyGlvUs4_2(.din(w_dff_B_AEgcHMBt7_2),.dout(w_dff_B_oJyGlvUs4_2),.clk(gclk));
	jdff dff_B_oYAFx4dZ2_2(.din(w_dff_B_oJyGlvUs4_2),.dout(w_dff_B_oYAFx4dZ2_2),.clk(gclk));
	jdff dff_B_pUjFk1WI7_2(.din(w_dff_B_oYAFx4dZ2_2),.dout(w_dff_B_pUjFk1WI7_2),.clk(gclk));
	jdff dff_B_8zzSTvs93_2(.din(w_dff_B_pUjFk1WI7_2),.dout(w_dff_B_8zzSTvs93_2),.clk(gclk));
	jdff dff_B_HZ1MYFKA4_2(.din(w_dff_B_8zzSTvs93_2),.dout(w_dff_B_HZ1MYFKA4_2),.clk(gclk));
	jdff dff_B_70V6dmNT8_2(.din(w_dff_B_HZ1MYFKA4_2),.dout(w_dff_B_70V6dmNT8_2),.clk(gclk));
	jdff dff_B_4YMXx4vV4_2(.din(w_dff_B_70V6dmNT8_2),.dout(w_dff_B_4YMXx4vV4_2),.clk(gclk));
	jdff dff_B_sKToEarR1_2(.din(w_dff_B_4YMXx4vV4_2),.dout(w_dff_B_sKToEarR1_2),.clk(gclk));
	jdff dff_B_tsfA4iAg5_2(.din(w_dff_B_sKToEarR1_2),.dout(w_dff_B_tsfA4iAg5_2),.clk(gclk));
	jdff dff_B_qX6Vr7g68_2(.din(w_dff_B_tsfA4iAg5_2),.dout(w_dff_B_qX6Vr7g68_2),.clk(gclk));
	jdff dff_B_2da2878j4_2(.din(w_dff_B_qX6Vr7g68_2),.dout(w_dff_B_2da2878j4_2),.clk(gclk));
	jdff dff_B_1nLpnGve6_2(.din(w_dff_B_2da2878j4_2),.dout(w_dff_B_1nLpnGve6_2),.clk(gclk));
	jdff dff_B_4t2jPIFm1_2(.din(w_dff_B_1nLpnGve6_2),.dout(w_dff_B_4t2jPIFm1_2),.clk(gclk));
	jdff dff_B_aWmcrJ1x8_2(.din(w_dff_B_4t2jPIFm1_2),.dout(w_dff_B_aWmcrJ1x8_2),.clk(gclk));
	jdff dff_B_zUJELoid4_2(.din(w_dff_B_aWmcrJ1x8_2),.dout(w_dff_B_zUJELoid4_2),.clk(gclk));
	jdff dff_B_nslbwkcb9_2(.din(w_dff_B_zUJELoid4_2),.dout(w_dff_B_nslbwkcb9_2),.clk(gclk));
	jdff dff_B_qiGqY5316_2(.din(w_dff_B_nslbwkcb9_2),.dout(w_dff_B_qiGqY5316_2),.clk(gclk));
	jdff dff_B_RaaEakny6_2(.din(w_dff_B_qiGqY5316_2),.dout(w_dff_B_RaaEakny6_2),.clk(gclk));
	jdff dff_B_CT3WHjNg5_2(.din(n1530),.dout(w_dff_B_CT3WHjNg5_2),.clk(gclk));
	jdff dff_B_0LPPkpTF8_1(.din(n1528),.dout(w_dff_B_0LPPkpTF8_1),.clk(gclk));
	jdff dff_B_ro4fgAqA8_2(.din(n1456),.dout(w_dff_B_ro4fgAqA8_2),.clk(gclk));
	jdff dff_B_HxMFnHtK6_2(.din(w_dff_B_ro4fgAqA8_2),.dout(w_dff_B_HxMFnHtK6_2),.clk(gclk));
	jdff dff_B_RU535DrL4_2(.din(w_dff_B_HxMFnHtK6_2),.dout(w_dff_B_RU535DrL4_2),.clk(gclk));
	jdff dff_B_VVHSkZ501_2(.din(w_dff_B_RU535DrL4_2),.dout(w_dff_B_VVHSkZ501_2),.clk(gclk));
	jdff dff_B_MjfSUJft1_2(.din(w_dff_B_VVHSkZ501_2),.dout(w_dff_B_MjfSUJft1_2),.clk(gclk));
	jdff dff_B_zuInLHpI9_2(.din(w_dff_B_MjfSUJft1_2),.dout(w_dff_B_zuInLHpI9_2),.clk(gclk));
	jdff dff_B_jVXcfI5U1_2(.din(w_dff_B_zuInLHpI9_2),.dout(w_dff_B_jVXcfI5U1_2),.clk(gclk));
	jdff dff_B_IJvuMKKD6_2(.din(w_dff_B_jVXcfI5U1_2),.dout(w_dff_B_IJvuMKKD6_2),.clk(gclk));
	jdff dff_B_KKRfMiwM5_2(.din(w_dff_B_IJvuMKKD6_2),.dout(w_dff_B_KKRfMiwM5_2),.clk(gclk));
	jdff dff_B_H35ZoJAT4_2(.din(w_dff_B_KKRfMiwM5_2),.dout(w_dff_B_H35ZoJAT4_2),.clk(gclk));
	jdff dff_B_ZHDQzUp84_2(.din(w_dff_B_H35ZoJAT4_2),.dout(w_dff_B_ZHDQzUp84_2),.clk(gclk));
	jdff dff_B_QrQq3D3c4_2(.din(w_dff_B_ZHDQzUp84_2),.dout(w_dff_B_QrQq3D3c4_2),.clk(gclk));
	jdff dff_B_6b2pPNmg5_2(.din(w_dff_B_QrQq3D3c4_2),.dout(w_dff_B_6b2pPNmg5_2),.clk(gclk));
	jdff dff_B_UfrgNYyG2_2(.din(w_dff_B_6b2pPNmg5_2),.dout(w_dff_B_UfrgNYyG2_2),.clk(gclk));
	jdff dff_B_9bSCueTo5_2(.din(w_dff_B_UfrgNYyG2_2),.dout(w_dff_B_9bSCueTo5_2),.clk(gclk));
	jdff dff_B_45HiwsA46_2(.din(w_dff_B_9bSCueTo5_2),.dout(w_dff_B_45HiwsA46_2),.clk(gclk));
	jdff dff_B_cbzno6ca3_2(.din(w_dff_B_45HiwsA46_2),.dout(w_dff_B_cbzno6ca3_2),.clk(gclk));
	jdff dff_B_ijZyGR887_2(.din(w_dff_B_cbzno6ca3_2),.dout(w_dff_B_ijZyGR887_2),.clk(gclk));
	jdff dff_B_KEqVdexm6_2(.din(w_dff_B_ijZyGR887_2),.dout(w_dff_B_KEqVdexm6_2),.clk(gclk));
	jdff dff_B_ppiFikWv1_2(.din(w_dff_B_KEqVdexm6_2),.dout(w_dff_B_ppiFikWv1_2),.clk(gclk));
	jdff dff_B_kU5hk7Wz5_2(.din(w_dff_B_ppiFikWv1_2),.dout(w_dff_B_kU5hk7Wz5_2),.clk(gclk));
	jdff dff_B_4CfiHYsM2_1(.din(n1462),.dout(w_dff_B_4CfiHYsM2_1),.clk(gclk));
	jdff dff_B_zYK4DSNq2_1(.din(w_dff_B_4CfiHYsM2_1),.dout(w_dff_B_zYK4DSNq2_1),.clk(gclk));
	jdff dff_B_NygoV7GR9_2(.din(n1461),.dout(w_dff_B_NygoV7GR9_2),.clk(gclk));
	jdff dff_B_PpOnQ7r68_2(.din(w_dff_B_NygoV7GR9_2),.dout(w_dff_B_PpOnQ7r68_2),.clk(gclk));
	jdff dff_B_6OGf1WYy6_2(.din(w_dff_B_PpOnQ7r68_2),.dout(w_dff_B_6OGf1WYy6_2),.clk(gclk));
	jdff dff_B_seqL7K5u9_2(.din(w_dff_B_6OGf1WYy6_2),.dout(w_dff_B_seqL7K5u9_2),.clk(gclk));
	jdff dff_B_vWRcOAUg8_2(.din(w_dff_B_seqL7K5u9_2),.dout(w_dff_B_vWRcOAUg8_2),.clk(gclk));
	jdff dff_B_AZUq8oyp9_2(.din(w_dff_B_vWRcOAUg8_2),.dout(w_dff_B_AZUq8oyp9_2),.clk(gclk));
	jdff dff_B_YZTjUDOJ7_2(.din(w_dff_B_AZUq8oyp9_2),.dout(w_dff_B_YZTjUDOJ7_2),.clk(gclk));
	jdff dff_B_p9zWEvwv3_2(.din(w_dff_B_YZTjUDOJ7_2),.dout(w_dff_B_p9zWEvwv3_2),.clk(gclk));
	jdff dff_B_6ZL7mFoF1_2(.din(w_dff_B_p9zWEvwv3_2),.dout(w_dff_B_6ZL7mFoF1_2),.clk(gclk));
	jdff dff_B_fwnuFRtw0_2(.din(w_dff_B_6ZL7mFoF1_2),.dout(w_dff_B_fwnuFRtw0_2),.clk(gclk));
	jdff dff_B_vLF1sW0w2_2(.din(w_dff_B_fwnuFRtw0_2),.dout(w_dff_B_vLF1sW0w2_2),.clk(gclk));
	jdff dff_B_B6bilmLw3_2(.din(w_dff_B_vLF1sW0w2_2),.dout(w_dff_B_B6bilmLw3_2),.clk(gclk));
	jdff dff_B_o85svmNf2_2(.din(w_dff_B_B6bilmLw3_2),.dout(w_dff_B_o85svmNf2_2),.clk(gclk));
	jdff dff_B_H3ektXat2_2(.din(w_dff_B_o85svmNf2_2),.dout(w_dff_B_H3ektXat2_2),.clk(gclk));
	jdff dff_B_YJSIwh8n5_2(.din(w_dff_B_H3ektXat2_2),.dout(w_dff_B_YJSIwh8n5_2),.clk(gclk));
	jdff dff_B_msx7xnt23_2(.din(w_dff_B_YJSIwh8n5_2),.dout(w_dff_B_msx7xnt23_2),.clk(gclk));
	jdff dff_B_JBteyBSG0_2(.din(w_dff_B_msx7xnt23_2),.dout(w_dff_B_JBteyBSG0_2),.clk(gclk));
	jdff dff_B_NAN3wn5C2_2(.din(w_dff_B_JBteyBSG0_2),.dout(w_dff_B_NAN3wn5C2_2),.clk(gclk));
	jdff dff_B_9b31hflg2_2(.din(n1460),.dout(w_dff_B_9b31hflg2_2),.clk(gclk));
	jdff dff_B_bn4XXQ5L1_2(.din(w_dff_B_9b31hflg2_2),.dout(w_dff_B_bn4XXQ5L1_2),.clk(gclk));
	jdff dff_B_uvPZUm570_2(.din(w_dff_B_bn4XXQ5L1_2),.dout(w_dff_B_uvPZUm570_2),.clk(gclk));
	jdff dff_B_RksPpFYX7_2(.din(w_dff_B_uvPZUm570_2),.dout(w_dff_B_RksPpFYX7_2),.clk(gclk));
	jdff dff_B_JxM20JC14_2(.din(w_dff_B_RksPpFYX7_2),.dout(w_dff_B_JxM20JC14_2),.clk(gclk));
	jdff dff_B_M9ak3Kws1_2(.din(w_dff_B_JxM20JC14_2),.dout(w_dff_B_M9ak3Kws1_2),.clk(gclk));
	jdff dff_B_ZsqlUFPP8_2(.din(w_dff_B_M9ak3Kws1_2),.dout(w_dff_B_ZsqlUFPP8_2),.clk(gclk));
	jdff dff_B_MK1w0YYY3_2(.din(w_dff_B_ZsqlUFPP8_2),.dout(w_dff_B_MK1w0YYY3_2),.clk(gclk));
	jdff dff_B_gioAlult0_2(.din(w_dff_B_MK1w0YYY3_2),.dout(w_dff_B_gioAlult0_2),.clk(gclk));
	jdff dff_B_Gx76qa393_2(.din(w_dff_B_gioAlult0_2),.dout(w_dff_B_Gx76qa393_2),.clk(gclk));
	jdff dff_B_kazSnlUS4_2(.din(w_dff_B_Gx76qa393_2),.dout(w_dff_B_kazSnlUS4_2),.clk(gclk));
	jdff dff_B_pMtSoTl52_2(.din(w_dff_B_kazSnlUS4_2),.dout(w_dff_B_pMtSoTl52_2),.clk(gclk));
	jdff dff_B_0t1rKXzn2_2(.din(w_dff_B_pMtSoTl52_2),.dout(w_dff_B_0t1rKXzn2_2),.clk(gclk));
	jdff dff_B_yEeBVL2n2_2(.din(w_dff_B_0t1rKXzn2_2),.dout(w_dff_B_yEeBVL2n2_2),.clk(gclk));
	jdff dff_B_dl3Fhrn45_2(.din(w_dff_B_yEeBVL2n2_2),.dout(w_dff_B_dl3Fhrn45_2),.clk(gclk));
	jdff dff_B_01Mgn8cX3_2(.din(w_dff_B_dl3Fhrn45_2),.dout(w_dff_B_01Mgn8cX3_2),.clk(gclk));
	jdff dff_B_LVChLgIA8_2(.din(w_dff_B_01Mgn8cX3_2),.dout(w_dff_B_LVChLgIA8_2),.clk(gclk));
	jdff dff_B_ePEybjNl3_2(.din(w_dff_B_LVChLgIA8_2),.dout(w_dff_B_ePEybjNl3_2),.clk(gclk));
	jdff dff_B_SxlNqlx32_2(.din(w_dff_B_ePEybjNl3_2),.dout(w_dff_B_SxlNqlx32_2),.clk(gclk));
	jdff dff_B_mDRr7Giz8_2(.din(w_dff_B_SxlNqlx32_2),.dout(w_dff_B_mDRr7Giz8_2),.clk(gclk));
	jdff dff_B_t2KKPViJ5_2(.din(n1459),.dout(w_dff_B_t2KKPViJ5_2),.clk(gclk));
	jdff dff_B_85e2vVXL1_1(.din(n1457),.dout(w_dff_B_85e2vVXL1_1),.clk(gclk));
	jdff dff_B_0fauM9z03_2(.din(n1378),.dout(w_dff_B_0fauM9z03_2),.clk(gclk));
	jdff dff_B_6jgaNYdq6_2(.din(w_dff_B_0fauM9z03_2),.dout(w_dff_B_6jgaNYdq6_2),.clk(gclk));
	jdff dff_B_iimuTfWp8_2(.din(w_dff_B_6jgaNYdq6_2),.dout(w_dff_B_iimuTfWp8_2),.clk(gclk));
	jdff dff_B_0hgtJpuu2_2(.din(w_dff_B_iimuTfWp8_2),.dout(w_dff_B_0hgtJpuu2_2),.clk(gclk));
	jdff dff_B_aqNhh1yW0_2(.din(w_dff_B_0hgtJpuu2_2),.dout(w_dff_B_aqNhh1yW0_2),.clk(gclk));
	jdff dff_B_JHAjo6kM2_2(.din(w_dff_B_aqNhh1yW0_2),.dout(w_dff_B_JHAjo6kM2_2),.clk(gclk));
	jdff dff_B_OZWJKUHE3_2(.din(w_dff_B_JHAjo6kM2_2),.dout(w_dff_B_OZWJKUHE3_2),.clk(gclk));
	jdff dff_B_Do8llFkC3_2(.din(w_dff_B_OZWJKUHE3_2),.dout(w_dff_B_Do8llFkC3_2),.clk(gclk));
	jdff dff_B_ggfJMlwP0_2(.din(w_dff_B_Do8llFkC3_2),.dout(w_dff_B_ggfJMlwP0_2),.clk(gclk));
	jdff dff_B_ggkfeHJt8_2(.din(w_dff_B_ggfJMlwP0_2),.dout(w_dff_B_ggkfeHJt8_2),.clk(gclk));
	jdff dff_B_E2Wox0Cw8_2(.din(w_dff_B_ggkfeHJt8_2),.dout(w_dff_B_E2Wox0Cw8_2),.clk(gclk));
	jdff dff_B_FpCNkiiD7_2(.din(w_dff_B_E2Wox0Cw8_2),.dout(w_dff_B_FpCNkiiD7_2),.clk(gclk));
	jdff dff_B_1GCLjYcJ5_2(.din(w_dff_B_FpCNkiiD7_2),.dout(w_dff_B_1GCLjYcJ5_2),.clk(gclk));
	jdff dff_B_sSXmnpaj4_2(.din(w_dff_B_1GCLjYcJ5_2),.dout(w_dff_B_sSXmnpaj4_2),.clk(gclk));
	jdff dff_B_xWS4CZJz3_2(.din(w_dff_B_sSXmnpaj4_2),.dout(w_dff_B_xWS4CZJz3_2),.clk(gclk));
	jdff dff_B_kmkDCwf04_2(.din(w_dff_B_xWS4CZJz3_2),.dout(w_dff_B_kmkDCwf04_2),.clk(gclk));
	jdff dff_B_3HXppIed7_2(.din(w_dff_B_kmkDCwf04_2),.dout(w_dff_B_3HXppIed7_2),.clk(gclk));
	jdff dff_B_L60jpsp08_2(.din(w_dff_B_3HXppIed7_2),.dout(w_dff_B_L60jpsp08_2),.clk(gclk));
	jdff dff_B_vNIMQ7pO9_1(.din(n1384),.dout(w_dff_B_vNIMQ7pO9_1),.clk(gclk));
	jdff dff_B_Oa0pA2St3_1(.din(w_dff_B_vNIMQ7pO9_1),.dout(w_dff_B_Oa0pA2St3_1),.clk(gclk));
	jdff dff_B_VPvmGoH24_2(.din(n1383),.dout(w_dff_B_VPvmGoH24_2),.clk(gclk));
	jdff dff_B_8FBpPTDB6_2(.din(w_dff_B_VPvmGoH24_2),.dout(w_dff_B_8FBpPTDB6_2),.clk(gclk));
	jdff dff_B_jmc6jy0Q9_2(.din(w_dff_B_8FBpPTDB6_2),.dout(w_dff_B_jmc6jy0Q9_2),.clk(gclk));
	jdff dff_B_ya44IFzw8_2(.din(w_dff_B_jmc6jy0Q9_2),.dout(w_dff_B_ya44IFzw8_2),.clk(gclk));
	jdff dff_B_6rUjq6ZQ4_2(.din(w_dff_B_ya44IFzw8_2),.dout(w_dff_B_6rUjq6ZQ4_2),.clk(gclk));
	jdff dff_B_rVlMZDtL8_2(.din(w_dff_B_6rUjq6ZQ4_2),.dout(w_dff_B_rVlMZDtL8_2),.clk(gclk));
	jdff dff_B_SVnO8GHo7_2(.din(w_dff_B_rVlMZDtL8_2),.dout(w_dff_B_SVnO8GHo7_2),.clk(gclk));
	jdff dff_B_yxSeJoTe5_2(.din(w_dff_B_SVnO8GHo7_2),.dout(w_dff_B_yxSeJoTe5_2),.clk(gclk));
	jdff dff_B_TTzUi0Sw7_2(.din(w_dff_B_yxSeJoTe5_2),.dout(w_dff_B_TTzUi0Sw7_2),.clk(gclk));
	jdff dff_B_BLNBaMqb2_2(.din(w_dff_B_TTzUi0Sw7_2),.dout(w_dff_B_BLNBaMqb2_2),.clk(gclk));
	jdff dff_B_qXrdNVGE2_2(.din(w_dff_B_BLNBaMqb2_2),.dout(w_dff_B_qXrdNVGE2_2),.clk(gclk));
	jdff dff_B_5f7cjCv48_2(.din(w_dff_B_qXrdNVGE2_2),.dout(w_dff_B_5f7cjCv48_2),.clk(gclk));
	jdff dff_B_KeOJ60LY6_2(.din(w_dff_B_5f7cjCv48_2),.dout(w_dff_B_KeOJ60LY6_2),.clk(gclk));
	jdff dff_B_XIIP9E6T4_2(.din(w_dff_B_KeOJ60LY6_2),.dout(w_dff_B_XIIP9E6T4_2),.clk(gclk));
	jdff dff_B_e44LNbve0_2(.din(w_dff_B_XIIP9E6T4_2),.dout(w_dff_B_e44LNbve0_2),.clk(gclk));
	jdff dff_B_pSTBK2IA9_2(.din(n1382),.dout(w_dff_B_pSTBK2IA9_2),.clk(gclk));
	jdff dff_B_gUWPyqyB6_2(.din(w_dff_B_pSTBK2IA9_2),.dout(w_dff_B_gUWPyqyB6_2),.clk(gclk));
	jdff dff_B_1xTkYIv49_2(.din(w_dff_B_gUWPyqyB6_2),.dout(w_dff_B_1xTkYIv49_2),.clk(gclk));
	jdff dff_B_EnfHMm6L9_2(.din(w_dff_B_1xTkYIv49_2),.dout(w_dff_B_EnfHMm6L9_2),.clk(gclk));
	jdff dff_B_sFJ9tXPQ9_2(.din(w_dff_B_EnfHMm6L9_2),.dout(w_dff_B_sFJ9tXPQ9_2),.clk(gclk));
	jdff dff_B_vp5o16l02_2(.din(w_dff_B_sFJ9tXPQ9_2),.dout(w_dff_B_vp5o16l02_2),.clk(gclk));
	jdff dff_B_DlAJR0Oy0_2(.din(w_dff_B_vp5o16l02_2),.dout(w_dff_B_DlAJR0Oy0_2),.clk(gclk));
	jdff dff_B_VCfUbysu6_2(.din(w_dff_B_DlAJR0Oy0_2),.dout(w_dff_B_VCfUbysu6_2),.clk(gclk));
	jdff dff_B_lrtzWRUR1_2(.din(w_dff_B_VCfUbysu6_2),.dout(w_dff_B_lrtzWRUR1_2),.clk(gclk));
	jdff dff_B_rpekBJZO8_2(.din(w_dff_B_lrtzWRUR1_2),.dout(w_dff_B_rpekBJZO8_2),.clk(gclk));
	jdff dff_B_VvlGChyo2_2(.din(w_dff_B_rpekBJZO8_2),.dout(w_dff_B_VvlGChyo2_2),.clk(gclk));
	jdff dff_B_82CmETf92_2(.din(w_dff_B_VvlGChyo2_2),.dout(w_dff_B_82CmETf92_2),.clk(gclk));
	jdff dff_B_YIzQmC5H5_2(.din(w_dff_B_82CmETf92_2),.dout(w_dff_B_YIzQmC5H5_2),.clk(gclk));
	jdff dff_B_aydLwHWl5_2(.din(w_dff_B_YIzQmC5H5_2),.dout(w_dff_B_aydLwHWl5_2),.clk(gclk));
	jdff dff_B_EmJgA1MC3_2(.din(w_dff_B_aydLwHWl5_2),.dout(w_dff_B_EmJgA1MC3_2),.clk(gclk));
	jdff dff_B_lqajwhXR8_2(.din(w_dff_B_EmJgA1MC3_2),.dout(w_dff_B_lqajwhXR8_2),.clk(gclk));
	jdff dff_B_GjFxFVhf7_2(.din(w_dff_B_lqajwhXR8_2),.dout(w_dff_B_GjFxFVhf7_2),.clk(gclk));
	jdff dff_B_D4V5DroH4_2(.din(n1381),.dout(w_dff_B_D4V5DroH4_2),.clk(gclk));
	jdff dff_B_JkXbNzCC9_1(.din(n1379),.dout(w_dff_B_JkXbNzCC9_1),.clk(gclk));
	jdff dff_B_hYkSZRMO2_2(.din(n1293),.dout(w_dff_B_hYkSZRMO2_2),.clk(gclk));
	jdff dff_B_kk2dACGn6_2(.din(w_dff_B_hYkSZRMO2_2),.dout(w_dff_B_kk2dACGn6_2),.clk(gclk));
	jdff dff_B_a37rvPZh4_2(.din(w_dff_B_kk2dACGn6_2),.dout(w_dff_B_a37rvPZh4_2),.clk(gclk));
	jdff dff_B_nlY0VBjh2_2(.din(w_dff_B_a37rvPZh4_2),.dout(w_dff_B_nlY0VBjh2_2),.clk(gclk));
	jdff dff_B_vUYkJgk47_2(.din(w_dff_B_nlY0VBjh2_2),.dout(w_dff_B_vUYkJgk47_2),.clk(gclk));
	jdff dff_B_lwe0PPRo7_2(.din(w_dff_B_vUYkJgk47_2),.dout(w_dff_B_lwe0PPRo7_2),.clk(gclk));
	jdff dff_B_ojwBDWI14_2(.din(w_dff_B_lwe0PPRo7_2),.dout(w_dff_B_ojwBDWI14_2),.clk(gclk));
	jdff dff_B_1NxNfpFi0_2(.din(w_dff_B_ojwBDWI14_2),.dout(w_dff_B_1NxNfpFi0_2),.clk(gclk));
	jdff dff_B_u11dyIK55_2(.din(w_dff_B_1NxNfpFi0_2),.dout(w_dff_B_u11dyIK55_2),.clk(gclk));
	jdff dff_B_iRMJOcA28_2(.din(w_dff_B_u11dyIK55_2),.dout(w_dff_B_iRMJOcA28_2),.clk(gclk));
	jdff dff_B_7NUR15Zs0_2(.din(w_dff_B_iRMJOcA28_2),.dout(w_dff_B_7NUR15Zs0_2),.clk(gclk));
	jdff dff_B_VtKaEXlg4_2(.din(w_dff_B_7NUR15Zs0_2),.dout(w_dff_B_VtKaEXlg4_2),.clk(gclk));
	jdff dff_B_3asc5Gvr4_2(.din(w_dff_B_VtKaEXlg4_2),.dout(w_dff_B_3asc5Gvr4_2),.clk(gclk));
	jdff dff_B_IjuRj1ww2_2(.din(w_dff_B_3asc5Gvr4_2),.dout(w_dff_B_IjuRj1ww2_2),.clk(gclk));
	jdff dff_B_rKVR8sWE1_2(.din(w_dff_B_IjuRj1ww2_2),.dout(w_dff_B_rKVR8sWE1_2),.clk(gclk));
	jdff dff_B_crnr4qrw6_1(.din(n1299),.dout(w_dff_B_crnr4qrw6_1),.clk(gclk));
	jdff dff_B_moMeQzNZ4_1(.din(w_dff_B_crnr4qrw6_1),.dout(w_dff_B_moMeQzNZ4_1),.clk(gclk));
	jdff dff_B_jArypyh02_2(.din(n1298),.dout(w_dff_B_jArypyh02_2),.clk(gclk));
	jdff dff_B_3EbBvGA42_2(.din(w_dff_B_jArypyh02_2),.dout(w_dff_B_3EbBvGA42_2),.clk(gclk));
	jdff dff_B_afahBYJG0_2(.din(w_dff_B_3EbBvGA42_2),.dout(w_dff_B_afahBYJG0_2),.clk(gclk));
	jdff dff_B_k2p4wguJ8_2(.din(w_dff_B_afahBYJG0_2),.dout(w_dff_B_k2p4wguJ8_2),.clk(gclk));
	jdff dff_B_NR3jfjt91_2(.din(w_dff_B_k2p4wguJ8_2),.dout(w_dff_B_NR3jfjt91_2),.clk(gclk));
	jdff dff_B_aPVnDS1Z4_2(.din(w_dff_B_NR3jfjt91_2),.dout(w_dff_B_aPVnDS1Z4_2),.clk(gclk));
	jdff dff_B_YXuXaoNM9_2(.din(w_dff_B_aPVnDS1Z4_2),.dout(w_dff_B_YXuXaoNM9_2),.clk(gclk));
	jdff dff_B_g6RJ1NVC7_2(.din(w_dff_B_YXuXaoNM9_2),.dout(w_dff_B_g6RJ1NVC7_2),.clk(gclk));
	jdff dff_B_gx6K9Wow9_2(.din(w_dff_B_g6RJ1NVC7_2),.dout(w_dff_B_gx6K9Wow9_2),.clk(gclk));
	jdff dff_B_TwhgTcSW8_2(.din(w_dff_B_gx6K9Wow9_2),.dout(w_dff_B_TwhgTcSW8_2),.clk(gclk));
	jdff dff_B_4g2faHve1_2(.din(w_dff_B_TwhgTcSW8_2),.dout(w_dff_B_4g2faHve1_2),.clk(gclk));
	jdff dff_B_Ki1nZEhn6_2(.din(w_dff_B_4g2faHve1_2),.dout(w_dff_B_Ki1nZEhn6_2),.clk(gclk));
	jdff dff_B_tegQGoKM7_2(.din(n1297),.dout(w_dff_B_tegQGoKM7_2),.clk(gclk));
	jdff dff_B_UgIDderV0_2(.din(w_dff_B_tegQGoKM7_2),.dout(w_dff_B_UgIDderV0_2),.clk(gclk));
	jdff dff_B_NXH9GbrM0_2(.din(w_dff_B_UgIDderV0_2),.dout(w_dff_B_NXH9GbrM0_2),.clk(gclk));
	jdff dff_B_Twdf0ORp8_2(.din(w_dff_B_NXH9GbrM0_2),.dout(w_dff_B_Twdf0ORp8_2),.clk(gclk));
	jdff dff_B_coGlQVZF5_2(.din(w_dff_B_Twdf0ORp8_2),.dout(w_dff_B_coGlQVZF5_2),.clk(gclk));
	jdff dff_B_4d6xiDjR5_2(.din(w_dff_B_coGlQVZF5_2),.dout(w_dff_B_4d6xiDjR5_2),.clk(gclk));
	jdff dff_B_9w8S3GlZ9_2(.din(w_dff_B_4d6xiDjR5_2),.dout(w_dff_B_9w8S3GlZ9_2),.clk(gclk));
	jdff dff_B_4pyJrmRF8_2(.din(w_dff_B_9w8S3GlZ9_2),.dout(w_dff_B_4pyJrmRF8_2),.clk(gclk));
	jdff dff_B_4EOU09hD8_2(.din(w_dff_B_4pyJrmRF8_2),.dout(w_dff_B_4EOU09hD8_2),.clk(gclk));
	jdff dff_B_POmBTAvC7_2(.din(w_dff_B_4EOU09hD8_2),.dout(w_dff_B_POmBTAvC7_2),.clk(gclk));
	jdff dff_B_WxnuOMZF6_2(.din(w_dff_B_POmBTAvC7_2),.dout(w_dff_B_WxnuOMZF6_2),.clk(gclk));
	jdff dff_B_BmwIfJcz5_2(.din(w_dff_B_WxnuOMZF6_2),.dout(w_dff_B_BmwIfJcz5_2),.clk(gclk));
	jdff dff_B_cab2Nc215_2(.din(w_dff_B_BmwIfJcz5_2),.dout(w_dff_B_cab2Nc215_2),.clk(gclk));
	jdff dff_B_QhMgLiIT7_2(.din(w_dff_B_cab2Nc215_2),.dout(w_dff_B_QhMgLiIT7_2),.clk(gclk));
	jdff dff_B_JjO1MDJb9_2(.din(n1296),.dout(w_dff_B_JjO1MDJb9_2),.clk(gclk));
	jdff dff_B_6OoSuzZF7_1(.din(n1294),.dout(w_dff_B_6OoSuzZF7_1),.clk(gclk));
	jdff dff_B_fX8bTeqw0_2(.din(n1203),.dout(w_dff_B_fX8bTeqw0_2),.clk(gclk));
	jdff dff_B_vpfPPq250_2(.din(w_dff_B_fX8bTeqw0_2),.dout(w_dff_B_vpfPPq250_2),.clk(gclk));
	jdff dff_B_BQqIShCe6_2(.din(w_dff_B_vpfPPq250_2),.dout(w_dff_B_BQqIShCe6_2),.clk(gclk));
	jdff dff_B_lRZTpFWs1_2(.din(w_dff_B_BQqIShCe6_2),.dout(w_dff_B_lRZTpFWs1_2),.clk(gclk));
	jdff dff_B_x1YsHaaj2_2(.din(w_dff_B_lRZTpFWs1_2),.dout(w_dff_B_x1YsHaaj2_2),.clk(gclk));
	jdff dff_B_TuaFXoE17_2(.din(w_dff_B_x1YsHaaj2_2),.dout(w_dff_B_TuaFXoE17_2),.clk(gclk));
	jdff dff_B_pPON8ijK0_2(.din(w_dff_B_TuaFXoE17_2),.dout(w_dff_B_pPON8ijK0_2),.clk(gclk));
	jdff dff_B_3bezBXOB5_2(.din(w_dff_B_pPON8ijK0_2),.dout(w_dff_B_3bezBXOB5_2),.clk(gclk));
	jdff dff_B_6NHPVkwv5_2(.din(w_dff_B_3bezBXOB5_2),.dout(w_dff_B_6NHPVkwv5_2),.clk(gclk));
	jdff dff_B_rBMRZ5Du1_2(.din(w_dff_B_6NHPVkwv5_2),.dout(w_dff_B_rBMRZ5Du1_2),.clk(gclk));
	jdff dff_B_Sa5id6kp7_2(.din(w_dff_B_rBMRZ5Du1_2),.dout(w_dff_B_Sa5id6kp7_2),.clk(gclk));
	jdff dff_B_eGtqjqZM3_2(.din(w_dff_B_Sa5id6kp7_2),.dout(w_dff_B_eGtqjqZM3_2),.clk(gclk));
	jdff dff_B_xrv1WuOu5_2(.din(n1208),.dout(w_dff_B_xrv1WuOu5_2),.clk(gclk));
	jdff dff_B_Voje3uex4_2(.din(w_dff_B_xrv1WuOu5_2),.dout(w_dff_B_Voje3uex4_2),.clk(gclk));
	jdff dff_B_XAc0eTrz4_2(.din(w_dff_B_Voje3uex4_2),.dout(w_dff_B_XAc0eTrz4_2),.clk(gclk));
	jdff dff_B_KwLOO7oH1_2(.din(w_dff_B_XAc0eTrz4_2),.dout(w_dff_B_KwLOO7oH1_2),.clk(gclk));
	jdff dff_B_IdU6J5MB4_2(.din(w_dff_B_KwLOO7oH1_2),.dout(w_dff_B_IdU6J5MB4_2),.clk(gclk));
	jdff dff_B_iExQuYZR4_2(.din(w_dff_B_IdU6J5MB4_2),.dout(w_dff_B_iExQuYZR4_2),.clk(gclk));
	jdff dff_B_3brHcHxm4_2(.din(w_dff_B_iExQuYZR4_2),.dout(w_dff_B_3brHcHxm4_2),.clk(gclk));
	jdff dff_B_4wJbf1jX4_2(.din(w_dff_B_3brHcHxm4_2),.dout(w_dff_B_4wJbf1jX4_2),.clk(gclk));
	jdff dff_B_v33DHjVQ4_2(.din(w_dff_B_4wJbf1jX4_2),.dout(w_dff_B_v33DHjVQ4_2),.clk(gclk));
	jdff dff_B_RhBT1oab0_2(.din(n1207),.dout(w_dff_B_RhBT1oab0_2),.clk(gclk));
	jdff dff_B_Pc6OwOEA5_2(.din(w_dff_B_RhBT1oab0_2),.dout(w_dff_B_Pc6OwOEA5_2),.clk(gclk));
	jdff dff_B_cPFS5UMl9_2(.din(w_dff_B_Pc6OwOEA5_2),.dout(w_dff_B_cPFS5UMl9_2),.clk(gclk));
	jdff dff_B_Mb4y08Yj5_2(.din(w_dff_B_cPFS5UMl9_2),.dout(w_dff_B_Mb4y08Yj5_2),.clk(gclk));
	jdff dff_B_RGmyYYux5_2(.din(w_dff_B_Mb4y08Yj5_2),.dout(w_dff_B_RGmyYYux5_2),.clk(gclk));
	jdff dff_B_fQ1m8iJV7_2(.din(w_dff_B_RGmyYYux5_2),.dout(w_dff_B_fQ1m8iJV7_2),.clk(gclk));
	jdff dff_B_lfb3DuC96_2(.din(w_dff_B_fQ1m8iJV7_2),.dout(w_dff_B_lfb3DuC96_2),.clk(gclk));
	jdff dff_B_LWfmRrg24_2(.din(w_dff_B_lfb3DuC96_2),.dout(w_dff_B_LWfmRrg24_2),.clk(gclk));
	jdff dff_B_cbHGpwvu8_2(.din(w_dff_B_LWfmRrg24_2),.dout(w_dff_B_cbHGpwvu8_2),.clk(gclk));
	jdff dff_B_DOCHpHWC7_2(.din(w_dff_B_cbHGpwvu8_2),.dout(w_dff_B_DOCHpHWC7_2),.clk(gclk));
	jdff dff_B_PtBSenI71_2(.din(w_dff_B_DOCHpHWC7_2),.dout(w_dff_B_PtBSenI71_2),.clk(gclk));
	jdff dff_B_qtCwMmqV7_2(.din(n1206),.dout(w_dff_B_qtCwMmqV7_2),.clk(gclk));
	jdff dff_B_1JPldOdX0_1(.din(n1204),.dout(w_dff_B_1JPldOdX0_1),.clk(gclk));
	jdff dff_B_t2RQxvvt5_2(.din(n1099),.dout(w_dff_B_t2RQxvvt5_2),.clk(gclk));
	jdff dff_B_E9dEHnKE3_2(.din(w_dff_B_t2RQxvvt5_2),.dout(w_dff_B_E9dEHnKE3_2),.clk(gclk));
	jdff dff_B_46rKKUJs4_2(.din(w_dff_B_E9dEHnKE3_2),.dout(w_dff_B_46rKKUJs4_2),.clk(gclk));
	jdff dff_B_Q9fo6tvq9_2(.din(w_dff_B_46rKKUJs4_2),.dout(w_dff_B_Q9fo6tvq9_2),.clk(gclk));
	jdff dff_B_vmcLBHZa6_2(.din(w_dff_B_Q9fo6tvq9_2),.dout(w_dff_B_vmcLBHZa6_2),.clk(gclk));
	jdff dff_B_M1cT6BMY3_2(.din(w_dff_B_vmcLBHZa6_2),.dout(w_dff_B_M1cT6BMY3_2),.clk(gclk));
	jdff dff_B_tE1xEeXB1_2(.din(w_dff_B_M1cT6BMY3_2),.dout(w_dff_B_tE1xEeXB1_2),.clk(gclk));
	jdff dff_B_ZocsiWzv7_2(.din(w_dff_B_tE1xEeXB1_2),.dout(w_dff_B_ZocsiWzv7_2),.clk(gclk));
	jdff dff_B_tmJgp1tV3_2(.din(w_dff_B_ZocsiWzv7_2),.dout(w_dff_B_tmJgp1tV3_2),.clk(gclk));
	jdff dff_A_Bpoorvzm5_0(.dout(w_n1110_0[0]),.din(w_dff_A_Bpoorvzm5_0),.clk(gclk));
	jdff dff_A_vg1N7GSx6_0(.dout(w_dff_A_Bpoorvzm5_0),.din(w_dff_A_vg1N7GSx6_0),.clk(gclk));
	jdff dff_B_BjpRqFhs3_2(.din(n1110),.dout(w_dff_B_BjpRqFhs3_2),.clk(gclk));
	jdff dff_B_LsD0lV718_2(.din(w_dff_B_BjpRqFhs3_2),.dout(w_dff_B_LsD0lV718_2),.clk(gclk));
	jdff dff_B_VC3sdodO5_1(.din(n1104),.dout(w_dff_B_VC3sdodO5_1),.clk(gclk));
	jdff dff_B_AQKaMuAp6_1(.din(w_dff_B_VC3sdodO5_1),.dout(w_dff_B_AQKaMuAp6_1),.clk(gclk));
	jdff dff_B_jPNVT33D5_1(.din(w_dff_B_AQKaMuAp6_1),.dout(w_dff_B_jPNVT33D5_1),.clk(gclk));
	jdff dff_B_bUMTWNEB1_1(.din(w_dff_B_jPNVT33D5_1),.dout(w_dff_B_bUMTWNEB1_1),.clk(gclk));
	jdff dff_B_eo89BVpV8_1(.din(n1105),.dout(w_dff_B_eo89BVpV8_1),.clk(gclk));
	jdff dff_A_MpFN9kOz1_1(.dout(w_G307gat_2[1]),.din(w_dff_A_MpFN9kOz1_1),.clk(gclk));
	jdff dff_A_Dnggmsxb1_1(.dout(w_dff_A_MpFN9kOz1_1),.din(w_dff_A_Dnggmsxb1_1),.clk(gclk));
	jdff dff_A_RD7anr8l3_1(.dout(w_dff_A_Dnggmsxb1_1),.din(w_dff_A_RD7anr8l3_1),.clk(gclk));
	jdff dff_A_OX52VQV68_1(.dout(w_dff_A_RD7anr8l3_1),.din(w_dff_A_OX52VQV68_1),.clk(gclk));
	jdff dff_A_D8rU4KIX2_1(.dout(w_dff_A_OX52VQV68_1),.din(w_dff_A_D8rU4KIX2_1),.clk(gclk));
	jdff dff_B_unvMkBRI7_2(.din(n1103),.dout(w_dff_B_unvMkBRI7_2),.clk(gclk));
	jdff dff_B_GzSO49xg9_2(.din(w_dff_B_unvMkBRI7_2),.dout(w_dff_B_GzSO49xg9_2),.clk(gclk));
	jdff dff_B_3SvcwYWA5_2(.din(w_dff_B_GzSO49xg9_2),.dout(w_dff_B_3SvcwYWA5_2),.clk(gclk));
	jdff dff_B_xoYT6RqI5_2(.din(w_dff_B_3SvcwYWA5_2),.dout(w_dff_B_xoYT6RqI5_2),.clk(gclk));
	jdff dff_B_Lo8sqDnR7_2(.din(w_dff_B_xoYT6RqI5_2),.dout(w_dff_B_Lo8sqDnR7_2),.clk(gclk));
	jdff dff_B_cYi2rSmd7_2(.din(w_dff_B_Lo8sqDnR7_2),.dout(w_dff_B_cYi2rSmd7_2),.clk(gclk));
	jdff dff_B_d8c3X7ZS7_2(.din(w_dff_B_cYi2rSmd7_2),.dout(w_dff_B_d8c3X7ZS7_2),.clk(gclk));
	jdff dff_B_Rw9ReYqf4_2(.din(w_dff_B_d8c3X7ZS7_2),.dout(w_dff_B_Rw9ReYqf4_2),.clk(gclk));
	jdff dff_B_8Y9hUj1G5_2(.din(n1102),.dout(w_dff_B_8Y9hUj1G5_2),.clk(gclk));
	jdff dff_B_04222BGw5_1(.din(n1100),.dout(w_dff_B_04222BGw5_1),.clk(gclk));
	jdff dff_B_6f8sRSvr3_2(.din(n1001),.dout(w_dff_B_6f8sRSvr3_2),.clk(gclk));
	jdff dff_B_jGOQpKDW6_2(.din(w_dff_B_6f8sRSvr3_2),.dout(w_dff_B_jGOQpKDW6_2),.clk(gclk));
	jdff dff_B_9LZahrSn2_2(.din(w_dff_B_jGOQpKDW6_2),.dout(w_dff_B_9LZahrSn2_2),.clk(gclk));
	jdff dff_B_VUMRSgNd1_2(.din(w_dff_B_9LZahrSn2_2),.dout(w_dff_B_VUMRSgNd1_2),.clk(gclk));
	jdff dff_B_UPPjNxRn4_2(.din(w_dff_B_VUMRSgNd1_2),.dout(w_dff_B_UPPjNxRn4_2),.clk(gclk));
	jdff dff_B_ImuegOsW8_2(.din(w_dff_B_UPPjNxRn4_2),.dout(w_dff_B_ImuegOsW8_2),.clk(gclk));
	jdff dff_B_qsysMGag1_2(.din(n1010),.dout(w_dff_B_qsysMGag1_2),.clk(gclk));
	jdff dff_B_PYu0KVco4_2(.din(w_dff_B_qsysMGag1_2),.dout(w_dff_B_PYu0KVco4_2),.clk(gclk));
	jdff dff_B_fl1OZwDh9_2(.din(w_dff_B_PYu0KVco4_2),.dout(w_dff_B_fl1OZwDh9_2),.clk(gclk));
	jdff dff_B_RUO3PTNq1_2(.din(w_dff_B_fl1OZwDh9_2),.dout(w_dff_B_RUO3PTNq1_2),.clk(gclk));
	jdff dff_A_G8AbBSSj2_0(.dout(w_n1008_0[0]),.din(w_dff_A_G8AbBSSj2_0),.clk(gclk));
	jdff dff_A_CBBvRGVn6_0(.dout(w_dff_A_G8AbBSSj2_0),.din(w_dff_A_CBBvRGVn6_0),.clk(gclk));
	jdff dff_A_be4tAm5B8_0(.dout(w_n793_0[0]),.din(w_dff_A_be4tAm5B8_0),.clk(gclk));
	jdff dff_A_oqTUZVoI6_1(.dout(w_n1006_0[1]),.din(w_dff_A_oqTUZVoI6_1),.clk(gclk));
	jdff dff_B_w8bbQZS44_1(.din(n1002),.dout(w_dff_B_w8bbQZS44_1),.clk(gclk));
	jdff dff_B_gOLdFHBa4_1(.din(w_dff_B_w8bbQZS44_1),.dout(w_dff_B_gOLdFHBa4_1),.clk(gclk));
	jdff dff_B_TVSLvhh41_1(.din(w_dff_B_gOLdFHBa4_1),.dout(w_dff_B_TVSLvhh41_1),.clk(gclk));
	jdff dff_B_NWt7fI1i0_1(.din(w_dff_B_TVSLvhh41_1),.dout(w_dff_B_NWt7fI1i0_1),.clk(gclk));
	jdff dff_B_rAaU6uUB6_0(.din(n905),.dout(w_dff_B_rAaU6uUB6_0),.clk(gclk));
	jdff dff_A_nbVdUsEx9_0(.dout(w_n903_0[0]),.din(w_dff_A_nbVdUsEx9_0),.clk(gclk));
	jdff dff_A_zLgoNo255_0(.dout(w_dff_A_nbVdUsEx9_0),.din(w_dff_A_zLgoNo255_0),.clk(gclk));
	jdff dff_A_6V0MbwZf0_1(.dout(w_n901_0[1]),.din(w_dff_A_6V0MbwZf0_1),.clk(gclk));
	jdff dff_A_idjRVIPl0_0(.dout(w_n695_0[0]),.din(w_dff_A_idjRVIPl0_0),.clk(gclk));
	jdff dff_A_r6vr8Qko8_0(.dout(w_dff_A_idjRVIPl0_0),.din(w_dff_A_r6vr8Qko8_0),.clk(gclk));
	jdff dff_B_PZUfM55S1_2(.din(n898),.dout(w_dff_B_PZUfM55S1_2),.clk(gclk));
	jdff dff_A_BXoSWlfi3_1(.dout(w_n896_0[1]),.din(w_dff_A_BXoSWlfi3_1),.clk(gclk));
	jdff dff_A_ztGCcWEc3_1(.dout(w_dff_A_BXoSWlfi3_1),.din(w_dff_A_ztGCcWEc3_1),.clk(gclk));
	jdff dff_A_1eNyPkSg7_1(.dout(w_dff_A_ztGCcWEc3_1),.din(w_dff_A_1eNyPkSg7_1),.clk(gclk));
	jdff dff_A_WQZtJbXd3_1(.dout(w_dff_A_1eNyPkSg7_1),.din(w_dff_A_WQZtJbXd3_1),.clk(gclk));
endmodule

