// Benchmark "c6288" written by ABC on Sun May 24 21:38:16 2020

module rf_c6288 ( 
    G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat,
    G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat,
    G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat,
    G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat,
    G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat,
    G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat,
    G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat,
    G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat,
    G6270gat, G6280gat, G6287gat, G6288gat  );
  input  G1gat, G18gat, G35gat, G52gat, G69gat, G86gat, G103gat, G120gat,
    G137gat, G154gat, G171gat, G188gat, G205gat, G222gat, G239gat, G256gat,
    G273gat, G290gat, G307gat, G324gat, G341gat, G358gat, G375gat, G392gat,
    G409gat, G426gat, G443gat, G460gat, G477gat, G494gat, G511gat, G528gat;
  output G545gat, G1581gat, G1901gat, G2223gat, G2548gat, G2877gat, G3211gat,
    G3552gat, G3895gat, G4241gat, G4591gat, G4946gat, G5308gat, G5672gat,
    G5971gat, G6123gat, G6150gat, G6160gat, G6170gat, G6180gat, G6190gat,
    G6200gat, G6210gat, G6220gat, G6230gat, G6240gat, G6250gat, G6260gat,
    G6270gat, G6280gat, G6287gat, G6288gat;
  wire n65, n66, n67, n68, n69, n70, n72, n73, n74, n75, n76, n77, n78, n79,
    n80, n81, n82, n83, n84, n85, n86, n87, n89, n90, n91, n92, n93, n94,
    n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
    n107, n108, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119,
    n120, n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
    n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
    n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
    n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
    n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
    n181, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
    n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
    n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
    n218, n219, n220, n221, n222, n223, n224, n226, n227, n228, n229, n230,
    n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
    n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
    n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
    n267, n268, n269, n270, n271, n272, n273, n274, n275, n277, n278, n279,
    n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
    n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
    n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
    n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
    n328, n329, n330, n331, n332, n333, n335, n336, n337, n338, n339, n340,
    n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
    n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
    n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
    n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387, n388,
    n389, n390, n391, n392, n393, n394, n395, n396, n397, n399, n400, n401,
    n402, n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
    n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
    n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
    n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448, n449,
    n450, n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
    n462, n463, n464, n465, n466, n467, n468, n469, n471, n472, n473, n474,
    n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
    n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497, n498,
    n499, n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
    n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521, n522,
    n523, n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
    n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
    n547, n548, n550, n551, n552, n553, n554, n555, n556, n557, n558, n559,
    n560, n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
    n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
    n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
    n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
    n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618, n619,
    n620, n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
    n632, n633, n634, n636, n637, n638, n639, n640, n641, n642, n643, n644,
    n645, n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
    n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
    n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679, n680,
    n681, n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
    n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
    n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
    n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n729,
    n730, n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
    n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752, n753,
    n754, n755, n756, n757, n758, n759, n760, n761, n762, n763, n764, n765,
    n766, n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
    n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
    n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800, n801,
    n802, n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
    n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
    n826, n827, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
    n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849, n850,
    n851, n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
    n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
    n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885, n886,
    n887, n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
    n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
    n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921, n922,
    n923, n924, n925, n926, n927, n928, n929, n930, n931, n932, n934, n935,
    n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
    n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
    n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970, n971,
    n972, n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
    n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
    n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
    n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
    n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
    n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
    n1036, n1037, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
    n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
    n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
    n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
    n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
    n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
    n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
    n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
    n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
    n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
    n1137, n1138, n1139, n1140, n1141, n1142, n1144, n1145, n1146, n1147,
    n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
    n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
    n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
    n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
    n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
    n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
    n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
    n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
    n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
    n1238, n1239, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
    n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
    n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
    n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
    n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
    n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
    n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
    n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
    n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1329,
    n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
    n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
    n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
    n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
    n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
    n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
    n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
    n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
    n1410, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
    n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
    n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
    n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
    n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
    n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
    n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
    n1481, n1482, n1483, n1484, n1485, n1486, n1488, n1489, n1490, n1491,
    n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
    n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
    n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
    n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
    n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
    n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
    n1552, n1553, n1554, n1555, n1557, n1558, n1559, n1560, n1561, n1562,
    n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
    n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
    n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
    n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
    n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
    n1613, n1614, n1615, n1616, n1617, n1619, n1620, n1621, n1622, n1623,
    n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
    n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
    n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
    n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
    n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1674,
    n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
    n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
    n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
    n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
    n1715, n1716, n1717, n1718, n1719, n1720, n1722, n1723, n1724, n1725,
    n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
    n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
    n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
    n1756, n1757, n1758, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
    n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
    n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
    n1787, n1788, n1789, n1790, n1791, n1793, n1794, n1795, n1796, n1797,
    n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
    n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
    n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
    n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1838, n1839,
    n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
    n1850, n1851;
  jand g0000(.dina(G273gat), .dinb(G1gat), .dout(G545gat));
  jand g0001(.dina(G273gat), .dinb(G18gat), .dout(n65));
  jand g0002(.dina(G290gat), .dinb(G1gat), .dout(n66));
  jor  g0003(.dina(n66), .dinb(n65), .dout(n67));
  jand g0004(.dina(G290gat), .dinb(G18gat), .dout(n68));
  jand g0005(.dina(n68), .dinb(G545gat), .dout(n69));
  jnot g0006(.din(n69), .dout(n70));
  jand g0007(.dina(n70), .dinb(n67), .dout(G1581gat));
  jand g0008(.dina(G307gat), .dinb(G1gat), .dout(n72));
  jnot g0009(.din(n72), .dout(n73));
  jnot g0010(.din(G18gat), .dout(n74));
  jnot g0011(.din(G290gat), .dout(n75));
  jor  g0012(.dina(n75), .dinb(n74), .dout(n76));
  jnot g0013(.din(G35gat), .dout(n77));
  jnot g0014(.din(G273gat), .dout(n78));
  jor  g0015(.dina(n78), .dinb(n77), .dout(n79));
  jand g0016(.dina(n79), .dinb(n76), .dout(n80));
  jand g0017(.dina(G290gat), .dinb(G35gat), .dout(n81));
  jand g0018(.dina(n81), .dinb(n65), .dout(n82));
  jor  g0019(.dina(n82), .dinb(n80), .dout(n83));
  jand g0020(.dina(n83), .dinb(n70), .dout(n84));
  jnot g0021(.din(n82), .dout(n85));
  jand g0022(.dina(n85), .dinb(n69), .dout(n86));
  jor  g0023(.dina(n86), .dinb(n84), .dout(n87));
  jxor g0024(.dina(n87), .dinb(n73), .dout(G1901gat));
  jand g0025(.dina(G324gat), .dinb(G1gat), .dout(n89));
  jnot g0026(.din(n89), .dout(n90));
  jnot g0027(.din(n84), .dout(n91));
  jor  g0028(.dina(n87), .dinb(n72), .dout(n92));
  jand g0029(.dina(n92), .dinb(n91), .dout(n93));
  jand g0030(.dina(G307gat), .dinb(G18gat), .dout(n94));
  jnot g0031(.din(n94), .dout(n95));
  jand g0032(.dina(G273gat), .dinb(G52gat), .dout(n96));
  jor  g0033(.dina(n96), .dinb(n81), .dout(n97));
  jand g0034(.dina(G273gat), .dinb(G35gat), .dout(n98));
  jand g0035(.dina(G290gat), .dinb(G52gat), .dout(n99));
  jand g0036(.dina(n99), .dinb(n98), .dout(n100));
  jnot g0037(.din(n100), .dout(n101));
  jand g0038(.dina(n101), .dinb(n97), .dout(n102));
  jor  g0039(.dina(n102), .dinb(n82), .dout(n103));
  jand g0040(.dina(n101), .dinb(n82), .dout(n104));
  jnot g0041(.din(n104), .dout(n105));
  jand g0042(.dina(n105), .dinb(n103), .dout(n106));
  jxor g0043(.dina(n106), .dinb(n95), .dout(n107));
  jxor g0044(.dina(n107), .dinb(n93), .dout(n108));
  jxor g0045(.dina(n108), .dinb(n90), .dout(G2223gat));
  jand g0046(.dina(G341gat), .dinb(G1gat), .dout(n110));
  jnot g0047(.din(n110), .dout(n111));
  jnot g0048(.din(n107), .dout(n112));
  jor  g0049(.dina(n112), .dinb(n93), .dout(n113));
  jor  g0050(.dina(n108), .dinb(n89), .dout(n114));
  jand g0051(.dina(n114), .dinb(n113), .dout(n115));
  jand g0052(.dina(G324gat), .dinb(G18gat), .dout(n116));
  jnot g0053(.din(n116), .dout(n117));
  jor  g0054(.dina(n75), .dinb(n77), .dout(n118));
  jnot g0055(.din(G52gat), .dout(n119));
  jor  g0056(.dina(n78), .dinb(n119), .dout(n120));
  jand g0057(.dina(n120), .dinb(n118), .dout(n121));
  jor  g0058(.dina(n100), .dinb(n121), .dout(n122));
  jand g0059(.dina(n122), .dinb(n85), .dout(n123));
  jor  g0060(.dina(n104), .dinb(n123), .dout(n124));
  jor  g0061(.dina(n124), .dinb(n94), .dout(n125));
  jand g0062(.dina(n125), .dinb(n103), .dout(n126));
  jand g0063(.dina(G307gat), .dinb(G35gat), .dout(n127));
  jnot g0064(.din(n127), .dout(n128));
  jand g0065(.dina(G273gat), .dinb(G69gat), .dout(n129));
  jor  g0066(.dina(n129), .dinb(n99), .dout(n130));
  jand g0067(.dina(G290gat), .dinb(G69gat), .dout(n131));
  jand g0068(.dina(n131), .dinb(n96), .dout(n132));
  jnot g0069(.din(n132), .dout(n133));
  jand g0070(.dina(n133), .dinb(n130), .dout(n134));
  jor  g0071(.dina(n134), .dinb(n100), .dout(n135));
  jand g0072(.dina(n133), .dinb(n100), .dout(n136));
  jnot g0073(.din(n136), .dout(n137));
  jand g0074(.dina(n137), .dinb(n135), .dout(n138));
  jxor g0075(.dina(n138), .dinb(n128), .dout(n139));
  jnot g0076(.din(n139), .dout(n140));
  jxor g0077(.dina(n140), .dinb(n126), .dout(n141));
  jxor g0078(.dina(n141), .dinb(n117), .dout(n142));
  jxor g0079(.dina(n142), .dinb(n115), .dout(n143));
  jxor g0080(.dina(n143), .dinb(n111), .dout(G2548gat));
  jand g0081(.dina(G358gat), .dinb(G1gat), .dout(n145));
  jnot g0082(.din(n145), .dout(n146));
  jnot g0083(.din(n142), .dout(n147));
  jor  g0084(.dina(n147), .dinb(n115), .dout(n148));
  jor  g0085(.dina(n143), .dinb(n110), .dout(n149));
  jand g0086(.dina(n149), .dinb(n148), .dout(n150));
  jand g0087(.dina(G341gat), .dinb(G18gat), .dout(n151));
  jnot g0088(.din(n151), .dout(n152));
  jor  g0089(.dina(n140), .dinb(n126), .dout(n153));
  jxor g0090(.dina(n139), .dinb(n126), .dout(n154));
  jor  g0091(.dina(n154), .dinb(n116), .dout(n155));
  jand g0092(.dina(n155), .dinb(n153), .dout(n156));
  jand g0093(.dina(G324gat), .dinb(G35gat), .dout(n157));
  jnot g0094(.din(n157), .dout(n158));
  jnot g0095(.din(n130), .dout(n159));
  jor  g0096(.dina(n132), .dinb(n159), .dout(n160));
  jand g0097(.dina(n160), .dinb(n101), .dout(n161));
  jand g0098(.dina(n138), .dinb(n128), .dout(n162));
  jor  g0099(.dina(n162), .dinb(n161), .dout(n163));
  jand g0100(.dina(G307gat), .dinb(G52gat), .dout(n164));
  jnot g0101(.din(n164), .dout(n165));
  jand g0102(.dina(G273gat), .dinb(G86gat), .dout(n166));
  jor  g0103(.dina(n166), .dinb(n131), .dout(n167));
  jand g0104(.dina(G290gat), .dinb(G86gat), .dout(n168));
  jand g0105(.dina(n168), .dinb(n129), .dout(n169));
  jnot g0106(.din(n169), .dout(n170));
  jand g0107(.dina(n170), .dinb(n167), .dout(n171));
  jor  g0108(.dina(n171), .dinb(n132), .dout(n172));
  jor  g0109(.dina(n169), .dinb(n133), .dout(n173));
  jand g0110(.dina(n173), .dinb(n172), .dout(n174));
  jxor g0111(.dina(n174), .dinb(n165), .dout(n175));
  jxor g0112(.dina(n175), .dinb(n163), .dout(n176));
  jxor g0113(.dina(n176), .dinb(n158), .dout(n177));
  jnot g0114(.din(n177), .dout(n178));
  jxor g0115(.dina(n178), .dinb(n156), .dout(n179));
  jxor g0116(.dina(n179), .dinb(n152), .dout(n180));
  jxor g0117(.dina(n180), .dinb(n150), .dout(n181));
  jxor g0118(.dina(n181), .dinb(n146), .dout(G2877gat));
  jand g0119(.dina(G375gat), .dinb(G1gat), .dout(n183));
  jnot g0120(.din(n183), .dout(n184));
  jnot g0121(.din(n180), .dout(n185));
  jor  g0122(.dina(n185), .dinb(n150), .dout(n186));
  jor  g0123(.dina(n181), .dinb(n145), .dout(n187));
  jand g0124(.dina(n187), .dinb(n186), .dout(n188));
  jand g0125(.dina(G358gat), .dinb(G18gat), .dout(n189));
  jnot g0126(.din(n189), .dout(n190));
  jor  g0127(.dina(n178), .dinb(n156), .dout(n191));
  jxor g0128(.dina(n177), .dinb(n156), .dout(n192));
  jor  g0129(.dina(n192), .dinb(n151), .dout(n193));
  jand g0130(.dina(n193), .dinb(n191), .dout(n194));
  jand g0131(.dina(G341gat), .dinb(G35gat), .dout(n195));
  jnot g0132(.din(n195), .dout(n196));
  jand g0133(.dina(n175), .dinb(n163), .dout(n197));
  jand g0134(.dina(n176), .dinb(n158), .dout(n198));
  jor  g0135(.dina(n198), .dinb(n197), .dout(n199));
  jand g0136(.dina(G324gat), .dinb(G52gat), .dout(n200));
  jnot g0137(.din(n200), .dout(n201));
  jnot g0138(.din(n172), .dout(n202));
  jand g0139(.dina(n174), .dinb(n165), .dout(n203));
  jor  g0140(.dina(n203), .dinb(n202), .dout(n204));
  jand g0141(.dina(G307gat), .dinb(G69gat), .dout(n205));
  jnot g0142(.din(n205), .dout(n206));
  jand g0143(.dina(G273gat), .dinb(G103gat), .dout(n207));
  jor  g0144(.dina(n207), .dinb(n168), .dout(n208));
  jand g0145(.dina(G290gat), .dinb(G103gat), .dout(n209));
  jand g0146(.dina(n209), .dinb(n166), .dout(n210));
  jnot g0147(.din(n210), .dout(n211));
  jand g0148(.dina(n211), .dinb(n208), .dout(n212));
  jor  g0149(.dina(n212), .dinb(n169), .dout(n213));
  jor  g0150(.dina(n210), .dinb(n170), .dout(n214));
  jand g0151(.dina(n214), .dinb(n213), .dout(n215));
  jxor g0152(.dina(n215), .dinb(n206), .dout(n216));
  jxor g0153(.dina(n216), .dinb(n204), .dout(n217));
  jxor g0154(.dina(n217), .dinb(n201), .dout(n218));
  jxor g0155(.dina(n218), .dinb(n199), .dout(n219));
  jxor g0156(.dina(n219), .dinb(n196), .dout(n220));
  jnot g0157(.din(n220), .dout(n221));
  jxor g0158(.dina(n221), .dinb(n194), .dout(n222));
  jxor g0159(.dina(n222), .dinb(n190), .dout(n223));
  jxor g0160(.dina(n223), .dinb(n188), .dout(n224));
  jxor g0161(.dina(n224), .dinb(n184), .dout(G3211gat));
  jand g0162(.dina(G392gat), .dinb(G1gat), .dout(n226));
  jnot g0163(.din(n226), .dout(n227));
  jnot g0164(.din(n223), .dout(n228));
  jor  g0165(.dina(n228), .dinb(n188), .dout(n229));
  jor  g0166(.dina(n224), .dinb(n183), .dout(n230));
  jand g0167(.dina(n230), .dinb(n229), .dout(n231));
  jand g0168(.dina(G375gat), .dinb(G18gat), .dout(n232));
  jnot g0169(.din(n232), .dout(n233));
  jor  g0170(.dina(n221), .dinb(n194), .dout(n234));
  jxor g0171(.dina(n220), .dinb(n194), .dout(n235));
  jor  g0172(.dina(n235), .dinb(n189), .dout(n236));
  jand g0173(.dina(n236), .dinb(n234), .dout(n237));
  jand g0174(.dina(G358gat), .dinb(G35gat), .dout(n238));
  jnot g0175(.din(n238), .dout(n239));
  jand g0176(.dina(n218), .dinb(n199), .dout(n240));
  jand g0177(.dina(n219), .dinb(n196), .dout(n241));
  jor  g0178(.dina(n241), .dinb(n240), .dout(n242));
  jand g0179(.dina(G341gat), .dinb(G52gat), .dout(n243));
  jnot g0180(.din(n243), .dout(n244));
  jand g0181(.dina(n216), .dinb(n204), .dout(n245));
  jand g0182(.dina(n217), .dinb(n201), .dout(n246));
  jor  g0183(.dina(n246), .dinb(n245), .dout(n247));
  jand g0184(.dina(G324gat), .dinb(G69gat), .dout(n248));
  jnot g0185(.din(n248), .dout(n249));
  jnot g0186(.din(n213), .dout(n250));
  jand g0187(.dina(n215), .dinb(n206), .dout(n251));
  jor  g0188(.dina(n251), .dinb(n250), .dout(n252));
  jand g0189(.dina(G307gat), .dinb(G86gat), .dout(n253));
  jnot g0190(.din(n253), .dout(n254));
  jand g0191(.dina(G273gat), .dinb(G120gat), .dout(n255));
  jor  g0192(.dina(n255), .dinb(n209), .dout(n256));
  jand g0193(.dina(G290gat), .dinb(G120gat), .dout(n257));
  jand g0194(.dina(n257), .dinb(n207), .dout(n258));
  jnot g0195(.din(n258), .dout(n259));
  jand g0196(.dina(n259), .dinb(n256), .dout(n260));
  jor  g0197(.dina(n260), .dinb(n210), .dout(n261));
  jand g0198(.dina(n259), .dinb(n210), .dout(n262));
  jnot g0199(.din(n262), .dout(n263));
  jand g0200(.dina(n263), .dinb(n261), .dout(n264));
  jxor g0201(.dina(n264), .dinb(n254), .dout(n265));
  jxor g0202(.dina(n265), .dinb(n252), .dout(n266));
  jxor g0203(.dina(n266), .dinb(n249), .dout(n267));
  jxor g0204(.dina(n267), .dinb(n247), .dout(n268));
  jxor g0205(.dina(n268), .dinb(n244), .dout(n269));
  jxor g0206(.dina(n269), .dinb(n242), .dout(n270));
  jxor g0207(.dina(n270), .dinb(n239), .dout(n271));
  jnot g0208(.din(n271), .dout(n272));
  jxor g0209(.dina(n272), .dinb(n237), .dout(n273));
  jxor g0210(.dina(n273), .dinb(n233), .dout(n274));
  jxor g0211(.dina(n274), .dinb(n231), .dout(n275));
  jxor g0212(.dina(n275), .dinb(n227), .dout(G3552gat));
  jand g0213(.dina(G409gat), .dinb(G1gat), .dout(n277));
  jnot g0214(.din(n277), .dout(n278));
  jnot g0215(.din(n274), .dout(n279));
  jor  g0216(.dina(n279), .dinb(n231), .dout(n280));
  jor  g0217(.dina(n275), .dinb(n226), .dout(n281));
  jand g0218(.dina(n281), .dinb(n280), .dout(n282));
  jand g0219(.dina(G392gat), .dinb(G18gat), .dout(n283));
  jnot g0220(.din(n283), .dout(n284));
  jor  g0221(.dina(n272), .dinb(n237), .dout(n285));
  jxor g0222(.dina(n271), .dinb(n237), .dout(n286));
  jor  g0223(.dina(n286), .dinb(n232), .dout(n287));
  jand g0224(.dina(n287), .dinb(n285), .dout(n288));
  jand g0225(.dina(G375gat), .dinb(G35gat), .dout(n289));
  jnot g0226(.din(n289), .dout(n290));
  jand g0227(.dina(n269), .dinb(n242), .dout(n291));
  jand g0228(.dina(n270), .dinb(n239), .dout(n292));
  jor  g0229(.dina(n292), .dinb(n291), .dout(n293));
  jand g0230(.dina(G358gat), .dinb(G52gat), .dout(n294));
  jnot g0231(.din(n294), .dout(n295));
  jand g0232(.dina(n267), .dinb(n247), .dout(n296));
  jand g0233(.dina(n268), .dinb(n244), .dout(n297));
  jor  g0234(.dina(n297), .dinb(n296), .dout(n298));
  jand g0235(.dina(G341gat), .dinb(G69gat), .dout(n299));
  jnot g0236(.din(n299), .dout(n300));
  jand g0237(.dina(n265), .dinb(n252), .dout(n301));
  jand g0238(.dina(n266), .dinb(n249), .dout(n302));
  jor  g0239(.dina(n302), .dinb(n301), .dout(n303));
  jand g0240(.dina(G324gat), .dinb(G86gat), .dout(n304));
  jnot g0241(.din(n304), .dout(n305));
  jnot g0242(.din(n261), .dout(n306));
  jand g0243(.dina(n264), .dinb(n254), .dout(n307));
  jor  g0244(.dina(n307), .dinb(n306), .dout(n308));
  jand g0245(.dina(G307gat), .dinb(G103gat), .dout(n309));
  jnot g0246(.din(n309), .dout(n310));
  jand g0247(.dina(G273gat), .dinb(G137gat), .dout(n311));
  jor  g0248(.dina(n311), .dinb(n257), .dout(n312));
  jand g0249(.dina(G290gat), .dinb(G137gat), .dout(n313));
  jand g0250(.dina(n313), .dinb(n255), .dout(n314));
  jnot g0251(.din(n314), .dout(n315));
  jand g0252(.dina(n315), .dinb(n312), .dout(n316));
  jor  g0253(.dina(n316), .dinb(n258), .dout(n317));
  jand g0254(.dina(n315), .dinb(n258), .dout(n318));
  jnot g0255(.din(n318), .dout(n319));
  jand g0256(.dina(n319), .dinb(n317), .dout(n320));
  jxor g0257(.dina(n320), .dinb(n310), .dout(n321));
  jxor g0258(.dina(n321), .dinb(n308), .dout(n322));
  jxor g0259(.dina(n322), .dinb(n305), .dout(n323));
  jxor g0260(.dina(n323), .dinb(n303), .dout(n324));
  jxor g0261(.dina(n324), .dinb(n300), .dout(n325));
  jxor g0262(.dina(n325), .dinb(n298), .dout(n326));
  jxor g0263(.dina(n326), .dinb(n295), .dout(n327));
  jxor g0264(.dina(n327), .dinb(n293), .dout(n328));
  jxor g0265(.dina(n328), .dinb(n290), .dout(n329));
  jnot g0266(.din(n329), .dout(n330));
  jxor g0267(.dina(n330), .dinb(n288), .dout(n331));
  jxor g0268(.dina(n331), .dinb(n284), .dout(n332));
  jxor g0269(.dina(n332), .dinb(n282), .dout(n333));
  jxor g0270(.dina(n333), .dinb(n278), .dout(G3895gat));
  jand g0271(.dina(G426gat), .dinb(G1gat), .dout(n335));
  jnot g0272(.din(n335), .dout(n336));
  jnot g0273(.din(n332), .dout(n337));
  jor  g0274(.dina(n337), .dinb(n282), .dout(n338));
  jor  g0275(.dina(n333), .dinb(n277), .dout(n339));
  jand g0276(.dina(n339), .dinb(n338), .dout(n340));
  jand g0277(.dina(G409gat), .dinb(G18gat), .dout(n341));
  jnot g0278(.din(n341), .dout(n342));
  jor  g0279(.dina(n330), .dinb(n288), .dout(n343));
  jxor g0280(.dina(n329), .dinb(n288), .dout(n344));
  jor  g0281(.dina(n344), .dinb(n283), .dout(n345));
  jand g0282(.dina(n345), .dinb(n343), .dout(n346));
  jand g0283(.dina(G392gat), .dinb(G35gat), .dout(n347));
  jnot g0284(.din(n347), .dout(n348));
  jand g0285(.dina(n327), .dinb(n293), .dout(n349));
  jand g0286(.dina(n328), .dinb(n290), .dout(n350));
  jor  g0287(.dina(n350), .dinb(n349), .dout(n351));
  jand g0288(.dina(G375gat), .dinb(G52gat), .dout(n352));
  jnot g0289(.din(n352), .dout(n353));
  jand g0290(.dina(n325), .dinb(n298), .dout(n354));
  jand g0291(.dina(n326), .dinb(n295), .dout(n355));
  jor  g0292(.dina(n355), .dinb(n354), .dout(n356));
  jand g0293(.dina(G358gat), .dinb(G69gat), .dout(n357));
  jnot g0294(.din(n357), .dout(n358));
  jand g0295(.dina(n323), .dinb(n303), .dout(n359));
  jand g0296(.dina(n324), .dinb(n300), .dout(n360));
  jor  g0297(.dina(n360), .dinb(n359), .dout(n361));
  jand g0298(.dina(G341gat), .dinb(G86gat), .dout(n362));
  jnot g0299(.din(n362), .dout(n363));
  jand g0300(.dina(n321), .dinb(n308), .dout(n364));
  jand g0301(.dina(n322), .dinb(n305), .dout(n365));
  jor  g0302(.dina(n365), .dinb(n364), .dout(n366));
  jand g0303(.dina(G324gat), .dinb(G103gat), .dout(n367));
  jnot g0304(.din(n367), .dout(n368));
  jnot g0305(.din(n317), .dout(n369));
  jand g0306(.dina(n320), .dinb(n310), .dout(n370));
  jor  g0307(.dina(n370), .dinb(n369), .dout(n371));
  jand g0308(.dina(G307gat), .dinb(G120gat), .dout(n372));
  jand g0309(.dina(G273gat), .dinb(G154gat), .dout(n373));
  jor  g0310(.dina(n373), .dinb(n313), .dout(n374));
  jand g0311(.dina(G290gat), .dinb(G154gat), .dout(n375));
  jand g0312(.dina(n375), .dinb(n311), .dout(n376));
  jnot g0313(.din(n376), .dout(n377));
  jand g0314(.dina(n377), .dinb(n374), .dout(n378));
  jor  g0315(.dina(n378), .dinb(n314), .dout(n379));
  jnot g0316(.din(n379), .dout(n380));
  jand g0317(.dina(n377), .dinb(n314), .dout(n381));
  jor  g0318(.dina(n381), .dinb(n380), .dout(n382));
  jxor g0319(.dina(n382), .dinb(n372), .dout(n383));
  jxor g0320(.dina(n383), .dinb(n371), .dout(n384));
  jxor g0321(.dina(n384), .dinb(n368), .dout(n385));
  jxor g0322(.dina(n385), .dinb(n366), .dout(n386));
  jxor g0323(.dina(n386), .dinb(n363), .dout(n387));
  jxor g0324(.dina(n387), .dinb(n361), .dout(n388));
  jxor g0325(.dina(n388), .dinb(n358), .dout(n389));
  jxor g0326(.dina(n389), .dinb(n356), .dout(n390));
  jxor g0327(.dina(n390), .dinb(n353), .dout(n391));
  jxor g0328(.dina(n391), .dinb(n351), .dout(n392));
  jxor g0329(.dina(n392), .dinb(n348), .dout(n393));
  jnot g0330(.din(n393), .dout(n394));
  jxor g0331(.dina(n394), .dinb(n346), .dout(n395));
  jxor g0332(.dina(n395), .dinb(n342), .dout(n396));
  jxor g0333(.dina(n396), .dinb(n340), .dout(n397));
  jxor g0334(.dina(n397), .dinb(n336), .dout(G4241gat));
  jand g0335(.dina(G443gat), .dinb(G1gat), .dout(n399));
  jnot g0336(.din(n399), .dout(n400));
  jnot g0337(.din(n396), .dout(n401));
  jor  g0338(.dina(n401), .dinb(n340), .dout(n402));
  jor  g0339(.dina(n397), .dinb(n335), .dout(n403));
  jand g0340(.dina(n403), .dinb(n402), .dout(n404));
  jand g0341(.dina(G426gat), .dinb(G18gat), .dout(n405));
  jnot g0342(.din(n405), .dout(n406));
  jor  g0343(.dina(n394), .dinb(n346), .dout(n407));
  jxor g0344(.dina(n393), .dinb(n346), .dout(n408));
  jor  g0345(.dina(n408), .dinb(n341), .dout(n409));
  jand g0346(.dina(n409), .dinb(n407), .dout(n410));
  jand g0347(.dina(G409gat), .dinb(G35gat), .dout(n411));
  jnot g0348(.din(n411), .dout(n412));
  jand g0349(.dina(n391), .dinb(n351), .dout(n413));
  jand g0350(.dina(n392), .dinb(n348), .dout(n414));
  jor  g0351(.dina(n414), .dinb(n413), .dout(n415));
  jand g0352(.dina(G392gat), .dinb(G52gat), .dout(n416));
  jnot g0353(.din(n416), .dout(n417));
  jand g0354(.dina(n389), .dinb(n356), .dout(n418));
  jand g0355(.dina(n390), .dinb(n353), .dout(n419));
  jor  g0356(.dina(n419), .dinb(n418), .dout(n420));
  jand g0357(.dina(G375gat), .dinb(G69gat), .dout(n421));
  jnot g0358(.din(n421), .dout(n422));
  jand g0359(.dina(n387), .dinb(n361), .dout(n423));
  jand g0360(.dina(n388), .dinb(n358), .dout(n424));
  jor  g0361(.dina(n424), .dinb(n423), .dout(n425));
  jand g0362(.dina(G358gat), .dinb(G86gat), .dout(n426));
  jnot g0363(.din(n426), .dout(n427));
  jand g0364(.dina(n385), .dinb(n366), .dout(n428));
  jand g0365(.dina(n386), .dinb(n363), .dout(n429));
  jor  g0366(.dina(n429), .dinb(n428), .dout(n430));
  jand g0367(.dina(G341gat), .dinb(G103gat), .dout(n431));
  jnot g0368(.din(n431), .dout(n432));
  jand g0369(.dina(n383), .dinb(n371), .dout(n433));
  jand g0370(.dina(n384), .dinb(n368), .dout(n434));
  jor  g0371(.dina(n434), .dinb(n433), .dout(n435));
  jand g0372(.dina(G324gat), .dinb(G120gat), .dout(n436));
  jnot g0373(.din(n436), .dout(n437));
  jnot g0374(.din(n372), .dout(n438));
  jnot g0375(.din(n382), .dout(n439));
  jand g0376(.dina(n439), .dinb(n438), .dout(n440));
  jor  g0377(.dina(n440), .dinb(n380), .dout(n441));
  jand g0378(.dina(G307gat), .dinb(G137gat), .dout(n442));
  jand g0379(.dina(G273gat), .dinb(G171gat), .dout(n443));
  jor  g0380(.dina(n443), .dinb(n375), .dout(n444));
  jand g0381(.dina(G290gat), .dinb(G171gat), .dout(n445));
  jand g0382(.dina(n445), .dinb(n373), .dout(n446));
  jnot g0383(.din(n446), .dout(n447));
  jand g0384(.dina(n447), .dinb(n444), .dout(n448));
  jor  g0385(.dina(n448), .dinb(n376), .dout(n449));
  jnot g0386(.din(n449), .dout(n450));
  jand g0387(.dina(n447), .dinb(n376), .dout(n451));
  jor  g0388(.dina(n451), .dinb(n450), .dout(n452));
  jxor g0389(.dina(n452), .dinb(n442), .dout(n453));
  jxor g0390(.dina(n453), .dinb(n441), .dout(n454));
  jxor g0391(.dina(n454), .dinb(n437), .dout(n455));
  jxor g0392(.dina(n455), .dinb(n435), .dout(n456));
  jxor g0393(.dina(n456), .dinb(n432), .dout(n457));
  jxor g0394(.dina(n457), .dinb(n430), .dout(n458));
  jxor g0395(.dina(n458), .dinb(n427), .dout(n459));
  jxor g0396(.dina(n459), .dinb(n425), .dout(n460));
  jxor g0397(.dina(n460), .dinb(n422), .dout(n461));
  jxor g0398(.dina(n461), .dinb(n420), .dout(n462));
  jxor g0399(.dina(n462), .dinb(n417), .dout(n463));
  jxor g0400(.dina(n463), .dinb(n415), .dout(n464));
  jxor g0401(.dina(n464), .dinb(n412), .dout(n465));
  jnot g0402(.din(n465), .dout(n466));
  jxor g0403(.dina(n466), .dinb(n410), .dout(n467));
  jxor g0404(.dina(n467), .dinb(n406), .dout(n468));
  jxor g0405(.dina(n468), .dinb(n404), .dout(n469));
  jxor g0406(.dina(n469), .dinb(n400), .dout(G4591gat));
  jand g0407(.dina(G460gat), .dinb(G1gat), .dout(n471));
  jnot g0408(.din(n471), .dout(n472));
  jnot g0409(.din(n468), .dout(n473));
  jor  g0410(.dina(n473), .dinb(n404), .dout(n474));
  jor  g0411(.dina(n469), .dinb(n399), .dout(n475));
  jand g0412(.dina(n475), .dinb(n474), .dout(n476));
  jand g0413(.dina(G443gat), .dinb(G18gat), .dout(n477));
  jnot g0414(.din(n477), .dout(n478));
  jor  g0415(.dina(n466), .dinb(n410), .dout(n479));
  jxor g0416(.dina(n465), .dinb(n410), .dout(n480));
  jor  g0417(.dina(n480), .dinb(n405), .dout(n481));
  jand g0418(.dina(n481), .dinb(n479), .dout(n482));
  jand g0419(.dina(G426gat), .dinb(G35gat), .dout(n483));
  jnot g0420(.din(n483), .dout(n484));
  jand g0421(.dina(n463), .dinb(n415), .dout(n485));
  jand g0422(.dina(n464), .dinb(n412), .dout(n486));
  jor  g0423(.dina(n486), .dinb(n485), .dout(n487));
  jand g0424(.dina(G409gat), .dinb(G52gat), .dout(n488));
  jnot g0425(.din(n488), .dout(n489));
  jand g0426(.dina(n461), .dinb(n420), .dout(n490));
  jand g0427(.dina(n462), .dinb(n417), .dout(n491));
  jor  g0428(.dina(n491), .dinb(n490), .dout(n492));
  jand g0429(.dina(G392gat), .dinb(G69gat), .dout(n493));
  jnot g0430(.din(n493), .dout(n494));
  jand g0431(.dina(n459), .dinb(n425), .dout(n495));
  jand g0432(.dina(n460), .dinb(n422), .dout(n496));
  jor  g0433(.dina(n496), .dinb(n495), .dout(n497));
  jand g0434(.dina(G375gat), .dinb(G86gat), .dout(n498));
  jnot g0435(.din(n498), .dout(n499));
  jand g0436(.dina(n457), .dinb(n430), .dout(n500));
  jand g0437(.dina(n458), .dinb(n427), .dout(n501));
  jor  g0438(.dina(n501), .dinb(n500), .dout(n502));
  jand g0439(.dina(G358gat), .dinb(G103gat), .dout(n503));
  jnot g0440(.din(n503), .dout(n504));
  jand g0441(.dina(n455), .dinb(n435), .dout(n505));
  jand g0442(.dina(n456), .dinb(n432), .dout(n506));
  jor  g0443(.dina(n506), .dinb(n505), .dout(n507));
  jand g0444(.dina(G341gat), .dinb(G120gat), .dout(n508));
  jnot g0445(.din(n508), .dout(n509));
  jand g0446(.dina(n453), .dinb(n441), .dout(n510));
  jand g0447(.dina(n454), .dinb(n437), .dout(n511));
  jor  g0448(.dina(n511), .dinb(n510), .dout(n512));
  jand g0449(.dina(G324gat), .dinb(G137gat), .dout(n513));
  jnot g0450(.din(n513), .dout(n514));
  jnot g0451(.din(n442), .dout(n515));
  jnot g0452(.din(n452), .dout(n516));
  jand g0453(.dina(n516), .dinb(n515), .dout(n517));
  jor  g0454(.dina(n517), .dinb(n450), .dout(n518));
  jand g0455(.dina(G307gat), .dinb(G154gat), .dout(n519));
  jand g0456(.dina(G273gat), .dinb(G188gat), .dout(n520));
  jor  g0457(.dina(n520), .dinb(n445), .dout(n521));
  jand g0458(.dina(G290gat), .dinb(G188gat), .dout(n522));
  jand g0459(.dina(n522), .dinb(n443), .dout(n523));
  jnot g0460(.din(n523), .dout(n524));
  jand g0461(.dina(n524), .dinb(n521), .dout(n525));
  jor  g0462(.dina(n525), .dinb(n446), .dout(n526));
  jnot g0463(.din(n526), .dout(n527));
  jand g0464(.dina(n524), .dinb(n446), .dout(n528));
  jor  g0465(.dina(n528), .dinb(n527), .dout(n529));
  jxor g0466(.dina(n529), .dinb(n519), .dout(n530));
  jxor g0467(.dina(n530), .dinb(n518), .dout(n531));
  jxor g0468(.dina(n531), .dinb(n514), .dout(n532));
  jxor g0469(.dina(n532), .dinb(n512), .dout(n533));
  jxor g0470(.dina(n533), .dinb(n509), .dout(n534));
  jxor g0471(.dina(n534), .dinb(n507), .dout(n535));
  jxor g0472(.dina(n535), .dinb(n504), .dout(n536));
  jxor g0473(.dina(n536), .dinb(n502), .dout(n537));
  jxor g0474(.dina(n537), .dinb(n499), .dout(n538));
  jxor g0475(.dina(n538), .dinb(n497), .dout(n539));
  jxor g0476(.dina(n539), .dinb(n494), .dout(n540));
  jxor g0477(.dina(n540), .dinb(n492), .dout(n541));
  jxor g0478(.dina(n541), .dinb(n489), .dout(n542));
  jxor g0479(.dina(n542), .dinb(n487), .dout(n543));
  jxor g0480(.dina(n543), .dinb(n484), .dout(n544));
  jnot g0481(.din(n544), .dout(n545));
  jxor g0482(.dina(n545), .dinb(n482), .dout(n546));
  jxor g0483(.dina(n546), .dinb(n478), .dout(n547));
  jxor g0484(.dina(n547), .dinb(n476), .dout(n548));
  jxor g0485(.dina(n548), .dinb(n472), .dout(G4946gat));
  jand g0486(.dina(G477gat), .dinb(G1gat), .dout(n550));
  jnot g0487(.din(n550), .dout(n551));
  jnot g0488(.din(n547), .dout(n552));
  jor  g0489(.dina(n552), .dinb(n476), .dout(n553));
  jor  g0490(.dina(n548), .dinb(n471), .dout(n554));
  jand g0491(.dina(n554), .dinb(n553), .dout(n555));
  jand g0492(.dina(G460gat), .dinb(G18gat), .dout(n556));
  jnot g0493(.din(n556), .dout(n557));
  jor  g0494(.dina(n545), .dinb(n482), .dout(n558));
  jxor g0495(.dina(n544), .dinb(n482), .dout(n559));
  jor  g0496(.dina(n559), .dinb(n477), .dout(n560));
  jand g0497(.dina(n560), .dinb(n558), .dout(n561));
  jand g0498(.dina(G443gat), .dinb(G35gat), .dout(n562));
  jnot g0499(.din(n562), .dout(n563));
  jand g0500(.dina(n542), .dinb(n487), .dout(n564));
  jand g0501(.dina(n543), .dinb(n484), .dout(n565));
  jor  g0502(.dina(n565), .dinb(n564), .dout(n566));
  jand g0503(.dina(G426gat), .dinb(G52gat), .dout(n567));
  jnot g0504(.din(n567), .dout(n568));
  jand g0505(.dina(n540), .dinb(n492), .dout(n569));
  jand g0506(.dina(n541), .dinb(n489), .dout(n570));
  jor  g0507(.dina(n570), .dinb(n569), .dout(n571));
  jand g0508(.dina(G409gat), .dinb(G69gat), .dout(n572));
  jnot g0509(.din(n572), .dout(n573));
  jand g0510(.dina(n538), .dinb(n497), .dout(n574));
  jand g0511(.dina(n539), .dinb(n494), .dout(n575));
  jor  g0512(.dina(n575), .dinb(n574), .dout(n576));
  jand g0513(.dina(G392gat), .dinb(G86gat), .dout(n577));
  jnot g0514(.din(n577), .dout(n578));
  jand g0515(.dina(n536), .dinb(n502), .dout(n579));
  jand g0516(.dina(n537), .dinb(n499), .dout(n580));
  jor  g0517(.dina(n580), .dinb(n579), .dout(n581));
  jand g0518(.dina(G375gat), .dinb(G103gat), .dout(n582));
  jnot g0519(.din(n582), .dout(n583));
  jand g0520(.dina(n534), .dinb(n507), .dout(n584));
  jand g0521(.dina(n535), .dinb(n504), .dout(n585));
  jor  g0522(.dina(n585), .dinb(n584), .dout(n586));
  jand g0523(.dina(G358gat), .dinb(G120gat), .dout(n587));
  jnot g0524(.din(n587), .dout(n588));
  jand g0525(.dina(n532), .dinb(n512), .dout(n589));
  jand g0526(.dina(n533), .dinb(n509), .dout(n590));
  jor  g0527(.dina(n590), .dinb(n589), .dout(n591));
  jand g0528(.dina(G341gat), .dinb(G137gat), .dout(n592));
  jnot g0529(.din(n592), .dout(n593));
  jand g0530(.dina(n530), .dinb(n518), .dout(n594));
  jand g0531(.dina(n531), .dinb(n514), .dout(n595));
  jor  g0532(.dina(n595), .dinb(n594), .dout(n596));
  jand g0533(.dina(G324gat), .dinb(G154gat), .dout(n597));
  jnot g0534(.din(n597), .dout(n598));
  jnot g0535(.din(n519), .dout(n599));
  jnot g0536(.din(n529), .dout(n600));
  jand g0537(.dina(n600), .dinb(n599), .dout(n601));
  jor  g0538(.dina(n601), .dinb(n527), .dout(n602));
  jand g0539(.dina(G307gat), .dinb(G171gat), .dout(n603));
  jand g0540(.dina(G273gat), .dinb(G205gat), .dout(n604));
  jor  g0541(.dina(n604), .dinb(n522), .dout(n605));
  jand g0542(.dina(G290gat), .dinb(G205gat), .dout(n606));
  jand g0543(.dina(n606), .dinb(n520), .dout(n607));
  jnot g0544(.din(n607), .dout(n608));
  jand g0545(.dina(n608), .dinb(n605), .dout(n609));
  jor  g0546(.dina(n609), .dinb(n523), .dout(n610));
  jnot g0547(.din(n610), .dout(n611));
  jand g0548(.dina(n608), .dinb(n523), .dout(n612));
  jor  g0549(.dina(n612), .dinb(n611), .dout(n613));
  jxor g0550(.dina(n613), .dinb(n603), .dout(n614));
  jxor g0551(.dina(n614), .dinb(n602), .dout(n615));
  jxor g0552(.dina(n615), .dinb(n598), .dout(n616));
  jxor g0553(.dina(n616), .dinb(n596), .dout(n617));
  jxor g0554(.dina(n617), .dinb(n593), .dout(n618));
  jxor g0555(.dina(n618), .dinb(n591), .dout(n619));
  jxor g0556(.dina(n619), .dinb(n588), .dout(n620));
  jxor g0557(.dina(n620), .dinb(n586), .dout(n621));
  jxor g0558(.dina(n621), .dinb(n583), .dout(n622));
  jxor g0559(.dina(n622), .dinb(n581), .dout(n623));
  jxor g0560(.dina(n623), .dinb(n578), .dout(n624));
  jxor g0561(.dina(n624), .dinb(n576), .dout(n625));
  jxor g0562(.dina(n625), .dinb(n573), .dout(n626));
  jxor g0563(.dina(n626), .dinb(n571), .dout(n627));
  jxor g0564(.dina(n627), .dinb(n568), .dout(n628));
  jxor g0565(.dina(n628), .dinb(n566), .dout(n629));
  jxor g0566(.dina(n629), .dinb(n563), .dout(n630));
  jnot g0567(.din(n630), .dout(n631));
  jxor g0568(.dina(n631), .dinb(n561), .dout(n632));
  jxor g0569(.dina(n632), .dinb(n557), .dout(n633));
  jxor g0570(.dina(n633), .dinb(n555), .dout(n634));
  jxor g0571(.dina(n634), .dinb(n551), .dout(G5308gat));
  jand g0572(.dina(G494gat), .dinb(G1gat), .dout(n636));
  jnot g0573(.din(n636), .dout(n637));
  jnot g0574(.din(n633), .dout(n638));
  jor  g0575(.dina(n638), .dinb(n555), .dout(n639));
  jor  g0576(.dina(n634), .dinb(n550), .dout(n640));
  jand g0577(.dina(n640), .dinb(n639), .dout(n641));
  jand g0578(.dina(G477gat), .dinb(G18gat), .dout(n642));
  jnot g0579(.din(n642), .dout(n643));
  jor  g0580(.dina(n631), .dinb(n561), .dout(n644));
  jxor g0581(.dina(n630), .dinb(n561), .dout(n645));
  jor  g0582(.dina(n645), .dinb(n556), .dout(n646));
  jand g0583(.dina(n646), .dinb(n644), .dout(n647));
  jand g0584(.dina(G460gat), .dinb(G35gat), .dout(n648));
  jnot g0585(.din(n648), .dout(n649));
  jand g0586(.dina(n628), .dinb(n566), .dout(n650));
  jand g0587(.dina(n629), .dinb(n563), .dout(n651));
  jor  g0588(.dina(n651), .dinb(n650), .dout(n652));
  jand g0589(.dina(G443gat), .dinb(G52gat), .dout(n653));
  jnot g0590(.din(n653), .dout(n654));
  jand g0591(.dina(n626), .dinb(n571), .dout(n655));
  jand g0592(.dina(n627), .dinb(n568), .dout(n656));
  jor  g0593(.dina(n656), .dinb(n655), .dout(n657));
  jand g0594(.dina(G426gat), .dinb(G69gat), .dout(n658));
  jnot g0595(.din(n658), .dout(n659));
  jand g0596(.dina(n624), .dinb(n576), .dout(n660));
  jand g0597(.dina(n625), .dinb(n573), .dout(n661));
  jor  g0598(.dina(n661), .dinb(n660), .dout(n662));
  jand g0599(.dina(G409gat), .dinb(G86gat), .dout(n663));
  jnot g0600(.din(n663), .dout(n664));
  jand g0601(.dina(n622), .dinb(n581), .dout(n665));
  jand g0602(.dina(n623), .dinb(n578), .dout(n666));
  jor  g0603(.dina(n666), .dinb(n665), .dout(n667));
  jand g0604(.dina(G392gat), .dinb(G103gat), .dout(n668));
  jnot g0605(.din(n668), .dout(n669));
  jand g0606(.dina(n620), .dinb(n586), .dout(n670));
  jand g0607(.dina(n621), .dinb(n583), .dout(n671));
  jor  g0608(.dina(n671), .dinb(n670), .dout(n672));
  jand g0609(.dina(G375gat), .dinb(G120gat), .dout(n673));
  jnot g0610(.din(n673), .dout(n674));
  jand g0611(.dina(n618), .dinb(n591), .dout(n675));
  jand g0612(.dina(n619), .dinb(n588), .dout(n676));
  jor  g0613(.dina(n676), .dinb(n675), .dout(n677));
  jand g0614(.dina(G358gat), .dinb(G137gat), .dout(n678));
  jnot g0615(.din(n678), .dout(n679));
  jand g0616(.dina(n616), .dinb(n596), .dout(n680));
  jand g0617(.dina(n617), .dinb(n593), .dout(n681));
  jor  g0618(.dina(n681), .dinb(n680), .dout(n682));
  jand g0619(.dina(G341gat), .dinb(G154gat), .dout(n683));
  jnot g0620(.din(n683), .dout(n684));
  jand g0621(.dina(n614), .dinb(n602), .dout(n685));
  jand g0622(.dina(n615), .dinb(n598), .dout(n686));
  jor  g0623(.dina(n686), .dinb(n685), .dout(n687));
  jand g0624(.dina(G324gat), .dinb(G171gat), .dout(n688));
  jnot g0625(.din(n688), .dout(n689));
  jnot g0626(.din(n603), .dout(n690));
  jnot g0627(.din(n613), .dout(n691));
  jand g0628(.dina(n691), .dinb(n690), .dout(n692));
  jor  g0629(.dina(n692), .dinb(n611), .dout(n693));
  jand g0630(.dina(G307gat), .dinb(G188gat), .dout(n694));
  jand g0631(.dina(G273gat), .dinb(G222gat), .dout(n695));
  jor  g0632(.dina(n695), .dinb(n606), .dout(n696));
  jand g0633(.dina(G290gat), .dinb(G222gat), .dout(n697));
  jand g0634(.dina(n697), .dinb(n604), .dout(n698));
  jnot g0635(.din(n698), .dout(n699));
  jand g0636(.dina(n699), .dinb(n696), .dout(n700));
  jor  g0637(.dina(n700), .dinb(n607), .dout(n701));
  jnot g0638(.din(n701), .dout(n702));
  jand g0639(.dina(n699), .dinb(n607), .dout(n703));
  jor  g0640(.dina(n703), .dinb(n702), .dout(n704));
  jxor g0641(.dina(n704), .dinb(n694), .dout(n705));
  jxor g0642(.dina(n705), .dinb(n693), .dout(n706));
  jxor g0643(.dina(n706), .dinb(n689), .dout(n707));
  jxor g0644(.dina(n707), .dinb(n687), .dout(n708));
  jxor g0645(.dina(n708), .dinb(n684), .dout(n709));
  jxor g0646(.dina(n709), .dinb(n682), .dout(n710));
  jxor g0647(.dina(n710), .dinb(n679), .dout(n711));
  jxor g0648(.dina(n711), .dinb(n677), .dout(n712));
  jxor g0649(.dina(n712), .dinb(n674), .dout(n713));
  jxor g0650(.dina(n713), .dinb(n672), .dout(n714));
  jxor g0651(.dina(n714), .dinb(n669), .dout(n715));
  jxor g0652(.dina(n715), .dinb(n667), .dout(n716));
  jxor g0653(.dina(n716), .dinb(n664), .dout(n717));
  jxor g0654(.dina(n717), .dinb(n662), .dout(n718));
  jxor g0655(.dina(n718), .dinb(n659), .dout(n719));
  jxor g0656(.dina(n719), .dinb(n657), .dout(n720));
  jxor g0657(.dina(n720), .dinb(n654), .dout(n721));
  jxor g0658(.dina(n721), .dinb(n652), .dout(n722));
  jxor g0659(.dina(n722), .dinb(n649), .dout(n723));
  jnot g0660(.din(n723), .dout(n724));
  jxor g0661(.dina(n724), .dinb(n647), .dout(n725));
  jxor g0662(.dina(n725), .dinb(n643), .dout(n726));
  jxor g0663(.dina(n726), .dinb(n641), .dout(n727));
  jxor g0664(.dina(n727), .dinb(n637), .dout(G5672gat));
  jand g0665(.dina(G511gat), .dinb(G1gat), .dout(n729));
  jnot g0666(.din(n729), .dout(n730));
  jnot g0667(.din(n726), .dout(n731));
  jor  g0668(.dina(n731), .dinb(n641), .dout(n732));
  jor  g0669(.dina(n727), .dinb(n636), .dout(n733));
  jand g0670(.dina(n733), .dinb(n732), .dout(n734));
  jand g0671(.dina(G494gat), .dinb(G18gat), .dout(n735));
  jnot g0672(.din(n735), .dout(n736));
  jor  g0673(.dina(n724), .dinb(n647), .dout(n737));
  jxor g0674(.dina(n723), .dinb(n647), .dout(n738));
  jor  g0675(.dina(n738), .dinb(n642), .dout(n739));
  jand g0676(.dina(n739), .dinb(n737), .dout(n740));
  jand g0677(.dina(G477gat), .dinb(G35gat), .dout(n741));
  jnot g0678(.din(n741), .dout(n742));
  jand g0679(.dina(n721), .dinb(n652), .dout(n743));
  jand g0680(.dina(n722), .dinb(n649), .dout(n744));
  jor  g0681(.dina(n744), .dinb(n743), .dout(n745));
  jand g0682(.dina(G460gat), .dinb(G52gat), .dout(n746));
  jnot g0683(.din(n746), .dout(n747));
  jand g0684(.dina(n719), .dinb(n657), .dout(n748));
  jand g0685(.dina(n720), .dinb(n654), .dout(n749));
  jor  g0686(.dina(n749), .dinb(n748), .dout(n750));
  jand g0687(.dina(G443gat), .dinb(G69gat), .dout(n751));
  jnot g0688(.din(n751), .dout(n752));
  jand g0689(.dina(n717), .dinb(n662), .dout(n753));
  jand g0690(.dina(n718), .dinb(n659), .dout(n754));
  jor  g0691(.dina(n754), .dinb(n753), .dout(n755));
  jand g0692(.dina(G426gat), .dinb(G86gat), .dout(n756));
  jnot g0693(.din(n756), .dout(n757));
  jand g0694(.dina(n715), .dinb(n667), .dout(n758));
  jand g0695(.dina(n716), .dinb(n664), .dout(n759));
  jor  g0696(.dina(n759), .dinb(n758), .dout(n760));
  jand g0697(.dina(G409gat), .dinb(G103gat), .dout(n761));
  jnot g0698(.din(n761), .dout(n762));
  jand g0699(.dina(n713), .dinb(n672), .dout(n763));
  jand g0700(.dina(n714), .dinb(n669), .dout(n764));
  jor  g0701(.dina(n764), .dinb(n763), .dout(n765));
  jand g0702(.dina(G392gat), .dinb(G120gat), .dout(n766));
  jnot g0703(.din(n766), .dout(n767));
  jand g0704(.dina(n711), .dinb(n677), .dout(n768));
  jand g0705(.dina(n712), .dinb(n674), .dout(n769));
  jor  g0706(.dina(n769), .dinb(n768), .dout(n770));
  jand g0707(.dina(G375gat), .dinb(G137gat), .dout(n771));
  jnot g0708(.din(n771), .dout(n772));
  jand g0709(.dina(n709), .dinb(n682), .dout(n773));
  jand g0710(.dina(n710), .dinb(n679), .dout(n774));
  jor  g0711(.dina(n774), .dinb(n773), .dout(n775));
  jand g0712(.dina(G358gat), .dinb(G154gat), .dout(n776));
  jnot g0713(.din(n776), .dout(n777));
  jand g0714(.dina(n707), .dinb(n687), .dout(n778));
  jand g0715(.dina(n708), .dinb(n684), .dout(n779));
  jor  g0716(.dina(n779), .dinb(n778), .dout(n780));
  jand g0717(.dina(G341gat), .dinb(G171gat), .dout(n781));
  jnot g0718(.din(n781), .dout(n782));
  jand g0719(.dina(n705), .dinb(n693), .dout(n783));
  jand g0720(.dina(n706), .dinb(n689), .dout(n784));
  jor  g0721(.dina(n784), .dinb(n783), .dout(n785));
  jand g0722(.dina(G324gat), .dinb(G188gat), .dout(n786));
  jnot g0723(.din(n786), .dout(n787));
  jnot g0724(.din(n694), .dout(n788));
  jnot g0725(.din(n704), .dout(n789));
  jand g0726(.dina(n789), .dinb(n788), .dout(n790));
  jor  g0727(.dina(n790), .dinb(n702), .dout(n791));
  jand g0728(.dina(G307gat), .dinb(G205gat), .dout(n792));
  jand g0729(.dina(G273gat), .dinb(G239gat), .dout(n793));
  jor  g0730(.dina(n793), .dinb(n697), .dout(n794));
  jand g0731(.dina(G290gat), .dinb(G239gat), .dout(n795));
  jand g0732(.dina(n795), .dinb(n695), .dout(n796));
  jnot g0733(.din(n796), .dout(n797));
  jand g0734(.dina(n797), .dinb(n794), .dout(n798));
  jor  g0735(.dina(n798), .dinb(n698), .dout(n799));
  jnot g0736(.din(n799), .dout(n800));
  jand g0737(.dina(n797), .dinb(n698), .dout(n801));
  jor  g0738(.dina(n801), .dinb(n800), .dout(n802));
  jxor g0739(.dina(n802), .dinb(n792), .dout(n803));
  jxor g0740(.dina(n803), .dinb(n791), .dout(n804));
  jxor g0741(.dina(n804), .dinb(n787), .dout(n805));
  jxor g0742(.dina(n805), .dinb(n785), .dout(n806));
  jxor g0743(.dina(n806), .dinb(n782), .dout(n807));
  jxor g0744(.dina(n807), .dinb(n780), .dout(n808));
  jxor g0745(.dina(n808), .dinb(n777), .dout(n809));
  jxor g0746(.dina(n809), .dinb(n775), .dout(n810));
  jxor g0747(.dina(n810), .dinb(n772), .dout(n811));
  jxor g0748(.dina(n811), .dinb(n770), .dout(n812));
  jxor g0749(.dina(n812), .dinb(n767), .dout(n813));
  jxor g0750(.dina(n813), .dinb(n765), .dout(n814));
  jxor g0751(.dina(n814), .dinb(n762), .dout(n815));
  jxor g0752(.dina(n815), .dinb(n760), .dout(n816));
  jxor g0753(.dina(n816), .dinb(n757), .dout(n817));
  jxor g0754(.dina(n817), .dinb(n755), .dout(n818));
  jxor g0755(.dina(n818), .dinb(n752), .dout(n819));
  jxor g0756(.dina(n819), .dinb(n750), .dout(n820));
  jxor g0757(.dina(n820), .dinb(n747), .dout(n821));
  jxor g0758(.dina(n821), .dinb(n745), .dout(n822));
  jxor g0759(.dina(n822), .dinb(n742), .dout(n823));
  jnot g0760(.din(n823), .dout(n824));
  jxor g0761(.dina(n824), .dinb(n740), .dout(n825));
  jxor g0762(.dina(n825), .dinb(n736), .dout(n826));
  jxor g0763(.dina(n826), .dinb(n734), .dout(n827));
  jxor g0764(.dina(n827), .dinb(n730), .dout(G5971gat));
  jand g0765(.dina(G528gat), .dinb(G1gat), .dout(n829));
  jnot g0766(.din(n829), .dout(n830));
  jnot g0767(.din(n826), .dout(n831));
  jor  g0768(.dina(n831), .dinb(n734), .dout(n832));
  jor  g0769(.dina(n827), .dinb(n729), .dout(n833));
  jand g0770(.dina(n833), .dinb(n832), .dout(n834));
  jand g0771(.dina(G511gat), .dinb(G18gat), .dout(n835));
  jor  g0772(.dina(n824), .dinb(n740), .dout(n836));
  jxor g0773(.dina(n823), .dinb(n740), .dout(n837));
  jor  g0774(.dina(n837), .dinb(n735), .dout(n838));
  jand g0775(.dina(n838), .dinb(n836), .dout(n839));
  jand g0776(.dina(G494gat), .dinb(G35gat), .dout(n840));
  jnot g0777(.din(n840), .dout(n841));
  jand g0778(.dina(n821), .dinb(n745), .dout(n842));
  jand g0779(.dina(n822), .dinb(n742), .dout(n843));
  jor  g0780(.dina(n843), .dinb(n842), .dout(n844));
  jand g0781(.dina(G477gat), .dinb(G52gat), .dout(n845));
  jnot g0782(.din(n845), .dout(n846));
  jand g0783(.dina(n819), .dinb(n750), .dout(n847));
  jand g0784(.dina(n820), .dinb(n747), .dout(n848));
  jor  g0785(.dina(n848), .dinb(n847), .dout(n849));
  jand g0786(.dina(G460gat), .dinb(G69gat), .dout(n850));
  jnot g0787(.din(n850), .dout(n851));
  jand g0788(.dina(n817), .dinb(n755), .dout(n852));
  jand g0789(.dina(n818), .dinb(n752), .dout(n853));
  jor  g0790(.dina(n853), .dinb(n852), .dout(n854));
  jand g0791(.dina(G443gat), .dinb(G86gat), .dout(n855));
  jnot g0792(.din(n855), .dout(n856));
  jand g0793(.dina(n815), .dinb(n760), .dout(n857));
  jand g0794(.dina(n816), .dinb(n757), .dout(n858));
  jor  g0795(.dina(n858), .dinb(n857), .dout(n859));
  jand g0796(.dina(G426gat), .dinb(G103gat), .dout(n860));
  jnot g0797(.din(n860), .dout(n861));
  jand g0798(.dina(n813), .dinb(n765), .dout(n862));
  jand g0799(.dina(n814), .dinb(n762), .dout(n863));
  jor  g0800(.dina(n863), .dinb(n862), .dout(n864));
  jand g0801(.dina(G409gat), .dinb(G120gat), .dout(n865));
  jnot g0802(.din(n865), .dout(n866));
  jand g0803(.dina(n811), .dinb(n770), .dout(n867));
  jand g0804(.dina(n812), .dinb(n767), .dout(n868));
  jor  g0805(.dina(n868), .dinb(n867), .dout(n869));
  jand g0806(.dina(G392gat), .dinb(G137gat), .dout(n870));
  jnot g0807(.din(n870), .dout(n871));
  jand g0808(.dina(n809), .dinb(n775), .dout(n872));
  jand g0809(.dina(n810), .dinb(n772), .dout(n873));
  jor  g0810(.dina(n873), .dinb(n872), .dout(n874));
  jand g0811(.dina(G375gat), .dinb(G154gat), .dout(n875));
  jnot g0812(.din(n875), .dout(n876));
  jand g0813(.dina(n807), .dinb(n780), .dout(n877));
  jand g0814(.dina(n808), .dinb(n777), .dout(n878));
  jor  g0815(.dina(n878), .dinb(n877), .dout(n879));
  jand g0816(.dina(G358gat), .dinb(G171gat), .dout(n880));
  jnot g0817(.din(n880), .dout(n881));
  jand g0818(.dina(n805), .dinb(n785), .dout(n882));
  jand g0819(.dina(n806), .dinb(n782), .dout(n883));
  jor  g0820(.dina(n883), .dinb(n882), .dout(n884));
  jand g0821(.dina(G341gat), .dinb(G188gat), .dout(n885));
  jnot g0822(.din(n885), .dout(n886));
  jand g0823(.dina(n803), .dinb(n791), .dout(n887));
  jand g0824(.dina(n804), .dinb(n787), .dout(n888));
  jor  g0825(.dina(n888), .dinb(n887), .dout(n889));
  jand g0826(.dina(G324gat), .dinb(G205gat), .dout(n890));
  jnot g0827(.din(n890), .dout(n891));
  jnot g0828(.din(n792), .dout(n892));
  jnot g0829(.din(n802), .dout(n893));
  jand g0830(.dina(n893), .dinb(n892), .dout(n894));
  jor  g0831(.dina(n894), .dinb(n800), .dout(n895));
  jand g0832(.dina(G307gat), .dinb(G222gat), .dout(n896));
  jnot g0833(.din(n795), .dout(n897));
  jand g0834(.dina(G273gat), .dinb(G256gat), .dout(n898));
  jand g0835(.dina(n898), .dinb(n897), .dout(n899));
  jnot g0836(.din(n899), .dout(n900));
  jor  g0837(.dina(n898), .dinb(n897), .dout(n901));
  jand g0838(.dina(n901), .dinb(n797), .dout(n902));
  jand g0839(.dina(n902), .dinb(n900), .dout(n903));
  jnot g0840(.din(n901), .dout(n904));
  jand g0841(.dina(n904), .dinb(n695), .dout(n905));
  jor  g0842(.dina(n905), .dinb(n903), .dout(n906));
  jxor g0843(.dina(n906), .dinb(n896), .dout(n907));
  jxor g0844(.dina(n907), .dinb(n895), .dout(n908));
  jxor g0845(.dina(n908), .dinb(n891), .dout(n909));
  jxor g0846(.dina(n909), .dinb(n889), .dout(n910));
  jxor g0847(.dina(n910), .dinb(n886), .dout(n911));
  jxor g0848(.dina(n911), .dinb(n884), .dout(n912));
  jxor g0849(.dina(n912), .dinb(n881), .dout(n913));
  jxor g0850(.dina(n913), .dinb(n879), .dout(n914));
  jxor g0851(.dina(n914), .dinb(n876), .dout(n915));
  jxor g0852(.dina(n915), .dinb(n874), .dout(n916));
  jxor g0853(.dina(n916), .dinb(n871), .dout(n917));
  jxor g0854(.dina(n917), .dinb(n869), .dout(n918));
  jxor g0855(.dina(n918), .dinb(n866), .dout(n919));
  jxor g0856(.dina(n919), .dinb(n864), .dout(n920));
  jxor g0857(.dina(n920), .dinb(n861), .dout(n921));
  jxor g0858(.dina(n921), .dinb(n859), .dout(n922));
  jxor g0859(.dina(n922), .dinb(n856), .dout(n923));
  jxor g0860(.dina(n923), .dinb(n854), .dout(n924));
  jxor g0861(.dina(n924), .dinb(n851), .dout(n925));
  jxor g0862(.dina(n925), .dinb(n849), .dout(n926));
  jxor g0863(.dina(n926), .dinb(n846), .dout(n927));
  jxor g0864(.dina(n927), .dinb(n844), .dout(n928));
  jxor g0865(.dina(n928), .dinb(n841), .dout(n929));
  jxor g0866(.dina(n929), .dinb(n839), .dout(n930));
  jxor g0867(.dina(n930), .dinb(n835), .dout(n931));
  jxor g0868(.dina(n931), .dinb(n834), .dout(n932));
  jxor g0869(.dina(n932), .dinb(n830), .dout(G6123gat));
  jnot g0870(.din(n931), .dout(n934));
  jor  g0871(.dina(n934), .dinb(n834), .dout(n935));
  jor  g0872(.dina(n932), .dinb(n829), .dout(n936));
  jand g0873(.dina(n936), .dinb(n935), .dout(n937));
  jand g0874(.dina(G528gat), .dinb(G18gat), .dout(n938));
  jnot g0875(.din(n929), .dout(n939));
  jor  g0876(.dina(n939), .dinb(n839), .dout(n940));
  jor  g0877(.dina(n930), .dinb(n835), .dout(n941));
  jand g0878(.dina(n941), .dinb(n940), .dout(n942));
  jand g0879(.dina(G511gat), .dinb(G35gat), .dout(n943));
  jand g0880(.dina(n927), .dinb(n844), .dout(n944));
  jnot g0881(.din(n944), .dout(n945));
  jnot g0882(.din(n927), .dout(n946));
  jxor g0883(.dina(n946), .dinb(n844), .dout(n947));
  jor  g0884(.dina(n947), .dinb(n840), .dout(n948));
  jand g0885(.dina(n948), .dinb(n945), .dout(n949));
  jand g0886(.dina(G494gat), .dinb(G52gat), .dout(n950));
  jnot g0887(.din(n950), .dout(n951));
  jand g0888(.dina(n925), .dinb(n849), .dout(n952));
  jand g0889(.dina(n926), .dinb(n846), .dout(n953));
  jor  g0890(.dina(n953), .dinb(n952), .dout(n954));
  jand g0891(.dina(G477gat), .dinb(G69gat), .dout(n955));
  jnot g0892(.din(n955), .dout(n956));
  jand g0893(.dina(n923), .dinb(n854), .dout(n957));
  jand g0894(.dina(n924), .dinb(n851), .dout(n958));
  jor  g0895(.dina(n958), .dinb(n957), .dout(n959));
  jand g0896(.dina(G460gat), .dinb(G86gat), .dout(n960));
  jnot g0897(.din(n960), .dout(n961));
  jand g0898(.dina(n921), .dinb(n859), .dout(n962));
  jand g0899(.dina(n922), .dinb(n856), .dout(n963));
  jor  g0900(.dina(n963), .dinb(n962), .dout(n964));
  jand g0901(.dina(G443gat), .dinb(G103gat), .dout(n965));
  jnot g0902(.din(n965), .dout(n966));
  jand g0903(.dina(n919), .dinb(n864), .dout(n967));
  jand g0904(.dina(n920), .dinb(n861), .dout(n968));
  jor  g0905(.dina(n968), .dinb(n967), .dout(n969));
  jand g0906(.dina(G426gat), .dinb(G120gat), .dout(n970));
  jnot g0907(.din(n970), .dout(n971));
  jand g0908(.dina(n917), .dinb(n869), .dout(n972));
  jand g0909(.dina(n918), .dinb(n866), .dout(n973));
  jor  g0910(.dina(n973), .dinb(n972), .dout(n974));
  jand g0911(.dina(G409gat), .dinb(G137gat), .dout(n975));
  jnot g0912(.din(n975), .dout(n976));
  jand g0913(.dina(n915), .dinb(n874), .dout(n977));
  jand g0914(.dina(n916), .dinb(n871), .dout(n978));
  jor  g0915(.dina(n978), .dinb(n977), .dout(n979));
  jand g0916(.dina(G392gat), .dinb(G154gat), .dout(n980));
  jnot g0917(.din(n980), .dout(n981));
  jand g0918(.dina(n913), .dinb(n879), .dout(n982));
  jand g0919(.dina(n914), .dinb(n876), .dout(n983));
  jor  g0920(.dina(n983), .dinb(n982), .dout(n984));
  jand g0921(.dina(G375gat), .dinb(G171gat), .dout(n985));
  jnot g0922(.din(n985), .dout(n986));
  jand g0923(.dina(n911), .dinb(n884), .dout(n987));
  jand g0924(.dina(n912), .dinb(n881), .dout(n988));
  jor  g0925(.dina(n988), .dinb(n987), .dout(n989));
  jand g0926(.dina(G358gat), .dinb(G188gat), .dout(n990));
  jnot g0927(.din(n990), .dout(n991));
  jand g0928(.dina(n909), .dinb(n889), .dout(n992));
  jand g0929(.dina(n910), .dinb(n886), .dout(n993));
  jor  g0930(.dina(n993), .dinb(n992), .dout(n994));
  jand g0931(.dina(G341gat), .dinb(G205gat), .dout(n995));
  jnot g0932(.din(n995), .dout(n996));
  jand g0933(.dina(n907), .dinb(n895), .dout(n997));
  jand g0934(.dina(n908), .dinb(n891), .dout(n998));
  jor  g0935(.dina(n998), .dinb(n997), .dout(n999));
  jand g0936(.dina(G324gat), .dinb(G222gat), .dout(n1000));
  jnot g0937(.din(n1000), .dout(n1001));
  jnot g0938(.din(n896), .dout(n1002));
  jnot g0939(.din(n906), .dout(n1003));
  jand g0940(.dina(n1003), .dinb(n1002), .dout(n1004));
  jor  g0941(.dina(n1004), .dinb(n903), .dout(n1005));
  jand g0942(.dina(G307gat), .dinb(G239gat), .dout(n1006));
  jand g0943(.dina(G290gat), .dinb(G256gat), .dout(n1007));
  jnot g0944(.din(n1007), .dout(n1008));
  jor  g0945(.dina(n1008), .dinb(n793), .dout(n1009));
  jxor g0946(.dina(n1009), .dinb(n1006), .dout(n1010));
  jxor g0947(.dina(n1010), .dinb(n1005), .dout(n1011));
  jxor g0948(.dina(n1011), .dinb(n1001), .dout(n1012));
  jxor g0949(.dina(n1012), .dinb(n999), .dout(n1013));
  jxor g0950(.dina(n1013), .dinb(n996), .dout(n1014));
  jxor g0951(.dina(n1014), .dinb(n994), .dout(n1015));
  jxor g0952(.dina(n1015), .dinb(n991), .dout(n1016));
  jxor g0953(.dina(n1016), .dinb(n989), .dout(n1017));
  jxor g0954(.dina(n1017), .dinb(n986), .dout(n1018));
  jxor g0955(.dina(n1018), .dinb(n984), .dout(n1019));
  jxor g0956(.dina(n1019), .dinb(n981), .dout(n1020));
  jxor g0957(.dina(n1020), .dinb(n979), .dout(n1021));
  jxor g0958(.dina(n1021), .dinb(n976), .dout(n1022));
  jxor g0959(.dina(n1022), .dinb(n974), .dout(n1023));
  jxor g0960(.dina(n1023), .dinb(n971), .dout(n1024));
  jxor g0961(.dina(n1024), .dinb(n969), .dout(n1025));
  jxor g0962(.dina(n1025), .dinb(n966), .dout(n1026));
  jxor g0963(.dina(n1026), .dinb(n964), .dout(n1027));
  jxor g0964(.dina(n1027), .dinb(n961), .dout(n1028));
  jxor g0965(.dina(n1028), .dinb(n959), .dout(n1029));
  jxor g0966(.dina(n1029), .dinb(n956), .dout(n1030));
  jxor g0967(.dina(n1030), .dinb(n954), .dout(n1031));
  jxor g0968(.dina(n1031), .dinb(n951), .dout(n1032));
  jxor g0969(.dina(n1032), .dinb(n949), .dout(n1033));
  jxor g0970(.dina(n1033), .dinb(n943), .dout(n1034));
  jnot g0971(.din(n1034), .dout(n1035));
  jxor g0972(.dina(n1035), .dinb(n942), .dout(n1036));
  jxor g0973(.dina(n1036), .dinb(n938), .dout(n1037));
  jxor g0974(.dina(n1037), .dinb(n937), .dout(G6150gat));
  jand g0975(.dina(n1037), .dinb(n937), .dout(n1039));
  jor  g0976(.dina(n1035), .dinb(n942), .dout(n1040));
  jxor g0977(.dina(n1034), .dinb(n942), .dout(n1041));
  jor  g0978(.dina(n1041), .dinb(n938), .dout(n1042));
  jand g0979(.dina(n1042), .dinb(n1040), .dout(n1043));
  jand g0980(.dina(G528gat), .dinb(G35gat), .dout(n1044));
  jnot g0981(.din(n1032), .dout(n1045));
  jor  g0982(.dina(n1045), .dinb(n949), .dout(n1046));
  jor  g0983(.dina(n1033), .dinb(n943), .dout(n1047));
  jand g0984(.dina(n1047), .dinb(n1046), .dout(n1048));
  jand g0985(.dina(G511gat), .dinb(G52gat), .dout(n1049));
  jand g0986(.dina(n1030), .dinb(n954), .dout(n1050));
  jand g0987(.dina(n1031), .dinb(n951), .dout(n1051));
  jor  g0988(.dina(n1051), .dinb(n1050), .dout(n1052));
  jand g0989(.dina(G494gat), .dinb(G69gat), .dout(n1053));
  jnot g0990(.din(n1053), .dout(n1054));
  jand g0991(.dina(n1028), .dinb(n959), .dout(n1055));
  jand g0992(.dina(n1029), .dinb(n956), .dout(n1056));
  jor  g0993(.dina(n1056), .dinb(n1055), .dout(n1057));
  jand g0994(.dina(G477gat), .dinb(G86gat), .dout(n1058));
  jnot g0995(.din(n1058), .dout(n1059));
  jand g0996(.dina(n1026), .dinb(n964), .dout(n1060));
  jand g0997(.dina(n1027), .dinb(n961), .dout(n1061));
  jor  g0998(.dina(n1061), .dinb(n1060), .dout(n1062));
  jand g0999(.dina(G460gat), .dinb(G103gat), .dout(n1063));
  jnot g1000(.din(n1063), .dout(n1064));
  jand g1001(.dina(n1024), .dinb(n969), .dout(n1065));
  jand g1002(.dina(n1025), .dinb(n966), .dout(n1066));
  jor  g1003(.dina(n1066), .dinb(n1065), .dout(n1067));
  jand g1004(.dina(G443gat), .dinb(G120gat), .dout(n1068));
  jnot g1005(.din(n1068), .dout(n1069));
  jand g1006(.dina(n1022), .dinb(n974), .dout(n1070));
  jand g1007(.dina(n1023), .dinb(n971), .dout(n1071));
  jor  g1008(.dina(n1071), .dinb(n1070), .dout(n1072));
  jand g1009(.dina(G426gat), .dinb(G137gat), .dout(n1073));
  jnot g1010(.din(n1073), .dout(n1074));
  jand g1011(.dina(n1020), .dinb(n979), .dout(n1075));
  jand g1012(.dina(n1021), .dinb(n976), .dout(n1076));
  jor  g1013(.dina(n1076), .dinb(n1075), .dout(n1077));
  jand g1014(.dina(G409gat), .dinb(G154gat), .dout(n1078));
  jnot g1015(.din(n1078), .dout(n1079));
  jand g1016(.dina(n1018), .dinb(n984), .dout(n1080));
  jand g1017(.dina(n1019), .dinb(n981), .dout(n1081));
  jor  g1018(.dina(n1081), .dinb(n1080), .dout(n1082));
  jand g1019(.dina(G392gat), .dinb(G171gat), .dout(n1083));
  jnot g1020(.din(n1083), .dout(n1084));
  jand g1021(.dina(n1016), .dinb(n989), .dout(n1085));
  jand g1022(.dina(n1017), .dinb(n986), .dout(n1086));
  jor  g1023(.dina(n1086), .dinb(n1085), .dout(n1087));
  jand g1024(.dina(G375gat), .dinb(G188gat), .dout(n1088));
  jnot g1025(.din(n1088), .dout(n1089));
  jand g1026(.dina(n1014), .dinb(n994), .dout(n1090));
  jand g1027(.dina(n1015), .dinb(n991), .dout(n1091));
  jor  g1028(.dina(n1091), .dinb(n1090), .dout(n1092));
  jand g1029(.dina(G358gat), .dinb(G205gat), .dout(n1093));
  jnot g1030(.din(n1093), .dout(n1094));
  jand g1031(.dina(n1012), .dinb(n999), .dout(n1095));
  jand g1032(.dina(n1013), .dinb(n996), .dout(n1096));
  jor  g1033(.dina(n1096), .dinb(n1095), .dout(n1097));
  jand g1034(.dina(G341gat), .dinb(G222gat), .dout(n1098));
  jnot g1035(.din(n1098), .dout(n1099));
  jand g1036(.dina(n1010), .dinb(n1005), .dout(n1100));
  jand g1037(.dina(n1011), .dinb(n1001), .dout(n1101));
  jor  g1038(.dina(n1101), .dinb(n1100), .dout(n1102));
  jand g1039(.dina(G324gat), .dinb(G239gat), .dout(n1103));
  jand g1040(.dina(G307gat), .dinb(G256gat), .dout(n1104));
  jnot g1041(.din(n1006), .dout(n1105));
  jnot g1042(.din(n1009), .dout(n1106));
  jand g1043(.dina(n1106), .dinb(n1105), .dout(n1107));
  jor  g1044(.dina(n1107), .dinb(n1008), .dout(n1108));
  jnot g1045(.din(n1108), .dout(n1109));
  jor  g1046(.dina(n1109), .dinb(n1104), .dout(n1110));
  jand g1047(.dina(n1109), .dinb(G307gat), .dout(n1111));
  jnot g1048(.din(n1111), .dout(n1112));
  jand g1049(.dina(n1112), .dinb(n1110), .dout(n1113));
  jnot g1050(.din(n1113), .dout(n1114));
  jxor g1051(.dina(n1114), .dinb(n1103), .dout(n1115));
  jxor g1052(.dina(n1115), .dinb(n1102), .dout(n1116));
  jxor g1053(.dina(n1116), .dinb(n1099), .dout(n1117));
  jxor g1054(.dina(n1117), .dinb(n1097), .dout(n1118));
  jxor g1055(.dina(n1118), .dinb(n1094), .dout(n1119));
  jxor g1056(.dina(n1119), .dinb(n1092), .dout(n1120));
  jxor g1057(.dina(n1120), .dinb(n1089), .dout(n1121));
  jxor g1058(.dina(n1121), .dinb(n1087), .dout(n1122));
  jxor g1059(.dina(n1122), .dinb(n1084), .dout(n1123));
  jxor g1060(.dina(n1123), .dinb(n1082), .dout(n1124));
  jxor g1061(.dina(n1124), .dinb(n1079), .dout(n1125));
  jxor g1062(.dina(n1125), .dinb(n1077), .dout(n1126));
  jxor g1063(.dina(n1126), .dinb(n1074), .dout(n1127));
  jxor g1064(.dina(n1127), .dinb(n1072), .dout(n1128));
  jxor g1065(.dina(n1128), .dinb(n1069), .dout(n1129));
  jxor g1066(.dina(n1129), .dinb(n1067), .dout(n1130));
  jxor g1067(.dina(n1130), .dinb(n1064), .dout(n1131));
  jxor g1068(.dina(n1131), .dinb(n1062), .dout(n1132));
  jxor g1069(.dina(n1132), .dinb(n1059), .dout(n1133));
  jxor g1070(.dina(n1133), .dinb(n1057), .dout(n1134));
  jxor g1071(.dina(n1134), .dinb(n1054), .dout(n1135));
  jxor g1072(.dina(n1135), .dinb(n1052), .dout(n1136));
  jnot g1073(.din(n1136), .dout(n1137));
  jxor g1074(.dina(n1137), .dinb(n1049), .dout(n1138));
  jxor g1075(.dina(n1138), .dinb(n1048), .dout(n1139));
  jxor g1076(.dina(n1139), .dinb(n1044), .dout(n1140));
  jxor g1077(.dina(n1140), .dinb(n1043), .dout(n1141));
  jnot g1078(.din(n1141), .dout(n1142));
  jxor g1079(.dina(n1142), .dinb(n1039), .dout(G6160gat));
  jnot g1080(.din(n1140), .dout(n1144));
  jor  g1081(.dina(n1144), .dinb(n1043), .dout(n1145));
  jor  g1082(.dina(n1141), .dinb(n1039), .dout(n1146));
  jand g1083(.dina(n1146), .dinb(n1145), .dout(n1147));
  jnot g1084(.din(n1138), .dout(n1148));
  jor  g1085(.dina(n1148), .dinb(n1048), .dout(n1149));
  jor  g1086(.dina(n1139), .dinb(n1044), .dout(n1150));
  jand g1087(.dina(n1150), .dinb(n1149), .dout(n1151));
  jand g1088(.dina(G528gat), .dinb(G52gat), .dout(n1152));
  jand g1089(.dina(n1135), .dinb(n1052), .dout(n1153));
  jnot g1090(.din(n1153), .dout(n1154));
  jor  g1091(.dina(n1137), .dinb(n1049), .dout(n1155));
  jand g1092(.dina(n1155), .dinb(n1154), .dout(n1156));
  jand g1093(.dina(G511gat), .dinb(G69gat), .dout(n1157));
  jnot g1094(.din(n1157), .dout(n1158));
  jand g1095(.dina(n1133), .dinb(n1057), .dout(n1159));
  jand g1096(.dina(n1134), .dinb(n1054), .dout(n1160));
  jor  g1097(.dina(n1160), .dinb(n1159), .dout(n1161));
  jand g1098(.dina(G494gat), .dinb(G86gat), .dout(n1162));
  jnot g1099(.din(n1162), .dout(n1163));
  jand g1100(.dina(n1131), .dinb(n1062), .dout(n1164));
  jand g1101(.dina(n1132), .dinb(n1059), .dout(n1165));
  jor  g1102(.dina(n1165), .dinb(n1164), .dout(n1166));
  jand g1103(.dina(G477gat), .dinb(G103gat), .dout(n1167));
  jnot g1104(.din(n1167), .dout(n1168));
  jand g1105(.dina(n1129), .dinb(n1067), .dout(n1169));
  jand g1106(.dina(n1130), .dinb(n1064), .dout(n1170));
  jor  g1107(.dina(n1170), .dinb(n1169), .dout(n1171));
  jand g1108(.dina(G460gat), .dinb(G120gat), .dout(n1172));
  jnot g1109(.din(n1172), .dout(n1173));
  jand g1110(.dina(n1127), .dinb(n1072), .dout(n1174));
  jand g1111(.dina(n1128), .dinb(n1069), .dout(n1175));
  jor  g1112(.dina(n1175), .dinb(n1174), .dout(n1176));
  jand g1113(.dina(G443gat), .dinb(G137gat), .dout(n1177));
  jnot g1114(.din(n1177), .dout(n1178));
  jand g1115(.dina(n1125), .dinb(n1077), .dout(n1179));
  jand g1116(.dina(n1126), .dinb(n1074), .dout(n1180));
  jor  g1117(.dina(n1180), .dinb(n1179), .dout(n1181));
  jand g1118(.dina(G426gat), .dinb(G154gat), .dout(n1182));
  jnot g1119(.din(n1182), .dout(n1183));
  jand g1120(.dina(n1123), .dinb(n1082), .dout(n1184));
  jand g1121(.dina(n1124), .dinb(n1079), .dout(n1185));
  jor  g1122(.dina(n1185), .dinb(n1184), .dout(n1186));
  jand g1123(.dina(G409gat), .dinb(G171gat), .dout(n1187));
  jnot g1124(.din(n1187), .dout(n1188));
  jand g1125(.dina(n1121), .dinb(n1087), .dout(n1189));
  jand g1126(.dina(n1122), .dinb(n1084), .dout(n1190));
  jor  g1127(.dina(n1190), .dinb(n1189), .dout(n1191));
  jand g1128(.dina(G392gat), .dinb(G188gat), .dout(n1192));
  jnot g1129(.din(n1192), .dout(n1193));
  jand g1130(.dina(n1119), .dinb(n1092), .dout(n1194));
  jand g1131(.dina(n1120), .dinb(n1089), .dout(n1195));
  jor  g1132(.dina(n1195), .dinb(n1194), .dout(n1196));
  jand g1133(.dina(G375gat), .dinb(G205gat), .dout(n1197));
  jnot g1134(.din(n1197), .dout(n1198));
  jand g1135(.dina(n1117), .dinb(n1097), .dout(n1199));
  jand g1136(.dina(n1118), .dinb(n1094), .dout(n1200));
  jor  g1137(.dina(n1200), .dinb(n1199), .dout(n1201));
  jand g1138(.dina(G358gat), .dinb(G222gat), .dout(n1202));
  jnot g1139(.din(n1202), .dout(n1203));
  jand g1140(.dina(n1115), .dinb(n1102), .dout(n1204));
  jand g1141(.dina(n1116), .dinb(n1099), .dout(n1205));
  jor  g1142(.dina(n1205), .dinb(n1204), .dout(n1206));
  jand g1143(.dina(G341gat), .dinb(G239gat), .dout(n1207));
  jand g1144(.dina(G324gat), .dinb(G256gat), .dout(n1208));
  jor  g1145(.dina(n1114), .dinb(n1103), .dout(n1209));
  jand g1146(.dina(n1209), .dinb(n1110), .dout(n1210));
  jxor g1147(.dina(n1210), .dinb(n1208), .dout(n1211));
  jnot g1148(.din(n1211), .dout(n1212));
  jxor g1149(.dina(n1212), .dinb(n1207), .dout(n1213));
  jxor g1150(.dina(n1213), .dinb(n1206), .dout(n1214));
  jxor g1151(.dina(n1214), .dinb(n1203), .dout(n1215));
  jxor g1152(.dina(n1215), .dinb(n1201), .dout(n1216));
  jxor g1153(.dina(n1216), .dinb(n1198), .dout(n1217));
  jxor g1154(.dina(n1217), .dinb(n1196), .dout(n1218));
  jxor g1155(.dina(n1218), .dinb(n1193), .dout(n1219));
  jxor g1156(.dina(n1219), .dinb(n1191), .dout(n1220));
  jxor g1157(.dina(n1220), .dinb(n1188), .dout(n1221));
  jxor g1158(.dina(n1221), .dinb(n1186), .dout(n1222));
  jxor g1159(.dina(n1222), .dinb(n1183), .dout(n1223));
  jxor g1160(.dina(n1223), .dinb(n1181), .dout(n1224));
  jxor g1161(.dina(n1224), .dinb(n1178), .dout(n1225));
  jxor g1162(.dina(n1225), .dinb(n1176), .dout(n1226));
  jxor g1163(.dina(n1226), .dinb(n1173), .dout(n1227));
  jxor g1164(.dina(n1227), .dinb(n1171), .dout(n1228));
  jxor g1165(.dina(n1228), .dinb(n1168), .dout(n1229));
  jxor g1166(.dina(n1229), .dinb(n1166), .dout(n1230));
  jxor g1167(.dina(n1230), .dinb(n1163), .dout(n1231));
  jxor g1168(.dina(n1231), .dinb(n1161), .dout(n1232));
  jxor g1169(.dina(n1232), .dinb(n1158), .dout(n1233));
  jnot g1170(.din(n1233), .dout(n1234));
  jxor g1171(.dina(n1234), .dinb(n1156), .dout(n1235));
  jnot g1172(.din(n1235), .dout(n1236));
  jxor g1173(.dina(n1236), .dinb(n1152), .dout(n1237));
  jxor g1174(.dina(n1237), .dinb(n1151), .dout(n1238));
  jnot g1175(.din(n1238), .dout(n1239));
  jxor g1176(.dina(n1239), .dinb(n1147), .dout(G6170gat));
  jnot g1177(.din(n1237), .dout(n1241));
  jor  g1178(.dina(n1241), .dinb(n1151), .dout(n1242));
  jor  g1179(.dina(n1238), .dinb(n1147), .dout(n1243));
  jand g1180(.dina(n1243), .dinb(n1242), .dout(n1244));
  jor  g1181(.dina(n1234), .dinb(n1156), .dout(n1245));
  jor  g1182(.dina(n1236), .dinb(n1152), .dout(n1246));
  jand g1183(.dina(n1246), .dinb(n1245), .dout(n1247));
  jand g1184(.dina(G528gat), .dinb(G69gat), .dout(n1248));
  jand g1185(.dina(n1231), .dinb(n1161), .dout(n1249));
  jand g1186(.dina(n1232), .dinb(n1158), .dout(n1250));
  jor  g1187(.dina(n1250), .dinb(n1249), .dout(n1251));
  jand g1188(.dina(G511gat), .dinb(G86gat), .dout(n1252));
  jnot g1189(.din(n1252), .dout(n1253));
  jand g1190(.dina(n1229), .dinb(n1166), .dout(n1254));
  jand g1191(.dina(n1230), .dinb(n1163), .dout(n1255));
  jor  g1192(.dina(n1255), .dinb(n1254), .dout(n1256));
  jand g1193(.dina(G494gat), .dinb(G103gat), .dout(n1257));
  jnot g1194(.din(n1257), .dout(n1258));
  jand g1195(.dina(n1227), .dinb(n1171), .dout(n1259));
  jand g1196(.dina(n1228), .dinb(n1168), .dout(n1260));
  jor  g1197(.dina(n1260), .dinb(n1259), .dout(n1261));
  jand g1198(.dina(G477gat), .dinb(G120gat), .dout(n1262));
  jnot g1199(.din(n1262), .dout(n1263));
  jand g1200(.dina(n1225), .dinb(n1176), .dout(n1264));
  jand g1201(.dina(n1226), .dinb(n1173), .dout(n1265));
  jor  g1202(.dina(n1265), .dinb(n1264), .dout(n1266));
  jand g1203(.dina(G460gat), .dinb(G137gat), .dout(n1267));
  jnot g1204(.din(n1267), .dout(n1268));
  jand g1205(.dina(n1223), .dinb(n1181), .dout(n1269));
  jand g1206(.dina(n1224), .dinb(n1178), .dout(n1270));
  jor  g1207(.dina(n1270), .dinb(n1269), .dout(n1271));
  jand g1208(.dina(G443gat), .dinb(G154gat), .dout(n1272));
  jnot g1209(.din(n1272), .dout(n1273));
  jand g1210(.dina(n1221), .dinb(n1186), .dout(n1274));
  jand g1211(.dina(n1222), .dinb(n1183), .dout(n1275));
  jor  g1212(.dina(n1275), .dinb(n1274), .dout(n1276));
  jand g1213(.dina(G426gat), .dinb(G171gat), .dout(n1277));
  jnot g1214(.din(n1277), .dout(n1278));
  jand g1215(.dina(n1219), .dinb(n1191), .dout(n1279));
  jand g1216(.dina(n1220), .dinb(n1188), .dout(n1280));
  jor  g1217(.dina(n1280), .dinb(n1279), .dout(n1281));
  jand g1218(.dina(G409gat), .dinb(G188gat), .dout(n1282));
  jnot g1219(.din(n1282), .dout(n1283));
  jand g1220(.dina(n1217), .dinb(n1196), .dout(n1284));
  jand g1221(.dina(n1218), .dinb(n1193), .dout(n1285));
  jor  g1222(.dina(n1285), .dinb(n1284), .dout(n1286));
  jand g1223(.dina(G392gat), .dinb(G205gat), .dout(n1287));
  jnot g1224(.din(n1287), .dout(n1288));
  jand g1225(.dina(n1215), .dinb(n1201), .dout(n1289));
  jand g1226(.dina(n1216), .dinb(n1198), .dout(n1290));
  jor  g1227(.dina(n1290), .dinb(n1289), .dout(n1291));
  jand g1228(.dina(G375gat), .dinb(G222gat), .dout(n1292));
  jnot g1229(.din(n1292), .dout(n1293));
  jand g1230(.dina(n1213), .dinb(n1206), .dout(n1294));
  jand g1231(.dina(n1214), .dinb(n1203), .dout(n1295));
  jor  g1232(.dina(n1295), .dinb(n1294), .dout(n1296));
  jand g1233(.dina(G358gat), .dinb(G239gat), .dout(n1297));
  jand g1234(.dina(G341gat), .dinb(G256gat), .dout(n1298));
  jor  g1235(.dina(n1210), .dinb(n1208), .dout(n1299));
  jor  g1236(.dina(n1212), .dinb(n1207), .dout(n1300));
  jand g1237(.dina(n1300), .dinb(n1299), .dout(n1301));
  jxor g1238(.dina(n1301), .dinb(n1298), .dout(n1302));
  jnot g1239(.din(n1302), .dout(n1303));
  jxor g1240(.dina(n1303), .dinb(n1297), .dout(n1304));
  jxor g1241(.dina(n1304), .dinb(n1296), .dout(n1305));
  jxor g1242(.dina(n1305), .dinb(n1293), .dout(n1306));
  jxor g1243(.dina(n1306), .dinb(n1291), .dout(n1307));
  jxor g1244(.dina(n1307), .dinb(n1288), .dout(n1308));
  jxor g1245(.dina(n1308), .dinb(n1286), .dout(n1309));
  jxor g1246(.dina(n1309), .dinb(n1283), .dout(n1310));
  jxor g1247(.dina(n1310), .dinb(n1281), .dout(n1311));
  jxor g1248(.dina(n1311), .dinb(n1278), .dout(n1312));
  jxor g1249(.dina(n1312), .dinb(n1276), .dout(n1313));
  jxor g1250(.dina(n1313), .dinb(n1273), .dout(n1314));
  jxor g1251(.dina(n1314), .dinb(n1271), .dout(n1315));
  jxor g1252(.dina(n1315), .dinb(n1268), .dout(n1316));
  jxor g1253(.dina(n1316), .dinb(n1266), .dout(n1317));
  jxor g1254(.dina(n1317), .dinb(n1263), .dout(n1318));
  jxor g1255(.dina(n1318), .dinb(n1261), .dout(n1319));
  jxor g1256(.dina(n1319), .dinb(n1258), .dout(n1320));
  jxor g1257(.dina(n1320), .dinb(n1256), .dout(n1321));
  jxor g1258(.dina(n1321), .dinb(n1253), .dout(n1322));
  jxor g1259(.dina(n1322), .dinb(n1251), .dout(n1323));
  jnot g1260(.din(n1323), .dout(n1324));
  jxor g1261(.dina(n1324), .dinb(n1248), .dout(n1325));
  jxor g1262(.dina(n1325), .dinb(n1247), .dout(n1326));
  jnot g1263(.din(n1326), .dout(n1327));
  jxor g1264(.dina(n1327), .dinb(n1244), .dout(G6180gat));
  jnot g1265(.din(n1325), .dout(n1329));
  jor  g1266(.dina(n1329), .dinb(n1247), .dout(n1330));
  jor  g1267(.dina(n1326), .dinb(n1244), .dout(n1331));
  jand g1268(.dina(n1331), .dinb(n1330), .dout(n1332));
  jnot g1269(.din(n1251), .dout(n1333));
  jnot g1270(.din(n1322), .dout(n1334));
  jor  g1271(.dina(n1334), .dinb(n1333), .dout(n1335));
  jor  g1272(.dina(n1324), .dinb(n1248), .dout(n1336));
  jand g1273(.dina(n1336), .dinb(n1335), .dout(n1337));
  jand g1274(.dina(G528gat), .dinb(G86gat), .dout(n1338));
  jand g1275(.dina(n1320), .dinb(n1256), .dout(n1339));
  jand g1276(.dina(n1321), .dinb(n1253), .dout(n1340));
  jor  g1277(.dina(n1340), .dinb(n1339), .dout(n1341));
  jand g1278(.dina(G511gat), .dinb(G103gat), .dout(n1342));
  jnot g1279(.din(n1342), .dout(n1343));
  jand g1280(.dina(n1318), .dinb(n1261), .dout(n1344));
  jand g1281(.dina(n1319), .dinb(n1258), .dout(n1345));
  jor  g1282(.dina(n1345), .dinb(n1344), .dout(n1346));
  jand g1283(.dina(G494gat), .dinb(G120gat), .dout(n1347));
  jnot g1284(.din(n1347), .dout(n1348));
  jand g1285(.dina(n1316), .dinb(n1266), .dout(n1349));
  jand g1286(.dina(n1317), .dinb(n1263), .dout(n1350));
  jor  g1287(.dina(n1350), .dinb(n1349), .dout(n1351));
  jand g1288(.dina(G477gat), .dinb(G137gat), .dout(n1352));
  jnot g1289(.din(n1352), .dout(n1353));
  jand g1290(.dina(n1314), .dinb(n1271), .dout(n1354));
  jand g1291(.dina(n1315), .dinb(n1268), .dout(n1355));
  jor  g1292(.dina(n1355), .dinb(n1354), .dout(n1356));
  jand g1293(.dina(G460gat), .dinb(G154gat), .dout(n1357));
  jnot g1294(.din(n1357), .dout(n1358));
  jand g1295(.dina(n1312), .dinb(n1276), .dout(n1359));
  jand g1296(.dina(n1313), .dinb(n1273), .dout(n1360));
  jor  g1297(.dina(n1360), .dinb(n1359), .dout(n1361));
  jand g1298(.dina(G443gat), .dinb(G171gat), .dout(n1362));
  jnot g1299(.din(n1362), .dout(n1363));
  jand g1300(.dina(n1310), .dinb(n1281), .dout(n1364));
  jand g1301(.dina(n1311), .dinb(n1278), .dout(n1365));
  jor  g1302(.dina(n1365), .dinb(n1364), .dout(n1366));
  jand g1303(.dina(G426gat), .dinb(G188gat), .dout(n1367));
  jnot g1304(.din(n1367), .dout(n1368));
  jand g1305(.dina(n1308), .dinb(n1286), .dout(n1369));
  jand g1306(.dina(n1309), .dinb(n1283), .dout(n1370));
  jor  g1307(.dina(n1370), .dinb(n1369), .dout(n1371));
  jand g1308(.dina(G409gat), .dinb(G205gat), .dout(n1372));
  jnot g1309(.din(n1372), .dout(n1373));
  jand g1310(.dina(n1306), .dinb(n1291), .dout(n1374));
  jand g1311(.dina(n1307), .dinb(n1288), .dout(n1375));
  jor  g1312(.dina(n1375), .dinb(n1374), .dout(n1376));
  jand g1313(.dina(G392gat), .dinb(G222gat), .dout(n1377));
  jnot g1314(.din(n1377), .dout(n1378));
  jand g1315(.dina(n1304), .dinb(n1296), .dout(n1379));
  jand g1316(.dina(n1305), .dinb(n1293), .dout(n1380));
  jor  g1317(.dina(n1380), .dinb(n1379), .dout(n1381));
  jand g1318(.dina(G375gat), .dinb(G239gat), .dout(n1382));
  jand g1319(.dina(G358gat), .dinb(G256gat), .dout(n1383));
  jor  g1320(.dina(n1301), .dinb(n1298), .dout(n1384));
  jor  g1321(.dina(n1303), .dinb(n1297), .dout(n1385));
  jand g1322(.dina(n1385), .dinb(n1384), .dout(n1386));
  jxor g1323(.dina(n1386), .dinb(n1383), .dout(n1387));
  jnot g1324(.din(n1387), .dout(n1388));
  jxor g1325(.dina(n1388), .dinb(n1382), .dout(n1389));
  jxor g1326(.dina(n1389), .dinb(n1381), .dout(n1390));
  jxor g1327(.dina(n1390), .dinb(n1378), .dout(n1391));
  jxor g1328(.dina(n1391), .dinb(n1376), .dout(n1392));
  jxor g1329(.dina(n1392), .dinb(n1373), .dout(n1393));
  jxor g1330(.dina(n1393), .dinb(n1371), .dout(n1394));
  jxor g1331(.dina(n1394), .dinb(n1368), .dout(n1395));
  jxor g1332(.dina(n1395), .dinb(n1366), .dout(n1396));
  jxor g1333(.dina(n1396), .dinb(n1363), .dout(n1397));
  jxor g1334(.dina(n1397), .dinb(n1361), .dout(n1398));
  jxor g1335(.dina(n1398), .dinb(n1358), .dout(n1399));
  jxor g1336(.dina(n1399), .dinb(n1356), .dout(n1400));
  jxor g1337(.dina(n1400), .dinb(n1353), .dout(n1401));
  jxor g1338(.dina(n1401), .dinb(n1351), .dout(n1402));
  jxor g1339(.dina(n1402), .dinb(n1348), .dout(n1403));
  jxor g1340(.dina(n1403), .dinb(n1346), .dout(n1404));
  jxor g1341(.dina(n1404), .dinb(n1343), .dout(n1405));
  jxor g1342(.dina(n1405), .dinb(n1341), .dout(n1406));
  jnot g1343(.din(n1406), .dout(n1407));
  jxor g1344(.dina(n1407), .dinb(n1338), .dout(n1408));
  jnot g1345(.din(n1408), .dout(n1409));
  jxor g1346(.dina(n1409), .dinb(n1337), .dout(n1410));
  jxor g1347(.dina(n1410), .dinb(n1332), .dout(G6190gat));
  jor  g1348(.dina(n1409), .dinb(n1337), .dout(n1412));
  jnot g1349(.din(n1410), .dout(n1413));
  jor  g1350(.dina(n1413), .dinb(n1332), .dout(n1414));
  jand g1351(.dina(n1414), .dinb(n1412), .dout(n1415));
  jnot g1352(.din(n1341), .dout(n1416));
  jnot g1353(.din(n1405), .dout(n1417));
  jor  g1354(.dina(n1417), .dinb(n1416), .dout(n1418));
  jor  g1355(.dina(n1407), .dinb(n1338), .dout(n1419));
  jand g1356(.dina(n1419), .dinb(n1418), .dout(n1420));
  jand g1357(.dina(G528gat), .dinb(G103gat), .dout(n1421));
  jand g1358(.dina(n1403), .dinb(n1346), .dout(n1422));
  jand g1359(.dina(n1404), .dinb(n1343), .dout(n1423));
  jor  g1360(.dina(n1423), .dinb(n1422), .dout(n1424));
  jand g1361(.dina(G511gat), .dinb(G120gat), .dout(n1425));
  jnot g1362(.din(n1425), .dout(n1426));
  jand g1363(.dina(n1401), .dinb(n1351), .dout(n1427));
  jand g1364(.dina(n1402), .dinb(n1348), .dout(n1428));
  jor  g1365(.dina(n1428), .dinb(n1427), .dout(n1429));
  jand g1366(.dina(G494gat), .dinb(G137gat), .dout(n1430));
  jnot g1367(.din(n1430), .dout(n1431));
  jand g1368(.dina(n1399), .dinb(n1356), .dout(n1432));
  jand g1369(.dina(n1400), .dinb(n1353), .dout(n1433));
  jor  g1370(.dina(n1433), .dinb(n1432), .dout(n1434));
  jand g1371(.dina(G477gat), .dinb(G154gat), .dout(n1435));
  jnot g1372(.din(n1435), .dout(n1436));
  jand g1373(.dina(n1397), .dinb(n1361), .dout(n1437));
  jand g1374(.dina(n1398), .dinb(n1358), .dout(n1438));
  jor  g1375(.dina(n1438), .dinb(n1437), .dout(n1439));
  jand g1376(.dina(G460gat), .dinb(G171gat), .dout(n1440));
  jnot g1377(.din(n1440), .dout(n1441));
  jand g1378(.dina(n1395), .dinb(n1366), .dout(n1442));
  jand g1379(.dina(n1396), .dinb(n1363), .dout(n1443));
  jor  g1380(.dina(n1443), .dinb(n1442), .dout(n1444));
  jand g1381(.dina(G443gat), .dinb(G188gat), .dout(n1445));
  jnot g1382(.din(n1445), .dout(n1446));
  jand g1383(.dina(n1393), .dinb(n1371), .dout(n1447));
  jand g1384(.dina(n1394), .dinb(n1368), .dout(n1448));
  jor  g1385(.dina(n1448), .dinb(n1447), .dout(n1449));
  jand g1386(.dina(G426gat), .dinb(G205gat), .dout(n1450));
  jnot g1387(.din(n1450), .dout(n1451));
  jand g1388(.dina(n1391), .dinb(n1376), .dout(n1452));
  jand g1389(.dina(n1392), .dinb(n1373), .dout(n1453));
  jor  g1390(.dina(n1453), .dinb(n1452), .dout(n1454));
  jand g1391(.dina(G409gat), .dinb(G222gat), .dout(n1455));
  jnot g1392(.din(n1455), .dout(n1456));
  jand g1393(.dina(n1389), .dinb(n1381), .dout(n1457));
  jand g1394(.dina(n1390), .dinb(n1378), .dout(n1458));
  jor  g1395(.dina(n1458), .dinb(n1457), .dout(n1459));
  jand g1396(.dina(G392gat), .dinb(G239gat), .dout(n1460));
  jand g1397(.dina(G375gat), .dinb(G256gat), .dout(n1461));
  jor  g1398(.dina(n1386), .dinb(n1383), .dout(n1462));
  jor  g1399(.dina(n1388), .dinb(n1382), .dout(n1463));
  jand g1400(.dina(n1463), .dinb(n1462), .dout(n1464));
  jxor g1401(.dina(n1464), .dinb(n1461), .dout(n1465));
  jnot g1402(.din(n1465), .dout(n1466));
  jxor g1403(.dina(n1466), .dinb(n1460), .dout(n1467));
  jxor g1404(.dina(n1467), .dinb(n1459), .dout(n1468));
  jxor g1405(.dina(n1468), .dinb(n1456), .dout(n1469));
  jxor g1406(.dina(n1469), .dinb(n1454), .dout(n1470));
  jxor g1407(.dina(n1470), .dinb(n1451), .dout(n1471));
  jxor g1408(.dina(n1471), .dinb(n1449), .dout(n1472));
  jxor g1409(.dina(n1472), .dinb(n1446), .dout(n1473));
  jxor g1410(.dina(n1473), .dinb(n1444), .dout(n1474));
  jxor g1411(.dina(n1474), .dinb(n1441), .dout(n1475));
  jxor g1412(.dina(n1475), .dinb(n1439), .dout(n1476));
  jxor g1413(.dina(n1476), .dinb(n1436), .dout(n1477));
  jxor g1414(.dina(n1477), .dinb(n1434), .dout(n1478));
  jxor g1415(.dina(n1478), .dinb(n1431), .dout(n1479));
  jxor g1416(.dina(n1479), .dinb(n1429), .dout(n1480));
  jxor g1417(.dina(n1480), .dinb(n1426), .dout(n1481));
  jxor g1418(.dina(n1481), .dinb(n1424), .dout(n1482));
  jnot g1419(.din(n1482), .dout(n1483));
  jxor g1420(.dina(n1483), .dinb(n1421), .dout(n1484));
  jnot g1421(.din(n1484), .dout(n1485));
  jxor g1422(.dina(n1485), .dinb(n1420), .dout(n1486));
  jxor g1423(.dina(n1486), .dinb(n1415), .dout(G6200gat));
  jor  g1424(.dina(n1485), .dinb(n1420), .dout(n1488));
  jnot g1425(.din(n1486), .dout(n1489));
  jor  g1426(.dina(n1489), .dinb(n1415), .dout(n1490));
  jand g1427(.dina(n1490), .dinb(n1488), .dout(n1491));
  jnot g1428(.din(n1424), .dout(n1492));
  jnot g1429(.din(n1481), .dout(n1493));
  jor  g1430(.dina(n1493), .dinb(n1492), .dout(n1494));
  jor  g1431(.dina(n1483), .dinb(n1421), .dout(n1495));
  jand g1432(.dina(n1495), .dinb(n1494), .dout(n1496));
  jand g1433(.dina(G528gat), .dinb(G120gat), .dout(n1497));
  jand g1434(.dina(n1479), .dinb(n1429), .dout(n1498));
  jand g1435(.dina(n1480), .dinb(n1426), .dout(n1499));
  jor  g1436(.dina(n1499), .dinb(n1498), .dout(n1500));
  jand g1437(.dina(G511gat), .dinb(G137gat), .dout(n1501));
  jnot g1438(.din(n1501), .dout(n1502));
  jand g1439(.dina(n1477), .dinb(n1434), .dout(n1503));
  jand g1440(.dina(n1478), .dinb(n1431), .dout(n1504));
  jor  g1441(.dina(n1504), .dinb(n1503), .dout(n1505));
  jand g1442(.dina(G494gat), .dinb(G154gat), .dout(n1506));
  jnot g1443(.din(n1506), .dout(n1507));
  jand g1444(.dina(n1475), .dinb(n1439), .dout(n1508));
  jand g1445(.dina(n1476), .dinb(n1436), .dout(n1509));
  jor  g1446(.dina(n1509), .dinb(n1508), .dout(n1510));
  jand g1447(.dina(G477gat), .dinb(G171gat), .dout(n1511));
  jnot g1448(.din(n1511), .dout(n1512));
  jand g1449(.dina(n1473), .dinb(n1444), .dout(n1513));
  jand g1450(.dina(n1474), .dinb(n1441), .dout(n1514));
  jor  g1451(.dina(n1514), .dinb(n1513), .dout(n1515));
  jand g1452(.dina(G460gat), .dinb(G188gat), .dout(n1516));
  jnot g1453(.din(n1516), .dout(n1517));
  jand g1454(.dina(n1471), .dinb(n1449), .dout(n1518));
  jand g1455(.dina(n1472), .dinb(n1446), .dout(n1519));
  jor  g1456(.dina(n1519), .dinb(n1518), .dout(n1520));
  jand g1457(.dina(G443gat), .dinb(G205gat), .dout(n1521));
  jnot g1458(.din(n1521), .dout(n1522));
  jand g1459(.dina(n1469), .dinb(n1454), .dout(n1523));
  jand g1460(.dina(n1470), .dinb(n1451), .dout(n1524));
  jor  g1461(.dina(n1524), .dinb(n1523), .dout(n1525));
  jand g1462(.dina(G426gat), .dinb(G222gat), .dout(n1526));
  jnot g1463(.din(n1526), .dout(n1527));
  jand g1464(.dina(n1467), .dinb(n1459), .dout(n1528));
  jand g1465(.dina(n1468), .dinb(n1456), .dout(n1529));
  jor  g1466(.dina(n1529), .dinb(n1528), .dout(n1530));
  jand g1467(.dina(G409gat), .dinb(G239gat), .dout(n1531));
  jand g1468(.dina(G392gat), .dinb(G256gat), .dout(n1532));
  jor  g1469(.dina(n1464), .dinb(n1461), .dout(n1533));
  jor  g1470(.dina(n1466), .dinb(n1460), .dout(n1534));
  jand g1471(.dina(n1534), .dinb(n1533), .dout(n1535));
  jxor g1472(.dina(n1535), .dinb(n1532), .dout(n1536));
  jnot g1473(.din(n1536), .dout(n1537));
  jxor g1474(.dina(n1537), .dinb(n1531), .dout(n1538));
  jxor g1475(.dina(n1538), .dinb(n1530), .dout(n1539));
  jxor g1476(.dina(n1539), .dinb(n1527), .dout(n1540));
  jxor g1477(.dina(n1540), .dinb(n1525), .dout(n1541));
  jxor g1478(.dina(n1541), .dinb(n1522), .dout(n1542));
  jxor g1479(.dina(n1542), .dinb(n1520), .dout(n1543));
  jxor g1480(.dina(n1543), .dinb(n1517), .dout(n1544));
  jxor g1481(.dina(n1544), .dinb(n1515), .dout(n1545));
  jxor g1482(.dina(n1545), .dinb(n1512), .dout(n1546));
  jxor g1483(.dina(n1546), .dinb(n1510), .dout(n1547));
  jxor g1484(.dina(n1547), .dinb(n1507), .dout(n1548));
  jxor g1485(.dina(n1548), .dinb(n1505), .dout(n1549));
  jxor g1486(.dina(n1549), .dinb(n1502), .dout(n1550));
  jxor g1487(.dina(n1550), .dinb(n1500), .dout(n1551));
  jnot g1488(.din(n1551), .dout(n1552));
  jxor g1489(.dina(n1552), .dinb(n1497), .dout(n1553));
  jnot g1490(.din(n1553), .dout(n1554));
  jxor g1491(.dina(n1554), .dinb(n1496), .dout(n1555));
  jxor g1492(.dina(n1555), .dinb(n1491), .dout(G6210gat));
  jor  g1493(.dina(n1554), .dinb(n1496), .dout(n1557));
  jnot g1494(.din(n1555), .dout(n1558));
  jor  g1495(.dina(n1558), .dinb(n1491), .dout(n1559));
  jand g1496(.dina(n1559), .dinb(n1557), .dout(n1560));
  jnot g1497(.din(n1500), .dout(n1561));
  jnot g1498(.din(n1550), .dout(n1562));
  jor  g1499(.dina(n1562), .dinb(n1561), .dout(n1563));
  jor  g1500(.dina(n1552), .dinb(n1497), .dout(n1564));
  jand g1501(.dina(n1564), .dinb(n1563), .dout(n1565));
  jand g1502(.dina(G528gat), .dinb(G137gat), .dout(n1566));
  jand g1503(.dina(n1548), .dinb(n1505), .dout(n1567));
  jand g1504(.dina(n1549), .dinb(n1502), .dout(n1568));
  jor  g1505(.dina(n1568), .dinb(n1567), .dout(n1569));
  jand g1506(.dina(G511gat), .dinb(G154gat), .dout(n1570));
  jnot g1507(.din(n1570), .dout(n1571));
  jand g1508(.dina(n1546), .dinb(n1510), .dout(n1572));
  jand g1509(.dina(n1547), .dinb(n1507), .dout(n1573));
  jor  g1510(.dina(n1573), .dinb(n1572), .dout(n1574));
  jand g1511(.dina(G494gat), .dinb(G171gat), .dout(n1575));
  jnot g1512(.din(n1575), .dout(n1576));
  jand g1513(.dina(n1544), .dinb(n1515), .dout(n1577));
  jand g1514(.dina(n1545), .dinb(n1512), .dout(n1578));
  jor  g1515(.dina(n1578), .dinb(n1577), .dout(n1579));
  jand g1516(.dina(G477gat), .dinb(G188gat), .dout(n1580));
  jnot g1517(.din(n1580), .dout(n1581));
  jand g1518(.dina(n1542), .dinb(n1520), .dout(n1582));
  jand g1519(.dina(n1543), .dinb(n1517), .dout(n1583));
  jor  g1520(.dina(n1583), .dinb(n1582), .dout(n1584));
  jand g1521(.dina(G460gat), .dinb(G205gat), .dout(n1585));
  jnot g1522(.din(n1585), .dout(n1586));
  jand g1523(.dina(n1540), .dinb(n1525), .dout(n1587));
  jand g1524(.dina(n1541), .dinb(n1522), .dout(n1588));
  jor  g1525(.dina(n1588), .dinb(n1587), .dout(n1589));
  jand g1526(.dina(G443gat), .dinb(G222gat), .dout(n1590));
  jnot g1527(.din(n1590), .dout(n1591));
  jand g1528(.dina(n1538), .dinb(n1530), .dout(n1592));
  jand g1529(.dina(n1539), .dinb(n1527), .dout(n1593));
  jor  g1530(.dina(n1593), .dinb(n1592), .dout(n1594));
  jand g1531(.dina(G426gat), .dinb(G239gat), .dout(n1595));
  jand g1532(.dina(G409gat), .dinb(G256gat), .dout(n1596));
  jor  g1533(.dina(n1535), .dinb(n1532), .dout(n1597));
  jor  g1534(.dina(n1537), .dinb(n1531), .dout(n1598));
  jand g1535(.dina(n1598), .dinb(n1597), .dout(n1599));
  jxor g1536(.dina(n1599), .dinb(n1596), .dout(n1600));
  jnot g1537(.din(n1600), .dout(n1601));
  jxor g1538(.dina(n1601), .dinb(n1595), .dout(n1602));
  jxor g1539(.dina(n1602), .dinb(n1594), .dout(n1603));
  jxor g1540(.dina(n1603), .dinb(n1591), .dout(n1604));
  jxor g1541(.dina(n1604), .dinb(n1589), .dout(n1605));
  jxor g1542(.dina(n1605), .dinb(n1586), .dout(n1606));
  jxor g1543(.dina(n1606), .dinb(n1584), .dout(n1607));
  jxor g1544(.dina(n1607), .dinb(n1581), .dout(n1608));
  jxor g1545(.dina(n1608), .dinb(n1579), .dout(n1609));
  jxor g1546(.dina(n1609), .dinb(n1576), .dout(n1610));
  jxor g1547(.dina(n1610), .dinb(n1574), .dout(n1611));
  jxor g1548(.dina(n1611), .dinb(n1571), .dout(n1612));
  jxor g1549(.dina(n1612), .dinb(n1569), .dout(n1613));
  jnot g1550(.din(n1613), .dout(n1614));
  jxor g1551(.dina(n1614), .dinb(n1566), .dout(n1615));
  jnot g1552(.din(n1615), .dout(n1616));
  jxor g1553(.dina(n1616), .dinb(n1565), .dout(n1617));
  jxor g1554(.dina(n1617), .dinb(n1560), .dout(G6220gat));
  jor  g1555(.dina(n1616), .dinb(n1565), .dout(n1619));
  jnot g1556(.din(n1617), .dout(n1620));
  jor  g1557(.dina(n1620), .dinb(n1560), .dout(n1621));
  jand g1558(.dina(n1621), .dinb(n1619), .dout(n1622));
  jnot g1559(.din(n1569), .dout(n1623));
  jnot g1560(.din(n1612), .dout(n1624));
  jor  g1561(.dina(n1624), .dinb(n1623), .dout(n1625));
  jor  g1562(.dina(n1614), .dinb(n1566), .dout(n1626));
  jand g1563(.dina(n1626), .dinb(n1625), .dout(n1627));
  jand g1564(.dina(G528gat), .dinb(G154gat), .dout(n1628));
  jand g1565(.dina(n1610), .dinb(n1574), .dout(n1629));
  jand g1566(.dina(n1611), .dinb(n1571), .dout(n1630));
  jor  g1567(.dina(n1630), .dinb(n1629), .dout(n1631));
  jand g1568(.dina(G511gat), .dinb(G171gat), .dout(n1632));
  jnot g1569(.din(n1632), .dout(n1633));
  jand g1570(.dina(n1608), .dinb(n1579), .dout(n1634));
  jand g1571(.dina(n1609), .dinb(n1576), .dout(n1635));
  jor  g1572(.dina(n1635), .dinb(n1634), .dout(n1636));
  jand g1573(.dina(G494gat), .dinb(G188gat), .dout(n1637));
  jnot g1574(.din(n1637), .dout(n1638));
  jand g1575(.dina(n1606), .dinb(n1584), .dout(n1639));
  jand g1576(.dina(n1607), .dinb(n1581), .dout(n1640));
  jor  g1577(.dina(n1640), .dinb(n1639), .dout(n1641));
  jand g1578(.dina(G477gat), .dinb(G205gat), .dout(n1642));
  jnot g1579(.din(n1642), .dout(n1643));
  jand g1580(.dina(n1604), .dinb(n1589), .dout(n1644));
  jand g1581(.dina(n1605), .dinb(n1586), .dout(n1645));
  jor  g1582(.dina(n1645), .dinb(n1644), .dout(n1646));
  jand g1583(.dina(G460gat), .dinb(G222gat), .dout(n1647));
  jnot g1584(.din(n1647), .dout(n1648));
  jand g1585(.dina(n1602), .dinb(n1594), .dout(n1649));
  jand g1586(.dina(n1603), .dinb(n1591), .dout(n1650));
  jor  g1587(.dina(n1650), .dinb(n1649), .dout(n1651));
  jand g1588(.dina(G443gat), .dinb(G239gat), .dout(n1652));
  jand g1589(.dina(G426gat), .dinb(G256gat), .dout(n1653));
  jor  g1590(.dina(n1599), .dinb(n1596), .dout(n1654));
  jor  g1591(.dina(n1601), .dinb(n1595), .dout(n1655));
  jand g1592(.dina(n1655), .dinb(n1654), .dout(n1656));
  jxor g1593(.dina(n1656), .dinb(n1653), .dout(n1657));
  jnot g1594(.din(n1657), .dout(n1658));
  jxor g1595(.dina(n1658), .dinb(n1652), .dout(n1659));
  jxor g1596(.dina(n1659), .dinb(n1651), .dout(n1660));
  jxor g1597(.dina(n1660), .dinb(n1648), .dout(n1661));
  jxor g1598(.dina(n1661), .dinb(n1646), .dout(n1662));
  jxor g1599(.dina(n1662), .dinb(n1643), .dout(n1663));
  jxor g1600(.dina(n1663), .dinb(n1641), .dout(n1664));
  jxor g1601(.dina(n1664), .dinb(n1638), .dout(n1665));
  jxor g1602(.dina(n1665), .dinb(n1636), .dout(n1666));
  jxor g1603(.dina(n1666), .dinb(n1633), .dout(n1667));
  jxor g1604(.dina(n1667), .dinb(n1631), .dout(n1668));
  jnot g1605(.din(n1668), .dout(n1669));
  jxor g1606(.dina(n1669), .dinb(n1628), .dout(n1670));
  jnot g1607(.din(n1670), .dout(n1671));
  jxor g1608(.dina(n1671), .dinb(n1627), .dout(n1672));
  jxor g1609(.dina(n1672), .dinb(n1622), .dout(G6230gat));
  jor  g1610(.dina(n1671), .dinb(n1627), .dout(n1674));
  jnot g1611(.din(n1672), .dout(n1675));
  jor  g1612(.dina(n1675), .dinb(n1622), .dout(n1676));
  jand g1613(.dina(n1676), .dinb(n1674), .dout(n1677));
  jnot g1614(.din(n1631), .dout(n1678));
  jnot g1615(.din(n1667), .dout(n1679));
  jor  g1616(.dina(n1679), .dinb(n1678), .dout(n1680));
  jor  g1617(.dina(n1669), .dinb(n1628), .dout(n1681));
  jand g1618(.dina(n1681), .dinb(n1680), .dout(n1682));
  jand g1619(.dina(G528gat), .dinb(G171gat), .dout(n1683));
  jnot g1620(.din(n1683), .dout(n1684));
  jand g1621(.dina(n1665), .dinb(n1636), .dout(n1685));
  jand g1622(.dina(n1666), .dinb(n1633), .dout(n1686));
  jor  g1623(.dina(n1686), .dinb(n1685), .dout(n1687));
  jand g1624(.dina(G511gat), .dinb(G188gat), .dout(n1688));
  jnot g1625(.din(n1688), .dout(n1689));
  jand g1626(.dina(n1663), .dinb(n1641), .dout(n1690));
  jand g1627(.dina(n1664), .dinb(n1638), .dout(n1691));
  jor  g1628(.dina(n1691), .dinb(n1690), .dout(n1692));
  jand g1629(.dina(G494gat), .dinb(G205gat), .dout(n1693));
  jnot g1630(.din(n1693), .dout(n1694));
  jand g1631(.dina(n1661), .dinb(n1646), .dout(n1695));
  jand g1632(.dina(n1662), .dinb(n1643), .dout(n1696));
  jor  g1633(.dina(n1696), .dinb(n1695), .dout(n1697));
  jand g1634(.dina(G477gat), .dinb(G222gat), .dout(n1698));
  jnot g1635(.din(n1698), .dout(n1699));
  jand g1636(.dina(n1659), .dinb(n1651), .dout(n1700));
  jand g1637(.dina(n1660), .dinb(n1648), .dout(n1701));
  jor  g1638(.dina(n1701), .dinb(n1700), .dout(n1702));
  jand g1639(.dina(G460gat), .dinb(G239gat), .dout(n1703));
  jand g1640(.dina(G443gat), .dinb(G256gat), .dout(n1704));
  jor  g1641(.dina(n1656), .dinb(n1653), .dout(n1705));
  jor  g1642(.dina(n1658), .dinb(n1652), .dout(n1706));
  jand g1643(.dina(n1706), .dinb(n1705), .dout(n1707));
  jxor g1644(.dina(n1707), .dinb(n1704), .dout(n1708));
  jnot g1645(.din(n1708), .dout(n1709));
  jxor g1646(.dina(n1709), .dinb(n1703), .dout(n1710));
  jxor g1647(.dina(n1710), .dinb(n1702), .dout(n1711));
  jxor g1648(.dina(n1711), .dinb(n1699), .dout(n1712));
  jxor g1649(.dina(n1712), .dinb(n1697), .dout(n1713));
  jxor g1650(.dina(n1713), .dinb(n1694), .dout(n1714));
  jxor g1651(.dina(n1714), .dinb(n1692), .dout(n1715));
  jxor g1652(.dina(n1715), .dinb(n1689), .dout(n1716));
  jxor g1653(.dina(n1716), .dinb(n1687), .dout(n1717));
  jxor g1654(.dina(n1717), .dinb(n1684), .dout(n1718));
  jnot g1655(.din(n1718), .dout(n1719));
  jxor g1656(.dina(n1719), .dinb(n1682), .dout(n1720));
  jxor g1657(.dina(n1720), .dinb(n1677), .dout(G6240gat));
  jor  g1658(.dina(n1719), .dinb(n1682), .dout(n1722));
  jnot g1659(.din(n1720), .dout(n1723));
  jor  g1660(.dina(n1723), .dinb(n1677), .dout(n1724));
  jand g1661(.dina(n1724), .dinb(n1722), .dout(n1725));
  jand g1662(.dina(n1716), .dinb(n1687), .dout(n1726));
  jand g1663(.dina(n1717), .dinb(n1684), .dout(n1727));
  jor  g1664(.dina(n1727), .dinb(n1726), .dout(n1728));
  jand g1665(.dina(G528gat), .dinb(G188gat), .dout(n1729));
  jnot g1666(.din(n1729), .dout(n1730));
  jand g1667(.dina(n1714), .dinb(n1692), .dout(n1731));
  jand g1668(.dina(n1715), .dinb(n1689), .dout(n1732));
  jor  g1669(.dina(n1732), .dinb(n1731), .dout(n1733));
  jand g1670(.dina(G511gat), .dinb(G205gat), .dout(n1734));
  jnot g1671(.din(n1734), .dout(n1735));
  jand g1672(.dina(n1712), .dinb(n1697), .dout(n1736));
  jand g1673(.dina(n1713), .dinb(n1694), .dout(n1737));
  jor  g1674(.dina(n1737), .dinb(n1736), .dout(n1738));
  jand g1675(.dina(G494gat), .dinb(G222gat), .dout(n1739));
  jnot g1676(.din(n1739), .dout(n1740));
  jand g1677(.dina(n1710), .dinb(n1702), .dout(n1741));
  jand g1678(.dina(n1711), .dinb(n1699), .dout(n1742));
  jor  g1679(.dina(n1742), .dinb(n1741), .dout(n1743));
  jand g1680(.dina(G477gat), .dinb(G239gat), .dout(n1744));
  jand g1681(.dina(G460gat), .dinb(G256gat), .dout(n1745));
  jor  g1682(.dina(n1707), .dinb(n1704), .dout(n1746));
  jor  g1683(.dina(n1709), .dinb(n1703), .dout(n1747));
  jand g1684(.dina(n1747), .dinb(n1746), .dout(n1748));
  jxor g1685(.dina(n1748), .dinb(n1745), .dout(n1749));
  jnot g1686(.din(n1749), .dout(n1750));
  jxor g1687(.dina(n1750), .dinb(n1744), .dout(n1751));
  jxor g1688(.dina(n1751), .dinb(n1743), .dout(n1752));
  jxor g1689(.dina(n1752), .dinb(n1740), .dout(n1753));
  jxor g1690(.dina(n1753), .dinb(n1738), .dout(n1754));
  jxor g1691(.dina(n1754), .dinb(n1735), .dout(n1755));
  jxor g1692(.dina(n1755), .dinb(n1733), .dout(n1756));
  jxor g1693(.dina(n1756), .dinb(n1730), .dout(n1757));
  jxor g1694(.dina(n1757), .dinb(n1728), .dout(n1758));
  jxor g1695(.dina(n1758), .dinb(n1725), .dout(G6250gat));
  jnot g1696(.din(n1728), .dout(n1760));
  jnot g1697(.din(n1757), .dout(n1761));
  jor  g1698(.dina(n1761), .dinb(n1760), .dout(n1762));
  jnot g1699(.din(n1758), .dout(n1763));
  jor  g1700(.dina(n1763), .dinb(n1725), .dout(n1764));
  jand g1701(.dina(n1764), .dinb(n1762), .dout(n1765));
  jand g1702(.dina(n1755), .dinb(n1733), .dout(n1766));
  jand g1703(.dina(n1756), .dinb(n1730), .dout(n1767));
  jor  g1704(.dina(n1767), .dinb(n1766), .dout(n1768));
  jand g1705(.dina(G528gat), .dinb(G205gat), .dout(n1769));
  jnot g1706(.din(n1769), .dout(n1770));
  jand g1707(.dina(n1753), .dinb(n1738), .dout(n1771));
  jand g1708(.dina(n1754), .dinb(n1735), .dout(n1772));
  jor  g1709(.dina(n1772), .dinb(n1771), .dout(n1773));
  jand g1710(.dina(G511gat), .dinb(G222gat), .dout(n1774));
  jnot g1711(.din(n1774), .dout(n1775));
  jand g1712(.dina(n1751), .dinb(n1743), .dout(n1776));
  jand g1713(.dina(n1752), .dinb(n1740), .dout(n1777));
  jor  g1714(.dina(n1777), .dinb(n1776), .dout(n1778));
  jand g1715(.dina(G494gat), .dinb(G239gat), .dout(n1779));
  jand g1716(.dina(G477gat), .dinb(G256gat), .dout(n1780));
  jor  g1717(.dina(n1748), .dinb(n1745), .dout(n1781));
  jor  g1718(.dina(n1750), .dinb(n1744), .dout(n1782));
  jand g1719(.dina(n1782), .dinb(n1781), .dout(n1783));
  jxor g1720(.dina(n1783), .dinb(n1780), .dout(n1784));
  jnot g1721(.din(n1784), .dout(n1785));
  jxor g1722(.dina(n1785), .dinb(n1779), .dout(n1786));
  jxor g1723(.dina(n1786), .dinb(n1778), .dout(n1787));
  jxor g1724(.dina(n1787), .dinb(n1775), .dout(n1788));
  jxor g1725(.dina(n1788), .dinb(n1773), .dout(n1789));
  jxor g1726(.dina(n1789), .dinb(n1770), .dout(n1790));
  jxor g1727(.dina(n1790), .dinb(n1768), .dout(n1791));
  jxor g1728(.dina(n1791), .dinb(n1765), .dout(G6260gat));
  jnot g1729(.din(n1768), .dout(n1793));
  jnot g1730(.din(n1790), .dout(n1794));
  jor  g1731(.dina(n1794), .dinb(n1793), .dout(n1795));
  jnot g1732(.din(n1791), .dout(n1796));
  jor  g1733(.dina(n1796), .dinb(n1765), .dout(n1797));
  jand g1734(.dina(n1797), .dinb(n1795), .dout(n1798));
  jand g1735(.dina(n1788), .dinb(n1773), .dout(n1799));
  jand g1736(.dina(n1789), .dinb(n1770), .dout(n1800));
  jor  g1737(.dina(n1800), .dinb(n1799), .dout(n1801));
  jand g1738(.dina(G528gat), .dinb(G222gat), .dout(n1802));
  jnot g1739(.din(n1802), .dout(n1803));
  jand g1740(.dina(n1786), .dinb(n1778), .dout(n1804));
  jand g1741(.dina(n1787), .dinb(n1775), .dout(n1805));
  jor  g1742(.dina(n1805), .dinb(n1804), .dout(n1806));
  jand g1743(.dina(G511gat), .dinb(G239gat), .dout(n1807));
  jand g1744(.dina(G494gat), .dinb(G256gat), .dout(n1808));
  jor  g1745(.dina(n1783), .dinb(n1780), .dout(n1809));
  jor  g1746(.dina(n1785), .dinb(n1779), .dout(n1810));
  jand g1747(.dina(n1810), .dinb(n1809), .dout(n1811));
  jxor g1748(.dina(n1811), .dinb(n1808), .dout(n1812));
  jnot g1749(.din(n1812), .dout(n1813));
  jxor g1750(.dina(n1813), .dinb(n1807), .dout(n1814));
  jxor g1751(.dina(n1814), .dinb(n1806), .dout(n1815));
  jxor g1752(.dina(n1815), .dinb(n1803), .dout(n1816));
  jxor g1753(.dina(n1816), .dinb(n1801), .dout(n1817));
  jxor g1754(.dina(n1817), .dinb(n1798), .dout(G6270gat));
  jnot g1755(.din(n1801), .dout(n1819));
  jnot g1756(.din(n1816), .dout(n1820));
  jor  g1757(.dina(n1820), .dinb(n1819), .dout(n1821));
  jnot g1758(.din(n1817), .dout(n1822));
  jor  g1759(.dina(n1822), .dinb(n1798), .dout(n1823));
  jand g1760(.dina(n1823), .dinb(n1821), .dout(n1824));
  jand g1761(.dina(n1814), .dinb(n1806), .dout(n1825));
  jand g1762(.dina(n1815), .dinb(n1803), .dout(n1826));
  jor  g1763(.dina(n1826), .dinb(n1825), .dout(n1827));
  jand g1764(.dina(G528gat), .dinb(G239gat), .dout(n1828));
  jand g1765(.dina(G511gat), .dinb(G256gat), .dout(n1829));
  jor  g1766(.dina(n1811), .dinb(n1808), .dout(n1830));
  jor  g1767(.dina(n1813), .dinb(n1807), .dout(n1831));
  jand g1768(.dina(n1831), .dinb(n1830), .dout(n1832));
  jxor g1769(.dina(n1832), .dinb(n1829), .dout(n1833));
  jnot g1770(.din(n1833), .dout(n1834));
  jxor g1771(.dina(n1834), .dinb(n1828), .dout(n1835));
  jxor g1772(.dina(n1835), .dinb(n1827), .dout(n1836));
  jxor g1773(.dina(n1836), .dinb(n1824), .dout(G6280gat));
  jand g1774(.dina(G528gat), .dinb(G256gat), .dout(n1838));
  jor  g1775(.dina(n1832), .dinb(n1829), .dout(n1839));
  jor  g1776(.dina(n1834), .dinb(n1828), .dout(n1840));
  jand g1777(.dina(n1840), .dinb(n1839), .dout(n1841));
  jor  g1778(.dina(n1841), .dinb(n1838), .dout(n1842));
  jnot g1779(.din(n1827), .dout(n1843));
  jnot g1780(.din(n1835), .dout(n1844));
  jor  g1781(.dina(n1844), .dinb(n1843), .dout(n1845));
  jnot g1782(.din(n1836), .dout(n1846));
  jor  g1783(.dina(n1846), .dinb(n1824), .dout(n1847));
  jand g1784(.dina(n1847), .dinb(n1845), .dout(n1848));
  jxor g1785(.dina(n1841), .dinb(n1838), .dout(n1849));
  jnot g1786(.din(n1849), .dout(n1850));
  jor  g1787(.dina(n1850), .dinb(n1848), .dout(n1851));
  jand g1788(.dina(n1851), .dinb(n1842), .dout(G6287gat));
  jxor g1789(.dina(n1849), .dinb(n1848), .dout(G6288gat));
endmodule


