/*
gf_c1355:
	jxor: 108
	jspl: 34
	jspl3: 68
	jnot: 17
	jdff: 509
	jand: 65
	jor: 6

Summary:
	jxor: 108
	jspl: 34
	jspl3: 68
	jnot: 17
	jdff: 509
	jand: 65
	jor: 6

The maximum logic level gap of any gate:
	gf_c1355: 11
*/

module gf_c1355(gclk, G1gat, G8gat, G15gat, G22gat, G29gat, G36gat, G43gat, G50gat, G57gat, G64gat, G71gat, G78gat, G85gat, G92gat, G99gat, G106gat, G113gat, G120gat, G127gat, G134gat, G141gat, G148gat, G155gat, G162gat, G169gat, G176gat, G183gat, G190gat, G197gat, G204gat, G211gat, G218gat, G225gat, G226gat, G227gat, G228gat, G229gat, G230gat, G231gat, G232gat, G233gat, G1324gat, G1325gat, G1326gat, G1327gat, G1328gat, G1329gat, G1330gat, G1331gat, G1332gat, G1333gat, G1334gat, G1335gat, G1336gat, G1337gat, G1338gat, G1339gat, G1340gat, G1341gat, G1342gat, G1343gat, G1344gat, G1345gat, G1346gat, G1347gat, G1348gat, G1349gat, G1350gat, G1351gat, G1352gat, G1353gat, G1354gat, G1355gat);
	input gclk;
	input G1gat;
	input G8gat;
	input G15gat;
	input G22gat;
	input G29gat;
	input G36gat;
	input G43gat;
	input G50gat;
	input G57gat;
	input G64gat;
	input G71gat;
	input G78gat;
	input G85gat;
	input G92gat;
	input G99gat;
	input G106gat;
	input G113gat;
	input G120gat;
	input G127gat;
	input G134gat;
	input G141gat;
	input G148gat;
	input G155gat;
	input G162gat;
	input G169gat;
	input G176gat;
	input G183gat;
	input G190gat;
	input G197gat;
	input G204gat;
	input G211gat;
	input G218gat;
	input G225gat;
	input G226gat;
	input G227gat;
	input G228gat;
	input G229gat;
	input G230gat;
	input G231gat;
	input G232gat;
	input G233gat;
	output G1324gat;
	output G1325gat;
	output G1326gat;
	output G1327gat;
	output G1328gat;
	output G1329gat;
	output G1330gat;
	output G1331gat;
	output G1332gat;
	output G1333gat;
	output G1334gat;
	output G1335gat;
	output G1336gat;
	output G1337gat;
	output G1338gat;
	output G1339gat;
	output G1340gat;
	output G1341gat;
	output G1342gat;
	output G1343gat;
	output G1344gat;
	output G1345gat;
	output G1346gat;
	output G1347gat;
	output G1348gat;
	output G1349gat;
	output G1350gat;
	output G1351gat;
	output G1352gat;
	output G1353gat;
	output G1354gat;
	output G1355gat;
	wire n73;
	wire n74;
	wire n75;
	wire n76;
	wire n77;
	wire n78;
	wire n79;
	wire n80;
	wire n81;
	wire n82;
	wire n83;
	wire n84;
	wire n85;
	wire n86;
	wire n87;
	wire n88;
	wire n89;
	wire n90;
	wire n91;
	wire n92;
	wire n93;
	wire n94;
	wire n95;
	wire n96;
	wire n97;
	wire n98;
	wire n99;
	wire n100;
	wire n101;
	wire n102;
	wire n103;
	wire n104;
	wire n105;
	wire n106;
	wire n107;
	wire n108;
	wire n109;
	wire n110;
	wire n111;
	wire n112;
	wire n113;
	wire n114;
	wire n115;
	wire n116;
	wire n117;
	wire n118;
	wire n119;
	wire n120;
	wire n121;
	wire n122;
	wire n123;
	wire n124;
	wire n125;
	wire n126;
	wire n127;
	wire n128;
	wire n129;
	wire n130;
	wire n131;
	wire n132;
	wire n133;
	wire n134;
	wire n135;
	wire n136;
	wire n137;
	wire n138;
	wire n139;
	wire n140;
	wire n141;
	wire n142;
	wire n143;
	wire n144;
	wire n145;
	wire n146;
	wire n147;
	wire n148;
	wire n149;
	wire n150;
	wire n151;
	wire n152;
	wire n153;
	wire n154;
	wire n155;
	wire n156;
	wire n157;
	wire n158;
	wire n159;
	wire n160;
	wire n161;
	wire n162;
	wire n163;
	wire n164;
	wire n165;
	wire n166;
	wire n167;
	wire n168;
	wire n169;
	wire n170;
	wire n171;
	wire n172;
	wire n173;
	wire n174;
	wire n175;
	wire n176;
	wire n178;
	wire n179;
	wire n181;
	wire n182;
	wire n184;
	wire n185;
	wire n187;
	wire n188;
	wire n189;
	wire n190;
	wire n191;
	wire n193;
	wire n195;
	wire n197;
	wire n199;
	wire n200;
	wire n201;
	wire n202;
	wire n203;
	wire n205;
	wire n207;
	wire n209;
	wire n211;
	wire n212;
	wire n214;
	wire n216;
	wire n218;
	wire n220;
	wire n221;
	wire n222;
	wire n223;
	wire n224;
	wire n225;
	wire n226;
	wire n227;
	wire n228;
	wire n229;
	wire n230;
	wire n231;
	wire n233;
	wire n235;
	wire n237;
	wire n239;
	wire n240;
	wire n241;
	wire n243;
	wire n245;
	wire n247;
	wire n249;
	wire n250;
	wire n251;
	wire n252;
	wire n254;
	wire n256;
	wire n258;
	wire n260;
	wire n261;
	wire n263;
	wire n265;
	wire n267;
	wire [2:0] w_G1gat_0;
	wire [2:0] w_G8gat_0;
	wire [2:0] w_G15gat_0;
	wire [2:0] w_G22gat_0;
	wire [2:0] w_G29gat_0;
	wire [2:0] w_G36gat_0;
	wire [2:0] w_G43gat_0;
	wire [2:0] w_G50gat_0;
	wire [2:0] w_G57gat_0;
	wire [2:0] w_G64gat_0;
	wire [2:0] w_G71gat_0;
	wire [2:0] w_G78gat_0;
	wire [2:0] w_G85gat_0;
	wire [2:0] w_G92gat_0;
	wire [2:0] w_G99gat_0;
	wire [2:0] w_G106gat_0;
	wire [2:0] w_G113gat_0;
	wire [2:0] w_G120gat_0;
	wire [2:0] w_G127gat_0;
	wire [2:0] w_G134gat_0;
	wire [2:0] w_G141gat_0;
	wire [2:0] w_G148gat_0;
	wire [2:0] w_G155gat_0;
	wire [2:0] w_G162gat_0;
	wire [2:0] w_G169gat_0;
	wire [2:0] w_G176gat_0;
	wire [2:0] w_G183gat_0;
	wire [2:0] w_G190gat_0;
	wire [2:0] w_G197gat_0;
	wire [2:0] w_G204gat_0;
	wire [2:0] w_G211gat_0;
	wire [2:0] w_G218gat_0;
	wire [2:0] w_G233gat_0;
	wire [2:0] w_G233gat_1;
	wire [1:0] w_n78_0;
	wire [1:0] w_n84_0;
	wire [2:0] w_n86_0;
	wire [1:0] w_n86_1;
	wire [2:0] w_n87_0;
	wire [2:0] w_n87_1;
	wire [1:0] w_n93_0;
	wire [2:0] w_n96_0;
	wire [1:0] w_n96_1;
	wire [1:0] w_n100_0;
	wire [2:0] w_n102_0;
	wire [1:0] w_n102_1;
	wire [1:0] w_n108_0;
	wire [1:0] w_n114_0;
	wire [2:0] w_n116_0;
	wire [1:0] w_n116_1;
	wire [2:0] w_n117_0;
	wire [2:0] w_n117_1;
	wire [1:0] w_n118_0;
	wire [1:0] w_n124_0;
	wire [1:0] w_n130_0;
	wire [2:0] w_n132_0;
	wire [1:0] w_n132_1;
	wire [2:0] w_n141_0;
	wire [1:0] w_n141_1;
	wire [2:0] w_n149_0;
	wire [1:0] w_n149_1;
	wire [2:0] w_n155_0;
	wire [2:0] w_n163_0;
	wire [1:0] w_n163_1;
	wire [2:0] w_n164_0;
	wire [2:0] w_n164_1;
	wire [2:0] w_n172_0;
	wire [1:0] w_n172_1;
	wire [1:0] w_n173_0;
	wire [2:0] w_n175_0;
	wire [1:0] w_n175_1;
	wire [2:0] w_n178_0;
	wire [2:0] w_n178_1;
	wire [2:0] w_n181_0;
	wire [2:0] w_n181_1;
	wire [2:0] w_n184_0;
	wire [2:0] w_n184_1;
	wire [2:0] w_n187_0;
	wire [2:0] w_n187_1;
	wire [1:0] w_n189_0;
	wire [2:0] w_n190_0;
	wire [1:0] w_n190_1;
	wire [2:0] w_n199_0;
	wire [2:0] w_n199_1;
	wire [1:0] w_n200_0;
	wire [2:0] w_n202_0;
	wire [1:0] w_n202_1;
	wire [2:0] w_n211_0;
	wire [1:0] w_n211_1;
	wire [1:0] w_n220_0;
	wire [1:0] w_n228_0;
	wire [1:0] w_n229_0;
	wire [2:0] w_n230_0;
	wire [1:0] w_n230_1;
	wire [1:0] w_n239_0;
	wire [2:0] w_n240_0;
	wire [1:0] w_n240_1;
	wire [1:0] w_n250_0;
	wire [2:0] w_n251_0;
	wire [1:0] w_n251_1;
	wire [2:0] w_n260_0;
	wire [1:0] w_n260_1;
	wire w_dff_A_g7fWtRC34_0;
	wire w_dff_B_UbdA9TpT0_2;
	wire w_dff_B_XLzfbrYo1_2;
	wire w_dff_A_XFMs5PF89_1;
	wire w_dff_B_C82Ol07Z2_2;
	wire w_dff_B_cMdmeUqR9_2;
	wire w_dff_B_oD2VeBYI1_2;
	wire w_dff_B_uXMssaTF3_2;
	wire w_dff_B_ictF7VVB8_2;
	wire w_dff_B_fEXmCUEr6_0;
	wire w_dff_B_qvVbhgQM2_0;
	wire w_dff_B_IfNW47ib0_1;
	wire w_dff_A_4kRfFieY2_0;
	wire w_dff_A_qvU4pT7M9_0;
	wire w_dff_A_w5BUOEI76_0;
	wire w_dff_A_WOeCCUnT6_0;
	wire w_dff_A_pjcl3KMO5_0;
	wire w_dff_A_bM5Ydb574_0;
	wire w_dff_A_FZGlmU2N4_0;
	wire w_dff_A_GY3GUQUV5_1;
	wire w_dff_A_bbxDdLtV6_1;
	wire w_dff_A_a0vgmC6X2_1;
	wire w_dff_A_xdfdtWBd6_1;
	wire w_dff_A_sFVdG6WN0_1;
	wire w_dff_A_qJ5zHxs81_0;
	wire w_dff_A_K1PQJV6P4_0;
	wire w_dff_A_Fo4NdyDl9_0;
	wire w_dff_A_cNwRv10B6_0;
	wire w_dff_A_iuTgCrL40_0;
	wire w_dff_A_0mjTla9J4_1;
	wire w_dff_A_MkIJKXmu7_1;
	wire w_dff_A_Br5tP2ke6_1;
	wire w_dff_A_kJVItLlC5_1;
	wire w_dff_A_pFx1qlrF2_1;
	wire w_dff_A_NyHcnITN2_0;
	wire w_dff_A_PjEsC2Nt6_0;
	wire w_dff_A_9hMNiwAr7_0;
	wire w_dff_A_3FNVJZ6b6_0;
	wire w_dff_A_BvcpixTz4_0;
	wire w_dff_A_OhMm5bUl1_1;
	wire w_dff_A_FNmPuiPJ4_1;
	wire w_dff_A_wzYEryQA7_1;
	wire w_dff_A_NlQU0y8n4_1;
	wire w_dff_A_ANbbw8Pr3_1;
	wire w_dff_B_I3NQ9kWv8_1;
	wire w_dff_B_X2Im87NO5_1;
	wire w_dff_A_nkRXkBK28_0;
	wire w_dff_A_y2E5kge90_0;
	wire w_dff_A_N0Qm4qx03_0;
	wire w_dff_A_KE3xKRPJ8_0;
	wire w_dff_A_HDvR5fGe3_0;
	wire w_dff_A_r5DYRlB56_2;
	wire w_dff_A_EXqygMbt8_2;
	wire w_dff_A_8TN8oAwb5_2;
	wire w_dff_A_kg3pIg939_2;
	wire w_dff_A_7DImgA5K9_2;
	wire w_dff_A_oCgw7TMx6_0;
	wire w_dff_A_I1aMf9ZZ5_0;
	wire w_dff_A_YeY29Oym9_0;
	wire w_dff_A_zBAy3kXJ3_0;
	wire w_dff_A_pFG4FcaY0_0;
	wire w_dff_A_OnF2YcdG6_1;
	wire w_dff_A_mPYlZrow8_1;
	wire w_dff_A_fx5E7a5D4_1;
	wire w_dff_A_CitHGTA41_1;
	wire w_dff_A_2DYJGpGs2_1;
	wire w_dff_B_Bvp8kghG2_2;
	wire w_dff_B_hw1dCfcE1_2;
	wire w_dff_B_ZnnCJ2u80_2;
	wire w_dff_A_tAxc8FNh3_0;
	wire w_dff_A_H9RAuYj59_0;
	wire w_dff_A_zhKE0ORh8_0;
	wire w_dff_A_978ixOg97_0;
	wire w_dff_A_Z09T7J496_0;
	wire w_dff_A_9vEsrmUR1_2;
	wire w_dff_A_3GTNAkxF1_2;
	wire w_dff_A_S26JRI2o8_2;
	wire w_dff_A_hf96O2073_2;
	wire w_dff_A_KepHnE5C4_2;
	wire w_dff_A_Pq1Q8flQ6_1;
	wire w_dff_A_tiXy71DX0_1;
	wire w_dff_A_J1RAxLIK9_1;
	wire w_dff_A_xA55UyWX5_1;
	wire w_dff_A_fiIPpVW66_1;
	wire w_dff_A_IZxkOlFJ1_2;
	wire w_dff_A_PRQAdJrd6_2;
	wire w_dff_A_ruYlIlni4_2;
	wire w_dff_A_OatywFOG1_2;
	wire w_dff_A_neoNnWwU3_2;
	wire w_dff_A_9woERz7Z9_0;
	wire w_dff_A_cI7o6xKU6_1;
	wire w_dff_A_p6IPhVq52_1;
	wire w_dff_A_x5ATtBGA0_1;
	wire w_dff_A_s89WmVE65_1;
	wire w_dff_A_Pt4jPtr59_1;
	wire w_dff_A_jw7x2tkw3_2;
	wire w_dff_A_6WsW1NfW8_2;
	wire w_dff_A_ShANqaSA1_2;
	wire w_dff_A_qOihlfpz6_2;
	wire w_dff_A_dDSIcMPD8_2;
	wire w_dff_A_Y51j7kVV7_1;
	wire w_dff_A_NqSOUP0c2_1;
	wire w_dff_A_G3ZB9A949_1;
	wire w_dff_A_chUHDdp50_1;
	wire w_dff_A_kjcJgFsq5_1;
	wire w_dff_A_C2tRsLlm2_1;
	wire w_dff_A_7ayfKDEO3_2;
	wire w_dff_A_2uRtdZbc2_2;
	wire w_dff_A_4uP4cjSF1_2;
	wire w_dff_A_grZsy7Tu6_2;
	wire w_dff_A_6rL5Wax43_2;
	wire w_dff_A_rIYE9OzL2_0;
	wire w_dff_B_qyGoOx4d0_1;
	wire w_dff_B_gMAT52TG0_1;
	wire w_dff_B_kBn5VUQX0_0;
	wire w_dff_A_xsODTihY7_2;
	wire w_dff_A_k2sYJBL53_2;
	wire w_dff_A_xz3I73mA6_2;
	wire w_dff_A_g5l9RMl53_0;
	wire w_dff_A_y8KyCeV62_0;
	wire w_dff_A_ifxEZZu00_0;
	wire w_dff_A_SBY2aqI75_0;
	wire w_dff_A_awOn1qiS3_0;
	wire w_dff_A_PzVgNCOy3_2;
	wire w_dff_A_kj68dVfq5_2;
	wire w_dff_A_BI0MT9n17_2;
	wire w_dff_A_45F2Wfbn4_2;
	wire w_dff_A_IBdGzWN69_2;
	wire w_dff_A_bOqX34r50_1;
	wire w_dff_A_nRDA2vYG6_0;
	wire w_dff_A_Mym3gcbE7_0;
	wire w_dff_A_gRCIq3DY7_0;
	wire w_dff_A_tfc7ibsH7_0;
	wire w_dff_A_pNPAEwfB1_0;
	wire w_dff_A_H3vghLHm2_0;
	wire w_dff_A_XkM3NqXz1_0;
	wire w_dff_A_UTLB9La62_0;
	wire w_dff_A_nvOZlLyp4_0;
	wire w_dff_A_eKpGKkJK3_0;
	wire w_dff_A_iq1FECP85_0;
	wire w_dff_A_LLwYrFqp7_0;
	wire w_dff_A_VMHuDbXW2_0;
	wire w_dff_A_6k0ZNcJS5_0;
	wire w_dff_A_MY4xu2Sr4_0;
	wire w_dff_A_d58reL1z1_0;
	wire w_dff_A_57UHzbkQ8_0;
	wire w_dff_A_817YCMfQ3_0;
	wire w_dff_A_IG27HCOo2_0;
	wire w_dff_A_p8E3sw4r8_0;
	wire w_dff_A_tEUrMgvT0_0;
	wire w_dff_A_D3IYoDKs3_0;
	wire w_dff_A_wHstNy2b2_1;
	wire w_dff_A_5WUuWzmE9_2;
	wire w_dff_A_aMsv7RJo4_0;
	wire w_dff_A_fqzMkq1x0_0;
	wire w_dff_A_mnjIAAwl1_0;
	wire w_dff_A_Q0rJsq7D2_0;
	wire w_dff_A_zwJqievP9_0;
	wire w_dff_A_8rcd7bQa7_0;
	wire w_dff_A_nXwlvstj8_0;
	wire w_dff_A_HLWbYNWE0_0;
	wire w_dff_A_FSgxPSWq7_0;
	wire w_dff_A_JCZNzEoJ9_0;
	wire w_dff_A_UcmzbQkh5_0;
	wire w_dff_A_B88P9Sez4_0;
	wire w_dff_A_FnxcZ3DO9_0;
	wire w_dff_A_46g3VgXk0_0;
	wire w_dff_A_e3Uxfk0L0_0;
	wire w_dff_A_D6pRyXT40_0;
	wire w_dff_A_AiXwK1vd9_0;
	wire w_dff_A_z5VEzgME0_0;
	wire w_dff_A_5sV6vwcA1_0;
	wire w_dff_A_8Uo2JvBy7_0;
	wire w_dff_A_sADhmOWS6_0;
	wire w_dff_A_l9rnSSI04_0;
	wire w_dff_B_HSHaE9Ih2_2;
	wire w_dff_B_XNRly9na4_2;
	wire w_dff_B_nHxscb9U4_2;
	wire w_dff_A_y1RUfWp32_0;
	wire w_dff_A_j7cpPJAr6_0;
	wire w_dff_A_YIskqoSz7_0;
	wire w_dff_A_mmKCDQrv0_0;
	wire w_dff_A_QkSzTCdN3_0;
	wire w_dff_A_M1aNCpEq0_2;
	wire w_dff_A_xxP5WCIH0_2;
	wire w_dff_A_5wqRAZPE4_2;
	wire w_dff_A_3ECLkrun6_2;
	wire w_dff_A_JKedJh0d4_2;
	wire w_dff_A_GSwAHdKK6_1;
	wire w_dff_A_ddD5a0Aw5_0;
	wire w_dff_A_hvyyoF785_0;
	wire w_dff_A_vOxg2hAo2_0;
	wire w_dff_A_ptyxYr8f2_0;
	wire w_dff_A_BSBT0qQK9_0;
	wire w_dff_A_7QY9nNvq6_0;
	wire w_dff_A_np3P7awH0_0;
	wire w_dff_A_gixtXHhu8_0;
	wire w_dff_A_16IA2rWe6_0;
	wire w_dff_A_XwxqnrD51_0;
	wire w_dff_A_rrqo86Nk9_0;
	wire w_dff_A_5ZT7LSoQ0_0;
	wire w_dff_A_bTiiKfGM2_0;
	wire w_dff_A_fZCFhG694_0;
	wire w_dff_A_sNfeIk8T6_0;
	wire w_dff_A_d1EHCy0X4_0;
	wire w_dff_A_7ulYWxJU5_0;
	wire w_dff_A_sRQ6aVyO3_0;
	wire w_dff_A_fDNR9epd3_0;
	wire w_dff_A_wBEH4Wj33_0;
	wire w_dff_A_DeyXqbRp9_0;
	wire w_dff_A_4US1ySSH8_0;
	wire w_dff_A_lnIce6xP3_0;
	wire w_dff_A_sic6zVz01_0;
	wire w_dff_A_rwoTpeUC7_0;
	wire w_dff_A_ZGUuCZRu1_0;
	wire w_dff_A_uamd48YW7_0;
	wire w_dff_A_8UeOxRJh2_0;
	wire w_dff_A_LNp6Muz40_0;
	wire w_dff_A_s02xCIfa1_0;
	wire w_dff_A_TKIVSopJ8_0;
	wire w_dff_A_U2BrVfOt1_0;
	wire w_dff_A_Q9CXhgde5_0;
	wire w_dff_A_53kmCpTX7_0;
	wire w_dff_A_hyBkMIIC4_0;
	wire w_dff_A_wiS5E5NZ3_0;
	wire w_dff_A_85Ht0P2y9_0;
	wire w_dff_A_rdvvKlaS2_0;
	wire w_dff_A_EDDOjM8Z0_0;
	wire w_dff_A_vDLbXTvY4_0;
	wire w_dff_A_qmiZIMVd8_0;
	wire w_dff_A_nv0TeVXs4_0;
	wire w_dff_A_8e3J57y30_0;
	wire w_dff_A_axs5ry7q1_0;
	wire w_dff_A_x43OYFnI8_0;
	wire w_dff_A_9WX8LZch9_0;
	wire w_dff_A_vkyOKHke5_0;
	wire w_dff_A_2NzI4PPC1_0;
	wire w_dff_A_W5cq667D0_0;
	wire w_dff_A_QDoA0WXj3_0;
	wire w_dff_A_bJzb9TiQ3_0;
	wire w_dff_A_KiDbmSMU7_0;
	wire w_dff_A_IRWXDphX8_0;
	wire w_dff_A_Rv7Ika1y6_0;
	wire w_dff_A_RaPgyqEB0_0;
	wire w_dff_A_8UClQlks9_0;
	wire w_dff_A_aDxvsTPX7_0;
	wire w_dff_A_oFeujOQt1_0;
	wire w_dff_A_10V6IQla6_0;
	wire w_dff_A_76AAjDM61_0;
	wire w_dff_A_4OFky0sv7_0;
	wire w_dff_A_DrSqs3n32_0;
	wire w_dff_A_AjUdYfVM5_0;
	wire w_dff_A_4tQryBox6_0;
	wire w_dff_A_zRUc7yJH0_0;
	wire w_dff_A_NpQuwQpU9_0;
	wire w_dff_A_0kag68kR1_0;
	wire w_dff_A_zjPOeu2C6_0;
	wire w_dff_A_Bc0fjxVV8_0;
	wire w_dff_A_VWomtTTY1_0;
	wire w_dff_A_RgvbKDty8_0;
	wire w_dff_A_EH6tmStE3_0;
	wire w_dff_A_2WpoxvPT7_0;
	wire w_dff_A_F3OywF0E2_0;
	wire w_dff_A_ZYFOHQcy8_0;
	wire w_dff_A_lVVieE0z3_0;
	wire w_dff_A_vfHsKIz05_0;
	wire w_dff_A_tUPJ8xBQ2_0;
	wire w_dff_A_qJpb2hhC9_0;
	wire w_dff_A_mZlViL2C3_0;
	wire w_dff_A_dIzhVf4v7_0;
	wire w_dff_A_JhQ1WFom2_0;
	wire w_dff_A_HrFpJHTX4_0;
	wire w_dff_A_i1uTj3yO9_0;
	wire w_dff_A_Kdk8Zcjt9_0;
	wire w_dff_A_zsblTJ4d8_0;
	wire w_dff_A_dU3kP5r20_0;
	wire w_dff_A_yreAeIPE7_0;
	wire w_dff_A_gx2kTY761_1;
	wire w_dff_A_KvbXou8D0_0;
	wire w_dff_A_RvvEEplq5_0;
	wire w_dff_A_RSoabOWz8_0;
	wire w_dff_A_A6blB7S96_0;
	wire w_dff_A_zNJAKhRu8_0;
	wire w_dff_A_ef7t8ovF2_0;
	wire w_dff_A_6EwLDQLU9_0;
	wire w_dff_A_GOkfIyGo4_0;
	wire w_dff_A_Pu10F1fI7_0;
	wire w_dff_A_VpVb5lPW9_0;
	wire w_dff_A_RNbr4DrG7_0;
	wire w_dff_A_Uvq2ISC13_0;
	wire w_dff_A_7NHM8MYj7_0;
	wire w_dff_A_2B33gQmD1_0;
	wire w_dff_A_VU7Wfq9c0_0;
	wire w_dff_A_E64gVZvF1_0;
	wire w_dff_A_oTj1Gib57_0;
	wire w_dff_A_3QTYpOlI5_0;
	wire w_dff_A_InFSudi49_0;
	wire w_dff_A_cckRExhv2_0;
	wire w_dff_A_FDtq2BbX6_0;
	wire w_dff_A_9ZJCqNHa9_0;
	wire w_dff_A_xLHFZHh25_0;
	wire w_dff_A_jH5hUEm57_0;
	wire w_dff_A_k2y2WbVO4_0;
	wire w_dff_A_KPvoMPps7_0;
	wire w_dff_A_zoXmEvjH7_0;
	wire w_dff_A_I9ltBUix1_0;
	wire w_dff_A_8rerxCpB2_0;
	wire w_dff_A_zOoOuxQo5_0;
	wire w_dff_A_dyUIIFQ78_0;
	wire w_dff_A_NW3saaZP9_0;
	wire w_dff_A_WzdV4eai8_0;
	wire w_dff_A_e4m04q3B9_0;
	wire w_dff_A_aJENA3Po1_0;
	wire w_dff_A_CnrwW58Q0_0;
	wire w_dff_A_aITPlvab5_0;
	wire w_dff_A_1UeYkWGW6_0;
	wire w_dff_A_mnYtbXEY3_0;
	wire w_dff_A_AfU7IXd18_0;
	wire w_dff_A_57nUM4lY3_0;
	wire w_dff_A_7qUonzYj2_0;
	wire w_dff_A_JAcdjA6v9_0;
	wire w_dff_A_DGF6gZJt9_0;
	wire w_dff_A_iWPGaqeT9_0;
	wire w_dff_A_tHhgsdKJ8_0;
	wire w_dff_A_XLpT9dqa2_0;
	wire w_dff_A_j4B1sx2o1_0;
	wire w_dff_A_AbQnepcZ1_0;
	wire w_dff_A_k9osiVcG7_0;
	wire w_dff_A_VFCyZIEE9_0;
	wire w_dff_A_QFLZhNPM4_0;
	wire w_dff_A_h6RqiRQ63_0;
	wire w_dff_A_tPOqLmLd3_0;
	wire w_dff_A_tVGFvDGq0_0;
	wire w_dff_A_V7659hYV8_0;
	wire w_dff_A_904aWuNT2_0;
	wire w_dff_A_dkWeLLyS6_0;
	wire w_dff_A_t7yj3dmV4_0;
	wire w_dff_A_tKFWOP2H5_0;
	wire w_dff_A_TcfeqVxa7_0;
	wire w_dff_A_0nMjYDmr2_0;
	wire w_dff_A_zret7jSo2_0;
	wire w_dff_A_YIBYXjAd8_0;
	wire w_dff_A_J88dYbRL2_0;
	wire w_dff_A_7v7dT4Ll9_0;
	wire w_dff_A_KjBgybxO9_0;
	wire w_dff_A_luIVE5603_0;
	wire w_dff_A_rTeWKTuK5_0;
	wire w_dff_A_UqGw2XlN2_0;
	wire w_dff_A_CENrdQJ84_0;
	wire w_dff_A_PmM4NndX9_0;
	wire w_dff_A_RHrH6hO82_0;
	wire w_dff_A_fue47tCg2_0;
	wire w_dff_A_8NznfdDM5_0;
	wire w_dff_A_CuWHA5Yp4_0;
	wire w_dff_A_M6HBiUCH5_0;
	wire w_dff_A_oJO62Rp16_0;
	wire w_dff_A_z7UbHL3d5_0;
	wire w_dff_A_1aYYLMj23_0;
	wire w_dff_A_ZyrqKgsj1_0;
	wire w_dff_A_Z1jwAMuK9_0;
	wire w_dff_A_tPPdVKKG0_0;
	wire w_dff_A_sfJWps624_0;
	wire w_dff_A_EJdh07eS4_0;
	wire w_dff_A_cJdhGI191_0;
	wire w_dff_A_ocWcBmRt3_0;
	wire w_dff_A_ZQIL4zOV3_0;
	wire w_dff_A_TnMHhmql2_1;
	wire w_dff_A_CxeUrvIJ4_1;
	wire w_dff_A_JCTjOkmL1_1;
	wire w_dff_A_PrT1bVMz2_1;
	wire w_dff_A_oKvAYkiG8_1;
	wire w_dff_A_DSe6qKbN2_2;
	wire w_dff_A_lkQsU6Fo1_2;
	wire w_dff_A_hFQ7RFzM3_2;
	wire w_dff_A_TYAYYZlu6_2;
	wire w_dff_A_oeYXzT0W7_2;
	wire w_dff_A_XXy1jOTI2_1;
	wire w_dff_A_JWYMyi2G2_0;
	wire w_dff_A_YhzLEPzi5_0;
	wire w_dff_A_laAcwvOq2_0;
	wire w_dff_A_HfW89dTG3_0;
	wire w_dff_A_uloYN7lo4_0;
	wire w_dff_A_Z1pFR60o7_0;
	wire w_dff_A_gOBFhiLk5_0;
	wire w_dff_A_Tih0hyYL3_0;
	wire w_dff_A_YgeUGz0u3_0;
	wire w_dff_A_952dId8H4_0;
	wire w_dff_A_drLvg0bw5_0;
	wire w_dff_A_8NgL0byW5_0;
	wire w_dff_A_jhBVRKmS9_0;
	wire w_dff_A_ajgQ6ECf4_0;
	wire w_dff_A_M3mEFDcA5_0;
	wire w_dff_A_xjhhtLpD2_0;
	wire w_dff_A_lgbpSjju5_0;
	wire w_dff_A_Xf7ek1yO6_0;
	wire w_dff_A_ZBlzI3ey8_0;
	wire w_dff_A_8fY33f0s7_0;
	wire w_dff_A_eBECbbOr7_0;
	wire w_dff_A_OB7GilfJ9_0;
	wire w_dff_A_PifLK1KF9_0;
	wire w_dff_A_lN9CVWBF2_0;
	wire w_dff_A_zcT3cTsb7_0;
	wire w_dff_A_E5vlx3Ay8_0;
	wire w_dff_A_c1PhGR751_0;
	wire w_dff_A_9QnLx7LZ2_0;
	wire w_dff_A_XFIyex0l2_0;
	wire w_dff_A_OGklGDSh0_0;
	wire w_dff_A_n8FL9cNI3_0;
	wire w_dff_A_Cry3SQuq9_0;
	wire w_dff_A_6CKFAuNy6_0;
	wire w_dff_A_tKZgqRDz6_0;
	wire w_dff_A_Hr4RJzin2_0;
	wire w_dff_A_jkxtHo3y3_0;
	wire w_dff_A_EagGbAgF2_0;
	wire w_dff_A_dBIHdzLw4_0;
	wire w_dff_A_mvr7PKmQ0_0;
	wire w_dff_A_vEymCU7L9_0;
	wire w_dff_A_iVB6eI8q1_0;
	wire w_dff_A_rXxZgoZN9_0;
	wire w_dff_A_W5moqzen2_0;
	wire w_dff_A_EWk6wSym1_0;
	wire w_dff_A_oghYpZ7M3_0;
	wire w_dff_A_4xUDPzTL8_0;
	wire w_dff_A_N5jH4jXA9_0;
	wire w_dff_A_N5Ot1bJF0_0;
	wire w_dff_A_33XygtPg9_0;
	wire w_dff_A_e6HsgDU97_0;
	wire w_dff_A_5qgA06l26_0;
	wire w_dff_A_4iVMijiM8_0;
	wire w_dff_A_8jt1bLpO0_0;
	wire w_dff_A_1WTtnRBD1_0;
	wire w_dff_A_fOGk2Zs59_0;
	wire w_dff_A_Pxm2Hynp3_0;
	wire w_dff_A_KIflMu126_0;
	wire w_dff_A_9WyYmbh25_0;
	wire w_dff_A_VJFhodmT2_0;
	wire w_dff_A_5cf0d9z87_0;
	wire w_dff_A_v9i7mDaN7_0;
	wire w_dff_A_7cCj6nXZ7_0;
	wire w_dff_A_yQ2U1kXz8_0;
	wire w_dff_A_Z5xDBAup9_0;
	wire w_dff_A_9v7HP2XB4_0;
	wire w_dff_A_ScOY6LQa6_0;
	wire w_dff_A_ptDHawF33_0;
	wire w_dff_A_LlqxGvMB3_0;
	wire w_dff_A_3bjSki6M1_0;
	wire w_dff_A_XMDCLix27_0;
	wire w_dff_A_0nrKv9xc9_0;
	wire w_dff_A_CqkDwW2h5_0;
	wire w_dff_A_avvZpOWE5_0;
	wire w_dff_A_AurYlREi0_0;
	wire w_dff_A_qcu5Rdl66_0;
	wire w_dff_A_iHtSzie08_0;
	wire w_dff_A_1TLSdQqz3_0;
	wire w_dff_A_qbVd0D6m1_0;
	wire w_dff_A_ekdPj6c14_0;
	wire w_dff_A_Qs8IxPQU4_0;
	wire w_dff_A_zG7HLKGw9_0;
	wire w_dff_A_JAZzS8LO5_0;
	wire w_dff_A_aRgEUGVX7_0;
	wire w_dff_A_MWMyUdxS1_0;
	wire w_dff_A_asTS1FeR3_0;
	wire w_dff_A_wxeVzPs08_0;
	wire w_dff_A_7rpyD8io6_0;
	wire w_dff_A_qsVz5g8R4_0;
	wire w_dff_A_8SAwAT9O2_0;
	wire w_dff_A_VWJb7aaj1_0;
	wire w_dff_A_uYZ9ddvD0_0;
	wire w_dff_A_lH4RvTb54_0;
	wire w_dff_A_5PlTz9Gj5_0;
	wire w_dff_A_7OnIDFpU2_0;
	wire w_dff_A_6iyMxZ369_0;
	wire w_dff_A_0Hk51g9W6_0;
	wire w_dff_A_XylOKzOO5_0;
	wire w_dff_A_9kXPIB2g0_0;
	wire w_dff_A_M94Wx5ES3_0;
	wire w_dff_A_6FqbQmRT9_0;
	wire w_dff_A_moTWRqlj4_0;
	wire w_dff_A_ydDsvXT58_0;
	wire w_dff_A_d7lTRz1w1_0;
	wire w_dff_A_S6I0eFoT7_0;
	wire w_dff_A_6S06bhx94_0;
	wire w_dff_A_o1QY7sx44_0;
	wire w_dff_A_XtmNMhD51_0;
	wire w_dff_A_nQYkzxOf3_0;
	wire w_dff_A_IjZ9WPvP0_0;
	wire w_dff_A_vKv8bSYv9_0;
	wire w_dff_A_deLr8FPU4_0;
	wire w_dff_A_wxcsNfRJ6_0;
	wire w_dff_A_Ckrg3HfM2_0;
	wire w_dff_A_3tq7bs351_0;
	wire w_dff_A_m43anPMI1_0;
	wire w_dff_A_YT6aLnYY2_0;
	wire w_dff_A_pkKkitfx9_0;
	wire w_dff_A_iIiGKZl39_0;
	wire w_dff_A_F1eypsoi6_0;
	wire w_dff_A_sRof27eR9_0;
	wire w_dff_A_jkYTbfyn8_0;
	wire w_dff_A_FapeOVY95_0;
	wire w_dff_A_uK1a1sii7_0;
	wire w_dff_A_FqwzPC3E8_0;
	wire w_dff_A_WtTdz0lC0_0;
	wire w_dff_A_PxWIvayd9_0;
	wire w_dff_A_HIZilLLr7_0;
	wire w_dff_A_metjIlrp0_0;
	wire w_dff_A_fMsTXQ4I3_0;
	wire w_dff_A_zZHpXqXw9_0;
	wire w_dff_A_ioNA677y0_0;
	wire w_dff_A_KQTvHfr49_0;
	jxor g000(.dina(w_G85gat_0[2]),.dinb(w_G57gat_0[2]),.dout(n73),.clk(gclk));
	jxor g001(.dina(w_G29gat_0[2]),.dinb(w_G1gat_0[2]),.dout(n74),.clk(gclk));
	jxor g002(.dina(n74),.dinb(n73),.dout(n75),.clk(gclk));
	jxor g003(.dina(w_G162gat_0[2]),.dinb(w_G155gat_0[2]),.dout(n76),.clk(gclk));
	jxor g004(.dina(w_G148gat_0[2]),.dinb(w_G141gat_0[2]),.dout(n77),.clk(gclk));
	jxor g005(.dina(n77),.dinb(n76),.dout(n78),.clk(gclk));
	jxor g006(.dina(w_n78_0[1]),.dinb(n75),.dout(n79),.clk(gclk));
	jand g007(.dina(w_G233gat_1[2]),.dinb(G225gat),.dout(n80),.clk(gclk));
	jnot g008(.din(n80),.dout(n81),.clk(gclk));
	jxor g009(.dina(w_G134gat_0[2]),.dinb(w_G127gat_0[2]),.dout(n82),.clk(gclk));
	jxor g010(.dina(w_G120gat_0[2]),.dinb(w_G113gat_0[2]),.dout(n83),.clk(gclk));
	jxor g011(.dina(n83),.dinb(n82),.dout(n84),.clk(gclk));
	jxor g012(.dina(w_n84_0[1]),.dinb(n81),.dout(n85),.clk(gclk));
	jxor g013(.dina(n85),.dinb(n79),.dout(n86),.clk(gclk));
	jnot g014(.din(w_n86_1[1]),.dout(n87),.clk(gclk));
	jxor g015(.dina(w_G218gat_0[2]),.dinb(w_G190gat_0[2]),.dout(n88),.clk(gclk));
	jxor g016(.dina(w_G162gat_0[1]),.dinb(w_G134gat_0[1]),.dout(n89),.clk(gclk));
	jxor g017(.dina(n89),.dinb(n88),.dout(n90),.clk(gclk));
	jxor g018(.dina(w_G106gat_0[2]),.dinb(w_G99gat_0[2]),.dout(n91),.clk(gclk));
	jxor g019(.dina(w_G92gat_0[2]),.dinb(w_G85gat_0[1]),.dout(n92),.clk(gclk));
	jxor g020(.dina(n92),.dinb(n91),.dout(n93),.clk(gclk));
	jxor g021(.dina(w_n93_0[1]),.dinb(n90),.dout(n94),.clk(gclk));
	jnot g022(.din(G232gat),.dout(n95),.clk(gclk));
	jnot g023(.din(w_G233gat_1[1]),.dout(n96),.clk(gclk));
	jor g024(.dina(w_n96_1[1]),.dinb(n95),.dout(n97),.clk(gclk));
	jxor g025(.dina(w_G50gat_0[2]),.dinb(w_G43gat_0[2]),.dout(n98),.clk(gclk));
	jxor g026(.dina(w_G36gat_0[2]),.dinb(w_G29gat_0[1]),.dout(n99),.clk(gclk));
	jxor g027(.dina(n99),.dinb(n98),.dout(n100),.clk(gclk));
	jxor g028(.dina(w_n100_0[1]),.dinb(n97),.dout(n101),.clk(gclk));
	jxor g029(.dina(n101),.dinb(n94),.dout(n102),.clk(gclk));
	jxor g030(.dina(w_G211gat_0[2]),.dinb(w_G183gat_0[2]),.dout(n103),.clk(gclk));
	jxor g031(.dina(w_G155gat_0[1]),.dinb(w_G127gat_0[1]),.dout(n104),.clk(gclk));
	jxor g032(.dina(n104),.dinb(n103),.dout(n105),.clk(gclk));
	jxor g033(.dina(w_G78gat_0[2]),.dinb(w_G71gat_0[2]),.dout(n106),.clk(gclk));
	jxor g034(.dina(w_G64gat_0[2]),.dinb(w_G57gat_0[1]),.dout(n107),.clk(gclk));
	jxor g035(.dina(n107),.dinb(n106),.dout(n108),.clk(gclk));
	jxor g036(.dina(w_n108_0[1]),.dinb(n105),.dout(n109),.clk(gclk));
	jnot g037(.din(G231gat),.dout(n110),.clk(gclk));
	jor g038(.dina(w_n96_1[0]),.dinb(n110),.dout(n111),.clk(gclk));
	jxor g039(.dina(w_G22gat_0[2]),.dinb(w_G15gat_0[2]),.dout(n112),.clk(gclk));
	jxor g040(.dina(w_G8gat_0[2]),.dinb(w_G1gat_0[1]),.dout(n113),.clk(gclk));
	jxor g041(.dina(n113),.dinb(n112),.dout(n114),.clk(gclk));
	jxor g042(.dina(w_n114_0[1]),.dinb(n111),.dout(n115),.clk(gclk));
	jxor g043(.dina(n115),.dinb(n109),.dout(n116),.clk(gclk));
	jnot g044(.din(w_n116_1[1]),.dout(n117),.clk(gclk));
	jand g045(.dina(w_n117_1[2]),.dinb(w_n102_1[1]),.dout(n118),.clk(gclk));
	jxor g046(.dina(w_G92gat_0[1]),.dinb(w_G64gat_0[1]),.dout(n119),.clk(gclk));
	jxor g047(.dina(w_G36gat_0[1]),.dinb(w_G8gat_0[1]),.dout(n120),.clk(gclk));
	jxor g048(.dina(n120),.dinb(n119),.dout(n121),.clk(gclk));
	jxor g049(.dina(w_G190gat_0[1]),.dinb(w_G183gat_0[1]),.dout(n122),.clk(gclk));
	jxor g050(.dina(w_G176gat_0[2]),.dinb(w_G169gat_0[2]),.dout(n123),.clk(gclk));
	jxor g051(.dina(n123),.dinb(n122),.dout(n124),.clk(gclk));
	jxor g052(.dina(w_n124_0[1]),.dinb(n121),.dout(n125),.clk(gclk));
	jand g053(.dina(w_G233gat_1[0]),.dinb(G226gat),.dout(n126),.clk(gclk));
	jnot g054(.din(n126),.dout(n127),.clk(gclk));
	jxor g055(.dina(w_G218gat_0[1]),.dinb(w_G211gat_0[1]),.dout(n128),.clk(gclk));
	jxor g056(.dina(w_G204gat_0[2]),.dinb(w_G197gat_0[2]),.dout(n129),.clk(gclk));
	jxor g057(.dina(n129),.dinb(n128),.dout(n130),.clk(gclk));
	jxor g058(.dina(w_n130_0[1]),.dinb(n127),.dout(n131),.clk(gclk));
	jxor g059(.dina(n131),.dinb(n125),.dout(n132),.clk(gclk));
	jxor g060(.dina(w_n132_1[1]),.dinb(w_n86_1[0]),.dout(n133),.clk(gclk));
	jxor g061(.dina(w_G99gat_0[1]),.dinb(w_G71gat_0[1]),.dout(n134),.clk(gclk));
	jxor g062(.dina(w_G43gat_0[1]),.dinb(w_G15gat_0[1]),.dout(n135),.clk(gclk));
	jxor g063(.dina(n135),.dinb(n134),.dout(n136),.clk(gclk));
	jxor g064(.dina(n136),.dinb(w_n124_0[0]),.dout(n137),.clk(gclk));
	jnot g065(.din(G227gat),.dout(n138),.clk(gclk));
	jor g066(.dina(w_n96_0[2]),.dinb(n138),.dout(n139),.clk(gclk));
	jxor g067(.dina(n139),.dinb(w_n84_0[0]),.dout(n140),.clk(gclk));
	jxor g068(.dina(n140),.dinb(n137),.dout(n141),.clk(gclk));
	jxor g069(.dina(w_G106gat_0[1]),.dinb(w_G78gat_0[1]),.dout(n142),.clk(gclk));
	jxor g070(.dina(w_G50gat_0[1]),.dinb(w_G22gat_0[1]),.dout(n143),.clk(gclk));
	jxor g071(.dina(n143),.dinb(n142),.dout(n144),.clk(gclk));
	jxor g072(.dina(n144),.dinb(w_n130_0[0]),.dout(n145),.clk(gclk));
	jnot g073(.din(G228gat),.dout(n146),.clk(gclk));
	jor g074(.dina(w_n96_0[1]),.dinb(n146),.dout(n147),.clk(gclk));
	jxor g075(.dina(n147),.dinb(w_n78_0[0]),.dout(n148),.clk(gclk));
	jxor g076(.dina(n148),.dinb(n145),.dout(n149),.clk(gclk));
	jand g077(.dina(w_n149_1[1]),.dinb(w_n141_1[1]),.dout(n150),.clk(gclk));
	jand g078(.dina(n150),.dinb(n133),.dout(n151),.clk(gclk));
	jxor g079(.dina(w_n149_1[0]),.dinb(w_n141_1[0]),.dout(n152),.clk(gclk));
	jand g080(.dina(n152),.dinb(w_n86_0[2]),.dout(n153),.clk(gclk));
	jand g081(.dina(n153),.dinb(w_n132_1[0]),.dout(n154),.clk(gclk));
	jor g082(.dina(n154),.dinb(w_dff_B_IfNW47ib0_1),.dout(n155),.clk(gclk));
	jxor g083(.dina(w_G197gat_0[1]),.dinb(w_G169gat_0[1]),.dout(n156),.clk(gclk));
	jxor g084(.dina(w_G141gat_0[1]),.dinb(w_G113gat_0[1]),.dout(n157),.clk(gclk));
	jxor g085(.dina(n157),.dinb(n156),.dout(n158),.clk(gclk));
	jxor g086(.dina(n158),.dinb(w_n114_0[0]),.dout(n159),.clk(gclk));
	jand g087(.dina(w_G233gat_0[2]),.dinb(G229gat),.dout(n160),.clk(gclk));
	jnot g088(.din(n160),.dout(n161),.clk(gclk));
	jxor g089(.dina(n161),.dinb(w_n100_0[0]),.dout(n162),.clk(gclk));
	jxor g090(.dina(n162),.dinb(n159),.dout(n163),.clk(gclk));
	jnot g091(.din(w_n163_1[1]),.dout(n164),.clk(gclk));
	jxor g092(.dina(w_G204gat_0[1]),.dinb(w_G176gat_0[1]),.dout(n165),.clk(gclk));
	jxor g093(.dina(w_G148gat_0[1]),.dinb(w_G120gat_0[1]),.dout(n166),.clk(gclk));
	jxor g094(.dina(n166),.dinb(n165),.dout(n167),.clk(gclk));
	jxor g095(.dina(n167),.dinb(w_n108_0[0]),.dout(n168),.clk(gclk));
	jand g096(.dina(w_G233gat_0[1]),.dinb(G230gat),.dout(n169),.clk(gclk));
	jnot g097(.din(n169),.dout(n170),.clk(gclk));
	jxor g098(.dina(n170),.dinb(w_n93_0[0]),.dout(n171),.clk(gclk));
	jxor g099(.dina(n171),.dinb(n168),.dout(n172),.clk(gclk));
	jand g100(.dina(w_n172_1[1]),.dinb(w_n164_1[2]),.dout(n173),.clk(gclk));
	jand g101(.dina(w_n173_0[1]),.dinb(w_n155_0[2]),.dout(n174),.clk(gclk));
	jand g102(.dina(n174),.dinb(w_n118_0[1]),.dout(n175),.clk(gclk));
	jand g103(.dina(w_n175_1[1]),.dinb(w_n87_1[2]),.dout(n176),.clk(gclk));
	jxor g104(.dina(n176),.dinb(w_G1gat_0[0]),.dout(G1324gat),.clk(gclk));
	jnot g105(.din(w_n132_0[2]),.dout(n178),.clk(gclk));
	jand g106(.dina(w_n175_1[0]),.dinb(w_n178_1[2]),.dout(n179),.clk(gclk));
	jxor g107(.dina(n179),.dinb(w_G8gat_0[0]),.dout(G1325gat),.clk(gclk));
	jnot g108(.din(w_n141_0[2]),.dout(n181),.clk(gclk));
	jand g109(.dina(w_n175_0[2]),.dinb(w_n181_1[2]),.dout(n182),.clk(gclk));
	jxor g110(.dina(n182),.dinb(w_G15gat_0[0]),.dout(G1326gat),.clk(gclk));
	jnot g111(.din(w_n149_0[2]),.dout(n184),.clk(gclk));
	jand g112(.dina(w_n175_0[1]),.dinb(w_n184_1[2]),.dout(n185),.clk(gclk));
	jxor g113(.dina(n185),.dinb(w_G22gat_0[0]),.dout(G1327gat),.clk(gclk));
	jnot g114(.din(w_n102_1[0]),.dout(n187),.clk(gclk));
	jand g115(.dina(w_n116_1[0]),.dinb(w_n187_1[2]),.dout(n188),.clk(gclk));
	jand g116(.dina(w_dff_B_qvVbhgQM2_0),.dinb(w_n155_0[1]),.dout(n189),.clk(gclk));
	jand g117(.dina(w_n189_0[1]),.dinb(w_n173_0[0]),.dout(n190),.clk(gclk));
	jand g118(.dina(w_n190_1[1]),.dinb(w_n87_1[1]),.dout(n191),.clk(gclk));
	jxor g119(.dina(n191),.dinb(w_G29gat_0[0]),.dout(G1328gat),.clk(gclk));
	jand g120(.dina(w_n190_1[0]),.dinb(w_n178_1[1]),.dout(n193),.clk(gclk));
	jxor g121(.dina(n193),.dinb(w_G36gat_0[0]),.dout(G1329gat),.clk(gclk));
	jand g122(.dina(w_n190_0[2]),.dinb(w_n181_1[1]),.dout(n195),.clk(gclk));
	jxor g123(.dina(n195),.dinb(w_G43gat_0[0]),.dout(G1330gat),.clk(gclk));
	jand g124(.dina(w_n190_0[1]),.dinb(w_n184_1[1]),.dout(n197),.clk(gclk));
	jxor g125(.dina(n197),.dinb(w_G50gat_0[0]),.dout(G1331gat),.clk(gclk));
	jnot g126(.din(w_n172_1[0]),.dout(n199),.clk(gclk));
	jand g127(.dina(w_n199_1[2]),.dinb(w_n163_1[0]),.dout(n200),.clk(gclk));
	jand g128(.dina(w_n155_0[0]),.dinb(w_n118_0[0]),.dout(n201),.clk(gclk));
	jand g129(.dina(n201),.dinb(w_n200_0[1]),.dout(n202),.clk(gclk));
	jand g130(.dina(w_n202_1[1]),.dinb(w_n87_1[0]),.dout(n203),.clk(gclk));
	jxor g131(.dina(n203),.dinb(w_G57gat_0[0]),.dout(G1332gat),.clk(gclk));
	jand g132(.dina(w_n202_1[0]),.dinb(w_n178_1[0]),.dout(n205),.clk(gclk));
	jxor g133(.dina(n205),.dinb(w_G64gat_0[0]),.dout(G1333gat),.clk(gclk));
	jand g134(.dina(w_n202_0[2]),.dinb(w_n181_1[0]),.dout(n207),.clk(gclk));
	jxor g135(.dina(n207),.dinb(w_G71gat_0[0]),.dout(G1334gat),.clk(gclk));
	jand g136(.dina(w_n202_0[1]),.dinb(w_n184_1[0]),.dout(n209),.clk(gclk));
	jxor g137(.dina(n209),.dinb(w_G78gat_0[0]),.dout(G1335gat),.clk(gclk));
	jand g138(.dina(w_n200_0[0]),.dinb(w_n189_0[0]),.dout(n211),.clk(gclk));
	jand g139(.dina(w_n211_1[1]),.dinb(w_n87_0[2]),.dout(n212),.clk(gclk));
	jxor g140(.dina(n212),.dinb(w_G85gat_0[0]),.dout(G1336gat),.clk(gclk));
	jand g141(.dina(w_n211_1[0]),.dinb(w_n178_0[2]),.dout(n214),.clk(gclk));
	jxor g142(.dina(n214),.dinb(w_G92gat_0[0]),.dout(G1337gat),.clk(gclk));
	jand g143(.dina(w_n211_0[2]),.dinb(w_n181_0[2]),.dout(n216),.clk(gclk));
	jxor g144(.dina(n216),.dinb(w_G99gat_0[0]),.dout(G1338gat),.clk(gclk));
	jand g145(.dina(w_n211_0[1]),.dinb(w_n184_0[2]),.dout(n218),.clk(gclk));
	jxor g146(.dina(n218),.dinb(w_G106gat_0[0]),.dout(G1339gat),.clk(gclk));
	jand g147(.dina(w_n149_0[1]),.dinb(w_n181_0[1]),.dout(n220),.clk(gclk));
	jand g148(.dina(w_n132_0[1]),.dinb(w_n87_0[1]),.dout(n221),.clk(gclk));
	jxor g149(.dina(w_n116_0[2]),.dinb(w_n102_0[2]),.dout(n222),.clk(gclk));
	jand g150(.dina(n222),.dinb(w_n163_0[2]),.dout(n223),.clk(gclk));
	jand g151(.dina(n223),.dinb(w_n172_0[2]),.dout(n224),.clk(gclk));
	jxor g152(.dina(w_n172_0[1]),.dinb(w_n163_0[1]),.dout(n225),.clk(gclk));
	jand g153(.dina(w_n116_0[1]),.dinb(w_n102_0[1]),.dout(n226),.clk(gclk));
	jand g154(.dina(n226),.dinb(n225),.dout(n227),.clk(gclk));
	jor g155(.dina(w_dff_B_kBn5VUQX0_0),.dinb(n224),.dout(n228),.clk(gclk));
	jand g156(.dina(w_n228_0[1]),.dinb(w_dff_B_X2Im87NO5_1),.dout(n229),.clk(gclk));
	jand g157(.dina(w_n229_0[1]),.dinb(w_n220_0[1]),.dout(n230),.clk(gclk));
	jand g158(.dina(w_n230_1[1]),.dinb(w_n164_1[1]),.dout(n231),.clk(gclk));
	jxor g159(.dina(n231),.dinb(w_G113gat_0[0]),.dout(G1340gat),.clk(gclk));
	jand g160(.dina(w_n230_1[0]),.dinb(w_n199_1[1]),.dout(n233),.clk(gclk));
	jxor g161(.dina(n233),.dinb(w_G120gat_0[0]),.dout(G1341gat),.clk(gclk));
	jand g162(.dina(w_n230_0[2]),.dinb(w_n117_1[1]),.dout(n235),.clk(gclk));
	jxor g163(.dina(n235),.dinb(w_G127gat_0[0]),.dout(G1342gat),.clk(gclk));
	jand g164(.dina(w_n230_0[1]),.dinb(w_n187_1[1]),.dout(n237),.clk(gclk));
	jxor g165(.dina(n237),.dinb(w_G134gat_0[0]),.dout(G1343gat),.clk(gclk));
	jand g166(.dina(w_n184_0[1]),.dinb(w_n141_0[1]),.dout(n239),.clk(gclk));
	jand g167(.dina(w_n229_0[0]),.dinb(w_n239_0[1]),.dout(n240),.clk(gclk));
	jand g168(.dina(w_n240_1[1]),.dinb(w_n164_1[0]),.dout(n241),.clk(gclk));
	jxor g169(.dina(n241),.dinb(w_G141gat_0[0]),.dout(G1344gat),.clk(gclk));
	jand g170(.dina(w_n240_1[0]),.dinb(w_n199_1[0]),.dout(n243),.clk(gclk));
	jxor g171(.dina(n243),.dinb(w_G148gat_0[0]),.dout(G1345gat),.clk(gclk));
	jand g172(.dina(w_n240_0[2]),.dinb(w_n117_1[0]),.dout(n245),.clk(gclk));
	jxor g173(.dina(n245),.dinb(w_G155gat_0[0]),.dout(G1346gat),.clk(gclk));
	jand g174(.dina(w_n240_0[1]),.dinb(w_n187_1[0]),.dout(n247),.clk(gclk));
	jxor g175(.dina(n247),.dinb(w_G162gat_0[0]),.dout(G1347gat),.clk(gclk));
	jand g176(.dina(w_n178_0[1]),.dinb(w_n86_0[1]),.dout(n249),.clk(gclk));
	jand g177(.dina(w_n228_0[0]),.dinb(w_dff_B_gMAT52TG0_1),.dout(n250),.clk(gclk));
	jand g178(.dina(w_n250_0[1]),.dinb(w_n220_0[0]),.dout(n251),.clk(gclk));
	jand g179(.dina(w_n251_1[1]),.dinb(w_n164_0[2]),.dout(n252),.clk(gclk));
	jxor g180(.dina(n252),.dinb(w_G169gat_0[0]),.dout(G1348gat),.clk(gclk));
	jand g181(.dina(w_n251_1[0]),.dinb(w_n199_0[2]),.dout(n254),.clk(gclk));
	jxor g182(.dina(n254),.dinb(w_G176gat_0[0]),.dout(G1349gat),.clk(gclk));
	jand g183(.dina(w_n251_0[2]),.dinb(w_n117_0[2]),.dout(n256),.clk(gclk));
	jxor g184(.dina(n256),.dinb(w_G183gat_0[0]),.dout(G1350gat),.clk(gclk));
	jand g185(.dina(w_n251_0[1]),.dinb(w_n187_0[2]),.dout(n258),.clk(gclk));
	jxor g186(.dina(n258),.dinb(w_G190gat_0[0]),.dout(G1351gat),.clk(gclk));
	jand g187(.dina(w_n250_0[0]),.dinb(w_n239_0[0]),.dout(n260),.clk(gclk));
	jand g188(.dina(w_n260_1[1]),.dinb(w_n164_0[1]),.dout(n261),.clk(gclk));
	jxor g189(.dina(n261),.dinb(w_G197gat_0[0]),.dout(G1352gat),.clk(gclk));
	jand g190(.dina(w_n260_1[0]),.dinb(w_n199_0[1]),.dout(n263),.clk(gclk));
	jxor g191(.dina(n263),.dinb(w_G204gat_0[0]),.dout(G1353gat),.clk(gclk));
	jand g192(.dina(w_n260_0[2]),.dinb(w_n117_0[1]),.dout(n265),.clk(gclk));
	jxor g193(.dina(n265),.dinb(w_G211gat_0[0]),.dout(G1354gat),.clk(gclk));
	jand g194(.dina(w_n260_0[1]),.dinb(w_n187_0[1]),.dout(n267),.clk(gclk));
	jxor g195(.dina(n267),.dinb(w_G218gat_0[0]),.dout(G1355gat),.clk(gclk));
	jspl3 jspl3_w_G1gat_0(.douta(w_dff_A_UcmzbQkh5_0),.doutb(w_G1gat_0[1]),.doutc(w_G1gat_0[2]),.din(G1gat));
	jspl3 jspl3_w_G8gat_0(.douta(w_dff_A_iq1FECP85_0),.doutb(w_G8gat_0[1]),.doutc(w_G8gat_0[2]),.din(G8gat));
	jspl3 jspl3_w_G15gat_0(.douta(w_dff_A_DGF6gZJt9_0),.doutb(w_G15gat_0[1]),.doutc(w_G15gat_0[2]),.din(G15gat));
	jspl3 jspl3_w_G22gat_0(.douta(w_dff_A_axs5ry7q1_0),.doutb(w_G22gat_0[1]),.doutc(w_G22gat_0[2]),.din(G22gat));
	jspl3 jspl3_w_G29gat_0(.douta(w_dff_A_OB7GilfJ9_0),.doutb(w_G29gat_0[1]),.doutc(w_G29gat_0[2]),.din(G29gat));
	jspl3 jspl3_w_G36gat_0(.douta(w_dff_A_drLvg0bw5_0),.doutb(w_G36gat_0[1]),.doutc(w_G36gat_0[2]),.din(G36gat));
	jspl3 jspl3_w_G43gat_0(.douta(w_dff_A_EWk6wSym1_0),.doutb(w_G43gat_0[1]),.doutc(w_G43gat_0[2]),.din(G43gat));
	jspl3 jspl3_w_G50gat_0(.douta(w_dff_A_6CKFAuNy6_0),.doutb(w_G50gat_0[1]),.doutc(w_G50gat_0[2]),.din(G50gat));
	jspl3 jspl3_w_G57gat_0(.douta(w_dff_A_l9rnSSI04_0),.doutb(w_G57gat_0[1]),.doutc(w_G57gat_0[2]),.din(G57gat));
	jspl3 jspl3_w_G64gat_0(.douta(w_dff_A_D3IYoDKs3_0),.doutb(w_G64gat_0[1]),.doutc(w_G64gat_0[2]),.din(G64gat));
	jspl3 jspl3_w_G71gat_0(.douta(w_dff_A_tVGFvDGq0_0),.doutb(w_G71gat_0[1]),.doutc(w_G71gat_0[2]),.din(G71gat));
	jspl3 jspl3_w_G78gat_0(.douta(w_dff_A_RaPgyqEB0_0),.doutb(w_G78gat_0[1]),.doutc(w_G78gat_0[2]),.din(G78gat));
	jspl3 jspl3_w_G85gat_0(.douta(w_dff_A_ScOY6LQa6_0),.doutb(w_G85gat_0[1]),.doutc(w_G85gat_0[2]),.din(G85gat));
	jspl3 jspl3_w_G92gat_0(.douta(w_dff_A_fOGk2Zs59_0),.doutb(w_G92gat_0[1]),.doutc(w_G92gat_0[2]),.din(G92gat));
	jspl3 jspl3_w_G99gat_0(.douta(w_dff_A_qsVz5g8R4_0),.doutb(w_G99gat_0[1]),.doutc(w_G99gat_0[2]),.din(G99gat));
	jspl3 jspl3_w_G106gat_0(.douta(w_dff_A_1TLSdQqz3_0),.doutb(w_G106gat_0[1]),.doutc(w_G106gat_0[2]),.din(G106gat));
	jspl3 jspl3_w_G113gat_0(.douta(w_dff_A_9ZJCqNHa9_0),.doutb(w_G113gat_0[1]),.doutc(w_G113gat_0[2]),.din(G113gat));
	jspl3 jspl3_w_G120gat_0(.douta(w_dff_A_RNbr4DrG7_0),.doutb(w_G120gat_0[1]),.doutc(w_G120gat_0[2]),.din(G120gat));
	jspl3 jspl3_w_G127gat_0(.douta(w_dff_A_WzdV4eai8_0),.doutb(w_G127gat_0[1]),.doutc(w_G127gat_0[2]),.din(G127gat));
	jspl3 jspl3_w_G134gat_0(.douta(w_dff_A_vKv8bSYv9_0),.doutb(w_G134gat_0[1]),.doutc(w_G134gat_0[2]),.din(G134gat));
	jspl3 jspl3_w_G141gat_0(.douta(w_dff_A_4US1ySSH8_0),.doutb(w_G141gat_0[1]),.doutc(w_G141gat_0[2]),.din(G141gat));
	jspl3 jspl3_w_G148gat_0(.douta(w_dff_A_rrqo86Nk9_0),.doutb(w_G148gat_0[1]),.doutc(w_G148gat_0[2]),.din(G148gat));
	jspl3 jspl3_w_G155gat_0(.douta(w_dff_A_Q9CXhgde5_0),.doutb(w_G155gat_0[1]),.doutc(w_G155gat_0[2]),.din(G155gat));
	jspl3 jspl3_w_G162gat_0(.douta(w_dff_A_M94Wx5ES3_0),.doutb(w_G162gat_0[1]),.doutc(w_G162gat_0[2]),.din(G162gat));
	jspl3 jspl3_w_G169gat_0(.douta(w_dff_A_M6HBiUCH5_0),.doutb(w_G169gat_0[1]),.doutc(w_G169gat_0[2]),.din(G169gat));
	jspl3 jspl3_w_G176gat_0(.douta(w_dff_A_7v7dT4Ll9_0),.doutb(w_G176gat_0[1]),.doutc(w_G176gat_0[2]),.din(G176gat));
	jspl3 jspl3_w_G183gat_0(.douta(w_dff_A_ZQIL4zOV3_0),.doutb(w_G183gat_0[1]),.doutc(w_G183gat_0[2]),.din(G183gat));
	jspl3 jspl3_w_G190gat_0(.douta(w_dff_A_KQTvHfr49_0),.doutb(w_G190gat_0[1]),.doutc(w_G190gat_0[2]),.din(G190gat));
	jspl3 jspl3_w_G197gat_0(.douta(w_dff_A_vfHsKIz05_0),.doutb(w_G197gat_0[1]),.doutc(w_G197gat_0[2]),.din(G197gat));
	jspl3 jspl3_w_G204gat_0(.douta(w_dff_A_NpQuwQpU9_0),.doutb(w_G204gat_0[1]),.doutc(w_G204gat_0[2]),.din(G204gat));
	jspl3 jspl3_w_G211gat_0(.douta(w_dff_A_yreAeIPE7_0),.doutb(w_G211gat_0[1]),.doutc(w_G211gat_0[2]),.din(G211gat));
	jspl3 jspl3_w_G218gat_0(.douta(w_dff_A_jkYTbfyn8_0),.doutb(w_G218gat_0[1]),.doutc(w_G218gat_0[2]),.din(G218gat));
	jspl3 jspl3_w_G233gat_0(.douta(w_G233gat_0[0]),.doutb(w_G233gat_0[1]),.doutc(w_G233gat_0[2]),.din(G233gat));
	jspl3 jspl3_w_G233gat_1(.douta(w_G233gat_1[0]),.doutb(w_G233gat_1[1]),.doutc(w_G233gat_1[2]),.din(w_G233gat_0[0]));
	jspl jspl_w_n78_0(.douta(w_n78_0[0]),.doutb(w_n78_0[1]),.din(n78));
	jspl jspl_w_n84_0(.douta(w_n84_0[0]),.doutb(w_n84_0[1]),.din(n84));
	jspl3 jspl3_w_n86_0(.douta(w_n86_0[0]),.doutb(w_dff_A_wHstNy2b2_1),.doutc(w_dff_A_5WUuWzmE9_2),.din(n86));
	jspl jspl_w_n86_1(.douta(w_n86_1[0]),.doutb(w_n86_1[1]),.din(w_n86_0[0]));
	jspl3 jspl3_w_n87_0(.douta(w_dff_A_HDvR5fGe3_0),.doutb(w_n87_0[1]),.doutc(w_dff_A_7DImgA5K9_2),.din(n87));
	jspl3 jspl3_w_n87_1(.douta(w_n87_1[0]),.doutb(w_n87_1[1]),.doutc(w_n87_1[2]),.din(w_n87_0[0]));
	jspl jspl_w_n93_0(.douta(w_n93_0[0]),.doutb(w_n93_0[1]),.din(n93));
	jspl3 jspl3_w_n96_0(.douta(w_n96_0[0]),.doutb(w_n96_0[1]),.doutc(w_n96_0[2]),.din(n96));
	jspl jspl_w_n96_1(.douta(w_n96_1[0]),.doutb(w_n96_1[1]),.din(w_n96_0[0]));
	jspl jspl_w_n100_0(.douta(w_n100_0[0]),.doutb(w_n100_0[1]),.din(n100));
	jspl3 jspl3_w_n102_0(.douta(w_n102_0[0]),.doutb(w_n102_0[1]),.doutc(w_n102_0[2]),.din(n102));
	jspl jspl_w_n102_1(.douta(w_n102_1[0]),.doutb(w_dff_A_XXy1jOTI2_1),.din(w_n102_0[0]));
	jspl jspl_w_n108_0(.douta(w_n108_0[0]),.doutb(w_n108_0[1]),.din(n108));
	jspl jspl_w_n114_0(.douta(w_n114_0[0]),.doutb(w_n114_0[1]),.din(n114));
	jspl3 jspl3_w_n116_0(.douta(w_n116_0[0]),.doutb(w_n116_0[1]),.doutc(w_n116_0[2]),.din(n116));
	jspl jspl_w_n116_1(.douta(w_dff_A_rIYE9OzL2_0),.doutb(w_n116_1[1]),.din(w_n116_0[0]));
	jspl3 jspl3_w_n117_0(.douta(w_n117_0[0]),.doutb(w_dff_A_C2tRsLlm2_1),.doutc(w_dff_A_6rL5Wax43_2),.din(n117));
	jspl3 jspl3_w_n117_1(.douta(w_dff_A_BvcpixTz4_0),.doutb(w_dff_A_ANbbw8Pr3_1),.doutc(w_n117_1[2]),.din(w_n117_0[0]));
	jspl jspl_w_n118_0(.douta(w_n118_0[0]),.doutb(w_dff_A_XFMs5PF89_1),.din(w_dff_B_cMdmeUqR9_2));
	jspl jspl_w_n124_0(.douta(w_n124_0[0]),.doutb(w_n124_0[1]),.din(n124));
	jspl jspl_w_n130_0(.douta(w_n130_0[0]),.doutb(w_n130_0[1]),.din(n130));
	jspl3 jspl3_w_n132_0(.douta(w_n132_0[0]),.doutb(w_dff_A_bOqX34r50_1),.doutc(w_n132_0[2]),.din(n132));
	jspl jspl_w_n132_1(.douta(w_dff_A_qvU4pT7M9_0),.doutb(w_n132_1[1]),.din(w_n132_0[0]));
	jspl3 jspl3_w_n141_0(.douta(w_n141_0[0]),.doutb(w_dff_A_gx2kTY761_1),.doutc(w_n141_0[2]),.din(n141));
	jspl jspl_w_n141_1(.douta(w_n141_1[0]),.doutb(w_n141_1[1]),.din(w_n141_0[0]));
	jspl3 jspl3_w_n149_0(.douta(w_n149_0[0]),.doutb(w_dff_A_GSwAHdKK6_1),.doutc(w_n149_0[2]),.din(n149));
	jspl jspl_w_n149_1(.douta(w_n149_1[0]),.doutb(w_n149_1[1]),.din(w_n149_0[0]));
	jspl3 jspl3_w_n155_0(.douta(w_n155_0[0]),.doutb(w_n155_0[1]),.doutc(w_n155_0[2]),.din(n155));
	jspl3 jspl3_w_n163_0(.douta(w_n163_0[0]),.doutb(w_n163_0[1]),.doutc(w_dff_A_xsODTihY7_2),.din(n163));
	jspl jspl_w_n163_1(.douta(w_dff_A_9woERz7Z9_0),.doutb(w_n163_1[1]),.din(w_n163_0[0]));
	jspl3 jspl3_w_n164_0(.douta(w_n164_0[0]),.doutb(w_dff_A_fiIPpVW66_1),.doutc(w_dff_A_neoNnWwU3_2),.din(n164));
	jspl3 jspl3_w_n164_1(.douta(w_dff_A_FZGlmU2N4_0),.doutb(w_dff_A_sFVdG6WN0_1),.doutc(w_n164_1[2]),.din(w_n164_0[0]));
	jspl3 jspl3_w_n172_0(.douta(w_n172_0[0]),.doutb(w_n172_0[1]),.doutc(w_dff_A_xz3I73mA6_2),.din(n172));
	jspl jspl_w_n172_1(.douta(w_n172_1[0]),.doutb(w_dff_A_Y51j7kVV7_1),.din(w_n172_0[0]));
	jspl jspl_w_n173_0(.douta(w_dff_A_g7fWtRC34_0),.doutb(w_n173_0[1]),.din(w_dff_B_XLzfbrYo1_2));
	jspl3 jspl3_w_n175_0(.douta(w_n175_0[0]),.doutb(w_n175_0[1]),.doutc(w_n175_0[2]),.din(n175));
	jspl jspl_w_n175_1(.douta(w_n175_1[0]),.doutb(w_n175_1[1]),.din(w_n175_0[0]));
	jspl3 jspl3_w_n178_0(.douta(w_dff_A_awOn1qiS3_0),.doutb(w_n178_0[1]),.doutc(w_dff_A_IBdGzWN69_2),.din(n178));
	jspl3 jspl3_w_n178_1(.douta(w_n178_1[0]),.doutb(w_n178_1[1]),.doutc(w_n178_1[2]),.din(w_n178_0[0]));
	jspl3 jspl3_w_n181_0(.douta(w_dff_A_Z09T7J496_0),.doutb(w_n181_0[1]),.doutc(w_dff_A_KepHnE5C4_2),.din(n181));
	jspl3 jspl3_w_n181_1(.douta(w_n181_1[0]),.doutb(w_n181_1[1]),.doutc(w_n181_1[2]),.din(w_n181_0[0]));
	jspl3 jspl3_w_n184_0(.douta(w_dff_A_QkSzTCdN3_0),.doutb(w_n184_0[1]),.doutc(w_dff_A_JKedJh0d4_2),.din(n184));
	jspl3 jspl3_w_n184_1(.douta(w_n184_1[0]),.doutb(w_n184_1[1]),.doutc(w_n184_1[2]),.din(w_n184_0[0]));
	jspl3 jspl3_w_n187_0(.douta(w_n187_0[0]),.doutb(w_dff_A_oKvAYkiG8_1),.doutc(w_dff_A_oeYXzT0W7_2),.din(n187));
	jspl3 jspl3_w_n187_1(.douta(w_dff_A_pFG4FcaY0_0),.doutb(w_dff_A_2DYJGpGs2_1),.doutc(w_n187_1[2]),.din(w_n187_0[0]));
	jspl jspl_w_n189_0(.douta(w_n189_0[0]),.doutb(w_n189_0[1]),.din(n189));
	jspl3 jspl3_w_n190_0(.douta(w_n190_0[0]),.doutb(w_n190_0[1]),.doutc(w_n190_0[2]),.din(n190));
	jspl jspl_w_n190_1(.douta(w_n190_1[0]),.doutb(w_n190_1[1]),.din(w_n190_0[0]));
	jspl3 jspl3_w_n199_0(.douta(w_n199_0[0]),.doutb(w_dff_A_Pt4jPtr59_1),.doutc(w_dff_A_dDSIcMPD8_2),.din(n199));
	jspl3 jspl3_w_n199_1(.douta(w_dff_A_iuTgCrL40_0),.doutb(w_dff_A_pFx1qlrF2_1),.doutc(w_n199_1[2]),.din(w_n199_0[0]));
	jspl jspl_w_n200_0(.douta(w_n200_0[0]),.doutb(w_n200_0[1]),.din(w_dff_B_ictF7VVB8_2));
	jspl3 jspl3_w_n202_0(.douta(w_n202_0[0]),.doutb(w_n202_0[1]),.doutc(w_n202_0[2]),.din(n202));
	jspl jspl_w_n202_1(.douta(w_n202_1[0]),.doutb(w_n202_1[1]),.din(w_n202_0[0]));
	jspl3 jspl3_w_n211_0(.douta(w_n211_0[0]),.doutb(w_n211_0[1]),.doutc(w_n211_0[2]),.din(n211));
	jspl jspl_w_n211_1(.douta(w_n211_1[0]),.doutb(w_n211_1[1]),.din(w_n211_0[0]));
	jspl jspl_w_n220_0(.douta(w_n220_0[0]),.doutb(w_n220_0[1]),.din(w_dff_B_ZnnCJ2u80_2));
	jspl jspl_w_n228_0(.douta(w_n228_0[0]),.doutb(w_n228_0[1]),.din(n228));
	jspl jspl_w_n229_0(.douta(w_n229_0[0]),.doutb(w_n229_0[1]),.din(n229));
	jspl3 jspl3_w_n230_0(.douta(w_n230_0[0]),.doutb(w_n230_0[1]),.doutc(w_n230_0[2]),.din(n230));
	jspl jspl_w_n230_1(.douta(w_n230_1[0]),.doutb(w_n230_1[1]),.din(w_n230_0[0]));
	jspl jspl_w_n239_0(.douta(w_n239_0[0]),.doutb(w_n239_0[1]),.din(w_dff_B_nHxscb9U4_2));
	jspl3 jspl3_w_n240_0(.douta(w_n240_0[0]),.doutb(w_n240_0[1]),.doutc(w_n240_0[2]),.din(n240));
	jspl jspl_w_n240_1(.douta(w_n240_1[0]),.doutb(w_n240_1[1]),.din(w_n240_0[0]));
	jspl jspl_w_n250_0(.douta(w_n250_0[0]),.doutb(w_n250_0[1]),.din(n250));
	jspl3 jspl3_w_n251_0(.douta(w_n251_0[0]),.doutb(w_n251_0[1]),.doutc(w_n251_0[2]),.din(n251));
	jspl jspl_w_n251_1(.douta(w_n251_1[0]),.doutb(w_n251_1[1]),.din(w_n251_0[0]));
	jspl3 jspl3_w_n260_0(.douta(w_n260_0[0]),.doutb(w_n260_0[1]),.doutc(w_n260_0[2]),.din(n260));
	jspl jspl_w_n260_1(.douta(w_n260_1[0]),.doutb(w_n260_1[1]),.din(w_n260_0[0]));
	jdff dff_A_g7fWtRC34_0(.dout(w_n173_0[0]),.din(w_dff_A_g7fWtRC34_0),.clk(gclk));
	jdff dff_B_UbdA9TpT0_2(.din(n173),.dout(w_dff_B_UbdA9TpT0_2),.clk(gclk));
	jdff dff_B_XLzfbrYo1_2(.din(w_dff_B_UbdA9TpT0_2),.dout(w_dff_B_XLzfbrYo1_2),.clk(gclk));
	jdff dff_A_XFMs5PF89_1(.dout(w_n118_0[1]),.din(w_dff_A_XFMs5PF89_1),.clk(gclk));
	jdff dff_B_C82Ol07Z2_2(.din(n118),.dout(w_dff_B_C82Ol07Z2_2),.clk(gclk));
	jdff dff_B_cMdmeUqR9_2(.din(w_dff_B_C82Ol07Z2_2),.dout(w_dff_B_cMdmeUqR9_2),.clk(gclk));
	jdff dff_B_oD2VeBYI1_2(.din(n200),.dout(w_dff_B_oD2VeBYI1_2),.clk(gclk));
	jdff dff_B_uXMssaTF3_2(.din(w_dff_B_oD2VeBYI1_2),.dout(w_dff_B_uXMssaTF3_2),.clk(gclk));
	jdff dff_B_ictF7VVB8_2(.din(w_dff_B_uXMssaTF3_2),.dout(w_dff_B_ictF7VVB8_2),.clk(gclk));
	jdff dff_B_fEXmCUEr6_0(.din(n188),.dout(w_dff_B_fEXmCUEr6_0),.clk(gclk));
	jdff dff_B_qvVbhgQM2_0(.din(w_dff_B_fEXmCUEr6_0),.dout(w_dff_B_qvVbhgQM2_0),.clk(gclk));
	jdff dff_B_IfNW47ib0_1(.din(n151),.dout(w_dff_B_IfNW47ib0_1),.clk(gclk));
	jdff dff_A_4kRfFieY2_0(.dout(w_n132_1[0]),.din(w_dff_A_4kRfFieY2_0),.clk(gclk));
	jdff dff_A_qvU4pT7M9_0(.dout(w_dff_A_4kRfFieY2_0),.din(w_dff_A_qvU4pT7M9_0),.clk(gclk));
	jdff dff_A_w5BUOEI76_0(.dout(w_n164_1[0]),.din(w_dff_A_w5BUOEI76_0),.clk(gclk));
	jdff dff_A_WOeCCUnT6_0(.dout(w_dff_A_w5BUOEI76_0),.din(w_dff_A_WOeCCUnT6_0),.clk(gclk));
	jdff dff_A_pjcl3KMO5_0(.dout(w_dff_A_WOeCCUnT6_0),.din(w_dff_A_pjcl3KMO5_0),.clk(gclk));
	jdff dff_A_bM5Ydb574_0(.dout(w_dff_A_pjcl3KMO5_0),.din(w_dff_A_bM5Ydb574_0),.clk(gclk));
	jdff dff_A_FZGlmU2N4_0(.dout(w_dff_A_bM5Ydb574_0),.din(w_dff_A_FZGlmU2N4_0),.clk(gclk));
	jdff dff_A_GY3GUQUV5_1(.dout(w_n164_1[1]),.din(w_dff_A_GY3GUQUV5_1),.clk(gclk));
	jdff dff_A_bbxDdLtV6_1(.dout(w_dff_A_GY3GUQUV5_1),.din(w_dff_A_bbxDdLtV6_1),.clk(gclk));
	jdff dff_A_a0vgmC6X2_1(.dout(w_dff_A_bbxDdLtV6_1),.din(w_dff_A_a0vgmC6X2_1),.clk(gclk));
	jdff dff_A_xdfdtWBd6_1(.dout(w_dff_A_a0vgmC6X2_1),.din(w_dff_A_xdfdtWBd6_1),.clk(gclk));
	jdff dff_A_sFVdG6WN0_1(.dout(w_dff_A_xdfdtWBd6_1),.din(w_dff_A_sFVdG6WN0_1),.clk(gclk));
	jdff dff_A_qJ5zHxs81_0(.dout(w_n199_1[0]),.din(w_dff_A_qJ5zHxs81_0),.clk(gclk));
	jdff dff_A_K1PQJV6P4_0(.dout(w_dff_A_qJ5zHxs81_0),.din(w_dff_A_K1PQJV6P4_0),.clk(gclk));
	jdff dff_A_Fo4NdyDl9_0(.dout(w_dff_A_K1PQJV6P4_0),.din(w_dff_A_Fo4NdyDl9_0),.clk(gclk));
	jdff dff_A_cNwRv10B6_0(.dout(w_dff_A_Fo4NdyDl9_0),.din(w_dff_A_cNwRv10B6_0),.clk(gclk));
	jdff dff_A_iuTgCrL40_0(.dout(w_dff_A_cNwRv10B6_0),.din(w_dff_A_iuTgCrL40_0),.clk(gclk));
	jdff dff_A_0mjTla9J4_1(.dout(w_n199_1[1]),.din(w_dff_A_0mjTla9J4_1),.clk(gclk));
	jdff dff_A_MkIJKXmu7_1(.dout(w_dff_A_0mjTla9J4_1),.din(w_dff_A_MkIJKXmu7_1),.clk(gclk));
	jdff dff_A_Br5tP2ke6_1(.dout(w_dff_A_MkIJKXmu7_1),.din(w_dff_A_Br5tP2ke6_1),.clk(gclk));
	jdff dff_A_kJVItLlC5_1(.dout(w_dff_A_Br5tP2ke6_1),.din(w_dff_A_kJVItLlC5_1),.clk(gclk));
	jdff dff_A_pFx1qlrF2_1(.dout(w_dff_A_kJVItLlC5_1),.din(w_dff_A_pFx1qlrF2_1),.clk(gclk));
	jdff dff_A_NyHcnITN2_0(.dout(w_n117_1[0]),.din(w_dff_A_NyHcnITN2_0),.clk(gclk));
	jdff dff_A_PjEsC2Nt6_0(.dout(w_dff_A_NyHcnITN2_0),.din(w_dff_A_PjEsC2Nt6_0),.clk(gclk));
	jdff dff_A_9hMNiwAr7_0(.dout(w_dff_A_PjEsC2Nt6_0),.din(w_dff_A_9hMNiwAr7_0),.clk(gclk));
	jdff dff_A_3FNVJZ6b6_0(.dout(w_dff_A_9hMNiwAr7_0),.din(w_dff_A_3FNVJZ6b6_0),.clk(gclk));
	jdff dff_A_BvcpixTz4_0(.dout(w_dff_A_3FNVJZ6b6_0),.din(w_dff_A_BvcpixTz4_0),.clk(gclk));
	jdff dff_A_OhMm5bUl1_1(.dout(w_n117_1[1]),.din(w_dff_A_OhMm5bUl1_1),.clk(gclk));
	jdff dff_A_FNmPuiPJ4_1(.dout(w_dff_A_OhMm5bUl1_1),.din(w_dff_A_FNmPuiPJ4_1),.clk(gclk));
	jdff dff_A_wzYEryQA7_1(.dout(w_dff_A_FNmPuiPJ4_1),.din(w_dff_A_wzYEryQA7_1),.clk(gclk));
	jdff dff_A_NlQU0y8n4_1(.dout(w_dff_A_wzYEryQA7_1),.din(w_dff_A_NlQU0y8n4_1),.clk(gclk));
	jdff dff_A_ANbbw8Pr3_1(.dout(w_dff_A_NlQU0y8n4_1),.din(w_dff_A_ANbbw8Pr3_1),.clk(gclk));
	jdff dff_B_I3NQ9kWv8_1(.din(n221),.dout(w_dff_B_I3NQ9kWv8_1),.clk(gclk));
	jdff dff_B_X2Im87NO5_1(.din(w_dff_B_I3NQ9kWv8_1),.dout(w_dff_B_X2Im87NO5_1),.clk(gclk));
	jdff dff_A_nkRXkBK28_0(.dout(w_n87_0[0]),.din(w_dff_A_nkRXkBK28_0),.clk(gclk));
	jdff dff_A_y2E5kge90_0(.dout(w_dff_A_nkRXkBK28_0),.din(w_dff_A_y2E5kge90_0),.clk(gclk));
	jdff dff_A_N0Qm4qx03_0(.dout(w_dff_A_y2E5kge90_0),.din(w_dff_A_N0Qm4qx03_0),.clk(gclk));
	jdff dff_A_KE3xKRPJ8_0(.dout(w_dff_A_N0Qm4qx03_0),.din(w_dff_A_KE3xKRPJ8_0),.clk(gclk));
	jdff dff_A_HDvR5fGe3_0(.dout(w_dff_A_KE3xKRPJ8_0),.din(w_dff_A_HDvR5fGe3_0),.clk(gclk));
	jdff dff_A_r5DYRlB56_2(.dout(w_n87_0[2]),.din(w_dff_A_r5DYRlB56_2),.clk(gclk));
	jdff dff_A_EXqygMbt8_2(.dout(w_dff_A_r5DYRlB56_2),.din(w_dff_A_EXqygMbt8_2),.clk(gclk));
	jdff dff_A_8TN8oAwb5_2(.dout(w_dff_A_EXqygMbt8_2),.din(w_dff_A_8TN8oAwb5_2),.clk(gclk));
	jdff dff_A_kg3pIg939_2(.dout(w_dff_A_8TN8oAwb5_2),.din(w_dff_A_kg3pIg939_2),.clk(gclk));
	jdff dff_A_7DImgA5K9_2(.dout(w_dff_A_kg3pIg939_2),.din(w_dff_A_7DImgA5K9_2),.clk(gclk));
	jdff dff_A_oCgw7TMx6_0(.dout(w_n187_1[0]),.din(w_dff_A_oCgw7TMx6_0),.clk(gclk));
	jdff dff_A_I1aMf9ZZ5_0(.dout(w_dff_A_oCgw7TMx6_0),.din(w_dff_A_I1aMf9ZZ5_0),.clk(gclk));
	jdff dff_A_YeY29Oym9_0(.dout(w_dff_A_I1aMf9ZZ5_0),.din(w_dff_A_YeY29Oym9_0),.clk(gclk));
	jdff dff_A_zBAy3kXJ3_0(.dout(w_dff_A_YeY29Oym9_0),.din(w_dff_A_zBAy3kXJ3_0),.clk(gclk));
	jdff dff_A_pFG4FcaY0_0(.dout(w_dff_A_zBAy3kXJ3_0),.din(w_dff_A_pFG4FcaY0_0),.clk(gclk));
	jdff dff_A_OnF2YcdG6_1(.dout(w_n187_1[1]),.din(w_dff_A_OnF2YcdG6_1),.clk(gclk));
	jdff dff_A_mPYlZrow8_1(.dout(w_dff_A_OnF2YcdG6_1),.din(w_dff_A_mPYlZrow8_1),.clk(gclk));
	jdff dff_A_fx5E7a5D4_1(.dout(w_dff_A_mPYlZrow8_1),.din(w_dff_A_fx5E7a5D4_1),.clk(gclk));
	jdff dff_A_CitHGTA41_1(.dout(w_dff_A_fx5E7a5D4_1),.din(w_dff_A_CitHGTA41_1),.clk(gclk));
	jdff dff_A_2DYJGpGs2_1(.dout(w_dff_A_CitHGTA41_1),.din(w_dff_A_2DYJGpGs2_1),.clk(gclk));
	jdff dff_B_Bvp8kghG2_2(.din(n220),.dout(w_dff_B_Bvp8kghG2_2),.clk(gclk));
	jdff dff_B_hw1dCfcE1_2(.din(w_dff_B_Bvp8kghG2_2),.dout(w_dff_B_hw1dCfcE1_2),.clk(gclk));
	jdff dff_B_ZnnCJ2u80_2(.din(w_dff_B_hw1dCfcE1_2),.dout(w_dff_B_ZnnCJ2u80_2),.clk(gclk));
	jdff dff_A_tAxc8FNh3_0(.dout(w_n181_0[0]),.din(w_dff_A_tAxc8FNh3_0),.clk(gclk));
	jdff dff_A_H9RAuYj59_0(.dout(w_dff_A_tAxc8FNh3_0),.din(w_dff_A_H9RAuYj59_0),.clk(gclk));
	jdff dff_A_zhKE0ORh8_0(.dout(w_dff_A_H9RAuYj59_0),.din(w_dff_A_zhKE0ORh8_0),.clk(gclk));
	jdff dff_A_978ixOg97_0(.dout(w_dff_A_zhKE0ORh8_0),.din(w_dff_A_978ixOg97_0),.clk(gclk));
	jdff dff_A_Z09T7J496_0(.dout(w_dff_A_978ixOg97_0),.din(w_dff_A_Z09T7J496_0),.clk(gclk));
	jdff dff_A_9vEsrmUR1_2(.dout(w_n181_0[2]),.din(w_dff_A_9vEsrmUR1_2),.clk(gclk));
	jdff dff_A_3GTNAkxF1_2(.dout(w_dff_A_9vEsrmUR1_2),.din(w_dff_A_3GTNAkxF1_2),.clk(gclk));
	jdff dff_A_S26JRI2o8_2(.dout(w_dff_A_3GTNAkxF1_2),.din(w_dff_A_S26JRI2o8_2),.clk(gclk));
	jdff dff_A_hf96O2073_2(.dout(w_dff_A_S26JRI2o8_2),.din(w_dff_A_hf96O2073_2),.clk(gclk));
	jdff dff_A_KepHnE5C4_2(.dout(w_dff_A_hf96O2073_2),.din(w_dff_A_KepHnE5C4_2),.clk(gclk));
	jdff dff_A_Pq1Q8flQ6_1(.dout(w_n164_0[1]),.din(w_dff_A_Pq1Q8flQ6_1),.clk(gclk));
	jdff dff_A_tiXy71DX0_1(.dout(w_dff_A_Pq1Q8flQ6_1),.din(w_dff_A_tiXy71DX0_1),.clk(gclk));
	jdff dff_A_J1RAxLIK9_1(.dout(w_dff_A_tiXy71DX0_1),.din(w_dff_A_J1RAxLIK9_1),.clk(gclk));
	jdff dff_A_xA55UyWX5_1(.dout(w_dff_A_J1RAxLIK9_1),.din(w_dff_A_xA55UyWX5_1),.clk(gclk));
	jdff dff_A_fiIPpVW66_1(.dout(w_dff_A_xA55UyWX5_1),.din(w_dff_A_fiIPpVW66_1),.clk(gclk));
	jdff dff_A_IZxkOlFJ1_2(.dout(w_n164_0[2]),.din(w_dff_A_IZxkOlFJ1_2),.clk(gclk));
	jdff dff_A_PRQAdJrd6_2(.dout(w_dff_A_IZxkOlFJ1_2),.din(w_dff_A_PRQAdJrd6_2),.clk(gclk));
	jdff dff_A_ruYlIlni4_2(.dout(w_dff_A_PRQAdJrd6_2),.din(w_dff_A_ruYlIlni4_2),.clk(gclk));
	jdff dff_A_OatywFOG1_2(.dout(w_dff_A_ruYlIlni4_2),.din(w_dff_A_OatywFOG1_2),.clk(gclk));
	jdff dff_A_neoNnWwU3_2(.dout(w_dff_A_OatywFOG1_2),.din(w_dff_A_neoNnWwU3_2),.clk(gclk));
	jdff dff_A_9woERz7Z9_0(.dout(w_n163_1[0]),.din(w_dff_A_9woERz7Z9_0),.clk(gclk));
	jdff dff_A_cI7o6xKU6_1(.dout(w_n199_0[1]),.din(w_dff_A_cI7o6xKU6_1),.clk(gclk));
	jdff dff_A_p6IPhVq52_1(.dout(w_dff_A_cI7o6xKU6_1),.din(w_dff_A_p6IPhVq52_1),.clk(gclk));
	jdff dff_A_x5ATtBGA0_1(.dout(w_dff_A_p6IPhVq52_1),.din(w_dff_A_x5ATtBGA0_1),.clk(gclk));
	jdff dff_A_s89WmVE65_1(.dout(w_dff_A_x5ATtBGA0_1),.din(w_dff_A_s89WmVE65_1),.clk(gclk));
	jdff dff_A_Pt4jPtr59_1(.dout(w_dff_A_s89WmVE65_1),.din(w_dff_A_Pt4jPtr59_1),.clk(gclk));
	jdff dff_A_jw7x2tkw3_2(.dout(w_n199_0[2]),.din(w_dff_A_jw7x2tkw3_2),.clk(gclk));
	jdff dff_A_6WsW1NfW8_2(.dout(w_dff_A_jw7x2tkw3_2),.din(w_dff_A_6WsW1NfW8_2),.clk(gclk));
	jdff dff_A_ShANqaSA1_2(.dout(w_dff_A_6WsW1NfW8_2),.din(w_dff_A_ShANqaSA1_2),.clk(gclk));
	jdff dff_A_qOihlfpz6_2(.dout(w_dff_A_ShANqaSA1_2),.din(w_dff_A_qOihlfpz6_2),.clk(gclk));
	jdff dff_A_dDSIcMPD8_2(.dout(w_dff_A_qOihlfpz6_2),.din(w_dff_A_dDSIcMPD8_2),.clk(gclk));
	jdff dff_A_Y51j7kVV7_1(.dout(w_n172_1[1]),.din(w_dff_A_Y51j7kVV7_1),.clk(gclk));
	jdff dff_A_NqSOUP0c2_1(.dout(w_n117_0[1]),.din(w_dff_A_NqSOUP0c2_1),.clk(gclk));
	jdff dff_A_G3ZB9A949_1(.dout(w_dff_A_NqSOUP0c2_1),.din(w_dff_A_G3ZB9A949_1),.clk(gclk));
	jdff dff_A_chUHDdp50_1(.dout(w_dff_A_G3ZB9A949_1),.din(w_dff_A_chUHDdp50_1),.clk(gclk));
	jdff dff_A_kjcJgFsq5_1(.dout(w_dff_A_chUHDdp50_1),.din(w_dff_A_kjcJgFsq5_1),.clk(gclk));
	jdff dff_A_C2tRsLlm2_1(.dout(w_dff_A_kjcJgFsq5_1),.din(w_dff_A_C2tRsLlm2_1),.clk(gclk));
	jdff dff_A_7ayfKDEO3_2(.dout(w_n117_0[2]),.din(w_dff_A_7ayfKDEO3_2),.clk(gclk));
	jdff dff_A_2uRtdZbc2_2(.dout(w_dff_A_7ayfKDEO3_2),.din(w_dff_A_2uRtdZbc2_2),.clk(gclk));
	jdff dff_A_4uP4cjSF1_2(.dout(w_dff_A_2uRtdZbc2_2),.din(w_dff_A_4uP4cjSF1_2),.clk(gclk));
	jdff dff_A_grZsy7Tu6_2(.dout(w_dff_A_4uP4cjSF1_2),.din(w_dff_A_grZsy7Tu6_2),.clk(gclk));
	jdff dff_A_6rL5Wax43_2(.dout(w_dff_A_grZsy7Tu6_2),.din(w_dff_A_6rL5Wax43_2),.clk(gclk));
	jdff dff_A_rIYE9OzL2_0(.dout(w_n116_1[0]),.din(w_dff_A_rIYE9OzL2_0),.clk(gclk));
	jdff dff_B_qyGoOx4d0_1(.din(n249),.dout(w_dff_B_qyGoOx4d0_1),.clk(gclk));
	jdff dff_B_gMAT52TG0_1(.din(w_dff_B_qyGoOx4d0_1),.dout(w_dff_B_gMAT52TG0_1),.clk(gclk));
	jdff dff_B_kBn5VUQX0_0(.din(n227),.dout(w_dff_B_kBn5VUQX0_0),.clk(gclk));
	jdff dff_A_xsODTihY7_2(.dout(w_n163_0[2]),.din(w_dff_A_xsODTihY7_2),.clk(gclk));
	jdff dff_A_k2sYJBL53_2(.dout(w_n172_0[2]),.din(w_dff_A_k2sYJBL53_2),.clk(gclk));
	jdff dff_A_xz3I73mA6_2(.dout(w_dff_A_k2sYJBL53_2),.din(w_dff_A_xz3I73mA6_2),.clk(gclk));
	jdff dff_A_g5l9RMl53_0(.dout(w_n178_0[0]),.din(w_dff_A_g5l9RMl53_0),.clk(gclk));
	jdff dff_A_y8KyCeV62_0(.dout(w_dff_A_g5l9RMl53_0),.din(w_dff_A_y8KyCeV62_0),.clk(gclk));
	jdff dff_A_ifxEZZu00_0(.dout(w_dff_A_y8KyCeV62_0),.din(w_dff_A_ifxEZZu00_0),.clk(gclk));
	jdff dff_A_SBY2aqI75_0(.dout(w_dff_A_ifxEZZu00_0),.din(w_dff_A_SBY2aqI75_0),.clk(gclk));
	jdff dff_A_awOn1qiS3_0(.dout(w_dff_A_SBY2aqI75_0),.din(w_dff_A_awOn1qiS3_0),.clk(gclk));
	jdff dff_A_PzVgNCOy3_2(.dout(w_n178_0[2]),.din(w_dff_A_PzVgNCOy3_2),.clk(gclk));
	jdff dff_A_kj68dVfq5_2(.dout(w_dff_A_PzVgNCOy3_2),.din(w_dff_A_kj68dVfq5_2),.clk(gclk));
	jdff dff_A_BI0MT9n17_2(.dout(w_dff_A_kj68dVfq5_2),.din(w_dff_A_BI0MT9n17_2),.clk(gclk));
	jdff dff_A_45F2Wfbn4_2(.dout(w_dff_A_BI0MT9n17_2),.din(w_dff_A_45F2Wfbn4_2),.clk(gclk));
	jdff dff_A_IBdGzWN69_2(.dout(w_dff_A_45F2Wfbn4_2),.din(w_dff_A_IBdGzWN69_2),.clk(gclk));
	jdff dff_A_bOqX34r50_1(.dout(w_n132_0[1]),.din(w_dff_A_bOqX34r50_1),.clk(gclk));
	jdff dff_A_nRDA2vYG6_0(.dout(w_G8gat_0[0]),.din(w_dff_A_nRDA2vYG6_0),.clk(gclk));
	jdff dff_A_Mym3gcbE7_0(.dout(w_dff_A_nRDA2vYG6_0),.din(w_dff_A_Mym3gcbE7_0),.clk(gclk));
	jdff dff_A_gRCIq3DY7_0(.dout(w_dff_A_Mym3gcbE7_0),.din(w_dff_A_gRCIq3DY7_0),.clk(gclk));
	jdff dff_A_tfc7ibsH7_0(.dout(w_dff_A_gRCIq3DY7_0),.din(w_dff_A_tfc7ibsH7_0),.clk(gclk));
	jdff dff_A_pNPAEwfB1_0(.dout(w_dff_A_tfc7ibsH7_0),.din(w_dff_A_pNPAEwfB1_0),.clk(gclk));
	jdff dff_A_H3vghLHm2_0(.dout(w_dff_A_pNPAEwfB1_0),.din(w_dff_A_H3vghLHm2_0),.clk(gclk));
	jdff dff_A_XkM3NqXz1_0(.dout(w_dff_A_H3vghLHm2_0),.din(w_dff_A_XkM3NqXz1_0),.clk(gclk));
	jdff dff_A_UTLB9La62_0(.dout(w_dff_A_XkM3NqXz1_0),.din(w_dff_A_UTLB9La62_0),.clk(gclk));
	jdff dff_A_nvOZlLyp4_0(.dout(w_dff_A_UTLB9La62_0),.din(w_dff_A_nvOZlLyp4_0),.clk(gclk));
	jdff dff_A_eKpGKkJK3_0(.dout(w_dff_A_nvOZlLyp4_0),.din(w_dff_A_eKpGKkJK3_0),.clk(gclk));
	jdff dff_A_iq1FECP85_0(.dout(w_dff_A_eKpGKkJK3_0),.din(w_dff_A_iq1FECP85_0),.clk(gclk));
	jdff dff_A_LLwYrFqp7_0(.dout(w_G64gat_0[0]),.din(w_dff_A_LLwYrFqp7_0),.clk(gclk));
	jdff dff_A_VMHuDbXW2_0(.dout(w_dff_A_LLwYrFqp7_0),.din(w_dff_A_VMHuDbXW2_0),.clk(gclk));
	jdff dff_A_6k0ZNcJS5_0(.dout(w_dff_A_VMHuDbXW2_0),.din(w_dff_A_6k0ZNcJS5_0),.clk(gclk));
	jdff dff_A_MY4xu2Sr4_0(.dout(w_dff_A_6k0ZNcJS5_0),.din(w_dff_A_MY4xu2Sr4_0),.clk(gclk));
	jdff dff_A_d58reL1z1_0(.dout(w_dff_A_MY4xu2Sr4_0),.din(w_dff_A_d58reL1z1_0),.clk(gclk));
	jdff dff_A_57UHzbkQ8_0(.dout(w_dff_A_d58reL1z1_0),.din(w_dff_A_57UHzbkQ8_0),.clk(gclk));
	jdff dff_A_817YCMfQ3_0(.dout(w_dff_A_57UHzbkQ8_0),.din(w_dff_A_817YCMfQ3_0),.clk(gclk));
	jdff dff_A_IG27HCOo2_0(.dout(w_dff_A_817YCMfQ3_0),.din(w_dff_A_IG27HCOo2_0),.clk(gclk));
	jdff dff_A_p8E3sw4r8_0(.dout(w_dff_A_IG27HCOo2_0),.din(w_dff_A_p8E3sw4r8_0),.clk(gclk));
	jdff dff_A_tEUrMgvT0_0(.dout(w_dff_A_p8E3sw4r8_0),.din(w_dff_A_tEUrMgvT0_0),.clk(gclk));
	jdff dff_A_D3IYoDKs3_0(.dout(w_dff_A_tEUrMgvT0_0),.din(w_dff_A_D3IYoDKs3_0),.clk(gclk));
	jdff dff_A_wHstNy2b2_1(.dout(w_n86_0[1]),.din(w_dff_A_wHstNy2b2_1),.clk(gclk));
	jdff dff_A_5WUuWzmE9_2(.dout(w_n86_0[2]),.din(w_dff_A_5WUuWzmE9_2),.clk(gclk));
	jdff dff_A_aMsv7RJo4_0(.dout(w_G1gat_0[0]),.din(w_dff_A_aMsv7RJo4_0),.clk(gclk));
	jdff dff_A_fqzMkq1x0_0(.dout(w_dff_A_aMsv7RJo4_0),.din(w_dff_A_fqzMkq1x0_0),.clk(gclk));
	jdff dff_A_mnjIAAwl1_0(.dout(w_dff_A_fqzMkq1x0_0),.din(w_dff_A_mnjIAAwl1_0),.clk(gclk));
	jdff dff_A_Q0rJsq7D2_0(.dout(w_dff_A_mnjIAAwl1_0),.din(w_dff_A_Q0rJsq7D2_0),.clk(gclk));
	jdff dff_A_zwJqievP9_0(.dout(w_dff_A_Q0rJsq7D2_0),.din(w_dff_A_zwJqievP9_0),.clk(gclk));
	jdff dff_A_8rcd7bQa7_0(.dout(w_dff_A_zwJqievP9_0),.din(w_dff_A_8rcd7bQa7_0),.clk(gclk));
	jdff dff_A_nXwlvstj8_0(.dout(w_dff_A_8rcd7bQa7_0),.din(w_dff_A_nXwlvstj8_0),.clk(gclk));
	jdff dff_A_HLWbYNWE0_0(.dout(w_dff_A_nXwlvstj8_0),.din(w_dff_A_HLWbYNWE0_0),.clk(gclk));
	jdff dff_A_FSgxPSWq7_0(.dout(w_dff_A_HLWbYNWE0_0),.din(w_dff_A_FSgxPSWq7_0),.clk(gclk));
	jdff dff_A_JCZNzEoJ9_0(.dout(w_dff_A_FSgxPSWq7_0),.din(w_dff_A_JCZNzEoJ9_0),.clk(gclk));
	jdff dff_A_UcmzbQkh5_0(.dout(w_dff_A_JCZNzEoJ9_0),.din(w_dff_A_UcmzbQkh5_0),.clk(gclk));
	jdff dff_A_B88P9Sez4_0(.dout(w_G57gat_0[0]),.din(w_dff_A_B88P9Sez4_0),.clk(gclk));
	jdff dff_A_FnxcZ3DO9_0(.dout(w_dff_A_B88P9Sez4_0),.din(w_dff_A_FnxcZ3DO9_0),.clk(gclk));
	jdff dff_A_46g3VgXk0_0(.dout(w_dff_A_FnxcZ3DO9_0),.din(w_dff_A_46g3VgXk0_0),.clk(gclk));
	jdff dff_A_e3Uxfk0L0_0(.dout(w_dff_A_46g3VgXk0_0),.din(w_dff_A_e3Uxfk0L0_0),.clk(gclk));
	jdff dff_A_D6pRyXT40_0(.dout(w_dff_A_e3Uxfk0L0_0),.din(w_dff_A_D6pRyXT40_0),.clk(gclk));
	jdff dff_A_AiXwK1vd9_0(.dout(w_dff_A_D6pRyXT40_0),.din(w_dff_A_AiXwK1vd9_0),.clk(gclk));
	jdff dff_A_z5VEzgME0_0(.dout(w_dff_A_AiXwK1vd9_0),.din(w_dff_A_z5VEzgME0_0),.clk(gclk));
	jdff dff_A_5sV6vwcA1_0(.dout(w_dff_A_z5VEzgME0_0),.din(w_dff_A_5sV6vwcA1_0),.clk(gclk));
	jdff dff_A_8Uo2JvBy7_0(.dout(w_dff_A_5sV6vwcA1_0),.din(w_dff_A_8Uo2JvBy7_0),.clk(gclk));
	jdff dff_A_sADhmOWS6_0(.dout(w_dff_A_8Uo2JvBy7_0),.din(w_dff_A_sADhmOWS6_0),.clk(gclk));
	jdff dff_A_l9rnSSI04_0(.dout(w_dff_A_sADhmOWS6_0),.din(w_dff_A_l9rnSSI04_0),.clk(gclk));
	jdff dff_B_HSHaE9Ih2_2(.din(n239),.dout(w_dff_B_HSHaE9Ih2_2),.clk(gclk));
	jdff dff_B_XNRly9na4_2(.din(w_dff_B_HSHaE9Ih2_2),.dout(w_dff_B_XNRly9na4_2),.clk(gclk));
	jdff dff_B_nHxscb9U4_2(.din(w_dff_B_XNRly9na4_2),.dout(w_dff_B_nHxscb9U4_2),.clk(gclk));
	jdff dff_A_y1RUfWp32_0(.dout(w_n184_0[0]),.din(w_dff_A_y1RUfWp32_0),.clk(gclk));
	jdff dff_A_j7cpPJAr6_0(.dout(w_dff_A_y1RUfWp32_0),.din(w_dff_A_j7cpPJAr6_0),.clk(gclk));
	jdff dff_A_YIskqoSz7_0(.dout(w_dff_A_j7cpPJAr6_0),.din(w_dff_A_YIskqoSz7_0),.clk(gclk));
	jdff dff_A_mmKCDQrv0_0(.dout(w_dff_A_YIskqoSz7_0),.din(w_dff_A_mmKCDQrv0_0),.clk(gclk));
	jdff dff_A_QkSzTCdN3_0(.dout(w_dff_A_mmKCDQrv0_0),.din(w_dff_A_QkSzTCdN3_0),.clk(gclk));
	jdff dff_A_M1aNCpEq0_2(.dout(w_n184_0[2]),.din(w_dff_A_M1aNCpEq0_2),.clk(gclk));
	jdff dff_A_xxP5WCIH0_2(.dout(w_dff_A_M1aNCpEq0_2),.din(w_dff_A_xxP5WCIH0_2),.clk(gclk));
	jdff dff_A_5wqRAZPE4_2(.dout(w_dff_A_xxP5WCIH0_2),.din(w_dff_A_5wqRAZPE4_2),.clk(gclk));
	jdff dff_A_3ECLkrun6_2(.dout(w_dff_A_5wqRAZPE4_2),.din(w_dff_A_3ECLkrun6_2),.clk(gclk));
	jdff dff_A_JKedJh0d4_2(.dout(w_dff_A_3ECLkrun6_2),.din(w_dff_A_JKedJh0d4_2),.clk(gclk));
	jdff dff_A_GSwAHdKK6_1(.dout(w_n149_0[1]),.din(w_dff_A_GSwAHdKK6_1),.clk(gclk));
	jdff dff_A_ddD5a0Aw5_0(.dout(w_G148gat_0[0]),.din(w_dff_A_ddD5a0Aw5_0),.clk(gclk));
	jdff dff_A_hvyyoF785_0(.dout(w_dff_A_ddD5a0Aw5_0),.din(w_dff_A_hvyyoF785_0),.clk(gclk));
	jdff dff_A_vOxg2hAo2_0(.dout(w_dff_A_hvyyoF785_0),.din(w_dff_A_vOxg2hAo2_0),.clk(gclk));
	jdff dff_A_ptyxYr8f2_0(.dout(w_dff_A_vOxg2hAo2_0),.din(w_dff_A_ptyxYr8f2_0),.clk(gclk));
	jdff dff_A_BSBT0qQK9_0(.dout(w_dff_A_ptyxYr8f2_0),.din(w_dff_A_BSBT0qQK9_0),.clk(gclk));
	jdff dff_A_7QY9nNvq6_0(.dout(w_dff_A_BSBT0qQK9_0),.din(w_dff_A_7QY9nNvq6_0),.clk(gclk));
	jdff dff_A_np3P7awH0_0(.dout(w_dff_A_7QY9nNvq6_0),.din(w_dff_A_np3P7awH0_0),.clk(gclk));
	jdff dff_A_gixtXHhu8_0(.dout(w_dff_A_np3P7awH0_0),.din(w_dff_A_gixtXHhu8_0),.clk(gclk));
	jdff dff_A_16IA2rWe6_0(.dout(w_dff_A_gixtXHhu8_0),.din(w_dff_A_16IA2rWe6_0),.clk(gclk));
	jdff dff_A_XwxqnrD51_0(.dout(w_dff_A_16IA2rWe6_0),.din(w_dff_A_XwxqnrD51_0),.clk(gclk));
	jdff dff_A_rrqo86Nk9_0(.dout(w_dff_A_XwxqnrD51_0),.din(w_dff_A_rrqo86Nk9_0),.clk(gclk));
	jdff dff_A_5ZT7LSoQ0_0(.dout(w_G141gat_0[0]),.din(w_dff_A_5ZT7LSoQ0_0),.clk(gclk));
	jdff dff_A_bTiiKfGM2_0(.dout(w_dff_A_5ZT7LSoQ0_0),.din(w_dff_A_bTiiKfGM2_0),.clk(gclk));
	jdff dff_A_fZCFhG694_0(.dout(w_dff_A_bTiiKfGM2_0),.din(w_dff_A_fZCFhG694_0),.clk(gclk));
	jdff dff_A_sNfeIk8T6_0(.dout(w_dff_A_fZCFhG694_0),.din(w_dff_A_sNfeIk8T6_0),.clk(gclk));
	jdff dff_A_d1EHCy0X4_0(.dout(w_dff_A_sNfeIk8T6_0),.din(w_dff_A_d1EHCy0X4_0),.clk(gclk));
	jdff dff_A_7ulYWxJU5_0(.dout(w_dff_A_d1EHCy0X4_0),.din(w_dff_A_7ulYWxJU5_0),.clk(gclk));
	jdff dff_A_sRQ6aVyO3_0(.dout(w_dff_A_7ulYWxJU5_0),.din(w_dff_A_sRQ6aVyO3_0),.clk(gclk));
	jdff dff_A_fDNR9epd3_0(.dout(w_dff_A_sRQ6aVyO3_0),.din(w_dff_A_fDNR9epd3_0),.clk(gclk));
	jdff dff_A_wBEH4Wj33_0(.dout(w_dff_A_fDNR9epd3_0),.din(w_dff_A_wBEH4Wj33_0),.clk(gclk));
	jdff dff_A_DeyXqbRp9_0(.dout(w_dff_A_wBEH4Wj33_0),.din(w_dff_A_DeyXqbRp9_0),.clk(gclk));
	jdff dff_A_4US1ySSH8_0(.dout(w_dff_A_DeyXqbRp9_0),.din(w_dff_A_4US1ySSH8_0),.clk(gclk));
	jdff dff_A_lnIce6xP3_0(.dout(w_G155gat_0[0]),.din(w_dff_A_lnIce6xP3_0),.clk(gclk));
	jdff dff_A_sic6zVz01_0(.dout(w_dff_A_lnIce6xP3_0),.din(w_dff_A_sic6zVz01_0),.clk(gclk));
	jdff dff_A_rwoTpeUC7_0(.dout(w_dff_A_sic6zVz01_0),.din(w_dff_A_rwoTpeUC7_0),.clk(gclk));
	jdff dff_A_ZGUuCZRu1_0(.dout(w_dff_A_rwoTpeUC7_0),.din(w_dff_A_ZGUuCZRu1_0),.clk(gclk));
	jdff dff_A_uamd48YW7_0(.dout(w_dff_A_ZGUuCZRu1_0),.din(w_dff_A_uamd48YW7_0),.clk(gclk));
	jdff dff_A_8UeOxRJh2_0(.dout(w_dff_A_uamd48YW7_0),.din(w_dff_A_8UeOxRJh2_0),.clk(gclk));
	jdff dff_A_LNp6Muz40_0(.dout(w_dff_A_8UeOxRJh2_0),.din(w_dff_A_LNp6Muz40_0),.clk(gclk));
	jdff dff_A_s02xCIfa1_0(.dout(w_dff_A_LNp6Muz40_0),.din(w_dff_A_s02xCIfa1_0),.clk(gclk));
	jdff dff_A_TKIVSopJ8_0(.dout(w_dff_A_s02xCIfa1_0),.din(w_dff_A_TKIVSopJ8_0),.clk(gclk));
	jdff dff_A_U2BrVfOt1_0(.dout(w_dff_A_TKIVSopJ8_0),.din(w_dff_A_U2BrVfOt1_0),.clk(gclk));
	jdff dff_A_Q9CXhgde5_0(.dout(w_dff_A_U2BrVfOt1_0),.din(w_dff_A_Q9CXhgde5_0),.clk(gclk));
	jdff dff_A_53kmCpTX7_0(.dout(w_G22gat_0[0]),.din(w_dff_A_53kmCpTX7_0),.clk(gclk));
	jdff dff_A_hyBkMIIC4_0(.dout(w_dff_A_53kmCpTX7_0),.din(w_dff_A_hyBkMIIC4_0),.clk(gclk));
	jdff dff_A_wiS5E5NZ3_0(.dout(w_dff_A_hyBkMIIC4_0),.din(w_dff_A_wiS5E5NZ3_0),.clk(gclk));
	jdff dff_A_85Ht0P2y9_0(.dout(w_dff_A_wiS5E5NZ3_0),.din(w_dff_A_85Ht0P2y9_0),.clk(gclk));
	jdff dff_A_rdvvKlaS2_0(.dout(w_dff_A_85Ht0P2y9_0),.din(w_dff_A_rdvvKlaS2_0),.clk(gclk));
	jdff dff_A_EDDOjM8Z0_0(.dout(w_dff_A_rdvvKlaS2_0),.din(w_dff_A_EDDOjM8Z0_0),.clk(gclk));
	jdff dff_A_vDLbXTvY4_0(.dout(w_dff_A_EDDOjM8Z0_0),.din(w_dff_A_vDLbXTvY4_0),.clk(gclk));
	jdff dff_A_qmiZIMVd8_0(.dout(w_dff_A_vDLbXTvY4_0),.din(w_dff_A_qmiZIMVd8_0),.clk(gclk));
	jdff dff_A_nv0TeVXs4_0(.dout(w_dff_A_qmiZIMVd8_0),.din(w_dff_A_nv0TeVXs4_0),.clk(gclk));
	jdff dff_A_8e3J57y30_0(.dout(w_dff_A_nv0TeVXs4_0),.din(w_dff_A_8e3J57y30_0),.clk(gclk));
	jdff dff_A_axs5ry7q1_0(.dout(w_dff_A_8e3J57y30_0),.din(w_dff_A_axs5ry7q1_0),.clk(gclk));
	jdff dff_A_x43OYFnI8_0(.dout(w_G78gat_0[0]),.din(w_dff_A_x43OYFnI8_0),.clk(gclk));
	jdff dff_A_9WX8LZch9_0(.dout(w_dff_A_x43OYFnI8_0),.din(w_dff_A_9WX8LZch9_0),.clk(gclk));
	jdff dff_A_vkyOKHke5_0(.dout(w_dff_A_9WX8LZch9_0),.din(w_dff_A_vkyOKHke5_0),.clk(gclk));
	jdff dff_A_2NzI4PPC1_0(.dout(w_dff_A_vkyOKHke5_0),.din(w_dff_A_2NzI4PPC1_0),.clk(gclk));
	jdff dff_A_W5cq667D0_0(.dout(w_dff_A_2NzI4PPC1_0),.din(w_dff_A_W5cq667D0_0),.clk(gclk));
	jdff dff_A_QDoA0WXj3_0(.dout(w_dff_A_W5cq667D0_0),.din(w_dff_A_QDoA0WXj3_0),.clk(gclk));
	jdff dff_A_bJzb9TiQ3_0(.dout(w_dff_A_QDoA0WXj3_0),.din(w_dff_A_bJzb9TiQ3_0),.clk(gclk));
	jdff dff_A_KiDbmSMU7_0(.dout(w_dff_A_bJzb9TiQ3_0),.din(w_dff_A_KiDbmSMU7_0),.clk(gclk));
	jdff dff_A_IRWXDphX8_0(.dout(w_dff_A_KiDbmSMU7_0),.din(w_dff_A_IRWXDphX8_0),.clk(gclk));
	jdff dff_A_Rv7Ika1y6_0(.dout(w_dff_A_IRWXDphX8_0),.din(w_dff_A_Rv7Ika1y6_0),.clk(gclk));
	jdff dff_A_RaPgyqEB0_0(.dout(w_dff_A_Rv7Ika1y6_0),.din(w_dff_A_RaPgyqEB0_0),.clk(gclk));
	jdff dff_A_8UClQlks9_0(.dout(w_G204gat_0[0]),.din(w_dff_A_8UClQlks9_0),.clk(gclk));
	jdff dff_A_aDxvsTPX7_0(.dout(w_dff_A_8UClQlks9_0),.din(w_dff_A_aDxvsTPX7_0),.clk(gclk));
	jdff dff_A_oFeujOQt1_0(.dout(w_dff_A_aDxvsTPX7_0),.din(w_dff_A_oFeujOQt1_0),.clk(gclk));
	jdff dff_A_10V6IQla6_0(.dout(w_dff_A_oFeujOQt1_0),.din(w_dff_A_10V6IQla6_0),.clk(gclk));
	jdff dff_A_76AAjDM61_0(.dout(w_dff_A_10V6IQla6_0),.din(w_dff_A_76AAjDM61_0),.clk(gclk));
	jdff dff_A_4OFky0sv7_0(.dout(w_dff_A_76AAjDM61_0),.din(w_dff_A_4OFky0sv7_0),.clk(gclk));
	jdff dff_A_DrSqs3n32_0(.dout(w_dff_A_4OFky0sv7_0),.din(w_dff_A_DrSqs3n32_0),.clk(gclk));
	jdff dff_A_AjUdYfVM5_0(.dout(w_dff_A_DrSqs3n32_0),.din(w_dff_A_AjUdYfVM5_0),.clk(gclk));
	jdff dff_A_4tQryBox6_0(.dout(w_dff_A_AjUdYfVM5_0),.din(w_dff_A_4tQryBox6_0),.clk(gclk));
	jdff dff_A_zRUc7yJH0_0(.dout(w_dff_A_4tQryBox6_0),.din(w_dff_A_zRUc7yJH0_0),.clk(gclk));
	jdff dff_A_NpQuwQpU9_0(.dout(w_dff_A_zRUc7yJH0_0),.din(w_dff_A_NpQuwQpU9_0),.clk(gclk));
	jdff dff_A_0kag68kR1_0(.dout(w_G197gat_0[0]),.din(w_dff_A_0kag68kR1_0),.clk(gclk));
	jdff dff_A_zjPOeu2C6_0(.dout(w_dff_A_0kag68kR1_0),.din(w_dff_A_zjPOeu2C6_0),.clk(gclk));
	jdff dff_A_Bc0fjxVV8_0(.dout(w_dff_A_zjPOeu2C6_0),.din(w_dff_A_Bc0fjxVV8_0),.clk(gclk));
	jdff dff_A_VWomtTTY1_0(.dout(w_dff_A_Bc0fjxVV8_0),.din(w_dff_A_VWomtTTY1_0),.clk(gclk));
	jdff dff_A_RgvbKDty8_0(.dout(w_dff_A_VWomtTTY1_0),.din(w_dff_A_RgvbKDty8_0),.clk(gclk));
	jdff dff_A_EH6tmStE3_0(.dout(w_dff_A_RgvbKDty8_0),.din(w_dff_A_EH6tmStE3_0),.clk(gclk));
	jdff dff_A_2WpoxvPT7_0(.dout(w_dff_A_EH6tmStE3_0),.din(w_dff_A_2WpoxvPT7_0),.clk(gclk));
	jdff dff_A_F3OywF0E2_0(.dout(w_dff_A_2WpoxvPT7_0),.din(w_dff_A_F3OywF0E2_0),.clk(gclk));
	jdff dff_A_ZYFOHQcy8_0(.dout(w_dff_A_F3OywF0E2_0),.din(w_dff_A_ZYFOHQcy8_0),.clk(gclk));
	jdff dff_A_lVVieE0z3_0(.dout(w_dff_A_ZYFOHQcy8_0),.din(w_dff_A_lVVieE0z3_0),.clk(gclk));
	jdff dff_A_vfHsKIz05_0(.dout(w_dff_A_lVVieE0z3_0),.din(w_dff_A_vfHsKIz05_0),.clk(gclk));
	jdff dff_A_tUPJ8xBQ2_0(.dout(w_G211gat_0[0]),.din(w_dff_A_tUPJ8xBQ2_0),.clk(gclk));
	jdff dff_A_qJpb2hhC9_0(.dout(w_dff_A_tUPJ8xBQ2_0),.din(w_dff_A_qJpb2hhC9_0),.clk(gclk));
	jdff dff_A_mZlViL2C3_0(.dout(w_dff_A_qJpb2hhC9_0),.din(w_dff_A_mZlViL2C3_0),.clk(gclk));
	jdff dff_A_dIzhVf4v7_0(.dout(w_dff_A_mZlViL2C3_0),.din(w_dff_A_dIzhVf4v7_0),.clk(gclk));
	jdff dff_A_JhQ1WFom2_0(.dout(w_dff_A_dIzhVf4v7_0),.din(w_dff_A_JhQ1WFom2_0),.clk(gclk));
	jdff dff_A_HrFpJHTX4_0(.dout(w_dff_A_JhQ1WFom2_0),.din(w_dff_A_HrFpJHTX4_0),.clk(gclk));
	jdff dff_A_i1uTj3yO9_0(.dout(w_dff_A_HrFpJHTX4_0),.din(w_dff_A_i1uTj3yO9_0),.clk(gclk));
	jdff dff_A_Kdk8Zcjt9_0(.dout(w_dff_A_i1uTj3yO9_0),.din(w_dff_A_Kdk8Zcjt9_0),.clk(gclk));
	jdff dff_A_zsblTJ4d8_0(.dout(w_dff_A_Kdk8Zcjt9_0),.din(w_dff_A_zsblTJ4d8_0),.clk(gclk));
	jdff dff_A_dU3kP5r20_0(.dout(w_dff_A_zsblTJ4d8_0),.din(w_dff_A_dU3kP5r20_0),.clk(gclk));
	jdff dff_A_yreAeIPE7_0(.dout(w_dff_A_dU3kP5r20_0),.din(w_dff_A_yreAeIPE7_0),.clk(gclk));
	jdff dff_A_gx2kTY761_1(.dout(w_n141_0[1]),.din(w_dff_A_gx2kTY761_1),.clk(gclk));
	jdff dff_A_KvbXou8D0_0(.dout(w_G120gat_0[0]),.din(w_dff_A_KvbXou8D0_0),.clk(gclk));
	jdff dff_A_RvvEEplq5_0(.dout(w_dff_A_KvbXou8D0_0),.din(w_dff_A_RvvEEplq5_0),.clk(gclk));
	jdff dff_A_RSoabOWz8_0(.dout(w_dff_A_RvvEEplq5_0),.din(w_dff_A_RSoabOWz8_0),.clk(gclk));
	jdff dff_A_A6blB7S96_0(.dout(w_dff_A_RSoabOWz8_0),.din(w_dff_A_A6blB7S96_0),.clk(gclk));
	jdff dff_A_zNJAKhRu8_0(.dout(w_dff_A_A6blB7S96_0),.din(w_dff_A_zNJAKhRu8_0),.clk(gclk));
	jdff dff_A_ef7t8ovF2_0(.dout(w_dff_A_zNJAKhRu8_0),.din(w_dff_A_ef7t8ovF2_0),.clk(gclk));
	jdff dff_A_6EwLDQLU9_0(.dout(w_dff_A_ef7t8ovF2_0),.din(w_dff_A_6EwLDQLU9_0),.clk(gclk));
	jdff dff_A_GOkfIyGo4_0(.dout(w_dff_A_6EwLDQLU9_0),.din(w_dff_A_GOkfIyGo4_0),.clk(gclk));
	jdff dff_A_Pu10F1fI7_0(.dout(w_dff_A_GOkfIyGo4_0),.din(w_dff_A_Pu10F1fI7_0),.clk(gclk));
	jdff dff_A_VpVb5lPW9_0(.dout(w_dff_A_Pu10F1fI7_0),.din(w_dff_A_VpVb5lPW9_0),.clk(gclk));
	jdff dff_A_RNbr4DrG7_0(.dout(w_dff_A_VpVb5lPW9_0),.din(w_dff_A_RNbr4DrG7_0),.clk(gclk));
	jdff dff_A_Uvq2ISC13_0(.dout(w_G113gat_0[0]),.din(w_dff_A_Uvq2ISC13_0),.clk(gclk));
	jdff dff_A_7NHM8MYj7_0(.dout(w_dff_A_Uvq2ISC13_0),.din(w_dff_A_7NHM8MYj7_0),.clk(gclk));
	jdff dff_A_2B33gQmD1_0(.dout(w_dff_A_7NHM8MYj7_0),.din(w_dff_A_2B33gQmD1_0),.clk(gclk));
	jdff dff_A_VU7Wfq9c0_0(.dout(w_dff_A_2B33gQmD1_0),.din(w_dff_A_VU7Wfq9c0_0),.clk(gclk));
	jdff dff_A_E64gVZvF1_0(.dout(w_dff_A_VU7Wfq9c0_0),.din(w_dff_A_E64gVZvF1_0),.clk(gclk));
	jdff dff_A_oTj1Gib57_0(.dout(w_dff_A_E64gVZvF1_0),.din(w_dff_A_oTj1Gib57_0),.clk(gclk));
	jdff dff_A_3QTYpOlI5_0(.dout(w_dff_A_oTj1Gib57_0),.din(w_dff_A_3QTYpOlI5_0),.clk(gclk));
	jdff dff_A_InFSudi49_0(.dout(w_dff_A_3QTYpOlI5_0),.din(w_dff_A_InFSudi49_0),.clk(gclk));
	jdff dff_A_cckRExhv2_0(.dout(w_dff_A_InFSudi49_0),.din(w_dff_A_cckRExhv2_0),.clk(gclk));
	jdff dff_A_FDtq2BbX6_0(.dout(w_dff_A_cckRExhv2_0),.din(w_dff_A_FDtq2BbX6_0),.clk(gclk));
	jdff dff_A_9ZJCqNHa9_0(.dout(w_dff_A_FDtq2BbX6_0),.din(w_dff_A_9ZJCqNHa9_0),.clk(gclk));
	jdff dff_A_xLHFZHh25_0(.dout(w_G127gat_0[0]),.din(w_dff_A_xLHFZHh25_0),.clk(gclk));
	jdff dff_A_jH5hUEm57_0(.dout(w_dff_A_xLHFZHh25_0),.din(w_dff_A_jH5hUEm57_0),.clk(gclk));
	jdff dff_A_k2y2WbVO4_0(.dout(w_dff_A_jH5hUEm57_0),.din(w_dff_A_k2y2WbVO4_0),.clk(gclk));
	jdff dff_A_KPvoMPps7_0(.dout(w_dff_A_k2y2WbVO4_0),.din(w_dff_A_KPvoMPps7_0),.clk(gclk));
	jdff dff_A_zoXmEvjH7_0(.dout(w_dff_A_KPvoMPps7_0),.din(w_dff_A_zoXmEvjH7_0),.clk(gclk));
	jdff dff_A_I9ltBUix1_0(.dout(w_dff_A_zoXmEvjH7_0),.din(w_dff_A_I9ltBUix1_0),.clk(gclk));
	jdff dff_A_8rerxCpB2_0(.dout(w_dff_A_I9ltBUix1_0),.din(w_dff_A_8rerxCpB2_0),.clk(gclk));
	jdff dff_A_zOoOuxQo5_0(.dout(w_dff_A_8rerxCpB2_0),.din(w_dff_A_zOoOuxQo5_0),.clk(gclk));
	jdff dff_A_dyUIIFQ78_0(.dout(w_dff_A_zOoOuxQo5_0),.din(w_dff_A_dyUIIFQ78_0),.clk(gclk));
	jdff dff_A_NW3saaZP9_0(.dout(w_dff_A_dyUIIFQ78_0),.din(w_dff_A_NW3saaZP9_0),.clk(gclk));
	jdff dff_A_WzdV4eai8_0(.dout(w_dff_A_NW3saaZP9_0),.din(w_dff_A_WzdV4eai8_0),.clk(gclk));
	jdff dff_A_e4m04q3B9_0(.dout(w_G15gat_0[0]),.din(w_dff_A_e4m04q3B9_0),.clk(gclk));
	jdff dff_A_aJENA3Po1_0(.dout(w_dff_A_e4m04q3B9_0),.din(w_dff_A_aJENA3Po1_0),.clk(gclk));
	jdff dff_A_CnrwW58Q0_0(.dout(w_dff_A_aJENA3Po1_0),.din(w_dff_A_CnrwW58Q0_0),.clk(gclk));
	jdff dff_A_aITPlvab5_0(.dout(w_dff_A_CnrwW58Q0_0),.din(w_dff_A_aITPlvab5_0),.clk(gclk));
	jdff dff_A_1UeYkWGW6_0(.dout(w_dff_A_aITPlvab5_0),.din(w_dff_A_1UeYkWGW6_0),.clk(gclk));
	jdff dff_A_mnYtbXEY3_0(.dout(w_dff_A_1UeYkWGW6_0),.din(w_dff_A_mnYtbXEY3_0),.clk(gclk));
	jdff dff_A_AfU7IXd18_0(.dout(w_dff_A_mnYtbXEY3_0),.din(w_dff_A_AfU7IXd18_0),.clk(gclk));
	jdff dff_A_57nUM4lY3_0(.dout(w_dff_A_AfU7IXd18_0),.din(w_dff_A_57nUM4lY3_0),.clk(gclk));
	jdff dff_A_7qUonzYj2_0(.dout(w_dff_A_57nUM4lY3_0),.din(w_dff_A_7qUonzYj2_0),.clk(gclk));
	jdff dff_A_JAcdjA6v9_0(.dout(w_dff_A_7qUonzYj2_0),.din(w_dff_A_JAcdjA6v9_0),.clk(gclk));
	jdff dff_A_DGF6gZJt9_0(.dout(w_dff_A_JAcdjA6v9_0),.din(w_dff_A_DGF6gZJt9_0),.clk(gclk));
	jdff dff_A_iWPGaqeT9_0(.dout(w_G71gat_0[0]),.din(w_dff_A_iWPGaqeT9_0),.clk(gclk));
	jdff dff_A_tHhgsdKJ8_0(.dout(w_dff_A_iWPGaqeT9_0),.din(w_dff_A_tHhgsdKJ8_0),.clk(gclk));
	jdff dff_A_XLpT9dqa2_0(.dout(w_dff_A_tHhgsdKJ8_0),.din(w_dff_A_XLpT9dqa2_0),.clk(gclk));
	jdff dff_A_j4B1sx2o1_0(.dout(w_dff_A_XLpT9dqa2_0),.din(w_dff_A_j4B1sx2o1_0),.clk(gclk));
	jdff dff_A_AbQnepcZ1_0(.dout(w_dff_A_j4B1sx2o1_0),.din(w_dff_A_AbQnepcZ1_0),.clk(gclk));
	jdff dff_A_k9osiVcG7_0(.dout(w_dff_A_AbQnepcZ1_0),.din(w_dff_A_k9osiVcG7_0),.clk(gclk));
	jdff dff_A_VFCyZIEE9_0(.dout(w_dff_A_k9osiVcG7_0),.din(w_dff_A_VFCyZIEE9_0),.clk(gclk));
	jdff dff_A_QFLZhNPM4_0(.dout(w_dff_A_VFCyZIEE9_0),.din(w_dff_A_QFLZhNPM4_0),.clk(gclk));
	jdff dff_A_h6RqiRQ63_0(.dout(w_dff_A_QFLZhNPM4_0),.din(w_dff_A_h6RqiRQ63_0),.clk(gclk));
	jdff dff_A_tPOqLmLd3_0(.dout(w_dff_A_h6RqiRQ63_0),.din(w_dff_A_tPOqLmLd3_0),.clk(gclk));
	jdff dff_A_tVGFvDGq0_0(.dout(w_dff_A_tPOqLmLd3_0),.din(w_dff_A_tVGFvDGq0_0),.clk(gclk));
	jdff dff_A_V7659hYV8_0(.dout(w_G176gat_0[0]),.din(w_dff_A_V7659hYV8_0),.clk(gclk));
	jdff dff_A_904aWuNT2_0(.dout(w_dff_A_V7659hYV8_0),.din(w_dff_A_904aWuNT2_0),.clk(gclk));
	jdff dff_A_dkWeLLyS6_0(.dout(w_dff_A_904aWuNT2_0),.din(w_dff_A_dkWeLLyS6_0),.clk(gclk));
	jdff dff_A_t7yj3dmV4_0(.dout(w_dff_A_dkWeLLyS6_0),.din(w_dff_A_t7yj3dmV4_0),.clk(gclk));
	jdff dff_A_tKFWOP2H5_0(.dout(w_dff_A_t7yj3dmV4_0),.din(w_dff_A_tKFWOP2H5_0),.clk(gclk));
	jdff dff_A_TcfeqVxa7_0(.dout(w_dff_A_tKFWOP2H5_0),.din(w_dff_A_TcfeqVxa7_0),.clk(gclk));
	jdff dff_A_0nMjYDmr2_0(.dout(w_dff_A_TcfeqVxa7_0),.din(w_dff_A_0nMjYDmr2_0),.clk(gclk));
	jdff dff_A_zret7jSo2_0(.dout(w_dff_A_0nMjYDmr2_0),.din(w_dff_A_zret7jSo2_0),.clk(gclk));
	jdff dff_A_YIBYXjAd8_0(.dout(w_dff_A_zret7jSo2_0),.din(w_dff_A_YIBYXjAd8_0),.clk(gclk));
	jdff dff_A_J88dYbRL2_0(.dout(w_dff_A_YIBYXjAd8_0),.din(w_dff_A_J88dYbRL2_0),.clk(gclk));
	jdff dff_A_7v7dT4Ll9_0(.dout(w_dff_A_J88dYbRL2_0),.din(w_dff_A_7v7dT4Ll9_0),.clk(gclk));
	jdff dff_A_KjBgybxO9_0(.dout(w_G169gat_0[0]),.din(w_dff_A_KjBgybxO9_0),.clk(gclk));
	jdff dff_A_luIVE5603_0(.dout(w_dff_A_KjBgybxO9_0),.din(w_dff_A_luIVE5603_0),.clk(gclk));
	jdff dff_A_rTeWKTuK5_0(.dout(w_dff_A_luIVE5603_0),.din(w_dff_A_rTeWKTuK5_0),.clk(gclk));
	jdff dff_A_UqGw2XlN2_0(.dout(w_dff_A_rTeWKTuK5_0),.din(w_dff_A_UqGw2XlN2_0),.clk(gclk));
	jdff dff_A_CENrdQJ84_0(.dout(w_dff_A_UqGw2XlN2_0),.din(w_dff_A_CENrdQJ84_0),.clk(gclk));
	jdff dff_A_PmM4NndX9_0(.dout(w_dff_A_CENrdQJ84_0),.din(w_dff_A_PmM4NndX9_0),.clk(gclk));
	jdff dff_A_RHrH6hO82_0(.dout(w_dff_A_PmM4NndX9_0),.din(w_dff_A_RHrH6hO82_0),.clk(gclk));
	jdff dff_A_fue47tCg2_0(.dout(w_dff_A_RHrH6hO82_0),.din(w_dff_A_fue47tCg2_0),.clk(gclk));
	jdff dff_A_8NznfdDM5_0(.dout(w_dff_A_fue47tCg2_0),.din(w_dff_A_8NznfdDM5_0),.clk(gclk));
	jdff dff_A_CuWHA5Yp4_0(.dout(w_dff_A_8NznfdDM5_0),.din(w_dff_A_CuWHA5Yp4_0),.clk(gclk));
	jdff dff_A_M6HBiUCH5_0(.dout(w_dff_A_CuWHA5Yp4_0),.din(w_dff_A_M6HBiUCH5_0),.clk(gclk));
	jdff dff_A_oJO62Rp16_0(.dout(w_G183gat_0[0]),.din(w_dff_A_oJO62Rp16_0),.clk(gclk));
	jdff dff_A_z7UbHL3d5_0(.dout(w_dff_A_oJO62Rp16_0),.din(w_dff_A_z7UbHL3d5_0),.clk(gclk));
	jdff dff_A_1aYYLMj23_0(.dout(w_dff_A_z7UbHL3d5_0),.din(w_dff_A_1aYYLMj23_0),.clk(gclk));
	jdff dff_A_ZyrqKgsj1_0(.dout(w_dff_A_1aYYLMj23_0),.din(w_dff_A_ZyrqKgsj1_0),.clk(gclk));
	jdff dff_A_Z1jwAMuK9_0(.dout(w_dff_A_ZyrqKgsj1_0),.din(w_dff_A_Z1jwAMuK9_0),.clk(gclk));
	jdff dff_A_tPPdVKKG0_0(.dout(w_dff_A_Z1jwAMuK9_0),.din(w_dff_A_tPPdVKKG0_0),.clk(gclk));
	jdff dff_A_sfJWps624_0(.dout(w_dff_A_tPPdVKKG0_0),.din(w_dff_A_sfJWps624_0),.clk(gclk));
	jdff dff_A_EJdh07eS4_0(.dout(w_dff_A_sfJWps624_0),.din(w_dff_A_EJdh07eS4_0),.clk(gclk));
	jdff dff_A_cJdhGI191_0(.dout(w_dff_A_EJdh07eS4_0),.din(w_dff_A_cJdhGI191_0),.clk(gclk));
	jdff dff_A_ocWcBmRt3_0(.dout(w_dff_A_cJdhGI191_0),.din(w_dff_A_ocWcBmRt3_0),.clk(gclk));
	jdff dff_A_ZQIL4zOV3_0(.dout(w_dff_A_ocWcBmRt3_0),.din(w_dff_A_ZQIL4zOV3_0),.clk(gclk));
	jdff dff_A_TnMHhmql2_1(.dout(w_n187_0[1]),.din(w_dff_A_TnMHhmql2_1),.clk(gclk));
	jdff dff_A_CxeUrvIJ4_1(.dout(w_dff_A_TnMHhmql2_1),.din(w_dff_A_CxeUrvIJ4_1),.clk(gclk));
	jdff dff_A_JCTjOkmL1_1(.dout(w_dff_A_CxeUrvIJ4_1),.din(w_dff_A_JCTjOkmL1_1),.clk(gclk));
	jdff dff_A_PrT1bVMz2_1(.dout(w_dff_A_JCTjOkmL1_1),.din(w_dff_A_PrT1bVMz2_1),.clk(gclk));
	jdff dff_A_oKvAYkiG8_1(.dout(w_dff_A_PrT1bVMz2_1),.din(w_dff_A_oKvAYkiG8_1),.clk(gclk));
	jdff dff_A_DSe6qKbN2_2(.dout(w_n187_0[2]),.din(w_dff_A_DSe6qKbN2_2),.clk(gclk));
	jdff dff_A_lkQsU6Fo1_2(.dout(w_dff_A_DSe6qKbN2_2),.din(w_dff_A_lkQsU6Fo1_2),.clk(gclk));
	jdff dff_A_hFQ7RFzM3_2(.dout(w_dff_A_lkQsU6Fo1_2),.din(w_dff_A_hFQ7RFzM3_2),.clk(gclk));
	jdff dff_A_TYAYYZlu6_2(.dout(w_dff_A_hFQ7RFzM3_2),.din(w_dff_A_TYAYYZlu6_2),.clk(gclk));
	jdff dff_A_oeYXzT0W7_2(.dout(w_dff_A_TYAYYZlu6_2),.din(w_dff_A_oeYXzT0W7_2),.clk(gclk));
	jdff dff_A_XXy1jOTI2_1(.dout(w_n102_1[1]),.din(w_dff_A_XXy1jOTI2_1),.clk(gclk));
	jdff dff_A_JWYMyi2G2_0(.dout(w_G36gat_0[0]),.din(w_dff_A_JWYMyi2G2_0),.clk(gclk));
	jdff dff_A_YhzLEPzi5_0(.dout(w_dff_A_JWYMyi2G2_0),.din(w_dff_A_YhzLEPzi5_0),.clk(gclk));
	jdff dff_A_laAcwvOq2_0(.dout(w_dff_A_YhzLEPzi5_0),.din(w_dff_A_laAcwvOq2_0),.clk(gclk));
	jdff dff_A_HfW89dTG3_0(.dout(w_dff_A_laAcwvOq2_0),.din(w_dff_A_HfW89dTG3_0),.clk(gclk));
	jdff dff_A_uloYN7lo4_0(.dout(w_dff_A_HfW89dTG3_0),.din(w_dff_A_uloYN7lo4_0),.clk(gclk));
	jdff dff_A_Z1pFR60o7_0(.dout(w_dff_A_uloYN7lo4_0),.din(w_dff_A_Z1pFR60o7_0),.clk(gclk));
	jdff dff_A_gOBFhiLk5_0(.dout(w_dff_A_Z1pFR60o7_0),.din(w_dff_A_gOBFhiLk5_0),.clk(gclk));
	jdff dff_A_Tih0hyYL3_0(.dout(w_dff_A_gOBFhiLk5_0),.din(w_dff_A_Tih0hyYL3_0),.clk(gclk));
	jdff dff_A_YgeUGz0u3_0(.dout(w_dff_A_Tih0hyYL3_0),.din(w_dff_A_YgeUGz0u3_0),.clk(gclk));
	jdff dff_A_952dId8H4_0(.dout(w_dff_A_YgeUGz0u3_0),.din(w_dff_A_952dId8H4_0),.clk(gclk));
	jdff dff_A_drLvg0bw5_0(.dout(w_dff_A_952dId8H4_0),.din(w_dff_A_drLvg0bw5_0),.clk(gclk));
	jdff dff_A_8NgL0byW5_0(.dout(w_G29gat_0[0]),.din(w_dff_A_8NgL0byW5_0),.clk(gclk));
	jdff dff_A_jhBVRKmS9_0(.dout(w_dff_A_8NgL0byW5_0),.din(w_dff_A_jhBVRKmS9_0),.clk(gclk));
	jdff dff_A_ajgQ6ECf4_0(.dout(w_dff_A_jhBVRKmS9_0),.din(w_dff_A_ajgQ6ECf4_0),.clk(gclk));
	jdff dff_A_M3mEFDcA5_0(.dout(w_dff_A_ajgQ6ECf4_0),.din(w_dff_A_M3mEFDcA5_0),.clk(gclk));
	jdff dff_A_xjhhtLpD2_0(.dout(w_dff_A_M3mEFDcA5_0),.din(w_dff_A_xjhhtLpD2_0),.clk(gclk));
	jdff dff_A_lgbpSjju5_0(.dout(w_dff_A_xjhhtLpD2_0),.din(w_dff_A_lgbpSjju5_0),.clk(gclk));
	jdff dff_A_Xf7ek1yO6_0(.dout(w_dff_A_lgbpSjju5_0),.din(w_dff_A_Xf7ek1yO6_0),.clk(gclk));
	jdff dff_A_ZBlzI3ey8_0(.dout(w_dff_A_Xf7ek1yO6_0),.din(w_dff_A_ZBlzI3ey8_0),.clk(gclk));
	jdff dff_A_8fY33f0s7_0(.dout(w_dff_A_ZBlzI3ey8_0),.din(w_dff_A_8fY33f0s7_0),.clk(gclk));
	jdff dff_A_eBECbbOr7_0(.dout(w_dff_A_8fY33f0s7_0),.din(w_dff_A_eBECbbOr7_0),.clk(gclk));
	jdff dff_A_OB7GilfJ9_0(.dout(w_dff_A_eBECbbOr7_0),.din(w_dff_A_OB7GilfJ9_0),.clk(gclk));
	jdff dff_A_PifLK1KF9_0(.dout(w_G50gat_0[0]),.din(w_dff_A_PifLK1KF9_0),.clk(gclk));
	jdff dff_A_lN9CVWBF2_0(.dout(w_dff_A_PifLK1KF9_0),.din(w_dff_A_lN9CVWBF2_0),.clk(gclk));
	jdff dff_A_zcT3cTsb7_0(.dout(w_dff_A_lN9CVWBF2_0),.din(w_dff_A_zcT3cTsb7_0),.clk(gclk));
	jdff dff_A_E5vlx3Ay8_0(.dout(w_dff_A_zcT3cTsb7_0),.din(w_dff_A_E5vlx3Ay8_0),.clk(gclk));
	jdff dff_A_c1PhGR751_0(.dout(w_dff_A_E5vlx3Ay8_0),.din(w_dff_A_c1PhGR751_0),.clk(gclk));
	jdff dff_A_9QnLx7LZ2_0(.dout(w_dff_A_c1PhGR751_0),.din(w_dff_A_9QnLx7LZ2_0),.clk(gclk));
	jdff dff_A_XFIyex0l2_0(.dout(w_dff_A_9QnLx7LZ2_0),.din(w_dff_A_XFIyex0l2_0),.clk(gclk));
	jdff dff_A_OGklGDSh0_0(.dout(w_dff_A_XFIyex0l2_0),.din(w_dff_A_OGklGDSh0_0),.clk(gclk));
	jdff dff_A_n8FL9cNI3_0(.dout(w_dff_A_OGklGDSh0_0),.din(w_dff_A_n8FL9cNI3_0),.clk(gclk));
	jdff dff_A_Cry3SQuq9_0(.dout(w_dff_A_n8FL9cNI3_0),.din(w_dff_A_Cry3SQuq9_0),.clk(gclk));
	jdff dff_A_6CKFAuNy6_0(.dout(w_dff_A_Cry3SQuq9_0),.din(w_dff_A_6CKFAuNy6_0),.clk(gclk));
	jdff dff_A_tKZgqRDz6_0(.dout(w_G43gat_0[0]),.din(w_dff_A_tKZgqRDz6_0),.clk(gclk));
	jdff dff_A_Hr4RJzin2_0(.dout(w_dff_A_tKZgqRDz6_0),.din(w_dff_A_Hr4RJzin2_0),.clk(gclk));
	jdff dff_A_jkxtHo3y3_0(.dout(w_dff_A_Hr4RJzin2_0),.din(w_dff_A_jkxtHo3y3_0),.clk(gclk));
	jdff dff_A_EagGbAgF2_0(.dout(w_dff_A_jkxtHo3y3_0),.din(w_dff_A_EagGbAgF2_0),.clk(gclk));
	jdff dff_A_dBIHdzLw4_0(.dout(w_dff_A_EagGbAgF2_0),.din(w_dff_A_dBIHdzLw4_0),.clk(gclk));
	jdff dff_A_mvr7PKmQ0_0(.dout(w_dff_A_dBIHdzLw4_0),.din(w_dff_A_mvr7PKmQ0_0),.clk(gclk));
	jdff dff_A_vEymCU7L9_0(.dout(w_dff_A_mvr7PKmQ0_0),.din(w_dff_A_vEymCU7L9_0),.clk(gclk));
	jdff dff_A_iVB6eI8q1_0(.dout(w_dff_A_vEymCU7L9_0),.din(w_dff_A_iVB6eI8q1_0),.clk(gclk));
	jdff dff_A_rXxZgoZN9_0(.dout(w_dff_A_iVB6eI8q1_0),.din(w_dff_A_rXxZgoZN9_0),.clk(gclk));
	jdff dff_A_W5moqzen2_0(.dout(w_dff_A_rXxZgoZN9_0),.din(w_dff_A_W5moqzen2_0),.clk(gclk));
	jdff dff_A_EWk6wSym1_0(.dout(w_dff_A_W5moqzen2_0),.din(w_dff_A_EWk6wSym1_0),.clk(gclk));
	jdff dff_A_oghYpZ7M3_0(.dout(w_G92gat_0[0]),.din(w_dff_A_oghYpZ7M3_0),.clk(gclk));
	jdff dff_A_4xUDPzTL8_0(.dout(w_dff_A_oghYpZ7M3_0),.din(w_dff_A_4xUDPzTL8_0),.clk(gclk));
	jdff dff_A_N5jH4jXA9_0(.dout(w_dff_A_4xUDPzTL8_0),.din(w_dff_A_N5jH4jXA9_0),.clk(gclk));
	jdff dff_A_N5Ot1bJF0_0(.dout(w_dff_A_N5jH4jXA9_0),.din(w_dff_A_N5Ot1bJF0_0),.clk(gclk));
	jdff dff_A_33XygtPg9_0(.dout(w_dff_A_N5Ot1bJF0_0),.din(w_dff_A_33XygtPg9_0),.clk(gclk));
	jdff dff_A_e6HsgDU97_0(.dout(w_dff_A_33XygtPg9_0),.din(w_dff_A_e6HsgDU97_0),.clk(gclk));
	jdff dff_A_5qgA06l26_0(.dout(w_dff_A_e6HsgDU97_0),.din(w_dff_A_5qgA06l26_0),.clk(gclk));
	jdff dff_A_4iVMijiM8_0(.dout(w_dff_A_5qgA06l26_0),.din(w_dff_A_4iVMijiM8_0),.clk(gclk));
	jdff dff_A_8jt1bLpO0_0(.dout(w_dff_A_4iVMijiM8_0),.din(w_dff_A_8jt1bLpO0_0),.clk(gclk));
	jdff dff_A_1WTtnRBD1_0(.dout(w_dff_A_8jt1bLpO0_0),.din(w_dff_A_1WTtnRBD1_0),.clk(gclk));
	jdff dff_A_fOGk2Zs59_0(.dout(w_dff_A_1WTtnRBD1_0),.din(w_dff_A_fOGk2Zs59_0),.clk(gclk));
	jdff dff_A_Pxm2Hynp3_0(.dout(w_G85gat_0[0]),.din(w_dff_A_Pxm2Hynp3_0),.clk(gclk));
	jdff dff_A_KIflMu126_0(.dout(w_dff_A_Pxm2Hynp3_0),.din(w_dff_A_KIflMu126_0),.clk(gclk));
	jdff dff_A_9WyYmbh25_0(.dout(w_dff_A_KIflMu126_0),.din(w_dff_A_9WyYmbh25_0),.clk(gclk));
	jdff dff_A_VJFhodmT2_0(.dout(w_dff_A_9WyYmbh25_0),.din(w_dff_A_VJFhodmT2_0),.clk(gclk));
	jdff dff_A_5cf0d9z87_0(.dout(w_dff_A_VJFhodmT2_0),.din(w_dff_A_5cf0d9z87_0),.clk(gclk));
	jdff dff_A_v9i7mDaN7_0(.dout(w_dff_A_5cf0d9z87_0),.din(w_dff_A_v9i7mDaN7_0),.clk(gclk));
	jdff dff_A_7cCj6nXZ7_0(.dout(w_dff_A_v9i7mDaN7_0),.din(w_dff_A_7cCj6nXZ7_0),.clk(gclk));
	jdff dff_A_yQ2U1kXz8_0(.dout(w_dff_A_7cCj6nXZ7_0),.din(w_dff_A_yQ2U1kXz8_0),.clk(gclk));
	jdff dff_A_Z5xDBAup9_0(.dout(w_dff_A_yQ2U1kXz8_0),.din(w_dff_A_Z5xDBAup9_0),.clk(gclk));
	jdff dff_A_9v7HP2XB4_0(.dout(w_dff_A_Z5xDBAup9_0),.din(w_dff_A_9v7HP2XB4_0),.clk(gclk));
	jdff dff_A_ScOY6LQa6_0(.dout(w_dff_A_9v7HP2XB4_0),.din(w_dff_A_ScOY6LQa6_0),.clk(gclk));
	jdff dff_A_ptDHawF33_0(.dout(w_G106gat_0[0]),.din(w_dff_A_ptDHawF33_0),.clk(gclk));
	jdff dff_A_LlqxGvMB3_0(.dout(w_dff_A_ptDHawF33_0),.din(w_dff_A_LlqxGvMB3_0),.clk(gclk));
	jdff dff_A_3bjSki6M1_0(.dout(w_dff_A_LlqxGvMB3_0),.din(w_dff_A_3bjSki6M1_0),.clk(gclk));
	jdff dff_A_XMDCLix27_0(.dout(w_dff_A_3bjSki6M1_0),.din(w_dff_A_XMDCLix27_0),.clk(gclk));
	jdff dff_A_0nrKv9xc9_0(.dout(w_dff_A_XMDCLix27_0),.din(w_dff_A_0nrKv9xc9_0),.clk(gclk));
	jdff dff_A_CqkDwW2h5_0(.dout(w_dff_A_0nrKv9xc9_0),.din(w_dff_A_CqkDwW2h5_0),.clk(gclk));
	jdff dff_A_avvZpOWE5_0(.dout(w_dff_A_CqkDwW2h5_0),.din(w_dff_A_avvZpOWE5_0),.clk(gclk));
	jdff dff_A_AurYlREi0_0(.dout(w_dff_A_avvZpOWE5_0),.din(w_dff_A_AurYlREi0_0),.clk(gclk));
	jdff dff_A_qcu5Rdl66_0(.dout(w_dff_A_AurYlREi0_0),.din(w_dff_A_qcu5Rdl66_0),.clk(gclk));
	jdff dff_A_iHtSzie08_0(.dout(w_dff_A_qcu5Rdl66_0),.din(w_dff_A_iHtSzie08_0),.clk(gclk));
	jdff dff_A_1TLSdQqz3_0(.dout(w_dff_A_iHtSzie08_0),.din(w_dff_A_1TLSdQqz3_0),.clk(gclk));
	jdff dff_A_qbVd0D6m1_0(.dout(w_G99gat_0[0]),.din(w_dff_A_qbVd0D6m1_0),.clk(gclk));
	jdff dff_A_ekdPj6c14_0(.dout(w_dff_A_qbVd0D6m1_0),.din(w_dff_A_ekdPj6c14_0),.clk(gclk));
	jdff dff_A_Qs8IxPQU4_0(.dout(w_dff_A_ekdPj6c14_0),.din(w_dff_A_Qs8IxPQU4_0),.clk(gclk));
	jdff dff_A_zG7HLKGw9_0(.dout(w_dff_A_Qs8IxPQU4_0),.din(w_dff_A_zG7HLKGw9_0),.clk(gclk));
	jdff dff_A_JAZzS8LO5_0(.dout(w_dff_A_zG7HLKGw9_0),.din(w_dff_A_JAZzS8LO5_0),.clk(gclk));
	jdff dff_A_aRgEUGVX7_0(.dout(w_dff_A_JAZzS8LO5_0),.din(w_dff_A_aRgEUGVX7_0),.clk(gclk));
	jdff dff_A_MWMyUdxS1_0(.dout(w_dff_A_aRgEUGVX7_0),.din(w_dff_A_MWMyUdxS1_0),.clk(gclk));
	jdff dff_A_asTS1FeR3_0(.dout(w_dff_A_MWMyUdxS1_0),.din(w_dff_A_asTS1FeR3_0),.clk(gclk));
	jdff dff_A_wxeVzPs08_0(.dout(w_dff_A_asTS1FeR3_0),.din(w_dff_A_wxeVzPs08_0),.clk(gclk));
	jdff dff_A_7rpyD8io6_0(.dout(w_dff_A_wxeVzPs08_0),.din(w_dff_A_7rpyD8io6_0),.clk(gclk));
	jdff dff_A_qsVz5g8R4_0(.dout(w_dff_A_7rpyD8io6_0),.din(w_dff_A_qsVz5g8R4_0),.clk(gclk));
	jdff dff_A_8SAwAT9O2_0(.dout(w_G162gat_0[0]),.din(w_dff_A_8SAwAT9O2_0),.clk(gclk));
	jdff dff_A_VWJb7aaj1_0(.dout(w_dff_A_8SAwAT9O2_0),.din(w_dff_A_VWJb7aaj1_0),.clk(gclk));
	jdff dff_A_uYZ9ddvD0_0(.dout(w_dff_A_VWJb7aaj1_0),.din(w_dff_A_uYZ9ddvD0_0),.clk(gclk));
	jdff dff_A_lH4RvTb54_0(.dout(w_dff_A_uYZ9ddvD0_0),.din(w_dff_A_lH4RvTb54_0),.clk(gclk));
	jdff dff_A_5PlTz9Gj5_0(.dout(w_dff_A_lH4RvTb54_0),.din(w_dff_A_5PlTz9Gj5_0),.clk(gclk));
	jdff dff_A_7OnIDFpU2_0(.dout(w_dff_A_5PlTz9Gj5_0),.din(w_dff_A_7OnIDFpU2_0),.clk(gclk));
	jdff dff_A_6iyMxZ369_0(.dout(w_dff_A_7OnIDFpU2_0),.din(w_dff_A_6iyMxZ369_0),.clk(gclk));
	jdff dff_A_0Hk51g9W6_0(.dout(w_dff_A_6iyMxZ369_0),.din(w_dff_A_0Hk51g9W6_0),.clk(gclk));
	jdff dff_A_XylOKzOO5_0(.dout(w_dff_A_0Hk51g9W6_0),.din(w_dff_A_XylOKzOO5_0),.clk(gclk));
	jdff dff_A_9kXPIB2g0_0(.dout(w_dff_A_XylOKzOO5_0),.din(w_dff_A_9kXPIB2g0_0),.clk(gclk));
	jdff dff_A_M94Wx5ES3_0(.dout(w_dff_A_9kXPIB2g0_0),.din(w_dff_A_M94Wx5ES3_0),.clk(gclk));
	jdff dff_A_6FqbQmRT9_0(.dout(w_G134gat_0[0]),.din(w_dff_A_6FqbQmRT9_0),.clk(gclk));
	jdff dff_A_moTWRqlj4_0(.dout(w_dff_A_6FqbQmRT9_0),.din(w_dff_A_moTWRqlj4_0),.clk(gclk));
	jdff dff_A_ydDsvXT58_0(.dout(w_dff_A_moTWRqlj4_0),.din(w_dff_A_ydDsvXT58_0),.clk(gclk));
	jdff dff_A_d7lTRz1w1_0(.dout(w_dff_A_ydDsvXT58_0),.din(w_dff_A_d7lTRz1w1_0),.clk(gclk));
	jdff dff_A_S6I0eFoT7_0(.dout(w_dff_A_d7lTRz1w1_0),.din(w_dff_A_S6I0eFoT7_0),.clk(gclk));
	jdff dff_A_6S06bhx94_0(.dout(w_dff_A_S6I0eFoT7_0),.din(w_dff_A_6S06bhx94_0),.clk(gclk));
	jdff dff_A_o1QY7sx44_0(.dout(w_dff_A_6S06bhx94_0),.din(w_dff_A_o1QY7sx44_0),.clk(gclk));
	jdff dff_A_XtmNMhD51_0(.dout(w_dff_A_o1QY7sx44_0),.din(w_dff_A_XtmNMhD51_0),.clk(gclk));
	jdff dff_A_nQYkzxOf3_0(.dout(w_dff_A_XtmNMhD51_0),.din(w_dff_A_nQYkzxOf3_0),.clk(gclk));
	jdff dff_A_IjZ9WPvP0_0(.dout(w_dff_A_nQYkzxOf3_0),.din(w_dff_A_IjZ9WPvP0_0),.clk(gclk));
	jdff dff_A_vKv8bSYv9_0(.dout(w_dff_A_IjZ9WPvP0_0),.din(w_dff_A_vKv8bSYv9_0),.clk(gclk));
	jdff dff_A_deLr8FPU4_0(.dout(w_G218gat_0[0]),.din(w_dff_A_deLr8FPU4_0),.clk(gclk));
	jdff dff_A_wxcsNfRJ6_0(.dout(w_dff_A_deLr8FPU4_0),.din(w_dff_A_wxcsNfRJ6_0),.clk(gclk));
	jdff dff_A_Ckrg3HfM2_0(.dout(w_dff_A_wxcsNfRJ6_0),.din(w_dff_A_Ckrg3HfM2_0),.clk(gclk));
	jdff dff_A_3tq7bs351_0(.dout(w_dff_A_Ckrg3HfM2_0),.din(w_dff_A_3tq7bs351_0),.clk(gclk));
	jdff dff_A_m43anPMI1_0(.dout(w_dff_A_3tq7bs351_0),.din(w_dff_A_m43anPMI1_0),.clk(gclk));
	jdff dff_A_YT6aLnYY2_0(.dout(w_dff_A_m43anPMI1_0),.din(w_dff_A_YT6aLnYY2_0),.clk(gclk));
	jdff dff_A_pkKkitfx9_0(.dout(w_dff_A_YT6aLnYY2_0),.din(w_dff_A_pkKkitfx9_0),.clk(gclk));
	jdff dff_A_iIiGKZl39_0(.dout(w_dff_A_pkKkitfx9_0),.din(w_dff_A_iIiGKZl39_0),.clk(gclk));
	jdff dff_A_F1eypsoi6_0(.dout(w_dff_A_iIiGKZl39_0),.din(w_dff_A_F1eypsoi6_0),.clk(gclk));
	jdff dff_A_sRof27eR9_0(.dout(w_dff_A_F1eypsoi6_0),.din(w_dff_A_sRof27eR9_0),.clk(gclk));
	jdff dff_A_jkYTbfyn8_0(.dout(w_dff_A_sRof27eR9_0),.din(w_dff_A_jkYTbfyn8_0),.clk(gclk));
	jdff dff_A_FapeOVY95_0(.dout(w_G190gat_0[0]),.din(w_dff_A_FapeOVY95_0),.clk(gclk));
	jdff dff_A_uK1a1sii7_0(.dout(w_dff_A_FapeOVY95_0),.din(w_dff_A_uK1a1sii7_0),.clk(gclk));
	jdff dff_A_FqwzPC3E8_0(.dout(w_dff_A_uK1a1sii7_0),.din(w_dff_A_FqwzPC3E8_0),.clk(gclk));
	jdff dff_A_WtTdz0lC0_0(.dout(w_dff_A_FqwzPC3E8_0),.din(w_dff_A_WtTdz0lC0_0),.clk(gclk));
	jdff dff_A_PxWIvayd9_0(.dout(w_dff_A_WtTdz0lC0_0),.din(w_dff_A_PxWIvayd9_0),.clk(gclk));
	jdff dff_A_HIZilLLr7_0(.dout(w_dff_A_PxWIvayd9_0),.din(w_dff_A_HIZilLLr7_0),.clk(gclk));
	jdff dff_A_metjIlrp0_0(.dout(w_dff_A_HIZilLLr7_0),.din(w_dff_A_metjIlrp0_0),.clk(gclk));
	jdff dff_A_fMsTXQ4I3_0(.dout(w_dff_A_metjIlrp0_0),.din(w_dff_A_fMsTXQ4I3_0),.clk(gclk));
	jdff dff_A_zZHpXqXw9_0(.dout(w_dff_A_fMsTXQ4I3_0),.din(w_dff_A_zZHpXqXw9_0),.clk(gclk));
	jdff dff_A_ioNA677y0_0(.dout(w_dff_A_zZHpXqXw9_0),.din(w_dff_A_ioNA677y0_0),.clk(gclk));
	jdff dff_A_KQTvHfr49_0(.dout(w_dff_A_ioNA677y0_0),.din(w_dff_A_KQTvHfr49_0),.clk(gclk));
endmodule

