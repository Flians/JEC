/*

c5315:
	jxor: 109
	jspl: 308
	jspl3: 385
	jnot: 226
	jcb: 419
	jdff: 2028
	jand: 605

Summary:
	jxor: 109
	jspl: 308
	jspl3: 385
	jnot: 226
	jcb: 419
	jdff: 2028
	jand: 605
*/

module c5315(gclk, G1, G4, G11, G14, G17, G20, G23, G24, G25, G26, G27, G31, G34, G37, G40, G43, G46, G49, G52, G53, G54, G61, G64, G67, G70, G73, G76, G79, G80, G81, G82, G83, G86, G87, G88, G91, G94, G97, G100, G103, G106, G109, G112, G113, G114, G115, G116, G117, G118, G119, G120, G121, G122, G123, G126, G127, G128, G129, G130, G131, G132, G135, G136, G137, G140, G141, G145, G146, G149, G152, G155, G158, G161, G164, G167, G170, G173, G176, G179, G182, G185, G188, G191, G194, G197, G200, G203, G206, G209, G210, G217, G218, G225, G226, G233, G234, G241, G242, G245, G248, G251, G254, G257, G264, G265, G272, G273, G280, G281, G288, G289, G292, G293, G299, G302, G307, G308, G315, G316, G323, G324, G331, G332, G335, G338, G341, G348, G351, G358, G361, G366, G369, G372, G373, G374, G386, G389, G400, G411, G422, G435, G446, G457, G468, G479, G490, G503, G514, G523, G534, G545, G549, G552, G556, G559, G562, G1497, G1689, G1690, G1691, G1694, G2174, G2358, G2824, G3173, G3546, G3548, G3550, G3552, G3717, G3724, G4087, G4088, G4089, G4090, G4091, G4092, G4115, G144, G298, G973, G594, G599, G600, G601, G602, G603, G604, G611, G612, G810, G848, G849, G850, G851, G634, G815, G845, G847, G926, G923, G921, G892, G887, G606, G656, G809, G993, G978, G949, G939, G889, G593, G636, G704, G717, G820, G639, G673, G707, G715, G598, G610, G588, G615, G626, G632, G1002, G1004, G591, G618, G621, G629, G822, G838, G861, G623, G722, G832, G834, G836, G859, G871, G873, G875, G877, G998, G1000, G575, G585, G661, G693, G747, G752, G757, G762, G787, G792, G797, G802, G642, G664, G667, G670, G676, G696, G699, G702, G818, G813, G824, G826, G828, G830, G854, G863, G865, G867, G869, G712, G727, G732, G737, G742, G772, G777, G782, G645, G648, G651, G654, G679, G682, G685, G688, G843, G882, G767, G807, G658, G690);
	input gclk;
	input G1;
	input G4;
	input G11;
	input G14;
	input G17;
	input G20;
	input G23;
	input G24;
	input G25;
	input G26;
	input G27;
	input G31;
	input G34;
	input G37;
	input G40;
	input G43;
	input G46;
	input G49;
	input G52;
	input G53;
	input G54;
	input G61;
	input G64;
	input G67;
	input G70;
	input G73;
	input G76;
	input G79;
	input G80;
	input G81;
	input G82;
	input G83;
	input G86;
	input G87;
	input G88;
	input G91;
	input G94;
	input G97;
	input G100;
	input G103;
	input G106;
	input G109;
	input G112;
	input G113;
	input G114;
	input G115;
	input G116;
	input G117;
	input G118;
	input G119;
	input G120;
	input G121;
	input G122;
	input G123;
	input G126;
	input G127;
	input G128;
	input G129;
	input G130;
	input G131;
	input G132;
	input G135;
	input G136;
	input G137;
	input G140;
	input G141;
	input G145;
	input G146;
	input G149;
	input G152;
	input G155;
	input G158;
	input G161;
	input G164;
	input G167;
	input G170;
	input G173;
	input G176;
	input G179;
	input G182;
	input G185;
	input G188;
	input G191;
	input G194;
	input G197;
	input G200;
	input G203;
	input G206;
	input G209;
	input G210;
	input G217;
	input G218;
	input G225;
	input G226;
	input G233;
	input G234;
	input G241;
	input G242;
	input G245;
	input G248;
	input G251;
	input G254;
	input G257;
	input G264;
	input G265;
	input G272;
	input G273;
	input G280;
	input G281;
	input G288;
	input G289;
	input G292;
	input G293;
	input G299;
	input G302;
	input G307;
	input G308;
	input G315;
	input G316;
	input G323;
	input G324;
	input G331;
	input G332;
	input G335;
	input G338;
	input G341;
	input G348;
	input G351;
	input G358;
	input G361;
	input G366;
	input G369;
	input G372;
	input G373;
	input G374;
	input G386;
	input G389;
	input G400;
	input G411;
	input G422;
	input G435;
	input G446;
	input G457;
	input G468;
	input G479;
	input G490;
	input G503;
	input G514;
	input G523;
	input G534;
	input G545;
	input G549;
	input G552;
	input G556;
	input G559;
	input G562;
	input G1497;
	input G1689;
	input G1690;
	input G1691;
	input G1694;
	input G2174;
	input G2358;
	input G2824;
	input G3173;
	input G3546;
	input G3548;
	input G3550;
	input G3552;
	input G3717;
	input G3724;
	input G4087;
	input G4088;
	input G4089;
	input G4090;
	input G4091;
	input G4092;
	input G4115;
	output G144;
	output G298;
	output G973;
	output G594;
	output G599;
	output G600;
	output G601;
	output G602;
	output G603;
	output G604;
	output G611;
	output G612;
	output G810;
	output G848;
	output G849;
	output G850;
	output G851;
	output G634;
	output G815;
	output G845;
	output G847;
	output G926;
	output G923;
	output G921;
	output G892;
	output G887;
	output G606;
	output G656;
	output G809;
	output G993;
	output G978;
	output G949;
	output G939;
	output G889;
	output G593;
	output G636;
	output G704;
	output G717;
	output G820;
	output G639;
	output G673;
	output G707;
	output G715;
	output G598;
	output G610;
	output G588;
	output G615;
	output G626;
	output G632;
	output G1002;
	output G1004;
	output G591;
	output G618;
	output G621;
	output G629;
	output G822;
	output G838;
	output G861;
	output G623;
	output G722;
	output G832;
	output G834;
	output G836;
	output G859;
	output G871;
	output G873;
	output G875;
	output G877;
	output G998;
	output G1000;
	output G575;
	output G585;
	output G661;
	output G693;
	output G747;
	output G752;
	output G757;
	output G762;
	output G787;
	output G792;
	output G797;
	output G802;
	output G642;
	output G664;
	output G667;
	output G670;
	output G676;
	output G696;
	output G699;
	output G702;
	output G818;
	output G813;
	output G824;
	output G826;
	output G828;
	output G830;
	output G854;
	output G863;
	output G865;
	output G867;
	output G869;
	output G712;
	output G727;
	output G732;
	output G737;
	output G742;
	output G772;
	output G777;
	output G782;
	output G645;
	output G648;
	output G651;
	output G654;
	output G679;
	output G682;
	output G685;
	output G688;
	output G843;
	output G882;
	output G767;
	output G807;
	output G658;
	output G690;
	wire n314;
	wire n316;
	wire n318;
	wire n320;
	wire n321;
	wire n325;
	wire n326;
	wire n327;
	wire n328;
	wire n329;
	wire n330;
	wire n332;
	wire n333;
	wire n334;
	wire n335;
	wire n336;
	wire n338;
	wire n340;
	wire n341;
	wire n342;
	wire n343;
	wire n345;
	wire n346;
	wire n347;
	wire n348;
	wire n350;
	wire n351;
	wire n352;
	wire n353;
	wire n355;
	wire n356;
	wire n357;
	wire n358;
	wire n360;
	wire n361;
	wire n362;
	wire n363;
	wire n364;
	wire n365;
	wire n366;
	wire n367;
	wire n368;
	wire n369;
	wire n370;
	wire n371;
	wire n372;
	wire n373;
	wire n374;
	wire n375;
	wire n376;
	wire n377;
	wire n378;
	wire n379;
	wire n380;
	wire n381;
	wire n382;
	wire n383;
	wire n384;
	wire n385;
	wire n386;
	wire n387;
	wire n388;
	wire n389;
	wire n390;
	wire n391;
	wire n392;
	wire n393;
	wire n394;
	wire n395;
	wire n396;
	wire n397;
	wire n398;
	wire n399;
	wire n400;
	wire n401;
	wire n402;
	wire n403;
	wire n404;
	wire n405;
	wire n406;
	wire n407;
	wire n408;
	wire n409;
	wire n410;
	wire n411;
	wire n412;
	wire n413;
	wire n414;
	wire n415;
	wire n416;
	wire n417;
	wire n418;
	wire n419;
	wire n420;
	wire n421;
	wire n422;
	wire n423;
	wire n424;
	wire n425;
	wire n426;
	wire n427;
	wire n428;
	wire n429;
	wire n430;
	wire n431;
	wire n432;
	wire n433;
	wire n434;
	wire n435;
	wire n436;
	wire n437;
	wire n438;
	wire n439;
	wire n440;
	wire n441;
	wire n442;
	wire n443;
	wire n444;
	wire n445;
	wire n446;
	wire n447;
	wire n449;
	wire n450;
	wire n451;
	wire n452;
	wire n453;
	wire n454;
	wire n455;
	wire n456;
	wire n457;
	wire n458;
	wire n459;
	wire n460;
	wire n461;
	wire n462;
	wire n463;
	wire n464;
	wire n465;
	wire n466;
	wire n467;
	wire n468;
	wire n469;
	wire n470;
	wire n471;
	wire n472;
	wire n473;
	wire n474;
	wire n475;
	wire n476;
	wire n477;
	wire n478;
	wire n479;
	wire n480;
	wire n481;
	wire n482;
	wire n483;
	wire n484;
	wire n485;
	wire n486;
	wire n487;
	wire n488;
	wire n489;
	wire n490;
	wire n491;
	wire n492;
	wire n493;
	wire n494;
	wire n495;
	wire n496;
	wire n497;
	wire n498;
	wire n499;
	wire n500;
	wire n501;
	wire n502;
	wire n503;
	wire n504;
	wire n505;
	wire n506;
	wire n507;
	wire n508;
	wire n509;
	wire n510;
	wire n511;
	wire n512;
	wire n513;
	wire n514;
	wire n515;
	wire n516;
	wire n517;
	wire n518;
	wire n519;
	wire n520;
	wire n521;
	wire n522;
	wire n523;
	wire n524;
	wire n525;
	wire n526;
	wire n527;
	wire n528;
	wire n529;
	wire n530;
	wire n531;
	wire n532;
	wire n533;
	wire n534;
	wire n535;
	wire n536;
	wire n537;
	wire n538;
	wire n539;
	wire n540;
	wire n541;
	wire n542;
	wire n543;
	wire n544;
	wire n545;
	wire n546;
	wire n547;
	wire n548;
	wire n549;
	wire n550;
	wire n551;
	wire n552;
	wire n553;
	wire n554;
	wire n556;
	wire n557;
	wire n558;
	wire n559;
	wire n560;
	wire n561;
	wire n562;
	wire n563;
	wire n564;
	wire n565;
	wire n566;
	wire n567;
	wire n568;
	wire n569;
	wire n570;
	wire n571;
	wire n572;
	wire n573;
	wire n574;
	wire n575;
	wire n576;
	wire n577;
	wire n578;
	wire n579;
	wire n580;
	wire n581;
	wire n582;
	wire n583;
	wire n584;
	wire n585;
	wire n586;
	wire n587;
	wire n588;
	wire n589;
	wire n590;
	wire n591;
	wire n592;
	wire n593;
	wire n594;
	wire n595;
	wire n596;
	wire n597;
	wire n598;
	wire n599;
	wire n600;
	wire n601;
	wire n602;
	wire n603;
	wire n604;
	wire n605;
	wire n606;
	wire n607;
	wire n609;
	wire n610;
	wire n611;
	wire n612;
	wire n613;
	wire n614;
	wire n615;
	wire n616;
	wire n617;
	wire n618;
	wire n619;
	wire n620;
	wire n621;
	wire n622;
	wire n623;
	wire n624;
	wire n625;
	wire n626;
	wire n627;
	wire n628;
	wire n629;
	wire n630;
	wire n631;
	wire n632;
	wire n633;
	wire n634;
	wire n635;
	wire n636;
	wire n637;
	wire n638;
	wire n639;
	wire n640;
	wire n641;
	wire n642;
	wire n643;
	wire n644;
	wire n645;
	wire n646;
	wire n647;
	wire n648;
	wire n649;
	wire n650;
	wire n651;
	wire n652;
	wire n654;
	wire n655;
	wire n656;
	wire n657;
	wire n658;
	wire n659;
	wire n660;
	wire n661;
	wire n663;
	wire n664;
	wire n665;
	wire n666;
	wire n667;
	wire n668;
	wire n669;
	wire n670;
	wire n671;
	wire n673;
	wire n674;
	wire n675;
	wire n676;
	wire n677;
	wire n678;
	wire n679;
	wire n680;
	wire n681;
	wire n682;
	wire n683;
	wire n684;
	wire n685;
	wire n686;
	wire n687;
	wire n688;
	wire n689;
	wire n690;
	wire n691;
	wire n692;
	wire n693;
	wire n694;
	wire n695;
	wire n696;
	wire n697;
	wire n698;
	wire n699;
	wire n700;
	wire n701;
	wire n702;
	wire n703;
	wire n704;
	wire n705;
	wire n706;
	wire n707;
	wire n708;
	wire n709;
	wire n711;
	wire n712;
	wire n713;
	wire n714;
	wire n715;
	wire n716;
	wire n717;
	wire n718;
	wire n719;
	wire n720;
	wire n721;
	wire n722;
	wire n723;
	wire n724;
	wire n725;
	wire n726;
	wire n727;
	wire n728;
	wire n729;
	wire n730;
	wire n731;
	wire n732;
	wire n733;
	wire n734;
	wire n735;
	wire n736;
	wire n737;
	wire n738;
	wire n739;
	wire n740;
	wire n741;
	wire n742;
	wire n744;
	wire n745;
	wire n746;
	wire n747;
	wire n748;
	wire n749;
	wire n750;
	wire n751;
	wire n752;
	wire n753;
	wire n754;
	wire n755;
	wire n756;
	wire n758;
	wire n759;
	wire n760;
	wire n761;
	wire n762;
	wire n763;
	wire n764;
	wire n765;
	wire n766;
	wire n767;
	wire n768;
	wire n769;
	wire n771;
	wire n772;
	wire n773;
	wire n774;
	wire n775;
	wire n776;
	wire n777;
	wire n779;
	wire n780;
	wire n781;
	wire n782;
	wire n783;
	wire n784;
	wire n785;
	wire n786;
	wire n787;
	wire n788;
	wire n789;
	wire n791;
	wire n792;
	wire n793;
	wire n794;
	wire n795;
	wire n796;
	wire n797;
	wire n798;
	wire n799;
	wire n800;
	wire n801;
	wire n802;
	wire n803;
	wire n804;
	wire n806;
	wire n807;
	wire n808;
	wire n809;
	wire n810;
	wire n811;
	wire n812;
	wire n813;
	wire n814;
	wire n816;
	wire n817;
	wire n818;
	wire n819;
	wire n820;
	wire n821;
	wire n822;
	wire n823;
	wire n824;
	wire n825;
	wire n826;
	wire n828;
	wire n829;
	wire n830;
	wire n831;
	wire n832;
	wire n833;
	wire n834;
	wire n835;
	wire n836;
	wire n837;
	wire n839;
	wire n840;
	wire n841;
	wire n842;
	wire n843;
	wire n844;
	wire n845;
	wire n846;
	wire n847;
	wire n848;
	wire n849;
	wire n850;
	wire n852;
	wire n853;
	wire n854;
	wire n855;
	wire n856;
	wire n857;
	wire n858;
	wire n859;
	wire n860;
	wire n861;
	wire n862;
	wire n863;
	wire n864;
	wire n865;
	wire n866;
	wire n867;
	wire n869;
	wire n870;
	wire n871;
	wire n872;
	wire n873;
	wire n874;
	wire n876;
	wire n877;
	wire n878;
	wire n879;
	wire n880;
	wire n881;
	wire n882;
	wire n883;
	wire n884;
	wire n885;
	wire n886;
	wire n887;
	wire n889;
	wire n890;
	wire n891;
	wire n892;
	wire n893;
	wire n894;
	wire n895;
	wire n896;
	wire n897;
	wire n898;
	wire n900;
	wire n901;
	wire n902;
	wire n903;
	wire n904;
	wire n905;
	wire n906;
	wire n907;
	wire n908;
	wire n909;
	wire n910;
	wire n911;
	wire n912;
	wire n913;
	wire n914;
	wire n916;
	wire n917;
	wire n918;
	wire n919;
	wire n920;
	wire n921;
	wire n922;
	wire n923;
	wire n924;
	wire n925;
	wire n926;
	wire n928;
	wire n929;
	wire n930;
	wire n931;
	wire n932;
	wire n933;
	wire n934;
	wire n935;
	wire n936;
	wire n937;
	wire n938;
	wire n939;
	wire n940;
	wire n941;
	wire n942;
	wire n943;
	wire n944;
	wire n945;
	wire n946;
	wire n947;
	wire n948;
	wire n949;
	wire n950;
	wire n951;
	wire n952;
	wire n953;
	wire n954;
	wire n955;
	wire n956;
	wire n957;
	wire n958;
	wire n959;
	wire n960;
	wire n961;
	wire n962;
	wire n963;
	wire n964;
	wire n965;
	wire n967;
	wire n968;
	wire n969;
	wire n970;
	wire n971;
	wire n972;
	wire n973;
	wire n974;
	wire n975;
	wire n976;
	wire n977;
	wire n978;
	wire n979;
	wire n980;
	wire n981;
	wire n982;
	wire n984;
	wire n985;
	wire n986;
	wire n987;
	wire n988;
	wire n989;
	wire n990;
	wire n991;
	wire n992;
	wire n993;
	wire n994;
	wire n995;
	wire n996;
	wire n998;
	wire n999;
	wire n1000;
	wire n1001;
	wire n1002;
	wire n1003;
	wire n1004;
	wire n1005;
	wire n1006;
	wire n1007;
	wire n1008;
	wire n1009;
	wire n1010;
	wire n1012;
	wire n1013;
	wire n1014;
	wire n1015;
	wire n1016;
	wire n1017;
	wire n1018;
	wire n1019;
	wire n1021;
	wire n1022;
	wire n1023;
	wire n1024;
	wire n1025;
	wire n1026;
	wire n1027;
	wire n1028;
	wire n1030;
	wire n1031;
	wire n1032;
	wire n1033;
	wire n1034;
	wire n1035;
	wire n1036;
	wire n1037;
	wire n1039;
	wire n1040;
	wire n1041;
	wire n1042;
	wire n1043;
	wire n1044;
	wire n1045;
	wire n1046;
	wire n1048;
	wire n1049;
	wire n1050;
	wire n1051;
	wire n1052;
	wire n1053;
	wire n1055;
	wire n1056;
	wire n1057;
	wire n1058;
	wire n1059;
	wire n1060;
	wire n1062;
	wire n1063;
	wire n1064;
	wire n1065;
	wire n1066;
	wire n1067;
	wire n1069;
	wire n1070;
	wire n1071;
	wire n1072;
	wire n1073;
	wire n1074;
	wire n1076;
	wire n1077;
	wire n1078;
	wire n1079;
	wire n1080;
	wire n1081;
	wire n1082;
	wire n1084;
	wire n1085;
	wire n1086;
	wire n1087;
	wire n1088;
	wire n1089;
	wire n1090;
	wire n1092;
	wire n1093;
	wire n1094;
	wire n1095;
	wire n1096;
	wire n1097;
	wire n1098;
	wire n1100;
	wire n1101;
	wire n1102;
	wire n1103;
	wire n1104;
	wire n1105;
	wire n1106;
	wire n1108;
	wire n1109;
	wire n1110;
	wire n1111;
	wire n1112;
	wire n1113;
	wire n1114;
	wire n1116;
	wire n1117;
	wire n1118;
	wire n1119;
	wire n1120;
	wire n1121;
	wire n1122;
	wire n1124;
	wire n1125;
	wire n1126;
	wire n1127;
	wire n1128;
	wire n1129;
	wire n1130;
	wire n1132;
	wire n1133;
	wire n1134;
	wire n1135;
	wire n1136;
	wire n1137;
	wire n1138;
	wire n1140;
	wire n1141;
	wire n1142;
	wire n1143;
	wire n1144;
	wire n1145;
	wire n1146;
	wire n1147;
	wire n1148;
	wire n1149;
	wire n1150;
	wire n1151;
	wire n1152;
	wire n1153;
	wire n1154;
	wire n1155;
	wire n1157;
	wire n1159;
	wire n1160;
	wire n1161;
	wire n1162;
	wire n1163;
	wire n1165;
	wire n1166;
	wire n1167;
	wire n1168;
	wire n1169;
	wire n1171;
	wire n1172;
	wire n1173;
	wire n1174;
	wire n1175;
	wire n1177;
	wire n1178;
	wire n1179;
	wire n1180;
	wire n1181;
	wire n1182;
	wire n1184;
	wire n1185;
	wire n1186;
	wire n1187;
	wire n1188;
	wire n1189;
	wire n1190;
	wire n1192;
	wire n1193;
	wire n1194;
	wire n1195;
	wire n1196;
	wire n1197;
	wire n1199;
	wire n1200;
	wire n1201;
	wire n1202;
	wire n1203;
	wire n1204;
	wire n1205;
	wire n1207;
	wire n1208;
	wire n1209;
	wire n1210;
	wire n1211;
	wire n1213;
	wire n1214;
	wire n1215;
	wire n1216;
	wire n1217;
	wire n1218;
	wire n1220;
	wire n1221;
	wire n1222;
	wire n1223;
	wire n1224;
	wire n1225;
	wire n1227;
	wire n1228;
	wire n1229;
	wire n1230;
	wire n1231;
	wire n1232;
	wire n1234;
	wire n1235;
	wire n1236;
	wire n1237;
	wire n1238;
	wire n1239;
	wire n1240;
	wire n1242;
	wire n1243;
	wire n1244;
	wire n1245;
	wire n1246;
	wire n1247;
	wire n1248;
	wire n1249;
	wire n1251;
	wire n1252;
	wire n1253;
	wire n1254;
	wire n1255;
	wire n1256;
	wire n1257;
	wire n1258;
	wire n1260;
	wire n1261;
	wire n1262;
	wire n1263;
	wire n1264;
	wire n1265;
	wire n1267;
	wire n1268;
	wire n1269;
	wire n1270;
	wire n1271;
	wire n1272;
	wire n1274;
	wire n1275;
	wire n1276;
	wire n1277;
	wire n1278;
	wire n1279;
	wire n1281;
	wire n1282;
	wire n1283;
	wire n1284;
	wire n1285;
	wire n1286;
	wire n1287;
	wire n1289;
	wire n1290;
	wire n1291;
	wire n1292;
	wire n1293;
	wire n1294;
	wire n1295;
	wire n1297;
	wire n1298;
	wire n1299;
	wire n1300;
	wire n1301;
	wire n1302;
	wire n1303;
	wire n1305;
	wire n1306;
	wire n1307;
	wire n1308;
	wire n1309;
	wire n1310;
	wire n1311;
	wire n1313;
	wire n1314;
	wire n1315;
	wire n1316;
	wire n1317;
	wire n1318;
	wire n1319;
	wire n1321;
	wire n1322;
	wire n1323;
	wire n1324;
	wire n1325;
	wire n1326;
	wire n1327;
	wire n1329;
	wire n1330;
	wire n1331;
	wire n1332;
	wire n1333;
	wire n1334;
	wire n1335;
	wire n1337;
	wire n1338;
	wire n1339;
	wire n1340;
	wire n1341;
	wire n1342;
	wire n1343;
	wire n1345;
	wire n1346;
	wire n1347;
	wire n1348;
	wire n1349;
	wire n1350;
	wire n1351;
	wire n1352;
	wire n1353;
	wire n1354;
	wire n1355;
	wire n1356;
	wire n1357;
	wire n1358;
	wire n1359;
	wire n1360;
	wire n1361;
	wire n1362;
	wire n1363;
	wire n1364;
	wire n1365;
	wire n1366;
	wire n1367;
	wire n1368;
	wire n1369;
	wire n1370;
	wire n1371;
	wire n1372;
	wire n1373;
	wire n1374;
	wire n1375;
	wire n1376;
	wire n1377;
	wire n1378;
	wire n1379;
	wire n1380;
	wire n1381;
	wire n1382;
	wire n1383;
	wire n1384;
	wire n1385;
	wire n1386;
	wire n1388;
	wire n1389;
	wire n1390;
	wire n1391;
	wire n1392;
	wire n1393;
	wire n1394;
	wire n1395;
	wire n1396;
	wire n1397;
	wire n1398;
	wire n1399;
	wire n1400;
	wire n1401;
	wire n1402;
	wire n1403;
	wire n1404;
	wire n1405;
	wire n1406;
	wire n1407;
	wire n1408;
	wire n1409;
	wire n1410;
	wire n1411;
	wire n1412;
	wire n1413;
	wire n1414;
	wire n1415;
	wire n1416;
	wire n1417;
	wire n1418;
	wire n1419;
	wire n1420;
	wire n1421;
	wire n1422;
	wire n1423;
	wire n1424;
	wire n1425;
	wire n1426;
	wire n1427;
	wire n1428;
	wire n1429;
	wire n1430;
	wire n1431;
	wire n1432;
	wire n1433;
	wire n1434;
	wire n1435;
	wire n1436;
	wire n1437;
	wire n1438;
	wire n1439;
	wire n1440;
	wire n1441;
	wire n1442;
	wire n1443;
	wire n1444;
	wire n1445;
	wire n1446;
	wire n1447;
	wire n1448;
	wire n1449;
	wire n1450;
	wire n1451;
	wire n1452;
	wire n1454;
	wire n1455;
	wire n1456;
	wire n1457;
	wire n1458;
	wire n1459;
	wire n1460;
	wire n1461;
	wire n1462;
	wire n1463;
	wire n1464;
	wire n1465;
	wire n1466;
	wire n1467;
	wire n1468;
	wire n1469;
	wire n1470;
	wire n1471;
	wire n1472;
	wire n1473;
	wire n1474;
	wire n1475;
	wire n1476;
	wire n1477;
	wire n1478;
	wire n1479;
	wire n1480;
	wire n1481;
	wire n1482;
	wire n1483;
	wire n1484;
	wire n1485;
	wire n1486;
	wire n1487;
	wire n1488;
	wire n1489;
	wire n1490;
	wire n1491;
	wire n1492;
	wire n1493;
	wire n1494;
	wire n1495;
	wire n1496;
	wire n1497;
	wire n1498;
	wire n1499;
	wire n1500;
	wire n1501;
	wire n1502;
	wire n1503;
	wire n1504;
	wire n1505;
	wire n1506;
	wire n1507;
	wire n1508;
	wire n1509;
	wire n1510;
	wire n1511;
	wire n1512;
	wire n1513;
	wire n1514;
	wire n1515;
	wire n1516;
	wire n1517;
	wire n1518;
	wire n1519;
	wire n1520;
	wire n1521;
	wire n1522;
	wire n1523;
	wire n1524;
	wire n1525;
	wire n1526;
	wire n1527;
	wire n1528;
	wire n1529;
	wire n1530;
	wire n1531;
	wire n1532;
	wire n1533;
	wire n1534;
	wire n1535;
	wire n1536;
	wire n1537;
	wire n1538;
	wire n1539;
	wire n1540;
	wire n1541;
	wire n1542;
	wire n1543;
	wire n1544;
	wire n1545;
	wire n1546;
	wire n1547;
	wire n1548;
	wire n1549;
	wire n1550;
	wire n1551;
	wire n1552;
	wire n1553;
	wire n1554;
	wire n1555;
	wire n1556;
	wire n1557;
	wire n1558;
	wire n1559;
	wire n1560;
	wire n1561;
	wire n1562;
	wire n1563;
	wire n1564;
	wire n1565;
	wire n1566;
	wire n1567;
	wire n1568;
	wire n1569;
	wire n1570;
	wire n1571;
	wire n1572;
	wire n1573;
	wire n1574;
	wire n1575;
	wire n1576;
	wire n1577;
	wire n1578;
	wire n1579;
	wire n1580;
	wire n1581;
	wire n1582;
	wire n1583;
	wire n1584;
	wire n1585;
	wire n1586;
	wire n1587;
	wire n1588;
	wire n1589;
	wire n1590;
	wire n1591;
	wire n1592;
	wire n1593;
	wire n1594;
	wire n1595;
	wire n1596;
	wire n1597;
	wire n1599;
	wire n1600;
	wire n1601;
	wire n1602;
	wire n1603;
	wire n1604;
	wire n1605;
	wire n1606;
	wire n1607;
	wire n1608;
	wire n1609;
	wire n1610;
	wire n1611;
	wire n1612;
	wire n1613;
	wire n1614;
	wire n1615;
	wire n1617;
	wire n1618;
	wire n1619;
	wire n1620;
	wire n1621;
	wire n1622;
	wire n1624;
	wire n1625;
	wire n1626;
	wire n1627;
	wire n1628;
	wire n1629;
	wire n1630;
	wire n1631;
	wire n1632;
	wire n1633;
	wire n1634;
	wire n1635;
	wire n1636;
	wire n1637;
	wire n1638;
	wire n1639;
	wire n1641;
	wire n1642;
	wire n1643;
	wire n1644;
	wire n1645;
	wire n1646;
	wire n1647;
	wire n1648;
	wire n1649;
	wire n1650;
	wire n1651;
	wire [2:0] w_G1_0;
	wire [2:0] w_G1_1;
	wire [1:0] w_G1_2;
	wire [2:0] w_G4_0;
	wire [1:0] w_G4_1;
	wire [1:0] w_G11_0;
	wire [1:0] w_G14_0;
	wire [1:0] w_G17_0;
	wire [1:0] w_G20_0;
	wire [1:0] w_G37_0;
	wire [1:0] w_G40_0;
	wire [1:0] w_G43_0;
	wire [1:0] w_G46_0;
	wire [1:0] w_G49_0;
	wire [1:0] w_G54_0;
	wire [1:0] w_G61_0;
	wire [1:0] w_G64_0;
	wire [1:0] w_G67_0;
	wire [1:0] w_G70_0;
	wire [1:0] w_G73_0;
	wire [1:0] w_G76_0;
	wire [1:0] w_G91_0;
	wire [1:0] w_G100_0;
	wire [1:0] w_G103_0;
	wire [1:0] w_G106_0;
	wire [1:0] w_G109_0;
	wire [1:0] w_G123_0;
	wire [1:0] w_G132_0;
	wire [2:0] w_G137_0;
	wire [2:0] w_G137_1;
	wire [2:0] w_G137_2;
	wire [2:0] w_G137_3;
	wire [2:0] w_G137_4;
	wire [2:0] w_G137_5;
	wire [2:0] w_G137_6;
	wire [2:0] w_G137_7;
	wire [2:0] w_G137_8;
	wire [1:0] w_G137_9;
	wire [2:0] w_G141_0;
	wire [2:0] w_G141_1;
	wire [2:0] w_G141_2;
	wire [1:0] w_G146_0;
	wire [1:0] w_G149_0;
	wire [1:0] w_G152_0;
	wire [1:0] w_G155_0;
	wire [1:0] w_G158_0;
	wire [1:0] w_G161_0;
	wire [1:0] w_G164_0;
	wire [1:0] w_G167_0;
	wire [1:0] w_G170_0;
	wire [1:0] w_G173_0;
	wire [1:0] w_G182_0;
	wire [1:0] w_G185_0;
	wire [1:0] w_G188_0;
	wire [1:0] w_G191_0;
	wire [1:0] w_G194_0;
	wire [1:0] w_G197_0;
	wire [1:0] w_G200_0;
	wire [1:0] w_G203_0;
	wire [2:0] w_G206_0;
	wire [2:0] w_G210_0;
	wire [2:0] w_G210_1;
	wire [2:0] w_G210_2;
	wire [2:0] w_G218_0;
	wire [2:0] w_G218_1;
	wire [2:0] w_G218_2;
	wire [2:0] w_G226_0;
	wire [2:0] w_G226_1;
	wire [2:0] w_G226_2;
	wire [2:0] w_G234_0;
	wire [2:0] w_G234_1;
	wire [1:0] w_G234_2;
	wire [2:0] w_G242_0;
	wire [2:0] w_G242_1;
	wire [1:0] w_G245_0;
	wire [2:0] w_G248_0;
	wire [2:0] w_G248_1;
	wire [2:0] w_G248_2;
	wire [2:0] w_G248_3;
	wire [2:0] w_G248_4;
	wire [1:0] w_G248_5;
	wire [2:0] w_G251_0;
	wire [2:0] w_G251_1;
	wire [2:0] w_G251_2;
	wire [2:0] w_G251_3;
	wire [2:0] w_G251_4;
	wire [2:0] w_G254_0;
	wire [2:0] w_G254_1;
	wire [2:0] w_G257_0;
	wire [2:0] w_G257_1;
	wire [2:0] w_G257_2;
	wire [2:0] w_G265_0;
	wire [2:0] w_G265_1;
	wire [1:0] w_G265_2;
	wire [2:0] w_G273_0;
	wire [2:0] w_G273_1;
	wire [2:0] w_G273_2;
	wire [1:0] w_G280_0;
	wire [2:0] w_G281_0;
	wire [2:0] w_G281_1;
	wire [1:0] w_G281_2;
	wire [1:0] w_G289_0;
	wire [2:0] w_G293_0;
	wire [2:0] w_G299_0;
	wire [2:0] w_G302_0;
	wire [2:0] w_G308_0;
	wire [2:0] w_G308_1;
	wire [2:0] w_G316_0;
	wire [2:0] w_G316_1;
	wire [2:0] w_G324_0;
	wire [2:0] w_G324_1;
	wire [1:0] w_G331_0;
	wire [2:0] w_G332_0;
	wire [2:0] w_G332_1;
	wire [2:0] w_G332_2;
	wire [2:0] w_G332_3;
	wire [2:0] w_G332_4;
	wire [2:0] w_G335_0;
	wire [2:0] w_G335_1;
	wire [2:0] w_G335_2;
	wire [2:0] w_G335_3;
	wire [1:0] w_G335_4;
	wire [2:0] w_G341_0;
	wire [2:0] w_G341_1;
	wire [2:0] w_G341_2;
	wire [1:0] w_G348_0;
	wire [2:0] w_G351_0;
	wire [2:0] w_G351_1;
	wire [2:0] w_G351_2;
	wire [1:0] w_G358_0;
	wire [2:0] w_G361_0;
	wire [1:0] w_G369_0;
	wire [2:0] w_G374_0;
	wire [2:0] w_G389_0;
	wire [2:0] w_G400_0;
	wire [1:0] w_G400_1;
	wire [2:0] w_G411_0;
	wire [2:0] w_G422_0;
	wire [2:0] w_G422_1;
	wire [1:0] w_G422_2;
	wire [2:0] w_G435_0;
	wire [2:0] w_G435_1;
	wire [2:0] w_G446_0;
	wire [2:0] w_G446_1;
	wire [2:0] w_G457_0;
	wire [2:0] w_G457_1;
	wire [1:0] w_G457_2;
	wire [2:0] w_G468_0;
	wire [2:0] w_G468_1;
	wire [2:0] w_G479_0;
	wire [1:0] w_G479_1;
	wire [2:0] w_G490_0;
	wire [2:0] w_G490_1;
	wire [2:0] w_G503_0;
	wire [2:0] w_G503_1;
	wire [2:0] w_G514_0;
	wire [1:0] w_G514_1;
	wire [2:0] w_G523_0;
	wire [1:0] w_G523_1;
	wire [2:0] w_G534_0;
	wire [2:0] w_G534_1;
	wire [2:0] w_G545_0;
	wire [2:0] w_G549_0;
	wire [1:0] w_G552_0;
	wire [1:0] w_G559_0;
	wire [1:0] w_G562_0;
	wire [2:0] w_G1497_0;
	wire [2:0] w_G1689_0;
	wire [2:0] w_G1690_0;
	wire [2:0] w_G1691_0;
	wire [2:0] w_G1694_0;
	wire [2:0] w_G2174_0;
	wire [2:0] w_G2358_0;
	wire [2:0] w_G2358_1;
	wire [2:0] w_G2358_2;
	wire [1:0] w_G3173_0;
	wire [2:0] w_G3546_0;
	wire [2:0] w_G3546_1;
	wire [2:0] w_G3546_2;
	wire [2:0] w_G3546_3;
	wire [2:0] w_G3546_4;
	wire [1:0] w_G3546_5;
	wire [2:0] w_G3548_0;
	wire [2:0] w_G3548_1;
	wire [2:0] w_G3548_2;
	wire [2:0] w_G3548_3;
	wire [2:0] w_G3548_4;
	wire [1:0] w_G3552_0;
	wire [1:0] w_G3717_0;
	wire [2:0] w_G3724_0;
	wire [2:0] w_G4087_0;
	wire [2:0] w_G4088_0;
	wire [2:0] w_G4089_0;
	wire [2:0] w_G4090_0;
	wire [2:0] w_G4091_0;
	wire [2:0] w_G4091_1;
	wire [2:0] w_G4091_2;
	wire [2:0] w_G4092_0;
	wire [2:0] w_G4092_1;
	wire w_G599_0;
	wire G599_fa_;
	wire w_G600_0;
	wire G600_fa_;
	wire w_G601_0;
	wire G601_fa_;
	wire w_G611_0;
	wire G611_fa_;
	wire w_G612_0;
	wire G612_fa_;
	wire [2:0] w_G809_0;
	wire [2:0] w_G809_1;
	wire [2:0] w_G809_2;
	wire [1:0] w_G809_3;
	wire G809_fa_;
	wire w_G593_0;
	wire G593_fa_;
	wire w_G822_0;
	wire G822_fa_;
	wire w_G838_0;
	wire G838_fa_;
	wire w_G861_0;
	wire G861_fa_;
	wire w_G832_0;
	wire G832_fa_;
	wire w_G834_0;
	wire G834_fa_;
	wire w_G836_0;
	wire G836_fa_;
	wire w_G871_0;
	wire G871_fa_;
	wire w_G873_0;
	wire G873_fa_;
	wire w_G875_0;
	wire G875_fa_;
	wire w_G877_0;
	wire G877_fa_;
	wire w_G1000_0;
	wire G1000_fa_;
	wire w_G826_0;
	wire G826_fa_;
	wire w_G828_0;
	wire G828_fa_;
	wire w_G830_0;
	wire G830_fa_;
	wire w_G867_0;
	wire G867_fa_;
	wire w_G869_0;
	wire G869_fa_;
	wire [1:0] w_n316_0;
	wire [1:0] w_n318_0;
	wire [2:0] w_n326_0;
	wire [2:0] w_n326_1;
	wire [1:0] w_n326_2;
	wire [1:0] w_n333_0;
	wire [1:0] w_n336_0;
	wire [1:0] w_n360_0;
	wire [1:0] w_n362_0;
	wire [2:0] w_n366_0;
	wire [2:0] w_n366_1;
	wire [2:0] w_n366_2;
	wire [2:0] w_n366_3;
	wire [2:0] w_n366_4;
	wire [2:0] w_n368_0;
	wire [2:0] w_n368_1;
	wire [2:0] w_n368_2;
	wire [2:0] w_n368_3;
	wire [2:0] w_n368_4;
	wire [1:0] w_n368_5;
	wire [2:0] w_n372_0;
	wire [1:0] w_n373_0;
	wire [2:0] w_n383_0;
	wire [2:0] w_n385_0;
	wire [2:0] w_n385_1;
	wire [2:0] w_n386_0;
	wire [2:0] w_n386_1;
	wire [2:0] w_n386_2;
	wire [2:0] w_n386_3;
	wire [2:0] w_n386_4;
	wire [2:0] w_n388_0;
	wire [2:0] w_n388_1;
	wire [2:0] w_n389_0;
	wire [2:0] w_n389_1;
	wire [2:0] w_n389_2;
	wire [2:0] w_n389_3;
	wire [2:0] w_n389_4;
	wire [1:0] w_n397_0;
	wire [2:0] w_n398_0;
	wire [2:0] w_n401_0;
	wire [2:0] w_n402_0;
	wire [2:0] w_n402_1;
	wire [1:0] w_n402_2;
	wire [1:0] w_n403_0;
	wire [2:0] w_n405_0;
	wire [2:0] w_n405_1;
	wire [1:0] w_n405_2;
	wire [1:0] w_n407_0;
	wire [1:0] w_n408_0;
	wire [2:0] w_n410_0;
	wire [1:0] w_n410_1;
	wire [1:0] w_n414_0;
	wire [1:0] w_n416_0;
	wire [2:0] w_n419_0;
	wire [2:0] w_n424_0;
	wire [2:0] w_n424_1;
	wire [1:0] w_n424_2;
	wire [1:0] w_n426_0;
	wire [1:0] w_n434_0;
	wire [2:0] w_n435_0;
	wire [2:0] w_n435_1;
	wire [2:0] w_n437_0;
	wire [2:0] w_n437_1;
	wire [1:0] w_n445_0;
	wire [2:0] w_n449_0;
	wire [2:0] w_n449_1;
	wire [2:0] w_n451_0;
	wire [1:0] w_n451_1;
	wire [1:0] w_n459_0;
	wire [2:0] w_n460_0;
	wire [2:0] w_n460_1;
	wire [2:0] w_n462_0;
	wire [1:0] w_n470_0;
	wire [2:0] w_n471_0;
	wire [1:0] w_n471_1;
	wire [2:0] w_n473_0;
	wire [2:0] w_n473_1;
	wire [1:0] w_n481_0;
	wire [2:0] w_n484_0;
	wire [1:0] w_n484_1;
	wire [2:0] w_n486_0;
	wire [1:0] w_n486_1;
	wire [1:0] w_n494_0;
	wire [2:0] w_n495_0;
	wire [2:0] w_n495_1;
	wire [2:0] w_n497_0;
	wire [1:0] w_n497_1;
	wire [1:0] w_n505_0;
	wire [2:0] w_n507_0;
	wire [1:0] w_n507_1;
	wire [1:0] w_n509_0;
	wire [1:0] w_n517_0;
	wire [2:0] w_n518_0;
	wire [1:0] w_n518_1;
	wire [2:0] w_n528_0;
	wire [2:0] w_n530_0;
	wire [1:0] w_n530_1;
	wire [1:0] w_n532_0;
	wire [1:0] w_n540_0;
	wire [2:0] w_n541_0;
	wire [1:0] w_n541_1;
	wire [1:0] w_n543_0;
	wire [1:0] w_n551_0;
	wire [2:0] w_n556_0;
	wire [2:0] w_n556_1;
	wire [2:0] w_n556_2;
	wire [2:0] w_n556_3;
	wire [2:0] w_n556_4;
	wire [1:0] w_n556_5;
	wire [2:0] w_n560_0;
	wire [1:0] w_n560_1;
	wire [2:0] w_n561_0;
	wire [1:0] w_n562_0;
	wire [2:0] w_n566_0;
	wire [2:0] w_n567_0;
	wire [1:0] w_n567_1;
	wire [1:0] w_n569_0;
	wire [1:0] w_n570_0;
	wire [2:0] w_n571_0;
	wire [1:0] w_n571_1;
	wire [2:0] w_n572_0;
	wire [2:0] w_n574_0;
	wire [2:0] w_n577_0;
	wire [2:0] w_n578_0;
	wire [2:0] w_n582_0;
	wire [1:0] w_n582_1;
	wire [2:0] w_n583_0;
	wire [1:0] w_n583_1;
	wire [1:0] w_n585_0;
	wire [2:0] w_n587_0;
	wire [1:0] w_n587_1;
	wire [2:0] w_n590_0;
	wire [1:0] w_n590_1;
	wire [1:0] w_n591_0;
	wire [2:0] w_n595_0;
	wire [1:0] w_n595_1;
	wire [2:0] w_n596_0;
	wire [2:0] w_n600_0;
	wire [1:0] w_n600_1;
	wire [1:0] w_n601_0;
	wire [2:0] w_n604_0;
	wire [2:0] w_n605_0;
	wire [2:0] w_n605_1;
	wire [2:0] w_n605_2;
	wire [2:0] w_n607_0;
	wire [2:0] w_n609_0;
	wire [2:0] w_n609_1;
	wire [2:0] w_n609_2;
	wire [2:0] w_n609_3;
	wire [2:0] w_n609_4;
	wire [2:0] w_n609_5;
	wire [2:0] w_n613_0;
	wire [2:0] w_n614_0;
	wire [2:0] w_n614_1;
	wire [1:0] w_n614_2;
	wire [2:0] w_n617_0;
	wire [1:0] w_n617_1;
	wire [2:0] w_n618_0;
	wire [1:0] w_n618_1;
	wire [2:0] w_n621_0;
	wire [2:0] w_n621_1;
	wire [1:0] w_n621_2;
	wire [2:0] w_n622_0;
	wire [1:0] w_n622_1;
	wire [1:0] w_n623_0;
	wire [2:0] w_n624_0;
	wire [2:0] w_n624_1;
	wire [2:0] w_n625_0;
	wire [2:0] w_n628_0;
	wire [2:0] w_n629_0;
	wire [1:0] w_n631_0;
	wire [2:0] w_n633_0;
	wire [1:0] w_n633_1;
	wire [2:0] w_n636_0;
	wire [1:0] w_n636_1;
	wire [2:0] w_n640_0;
	wire [2:0] w_n640_1;
	wire [1:0] w_n641_0;
	wire [1:0] w_n642_0;
	wire [2:0] w_n645_0;
	wire [2:0] w_n646_0;
	wire [2:0] w_n649_0;
	wire [1:0] w_n649_1;
	wire [1:0] w_n650_0;
	wire [2:0] w_n651_0;
	wire [1:0] w_n651_1;
	wire [1:0] w_n652_0;
	wire [1:0] w_n661_0;
	wire [1:0] w_n671_0;
	wire [1:0] w_n677_0;
	wire [1:0] w_n678_0;
	wire [1:0] w_n679_0;
	wire [1:0] w_n680_0;
	wire [2:0] w_n681_0;
	wire [2:0] w_n681_1;
	wire [1:0] w_n681_2;
	wire [1:0] w_n682_0;
	wire [2:0] w_n687_0;
	wire [1:0] w_n689_0;
	wire [2:0] w_n691_0;
	wire [2:0] w_n693_0;
	wire [2:0] w_n696_0;
	wire [1:0] w_n697_0;
	wire [1:0] w_n700_0;
	wire [1:0] w_n702_0;
	wire [2:0] w_n703_0;
	wire [1:0] w_n705_0;
	wire [1:0] w_n706_0;
	wire [2:0] w_n707_0;
	wire [1:0] w_n709_0;
	wire [1:0] w_n716_0;
	wire [2:0] w_n717_0;
	wire [1:0] w_n720_0;
	wire [2:0] w_n721_0;
	wire [1:0] w_n723_0;
	wire [1:0] w_n726_0;
	wire [2:0] w_n727_0;
	wire [2:0] w_n729_0;
	wire [1:0] w_n729_1;
	wire [2:0] w_n732_0;
	wire [1:0] w_n733_0;
	wire [1:0] w_n735_0;
	wire [1:0] w_n736_0;
	wire [2:0] w_n739_0;
	wire [1:0] w_n739_1;
	wire [1:0] w_n740_0;
	wire [1:0] w_n741_0;
	wire [1:0] w_n742_0;
	wire [2:0] w_n744_0;
	wire [2:0] w_n744_1;
	wire [2:0] w_n746_0;
	wire [2:0] w_n746_1;
	wire [2:0] w_n747_0;
	wire [2:0] w_n747_1;
	wire [2:0] w_n747_2;
	wire [2:0] w_n747_3;
	wire [2:0] w_n748_0;
	wire [2:0] w_n748_1;
	wire [2:0] w_n748_2;
	wire [2:0] w_n748_3;
	wire [1:0] w_n748_4;
	wire [2:0] w_n750_0;
	wire [1:0] w_n750_1;
	wire [2:0] w_n751_0;
	wire [2:0] w_n751_1;
	wire [1:0] w_n751_2;
	wire [2:0] w_n753_0;
	wire [2:0] w_n753_1;
	wire [2:0] w_n753_2;
	wire [2:0] w_n753_3;
	wire [2:0] w_n753_4;
	wire [2:0] w_n753_5;
	wire [2:0] w_n753_6;
	wire [2:0] w_n753_7;
	wire [1:0] w_n753_8;
	wire [1:0] w_n759_0;
	wire [1:0] w_n760_0;
	wire [1:0] w_n761_0;
	wire [2:0] w_n765_0;
	wire [2:0] w_n765_1;
	wire [2:0] w_n765_2;
	wire [2:0] w_n765_3;
	wire [2:0] w_n765_4;
	wire [2:0] w_n765_5;
	wire [1:0] w_n771_0;
	wire [1:0] w_n779_0;
	wire [2:0] w_n781_0;
	wire [2:0] w_n783_0;
	wire [1:0] w_n783_1;
	wire [1:0] w_n786_0;
	wire [1:0] w_n787_0;
	wire [2:0] w_n789_0;
	wire [2:0] w_n791_0;
	wire [1:0] w_n791_1;
	wire [1:0] w_n792_0;
	wire [2:0] w_n793_0;
	wire [2:0] w_n793_1;
	wire [2:0] w_n793_2;
	wire [2:0] w_n793_3;
	wire [1:0] w_n793_4;
	wire [2:0] w_n795_0;
	wire [1:0] w_n795_1;
	wire [1:0] w_n796_0;
	wire [2:0] w_n797_0;
	wire [2:0] w_n797_1;
	wire [2:0] w_n797_2;
	wire [2:0] w_n797_3;
	wire [1:0] w_n797_4;
	wire [2:0] w_n799_0;
	wire [2:0] w_n799_1;
	wire [2:0] w_n799_2;
	wire [2:0] w_n799_3;
	wire [1:0] w_n799_4;
	wire [2:0] w_n801_0;
	wire [2:0] w_n801_1;
	wire [2:0] w_n801_2;
	wire [2:0] w_n801_3;
	wire [1:0] w_n801_4;
	wire [2:0] w_n806_0;
	wire [1:0] w_n809_0;
	wire [1:0] w_n819_0;
	wire [1:0] w_n821_0;
	wire [2:0] w_n828_0;
	wire [1:0] w_n829_0;
	wire [1:0] w_n832_0;
	wire [1:0] w_n839_0;
	wire [2:0] w_n840_0;
	wire [2:0] w_n840_1;
	wire [2:0] w_n840_2;
	wire [2:0] w_n840_3;
	wire [1:0] w_n840_4;
	wire [1:0] w_n842_0;
	wire [2:0] w_n843_0;
	wire [2:0] w_n843_1;
	wire [2:0] w_n843_2;
	wire [2:0] w_n843_3;
	wire [1:0] w_n843_4;
	wire [2:0] w_n845_0;
	wire [2:0] w_n845_1;
	wire [2:0] w_n845_2;
	wire [2:0] w_n845_3;
	wire [1:0] w_n845_4;
	wire [2:0] w_n847_0;
	wire [2:0] w_n847_1;
	wire [2:0] w_n847_2;
	wire [2:0] w_n847_3;
	wire [1:0] w_n847_4;
	wire [1:0] w_n853_0;
	wire [1:0] w_n855_0;
	wire [1:0] w_n856_0;
	wire [1:0] w_n857_0;
	wire [1:0] w_n859_0;
	wire [1:0] w_n862_0;
	wire [1:0] w_n869_0;
	wire [1:0] w_n877_0;
	wire [1:0] w_n879_0;
	wire [1:0] w_n881_0;
	wire [1:0] w_n892_0;
	wire [1:0] w_n914_0;
	wire [1:0] w_n928_0;
	wire [2:0] w_n930_0;
	wire [1:0] w_n932_0;
	wire [2:0] w_n936_0;
	wire [1:0] w_n938_0;
	wire [1:0] w_n941_0;
	wire [1:0] w_n943_0;
	wire [1:0] w_n944_0;
	wire [1:0] w_n946_0;
	wire [2:0] w_n948_0;
	wire [1:0] w_n953_0;
	wire [1:0] w_n954_0;
	wire [1:0] w_n968_0;
	wire [1:0] w_n971_0;
	wire [1:0] w_n972_0;
	wire [1:0] w_n973_0;
	wire [1:0] w_n984_0;
	wire [2:0] w_n985_0;
	wire [2:0] w_n985_1;
	wire [2:0] w_n985_2;
	wire [2:0] w_n985_3;
	wire [1:0] w_n985_4;
	wire [1:0] w_n987_0;
	wire [2:0] w_n988_0;
	wire [2:0] w_n988_1;
	wire [2:0] w_n988_2;
	wire [2:0] w_n988_3;
	wire [1:0] w_n988_4;
	wire [2:0] w_n990_0;
	wire [2:0] w_n990_1;
	wire [2:0] w_n990_2;
	wire [2:0] w_n990_3;
	wire [1:0] w_n990_4;
	wire [2:0] w_n992_0;
	wire [2:0] w_n992_1;
	wire [2:0] w_n992_2;
	wire [2:0] w_n992_3;
	wire [1:0] w_n992_4;
	wire [1:0] w_n998_0;
	wire [2:0] w_n999_0;
	wire [2:0] w_n999_1;
	wire [2:0] w_n999_2;
	wire [2:0] w_n999_3;
	wire [1:0] w_n999_4;
	wire [1:0] w_n1001_0;
	wire [2:0] w_n1002_0;
	wire [2:0] w_n1002_1;
	wire [2:0] w_n1002_2;
	wire [2:0] w_n1002_3;
	wire [1:0] w_n1002_4;
	wire [2:0] w_n1004_0;
	wire [2:0] w_n1004_1;
	wire [2:0] w_n1004_2;
	wire [2:0] w_n1004_3;
	wire [1:0] w_n1004_4;
	wire [2:0] w_n1006_0;
	wire [2:0] w_n1006_1;
	wire [2:0] w_n1006_2;
	wire [2:0] w_n1006_3;
	wire [1:0] w_n1006_4;
	wire [2:0] w_n1012_0;
	wire [1:0] w_n1012_1;
	wire [2:0] w_n1014_0;
	wire [1:0] w_n1014_1;
	wire [2:0] w_n1021_0;
	wire [1:0] w_n1021_1;
	wire [2:0] w_n1023_0;
	wire [1:0] w_n1023_1;
	wire [2:0] w_n1030_0;
	wire [1:0] w_n1030_1;
	wire [2:0] w_n1032_0;
	wire [1:0] w_n1032_1;
	wire [2:0] w_n1039_0;
	wire [1:0] w_n1039_1;
	wire [2:0] w_n1041_0;
	wire [1:0] w_n1041_1;
	wire [1:0] w_n1142_0;
	wire [1:0] w_n1151_0;
	wire [2:0] w_n1163_0;
	wire [2:0] w_n1163_1;
	wire [2:0] w_n1197_0;
	wire [2:0] w_n1197_1;
	wire [2:0] w_n1205_0;
	wire [2:0] w_n1205_1;
	wire [2:0] w_n1235_0;
	wire [1:0] w_n1235_1;
	wire [2:0] w_n1242_0;
	wire [1:0] w_n1242_1;
	wire [2:0] w_n1244_0;
	wire [1:0] w_n1244_1;
	wire [2:0] w_n1251_0;
	wire [1:0] w_n1251_1;
	wire [2:0] w_n1253_0;
	wire [1:0] w_n1253_1;
	wire [1:0] w_n1358_0;
	wire [1:0] w_n1383_0;
	wire [1:0] w_n1391_0;
	wire [1:0] w_n1394_0;
	wire [1:0] w_n1398_0;
	wire [1:0] w_n1399_0;
	wire [1:0] w_n1409_0;
	wire [1:0] w_n1410_0;
	wire [1:0] w_n1411_0;
	wire [1:0] w_n1421_0;
	wire [1:0] w_n1425_0;
	wire [1:0] w_n1434_0;
	wire [1:0] w_n1438_0;
	wire [1:0] w_n1445_0;
	wire [1:0] w_n1446_0;
	wire [1:0] w_n1447_0;
	wire [1:0] w_n1452_0;
	wire [1:0] w_n1494_0;
	wire [1:0] w_n1533_0;
	wire [1:0] w_n1543_0;
	wire [1:0] w_n1545_0;
	wire [1:0] w_n1553_0;
	wire [1:0] w_n1555_0;
	wire [1:0] w_n1560_0;
	wire [1:0] w_n1568_0;
	wire [1:0] w_n1591_0;
	wire [1:0] w_n1597_0;
	wire [2:0] w_n1601_0;
	wire [1:0] w_n1602_0;
	wire [1:0] w_n1609_0;
	wire [1:0] w_n1610_0;
	wire [1:0] w_n1624_0;
	wire [1:0] w_n1629_0;
	wire [1:0] w_n1631_0;
	wire [1:0] w_n1634_0;
	wire w_dff_B_WGdD0rVS3_1;
	wire w_dff_B_f0LYeUl25_0;
	wire w_dff_A_BFIIhYPO2_0;
	wire w_dff_B_VJcHhuhL0_0;
	wire w_dff_A_YBhqqeWI3_2;
	wire w_dff_B_BlANR4eP3_1;
	wire w_dff_B_JCFpbHak3_0;
	wire w_dff_B_q4l2q9D84_1;
	wire w_dff_A_p8cfZKe11_0;
	wire w_dff_A_mDj9H6QG7_0;
	wire w_dff_A_I6kXeqgr8_1;
	wire w_dff_A_AkhK1X9s5_1;
	wire w_dff_B_8ew7en6g4_0;
	wire w_dff_B_WJPsYA0z2_1;
	wire w_dff_B_eOyn8kPV5_0;
	wire w_dff_B_nZ4R98sA0_1;
	wire w_dff_A_UZf91e0e1_0;
	wire w_dff_A_kvAw0xGb1_1;
	wire w_dff_A_cmdfPIZp2_1;
	wire w_dff_A_3bTWSZ4q7_1;
	wire w_dff_A_Oq6xX8ZF7_2;
	wire w_dff_A_gGbZoHhG3_2;
	wire w_dff_B_eCm3PMS85_1;
	wire w_dff_B_e4aO8TUb8_1;
	wire w_dff_B_QKD54ivv8_1;
	wire w_dff_B_8ntSLRtx1_0;
	wire w_dff_B_905voHzG3_0;
	wire w_dff_B_gU6HXDMJ4_1;
	wire w_dff_B_yw7XDC1h4_1;
	wire w_dff_B_DSVEcvlF0_2;
	wire w_dff_B_yBanOqkZ1_2;
	wire w_dff_B_yCe85Kji7_2;
	wire w_dff_B_tml5FdyV9_1;
	wire w_dff_B_F8cqQGOc6_1;
	wire w_dff_A_Y58LOX3i0_1;
	wire w_dff_B_VSrcI6kO7_0;
	wire w_dff_B_W1C3vtJh6_0;
	wire w_dff_B_GqvEaJZe2_2;
	wire w_dff_A_n5t01ZQF1_0;
	wire w_dff_B_PhSDkhuw2_0;
	wire w_dff_B_w4igoQQ31_0;
	wire w_dff_B_Vzbf7DTq3_0;
	wire w_dff_B_8H1wQF9T7_0;
	wire w_dff_B_yjg5KfqY6_0;
	wire w_dff_B_TeOv1NbB9_0;
	wire w_dff_B_F722iPpp8_0;
	wire w_dff_B_2cN4VASt5_0;
	wire w_dff_B_Y4WLp8Fb2_0;
	wire w_dff_B_9BhNk8EB2_0;
	wire w_dff_B_SR0lf29E3_0;
	wire w_dff_B_z1phqwup6_0;
	wire w_dff_B_rySoRXaP3_0;
	wire w_dff_B_Mw5zA2y87_0;
	wire w_dff_B_OBQcQGTx9_2;
	wire w_dff_B_aHqIICak1_2;
	wire w_dff_B_BiD5EdXq3_2;
	wire w_dff_B_FwBDmWms0_1;
	wire w_dff_B_9Xrlp8t79_1;
	wire w_dff_B_FLk7yXTK9_1;
	wire w_dff_B_I6hnxsZq9_1;
	wire w_dff_B_dSMLp7Iu5_1;
	wire w_dff_B_aGPEn6zR7_1;
	wire w_dff_B_DxRhincp4_1;
	wire w_dff_B_5hBGFDgg4_1;
	wire w_dff_B_lMCtFf5v0_1;
	wire w_dff_B_Hs2jrfC70_1;
	wire w_dff_B_Cc4JLWJc2_1;
	wire w_dff_B_pastvOPG7_0;
	wire w_dff_B_PlStXqfk4_0;
	wire w_dff_B_TxdIXZpt4_0;
	wire w_dff_B_2u3sRBDv6_0;
	wire w_dff_B_dZxZuFOa6_0;
	wire w_dff_B_za3o7y3d3_0;
	wire w_dff_B_8Q2p3NVF7_0;
	wire w_dff_B_tOz9RWR58_0;
	wire w_dff_B_4xQBvl2r0_0;
	wire w_dff_B_lXhl7vWC1_0;
	wire w_dff_B_KpZXeaHc9_0;
	wire w_dff_B_qC6oRdRK1_0;
	wire w_dff_B_e0WHgypv3_0;
	wire w_dff_B_sZWv7KcA3_0;
	wire w_dff_B_IB2lwABJ2_0;
	wire w_dff_B_Slzp9vaC8_0;
	wire w_dff_B_8Yt5X2SC2_2;
	wire w_dff_B_f8KbmwrY8_2;
	wire w_dff_B_y7pSZth39_2;
	wire w_dff_B_eSJT5Mt21_1;
	wire w_dff_B_Vtl8R2nH1_1;
	wire w_dff_B_26hfeWVD4_1;
	wire w_dff_B_2OZpruAF3_0;
	wire w_dff_B_nYzCmORx9_1;
	wire w_dff_B_gyx2IgSc9_1;
	wire w_dff_B_gMgEU3kz8_1;
	wire w_dff_B_1pMomV046_0;
	wire w_dff_B_Mw9bT7h82_0;
	wire w_dff_B_WWtYwvnd6_0;
	wire w_dff_B_jLsh2peL3_0;
	wire w_dff_B_TBw81uok5_0;
	wire w_dff_B_JVjiMPN85_0;
	wire w_dff_B_X97uTZ773_0;
	wire w_dff_B_goH244bY6_0;
	wire w_dff_B_G8RuqwgS0_0;
	wire w_dff_B_Aaqk6xgn3_0;
	wire w_dff_B_hjjrRSHq0_0;
	wire w_dff_B_QwYmrZtN6_0;
	wire w_dff_B_yzh2W3DX2_0;
	wire w_dff_A_VAD0TqVh9_0;
	wire w_dff_A_4h6dq7J39_0;
	wire w_dff_A_Izq4Ek8W1_0;
	wire w_dff_A_rFYTqiN56_0;
	wire w_dff_A_Q5vjTzVR8_0;
	wire w_dff_A_Vk6xNNQ11_0;
	wire w_dff_A_xdg5shdo1_0;
	wire w_dff_A_ZCK0Bsrp4_0;
	wire w_dff_B_Gx18M9zT8_0;
	wire w_dff_B_3yp9MbZK8_0;
	wire w_dff_B_pBpLQpd10_0;
	wire w_dff_B_SYCIhiJY9_0;
	wire w_dff_B_7I729Ujb7_0;
	wire w_dff_B_2uBfnEDK1_0;
	wire w_dff_B_5ouMzg7U1_0;
	wire w_dff_B_8cuKNfSZ2_0;
	wire w_dff_B_LnPLsUzR2_0;
	wire w_dff_B_0l4ExStx1_0;
	wire w_dff_B_EFOHvvMd4_0;
	wire w_dff_B_khimyeJF9_0;
	wire w_dff_B_AdtNkSCw9_0;
	wire w_dff_B_MaPgAzdj1_0;
	wire w_dff_B_CTXroHMd3_0;
	wire w_dff_B_J6wrzi0i8_0;
	wire w_dff_B_RYV23nIl2_0;
	wire w_dff_B_eZrPI4Qr5_0;
	wire w_dff_B_KIUWV3WE9_0;
	wire w_dff_B_5gEmHFrd6_0;
	wire w_dff_B_Lr4O21im4_0;
	wire w_dff_B_1C1cxjdS6_0;
	wire w_dff_B_oY8yNrqq5_0;
	wire w_dff_B_8heiXQ8D1_0;
	wire w_dff_B_twzCbOZs0_0;
	wire w_dff_B_2A9yH7yX5_0;
	wire w_dff_B_c8kVFgYn3_0;
	wire w_dff_B_iFytHTv26_0;
	wire w_dff_B_LQ9cAgVa6_0;
	wire w_dff_B_MjDqlfFb8_0;
	wire w_dff_B_5ETUfBtl6_0;
	wire w_dff_B_XCdzVBk76_0;
	wire w_dff_B_Yr3r80KN9_0;
	wire w_dff_A_wcEwDFX14_1;
	wire w_dff_A_okWsnYcW0_2;
	wire w_dff_B_xtW8R4l04_0;
	wire w_dff_B_Hqj2BGyl6_0;
	wire w_dff_B_jJSd5e4E3_0;
	wire w_dff_B_oef3wOMR0_0;
	wire w_dff_B_9JNPfFuv2_0;
	wire w_dff_B_vwqSx1125_0;
	wire w_dff_B_VVhxjbwL1_0;
	wire w_dff_B_ElcNvPpo7_0;
	wire w_dff_B_ng7hVfxZ8_0;
	wire w_dff_B_a3Ht3qBZ7_0;
	wire w_dff_B_cQsrr4c32_0;
	wire w_dff_B_pW89VdJt3_0;
	wire w_dff_B_xxhTC5x54_2;
	wire w_dff_B_W2UJTWXX5_2;
	wire w_dff_B_jwtZKyDM4_2;
	wire w_dff_A_3wxzoUkB3_0;
	wire w_dff_A_NwY7EWSI2_0;
	wire w_dff_A_jbpOdlvy3_0;
	wire w_dff_A_KRCB5eEO6_0;
	wire w_dff_A_E6neABW57_0;
	wire w_dff_A_ZEZKEdrn9_0;
	wire w_dff_A_U9CsHbJj0_0;
	wire w_dff_A_fGW91Ct89_0;
	wire w_dff_B_idkaQGLg2_0;
	wire w_dff_B_BgSD60qq6_0;
	wire w_dff_B_jHgNWtvc9_0;
	wire w_dff_B_wNxtMbtO6_0;
	wire w_dff_B_YnJ1Yh5H7_0;
	wire w_dff_B_F0gT7RyK7_0;
	wire w_dff_B_QXDjpZVM0_0;
	wire w_dff_B_kmRSgUaW3_0;
	wire w_dff_B_YQI6wa8Z8_0;
	wire w_dff_B_TNC4Qb987_0;
	wire w_dff_B_GaCqMgtu1_0;
	wire w_dff_B_8T3VWiob3_2;
	wire w_dff_B_xTwIwzGE1_2;
	wire w_dff_B_hl6lL76m7_2;
	wire w_dff_B_OTb1d4NB6_0;
	wire w_dff_B_02LvlSIN4_0;
	wire w_dff_B_2jnld2Lr1_0;
	wire w_dff_B_59nKBC3D3_0;
	wire w_dff_B_iy8RiUN58_0;
	wire w_dff_B_7NWbyQmR1_0;
	wire w_dff_B_yloQAErT0_0;
	wire w_dff_B_Daw1tBii1_0;
	wire w_dff_B_k9DmYLW29_0;
	wire w_dff_B_JurtH47K4_0;
	wire w_dff_B_9FV3cLIM8_0;
	wire w_dff_B_933tUGNJ1_2;
	wire w_dff_B_yoWYvQti6_2;
	wire w_dff_B_9UiXsHup0_2;
	wire w_dff_B_Rlcf1GDx5_0;
	wire w_dff_B_XDV9kWAm9_0;
	wire w_dff_B_qBWSZGAX7_0;
	wire w_dff_B_brjs7dzY8_0;
	wire w_dff_B_Wv0NtsIA4_0;
	wire w_dff_B_l5Uh0TeI7_0;
	wire w_dff_B_r48g0MKq6_0;
	wire w_dff_B_8aRDAa4P7_0;
	wire w_dff_B_nNKbKmfi0_0;
	wire w_dff_B_wBIa7dao0_0;
	wire w_dff_B_mvLIU5Ui7_0;
	wire w_dff_B_evZZUxAQ6_2;
	wire w_dff_B_Sr0Z6q3F9_2;
	wire w_dff_B_ebTHCX9D8_2;
	wire w_dff_A_9OgRyhsy3_1;
	wire w_dff_A_X0jYu4GN5_2;
	wire w_dff_B_De6HjeTr5_0;
	wire w_dff_B_1pC0sKdg5_0;
	wire w_dff_B_JFXFQfai5_0;
	wire w_dff_B_1IWmYF6w0_0;
	wire w_dff_B_7p7zo9qH2_0;
	wire w_dff_B_AfJ0b24G1_0;
	wire w_dff_B_gwLsbmn47_0;
	wire w_dff_B_gfgEgEin8_0;
	wire w_dff_B_BkkvnJa04_0;
	wire w_dff_B_pi3bOMe96_0;
	wire w_dff_B_Gf4T2pe65_0;
	wire w_dff_B_1b6BJ2b44_0;
	wire w_dff_A_Ga6sOL0g0_0;
	wire w_dff_A_AmZchLaN3_0;
	wire w_dff_A_5DV6LkPy1_0;
	wire w_dff_A_bB5nYlHV7_0;
	wire w_dff_A_lTP63Spd9_0;
	wire w_dff_A_YDMzKWpx9_0;
	wire w_dff_A_QD945d3m7_0;
	wire w_dff_A_lbsv0ReK6_0;
	wire w_dff_B_c86NDLmv7_0;
	wire w_dff_B_llIEBgxY1_0;
	wire w_dff_B_mgGvZFKz3_0;
	wire w_dff_B_DKuPd3Q95_0;
	wire w_dff_B_x8TsiQby5_0;
	wire w_dff_B_WY0rg8lq3_0;
	wire w_dff_B_N8nNB1em7_0;
	wire w_dff_B_wgb1a7W06_0;
	wire w_dff_B_SjL1xJhq7_0;
	wire w_dff_B_fXQYtvhd2_0;
	wire w_dff_B_Pwkrnbqn8_0;
	wire w_dff_B_mPKyzr5A0_0;
	wire w_dff_B_OmmcV7zM7_0;
	wire w_dff_B_8uskkqVH8_0;
	wire w_dff_B_9GS9SIJm4_0;
	wire w_dff_B_BxP2vLRX4_0;
	wire w_dff_B_bfCgYGGY8_0;
	wire w_dff_B_XBCxwza53_0;
	wire w_dff_B_7z8UO4ak4_0;
	wire w_dff_B_TMykp1pR1_0;
	wire w_dff_B_o59bURzk6_0;
	wire w_dff_B_C4GUCiLi4_0;
	wire w_dff_A_etCgCDAc9_2;
	wire w_dff_B_QXbdTfSC4_0;
	wire w_dff_B_yDMjWOG83_0;
	wire w_dff_B_A7VHVmSN2_0;
	wire w_dff_B_FJNmdIq07_0;
	wire w_dff_B_KEzPG80v8_0;
	wire w_dff_B_Z3nKmgEY0_0;
	wire w_dff_B_yPKn7UWd1_0;
	wire w_dff_B_HDBGGIma9_0;
	wire w_dff_B_gh5w2VDO3_0;
	wire w_dff_B_1CYes5n85_0;
	wire w_dff_B_JcqG57Ro5_0;
	wire w_dff_A_r7GzCRg66_0;
	wire w_dff_A_uLwnQKui8_1;
	wire w_dff_B_SbPu66re4_0;
	wire w_dff_B_Zf9fuJPj0_0;
	wire w_dff_B_2YVle0hT3_0;
	wire w_dff_B_43EMR9wJ7_0;
	wire w_dff_B_dTkXopeo5_0;
	wire w_dff_B_8kSi8rGV7_0;
	wire w_dff_B_uMNth0T19_0;
	wire w_dff_B_bTZDVqR75_0;
	wire w_dff_B_wkyzqvan1_0;
	wire w_dff_B_7IdryhxC2_0;
	wire w_dff_B_c47yMk2V7_0;
	wire w_dff_B_tRGiG3Pb4_0;
	wire w_dff_B_IHVmLyWb3_2;
	wire w_dff_B_UaLU43c64_2;
	wire w_dff_B_NPBlv3NP1_2;
	wire w_dff_A_LpkRCZlm5_0;
	wire w_dff_A_1Rm34mUJ6_0;
	wire w_dff_A_TExLgcsK5_0;
	wire w_dff_B_z2ueqf6J2_0;
	wire w_dff_B_RP8ZKKAf4_0;
	wire w_dff_B_mZBKS0aB4_1;
	wire w_dff_B_woAQXQKr3_1;
	wire w_dff_B_g8h89HDW9_1;
	wire w_dff_B_cRPOVfjX1_0;
	wire w_dff_A_kiedNMSw1_0;
	wire w_dff_A_hn1tQkK67_0;
	wire w_dff_A_WGusxvTa4_0;
	wire w_dff_A_3nXvSp6U4_0;
	wire w_dff_A_696SBWZe9_0;
	wire w_dff_A_PyIf5qVQ1_0;
	wire w_dff_B_Jp14vPOY8_0;
	wire w_dff_B_Grvczgnb2_0;
	wire w_dff_B_9QgfQnwM9_0;
	wire w_dff_B_E90BmrV45_0;
	wire w_dff_B_LHxyY0hH1_0;
	wire w_dff_B_HpKf3Jb22_0;
	wire w_dff_B_HM2nPqvS0_1;
	wire w_dff_B_4XQltSQF7_1;
	wire w_dff_B_X0msDUlY1_1;
	wire w_dff_B_bxr6B7Pd8_0;
	wire w_dff_A_kqaLlRCo8_0;
	wire w_dff_B_QRZS0TQ75_1;
	wire w_dff_B_nxN2Esor1_1;
	wire w_dff_B_wtqKpTH95_1;
	wire w_dff_B_4Us65xLQ6_1;
	wire w_dff_B_SeCdQpjF7_0;
	wire w_dff_B_GsZTZZTF3_0;
	wire w_dff_B_DoSOZjuk2_0;
	wire w_dff_B_oGIWPZO36_0;
	wire w_dff_B_GVcn3f3y3_0;
	wire w_dff_B_blczhI4C9_0;
	wire w_dff_B_BtGuEXDp7_0;
	wire w_dff_B_nPwJ4cy59_0;
	wire w_dff_B_Cv6Jnwn13_0;
	wire w_dff_B_ICQv7vJ08_0;
	wire w_dff_B_HXNCn4GD1_0;
	wire w_dff_B_iHtaYKnk5_2;
	wire w_dff_B_IIOCkE468_2;
	wire w_dff_B_NXJzxM3B9_2;
	wire w_dff_B_2i2NURNA2_1;
	wire w_dff_B_R4LcYWub1_1;
	wire w_dff_B_NZQc0blX1_1;
	wire w_dff_A_nclew3Bq1_1;
	wire w_dff_A_dMEordML7_1;
	wire w_dff_B_F0IHH1581_0;
	wire w_dff_B_ndd83xYU6_0;
	wire w_dff_A_Q1pMjrZr8_0;
	wire w_dff_B_hkjOxdZj3_0;
	wire w_dff_B_5M6LyKYf2_0;
	wire w_dff_B_06dd8j4n1_0;
	wire w_dff_B_eM3WcKdS2_0;
	wire w_dff_B_OfAy3uSm0_0;
	wire w_dff_B_eT3Orvrj8_1;
	wire w_dff_B_2Nbdvzzq5_1;
	wire w_dff_B_4LuH5Jpo9_1;
	wire w_dff_B_HTcQ0nIP8_0;
	wire w_dff_B_fSP7FxFs7_0;
	wire w_dff_A_mZmQW8xh3_1;
	wire w_dff_A_h9YeP2SC0_0;
	wire w_dff_A_GBysIiG21_0;
	wire w_dff_A_2G2UlGTq2_0;
	wire w_dff_A_ixpkdBVh1_0;
	wire w_dff_A_h27SHOlY8_1;
	wire w_dff_A_cSz0DHgh1_1;
	wire w_dff_A_eqRDN5xA8_1;
	wire w_dff_A_brxb91Nl9_1;
	wire w_dff_B_jXja1grm6_0;
	wire w_dff_B_qQQQr57e4_0;
	wire w_dff_B_ChStDK2h5_0;
	wire w_dff_B_i1TJoECv1_0;
	wire w_dff_B_9UhDffR76_0;
	wire w_dff_B_hyVTKsxV8_0;
	wire w_dff_B_43etQwju5_0;
	wire w_dff_B_dmuBxmgh2_0;
	wire w_dff_B_n35d1YZH7_0;
	wire w_dff_B_wtTfk3g40_0;
	wire w_dff_B_lGjRA1MP6_0;
	wire w_dff_B_F85S2bmz5_2;
	wire w_dff_B_brbJCPoz3_2;
	wire w_dff_B_tDQP5nyd7_2;
	wire w_dff_B_B4AvEkKb9_0;
	wire w_dff_B_AIv8lL129_1;
	wire w_dff_B_9j0d0Nud2_1;
	wire w_dff_B_UnolPSSa7_1;
	wire w_dff_B_JsUpw6qs3_0;
	wire w_dff_A_mrTqWM7Y8_0;
	wire w_dff_A_7dbIcJVQ6_0;
	wire w_dff_A_lJ4K7l0o8_0;
	wire w_dff_B_loTIAKmz0_0;
	wire w_dff_B_932T30un2_0;
	wire w_dff_B_xnOx4Plp4_0;
	wire w_dff_B_ZxEwx3is0_0;
	wire w_dff_B_cPsXwyo38_0;
	wire w_dff_B_UhDPWxwS4_1;
	wire w_dff_B_h5xBjHl44_1;
	wire w_dff_B_oY61uKLk2_1;
	wire w_dff_A_eGdNV9IC6_1;
	wire w_dff_B_ADAxB4i80_0;
	wire w_dff_A_MkzCM3QZ5_0;
	wire w_dff_B_AemQpIVj9_0;
	wire w_dff_B_xK6VGpEU5_0;
	wire w_dff_B_YWZeFU5n3_0;
	wire w_dff_B_d6uNA6YY6_0;
	wire w_dff_B_EXi4GZeS8_0;
	wire w_dff_B_vD5Fk35Y5_0;
	wire w_dff_B_t9tYVirr1_0;
	wire w_dff_B_VziqwfyY0_0;
	wire w_dff_B_uMuZL7Bd4_0;
	wire w_dff_B_Uf2LOJKb1_0;
	wire w_dff_B_AdB8vm2y9_0;
	wire w_dff_B_uA3DEimy4_2;
	wire w_dff_B_HDXzGdZK7_2;
	wire w_dff_B_EHofCk4u4_2;
	wire w_dff_A_dpCZoQk20_0;
	wire w_dff_A_7luvimY03_1;
	wire w_dff_B_mE0h48r77_0;
	wire w_dff_B_IGABrCwK7_0;
	wire w_dff_B_pNgu8r555_1;
	wire w_dff_B_H8s9gCkA2_1;
	wire w_dff_B_1BQvMScw8_0;
	wire w_dff_A_tduSDlpK3_0;
	wire w_dff_B_4emycJed9_1;
	wire w_dff_A_iBioveLm8_2;
	wire w_dff_A_UOES35z51_2;
	wire w_dff_B_luKw20Og5_3;
	wire w_dff_A_scjTpqwT0_2;
	wire w_dff_B_m6qwZRr16_0;
	wire w_dff_B_3R4wQPxn7_0;
	wire w_dff_B_c5I1m2YB9_0;
	wire w_dff_B_Lo8OStMm4_0;
	wire w_dff_B_I14rXkob3_0;
	wire w_dff_B_VWz7lHXZ8_1;
	wire w_dff_B_O9QHLiIa6_1;
	wire w_dff_B_HRMR7rpT2_1;
	wire w_dff_B_99e8Gtle2_0;
	wire w_dff_A_cp2V9q6e7_0;
	wire w_dff_B_epkIxhZs3_0;
	wire w_dff_B_3B64H4dF4_0;
	wire w_dff_B_sGff82Uf3_0;
	wire w_dff_A_CocBSnos7_0;
	wire w_dff_A_xUYhHAIk5_0;
	wire w_dff_B_SSfT7VwG3_0;
	wire w_dff_B_t67Rp19n4_0;
	wire w_dff_B_Z8j8lMpG2_0;
	wire w_dff_B_DcnYlsUl8_0;
	wire w_dff_B_WPf4cHkf0_0;
	wire w_dff_B_WNZNiIJS5_0;
	wire w_dff_B_9alznzrA7_1;
	wire w_dff_B_iXCOEUcA2_1;
	wire w_dff_B_8iUufvxb4_1;
	wire w_dff_B_9Rj5hHeL6_0;
	wire w_dff_B_BDmvZIaY5_0;
	wire w_dff_B_evefBOMY8_0;
	wire w_dff_B_cezlCk7Y4_0;
	wire w_dff_B_MIcPi9al6_0;
	wire w_dff_B_tnAQ7MbG3_0;
	wire w_dff_B_zqUFj38Q5_0;
	wire w_dff_B_QikZCtSI9_0;
	wire w_dff_B_ROAuJexP8_0;
	wire w_dff_B_skaBgWq53_1;
	wire w_dff_A_gaSKnasO8_0;
	wire w_dff_A_EI7ad8R13_0;
	wire w_dff_A_WrcUgB0F1_0;
	wire w_dff_A_67RcbT2e6_0;
	wire w_dff_A_c1SIEnVh5_0;
	wire w_dff_A_FvB3tIyx2_0;
	wire w_dff_A_ySM5rlIz0_0;
	wire w_dff_A_GycpXLU83_0;
	wire w_dff_A_629NqC8a0_0;
	wire w_dff_A_YnPLfKPy1_2;
	wire w_dff_A_DGr94NIX6_2;
	wire w_dff_A_55gpo2Ti6_2;
	wire w_dff_A_Rz7TMaaL4_2;
	wire w_dff_A_h6fIR9He3_2;
	wire w_dff_A_hqjnQ6OE8_2;
	wire w_dff_A_Ju0cGdxc2_2;
	wire w_dff_A_0meZ6t1G5_2;
	wire w_dff_A_jO3GpOIl5_2;
	wire w_dff_A_YCUoHJmc3_2;
	wire w_dff_A_qfKdnG4t3_0;
	wire w_dff_A_A3E73v3x3_0;
	wire w_dff_A_zQxJxC6H6_0;
	wire w_dff_A_arJIqD5j3_0;
	wire w_dff_A_m80uWGCS8_0;
	wire w_dff_A_F3dasG4b4_0;
	wire w_dff_B_88yunF5y9_2;
	wire w_dff_B_UOzhcatG6_2;
	wire w_dff_B_OsXxBvxJ0_1;
	wire w_dff_B_cIa0RRGx9_0;
	wire w_dff_B_myBjpaiO4_0;
	wire w_dff_B_ryzSXgLC1_0;
	wire w_dff_A_OpW0ntUi9_0;
	wire w_dff_B_1wrzx3hs6_1;
	wire w_dff_A_GfxdPqk05_0;
	wire w_dff_B_PK1nw0l90_1;
	wire w_dff_B_Qqtg0nxm7_0;
	wire w_dff_B_KLnd0Szl5_1;
	wire w_dff_B_ImVXIuGq5_1;
	wire w_dff_B_XFaalHQD9_1;
	wire w_dff_B_9t3Iv5XK3_0;
	wire w_dff_B_mqvQ6SXx6_1;
	wire w_dff_B_F4wIN6jS5_0;
	wire w_dff_A_6gJRWWHu3_0;
	wire w_dff_B_VurSCaJD9_0;
	wire w_dff_A_5cIVWmKE3_0;
	wire w_dff_A_8SlZqIuw7_0;
	wire w_dff_A_oLBtXOd74_0;
	wire w_dff_A_ZzUXv6Dg6_0;
	wire w_dff_B_mfm0ebpX6_1;
	wire w_dff_B_lpWqvyMa2_0;
	wire w_dff_B_c1NEaN4f0_0;
	wire w_dff_A_wLOdru9x4_0;
	wire w_dff_B_0HVgotjO2_0;
	wire w_dff_B_nAmKSWzQ8_0;
	wire w_dff_B_pwZfNd2I0_0;
	wire w_dff_B_T5Qe86438_0;
	wire w_dff_B_SyZgZmfS3_0;
	wire w_dff_B_sJ1EqXTQ3_0;
	wire w_dff_B_F0CJDHJM1_0;
	wire w_dff_B_n1ggcqH11_0;
	wire w_dff_B_95K4cv8e4_0;
	wire w_dff_B_S8poXftF0_0;
	wire w_dff_B_lcRHJFF64_0;
	wire w_dff_B_e8e7yQGH2_0;
	wire w_dff_B_XuaI41C61_0;
	wire w_dff_B_YVGo4UPM2_0;
	wire w_dff_B_Fb5Ls2ud3_0;
	wire w_dff_B_20IF8xx75_0;
	wire w_dff_B_aUdnxN211_0;
	wire w_dff_B_baLZapjS5_0;
	wire w_dff_B_ubwNbGnP8_0;
	wire w_dff_B_K8fPladJ7_0;
	wire w_dff_B_ydNagheH1_0;
	wire w_dff_B_B8ShOeCI8_0;
	wire w_dff_B_lBEKmMGR7_0;
	wire w_dff_B_D1GTF7xj2_0;
	wire w_dff_B_9zaiP92j1_2;
	wire w_dff_B_UnAOanOz8_2;
	wire w_dff_B_THH2YkVh9_2;
	wire w_dff_B_gsB4FoXm1_0;
	wire w_dff_B_4kLkfKo12_0;
	wire w_dff_B_21ZpFLLb4_0;
	wire w_dff_B_CMEIqyEC2_0;
	wire w_dff_B_IZhbXuXO6_0;
	wire w_dff_B_CHzR3QmG2_0;
	wire w_dff_B_PtJene9p6_0;
	wire w_dff_B_7UMCqO7y1_0;
	wire w_dff_B_3ZkuFiEy8_0;
	wire w_dff_B_bNuuCorj1_0;
	wire w_dff_B_9lyVfhjn2_0;
	wire w_dff_B_jdyTFGON9_0;
	wire w_dff_B_f93g6uv19_0;
	wire w_dff_B_K6eGth8v6_0;
	wire w_dff_B_KEvTavOV0_0;
	wire w_dff_B_6ZmFjkKK2_0;
	wire w_dff_B_XSqPl3ZV0_0;
	wire w_dff_B_zBWmmBda7_0;
	wire w_dff_B_RUW842451_0;
	wire w_dff_B_8pYaD5ov0_0;
	wire w_dff_B_QArQyq8Q0_0;
	wire w_dff_B_EXBGyFM30_0;
	wire w_dff_B_xfouMmUx8_0;
	wire w_dff_B_YBXa6sB24_0;
	wire w_dff_B_8J0lArrZ8_0;
	wire w_dff_A_2X5lSC9C7_0;
	wire w_dff_B_wrLMei2Q8_0;
	wire w_dff_B_YxTIEnT70_0;
	wire w_dff_B_XS8AGY9p0_0;
	wire w_dff_B_YT8gJEJV1_0;
	wire w_dff_B_hn1epTdc7_0;
	wire w_dff_B_WCGhpb738_0;
	wire w_dff_B_Sr29IMGI0_0;
	wire w_dff_B_OAWvXCb19_0;
	wire w_dff_B_W7QiUbOv5_0;
	wire w_dff_B_c5Wf58tx4_0;
	wire w_dff_B_8H9Nxs8R9_0;
	wire w_dff_B_zrm5P10X0_0;
	wire w_dff_B_6M8cMGMJ4_0;
	wire w_dff_B_By08MlUX8_0;
	wire w_dff_B_bfR9spID6_0;
	wire w_dff_B_5NMMGf1M8_0;
	wire w_dff_B_SuUkj5c21_0;
	wire w_dff_B_OENpHhtD4_0;
	wire w_dff_B_uXsAf7yt8_0;
	wire w_dff_B_so6IUW984_0;
	wire w_dff_B_xRaaIIR30_0;
	wire w_dff_B_GPFUh6Jo5_0;
	wire w_dff_B_hDZQT4wf6_0;
	wire w_dff_B_5zdEAoKI9_0;
	wire w_dff_B_eTqwgJac6_0;
	wire w_dff_B_V3RaC9xA7_0;
	wire w_dff_B_NNNAuk3Y0_2;
	wire w_dff_B_nGik8l1A5_2;
	wire w_dff_B_19FnkAzX5_2;
	wire w_dff_B_NNKyvdJ29_0;
	wire w_dff_B_5Tx3Shrb9_0;
	wire w_dff_B_LqaCsD8p8_0;
	wire w_dff_B_mO9xCXNt0_0;
	wire w_dff_B_7lA60dox5_0;
	wire w_dff_B_LRZkUum75_0;
	wire w_dff_B_9at1ByCj6_0;
	wire w_dff_B_LR86h8DS1_0;
	wire w_dff_B_hfsJQ9OX6_0;
	wire w_dff_B_MyhW5Q118_0;
	wire w_dff_B_ZMGHqk8a6_0;
	wire w_dff_B_qLP4lseT5_0;
	wire w_dff_B_f6ms2hRU9_0;
	wire w_dff_B_jRX7vECG9_2;
	wire w_dff_B_O70naEaZ5_2;
	wire w_dff_B_8Yyyj7RI1_2;
	wire w_dff_A_SjmIzxNS3_0;
	wire w_dff_B_oEHMjoZM4_0;
	wire w_dff_B_0UVXI1LF8_0;
	wire w_dff_B_1JF1dcMV9_0;
	wire w_dff_B_qlGZLACm0_0;
	wire w_dff_B_o3RAEwwq5_0;
	wire w_dff_B_GIm0chOL1_0;
	wire w_dff_B_m7Qul1kx6_0;
	wire w_dff_B_QU5O1tk84_0;
	wire w_dff_B_blxjcLSa4_0;
	wire w_dff_B_ojJnp0J70_0;
	wire w_dff_B_kBUkPofw5_0;
	wire w_dff_B_T1l0oZsW6_0;
	wire w_dff_B_d8DnDGOF9_0;
	wire w_dff_B_q20txiL02_0;
	wire w_dff_B_zXfMPo1R6_2;
	wire w_dff_B_MQq2MLku5_2;
	wire w_dff_B_kYuYIcMt3_2;
	wire w_dff_B_ZOzHQm2o8_0;
	wire w_dff_B_ERsYOr3c9_0;
	wire w_dff_B_m3koI63o4_0;
	wire w_dff_B_uzBL3Vhi0_0;
	wire w_dff_B_5xB5dWrk5_0;
	wire w_dff_B_5xbZSuV02_0;
	wire w_dff_B_ICvipmzU5_0;
	wire w_dff_B_wmcbES5X2_0;
	wire w_dff_B_5jxlTNV85_0;
	wire w_dff_B_njHTkLKH5_0;
	wire w_dff_B_2dSk21kk0_0;
	wire w_dff_B_6swa5yUS6_0;
	wire w_dff_B_Lv9JQ9Y06_0;
	wire w_dff_B_Cx88I4iO0_0;
	wire w_dff_A_vITD7vPb0_0;
	wire w_dff_A_WbwDnkIO3_0;
	wire w_dff_A_8JoHe52a3_0;
	wire w_dff_B_lbHHsTzM8_0;
	wire w_dff_B_b5kwYdD60_0;
	wire w_dff_B_Uw33huRr7_0;
	wire w_dff_B_vLBJNzGY0_0;
	wire w_dff_B_iA9bVtkV3_0;
	wire w_dff_B_NsB6g8zc0_0;
	wire w_dff_B_4wiyKpNu5_0;
	wire w_dff_B_0rJSfrYf8_0;
	wire w_dff_B_Wue1VuDB7_0;
	wire w_dff_B_DbWznKL27_0;
	wire w_dff_B_gPUORSrF9_0;
	wire w_dff_B_xcUtQedf4_0;
	wire w_dff_B_BgYH8FIF4_0;
	wire w_dff_B_Ng6Rn8W99_0;
	wire w_dff_B_U6uAs9no9_0;
	wire w_dff_B_7Wj7KvJt5_0;
	wire w_dff_B_V0vbzK4e1_0;
	wire w_dff_B_NsRBJ3iU3_0;
	wire w_dff_B_zNKGFW5e9_0;
	wire w_dff_B_zV1Q3ny67_0;
	wire w_dff_B_TQMcUYh46_0;
	wire w_dff_B_9i2GNllg1_0;
	wire w_dff_B_XGpEbwUZ0_0;
	wire w_dff_B_fdPo0AZw9_0;
	wire w_dff_B_2NvQOqmD9_0;
	wire w_dff_A_rrTVTbpo5_2;
	wire w_dff_A_BdZzNksn6_1;
	wire w_dff_A_BWQGC92m1_2;
	wire w_dff_A_ECbPHj9f5_2;
	wire w_dff_B_gOi5EzOj8_0;
	wire w_dff_B_EtmPvepO1_0;
	wire w_dff_B_G2h9uHxD4_0;
	wire w_dff_B_F4yeVIzN2_0;
	wire w_dff_B_ayUldVDk7_0;
	wire w_dff_B_weEEwUjX6_0;
	wire w_dff_B_A0rIVWEu8_0;
	wire w_dff_B_8KsF5R416_0;
	wire w_dff_B_yoXsPQ4H1_0;
	wire w_dff_B_Lu8lYJLh5_0;
	wire w_dff_B_iU3KJzgu0_0;
	wire w_dff_B_o5e6IOru5_0;
	wire w_dff_A_8i5JmseF1_2;
	wire w_dff_B_oedsz4iZ2_0;
	wire w_dff_B_hw9IJ1Bl2_0;
	wire w_dff_B_x5UCoTEU2_0;
	wire w_dff_B_NLSYKpBl1_0;
	wire w_dff_B_plyQ8HPL6_0;
	wire w_dff_B_1U7ck2i94_0;
	wire w_dff_B_feDNCScj2_0;
	wire w_dff_B_yefaxNen0_0;
	wire w_dff_B_visyYMWp4_0;
	wire w_dff_B_j9G7auJy6_0;
	wire w_dff_B_NgGmCUIL6_0;
	wire w_dff_B_Krh0mYAU6_0;
	wire w_dff_B_tiqgSRIB6_0;
	wire w_dff_B_4PSQfdGY6_0;
	wire w_dff_B_YPRdsmVb0_2;
	wire w_dff_B_kI74GGDN6_2;
	wire w_dff_B_dLHRqh202_2;
	wire w_dff_B_eFZn4Thj1_0;
	wire w_dff_B_LJAJG16A1_0;
	wire w_dff_B_JeW58ZwZ2_0;
	wire w_dff_B_AMqtIJq76_0;
	wire w_dff_B_SiShHYSa7_0;
	wire w_dff_B_rriyiCdb7_1;
	wire w_dff_B_QskXEO8H8_1;
	wire w_dff_B_E0lFfosK4_1;
	wire w_dff_B_Vz1ntBHV2_0;
	wire w_dff_B_6B5mhpyF8_0;
	wire w_dff_B_zhPGh3cK0_0;
	wire w_dff_B_eAaYpwze3_0;
	wire w_dff_B_COuRIf2v1_0;
	wire w_dff_B_dtmJ3N519_0;
	wire w_dff_B_ISnxJlzE9_0;
	wire w_dff_B_LaggcDo98_0;
	wire w_dff_B_1XCOXLIU0_1;
	wire w_dff_B_PYLWk6ka0_1;
	wire w_dff_B_JdJmN8DZ9_1;
	wire w_dff_B_SlI5zjop1_0;
	wire w_dff_B_acpYoPnv5_0;
	wire w_dff_B_fzyS4ZHU6_0;
	wire w_dff_B_faGCYL2X9_0;
	wire w_dff_B_whRg3B451_0;
	wire w_dff_B_WqSqG6bc3_0;
	wire w_dff_B_YmxtpP3m7_0;
	wire w_dff_B_5eds7RG33_0;
	wire w_dff_B_udGgoTHc8_0;
	wire w_dff_B_hERHpCd72_0;
	wire w_dff_B_Gh8s5APZ8_0;
	wire w_dff_B_PCWCeHBx3_0;
	wire w_dff_B_Eeolb1wv2_0;
	wire w_dff_B_vy9ULEa11_0;
	wire w_dff_B_hpxdS3QY5_2;
	wire w_dff_B_MFi49ebU8_2;
	wire w_dff_B_rCprmroI2_2;
	wire w_dff_B_GMkp0s0z6_0;
	wire w_dff_B_Pp4FAqis2_0;
	wire w_dff_B_mhjMIrs43_0;
	wire w_dff_B_D43eyW007_0;
	wire w_dff_B_lyCXxF103_1;
	wire w_dff_B_Olgdvryu5_1;
	wire w_dff_B_R5eMOqaD7_1;
	wire w_dff_A_rIWRxbCO5_1;
	wire w_dff_A_05jXUVYb5_1;
	wire w_dff_B_AbC2ilUe7_1;
	wire w_dff_B_JRvU0wqr5_1;
	wire w_dff_B_KRYrmHnS6_1;
	wire w_dff_B_jfGC3CN29_1;
	wire w_dff_B_raw05elo1_0;
	wire w_dff_B_HH4FIpVi3_0;
	wire w_dff_B_IEpRikXA7_0;
	wire w_dff_B_3pjLBGFh6_0;
	wire w_dff_B_nXu5OdZo0_0;
	wire w_dff_B_3iC6jjnK9_0;
	wire w_dff_B_XiAZqJNi4_0;
	wire w_dff_B_UrrZoGXb3_1;
	wire w_dff_B_8aI5nUHz3_1;
	wire w_dff_B_EreY5MCq2_1;
	wire w_dff_B_VcxDnBYM0_0;
	wire w_dff_A_jmZ7L2ae0_1;
	wire w_dff_A_wjn5Vn6R9_1;
	wire w_dff_B_Dgj4G4vl7_1;
	wire w_dff_B_zWvbwJsk7_1;
	wire w_dff_B_fjTAuQFX2_1;
	wire w_dff_B_p7N3tSMZ1_1;
	wire w_dff_B_1B5dW4gv3_1;
	wire w_dff_B_U8qdlVqH8_1;
	wire w_dff_B_B2VgIguc1_1;
	wire w_dff_B_0RClE1oJ5_1;
	wire w_dff_B_5MI8Awnl5_1;
	wire w_dff_B_5Z2NNARz1_1;
	wire w_dff_B_z4wiDlmQ1_1;
	wire w_dff_B_WREghjRO3_1;
	wire w_dff_B_Tmuo6mTq9_1;
	wire w_dff_B_rNTWf0vb8_1;
	wire w_dff_A_WqzXDVaw3_1;
	wire w_dff_A_6XXnUosv2_1;
	wire w_dff_A_mOrcPzMO3_1;
	wire w_dff_A_xnKGH3WI2_1;
	wire w_dff_A_fr2wMieK9_1;
	wire w_dff_A_PhT7RjdB1_1;
	wire w_dff_A_Hl0Q5VCh0_1;
	wire w_dff_A_z36PlgSe5_1;
	wire w_dff_A_fXiwjX984_1;
	wire w_dff_A_WRWLsXku9_2;
	wire w_dff_A_MXDRsjqQ0_2;
	wire w_dff_A_KJjsWf3F7_2;
	wire w_dff_A_zEXBvlxm0_2;
	wire w_dff_A_TNNwyAnz4_2;
	wire w_dff_A_sWLOdO185_2;
	wire w_dff_B_22OVXIZw7_0;
	wire w_dff_B_OeLX3bdT2_0;
	wire w_dff_B_pq6GNIyG0_0;
	wire w_dff_B_iDlfVGcF8_0;
	wire w_dff_B_qJPRHBPH9_0;
	wire w_dff_B_yP90QQdN5_0;
	wire w_dff_B_yJYsWwSD7_0;
	wire w_dff_B_pJYulsn07_0;
	wire w_dff_B_pJF4Jypo6_0;
	wire w_dff_B_SFnz6RF04_0;
	wire w_dff_B_TeA0l5RY6_0;
	wire w_dff_B_q8GF83v79_0;
	wire w_dff_B_U9xFB3tu4_2;
	wire w_dff_B_Q4LtkL6W1_2;
	wire w_dff_B_4OU2SCCW1_2;
	wire w_dff_B_dUgtlIFV2_0;
	wire w_dff_B_9xqbSwPw2_0;
	wire w_dff_B_zHdPq9Yi6_0;
	wire w_dff_B_JtyCeYB62_0;
	wire w_dff_B_A49QF9CZ7_0;
	wire w_dff_B_OSHN10nK3_1;
	wire w_dff_B_cnWEupaI2_1;
	wire w_dff_A_EQbq1Jpa1_1;
	wire w_dff_A_Fh9xh3C97_1;
	wire w_dff_A_zTdByzIN4_2;
	wire w_dff_A_GzU8HWgG0_2;
	wire w_dff_A_1hnT5ZfW1_1;
	wire w_dff_A_YzYrO1eU3_1;
	wire w_dff_A_fKMKsLFO5_1;
	wire w_dff_A_1sHSKFOe3_1;
	wire w_dff_A_Ubk7zqdW1_1;
	wire w_dff_A_DAWyJfAl7_1;
	wire w_dff_A_9d8L8x0H4_2;
	wire w_dff_A_SjxSNAMP4_2;
	wire w_dff_A_wCrRRJR36_2;
	wire w_dff_A_r18v1tHD8_0;
	wire w_dff_A_x23Z2iOW2_0;
	wire w_dff_A_sFJ45rlF1_0;
	wire w_dff_A_0Ocy39pC6_0;
	wire w_dff_A_hjZUStJG5_0;
	wire w_dff_A_SS5FoYVk2_0;
	wire w_dff_A_Hw5wbg2B0_1;
	wire w_dff_A_1fLKU9vB1_1;
	wire w_dff_A_KzcxDb729_2;
	wire w_dff_B_li6rMYPd0_0;
	wire w_dff_B_ARaiKiPd6_0;
	wire w_dff_B_3qpbMsdT4_0;
	wire w_dff_B_hx5DLAU38_0;
	wire w_dff_B_FjyRfDIm0_0;
	wire w_dff_B_tYWbr3Pe8_0;
	wire w_dff_B_y5jcS6ZD3_0;
	wire w_dff_B_GDnjo22a3_1;
	wire w_dff_B_nDROfitL5_1;
	wire w_dff_B_nyZz9qgn8_1;
	wire w_dff_B_VQfTMgXa2_0;
	wire w_dff_B_slQjwQXb7_3;
	wire w_dff_A_SAJWWZnn5_1;
	wire w_dff_A_Id5oNvbB0_2;
	wire w_dff_A_4jcnKlLF8_2;
	wire w_dff_A_GSkyqbtI8_1;
	wire w_dff_A_XRpTZvDQ0_2;
	wire w_dff_A_ENGhT1wc6_2;
	wire w_dff_A_vm4mmnSs7_0;
	wire w_dff_A_LW3Zr75J1_1;
	wire w_dff_B_M7SHGnkw8_0;
	wire w_dff_B_qtFJrn8I0_0;
	wire w_dff_B_8cBj3oOq5_0;
	wire w_dff_B_5c0bILSV0_0;
	wire w_dff_B_oTNeUFKQ7_0;
	wire w_dff_B_e8YAPToP2_0;
	wire w_dff_B_M4zknGzF3_0;
	wire w_dff_B_p9MjM4yu6_0;
	wire w_dff_B_xf6O3MZo7_0;
	wire w_dff_B_YAPnp2Q61_0;
	wire w_dff_B_yy97jijI8_0;
	wire w_dff_B_VdR7OR9Q3_0;
	wire w_dff_B_2SbTkK094_2;
	wire w_dff_B_TiplbXo39_2;
	wire w_dff_B_cpaVajUF2_2;
	wire w_dff_B_HfFaPkC65_0;
	wire w_dff_B_8XrlRDYx1_0;
	wire w_dff_B_O1Otu4Kr7_0;
	wire w_dff_B_ZkgHXbfY0_0;
	wire w_dff_B_BNivMpSa4_0;
	wire w_dff_B_tiF4XvPQ7_0;
	wire w_dff_B_qUG4y7cK7_0;
	wire w_dff_B_OMwLOQoe0_1;
	wire w_dff_A_1tQJNjSy6_1;
	wire w_dff_A_Pny1KaRT0_0;
	wire w_dff_B_PL0GQhlg7_2;
	wire w_dff_B_4bhq2NKq5_0;
	wire w_dff_A_8ttTp3Vi9_1;
	wire w_dff_A_gJmCSXsn7_0;
	wire w_dff_A_StlX5KTO3_0;
	wire w_dff_A_fw76MlPt4_0;
	wire w_dff_A_2pMiESGr0_0;
	wire w_dff_A_ro6qKbEt7_0;
	wire w_dff_A_6Dvk6O510_0;
	wire w_dff_A_J5FJNJKh7_0;
	wire w_dff_B_jDCZofNF4_2;
	wire w_dff_A_llMijzDi0_1;
	wire w_dff_A_WSi3kZeY5_1;
	wire w_dff_B_kiRT4vhG2_0;
	wire w_dff_B_g3wjCMSv3_0;
	wire w_dff_B_rsSuToCT0_0;
	wire w_dff_B_3gfUOwFb5_0;
	wire w_dff_B_OZTkSiqQ5_0;
	wire w_dff_B_RiEGixy43_0;
	wire w_dff_B_W7HNd5l65_0;
	wire w_dff_B_J5kFLssw3_0;
	wire w_dff_B_RJFQge1i7_0;
	wire w_dff_B_e9P0BzYN6_0;
	wire w_dff_B_0I6h65H62_1;
	wire w_dff_B_wxWIjnjD9_1;
	wire w_dff_A_ggzm7CIh2_2;
	wire w_dff_A_SGJuPREI6_2;
	wire w_dff_B_KTjZAv1M5_1;
	wire w_dff_B_vex8H1gp2_1;
	wire w_dff_B_XZUn9BKN5_1;
	wire w_dff_B_nrpAOopt1_1;
	wire w_dff_B_9viapTLL6_1;
	wire w_dff_B_IjVSjQ8n3_1;
	wire w_dff_B_6o6s6cOq5_1;
	wire w_dff_B_zFkwWUqm1_1;
	wire w_dff_B_W6tnOw9y0_1;
	wire w_dff_B_fQWhak0j7_1;
	wire w_dff_A_W5XI0bWh9_1;
	wire w_dff_A_WCcbNtYi1_1;
	wire w_dff_A_9sdbsVg40_1;
	wire w_dff_A_MNXxV7ES6_1;
	wire w_dff_B_TibwFOW81_3;
	wire w_dff_B_pX7f7LqH6_3;
	wire w_dff_B_gTmA6XQD6_3;
	wire w_dff_B_QjCsz9SH9_2;
	wire w_dff_B_RcmgbfyC8_2;
	wire w_dff_B_9EKcqnJ09_2;
	wire w_dff_B_bzelxDXV2_2;
	wire w_dff_B_VIoBQoCF0_2;
	wire w_dff_B_N3N1Y1jD7_2;
	wire w_dff_A_DxmC90yB9_1;
	wire w_dff_A_7X10HfUW9_2;
	wire w_dff_A_mgsbhz6J6_0;
	wire w_dff_A_m7oKYewi8_0;
	wire w_dff_A_JUZSiVxA0_0;
	wire w_dff_A_7nP5QKik0_0;
	wire w_dff_A_mgfZHYHO8_0;
	wire w_dff_A_mxBuZMhX9_0;
	wire w_dff_A_6jB4SwTD5_0;
	wire w_dff_A_K7Di0Uvu6_0;
	wire w_dff_A_cENZyIIS1_0;
	wire w_dff_A_HlGmURBk0_1;
	wire w_dff_A_HKYxXTwe9_1;
	wire w_dff_A_fUcf2fqC9_1;
	wire w_dff_A_shtfT2Pp1_1;
	wire w_dff_A_93Tmmsg90_1;
	wire w_dff_A_RIpPmYAd8_1;
	wire w_dff_B_i3FsJUr95_1;
	wire w_dff_B_fFwXDLlc1_1;
	wire w_dff_B_E3RDMGLX3_1;
	wire w_dff_B_uOuoRYtZ2_1;
	wire w_dff_B_NUJRDPGh3_1;
	wire w_dff_B_mtu0Bx9L3_1;
	wire w_dff_B_UcVSyL2i5_1;
	wire w_dff_B_e4YOXTGO5_1;
	wire w_dff_B_yxfhv4Fa6_1;
	wire w_dff_B_5zC0WoXC2_1;
	wire w_dff_B_LgoqLde44_1;
	wire w_dff_B_zAIAJcVN6_1;
	wire w_dff_B_B99ennDR0_0;
	wire w_dff_B_bFOj7a0R4_1;
	wire w_dff_B_6sM8oGHm0_1;
	wire w_dff_B_B1UYFk2o4_1;
	wire w_dff_B_Nq54T7Ky9_1;
	wire w_dff_B_QPDnPbRd3_1;
	wire w_dff_B_RauW5Vu18_1;
	wire w_dff_B_MJdzDbaa6_1;
	wire w_dff_B_EBoRtQx52_1;
	wire w_dff_B_fuFAjgps1_1;
	wire w_dff_B_zgPyu6ru9_1;
	wire w_dff_B_pbz0Cmqh4_1;
	wire w_dff_B_FtthFBnC9_1;
	wire w_dff_B_fPpq6yDu9_1;
	wire w_dff_B_wicwbTDi0_1;
	wire w_dff_B_Pyyd8abY6_1;
	wire w_dff_B_htnjqMlm6_0;
	wire w_dff_B_BGFZewS63_0;
	wire w_dff_B_5ctXP9eo4_0;
	wire w_dff_B_VkhQF9W88_0;
	wire w_dff_B_hdMl9aRK1_0;
	wire w_dff_B_8sUGvrK17_0;
	wire w_dff_B_nCk8U6TP4_0;
	wire w_dff_B_PRMxhqAJ0_0;
	wire w_dff_B_sjSsXpMB5_0;
	wire w_dff_B_e6Z5c8AC5_0;
	wire w_dff_B_JTD7njZr3_0;
	wire w_dff_B_FZlu4RZA7_0;
	wire w_dff_B_1M3YZdXG6_0;
	wire w_dff_B_KHEGqgld8_0;
	wire w_dff_B_qVVUs1qO2_0;
	wire w_dff_B_7vOvb3sI0_0;
	wire w_dff_B_1A9Un1F09_0;
	wire w_dff_B_VGR9opvU0_0;
	wire w_dff_A_Rhc3tDM80_1;
	wire w_dff_A_H3oBqD3L7_1;
	wire w_dff_A_xerHdk6D7_1;
	wire w_dff_A_ZgTFHJnh9_1;
	wire w_dff_A_f3qoZ7Cz7_1;
	wire w_dff_A_MYL3Ibh64_1;
	wire w_dff_A_ZFvdDV6w3_1;
	wire w_dff_A_RfCGG9Om0_2;
	wire w_dff_A_wid5fOrc7_2;
	wire w_dff_A_nVSbX7wO5_2;
	wire w_dff_A_eTvjzC3E2_2;
	wire w_dff_A_llyazwr65_2;
	wire w_dff_A_bAjPhM2N9_2;
	wire w_dff_A_k3WV8kxG7_1;
	wire w_dff_A_OYUtI3739_1;
	wire w_dff_A_rwkBpeNA8_1;
	wire w_dff_A_XqzPCH1w8_1;
	wire w_dff_A_QS2IeYwS3_1;
	wire w_dff_A_Zckhoghx0_2;
	wire w_dff_B_YSXjY3xx5_3;
	wire w_dff_B_HB2DzWmL0_3;
	wire w_dff_B_vpIeW4oQ2_3;
	wire w_dff_B_7IGwgqcQ8_3;
	wire w_dff_A_iUZuXxWP7_1;
	wire w_dff_A_VanVvJhj2_1;
	wire w_dff_A_CxN3yo6u0_1;
	wire w_dff_A_rFFwgffD7_1;
	wire w_dff_A_I9MJSD190_1;
	wire w_dff_A_QlZOPNq30_1;
	wire w_dff_A_bHmzluzP8_1;
	wire w_dff_A_jpRvdR2a4_1;
	wire w_dff_A_OqdiTg7f4_1;
	wire w_dff_A_2W8pSPwQ6_1;
	wire w_dff_A_lnjU3B0F6_2;
	wire w_dff_A_iq8ABI189_2;
	wire w_dff_A_E4OTRdCl7_2;
	wire w_dff_A_Uo3QZuGO4_2;
	wire w_dff_A_jJ6AozAY6_2;
	wire w_dff_A_8pvUP4jg8_2;
	wire w_dff_A_j7BaaYgz3_2;
	wire w_dff_A_1cCJGC275_1;
	wire w_dff_A_tbNhpOKQ3_1;
	wire w_dff_A_XbVu0WMF1_1;
	wire w_dff_A_u2MqTlpg8_1;
	wire w_dff_A_CLCfiF5u8_1;
	wire w_dff_A_l6LMCiKm3_2;
	wire w_dff_A_8Mno0JcQ7_2;
	wire w_dff_A_PDsmLccJ7_2;
	wire w_dff_A_1vCY42P70_2;
	wire w_dff_B_YmYQRpHf4_3;
	wire w_dff_B_B6H4VXy27_3;
	wire w_dff_B_gqD19LCf9_3;
	wire w_dff_B_NpdFLm1V0_3;
	wire w_dff_B_r4PTKkIp0_3;
	wire w_dff_B_W0wuerbt5_3;
	wire w_dff_A_D88n27GW8_2;
	wire w_dff_A_PjTDWTfI7_1;
	wire w_dff_B_IyXlR4hY7_0;
	wire w_dff_B_ZLtLf6e24_0;
	wire w_dff_B_qNgk59pk6_0;
	wire w_dff_B_3WrV56Wd1_0;
	wire w_dff_B_hOPT3Yyh1_0;
	wire w_dff_B_wnElaByr2_0;
	wire w_dff_B_JxVXYiaX8_0;
	wire w_dff_B_GV2db3OD6_0;
	wire w_dff_B_V0ZsOrIP0_0;
	wire w_dff_B_pVj1v5wW0_0;
	wire w_dff_B_YYdSncrK0_0;
	wire w_dff_B_7ckjdnBU4_0;
	wire w_dff_B_Gwk3KFCt9_0;
	wire w_dff_B_p1sY2Bkz6_0;
	wire w_dff_B_AEdSkG510_0;
	wire w_dff_B_2ozSsQQ30_0;
	wire w_dff_B_TbPXMdHi8_0;
	wire w_dff_B_wYeNHq3I4_2;
	wire w_dff_B_goR4it6E5_2;
	wire w_dff_B_Vi4narfa5_2;
	wire w_dff_A_4D4LeZGo5_1;
	wire w_dff_A_zdEm43ho5_1;
	wire w_dff_A_aOjiNL5O2_1;
	wire w_dff_A_y6ed07EG4_1;
	wire w_dff_A_gaCAXaqN9_1;
	wire w_dff_A_fCefUJbV9_1;
	wire w_dff_A_i6yV8PVe8_1;
	wire w_dff_A_iYlu67LX7_2;
	wire w_dff_A_BalXCdcn6_2;
	wire w_dff_A_Gxfq656C7_2;
	wire w_dff_A_CoexmRvB7_2;
	wire w_dff_A_zJTbukgA4_2;
	wire w_dff_A_8m2i4gXb4_2;
	wire w_dff_A_4joDZmYv9_1;
	wire w_dff_A_HnYLLHG05_1;
	wire w_dff_A_7Qp7UjoB4_1;
	wire w_dff_A_bramFFDL0_1;
	wire w_dff_A_EWrfPdBv2_1;
	wire w_dff_A_pPhhY0IA6_2;
	wire w_dff_B_IiAysqFu4_3;
	wire w_dff_B_PYX2lF964_3;
	wire w_dff_B_p5nMLCf24_3;
	wire w_dff_B_otVDLEHT6_3;
	wire w_dff_A_7LYzfzSD1_1;
	wire w_dff_A_3lQP8ya17_1;
	wire w_dff_A_3kuZopJo7_1;
	wire w_dff_A_b5vc8FTZ1_1;
	wire w_dff_A_6fhnPVYK1_1;
	wire w_dff_A_OdWhSluN0_1;
	wire w_dff_A_HBrApsK97_1;
	wire w_dff_A_m2wipF8h2_1;
	wire w_dff_A_byVzplzN1_1;
	wire w_dff_A_OAmdyT2Q3_1;
	wire w_dff_A_V1sULonp0_2;
	wire w_dff_A_LDDCOmTK7_2;
	wire w_dff_A_STwPZpN01_2;
	wire w_dff_A_w7rRNa1K2_2;
	wire w_dff_A_k8BHUIRL0_2;
	wire w_dff_A_6l0cAnec7_2;
	wire w_dff_A_2csyo9hG7_2;
	wire w_dff_A_K2lEsZEX3_1;
	wire w_dff_A_rOGRVMiY5_1;
	wire w_dff_A_YLqsyOWq0_1;
	wire w_dff_A_qr0LnxOY1_1;
	wire w_dff_A_uFGO2QA43_1;
	wire w_dff_A_sCQiNn1o4_2;
	wire w_dff_A_KFFPcOaf4_2;
	wire w_dff_A_xGvSj7hy3_2;
	wire w_dff_A_225P8l8c2_2;
	wire w_dff_B_tBgkUl0I6_3;
	wire w_dff_B_hr7FeO4t4_3;
	wire w_dff_B_VSUl2bQH4_3;
	wire w_dff_B_SwqRqUfg5_3;
	wire w_dff_B_eS2njwbW0_3;
	wire w_dff_B_47vXz1si6_3;
	wire w_dff_A_oD4ZL31J1_1;
	wire w_dff_A_CfNDWJtS0_2;
	wire w_dff_B_sNBr3ATY3_0;
	wire w_dff_B_eBSRsZqY1_0;
	wire w_dff_B_okrWZa0i1_0;
	wire w_dff_B_OS5yAMzL9_0;
	wire w_dff_B_uzvCX6Ce6_0;
	wire w_dff_B_I8A9TEcj2_0;
	wire w_dff_B_mcHwpzJl9_0;
	wire w_dff_B_mawCYAhC3_0;
	wire w_dff_B_lzhpR4z89_0;
	wire w_dff_B_Y33MBaP45_0;
	wire w_dff_B_uGuT4d9i7_0;
	wire w_dff_B_7OXd0QYL8_0;
	wire w_dff_B_iLAdrS1b7_1;
	wire w_dff_B_BvUgjQVi0_1;
	wire w_dff_B_hZ2QxyWZ5_1;
	wire w_dff_B_maOVicp01_1;
	wire w_dff_B_ABCI4f7I3_1;
	wire w_dff_B_HWHU7TwK8_1;
	wire w_dff_B_f0LutFs85_1;
	wire w_dff_B_o2ZrxLxI2_1;
	wire w_dff_B_GfeBdrXb4_1;
	wire w_dff_B_e89mvSKZ7_1;
	wire w_dff_B_fWsQXXrF4_1;
	wire w_dff_B_VaxEOFz65_1;
	wire w_dff_A_2u9BSIhp7_0;
	wire w_dff_A_DdmFGqHt5_0;
	wire w_dff_A_dJaYxjqo6_0;
	wire w_dff_A_pWkXD5lq7_0;
	wire w_dff_A_YGRwvE6t0_2;
	wire w_dff_A_cw52e6LO7_2;
	wire w_dff_A_pBaM6wMA7_2;
	wire w_dff_A_z0Jg1tsc0_2;
	wire w_dff_A_TjEuZVEy3_2;
	wire w_dff_A_zWFcKXYn6_2;
	wire w_dff_A_82wkT1EN3_2;
	wire w_dff_A_QsdVDy8B5_2;
	wire w_dff_A_m3SICdOU5_2;
	wire w_dff_A_7RiZXL4r0_1;
	wire w_dff_A_ZItrffyO1_1;
	wire w_dff_A_Cm1cGdOU7_1;
	wire w_dff_A_5o8TgSOR1_1;
	wire w_dff_A_PknUmGKH2_1;
	wire w_dff_A_Pl6plcCR9_1;
	wire w_dff_A_Fo2TcyFP3_1;
	wire w_dff_A_eKpMuOXE5_1;
	wire w_dff_A_oWhN8KOx3_1;
	wire w_dff_A_052EMNkd0_2;
	wire w_dff_A_fknCMaa94_2;
	wire w_dff_A_4rJKj9vY1_2;
	wire w_dff_A_1KKrVCTr9_2;
	wire w_dff_A_rMbDKlHt8_2;
	wire w_dff_B_0KlNMVYb2_1;
	wire w_dff_B_aojd7tuv2_1;
	wire w_dff_B_trfTZQBd9_1;
	wire w_dff_B_wxInqJFz6_1;
	wire w_dff_B_00lEdccQ8_1;
	wire w_dff_B_tlznQ9Nw9_1;
	wire w_dff_B_o4aJ5EZ73_1;
	wire w_dff_B_72JzGlTT8_1;
	wire w_dff_B_QeCboIuJ4_1;
	wire w_dff_B_uKF5PvQs8_1;
	wire w_dff_B_Ft5VBjlW8_1;
	wire w_dff_B_VBe4Pi9L6_1;
	wire w_dff_B_41iV7Vct0_1;
	wire w_dff_B_jecj7M9W1_1;
	wire w_dff_A_adHWuCeE4_0;
	wire w_dff_A_leLUn6aC2_0;
	wire w_dff_A_NMvM3QNc1_0;
	wire w_dff_A_sHkldfAJ2_0;
	wire w_dff_A_kN3KSB2c5_0;
	wire w_dff_A_YSPdOOlB5_0;
	wire w_dff_A_oYXk3jmS2_2;
	wire w_dff_A_OwsF0eaN9_2;
	wire w_dff_A_hNECWQIm3_2;
	wire w_dff_A_GG3wOGg22_2;
	wire w_dff_A_dszaMtZc7_2;
	wire w_dff_A_NjS41Zuc0_2;
	wire w_dff_A_BOsRK9m87_2;
	wire w_dff_A_UclOCWtG6_2;
	wire w_dff_A_qiAxdV336_2;
	wire w_dff_A_pVUEcUwf2_2;
	wire w_dff_A_YrOEY4DL7_2;
	wire w_dff_A_U60A0pOU2_1;
	wire w_dff_A_ePAM0KZN2_1;
	wire w_dff_A_TbNVKSXl8_1;
	wire w_dff_A_czh8Ldbd9_1;
	wire w_dff_A_giM0K1t94_1;
	wire w_dff_A_RFGR9Min8_1;
	wire w_dff_A_uQhfEnFK9_1;
	wire w_dff_A_LPO3o2Em8_1;
	wire w_dff_A_4Kcgv1au1_1;
	wire w_dff_A_FcxtTaGY8_1;
	wire w_dff_A_PWutiuU86_1;
	wire w_dff_A_CHXxb75R2_2;
	wire w_dff_A_lhKde5el0_2;
	wire w_dff_A_fqSfXrmM9_2;
	wire w_dff_A_edZWuZD80_2;
	wire w_dff_A_0fzo63Xs3_2;
	wire w_dff_A_eDqHULD71_2;
	wire w_dff_A_zlirVD4t1_2;
	wire w_dff_A_hyaNnRaW1_2;
	wire w_dff_A_FKlsEDyB0_2;
	wire w_dff_A_AL1UiXwR6_2;
	wire w_dff_A_qzXADXbr4_1;
	wire w_dff_A_URGcx6v34_2;
	wire w_dff_B_fqWouHea6_0;
	wire w_dff_B_vBojNKb56_0;
	wire w_dff_B_WM1tHPGa7_0;
	wire w_dff_B_FaABieyl2_0;
	wire w_dff_B_u7LXajn30_0;
	wire w_dff_B_bbJzPE2w9_0;
	wire w_dff_B_UzxBI4C67_0;
	wire w_dff_B_agNzetIO5_0;
	wire w_dff_B_Tnf8RmDr2_0;
	wire w_dff_B_f8Xw0BPk7_0;
	wire w_dff_B_7l4zDyOq7_0;
	wire w_dff_B_c0kWm8PA4_0;
	wire w_dff_B_j1RoE3pl4_1;
	wire w_dff_B_OYLwbySd3_2;
	wire w_dff_B_IijeVrdw9_2;
	wire w_dff_B_yuVHT2KF9_2;
	wire w_dff_B_mfru56XC0_1;
	wire w_dff_B_rtdV5vk31_1;
	wire w_dff_B_5UTeVcWU8_1;
	wire w_dff_B_jHTfRm792_1;
	wire w_dff_B_sVg7GnU89_1;
	wire w_dff_B_fOBGt4Bz8_1;
	wire w_dff_B_ORhifE5o6_1;
	wire w_dff_B_0Aa7H1r13_1;
	wire w_dff_B_Z5BzX2Ir7_1;
	wire w_dff_B_So66SSTL9_1;
	wire w_dff_B_fOlDPyLf2_1;
	wire w_dff_B_jFTjUPkQ1_0;
	wire w_dff_B_t7aTVRiG7_0;
	wire w_dff_B_PUgWhadD3_0;
	wire w_dff_B_Qu0lJpbU3_0;
	wire w_dff_B_xGlEeWWG5_0;
	wire w_dff_B_ZnOInu1j7_0;
	wire w_dff_B_5lYKl7oa9_0;
	wire w_dff_B_hpEDnRyu5_0;
	wire w_dff_B_vcfHocrm7_0;
	wire w_dff_B_PpfcEzsH6_0;
	wire w_dff_B_YbeTSPWj2_0;
	wire w_dff_A_rCYBnmEg1_1;
	wire w_dff_A_lP26CVsM0_1;
	wire w_dff_A_AhLdy75s1_1;
	wire w_dff_A_MTiQNhBQ7_1;
	wire w_dff_A_Pmj0bQon5_1;
	wire w_dff_A_VDZLaOd94_1;
	wire w_dff_A_2ABTlY0k5_1;
	wire w_dff_A_SPpikRhb5_1;
	wire w_dff_A_FHEEx5ER8_1;
	wire w_dff_A_t8CA8yz12_1;
	wire w_dff_A_6nFD0VXw5_1;
	wire w_dff_A_DtNh0NaG6_1;
	wire w_dff_B_IaVweoaI3_1;
	wire w_dff_B_h1XvESGJ0_1;
	wire w_dff_B_Zd4hGI9Q4_1;
	wire w_dff_A_D7xd73bS1_1;
	wire w_dff_B_ydJ6yyv97_1;
	wire w_dff_B_6MrwQT9Q8_1;
	wire w_dff_B_QzR7Lzsn5_1;
	wire w_dff_B_3a1Rd7XP1_1;
	wire w_dff_B_ulOgNjix6_1;
	wire w_dff_B_F6BENzHa7_0;
	wire w_dff_A_pKuIPQC85_1;
	wire w_dff_A_OosqPwxe4_1;
	wire w_dff_B_d48WTmlE2_1;
	wire w_dff_B_PoG6LbAh5_1;
	wire w_dff_B_kcnU5YOQ8_1;
	wire w_dff_B_tyFSTSqR1_1;
	wire w_dff_B_n9yeWDR19_1;
	wire w_dff_B_nnw0AT4Z5_1;
	wire w_dff_B_M8LVzLZV3_1;
	wire w_dff_A_dKjpUH6t2_0;
	wire w_dff_B_kv5PswOs4_0;
	wire w_dff_A_NH7oi9Al9_1;
	wire w_dff_A_BQYkyJkX0_0;
	wire w_dff_A_M91kGm5M5_2;
	wire w_dff_A_Hr6ZOa831_1;
	wire w_dff_A_9UO06Igl5_1;
	wire w_dff_A_5tZlyRKT7_1;
	wire w_dff_A_IUNeA1Eq8_2;
	wire w_dff_B_uzq9ZczS6_3;
	wire w_dff_A_EFYaffDo5_0;
	wire w_dff_B_Zp6fleZK1_2;
	wire w_dff_B_uDLjX3Wb0_2;
	wire w_dff_A_OPaFR7er4_1;
	wire w_dff_A_hzaxWGKC6_1;
	wire w_dff_A_IeQOYRoV6_1;
	wire w_dff_A_94AJ8mIn3_1;
	wire w_dff_A_5khHNIqZ3_1;
	wire w_dff_B_t1yzHTb16_2;
	wire w_dff_A_zdmK2Fm59_1;
	wire w_dff_A_9glmY7mj1_1;
	wire w_dff_A_Hf5VxlTZ1_1;
	wire w_dff_A_Kt22aKLs3_0;
	wire w_dff_A_9KwEno5i5_0;
	wire w_dff_A_RCY82oFT2_0;
	wire w_dff_A_rgjTPVoo8_0;
	wire w_dff_A_Km3aMFaw3_0;
	wire w_dff_A_1QglDTsf6_0;
	wire w_dff_B_KpRwIewu3_2;
	wire w_dff_A_ixjBq7ey4_0;
	wire w_dff_A_0EqgIHIf3_0;
	wire w_dff_B_w1DKnOjX2_2;
	wire w_dff_B_Ocovon7m7_2;
	wire w_dff_B_BeqW3IrJ0_2;
	wire w_dff_B_O8BSADvy1_2;
	wire w_dff_B_4snys8hk0_2;
	wire w_dff_B_NI9LZYTr6_0;
	wire w_dff_B_qJMIxHQY4_1;
	wire w_dff_B_rufnpOUb5_1;
	wire w_dff_A_bmnWK5Td5_1;
	wire w_dff_A_u4jsXSRD5_2;
	wire w_dff_B_i8UCO9ug3_3;
	wire w_dff_B_dnF49iJf3_3;
	wire w_dff_A_CDRu5jLO8_0;
	wire w_dff_A_9amyVOl78_0;
	wire w_dff_A_GUVM0xNJ5_0;
	wire w_dff_A_0ufqH2QY2_0;
	wire w_dff_B_PnB00RFh4_1;
	wire w_dff_B_cSHY93X78_2;
	wire w_dff_B_kFnoWgK29_2;
	wire w_dff_A_K7OHIxSs5_0;
	wire w_dff_A_UNWT6EtT7_0;
	wire w_dff_A_coU1vn0C6_0;
	wire w_dff_A_etJHdBC44_0;
	wire w_dff_A_v1RVEhNo4_2;
	wire w_dff_A_BoGRGPrV2_2;
	wire w_dff_A_G3Y4nvfc4_2;
	wire w_dff_A_EfhrMbP10_2;
	wire w_dff_A_EvXNODuB0_2;
	wire w_dff_B_QqwOgu0G4_0;
	wire w_dff_B_78eIDvzX2_1;
	wire w_dff_A_mKm665x34_0;
	wire w_dff_A_Jr12Bcpi8_0;
	wire w_dff_A_LPSyP4Pt9_0;
	wire w_dff_A_AmHetrVC6_0;
	wire w_dff_A_XFlxTCG45_0;
	wire w_dff_A_4xVxefcF9_0;
	wire w_dff_B_2JsLxuzT3_0;
	wire w_dff_B_qtjpYBK03_1;
	wire w_dff_A_wcmYu4qH4_2;
	wire w_dff_A_QSWmYASL9_2;
	wire w_dff_A_cXeHmrsK1_2;
	wire w_dff_A_N2Dbv83U3_2;
	wire w_dff_B_PtTfgjsn3_1;
	wire w_dff_B_L47W1YaZ0_1;
	wire w_dff_B_AUXkLHfA1_1;
	wire w_dff_A_1ROaP6aB5_1;
	wire w_dff_A_Nx4u9VHS9_1;
	wire w_dff_B_N09eC2bC1_0;
	wire w_dff_A_MyLlQ7YH5_0;
	wire w_dff_A_d1F1DZWd3_0;
	wire w_dff_A_DUWzhjT65_1;
	wire w_dff_A_EW7Myzab6_1;
	wire w_dff_A_HsDMthT51_1;
	wire w_dff_B_eHBdsIik4_0;
	wire w_dff_A_JgTALPGG5_0;
	wire w_dff_B_IY0qRKJx2_0;
	wire w_dff_A_hwNTQuYx7_0;
	wire w_dff_A_63dm3p8a8_0;
	wire w_dff_A_tfA75Vlz0_0;
	wire w_dff_A_TXkRm9yv3_0;
	wire w_dff_A_MYJX4VXo0_0;
	wire w_dff_A_lwdxxGTz4_0;
	wire w_dff_A_STo9Voqn1_0;
	wire w_dff_A_2jpO3pqG4_2;
	wire w_dff_A_45eAnUZd1_2;
	wire w_dff_A_kUPfPcNI0_2;
	wire w_dff_A_YbhPx2op1_2;
	wire w_dff_A_WmAB5ocj6_2;
	wire w_dff_A_AAsaCbbk5_2;
	wire w_dff_B_apOsHt3m3_1;
	wire w_dff_B_uC2qMyA97_1;
	wire w_dff_B_ahL5F1aQ9_1;
	wire w_dff_B_TEmQKGRc4_1;
	wire w_dff_B_1ge2BBjr5_1;
	wire w_dff_A_cs8aPMXM3_0;
	wire w_dff_A_HGohNdA72_0;
	wire w_dff_A_ry2AKRK42_1;
	wire w_dff_A_DrPWSbRu9_1;
	wire w_dff_A_y2ad8xAP5_1;
	wire w_dff_A_vPdbNkDr1_0;
	wire w_dff_A_MLsveOjQ4_1;
	wire w_dff_A_qauZ8gI89_1;
	wire w_dff_A_2YaYhArt2_2;
	wire w_dff_A_mQjqQizc4_0;
	wire w_dff_A_C1ZAZGdu3_0;
	wire w_dff_A_Qh9JfHui7_0;
	wire w_dff_A_SQnpHEaN0_2;
	wire w_dff_A_GJhqp7rA4_0;
	wire w_dff_A_BNmdF2OE6_0;
	wire w_dff_B_qSdA76el8_1;
	wire w_dff_B_bBt0olEp2_1;
	wire w_dff_A_XLxZLxTv8_0;
	wire w_dff_A_GdXNJ0p72_2;
	wire w_dff_A_ad3WK7eX1_1;
	wire w_dff_A_xq5uLGyz1_0;
	wire w_dff_A_eQP8c7Jd2_0;
	wire w_dff_A_o4GHBTC55_0;
	wire w_dff_B_ERBCSkDC7_1;
	wire w_dff_A_XdoSacvi2_1;
	wire w_dff_A_fCXREFVt6_1;
	wire w_dff_A_RZM6XJEj9_1;
	wire w_dff_A_QxuUtuVM6_1;
	wire w_dff_A_DbdoA8zo3_1;
	wire w_dff_A_0fg3PRYx0_1;
	wire w_dff_A_vPlwieRL3_1;
	wire w_dff_A_mFCRSRPz5_1;
	wire w_dff_A_pwgMBxzc3_1;
	wire w_dff_A_rNNYK3CC2_1;
	wire w_dff_A_GsGWKxYK5_1;
	wire w_dff_A_B3StbEzu5_2;
	wire w_dff_A_hAVoL98k3_2;
	wire w_dff_A_wLE58KEQ9_2;
	wire w_dff_A_qB8LxgmY1_2;
	wire w_dff_A_AJ0pjxUi0_2;
	wire w_dff_A_If7em4U27_2;
	wire w_dff_A_EMgxuTUe0_2;
	wire w_dff_A_thHBqV6D1_2;
	wire w_dff_A_qJ8L9seo0_0;
	wire w_dff_A_6wIWtBnV1_0;
	wire w_dff_B_Q4zcJ1XI4_1;
	wire w_dff_B_5NGtMF6T2_0;
	wire w_dff_A_CDFLFID79_1;
	wire w_dff_A_kUrqyGKP4_0;
	wire w_dff_A_Lwvf9oX12_0;
	wire w_dff_A_pBdrQaSq8_0;
	wire w_dff_A_FnOpcfzC2_0;
	wire w_dff_A_yCbNsVp33_1;
	wire w_dff_A_iPQ35uet1_1;
	wire w_dff_A_2TZ0HTV80_1;
	wire w_dff_A_6NnNjB6v3_2;
	wire w_dff_A_fbYWB9YI0_2;
	wire w_dff_A_RNhbJnaP4_2;
	wire w_dff_A_QtjbEeNI5_2;
	wire w_dff_A_na05WsST4_1;
	wire w_dff_A_0MXc5Cex0_1;
	wire w_dff_B_MWMKD1DM0_1;
	wire w_dff_B_mWIbgAuX5_1;
	wire w_dff_A_gxRtB9es3_0;
	wire w_dff_A_cLtBuRqT4_2;
	wire w_dff_A_GcIbqoCF5_0;
	wire w_dff_A_h3pchY909_0;
	wire w_dff_A_sd7fZ1847_1;
	wire w_dff_B_aVuxNvvi6_1;
	wire w_dff_A_5PM0iRLc9_1;
	wire w_dff_A_gVDVdBJY9_1;
	wire w_dff_A_2mwCsm4j6_2;
	wire w_dff_A_NIGnlWba9_2;
	wire w_dff_A_OGSlSAjg7_0;
	wire w_dff_A_AnvJjx9h2_2;
	wire w_dff_A_TQfhw9Mw6_1;
	wire w_dff_A_K6TAvHT69_2;
	wire w_dff_A_MLS9kANA5_2;
	wire w_dff_A_kj64doxa1_1;
	wire w_dff_B_0n2IaQjd2_1;
	wire w_dff_B_BboVEPTk3_1;
	wire w_dff_B_MHBdHR0n1_0;
	wire w_dff_A_3hOdmrop4_0;
	wire w_dff_A_DyUcskyR5_0;
	wire w_dff_A_cO9Gr6OZ1_1;
	wire w_dff_A_F0OTlOFe7_1;
	wire w_dff_A_Ac2yJfaK8_1;
	wire w_dff_A_MKWq9gVH1_1;
	wire w_dff_A_P03s7JlX1_2;
	wire w_dff_A_atVKGEcb4_2;
	wire w_dff_A_0ZhmUMim8_0;
	wire w_dff_B_e1go9qx96_0;
	wire w_dff_A_oXlSBaSx5_0;
	wire w_dff_A_d5VI5gxX9_0;
	wire w_dff_A_6R23NZgw3_0;
	wire w_dff_A_gVYY9rGg0_0;
	wire w_dff_A_eEayZ6AJ4_1;
	wire w_dff_A_fMXpPf7C0_1;
	wire w_dff_A_FHY5TT1y0_2;
	wire w_dff_A_0x3qhw4g3_2;
	wire w_dff_A_bZHPyQTY7_0;
	wire w_dff_A_Jnph24Rg6_0;
	wire w_dff_A_TNwFbmIf5_1;
	wire w_dff_A_5kixj4V24_0;
	wire w_dff_A_XsN8yS8u2_2;
	wire w_dff_A_W8Mlyg2V4_1;
	wire w_dff_B_aHlrTtf12_0;
	wire w_dff_A_6dzRm1Bg9_0;
	wire w_dff_A_fDbBMFjd2_2;
	wire w_dff_A_SM2qFWos7_0;
	wire w_dff_A_cu79otYr7_1;
	wire w_dff_A_OzvjWbRM9_1;
	wire w_dff_A_KozyfIKl5_2;
	wire w_dff_A_jAj800uz2_2;
	wire w_dff_A_S7x97lQ49_1;
	wire w_dff_A_Yk7dySkI4_2;
	wire w_dff_A_TnGIPudw5_2;
	wire w_dff_A_6EVykQ313_2;
	wire w_dff_A_1ajh71Lv4_2;
	wire w_dff_A_asEazgg44_2;
	wire w_dff_A_9WMDtgRQ9_2;
	wire w_dff_A_YSMGR71D3_2;
	wire w_dff_A_MWIaVXE52_2;
	wire w_dff_A_7j0KxMEI6_0;
	wire w_dff_A_qzgnXvTw3_0;
	wire w_dff_A_SzPMDIlA3_0;
	wire w_dff_A_HgKl2ejf3_0;
	wire w_dff_A_hpWNJz8J2_2;
	wire w_dff_A_yUafKato1_2;
	wire w_dff_A_OJM2wDhK4_2;
	wire w_dff_A_8pQ9if736_2;
	wire w_dff_A_9EOsrfw04_2;
	wire w_dff_A_ACt647wx5_2;
	wire w_dff_A_pmETJqGf8_2;
	wire w_dff_A_23xNqoGD4_2;
	wire w_dff_A_qqem33b11_2;
	wire w_dff_A_WcsxV8R50_1;
	wire w_dff_A_MbGbA55Z6_1;
	wire w_dff_A_IecQwGAt9_1;
	wire w_dff_A_4w7RLAhu3_1;
	wire w_dff_A_XMJJW0tL8_1;
	wire w_dff_A_nATH1QcU2_1;
	wire w_dff_A_0abN5IuP0_1;
	wire w_dff_A_AlwHnu960_1;
	wire w_dff_A_06tVJ6yW9_1;
	wire w_dff_A_M5ypYtmO1_2;
	wire w_dff_A_iXloacdp9_2;
	wire w_dff_A_LedMmay24_2;
	wire w_dff_A_GeOtFvMz8_2;
	wire w_dff_A_XrIU7Ouo9_2;
	wire w_dff_B_a7NpkydQ0_1;
	wire w_dff_B_TYsxJWRF4_1;
	wire w_dff_B_9wK0nXUx1_1;
	wire w_dff_B_hZbVmIT35_1;
	wire w_dff_B_yrHkSmoJ3_1;
	wire w_dff_B_7Y4A6LGo2_1;
	wire w_dff_B_NghpbNt44_1;
	wire w_dff_B_TPpiuW7q6_1;
	wire w_dff_B_Lmmcwpge6_1;
	wire w_dff_B_ce0KwDZg2_1;
	wire w_dff_B_60oi5j988_1;
	wire w_dff_B_J4oyQ6Tf1_1;
	wire w_dff_B_vd96JV3q7_1;
	wire w_dff_B_r8TMHfw99_1;
	wire w_dff_B_puD2XYxx4_0;
	wire w_dff_B_EYBxdOib0_0;
	wire w_dff_B_rqj1dBHn1_0;
	wire w_dff_B_Vk5lW8kJ2_0;
	wire w_dff_B_mEW6uHnO7_0;
	wire w_dff_B_W0Xf4Z5O5_0;
	wire w_dff_B_gPz1QXqV5_0;
	wire w_dff_B_3neDW6fj7_0;
	wire w_dff_B_Nt2c5WbK8_0;
	wire w_dff_B_AenvPhnV0_0;
	wire w_dff_B_ZbWxVY6Z8_0;
	wire w_dff_B_BYbj11AS2_0;
	wire w_dff_B_uKJRfvDV7_0;
	wire w_dff_B_Oddba9KG5_0;
	wire w_dff_B_lyNzQbrW4_1;
	wire w_dff_B_fVY8S10L6_1;
	wire w_dff_B_fzbEwBZS2_1;
	wire w_dff_B_Jl7gnC2Q1_1;
	wire w_dff_B_OFt7BEtg6_1;
	wire w_dff_B_KkBBRbQw1_1;
	wire w_dff_B_ruE9ChaX7_1;
	wire w_dff_B_AcB2ERIg3_0;
	wire w_dff_B_Xe7C2mQ81_1;
	wire w_dff_B_9sqnuwhk9_1;
	wire w_dff_B_28Ijl9f45_0;
	wire w_dff_B_AiB4gh4m8_0;
	wire w_dff_B_MMoHMBXD7_0;
	wire w_dff_B_g3O8EnKR9_1;
	wire w_dff_B_PwDiaseQ0_0;
	wire w_dff_B_vmJBUhKe9_1;
	wire w_dff_B_B1P9dUjr7_1;
	wire w_dff_B_dS49bua96_1;
	wire w_dff_B_8sHUGYlX8_1;
	wire w_dff_B_rbRekOsa1_1;
	wire w_dff_B_cFzSoUsO2_1;
	wire w_dff_B_vIv3LLS91_1;
	wire w_dff_B_o40UGd8j8_1;
	wire w_dff_B_VkAZvjam5_1;
	wire w_dff_B_BMknLLvv6_1;
	wire w_dff_B_kgYAeSDA7_1;
	wire w_dff_B_903H55d30_1;
	wire w_dff_B_Glpa9uIe1_1;
	wire w_dff_B_hvNLbXMv0_1;
	wire w_dff_B_iCKgjrF94_1;
	wire w_dff_B_4PpQDkje0_1;
	wire w_dff_B_ZkE0SPhO5_0;
	wire w_dff_A_pddUHG9k4_1;
	wire w_dff_B_h7Crkwla2_2;
	wire w_dff_B_ID5YT5Fh9_2;
	wire w_dff_B_E3ZWldZh9_2;
	wire w_dff_B_WzfnIOVU6_2;
	wire w_dff_A_mVU5x45s0_0;
	wire w_dff_A_2ebXTWkX1_0;
	wire w_dff_A_50lyW5Wd4_1;
	wire w_dff_A_DmbG28e35_1;
	wire w_dff_B_vMN4xilR7_2;
	wire w_dff_B_VBxjGP5o5_0;
	wire w_dff_A_JfvCvCPd3_0;
	wire w_dff_B_OmSN4Hff7_2;
	wire w_dff_B_IJ6EX7S53_2;
	wire w_dff_B_3dRmf2ut7_2;
	wire w_dff_B_3OqlOmy05_0;
	wire w_dff_B_8pmLg6vj4_0;
	wire w_dff_B_O4SYiGmJ5_0;
	wire w_dff_B_ULwlZ6nV6_0;
	wire w_dff_A_fMprN1J51_2;
	wire w_dff_A_en7ad1Kn4_2;
	wire w_dff_A_WLOZ7s6Q0_2;
	wire w_dff_A_BuNbo8jw9_2;
	wire w_dff_A_56x25ONW9_2;
	wire w_dff_A_c6TOSdvJ3_2;
	wire w_dff_A_56NzQtJd9_2;
	wire w_dff_A_GhjW42Og9_2;
	wire w_dff_A_GZztyjC65_0;
	wire w_dff_A_o9kwGvjU0_1;
	wire w_dff_A_RgqKSrrU3_1;
	wire w_dff_A_mq9RuaIy5_1;
	wire w_dff_A_raj9x4Dl2_1;
	wire w_dff_A_9AA4jxtz7_1;
	wire w_dff_A_qTwRcuC64_1;
	wire w_dff_A_t5vzpAcD6_2;
	wire w_dff_A_XqPQdzNs6_2;
	wire w_dff_A_5hchiyYo2_2;
	wire w_dff_A_DzwLaq156_2;
	wire w_dff_A_iFfrMLOE4_2;
	wire w_dff_B_zYtFHTP31_3;
	wire w_dff_B_E3phhCox2_3;
	wire w_dff_A_zfuHo9Re4_1;
	wire w_dff_A_K4XQ6b8l3_1;
	wire w_dff_A_QuPSF2du9_0;
	wire w_dff_B_dsPbd1ZL5_1;
	wire w_dff_B_G7uNY9om7_0;
	wire w_dff_B_sWj5ZqZw4_1;
	wire w_dff_B_c7Q5rMIL4_2;
	wire w_dff_A_0QktJ4318_0;
	wire w_dff_A_X9guJ0Ki5_0;
	wire w_dff_B_IEvps7dX4_0;
	wire w_dff_B_RwvYYWHM3_1;
	wire w_dff_A_JhNsed8J2_1;
	wire w_dff_A_9po5nfMh2_1;
	wire w_dff_A_fRsPcMSn4_1;
	wire w_dff_A_kzBFYKwr1_1;
	wire w_dff_A_ElfGvmoY0_1;
	wire w_dff_A_Vrj1WP1J8_0;
	wire w_dff_B_w4lX7e4x9_1;
	wire w_dff_B_DFcrzi0Y8_1;
	wire w_dff_B_MxggyYSc5_1;
	wire w_dff_B_ZZh5tCdu9_0;
	wire w_dff_B_OHyepcNP0_0;
	wire w_dff_B_U8qwk8bP1_0;
	wire w_dff_A_MnCHQddv6_0;
	wire w_dff_A_kCz2zH7F5_0;
	wire w_dff_A_f2LfcUUq5_0;
	wire w_dff_A_jG3uHNL70_0;
	wire w_dff_A_O923MLma9_1;
	wire w_dff_A_JgZzs1jo2_0;
	wire w_dff_A_XWnsyk0Z9_0;
	wire w_dff_A_zgU2YMnZ9_0;
	wire w_dff_A_Z9CoqXJ94_0;
	wire w_dff_A_nEV5xnJU2_1;
	wire w_dff_A_khti5bYU3_1;
	wire w_dff_A_2P0wzb8F8_0;
	wire w_dff_A_LEr7TiXz9_0;
	wire w_dff_A_7oiQ3gwa3_0;
	wire w_dff_A_qaAvJrj08_0;
	wire w_dff_A_vgJ2DXI13_0;
	wire w_dff_A_Zf7vTtPH2_0;
	wire w_dff_A_9ov1B3Sl8_0;
	wire w_dff_A_kdJh28BH4_0;
	wire w_dff_A_8BUd6CkQ8_2;
	wire w_dff_A_jlzzTimf3_2;
	wire w_dff_A_eH6lPn1M8_2;
	wire w_dff_A_VnWqJ54o4_2;
	wire w_dff_A_02evRjqD3_2;
	wire w_dff_A_h8mlJ5ry7_2;
	wire w_dff_A_G5zBqwwm1_2;
	wire w_dff_B_1EgBCTye7_0;
	wire w_dff_B_cLKal65A0_1;
	wire w_dff_A_dhh6kTWW6_1;
	wire w_dff_A_xtYlC6vM0_1;
	wire w_dff_A_yUFvQGBe4_1;
	wire w_dff_A_kiTgCdMK9_0;
	wire w_dff_A_ns7p0HW69_1;
	wire w_dff_A_tub42awF6_1;
	wire w_dff_A_yPXAgVCv6_1;
	wire w_dff_A_qh2rtEy50_1;
	wire w_dff_B_Q9etFRNv5_0;
	wire w_dff_A_KhdVihu96_2;
	wire w_dff_A_jVOsbSPk5_2;
	wire w_dff_A_TzhCfWqV9_2;
	wire w_dff_A_p5UUECnV1_1;
	wire w_dff_A_ukhumN2q9_1;
	wire w_dff_A_1sgg50Vh5_0;
	wire w_dff_A_FjXNNgSc6_0;
	wire w_dff_A_u58kNjAx0_0;
	wire w_dff_A_ejRfFmEt0_1;
	wire w_dff_A_dN1kmbjE3_1;
	wire w_dff_A_aMAMcnaI2_1;
	wire w_dff_A_OWasprSn8_1;
	wire w_dff_B_e8L57UDN4_1;
	wire w_dff_B_aLPQmUoB9_1;
	wire w_dff_B_KBLk7vCb4_1;
	wire w_dff_B_JVOrBYxW0_2;
	wire w_dff_B_fNYVBgIL5_2;
	wire w_dff_B_Y6TYRwuO0_2;
	wire w_dff_B_JiSN9Gy68_2;
	wire w_dff_B_xUG6aHmB6_2;
	wire w_dff_B_vtY4jYEU8_2;
	wire w_dff_B_hPZshaVc0_2;
	wire w_dff_A_f79kWhbe5_2;
	wire w_dff_A_pWeJZXtu1_2;
	wire w_dff_A_bRfgWAj95_2;
	wire w_dff_A_Yf2qE8Lp4_2;
	wire w_dff_A_tIC1BynL9_1;
	wire w_dff_A_i76LOC2U0_1;
	wire w_dff_A_1Ub2jJXa3_1;
	wire w_dff_A_QykfMVeT2_1;
	wire w_dff_A_3ADiFjjj6_1;
	wire w_dff_A_Vqq2KzBu3_1;
	wire w_dff_B_pJf8iC144_0;
	wire w_dff_A_Osos0htW4_0;
	wire w_dff_B_tcW54GU74_1;
	wire w_dff_A_p4y39Lw87_0;
	wire w_dff_A_vLeUpb2s1_1;
	wire w_dff_A_9qwxkvpO9_1;
	wire w_dff_A_WSYdpcS13_1;
	wire w_dff_A_clTPiQcX1_1;
	wire w_dff_A_6tWZHaJc8_1;
	wire w_dff_A_KEeEvvGT0_1;
	wire w_dff_A_sk2iuow46_1;
	wire w_dff_A_c8k55u2I4_1;
	wire w_dff_A_ivFqTZDA0_1;
	wire w_dff_A_vCI94uB73_1;
	wire w_dff_A_zWJzag0i3_1;
	wire w_dff_B_FFemuDfY4_0;
	wire w_dff_B_BES1QqrZ5_1;
	wire w_dff_A_yd3URyCi7_0;
	wire w_dff_A_bjbwUG7M0_2;
	wire w_dff_B_fZBBz8PT9_0;
	wire w_dff_A_wUBAaK9o5_1;
	wire w_dff_A_IRGXz4DO5_1;
	wire w_dff_A_99mLvw3T2_1;
	wire w_dff_A_yfizk2VW9_1;
	wire w_dff_A_0tA7cmZF9_1;
	wire w_dff_A_rUUA4veq5_1;
	wire w_dff_A_3iL3Rmpg0_1;
	wire w_dff_A_sl7mnM717_1;
	wire w_dff_A_klDAUInG2_1;
	wire w_dff_A_9CJp5tTw1_1;
	wire w_dff_A_ABuFr46p9_1;
	wire w_dff_A_9MIa6QAY4_2;
	wire w_dff_A_xYW9Q1cW3_2;
	wire w_dff_A_w7fSKZSl7_2;
	wire w_dff_A_wp8DNQnT5_2;
	wire w_dff_A_Lsd8e2ir4_2;
	wire w_dff_A_vKBiK2D37_2;
	wire w_dff_A_YIaTwVTq4_2;
	wire w_dff_A_H6bIqRMJ3_2;
	wire w_dff_A_OXVi1ln21_2;
	wire w_dff_A_1YgcUGKM0_2;
	wire w_dff_A_LEkVKVBX8_2;
	wire w_dff_A_aLyJPXB60_2;
	wire w_dff_A_1WXVIlvZ0_2;
	wire w_dff_A_5aFFldOM1_2;
	wire w_dff_A_lYniwzhv0_2;
	wire w_dff_A_0WzQkEuT8_2;
	wire w_dff_A_6AbCe3U21_2;
	wire w_dff_A_yBX3zBhB4_2;
	wire w_dff_A_LQkLYlbU9_2;
	wire w_dff_B_MCAgvn5H2_2;
	wire w_dff_B_nuDczt3V7_0;
	wire w_dff_A_LAvEutKN7_0;
	wire w_dff_A_t4Wy8jsh4_2;
	wire w_dff_A_lofmVhhj3_0;
	wire w_dff_A_7sr0iuu30_0;
	wire w_dff_A_1Hs6LHY27_1;
	wire w_dff_A_Fsw5FWWf3_1;
	wire w_dff_A_oG5mlAkU3_2;
	wire w_dff_B_QpVmftZ76_1;
	wire w_dff_B_gegiqUQb2_1;
	wire w_dff_A_hd0J9uOv7_0;
	wire w_dff_A_mYCOLQWJ5_2;
	wire w_dff_A_Cds4j2RZ3_2;
	wire w_dff_B_qAzlFbbr0_1;
	wire w_dff_A_itVy6ivB7_1;
	wire w_dff_A_dVCXe1m09_0;
	wire w_dff_A_bMCTS3lh5_1;
	wire w_dff_A_uLwLcYkQ5_0;
	wire w_dff_B_c7KuWy6q2_0;
	wire w_dff_A_aX7Q3r0A3_0;
	wire w_dff_A_SIaOqvhL3_2;
	wire w_dff_A_TIbKSzWp7_0;
	wire w_dff_A_BDi6pTbm8_1;
	wire w_dff_A_6BxukAJX7_1;
	wire w_dff_A_Dkuju8IF0_2;
	wire w_dff_A_2ZmmhUZk7_2;
	wire w_dff_A_nh5h3Tpz4_0;
	wire w_dff_A_HsHNtB4R8_2;
	wire w_dff_B_bIs2Ifyb2_0;
	wire w_dff_A_Gyr6Xdi39_0;
	wire w_dff_A_rUqn3KEZ1_2;
	wire w_dff_A_ywFPaaCB1_0;
	wire w_dff_A_DU9og2s62_0;
	wire w_dff_A_IFGuyCP12_1;
	wire w_dff_A_x9Mga5Vo5_0;
	wire w_dff_A_92zf0YJc9_2;
	wire w_dff_B_qxKn9S912_1;
	wire w_dff_B_1gVAaMPB9_1;
	wire w_dff_B_4jxE2WRh1_0;
	wire w_dff_A_LRGG1Bdy9_1;
	wire w_dff_A_rQBGozHr8_1;
	wire w_dff_A_UjyjVKCa7_0;
	wire w_dff_A_t7kWPFrr4_0;
	wire w_dff_A_FTBFJaf07_0;
	wire w_dff_A_am9HuM5N3_2;
	wire w_dff_A_XdkzTyra1_2;
	wire w_dff_A_oO8qcMEs4_1;
	wire w_dff_A_dBgxT8vC6_2;
	wire w_dff_B_UWRsh97v6_1;
	wire w_dff_B_ufvP6d3X3_1;
	wire w_dff_A_kGhS7hCR3_1;
	wire w_dff_A_OYzD7mj43_0;
	wire w_dff_A_vXbNci8I3_0;
	wire w_dff_A_Rwtbp0hX3_1;
	wire w_dff_B_rPkfXDut9_1;
	wire w_dff_A_7GTAHaeJ5_1;
	wire w_dff_A_jHQrua3D1_1;
	wire w_dff_A_pyWdyymZ4_2;
	wire w_dff_A_Arb3f7to5_2;
	wire w_dff_A_aMxlNGir1_0;
	wire w_dff_B_Wl0mEALJ0_1;
	wire w_dff_B_weVoAiYu5_1;
	wire w_dff_A_5h5lW8da8_1;
	wire w_dff_A_VqUJsa6V0_0;
	wire w_dff_B_P4UFu9w18_1;
	wire w_dff_A_an3LtqQN4_1;
	wire w_dff_A_QTvnrDK57_0;
	wire w_dff_A_G3VvcAxt0_0;
	wire w_dff_A_IKwuN2PV3_2;
	wire w_dff_A_wyHVClMG1_1;
	wire w_dff_A_mssGpBpw2_2;
	wire w_dff_A_A6waiVFy5_1;
	wire w_dff_A_KqWzSVqx9_2;
	wire w_dff_A_DvF0fMCl5_0;
	wire w_dff_B_BcV4qtdl5_0;
	wire w_dff_A_Hu0gcDYA1_0;
	wire w_dff_A_jgz4A8ZC0_0;
	wire w_dff_A_GOsOZ2FX8_0;
	wire w_dff_A_8flNOkE21_0;
	wire w_dff_A_JRghSMkZ4_1;
	wire w_dff_A_iKiEC3sc5_1;
	wire w_dff_A_iaeHegeY5_1;
	wire w_dff_A_bmLrmGfX2_1;
	wire w_dff_A_Tp4monOj8_1;
	wire w_dff_A_oi8BN86S2_1;
	wire w_dff_A_UaTz9xX71_2;
	wire w_dff_A_akMWDiC57_2;
	wire w_dff_A_DG9GqePC8_2;
	wire w_dff_A_kfmutEPO3_2;
	wire w_dff_A_27FkoB2q8_0;
	wire w_dff_A_qoxOJcP88_0;
	wire w_dff_A_hmdwoiRC5_1;
	wire w_dff_A_eq9gA4NK7_1;
	wire w_dff_A_uf7O1jrH4_2;
	wire w_dff_B_EYGPxgol6_0;
	wire w_dff_A_yj6NuqGK2_2;
	wire w_dff_A_ZQjdUpdm1_1;
	wire w_dff_A_2qaOPaK74_1;
	wire w_dff_A_r5cUzes00_1;
	wire w_dff_A_cXlOgeUS3_1;
	wire w_dff_A_tzs6aVif1_2;
	wire w_dff_A_ynQu8YKB0_0;
	wire w_dff_A_VdwvlNOa8_0;
	wire w_dff_A_fSkY3zGm9_0;
	wire w_dff_A_olwED41o7_0;
	wire w_dff_A_42D1ZSQZ3_1;
	wire w_dff_A_68LXjsIP1_1;
	wire w_dff_A_35cJy9Fu7_1;
	wire w_dff_A_ZF4JHgGb1_2;
	wire w_dff_A_hXTgRgpi5_2;
	wire w_dff_A_QQpdEMIz9_2;
	wire w_dff_A_bVfatrKy2_2;
	wire w_dff_A_mImFSVqW2_1;
	wire w_dff_A_GOTqrNDj2_2;
	wire w_dff_A_Qzss2TnV3_0;
	wire w_dff_A_B2BOyBS42_2;
	wire w_dff_A_h6Bje0u85_0;
	wire w_dff_A_8dtHPSLt3_0;
	wire w_dff_A_0IBeB7vB8_0;
	wire w_dff_A_menPV4hY9_0;
	wire w_dff_A_qoCehplD0_0;
	wire w_dff_A_yJIV1UTL6_0;
	wire w_dff_A_DCktl07W6_0;
	wire w_dff_A_PqJjzx568_0;
	wire w_dff_A_Tka5TvuH0_0;
	wire w_dff_A_rRft9HIC6_1;
	wire w_dff_A_jrDNxaWR0_0;
	wire w_dff_A_pWVrn1Ru0_0;
	wire w_dff_A_SqyQK0Um1_0;
	wire w_dff_A_YaQijCGJ1_0;
	wire w_dff_A_xhZzeUGE6_0;
	wire w_dff_A_C7kY2QMG8_0;
	wire w_dff_A_GTWccmwW1_2;
	wire w_dff_A_SRr5tQVE7_2;
	wire w_dff_A_KzBGOplm6_2;
	wire w_dff_A_XEBab9VM6_2;
	wire w_dff_A_ZPP8Z6Ok2_2;
	wire w_dff_A_wOz1qlpK5_2;
	wire w_dff_A_68Ycn3WV1_2;
	wire w_dff_A_oekBM2LI9_2;
	wire w_dff_A_NMinA4VU9_2;
	wire w_dff_A_hzACrLF68_2;
	wire w_dff_A_BW1HhNof2_2;
	wire w_dff_A_2vzhdSBC8_1;
	wire w_dff_A_yOFZhdsY9_1;
	wire w_dff_A_EOOm8Zae7_1;
	wire w_dff_A_W6SOQCUV2_1;
	wire w_dff_A_8zyiSCVZ6_1;
	wire w_dff_A_73FL0xGj1_1;
	wire w_dff_A_i51OnKUc9_1;
	wire w_dff_A_roWUZvzK1_1;
	wire w_dff_A_nEMLz3Xv9_1;
	wire w_dff_A_3QYF7sbO8_1;
	wire w_dff_A_fE3PXaSr1_1;
	wire w_dff_A_lVagmxix5_2;
	wire w_dff_A_mseKgEfw7_2;
	wire w_dff_A_hyrXHCH65_2;
	wire w_dff_A_4RrNPMzp2_2;
	wire w_dff_A_Y3eirACm9_2;
	wire w_dff_A_rfJtINS35_2;
	wire w_dff_A_aNJli9L43_2;
	wire w_dff_A_15yWLHBU3_2;
	wire w_dff_A_CzxrGben0_2;
	wire w_dff_A_4Xqc6g2q8_2;
	wire w_dff_A_RoRRi9D51_1;
	wire w_dff_A_YqYBMRA82_2;
	wire w_dff_B_hAsW1QNe5_2;
	wire w_dff_B_e8lsLn8v4_2;
	wire w_dff_B_GhCQXu828_2;
	wire w_dff_B_DdSWIOmF9_2;
	wire w_dff_B_LE69BYv77_2;
	wire w_dff_B_ex6DH80C1_2;
	wire w_dff_B_yFtCufYV9_2;
	wire w_dff_B_IOQQV4z05_2;
	wire w_dff_B_HYMfqDBi5_2;
	wire w_dff_B_MfX2NhZT2_2;
	wire w_dff_B_E7iF19gs1_2;
	wire w_dff_B_Vdc2STjF8_2;
	wire w_dff_B_XJnI6Mjh4_2;
	wire w_dff_B_TIr9kou64_2;
	wire w_dff_B_O1MltaaW7_2;
	wire w_dff_B_2TonRPCs2_2;
	wire w_dff_B_Zp36ZbYQ3_2;
	wire w_dff_A_pSl7gS7l5_2;
	wire w_dff_A_7tP8I1sh3_2;
	wire w_dff_A_aRuwM3Bt5_2;
	wire w_dff_A_umpHbgv29_2;
	wire w_dff_A_SCuXrD4p4_2;
	wire w_dff_A_al0XeZAo5_2;
	wire w_dff_A_ULJw2YN13_2;
	wire w_dff_A_vJgwuPfK8_2;
	wire w_dff_A_nOoVUVcn4_2;
	wire w_dff_A_oLSzWvxp9_2;
	wire w_dff_A_9Sn4SKqe4_2;
	wire w_dff_A_IrsfRMPU8_2;
	wire w_dff_A_uOeiWLTT8_2;
	wire w_dff_A_F3DBGDKX0_2;
	wire w_dff_A_OuvWcien5_0;
	wire w_dff_A_AzByg08a7_0;
	wire w_dff_A_nu0SSnYp0_0;
	wire w_dff_A_hnC9rVHO7_0;
	wire w_dff_A_4jFUwV7r7_0;
	wire w_dff_A_TLgGqsiv1_0;
	wire w_dff_A_798Txwvh4_0;
	wire w_dff_A_nc50f9tC2_0;
	wire w_dff_A_mHr5OAWm1_0;
	wire w_dff_A_EP1eZVSK3_0;
	wire w_dff_A_jrhmiOFV1_0;
	wire w_dff_A_fhfniE1w6_0;
	wire w_dff_A_a8ZdlOSK8_0;
	wire w_dff_A_tQ26enkn1_1;
	wire w_dff_A_9mTtV3JI1_1;
	wire w_dff_A_hSn8K9yg3_1;
	wire w_dff_A_vf2EN9pX1_1;
	wire w_dff_A_S5OQd7Ct9_1;
	wire w_dff_A_USVXLc106_1;
	wire w_dff_A_ipof18BS6_1;
	wire w_dff_A_f3QZiukM0_1;
	wire w_dff_A_WjS2D61k4_1;
	jnot g0000(.din(w_G545_0[2]),.dout(G594),.clk(gclk));
	jnot g0001(.din(w_G348_0[1]),.dout(G599_fa_),.clk(gclk));
	jnot g0002(.din(G366),.dout(G600_fa_),.clk(gclk));
	jand g0003(.dina(w_G562_0[1]),.dinb(w_G552_0[1]),.dout(G601_fa_),.clk(gclk));
	jnot g0004(.din(w_G549_0[2]),.dout(G602),.clk(gclk));
	jnot g0005(.din(G338),.dout(G611_fa_),.clk(gclk));
	jnot g0006(.din(w_G358_0[1]),.dout(G612_fa_),.clk(gclk));
	jand g0007(.dina(G145),.dinb(w_G141_2[2]),.dout(G810),.clk(gclk));
	jnot g0008(.din(w_G245_0[1]),.dout(G848),.clk(gclk));
	jnot g0009(.din(w_G552_0[0]),.dout(G849),.clk(gclk));
	jnot g0010(.din(w_G562_0[0]),.dout(G850),.clk(gclk));
	jnot g0011(.din(w_G559_0[1]),.dout(G851),.clk(gclk));
	jand g0012(.dina(G373),.dinb(w_G1_2[1]),.dout(G634),.clk(gclk));
	jnot g0013(.din(w_G3173_0[1]),.dout(n314),.clk(gclk));
	jand g0014(.dina(n314),.dinb(w_dff_B_WGdD0rVS3_1),.dout(G815),.clk(gclk));
	jnot g0015(.din(G27),.dout(n316),.clk(gclk));
	jcb g0016(.dina(w_dff_B_f0LYeUl25_0),.dinb(w_n316_0[1]),.dout(G845));
	jand g0017(.dina(G556),.dinb(G386),.dout(n318),.clk(gclk));
	jnot g0018(.din(w_n318_0[1]),.dout(G847),.clk(gclk));
	jnot g0019(.din(G140),.dout(n320),.clk(gclk));
	jnot g0020(.din(G31),.dout(n321),.clk(gclk));
	jcb g0021(.dina(n321),.dinb(w_n316_0[0]),.dout(G809_fa_));
	jcb g0022(.dina(w_G809_3[1]),.dinb(n320),.dout(G656));
	jnot g0023(.din(w_G299_0[2]),.dout(G593_fa_),.clk(gclk));
	jnot g0024(.din(G86),.dout(n325),.clk(gclk));
	jnot g0025(.din(w_G2358_2[2]),.dout(n326),.clk(gclk));
	jand g0026(.dina(w_n326_2[1]),.dinb(n325),.dout(n327),.clk(gclk));
	jnot g0027(.din(G87),.dout(n328),.clk(gclk));
	jand g0028(.dina(w_G2358_2[1]),.dinb(n328),.dout(n329),.clk(gclk));
	jcb g0029(.dina(n329),.dinb(w_G809_3[0]),.dout(n330));
	jcb g0030(.dina(n330),.dinb(n327),.dout(G636));
	jnot g0031(.din(G88),.dout(n332),.clk(gclk));
	jand g0032(.dina(w_n326_2[0]),.dinb(n332),.dout(n333),.clk(gclk));
	jnot g0033(.din(G34),.dout(n334),.clk(gclk));
	jand g0034(.dina(w_G2358_2[0]),.dinb(n334),.dout(n335),.clk(gclk));
	jcb g0035(.dina(n335),.dinb(w_G809_2[2]),.dout(n336));
	jcb g0036(.dina(w_n336_0[1]),.dinb(w_n333_0[1]),.dout(G704));
	jnot g0037(.din(G83),.dout(n338),.clk(gclk));
	jcb g0038(.dina(w_G809_2[1]),.dinb(n338),.dout(G820));
	jand g0039(.dina(w_n326_1[2]),.dinb(w_dff_B_BlANR4eP3_1),.dout(n340),.clk(gclk));
	jand g0040(.dina(w_G2358_1[2]),.dinb(G25),.dout(n341),.clk(gclk));
	jcb g0041(.dina(n341),.dinb(w_G809_2[0]),.dout(n342));
	jcb g0042(.dina(w_dff_B_VJcHhuhL0_0),.dinb(n340),.dout(n343));
	jand g0043(.dina(n343),.dinb(w_G141_2[1]),.dout(G639),.clk(gclk));
	jand g0044(.dina(w_n326_1[1]),.dinb(w_dff_B_q4l2q9D84_1),.dout(n345),.clk(gclk));
	jand g0045(.dina(w_G2358_1[1]),.dinb(G81),.dout(n346),.clk(gclk));
	jcb g0046(.dina(n346),.dinb(w_G809_1[2]),.dout(n347));
	jcb g0047(.dina(w_dff_B_JCFpbHak3_0),.dinb(n345),.dout(n348));
	jand g0048(.dina(n348),.dinb(w_G141_2[0]),.dout(G673),.clk(gclk));
	jand g0049(.dina(w_n326_1[0]),.dinb(w_dff_B_WJPsYA0z2_1),.dout(n350),.clk(gclk));
	jand g0050(.dina(w_G2358_1[0]),.dinb(G23),.dout(n351),.clk(gclk));
	jcb g0051(.dina(n351),.dinb(w_G809_1[1]),.dout(n352));
	jcb g0052(.dina(w_dff_B_8ew7en6g4_0),.dinb(n350),.dout(n353));
	jand g0053(.dina(n353),.dinb(w_G141_1[2]),.dout(G707),.clk(gclk));
	jand g0054(.dina(w_n326_0[2]),.dinb(w_dff_B_nZ4R98sA0_1),.dout(n355),.clk(gclk));
	jand g0055(.dina(w_G2358_0[2]),.dinb(G80),.dout(n356),.clk(gclk));
	jcb g0056(.dina(n356),.dinb(w_G809_1[0]),.dout(n357));
	jcb g0057(.dina(w_dff_B_eOyn8kPV5_0),.dinb(n355),.dout(n358));
	jand g0058(.dina(n358),.dinb(w_G141_1[1]),.dout(G715),.clk(gclk));
	jnot g0059(.din(w_G308_1[2]),.dout(n360),.clk(gclk));
	jand g0060(.dina(w_n360_0[1]),.dinb(w_G251_4[2]),.dout(n361),.clk(gclk));
	jnot g0061(.din(w_G479_1[1]),.dout(n362),.clk(gclk));
	jand g0062(.dina(w_G308_1[1]),.dinb(w_G248_5[1]),.dout(n363),.clk(gclk));
	jcb g0063(.dina(n363),.dinb(w_n362_0[1]),.dout(n364));
	jcb g0064(.dina(w_dff_B_e1go9qx96_0),.dinb(n361),.dout(n365));
	jnot g0065(.din(w_G254_1[2]),.dout(n366),.clk(gclk));
	jand g0066(.dina(w_n360_0[0]),.dinb(w_n366_4[2]),.dout(n367),.clk(gclk));
	jnot g0067(.din(w_G242_1[2]),.dout(n368),.clk(gclk));
	jand g0068(.dina(w_G308_1[0]),.dinb(w_n368_5[1]),.dout(n369),.clk(gclk));
	jcb g0069(.dina(n369),.dinb(w_G479_1[0]),.dout(n370));
	jcb g0070(.dina(n370),.dinb(n367),.dout(n371));
	jand g0071(.dina(n371),.dinb(n365),.dout(n372),.clk(gclk));
	jnot g0072(.din(w_G316_1[2]),.dout(n373),.clk(gclk));
	jand g0073(.dina(w_n373_0[1]),.dinb(w_G251_4[1]),.dout(n374),.clk(gclk));
	jnot g0074(.din(w_G490_1[2]),.dout(n375),.clk(gclk));
	jand g0075(.dina(w_G316_1[1]),.dinb(w_G248_5[0]),.dout(n376),.clk(gclk));
	jcb g0076(.dina(n376),.dinb(n375),.dout(n377));
	jcb g0077(.dina(w_dff_B_MHBdHR0n1_0),.dinb(n374),.dout(n378));
	jand g0078(.dina(w_n373_0[0]),.dinb(w_n366_4[1]),.dout(n379),.clk(gclk));
	jand g0079(.dina(w_G316_1[0]),.dinb(w_n368_5[0]),.dout(n380),.clk(gclk));
	jcb g0080(.dina(n380),.dinb(w_G490_1[1]),.dout(n381));
	jcb g0081(.dina(n381),.dinb(n379),.dout(n382));
	jand g0082(.dina(n382),.dinb(n378),.dout(n383),.clk(gclk));
	jand g0083(.dina(w_n383_0[2]),.dinb(w_n372_0[2]),.dout(n384),.clk(gclk));
	jnot g0084(.din(w_G351_2[2]),.dout(n385),.clk(gclk));
	jnot g0085(.din(G3550),.dout(n386),.clk(gclk));
	jand g0086(.dina(w_n386_4[2]),.dinb(w_n385_1[2]),.dout(n387),.clk(gclk));
	jnot g0087(.din(w_G534_1[2]),.dout(n388),.clk(gclk));
	jnot g0088(.din(w_G3552_0[1]),.dout(n389),.clk(gclk));
	jand g0089(.dina(w_n389_4[2]),.dinb(w_G351_2[1]),.dout(n390),.clk(gclk));
	jcb g0090(.dina(n390),.dinb(w_n388_1[2]),.dout(n391));
	jcb g0091(.dina(n391),.dinb(n387),.dout(n392));
	jand g0092(.dina(w_G3548_4[2]),.dinb(w_n385_1[1]),.dout(n393),.clk(gclk));
	jand g0093(.dina(w_G3546_5[1]),.dinb(w_G351_2[0]),.dout(n394),.clk(gclk));
	jcb g0094(.dina(n394),.dinb(w_G534_1[1]),.dout(n395));
	jcb g0095(.dina(w_dff_B_F0IHH1581_0),.dinb(n393),.dout(n396));
	jand g0096(.dina(n396),.dinb(n392),.dout(n397),.clk(gclk));
	jnot g0097(.din(w_G293_0[2]),.dout(n398),.clk(gclk));
	jand g0098(.dina(w_n398_0[2]),.dinb(w_n366_4[0]),.dout(n399),.clk(gclk));
	jand g0099(.dina(w_G293_0[1]),.dinb(w_n368_4[2]),.dout(n400),.clk(gclk));
	jcb g0100(.dina(n400),.dinb(n399),.dout(n401));
	jnot g0101(.din(w_G251_4[0]),.dout(n402),.clk(gclk));
	jnot g0102(.din(w_G302_0[2]),.dout(n403),.clk(gclk));
	jand g0103(.dina(w_n403_0[1]),.dinb(w_n402_2[1]),.dout(n404),.clk(gclk));
	jnot g0104(.din(w_G248_4[2]),.dout(n405),.clk(gclk));
	jand g0105(.dina(w_G302_0[1]),.dinb(w_n405_2[1]),.dout(n406),.clk(gclk));
	jcb g0106(.dina(n406),.dinb(n404),.dout(n407));
	jnot g0107(.din(w_n407_0[1]),.dout(n408),.clk(gclk));
	jand g0108(.dina(w_n408_0[1]),.dinb(w_n401_0[2]),.dout(n409),.clk(gclk));
	jnot g0109(.din(w_G514_1[1]),.dout(n410),.clk(gclk));
	jnot g0110(.din(w_G3546_5[0]),.dout(n411),.clk(gclk));
	jand g0111(.dina(n411),.dinb(w_n410_1[1]),.dout(n412),.clk(gclk));
	jand g0112(.dina(w_G3552_0[0]),.dinb(w_G514_1[0]),.dout(n413),.clk(gclk));
	jcb g0113(.dina(w_dff_B_1BQvMScw8_0),.dinb(n412),.dout(n414));
	jnot g0114(.din(w_n414_0[1]),.dout(n415),.clk(gclk));
	jnot g0115(.din(w_G361_0[2]),.dout(n416),.clk(gclk));
	jand g0116(.dina(w_n416_0[1]),.dinb(w_n402_2[0]),.dout(n417),.clk(gclk));
	jand g0117(.dina(w_G361_0[1]),.dinb(w_n405_2[0]),.dout(n418),.clk(gclk));
	jcb g0118(.dina(n418),.dinb(n417),.dout(n419));
	jnot g0119(.din(w_n419_0[2]),.dout(n420),.clk(gclk));
	jand g0120(.dina(n420),.dinb(n415),.dout(n421),.clk(gclk));
	jand g0121(.dina(n421),.dinb(n409),.dout(n422),.clk(gclk));
	jand g0122(.dina(n422),.dinb(w_n397_0[1]),.dout(n423),.clk(gclk));
	jnot g0123(.din(w_G324_1[2]),.dout(n424),.clk(gclk));
	jand g0124(.dina(w_n386_4[1]),.dinb(w_n424_2[1]),.dout(n425),.clk(gclk));
	jnot g0125(.din(w_G503_1[2]),.dout(n426),.clk(gclk));
	jand g0126(.dina(w_n389_4[1]),.dinb(w_G324_1[1]),.dout(n427),.clk(gclk));
	jcb g0127(.dina(n427),.dinb(w_n426_0[1]),.dout(n428));
	jcb g0128(.dina(n428),.dinb(n425),.dout(n429));
	jand g0129(.dina(w_G3548_4[1]),.dinb(w_n424_2[0]),.dout(n430),.clk(gclk));
	jand g0130(.dina(w_G3546_4[2]),.dinb(w_G324_1[0]),.dout(n431),.clk(gclk));
	jcb g0131(.dina(n431),.dinb(w_G503_1[1]),.dout(n432));
	jcb g0132(.dina(w_dff_B_cRPOVfjX1_0),.dinb(n430),.dout(n433));
	jand g0133(.dina(n433),.dinb(n429),.dout(n434),.clk(gclk));
	jnot g0134(.din(w_G341_2[2]),.dout(n435),.clk(gclk));
	jand g0135(.dina(w_n386_4[0]),.dinb(w_n435_1[2]),.dout(n436),.clk(gclk));
	jnot g0136(.din(w_G523_1[1]),.dout(n437),.clk(gclk));
	jand g0137(.dina(w_n389_4[0]),.dinb(w_G341_2[1]),.dout(n438),.clk(gclk));
	jcb g0138(.dina(n438),.dinb(w_n437_1[2]),.dout(n439));
	jcb g0139(.dina(n439),.dinb(n436),.dout(n440));
	jand g0140(.dina(w_G3548_4[0]),.dinb(w_n435_1[1]),.dout(n441),.clk(gclk));
	jand g0141(.dina(w_G3546_4[1]),.dinb(w_G341_2[0]),.dout(n442),.clk(gclk));
	jcb g0142(.dina(n442),.dinb(w_G523_1[0]),.dout(n443));
	jcb g0143(.dina(w_dff_B_JsUpw6qs3_0),.dinb(n441),.dout(n444));
	jand g0144(.dina(n444),.dinb(n440),.dout(n445),.clk(gclk));
	jand g0145(.dina(w_n445_0[1]),.dinb(w_n434_0[1]),.dout(n446),.clk(gclk));
	jand g0146(.dina(w_dff_B_905voHzG3_0),.dinb(n423),.dout(n447),.clk(gclk));
	jand g0147(.dina(n447),.dinb(w_dff_B_QKD54ivv8_1),.dout(G598),.clk(gclk));
	jnot g0148(.din(w_G265_2[1]),.dout(n449),.clk(gclk));
	jand g0149(.dina(w_n386_3[2]),.dinb(w_n449_1[2]),.dout(n450),.clk(gclk));
	jnot g0150(.din(w_G400_1[1]),.dout(n451),.clk(gclk));
	jand g0151(.dina(w_n389_3[2]),.dinb(w_G265_2[0]),.dout(n452),.clk(gclk));
	jcb g0152(.dina(n452),.dinb(w_n451_1[1]),.dout(n453));
	jcb g0153(.dina(n453),.dinb(n450),.dout(n454));
	jand g0154(.dina(w_G3548_3[2]),.dinb(w_n449_1[1]),.dout(n455),.clk(gclk));
	jand g0155(.dina(w_G3546_4[0]),.dinb(w_G265_1[2]),.dout(n456),.clk(gclk));
	jcb g0156(.dina(n456),.dinb(w_G400_1[0]),.dout(n457));
	jcb g0157(.dina(w_dff_B_ADAxB4i80_0),.dinb(n455),.dout(n458));
	jand g0158(.dina(n458),.dinb(n454),.dout(n459),.clk(gclk));
	jnot g0159(.din(w_G234_2[1]),.dout(n460),.clk(gclk));
	jand g0160(.dina(w_n386_3[1]),.dinb(w_n460_1[2]),.dout(n461),.clk(gclk));
	jnot g0161(.din(w_G435_1[2]),.dout(n462),.clk(gclk));
	jand g0162(.dina(w_n389_3[1]),.dinb(w_G234_2[0]),.dout(n463),.clk(gclk));
	jcb g0163(.dina(n463),.dinb(w_n462_0[2]),.dout(n464));
	jcb g0164(.dina(n464),.dinb(n461),.dout(n465));
	jand g0165(.dina(w_G3548_3[1]),.dinb(w_n460_1[1]),.dout(n466),.clk(gclk));
	jand g0166(.dina(w_G3546_3[2]),.dinb(w_G234_1[2]),.dout(n467),.clk(gclk));
	jcb g0167(.dina(n467),.dinb(w_G435_1[1]),.dout(n468));
	jcb g0168(.dina(w_dff_B_bxr6B7Pd8_0),.dinb(n466),.dout(n469));
	jand g0169(.dina(n469),.dinb(n465),.dout(n470),.clk(gclk));
	jnot g0170(.din(w_G257_2[2]),.dout(n471),.clk(gclk));
	jand g0171(.dina(w_n386_3[0]),.dinb(w_n471_1[1]),.dout(n472),.clk(gclk));
	jnot g0172(.din(w_G389_0[2]),.dout(n473),.clk(gclk));
	jand g0173(.dina(w_n389_3[0]),.dinb(w_G257_2[1]),.dout(n474),.clk(gclk));
	jcb g0174(.dina(n474),.dinb(w_n473_1[2]),.dout(n475));
	jcb g0175(.dina(n475),.dinb(n472),.dout(n476));
	jand g0176(.dina(w_G3548_3[0]),.dinb(w_n471_1[0]),.dout(n477),.clk(gclk));
	jand g0177(.dina(w_G3546_3[1]),.dinb(w_G257_2[0]),.dout(n478),.clk(gclk));
	jcb g0178(.dina(n478),.dinb(w_G389_0[1]),.dout(n479));
	jcb g0179(.dina(w_dff_B_99e8Gtle2_0),.dinb(n477),.dout(n480));
	jand g0180(.dina(n480),.dinb(n476),.dout(n481),.clk(gclk));
	jand g0181(.dina(w_n481_0[1]),.dinb(w_n470_0[1]),.dout(n482),.clk(gclk));
	jand g0182(.dina(n482),.dinb(w_n459_0[1]),.dout(n483),.clk(gclk));
	jnot g0183(.din(w_G273_2[2]),.dout(n484),.clk(gclk));
	jand g0184(.dina(w_n386_2[2]),.dinb(w_n484_1[1]),.dout(n485),.clk(gclk));
	jnot g0185(.din(w_G411_0[2]),.dout(n486),.clk(gclk));
	jand g0186(.dina(w_n389_2[2]),.dinb(w_G273_2[1]),.dout(n487),.clk(gclk));
	jcb g0187(.dina(n487),.dinb(w_n486_1[1]),.dout(n488));
	jcb g0188(.dina(n488),.dinb(n485),.dout(n489));
	jand g0189(.dina(w_G3548_2[2]),.dinb(w_n484_1[0]),.dout(n490),.clk(gclk));
	jand g0190(.dina(w_G3546_3[0]),.dinb(w_G273_2[0]),.dout(n491),.clk(gclk));
	jcb g0191(.dina(n491),.dinb(w_G411_0[1]),.dout(n492));
	jcb g0192(.dina(w_dff_B_HTcQ0nIP8_0),.dinb(n490),.dout(n493));
	jand g0193(.dina(n493),.dinb(n489),.dout(n494),.clk(gclk));
	jnot g0194(.din(w_G281_2[1]),.dout(n495),.clk(gclk));
	jand g0195(.dina(w_n386_2[1]),.dinb(w_n495_1[2]),.dout(n496),.clk(gclk));
	jnot g0196(.din(w_G374_0[2]),.dout(n497),.clk(gclk));
	jand g0197(.dina(w_n389_2[1]),.dinb(w_G281_2[0]),.dout(n498),.clk(gclk));
	jcb g0198(.dina(n498),.dinb(w_n497_1[1]),.dout(n499));
	jcb g0199(.dina(n499),.dinb(n496),.dout(n500));
	jand g0200(.dina(w_G3548_2[1]),.dinb(w_n495_1[1]),.dout(n501),.clk(gclk));
	jand g0201(.dina(w_G3546_2[2]),.dinb(w_G281_1[2]),.dout(n502),.clk(gclk));
	jcb g0202(.dina(n502),.dinb(w_G374_0[1]),.dout(n503));
	jcb g0203(.dina(w_dff_B_1pMomV046_0),.dinb(n501),.dout(n504));
	jand g0204(.dina(n504),.dinb(n500),.dout(n505),.clk(gclk));
	jand g0205(.dina(w_n505_0[1]),.dinb(w_n494_0[1]),.dout(n506),.clk(gclk));
	jnot g0206(.din(w_G218_2[2]),.dout(n507),.clk(gclk));
	jand g0207(.dina(w_n386_2[0]),.dinb(w_n507_1[1]),.dout(n508),.clk(gclk));
	jnot g0208(.din(w_G468_1[2]),.dout(n509),.clk(gclk));
	jand g0209(.dina(w_n389_2[0]),.dinb(w_G218_2[1]),.dout(n510),.clk(gclk));
	jcb g0210(.dina(n510),.dinb(w_n509_0[1]),.dout(n511));
	jcb g0211(.dina(n511),.dinb(n508),.dout(n512));
	jand g0212(.dina(w_G3548_2[0]),.dinb(w_n507_1[0]),.dout(n513),.clk(gclk));
	jand g0213(.dina(w_G3546_2[1]),.dinb(w_G218_2[0]),.dout(n514),.clk(gclk));
	jcb g0214(.dina(n514),.dinb(w_G468_1[1]),.dout(n515));
	jcb g0215(.dina(w_dff_B_VcxDnBYM0_0),.dinb(n513),.dout(n516));
	jand g0216(.dina(n516),.dinb(n512),.dout(n517),.clk(gclk));
	jnot g0217(.din(w_G206_0[2]),.dout(n518),.clk(gclk));
	jand g0218(.dina(w_G251_3[2]),.dinb(w_n518_1[1]),.dout(n519),.clk(gclk));
	jnot g0219(.din(w_G446_1[2]),.dout(n520),.clk(gclk));
	jand g0220(.dina(w_G248_4[1]),.dinb(w_G206_0[1]),.dout(n521),.clk(gclk));
	jcb g0221(.dina(n521),.dinb(n520),.dout(n522));
	jcb g0222(.dina(w_dff_B_BcV4qtdl5_0),.dinb(n519),.dout(n523));
	jand g0223(.dina(w_n366_3[2]),.dinb(w_n518_1[0]),.dout(n524),.clk(gclk));
	jand g0224(.dina(w_n368_4[1]),.dinb(w_G206_0[0]),.dout(n525),.clk(gclk));
	jcb g0225(.dina(n525),.dinb(w_G446_1[1]),.dout(n526));
	jcb g0226(.dina(n526),.dinb(n524),.dout(n527));
	jand g0227(.dina(n527),.dinb(n523),.dout(n528),.clk(gclk));
	jand g0228(.dina(w_n528_0[2]),.dinb(w_n517_0[1]),.dout(n529),.clk(gclk));
	jnot g0229(.din(w_G226_2[2]),.dout(n530),.clk(gclk));
	jand g0230(.dina(w_n386_1[2]),.dinb(w_n530_1[1]),.dout(n531),.clk(gclk));
	jnot g0231(.din(w_G422_2[1]),.dout(n532),.clk(gclk));
	jand g0232(.dina(w_n389_1[2]),.dinb(w_G226_2[1]),.dout(n533),.clk(gclk));
	jcb g0233(.dina(n533),.dinb(w_n532_0[1]),.dout(n534));
	jcb g0234(.dina(n534),.dinb(n531),.dout(n535));
	jand g0235(.dina(w_G3548_1[2]),.dinb(w_n530_1[0]),.dout(n536),.clk(gclk));
	jand g0236(.dina(w_G3546_2[0]),.dinb(w_G226_2[0]),.dout(n537),.clk(gclk));
	jcb g0237(.dina(n537),.dinb(w_G422_2[0]),.dout(n538));
	jcb g0238(.dina(w_dff_B_SlI5zjop1_0),.dinb(n536),.dout(n539));
	jand g0239(.dina(n539),.dinb(n535),.dout(n540),.clk(gclk));
	jnot g0240(.din(w_G210_2[2]),.dout(n541),.clk(gclk));
	jand g0241(.dina(w_n386_1[1]),.dinb(w_n541_1[1]),.dout(n542),.clk(gclk));
	jnot g0242(.din(w_G457_2[1]),.dout(n543),.clk(gclk));
	jand g0243(.dina(w_n389_1[1]),.dinb(w_G210_2[1]),.dout(n544),.clk(gclk));
	jcb g0244(.dina(n544),.dinb(w_n543_0[1]),.dout(n545));
	jcb g0245(.dina(n545),.dinb(n542),.dout(n546));
	jand g0246(.dina(w_G3548_1[1]),.dinb(w_n541_1[0]),.dout(n547),.clk(gclk));
	jand g0247(.dina(w_G3546_1[2]),.dinb(w_G210_2[0]),.dout(n548),.clk(gclk));
	jcb g0248(.dina(n548),.dinb(w_G457_2[0]),.dout(n549));
	jcb g0249(.dina(w_dff_B_VQfTMgXa2_0),.dinb(n547),.dout(n550));
	jand g0250(.dina(n550),.dinb(n546),.dout(n551),.clk(gclk));
	jand g0251(.dina(w_n551_0[1]),.dinb(w_n540_0[1]),.dout(n552),.clk(gclk));
	jand g0252(.dina(n552),.dinb(n529),.dout(n553),.clk(gclk));
	jand g0253(.dina(n553),.dinb(w_dff_B_yw7XDC1h4_1),.dout(n554),.clk(gclk));
	jand g0254(.dina(n554),.dinb(w_dff_B_gU6HXDMJ4_1),.dout(G610),.clk(gclk));
	jnot g0255(.din(w_G335_4[1]),.dout(n556),.clk(gclk));
	jcb g0256(.dina(w_n556_5[1]),.dinb(w_dff_B_KBLk7vCb4_1),.dout(n557));
	jand g0257(.dina(w_n556_5[0]),.dinb(w_n460_1[0]),.dout(n558),.clk(gclk));
	jnot g0258(.din(n558),.dout(n559),.clk(gclk));
	jand g0259(.dina(n559),.dinb(w_dff_B_aLPQmUoB9_1),.dout(n560),.clk(gclk));
	jxor g0260(.dina(w_n560_1[1]),.dinb(w_G435_1[0]),.dout(n561),.clk(gclk));
	jnot g0261(.din(w_n561_0[2]),.dout(n562),.clk(gclk));
	jnot g0262(.din(G288),.dout(n563),.clk(gclk));
	jand g0263(.dina(w_G335_4[0]),.dinb(n563),.dout(n564),.clk(gclk));
	jand g0264(.dina(w_n556_4[2]),.dinb(w_n495_1[0]),.dout(n565),.clk(gclk));
	jcb g0265(.dina(n565),.dinb(n564),.dout(n566));
	jxor g0266(.dina(w_n566_0[2]),.dinb(w_n497_1[0]),.dout(n567),.clk(gclk));
	jcb g0267(.dina(w_n556_4[1]),.dinb(w_G280_0[1]),.dout(n568));
	jcb g0268(.dina(w_G335_3[2]),.dinb(w_G273_1[2]),.dout(n569));
	jand g0269(.dina(w_n569_0[1]),.dinb(n568),.dout(n570),.clk(gclk));
	jxor g0270(.dina(w_n570_0[1]),.dinb(w_n486_1[0]),.dout(n571),.clk(gclk));
	jnot g0271(.din(w_n571_1[1]),.dout(n572),.clk(gclk));
	jand g0272(.dina(w_n572_0[2]),.dinb(w_n567_1[1]),.dout(n573),.clk(gclk));
	jnot g0273(.din(n573),.dout(n574),.clk(gclk));
	jcb g0274(.dina(w_n556_4[0]),.dinb(w_dff_B_tcW54GU74_1),.dout(n575));
	jcb g0275(.dina(w_G335_3[1]),.dinb(w_G257_1[2]),.dout(n576));
	jand g0276(.dina(w_dff_B_pJf8iC144_0),.dinb(n575),.dout(n577),.clk(gclk));
	jxor g0277(.dina(w_n577_0[2]),.dinb(w_n473_1[1]),.dout(n578),.clk(gclk));
	jnot g0278(.din(G272),.dout(n579),.clk(gclk));
	jand g0279(.dina(w_G335_3[0]),.dinb(n579),.dout(n580),.clk(gclk));
	jand g0280(.dina(w_n556_3[2]),.dinb(w_n449_1[0]),.dout(n581),.clk(gclk));
	jcb g0281(.dina(n581),.dinb(n580),.dout(n582));
	jxor g0282(.dina(w_n582_1[1]),.dinb(w_G400_0[2]),.dout(n583),.clk(gclk));
	jcb g0283(.dina(w_n583_1[1]),.dinb(w_n578_0[2]),.dout(n584));
	jcb g0284(.dina(w_dff_B_U8qwk8bP1_0),.dinb(w_n574_0[2]),.dout(n585));
	jcb g0285(.dina(w_n585_0[1]),.dinb(w_n562_0[1]),.dout(n586));
	jnot g0286(.din(n586),.dout(n587),.clk(gclk));
	jcb g0287(.dina(w_n556_3[1]),.dinb(w_dff_B_BES1QqrZ5_1),.dout(n588));
	jcb g0288(.dina(w_G335_2[2]),.dinb(w_G210_1[2]),.dout(n589));
	jand g0289(.dina(w_dff_B_FFemuDfY4_0),.dinb(n588),.dout(n590),.clk(gclk));
	jxor g0290(.dina(w_n590_1[1]),.dinb(w_G457_1[2]),.dout(n591),.clk(gclk));
	jcb g0291(.dina(w_n556_3[0]),.dinb(w_dff_B_MxggyYSc5_1),.dout(n592));
	jand g0292(.dina(w_n556_2[2]),.dinb(w_n518_0[2]),.dout(n593),.clk(gclk));
	jnot g0293(.din(n593),.dout(n594),.clk(gclk));
	jand g0294(.dina(n594),.dinb(w_dff_B_DFcrzi0Y8_1),.dout(n595),.clk(gclk));
	jxor g0295(.dina(w_n595_1[1]),.dinb(w_G446_1[0]),.dout(n596),.clk(gclk));
	jand g0296(.dina(w_n596_0[2]),.dinb(w_n591_0[1]),.dout(n597),.clk(gclk));
	jcb g0297(.dina(w_n556_2[1]),.dinb(w_dff_B_sWj5ZqZw4_1),.dout(n598));
	jcb g0298(.dina(w_G335_2[1]),.dinb(w_G226_1[2]),.dout(n599));
	jand g0299(.dina(w_dff_B_G7uNY9om7_0),.dinb(n598),.dout(n600),.clk(gclk));
	jxor g0300(.dina(w_n600_1[1]),.dinb(w_G422_1[2]),.dout(n601),.clk(gclk));
	jcb g0301(.dina(w_n556_2[0]),.dinb(w_dff_B_RwvYYWHM3_1),.dout(n602));
	jcb g0302(.dina(w_G335_2[0]),.dinb(w_G218_1[2]),.dout(n603));
	jand g0303(.dina(w_dff_B_IEvps7dX4_0),.dinb(n602),.dout(n604),.clk(gclk));
	jxor g0304(.dina(w_n604_0[2]),.dinb(w_G468_1[0]),.dout(n605),.clk(gclk));
	jand g0305(.dina(w_n605_2[2]),.dinb(w_n601_0[1]),.dout(n606),.clk(gclk));
	jand g0306(.dina(w_dff_B_W1C3vtJh6_0),.dinb(n597),.dout(n607),.clk(gclk));
	jand g0307(.dina(w_n607_0[2]),.dinb(w_n587_1[1]),.dout(G588),.clk(gclk));
	jnot g0308(.din(w_G332_4[2]),.dout(n609),.clk(gclk));
	jcb g0309(.dina(w_n609_5[2]),.dinb(w_G331_0[1]),.dout(n610));
	jand g0310(.dina(w_n609_5[1]),.dinb(w_n424_1[2]),.dout(n611),.clk(gclk));
	jnot g0311(.din(n611),.dout(n612),.clk(gclk));
	jand g0312(.dina(n612),.dinb(w_dff_B_bBt0olEp2_1),.dout(n613),.clk(gclk));
	jxor g0313(.dina(w_n613_0[2]),.dinb(w_G503_1[0]),.dout(n614),.clk(gclk));
	jcb g0314(.dina(w_G358_0[0]),.dinb(w_n609_5[0]),.dout(n615));
	jcb g0315(.dina(w_G351_1[2]),.dinb(w_G332_4[1]),.dout(n616));
	jand g0316(.dina(w_dff_B_IY0qRKJx2_0),.dinb(n615),.dout(n617),.clk(gclk));
	jxor g0317(.dina(w_n617_1[1]),.dinb(w_n388_1[1]),.dout(n618),.clk(gclk));
	jand g0318(.dina(w_G600_0),.dinb(w_G332_4[0]),.dout(n619),.clk(gclk));
	jand g0319(.dina(w_n416_0[0]),.dinb(w_n609_4[2]),.dout(n620),.clk(gclk));
	jcb g0320(.dina(n620),.dinb(n619),.dout(n621));
	jnot g0321(.din(w_n621_2[1]),.dout(n622),.clk(gclk));
	jcb g0322(.dina(w_n622_1[1]),.dinb(w_n618_1[1]),.dout(n623));
	jand g0323(.dina(w_G611_0),.dinb(w_G332_3[2]),.dout(n624),.clk(gclk));
	jxor g0324(.dina(w_n624_1[2]),.dinb(w_G514_0[2]),.dout(n625),.clk(gclk));
	jcb g0325(.dina(w_G348_0[0]),.dinb(w_n609_4[1]),.dout(n626));
	jcb g0326(.dina(w_G341_1[2]),.dinb(w_G332_3[1]),.dout(n627));
	jand g0327(.dina(w_dff_B_eHBdsIik4_0),.dinb(n626),.dout(n628),.clk(gclk));
	jxor g0328(.dina(w_n628_0[2]),.dinb(w_n437_1[1]),.dout(n629),.clk(gclk));
	jcb g0329(.dina(w_n629_0[2]),.dinb(w_n625_0[2]),.dout(n630));
	jcb g0330(.dina(n630),.dinb(w_n623_0[1]),.dout(n631));
	jnot g0331(.din(w_n631_0[1]),.dout(n632),.clk(gclk));
	jand g0332(.dina(w_dff_B_N09eC2bC1_0),.dinb(w_n614_2[1]),.dout(n633),.clk(gclk));
	jand g0333(.dina(w_G332_3[0]),.dinb(w_G593_0),.dout(n634),.clk(gclk));
	jand g0334(.dina(w_n609_4[0]),.dinb(w_n398_0[1]),.dout(n635),.clk(gclk));
	jcb g0335(.dina(n635),.dinb(n634),.dout(n636));
	jcb g0336(.dina(w_n609_3[2]),.dinb(w_dff_B_AUXkLHfA1_1),.dout(n637));
	jand g0337(.dina(w_n609_3[1]),.dinb(w_n403_0[0]),.dout(n638),.clk(gclk));
	jnot g0338(.din(n638),.dout(n639),.clk(gclk));
	jand g0339(.dina(n639),.dinb(w_dff_B_L47W1YaZ0_1),.dout(n640),.clk(gclk));
	jnot g0340(.din(w_n640_1[2]),.dout(n641),.clk(gclk));
	jand g0341(.dina(w_n641_0[1]),.dinb(w_n636_1[1]),.dout(n642),.clk(gclk));
	jcb g0342(.dina(w_n609_3[0]),.dinb(w_dff_B_qtjpYBK03_1),.dout(n643));
	jcb g0343(.dina(w_G332_2[2]),.dinb(w_G308_0[2]),.dout(n644));
	jand g0344(.dina(w_dff_B_2JsLxuzT3_0),.dinb(n643),.dout(n645),.clk(gclk));
	jxor g0345(.dina(w_n645_0[2]),.dinb(w_G479_0[2]),.dout(n646),.clk(gclk));
	jcb g0346(.dina(w_n609_2[2]),.dinb(w_dff_B_78eIDvzX2_1),.dout(n647));
	jcb g0347(.dina(w_G332_2[1]),.dinb(w_G316_0[2]),.dout(n648));
	jand g0348(.dina(w_dff_B_QqwOgu0G4_0),.dinb(n647),.dout(n649),.clk(gclk));
	jxor g0349(.dina(w_n649_1[1]),.dinb(w_G490_1[0]),.dout(n650),.clk(gclk));
	jand g0350(.dina(w_n650_0[1]),.dinb(w_n646_0[2]),.dout(n651),.clk(gclk));
	jand g0351(.dina(w_n651_1[1]),.dinb(w_n642_0[1]),.dout(n652),.clk(gclk));
	jand g0352(.dina(w_n652_0[1]),.dinb(w_n633_1[1]),.dout(G615),.clk(gclk));
	jxor g0353(.dina(w_G316_0[1]),.dinb(w_G308_0[1]),.dout(n654),.clk(gclk));
	jxor g0354(.dina(w_G351_1[1]),.dinb(w_G341_1[1]),.dout(n655),.clk(gclk));
	jxor g0355(.dina(n655),.dinb(n654),.dout(n656),.clk(gclk));
	jxor g0356(.dina(w_G369_0[1]),.dinb(w_G361_0[0]),.dout(n657),.clk(gclk));
	jxor g0357(.dina(n657),.dinb(w_n424_1[1]),.dout(n658),.clk(gclk));
	jxor g0358(.dina(w_G302_0[0]),.dinb(w_n398_0[0]),.dout(n659),.clk(gclk));
	jxor g0359(.dina(n659),.dinb(n658),.dout(n660),.clk(gclk));
	jxor g0360(.dina(n660),.dinb(w_dff_B_1wrzx3hs6_1),.dout(n661),.clk(gclk));
	jnot g0361(.din(w_n661_0[1]),.dout(G1002),.clk(gclk));
	jxor g0362(.dina(w_G226_1[1]),.dinb(w_G218_1[1]),.dout(n663),.clk(gclk));
	jxor g0363(.dina(w_G273_1[1]),.dinb(w_G265_1[1]),.dout(n664),.clk(gclk));
	jxor g0364(.dina(n664),.dinb(n663),.dout(n665),.clk(gclk));
	jxor g0365(.dina(w_G289_0[1]),.dinb(w_G281_1[1]),.dout(n666),.clk(gclk));
	jxor g0366(.dina(w_G257_1[1]),.dinb(w_G234_1[1]),.dout(n667),.clk(gclk));
	jxor g0367(.dina(n667),.dinb(n666),.dout(n668),.clk(gclk));
	jxor g0368(.dina(w_G210_1[1]),.dinb(w_n518_0[1]),.dout(n669),.clk(gclk));
	jxor g0369(.dina(n669),.dinb(n668),.dout(n670),.clk(gclk));
	jxor g0370(.dina(n670),.dinb(w_dff_B_PK1nw0l90_1),.dout(n671),.clk(gclk));
	jnot g0371(.din(w_n671_0[1]),.dout(G1004),.clk(gclk));
	jnot g0372(.din(w_n560_1[0]),.dout(n673),.clk(gclk));
	jand g0373(.dina(n673),.dinb(w_n462_0[1]),.dout(n674),.clk(gclk));
	jnot g0374(.din(n674),.dout(n675),.clk(gclk));
	jand g0375(.dina(w_n560_0[2]),.dinb(w_G435_0[2]),.dout(n676),.clk(gclk));
	jnot g0376(.din(w_n577_0[1]),.dout(n677),.clk(gclk));
	jand g0377(.dina(w_n677_0[1]),.dinb(w_n473_1[0]),.dout(n678),.clk(gclk));
	jcb g0378(.dina(w_n677_0[0]),.dinb(w_n473_0[2]),.dout(n679));
	jand g0379(.dina(w_n582_1[0]),.dinb(w_n451_1[0]),.dout(n680),.clk(gclk));
	jcb g0380(.dina(w_n566_0[1]),.dinb(w_n497_0[2]),.dout(n681));
	jcb g0381(.dina(w_n571_1[0]),.dinb(w_n681_2[1]),.dout(n682));
	jnot g0382(.din(w_G280_0[0]),.dout(n683),.clk(gclk));
	jand g0383(.dina(w_G335_1[2]),.dinb(n683),.dout(n684),.clk(gclk));
	jnot g0384(.din(w_n569_0[0]),.dout(n685),.clk(gclk));
	jcb g0385(.dina(w_dff_B_Q9etFRNv5_0),.dinb(n684),.dout(n686));
	jcb g0386(.dina(n686),.dinb(w_n486_0[2]),.dout(n687));
	jcb g0387(.dina(w_n582_0[2]),.dinb(w_n451_0[2]),.dout(n688));
	jand g0388(.dina(n688),.dinb(w_n687_0[2]),.dout(n689),.clk(gclk));
	jand g0389(.dina(w_n689_0[1]),.dinb(w_n682_0[1]),.dout(n690),.clk(gclk));
	jcb g0390(.dina(n690),.dinb(w_n680_0[1]),.dout(n691));
	jand g0391(.dina(w_n691_0[2]),.dinb(w_n679_0[1]),.dout(n692),.clk(gclk));
	jcb g0392(.dina(n692),.dinb(w_n678_0[1]),.dout(n693));
	jnot g0393(.din(w_n693_0[2]),.dout(n694),.clk(gclk));
	jcb g0394(.dina(n694),.dinb(w_dff_B_cLKal65A0_1),.dout(n695));
	jand g0395(.dina(w_dff_B_1EgBCTye7_0),.dinb(n675),.dout(n696),.clk(gclk));
	jand g0396(.dina(w_n696_0[2]),.dinb(w_n607_0[1]),.dout(n697),.clk(gclk));
	jand g0397(.dina(w_n595_1[0]),.dinb(w_G446_0[2]),.dout(n698),.clk(gclk));
	jcb g0398(.dina(w_n595_0[2]),.dinb(w_G446_0[1]),.dout(n699));
	jcb g0399(.dina(w_n590_1[0]),.dinb(w_G457_1[1]),.dout(n700));
	jand g0400(.dina(w_n590_0[2]),.dinb(w_G457_1[0]),.dout(n701),.clk(gclk));
	jand g0401(.dina(w_n604_0[1]),.dinb(w_G468_0[2]),.dout(n702),.clk(gclk));
	jand g0402(.dina(w_n600_1[0]),.dinb(w_G422_1[1]),.dout(n703),.clk(gclk));
	jand g0403(.dina(w_n605_2[1]),.dinb(w_n703_0[2]),.dout(n704),.clk(gclk));
	jcb g0404(.dina(n704),.dinb(w_n702_0[1]),.dout(n705));
	jcb g0405(.dina(w_n705_0[1]),.dinb(w_dff_B_dsPbd1ZL5_1),.dout(n706));
	jand g0406(.dina(w_n706_0[1]),.dinb(w_n700_0[1]),.dout(n707),.clk(gclk));
	jand g0407(.dina(w_n707_0[2]),.dinb(w_dff_B_F8cqQGOc6_1),.dout(n708),.clk(gclk));
	jcb g0408(.dina(n708),.dinb(w_dff_B_tml5FdyV9_1),.dout(n709));
	jcb g0409(.dina(w_n709_0[1]),.dinb(w_n697_0[1]),.dout(G591));
	jand g0410(.dina(w_n613_0[1]),.dinb(w_G503_0[2]),.dout(n711),.clk(gclk));
	jcb g0411(.dina(w_n624_1[1]),.dinb(w_n410_1[0]),.dout(n712));
	jand g0412(.dina(w_n624_1[0]),.dinb(w_n410_0[2]),.dout(n713),.clk(gclk));
	jand g0413(.dina(w_G599_0),.dinb(w_G332_2[0]),.dout(n714),.clk(gclk));
	jand g0414(.dina(w_n435_1[0]),.dinb(w_n609_2[1]),.dout(n715),.clk(gclk));
	jcb g0415(.dina(n715),.dinb(n714),.dout(n716));
	jand g0416(.dina(w_n716_0[1]),.dinb(w_n437_1[0]),.dout(n717),.clk(gclk));
	jand g0417(.dina(w_G612_0),.dinb(w_G332_1[2]),.dout(n718),.clk(gclk));
	jand g0418(.dina(w_n385_1[0]),.dinb(w_n609_2[0]),.dout(n719),.clk(gclk));
	jcb g0419(.dina(n719),.dinb(n718),.dout(n720));
	jand g0420(.dina(w_n720_0[1]),.dinb(w_n388_1[0]),.dout(n721),.clk(gclk));
	jcb g0421(.dina(w_n621_2[0]),.dinb(w_n721_0[2]),.dout(n722));
	jcb g0422(.dina(w_n720_0[0]),.dinb(w_n388_0[2]),.dout(n723));
	jcb g0423(.dina(w_n716_0[0]),.dinb(w_n437_0[2]),.dout(n724));
	jand g0424(.dina(n724),.dinb(w_n723_0[1]),.dout(n725),.clk(gclk));
	jand g0425(.dina(n725),.dinb(n722),.dout(n726),.clk(gclk));
	jcb g0426(.dina(w_n726_0[1]),.dinb(w_n717_0[2]),.dout(n727));
	jcb g0427(.dina(w_n727_0[2]),.dinb(w_dff_B_1ge2BBjr5_1),.dout(n728));
	jand g0428(.dina(n728),.dinb(w_dff_B_TEmQKGRc4_1),.dout(n729),.clk(gclk));
	jnot g0429(.din(w_n729_1[1]),.dout(n730),.clk(gclk));
	jand g0430(.dina(n730),.dinb(w_n614_2[0]),.dout(n731),.clk(gclk));
	jcb g0431(.dina(n731),.dinb(w_dff_B_uC2qMyA97_1),.dout(n732));
	jand g0432(.dina(w_n732_0[2]),.dinb(w_n651_1[0]),.dout(n733),.clk(gclk));
	jnot g0433(.din(w_n642_0[0]),.dout(n734),.clk(gclk));
	jnot g0434(.din(w_n645_0[1]),.dout(n735),.clk(gclk));
	jand g0435(.dina(w_n735_0[1]),.dinb(w_n362_0[0]),.dout(n736),.clk(gclk));
	jnot g0436(.din(w_n736_0[1]),.dout(n737),.clk(gclk));
	jand g0437(.dina(w_n645_0[0]),.dinb(w_G479_0[1]),.dout(n738),.clk(gclk));
	jand g0438(.dina(w_n649_1[0]),.dinb(w_G490_0[2]),.dout(n739),.clk(gclk));
	jcb g0439(.dina(w_n739_1[1]),.dinb(n738),.dout(n740));
	jand g0440(.dina(w_n740_0[1]),.dinb(n737),.dout(n741),.clk(gclk));
	jcb g0441(.dina(w_n741_0[1]),.dinb(n734),.dout(n742));
	jcb g0442(.dina(w_n742_0[1]),.dinb(w_n733_0[1]),.dout(G618));
	jnot g0443(.din(w_G54_0[1]),.dout(n744),.clk(gclk));
	jxor g0444(.dina(w_n621_1[2]),.dinb(w_n744_1[2]),.dout(n745),.clk(gclk));
	jnot g0445(.din(w_G4092_1[2]),.dout(n746),.clk(gclk));
	jand g0446(.dina(w_n746_1[2]),.dinb(w_G4091_2[2]),.dout(n747),.clk(gclk));
	jnot g0447(.din(w_n747_3[2]),.dout(n748),.clk(gclk));
	jcb g0448(.dina(w_n748_4[1]),.dinb(n745),.dout(n749));
	jnot g0449(.din(w_G4091_2[1]),.dout(n750),.clk(gclk));
	jand g0450(.dina(w_n746_1[1]),.dinb(w_n750_1[1]),.dout(n751),.clk(gclk));
	jand g0451(.dina(w_n751_2[1]),.dinb(w_n419_0[1]),.dout(n752),.clk(gclk));
	jand g0452(.dina(w_G4092_1[1]),.dinb(w_n750_1[0]),.dout(n753),.clk(gclk));
	jand g0453(.dina(w_n753_8[1]),.dinb(w_dff_B_26hfeWVD4_1),.dout(n754),.clk(gclk));
	jcb g0454(.dina(n754),.dinb(n752),.dout(n755));
	jnot g0455(.din(n755),.dout(n756),.clk(gclk));
	jand g0456(.dina(n756),.dinb(w_dff_B_eSJT5Mt21_1),.dout(G822_fa_),.clk(gclk));
	jnot g0457(.din(w_n618_1[0]),.dout(n758),.clk(gclk));
	jand g0458(.dina(w_n621_1[1]),.dinb(w_n744_1[1]),.dout(n759),.clk(gclk));
	jnot g0459(.din(w_n759_0[1]),.dout(n760),.clk(gclk));
	jand g0460(.dina(w_n760_0[1]),.dinb(n758),.dout(n761),.clk(gclk));
	jand g0461(.dina(w_n759_0[0]),.dinb(w_n618_0[2]),.dout(n762),.clk(gclk));
	jcb g0462(.dina(n762),.dinb(w_n748_4[0]),.dout(n763));
	jcb g0463(.dina(w_dff_B_ndd83xYU6_0),.dinb(w_n761_0[1]),.dout(n764));
	jnot g0464(.din(w_n751_2[0]),.dout(n765),.clk(gclk));
	jcb g0465(.dina(w_n765_5[2]),.dinb(w_n397_0[0]),.dout(n766));
	jand g0466(.dina(w_n753_8[0]),.dinb(w_dff_B_NZQc0blX1_1),.dout(n767),.clk(gclk));
	jnot g0467(.din(n767),.dout(n768),.clk(gclk));
	jand g0468(.dina(n768),.dinb(w_dff_B_2i2NURNA2_1),.dout(n769),.clk(gclk));
	jand g0469(.dina(n769),.dinb(n764),.dout(G838_fa_),.clk(gclk));
	jxor g0470(.dina(w_n567_1[0]),.dinb(w_G4_1[1]),.dout(n771),.clk(gclk));
	jand g0471(.dina(w_n771_0[1]),.dinb(w_n747_3[1]),.dout(n772),.clk(gclk));
	jnot g0472(.din(n772),.dout(n773),.clk(gclk));
	jcb g0473(.dina(w_n765_5[1]),.dinb(w_n505_0[0]),.dout(n774));
	jand g0474(.dina(w_n753_7[2]),.dinb(w_dff_B_gMgEU3kz8_1),.dout(n775),.clk(gclk));
	jnot g0475(.din(n775),.dout(n776),.clk(gclk));
	jand g0476(.dina(n776),.dinb(w_dff_B_nYzCmORx9_1),.dout(n777),.clk(gclk));
	jand g0477(.dina(w_dff_B_2OZpruAF3_0),.dinb(n773),.dout(G861_fa_),.clk(gclk));
	jnot g0478(.din(w_n636_1[0]),.dout(n779),.clk(gclk));
	jand g0479(.dina(w_n633_1[0]),.dinb(w_G54_0[0]),.dout(n780),.clk(gclk));
	jcb g0480(.dina(n780),.dinb(w_n732_0[1]),.dout(n781));
	jand g0481(.dina(w_n781_0[2]),.dinb(w_n651_0[2]),.dout(n782),.clk(gclk));
	jcb g0482(.dina(n782),.dinb(w_n741_0[0]),.dout(n783));
	jnot g0483(.din(w_n783_1[1]),.dout(n784),.clk(gclk));
	jcb g0484(.dina(n784),.dinb(w_n779_0[1]),.dout(n785));
	jxor g0485(.dina(w_n640_1[1]),.dinb(w_n779_0[0]),.dout(n786),.clk(gclk));
	jnot g0486(.din(w_n786_0[1]),.dout(n787),.clk(gclk));
	jcb g0487(.dina(w_n787_0[1]),.dinb(w_n783_1[0]),.dout(n788));
	jand g0488(.dina(w_dff_B_4bhq2NKq5_0),.dinb(n785),.dout(n789),.clk(gclk));
	jnot g0489(.din(w_n789_0[2]),.dout(G623),.clk(gclk));
	jnot g0490(.din(w_G861_0),.dout(n791),.clk(gclk));
	jnot g0491(.din(w_G4087_0[2]),.dout(n792),.clk(gclk));
	jand g0492(.dina(w_G4088_0[2]),.dinb(w_n792_0[1]),.dout(n793),.clk(gclk));
	jand g0493(.dina(w_n793_4[1]),.dinb(w_n791_1[1]),.dout(n794),.clk(gclk));
	jnot g0494(.din(w_G822_0),.dout(n795),.clk(gclk));
	jnot g0495(.din(w_G4088_0[1]),.dout(n796),.clk(gclk));
	jand g0496(.dina(w_n796_0[1]),.dinb(w_n792_0[0]),.dout(n797),.clk(gclk));
	jand g0497(.dina(w_n797_4[1]),.dinb(w_n795_1[1]),.dout(n798),.clk(gclk));
	jand g0498(.dina(w_n796_0[0]),.dinb(w_G4087_0[1]),.dout(n799),.clk(gclk));
	jand g0499(.dina(w_n799_4[1]),.dinb(w_G11_0[1]),.dout(n800),.clk(gclk));
	jand g0500(.dina(w_G4088_0[0]),.dinb(w_G4087_0[0]),.dout(n801),.clk(gclk));
	jand g0501(.dina(w_n801_4[1]),.dinb(w_G61_0[1]),.dout(n802),.clk(gclk));
	jcb g0502(.dina(w_dff_B_F722iPpp8_0),.dinb(n800),.dout(n803));
	jcb g0503(.dina(w_dff_B_TeOv1NbB9_0),.dinb(n798),.dout(n804));
	jcb g0504(.dina(w_dff_B_w4igoQQ31_0),.dinb(n794),.dout(G722));
	jand g0505(.dina(w_n729_1[0]),.dinb(w_n631_0[0]),.dout(n806),.clk(gclk));
	jand g0506(.dina(w_n729_0[2]),.dinb(w_n744_1[0]),.dout(n807),.clk(gclk));
	jcb g0507(.dina(n807),.dinb(w_n806_0[2]),.dout(n808));
	jxor g0508(.dina(n808),.dinb(w_n614_1[2]),.dout(n809),.clk(gclk));
	jcb g0509(.dina(w_n809_0[1]),.dinb(w_n748_3[2]),.dout(n810));
	jcb g0510(.dina(w_n765_5[0]),.dinb(w_n434_0[0]),.dout(n811));
	jand g0511(.dina(w_n753_7[1]),.dinb(w_dff_B_g8h89HDW9_1),.dout(n812),.clk(gclk));
	jnot g0512(.din(n812),.dout(n813),.clk(gclk));
	jand g0513(.dina(n813),.dinb(w_dff_B_mZBKS0aB4_1),.dout(n814),.clk(gclk));
	jand g0514(.dina(w_dff_B_RP8ZKKAf4_0),.dinb(n810),.dout(G832_fa_),.clk(gclk));
	jnot g0515(.din(w_n625_0[1]),.dout(n816),.clk(gclk));
	jand g0516(.dina(w_n727_0[1]),.dinb(w_n744_0[2]),.dout(n817),.clk(gclk));
	jand g0517(.dina(w_n726_0[0]),.dinb(w_n623_0[0]),.dout(n818),.clk(gclk));
	jcb g0518(.dina(n818),.dinb(w_n717_0[1]),.dout(n819));
	jcb g0519(.dina(w_n819_0[1]),.dinb(n817),.dout(n820));
	jxor g0520(.dina(n820),.dinb(w_dff_B_4emycJed9_1),.dout(n821),.clk(gclk));
	jcb g0521(.dina(w_n821_0[1]),.dinb(w_n748_3[1]),.dout(n822));
	jand g0522(.dina(w_n751_1[2]),.dinb(w_n414_0[0]),.dout(n823),.clk(gclk));
	jand g0523(.dina(w_n753_7[0]),.dinb(w_dff_B_H8s9gCkA2_1),.dout(n824),.clk(gclk));
	jcb g0524(.dina(n824),.dinb(n823),.dout(n825));
	jnot g0525(.din(n825),.dout(n826),.clk(gclk));
	jand g0526(.dina(w_dff_B_IGABrCwK7_0),.dinb(n822),.dout(G834_fa_),.clk(gclk));
	jcb g0527(.dina(w_n617_1[0]),.dinb(w_G534_1[0]),.dout(n828));
	jand g0528(.dina(w_n617_0[2]),.dinb(w_G534_0[2]),.dout(n829),.clk(gclk));
	jcb g0529(.dina(w_n760_0[0]),.dinb(w_n829_0[1]),.dout(n830));
	jand g0530(.dina(n830),.dinb(w_n828_0[2]),.dout(n831),.clk(gclk));
	jxor g0531(.dina(n831),.dinb(w_n629_0[1]),.dout(n832),.clk(gclk));
	jcb g0532(.dina(w_n832_0[1]),.dinb(w_n748_3[0]),.dout(n833));
	jcb g0533(.dina(w_n765_4[2]),.dinb(w_n445_0[0]),.dout(n834));
	jand g0534(.dina(w_n753_6[2]),.dinb(w_dff_B_UnolPSSa7_1),.dout(n835),.clk(gclk));
	jnot g0535(.din(n835),.dout(n836),.clk(gclk));
	jand g0536(.dina(n836),.dinb(w_dff_B_AIv8lL129_1),.dout(n837),.clk(gclk));
	jand g0537(.dina(w_dff_B_B4AvEkKb9_0),.dinb(n833),.dout(G836_fa_),.clk(gclk));
	jnot g0538(.din(w_G4090_0[2]),.dout(n839),.clk(gclk));
	jand g0539(.dina(w_n839_0[1]),.dinb(w_G4089_0[2]),.dout(n840),.clk(gclk));
	jand g0540(.dina(w_n840_4[1]),.dinb(w_n791_1[0]),.dout(n841),.clk(gclk));
	jnot g0541(.din(w_G4089_0[1]),.dout(n842),.clk(gclk));
	jand g0542(.dina(w_n839_0[0]),.dinb(w_n842_0[1]),.dout(n843),.clk(gclk));
	jand g0543(.dina(w_n843_4[1]),.dinb(w_n795_1[0]),.dout(n844),.clk(gclk));
	jand g0544(.dina(w_G4090_0[1]),.dinb(w_n842_0[0]),.dout(n845),.clk(gclk));
	jand g0545(.dina(w_n845_4[1]),.dinb(w_G11_0[0]),.dout(n846),.clk(gclk));
	jand g0546(.dina(w_G4090_0[0]),.dinb(w_G4089_0[0]),.dout(n847),.clk(gclk));
	jand g0547(.dina(w_n847_4[1]),.dinb(w_G61_0[0]),.dout(n848),.clk(gclk));
	jcb g0548(.dina(w_dff_B_Mw5zA2y87_0),.dinb(n846),.dout(n849));
	jcb g0549(.dina(w_dff_B_rySoRXaP3_0),.dinb(n844),.dout(n850));
	jcb g0550(.dina(w_dff_B_Y4WLp8Fb2_0),.dinb(n841),.dout(G859));
	jnot g0551(.din(w_n678_0[0]),.dout(n852),.clk(gclk));
	jnot g0552(.din(w_n679_0[0]),.dout(n853),.clk(gclk));
	jcb g0553(.dina(w_n583_1[0]),.dinb(w_n574_0[1]),.dout(n854));
	jand g0554(.dina(n854),.dinb(w_n691_0[1]),.dout(n855),.clk(gclk));
	jnot g0555(.din(w_n855_0[1]),.dout(n856),.clk(gclk));
	jnot g0556(.din(w_n691_0[0]),.dout(n857),.clk(gclk));
	jcb g0557(.dina(w_n857_0[1]),.dinb(w_G4_1[0]),.dout(n858));
	jand g0558(.dina(w_dff_B_sGff82Uf3_0),.dinb(w_n856_0[1]),.dout(n859),.clk(gclk));
	jcb g0559(.dina(w_n859_0[1]),.dinb(w_n853_0[1]),.dout(n860));
	jand g0560(.dina(n860),.dinb(w_dff_B_4Us65xLQ6_1),.dout(n861),.clk(gclk));
	jxor g0561(.dina(n861),.dinb(w_n562_0[0]),.dout(n862),.clk(gclk));
	jcb g0562(.dina(w_n862_0[1]),.dinb(w_n748_2[2]),.dout(n863));
	jcb g0563(.dina(w_n765_4[1]),.dinb(w_n470_0[0]),.dout(n864));
	jand g0564(.dina(w_n753_6[1]),.dinb(w_dff_B_X0msDUlY1_1),.dout(n865),.clk(gclk));
	jnot g0565(.din(n865),.dout(n866),.clk(gclk));
	jand g0566(.dina(n866),.dinb(w_dff_B_HM2nPqvS0_1),.dout(n867),.clk(gclk));
	jand g0567(.dina(w_dff_B_HpKf3Jb22_0),.dinb(n863),.dout(G871_fa_),.clk(gclk));
	jxor g0568(.dina(w_n859_0[0]),.dinb(w_n578_0[1]),.dout(n869),.clk(gclk));
	jcb g0569(.dina(w_n869_0[1]),.dinb(w_n748_2[1]),.dout(n870));
	jcb g0570(.dina(w_n765_4[0]),.dinb(w_n481_0[0]),.dout(n871));
	jand g0571(.dina(w_n753_6[0]),.dinb(w_dff_B_HRMR7rpT2_1),.dout(n872),.clk(gclk));
	jnot g0572(.din(n872),.dout(n873),.clk(gclk));
	jand g0573(.dina(n873),.dinb(w_dff_B_VWz7lHXZ8_1),.dout(n874),.clk(gclk));
	jand g0574(.dina(w_dff_B_I14rXkob3_0),.dinb(n870),.dout(G873_fa_),.clk(gclk));
	jand g0575(.dina(w_n567_0[2]),.dinb(w_G4_0[2]),.dout(n876),.clk(gclk));
	jnot g0576(.din(n876),.dout(n877),.clk(gclk));
	jand g0577(.dina(w_n877_0[1]),.dinb(w_n681_2[0]),.dout(n878),.clk(gclk));
	jcb g0578(.dina(n878),.dinb(w_n571_0[2]),.dout(n879));
	jand g0579(.dina(w_n879_0[1]),.dinb(w_n687_0[1]),.dout(n880),.clk(gclk));
	jxor g0580(.dina(n880),.dinb(w_n583_0[2]),.dout(n881),.clk(gclk));
	jand g0581(.dina(w_n881_0[1]),.dinb(w_n747_3[0]),.dout(n882),.clk(gclk));
	jnot g0582(.din(n882),.dout(n883),.clk(gclk));
	jcb g0583(.dina(w_n765_3[2]),.dinb(w_n459_0[0]),.dout(n884));
	jand g0584(.dina(w_n753_5[2]),.dinb(w_dff_B_oY61uKLk2_1),.dout(n885),.clk(gclk));
	jnot g0585(.din(n885),.dout(n886),.clk(gclk));
	jand g0586(.dina(n886),.dinb(w_dff_B_UhDPWxwS4_1),.dout(n887),.clk(gclk));
	jand g0587(.dina(w_dff_B_cPsXwyo38_0),.dinb(n883),.dout(G875_fa_),.clk(gclk));
	jand g0588(.dina(w_n571_0[1]),.dinb(w_n681_1[2]),.dout(n889),.clk(gclk));
	jand g0589(.dina(w_dff_B_fSP7FxFs7_0),.dinb(w_n877_0[0]),.dout(n890),.clk(gclk));
	jnot g0590(.din(n890),.dout(n891),.clk(gclk));
	jand g0591(.dina(n891),.dinb(w_n879_0[0]),.dout(n892),.clk(gclk));
	jand g0592(.dina(w_n892_0[1]),.dinb(w_n747_2[2]),.dout(n893),.clk(gclk));
	jnot g0593(.din(n893),.dout(n894),.clk(gclk));
	jcb g0594(.dina(w_n765_3[1]),.dinb(w_n494_0[0]),.dout(n895));
	jand g0595(.dina(w_n753_5[1]),.dinb(w_dff_B_4LuH5Jpo9_1),.dout(n896),.clk(gclk));
	jnot g0596(.din(n896),.dout(n897),.clk(gclk));
	jand g0597(.dina(n897),.dinb(w_dff_B_eT3Orvrj8_1),.dout(n898),.clk(gclk));
	jand g0598(.dina(w_dff_B_OfAy3uSm0_0),.dinb(n894),.dout(G877_fa_),.clk(gclk));
	jxor g0599(.dina(w_n649_0[2]),.dinb(w_n735_0[0]),.dout(n900),.clk(gclk));
	jxor g0600(.dina(w_dff_B_VurSCaJD9_0),.dinb(w_n786_0[0]),.dout(n901),.clk(gclk));
	jxor g0601(.dina(n901),.dinb(w_n621_1[0]),.dout(n902),.clk(gclk));
	jand g0602(.dina(w_G369_0[0]),.dinb(w_n609_1[2]),.dout(n903),.clk(gclk));
	jand g0603(.dina(G372),.dinb(w_G332_1[1]),.dout(n904),.clk(gclk));
	jcb g0604(.dina(w_dff_B_F4wIN6jS5_0),.dinb(n903),.dout(n905));
	jxor g0605(.dina(n905),.dinb(w_n617_0[1]),.dout(n906),.clk(gclk));
	jxor g0606(.dina(n906),.dinb(w_n628_0[1]),.dout(n907),.clk(gclk));
	jnot g0607(.din(w_G331_0[0]),.dout(n908),.clk(gclk));
	jand g0608(.dina(w_n624_0[2]),.dinb(w_dff_B_mqvQ6SXx6_1),.dout(n909),.clk(gclk));
	jnot g0609(.din(w_n624_0[1]),.dout(n910),.clk(gclk));
	jand g0610(.dina(w_dff_B_9t3Iv5XK3_0),.dinb(w_n613_0[0]),.dout(n911),.clk(gclk));
	jcb g0611(.dina(n911),.dinb(w_dff_B_XFaalHQD9_1),.dout(n912));
	jxor g0612(.dina(n912),.dinb(w_dff_B_KLnd0Szl5_1),.dout(n913),.clk(gclk));
	jxor g0613(.dina(w_dff_B_Qqtg0nxm7_0),.dinb(n902),.dout(n914),.clk(gclk));
	jnot g0614(.din(w_n914_0[1]),.dout(G998),.clk(gclk));
	jxor g0615(.dina(w_n577_0[0]),.dinb(w_n566_0[0]),.dout(n916),.clk(gclk));
	jxor g0616(.dina(w_n582_0[1]),.dinb(w_n570_0[0]),.dout(n917),.clk(gclk));
	jxor g0617(.dina(n917),.dinb(n916),.dout(n918),.clk(gclk));
	jxor g0618(.dina(n918),.dinb(w_n590_0[1]),.dout(n919),.clk(gclk));
	jand g0619(.dina(w_n556_1[2]),.dinb(w_G289_0[0]),.dout(n920),.clk(gclk));
	jand g0620(.dina(w_G335_1[1]),.dinb(G292),.dout(n921),.clk(gclk));
	jcb g0621(.dina(w_dff_B_c1NEaN4f0_0),.dinb(n920),.dout(n922));
	jxor g0622(.dina(n922),.dinb(w_n600_0[2]),.dout(n923),.clk(gclk));
	jxor g0623(.dina(w_dff_B_lpWqvyMa2_0),.dinb(w_n560_0[1]),.dout(n924),.clk(gclk));
	jxor g0624(.dina(w_n604_0[0]),.dinb(w_n595_0[1]),.dout(n925),.clk(gclk));
	jxor g0625(.dina(n925),.dinb(n924),.dout(n926),.clk(gclk));
	jxor g0626(.dina(n926),.dinb(w_dff_B_mfm0ebpX6_1),.dout(G1000_fa_),.clk(gclk));
	jnot g0627(.din(w_n596_0[1]),.dout(n928),.clk(gclk));
	jnot g0628(.din(w_n707_0[1]),.dout(n929),.clk(gclk));
	jnot g0629(.din(w_n700_0[0]),.dout(n930),.clk(gclk));
	jnot g0630(.din(w_n605_2[0]),.dout(n931),.clk(gclk));
	jnot g0631(.din(w_n601_0[0]),.dout(n932),.clk(gclk));
	jnot g0632(.din(w_n696_0[1]),.dout(n933),.clk(gclk));
	jand g0633(.dina(w_n587_1[0]),.dinb(w_G4_0[1]),.dout(n934),.clk(gclk));
	jnot g0634(.din(n934),.dout(n935),.clk(gclk));
	jand g0635(.dina(n935),.dinb(n933),.dout(n936),.clk(gclk));
	jcb g0636(.dina(w_n936_0[2]),.dinb(w_n932_0[1]),.dout(n937));
	jcb g0637(.dina(n937),.dinb(w_dff_B_fQWhak0j7_1),.dout(n938));
	jcb g0638(.dina(w_n938_0[1]),.dinb(w_n930_0[2]),.dout(n939));
	jand g0639(.dina(n939),.dinb(w_dff_B_nrpAOopt1_1),.dout(n940),.clk(gclk));
	jxor g0640(.dina(n940),.dinb(w_n928_0[1]),.dout(n941),.clk(gclk));
	jnot g0641(.din(w_n941_0[1]),.dout(n942),.clk(gclk));
	jnot g0642(.din(w_n591_0[0]),.dout(n943),.clk(gclk));
	jnot g0643(.din(w_n705_0[0]),.dout(n944),.clk(gclk));
	jand g0644(.dina(w_n938_0[0]),.dinb(w_n944_0[1]),.dout(n945),.clk(gclk));
	jxor g0645(.dina(n945),.dinb(w_n943_0[1]),.dout(n946),.clk(gclk));
	jnot g0646(.din(w_n946_0[1]),.dout(n947),.clk(gclk));
	jcb g0647(.dina(w_n600_0[1]),.dinb(w_G422_1[0]),.dout(n948));
	jnot g0648(.din(w_n948_0[2]),.dout(n949),.clk(gclk));
	jnot g0649(.din(w_n703_0[1]),.dout(n950),.clk(gclk));
	jand g0650(.dina(w_n936_0[1]),.dinb(w_dff_B_rNTWf0vb8_1),.dout(n951),.clk(gclk));
	jcb g0651(.dina(n951),.dinb(w_dff_B_0RClE1oJ5_1),.dout(n952));
	jxor g0652(.dina(n952),.dinb(w_n605_1[2]),.dout(n953),.clk(gclk));
	jxor g0653(.dina(w_n936_0[0]),.dinb(w_n932_0[0]),.dout(n954),.clk(gclk));
	jnot g0654(.din(w_n954_0[1]),.dout(n955),.clk(gclk));
	jnot g0655(.din(w_n881_0[0]),.dout(n956),.clk(gclk));
	jnot g0656(.din(w_n771_0[0]),.dout(n957),.clk(gclk));
	jnot g0657(.din(w_n892_0[0]),.dout(n958),.clk(gclk));
	jand g0658(.dina(n958),.dinb(w_dff_B_Cc4JLWJc2_1),.dout(n959),.clk(gclk));
	jand g0659(.dina(n959),.dinb(w_dff_B_DxRhincp4_1),.dout(n960),.clk(gclk));
	jand g0660(.dina(n960),.dinb(w_n869_0[0]),.dout(n961),.clk(gclk));
	jand g0661(.dina(n961),.dinb(w_n862_0[0]),.dout(n962),.clk(gclk));
	jand g0662(.dina(n962),.dinb(w_dff_B_aGPEn6zR7_1),.dout(n963),.clk(gclk));
	jand g0663(.dina(n963),.dinb(w_n953_0[1]),.dout(n964),.clk(gclk));
	jand g0664(.dina(n964),.dinb(w_dff_B_dSMLp7Iu5_1),.dout(n965),.clk(gclk));
	jand g0665(.dina(n965),.dinb(w_dff_B_FLk7yXTK9_1),.dout(G575),.clk(gclk));
	jnot g0666(.din(w_n646_0[1]),.dout(n967),.clk(gclk));
	jcb g0667(.dina(w_n649_0[1]),.dinb(w_G490_0[1]),.dout(n968));
	jcb g0668(.dina(w_n781_0[1]),.dinb(w_n739_1[0]),.dout(n969));
	jand g0669(.dina(n969),.dinb(w_n968_0[1]),.dout(n970),.clk(gclk));
	jxor g0670(.dina(n970),.dinb(w_dff_B_jfGC3CN29_1),.dout(n971),.clk(gclk));
	jxor g0671(.dina(w_n783_0[2]),.dinb(w_n640_1[0]),.dout(n972),.clk(gclk));
	jxor g0672(.dina(w_n781_0[0]),.dinb(w_n650_0[0]),.dout(n973),.clk(gclk));
	jnot g0673(.din(w_n973_0[1]),.dout(n974),.clk(gclk));
	jcb g0674(.dina(w_n621_0[2]),.dinb(w_n744_0[1]),.dout(n975));
	jand g0675(.dina(n975),.dinb(w_n636_0[2]),.dout(n976),.clk(gclk));
	jand g0676(.dina(w_dff_B_PlStXqfk4_0),.dinb(w_n761_0[0]),.dout(n977),.clk(gclk));
	jand g0677(.dina(n977),.dinb(w_n832_0[0]),.dout(n978),.clk(gclk));
	jand g0678(.dina(n978),.dinb(w_n821_0[0]),.dout(n979),.clk(gclk));
	jand g0679(.dina(n979),.dinb(w_n809_0[0]),.dout(n980),.clk(gclk));
	jand g0680(.dina(n980),.dinb(n974),.dout(n981),.clk(gclk));
	jand g0681(.dina(n981),.dinb(w_n972_0[1]),.dout(n982),.clk(gclk));
	jand g0682(.dina(n982),.dinb(w_n971_0[1]),.dout(G585),.clk(gclk));
	jnot g0683(.din(w_G1690_0[2]),.dout(n984),.clk(gclk));
	jand g0684(.dina(w_n984_0[1]),.dinb(w_G1689_0[2]),.dout(n985),.clk(gclk));
	jand g0685(.dina(w_n985_4[1]),.dinb(w_n791_0[2]),.dout(n986),.clk(gclk));
	jnot g0686(.din(w_G1689_0[1]),.dout(n987),.clk(gclk));
	jand g0687(.dina(w_n984_0[0]),.dinb(w_n987_0[1]),.dout(n988),.clk(gclk));
	jand g0688(.dina(w_n988_4[1]),.dinb(w_n795_0[2]),.dout(n989),.clk(gclk));
	jand g0689(.dina(w_G1690_0[1]),.dinb(w_n987_0[0]),.dout(n990),.clk(gclk));
	jand g0690(.dina(w_n990_4[1]),.dinb(w_G182_0[1]),.dout(n991),.clk(gclk));
	jand g0691(.dina(w_G1690_0[0]),.dinb(w_G1689_0[0]),.dout(n992),.clk(gclk));
	jand g0692(.dina(w_n992_4[1]),.dinb(w_G185_0[1]),.dout(n993),.clk(gclk));
	jcb g0693(.dina(w_dff_B_4xQBvl2r0_0),.dinb(n991),.dout(n994));
	jcb g0694(.dina(w_dff_B_tOz9RWR58_0),.dinb(n989),.dout(n995));
	jcb g0695(.dina(w_dff_B_2u3sRBDv6_0),.dinb(n986),.dout(n996));
	jand g0696(.dina(n996),.dinb(w_G137_9[1]),.dout(G661),.clk(gclk));
	jnot g0697(.din(w_G1694_0[2]),.dout(n998),.clk(gclk));
	jand g0698(.dina(w_n998_0[1]),.dinb(w_G1691_0[2]),.dout(n999),.clk(gclk));
	jand g0699(.dina(w_n999_4[1]),.dinb(w_n791_0[1]),.dout(n1000),.clk(gclk));
	jnot g0700(.din(w_G1691_0[1]),.dout(n1001),.clk(gclk));
	jand g0701(.dina(w_n998_0[0]),.dinb(w_n1001_0[1]),.dout(n1002),.clk(gclk));
	jand g0702(.dina(w_n1002_4[1]),.dinb(w_n795_0[1]),.dout(n1003),.clk(gclk));
	jand g0703(.dina(w_G1694_0[1]),.dinb(w_n1001_0[0]),.dout(n1004),.clk(gclk));
	jand g0704(.dina(w_n1004_4[1]),.dinb(w_G182_0[0]),.dout(n1005),.clk(gclk));
	jand g0705(.dina(w_G1694_0[0]),.dinb(w_G1691_0[0]),.dout(n1006),.clk(gclk));
	jand g0706(.dina(w_n1006_4[1]),.dinb(w_G185_0[0]),.dout(n1007),.clk(gclk));
	jcb g0707(.dina(w_dff_B_Slzp9vaC8_0),.dinb(n1005),.dout(n1008));
	jcb g0708(.dina(w_dff_B_IB2lwABJ2_0),.dinb(n1003),.dout(n1009));
	jcb g0709(.dina(w_dff_B_KpZXeaHc9_0),.dinb(n1000),.dout(n1010));
	jand g0710(.dina(n1010),.dinb(w_G137_9[0]),.dout(G693),.clk(gclk));
	jnot g0711(.din(w_G871_0),.dout(n1012),.clk(gclk));
	jand g0712(.dina(w_n1012_1[1]),.dinb(w_n793_4[0]),.dout(n1013),.clk(gclk));
	jnot g0713(.din(w_G832_0),.dout(n1014),.clk(gclk));
	jand g0714(.dina(w_n1014_1[1]),.dinb(w_n797_4[0]),.dout(n1015),.clk(gclk));
	jand g0715(.dina(w_n799_4[0]),.dinb(w_G43_0[1]),.dout(n1016),.clk(gclk));
	jand g0716(.dina(w_n801_4[0]),.dinb(w_G37_0[1]),.dout(n1017),.clk(gclk));
	jcb g0717(.dina(w_dff_B_yzh2W3DX2_0),.dinb(n1016),.dout(n1018));
	jcb g0718(.dina(w_dff_B_QwYmrZtN6_0),.dinb(n1015),.dout(n1019));
	jcb g0719(.dina(w_dff_B_TBw81uok5_0),.dinb(n1013),.dout(G747));
	jnot g0720(.din(w_G873_0),.dout(n1021),.clk(gclk));
	jand g0721(.dina(w_n1021_1[1]),.dinb(w_n793_3[2]),.dout(n1022),.clk(gclk));
	jnot g0722(.din(w_G834_0),.dout(n1023),.clk(gclk));
	jand g0723(.dina(w_n1023_1[1]),.dinb(w_n797_3[2]),.dout(n1024),.clk(gclk));
	jand g0724(.dina(w_n799_3[2]),.dinb(w_G76_0[1]),.dout(n1025),.clk(gclk));
	jand g0725(.dina(w_n801_3[2]),.dinb(w_G20_0[1]),.dout(n1026),.clk(gclk));
	jcb g0726(.dina(w_dff_B_EFOHvvMd4_0),.dinb(n1025),.dout(n1027));
	jcb g0727(.dina(w_dff_B_0l4ExStx1_0),.dinb(n1024),.dout(n1028));
	jcb g0728(.dina(w_dff_B_SYCIhiJY9_0),.dinb(n1022),.dout(G752));
	jnot g0729(.din(w_G875_0),.dout(n1030),.clk(gclk));
	jand g0730(.dina(w_n1030_1[1]),.dinb(w_n793_3[1]),.dout(n1031),.clk(gclk));
	jnot g0731(.din(w_G836_0),.dout(n1032),.clk(gclk));
	jand g0732(.dina(w_n1032_1[1]),.dinb(w_n797_3[1]),.dout(n1033),.clk(gclk));
	jand g0733(.dina(w_n799_3[1]),.dinb(w_G73_0[1]),.dout(n1034),.clk(gclk));
	jand g0734(.dina(w_n801_3[1]),.dinb(w_G17_0[1]),.dout(n1035),.clk(gclk));
	jcb g0735(.dina(w_dff_B_1C1cxjdS6_0),.dinb(n1034),.dout(n1036));
	jcb g0736(.dina(w_dff_B_Lr4O21im4_0),.dinb(n1033),.dout(n1037));
	jcb g0737(.dina(w_dff_B_CTXroHMd3_0),.dinb(n1031),.dout(G757));
	jnot g0738(.din(w_G877_0),.dout(n1039),.clk(gclk));
	jand g0739(.dina(w_n1039_1[1]),.dinb(w_n793_3[0]),.dout(n1040),.clk(gclk));
	jnot g0740(.din(w_G838_0),.dout(n1041),.clk(gclk));
	jand g0741(.dina(w_n797_3[0]),.dinb(w_n1041_1[1]),.dout(n1042),.clk(gclk));
	jand g0742(.dina(w_n799_3[0]),.dinb(w_G67_0[1]),.dout(n1043),.clk(gclk));
	jand g0743(.dina(w_n801_3[0]),.dinb(w_G70_0[1]),.dout(n1044),.clk(gclk));
	jcb g0744(.dina(w_dff_B_Yr3r80KN9_0),.dinb(n1043),.dout(n1045));
	jcb g0745(.dina(w_dff_B_XCdzVBk76_0),.dinb(n1042),.dout(n1046));
	jcb g0746(.dina(w_dff_B_c8kVFgYn3_0),.dinb(n1040),.dout(G762));
	jand g0747(.dina(w_n1012_1[0]),.dinb(w_n840_4[0]),.dout(n1048),.clk(gclk));
	jand g0748(.dina(w_n843_4[0]),.dinb(w_n1014_1[0]),.dout(n1049),.clk(gclk));
	jand g0749(.dina(w_n845_4[0]),.dinb(w_G43_0[0]),.dout(n1050),.clk(gclk));
	jand g0750(.dina(w_n847_4[0]),.dinb(w_G37_0[0]),.dout(n1051),.clk(gclk));
	jcb g0751(.dina(w_dff_B_pW89VdJt3_0),.dinb(n1050),.dout(n1052));
	jcb g0752(.dina(w_dff_B_cQsrr4c32_0),.dinb(n1049),.dout(n1053));
	jcb g0753(.dina(w_dff_B_oef3wOMR0_0),.dinb(n1048),.dout(G787));
	jand g0754(.dina(w_n1021_1[0]),.dinb(w_n840_3[2]),.dout(n1055),.clk(gclk));
	jand g0755(.dina(w_n843_3[2]),.dinb(w_n1023_1[0]),.dout(n1056),.clk(gclk));
	jand g0756(.dina(w_n845_3[2]),.dinb(w_G76_0[0]),.dout(n1057),.clk(gclk));
	jand g0757(.dina(w_n847_3[2]),.dinb(w_G20_0[0]),.dout(n1058),.clk(gclk));
	jcb g0758(.dina(w_dff_B_GaCqMgtu1_0),.dinb(n1057),.dout(n1059));
	jcb g0759(.dina(w_dff_B_TNC4Qb987_0),.dinb(n1056),.dout(n1060));
	jcb g0760(.dina(w_dff_B_wNxtMbtO6_0),.dinb(n1055),.dout(G792));
	jand g0761(.dina(w_n1030_1[0]),.dinb(w_n840_3[1]),.dout(n1062),.clk(gclk));
	jand g0762(.dina(w_n843_3[1]),.dinb(w_n1032_1[0]),.dout(n1063),.clk(gclk));
	jand g0763(.dina(w_n845_3[1]),.dinb(w_G73_0[0]),.dout(n1064),.clk(gclk));
	jand g0764(.dina(w_n847_3[1]),.dinb(w_G17_0[0]),.dout(n1065),.clk(gclk));
	jcb g0765(.dina(w_dff_B_9FV3cLIM8_0),.dinb(n1064),.dout(n1066));
	jcb g0766(.dina(w_dff_B_JurtH47K4_0),.dinb(n1063),.dout(n1067));
	jcb g0767(.dina(w_dff_B_59nKBC3D3_0),.dinb(n1062),.dout(G797));
	jand g0768(.dina(w_n1039_1[0]),.dinb(w_n840_3[0]),.dout(n1069),.clk(gclk));
	jand g0769(.dina(w_n843_3[0]),.dinb(w_n1041_1[0]),.dout(n1070),.clk(gclk));
	jand g0770(.dina(w_n845_3[0]),.dinb(w_G67_0[0]),.dout(n1071),.clk(gclk));
	jand g0771(.dina(w_n847_3[0]),.dinb(w_G70_0[0]),.dout(n1072),.clk(gclk));
	jcb g0772(.dina(w_dff_B_mvLIU5Ui7_0),.dinb(n1071),.dout(n1073));
	jcb g0773(.dina(w_dff_B_wBIa7dao0_0),.dinb(n1070),.dout(n1074));
	jcb g0774(.dina(w_dff_B_Wv0NtsIA4_0),.dinb(n1069),.dout(G802));
	jand g0775(.dina(w_n985_4[0]),.dinb(w_n1012_0[2]),.dout(n1076),.clk(gclk));
	jand g0776(.dina(w_n988_4[0]),.dinb(w_n1014_0[2]),.dout(n1077),.clk(gclk));
	jand g0777(.dina(w_n990_4[0]),.dinb(w_G200_0[1]),.dout(n1078),.clk(gclk));
	jand g0778(.dina(w_n992_4[0]),.dinb(w_G170_0[1]),.dout(n1079),.clk(gclk));
	jcb g0779(.dina(w_dff_B_1b6BJ2b44_0),.dinb(n1078),.dout(n1080));
	jcb g0780(.dina(w_dff_B_Gf4T2pe65_0),.dinb(n1077),.dout(n1081));
	jcb g0781(.dina(w_dff_B_1IWmYF6w0_0),.dinb(n1076),.dout(n1082));
	jand g0782(.dina(n1082),.dinb(w_G137_8[2]),.dout(G642),.clk(gclk));
	jand g0783(.dina(w_n985_3[2]),.dinb(w_n1039_0[2]),.dout(n1084),.clk(gclk));
	jand g0784(.dina(w_n988_3[2]),.dinb(w_n1041_0[2]),.dout(n1085),.clk(gclk));
	jand g0785(.dina(w_n990_3[2]),.dinb(w_G188_0[1]),.dout(n1086),.clk(gclk));
	jand g0786(.dina(w_n992_3[2]),.dinb(w_G158_0[1]),.dout(n1087),.clk(gclk));
	jcb g0787(.dina(w_dff_B_Pwkrnbqn8_0),.dinb(n1086),.dout(n1088));
	jcb g0788(.dina(w_dff_B_fXQYtvhd2_0),.dinb(n1085),.dout(n1089));
	jcb g0789(.dina(w_dff_B_x8TsiQby5_0),.dinb(n1084),.dout(n1090));
	jand g0790(.dina(n1090),.dinb(w_G137_8[1]),.dout(G664),.clk(gclk));
	jand g0791(.dina(w_n985_3[1]),.dinb(w_n1030_0[2]),.dout(n1092),.clk(gclk));
	jand g0792(.dina(w_n988_3[1]),.dinb(w_n1032_0[2]),.dout(n1093),.clk(gclk));
	jand g0793(.dina(w_n990_3[1]),.dinb(w_G155_0[1]),.dout(n1094),.clk(gclk));
	jand g0794(.dina(w_n992_3[1]),.dinb(w_G152_0[1]),.dout(n1095),.clk(gclk));
	jcb g0795(.dina(w_dff_B_C4GUCiLi4_0),.dinb(n1094),.dout(n1096));
	jcb g0796(.dina(w_dff_B_o59bURzk6_0),.dinb(n1093),.dout(n1097));
	jcb g0797(.dina(w_dff_B_9GS9SIJm4_0),.dinb(n1092),.dout(n1098));
	jand g0798(.dina(n1098),.dinb(w_G137_8[0]),.dout(G667),.clk(gclk));
	jand g0799(.dina(w_n985_3[0]),.dinb(w_n1021_0[2]),.dout(n1100),.clk(gclk));
	jand g0800(.dina(w_n988_3[0]),.dinb(w_n1023_0[2]),.dout(n1101),.clk(gclk));
	jand g0801(.dina(w_n990_3[0]),.dinb(w_G149_0[1]),.dout(n1102),.clk(gclk));
	jand g0802(.dina(w_n992_3[0]),.dinb(w_G146_0[1]),.dout(n1103),.clk(gclk));
	jcb g0803(.dina(w_dff_B_JcqG57Ro5_0),.dinb(n1102),.dout(n1104));
	jcb g0804(.dina(w_dff_B_1CYes5n85_0),.dinb(n1101),.dout(n1105));
	jcb g0805(.dina(w_dff_B_FJNmdIq07_0),.dinb(n1100),.dout(n1106));
	jand g0806(.dina(n1106),.dinb(w_G137_7[2]),.dout(G670),.clk(gclk));
	jand g0807(.dina(w_n999_4[0]),.dinb(w_n1012_0[1]),.dout(n1108),.clk(gclk));
	jand g0808(.dina(w_n1002_4[0]),.dinb(w_n1014_0[1]),.dout(n1109),.clk(gclk));
	jand g0809(.dina(w_n1004_4[0]),.dinb(w_G200_0[0]),.dout(n1110),.clk(gclk));
	jand g0810(.dina(w_n1006_4[0]),.dinb(w_G170_0[0]),.dout(n1111),.clk(gclk));
	jcb g0811(.dina(w_dff_B_tRGiG3Pb4_0),.dinb(n1110),.dout(n1112));
	jcb g0812(.dina(w_dff_B_c47yMk2V7_0),.dinb(n1109),.dout(n1113));
	jcb g0813(.dina(w_dff_B_43EMR9wJ7_0),.dinb(n1108),.dout(n1114));
	jand g0814(.dina(n1114),.dinb(w_G137_7[1]),.dout(G676),.clk(gclk));
	jand g0815(.dina(w_n999_3[2]),.dinb(w_n1039_0[1]),.dout(n1116),.clk(gclk));
	jand g0816(.dina(w_n1002_3[2]),.dinb(w_n1041_0[1]),.dout(n1117),.clk(gclk));
	jand g0817(.dina(w_n1004_3[2]),.dinb(w_G188_0[0]),.dout(n1118),.clk(gclk));
	jand g0818(.dina(w_n1006_3[2]),.dinb(w_G158_0[0]),.dout(n1119),.clk(gclk));
	jcb g0819(.dina(w_dff_B_HXNCn4GD1_0),.dinb(n1118),.dout(n1120));
	jcb g0820(.dina(w_dff_B_ICQv7vJ08_0),.dinb(n1117),.dout(n1121));
	jcb g0821(.dina(w_dff_B_GVcn3f3y3_0),.dinb(n1116),.dout(n1122));
	jand g0822(.dina(n1122),.dinb(w_G137_7[0]),.dout(G696),.clk(gclk));
	jand g0823(.dina(w_n999_3[1]),.dinb(w_n1030_0[1]),.dout(n1124),.clk(gclk));
	jand g0824(.dina(w_n1002_3[1]),.dinb(w_n1032_0[1]),.dout(n1125),.clk(gclk));
	jand g0825(.dina(w_n1004_3[1]),.dinb(w_G155_0[0]),.dout(n1126),.clk(gclk));
	jand g0826(.dina(w_n1006_3[1]),.dinb(w_G152_0[0]),.dout(n1127),.clk(gclk));
	jcb g0827(.dina(w_dff_B_lGjRA1MP6_0),.dinb(n1126),.dout(n1128));
	jcb g0828(.dina(w_dff_B_wtTfk3g40_0),.dinb(n1125),.dout(n1129));
	jcb g0829(.dina(w_dff_B_i1TJoECv1_0),.dinb(n1124),.dout(n1130));
	jand g0830(.dina(n1130),.dinb(w_G137_6[2]),.dout(G699),.clk(gclk));
	jand g0831(.dina(w_n999_3[0]),.dinb(w_n1021_0[1]),.dout(n1132),.clk(gclk));
	jand g0832(.dina(w_n1002_3[0]),.dinb(w_n1023_0[1]),.dout(n1133),.clk(gclk));
	jand g0833(.dina(w_n1004_3[0]),.dinb(w_G149_0[0]),.dout(n1134),.clk(gclk));
	jand g0834(.dina(w_n1006_3[0]),.dinb(w_G146_0[0]),.dout(n1135),.clk(gclk));
	jcb g0835(.dina(w_dff_B_AdB8vm2y9_0),.dinb(n1134),.dout(n1136));
	jcb g0836(.dina(w_dff_B_Uf2LOJKb1_0),.dinb(n1133),.dout(n1137));
	jcb g0837(.dina(w_dff_B_d6uNA6YY6_0),.dinb(n1132),.dout(n1138));
	jand g0838(.dina(n1138),.dinb(w_G137_6[1]),.dout(G702),.clk(gclk));
	jand g0839(.dina(w_n789_0[1]),.dinb(w_G3724_0[2]),.dout(n1140),.clk(gclk));
	jnot g0840(.din(w_G3717_0[1]),.dout(n1141),.clk(gclk));
	jnot g0841(.din(w_G3724_0[1]),.dout(n1142),.clk(gclk));
	jand g0842(.dina(w_n1142_0[1]),.dinb(w_G123_0[1]),.dout(n1143),.clk(gclk));
	jcb g0843(.dina(n1143),.dinb(w_dff_B_skaBgWq53_1),.dout(n1144));
	jcb g0844(.dina(w_dff_B_ROAuJexP8_0),.dinb(n1140),.dout(n1145));
	jnot g0845(.din(G135),.dout(n1146),.clk(gclk));
	jnot g0846(.din(G4115),.dout(n1147),.clk(gclk));
	jcb g0847(.dina(n1147),.dinb(n1146),.dout(n1148));
	jxor g0848(.dina(w_n636_0[1]),.dinb(w_G132_0[1]),.dout(n1149),.clk(gclk));
	jand g0849(.dina(n1149),.dinb(w_G3724_0[0]),.dout(n1150),.clk(gclk));
	jnot g0850(.din(w_n401_0[1]),.dout(n1151),.clk(gclk));
	jand g0851(.dina(w_n1151_0[1]),.dinb(w_n1142_0[0]),.dout(n1152),.clk(gclk));
	jcb g0852(.dina(n1152),.dinb(w_G3717_0[0]),.dout(n1153));
	jcb g0853(.dina(n1153),.dinb(n1150),.dout(n1154));
	jand g0854(.dina(n1154),.dinb(w_dff_B_8iUufvxb4_1),.dout(n1155),.clk(gclk));
	jand g0855(.dina(w_dff_B_WNZNiIJS5_0),.dinb(n1145),.dout(G818),.clk(gclk));
	jcb g0856(.dina(w_n783_0[1]),.dinb(w_n640_0[2]),.dout(n1157));
	jxor g0857(.dina(n1157),.dinb(w_G132_0[0]),.dout(G813),.clk(gclk));
	jand g0858(.dina(w_n789_0[0]),.dinb(w_n747_2[1]),.dout(n1159),.clk(gclk));
	jand g0859(.dina(w_n753_5[0]),.dinb(w_G123_0[0]),.dout(n1160),.clk(gclk));
	jand g0860(.dina(w_n751_1[1]),.dinb(w_n1151_0[0]),.dout(n1161),.clk(gclk));
	jcb g0861(.dina(n1161),.dinb(w_dff_B_OMwLOQoe0_1),.dout(n1162));
	jcb g0862(.dina(w_dff_B_qUG4y7cK7_0),.dinb(n1159),.dout(n1163));
	jnot g0863(.din(w_n1163_1[2]),.dout(G824),.clk(gclk));
	jcb g0864(.dina(w_n972_0[0]),.dinb(w_n748_2[0]),.dout(n1165));
	jand g0865(.dina(w_n751_1[0]),.dinb(w_n407_0[0]),.dout(n1166),.clk(gclk));
	jand g0866(.dina(w_n753_4[2]),.dinb(w_dff_B_cnWEupaI2_1),.dout(n1167),.clk(gclk));
	jcb g0867(.dina(n1167),.dinb(n1166),.dout(n1168));
	jnot g0868(.din(n1168),.dout(n1169),.clk(gclk));
	jand g0869(.dina(w_dff_B_A49QF9CZ7_0),.dinb(n1165),.dout(G826_fa_),.clk(gclk));
	jcb g0870(.dina(w_n971_0[0]),.dinb(w_n748_1[2]),.dout(n1171));
	jcb g0871(.dina(w_n765_3[0]),.dinb(w_n372_0[1]),.dout(n1172));
	jand g0872(.dina(w_n753_4[1]),.dinb(w_dff_B_R5eMOqaD7_1),.dout(n1173),.clk(gclk));
	jnot g0873(.din(n1173),.dout(n1174),.clk(gclk));
	jand g0874(.dina(n1174),.dinb(w_dff_B_lyCXxF103_1),.dout(n1175),.clk(gclk));
	jand g0875(.dina(w_dff_B_D43eyW007_0),.dinb(n1171),.dout(G828_fa_),.clk(gclk));
	jand g0876(.dina(w_n973_0[0]),.dinb(w_n747_2[0]),.dout(n1177),.clk(gclk));
	jnot g0877(.din(n1177),.dout(n1178),.clk(gclk));
	jcb g0878(.dina(w_n765_2[2]),.dinb(w_n383_0[1]),.dout(n1179));
	jand g0879(.dina(w_n753_4[0]),.dinb(w_dff_B_E0lFfosK4_1),.dout(n1180),.clk(gclk));
	jnot g0880(.din(n1180),.dout(n1181),.clk(gclk));
	jand g0881(.dina(n1181),.dinb(w_dff_B_rriyiCdb7_1),.dout(n1182),.clk(gclk));
	jand g0882(.dina(w_dff_B_SiShHYSa7_0),.dinb(n1178),.dout(G830_fa_),.clk(gclk));
	jnot g0883(.din(w_G1000_0),.dout(n1184),.clk(gclk));
	jand g0884(.dina(w_G559_0[0]),.dinb(w_G245_0[0]),.dout(n1185),.clk(gclk));
	jand g0885(.dina(n1185),.dinb(w_n318_0[0]),.dout(n1186),.clk(gclk));
	jand g0886(.dina(n1186),.dinb(w_G601_0),.dout(n1187),.clk(gclk));
	jand g0887(.dina(w_dff_B_ryzSXgLC1_0),.dinb(w_n661_0[0]),.dout(n1188),.clk(gclk));
	jand g0888(.dina(n1188),.dinb(w_n671_0[0]),.dout(n1189),.clk(gclk));
	jand g0889(.dina(w_dff_B_myBjpaiO4_0),.dinb(w_n914_0[0]),.dout(n1190),.clk(gclk));
	jand g0890(.dina(n1190),.dinb(w_dff_B_OsXxBvxJ0_1),.dout(G854),.clk(gclk));
	jand g0891(.dina(w_n941_0[0]),.dinb(w_n747_1[2]),.dout(n1192),.clk(gclk));
	jnot g0892(.din(w_n528_0[1]),.dout(n1193),.clk(gclk));
	jand g0893(.dina(w_n751_0[2]),.dinb(n1193),.dout(n1194),.clk(gclk));
	jand g0894(.dina(w_n753_3[2]),.dinb(w_dff_B_wxWIjnjD9_1),.dout(n1195),.clk(gclk));
	jcb g0895(.dina(w_dff_B_e9P0BzYN6_0),.dinb(n1194),.dout(n1196));
	jcb g0896(.dina(w_dff_B_J5kFLssw3_0),.dinb(n1192),.dout(n1197));
	jnot g0897(.din(w_n1197_1[2]),.dout(G863),.clk(gclk));
	jand g0898(.dina(w_n946_0[0]),.dinb(w_n747_1[1]),.dout(n1199),.clk(gclk));
	jcb g0899(.dina(w_n765_2[1]),.dinb(w_n551_0[0]),.dout(n1200));
	jand g0900(.dina(w_n753_3[1]),.dinb(w_dff_B_nyZz9qgn8_1),.dout(n1201),.clk(gclk));
	jnot g0901(.din(n1201),.dout(n1202),.clk(gclk));
	jand g0902(.dina(n1202),.dinb(w_dff_B_GDnjo22a3_1),.dout(n1203),.clk(gclk));
	jnot g0903(.din(n1203),.dout(n1204),.clk(gclk));
	jcb g0904(.dina(w_dff_B_y5jcS6ZD3_0),.dinb(n1199),.dout(n1205));
	jnot g0905(.din(w_n1205_1[2]),.dout(G865),.clk(gclk));
	jcb g0906(.dina(w_n953_0[0]),.dinb(w_n748_1[1]),.dout(n1207));
	jcb g0907(.dina(w_n765_2[0]),.dinb(w_n517_0[0]),.dout(n1208));
	jand g0908(.dina(w_n753_3[0]),.dinb(w_dff_B_EreY5MCq2_1),.dout(n1209),.clk(gclk));
	jnot g0909(.din(n1209),.dout(n1210),.clk(gclk));
	jand g0910(.dina(n1210),.dinb(w_dff_B_UrrZoGXb3_1),.dout(n1211),.clk(gclk));
	jand g0911(.dina(w_dff_B_XiAZqJNi4_0),.dinb(n1207),.dout(G867_fa_),.clk(gclk));
	jand g0912(.dina(w_n954_0[0]),.dinb(w_n747_1[0]),.dout(n1213),.clk(gclk));
	jnot g0913(.din(n1213),.dout(n1214),.clk(gclk));
	jcb g0914(.dina(w_n765_1[2]),.dinb(w_n540_0[0]),.dout(n1215));
	jand g0915(.dina(w_n753_2[2]),.dinb(w_dff_B_JdJmN8DZ9_1),.dout(n1216),.clk(gclk));
	jnot g0916(.din(n1216),.dout(n1217),.clk(gclk));
	jand g0917(.dina(n1217),.dinb(w_dff_B_1XCOXLIU0_1),.dout(n1218),.clk(gclk));
	jand g0918(.dina(w_dff_B_LaggcDo98_0),.dinb(n1214),.dout(G869_fa_),.clk(gclk));
	jand g0919(.dina(w_n1197_1[1]),.dinb(w_n840_2[2]),.dout(n1220),.clk(gclk));
	jand g0920(.dina(w_n1163_1[1]),.dinb(w_n843_2[2]),.dout(n1221),.clk(gclk));
	jand g0921(.dina(w_n845_2[2]),.dinb(w_G109_0[1]),.dout(n1222),.clk(gclk));
	jand g0922(.dina(w_n847_2[2]),.dinb(w_G106_0[1]),.dout(n1223),.clk(gclk));
	jcb g0923(.dina(w_dff_B_e8e7yQGH2_0),.dinb(n1222),.dout(n1224));
	jcb g0924(.dina(w_dff_B_lcRHJFF64_0),.dinb(n1221),.dout(n1225));
	jcb g0925(.dina(w_dff_B_nAmKSWzQ8_0),.dinb(n1220),.dout(G712));
	jand g0926(.dina(w_n1197_1[0]),.dinb(w_n793_2[2]),.dout(n1227),.clk(gclk));
	jand g0927(.dina(w_n1163_1[0]),.dinb(w_n797_2[2]),.dout(n1228),.clk(gclk));
	jand g0928(.dina(w_n799_2[2]),.dinb(w_G109_0[0]),.dout(n1229),.clk(gclk));
	jand g0929(.dina(w_n801_2[2]),.dinb(w_G106_0[0]),.dout(n1230),.clk(gclk));
	jcb g0930(.dina(w_dff_B_D1GTF7xj2_0),.dinb(n1229),.dout(n1231));
	jcb g0931(.dina(w_dff_B_lBEKmMGR7_0),.dinb(n1228),.dout(n1232));
	jcb g0932(.dina(w_dff_B_YVGo4UPM2_0),.dinb(n1227),.dout(G727));
	jand g0933(.dina(w_n1205_1[1]),.dinb(w_n793_2[1]),.dout(n1234),.clk(gclk));
	jnot g0934(.din(w_G826_0),.dout(n1235),.clk(gclk));
	jand g0935(.dina(w_n1235_1[1]),.dinb(w_n797_2[1]),.dout(n1236),.clk(gclk));
	jand g0936(.dina(w_n799_2[1]),.dinb(w_G46_0[1]),.dout(n1237),.clk(gclk));
	jand g0937(.dina(w_n801_2[1]),.dinb(w_G49_0[1]),.dout(n1238),.clk(gclk));
	jcb g0938(.dina(w_dff_B_jdyTFGON9_0),.dinb(n1237),.dout(n1239));
	jcb g0939(.dina(w_dff_B_9lyVfhjn2_0),.dinb(n1236),.dout(n1240));
	jcb g0940(.dina(w_dff_B_4kLkfKo12_0),.dinb(n1234),.dout(G732));
	jnot g0941(.din(w_G867_0),.dout(n1242),.clk(gclk));
	jand g0942(.dina(w_n1242_1[1]),.dinb(w_n793_2[0]),.dout(n1243),.clk(gclk));
	jnot g0943(.din(w_G828_0),.dout(n1244),.clk(gclk));
	jand g0944(.dina(w_n1244_1[1]),.dinb(w_n797_2[0]),.dout(n1245),.clk(gclk));
	jand g0945(.dina(w_n799_2[0]),.dinb(w_G100_0[1]),.dout(n1246),.clk(gclk));
	jand g0946(.dina(w_n801_2[0]),.dinb(w_G103_0[1]),.dout(n1247),.clk(gclk));
	jcb g0947(.dina(w_dff_B_8J0lArrZ8_0),.dinb(n1246),.dout(n1248));
	jcb g0948(.dina(w_dff_B_YBXa6sB24_0),.dinb(n1245),.dout(n1249));
	jcb g0949(.dina(w_dff_B_KEvTavOV0_0),.dinb(n1243),.dout(G737));
	jnot g0950(.din(w_G869_0),.dout(n1251),.clk(gclk));
	jand g0951(.dina(w_n1251_1[1]),.dinb(w_n793_1[2]),.dout(n1252),.clk(gclk));
	jnot g0952(.din(w_G830_0),.dout(n1253),.clk(gclk));
	jand g0953(.dina(w_n1253_1[1]),.dinb(w_n797_1[2]),.dout(n1254),.clk(gclk));
	jand g0954(.dina(w_n799_1[2]),.dinb(w_G91_0[1]),.dout(n1255),.clk(gclk));
	jand g0955(.dina(w_n801_1[2]),.dinb(w_G40_0[1]),.dout(n1256),.clk(gclk));
	jcb g0956(.dina(w_dff_B_By08MlUX8_0),.dinb(n1255),.dout(n1257));
	jcb g0957(.dina(w_dff_B_6M8cMGMJ4_0),.dinb(n1254),.dout(n1258));
	jcb g0958(.dina(w_dff_B_XS8AGY9p0_0),.dinb(n1252),.dout(G742));
	jand g0959(.dina(w_n1205_1[0]),.dinb(w_n840_2[1]),.dout(n1260),.clk(gclk));
	jand g0960(.dina(w_n1235_1[0]),.dinb(w_n843_2[1]),.dout(n1261),.clk(gclk));
	jand g0961(.dina(w_n845_2[1]),.dinb(w_G46_0[0]),.dout(n1262),.clk(gclk));
	jand g0962(.dina(w_n847_2[1]),.dinb(w_G49_0[0]),.dout(n1263),.clk(gclk));
	jcb g0963(.dina(w_dff_B_V3RaC9xA7_0),.dinb(n1262),.dout(n1264));
	jcb g0964(.dina(w_dff_B_eTqwgJac6_0),.dinb(n1261),.dout(n1265));
	jcb g0965(.dina(w_dff_B_5NMMGf1M8_0),.dinb(n1260),.dout(G772));
	jand g0966(.dina(w_n1242_1[0]),.dinb(w_n840_2[0]),.dout(n1267),.clk(gclk));
	jand g0967(.dina(w_n1244_1[0]),.dinb(w_n843_2[0]),.dout(n1268),.clk(gclk));
	jand g0968(.dina(w_n845_2[0]),.dinb(w_G100_0[0]),.dout(n1269),.clk(gclk));
	jand g0969(.dina(w_n847_2[0]),.dinb(w_G103_0[0]),.dout(n1270),.clk(gclk));
	jcb g0970(.dina(w_dff_B_f6ms2hRU9_0),.dinb(n1269),.dout(n1271));
	jcb g0971(.dina(w_dff_B_qLP4lseT5_0),.dinb(n1268),.dout(n1272));
	jcb g0972(.dina(w_dff_B_LqaCsD8p8_0),.dinb(n1267),.dout(G777));
	jand g0973(.dina(w_n1251_1[0]),.dinb(w_n840_1[2]),.dout(n1274),.clk(gclk));
	jand g0974(.dina(w_n1253_1[0]),.dinb(w_n843_1[2]),.dout(n1275),.clk(gclk));
	jand g0975(.dina(w_n845_1[2]),.dinb(w_G91_0[0]),.dout(n1276),.clk(gclk));
	jand g0976(.dina(w_n847_1[2]),.dinb(w_G40_0[0]),.dout(n1277),.clk(gclk));
	jcb g0977(.dina(w_dff_B_q20txiL02_0),.dinb(n1276),.dout(n1278));
	jcb g0978(.dina(w_dff_B_d8DnDGOF9_0),.dinb(n1275),.dout(n1279));
	jcb g0979(.dina(w_dff_B_1JF1dcMV9_0),.dinb(n1274),.dout(G782));
	jand g0980(.dina(w_n1251_0[2]),.dinb(w_n985_2[2]),.dout(n1281),.clk(gclk));
	jand g0981(.dina(w_n1253_0[2]),.dinb(w_n988_2[2]),.dout(n1282),.clk(gclk));
	jand g0982(.dina(w_n990_2[2]),.dinb(w_G203_0[1]),.dout(n1283),.clk(gclk));
	jand g0983(.dina(w_n992_2[2]),.dinb(w_G173_0[1]),.dout(n1284),.clk(gclk));
	jcb g0984(.dina(w_dff_B_Cx88I4iO0_0),.dinb(n1283),.dout(n1285));
	jcb g0985(.dina(w_dff_B_Lv9JQ9Y06_0),.dinb(n1282),.dout(n1286));
	jcb g0986(.dina(w_dff_B_m3koI63o4_0),.dinb(n1281),.dout(n1287));
	jand g0987(.dina(n1287),.dinb(w_G137_6[0]),.dout(G645),.clk(gclk));
	jand g0988(.dina(w_n1242_0[2]),.dinb(w_n985_2[1]),.dout(n1289),.clk(gclk));
	jand g0989(.dina(w_n1244_0[2]),.dinb(w_n988_2[1]),.dout(n1290),.clk(gclk));
	jand g0990(.dina(w_n990_2[1]),.dinb(w_G197_0[1]),.dout(n1291),.clk(gclk));
	jand g0991(.dina(w_n992_2[1]),.dinb(w_G167_0[1]),.dout(n1292),.clk(gclk));
	jcb g0992(.dina(w_dff_B_BgYH8FIF4_0),.dinb(n1291),.dout(n1293));
	jcb g0993(.dina(w_dff_B_xcUtQedf4_0),.dinb(n1290),.dout(n1294));
	jcb g0994(.dina(w_dff_B_Uw33huRr7_0),.dinb(n1289),.dout(n1295));
	jand g0995(.dina(n1295),.dinb(w_G137_5[2]),.dout(G648),.clk(gclk));
	jand g0996(.dina(w_n1205_0[2]),.dinb(w_n985_2[0]),.dout(n1297),.clk(gclk));
	jand g0997(.dina(w_n1235_0[2]),.dinb(w_n988_2[0]),.dout(n1298),.clk(gclk));
	jand g0998(.dina(w_n990_2[0]),.dinb(w_G194_0[1]),.dout(n1299),.clk(gclk));
	jand g0999(.dina(w_n992_2[0]),.dinb(w_G164_0[1]),.dout(n1300),.clk(gclk));
	jcb g1000(.dina(w_dff_B_2NvQOqmD9_0),.dinb(n1299),.dout(n1301));
	jcb g1001(.dina(w_dff_B_fdPo0AZw9_0),.dinb(n1298),.dout(n1302));
	jcb g1002(.dina(w_dff_B_U6uAs9no9_0),.dinb(n1297),.dout(n1303));
	jand g1003(.dina(n1303),.dinb(w_G137_5[1]),.dout(G651),.clk(gclk));
	jand g1004(.dina(w_n1197_0[2]),.dinb(w_n985_1[2]),.dout(n1305),.clk(gclk));
	jand g1005(.dina(w_n1163_0[2]),.dinb(w_n988_1[2]),.dout(n1306),.clk(gclk));
	jand g1006(.dina(w_n990_1[2]),.dinb(w_G191_0[1]),.dout(n1307),.clk(gclk));
	jand g1007(.dina(w_n992_1[2]),.dinb(w_G161_0[1]),.dout(n1308),.clk(gclk));
	jcb g1008(.dina(w_dff_B_o5e6IOru5_0),.dinb(n1307),.dout(n1309));
	jcb g1009(.dina(w_dff_B_iU3KJzgu0_0),.dinb(n1306),.dout(n1310));
	jcb g1010(.dina(w_dff_B_EtmPvepO1_0),.dinb(n1305),.dout(n1311));
	jand g1011(.dina(n1311),.dinb(w_G137_5[0]),.dout(G654),.clk(gclk));
	jand g1012(.dina(w_n1251_0[1]),.dinb(w_n999_2[2]),.dout(n1313),.clk(gclk));
	jand g1013(.dina(w_n1253_0[1]),.dinb(w_n1002_2[2]),.dout(n1314),.clk(gclk));
	jand g1014(.dina(w_n1004_2[2]),.dinb(w_G203_0[0]),.dout(n1315),.clk(gclk));
	jand g1015(.dina(w_n1006_2[2]),.dinb(w_G173_0[0]),.dout(n1316),.clk(gclk));
	jcb g1016(.dina(w_dff_B_4PSQfdGY6_0),.dinb(n1315),.dout(n1317));
	jcb g1017(.dina(w_dff_B_tiqgSRIB6_0),.dinb(n1314),.dout(n1318));
	jcb g1018(.dina(w_dff_B_x5UCoTEU2_0),.dinb(n1313),.dout(n1319));
	jand g1019(.dina(n1319),.dinb(w_G137_4[2]),.dout(G679),.clk(gclk));
	jand g1020(.dina(w_n1242_0[1]),.dinb(w_n999_2[1]),.dout(n1321),.clk(gclk));
	jand g1021(.dina(w_n1244_0[1]),.dinb(w_n1002_2[1]),.dout(n1322),.clk(gclk));
	jand g1022(.dina(w_n1004_2[1]),.dinb(w_G197_0[0]),.dout(n1323),.clk(gclk));
	jand g1023(.dina(w_n1006_2[1]),.dinb(w_G167_0[0]),.dout(n1324),.clk(gclk));
	jcb g1024(.dina(w_dff_B_vy9ULEa11_0),.dinb(n1323),.dout(n1325));
	jcb g1025(.dina(w_dff_B_Eeolb1wv2_0),.dinb(n1322),.dout(n1326));
	jcb g1026(.dina(w_dff_B_faGCYL2X9_0),.dinb(n1321),.dout(n1327));
	jand g1027(.dina(n1327),.dinb(w_G137_4[1]),.dout(G682),.clk(gclk));
	jand g1028(.dina(w_n1205_0[1]),.dinb(w_n999_2[0]),.dout(n1329),.clk(gclk));
	jand g1029(.dina(w_n1235_0[1]),.dinb(w_n1002_2[0]),.dout(n1330),.clk(gclk));
	jand g1030(.dina(w_n1004_2[0]),.dinb(w_G194_0[0]),.dout(n1331),.clk(gclk));
	jand g1031(.dina(w_n1006_2[0]),.dinb(w_G164_0[0]),.dout(n1332),.clk(gclk));
	jcb g1032(.dina(w_dff_B_q8GF83v79_0),.dinb(n1331),.dout(n1333));
	jcb g1033(.dina(w_dff_B_TeA0l5RY6_0),.dinb(n1330),.dout(n1334));
	jcb g1034(.dina(w_dff_B_OeLX3bdT2_0),.dinb(n1329),.dout(n1335));
	jand g1035(.dina(n1335),.dinb(w_G137_4[0]),.dout(G685),.clk(gclk));
	jand g1036(.dina(w_n1197_0[1]),.dinb(w_n999_1[2]),.dout(n1337),.clk(gclk));
	jand g1037(.dina(w_n1163_0[1]),.dinb(w_n1002_1[2]),.dout(n1338),.clk(gclk));
	jand g1038(.dina(w_n1004_1[2]),.dinb(w_G191_0[0]),.dout(n1339),.clk(gclk));
	jand g1039(.dina(w_n1006_1[2]),.dinb(w_G161_0[0]),.dout(n1340),.clk(gclk));
	jcb g1040(.dina(w_dff_B_VdR7OR9Q3_0),.dinb(n1339),.dout(n1341));
	jcb g1041(.dina(w_dff_B_yy97jijI8_0),.dinb(n1338),.dout(n1342));
	jcb g1042(.dina(w_dff_B_qtFJrn8I0_0),.dinb(n1337),.dout(n1343));
	jand g1043(.dina(n1343),.dinb(w_G137_3[2]),.dout(G688),.clk(gclk));
	jcb g1044(.dina(w_G4091_2[0]),.dinb(G120),.dout(n1345));
	jand g1045(.dina(w_n435_0[2]),.dinb(w_G251_3[1]),.dout(n1346),.clk(gclk));
	jand g1046(.dina(w_G341_1[0]),.dinb(w_G248_4[0]),.dout(n1347),.clk(gclk));
	jcb g1047(.dina(n1347),.dinb(w_n437_0[1]),.dout(n1348));
	jcb g1048(.dina(w_dff_B_aHlrTtf12_0),.dinb(n1346),.dout(n1349));
	jand g1049(.dina(w_n435_0[1]),.dinb(w_n366_3[1]),.dout(n1350),.clk(gclk));
	jand g1050(.dina(w_G341_0[2]),.dinb(w_n368_4[0]),.dout(n1351),.clk(gclk));
	jcb g1051(.dina(n1351),.dinb(w_G523_0[2]),.dout(n1352));
	jcb g1052(.dina(n1352),.dinb(n1350),.dout(n1353));
	jand g1053(.dina(n1353),.dinb(n1349),.dout(n1354),.clk(gclk));
	jxor g1054(.dina(w_n408_0[0]),.dinb(w_n401_0[0]),.dout(n1355),.clk(gclk));
	jxor g1055(.dina(w_n383_0[0]),.dinb(w_n372_0[0]),.dout(n1356),.clk(gclk));
	jxor g1056(.dina(n1356),.dinb(n1355),.dout(n1357),.clk(gclk));
	jxor g1057(.dina(n1357),.dinb(w_dff_B_BboVEPTk3_1),.dout(n1358),.clk(gclk));
	jnot g1058(.din(w_n1358_0[1]),.dout(n1359),.clk(gclk));
	jcb g1059(.dina(w_n410_0[1]),.dinb(w_G248_3[2]),.dout(n1360));
	jcb g1060(.dina(w_G514_0[1]),.dinb(w_n368_3[2]),.dout(n1361));
	jand g1061(.dina(n1361),.dinb(n1360),.dout(n1362),.clk(gclk));
	jxor g1062(.dina(n1362),.dinb(w_n419_0[0]),.dout(n1363),.clk(gclk));
	jcb g1063(.dina(w_G351_1[0]),.dinb(w_n402_1[2]),.dout(n1364));
	jcb g1064(.dina(w_n385_0[2]),.dinb(w_n405_1[2]),.dout(n1365));
	jand g1065(.dina(n1365),.dinb(w_G534_0[1]),.dout(n1366),.clk(gclk));
	jand g1066(.dina(n1366),.dinb(w_dff_B_aVuxNvvi6_1),.dout(n1367),.clk(gclk));
	jcb g1067(.dina(w_G351_0[2]),.dinb(w_G254_1[1]),.dout(n1368));
	jcb g1068(.dina(w_n385_0[1]),.dinb(w_G242_1[1]),.dout(n1369));
	jand g1069(.dina(n1369),.dinb(w_n388_0[1]),.dout(n1370),.clk(gclk));
	jand g1070(.dina(n1370),.dinb(w_dff_B_mWIbgAuX5_1),.dout(n1371),.clk(gclk));
	jcb g1071(.dina(n1371),.dinb(n1367),.dout(n1372));
	jand g1072(.dina(w_n424_1[0]),.dinb(w_G251_3[0]),.dout(n1373),.clk(gclk));
	jand g1073(.dina(w_G324_0[2]),.dinb(w_G248_3[1]),.dout(n1374),.clk(gclk));
	jcb g1074(.dina(n1374),.dinb(w_n426_0[0]),.dout(n1375));
	jcb g1075(.dina(w_dff_B_5NGtMF6T2_0),.dinb(n1373),.dout(n1376));
	jand g1076(.dina(w_n424_0[2]),.dinb(w_n366_3[0]),.dout(n1377),.clk(gclk));
	jand g1077(.dina(w_G324_0[1]),.dinb(w_n368_3[1]),.dout(n1378),.clk(gclk));
	jcb g1078(.dina(n1378),.dinb(w_G503_0[1]),.dout(n1379));
	jcb g1079(.dina(n1379),.dinb(n1377),.dout(n1380));
	jand g1080(.dina(n1380),.dinb(n1376),.dout(n1381),.clk(gclk));
	jxor g1081(.dina(n1381),.dinb(n1372),.dout(n1382),.clk(gclk));
	jxor g1082(.dina(n1382),.dinb(w_dff_B_Q4zcJ1XI4_1),.dout(n1383),.clk(gclk));
	jnot g1083(.din(w_n1383_0[1]),.dout(n1384),.clk(gclk));
	jand g1084(.dina(w_n1383_0[0]),.dinb(n1359),.dout(n1385),.clk(gclk));
	jcb g1085(.dina(n1385),.dinb(w_G4091_1[2]),.dout(n1386));
	jcb g1086(.dina(w_dff_B_B99ennDR0_0),.dinb(w_n746_1[0]),.dout(n1388));
	jand g1087(.dina(n1384),.dinb(w_n1358_0[0]),.dout(n1389),.clk(gclk));
	jcb g1088(.dina(n1386),.dinb(w_dff_B_ERBCSkDC7_1),.dout(n1390));
	jand g1089(.dina(n1390),.dinb(w_n746_0[2]),.dout(n1391),.clk(gclk));
	jnot g1090(.din(w_n1391_0[1]),.dout(n1392),.clk(gclk));
	jand g1091(.dina(w_n633_0[2]),.dinb(w_G2174_0[2]),.dout(n1393),.clk(gclk));
	jcb g1092(.dina(n1393),.dinb(w_n732_0[0]),.dout(n1394));
	jand g1093(.dina(w_n736_0[0]),.dinb(w_n640_0[1]),.dout(n1395),.clk(gclk));
	jcb g1094(.dina(w_n740_0[0]),.dinb(w_n641_0[0]),.dout(n1396));
	jand g1095(.dina(n1396),.dinb(w_n646_0[0]),.dout(n1397),.clk(gclk));
	jcb g1096(.dina(n1397),.dinb(w_dff_B_PnB00RFh4_1),.dout(n1398));
	jnot g1097(.din(w_n1398_0[1]),.dout(n1399),.clk(gclk));
	jand g1098(.dina(w_n1399_0[1]),.dinb(w_n739_0[2]),.dout(n1400),.clk(gclk));
	jnot g1099(.din(w_n739_0[1]),.dout(n1401),.clk(gclk));
	jand g1100(.dina(w_n1398_0[0]),.dinb(w_dff_B_rufnpOUb5_1),.dout(n1402),.clk(gclk));
	jcb g1101(.dina(n1402),.dinb(w_n651_0[1]),.dout(n1403));
	jcb g1102(.dina(w_dff_B_NI9LZYTr6_0),.dinb(n1400),.dout(n1404));
	jand g1103(.dina(n1404),.dinb(w_n1394_0[1]),.dout(n1405),.clk(gclk));
	jnot g1104(.din(w_n1394_0[0]),.dout(n1406),.clk(gclk));
	jxor g1105(.dina(w_n1399_0[0]),.dinb(w_n968_0[0]),.dout(n1407),.clk(gclk));
	jand g1106(.dina(n1407),.dinb(n1406),.dout(n1408),.clk(gclk));
	jcb g1107(.dina(n1408),.dinb(n1405),.dout(n1409));
	jnot g1108(.din(w_n1409_0[1]),.dout(n1410),.clk(gclk));
	jxor g1109(.dina(w_n629_0[0]),.dinb(w_n625_0[0]),.dout(n1411),.clk(gclk));
	jnot g1110(.din(w_n1411_0[1]),.dout(n1412),.clk(gclk));
	jxor g1111(.dina(w_n806_0[1]),.dinb(w_n828_0[1]),.dout(n1413),.clk(gclk));
	jnot g1112(.din(w_n614_1[1]),.dout(n1414),.clk(gclk));
	jnot g1113(.din(w_n717_0[0]),.dout(n1415),.clk(gclk));
	jand g1114(.dina(w_n622_1[0]),.dinb(w_n828_0[0]),.dout(n1416),.clk(gclk));
	jand g1115(.dina(w_n628_0[0]),.dinb(w_G523_0[1]),.dout(n1417),.clk(gclk));
	jcb g1116(.dina(n1417),.dinb(w_n829_0[0]),.dout(n1418));
	jcb g1117(.dina(w_dff_B_kv5PswOs4_0),.dinb(n1416),.dout(n1419));
	jand g1118(.dina(n1419),.dinb(n1415),.dout(n1420),.clk(gclk));
	jxor g1119(.dina(w_n622_0[2]),.dinb(w_n618_0[1]),.dout(n1421),.clk(gclk));
	jnot g1120(.din(w_n1421_0[1]),.dout(n1422),.clk(gclk));
	jcb g1121(.dina(n1422),.dinb(n1420),.dout(n1423));
	jcb g1122(.dina(w_n1421_0[0]),.dinb(w_n819_0[0]),.dout(n1424));
	jand g1123(.dina(n1424),.dinb(n1423),.dout(n1425),.clk(gclk));
	jxor g1124(.dina(w_n1425_0[1]),.dinb(n1414),.dout(n1426),.clk(gclk));
	jand g1125(.dina(n1426),.dinb(n1413),.dout(n1427),.clk(gclk));
	jnot g1126(.din(w_G2174_0[1]),.dout(n1428),.clk(gclk));
	jxor g1127(.dina(w_n806_0[0]),.dinb(w_n721_0[1]),.dout(n1429),.clk(gclk));
	jxor g1128(.dina(w_n1425_0[0]),.dinb(w_n614_1[0]),.dout(n1430),.clk(gclk));
	jand g1129(.dina(n1430),.dinb(n1429),.dout(n1431),.clk(gclk));
	jcb g1130(.dina(n1431),.dinb(w_dff_B_M8LVzLZV3_1),.dout(n1432));
	jcb g1131(.dina(n1432),.dinb(n1427),.dout(n1433));
	jxor g1132(.dina(w_n729_0[1]),.dinb(w_n614_0[2]),.dout(n1434),.clk(gclk));
	jnot g1133(.din(w_n1434_0[1]),.dout(n1435),.clk(gclk));
	jcb g1134(.dina(w_n622_0[1]),.dinb(w_n721_0[0]),.dout(n1436));
	jand g1135(.dina(n1436),.dinb(w_n723_0[0]),.dout(n1437),.clk(gclk));
	jxor g1136(.dina(n1437),.dinb(w_n727_0[0]),.dout(n1438),.clk(gclk));
	jand g1137(.dina(w_n1438_0[1]),.dinb(n1435),.dout(n1439),.clk(gclk));
	jnot g1138(.din(w_n1438_0[0]),.dout(n1440),.clk(gclk));
	jand g1139(.dina(n1440),.dinb(w_n1434_0[0]),.dout(n1441),.clk(gclk));
	jcb g1140(.dina(n1441),.dinb(w_G2174_0[0]),.dout(n1442));
	jcb g1141(.dina(w_dff_B_F6BENzHa7_0),.dinb(n1439),.dout(n1443));
	jand g1142(.dina(n1443),.dinb(n1433),.dout(n1444),.clk(gclk));
	jxor g1143(.dina(n1444),.dinb(w_n787_0[0]),.dout(n1445),.clk(gclk));
	jxor g1144(.dina(w_n1445_0[1]),.dinb(w_dff_B_ulOgNjix6_1),.dout(n1446),.clk(gclk));
	jcb g1145(.dina(w_n1446_0[1]),.dinb(w_n1410_0[1]),.dout(n1447));
	jxor g1146(.dina(w_n1445_0[0]),.dinb(w_n1411_0[0]),.dout(n1448),.clk(gclk));
	jcb g1147(.dina(n1448),.dinb(w_n1409_0[0]),.dout(n1449));
	jand g1148(.dina(n1449),.dinb(w_G4091_1[1]),.dout(n1450),.clk(gclk));
	jand g1149(.dina(n1450),.dinb(w_n1447_0[1]),.dout(n1451),.clk(gclk));
	jcb g1150(.dina(n1451),.dinb(w_dff_B_Zd4hGI9Q4_1),.dout(n1452));
	jand g1151(.dina(w_n1452_0[1]),.dinb(w_dff_B_zAIAJcVN6_1),.dout(G843),.clk(gclk));
	jcb g1152(.dina(w_G4091_1[0]),.dinb(G118),.dout(n1454));
	jand g1153(.dina(w_G251_2[2]),.dinb(w_n460_0[2]),.dout(n1455),.clk(gclk));
	jand g1154(.dina(w_G248_3[0]),.dinb(w_G234_1[0]),.dout(n1456),.clk(gclk));
	jcb g1155(.dina(n1456),.dinb(w_n462_0[0]),.dout(n1457));
	jcb g1156(.dina(w_dff_B_EYGPxgol6_0),.dinb(n1455),.dout(n1458));
	jand g1157(.dina(w_n366_2[2]),.dinb(w_n460_0[1]),.dout(n1459),.clk(gclk));
	jand g1158(.dina(w_n368_3[0]),.dinb(w_G234_0[2]),.dout(n1460),.clk(gclk));
	jcb g1159(.dina(n1460),.dinb(w_G435_0[1]),.dout(n1461));
	jcb g1160(.dina(n1461),.dinb(n1459),.dout(n1462));
	jand g1161(.dina(n1462),.dinb(n1458),.dout(n1463),.clk(gclk));
	jcb g1162(.dina(w_n402_1[1]),.dinb(w_G226_1[0]),.dout(n1464));
	jcb g1163(.dina(w_n405_1[1]),.dinb(w_n530_0[2]),.dout(n1465));
	jand g1164(.dina(n1465),.dinb(w_G422_0[2]),.dout(n1466),.clk(gclk));
	jand g1165(.dina(n1466),.dinb(w_dff_B_P4UFu9w18_1),.dout(n1467),.clk(gclk));
	jcb g1166(.dina(w_G254_1[0]),.dinb(w_G226_0[2]),.dout(n1468));
	jcb g1167(.dina(w_G242_1[0]),.dinb(w_n530_0[1]),.dout(n1469));
	jand g1168(.dina(n1469),.dinb(w_n532_0[0]),.dout(n1470),.clk(gclk));
	jand g1169(.dina(n1470),.dinb(w_dff_B_weVoAiYu5_1),.dout(n1471),.clk(gclk));
	jcb g1170(.dina(n1471),.dinb(n1467),.dout(n1472));
	jxor g1171(.dina(n1472),.dinb(w_n528_0[0]),.dout(n1473),.clk(gclk));
	jcb g1172(.dina(w_n402_1[0]),.dinb(w_G218_1[0]),.dout(n1474));
	jcb g1173(.dina(w_n405_1[0]),.dinb(w_n507_0[2]),.dout(n1475));
	jand g1174(.dina(n1475),.dinb(w_G468_0[1]),.dout(n1476),.clk(gclk));
	jand g1175(.dina(n1476),.dinb(w_dff_B_rPkfXDut9_1),.dout(n1477),.clk(gclk));
	jcb g1176(.dina(w_G254_0[2]),.dinb(w_G218_0[2]),.dout(n1478));
	jcb g1177(.dina(w_G242_0[2]),.dinb(w_n507_0[1]),.dout(n1479));
	jand g1178(.dina(n1479),.dinb(w_n509_0[0]),.dout(n1480),.clk(gclk));
	jand g1179(.dina(n1480),.dinb(w_dff_B_ufvP6d3X3_1),.dout(n1481),.clk(gclk));
	jcb g1180(.dina(n1481),.dinb(n1477),.dout(n1482));
	jand g1181(.dina(w_G251_2[1]),.dinb(w_n541_0[2]),.dout(n1483),.clk(gclk));
	jand g1182(.dina(w_G248_2[2]),.dinb(w_G210_1[0]),.dout(n1484),.clk(gclk));
	jcb g1183(.dina(n1484),.dinb(w_n543_0[0]),.dout(n1485));
	jcb g1184(.dina(w_dff_B_4jxE2WRh1_0),.dinb(n1483),.dout(n1486));
	jand g1185(.dina(w_n366_2[1]),.dinb(w_n541_0[1]),.dout(n1487),.clk(gclk));
	jand g1186(.dina(w_n368_2[2]),.dinb(w_G210_0[2]),.dout(n1488),.clk(gclk));
	jcb g1187(.dina(n1488),.dinb(w_G457_0[2]),.dout(n1489));
	jcb g1188(.dina(n1489),.dinb(n1487),.dout(n1490));
	jand g1189(.dina(n1490),.dinb(n1486),.dout(n1491),.clk(gclk));
	jxor g1190(.dina(n1491),.dinb(n1482),.dout(n1492),.clk(gclk));
	jxor g1191(.dina(n1492),.dinb(n1473),.dout(n1493),.clk(gclk));
	jxor g1192(.dina(n1493),.dinb(w_dff_B_1gVAaMPB9_1),.dout(n1494),.clk(gclk));
	jand g1193(.dina(w_n495_0[2]),.dinb(w_G251_2[0]),.dout(n1495),.clk(gclk));
	jand g1194(.dina(w_G281_1[0]),.dinb(w_G248_2[1]),.dout(n1496),.clk(gclk));
	jcb g1195(.dina(n1496),.dinb(w_n497_0[1]),.dout(n1497));
	jcb g1196(.dina(w_dff_B_bIs2Ifyb2_0),.dinb(n1495),.dout(n1498));
	jand g1197(.dina(w_n495_0[1]),.dinb(w_n366_2[0]),.dout(n1499),.clk(gclk));
	jand g1198(.dina(w_G281_0[2]),.dinb(w_n368_2[1]),.dout(n1500),.clk(gclk));
	jcb g1199(.dina(n1500),.dinb(w_G374_0[0]),.dout(n1501));
	jcb g1200(.dina(n1501),.dinb(n1499),.dout(n1502));
	jand g1201(.dina(n1502),.dinb(n1498),.dout(n1503),.clk(gclk));
	jand g1202(.dina(w_n449_0[2]),.dinb(w_G251_1[2]),.dout(n1504),.clk(gclk));
	jand g1203(.dina(w_G265_1[0]),.dinb(w_G248_2[0]),.dout(n1505),.clk(gclk));
	jcb g1204(.dina(n1505),.dinb(w_n451_0[1]),.dout(n1506));
	jcb g1205(.dina(w_dff_B_c7KuWy6q2_0),.dinb(n1504),.dout(n1507));
	jand g1206(.dina(w_n449_0[1]),.dinb(w_n366_1[2]),.dout(n1508),.clk(gclk));
	jand g1207(.dina(w_G265_0[2]),.dinb(w_n368_2[0]),.dout(n1509),.clk(gclk));
	jcb g1208(.dina(n1509),.dinb(w_G400_0[1]),.dout(n1510));
	jcb g1209(.dina(n1510),.dinb(n1508),.dout(n1511));
	jand g1210(.dina(n1511),.dinb(n1507),.dout(n1512),.clk(gclk));
	jxor g1211(.dina(n1512),.dinb(n1503),.dout(n1513),.clk(gclk));
	jcb g1212(.dina(w_G257_1[0]),.dinb(w_n402_0[2]),.dout(n1514));
	jcb g1213(.dina(w_n471_0[2]),.dinb(w_n405_0[2]),.dout(n1515));
	jand g1214(.dina(n1515),.dinb(w_G389_0[0]),.dout(n1516),.clk(gclk));
	jand g1215(.dina(n1516),.dinb(w_dff_B_qAzlFbbr0_1),.dout(n1517),.clk(gclk));
	jcb g1216(.dina(w_G257_0[2]),.dinb(w_G254_0[1]),.dout(n1518));
	jcb g1217(.dina(w_n471_0[1]),.dinb(w_G242_0[1]),.dout(n1519));
	jand g1218(.dina(n1519),.dinb(w_n473_0[1]),.dout(n1520),.clk(gclk));
	jand g1219(.dina(n1520),.dinb(w_dff_B_gegiqUQb2_1),.dout(n1521),.clk(gclk));
	jcb g1220(.dina(n1521),.dinb(n1517),.dout(n1522));
	jand g1221(.dina(w_n484_0[2]),.dinb(w_G251_1[1]),.dout(n1523),.clk(gclk));
	jand g1222(.dina(w_G273_1[0]),.dinb(w_G248_1[2]),.dout(n1524),.clk(gclk));
	jcb g1223(.dina(n1524),.dinb(w_n486_0[1]),.dout(n1525));
	jcb g1224(.dina(w_dff_B_nuDczt3V7_0),.dinb(n1523),.dout(n1526));
	jand g1225(.dina(w_n484_0[1]),.dinb(w_n366_1[1]),.dout(n1527),.clk(gclk));
	jand g1226(.dina(w_G273_0[2]),.dinb(w_n368_1[2]),.dout(n1528),.clk(gclk));
	jcb g1227(.dina(n1528),.dinb(w_G411_0[0]),.dout(n1529));
	jcb g1228(.dina(n1529),.dinb(n1527),.dout(n1530));
	jand g1229(.dina(n1530),.dinb(n1526),.dout(n1531),.clk(gclk));
	jxor g1230(.dina(n1531),.dinb(n1522),.dout(n1532),.clk(gclk));
	jxor g1231(.dina(n1532),.dinb(n1513),.dout(n1533),.clk(gclk));
	jand g1232(.dina(w_n1533_0[1]),.dinb(w_n1494_0[1]),.dout(n1534),.clk(gclk));
	jnot g1233(.din(n1534),.dout(n1535),.clk(gclk));
	jcb g1234(.dina(w_n1533_0[0]),.dinb(w_n1494_0[0]),.dout(n1536));
	jand g1235(.dina(n1536),.dinb(w_n750_0[2]),.dout(n1537),.clk(gclk));
	jand g1236(.dina(w_dff_B_fZBBz8PT9_0),.dinb(n1535),.dout(n1538),.clk(gclk));
	jcb g1237(.dina(w_dff_B_htnjqMlm6_0),.dinb(w_n746_0[1]),.dout(n1539));
	jcb g1238(.dina(n1538),.dinb(w_G4092_1[0]),.dout(n1540));
	jxor g1239(.dina(w_n583_0[1]),.dinb(w_n578_0[0]),.dout(n1541),.clk(gclk));
	jxor g1240(.dina(n1541),.dinb(w_n943_0[0]),.dout(n1542),.clk(gclk));
	jnot g1241(.din(n1542),.dout(n1543),.clk(gclk));
	jand g1242(.dina(w_n587_0[2]),.dinb(w_G1497_0[2]),.dout(n1544),.clk(gclk));
	jcb g1243(.dina(n1544),.dinb(w_n696_0[0]),.dout(n1545));
	jnot g1244(.din(w_n1545_0[1]),.dout(n1546),.clk(gclk));
	jcb g1245(.dina(w_n944_0[0]),.dinb(w_n930_0[1]),.dout(n1547));
	jand g1246(.dina(n1547),.dinb(w_n706_0[0]),.dout(n1548),.clk(gclk));
	jxor g1247(.dina(n1548),.dinb(w_n928_0[0]),.dout(n1549),.clk(gclk));
	jxor g1248(.dina(w_n605_1[1]),.dinb(w_n948_0[1]),.dout(n1550),.clk(gclk));
	jxor g1249(.dina(w_dff_B_ULwlZ6nV6_0),.dinb(n1549),.dout(n1551),.clk(gclk));
	jand g1250(.dina(w_dff_B_3OqlOmy05_0),.dinb(n1546),.dout(n1552),.clk(gclk));
	jxor g1251(.dina(w_n605_1[0]),.dinb(w_n703_0[0]),.dout(n1553),.clk(gclk));
	jand g1252(.dina(w_n605_0[2]),.dinb(w_n948_0[0]),.dout(n1554),.clk(gclk));
	jcb g1253(.dina(n1554),.dinb(w_n702_0[0]),.dout(n1555));
	jnot g1254(.din(w_n1555_0[1]),.dout(n1556),.clk(gclk));
	jcb g1255(.dina(n1556),.dinb(w_n930_0[0]),.dout(n1557));
	jcb g1256(.dina(w_n1555_0[0]),.dinb(w_n707_0[0]),.dout(n1558));
	jand g1257(.dina(n1558),.dinb(n1557),.dout(n1559),.clk(gclk));
	jxor g1258(.dina(n1559),.dinb(w_n596_0[0]),.dout(n1560),.clk(gclk));
	jand g1259(.dina(w_n1560_0[1]),.dinb(w_n1553_0[1]),.dout(n1561),.clk(gclk));
	jnot g1260(.din(n1561),.dout(n1562),.clk(gclk));
	jcb g1261(.dina(w_n1560_0[0]),.dinb(w_n1553_0[0]),.dout(n1563));
	jand g1262(.dina(w_dff_B_VBxjGP5o5_0),.dinb(w_n1545_0[0]),.dout(n1564),.clk(gclk));
	jand g1263(.dina(n1564),.dinb(n1562),.dout(n1565),.clk(gclk));
	jcb g1264(.dina(n1565),.dinb(n1552),.dout(n1566));
	jnot g1265(.din(w_G1497_0[1]),.dout(n1567),.clk(gclk));
	jand g1266(.dina(w_n682_0[0]),.dinb(w_n687_0[0]),.dout(n1568),.clk(gclk));
	jand g1267(.dina(w_n1568_0[1]),.dinb(w_n574_0[0]),.dout(n1569),.clk(gclk));
	jxor g1268(.dina(n1569),.dinb(w_n561_0[1]),.dout(n1570),.clk(gclk));
	jxor g1269(.dina(w_n572_0[1]),.dinb(w_n681_1[1]),.dout(n1571),.clk(gclk));
	jcb g1270(.dina(w_n856_0[0]),.dinb(w_n853_0[0]),.dout(n1572));
	jand g1271(.dina(w_n693_0[1]),.dinb(w_n585_0[0]),.dout(n1573),.clk(gclk));
	jcb g1272(.dina(n1573),.dinb(w_n855_0[0]),.dout(n1574));
	jand g1273(.dina(w_dff_B_ZkE0SPhO5_0),.dinb(n1572),.dout(n1575),.clk(gclk));
	jxor g1274(.dina(n1575),.dinb(w_dff_B_4PpQDkje0_1),.dout(n1576),.clk(gclk));
	jxor g1275(.dina(n1576),.dinb(w_dff_B_903H55d30_1),.dout(n1577),.clk(gclk));
	jcb g1276(.dina(n1577),.dinb(w_dff_B_BMknLLvv6_1),.dout(n1578));
	jxor g1277(.dina(w_n693_0[0]),.dinb(w_n572_0[0]),.dout(n1579),.clk(gclk));
	jcb g1278(.dina(w_n857_0[0]),.dinb(w_n681_1[0]),.dout(n1580));
	jnot g1279(.din(w_n681_0[2]),.dout(n1581),.clk(gclk));
	jcb g1280(.dina(w_n680_0[0]),.dinb(n1581),.dout(n1582));
	jcb g1281(.dina(n1582),.dinb(w_n689_0[0]),.dout(n1583));
	jxor g1282(.dina(n1583),.dinb(w_n567_0[1]),.dout(n1584),.clk(gclk));
	jand g1283(.dina(w_dff_B_PwDiaseQ0_0),.dinb(n1580),.dout(n1585),.clk(gclk));
	jxor g1284(.dina(w_n1568_0[0]),.dinb(w_n561_0[0]),.dout(n1586),.clk(gclk));
	jxor g1285(.dina(n1586),.dinb(n1585),.dout(n1587),.clk(gclk));
	jxor g1286(.dina(n1587),.dinb(w_dff_B_g3O8EnKR9_1),.dout(n1588),.clk(gclk));
	jcb g1287(.dina(n1588),.dinb(w_G1497_0[0]),.dout(n1589));
	jand g1288(.dina(w_dff_B_MMoHMBXD7_0),.dinb(n1578),.dout(n1590),.clk(gclk));
	jxor g1289(.dina(n1590),.dinb(w_dff_B_9sqnuwhk9_1),.dout(n1591),.clk(gclk));
	jand g1290(.dina(w_n1591_0[1]),.dinb(w_n1543_0[1]),.dout(n1592),.clk(gclk));
	jnot g1291(.din(n1592),.dout(n1593),.clk(gclk));
	jcb g1292(.dina(w_n1591_0[0]),.dinb(w_n1543_0[0]),.dout(n1594));
	jand g1293(.dina(n1594),.dinb(w_G4091_0[2]),.dout(n1595),.clk(gclk));
	jand g1294(.dina(w_dff_B_AcB2ERIg3_0),.dinb(n1593),.dout(n1596),.clk(gclk));
	jcb g1295(.dina(n1596),.dinb(w_dff_B_ruE9ChaX7_1),.dout(n1597));
	jand g1296(.dina(w_n1597_0[1]),.dinb(w_dff_B_Pyyd8abY6_1),.dout(G882),.clk(gclk));
	jand g1297(.dina(w_G4092_0[2]),.dinb(G97),.dout(n1599),.clk(gclk));
	jnot g1298(.din(n1599),.dout(n1600),.clk(gclk));
	jand g1299(.dina(w_dff_B_Oddba9KG5_0),.dinb(w_n1597_0[0]),.dout(n1601),.clk(gclk));
	jnot g1300(.din(w_n1601_0[2]),.dout(n1602),.clk(gclk));
	jand g1301(.dina(w_n1602_0[1]),.dinb(w_n793_1[1]),.dout(n1603),.clk(gclk));
	jnot g1302(.din(w_n1447_0[0]),.dout(n1604),.clk(gclk));
	jand g1303(.dina(w_n1446_0[0]),.dinb(w_n1410_0[0]),.dout(n1605),.clk(gclk));
	jcb g1304(.dina(n1605),.dinb(w_n750_0[1]),.dout(n1606));
	jcb g1305(.dina(n1606),.dinb(n1604),.dout(n1607));
	jand g1306(.dina(n1607),.dinb(w_n1391_0[0]),.dout(n1608),.clk(gclk));
	jand g1307(.dina(w_G4092_0[1]),.dinb(G94),.dout(n1609),.clk(gclk));
	jcb g1308(.dina(w_n1609_0[1]),.dinb(n1608),.dout(n1610));
	jand g1309(.dina(w_n1610_0[1]),.dinb(w_n797_1[1]),.dout(n1611),.clk(gclk));
	jand g1310(.dina(w_n799_1[1]),.dinb(w_G14_0[1]),.dout(n1612),.clk(gclk));
	jand g1311(.dina(w_n801_1[1]),.dinb(w_G64_0[1]),.dout(n1613),.clk(gclk));
	jcb g1312(.dina(w_dff_B_VGR9opvU0_0),.dinb(n1612),.dout(n1614));
	jcb g1313(.dina(w_dff_B_1A9Un1F09_0),.dinb(n1611),.dout(n1615));
	jcb g1314(.dina(w_dff_B_8sUGvrK17_0),.dinb(n1603),.dout(G767));
	jand g1315(.dina(w_n1602_0[0]),.dinb(w_n840_1[1]),.dout(n1617),.clk(gclk));
	jand g1316(.dina(w_n1610_0[0]),.dinb(w_n843_1[1]),.dout(n1618),.clk(gclk));
	jand g1317(.dina(w_n845_1[1]),.dinb(w_G14_0[0]),.dout(n1619),.clk(gclk));
	jand g1318(.dina(w_n847_1[1]),.dinb(w_G64_0[0]),.dout(n1620),.clk(gclk));
	jcb g1319(.dina(w_dff_B_TbPXMdHi8_0),.dinb(n1619),.dout(n1621));
	jcb g1320(.dina(w_dff_B_2ozSsQQ30_0),.dinb(n1618),.dout(n1622));
	jcb g1321(.dina(w_dff_B_hOPT3Yyh1_0),.dinb(n1617),.dout(G807));
	jnot g1322(.din(w_G137_3[1]),.dout(n1624),.clk(gclk));
	jnot g1323(.din(w_n985_1[1]),.dout(n1625),.clk(gclk));
	jcb g1324(.dina(w_n1601_0[1]),.dinb(w_dff_B_jecj7M9W1_1),.dout(n1626));
	jnot g1325(.din(w_n988_1[1]),.dout(n1627),.clk(gclk));
	jnot g1326(.din(w_n1609_0[0]),.dout(n1628),.clk(gclk));
	jand g1327(.dina(w_dff_B_YbeTSPWj2_0),.dinb(w_n1452_0[0]),.dout(n1629),.clk(gclk));
	jcb g1328(.dina(w_n1629_0[1]),.dinb(w_dff_B_VaxEOFz65_1),.dout(n1630));
	jnot g1329(.din(G179),.dout(n1631),.clk(gclk));
	jnot g1330(.din(w_n992_1[1]),.dout(n1632),.clk(gclk));
	jcb g1331(.dina(n1632),.dinb(w_n1631_0[1]),.dout(n1633));
	jnot g1332(.din(G176),.dout(n1634),.clk(gclk));
	jnot g1333(.din(w_n990_1[1]),.dout(n1635),.clk(gclk));
	jcb g1334(.dina(n1635),.dinb(w_n1634_0[1]),.dout(n1636));
	jand g1335(.dina(n1636),.dinb(w_dff_B_iLAdrS1b7_1),.dout(n1637),.clk(gclk));
	jand g1336(.dina(w_dff_B_7OXd0QYL8_0),.dinb(n1630),.dout(n1638),.clk(gclk));
	jand g1337(.dina(w_dff_B_eBSRsZqY1_0),.dinb(n1626),.dout(n1639),.clk(gclk));
	jcb g1338(.dina(n1639),.dinb(w_n1624_0[1]),.dout(G658));
	jnot g1339(.din(w_n999_1[1]),.dout(n1641),.clk(gclk));
	jcb g1340(.dina(w_n1601_0[0]),.dinb(w_dff_B_r8TMHfw99_1),.dout(n1642));
	jnot g1341(.din(w_n1002_1[1]),.dout(n1643),.clk(gclk));
	jcb g1342(.dina(w_n1629_0[0]),.dinb(w_dff_B_fOlDPyLf2_1),.dout(n1644));
	jnot g1343(.din(w_n1006_1[1]),.dout(n1645),.clk(gclk));
	jcb g1344(.dina(n1645),.dinb(w_n1631_0[0]),.dout(n1646));
	jnot g1345(.din(w_n1004_1[1]),.dout(n1647),.clk(gclk));
	jcb g1346(.dina(n1647),.dinb(w_n1634_0[0]),.dout(n1648));
	jand g1347(.dina(n1648),.dinb(w_dff_B_j1RoE3pl4_1),.dout(n1649),.clk(gclk));
	jand g1348(.dina(w_dff_B_c0kWm8PA4_0),.dinb(n1644),.dout(n1650),.clk(gclk));
	jand g1349(.dina(w_dff_B_vBojNKb56_0),.dinb(n1642),.dout(n1651),.clk(gclk));
	jcb g1350(.dina(n1651),.dinb(w_n1624_0[0]),.dout(G690));
	jdff g1351(.din(w_G141_1[0]),.dout(G144));
	jdff g1352(.din(w_G293_0[0]),.dout(G298));
	jdff g1353(.din(w_G3173_0[0]),.dout(G973));
	jnot g1354(.din(w_G545_0[1]),.dout(G603),.clk(gclk));
	jnot g1355(.din(w_G545_0[0]),.dout(G604),.clk(gclk));
	jdff g1356(.din(w_G137_3[0]),.dout(G926));
	jdff g1357(.din(w_G141_0[2]),.dout(G923));
	jdff g1358(.din(w_G1_2[0]),.dout(G921));
	jdff g1359(.din(w_G549_0[1]),.dout(G892));
	jdff g1360(.din(w_G299_0[1]),.dout(G887));
	jnot g1361(.din(w_G549_0[0]),.dout(G606),.clk(gclk));
	jdff g1362(.din(w_G1_1[2]),.dout(G993));
	jdff g1363(.din(w_G1_1[1]),.dout(G978));
	jdff g1364(.din(w_G1_1[0]),.dout(G949));
	jdff g1365(.din(w_G1_0[2]),.dout(G939));
	jdff g1366(.din(w_G299_0[0]),.dout(G889));
	jcb g1367(.dina(w_n336_0[0]),.dinb(w_n333_0[0]),.dout(G717));
	jand g1368(.dina(w_n652_0[0]),.dinb(w_n633_0[1]),.dout(G626),.clk(gclk));
	jand g1369(.dina(w_n607_0[0]),.dinb(w_n587_0[1]),.dout(G632),.clk(gclk));
	jcb g1370(.dina(w_n709_0[0]),.dinb(w_n697_0[0]),.dout(G621));
	jcb g1371(.dina(w_n742_0[0]),.dinb(w_n733_0[0]),.dout(G629));
	jspl3 jspl3_w_G1_0(.douta(w_G1_0[0]),.doutb(w_G1_0[1]),.doutc(w_G1_0[2]),.din(G1));
	jspl3 jspl3_w_G1_1(.douta(w_G1_1[0]),.doutb(w_G1_1[1]),.doutc(w_G1_1[2]),.din(w_G1_0[0]));
	jspl jspl_w_G1_2(.douta(w_G1_2[0]),.doutb(w_G1_2[1]),.din(w_G1_0[1]));
	jspl3 jspl3_w_G4_0(.douta(w_G4_0[0]),.doutb(w_dff_A_MNXxV7ES6_1),.doutc(w_G4_0[2]),.din(w_dff_B_gTmA6XQD6_3));
	jspl jspl_w_G4_1(.douta(w_dff_A_xUYhHAIk5_0),.doutb(w_G4_1[1]),.din(w_G4_0[0]));
	jspl jspl_w_G11_0(.douta(w_G11_0[0]),.doutb(w_G11_0[1]),.din(w_dff_B_BiD5EdXq3_2));
	jspl jspl_w_G14_0(.douta(w_G14_0[0]),.doutb(w_G14_0[1]),.din(w_dff_B_Vi4narfa5_2));
	jspl jspl_w_G17_0(.douta(w_G17_0[0]),.doutb(w_G17_0[1]),.din(w_dff_B_933tUGNJ1_2));
	jspl jspl_w_G20_0(.douta(w_G20_0[0]),.doutb(w_G20_0[1]),.din(w_dff_B_8T3VWiob3_2));
	jspl jspl_w_G37_0(.douta(w_G37_0[0]),.doutb(w_G37_0[1]),.din(w_dff_B_xxhTC5x54_2));
	jspl jspl_w_G40_0(.douta(w_G40_0[0]),.doutb(w_G40_0[1]),.din(w_dff_B_zXfMPo1R6_2));
	jspl jspl_w_G43_0(.douta(w_G43_0[0]),.doutb(w_G43_0[1]),.din(w_dff_B_jwtZKyDM4_2));
	jspl jspl_w_G46_0(.douta(w_G46_0[0]),.doutb(w_G46_0[1]),.din(w_dff_B_19FnkAzX5_2));
	jspl jspl_w_G49_0(.douta(w_G49_0[0]),.doutb(w_G49_0[1]),.din(w_dff_B_NNNAuk3Y0_2));
	jspl jspl_w_G54_0(.douta(w_dff_A_6Dvk6O510_0),.doutb(w_G54_0[1]),.din(G54));
	jspl jspl_w_G61_0(.douta(w_G61_0[0]),.doutb(w_G61_0[1]),.din(w_dff_B_OBQcQGTx9_2));
	jspl jspl_w_G64_0(.douta(w_G64_0[0]),.doutb(w_G64_0[1]),.din(w_dff_B_wYeNHq3I4_2));
	jspl jspl_w_G67_0(.douta(w_G67_0[0]),.doutb(w_G67_0[1]),.din(w_dff_B_ebTHCX9D8_2));
	jspl jspl_w_G70_0(.douta(w_G70_0[0]),.doutb(w_G70_0[1]),.din(w_dff_B_evZZUxAQ6_2));
	jspl jspl_w_G73_0(.douta(w_G73_0[0]),.doutb(w_G73_0[1]),.din(w_dff_B_9UiXsHup0_2));
	jspl jspl_w_G76_0(.douta(w_G76_0[0]),.doutb(w_G76_0[1]),.din(w_dff_B_hl6lL76m7_2));
	jspl jspl_w_G91_0(.douta(w_G91_0[0]),.doutb(w_G91_0[1]),.din(w_dff_B_kYuYIcMt3_2));
	jspl jspl_w_G100_0(.douta(w_G100_0[0]),.doutb(w_G100_0[1]),.din(w_dff_B_8Yyyj7RI1_2));
	jspl jspl_w_G103_0(.douta(w_G103_0[0]),.doutb(w_G103_0[1]),.din(w_dff_B_jRX7vECG9_2));
	jspl jspl_w_G106_0(.douta(w_G106_0[0]),.doutb(w_G106_0[1]),.din(w_dff_B_9zaiP92j1_2));
	jspl jspl_w_G109_0(.douta(w_G109_0[0]),.doutb(w_G109_0[1]),.din(w_dff_B_THH2YkVh9_2));
	jspl jspl_w_G123_0(.douta(w_dff_A_Pny1KaRT0_0),.doutb(w_G123_0[1]),.din(w_dff_B_PL0GQhlg7_2));
	jspl jspl_w_G132_0(.douta(w_dff_A_F3dasG4b4_0),.doutb(w_G132_0[1]),.din(w_dff_B_UOzhcatG6_2));
	jspl3 jspl3_w_G137_0(.douta(w_dff_A_a8ZdlOSK8_0),.doutb(w_dff_A_WjS2D61k4_1),.doutc(w_G137_0[2]),.din(G137));
	jspl3 jspl3_w_G137_1(.douta(w_dff_A_vm4mmnSs7_0),.doutb(w_dff_A_LW3Zr75J1_1),.doutc(w_G137_1[2]),.din(w_G137_0[0]));
	jspl3 jspl3_w_G137_2(.douta(w_dff_A_ixpkdBVh1_0),.doutb(w_dff_A_brxb91Nl9_1),.doutc(w_G137_2[2]),.din(w_G137_0[1]));
	jspl3 jspl3_w_G137_3(.douta(w_G137_3[0]),.doutb(w_G137_3[1]),.doutc(w_dff_A_F3DBGDKX0_2),.din(w_G137_0[2]));
	jspl3 jspl3_w_G137_4(.douta(w_G137_4[0]),.doutb(w_dff_A_GSkyqbtI8_1),.doutc(w_dff_A_ENGhT1wc6_2),.din(w_G137_1[0]));
	jspl3 jspl3_w_G137_5(.douta(w_G137_5[0]),.doutb(w_G137_5[1]),.doutc(w_dff_A_8i5JmseF1_2),.din(w_G137_1[1]));
	jspl3 jspl3_w_G137_6(.douta(w_dff_A_8JoHe52a3_0),.doutb(w_G137_6[1]),.doutc(w_G137_6[2]),.din(w_G137_1[2]));
	jspl3 jspl3_w_G137_7(.douta(w_G137_7[0]),.doutb(w_dff_A_mZmQW8xh3_1),.doutc(w_G137_7[2]),.din(w_G137_2[0]));
	jspl3 jspl3_w_G137_8(.douta(w_G137_8[0]),.doutb(w_G137_8[1]),.doutc(w_dff_A_etCgCDAc9_2),.din(w_G137_2[1]));
	jspl jspl_w_G137_9(.douta(w_G137_9[0]),.doutb(w_G137_9[1]),.din(w_G137_2[2]));
	jspl3 jspl3_w_G141_0(.douta(w_G141_0[0]),.doutb(w_G141_0[1]),.doutc(w_G141_0[2]),.din(G141));
	jspl3 jspl3_w_G141_1(.douta(w_G141_1[0]),.doutb(w_dff_A_3bTWSZ4q7_1),.doutc(w_dff_A_gGbZoHhG3_2),.din(w_G141_0[0]));
	jspl3 jspl3_w_G141_2(.douta(w_dff_A_mDj9H6QG7_0),.doutb(w_dff_A_AkhK1X9s5_1),.doutc(w_G141_2[2]),.din(w_G141_0[1]));
	jspl jspl_w_G146_0(.douta(w_G146_0[0]),.doutb(w_G146_0[1]),.din(w_dff_B_uA3DEimy4_2));
	jspl jspl_w_G149_0(.douta(w_G149_0[0]),.doutb(w_G149_0[1]),.din(w_dff_B_EHofCk4u4_2));
	jspl jspl_w_G152_0(.douta(w_G152_0[0]),.doutb(w_G152_0[1]),.din(w_dff_B_F85S2bmz5_2));
	jspl jspl_w_G155_0(.douta(w_G155_0[0]),.doutb(w_G155_0[1]),.din(w_dff_B_tDQP5nyd7_2));
	jspl jspl_w_G158_0(.douta(w_G158_0[0]),.doutb(w_G158_0[1]),.din(w_dff_B_iHtaYKnk5_2));
	jspl jspl_w_G161_0(.douta(w_G161_0[0]),.doutb(w_G161_0[1]),.din(w_dff_B_2SbTkK094_2));
	jspl jspl_w_G164_0(.douta(w_G164_0[0]),.doutb(w_G164_0[1]),.din(w_dff_B_U9xFB3tu4_2));
	jspl jspl_w_G167_0(.douta(w_G167_0[0]),.doutb(w_G167_0[1]),.din(w_dff_B_hpxdS3QY5_2));
	jspl jspl_w_G170_0(.douta(w_G170_0[0]),.doutb(w_G170_0[1]),.din(w_dff_B_IHVmLyWb3_2));
	jspl jspl_w_G173_0(.douta(w_G173_0[0]),.doutb(w_G173_0[1]),.din(w_dff_B_YPRdsmVb0_2));
	jspl jspl_w_G182_0(.douta(w_G182_0[0]),.doutb(w_G182_0[1]),.din(w_dff_B_y7pSZth39_2));
	jspl jspl_w_G185_0(.douta(w_G185_0[0]),.doutb(w_G185_0[1]),.din(w_dff_B_8Yt5X2SC2_2));
	jspl jspl_w_G188_0(.douta(w_G188_0[0]),.doutb(w_G188_0[1]),.din(w_dff_B_NXJzxM3B9_2));
	jspl jspl_w_G191_0(.douta(w_G191_0[0]),.doutb(w_G191_0[1]),.din(w_dff_B_cpaVajUF2_2));
	jspl jspl_w_G194_0(.douta(w_G194_0[0]),.doutb(w_G194_0[1]),.din(w_dff_B_4OU2SCCW1_2));
	jspl jspl_w_G197_0(.douta(w_G197_0[0]),.doutb(w_G197_0[1]),.din(w_dff_B_rCprmroI2_2));
	jspl jspl_w_G200_0(.douta(w_G200_0[0]),.doutb(w_G200_0[1]),.din(w_dff_B_NPBlv3NP1_2));
	jspl jspl_w_G203_0(.douta(w_G203_0[0]),.doutb(w_G203_0[1]),.din(w_dff_B_dLHRqh202_2));
	jspl3 jspl3_w_G206_0(.douta(w_dff_A_27FkoB2q8_0),.doutb(w_G206_0[1]),.doutc(w_G206_0[2]),.din(G206));
	jspl3 jspl3_w_G210_0(.douta(w_G210_0[0]),.doutb(w_G210_0[1]),.doutc(w_dff_A_dBgxT8vC6_2),.din(G210));
	jspl3 jspl3_w_G210_1(.douta(w_G210_1[0]),.doutb(w_dff_A_LRGG1Bdy9_1),.doutc(w_G210_1[2]),.din(w_G210_0[0]));
	jspl3 jspl3_w_G210_2(.douta(w_G210_2[0]),.doutb(w_dff_A_oO8qcMEs4_1),.doutc(w_G210_2[2]),.din(w_G210_0[1]));
	jspl3 jspl3_w_G218_0(.douta(w_G218_0[0]),.doutb(w_G218_0[1]),.doutc(w_G218_0[2]),.din(G218));
	jspl3 jspl3_w_G218_1(.douta(w_dff_A_aMxlNGir1_0),.doutb(w_G218_1[1]),.doutc(w_G218_1[2]),.din(w_G218_0[0]));
	jspl3 jspl3_w_G218_2(.douta(w_G218_2[0]),.doutb(w_dff_A_7GTAHaeJ5_1),.doutc(w_G218_2[2]),.din(w_G218_0[1]));
	jspl3 jspl3_w_G226_0(.douta(w_G226_0[0]),.doutb(w_G226_0[1]),.doutc(w_G226_0[2]),.din(G226));
	jspl3 jspl3_w_G226_1(.douta(w_dff_A_DvF0fMCl5_0),.doutb(w_G226_1[1]),.doutc(w_G226_1[2]),.din(w_G226_0[0]));
	jspl3 jspl3_w_G226_2(.douta(w_G226_2[0]),.doutb(w_dff_A_an3LtqQN4_1),.doutc(w_G226_2[2]),.din(w_G226_0[1]));
	jspl3 jspl3_w_G234_0(.douta(w_G234_0[0]),.doutb(w_G234_0[1]),.doutc(w_dff_A_B2BOyBS42_2),.din(G234));
	jspl3 jspl3_w_G234_1(.douta(w_G234_1[0]),.doutb(w_G234_1[1]),.doutc(w_G234_1[2]),.din(w_G234_0[0]));
	jspl jspl_w_G234_2(.douta(w_dff_A_Qzss2TnV3_0),.doutb(w_G234_2[1]),.din(w_G234_0[1]));
	jspl3 jspl3_w_G242_0(.douta(w_G242_0[0]),.doutb(w_dff_A_eq9gA4NK7_1),.doutc(w_dff_A_uf7O1jrH4_2),.din(G242));
	jspl3 jspl3_w_G242_1(.douta(w_dff_A_qoxOJcP88_0),.doutb(w_dff_A_hmdwoiRC5_1),.doutc(w_G242_1[2]),.din(w_G242_0[0]));
	jspl jspl_w_G245_0(.douta(w_G245_0[0]),.doutb(w_G245_0[1]),.din(G245));
	jspl3 jspl3_w_G248_0(.douta(w_G248_0[0]),.doutb(w_G248_0[1]),.doutc(w_G248_0[2]),.din(G248));
	jspl3 jspl3_w_G248_1(.douta(w_G248_1[0]),.doutb(w_G248_1[1]),.doutc(w_G248_1[2]),.din(w_G248_0[0]));
	jspl3 jspl3_w_G248_2(.douta(w_G248_2[0]),.doutb(w_G248_2[1]),.doutc(w_G248_2[2]),.din(w_G248_0[1]));
	jspl3 jspl3_w_G248_3(.douta(w_G248_3[0]),.doutb(w_G248_3[1]),.doutc(w_dff_A_yj6NuqGK2_2),.din(w_G248_0[2]));
	jspl3 jspl3_w_G248_4(.douta(w_G248_4[0]),.doutb(w_G248_4[1]),.doutc(w_G248_4[2]),.din(w_G248_1[0]));
	jspl jspl_w_G248_5(.douta(w_G248_5[0]),.doutb(w_G248_5[1]),.din(w_G248_1[1]));
	jspl3 jspl3_w_G251_0(.douta(w_G251_0[0]),.doutb(w_dff_A_mImFSVqW2_1),.doutc(w_dff_A_GOTqrNDj2_2),.din(G251));
	jspl3 jspl3_w_G251_1(.douta(w_G251_1[0]),.doutb(w_dff_A_A6waiVFy5_1),.doutc(w_dff_A_KqWzSVqx9_2),.din(w_G251_0[0]));
	jspl3 jspl3_w_G251_2(.douta(w_G251_2[0]),.doutb(w_G251_2[1]),.doutc(w_G251_2[2]),.din(w_G251_0[1]));
	jspl3 jspl3_w_G251_3(.douta(w_G251_3[0]),.doutb(w_G251_3[1]),.doutc(w_G251_3[2]),.din(w_G251_0[2]));
	jspl3 jspl3_w_G251_4(.douta(w_G251_4[0]),.doutb(w_dff_A_wyHVClMG1_1),.doutc(w_dff_A_mssGpBpw2_2),.din(w_G251_1[0]));
	jspl3 jspl3_w_G254_0(.douta(w_G254_0[0]),.doutb(w_G254_0[1]),.doutc(w_G254_0[2]),.din(G254));
	jspl3 jspl3_w_G254_1(.douta(w_G254_1[0]),.doutb(w_G254_1[1]),.doutc(w_G254_1[2]),.din(w_G254_0[0]));
	jspl3 jspl3_w_G257_0(.douta(w_G257_0[0]),.doutb(w_G257_0[1]),.doutc(w_G257_0[2]),.din(G257));
	jspl3 jspl3_w_G257_1(.douta(w_dff_A_uLwLcYkQ5_0),.doutb(w_G257_1[1]),.doutc(w_G257_1[2]),.din(w_G257_0[0]));
	jspl3 jspl3_w_G257_2(.douta(w_G257_2[0]),.doutb(w_dff_A_itVy6ivB7_1),.doutc(w_G257_2[2]),.din(w_G257_0[1]));
	jspl3 jspl3_w_G265_0(.douta(w_G265_0[0]),.doutb(w_G265_0[1]),.doutc(w_dff_A_HsHNtB4R8_2),.din(G265));
	jspl3 jspl3_w_G265_1(.douta(w_G265_1[0]),.doutb(w_G265_1[1]),.doutc(w_G265_1[2]),.din(w_G265_0[0]));
	jspl jspl_w_G265_2(.douta(w_dff_A_nh5h3Tpz4_0),.doutb(w_G265_2[1]),.din(w_G265_0[1]));
	jspl3 jspl3_w_G273_0(.douta(w_G273_0[0]),.doutb(w_G273_0[1]),.doutc(w_dff_A_oG5mlAkU3_2),.din(G273));
	jspl3 jspl3_w_G273_1(.douta(w_G273_1[0]),.doutb(w_G273_1[1]),.doutc(w_G273_1[2]),.din(w_G273_0[0]));
	jspl3 jspl3_w_G273_2(.douta(w_G273_2[0]),.doutb(w_dff_A_Fsw5FWWf3_1),.doutc(w_G273_2[2]),.din(w_G273_0[1]));
	jspl jspl_w_G280_0(.douta(w_G280_0[0]),.doutb(w_dff_A_ukhumN2q9_1),.din(G280));
	jspl3 jspl3_w_G281_0(.douta(w_G281_0[0]),.doutb(w_G281_0[1]),.doutc(w_dff_A_92zf0YJc9_2),.din(G281));
	jspl3 jspl3_w_G281_1(.douta(w_G281_1[0]),.doutb(w_G281_1[1]),.doutc(w_G281_1[2]),.din(w_G281_0[0]));
	jspl jspl_w_G281_2(.douta(w_dff_A_x9Mga5Vo5_0),.doutb(w_G281_2[1]),.din(w_G281_0[1]));
	jspl jspl_w_G289_0(.douta(w_dff_A_wLOdru9x4_0),.doutb(w_G289_0[1]),.din(G289));
	jspl3 jspl3_w_G293_0(.douta(w_G293_0[0]),.doutb(w_dff_A_W8Mlyg2V4_1),.doutc(w_G293_0[2]),.din(G293));
	jspl3 jspl3_w_G299_0(.douta(w_G299_0[0]),.doutb(w_G299_0[1]),.doutc(w_G299_0[2]),.din(G299));
	jspl3 jspl3_w_G302_0(.douta(w_dff_A_Jnph24Rg6_0),.doutb(w_dff_A_TNwFbmIf5_1),.doutc(w_G302_0[2]),.din(G302));
	jspl3 jspl3_w_G308_0(.douta(w_G308_0[0]),.doutb(w_G308_0[1]),.doutc(w_G308_0[2]),.din(G308));
	jspl3 jspl3_w_G308_1(.douta(w_dff_A_bZHPyQTY7_0),.doutb(w_G308_1[1]),.doutc(w_G308_1[2]),.din(w_G308_0[0]));
	jspl3 jspl3_w_G316_0(.douta(w_G316_0[0]),.doutb(w_G316_0[1]),.doutc(w_G316_0[2]),.din(G316));
	jspl3 jspl3_w_G316_1(.douta(w_dff_A_0ZhmUMim8_0),.doutb(w_G316_1[1]),.doutc(w_G316_1[2]),.din(w_G316_0[0]));
	jspl3 jspl3_w_G324_0(.douta(w_G324_0[0]),.doutb(w_dff_A_0MXc5Cex0_1),.doutc(w_G324_0[2]),.din(G324));
	jspl3 jspl3_w_G324_1(.douta(w_G324_1[0]),.doutb(w_dff_A_na05WsST4_1),.doutc(w_G324_1[2]),.din(w_G324_0[0]));
	jspl jspl_w_G331_0(.douta(w_G331_0[0]),.doutb(w_dff_A_ad3WK7eX1_1),.din(G331));
	jspl3 jspl3_w_G332_0(.douta(w_G332_0[0]),.doutb(w_G332_0[1]),.doutc(w_G332_0[2]),.din(G332));
	jspl3 jspl3_w_G332_1(.douta(w_G332_1[0]),.doutb(w_G332_1[1]),.doutc(w_dff_A_GdXNJ0p72_2),.din(w_G332_0[0]));
	jspl3 jspl3_w_G332_2(.douta(w_dff_A_C1ZAZGdu3_0),.doutb(w_G332_2[1]),.doutc(w_G332_2[2]),.din(w_G332_0[1]));
	jspl3 jspl3_w_G332_3(.douta(w_dff_A_Qh9JfHui7_0),.doutb(w_G332_3[1]),.doutc(w_dff_A_SQnpHEaN0_2),.din(w_G332_0[2]));
	jspl3 jspl3_w_G332_4(.douta(w_dff_A_XLxZLxTv8_0),.doutb(w_G332_4[1]),.doutc(w_G332_4[2]),.din(w_G332_1[0]));
	jspl3 jspl3_w_G335_0(.douta(w_G335_0[0]),.doutb(w_G335_0[1]),.doutc(w_G335_0[2]),.din(G335));
	jspl3 jspl3_w_G335_1(.douta(w_G335_1[0]),.doutb(w_G335_1[1]),.doutc(w_dff_A_bjbwUG7M0_2),.din(w_G335_0[0]));
	jspl3 jspl3_w_G335_2(.douta(w_G335_2[0]),.doutb(w_G335_2[1]),.doutc(w_G335_2[2]),.din(w_G335_0[1]));
	jspl3 jspl3_w_G335_3(.douta(w_dff_A_Osos0htW4_0),.doutb(w_G335_3[1]),.doutc(w_G335_3[2]),.din(w_G335_0[2]));
	jspl jspl_w_G335_4(.douta(w_dff_A_yd3URyCi7_0),.doutb(w_G335_4[1]),.din(w_G335_1[0]));
	jspl3 jspl3_w_G341_0(.douta(w_G341_0[0]),.doutb(w_G341_0[1]),.doutc(w_dff_A_Yk7dySkI4_2),.din(G341));
	jspl3 jspl3_w_G341_1(.douta(w_G341_1[0]),.doutb(w_G341_1[1]),.doutc(w_G341_1[2]),.din(w_G341_0[0]));
	jspl3 jspl3_w_G341_2(.douta(w_G341_2[0]),.doutb(w_dff_A_S7x97lQ49_1),.doutc(w_G341_2[2]),.din(w_G341_0[1]));
	jspl jspl_w_G348_0(.douta(w_dff_A_mQjqQizc4_0),.doutb(w_G348_0[1]),.din(G348));
	jspl3 jspl3_w_G351_0(.douta(w_G351_0[0]),.doutb(w_G351_0[1]),.doutc(w_G351_0[2]),.din(G351));
	jspl3 jspl3_w_G351_1(.douta(w_dff_A_OGSlSAjg7_0),.doutb(w_G351_1[1]),.doutc(w_G351_1[2]),.din(w_G351_0[0]));
	jspl3 jspl3_w_G351_2(.douta(w_G351_2[0]),.doutb(w_dff_A_5PM0iRLc9_1),.doutc(w_G351_2[2]),.din(w_G351_0[1]));
	jspl jspl_w_G358_0(.douta(w_dff_A_vPdbNkDr1_0),.doutb(w_G358_0[1]),.din(G358));
	jspl3 jspl3_w_G361_0(.douta(w_G361_0[0]),.doutb(w_dff_A_kj64doxa1_1),.doutc(w_G361_0[2]),.din(G361));
	jspl jspl_w_G369_0(.douta(w_dff_A_6gJRWWHu3_0),.doutb(w_G369_0[1]),.din(G369));
	jspl3 jspl3_w_G374_0(.douta(w_dff_A_DU9og2s62_0),.doutb(w_dff_A_IFGuyCP12_1),.doutc(w_G374_0[2]),.din(G374));
	jspl3 jspl3_w_G389_0(.douta(w_dff_A_dVCXe1m09_0),.doutb(w_dff_A_bMCTS3lh5_1),.doutc(w_G389_0[2]),.din(G389));
	jspl3 jspl3_w_G400_0(.douta(w_G400_0[0]),.doutb(w_dff_A_6BxukAJX7_1),.doutc(w_dff_A_2ZmmhUZk7_2),.din(G400));
	jspl jspl_w_G400_1(.douta(w_dff_A_TIbKSzWp7_0),.doutb(w_G400_1[1]),.din(w_G400_0[0]));
	jspl3 jspl3_w_G411_0(.douta(w_dff_A_7sr0iuu30_0),.doutb(w_dff_A_1Hs6LHY27_1),.doutc(w_G411_0[2]),.din(G411));
	jspl3 jspl3_w_G422_0(.douta(w_dff_A_G3VvcAxt0_0),.doutb(w_G422_0[1]),.doutc(w_dff_A_IKwuN2PV3_2),.din(G422));
	jspl3 jspl3_w_G422_1(.douta(w_G422_1[0]),.doutb(w_G422_1[1]),.doutc(w_G422_1[2]),.din(w_G422_0[0]));
	jspl jspl_w_G422_2(.douta(w_dff_A_VqUJsa6V0_0),.doutb(w_G422_2[1]),.din(w_G422_0[1]));
	jspl3 jspl3_w_G435_0(.douta(w_G435_0[0]),.doutb(w_dff_A_35cJy9Fu7_1),.doutc(w_dff_A_bVfatrKy2_2),.din(G435));
	jspl3 jspl3_w_G435_1(.douta(w_dff_A_olwED41o7_0),.doutb(w_dff_A_42D1ZSQZ3_1),.doutc(w_G435_1[2]),.din(w_G435_0[0]));
	jspl3 jspl3_w_G446_0(.douta(w_G446_0[0]),.doutb(w_dff_A_oi8BN86S2_1),.doutc(w_dff_A_kfmutEPO3_2),.din(G446));
	jspl3 jspl3_w_G446_1(.douta(w_dff_A_8flNOkE21_0),.doutb(w_dff_A_iKiEC3sc5_1),.doutc(w_G446_1[2]),.din(w_G446_0[0]));
	jspl3 jspl3_w_G457_0(.douta(w_dff_A_FTBFJaf07_0),.doutb(w_G457_0[1]),.doutc(w_dff_A_XdkzTyra1_2),.din(G457));
	jspl3 jspl3_w_G457_1(.douta(w_G457_1[0]),.doutb(w_G457_1[1]),.doutc(w_G457_1[2]),.din(w_G457_0[0]));
	jspl jspl_w_G457_2(.douta(w_dff_A_UjyjVKCa7_0),.doutb(w_G457_2[1]),.din(w_G457_0[1]));
	jspl3 jspl3_w_G468_0(.douta(w_G468_0[0]),.doutb(w_dff_A_jHQrua3D1_1),.doutc(w_dff_A_Arb3f7to5_2),.din(G468));
	jspl3 jspl3_w_G468_1(.douta(w_dff_A_vXbNci8I3_0),.doutb(w_dff_A_Rwtbp0hX3_1),.doutc(w_G468_1[2]),.din(w_G468_0[0]));
	jspl3 jspl3_w_G479_0(.douta(w_G479_0[0]),.doutb(w_dff_A_fMXpPf7C0_1),.doutc(w_dff_A_0x3qhw4g3_2),.din(G479));
	jspl jspl_w_G479_1(.douta(w_dff_A_gVYY9rGg0_0),.doutb(w_G479_1[1]),.din(w_G479_0[0]));
	jspl3 jspl3_w_G490_0(.douta(w_G490_0[0]),.doutb(w_dff_A_MKWq9gVH1_1),.doutc(w_dff_A_atVKGEcb4_2),.din(G490));
	jspl3 jspl3_w_G490_1(.douta(w_dff_A_DyUcskyR5_0),.doutb(w_dff_A_F0OTlOFe7_1),.doutc(w_G490_1[2]),.din(w_G490_0[0]));
	jspl3 jspl3_w_G503_0(.douta(w_G503_0[0]),.doutb(w_dff_A_2TZ0HTV80_1),.doutc(w_dff_A_QtjbEeNI5_2),.din(G503));
	jspl3 jspl3_w_G503_1(.douta(w_dff_A_FnOpcfzC2_0),.doutb(w_dff_A_yCbNsVp33_1),.doutc(w_G503_1[2]),.din(w_G503_0[0]));
	jspl3 jspl3_w_G514_0(.douta(w_G514_0[0]),.doutb(w_dff_A_TQfhw9Mw6_1),.doutc(w_dff_A_MLS9kANA5_2),.din(G514));
	jspl jspl_w_G514_1(.douta(w_G514_1[0]),.doutb(w_G514_1[1]),.din(w_G514_0[0]));
	jspl3 jspl3_w_G523_0(.douta(w_G523_0[0]),.doutb(w_dff_A_OzvjWbRM9_1),.doutc(w_dff_A_jAj800uz2_2),.din(G523));
	jspl jspl_w_G523_1(.douta(w_dff_A_SM2qFWos7_0),.doutb(w_G523_1[1]),.din(w_G523_0[0]));
	jspl3 jspl3_w_G534_0(.douta(w_G534_0[0]),.doutb(w_dff_A_gVDVdBJY9_1),.doutc(w_dff_A_NIGnlWba9_2),.din(G534));
	jspl3 jspl3_w_G534_1(.douta(w_dff_A_h3pchY909_0),.doutb(w_dff_A_sd7fZ1847_1),.doutc(w_G534_1[2]),.din(w_G534_0[0]));
	jspl3 jspl3_w_G545_0(.douta(w_G545_0[0]),.doutb(w_G545_0[1]),.doutc(w_G545_0[2]),.din(G545));
	jspl3 jspl3_w_G549_0(.douta(w_G549_0[0]),.doutb(w_G549_0[1]),.doutc(w_G549_0[2]),.din(G549));
	jspl jspl_w_G552_0(.douta(w_G552_0[0]),.doutb(w_G552_0[1]),.din(G552));
	jspl jspl_w_G559_0(.douta(w_G559_0[0]),.doutb(w_G559_0[1]),.din(G559));
	jspl jspl_w_G562_0(.douta(w_G562_0[0]),.doutb(w_G562_0[1]),.din(G562));
	jspl3 jspl3_w_G1497_0(.douta(w_dff_A_kdJh28BH4_0),.doutb(w_G1497_0[1]),.doutc(w_dff_A_G5zBqwwm1_2),.din(G1497));
	jspl3 jspl3_w_G1689_0(.douta(w_G1689_0[0]),.doutb(w_G1689_0[1]),.doutc(w_dff_A_URGcx6v34_2),.din(G1689));
	jspl3 jspl3_w_G1690_0(.douta(w_G1690_0[0]),.doutb(w_dff_A_qzXADXbr4_1),.doutc(w_G1690_0[2]),.din(G1690));
	jspl3 jspl3_w_G1691_0(.douta(w_G1691_0[0]),.doutb(w_G1691_0[1]),.doutc(w_dff_A_YqYBMRA82_2),.din(G1691));
	jspl3 jspl3_w_G1694_0(.douta(w_G1694_0[0]),.doutb(w_dff_A_RoRRi9D51_1),.doutc(w_G1694_0[2]),.din(G1694));
	jspl3 jspl3_w_G2174_0(.douta(w_dff_A_STo9Voqn1_0),.doutb(w_G2174_0[1]),.doutc(w_dff_A_AAsaCbbk5_2),.din(G2174));
	jspl3 jspl3_w_G2358_0(.douta(w_G2358_0[0]),.doutb(w_G2358_0[1]),.doutc(w_G2358_0[2]),.din(G2358));
	jspl3 jspl3_w_G2358_1(.douta(w_G2358_1[0]),.doutb(w_G2358_1[1]),.doutc(w_G2358_1[2]),.din(w_G2358_0[0]));
	jspl3 jspl3_w_G2358_2(.douta(w_dff_A_UZf91e0e1_0),.doutb(w_dff_A_kvAw0xGb1_1),.doutc(w_G2358_2[2]),.din(w_G2358_0[1]));
	jspl jspl_w_G3173_0(.douta(w_G3173_0[0]),.doutb(w_G3173_0[1]),.din(G3173));
	jspl3 jspl3_w_G3546_0(.douta(w_G3546_0[0]),.doutb(w_G3546_0[1]),.doutc(w_G3546_0[2]),.din(G3546));
	jspl3 jspl3_w_G3546_1(.douta(w_G3546_1[0]),.doutb(w_G3546_1[1]),.doutc(w_G3546_1[2]),.din(w_G3546_0[0]));
	jspl3 jspl3_w_G3546_2(.douta(w_G3546_2[0]),.doutb(w_G3546_2[1]),.doutc(w_G3546_2[2]),.din(w_G3546_0[1]));
	jspl3 jspl3_w_G3546_3(.douta(w_G3546_3[0]),.doutb(w_G3546_3[1]),.doutc(w_G3546_3[2]),.din(w_G3546_0[2]));
	jspl3 jspl3_w_G3546_4(.douta(w_G3546_4[0]),.doutb(w_G3546_4[1]),.doutc(w_G3546_4[2]),.din(w_G3546_1[0]));
	jspl jspl_w_G3546_5(.douta(w_G3546_5[0]),.doutb(w_G3546_5[1]),.din(w_G3546_1[1]));
	jspl3 jspl3_w_G3548_0(.douta(w_G3548_0[0]),.doutb(w_G3548_0[1]),.doutc(w_G3548_0[2]),.din(w_dff_B_slQjwQXb7_3));
	jspl3 jspl3_w_G3548_1(.douta(w_G3548_1[0]),.doutb(w_G3548_1[1]),.doutc(w_G3548_1[2]),.din(w_G3548_0[0]));
	jspl3 jspl3_w_G3548_2(.douta(w_G3548_2[0]),.doutb(w_G3548_2[1]),.doutc(w_G3548_2[2]),.din(w_G3548_0[1]));
	jspl3 jspl3_w_G3548_3(.douta(w_G3548_3[0]),.doutb(w_G3548_3[1]),.doutc(w_G3548_3[2]),.din(w_G3548_0[2]));
	jspl3 jspl3_w_G3548_4(.douta(w_G3548_4[0]),.doutb(w_G3548_4[1]),.doutc(w_G3548_4[2]),.din(w_G3548_1[0]));
	jspl jspl_w_G3552_0(.douta(w_G3552_0[0]),.doutb(w_G3552_0[1]),.din(G3552));
	jspl jspl_w_G3717_0(.douta(w_dff_A_FvB3tIyx2_0),.doutb(w_G3717_0[1]),.din(G3717));
	jspl3 jspl3_w_G3724_0(.douta(w_dff_A_629NqC8a0_0),.doutb(w_G3724_0[1]),.doutc(w_dff_A_YCUoHJmc3_2),.din(G3724));
	jspl3 jspl3_w_G4087_0(.douta(w_G4087_0[0]),.doutb(w_dff_A_PjTDWTfI7_1),.doutc(w_G4087_0[2]),.din(G4087));
	jspl3 jspl3_w_G4088_0(.douta(w_G4088_0[0]),.doutb(w_G4088_0[1]),.doutc(w_dff_A_D88n27GW8_2),.din(G4088));
	jspl3 jspl3_w_G4089_0(.douta(w_G4089_0[0]),.doutb(w_G4089_0[1]),.doutc(w_dff_A_CfNDWJtS0_2),.din(G4089));
	jspl3 jspl3_w_G4090_0(.douta(w_G4090_0[0]),.doutb(w_dff_A_oD4ZL31J1_1),.doutc(w_G4090_0[2]),.din(G4090));
	jspl3 jspl3_w_G4091_0(.douta(w_G4091_0[0]),.doutb(w_G4091_0[1]),.doutc(w_dff_A_LQkLYlbU9_2),.din(G4091));
	jspl3 jspl3_w_G4091_1(.douta(w_G4091_1[0]),.doutb(w_dff_A_GsGWKxYK5_1),.doutc(w_dff_A_thHBqV6D1_2),.din(w_G4091_0[0]));
	jspl3 jspl3_w_G4091_2(.douta(w_G4091_2[0]),.doutb(w_G4091_2[1]),.doutc(w_dff_A_vKBiK2D37_2),.din(w_G4091_0[1]));
	jspl3 jspl3_w_G4092_0(.douta(w_G4092_0[0]),.doutb(w_G4092_0[1]),.doutc(w_G4092_0[2]),.din(G4092));
	jspl3 jspl3_w_G4092_1(.douta(w_dff_A_Tka5TvuH0_0),.doutb(w_dff_A_rRft9HIC6_1),.doutc(w_G4092_1[2]),.din(w_G4092_0[0]));
	jspl jspl_w_G599_0(.douta(w_G599_0),.doutb(G599),.din(G599_fa_));
	jspl jspl_w_G600_0(.douta(w_G600_0),.doutb(G600),.din(G600_fa_));
	jspl jspl_w_G601_0(.douta(w_dff_A_OpW0ntUi9_0),.doutb(G601),.din(G601_fa_));
	jspl jspl_w_G611_0(.douta(w_G611_0),.doutb(G611),.din(G611_fa_));
	jspl jspl_w_G612_0(.douta(w_G612_0),.doutb(G612),.din(G612_fa_));
	jspl3 jspl3_w_G809_0(.douta(w_G809_0[0]),.doutb(w_G809_0[1]),.doutc(w_G809_0[2]),.din(G809_fa_));
	jspl3 jspl3_w_G809_1(.douta(w_G809_1[0]),.doutb(w_G809_1[1]),.doutc(w_G809_1[2]),.din(w_G809_0[0]));
	jspl3 jspl3_w_G809_2(.douta(w_G809_2[0]),.doutb(w_G809_2[1]),.doutc(w_dff_A_YBhqqeWI3_2),.din(w_G809_0[1]));
	jspl3 jspl3_w_G809_3(.douta(w_dff_A_BFIIhYPO2_0),.doutb(w_G809_3[1]),.doutc(G809),.din(w_G809_0[2]));
	jspl jspl_w_G593_0(.douta(w_G593_0),.doutb(G593),.din(G593_fa_));
	jspl jspl_w_G822_0(.douta(w_G822_0),.doutb(G822),.din(G822_fa_));
	jspl jspl_w_G838_0(.douta(w_G838_0),.doutb(G838),.din(G838_fa_));
	jspl jspl_w_G861_0(.douta(w_G861_0),.doutb(G861),.din(G861_fa_));
	jspl jspl_w_G832_0(.douta(w_G832_0),.doutb(G832),.din(G832_fa_));
	jspl jspl_w_G834_0(.douta(w_G834_0),.doutb(G834),.din(G834_fa_));
	jspl jspl_w_G836_0(.douta(w_G836_0),.doutb(G836),.din(G836_fa_));
	jspl jspl_w_G871_0(.douta(w_G871_0),.doutb(G871),.din(G871_fa_));
	jspl jspl_w_G873_0(.douta(w_G873_0),.doutb(G873),.din(G873_fa_));
	jspl jspl_w_G875_0(.douta(w_G875_0),.doutb(G875),.din(G875_fa_));
	jspl jspl_w_G877_0(.douta(w_G877_0),.doutb(G877),.din(G877_fa_));
	jspl jspl_w_G1000_0(.douta(w_G1000_0),.doutb(G1000),.din(G1000_fa_));
	jspl jspl_w_G826_0(.douta(w_G826_0),.doutb(G826),.din(G826_fa_));
	jspl jspl_w_G828_0(.douta(w_G828_0),.doutb(G828),.din(G828_fa_));
	jspl jspl_w_G830_0(.douta(w_G830_0),.doutb(G830),.din(G830_fa_));
	jspl jspl_w_G867_0(.douta(w_G867_0),.doutb(G867),.din(G867_fa_));
	jspl jspl_w_G869_0(.douta(w_G869_0),.doutb(G869),.din(G869_fa_));
	jspl jspl_w_n316_0(.douta(w_n316_0[0]),.doutb(w_n316_0[1]),.din(n316));
	jspl jspl_w_n318_0(.douta(w_n318_0[0]),.doutb(w_n318_0[1]),.din(n318));
	jspl3 jspl3_w_n326_0(.douta(w_n326_0[0]),.doutb(w_n326_0[1]),.doutc(w_n326_0[2]),.din(n326));
	jspl3 jspl3_w_n326_1(.douta(w_n326_1[0]),.doutb(w_n326_1[1]),.doutc(w_n326_1[2]),.din(w_n326_0[0]));
	jspl jspl_w_n326_2(.douta(w_n326_2[0]),.doutb(w_n326_2[1]),.din(w_n326_0[1]));
	jspl jspl_w_n333_0(.douta(w_n333_0[0]),.doutb(w_n333_0[1]),.din(n333));
	jspl jspl_w_n336_0(.douta(w_n336_0[0]),.doutb(w_n336_0[1]),.din(n336));
	jspl jspl_w_n360_0(.douta(w_n360_0[0]),.doutb(w_n360_0[1]),.din(n360));
	jspl jspl_w_n362_0(.douta(w_dff_A_d5VI5gxX9_0),.doutb(w_n362_0[1]),.din(n362));
	jspl3 jspl3_w_n366_0(.douta(w_n366_0[0]),.doutb(w_n366_0[1]),.doutc(w_n366_0[2]),.din(n366));
	jspl3 jspl3_w_n366_1(.douta(w_n366_1[0]),.doutb(w_n366_1[1]),.doutc(w_n366_1[2]),.din(w_n366_0[0]));
	jspl3 jspl3_w_n366_2(.douta(w_n366_2[0]),.doutb(w_n366_2[1]),.doutc(w_n366_2[2]),.din(w_n366_0[1]));
	jspl3 jspl3_w_n366_3(.douta(w_n366_3[0]),.doutb(w_n366_3[1]),.doutc(w_n366_3[2]),.din(w_n366_0[2]));
	jspl3 jspl3_w_n366_4(.douta(w_n366_4[0]),.doutb(w_n366_4[1]),.doutc(w_n366_4[2]),.din(w_n366_1[0]));
	jspl3 jspl3_w_n368_0(.douta(w_n368_0[0]),.doutb(w_n368_0[1]),.doutc(w_n368_0[2]),.din(n368));
	jspl3 jspl3_w_n368_1(.douta(w_n368_1[0]),.doutb(w_n368_1[1]),.doutc(w_n368_1[2]),.din(w_n368_0[0]));
	jspl3 jspl3_w_n368_2(.douta(w_n368_2[0]),.doutb(w_n368_2[1]),.doutc(w_n368_2[2]),.din(w_n368_0[1]));
	jspl3 jspl3_w_n368_3(.douta(w_n368_3[0]),.doutb(w_n368_3[1]),.doutc(w_n368_3[2]),.din(w_n368_0[2]));
	jspl3 jspl3_w_n368_4(.douta(w_n368_4[0]),.doutb(w_n368_4[1]),.doutc(w_n368_4[2]),.din(w_n368_1[0]));
	jspl jspl_w_n368_5(.douta(w_n368_5[0]),.doutb(w_n368_5[1]),.din(w_n368_1[1]));
	jspl3 jspl3_w_n372_0(.douta(w_n372_0[0]),.doutb(w_n372_0[1]),.doutc(w_n372_0[2]),.din(n372));
	jspl jspl_w_n373_0(.douta(w_n373_0[0]),.doutb(w_n373_0[1]),.din(n373));
	jspl3 jspl3_w_n383_0(.douta(w_n383_0[0]),.doutb(w_n383_0[1]),.doutc(w_n383_0[2]),.din(n383));
	jspl3 jspl3_w_n385_0(.douta(w_n385_0[0]),.doutb(w_n385_0[1]),.doutc(w_n385_0[2]),.din(n385));
	jspl3 jspl3_w_n385_1(.douta(w_n385_1[0]),.doutb(w_n385_1[1]),.doutc(w_n385_1[2]),.din(w_n385_0[0]));
	jspl3 jspl3_w_n386_0(.douta(w_n386_0[0]),.doutb(w_n386_0[1]),.doutc(w_n386_0[2]),.din(n386));
	jspl3 jspl3_w_n386_1(.douta(w_n386_1[0]),.doutb(w_n386_1[1]),.doutc(w_n386_1[2]),.din(w_n386_0[0]));
	jspl3 jspl3_w_n386_2(.douta(w_n386_2[0]),.doutb(w_n386_2[1]),.doutc(w_n386_2[2]),.din(w_n386_0[1]));
	jspl3 jspl3_w_n386_3(.douta(w_n386_3[0]),.doutb(w_n386_3[1]),.doutc(w_n386_3[2]),.din(w_n386_0[2]));
	jspl3 jspl3_w_n386_4(.douta(w_n386_4[0]),.doutb(w_n386_4[1]),.doutc(w_n386_4[2]),.din(w_n386_1[0]));
	jspl3 jspl3_w_n388_0(.douta(w_dff_A_gxRtB9es3_0),.doutb(w_n388_0[1]),.doutc(w_dff_A_cLtBuRqT4_2),.din(n388));
	jspl3 jspl3_w_n388_1(.douta(w_n388_1[0]),.doutb(w_n388_1[1]),.doutc(w_n388_1[2]),.din(w_n388_0[0]));
	jspl3 jspl3_w_n389_0(.douta(w_n389_0[0]),.doutb(w_n389_0[1]),.doutc(w_n389_0[2]),.din(n389));
	jspl3 jspl3_w_n389_1(.douta(w_n389_1[0]),.doutb(w_n389_1[1]),.doutc(w_n389_1[2]),.din(w_n389_0[0]));
	jspl3 jspl3_w_n389_2(.douta(w_n389_2[0]),.doutb(w_n389_2[1]),.doutc(w_n389_2[2]),.din(w_n389_0[1]));
	jspl3 jspl3_w_n389_3(.douta(w_n389_3[0]),.doutb(w_n389_3[1]),.doutc(w_n389_3[2]),.din(w_n389_0[2]));
	jspl3 jspl3_w_n389_4(.douta(w_n389_4[0]),.doutb(w_n389_4[1]),.doutc(w_n389_4[2]),.din(w_n389_1[0]));
	jspl jspl_w_n397_0(.douta(w_n397_0[0]),.doutb(w_dff_A_dMEordML7_1),.din(n397));
	jspl3 jspl3_w_n398_0(.douta(w_n398_0[0]),.doutb(w_n398_0[1]),.doutc(w_n398_0[2]),.din(n398));
	jspl3 jspl3_w_n401_0(.douta(w_dff_A_5kixj4V24_0),.doutb(w_n401_0[1]),.doutc(w_dff_A_XsN8yS8u2_2),.din(n401));
	jspl3 jspl3_w_n402_0(.douta(w_n402_0[0]),.doutb(w_n402_0[1]),.doutc(w_n402_0[2]),.din(n402));
	jspl3 jspl3_w_n402_1(.douta(w_n402_1[0]),.doutb(w_n402_1[1]),.doutc(w_n402_1[2]),.din(w_n402_0[0]));
	jspl jspl_w_n402_2(.douta(w_n402_2[0]),.doutb(w_n402_2[1]),.din(w_n402_0[1]));
	jspl jspl_w_n403_0(.douta(w_n403_0[0]),.doutb(w_n403_0[1]),.din(n403));
	jspl3 jspl3_w_n405_0(.douta(w_n405_0[0]),.doutb(w_n405_0[1]),.doutc(w_n405_0[2]),.din(n405));
	jspl3 jspl3_w_n405_1(.douta(w_n405_1[0]),.doutb(w_n405_1[1]),.doutc(w_n405_1[2]),.din(w_n405_0[0]));
	jspl jspl_w_n405_2(.douta(w_n405_2[0]),.doutb(w_n405_2[1]),.din(w_n405_0[1]));
	jspl jspl_w_n407_0(.douta(w_n407_0[0]),.doutb(w_n407_0[1]),.din(n407));
	jspl jspl_w_n408_0(.douta(w_n408_0[0]),.doutb(w_n408_0[1]),.din(n408));
	jspl3 jspl3_w_n410_0(.douta(w_n410_0[0]),.doutb(w_n410_0[1]),.doutc(w_dff_A_AnvJjx9h2_2),.din(n410));
	jspl jspl_w_n410_1(.douta(w_dff_A_GJhqp7rA4_0),.doutb(w_n410_1[1]),.din(w_n410_0[0]));
	jspl jspl_w_n414_0(.douta(w_n414_0[0]),.doutb(w_n414_0[1]),.din(n414));
	jspl jspl_w_n416_0(.douta(w_n416_0[0]),.doutb(w_n416_0[1]),.din(n416));
	jspl3 jspl3_w_n419_0(.douta(w_n419_0[0]),.doutb(w_n419_0[1]),.doutc(w_n419_0[2]),.din(n419));
	jspl3 jspl3_w_n424_0(.douta(w_n424_0[0]),.doutb(w_n424_0[1]),.doutc(w_n424_0[2]),.din(n424));
	jspl3 jspl3_w_n424_1(.douta(w_n424_1[0]),.doutb(w_n424_1[1]),.doutc(w_n424_1[2]),.din(w_n424_0[0]));
	jspl jspl_w_n424_2(.douta(w_n424_2[0]),.doutb(w_n424_2[1]),.din(w_n424_0[1]));
	jspl jspl_w_n426_0(.douta(w_n426_0[0]),.doutb(w_dff_A_CDFLFID79_1),.din(n426));
	jspl jspl_w_n434_0(.douta(w_n434_0[0]),.doutb(w_n434_0[1]),.din(n434));
	jspl3 jspl3_w_n435_0(.douta(w_n435_0[0]),.doutb(w_n435_0[1]),.doutc(w_n435_0[2]),.din(n435));
	jspl3 jspl3_w_n435_1(.douta(w_n435_1[0]),.doutb(w_n435_1[1]),.doutc(w_n435_1[2]),.din(w_n435_0[0]));
	jspl3 jspl3_w_n437_0(.douta(w_dff_A_6dzRm1Bg9_0),.doutb(w_n437_0[1]),.doutc(w_dff_A_fDbBMFjd2_2),.din(n437));
	jspl3 jspl3_w_n437_1(.douta(w_n437_1[0]),.doutb(w_n437_1[1]),.doutc(w_n437_1[2]),.din(w_n437_0[0]));
	jspl jspl_w_n445_0(.douta(w_n445_0[0]),.doutb(w_n445_0[1]),.din(n445));
	jspl3 jspl3_w_n449_0(.douta(w_n449_0[0]),.doutb(w_n449_0[1]),.doutc(w_n449_0[2]),.din(n449));
	jspl3 jspl3_w_n449_1(.douta(w_n449_1[0]),.doutb(w_n449_1[1]),.doutc(w_n449_1[2]),.din(w_n449_0[0]));
	jspl3 jspl3_w_n451_0(.douta(w_dff_A_aX7Q3r0A3_0),.doutb(w_n451_0[1]),.doutc(w_dff_A_SIaOqvhL3_2),.din(n451));
	jspl jspl_w_n451_1(.douta(w_n451_1[0]),.doutb(w_n451_1[1]),.din(w_n451_0[0]));
	jspl jspl_w_n459_0(.douta(w_n459_0[0]),.doutb(w_dff_A_eGdNV9IC6_1),.din(n459));
	jspl3 jspl3_w_n460_0(.douta(w_n460_0[0]),.doutb(w_n460_0[1]),.doutc(w_n460_0[2]),.din(n460));
	jspl3 jspl3_w_n460_1(.douta(w_n460_1[0]),.doutb(w_n460_1[1]),.doutc(w_n460_1[2]),.din(w_n460_0[0]));
	jspl3 jspl3_w_n462_0(.douta(w_n462_0[0]),.doutb(w_dff_A_cXlOgeUS3_1),.doutc(w_dff_A_tzs6aVif1_2),.din(n462));
	jspl jspl_w_n470_0(.douta(w_n470_0[0]),.doutb(w_n470_0[1]),.din(n470));
	jspl3 jspl3_w_n471_0(.douta(w_n471_0[0]),.doutb(w_n471_0[1]),.doutc(w_n471_0[2]),.din(n471));
	jspl jspl_w_n471_1(.douta(w_n471_1[0]),.doutb(w_n471_1[1]),.din(w_n471_0[0]));
	jspl3 jspl3_w_n473_0(.douta(w_dff_A_hd0J9uOv7_0),.doutb(w_n473_0[1]),.doutc(w_dff_A_Cds4j2RZ3_2),.din(n473));
	jspl3 jspl3_w_n473_1(.douta(w_dff_A_p4y39Lw87_0),.doutb(w_n473_1[1]),.doutc(w_n473_1[2]),.din(w_n473_0[0]));
	jspl jspl_w_n481_0(.douta(w_n481_0[0]),.doutb(w_n481_0[1]),.din(n481));
	jspl3 jspl3_w_n484_0(.douta(w_n484_0[0]),.doutb(w_n484_0[1]),.doutc(w_n484_0[2]),.din(n484));
	jspl jspl_w_n484_1(.douta(w_n484_1[0]),.doutb(w_n484_1[1]),.din(w_n484_0[0]));
	jspl3 jspl3_w_n486_0(.douta(w_dff_A_LAvEutKN7_0),.doutb(w_n486_0[1]),.doutc(w_dff_A_t4Wy8jsh4_2),.din(n486));
	jspl jspl_w_n486_1(.douta(w_n486_1[0]),.doutb(w_n486_1[1]),.din(w_n486_0[0]));
	jspl jspl_w_n494_0(.douta(w_n494_0[0]),.doutb(w_n494_0[1]),.din(n494));
	jspl3 jspl3_w_n495_0(.douta(w_n495_0[0]),.doutb(w_n495_0[1]),.doutc(w_n495_0[2]),.din(n495));
	jspl3 jspl3_w_n495_1(.douta(w_n495_1[0]),.doutb(w_n495_1[1]),.doutc(w_n495_1[2]),.din(w_n495_0[0]));
	jspl3 jspl3_w_n497_0(.douta(w_dff_A_Gyr6Xdi39_0),.doutb(w_n497_0[1]),.doutc(w_dff_A_rUqn3KEZ1_2),.din(n497));
	jspl jspl_w_n497_1(.douta(w_n497_1[0]),.doutb(w_n497_1[1]),.din(w_n497_0[0]));
	jspl jspl_w_n505_0(.douta(w_n505_0[0]),.doutb(w_n505_0[1]),.din(n505));
	jspl3 jspl3_w_n507_0(.douta(w_n507_0[0]),.doutb(w_n507_0[1]),.doutc(w_n507_0[2]),.din(n507));
	jspl jspl_w_n507_1(.douta(w_n507_1[0]),.doutb(w_n507_1[1]),.din(w_n507_0[0]));
	jspl jspl_w_n509_0(.douta(w_n509_0[0]),.doutb(w_dff_A_kGhS7hCR3_1),.din(n509));
	jspl jspl_w_n517_0(.douta(w_n517_0[0]),.doutb(w_n517_0[1]),.din(n517));
	jspl3 jspl3_w_n518_0(.douta(w_n518_0[0]),.doutb(w_n518_0[1]),.doutc(w_n518_0[2]),.din(n518));
	jspl jspl_w_n518_1(.douta(w_n518_1[0]),.doutb(w_n518_1[1]),.din(w_n518_0[0]));
	jspl3 jspl3_w_n528_0(.douta(w_n528_0[0]),.doutb(w_n528_0[1]),.doutc(w_n528_0[2]),.din(n528));
	jspl3 jspl3_w_n530_0(.douta(w_n530_0[0]),.doutb(w_n530_0[1]),.doutc(w_n530_0[2]),.din(n530));
	jspl jspl_w_n530_1(.douta(w_n530_1[0]),.doutb(w_n530_1[1]),.din(w_n530_0[0]));
	jspl jspl_w_n532_0(.douta(w_n532_0[0]),.doutb(w_dff_A_5h5lW8da8_1),.din(n532));
	jspl jspl_w_n540_0(.douta(w_n540_0[0]),.doutb(w_n540_0[1]),.din(n540));
	jspl3 jspl3_w_n541_0(.douta(w_n541_0[0]),.doutb(w_n541_0[1]),.doutc(w_n541_0[2]),.din(n541));
	jspl jspl_w_n541_1(.douta(w_n541_1[0]),.doutb(w_n541_1[1]),.din(w_n541_0[0]));
	jspl jspl_w_n543_0(.douta(w_n543_0[0]),.doutb(w_dff_A_rQBGozHr8_1),.din(n543));
	jspl jspl_w_n551_0(.douta(w_n551_0[0]),.doutb(w_n551_0[1]),.din(n551));
	jspl3 jspl3_w_n556_0(.douta(w_n556_0[0]),.doutb(w_n556_0[1]),.doutc(w_n556_0[2]),.din(n556));
	jspl3 jspl3_w_n556_1(.douta(w_n556_1[0]),.doutb(w_n556_1[1]),.doutc(w_n556_1[2]),.din(w_n556_0[0]));
	jspl3 jspl3_w_n556_2(.douta(w_n556_2[0]),.doutb(w_n556_2[1]),.doutc(w_n556_2[2]),.din(w_n556_0[1]));
	jspl3 jspl3_w_n556_3(.douta(w_n556_3[0]),.doutb(w_n556_3[1]),.doutc(w_n556_3[2]),.din(w_n556_0[2]));
	jspl3 jspl3_w_n556_4(.douta(w_n556_4[0]),.doutb(w_n556_4[1]),.doutc(w_n556_4[2]),.din(w_n556_1[0]));
	jspl jspl_w_n556_5(.douta(w_n556_5[0]),.doutb(w_n556_5[1]),.din(w_n556_1[1]));
	jspl3 jspl3_w_n560_0(.douta(w_n560_0[0]),.doutb(w_n560_0[1]),.doutc(w_n560_0[2]),.din(n560));
	jspl jspl_w_n560_1(.douta(w_n560_1[0]),.doutb(w_n560_1[1]),.din(w_n560_0[0]));
	jspl3 jspl3_w_n561_0(.douta(w_n561_0[0]),.doutb(w_dff_A_khti5bYU3_1),.doutc(w_n561_0[2]),.din(n561));
	jspl jspl_w_n562_0(.douta(w_dff_A_Z9CoqXJ94_0),.doutb(w_n562_0[1]),.din(n562));
	jspl3 jspl3_w_n566_0(.douta(w_n566_0[0]),.doutb(w_n566_0[1]),.doutc(w_n566_0[2]),.din(n566));
	jspl3 jspl3_w_n567_0(.douta(w_n567_0[0]),.doutb(w_n567_0[1]),.doutc(w_n567_0[2]),.din(n567));
	jspl jspl_w_n567_1(.douta(w_n567_1[0]),.doutb(w_dff_A_O923MLma9_1),.din(w_n567_0[0]));
	jspl jspl_w_n569_0(.douta(w_n569_0[0]),.doutb(w_dff_A_p5UUECnV1_1),.din(n569));
	jspl jspl_w_n570_0(.douta(w_n570_0[0]),.doutb(w_n570_0[1]),.din(n570));
	jspl3 jspl3_w_n571_0(.douta(w_n571_0[0]),.doutb(w_n571_0[1]),.doutc(w_dff_A_TzhCfWqV9_2),.din(n571));
	jspl jspl_w_n571_1(.douta(w_n571_1[0]),.doutb(w_n571_1[1]),.din(w_n571_0[0]));
	jspl3 jspl3_w_n572_0(.douta(w_dff_A_jG3uHNL70_0),.doutb(w_n572_0[1]),.doutc(w_n572_0[2]),.din(n572));
	jspl3 jspl3_w_n574_0(.douta(w_n574_0[0]),.doutb(w_n574_0[1]),.doutc(w_n574_0[2]),.din(n574));
	jspl3 jspl3_w_n577_0(.douta(w_n577_0[0]),.doutb(w_n577_0[1]),.doutc(w_n577_0[2]),.din(n577));
	jspl3 jspl3_w_n578_0(.douta(w_n578_0[0]),.doutb(w_dff_A_Vqq2KzBu3_1),.doutc(w_n578_0[2]),.din(n578));
	jspl3 jspl3_w_n582_0(.douta(w_n582_0[0]),.doutb(w_n582_0[1]),.doutc(w_n582_0[2]),.din(n582));
	jspl jspl_w_n582_1(.douta(w_n582_1[0]),.doutb(w_n582_1[1]),.din(w_n582_0[0]));
	jspl3 jspl3_w_n583_0(.douta(w_n583_0[0]),.doutb(w_n583_0[1]),.doutc(w_dff_A_Yf2qE8Lp4_2),.din(n583));
	jspl jspl_w_n583_1(.douta(w_dff_A_f2LfcUUq5_0),.doutb(w_n583_1[1]),.din(w_n583_0[0]));
	jspl jspl_w_n585_0(.douta(w_n585_0[0]),.doutb(w_n585_0[1]),.din(n585));
	jspl3 jspl3_w_n587_0(.douta(w_n587_0[0]),.doutb(w_n587_0[1]),.doutc(w_n587_0[2]),.din(n587));
	jspl jspl_w_n587_1(.douta(w_n587_1[0]),.doutb(w_n587_1[1]),.din(w_n587_0[0]));
	jspl3 jspl3_w_n590_0(.douta(w_n590_0[0]),.doutb(w_dff_A_zWJzag0i3_1),.doutc(w_n590_0[2]),.din(n590));
	jspl jspl_w_n590_1(.douta(w_n590_1[0]),.doutb(w_n590_1[1]),.din(w_n590_0[0]));
	jspl jspl_w_n591_0(.douta(w_n591_0[0]),.doutb(w_dff_A_ivFqTZDA0_1),.din(n591));
	jspl3 jspl3_w_n595_0(.douta(w_n595_0[0]),.doutb(w_n595_0[1]),.doutc(w_n595_0[2]),.din(n595));
	jspl jspl_w_n595_1(.douta(w_n595_1[0]),.doutb(w_n595_1[1]),.din(w_n595_0[0]));
	jspl3 jspl3_w_n596_0(.douta(w_dff_A_Vrj1WP1J8_0),.doutb(w_n596_0[1]),.doutc(w_n596_0[2]),.din(n596));
	jspl3 jspl3_w_n600_0(.douta(w_n600_0[0]),.doutb(w_n600_0[1]),.doutc(w_n600_0[2]),.din(n600));
	jspl jspl_w_n600_1(.douta(w_n600_1[0]),.doutb(w_n600_1[1]),.din(w_n600_0[0]));
	jspl jspl_w_n601_0(.douta(w_n601_0[0]),.doutb(w_n601_0[1]),.din(n601));
	jspl3 jspl3_w_n604_0(.douta(w_dff_A_X9guJ0Ki5_0),.doutb(w_n604_0[1]),.doutc(w_n604_0[2]),.din(n604));
	jspl3 jspl3_w_n605_0(.douta(w_n605_0[0]),.doutb(w_n605_0[1]),.doutc(w_n605_0[2]),.din(n605));
	jspl3 jspl3_w_n605_1(.douta(w_n605_1[0]),.doutb(w_n605_1[1]),.doutc(w_dff_A_GhjW42Og9_2),.din(w_n605_0[0]));
	jspl3 jspl3_w_n605_2(.douta(w_n605_2[0]),.doutb(w_n605_2[1]),.doutc(w_n605_2[2]),.din(w_n605_0[1]));
	jspl3 jspl3_w_n607_0(.douta(w_n607_0[0]),.doutb(w_dff_A_Y58LOX3i0_1),.doutc(w_n607_0[2]),.din(n607));
	jspl3 jspl3_w_n609_0(.douta(w_n609_0[0]),.doutb(w_n609_0[1]),.doutc(w_n609_0[2]),.din(n609));
	jspl3 jspl3_w_n609_1(.douta(w_n609_1[0]),.doutb(w_n609_1[1]),.doutc(w_n609_1[2]),.din(w_n609_0[0]));
	jspl3 jspl3_w_n609_2(.douta(w_n609_2[0]),.doutb(w_n609_2[1]),.doutc(w_n609_2[2]),.din(w_n609_0[1]));
	jspl3 jspl3_w_n609_3(.douta(w_n609_3[0]),.doutb(w_n609_3[1]),.doutc(w_n609_3[2]),.din(w_n609_0[2]));
	jspl3 jspl3_w_n609_4(.douta(w_n609_4[0]),.doutb(w_n609_4[1]),.doutc(w_n609_4[2]),.din(w_n609_1[0]));
	jspl3 jspl3_w_n609_5(.douta(w_n609_5[0]),.doutb(w_n609_5[1]),.doutc(w_n609_5[2]),.din(w_n609_1[1]));
	jspl3 jspl3_w_n613_0(.douta(w_n613_0[0]),.doutb(w_n613_0[1]),.doutc(w_n613_0[2]),.din(n613));
	jspl3 jspl3_w_n614_0(.douta(w_n614_0[0]),.doutb(w_n614_0[1]),.doutc(w_n614_0[2]),.din(n614));
	jspl3 jspl3_w_n614_1(.douta(w_dff_A_BQYkyJkX0_0),.doutb(w_n614_1[1]),.doutc(w_dff_A_M91kGm5M5_2),.din(w_n614_0[0]));
	jspl jspl_w_n614_2(.douta(w_dff_A_BNmdF2OE6_0),.doutb(w_n614_2[1]),.din(w_n614_0[1]));
	jspl3 jspl3_w_n617_0(.douta(w_n617_0[0]),.doutb(w_n617_0[1]),.doutc(w_n617_0[2]),.din(n617));
	jspl jspl_w_n617_1(.douta(w_n617_1[0]),.doutb(w_n617_1[1]),.din(w_n617_0[0]));
	jspl3 jspl3_w_n618_0(.douta(w_n618_0[0]),.doutb(w_n618_0[1]),.doutc(w_n618_0[2]),.din(n618));
	jspl jspl_w_n618_1(.douta(w_n618_1[0]),.doutb(w_n618_1[1]),.din(w_n618_0[0]));
	jspl3 jspl3_w_n621_0(.douta(w_n621_0[0]),.doutb(w_n621_0[1]),.doutc(w_n621_0[2]),.din(n621));
	jspl3 jspl3_w_n621_1(.douta(w_dff_A_ZzUXv6Dg6_0),.doutb(w_n621_1[1]),.doutc(w_n621_1[2]),.din(w_n621_0[0]));
	jspl jspl_w_n621_2(.douta(w_dff_A_HGohNdA72_0),.doutb(w_n621_2[1]),.din(w_n621_0[1]));
	jspl3 jspl3_w_n622_0(.douta(w_n622_0[0]),.doutb(w_n622_0[1]),.doutc(w_n622_0[2]),.din(n622));
	jspl jspl_w_n622_1(.douta(w_n622_1[0]),.doutb(w_n622_1[1]),.din(w_n622_0[0]));
	jspl jspl_w_n623_0(.douta(w_dff_A_JgTALPGG5_0),.doutb(w_n623_0[1]),.din(n623));
	jspl3 jspl3_w_n624_0(.douta(w_n624_0[0]),.doutb(w_n624_0[1]),.doutc(w_n624_0[2]),.din(n624));
	jspl3 jspl3_w_n624_1(.douta(w_n624_1[0]),.doutb(w_n624_1[1]),.doutc(w_n624_1[2]),.din(w_n624_0[0]));
	jspl3 jspl3_w_n625_0(.douta(w_n625_0[0]),.doutb(w_n625_0[1]),.doutc(w_n625_0[2]),.din(n625));
	jspl3 jspl3_w_n628_0(.douta(w_n628_0[0]),.doutb(w_dff_A_HsDMthT51_1),.doutc(w_n628_0[2]),.din(n628));
	jspl3 jspl3_w_n629_0(.douta(w_n629_0[0]),.doutb(w_dff_A_EW7Myzab6_1),.doutc(w_n629_0[2]),.din(n629));
	jspl jspl_w_n631_0(.douta(w_dff_A_d1F1DZWd3_0),.doutb(w_n631_0[1]),.din(n631));
	jspl3 jspl3_w_n633_0(.douta(w_n633_0[0]),.doutb(w_dff_A_Nx4u9VHS9_1),.doutc(w_n633_0[2]),.din(n633));
	jspl jspl_w_n633_1(.douta(w_n633_1[0]),.doutb(w_dff_A_8ttTp3Vi9_1),.din(w_n633_0[0]));
	jspl3 jspl3_w_n636_0(.douta(w_n636_0[0]),.doutb(w_n636_0[1]),.doutc(w_n636_0[2]),.din(n636));
	jspl jspl_w_n636_1(.douta(w_n636_1[0]),.doutb(w_dff_A_Hf5VxlTZ1_1),.din(w_n636_0[0]));
	jspl3 jspl3_w_n640_0(.douta(w_n640_0[0]),.doutb(w_n640_0[1]),.doutc(w_dff_A_N2Dbv83U3_2),.din(n640));
	jspl3 jspl3_w_n640_1(.douta(w_dff_A_AmHetrVC6_0),.doutb(w_n640_1[1]),.doutc(w_n640_1[2]),.din(w_n640_0[0]));
	jspl jspl_w_n641_0(.douta(w_n641_0[0]),.doutb(w_n641_0[1]),.din(n641));
	jspl jspl_w_n642_0(.douta(w_n642_0[0]),.doutb(w_n642_0[1]),.din(n642));
	jspl3 jspl3_w_n645_0(.douta(w_n645_0[0]),.doutb(w_n645_0[1]),.doutc(w_n645_0[2]),.din(n645));
	jspl3 jspl3_w_n646_0(.douta(w_dff_A_4xVxefcF9_0),.doutb(w_n646_0[1]),.doutc(w_n646_0[2]),.din(n646));
	jspl3 jspl3_w_n649_0(.douta(w_n649_0[0]),.doutb(w_n649_0[1]),.doutc(w_dff_A_EvXNODuB0_2),.din(n649));
	jspl jspl_w_n649_1(.douta(w_n649_1[0]),.doutb(w_n649_1[1]),.din(w_n649_0[0]));
	jspl jspl_w_n650_0(.douta(w_dff_A_0ufqH2QY2_0),.doutb(w_n650_0[1]),.din(n650));
	jspl3 jspl3_w_n651_0(.douta(w_n651_0[0]),.doutb(w_dff_A_bmnWK5Td5_1),.doutc(w_dff_A_u4jsXSRD5_2),.din(w_dff_B_dnF49iJf3_3));
	jspl jspl_w_n651_1(.douta(w_dff_A_n5t01ZQF1_0),.doutb(w_n651_1[1]),.din(w_n651_0[0]));
	jspl jspl_w_n652_0(.douta(w_n652_0[0]),.doutb(w_n652_0[1]),.din(n652));
	jspl jspl_w_n661_0(.douta(w_n661_0[0]),.doutb(w_n661_0[1]),.din(n661));
	jspl jspl_w_n671_0(.douta(w_dff_A_GfxdPqk05_0),.doutb(w_n671_0[1]),.din(n671));
	jspl jspl_w_n677_0(.douta(w_n677_0[0]),.doutb(w_n677_0[1]),.din(n677));
	jspl jspl_w_n678_0(.douta(w_n678_0[0]),.doutb(w_dff_A_OWasprSn8_1),.din(n678));
	jspl jspl_w_n679_0(.douta(w_n679_0[0]),.doutb(w_dff_A_aMAMcnaI2_1),.din(n679));
	jspl jspl_w_n680_0(.douta(w_n680_0[0]),.doutb(w_dff_A_dN1kmbjE3_1),.din(n680));
	jspl3 jspl3_w_n681_0(.douta(w_dff_A_u58kNjAx0_0),.doutb(w_dff_A_ejRfFmEt0_1),.doutc(w_n681_0[2]),.din(n681));
	jspl3 jspl3_w_n681_1(.douta(w_dff_A_2ebXTWkX1_0),.doutb(w_dff_A_50lyW5Wd4_1),.doutc(w_n681_1[2]),.din(w_n681_0[0]));
	jspl jspl_w_n681_2(.douta(w_dff_A_FjXNNgSc6_0),.doutb(w_n681_2[1]),.din(w_n681_0[1]));
	jspl jspl_w_n682_0(.douta(w_n682_0[0]),.doutb(w_n682_0[1]),.din(n682));
	jspl3 jspl3_w_n687_0(.douta(w_dff_A_kiTgCdMK9_0),.doutb(w_dff_A_qh2rtEy50_1),.doutc(w_n687_0[2]),.din(n687));
	jspl jspl_w_n689_0(.douta(w_n689_0[0]),.doutb(w_n689_0[1]),.din(n689));
	jspl3 jspl3_w_n691_0(.douta(w_n691_0[0]),.doutb(w_dff_A_yUFvQGBe4_1),.doutc(w_n691_0[2]),.din(n691));
	jspl3 jspl3_w_n693_0(.douta(w_n693_0[0]),.doutb(w_dff_A_dhh6kTWW6_1),.doutc(w_n693_0[2]),.din(n693));
	jspl3 jspl3_w_n696_0(.douta(w_n696_0[0]),.doutb(w_n696_0[1]),.doutc(w_n696_0[2]),.din(n696));
	jspl jspl_w_n697_0(.douta(w_n697_0[0]),.doutb(w_n697_0[1]),.din(n697));
	jspl jspl_w_n700_0(.douta(w_n700_0[0]),.doutb(w_dff_A_K4XQ6b8l3_1),.din(n700));
	jspl jspl_w_n702_0(.douta(w_n702_0[0]),.doutb(w_n702_0[1]),.din(w_dff_B_c7Q5rMIL4_2));
	jspl3 jspl3_w_n703_0(.douta(w_n703_0[0]),.doutb(w_n703_0[1]),.doutc(w_n703_0[2]),.din(n703));
	jspl jspl_w_n705_0(.douta(w_n705_0[0]),.doutb(w_n705_0[1]),.din(n705));
	jspl jspl_w_n706_0(.douta(w_dff_A_QuPSF2du9_0),.doutb(w_n706_0[1]),.din(n706));
	jspl3 jspl3_w_n707_0(.douta(w_n707_0[0]),.doutb(w_n707_0[1]),.doutc(w_n707_0[2]),.din(n707));
	jspl jspl_w_n709_0(.douta(w_n709_0[0]),.doutb(w_n709_0[1]),.din(w_dff_B_yCe85Kji7_2));
	jspl jspl_w_n716_0(.douta(w_n716_0[0]),.doutb(w_n716_0[1]),.din(n716));
	jspl3 jspl3_w_n717_0(.douta(w_n717_0[0]),.doutb(w_dff_A_qauZ8gI89_1),.doutc(w_dff_A_2YaYhArt2_2),.din(n717));
	jspl jspl_w_n720_0(.douta(w_n720_0[0]),.doutb(w_n720_0[1]),.din(n720));
	jspl3 jspl3_w_n721_0(.douta(w_n721_0[0]),.doutb(w_dff_A_y2ad8xAP5_1),.doutc(w_n721_0[2]),.din(n721));
	jspl jspl_w_n723_0(.douta(w_dff_A_cs8aPMXM3_0),.doutb(w_n723_0[1]),.din(n723));
	jspl jspl_w_n726_0(.douta(w_n726_0[0]),.doutb(w_n726_0[1]),.din(n726));
	jspl3 jspl3_w_n727_0(.douta(w_n727_0[0]),.doutb(w_n727_0[1]),.doutc(w_n727_0[2]),.din(n727));
	jspl3 jspl3_w_n729_0(.douta(w_n729_0[0]),.doutb(w_n729_0[1]),.doutc(w_n729_0[2]),.din(n729));
	jspl jspl_w_n729_1(.douta(w_n729_1[0]),.doutb(w_n729_1[1]),.din(w_n729_0[0]));
	jspl3 jspl3_w_n732_0(.douta(w_n732_0[0]),.doutb(w_n732_0[1]),.doutc(w_n732_0[2]),.din(n732));
	jspl jspl_w_n733_0(.douta(w_n733_0[0]),.doutb(w_n733_0[1]),.din(n733));
	jspl jspl_w_n735_0(.douta(w_n735_0[0]),.doutb(w_n735_0[1]),.din(n735));
	jspl jspl_w_n736_0(.douta(w_n736_0[0]),.doutb(w_n736_0[1]),.din(n736));
	jspl3 jspl3_w_n739_0(.douta(w_n739_0[0]),.doutb(w_n739_0[1]),.doutc(w_dff_A_EfhrMbP10_2),.din(n739));
	jspl jspl_w_n739_1(.douta(w_dff_A_etJHdBC44_0),.doutb(w_n739_1[1]),.din(w_n739_0[0]));
	jspl jspl_w_n740_0(.douta(w_n740_0[0]),.doutb(w_n740_0[1]),.din(w_dff_B_kFnoWgK29_2));
	jspl jspl_w_n741_0(.douta(w_dff_A_J5FJNJKh7_0),.doutb(w_n741_0[1]),.din(w_dff_B_jDCZofNF4_2));
	jspl jspl_w_n742_0(.douta(w_n742_0[0]),.doutb(w_n742_0[1]),.din(w_dff_B_GqvEaJZe2_2));
	jspl3 jspl3_w_n744_0(.douta(w_n744_0[0]),.doutb(w_n744_0[1]),.doutc(w_dff_A_UOES35z51_2),.din(w_dff_B_luKw20Og5_3));
	jspl3 jspl3_w_n744_1(.douta(w_dff_A_lJ4K7l0o8_0),.doutb(w_n744_1[1]),.doutc(w_n744_1[2]),.din(w_n744_0[0]));
	jspl3 jspl3_w_n746_0(.douta(w_n746_0[0]),.doutb(w_n746_0[1]),.doutc(w_dff_A_MWIaVXE52_2),.din(n746));
	jspl3 jspl3_w_n746_1(.douta(w_n746_1[0]),.doutb(w_n746_1[1]),.doutc(w_n746_1[2]),.din(w_n746_0[0]));
	jspl3 jspl3_w_n747_0(.douta(w_dff_A_cENZyIIS1_0),.doutb(w_dff_A_RIpPmYAd8_1),.doutc(w_n747_0[2]),.din(n747));
	jspl3 jspl3_w_n747_1(.douta(w_n747_1[0]),.doutb(w_dff_A_DxmC90yB9_1),.doutc(w_dff_A_7X10HfUW9_2),.din(w_n747_0[0]));
	jspl3 jspl3_w_n747_2(.douta(w_n747_2[0]),.doutb(w_dff_A_WSi3kZeY5_1),.doutc(w_n747_2[2]),.din(w_n747_0[1]));
	jspl3 jspl3_w_n747_3(.douta(w_dff_A_SS5FoYVk2_0),.doutb(w_dff_A_1fLKU9vB1_1),.doutc(w_n747_3[2]),.din(w_n747_0[2]));
	jspl3 jspl3_w_n748_0(.douta(w_n748_0[0]),.doutb(w_dff_A_DAWyJfAl7_1),.doutc(w_dff_A_wCrRRJR36_2),.din(n748));
	jspl3 jspl3_w_n748_1(.douta(w_n748_1[0]),.doutb(w_dff_A_fXiwjX984_1),.doutc(w_dff_A_sWLOdO185_2),.din(w_n748_0[0]));
	jspl3 jspl3_w_n748_2(.douta(w_n748_2[0]),.doutb(w_dff_A_Fh9xh3C97_1),.doutc(w_dff_A_GzU8HWgG0_2),.din(w_n748_0[1]));
	jspl3 jspl3_w_n748_3(.douta(w_n748_3[0]),.doutb(w_n748_3[1]),.doutc(w_dff_A_scjTpqwT0_2),.din(w_n748_0[2]));
	jspl jspl_w_n748_4(.douta(w_dff_A_Q1pMjrZr8_0),.doutb(w_n748_4[1]),.din(w_n748_1[0]));
	jspl3 jspl3_w_n750_0(.douta(w_n750_0[0]),.doutb(w_dff_A_ABuFr46p9_1),.doutc(w_dff_A_Lsd8e2ir4_2),.din(n750));
	jspl jspl_w_n750_1(.douta(w_n750_1[0]),.doutb(w_n750_1[1]),.din(w_n750_0[0]));
	jspl3 jspl3_w_n751_0(.douta(w_n751_0[0]),.doutb(w_n751_0[1]),.doutc(w_dff_A_SGJuPREI6_2),.din(n751));
	jspl3 jspl3_w_n751_1(.douta(w_n751_1[0]),.doutb(w_dff_A_1tQJNjSy6_1),.doutc(w_n751_1[2]),.din(w_n751_0[0]));
	jspl jspl_w_n751_2(.douta(w_n751_2[0]),.doutb(w_n751_2[1]),.din(w_n751_0[1]));
	jspl3 jspl3_w_n753_0(.douta(w_n753_0[0]),.doutb(w_n753_0[1]),.doutc(w_n753_0[2]),.din(n753));
	jspl3 jspl3_w_n753_1(.douta(w_n753_1[0]),.doutb(w_n753_1[1]),.doutc(w_n753_1[2]),.din(w_n753_0[0]));
	jspl3 jspl3_w_n753_2(.douta(w_n753_2[0]),.doutb(w_n753_2[1]),.doutc(w_n753_2[2]),.din(w_n753_0[1]));
	jspl3 jspl3_w_n753_3(.douta(w_n753_3[0]),.doutb(w_n753_3[1]),.doutc(w_n753_3[2]),.din(w_n753_0[2]));
	jspl3 jspl3_w_n753_4(.douta(w_n753_4[0]),.doutb(w_n753_4[1]),.doutc(w_n753_4[2]),.din(w_n753_1[0]));
	jspl3 jspl3_w_n753_5(.douta(w_n753_5[0]),.doutb(w_n753_5[1]),.doutc(w_n753_5[2]),.din(w_n753_1[1]));
	jspl3 jspl3_w_n753_6(.douta(w_n753_6[0]),.doutb(w_n753_6[1]),.doutc(w_n753_6[2]),.din(w_n753_1[2]));
	jspl3 jspl3_w_n753_7(.douta(w_n753_7[0]),.doutb(w_n753_7[1]),.doutc(w_n753_7[2]),.din(w_n753_2[0]));
	jspl jspl_w_n753_8(.douta(w_n753_8[0]),.doutb(w_n753_8[1]),.din(w_n753_2[1]));
	jspl jspl_w_n759_0(.douta(w_n759_0[0]),.doutb(w_n759_0[1]),.din(n759));
	jspl jspl_w_n760_0(.douta(w_n760_0[0]),.doutb(w_n760_0[1]),.din(n760));
	jspl jspl_w_n761_0(.douta(w_n761_0[0]),.doutb(w_n761_0[1]),.din(n761));
	jspl3 jspl3_w_n765_0(.douta(w_n765_0[0]),.doutb(w_n765_0[1]),.doutc(w_n765_0[2]),.din(n765));
	jspl3 jspl3_w_n765_1(.douta(w_n765_1[0]),.doutb(w_n765_1[1]),.doutc(w_n765_1[2]),.din(w_n765_0[0]));
	jspl3 jspl3_w_n765_2(.douta(w_n765_2[0]),.doutb(w_n765_2[1]),.doutc(w_n765_2[2]),.din(w_n765_0[1]));
	jspl3 jspl3_w_n765_3(.douta(w_n765_3[0]),.doutb(w_n765_3[1]),.doutc(w_n765_3[2]),.din(w_n765_0[2]));
	jspl3 jspl3_w_n765_4(.douta(w_n765_4[0]),.doutb(w_n765_4[1]),.doutc(w_n765_4[2]),.din(w_n765_1[0]));
	jspl3 jspl3_w_n765_5(.douta(w_n765_5[0]),.doutb(w_n765_5[1]),.doutc(w_n765_5[2]),.din(w_n765_1[1]));
	jspl jspl_w_n771_0(.douta(w_n771_0[0]),.doutb(w_n771_0[1]),.din(n771));
	jspl jspl_w_n779_0(.douta(w_n779_0[0]),.doutb(w_dff_A_5khHNIqZ3_1),.din(w_dff_B_t1yzHTb16_2));
	jspl3 jspl3_w_n781_0(.douta(w_n781_0[0]),.doutb(w_n781_0[1]),.doutc(w_n781_0[2]),.din(n781));
	jspl3 jspl3_w_n783_0(.douta(w_n783_0[0]),.doutb(w_n783_0[1]),.doutc(w_n783_0[2]),.din(n783));
	jspl jspl_w_n783_1(.douta(w_n783_1[0]),.doutb(w_n783_1[1]),.din(w_n783_0[0]));
	jspl jspl_w_n786_0(.douta(w_n786_0[0]),.doutb(w_n786_0[1]),.din(n786));
	jspl jspl_w_n787_0(.douta(w_dff_A_EFYaffDo5_0),.doutb(w_n787_0[1]),.din(w_dff_B_uDLjX3Wb0_2));
	jspl3 jspl3_w_n789_0(.douta(w_n789_0[0]),.doutb(w_n789_0[1]),.doutc(w_n789_0[2]),.din(n789));
	jspl3 jspl3_w_n791_0(.douta(w_n791_0[0]),.doutb(w_n791_0[1]),.doutc(w_n791_0[2]),.din(n791));
	jspl jspl_w_n791_1(.douta(w_n791_1[0]),.doutb(w_n791_1[1]),.din(w_n791_0[0]));
	jspl jspl_w_n792_0(.douta(w_n792_0[0]),.doutb(w_n792_0[1]),.din(n792));
	jspl3 jspl3_w_n793_0(.douta(w_n793_0[0]),.doutb(w_dff_A_CLCfiF5u8_1),.doutc(w_dff_A_1vCY42P70_2),.din(w_dff_B_W0wuerbt5_3));
	jspl3 jspl3_w_n793_1(.douta(w_n793_1[0]),.doutb(w_dff_A_2W8pSPwQ6_1),.doutc(w_dff_A_j7BaaYgz3_2),.din(w_n793_0[0]));
	jspl3 jspl3_w_n793_2(.douta(w_dff_A_2X5lSC9C7_0),.doutb(w_n793_2[1]),.doutc(w_n793_2[2]),.din(w_n793_0[1]));
	jspl3 jspl3_w_n793_3(.douta(w_n793_3[0]),.doutb(w_n793_3[1]),.doutc(w_n793_3[2]),.din(w_n793_0[2]));
	jspl jspl_w_n793_4(.douta(w_dff_A_ZCK0Bsrp4_0),.doutb(w_n793_4[1]),.din(w_n793_1[0]));
	jspl3 jspl3_w_n795_0(.douta(w_n795_0[0]),.doutb(w_n795_0[1]),.doutc(w_n795_0[2]),.din(n795));
	jspl jspl_w_n795_1(.douta(w_n795_1[0]),.doutb(w_n795_1[1]),.din(w_n795_0[0]));
	jspl jspl_w_n796_0(.douta(w_n796_0[0]),.doutb(w_n796_0[1]),.din(n796));
	jspl3 jspl3_w_n797_0(.douta(w_n797_0[0]),.doutb(w_dff_A_QS2IeYwS3_1),.doutc(w_dff_A_Zckhoghx0_2),.din(w_dff_B_7IGwgqcQ8_3));
	jspl3 jspl3_w_n797_1(.douta(w_n797_1[0]),.doutb(w_dff_A_ZFvdDV6w3_1),.doutc(w_dff_A_bAjPhM2N9_2),.din(w_n797_0[0]));
	jspl3 jspl3_w_n797_2(.douta(w_n797_2[0]),.doutb(w_n797_2[1]),.doutc(w_n797_2[2]),.din(w_n797_0[1]));
	jspl3 jspl3_w_n797_3(.douta(w_n797_3[0]),.doutb(w_dff_A_wcEwDFX14_1),.doutc(w_dff_A_okWsnYcW0_2),.din(w_n797_0[2]));
	jspl jspl_w_n797_4(.douta(w_dff_A_Izq4Ek8W1_0),.doutb(w_n797_4[1]),.din(w_n797_1[0]));
	jspl3 jspl3_w_n799_0(.douta(w_n799_0[0]),.doutb(w_n799_0[1]),.doutc(w_n799_0[2]),.din(n799));
	jspl3 jspl3_w_n799_1(.douta(w_n799_1[0]),.doutb(w_n799_1[1]),.doutc(w_n799_1[2]),.din(w_n799_0[0]));
	jspl3 jspl3_w_n799_2(.douta(w_n799_2[0]),.doutb(w_n799_2[1]),.doutc(w_n799_2[2]),.din(w_n799_0[1]));
	jspl3 jspl3_w_n799_3(.douta(w_n799_3[0]),.doutb(w_n799_3[1]),.doutc(w_n799_3[2]),.din(w_n799_0[2]));
	jspl jspl_w_n799_4(.douta(w_n799_4[0]),.doutb(w_n799_4[1]),.din(w_n799_1[0]));
	jspl3 jspl3_w_n801_0(.douta(w_n801_0[0]),.doutb(w_n801_0[1]),.doutc(w_n801_0[2]),.din(n801));
	jspl3 jspl3_w_n801_1(.douta(w_n801_1[0]),.doutb(w_n801_1[1]),.doutc(w_n801_1[2]),.din(w_n801_0[0]));
	jspl3 jspl3_w_n801_2(.douta(w_n801_2[0]),.doutb(w_n801_2[1]),.doutc(w_n801_2[2]),.din(w_n801_0[1]));
	jspl3 jspl3_w_n801_3(.douta(w_n801_3[0]),.doutb(w_n801_3[1]),.doutc(w_n801_3[2]),.din(w_n801_0[2]));
	jspl jspl_w_n801_4(.douta(w_n801_4[0]),.doutb(w_n801_4[1]),.din(w_n801_1[0]));
	jspl3 jspl3_w_n806_0(.douta(w_n806_0[0]),.doutb(w_n806_0[1]),.doutc(w_n806_0[2]),.din(n806));
	jspl jspl_w_n809_0(.douta(w_dff_A_kiedNMSw1_0),.doutb(w_n809_0[1]),.din(n809));
	jspl jspl_w_n819_0(.douta(w_n819_0[0]),.doutb(w_n819_0[1]),.din(n819));
	jspl jspl_w_n821_0(.douta(w_dff_A_tduSDlpK3_0),.doutb(w_n821_0[1]),.din(n821));
	jspl3 jspl3_w_n828_0(.douta(w_n828_0[0]),.doutb(w_dff_A_5tZlyRKT7_1),.doutc(w_dff_A_IUNeA1Eq8_2),.din(w_dff_B_uzq9ZczS6_3));
	jspl jspl_w_n829_0(.douta(w_n829_0[0]),.doutb(w_dff_A_NH7oi9Al9_1),.din(n829));
	jspl jspl_w_n832_0(.douta(w_n832_0[0]),.doutb(w_n832_0[1]),.din(n832));
	jspl jspl_w_n839_0(.douta(w_n839_0[0]),.doutb(w_n839_0[1]),.din(n839));
	jspl3 jspl3_w_n840_0(.douta(w_n840_0[0]),.doutb(w_dff_A_uFGO2QA43_1),.doutc(w_dff_A_225P8l8c2_2),.din(w_dff_B_47vXz1si6_3));
	jspl3 jspl3_w_n840_1(.douta(w_n840_1[0]),.doutb(w_dff_A_OAmdyT2Q3_1),.doutc(w_dff_A_2csyo9hG7_2),.din(w_n840_0[0]));
	jspl3 jspl3_w_n840_2(.douta(w_dff_A_SjmIzxNS3_0),.doutb(w_n840_2[1]),.doutc(w_n840_2[2]),.din(w_n840_0[1]));
	jspl3 jspl3_w_n840_3(.douta(w_n840_3[0]),.doutb(w_n840_3[1]),.doutc(w_n840_3[2]),.din(w_n840_0[2]));
	jspl jspl_w_n840_4(.douta(w_dff_A_fGW91Ct89_0),.doutb(w_n840_4[1]),.din(w_n840_1[0]));
	jspl jspl_w_n842_0(.douta(w_n842_0[0]),.doutb(w_n842_0[1]),.din(n842));
	jspl3 jspl3_w_n843_0(.douta(w_n843_0[0]),.doutb(w_dff_A_EWrfPdBv2_1),.doutc(w_dff_A_pPhhY0IA6_2),.din(w_dff_B_otVDLEHT6_3));
	jspl3 jspl3_w_n843_1(.douta(w_n843_1[0]),.doutb(w_dff_A_i6yV8PVe8_1),.doutc(w_dff_A_8m2i4gXb4_2),.din(w_n843_0[0]));
	jspl3 jspl3_w_n843_2(.douta(w_n843_2[0]),.doutb(w_n843_2[1]),.doutc(w_n843_2[2]),.din(w_n843_0[1]));
	jspl3 jspl3_w_n843_3(.douta(w_n843_3[0]),.doutb(w_dff_A_9OgRyhsy3_1),.doutc(w_dff_A_X0jYu4GN5_2),.din(w_n843_0[2]));
	jspl jspl_w_n843_4(.douta(w_dff_A_jbpOdlvy3_0),.doutb(w_n843_4[1]),.din(w_n843_1[0]));
	jspl3 jspl3_w_n845_0(.douta(w_n845_0[0]),.doutb(w_n845_0[1]),.doutc(w_n845_0[2]),.din(n845));
	jspl3 jspl3_w_n845_1(.douta(w_n845_1[0]),.doutb(w_n845_1[1]),.doutc(w_n845_1[2]),.din(w_n845_0[0]));
	jspl3 jspl3_w_n845_2(.douta(w_n845_2[0]),.doutb(w_n845_2[1]),.doutc(w_n845_2[2]),.din(w_n845_0[1]));
	jspl3 jspl3_w_n845_3(.douta(w_n845_3[0]),.doutb(w_n845_3[1]),.doutc(w_n845_3[2]),.din(w_n845_0[2]));
	jspl jspl_w_n845_4(.douta(w_n845_4[0]),.doutb(w_n845_4[1]),.din(w_n845_1[0]));
	jspl3 jspl3_w_n847_0(.douta(w_n847_0[0]),.doutb(w_n847_0[1]),.doutc(w_n847_0[2]),.din(n847));
	jspl3 jspl3_w_n847_1(.douta(w_n847_1[0]),.doutb(w_n847_1[1]),.doutc(w_n847_1[2]),.din(w_n847_0[0]));
	jspl3 jspl3_w_n847_2(.douta(w_n847_2[0]),.doutb(w_n847_2[1]),.doutc(w_n847_2[2]),.din(w_n847_0[1]));
	jspl3 jspl3_w_n847_3(.douta(w_n847_3[0]),.doutb(w_n847_3[1]),.doutc(w_n847_3[2]),.din(w_n847_0[2]));
	jspl jspl_w_n847_4(.douta(w_n847_4[0]),.doutb(w_n847_4[1]),.din(w_n847_1[0]));
	jspl jspl_w_n853_0(.douta(w_n853_0[0]),.doutb(w_dff_A_pddUHG9k4_1),.din(w_dff_B_WzfnIOVU6_2));
	jspl jspl_w_n855_0(.douta(w_n855_0[0]),.doutb(w_n855_0[1]),.din(n855));
	jspl jspl_w_n856_0(.douta(w_n856_0[0]),.doutb(w_n856_0[1]),.din(n856));
	jspl jspl_w_n857_0(.douta(w_n857_0[0]),.doutb(w_n857_0[1]),.din(n857));
	jspl jspl_w_n859_0(.douta(w_n859_0[0]),.doutb(w_n859_0[1]),.din(n859));
	jspl jspl_w_n862_0(.douta(w_dff_A_kqaLlRCo8_0),.doutb(w_n862_0[1]),.din(n862));
	jspl jspl_w_n869_0(.douta(w_dff_A_cp2V9q6e7_0),.doutb(w_n869_0[1]),.din(n869));
	jspl jspl_w_n877_0(.douta(w_n877_0[0]),.doutb(w_n877_0[1]),.din(n877));
	jspl jspl_w_n879_0(.douta(w_dff_A_MkzCM3QZ5_0),.doutb(w_n879_0[1]),.din(n879));
	jspl jspl_w_n881_0(.douta(w_n881_0[0]),.doutb(w_n881_0[1]),.din(n881));
	jspl jspl_w_n892_0(.douta(w_n892_0[0]),.doutb(w_n892_0[1]),.din(n892));
	jspl jspl_w_n914_0(.douta(w_n914_0[0]),.doutb(w_n914_0[1]),.din(n914));
	jspl jspl_w_n928_0(.douta(w_n928_0[0]),.doutb(w_dff_A_ElfGvmoY0_1),.din(n928));
	jspl3 jspl3_w_n930_0(.douta(w_n930_0[0]),.doutb(w_n930_0[1]),.doutc(w_dff_A_iFfrMLOE4_2),.din(w_dff_B_E3phhCox2_3));
	jspl jspl_w_n932_0(.douta(w_n932_0[0]),.doutb(w_n932_0[1]),.din(w_dff_B_N3N1Y1jD7_2));
	jspl3 jspl3_w_n936_0(.douta(w_n936_0[0]),.doutb(w_n936_0[1]),.doutc(w_n936_0[2]),.din(n936));
	jspl jspl_w_n938_0(.douta(w_n938_0[0]),.doutb(w_n938_0[1]),.din(n938));
	jspl jspl_w_n941_0(.douta(w_n941_0[0]),.doutb(w_n941_0[1]),.din(n941));
	jspl jspl_w_n943_0(.douta(w_n943_0[0]),.doutb(w_dff_A_sk2iuow46_1),.din(n943));
	jspl jspl_w_n944_0(.douta(w_n944_0[0]),.doutb(w_dff_A_qTwRcuC64_1),.din(n944));
	jspl jspl_w_n946_0(.douta(w_n946_0[0]),.doutb(w_n946_0[1]),.din(n946));
	jspl3 jspl3_w_n948_0(.douta(w_dff_A_GZztyjC65_0),.doutb(w_dff_A_o9kwGvjU0_1),.doutc(w_n948_0[2]),.din(n948));
	jspl jspl_w_n953_0(.douta(w_n953_0[0]),.doutb(w_dff_A_wjn5Vn6R9_1),.din(n953));
	jspl jspl_w_n954_0(.douta(w_n954_0[0]),.doutb(w_n954_0[1]),.din(n954));
	jspl jspl_w_n968_0(.douta(w_n968_0[0]),.doutb(w_n968_0[1]),.din(w_dff_B_4snys8hk0_2));
	jspl jspl_w_n971_0(.douta(w_n971_0[0]),.doutb(w_dff_A_05jXUVYb5_1),.din(n971));
	jspl jspl_w_n972_0(.douta(w_n972_0[0]),.doutb(w_dff_A_EQbq1Jpa1_1),.din(n972));
	jspl jspl_w_n973_0(.douta(w_n973_0[0]),.doutb(w_n973_0[1]),.din(n973));
	jspl jspl_w_n984_0(.douta(w_n984_0[0]),.doutb(w_n984_0[1]),.din(n984));
	jspl3 jspl3_w_n985_0(.douta(w_n985_0[0]),.doutb(w_dff_A_PWutiuU86_1),.doutc(w_dff_A_AL1UiXwR6_2),.din(n985));
	jspl3 jspl3_w_n985_1(.douta(w_dff_A_YSPdOOlB5_0),.doutb(w_n985_1[1]),.doutc(w_dff_A_YrOEY4DL7_2),.din(w_n985_0[0]));
	jspl3 jspl3_w_n985_2(.douta(w_n985_2[0]),.doutb(w_dff_A_BdZzNksn6_1),.doutc(w_dff_A_ECbPHj9f5_2),.din(w_n985_0[1]));
	jspl3 jspl3_w_n985_3(.douta(w_n985_3[0]),.doutb(w_n985_3[1]),.doutc(w_n985_3[2]),.din(w_n985_0[2]));
	jspl jspl_w_n985_4(.douta(w_dff_A_lbsv0ReK6_0),.doutb(w_n985_4[1]),.din(w_n985_1[0]));
	jspl jspl_w_n987_0(.douta(w_n987_0[0]),.doutb(w_n987_0[1]),.din(n987));
	jspl3 jspl3_w_n988_0(.douta(w_n988_0[0]),.doutb(w_dff_A_oWhN8KOx3_1),.doutc(w_dff_A_rMbDKlHt8_2),.din(n988));
	jspl3 jspl3_w_n988_1(.douta(w_dff_A_pWkXD5lq7_0),.doutb(w_n988_1[1]),.doutc(w_dff_A_m3SICdOU5_2),.din(w_n988_0[0]));
	jspl3 jspl3_w_n988_2(.douta(w_n988_2[0]),.doutb(w_n988_2[1]),.doutc(w_dff_A_rrTVTbpo5_2),.din(w_n988_0[1]));
	jspl3 jspl3_w_n988_3(.douta(w_dff_A_r7GzCRg66_0),.doutb(w_dff_A_uLwnQKui8_1),.doutc(w_n988_3[2]),.din(w_n988_0[2]));
	jspl jspl_w_n988_4(.douta(w_dff_A_5DV6LkPy1_0),.doutb(w_n988_4[1]),.din(w_n988_1[0]));
	jspl3 jspl3_w_n990_0(.douta(w_n990_0[0]),.doutb(w_n990_0[1]),.doutc(w_n990_0[2]),.din(n990));
	jspl3 jspl3_w_n990_1(.douta(w_n990_1[0]),.doutb(w_n990_1[1]),.doutc(w_n990_1[2]),.din(w_n990_0[0]));
	jspl3 jspl3_w_n990_2(.douta(w_n990_2[0]),.doutb(w_n990_2[1]),.doutc(w_n990_2[2]),.din(w_n990_0[1]));
	jspl3 jspl3_w_n990_3(.douta(w_n990_3[0]),.doutb(w_n990_3[1]),.doutc(w_n990_3[2]),.din(w_n990_0[2]));
	jspl jspl_w_n990_4(.douta(w_n990_4[0]),.doutb(w_n990_4[1]),.din(w_n990_1[0]));
	jspl3 jspl3_w_n992_0(.douta(w_n992_0[0]),.doutb(w_n992_0[1]),.doutc(w_n992_0[2]),.din(n992));
	jspl3 jspl3_w_n992_1(.douta(w_n992_1[0]),.doutb(w_n992_1[1]),.doutc(w_n992_1[2]),.din(w_n992_0[0]));
	jspl3 jspl3_w_n992_2(.douta(w_n992_2[0]),.doutb(w_n992_2[1]),.doutc(w_n992_2[2]),.din(w_n992_0[1]));
	jspl3 jspl3_w_n992_3(.douta(w_n992_3[0]),.doutb(w_n992_3[1]),.doutc(w_n992_3[2]),.din(w_n992_0[2]));
	jspl jspl_w_n992_4(.douta(w_n992_4[0]),.doutb(w_n992_4[1]),.din(w_n992_1[0]));
	jspl jspl_w_n998_0(.douta(w_n998_0[0]),.doutb(w_n998_0[1]),.din(n998));
	jspl3 jspl3_w_n999_0(.douta(w_n999_0[0]),.doutb(w_dff_A_fE3PXaSr1_1),.doutc(w_dff_A_4Xqc6g2q8_2),.din(n999));
	jspl3 jspl3_w_n999_1(.douta(w_dff_A_C7kY2QMG8_0),.doutb(w_n999_1[1]),.doutc(w_dff_A_BW1HhNof2_2),.din(w_n999_0[0]));
	jspl3 jspl3_w_n999_2(.douta(w_n999_2[0]),.doutb(w_dff_A_SAJWWZnn5_1),.doutc(w_dff_A_4jcnKlLF8_2),.din(w_n999_0[1]));
	jspl3 jspl3_w_n999_3(.douta(w_n999_3[0]),.doutb(w_n999_3[1]),.doutc(w_n999_3[2]),.din(w_n999_0[2]));
	jspl jspl_w_n999_4(.douta(w_dff_A_PyIf5qVQ1_0),.doutb(w_n999_4[1]),.din(w_n999_1[0]));
	jspl jspl_w_n1001_0(.douta(w_n1001_0[0]),.doutb(w_n1001_0[1]),.din(n1001));
	jspl3 jspl3_w_n1002_0(.douta(w_n1002_0[0]),.doutb(w_dff_A_06tVJ6yW9_1),.doutc(w_dff_A_XrIU7Ouo9_2),.din(n1002));
	jspl3 jspl3_w_n1002_1(.douta(w_dff_A_HgKl2ejf3_0),.doutb(w_n1002_1[1]),.doutc(w_dff_A_qqem33b11_2),.din(w_n1002_0[0]));
	jspl3 jspl3_w_n1002_2(.douta(w_n1002_2[0]),.doutb(w_n1002_2[1]),.doutc(w_dff_A_KzcxDb729_2),.din(w_n1002_0[1]));
	jspl3 jspl3_w_n1002_3(.douta(w_dff_A_dpCZoQk20_0),.doutb(w_dff_A_7luvimY03_1),.doutc(w_n1002_3[2]),.din(w_n1002_0[2]));
	jspl jspl_w_n1002_4(.douta(w_dff_A_TExLgcsK5_0),.doutb(w_n1002_4[1]),.din(w_n1002_1[0]));
	jspl3 jspl3_w_n1004_0(.douta(w_n1004_0[0]),.doutb(w_n1004_0[1]),.doutc(w_n1004_0[2]),.din(n1004));
	jspl3 jspl3_w_n1004_1(.douta(w_n1004_1[0]),.doutb(w_n1004_1[1]),.doutc(w_n1004_1[2]),.din(w_n1004_0[0]));
	jspl3 jspl3_w_n1004_2(.douta(w_n1004_2[0]),.doutb(w_n1004_2[1]),.doutc(w_n1004_2[2]),.din(w_n1004_0[1]));
	jspl3 jspl3_w_n1004_3(.douta(w_n1004_3[0]),.doutb(w_n1004_3[1]),.doutc(w_n1004_3[2]),.din(w_n1004_0[2]));
	jspl jspl_w_n1004_4(.douta(w_n1004_4[0]),.doutb(w_n1004_4[1]),.din(w_n1004_1[0]));
	jspl3 jspl3_w_n1006_0(.douta(w_n1006_0[0]),.doutb(w_n1006_0[1]),.doutc(w_n1006_0[2]),.din(n1006));
	jspl3 jspl3_w_n1006_1(.douta(w_n1006_1[0]),.doutb(w_n1006_1[1]),.doutc(w_n1006_1[2]),.din(w_n1006_0[0]));
	jspl3 jspl3_w_n1006_2(.douta(w_n1006_2[0]),.doutb(w_n1006_2[1]),.doutc(w_n1006_2[2]),.din(w_n1006_0[1]));
	jspl3 jspl3_w_n1006_3(.douta(w_n1006_3[0]),.doutb(w_n1006_3[1]),.doutc(w_n1006_3[2]),.din(w_n1006_0[2]));
	jspl jspl_w_n1006_4(.douta(w_n1006_4[0]),.doutb(w_n1006_4[1]),.din(w_n1006_1[0]));
	jspl3 jspl3_w_n1012_0(.douta(w_n1012_0[0]),.doutb(w_n1012_0[1]),.doutc(w_n1012_0[2]),.din(n1012));
	jspl jspl_w_n1012_1(.douta(w_n1012_1[0]),.doutb(w_n1012_1[1]),.din(w_n1012_0[0]));
	jspl3 jspl3_w_n1014_0(.douta(w_n1014_0[0]),.doutb(w_n1014_0[1]),.doutc(w_n1014_0[2]),.din(n1014));
	jspl jspl_w_n1014_1(.douta(w_n1014_1[0]),.doutb(w_n1014_1[1]),.din(w_n1014_0[0]));
	jspl3 jspl3_w_n1021_0(.douta(w_n1021_0[0]),.doutb(w_n1021_0[1]),.doutc(w_n1021_0[2]),.din(n1021));
	jspl jspl_w_n1021_1(.douta(w_n1021_1[0]),.doutb(w_n1021_1[1]),.din(w_n1021_0[0]));
	jspl3 jspl3_w_n1023_0(.douta(w_n1023_0[0]),.doutb(w_n1023_0[1]),.doutc(w_n1023_0[2]),.din(n1023));
	jspl jspl_w_n1023_1(.douta(w_n1023_1[0]),.doutb(w_n1023_1[1]),.din(w_n1023_0[0]));
	jspl3 jspl3_w_n1030_0(.douta(w_n1030_0[0]),.doutb(w_n1030_0[1]),.doutc(w_n1030_0[2]),.din(n1030));
	jspl jspl_w_n1030_1(.douta(w_n1030_1[0]),.doutb(w_n1030_1[1]),.din(w_n1030_0[0]));
	jspl3 jspl3_w_n1032_0(.douta(w_n1032_0[0]),.doutb(w_n1032_0[1]),.doutc(w_n1032_0[2]),.din(n1032));
	jspl jspl_w_n1032_1(.douta(w_n1032_1[0]),.doutb(w_n1032_1[1]),.din(w_n1032_0[0]));
	jspl3 jspl3_w_n1039_0(.douta(w_n1039_0[0]),.doutb(w_n1039_0[1]),.doutc(w_n1039_0[2]),.din(n1039));
	jspl jspl_w_n1039_1(.douta(w_n1039_1[0]),.doutb(w_n1039_1[1]),.din(w_n1039_0[0]));
	jspl3 jspl3_w_n1041_0(.douta(w_n1041_0[0]),.doutb(w_n1041_0[1]),.doutc(w_n1041_0[2]),.din(n1041));
	jspl jspl_w_n1041_1(.douta(w_n1041_1[0]),.doutb(w_n1041_1[1]),.din(w_n1041_0[0]));
	jspl jspl_w_n1142_0(.douta(w_dff_A_EI7ad8R13_0),.doutb(w_n1142_0[1]),.din(n1142));
	jspl jspl_w_n1151_0(.douta(w_n1151_0[0]),.doutb(w_n1151_0[1]),.din(n1151));
	jspl3 jspl3_w_n1163_0(.douta(w_n1163_0[0]),.doutb(w_n1163_0[1]),.doutc(w_n1163_0[2]),.din(n1163));
	jspl3 jspl3_w_n1163_1(.douta(w_n1163_1[0]),.doutb(w_n1163_1[1]),.doutc(w_n1163_1[2]),.din(w_n1163_0[0]));
	jspl3 jspl3_w_n1197_0(.douta(w_n1197_0[0]),.doutb(w_n1197_0[1]),.doutc(w_n1197_0[2]),.din(n1197));
	jspl3 jspl3_w_n1197_1(.douta(w_n1197_1[0]),.doutb(w_n1197_1[1]),.doutc(w_n1197_1[2]),.din(w_n1197_0[0]));
	jspl3 jspl3_w_n1205_0(.douta(w_n1205_0[0]),.doutb(w_n1205_0[1]),.doutc(w_n1205_0[2]),.din(n1205));
	jspl3 jspl3_w_n1205_1(.douta(w_n1205_1[0]),.doutb(w_n1205_1[1]),.doutc(w_n1205_1[2]),.din(w_n1205_0[0]));
	jspl3 jspl3_w_n1235_0(.douta(w_n1235_0[0]),.doutb(w_n1235_0[1]),.doutc(w_n1235_0[2]),.din(n1235));
	jspl jspl_w_n1235_1(.douta(w_n1235_1[0]),.doutb(w_n1235_1[1]),.din(w_n1235_0[0]));
	jspl3 jspl3_w_n1242_0(.douta(w_n1242_0[0]),.doutb(w_n1242_0[1]),.doutc(w_n1242_0[2]),.din(n1242));
	jspl jspl_w_n1242_1(.douta(w_n1242_1[0]),.doutb(w_n1242_1[1]),.din(w_n1242_0[0]));
	jspl3 jspl3_w_n1244_0(.douta(w_n1244_0[0]),.doutb(w_n1244_0[1]),.doutc(w_n1244_0[2]),.din(n1244));
	jspl jspl_w_n1244_1(.douta(w_n1244_1[0]),.doutb(w_n1244_1[1]),.din(w_n1244_0[0]));
	jspl3 jspl3_w_n1251_0(.douta(w_n1251_0[0]),.doutb(w_n1251_0[1]),.doutc(w_n1251_0[2]),.din(n1251));
	jspl jspl_w_n1251_1(.douta(w_n1251_1[0]),.doutb(w_n1251_1[1]),.din(w_n1251_0[0]));
	jspl3 jspl3_w_n1253_0(.douta(w_n1253_0[0]),.doutb(w_n1253_0[1]),.doutc(w_n1253_0[2]),.din(n1253));
	jspl jspl_w_n1253_1(.douta(w_n1253_1[0]),.doutb(w_n1253_1[1]),.din(w_n1253_0[0]));
	jspl jspl_w_n1358_0(.douta(w_n1358_0[0]),.doutb(w_n1358_0[1]),.din(n1358));
	jspl jspl_w_n1383_0(.douta(w_dff_A_6wIWtBnV1_0),.doutb(w_n1383_0[1]),.din(n1383));
	jspl jspl_w_n1391_0(.douta(w_dff_A_o4GHBTC55_0),.doutb(w_n1391_0[1]),.din(n1391));
	jspl jspl_w_n1394_0(.douta(w_n1394_0[0]),.doutb(w_dff_A_1ROaP6aB5_1),.din(n1394));
	jspl jspl_w_n1398_0(.douta(w_n1398_0[0]),.doutb(w_n1398_0[1]),.din(n1398));
	jspl jspl_w_n1399_0(.douta(w_n1399_0[0]),.doutb(w_n1399_0[1]),.din(n1399));
	jspl jspl_w_n1409_0(.douta(w_dff_A_0EqgIHIf3_0),.doutb(w_n1409_0[1]),.din(n1409));
	jspl jspl_w_n1410_0(.douta(w_n1410_0[0]),.doutb(w_n1410_0[1]),.din(w_dff_B_KpRwIewu3_2));
	jspl jspl_w_n1411_0(.douta(w_dff_A_1QglDTsf6_0),.doutb(w_n1411_0[1]),.din(n1411));
	jspl jspl_w_n1421_0(.douta(w_dff_A_dKjpUH6t2_0),.doutb(w_n1421_0[1]),.din(n1421));
	jspl jspl_w_n1425_0(.douta(w_n1425_0[0]),.doutb(w_n1425_0[1]),.din(n1425));
	jspl jspl_w_n1434_0(.douta(w_n1434_0[0]),.doutb(w_n1434_0[1]),.din(n1434));
	jspl jspl_w_n1438_0(.douta(w_n1438_0[0]),.doutb(w_dff_A_OosqPwxe4_1),.din(n1438));
	jspl jspl_w_n1445_0(.douta(w_n1445_0[0]),.doutb(w_n1445_0[1]),.din(n1445));
	jspl jspl_w_n1446_0(.douta(w_n1446_0[0]),.doutb(w_n1446_0[1]),.din(n1446));
	jspl jspl_w_n1447_0(.douta(w_n1447_0[0]),.doutb(w_dff_A_D7xd73bS1_1),.din(n1447));
	jspl jspl_w_n1452_0(.douta(w_n1452_0[0]),.doutb(w_n1452_0[1]),.din(n1452));
	jspl jspl_w_n1494_0(.douta(w_n1494_0[0]),.doutb(w_n1494_0[1]),.din(n1494));
	jspl jspl_w_n1533_0(.douta(w_n1533_0[0]),.doutb(w_n1533_0[1]),.din(w_dff_B_MCAgvn5H2_2));
	jspl jspl_w_n1543_0(.douta(w_n1543_0[0]),.doutb(w_n1543_0[1]),.din(w_dff_B_hPZshaVc0_2));
	jspl jspl_w_n1545_0(.douta(w_n1545_0[0]),.doutb(w_n1545_0[1]),.din(n1545));
	jspl jspl_w_n1553_0(.douta(w_n1553_0[0]),.doutb(w_n1553_0[1]),.din(w_dff_B_3dRmf2ut7_2));
	jspl jspl_w_n1555_0(.douta(w_dff_A_JfvCvCPd3_0),.doutb(w_n1555_0[1]),.din(n1555));
	jspl jspl_w_n1560_0(.douta(w_n1560_0[0]),.doutb(w_n1560_0[1]),.din(n1560));
	jspl jspl_w_n1568_0(.douta(w_n1568_0[0]),.doutb(w_dff_A_DmbG28e35_1),.din(w_dff_B_vMN4xilR7_2));
	jspl jspl_w_n1591_0(.douta(w_n1591_0[0]),.doutb(w_n1591_0[1]),.din(n1591));
	jspl jspl_w_n1597_0(.douta(w_n1597_0[0]),.doutb(w_n1597_0[1]),.din(n1597));
	jspl3 jspl3_w_n1601_0(.douta(w_n1601_0[0]),.doutb(w_n1601_0[1]),.doutc(w_n1601_0[2]),.din(n1601));
	jspl jspl_w_n1602_0(.douta(w_n1602_0[0]),.doutb(w_n1602_0[1]),.din(n1602));
	jspl jspl_w_n1609_0(.douta(w_n1609_0[0]),.doutb(w_dff_A_DtNh0NaG6_1),.din(n1609));
	jspl jspl_w_n1610_0(.douta(w_n1610_0[0]),.doutb(w_n1610_0[1]),.din(n1610));
	jspl jspl_w_n1624_0(.douta(w_n1624_0[0]),.doutb(w_n1624_0[1]),.din(w_dff_B_Zp36ZbYQ3_2));
	jspl jspl_w_n1629_0(.douta(w_n1629_0[0]),.doutb(w_n1629_0[1]),.din(n1629));
	jspl jspl_w_n1631_0(.douta(w_n1631_0[0]),.doutb(w_n1631_0[1]),.din(w_dff_B_yuVHT2KF9_2));
	jspl jspl_w_n1634_0(.douta(w_n1634_0[0]),.doutb(w_n1634_0[1]),.din(w_dff_B_IijeVrdw9_2));
	jdff dff_B_WGdD0rVS3_1(.din(G136),.dout(w_dff_B_WGdD0rVS3_1),.clk(gclk));
	jdff dff_B_f0LYeUl25_0(.din(G2824),.dout(w_dff_B_f0LYeUl25_0),.clk(gclk));
	jdff dff_A_BFIIhYPO2_0(.dout(w_G809_3[0]),.din(w_dff_A_BFIIhYPO2_0),.clk(gclk));
	jdff dff_B_VJcHhuhL0_0(.din(n342),.dout(w_dff_B_VJcHhuhL0_0),.clk(gclk));
	jdff dff_A_YBhqqeWI3_2(.dout(w_G809_2[2]),.din(w_dff_A_YBhqqeWI3_2),.clk(gclk));
	jdff dff_B_BlANR4eP3_1(.din(G24),.dout(w_dff_B_BlANR4eP3_1),.clk(gclk));
	jdff dff_B_JCFpbHak3_0(.din(n347),.dout(w_dff_B_JCFpbHak3_0),.clk(gclk));
	jdff dff_B_q4l2q9D84_1(.din(G26),.dout(w_dff_B_q4l2q9D84_1),.clk(gclk));
	jdff dff_A_p8cfZKe11_0(.dout(w_G141_2[0]),.din(w_dff_A_p8cfZKe11_0),.clk(gclk));
	jdff dff_A_mDj9H6QG7_0(.dout(w_dff_A_p8cfZKe11_0),.din(w_dff_A_mDj9H6QG7_0),.clk(gclk));
	jdff dff_A_I6kXeqgr8_1(.dout(w_G141_2[1]),.din(w_dff_A_I6kXeqgr8_1),.clk(gclk));
	jdff dff_A_AkhK1X9s5_1(.dout(w_dff_A_I6kXeqgr8_1),.din(w_dff_A_AkhK1X9s5_1),.clk(gclk));
	jdff dff_B_8ew7en6g4_0(.din(n352),.dout(w_dff_B_8ew7en6g4_0),.clk(gclk));
	jdff dff_B_WJPsYA0z2_1(.din(G79),.dout(w_dff_B_WJPsYA0z2_1),.clk(gclk));
	jdff dff_B_eOyn8kPV5_0(.din(n357),.dout(w_dff_B_eOyn8kPV5_0),.clk(gclk));
	jdff dff_B_nZ4R98sA0_1(.din(G82),.dout(w_dff_B_nZ4R98sA0_1),.clk(gclk));
	jdff dff_A_UZf91e0e1_0(.dout(w_G2358_2[0]),.din(w_dff_A_UZf91e0e1_0),.clk(gclk));
	jdff dff_A_kvAw0xGb1_1(.dout(w_G2358_2[1]),.din(w_dff_A_kvAw0xGb1_1),.clk(gclk));
	jdff dff_A_cmdfPIZp2_1(.dout(w_G141_1[1]),.din(w_dff_A_cmdfPIZp2_1),.clk(gclk));
	jdff dff_A_3bTWSZ4q7_1(.dout(w_dff_A_cmdfPIZp2_1),.din(w_dff_A_3bTWSZ4q7_1),.clk(gclk));
	jdff dff_A_Oq6xX8ZF7_2(.dout(w_G141_1[2]),.din(w_dff_A_Oq6xX8ZF7_2),.clk(gclk));
	jdff dff_A_gGbZoHhG3_2(.dout(w_dff_A_Oq6xX8ZF7_2),.din(w_dff_A_gGbZoHhG3_2),.clk(gclk));
	jdff dff_B_eCm3PMS85_1(.din(n384),.dout(w_dff_B_eCm3PMS85_1),.clk(gclk));
	jdff dff_B_e4aO8TUb8_1(.din(w_dff_B_eCm3PMS85_1),.dout(w_dff_B_e4aO8TUb8_1),.clk(gclk));
	jdff dff_B_QKD54ivv8_1(.din(w_dff_B_e4aO8TUb8_1),.dout(w_dff_B_QKD54ivv8_1),.clk(gclk));
	jdff dff_B_8ntSLRtx1_0(.din(n446),.dout(w_dff_B_8ntSLRtx1_0),.clk(gclk));
	jdff dff_B_905voHzG3_0(.din(w_dff_B_8ntSLRtx1_0),.dout(w_dff_B_905voHzG3_0),.clk(gclk));
	jdff dff_B_gU6HXDMJ4_1(.din(n483),.dout(w_dff_B_gU6HXDMJ4_1),.clk(gclk));
	jdff dff_B_yw7XDC1h4_1(.din(n506),.dout(w_dff_B_yw7XDC1h4_1),.clk(gclk));
	jdff dff_B_DSVEcvlF0_2(.din(n709),.dout(w_dff_B_DSVEcvlF0_2),.clk(gclk));
	jdff dff_B_yBanOqkZ1_2(.din(w_dff_B_DSVEcvlF0_2),.dout(w_dff_B_yBanOqkZ1_2),.clk(gclk));
	jdff dff_B_yCe85Kji7_2(.din(w_dff_B_yBanOqkZ1_2),.dout(w_dff_B_yCe85Kji7_2),.clk(gclk));
	jdff dff_B_tml5FdyV9_1(.din(n698),.dout(w_dff_B_tml5FdyV9_1),.clk(gclk));
	jdff dff_B_F8cqQGOc6_1(.din(n699),.dout(w_dff_B_F8cqQGOc6_1),.clk(gclk));
	jdff dff_A_Y58LOX3i0_1(.dout(w_n607_0[1]),.din(w_dff_A_Y58LOX3i0_1),.clk(gclk));
	jdff dff_B_VSrcI6kO7_0(.din(n606),.dout(w_dff_B_VSrcI6kO7_0),.clk(gclk));
	jdff dff_B_W1C3vtJh6_0(.din(w_dff_B_VSrcI6kO7_0),.dout(w_dff_B_W1C3vtJh6_0),.clk(gclk));
	jdff dff_B_GqvEaJZe2_2(.din(n742),.dout(w_dff_B_GqvEaJZe2_2),.clk(gclk));
	jdff dff_A_n5t01ZQF1_0(.dout(w_n651_1[0]),.din(w_dff_A_n5t01ZQF1_0),.clk(gclk));
	jdff dff_B_PhSDkhuw2_0(.din(n804),.dout(w_dff_B_PhSDkhuw2_0),.clk(gclk));
	jdff dff_B_w4igoQQ31_0(.din(w_dff_B_PhSDkhuw2_0),.dout(w_dff_B_w4igoQQ31_0),.clk(gclk));
	jdff dff_B_Vzbf7DTq3_0(.din(n803),.dout(w_dff_B_Vzbf7DTq3_0),.clk(gclk));
	jdff dff_B_8H1wQF9T7_0(.din(w_dff_B_Vzbf7DTq3_0),.dout(w_dff_B_8H1wQF9T7_0),.clk(gclk));
	jdff dff_B_yjg5KfqY6_0(.din(w_dff_B_8H1wQF9T7_0),.dout(w_dff_B_yjg5KfqY6_0),.clk(gclk));
	jdff dff_B_TeOv1NbB9_0(.din(w_dff_B_yjg5KfqY6_0),.dout(w_dff_B_TeOv1NbB9_0),.clk(gclk));
	jdff dff_B_F722iPpp8_0(.din(n802),.dout(w_dff_B_F722iPpp8_0),.clk(gclk));
	jdff dff_B_2cN4VASt5_0(.din(n850),.dout(w_dff_B_2cN4VASt5_0),.clk(gclk));
	jdff dff_B_Y4WLp8Fb2_0(.din(w_dff_B_2cN4VASt5_0),.dout(w_dff_B_Y4WLp8Fb2_0),.clk(gclk));
	jdff dff_B_9BhNk8EB2_0(.din(n849),.dout(w_dff_B_9BhNk8EB2_0),.clk(gclk));
	jdff dff_B_SR0lf29E3_0(.din(w_dff_B_9BhNk8EB2_0),.dout(w_dff_B_SR0lf29E3_0),.clk(gclk));
	jdff dff_B_z1phqwup6_0(.din(w_dff_B_SR0lf29E3_0),.dout(w_dff_B_z1phqwup6_0),.clk(gclk));
	jdff dff_B_rySoRXaP3_0(.din(w_dff_B_z1phqwup6_0),.dout(w_dff_B_rySoRXaP3_0),.clk(gclk));
	jdff dff_B_Mw5zA2y87_0(.din(n848),.dout(w_dff_B_Mw5zA2y87_0),.clk(gclk));
	jdff dff_B_OBQcQGTx9_2(.din(G61),.dout(w_dff_B_OBQcQGTx9_2),.clk(gclk));
	jdff dff_B_aHqIICak1_2(.din(G11),.dout(w_dff_B_aHqIICak1_2),.clk(gclk));
	jdff dff_B_BiD5EdXq3_2(.din(w_dff_B_aHqIICak1_2),.dout(w_dff_B_BiD5EdXq3_2),.clk(gclk));
	jdff dff_B_FwBDmWms0_1(.din(n942),.dout(w_dff_B_FwBDmWms0_1),.clk(gclk));
	jdff dff_B_9Xrlp8t79_1(.din(w_dff_B_FwBDmWms0_1),.dout(w_dff_B_9Xrlp8t79_1),.clk(gclk));
	jdff dff_B_FLk7yXTK9_1(.din(w_dff_B_9Xrlp8t79_1),.dout(w_dff_B_FLk7yXTK9_1),.clk(gclk));
	jdff dff_B_I6hnxsZq9_1(.din(n947),.dout(w_dff_B_I6hnxsZq9_1),.clk(gclk));
	jdff dff_B_dSMLp7Iu5_1(.din(w_dff_B_I6hnxsZq9_1),.dout(w_dff_B_dSMLp7Iu5_1),.clk(gclk));
	jdff dff_B_aGPEn6zR7_1(.din(n955),.dout(w_dff_B_aGPEn6zR7_1),.clk(gclk));
	jdff dff_B_DxRhincp4_1(.din(n956),.dout(w_dff_B_DxRhincp4_1),.clk(gclk));
	jdff dff_B_5hBGFDgg4_1(.din(n957),.dout(w_dff_B_5hBGFDgg4_1),.clk(gclk));
	jdff dff_B_lMCtFf5v0_1(.din(w_dff_B_5hBGFDgg4_1),.dout(w_dff_B_lMCtFf5v0_1),.clk(gclk));
	jdff dff_B_Hs2jrfC70_1(.din(w_dff_B_lMCtFf5v0_1),.dout(w_dff_B_Hs2jrfC70_1),.clk(gclk));
	jdff dff_B_Cc4JLWJc2_1(.din(w_dff_B_Hs2jrfC70_1),.dout(w_dff_B_Cc4JLWJc2_1),.clk(gclk));
	jdff dff_B_pastvOPG7_0(.din(n976),.dout(w_dff_B_pastvOPG7_0),.clk(gclk));
	jdff dff_B_PlStXqfk4_0(.din(w_dff_B_pastvOPG7_0),.dout(w_dff_B_PlStXqfk4_0),.clk(gclk));
	jdff dff_B_TxdIXZpt4_0(.din(n995),.dout(w_dff_B_TxdIXZpt4_0),.clk(gclk));
	jdff dff_B_2u3sRBDv6_0(.din(w_dff_B_TxdIXZpt4_0),.dout(w_dff_B_2u3sRBDv6_0),.clk(gclk));
	jdff dff_B_dZxZuFOa6_0(.din(n994),.dout(w_dff_B_dZxZuFOa6_0),.clk(gclk));
	jdff dff_B_za3o7y3d3_0(.din(w_dff_B_dZxZuFOa6_0),.dout(w_dff_B_za3o7y3d3_0),.clk(gclk));
	jdff dff_B_8Q2p3NVF7_0(.din(w_dff_B_za3o7y3d3_0),.dout(w_dff_B_8Q2p3NVF7_0),.clk(gclk));
	jdff dff_B_tOz9RWR58_0(.din(w_dff_B_8Q2p3NVF7_0),.dout(w_dff_B_tOz9RWR58_0),.clk(gclk));
	jdff dff_B_4xQBvl2r0_0(.din(n993),.dout(w_dff_B_4xQBvl2r0_0),.clk(gclk));
	jdff dff_B_lXhl7vWC1_0(.din(n1009),.dout(w_dff_B_lXhl7vWC1_0),.clk(gclk));
	jdff dff_B_KpZXeaHc9_0(.din(w_dff_B_lXhl7vWC1_0),.dout(w_dff_B_KpZXeaHc9_0),.clk(gclk));
	jdff dff_B_qC6oRdRK1_0(.din(n1008),.dout(w_dff_B_qC6oRdRK1_0),.clk(gclk));
	jdff dff_B_e0WHgypv3_0(.din(w_dff_B_qC6oRdRK1_0),.dout(w_dff_B_e0WHgypv3_0),.clk(gclk));
	jdff dff_B_sZWv7KcA3_0(.din(w_dff_B_e0WHgypv3_0),.dout(w_dff_B_sZWv7KcA3_0),.clk(gclk));
	jdff dff_B_IB2lwABJ2_0(.din(w_dff_B_sZWv7KcA3_0),.dout(w_dff_B_IB2lwABJ2_0),.clk(gclk));
	jdff dff_B_Slzp9vaC8_0(.din(n1007),.dout(w_dff_B_Slzp9vaC8_0),.clk(gclk));
	jdff dff_B_8Yt5X2SC2_2(.din(G185),.dout(w_dff_B_8Yt5X2SC2_2),.clk(gclk));
	jdff dff_B_f8KbmwrY8_2(.din(G182),.dout(w_dff_B_f8KbmwrY8_2),.clk(gclk));
	jdff dff_B_y7pSZth39_2(.din(w_dff_B_f8KbmwrY8_2),.dout(w_dff_B_y7pSZth39_2),.clk(gclk));
	jdff dff_B_eSJT5Mt21_1(.din(n749),.dout(w_dff_B_eSJT5Mt21_1),.clk(gclk));
	jdff dff_B_Vtl8R2nH1_1(.din(G131),.dout(w_dff_B_Vtl8R2nH1_1),.clk(gclk));
	jdff dff_B_26hfeWVD4_1(.din(w_dff_B_Vtl8R2nH1_1),.dout(w_dff_B_26hfeWVD4_1),.clk(gclk));
	jdff dff_B_2OZpruAF3_0(.din(n777),.dout(w_dff_B_2OZpruAF3_0),.clk(gclk));
	jdff dff_B_nYzCmORx9_1(.din(n774),.dout(w_dff_B_nYzCmORx9_1),.clk(gclk));
	jdff dff_B_gyx2IgSc9_1(.din(G117),.dout(w_dff_B_gyx2IgSc9_1),.clk(gclk));
	jdff dff_B_gMgEU3kz8_1(.din(w_dff_B_gyx2IgSc9_1),.dout(w_dff_B_gMgEU3kz8_1),.clk(gclk));
	jdff dff_B_1pMomV046_0(.din(n503),.dout(w_dff_B_1pMomV046_0),.clk(gclk));
	jdff dff_B_Mw9bT7h82_0(.din(n1019),.dout(w_dff_B_Mw9bT7h82_0),.clk(gclk));
	jdff dff_B_WWtYwvnd6_0(.din(w_dff_B_Mw9bT7h82_0),.dout(w_dff_B_WWtYwvnd6_0),.clk(gclk));
	jdff dff_B_jLsh2peL3_0(.din(w_dff_B_WWtYwvnd6_0),.dout(w_dff_B_jLsh2peL3_0),.clk(gclk));
	jdff dff_B_TBw81uok5_0(.din(w_dff_B_jLsh2peL3_0),.dout(w_dff_B_TBw81uok5_0),.clk(gclk));
	jdff dff_B_JVjiMPN85_0(.din(n1018),.dout(w_dff_B_JVjiMPN85_0),.clk(gclk));
	jdff dff_B_X97uTZ773_0(.din(w_dff_B_JVjiMPN85_0),.dout(w_dff_B_X97uTZ773_0),.clk(gclk));
	jdff dff_B_goH244bY6_0(.din(w_dff_B_X97uTZ773_0),.dout(w_dff_B_goH244bY6_0),.clk(gclk));
	jdff dff_B_G8RuqwgS0_0(.din(w_dff_B_goH244bY6_0),.dout(w_dff_B_G8RuqwgS0_0),.clk(gclk));
	jdff dff_B_Aaqk6xgn3_0(.din(w_dff_B_G8RuqwgS0_0),.dout(w_dff_B_Aaqk6xgn3_0),.clk(gclk));
	jdff dff_B_hjjrRSHq0_0(.din(w_dff_B_Aaqk6xgn3_0),.dout(w_dff_B_hjjrRSHq0_0),.clk(gclk));
	jdff dff_B_QwYmrZtN6_0(.din(w_dff_B_hjjrRSHq0_0),.dout(w_dff_B_QwYmrZtN6_0),.clk(gclk));
	jdff dff_B_yzh2W3DX2_0(.din(n1017),.dout(w_dff_B_yzh2W3DX2_0),.clk(gclk));
	jdff dff_A_VAD0TqVh9_0(.dout(w_n797_4[0]),.din(w_dff_A_VAD0TqVh9_0),.clk(gclk));
	jdff dff_A_4h6dq7J39_0(.dout(w_dff_A_VAD0TqVh9_0),.din(w_dff_A_4h6dq7J39_0),.clk(gclk));
	jdff dff_A_Izq4Ek8W1_0(.dout(w_dff_A_4h6dq7J39_0),.din(w_dff_A_Izq4Ek8W1_0),.clk(gclk));
	jdff dff_A_rFYTqiN56_0(.dout(w_n793_4[0]),.din(w_dff_A_rFYTqiN56_0),.clk(gclk));
	jdff dff_A_Q5vjTzVR8_0(.dout(w_dff_A_rFYTqiN56_0),.din(w_dff_A_Q5vjTzVR8_0),.clk(gclk));
	jdff dff_A_Vk6xNNQ11_0(.dout(w_dff_A_Q5vjTzVR8_0),.din(w_dff_A_Vk6xNNQ11_0),.clk(gclk));
	jdff dff_A_xdg5shdo1_0(.dout(w_dff_A_Vk6xNNQ11_0),.din(w_dff_A_xdg5shdo1_0),.clk(gclk));
	jdff dff_A_ZCK0Bsrp4_0(.dout(w_dff_A_xdg5shdo1_0),.din(w_dff_A_ZCK0Bsrp4_0),.clk(gclk));
	jdff dff_B_Gx18M9zT8_0(.din(n1028),.dout(w_dff_B_Gx18M9zT8_0),.clk(gclk));
	jdff dff_B_3yp9MbZK8_0(.din(w_dff_B_Gx18M9zT8_0),.dout(w_dff_B_3yp9MbZK8_0),.clk(gclk));
	jdff dff_B_pBpLQpd10_0(.din(w_dff_B_3yp9MbZK8_0),.dout(w_dff_B_pBpLQpd10_0),.clk(gclk));
	jdff dff_B_SYCIhiJY9_0(.din(w_dff_B_pBpLQpd10_0),.dout(w_dff_B_SYCIhiJY9_0),.clk(gclk));
	jdff dff_B_7I729Ujb7_0(.din(n1027),.dout(w_dff_B_7I729Ujb7_0),.clk(gclk));
	jdff dff_B_2uBfnEDK1_0(.din(w_dff_B_7I729Ujb7_0),.dout(w_dff_B_2uBfnEDK1_0),.clk(gclk));
	jdff dff_B_5ouMzg7U1_0(.din(w_dff_B_2uBfnEDK1_0),.dout(w_dff_B_5ouMzg7U1_0),.clk(gclk));
	jdff dff_B_8cuKNfSZ2_0(.din(w_dff_B_5ouMzg7U1_0),.dout(w_dff_B_8cuKNfSZ2_0),.clk(gclk));
	jdff dff_B_LnPLsUzR2_0(.din(w_dff_B_8cuKNfSZ2_0),.dout(w_dff_B_LnPLsUzR2_0),.clk(gclk));
	jdff dff_B_0l4ExStx1_0(.din(w_dff_B_LnPLsUzR2_0),.dout(w_dff_B_0l4ExStx1_0),.clk(gclk));
	jdff dff_B_EFOHvvMd4_0(.din(n1026),.dout(w_dff_B_EFOHvvMd4_0),.clk(gclk));
	jdff dff_B_khimyeJF9_0(.din(n1037),.dout(w_dff_B_khimyeJF9_0),.clk(gclk));
	jdff dff_B_AdtNkSCw9_0(.din(w_dff_B_khimyeJF9_0),.dout(w_dff_B_AdtNkSCw9_0),.clk(gclk));
	jdff dff_B_MaPgAzdj1_0(.din(w_dff_B_AdtNkSCw9_0),.dout(w_dff_B_MaPgAzdj1_0),.clk(gclk));
	jdff dff_B_CTXroHMd3_0(.din(w_dff_B_MaPgAzdj1_0),.dout(w_dff_B_CTXroHMd3_0),.clk(gclk));
	jdff dff_B_J6wrzi0i8_0(.din(n1036),.dout(w_dff_B_J6wrzi0i8_0),.clk(gclk));
	jdff dff_B_RYV23nIl2_0(.din(w_dff_B_J6wrzi0i8_0),.dout(w_dff_B_RYV23nIl2_0),.clk(gclk));
	jdff dff_B_eZrPI4Qr5_0(.din(w_dff_B_RYV23nIl2_0),.dout(w_dff_B_eZrPI4Qr5_0),.clk(gclk));
	jdff dff_B_KIUWV3WE9_0(.din(w_dff_B_eZrPI4Qr5_0),.dout(w_dff_B_KIUWV3WE9_0),.clk(gclk));
	jdff dff_B_5gEmHFrd6_0(.din(w_dff_B_KIUWV3WE9_0),.dout(w_dff_B_5gEmHFrd6_0),.clk(gclk));
	jdff dff_B_Lr4O21im4_0(.din(w_dff_B_5gEmHFrd6_0),.dout(w_dff_B_Lr4O21im4_0),.clk(gclk));
	jdff dff_B_1C1cxjdS6_0(.din(n1035),.dout(w_dff_B_1C1cxjdS6_0),.clk(gclk));
	jdff dff_B_oY8yNrqq5_0(.din(n1046),.dout(w_dff_B_oY8yNrqq5_0),.clk(gclk));
	jdff dff_B_8heiXQ8D1_0(.din(w_dff_B_oY8yNrqq5_0),.dout(w_dff_B_8heiXQ8D1_0),.clk(gclk));
	jdff dff_B_twzCbOZs0_0(.din(w_dff_B_8heiXQ8D1_0),.dout(w_dff_B_twzCbOZs0_0),.clk(gclk));
	jdff dff_B_2A9yH7yX5_0(.din(w_dff_B_twzCbOZs0_0),.dout(w_dff_B_2A9yH7yX5_0),.clk(gclk));
	jdff dff_B_c8kVFgYn3_0(.din(w_dff_B_2A9yH7yX5_0),.dout(w_dff_B_c8kVFgYn3_0),.clk(gclk));
	jdff dff_B_iFytHTv26_0(.din(n1045),.dout(w_dff_B_iFytHTv26_0),.clk(gclk));
	jdff dff_B_LQ9cAgVa6_0(.din(w_dff_B_iFytHTv26_0),.dout(w_dff_B_LQ9cAgVa6_0),.clk(gclk));
	jdff dff_B_MjDqlfFb8_0(.din(w_dff_B_LQ9cAgVa6_0),.dout(w_dff_B_MjDqlfFb8_0),.clk(gclk));
	jdff dff_B_5ETUfBtl6_0(.din(w_dff_B_MjDqlfFb8_0),.dout(w_dff_B_5ETUfBtl6_0),.clk(gclk));
	jdff dff_B_XCdzVBk76_0(.din(w_dff_B_5ETUfBtl6_0),.dout(w_dff_B_XCdzVBk76_0),.clk(gclk));
	jdff dff_B_Yr3r80KN9_0(.din(n1044),.dout(w_dff_B_Yr3r80KN9_0),.clk(gclk));
	jdff dff_A_wcEwDFX14_1(.dout(w_n797_3[1]),.din(w_dff_A_wcEwDFX14_1),.clk(gclk));
	jdff dff_A_okWsnYcW0_2(.dout(w_n797_3[2]),.din(w_dff_A_okWsnYcW0_2),.clk(gclk));
	jdff dff_B_xtW8R4l04_0(.din(n1053),.dout(w_dff_B_xtW8R4l04_0),.clk(gclk));
	jdff dff_B_Hqj2BGyl6_0(.din(w_dff_B_xtW8R4l04_0),.dout(w_dff_B_Hqj2BGyl6_0),.clk(gclk));
	jdff dff_B_jJSd5e4E3_0(.din(w_dff_B_Hqj2BGyl6_0),.dout(w_dff_B_jJSd5e4E3_0),.clk(gclk));
	jdff dff_B_oef3wOMR0_0(.din(w_dff_B_jJSd5e4E3_0),.dout(w_dff_B_oef3wOMR0_0),.clk(gclk));
	jdff dff_B_9JNPfFuv2_0(.din(n1052),.dout(w_dff_B_9JNPfFuv2_0),.clk(gclk));
	jdff dff_B_vwqSx1125_0(.din(w_dff_B_9JNPfFuv2_0),.dout(w_dff_B_vwqSx1125_0),.clk(gclk));
	jdff dff_B_VVhxjbwL1_0(.din(w_dff_B_vwqSx1125_0),.dout(w_dff_B_VVhxjbwL1_0),.clk(gclk));
	jdff dff_B_ElcNvPpo7_0(.din(w_dff_B_VVhxjbwL1_0),.dout(w_dff_B_ElcNvPpo7_0),.clk(gclk));
	jdff dff_B_ng7hVfxZ8_0(.din(w_dff_B_ElcNvPpo7_0),.dout(w_dff_B_ng7hVfxZ8_0),.clk(gclk));
	jdff dff_B_a3Ht3qBZ7_0(.din(w_dff_B_ng7hVfxZ8_0),.dout(w_dff_B_a3Ht3qBZ7_0),.clk(gclk));
	jdff dff_B_cQsrr4c32_0(.din(w_dff_B_a3Ht3qBZ7_0),.dout(w_dff_B_cQsrr4c32_0),.clk(gclk));
	jdff dff_B_pW89VdJt3_0(.din(n1051),.dout(w_dff_B_pW89VdJt3_0),.clk(gclk));
	jdff dff_B_xxhTC5x54_2(.din(G37),.dout(w_dff_B_xxhTC5x54_2),.clk(gclk));
	jdff dff_B_W2UJTWXX5_2(.din(G43),.dout(w_dff_B_W2UJTWXX5_2),.clk(gclk));
	jdff dff_B_jwtZKyDM4_2(.din(w_dff_B_W2UJTWXX5_2),.dout(w_dff_B_jwtZKyDM4_2),.clk(gclk));
	jdff dff_A_3wxzoUkB3_0(.dout(w_n843_4[0]),.din(w_dff_A_3wxzoUkB3_0),.clk(gclk));
	jdff dff_A_NwY7EWSI2_0(.dout(w_dff_A_3wxzoUkB3_0),.din(w_dff_A_NwY7EWSI2_0),.clk(gclk));
	jdff dff_A_jbpOdlvy3_0(.dout(w_dff_A_NwY7EWSI2_0),.din(w_dff_A_jbpOdlvy3_0),.clk(gclk));
	jdff dff_A_KRCB5eEO6_0(.dout(w_n840_4[0]),.din(w_dff_A_KRCB5eEO6_0),.clk(gclk));
	jdff dff_A_E6neABW57_0(.dout(w_dff_A_KRCB5eEO6_0),.din(w_dff_A_E6neABW57_0),.clk(gclk));
	jdff dff_A_ZEZKEdrn9_0(.dout(w_dff_A_E6neABW57_0),.din(w_dff_A_ZEZKEdrn9_0),.clk(gclk));
	jdff dff_A_U9CsHbJj0_0(.dout(w_dff_A_ZEZKEdrn9_0),.din(w_dff_A_U9CsHbJj0_0),.clk(gclk));
	jdff dff_A_fGW91Ct89_0(.dout(w_dff_A_U9CsHbJj0_0),.din(w_dff_A_fGW91Ct89_0),.clk(gclk));
	jdff dff_B_idkaQGLg2_0(.din(n1060),.dout(w_dff_B_idkaQGLg2_0),.clk(gclk));
	jdff dff_B_BgSD60qq6_0(.din(w_dff_B_idkaQGLg2_0),.dout(w_dff_B_BgSD60qq6_0),.clk(gclk));
	jdff dff_B_jHgNWtvc9_0(.din(w_dff_B_BgSD60qq6_0),.dout(w_dff_B_jHgNWtvc9_0),.clk(gclk));
	jdff dff_B_wNxtMbtO6_0(.din(w_dff_B_jHgNWtvc9_0),.dout(w_dff_B_wNxtMbtO6_0),.clk(gclk));
	jdff dff_B_YnJ1Yh5H7_0(.din(n1059),.dout(w_dff_B_YnJ1Yh5H7_0),.clk(gclk));
	jdff dff_B_F0gT7RyK7_0(.din(w_dff_B_YnJ1Yh5H7_0),.dout(w_dff_B_F0gT7RyK7_0),.clk(gclk));
	jdff dff_B_QXDjpZVM0_0(.din(w_dff_B_F0gT7RyK7_0),.dout(w_dff_B_QXDjpZVM0_0),.clk(gclk));
	jdff dff_B_kmRSgUaW3_0(.din(w_dff_B_QXDjpZVM0_0),.dout(w_dff_B_kmRSgUaW3_0),.clk(gclk));
	jdff dff_B_YQI6wa8Z8_0(.din(w_dff_B_kmRSgUaW3_0),.dout(w_dff_B_YQI6wa8Z8_0),.clk(gclk));
	jdff dff_B_TNC4Qb987_0(.din(w_dff_B_YQI6wa8Z8_0),.dout(w_dff_B_TNC4Qb987_0),.clk(gclk));
	jdff dff_B_GaCqMgtu1_0(.din(n1058),.dout(w_dff_B_GaCqMgtu1_0),.clk(gclk));
	jdff dff_B_8T3VWiob3_2(.din(G20),.dout(w_dff_B_8T3VWiob3_2),.clk(gclk));
	jdff dff_B_xTwIwzGE1_2(.din(G76),.dout(w_dff_B_xTwIwzGE1_2),.clk(gclk));
	jdff dff_B_hl6lL76m7_2(.din(w_dff_B_xTwIwzGE1_2),.dout(w_dff_B_hl6lL76m7_2),.clk(gclk));
	jdff dff_B_OTb1d4NB6_0(.din(n1067),.dout(w_dff_B_OTb1d4NB6_0),.clk(gclk));
	jdff dff_B_02LvlSIN4_0(.din(w_dff_B_OTb1d4NB6_0),.dout(w_dff_B_02LvlSIN4_0),.clk(gclk));
	jdff dff_B_2jnld2Lr1_0(.din(w_dff_B_02LvlSIN4_0),.dout(w_dff_B_2jnld2Lr1_0),.clk(gclk));
	jdff dff_B_59nKBC3D3_0(.din(w_dff_B_2jnld2Lr1_0),.dout(w_dff_B_59nKBC3D3_0),.clk(gclk));
	jdff dff_B_iy8RiUN58_0(.din(n1066),.dout(w_dff_B_iy8RiUN58_0),.clk(gclk));
	jdff dff_B_7NWbyQmR1_0(.din(w_dff_B_iy8RiUN58_0),.dout(w_dff_B_7NWbyQmR1_0),.clk(gclk));
	jdff dff_B_yloQAErT0_0(.din(w_dff_B_7NWbyQmR1_0),.dout(w_dff_B_yloQAErT0_0),.clk(gclk));
	jdff dff_B_Daw1tBii1_0(.din(w_dff_B_yloQAErT0_0),.dout(w_dff_B_Daw1tBii1_0),.clk(gclk));
	jdff dff_B_k9DmYLW29_0(.din(w_dff_B_Daw1tBii1_0),.dout(w_dff_B_k9DmYLW29_0),.clk(gclk));
	jdff dff_B_JurtH47K4_0(.din(w_dff_B_k9DmYLW29_0),.dout(w_dff_B_JurtH47K4_0),.clk(gclk));
	jdff dff_B_9FV3cLIM8_0(.din(n1065),.dout(w_dff_B_9FV3cLIM8_0),.clk(gclk));
	jdff dff_B_933tUGNJ1_2(.din(G17),.dout(w_dff_B_933tUGNJ1_2),.clk(gclk));
	jdff dff_B_yoWYvQti6_2(.din(G73),.dout(w_dff_B_yoWYvQti6_2),.clk(gclk));
	jdff dff_B_9UiXsHup0_2(.din(w_dff_B_yoWYvQti6_2),.dout(w_dff_B_9UiXsHup0_2),.clk(gclk));
	jdff dff_B_Rlcf1GDx5_0(.din(n1074),.dout(w_dff_B_Rlcf1GDx5_0),.clk(gclk));
	jdff dff_B_XDV9kWAm9_0(.din(w_dff_B_Rlcf1GDx5_0),.dout(w_dff_B_XDV9kWAm9_0),.clk(gclk));
	jdff dff_B_qBWSZGAX7_0(.din(w_dff_B_XDV9kWAm9_0),.dout(w_dff_B_qBWSZGAX7_0),.clk(gclk));
	jdff dff_B_brjs7dzY8_0(.din(w_dff_B_qBWSZGAX7_0),.dout(w_dff_B_brjs7dzY8_0),.clk(gclk));
	jdff dff_B_Wv0NtsIA4_0(.din(w_dff_B_brjs7dzY8_0),.dout(w_dff_B_Wv0NtsIA4_0),.clk(gclk));
	jdff dff_B_l5Uh0TeI7_0(.din(n1073),.dout(w_dff_B_l5Uh0TeI7_0),.clk(gclk));
	jdff dff_B_r48g0MKq6_0(.din(w_dff_B_l5Uh0TeI7_0),.dout(w_dff_B_r48g0MKq6_0),.clk(gclk));
	jdff dff_B_8aRDAa4P7_0(.din(w_dff_B_r48g0MKq6_0),.dout(w_dff_B_8aRDAa4P7_0),.clk(gclk));
	jdff dff_B_nNKbKmfi0_0(.din(w_dff_B_8aRDAa4P7_0),.dout(w_dff_B_nNKbKmfi0_0),.clk(gclk));
	jdff dff_B_wBIa7dao0_0(.din(w_dff_B_nNKbKmfi0_0),.dout(w_dff_B_wBIa7dao0_0),.clk(gclk));
	jdff dff_B_mvLIU5Ui7_0(.din(n1072),.dout(w_dff_B_mvLIU5Ui7_0),.clk(gclk));
	jdff dff_B_evZZUxAQ6_2(.din(G70),.dout(w_dff_B_evZZUxAQ6_2),.clk(gclk));
	jdff dff_B_Sr0Z6q3F9_2(.din(G67),.dout(w_dff_B_Sr0Z6q3F9_2),.clk(gclk));
	jdff dff_B_ebTHCX9D8_2(.din(w_dff_B_Sr0Z6q3F9_2),.dout(w_dff_B_ebTHCX9D8_2),.clk(gclk));
	jdff dff_A_9OgRyhsy3_1(.dout(w_n843_3[1]),.din(w_dff_A_9OgRyhsy3_1),.clk(gclk));
	jdff dff_A_X0jYu4GN5_2(.dout(w_n843_3[2]),.din(w_dff_A_X0jYu4GN5_2),.clk(gclk));
	jdff dff_B_De6HjeTr5_0(.din(n1081),.dout(w_dff_B_De6HjeTr5_0),.clk(gclk));
	jdff dff_B_1pC0sKdg5_0(.din(w_dff_B_De6HjeTr5_0),.dout(w_dff_B_1pC0sKdg5_0),.clk(gclk));
	jdff dff_B_JFXFQfai5_0(.din(w_dff_B_1pC0sKdg5_0),.dout(w_dff_B_JFXFQfai5_0),.clk(gclk));
	jdff dff_B_1IWmYF6w0_0(.din(w_dff_B_JFXFQfai5_0),.dout(w_dff_B_1IWmYF6w0_0),.clk(gclk));
	jdff dff_B_7p7zo9qH2_0(.din(n1080),.dout(w_dff_B_7p7zo9qH2_0),.clk(gclk));
	jdff dff_B_AfJ0b24G1_0(.din(w_dff_B_7p7zo9qH2_0),.dout(w_dff_B_AfJ0b24G1_0),.clk(gclk));
	jdff dff_B_gwLsbmn47_0(.din(w_dff_B_AfJ0b24G1_0),.dout(w_dff_B_gwLsbmn47_0),.clk(gclk));
	jdff dff_B_gfgEgEin8_0(.din(w_dff_B_gwLsbmn47_0),.dout(w_dff_B_gfgEgEin8_0),.clk(gclk));
	jdff dff_B_BkkvnJa04_0(.din(w_dff_B_gfgEgEin8_0),.dout(w_dff_B_BkkvnJa04_0),.clk(gclk));
	jdff dff_B_pi3bOMe96_0(.din(w_dff_B_BkkvnJa04_0),.dout(w_dff_B_pi3bOMe96_0),.clk(gclk));
	jdff dff_B_Gf4T2pe65_0(.din(w_dff_B_pi3bOMe96_0),.dout(w_dff_B_Gf4T2pe65_0),.clk(gclk));
	jdff dff_B_1b6BJ2b44_0(.din(n1079),.dout(w_dff_B_1b6BJ2b44_0),.clk(gclk));
	jdff dff_A_Ga6sOL0g0_0(.dout(w_n988_4[0]),.din(w_dff_A_Ga6sOL0g0_0),.clk(gclk));
	jdff dff_A_AmZchLaN3_0(.dout(w_dff_A_Ga6sOL0g0_0),.din(w_dff_A_AmZchLaN3_0),.clk(gclk));
	jdff dff_A_5DV6LkPy1_0(.dout(w_dff_A_AmZchLaN3_0),.din(w_dff_A_5DV6LkPy1_0),.clk(gclk));
	jdff dff_A_bB5nYlHV7_0(.dout(w_n985_4[0]),.din(w_dff_A_bB5nYlHV7_0),.clk(gclk));
	jdff dff_A_lTP63Spd9_0(.dout(w_dff_A_bB5nYlHV7_0),.din(w_dff_A_lTP63Spd9_0),.clk(gclk));
	jdff dff_A_YDMzKWpx9_0(.dout(w_dff_A_lTP63Spd9_0),.din(w_dff_A_YDMzKWpx9_0),.clk(gclk));
	jdff dff_A_QD945d3m7_0(.dout(w_dff_A_YDMzKWpx9_0),.din(w_dff_A_QD945d3m7_0),.clk(gclk));
	jdff dff_A_lbsv0ReK6_0(.dout(w_dff_A_QD945d3m7_0),.din(w_dff_A_lbsv0ReK6_0),.clk(gclk));
	jdff dff_B_c86NDLmv7_0(.din(n1089),.dout(w_dff_B_c86NDLmv7_0),.clk(gclk));
	jdff dff_B_llIEBgxY1_0(.din(w_dff_B_c86NDLmv7_0),.dout(w_dff_B_llIEBgxY1_0),.clk(gclk));
	jdff dff_B_mgGvZFKz3_0(.din(w_dff_B_llIEBgxY1_0),.dout(w_dff_B_mgGvZFKz3_0),.clk(gclk));
	jdff dff_B_DKuPd3Q95_0(.din(w_dff_B_mgGvZFKz3_0),.dout(w_dff_B_DKuPd3Q95_0),.clk(gclk));
	jdff dff_B_x8TsiQby5_0(.din(w_dff_B_DKuPd3Q95_0),.dout(w_dff_B_x8TsiQby5_0),.clk(gclk));
	jdff dff_B_WY0rg8lq3_0(.din(n1088),.dout(w_dff_B_WY0rg8lq3_0),.clk(gclk));
	jdff dff_B_N8nNB1em7_0(.din(w_dff_B_WY0rg8lq3_0),.dout(w_dff_B_N8nNB1em7_0),.clk(gclk));
	jdff dff_B_wgb1a7W06_0(.din(w_dff_B_N8nNB1em7_0),.dout(w_dff_B_wgb1a7W06_0),.clk(gclk));
	jdff dff_B_SjL1xJhq7_0(.din(w_dff_B_wgb1a7W06_0),.dout(w_dff_B_SjL1xJhq7_0),.clk(gclk));
	jdff dff_B_fXQYtvhd2_0(.din(w_dff_B_SjL1xJhq7_0),.dout(w_dff_B_fXQYtvhd2_0),.clk(gclk));
	jdff dff_B_Pwkrnbqn8_0(.din(n1087),.dout(w_dff_B_Pwkrnbqn8_0),.clk(gclk));
	jdff dff_B_mPKyzr5A0_0(.din(n1097),.dout(w_dff_B_mPKyzr5A0_0),.clk(gclk));
	jdff dff_B_OmmcV7zM7_0(.din(w_dff_B_mPKyzr5A0_0),.dout(w_dff_B_OmmcV7zM7_0),.clk(gclk));
	jdff dff_B_8uskkqVH8_0(.din(w_dff_B_OmmcV7zM7_0),.dout(w_dff_B_8uskkqVH8_0),.clk(gclk));
	jdff dff_B_9GS9SIJm4_0(.din(w_dff_B_8uskkqVH8_0),.dout(w_dff_B_9GS9SIJm4_0),.clk(gclk));
	jdff dff_B_BxP2vLRX4_0(.din(n1096),.dout(w_dff_B_BxP2vLRX4_0),.clk(gclk));
	jdff dff_B_bfCgYGGY8_0(.din(w_dff_B_BxP2vLRX4_0),.dout(w_dff_B_bfCgYGGY8_0),.clk(gclk));
	jdff dff_B_XBCxwza53_0(.din(w_dff_B_bfCgYGGY8_0),.dout(w_dff_B_XBCxwza53_0),.clk(gclk));
	jdff dff_B_7z8UO4ak4_0(.din(w_dff_B_XBCxwza53_0),.dout(w_dff_B_7z8UO4ak4_0),.clk(gclk));
	jdff dff_B_TMykp1pR1_0(.din(w_dff_B_7z8UO4ak4_0),.dout(w_dff_B_TMykp1pR1_0),.clk(gclk));
	jdff dff_B_o59bURzk6_0(.din(w_dff_B_TMykp1pR1_0),.dout(w_dff_B_o59bURzk6_0),.clk(gclk));
	jdff dff_B_C4GUCiLi4_0(.din(n1095),.dout(w_dff_B_C4GUCiLi4_0),.clk(gclk));
	jdff dff_A_etCgCDAc9_2(.dout(w_G137_8[2]),.din(w_dff_A_etCgCDAc9_2),.clk(gclk));
	jdff dff_B_QXbdTfSC4_0(.din(n1105),.dout(w_dff_B_QXbdTfSC4_0),.clk(gclk));
	jdff dff_B_yDMjWOG83_0(.din(w_dff_B_QXbdTfSC4_0),.dout(w_dff_B_yDMjWOG83_0),.clk(gclk));
	jdff dff_B_A7VHVmSN2_0(.din(w_dff_B_yDMjWOG83_0),.dout(w_dff_B_A7VHVmSN2_0),.clk(gclk));
	jdff dff_B_FJNmdIq07_0(.din(w_dff_B_A7VHVmSN2_0),.dout(w_dff_B_FJNmdIq07_0),.clk(gclk));
	jdff dff_B_KEzPG80v8_0(.din(n1104),.dout(w_dff_B_KEzPG80v8_0),.clk(gclk));
	jdff dff_B_Z3nKmgEY0_0(.din(w_dff_B_KEzPG80v8_0),.dout(w_dff_B_Z3nKmgEY0_0),.clk(gclk));
	jdff dff_B_yPKn7UWd1_0(.din(w_dff_B_Z3nKmgEY0_0),.dout(w_dff_B_yPKn7UWd1_0),.clk(gclk));
	jdff dff_B_HDBGGIma9_0(.din(w_dff_B_yPKn7UWd1_0),.dout(w_dff_B_HDBGGIma9_0),.clk(gclk));
	jdff dff_B_gh5w2VDO3_0(.din(w_dff_B_HDBGGIma9_0),.dout(w_dff_B_gh5w2VDO3_0),.clk(gclk));
	jdff dff_B_1CYes5n85_0(.din(w_dff_B_gh5w2VDO3_0),.dout(w_dff_B_1CYes5n85_0),.clk(gclk));
	jdff dff_B_JcqG57Ro5_0(.din(n1103),.dout(w_dff_B_JcqG57Ro5_0),.clk(gclk));
	jdff dff_A_r7GzCRg66_0(.dout(w_n988_3[0]),.din(w_dff_A_r7GzCRg66_0),.clk(gclk));
	jdff dff_A_uLwnQKui8_1(.dout(w_n988_3[1]),.din(w_dff_A_uLwnQKui8_1),.clk(gclk));
	jdff dff_B_SbPu66re4_0(.din(n1113),.dout(w_dff_B_SbPu66re4_0),.clk(gclk));
	jdff dff_B_Zf9fuJPj0_0(.din(w_dff_B_SbPu66re4_0),.dout(w_dff_B_Zf9fuJPj0_0),.clk(gclk));
	jdff dff_B_2YVle0hT3_0(.din(w_dff_B_Zf9fuJPj0_0),.dout(w_dff_B_2YVle0hT3_0),.clk(gclk));
	jdff dff_B_43EMR9wJ7_0(.din(w_dff_B_2YVle0hT3_0),.dout(w_dff_B_43EMR9wJ7_0),.clk(gclk));
	jdff dff_B_dTkXopeo5_0(.din(n1112),.dout(w_dff_B_dTkXopeo5_0),.clk(gclk));
	jdff dff_B_8kSi8rGV7_0(.din(w_dff_B_dTkXopeo5_0),.dout(w_dff_B_8kSi8rGV7_0),.clk(gclk));
	jdff dff_B_uMNth0T19_0(.din(w_dff_B_8kSi8rGV7_0),.dout(w_dff_B_uMNth0T19_0),.clk(gclk));
	jdff dff_B_bTZDVqR75_0(.din(w_dff_B_uMNth0T19_0),.dout(w_dff_B_bTZDVqR75_0),.clk(gclk));
	jdff dff_B_wkyzqvan1_0(.din(w_dff_B_bTZDVqR75_0),.dout(w_dff_B_wkyzqvan1_0),.clk(gclk));
	jdff dff_B_7IdryhxC2_0(.din(w_dff_B_wkyzqvan1_0),.dout(w_dff_B_7IdryhxC2_0),.clk(gclk));
	jdff dff_B_c47yMk2V7_0(.din(w_dff_B_7IdryhxC2_0),.dout(w_dff_B_c47yMk2V7_0),.clk(gclk));
	jdff dff_B_tRGiG3Pb4_0(.din(n1111),.dout(w_dff_B_tRGiG3Pb4_0),.clk(gclk));
	jdff dff_B_IHVmLyWb3_2(.din(G170),.dout(w_dff_B_IHVmLyWb3_2),.clk(gclk));
	jdff dff_B_UaLU43c64_2(.din(G200),.dout(w_dff_B_UaLU43c64_2),.clk(gclk));
	jdff dff_B_NPBlv3NP1_2(.din(w_dff_B_UaLU43c64_2),.dout(w_dff_B_NPBlv3NP1_2),.clk(gclk));
	jdff dff_A_LpkRCZlm5_0(.dout(w_n1002_4[0]),.din(w_dff_A_LpkRCZlm5_0),.clk(gclk));
	jdff dff_A_1Rm34mUJ6_0(.dout(w_dff_A_LpkRCZlm5_0),.din(w_dff_A_1Rm34mUJ6_0),.clk(gclk));
	jdff dff_A_TExLgcsK5_0(.dout(w_dff_A_1Rm34mUJ6_0),.din(w_dff_A_TExLgcsK5_0),.clk(gclk));
	jdff dff_B_z2ueqf6J2_0(.din(n814),.dout(w_dff_B_z2ueqf6J2_0),.clk(gclk));
	jdff dff_B_RP8ZKKAf4_0(.din(w_dff_B_z2ueqf6J2_0),.dout(w_dff_B_RP8ZKKAf4_0),.clk(gclk));
	jdff dff_B_mZBKS0aB4_1(.din(n811),.dout(w_dff_B_mZBKS0aB4_1),.clk(gclk));
	jdff dff_B_woAQXQKr3_1(.din(G52),.dout(w_dff_B_woAQXQKr3_1),.clk(gclk));
	jdff dff_B_g8h89HDW9_1(.din(w_dff_B_woAQXQKr3_1),.dout(w_dff_B_g8h89HDW9_1),.clk(gclk));
	jdff dff_B_cRPOVfjX1_0(.din(n432),.dout(w_dff_B_cRPOVfjX1_0),.clk(gclk));
	jdff dff_A_kiedNMSw1_0(.dout(w_n809_0[0]),.din(w_dff_A_kiedNMSw1_0),.clk(gclk));
	jdff dff_A_hn1tQkK67_0(.dout(w_n999_4[0]),.din(w_dff_A_hn1tQkK67_0),.clk(gclk));
	jdff dff_A_WGusxvTa4_0(.dout(w_dff_A_hn1tQkK67_0),.din(w_dff_A_WGusxvTa4_0),.clk(gclk));
	jdff dff_A_3nXvSp6U4_0(.dout(w_dff_A_WGusxvTa4_0),.din(w_dff_A_3nXvSp6U4_0),.clk(gclk));
	jdff dff_A_696SBWZe9_0(.dout(w_dff_A_3nXvSp6U4_0),.din(w_dff_A_696SBWZe9_0),.clk(gclk));
	jdff dff_A_PyIf5qVQ1_0(.dout(w_dff_A_696SBWZe9_0),.din(w_dff_A_PyIf5qVQ1_0),.clk(gclk));
	jdff dff_B_Jp14vPOY8_0(.din(n867),.dout(w_dff_B_Jp14vPOY8_0),.clk(gclk));
	jdff dff_B_Grvczgnb2_0(.din(w_dff_B_Jp14vPOY8_0),.dout(w_dff_B_Grvczgnb2_0),.clk(gclk));
	jdff dff_B_9QgfQnwM9_0(.din(w_dff_B_Grvczgnb2_0),.dout(w_dff_B_9QgfQnwM9_0),.clk(gclk));
	jdff dff_B_E90BmrV45_0(.din(w_dff_B_9QgfQnwM9_0),.dout(w_dff_B_E90BmrV45_0),.clk(gclk));
	jdff dff_B_LHxyY0hH1_0(.din(w_dff_B_E90BmrV45_0),.dout(w_dff_B_LHxyY0hH1_0),.clk(gclk));
	jdff dff_B_HpKf3Jb22_0(.din(w_dff_B_LHxyY0hH1_0),.dout(w_dff_B_HpKf3Jb22_0),.clk(gclk));
	jdff dff_B_HM2nPqvS0_1(.din(n864),.dout(w_dff_B_HM2nPqvS0_1),.clk(gclk));
	jdff dff_B_4XQltSQF7_1(.din(G122),.dout(w_dff_B_4XQltSQF7_1),.clk(gclk));
	jdff dff_B_X0msDUlY1_1(.din(w_dff_B_4XQltSQF7_1),.dout(w_dff_B_X0msDUlY1_1),.clk(gclk));
	jdff dff_B_bxr6B7Pd8_0(.din(n468),.dout(w_dff_B_bxr6B7Pd8_0),.clk(gclk));
	jdff dff_A_kqaLlRCo8_0(.dout(w_n862_0[0]),.din(w_dff_A_kqaLlRCo8_0),.clk(gclk));
	jdff dff_B_QRZS0TQ75_1(.din(n852),.dout(w_dff_B_QRZS0TQ75_1),.clk(gclk));
	jdff dff_B_nxN2Esor1_1(.din(w_dff_B_QRZS0TQ75_1),.dout(w_dff_B_nxN2Esor1_1),.clk(gclk));
	jdff dff_B_wtqKpTH95_1(.din(w_dff_B_nxN2Esor1_1),.dout(w_dff_B_wtqKpTH95_1),.clk(gclk));
	jdff dff_B_4Us65xLQ6_1(.din(w_dff_B_wtqKpTH95_1),.dout(w_dff_B_4Us65xLQ6_1),.clk(gclk));
	jdff dff_B_SeCdQpjF7_0(.din(n1121),.dout(w_dff_B_SeCdQpjF7_0),.clk(gclk));
	jdff dff_B_GsZTZZTF3_0(.din(w_dff_B_SeCdQpjF7_0),.dout(w_dff_B_GsZTZZTF3_0),.clk(gclk));
	jdff dff_B_DoSOZjuk2_0(.din(w_dff_B_GsZTZZTF3_0),.dout(w_dff_B_DoSOZjuk2_0),.clk(gclk));
	jdff dff_B_oGIWPZO36_0(.din(w_dff_B_DoSOZjuk2_0),.dout(w_dff_B_oGIWPZO36_0),.clk(gclk));
	jdff dff_B_GVcn3f3y3_0(.din(w_dff_B_oGIWPZO36_0),.dout(w_dff_B_GVcn3f3y3_0),.clk(gclk));
	jdff dff_B_blczhI4C9_0(.din(n1120),.dout(w_dff_B_blczhI4C9_0),.clk(gclk));
	jdff dff_B_BtGuEXDp7_0(.din(w_dff_B_blczhI4C9_0),.dout(w_dff_B_BtGuEXDp7_0),.clk(gclk));
	jdff dff_B_nPwJ4cy59_0(.din(w_dff_B_BtGuEXDp7_0),.dout(w_dff_B_nPwJ4cy59_0),.clk(gclk));
	jdff dff_B_Cv6Jnwn13_0(.din(w_dff_B_nPwJ4cy59_0),.dout(w_dff_B_Cv6Jnwn13_0),.clk(gclk));
	jdff dff_B_ICQv7vJ08_0(.din(w_dff_B_Cv6Jnwn13_0),.dout(w_dff_B_ICQv7vJ08_0),.clk(gclk));
	jdff dff_B_HXNCn4GD1_0(.din(n1119),.dout(w_dff_B_HXNCn4GD1_0),.clk(gclk));
	jdff dff_B_iHtaYKnk5_2(.din(G158),.dout(w_dff_B_iHtaYKnk5_2),.clk(gclk));
	jdff dff_B_IIOCkE468_2(.din(G188),.dout(w_dff_B_IIOCkE468_2),.clk(gclk));
	jdff dff_B_NXJzxM3B9_2(.din(w_dff_B_IIOCkE468_2),.dout(w_dff_B_NXJzxM3B9_2),.clk(gclk));
	jdff dff_B_2i2NURNA2_1(.din(n766),.dout(w_dff_B_2i2NURNA2_1),.clk(gclk));
	jdff dff_B_R4LcYWub1_1(.din(G129),.dout(w_dff_B_R4LcYWub1_1),.clk(gclk));
	jdff dff_B_NZQc0blX1_1(.din(w_dff_B_R4LcYWub1_1),.dout(w_dff_B_NZQc0blX1_1),.clk(gclk));
	jdff dff_A_nclew3Bq1_1(.dout(w_n397_0[1]),.din(w_dff_A_nclew3Bq1_1),.clk(gclk));
	jdff dff_A_dMEordML7_1(.dout(w_dff_A_nclew3Bq1_1),.din(w_dff_A_dMEordML7_1),.clk(gclk));
	jdff dff_B_F0IHH1581_0(.din(n395),.dout(w_dff_B_F0IHH1581_0),.clk(gclk));
	jdff dff_B_ndd83xYU6_0(.din(n763),.dout(w_dff_B_ndd83xYU6_0),.clk(gclk));
	jdff dff_A_Q1pMjrZr8_0(.dout(w_n748_4[0]),.din(w_dff_A_Q1pMjrZr8_0),.clk(gclk));
	jdff dff_B_hkjOxdZj3_0(.din(n898),.dout(w_dff_B_hkjOxdZj3_0),.clk(gclk));
	jdff dff_B_5M6LyKYf2_0(.din(w_dff_B_hkjOxdZj3_0),.dout(w_dff_B_5M6LyKYf2_0),.clk(gclk));
	jdff dff_B_06dd8j4n1_0(.din(w_dff_B_5M6LyKYf2_0),.dout(w_dff_B_06dd8j4n1_0),.clk(gclk));
	jdff dff_B_eM3WcKdS2_0(.din(w_dff_B_06dd8j4n1_0),.dout(w_dff_B_eM3WcKdS2_0),.clk(gclk));
	jdff dff_B_OfAy3uSm0_0(.din(w_dff_B_eM3WcKdS2_0),.dout(w_dff_B_OfAy3uSm0_0),.clk(gclk));
	jdff dff_B_eT3Orvrj8_1(.din(n895),.dout(w_dff_B_eT3Orvrj8_1),.clk(gclk));
	jdff dff_B_2Nbdvzzq5_1(.din(G126),.dout(w_dff_B_2Nbdvzzq5_1),.clk(gclk));
	jdff dff_B_4LuH5Jpo9_1(.din(w_dff_B_2Nbdvzzq5_1),.dout(w_dff_B_4LuH5Jpo9_1),.clk(gclk));
	jdff dff_B_HTcQ0nIP8_0(.din(n492),.dout(w_dff_B_HTcQ0nIP8_0),.clk(gclk));
	jdff dff_B_fSP7FxFs7_0(.din(n889),.dout(w_dff_B_fSP7FxFs7_0),.clk(gclk));
	jdff dff_A_mZmQW8xh3_1(.dout(w_G137_7[1]),.din(w_dff_A_mZmQW8xh3_1),.clk(gclk));
	jdff dff_A_h9YeP2SC0_0(.dout(w_G137_2[0]),.din(w_dff_A_h9YeP2SC0_0),.clk(gclk));
	jdff dff_A_GBysIiG21_0(.dout(w_dff_A_h9YeP2SC0_0),.din(w_dff_A_GBysIiG21_0),.clk(gclk));
	jdff dff_A_2G2UlGTq2_0(.dout(w_dff_A_GBysIiG21_0),.din(w_dff_A_2G2UlGTq2_0),.clk(gclk));
	jdff dff_A_ixpkdBVh1_0(.dout(w_dff_A_2G2UlGTq2_0),.din(w_dff_A_ixpkdBVh1_0),.clk(gclk));
	jdff dff_A_h27SHOlY8_1(.dout(w_G137_2[1]),.din(w_dff_A_h27SHOlY8_1),.clk(gclk));
	jdff dff_A_cSz0DHgh1_1(.dout(w_dff_A_h27SHOlY8_1),.din(w_dff_A_cSz0DHgh1_1),.clk(gclk));
	jdff dff_A_eqRDN5xA8_1(.dout(w_dff_A_cSz0DHgh1_1),.din(w_dff_A_eqRDN5xA8_1),.clk(gclk));
	jdff dff_A_brxb91Nl9_1(.dout(w_dff_A_eqRDN5xA8_1),.din(w_dff_A_brxb91Nl9_1),.clk(gclk));
	jdff dff_B_jXja1grm6_0(.din(n1129),.dout(w_dff_B_jXja1grm6_0),.clk(gclk));
	jdff dff_B_qQQQr57e4_0(.din(w_dff_B_jXja1grm6_0),.dout(w_dff_B_qQQQr57e4_0),.clk(gclk));
	jdff dff_B_ChStDK2h5_0(.din(w_dff_B_qQQQr57e4_0),.dout(w_dff_B_ChStDK2h5_0),.clk(gclk));
	jdff dff_B_i1TJoECv1_0(.din(w_dff_B_ChStDK2h5_0),.dout(w_dff_B_i1TJoECv1_0),.clk(gclk));
	jdff dff_B_9UhDffR76_0(.din(n1128),.dout(w_dff_B_9UhDffR76_0),.clk(gclk));
	jdff dff_B_hyVTKsxV8_0(.din(w_dff_B_9UhDffR76_0),.dout(w_dff_B_hyVTKsxV8_0),.clk(gclk));
	jdff dff_B_43etQwju5_0(.din(w_dff_B_hyVTKsxV8_0),.dout(w_dff_B_43etQwju5_0),.clk(gclk));
	jdff dff_B_dmuBxmgh2_0(.din(w_dff_B_43etQwju5_0),.dout(w_dff_B_dmuBxmgh2_0),.clk(gclk));
	jdff dff_B_n35d1YZH7_0(.din(w_dff_B_dmuBxmgh2_0),.dout(w_dff_B_n35d1YZH7_0),.clk(gclk));
	jdff dff_B_wtTfk3g40_0(.din(w_dff_B_n35d1YZH7_0),.dout(w_dff_B_wtTfk3g40_0),.clk(gclk));
	jdff dff_B_lGjRA1MP6_0(.din(n1127),.dout(w_dff_B_lGjRA1MP6_0),.clk(gclk));
	jdff dff_B_F85S2bmz5_2(.din(G152),.dout(w_dff_B_F85S2bmz5_2),.clk(gclk));
	jdff dff_B_brbJCPoz3_2(.din(G155),.dout(w_dff_B_brbJCPoz3_2),.clk(gclk));
	jdff dff_B_tDQP5nyd7_2(.din(w_dff_B_brbJCPoz3_2),.dout(w_dff_B_tDQP5nyd7_2),.clk(gclk));
	jdff dff_B_B4AvEkKb9_0(.din(n837),.dout(w_dff_B_B4AvEkKb9_0),.clk(gclk));
	jdff dff_B_AIv8lL129_1(.din(n834),.dout(w_dff_B_AIv8lL129_1),.clk(gclk));
	jdff dff_B_9j0d0Nud2_1(.din(G119),.dout(w_dff_B_9j0d0Nud2_1),.clk(gclk));
	jdff dff_B_UnolPSSa7_1(.din(w_dff_B_9j0d0Nud2_1),.dout(w_dff_B_UnolPSSa7_1),.clk(gclk));
	jdff dff_B_JsUpw6qs3_0(.din(n443),.dout(w_dff_B_JsUpw6qs3_0),.clk(gclk));
	jdff dff_A_mrTqWM7Y8_0(.dout(w_n744_1[0]),.din(w_dff_A_mrTqWM7Y8_0),.clk(gclk));
	jdff dff_A_7dbIcJVQ6_0(.dout(w_dff_A_mrTqWM7Y8_0),.din(w_dff_A_7dbIcJVQ6_0),.clk(gclk));
	jdff dff_A_lJ4K7l0o8_0(.dout(w_dff_A_7dbIcJVQ6_0),.din(w_dff_A_lJ4K7l0o8_0),.clk(gclk));
	jdff dff_B_loTIAKmz0_0(.din(n887),.dout(w_dff_B_loTIAKmz0_0),.clk(gclk));
	jdff dff_B_932T30un2_0(.din(w_dff_B_loTIAKmz0_0),.dout(w_dff_B_932T30un2_0),.clk(gclk));
	jdff dff_B_xnOx4Plp4_0(.din(w_dff_B_932T30un2_0),.dout(w_dff_B_xnOx4Plp4_0),.clk(gclk));
	jdff dff_B_ZxEwx3is0_0(.din(w_dff_B_xnOx4Plp4_0),.dout(w_dff_B_ZxEwx3is0_0),.clk(gclk));
	jdff dff_B_cPsXwyo38_0(.din(w_dff_B_ZxEwx3is0_0),.dout(w_dff_B_cPsXwyo38_0),.clk(gclk));
	jdff dff_B_UhDPWxwS4_1(.din(n884),.dout(w_dff_B_UhDPWxwS4_1),.clk(gclk));
	jdff dff_B_h5xBjHl44_1(.din(G127),.dout(w_dff_B_h5xBjHl44_1),.clk(gclk));
	jdff dff_B_oY61uKLk2_1(.din(w_dff_B_h5xBjHl44_1),.dout(w_dff_B_oY61uKLk2_1),.clk(gclk));
	jdff dff_A_eGdNV9IC6_1(.dout(w_n459_0[1]),.din(w_dff_A_eGdNV9IC6_1),.clk(gclk));
	jdff dff_B_ADAxB4i80_0(.din(n457),.dout(w_dff_B_ADAxB4i80_0),.clk(gclk));
	jdff dff_A_MkzCM3QZ5_0(.dout(w_n879_0[0]),.din(w_dff_A_MkzCM3QZ5_0),.clk(gclk));
	jdff dff_B_AemQpIVj9_0(.din(n1137),.dout(w_dff_B_AemQpIVj9_0),.clk(gclk));
	jdff dff_B_xK6VGpEU5_0(.din(w_dff_B_AemQpIVj9_0),.dout(w_dff_B_xK6VGpEU5_0),.clk(gclk));
	jdff dff_B_YWZeFU5n3_0(.din(w_dff_B_xK6VGpEU5_0),.dout(w_dff_B_YWZeFU5n3_0),.clk(gclk));
	jdff dff_B_d6uNA6YY6_0(.din(w_dff_B_YWZeFU5n3_0),.dout(w_dff_B_d6uNA6YY6_0),.clk(gclk));
	jdff dff_B_EXi4GZeS8_0(.din(n1136),.dout(w_dff_B_EXi4GZeS8_0),.clk(gclk));
	jdff dff_B_vD5Fk35Y5_0(.din(w_dff_B_EXi4GZeS8_0),.dout(w_dff_B_vD5Fk35Y5_0),.clk(gclk));
	jdff dff_B_t9tYVirr1_0(.din(w_dff_B_vD5Fk35Y5_0),.dout(w_dff_B_t9tYVirr1_0),.clk(gclk));
	jdff dff_B_VziqwfyY0_0(.din(w_dff_B_t9tYVirr1_0),.dout(w_dff_B_VziqwfyY0_0),.clk(gclk));
	jdff dff_B_uMuZL7Bd4_0(.din(w_dff_B_VziqwfyY0_0),.dout(w_dff_B_uMuZL7Bd4_0),.clk(gclk));
	jdff dff_B_Uf2LOJKb1_0(.din(w_dff_B_uMuZL7Bd4_0),.dout(w_dff_B_Uf2LOJKb1_0),.clk(gclk));
	jdff dff_B_AdB8vm2y9_0(.din(n1135),.dout(w_dff_B_AdB8vm2y9_0),.clk(gclk));
	jdff dff_B_uA3DEimy4_2(.din(G146),.dout(w_dff_B_uA3DEimy4_2),.clk(gclk));
	jdff dff_B_HDXzGdZK7_2(.din(G149),.dout(w_dff_B_HDXzGdZK7_2),.clk(gclk));
	jdff dff_B_EHofCk4u4_2(.din(w_dff_B_HDXzGdZK7_2),.dout(w_dff_B_EHofCk4u4_2),.clk(gclk));
	jdff dff_A_dpCZoQk20_0(.dout(w_n1002_3[0]),.din(w_dff_A_dpCZoQk20_0),.clk(gclk));
	jdff dff_A_7luvimY03_1(.dout(w_n1002_3[1]),.din(w_dff_A_7luvimY03_1),.clk(gclk));
	jdff dff_B_mE0h48r77_0(.din(n826),.dout(w_dff_B_mE0h48r77_0),.clk(gclk));
	jdff dff_B_IGABrCwK7_0(.din(w_dff_B_mE0h48r77_0),.dout(w_dff_B_IGABrCwK7_0),.clk(gclk));
	jdff dff_B_pNgu8r555_1(.din(G130),.dout(w_dff_B_pNgu8r555_1),.clk(gclk));
	jdff dff_B_H8s9gCkA2_1(.din(w_dff_B_pNgu8r555_1),.dout(w_dff_B_H8s9gCkA2_1),.clk(gclk));
	jdff dff_B_1BQvMScw8_0(.din(n413),.dout(w_dff_B_1BQvMScw8_0),.clk(gclk));
	jdff dff_A_tduSDlpK3_0(.dout(w_n821_0[0]),.din(w_dff_A_tduSDlpK3_0),.clk(gclk));
	jdff dff_B_4emycJed9_1(.din(n816),.dout(w_dff_B_4emycJed9_1),.clk(gclk));
	jdff dff_A_iBioveLm8_2(.dout(w_n744_0[2]),.din(w_dff_A_iBioveLm8_2),.clk(gclk));
	jdff dff_A_UOES35z51_2(.dout(w_dff_A_iBioveLm8_2),.din(w_dff_A_UOES35z51_2),.clk(gclk));
	jdff dff_B_luKw20Og5_3(.din(n744),.dout(w_dff_B_luKw20Og5_3),.clk(gclk));
	jdff dff_A_scjTpqwT0_2(.dout(w_n748_3[2]),.din(w_dff_A_scjTpqwT0_2),.clk(gclk));
	jdff dff_B_m6qwZRr16_0(.din(n874),.dout(w_dff_B_m6qwZRr16_0),.clk(gclk));
	jdff dff_B_3R4wQPxn7_0(.din(w_dff_B_m6qwZRr16_0),.dout(w_dff_B_3R4wQPxn7_0),.clk(gclk));
	jdff dff_B_c5I1m2YB9_0(.din(w_dff_B_3R4wQPxn7_0),.dout(w_dff_B_c5I1m2YB9_0),.clk(gclk));
	jdff dff_B_Lo8OStMm4_0(.din(w_dff_B_c5I1m2YB9_0),.dout(w_dff_B_Lo8OStMm4_0),.clk(gclk));
	jdff dff_B_I14rXkob3_0(.din(w_dff_B_Lo8OStMm4_0),.dout(w_dff_B_I14rXkob3_0),.clk(gclk));
	jdff dff_B_VWz7lHXZ8_1(.din(n871),.dout(w_dff_B_VWz7lHXZ8_1),.clk(gclk));
	jdff dff_B_O9QHLiIa6_1(.din(G128),.dout(w_dff_B_O9QHLiIa6_1),.clk(gclk));
	jdff dff_B_HRMR7rpT2_1(.din(w_dff_B_O9QHLiIa6_1),.dout(w_dff_B_HRMR7rpT2_1),.clk(gclk));
	jdff dff_B_99e8Gtle2_0(.din(n479),.dout(w_dff_B_99e8Gtle2_0),.clk(gclk));
	jdff dff_A_cp2V9q6e7_0(.dout(w_n869_0[0]),.din(w_dff_A_cp2V9q6e7_0),.clk(gclk));
	jdff dff_B_epkIxhZs3_0(.din(n858),.dout(w_dff_B_epkIxhZs3_0),.clk(gclk));
	jdff dff_B_3B64H4dF4_0(.din(w_dff_B_epkIxhZs3_0),.dout(w_dff_B_3B64H4dF4_0),.clk(gclk));
	jdff dff_B_sGff82Uf3_0(.din(w_dff_B_3B64H4dF4_0),.dout(w_dff_B_sGff82Uf3_0),.clk(gclk));
	jdff dff_A_CocBSnos7_0(.dout(w_G4_1[0]),.din(w_dff_A_CocBSnos7_0),.clk(gclk));
	jdff dff_A_xUYhHAIk5_0(.dout(w_dff_A_CocBSnos7_0),.din(w_dff_A_xUYhHAIk5_0),.clk(gclk));
	jdff dff_B_SSfT7VwG3_0(.din(n1155),.dout(w_dff_B_SSfT7VwG3_0),.clk(gclk));
	jdff dff_B_t67Rp19n4_0(.din(w_dff_B_SSfT7VwG3_0),.dout(w_dff_B_t67Rp19n4_0),.clk(gclk));
	jdff dff_B_Z8j8lMpG2_0(.din(w_dff_B_t67Rp19n4_0),.dout(w_dff_B_Z8j8lMpG2_0),.clk(gclk));
	jdff dff_B_DcnYlsUl8_0(.din(w_dff_B_Z8j8lMpG2_0),.dout(w_dff_B_DcnYlsUl8_0),.clk(gclk));
	jdff dff_B_WPf4cHkf0_0(.din(w_dff_B_DcnYlsUl8_0),.dout(w_dff_B_WPf4cHkf0_0),.clk(gclk));
	jdff dff_B_WNZNiIJS5_0(.din(w_dff_B_WPf4cHkf0_0),.dout(w_dff_B_WNZNiIJS5_0),.clk(gclk));
	jdff dff_B_9alznzrA7_1(.din(n1148),.dout(w_dff_B_9alznzrA7_1),.clk(gclk));
	jdff dff_B_iXCOEUcA2_1(.din(w_dff_B_9alznzrA7_1),.dout(w_dff_B_iXCOEUcA2_1),.clk(gclk));
	jdff dff_B_8iUufvxb4_1(.din(w_dff_B_iXCOEUcA2_1),.dout(w_dff_B_8iUufvxb4_1),.clk(gclk));
	jdff dff_B_9Rj5hHeL6_0(.din(n1144),.dout(w_dff_B_9Rj5hHeL6_0),.clk(gclk));
	jdff dff_B_BDmvZIaY5_0(.din(w_dff_B_9Rj5hHeL6_0),.dout(w_dff_B_BDmvZIaY5_0),.clk(gclk));
	jdff dff_B_evefBOMY8_0(.din(w_dff_B_BDmvZIaY5_0),.dout(w_dff_B_evefBOMY8_0),.clk(gclk));
	jdff dff_B_cezlCk7Y4_0(.din(w_dff_B_evefBOMY8_0),.dout(w_dff_B_cezlCk7Y4_0),.clk(gclk));
	jdff dff_B_MIcPi9al6_0(.din(w_dff_B_cezlCk7Y4_0),.dout(w_dff_B_MIcPi9al6_0),.clk(gclk));
	jdff dff_B_tnAQ7MbG3_0(.din(w_dff_B_MIcPi9al6_0),.dout(w_dff_B_tnAQ7MbG3_0),.clk(gclk));
	jdff dff_B_zqUFj38Q5_0(.din(w_dff_B_tnAQ7MbG3_0),.dout(w_dff_B_zqUFj38Q5_0),.clk(gclk));
	jdff dff_B_QikZCtSI9_0(.din(w_dff_B_zqUFj38Q5_0),.dout(w_dff_B_QikZCtSI9_0),.clk(gclk));
	jdff dff_B_ROAuJexP8_0(.din(w_dff_B_QikZCtSI9_0),.dout(w_dff_B_ROAuJexP8_0),.clk(gclk));
	jdff dff_B_skaBgWq53_1(.din(n1141),.dout(w_dff_B_skaBgWq53_1),.clk(gclk));
	jdff dff_A_gaSKnasO8_0(.dout(w_n1142_0[0]),.din(w_dff_A_gaSKnasO8_0),.clk(gclk));
	jdff dff_A_EI7ad8R13_0(.dout(w_dff_A_gaSKnasO8_0),.din(w_dff_A_EI7ad8R13_0),.clk(gclk));
	jdff dff_A_WrcUgB0F1_0(.dout(w_G3717_0[0]),.din(w_dff_A_WrcUgB0F1_0),.clk(gclk));
	jdff dff_A_67RcbT2e6_0(.dout(w_dff_A_WrcUgB0F1_0),.din(w_dff_A_67RcbT2e6_0),.clk(gclk));
	jdff dff_A_c1SIEnVh5_0(.dout(w_dff_A_67RcbT2e6_0),.din(w_dff_A_c1SIEnVh5_0),.clk(gclk));
	jdff dff_A_FvB3tIyx2_0(.dout(w_dff_A_c1SIEnVh5_0),.din(w_dff_A_FvB3tIyx2_0),.clk(gclk));
	jdff dff_A_ySM5rlIz0_0(.dout(w_G3724_0[0]),.din(w_dff_A_ySM5rlIz0_0),.clk(gclk));
	jdff dff_A_GycpXLU83_0(.dout(w_dff_A_ySM5rlIz0_0),.din(w_dff_A_GycpXLU83_0),.clk(gclk));
	jdff dff_A_629NqC8a0_0(.dout(w_dff_A_GycpXLU83_0),.din(w_dff_A_629NqC8a0_0),.clk(gclk));
	jdff dff_A_YnPLfKPy1_2(.dout(w_G3724_0[2]),.din(w_dff_A_YnPLfKPy1_2),.clk(gclk));
	jdff dff_A_DGr94NIX6_2(.dout(w_dff_A_YnPLfKPy1_2),.din(w_dff_A_DGr94NIX6_2),.clk(gclk));
	jdff dff_A_55gpo2Ti6_2(.dout(w_dff_A_DGr94NIX6_2),.din(w_dff_A_55gpo2Ti6_2),.clk(gclk));
	jdff dff_A_Rz7TMaaL4_2(.dout(w_dff_A_55gpo2Ti6_2),.din(w_dff_A_Rz7TMaaL4_2),.clk(gclk));
	jdff dff_A_h6fIR9He3_2(.dout(w_dff_A_Rz7TMaaL4_2),.din(w_dff_A_h6fIR9He3_2),.clk(gclk));
	jdff dff_A_hqjnQ6OE8_2(.dout(w_dff_A_h6fIR9He3_2),.din(w_dff_A_hqjnQ6OE8_2),.clk(gclk));
	jdff dff_A_Ju0cGdxc2_2(.dout(w_dff_A_hqjnQ6OE8_2),.din(w_dff_A_Ju0cGdxc2_2),.clk(gclk));
	jdff dff_A_0meZ6t1G5_2(.dout(w_dff_A_Ju0cGdxc2_2),.din(w_dff_A_0meZ6t1G5_2),.clk(gclk));
	jdff dff_A_jO3GpOIl5_2(.dout(w_dff_A_0meZ6t1G5_2),.din(w_dff_A_jO3GpOIl5_2),.clk(gclk));
	jdff dff_A_YCUoHJmc3_2(.dout(w_dff_A_jO3GpOIl5_2),.din(w_dff_A_YCUoHJmc3_2),.clk(gclk));
	jdff dff_A_qfKdnG4t3_0(.dout(w_G132_0[0]),.din(w_dff_A_qfKdnG4t3_0),.clk(gclk));
	jdff dff_A_A3E73v3x3_0(.dout(w_dff_A_qfKdnG4t3_0),.din(w_dff_A_A3E73v3x3_0),.clk(gclk));
	jdff dff_A_zQxJxC6H6_0(.dout(w_dff_A_A3E73v3x3_0),.din(w_dff_A_zQxJxC6H6_0),.clk(gclk));
	jdff dff_A_arJIqD5j3_0(.dout(w_dff_A_zQxJxC6H6_0),.din(w_dff_A_arJIqD5j3_0),.clk(gclk));
	jdff dff_A_m80uWGCS8_0(.dout(w_dff_A_arJIqD5j3_0),.din(w_dff_A_m80uWGCS8_0),.clk(gclk));
	jdff dff_A_F3dasG4b4_0(.dout(w_dff_A_m80uWGCS8_0),.din(w_dff_A_F3dasG4b4_0),.clk(gclk));
	jdff dff_B_88yunF5y9_2(.din(G132),.dout(w_dff_B_88yunF5y9_2),.clk(gclk));
	jdff dff_B_UOzhcatG6_2(.din(w_dff_B_88yunF5y9_2),.dout(w_dff_B_UOzhcatG6_2),.clk(gclk));
	jdff dff_B_OsXxBvxJ0_1(.din(n1184),.dout(w_dff_B_OsXxBvxJ0_1),.clk(gclk));
	jdff dff_B_cIa0RRGx9_0(.din(n1189),.dout(w_dff_B_cIa0RRGx9_0),.clk(gclk));
	jdff dff_B_myBjpaiO4_0(.din(w_dff_B_cIa0RRGx9_0),.dout(w_dff_B_myBjpaiO4_0),.clk(gclk));
	jdff dff_B_ryzSXgLC1_0(.din(n1187),.dout(w_dff_B_ryzSXgLC1_0),.clk(gclk));
	jdff dff_A_OpW0ntUi9_0(.dout(w_G601_0),.din(w_dff_A_OpW0ntUi9_0),.clk(gclk));
	jdff dff_B_1wrzx3hs6_1(.din(n656),.dout(w_dff_B_1wrzx3hs6_1),.clk(gclk));
	jdff dff_A_GfxdPqk05_0(.dout(w_n671_0[0]),.din(w_dff_A_GfxdPqk05_0),.clk(gclk));
	jdff dff_B_PK1nw0l90_1(.din(n665),.dout(w_dff_B_PK1nw0l90_1),.clk(gclk));
	jdff dff_B_Qqtg0nxm7_0(.din(n913),.dout(w_dff_B_Qqtg0nxm7_0),.clk(gclk));
	jdff dff_B_KLnd0Szl5_1(.din(n907),.dout(w_dff_B_KLnd0Szl5_1),.clk(gclk));
	jdff dff_B_ImVXIuGq5_1(.din(n909),.dout(w_dff_B_ImVXIuGq5_1),.clk(gclk));
	jdff dff_B_XFaalHQD9_1(.din(w_dff_B_ImVXIuGq5_1),.dout(w_dff_B_XFaalHQD9_1),.clk(gclk));
	jdff dff_B_9t3Iv5XK3_0(.din(n910),.dout(w_dff_B_9t3Iv5XK3_0),.clk(gclk));
	jdff dff_B_mqvQ6SXx6_1(.din(n908),.dout(w_dff_B_mqvQ6SXx6_1),.clk(gclk));
	jdff dff_B_F4wIN6jS5_0(.din(n904),.dout(w_dff_B_F4wIN6jS5_0),.clk(gclk));
	jdff dff_A_6gJRWWHu3_0(.dout(w_G369_0[0]),.din(w_dff_A_6gJRWWHu3_0),.clk(gclk));
	jdff dff_B_VurSCaJD9_0(.din(n900),.dout(w_dff_B_VurSCaJD9_0),.clk(gclk));
	jdff dff_A_5cIVWmKE3_0(.dout(w_n621_1[0]),.din(w_dff_A_5cIVWmKE3_0),.clk(gclk));
	jdff dff_A_8SlZqIuw7_0(.dout(w_dff_A_5cIVWmKE3_0),.din(w_dff_A_8SlZqIuw7_0),.clk(gclk));
	jdff dff_A_oLBtXOd74_0(.dout(w_dff_A_8SlZqIuw7_0),.din(w_dff_A_oLBtXOd74_0),.clk(gclk));
	jdff dff_A_ZzUXv6Dg6_0(.dout(w_dff_A_oLBtXOd74_0),.din(w_dff_A_ZzUXv6Dg6_0),.clk(gclk));
	jdff dff_B_mfm0ebpX6_1(.din(n919),.dout(w_dff_B_mfm0ebpX6_1),.clk(gclk));
	jdff dff_B_lpWqvyMa2_0(.din(n923),.dout(w_dff_B_lpWqvyMa2_0),.clk(gclk));
	jdff dff_B_c1NEaN4f0_0(.din(n921),.dout(w_dff_B_c1NEaN4f0_0),.clk(gclk));
	jdff dff_A_wLOdru9x4_0(.dout(w_G289_0[0]),.din(w_dff_A_wLOdru9x4_0),.clk(gclk));
	jdff dff_B_0HVgotjO2_0(.din(n1225),.dout(w_dff_B_0HVgotjO2_0),.clk(gclk));
	jdff dff_B_nAmKSWzQ8_0(.din(w_dff_B_0HVgotjO2_0),.dout(w_dff_B_nAmKSWzQ8_0),.clk(gclk));
	jdff dff_B_pwZfNd2I0_0(.din(n1224),.dout(w_dff_B_pwZfNd2I0_0),.clk(gclk));
	jdff dff_B_T5Qe86438_0(.din(w_dff_B_pwZfNd2I0_0),.dout(w_dff_B_T5Qe86438_0),.clk(gclk));
	jdff dff_B_SyZgZmfS3_0(.din(w_dff_B_T5Qe86438_0),.dout(w_dff_B_SyZgZmfS3_0),.clk(gclk));
	jdff dff_B_sJ1EqXTQ3_0(.din(w_dff_B_SyZgZmfS3_0),.dout(w_dff_B_sJ1EqXTQ3_0),.clk(gclk));
	jdff dff_B_F0CJDHJM1_0(.din(w_dff_B_sJ1EqXTQ3_0),.dout(w_dff_B_F0CJDHJM1_0),.clk(gclk));
	jdff dff_B_n1ggcqH11_0(.din(w_dff_B_F0CJDHJM1_0),.dout(w_dff_B_n1ggcqH11_0),.clk(gclk));
	jdff dff_B_95K4cv8e4_0(.din(w_dff_B_n1ggcqH11_0),.dout(w_dff_B_95K4cv8e4_0),.clk(gclk));
	jdff dff_B_S8poXftF0_0(.din(w_dff_B_95K4cv8e4_0),.dout(w_dff_B_S8poXftF0_0),.clk(gclk));
	jdff dff_B_lcRHJFF64_0(.din(w_dff_B_S8poXftF0_0),.dout(w_dff_B_lcRHJFF64_0),.clk(gclk));
	jdff dff_B_e8e7yQGH2_0(.din(n1223),.dout(w_dff_B_e8e7yQGH2_0),.clk(gclk));
	jdff dff_B_XuaI41C61_0(.din(n1232),.dout(w_dff_B_XuaI41C61_0),.clk(gclk));
	jdff dff_B_YVGo4UPM2_0(.din(w_dff_B_XuaI41C61_0),.dout(w_dff_B_YVGo4UPM2_0),.clk(gclk));
	jdff dff_B_Fb5Ls2ud3_0(.din(n1231),.dout(w_dff_B_Fb5Ls2ud3_0),.clk(gclk));
	jdff dff_B_20IF8xx75_0(.din(w_dff_B_Fb5Ls2ud3_0),.dout(w_dff_B_20IF8xx75_0),.clk(gclk));
	jdff dff_B_aUdnxN211_0(.din(w_dff_B_20IF8xx75_0),.dout(w_dff_B_aUdnxN211_0),.clk(gclk));
	jdff dff_B_baLZapjS5_0(.din(w_dff_B_aUdnxN211_0),.dout(w_dff_B_baLZapjS5_0),.clk(gclk));
	jdff dff_B_ubwNbGnP8_0(.din(w_dff_B_baLZapjS5_0),.dout(w_dff_B_ubwNbGnP8_0),.clk(gclk));
	jdff dff_B_K8fPladJ7_0(.din(w_dff_B_ubwNbGnP8_0),.dout(w_dff_B_K8fPladJ7_0),.clk(gclk));
	jdff dff_B_ydNagheH1_0(.din(w_dff_B_K8fPladJ7_0),.dout(w_dff_B_ydNagheH1_0),.clk(gclk));
	jdff dff_B_B8ShOeCI8_0(.din(w_dff_B_ydNagheH1_0),.dout(w_dff_B_B8ShOeCI8_0),.clk(gclk));
	jdff dff_B_lBEKmMGR7_0(.din(w_dff_B_B8ShOeCI8_0),.dout(w_dff_B_lBEKmMGR7_0),.clk(gclk));
	jdff dff_B_D1GTF7xj2_0(.din(n1230),.dout(w_dff_B_D1GTF7xj2_0),.clk(gclk));
	jdff dff_B_9zaiP92j1_2(.din(G106),.dout(w_dff_B_9zaiP92j1_2),.clk(gclk));
	jdff dff_B_UnAOanOz8_2(.din(G109),.dout(w_dff_B_UnAOanOz8_2),.clk(gclk));
	jdff dff_B_THH2YkVh9_2(.din(w_dff_B_UnAOanOz8_2),.dout(w_dff_B_THH2YkVh9_2),.clk(gclk));
	jdff dff_B_gsB4FoXm1_0(.din(n1240),.dout(w_dff_B_gsB4FoXm1_0),.clk(gclk));
	jdff dff_B_4kLkfKo12_0(.din(w_dff_B_gsB4FoXm1_0),.dout(w_dff_B_4kLkfKo12_0),.clk(gclk));
	jdff dff_B_21ZpFLLb4_0(.din(n1239),.dout(w_dff_B_21ZpFLLb4_0),.clk(gclk));
	jdff dff_B_CMEIqyEC2_0(.din(w_dff_B_21ZpFLLb4_0),.dout(w_dff_B_CMEIqyEC2_0),.clk(gclk));
	jdff dff_B_IZhbXuXO6_0(.din(w_dff_B_CMEIqyEC2_0),.dout(w_dff_B_IZhbXuXO6_0),.clk(gclk));
	jdff dff_B_CHzR3QmG2_0(.din(w_dff_B_IZhbXuXO6_0),.dout(w_dff_B_CHzR3QmG2_0),.clk(gclk));
	jdff dff_B_PtJene9p6_0(.din(w_dff_B_CHzR3QmG2_0),.dout(w_dff_B_PtJene9p6_0),.clk(gclk));
	jdff dff_B_7UMCqO7y1_0(.din(w_dff_B_PtJene9p6_0),.dout(w_dff_B_7UMCqO7y1_0),.clk(gclk));
	jdff dff_B_3ZkuFiEy8_0(.din(w_dff_B_7UMCqO7y1_0),.dout(w_dff_B_3ZkuFiEy8_0),.clk(gclk));
	jdff dff_B_bNuuCorj1_0(.din(w_dff_B_3ZkuFiEy8_0),.dout(w_dff_B_bNuuCorj1_0),.clk(gclk));
	jdff dff_B_9lyVfhjn2_0(.din(w_dff_B_bNuuCorj1_0),.dout(w_dff_B_9lyVfhjn2_0),.clk(gclk));
	jdff dff_B_jdyTFGON9_0(.din(n1238),.dout(w_dff_B_jdyTFGON9_0),.clk(gclk));
	jdff dff_B_f93g6uv19_0(.din(n1249),.dout(w_dff_B_f93g6uv19_0),.clk(gclk));
	jdff dff_B_K6eGth8v6_0(.din(w_dff_B_f93g6uv19_0),.dout(w_dff_B_K6eGth8v6_0),.clk(gclk));
	jdff dff_B_KEvTavOV0_0(.din(w_dff_B_K6eGth8v6_0),.dout(w_dff_B_KEvTavOV0_0),.clk(gclk));
	jdff dff_B_6ZmFjkKK2_0(.din(n1248),.dout(w_dff_B_6ZmFjkKK2_0),.clk(gclk));
	jdff dff_B_XSqPl3ZV0_0(.din(w_dff_B_6ZmFjkKK2_0),.dout(w_dff_B_XSqPl3ZV0_0),.clk(gclk));
	jdff dff_B_zBWmmBda7_0(.din(w_dff_B_XSqPl3ZV0_0),.dout(w_dff_B_zBWmmBda7_0),.clk(gclk));
	jdff dff_B_RUW842451_0(.din(w_dff_B_zBWmmBda7_0),.dout(w_dff_B_RUW842451_0),.clk(gclk));
	jdff dff_B_8pYaD5ov0_0(.din(w_dff_B_RUW842451_0),.dout(w_dff_B_8pYaD5ov0_0),.clk(gclk));
	jdff dff_B_QArQyq8Q0_0(.din(w_dff_B_8pYaD5ov0_0),.dout(w_dff_B_QArQyq8Q0_0),.clk(gclk));
	jdff dff_B_EXBGyFM30_0(.din(w_dff_B_QArQyq8Q0_0),.dout(w_dff_B_EXBGyFM30_0),.clk(gclk));
	jdff dff_B_xfouMmUx8_0(.din(w_dff_B_EXBGyFM30_0),.dout(w_dff_B_xfouMmUx8_0),.clk(gclk));
	jdff dff_B_YBXa6sB24_0(.din(w_dff_B_xfouMmUx8_0),.dout(w_dff_B_YBXa6sB24_0),.clk(gclk));
	jdff dff_B_8J0lArrZ8_0(.din(n1247),.dout(w_dff_B_8J0lArrZ8_0),.clk(gclk));
	jdff dff_A_2X5lSC9C7_0(.dout(w_n793_2[0]),.din(w_dff_A_2X5lSC9C7_0),.clk(gclk));
	jdff dff_B_wrLMei2Q8_0(.din(n1258),.dout(w_dff_B_wrLMei2Q8_0),.clk(gclk));
	jdff dff_B_YxTIEnT70_0(.din(w_dff_B_wrLMei2Q8_0),.dout(w_dff_B_YxTIEnT70_0),.clk(gclk));
	jdff dff_B_XS8AGY9p0_0(.din(w_dff_B_YxTIEnT70_0),.dout(w_dff_B_XS8AGY9p0_0),.clk(gclk));
	jdff dff_B_YT8gJEJV1_0(.din(n1257),.dout(w_dff_B_YT8gJEJV1_0),.clk(gclk));
	jdff dff_B_hn1epTdc7_0(.din(w_dff_B_YT8gJEJV1_0),.dout(w_dff_B_hn1epTdc7_0),.clk(gclk));
	jdff dff_B_WCGhpb738_0(.din(w_dff_B_hn1epTdc7_0),.dout(w_dff_B_WCGhpb738_0),.clk(gclk));
	jdff dff_B_Sr29IMGI0_0(.din(w_dff_B_WCGhpb738_0),.dout(w_dff_B_Sr29IMGI0_0),.clk(gclk));
	jdff dff_B_OAWvXCb19_0(.din(w_dff_B_Sr29IMGI0_0),.dout(w_dff_B_OAWvXCb19_0),.clk(gclk));
	jdff dff_B_W7QiUbOv5_0(.din(w_dff_B_OAWvXCb19_0),.dout(w_dff_B_W7QiUbOv5_0),.clk(gclk));
	jdff dff_B_c5Wf58tx4_0(.din(w_dff_B_W7QiUbOv5_0),.dout(w_dff_B_c5Wf58tx4_0),.clk(gclk));
	jdff dff_B_8H9Nxs8R9_0(.din(w_dff_B_c5Wf58tx4_0),.dout(w_dff_B_8H9Nxs8R9_0),.clk(gclk));
	jdff dff_B_zrm5P10X0_0(.din(w_dff_B_8H9Nxs8R9_0),.dout(w_dff_B_zrm5P10X0_0),.clk(gclk));
	jdff dff_B_6M8cMGMJ4_0(.din(w_dff_B_zrm5P10X0_0),.dout(w_dff_B_6M8cMGMJ4_0),.clk(gclk));
	jdff dff_B_By08MlUX8_0(.din(n1256),.dout(w_dff_B_By08MlUX8_0),.clk(gclk));
	jdff dff_B_bfR9spID6_0(.din(n1265),.dout(w_dff_B_bfR9spID6_0),.clk(gclk));
	jdff dff_B_5NMMGf1M8_0(.din(w_dff_B_bfR9spID6_0),.dout(w_dff_B_5NMMGf1M8_0),.clk(gclk));
	jdff dff_B_SuUkj5c21_0(.din(n1264),.dout(w_dff_B_SuUkj5c21_0),.clk(gclk));
	jdff dff_B_OENpHhtD4_0(.din(w_dff_B_SuUkj5c21_0),.dout(w_dff_B_OENpHhtD4_0),.clk(gclk));
	jdff dff_B_uXsAf7yt8_0(.din(w_dff_B_OENpHhtD4_0),.dout(w_dff_B_uXsAf7yt8_0),.clk(gclk));
	jdff dff_B_so6IUW984_0(.din(w_dff_B_uXsAf7yt8_0),.dout(w_dff_B_so6IUW984_0),.clk(gclk));
	jdff dff_B_xRaaIIR30_0(.din(w_dff_B_so6IUW984_0),.dout(w_dff_B_xRaaIIR30_0),.clk(gclk));
	jdff dff_B_GPFUh6Jo5_0(.din(w_dff_B_xRaaIIR30_0),.dout(w_dff_B_GPFUh6Jo5_0),.clk(gclk));
	jdff dff_B_hDZQT4wf6_0(.din(w_dff_B_GPFUh6Jo5_0),.dout(w_dff_B_hDZQT4wf6_0),.clk(gclk));
	jdff dff_B_5zdEAoKI9_0(.din(w_dff_B_hDZQT4wf6_0),.dout(w_dff_B_5zdEAoKI9_0),.clk(gclk));
	jdff dff_B_eTqwgJac6_0(.din(w_dff_B_5zdEAoKI9_0),.dout(w_dff_B_eTqwgJac6_0),.clk(gclk));
	jdff dff_B_V3RaC9xA7_0(.din(n1263),.dout(w_dff_B_V3RaC9xA7_0),.clk(gclk));
	jdff dff_B_NNNAuk3Y0_2(.din(G49),.dout(w_dff_B_NNNAuk3Y0_2),.clk(gclk));
	jdff dff_B_nGik8l1A5_2(.din(G46),.dout(w_dff_B_nGik8l1A5_2),.clk(gclk));
	jdff dff_B_19FnkAzX5_2(.din(w_dff_B_nGik8l1A5_2),.dout(w_dff_B_19FnkAzX5_2),.clk(gclk));
	jdff dff_B_NNKyvdJ29_0(.din(n1272),.dout(w_dff_B_NNKyvdJ29_0),.clk(gclk));
	jdff dff_B_5Tx3Shrb9_0(.din(w_dff_B_NNKyvdJ29_0),.dout(w_dff_B_5Tx3Shrb9_0),.clk(gclk));
	jdff dff_B_LqaCsD8p8_0(.din(w_dff_B_5Tx3Shrb9_0),.dout(w_dff_B_LqaCsD8p8_0),.clk(gclk));
	jdff dff_B_mO9xCXNt0_0(.din(n1271),.dout(w_dff_B_mO9xCXNt0_0),.clk(gclk));
	jdff dff_B_7lA60dox5_0(.din(w_dff_B_mO9xCXNt0_0),.dout(w_dff_B_7lA60dox5_0),.clk(gclk));
	jdff dff_B_LRZkUum75_0(.din(w_dff_B_7lA60dox5_0),.dout(w_dff_B_LRZkUum75_0),.clk(gclk));
	jdff dff_B_9at1ByCj6_0(.din(w_dff_B_LRZkUum75_0),.dout(w_dff_B_9at1ByCj6_0),.clk(gclk));
	jdff dff_B_LR86h8DS1_0(.din(w_dff_B_9at1ByCj6_0),.dout(w_dff_B_LR86h8DS1_0),.clk(gclk));
	jdff dff_B_hfsJQ9OX6_0(.din(w_dff_B_LR86h8DS1_0),.dout(w_dff_B_hfsJQ9OX6_0),.clk(gclk));
	jdff dff_B_MyhW5Q118_0(.din(w_dff_B_hfsJQ9OX6_0),.dout(w_dff_B_MyhW5Q118_0),.clk(gclk));
	jdff dff_B_ZMGHqk8a6_0(.din(w_dff_B_MyhW5Q118_0),.dout(w_dff_B_ZMGHqk8a6_0),.clk(gclk));
	jdff dff_B_qLP4lseT5_0(.din(w_dff_B_ZMGHqk8a6_0),.dout(w_dff_B_qLP4lseT5_0),.clk(gclk));
	jdff dff_B_f6ms2hRU9_0(.din(n1270),.dout(w_dff_B_f6ms2hRU9_0),.clk(gclk));
	jdff dff_B_jRX7vECG9_2(.din(G103),.dout(w_dff_B_jRX7vECG9_2),.clk(gclk));
	jdff dff_B_O70naEaZ5_2(.din(G100),.dout(w_dff_B_O70naEaZ5_2),.clk(gclk));
	jdff dff_B_8Yyyj7RI1_2(.din(w_dff_B_O70naEaZ5_2),.dout(w_dff_B_8Yyyj7RI1_2),.clk(gclk));
	jdff dff_A_SjmIzxNS3_0(.dout(w_n840_2[0]),.din(w_dff_A_SjmIzxNS3_0),.clk(gclk));
	jdff dff_B_oEHMjoZM4_0(.din(n1279),.dout(w_dff_B_oEHMjoZM4_0),.clk(gclk));
	jdff dff_B_0UVXI1LF8_0(.din(w_dff_B_oEHMjoZM4_0),.dout(w_dff_B_0UVXI1LF8_0),.clk(gclk));
	jdff dff_B_1JF1dcMV9_0(.din(w_dff_B_0UVXI1LF8_0),.dout(w_dff_B_1JF1dcMV9_0),.clk(gclk));
	jdff dff_B_qlGZLACm0_0(.din(n1278),.dout(w_dff_B_qlGZLACm0_0),.clk(gclk));
	jdff dff_B_o3RAEwwq5_0(.din(w_dff_B_qlGZLACm0_0),.dout(w_dff_B_o3RAEwwq5_0),.clk(gclk));
	jdff dff_B_GIm0chOL1_0(.din(w_dff_B_o3RAEwwq5_0),.dout(w_dff_B_GIm0chOL1_0),.clk(gclk));
	jdff dff_B_m7Qul1kx6_0(.din(w_dff_B_GIm0chOL1_0),.dout(w_dff_B_m7Qul1kx6_0),.clk(gclk));
	jdff dff_B_QU5O1tk84_0(.din(w_dff_B_m7Qul1kx6_0),.dout(w_dff_B_QU5O1tk84_0),.clk(gclk));
	jdff dff_B_blxjcLSa4_0(.din(w_dff_B_QU5O1tk84_0),.dout(w_dff_B_blxjcLSa4_0),.clk(gclk));
	jdff dff_B_ojJnp0J70_0(.din(w_dff_B_blxjcLSa4_0),.dout(w_dff_B_ojJnp0J70_0),.clk(gclk));
	jdff dff_B_kBUkPofw5_0(.din(w_dff_B_ojJnp0J70_0),.dout(w_dff_B_kBUkPofw5_0),.clk(gclk));
	jdff dff_B_T1l0oZsW6_0(.din(w_dff_B_kBUkPofw5_0),.dout(w_dff_B_T1l0oZsW6_0),.clk(gclk));
	jdff dff_B_d8DnDGOF9_0(.din(w_dff_B_T1l0oZsW6_0),.dout(w_dff_B_d8DnDGOF9_0),.clk(gclk));
	jdff dff_B_q20txiL02_0(.din(n1277),.dout(w_dff_B_q20txiL02_0),.clk(gclk));
	jdff dff_B_zXfMPo1R6_2(.din(G40),.dout(w_dff_B_zXfMPo1R6_2),.clk(gclk));
	jdff dff_B_MQq2MLku5_2(.din(G91),.dout(w_dff_B_MQq2MLku5_2),.clk(gclk));
	jdff dff_B_kYuYIcMt3_2(.din(w_dff_B_MQq2MLku5_2),.dout(w_dff_B_kYuYIcMt3_2),.clk(gclk));
	jdff dff_B_ZOzHQm2o8_0(.din(n1286),.dout(w_dff_B_ZOzHQm2o8_0),.clk(gclk));
	jdff dff_B_ERsYOr3c9_0(.din(w_dff_B_ZOzHQm2o8_0),.dout(w_dff_B_ERsYOr3c9_0),.clk(gclk));
	jdff dff_B_m3koI63o4_0(.din(w_dff_B_ERsYOr3c9_0),.dout(w_dff_B_m3koI63o4_0),.clk(gclk));
	jdff dff_B_uzBL3Vhi0_0(.din(n1285),.dout(w_dff_B_uzBL3Vhi0_0),.clk(gclk));
	jdff dff_B_5xB5dWrk5_0(.din(w_dff_B_uzBL3Vhi0_0),.dout(w_dff_B_5xB5dWrk5_0),.clk(gclk));
	jdff dff_B_5xbZSuV02_0(.din(w_dff_B_5xB5dWrk5_0),.dout(w_dff_B_5xbZSuV02_0),.clk(gclk));
	jdff dff_B_ICvipmzU5_0(.din(w_dff_B_5xbZSuV02_0),.dout(w_dff_B_ICvipmzU5_0),.clk(gclk));
	jdff dff_B_wmcbES5X2_0(.din(w_dff_B_ICvipmzU5_0),.dout(w_dff_B_wmcbES5X2_0),.clk(gclk));
	jdff dff_B_5jxlTNV85_0(.din(w_dff_B_wmcbES5X2_0),.dout(w_dff_B_5jxlTNV85_0),.clk(gclk));
	jdff dff_B_njHTkLKH5_0(.din(w_dff_B_5jxlTNV85_0),.dout(w_dff_B_njHTkLKH5_0),.clk(gclk));
	jdff dff_B_2dSk21kk0_0(.din(w_dff_B_njHTkLKH5_0),.dout(w_dff_B_2dSk21kk0_0),.clk(gclk));
	jdff dff_B_6swa5yUS6_0(.din(w_dff_B_2dSk21kk0_0),.dout(w_dff_B_6swa5yUS6_0),.clk(gclk));
	jdff dff_B_Lv9JQ9Y06_0(.din(w_dff_B_6swa5yUS6_0),.dout(w_dff_B_Lv9JQ9Y06_0),.clk(gclk));
	jdff dff_B_Cx88I4iO0_0(.din(n1284),.dout(w_dff_B_Cx88I4iO0_0),.clk(gclk));
	jdff dff_A_vITD7vPb0_0(.dout(w_G137_6[0]),.din(w_dff_A_vITD7vPb0_0),.clk(gclk));
	jdff dff_A_WbwDnkIO3_0(.dout(w_dff_A_vITD7vPb0_0),.din(w_dff_A_WbwDnkIO3_0),.clk(gclk));
	jdff dff_A_8JoHe52a3_0(.dout(w_dff_A_WbwDnkIO3_0),.din(w_dff_A_8JoHe52a3_0),.clk(gclk));
	jdff dff_B_lbHHsTzM8_0(.din(n1294),.dout(w_dff_B_lbHHsTzM8_0),.clk(gclk));
	jdff dff_B_b5kwYdD60_0(.din(w_dff_B_lbHHsTzM8_0),.dout(w_dff_B_b5kwYdD60_0),.clk(gclk));
	jdff dff_B_Uw33huRr7_0(.din(w_dff_B_b5kwYdD60_0),.dout(w_dff_B_Uw33huRr7_0),.clk(gclk));
	jdff dff_B_vLBJNzGY0_0(.din(n1293),.dout(w_dff_B_vLBJNzGY0_0),.clk(gclk));
	jdff dff_B_iA9bVtkV3_0(.din(w_dff_B_vLBJNzGY0_0),.dout(w_dff_B_iA9bVtkV3_0),.clk(gclk));
	jdff dff_B_NsB6g8zc0_0(.din(w_dff_B_iA9bVtkV3_0),.dout(w_dff_B_NsB6g8zc0_0),.clk(gclk));
	jdff dff_B_4wiyKpNu5_0(.din(w_dff_B_NsB6g8zc0_0),.dout(w_dff_B_4wiyKpNu5_0),.clk(gclk));
	jdff dff_B_0rJSfrYf8_0(.din(w_dff_B_4wiyKpNu5_0),.dout(w_dff_B_0rJSfrYf8_0),.clk(gclk));
	jdff dff_B_Wue1VuDB7_0(.din(w_dff_B_0rJSfrYf8_0),.dout(w_dff_B_Wue1VuDB7_0),.clk(gclk));
	jdff dff_B_DbWznKL27_0(.din(w_dff_B_Wue1VuDB7_0),.dout(w_dff_B_DbWznKL27_0),.clk(gclk));
	jdff dff_B_gPUORSrF9_0(.din(w_dff_B_DbWznKL27_0),.dout(w_dff_B_gPUORSrF9_0),.clk(gclk));
	jdff dff_B_xcUtQedf4_0(.din(w_dff_B_gPUORSrF9_0),.dout(w_dff_B_xcUtQedf4_0),.clk(gclk));
	jdff dff_B_BgYH8FIF4_0(.din(n1292),.dout(w_dff_B_BgYH8FIF4_0),.clk(gclk));
	jdff dff_B_Ng6Rn8W99_0(.din(n1302),.dout(w_dff_B_Ng6Rn8W99_0),.clk(gclk));
	jdff dff_B_U6uAs9no9_0(.din(w_dff_B_Ng6Rn8W99_0),.dout(w_dff_B_U6uAs9no9_0),.clk(gclk));
	jdff dff_B_7Wj7KvJt5_0(.din(n1301),.dout(w_dff_B_7Wj7KvJt5_0),.clk(gclk));
	jdff dff_B_V0vbzK4e1_0(.din(w_dff_B_7Wj7KvJt5_0),.dout(w_dff_B_V0vbzK4e1_0),.clk(gclk));
	jdff dff_B_NsRBJ3iU3_0(.din(w_dff_B_V0vbzK4e1_0),.dout(w_dff_B_NsRBJ3iU3_0),.clk(gclk));
	jdff dff_B_zNKGFW5e9_0(.din(w_dff_B_NsRBJ3iU3_0),.dout(w_dff_B_zNKGFW5e9_0),.clk(gclk));
	jdff dff_B_zV1Q3ny67_0(.din(w_dff_B_zNKGFW5e9_0),.dout(w_dff_B_zV1Q3ny67_0),.clk(gclk));
	jdff dff_B_TQMcUYh46_0(.din(w_dff_B_zV1Q3ny67_0),.dout(w_dff_B_TQMcUYh46_0),.clk(gclk));
	jdff dff_B_9i2GNllg1_0(.din(w_dff_B_TQMcUYh46_0),.dout(w_dff_B_9i2GNllg1_0),.clk(gclk));
	jdff dff_B_XGpEbwUZ0_0(.din(w_dff_B_9i2GNllg1_0),.dout(w_dff_B_XGpEbwUZ0_0),.clk(gclk));
	jdff dff_B_fdPo0AZw9_0(.din(w_dff_B_XGpEbwUZ0_0),.dout(w_dff_B_fdPo0AZw9_0),.clk(gclk));
	jdff dff_B_2NvQOqmD9_0(.din(n1300),.dout(w_dff_B_2NvQOqmD9_0),.clk(gclk));
	jdff dff_A_rrTVTbpo5_2(.dout(w_n988_2[2]),.din(w_dff_A_rrTVTbpo5_2),.clk(gclk));
	jdff dff_A_BdZzNksn6_1(.dout(w_n985_2[1]),.din(w_dff_A_BdZzNksn6_1),.clk(gclk));
	jdff dff_A_BWQGC92m1_2(.dout(w_n985_2[2]),.din(w_dff_A_BWQGC92m1_2),.clk(gclk));
	jdff dff_A_ECbPHj9f5_2(.dout(w_dff_A_BWQGC92m1_2),.din(w_dff_A_ECbPHj9f5_2),.clk(gclk));
	jdff dff_B_gOi5EzOj8_0(.din(n1310),.dout(w_dff_B_gOi5EzOj8_0),.clk(gclk));
	jdff dff_B_EtmPvepO1_0(.din(w_dff_B_gOi5EzOj8_0),.dout(w_dff_B_EtmPvepO1_0),.clk(gclk));
	jdff dff_B_G2h9uHxD4_0(.din(n1309),.dout(w_dff_B_G2h9uHxD4_0),.clk(gclk));
	jdff dff_B_F4yeVIzN2_0(.din(w_dff_B_G2h9uHxD4_0),.dout(w_dff_B_F4yeVIzN2_0),.clk(gclk));
	jdff dff_B_ayUldVDk7_0(.din(w_dff_B_F4yeVIzN2_0),.dout(w_dff_B_ayUldVDk7_0),.clk(gclk));
	jdff dff_B_weEEwUjX6_0(.din(w_dff_B_ayUldVDk7_0),.dout(w_dff_B_weEEwUjX6_0),.clk(gclk));
	jdff dff_B_A0rIVWEu8_0(.din(w_dff_B_weEEwUjX6_0),.dout(w_dff_B_A0rIVWEu8_0),.clk(gclk));
	jdff dff_B_8KsF5R416_0(.din(w_dff_B_A0rIVWEu8_0),.dout(w_dff_B_8KsF5R416_0),.clk(gclk));
	jdff dff_B_yoXsPQ4H1_0(.din(w_dff_B_8KsF5R416_0),.dout(w_dff_B_yoXsPQ4H1_0),.clk(gclk));
	jdff dff_B_Lu8lYJLh5_0(.din(w_dff_B_yoXsPQ4H1_0),.dout(w_dff_B_Lu8lYJLh5_0),.clk(gclk));
	jdff dff_B_iU3KJzgu0_0(.din(w_dff_B_Lu8lYJLh5_0),.dout(w_dff_B_iU3KJzgu0_0),.clk(gclk));
	jdff dff_B_o5e6IOru5_0(.din(n1308),.dout(w_dff_B_o5e6IOru5_0),.clk(gclk));
	jdff dff_A_8i5JmseF1_2(.dout(w_G137_5[2]),.din(w_dff_A_8i5JmseF1_2),.clk(gclk));
	jdff dff_B_oedsz4iZ2_0(.din(n1318),.dout(w_dff_B_oedsz4iZ2_0),.clk(gclk));
	jdff dff_B_hw9IJ1Bl2_0(.din(w_dff_B_oedsz4iZ2_0),.dout(w_dff_B_hw9IJ1Bl2_0),.clk(gclk));
	jdff dff_B_x5UCoTEU2_0(.din(w_dff_B_hw9IJ1Bl2_0),.dout(w_dff_B_x5UCoTEU2_0),.clk(gclk));
	jdff dff_B_NLSYKpBl1_0(.din(n1317),.dout(w_dff_B_NLSYKpBl1_0),.clk(gclk));
	jdff dff_B_plyQ8HPL6_0(.din(w_dff_B_NLSYKpBl1_0),.dout(w_dff_B_plyQ8HPL6_0),.clk(gclk));
	jdff dff_B_1U7ck2i94_0(.din(w_dff_B_plyQ8HPL6_0),.dout(w_dff_B_1U7ck2i94_0),.clk(gclk));
	jdff dff_B_feDNCScj2_0(.din(w_dff_B_1U7ck2i94_0),.dout(w_dff_B_feDNCScj2_0),.clk(gclk));
	jdff dff_B_yefaxNen0_0(.din(w_dff_B_feDNCScj2_0),.dout(w_dff_B_yefaxNen0_0),.clk(gclk));
	jdff dff_B_visyYMWp4_0(.din(w_dff_B_yefaxNen0_0),.dout(w_dff_B_visyYMWp4_0),.clk(gclk));
	jdff dff_B_j9G7auJy6_0(.din(w_dff_B_visyYMWp4_0),.dout(w_dff_B_j9G7auJy6_0),.clk(gclk));
	jdff dff_B_NgGmCUIL6_0(.din(w_dff_B_j9G7auJy6_0),.dout(w_dff_B_NgGmCUIL6_0),.clk(gclk));
	jdff dff_B_Krh0mYAU6_0(.din(w_dff_B_NgGmCUIL6_0),.dout(w_dff_B_Krh0mYAU6_0),.clk(gclk));
	jdff dff_B_tiqgSRIB6_0(.din(w_dff_B_Krh0mYAU6_0),.dout(w_dff_B_tiqgSRIB6_0),.clk(gclk));
	jdff dff_B_4PSQfdGY6_0(.din(n1316),.dout(w_dff_B_4PSQfdGY6_0),.clk(gclk));
	jdff dff_B_YPRdsmVb0_2(.din(G173),.dout(w_dff_B_YPRdsmVb0_2),.clk(gclk));
	jdff dff_B_kI74GGDN6_2(.din(G203),.dout(w_dff_B_kI74GGDN6_2),.clk(gclk));
	jdff dff_B_dLHRqh202_2(.din(w_dff_B_kI74GGDN6_2),.dout(w_dff_B_dLHRqh202_2),.clk(gclk));
	jdff dff_B_eFZn4Thj1_0(.din(n1182),.dout(w_dff_B_eFZn4Thj1_0),.clk(gclk));
	jdff dff_B_LJAJG16A1_0(.din(w_dff_B_eFZn4Thj1_0),.dout(w_dff_B_LJAJG16A1_0),.clk(gclk));
	jdff dff_B_JeW58ZwZ2_0(.din(w_dff_B_LJAJG16A1_0),.dout(w_dff_B_JeW58ZwZ2_0),.clk(gclk));
	jdff dff_B_AMqtIJq76_0(.din(w_dff_B_JeW58ZwZ2_0),.dout(w_dff_B_AMqtIJq76_0),.clk(gclk));
	jdff dff_B_SiShHYSa7_0(.din(w_dff_B_AMqtIJq76_0),.dout(w_dff_B_SiShHYSa7_0),.clk(gclk));
	jdff dff_B_rriyiCdb7_1(.din(n1179),.dout(w_dff_B_rriyiCdb7_1),.clk(gclk));
	jdff dff_B_QskXEO8H8_1(.din(G112),.dout(w_dff_B_QskXEO8H8_1),.clk(gclk));
	jdff dff_B_E0lFfosK4_1(.din(w_dff_B_QskXEO8H8_1),.dout(w_dff_B_E0lFfosK4_1),.clk(gclk));
	jdff dff_B_Vz1ntBHV2_0(.din(n1218),.dout(w_dff_B_Vz1ntBHV2_0),.clk(gclk));
	jdff dff_B_6B5mhpyF8_0(.din(w_dff_B_Vz1ntBHV2_0),.dout(w_dff_B_6B5mhpyF8_0),.clk(gclk));
	jdff dff_B_zhPGh3cK0_0(.din(w_dff_B_6B5mhpyF8_0),.dout(w_dff_B_zhPGh3cK0_0),.clk(gclk));
	jdff dff_B_eAaYpwze3_0(.din(w_dff_B_zhPGh3cK0_0),.dout(w_dff_B_eAaYpwze3_0),.clk(gclk));
	jdff dff_B_COuRIf2v1_0(.din(w_dff_B_eAaYpwze3_0),.dout(w_dff_B_COuRIf2v1_0),.clk(gclk));
	jdff dff_B_dtmJ3N519_0(.din(w_dff_B_COuRIf2v1_0),.dout(w_dff_B_dtmJ3N519_0),.clk(gclk));
	jdff dff_B_ISnxJlzE9_0(.din(w_dff_B_dtmJ3N519_0),.dout(w_dff_B_ISnxJlzE9_0),.clk(gclk));
	jdff dff_B_LaggcDo98_0(.din(w_dff_B_ISnxJlzE9_0),.dout(w_dff_B_LaggcDo98_0),.clk(gclk));
	jdff dff_B_1XCOXLIU0_1(.din(n1215),.dout(w_dff_B_1XCOXLIU0_1),.clk(gclk));
	jdff dff_B_PYLWk6ka0_1(.din(G113),.dout(w_dff_B_PYLWk6ka0_1),.clk(gclk));
	jdff dff_B_JdJmN8DZ9_1(.din(w_dff_B_PYLWk6ka0_1),.dout(w_dff_B_JdJmN8DZ9_1),.clk(gclk));
	jdff dff_B_SlI5zjop1_0(.din(n538),.dout(w_dff_B_SlI5zjop1_0),.clk(gclk));
	jdff dff_B_acpYoPnv5_0(.din(n1326),.dout(w_dff_B_acpYoPnv5_0),.clk(gclk));
	jdff dff_B_fzyS4ZHU6_0(.din(w_dff_B_acpYoPnv5_0),.dout(w_dff_B_fzyS4ZHU6_0),.clk(gclk));
	jdff dff_B_faGCYL2X9_0(.din(w_dff_B_fzyS4ZHU6_0),.dout(w_dff_B_faGCYL2X9_0),.clk(gclk));
	jdff dff_B_whRg3B451_0(.din(n1325),.dout(w_dff_B_whRg3B451_0),.clk(gclk));
	jdff dff_B_WqSqG6bc3_0(.din(w_dff_B_whRg3B451_0),.dout(w_dff_B_WqSqG6bc3_0),.clk(gclk));
	jdff dff_B_YmxtpP3m7_0(.din(w_dff_B_WqSqG6bc3_0),.dout(w_dff_B_YmxtpP3m7_0),.clk(gclk));
	jdff dff_B_5eds7RG33_0(.din(w_dff_B_YmxtpP3m7_0),.dout(w_dff_B_5eds7RG33_0),.clk(gclk));
	jdff dff_B_udGgoTHc8_0(.din(w_dff_B_5eds7RG33_0),.dout(w_dff_B_udGgoTHc8_0),.clk(gclk));
	jdff dff_B_hERHpCd72_0(.din(w_dff_B_udGgoTHc8_0),.dout(w_dff_B_hERHpCd72_0),.clk(gclk));
	jdff dff_B_Gh8s5APZ8_0(.din(w_dff_B_hERHpCd72_0),.dout(w_dff_B_Gh8s5APZ8_0),.clk(gclk));
	jdff dff_B_PCWCeHBx3_0(.din(w_dff_B_Gh8s5APZ8_0),.dout(w_dff_B_PCWCeHBx3_0),.clk(gclk));
	jdff dff_B_Eeolb1wv2_0(.din(w_dff_B_PCWCeHBx3_0),.dout(w_dff_B_Eeolb1wv2_0),.clk(gclk));
	jdff dff_B_vy9ULEa11_0(.din(n1324),.dout(w_dff_B_vy9ULEa11_0),.clk(gclk));
	jdff dff_B_hpxdS3QY5_2(.din(G167),.dout(w_dff_B_hpxdS3QY5_2),.clk(gclk));
	jdff dff_B_MFi49ebU8_2(.din(G197),.dout(w_dff_B_MFi49ebU8_2),.clk(gclk));
	jdff dff_B_rCprmroI2_2(.din(w_dff_B_MFi49ebU8_2),.dout(w_dff_B_rCprmroI2_2),.clk(gclk));
	jdff dff_B_GMkp0s0z6_0(.din(n1175),.dout(w_dff_B_GMkp0s0z6_0),.clk(gclk));
	jdff dff_B_Pp4FAqis2_0(.din(w_dff_B_GMkp0s0z6_0),.dout(w_dff_B_Pp4FAqis2_0),.clk(gclk));
	jdff dff_B_mhjMIrs43_0(.din(w_dff_B_Pp4FAqis2_0),.dout(w_dff_B_mhjMIrs43_0),.clk(gclk));
	jdff dff_B_D43eyW007_0(.din(w_dff_B_mhjMIrs43_0),.dout(w_dff_B_D43eyW007_0),.clk(gclk));
	jdff dff_B_lyCXxF103_1(.din(n1172),.dout(w_dff_B_lyCXxF103_1),.clk(gclk));
	jdff dff_B_Olgdvryu5_1(.din(G116),.dout(w_dff_B_Olgdvryu5_1),.clk(gclk));
	jdff dff_B_R5eMOqaD7_1(.din(w_dff_B_Olgdvryu5_1),.dout(w_dff_B_R5eMOqaD7_1),.clk(gclk));
	jdff dff_A_rIWRxbCO5_1(.dout(w_n971_0[1]),.din(w_dff_A_rIWRxbCO5_1),.clk(gclk));
	jdff dff_A_05jXUVYb5_1(.dout(w_dff_A_rIWRxbCO5_1),.din(w_dff_A_05jXUVYb5_1),.clk(gclk));
	jdff dff_B_AbC2ilUe7_1(.din(n967),.dout(w_dff_B_AbC2ilUe7_1),.clk(gclk));
	jdff dff_B_JRvU0wqr5_1(.din(w_dff_B_AbC2ilUe7_1),.dout(w_dff_B_JRvU0wqr5_1),.clk(gclk));
	jdff dff_B_KRYrmHnS6_1(.din(w_dff_B_JRvU0wqr5_1),.dout(w_dff_B_KRYrmHnS6_1),.clk(gclk));
	jdff dff_B_jfGC3CN29_1(.din(w_dff_B_KRYrmHnS6_1),.dout(w_dff_B_jfGC3CN29_1),.clk(gclk));
	jdff dff_B_raw05elo1_0(.din(n1211),.dout(w_dff_B_raw05elo1_0),.clk(gclk));
	jdff dff_B_HH4FIpVi3_0(.din(w_dff_B_raw05elo1_0),.dout(w_dff_B_HH4FIpVi3_0),.clk(gclk));
	jdff dff_B_IEpRikXA7_0(.din(w_dff_B_HH4FIpVi3_0),.dout(w_dff_B_IEpRikXA7_0),.clk(gclk));
	jdff dff_B_3pjLBGFh6_0(.din(w_dff_B_IEpRikXA7_0),.dout(w_dff_B_3pjLBGFh6_0),.clk(gclk));
	jdff dff_B_nXu5OdZo0_0(.din(w_dff_B_3pjLBGFh6_0),.dout(w_dff_B_nXu5OdZo0_0),.clk(gclk));
	jdff dff_B_3iC6jjnK9_0(.din(w_dff_B_nXu5OdZo0_0),.dout(w_dff_B_3iC6jjnK9_0),.clk(gclk));
	jdff dff_B_XiAZqJNi4_0(.din(w_dff_B_3iC6jjnK9_0),.dout(w_dff_B_XiAZqJNi4_0),.clk(gclk));
	jdff dff_B_UrrZoGXb3_1(.din(n1208),.dout(w_dff_B_UrrZoGXb3_1),.clk(gclk));
	jdff dff_B_8aI5nUHz3_1(.din(G53),.dout(w_dff_B_8aI5nUHz3_1),.clk(gclk));
	jdff dff_B_EreY5MCq2_1(.din(w_dff_B_8aI5nUHz3_1),.dout(w_dff_B_EreY5MCq2_1),.clk(gclk));
	jdff dff_B_VcxDnBYM0_0(.din(n515),.dout(w_dff_B_VcxDnBYM0_0),.clk(gclk));
	jdff dff_A_jmZ7L2ae0_1(.dout(w_n953_0[1]),.din(w_dff_A_jmZ7L2ae0_1),.clk(gclk));
	jdff dff_A_wjn5Vn6R9_1(.dout(w_dff_A_jmZ7L2ae0_1),.din(w_dff_A_wjn5Vn6R9_1),.clk(gclk));
	jdff dff_B_Dgj4G4vl7_1(.din(n949),.dout(w_dff_B_Dgj4G4vl7_1),.clk(gclk));
	jdff dff_B_zWvbwJsk7_1(.din(w_dff_B_Dgj4G4vl7_1),.dout(w_dff_B_zWvbwJsk7_1),.clk(gclk));
	jdff dff_B_fjTAuQFX2_1(.din(w_dff_B_zWvbwJsk7_1),.dout(w_dff_B_fjTAuQFX2_1),.clk(gclk));
	jdff dff_B_p7N3tSMZ1_1(.din(w_dff_B_fjTAuQFX2_1),.dout(w_dff_B_p7N3tSMZ1_1),.clk(gclk));
	jdff dff_B_1B5dW4gv3_1(.din(w_dff_B_p7N3tSMZ1_1),.dout(w_dff_B_1B5dW4gv3_1),.clk(gclk));
	jdff dff_B_U8qdlVqH8_1(.din(w_dff_B_1B5dW4gv3_1),.dout(w_dff_B_U8qdlVqH8_1),.clk(gclk));
	jdff dff_B_B2VgIguc1_1(.din(w_dff_B_U8qdlVqH8_1),.dout(w_dff_B_B2VgIguc1_1),.clk(gclk));
	jdff dff_B_0RClE1oJ5_1(.din(w_dff_B_B2VgIguc1_1),.dout(w_dff_B_0RClE1oJ5_1),.clk(gclk));
	jdff dff_B_5MI8Awnl5_1(.din(n950),.dout(w_dff_B_5MI8Awnl5_1),.clk(gclk));
	jdff dff_B_5Z2NNARz1_1(.din(w_dff_B_5MI8Awnl5_1),.dout(w_dff_B_5Z2NNARz1_1),.clk(gclk));
	jdff dff_B_z4wiDlmQ1_1(.din(w_dff_B_5Z2NNARz1_1),.dout(w_dff_B_z4wiDlmQ1_1),.clk(gclk));
	jdff dff_B_WREghjRO3_1(.din(w_dff_B_z4wiDlmQ1_1),.dout(w_dff_B_WREghjRO3_1),.clk(gclk));
	jdff dff_B_Tmuo6mTq9_1(.din(w_dff_B_WREghjRO3_1),.dout(w_dff_B_Tmuo6mTq9_1),.clk(gclk));
	jdff dff_B_rNTWf0vb8_1(.din(w_dff_B_Tmuo6mTq9_1),.dout(w_dff_B_rNTWf0vb8_1),.clk(gclk));
	jdff dff_A_WqzXDVaw3_1(.dout(w_n748_1[1]),.din(w_dff_A_WqzXDVaw3_1),.clk(gclk));
	jdff dff_A_6XXnUosv2_1(.dout(w_dff_A_WqzXDVaw3_1),.din(w_dff_A_6XXnUosv2_1),.clk(gclk));
	jdff dff_A_mOrcPzMO3_1(.dout(w_dff_A_6XXnUosv2_1),.din(w_dff_A_mOrcPzMO3_1),.clk(gclk));
	jdff dff_A_xnKGH3WI2_1(.dout(w_dff_A_mOrcPzMO3_1),.din(w_dff_A_xnKGH3WI2_1),.clk(gclk));
	jdff dff_A_fr2wMieK9_1(.dout(w_dff_A_xnKGH3WI2_1),.din(w_dff_A_fr2wMieK9_1),.clk(gclk));
	jdff dff_A_PhT7RjdB1_1(.dout(w_dff_A_fr2wMieK9_1),.din(w_dff_A_PhT7RjdB1_1),.clk(gclk));
	jdff dff_A_Hl0Q5VCh0_1(.dout(w_dff_A_PhT7RjdB1_1),.din(w_dff_A_Hl0Q5VCh0_1),.clk(gclk));
	jdff dff_A_z36PlgSe5_1(.dout(w_dff_A_Hl0Q5VCh0_1),.din(w_dff_A_z36PlgSe5_1),.clk(gclk));
	jdff dff_A_fXiwjX984_1(.dout(w_dff_A_z36PlgSe5_1),.din(w_dff_A_fXiwjX984_1),.clk(gclk));
	jdff dff_A_WRWLsXku9_2(.dout(w_n748_1[2]),.din(w_dff_A_WRWLsXku9_2),.clk(gclk));
	jdff dff_A_MXDRsjqQ0_2(.dout(w_dff_A_WRWLsXku9_2),.din(w_dff_A_MXDRsjqQ0_2),.clk(gclk));
	jdff dff_A_KJjsWf3F7_2(.dout(w_dff_A_MXDRsjqQ0_2),.din(w_dff_A_KJjsWf3F7_2),.clk(gclk));
	jdff dff_A_zEXBvlxm0_2(.dout(w_dff_A_KJjsWf3F7_2),.din(w_dff_A_zEXBvlxm0_2),.clk(gclk));
	jdff dff_A_TNNwyAnz4_2(.dout(w_dff_A_zEXBvlxm0_2),.din(w_dff_A_TNNwyAnz4_2),.clk(gclk));
	jdff dff_A_sWLOdO185_2(.dout(w_dff_A_TNNwyAnz4_2),.din(w_dff_A_sWLOdO185_2),.clk(gclk));
	jdff dff_B_22OVXIZw7_0(.din(n1334),.dout(w_dff_B_22OVXIZw7_0),.clk(gclk));
	jdff dff_B_OeLX3bdT2_0(.din(w_dff_B_22OVXIZw7_0),.dout(w_dff_B_OeLX3bdT2_0),.clk(gclk));
	jdff dff_B_pq6GNIyG0_0(.din(n1333),.dout(w_dff_B_pq6GNIyG0_0),.clk(gclk));
	jdff dff_B_iDlfVGcF8_0(.din(w_dff_B_pq6GNIyG0_0),.dout(w_dff_B_iDlfVGcF8_0),.clk(gclk));
	jdff dff_B_qJPRHBPH9_0(.din(w_dff_B_iDlfVGcF8_0),.dout(w_dff_B_qJPRHBPH9_0),.clk(gclk));
	jdff dff_B_yP90QQdN5_0(.din(w_dff_B_qJPRHBPH9_0),.dout(w_dff_B_yP90QQdN5_0),.clk(gclk));
	jdff dff_B_yJYsWwSD7_0(.din(w_dff_B_yP90QQdN5_0),.dout(w_dff_B_yJYsWwSD7_0),.clk(gclk));
	jdff dff_B_pJYulsn07_0(.din(w_dff_B_yJYsWwSD7_0),.dout(w_dff_B_pJYulsn07_0),.clk(gclk));
	jdff dff_B_pJF4Jypo6_0(.din(w_dff_B_pJYulsn07_0),.dout(w_dff_B_pJF4Jypo6_0),.clk(gclk));
	jdff dff_B_SFnz6RF04_0(.din(w_dff_B_pJF4Jypo6_0),.dout(w_dff_B_SFnz6RF04_0),.clk(gclk));
	jdff dff_B_TeA0l5RY6_0(.din(w_dff_B_SFnz6RF04_0),.dout(w_dff_B_TeA0l5RY6_0),.clk(gclk));
	jdff dff_B_q8GF83v79_0(.din(n1332),.dout(w_dff_B_q8GF83v79_0),.clk(gclk));
	jdff dff_B_U9xFB3tu4_2(.din(G164),.dout(w_dff_B_U9xFB3tu4_2),.clk(gclk));
	jdff dff_B_Q4LtkL6W1_2(.din(G194),.dout(w_dff_B_Q4LtkL6W1_2),.clk(gclk));
	jdff dff_B_4OU2SCCW1_2(.din(w_dff_B_Q4LtkL6W1_2),.dout(w_dff_B_4OU2SCCW1_2),.clk(gclk));
	jdff dff_B_dUgtlIFV2_0(.din(n1169),.dout(w_dff_B_dUgtlIFV2_0),.clk(gclk));
	jdff dff_B_9xqbSwPw2_0(.din(w_dff_B_dUgtlIFV2_0),.dout(w_dff_B_9xqbSwPw2_0),.clk(gclk));
	jdff dff_B_zHdPq9Yi6_0(.din(w_dff_B_9xqbSwPw2_0),.dout(w_dff_B_zHdPq9Yi6_0),.clk(gclk));
	jdff dff_B_JtyCeYB62_0(.din(w_dff_B_zHdPq9Yi6_0),.dout(w_dff_B_JtyCeYB62_0),.clk(gclk));
	jdff dff_B_A49QF9CZ7_0(.din(w_dff_B_JtyCeYB62_0),.dout(w_dff_B_A49QF9CZ7_0),.clk(gclk));
	jdff dff_B_OSHN10nK3_1(.din(G121),.dout(w_dff_B_OSHN10nK3_1),.clk(gclk));
	jdff dff_B_cnWEupaI2_1(.din(w_dff_B_OSHN10nK3_1),.dout(w_dff_B_cnWEupaI2_1),.clk(gclk));
	jdff dff_A_EQbq1Jpa1_1(.dout(w_n972_0[1]),.din(w_dff_A_EQbq1Jpa1_1),.clk(gclk));
	jdff dff_A_Fh9xh3C97_1(.dout(w_n748_2[1]),.din(w_dff_A_Fh9xh3C97_1),.clk(gclk));
	jdff dff_A_zTdByzIN4_2(.dout(w_n748_2[2]),.din(w_dff_A_zTdByzIN4_2),.clk(gclk));
	jdff dff_A_GzU8HWgG0_2(.dout(w_dff_A_zTdByzIN4_2),.din(w_dff_A_GzU8HWgG0_2),.clk(gclk));
	jdff dff_A_1hnT5ZfW1_1(.dout(w_n748_0[1]),.din(w_dff_A_1hnT5ZfW1_1),.clk(gclk));
	jdff dff_A_YzYrO1eU3_1(.dout(w_dff_A_1hnT5ZfW1_1),.din(w_dff_A_YzYrO1eU3_1),.clk(gclk));
	jdff dff_A_fKMKsLFO5_1(.dout(w_dff_A_YzYrO1eU3_1),.din(w_dff_A_fKMKsLFO5_1),.clk(gclk));
	jdff dff_A_1sHSKFOe3_1(.dout(w_dff_A_fKMKsLFO5_1),.din(w_dff_A_1sHSKFOe3_1),.clk(gclk));
	jdff dff_A_Ubk7zqdW1_1(.dout(w_dff_A_1sHSKFOe3_1),.din(w_dff_A_Ubk7zqdW1_1),.clk(gclk));
	jdff dff_A_DAWyJfAl7_1(.dout(w_dff_A_Ubk7zqdW1_1),.din(w_dff_A_DAWyJfAl7_1),.clk(gclk));
	jdff dff_A_9d8L8x0H4_2(.dout(w_n748_0[2]),.din(w_dff_A_9d8L8x0H4_2),.clk(gclk));
	jdff dff_A_SjxSNAMP4_2(.dout(w_dff_A_9d8L8x0H4_2),.din(w_dff_A_SjxSNAMP4_2),.clk(gclk));
	jdff dff_A_wCrRRJR36_2(.dout(w_dff_A_SjxSNAMP4_2),.din(w_dff_A_wCrRRJR36_2),.clk(gclk));
	jdff dff_A_r18v1tHD8_0(.dout(w_n747_3[0]),.din(w_dff_A_r18v1tHD8_0),.clk(gclk));
	jdff dff_A_x23Z2iOW2_0(.dout(w_dff_A_r18v1tHD8_0),.din(w_dff_A_x23Z2iOW2_0),.clk(gclk));
	jdff dff_A_sFJ45rlF1_0(.dout(w_dff_A_x23Z2iOW2_0),.din(w_dff_A_sFJ45rlF1_0),.clk(gclk));
	jdff dff_A_0Ocy39pC6_0(.dout(w_dff_A_sFJ45rlF1_0),.din(w_dff_A_0Ocy39pC6_0),.clk(gclk));
	jdff dff_A_hjZUStJG5_0(.dout(w_dff_A_0Ocy39pC6_0),.din(w_dff_A_hjZUStJG5_0),.clk(gclk));
	jdff dff_A_SS5FoYVk2_0(.dout(w_dff_A_hjZUStJG5_0),.din(w_dff_A_SS5FoYVk2_0),.clk(gclk));
	jdff dff_A_Hw5wbg2B0_1(.dout(w_n747_3[1]),.din(w_dff_A_Hw5wbg2B0_1),.clk(gclk));
	jdff dff_A_1fLKU9vB1_1(.dout(w_dff_A_Hw5wbg2B0_1),.din(w_dff_A_1fLKU9vB1_1),.clk(gclk));
	jdff dff_A_KzcxDb729_2(.dout(w_n1002_2[2]),.din(w_dff_A_KzcxDb729_2),.clk(gclk));
	jdff dff_B_li6rMYPd0_0(.din(n1204),.dout(w_dff_B_li6rMYPd0_0),.clk(gclk));
	jdff dff_B_ARaiKiPd6_0(.din(w_dff_B_li6rMYPd0_0),.dout(w_dff_B_ARaiKiPd6_0),.clk(gclk));
	jdff dff_B_3qpbMsdT4_0(.din(w_dff_B_ARaiKiPd6_0),.dout(w_dff_B_3qpbMsdT4_0),.clk(gclk));
	jdff dff_B_hx5DLAU38_0(.din(w_dff_B_3qpbMsdT4_0),.dout(w_dff_B_hx5DLAU38_0),.clk(gclk));
	jdff dff_B_FjyRfDIm0_0(.din(w_dff_B_hx5DLAU38_0),.dout(w_dff_B_FjyRfDIm0_0),.clk(gclk));
	jdff dff_B_tYWbr3Pe8_0(.din(w_dff_B_FjyRfDIm0_0),.dout(w_dff_B_tYWbr3Pe8_0),.clk(gclk));
	jdff dff_B_y5jcS6ZD3_0(.din(w_dff_B_tYWbr3Pe8_0),.dout(w_dff_B_y5jcS6ZD3_0),.clk(gclk));
	jdff dff_B_GDnjo22a3_1(.din(n1200),.dout(w_dff_B_GDnjo22a3_1),.clk(gclk));
	jdff dff_B_nDROfitL5_1(.din(G114),.dout(w_dff_B_nDROfitL5_1),.clk(gclk));
	jdff dff_B_nyZz9qgn8_1(.din(w_dff_B_nDROfitL5_1),.dout(w_dff_B_nyZz9qgn8_1),.clk(gclk));
	jdff dff_B_VQfTMgXa2_0(.din(n549),.dout(w_dff_B_VQfTMgXa2_0),.clk(gclk));
	jdff dff_B_slQjwQXb7_3(.din(G3548),.dout(w_dff_B_slQjwQXb7_3),.clk(gclk));
	jdff dff_A_SAJWWZnn5_1(.dout(w_n999_2[1]),.din(w_dff_A_SAJWWZnn5_1),.clk(gclk));
	jdff dff_A_Id5oNvbB0_2(.dout(w_n999_2[2]),.din(w_dff_A_Id5oNvbB0_2),.clk(gclk));
	jdff dff_A_4jcnKlLF8_2(.dout(w_dff_A_Id5oNvbB0_2),.din(w_dff_A_4jcnKlLF8_2),.clk(gclk));
	jdff dff_A_GSkyqbtI8_1(.dout(w_G137_4[1]),.din(w_dff_A_GSkyqbtI8_1),.clk(gclk));
	jdff dff_A_XRpTZvDQ0_2(.dout(w_G137_4[2]),.din(w_dff_A_XRpTZvDQ0_2),.clk(gclk));
	jdff dff_A_ENGhT1wc6_2(.dout(w_dff_A_XRpTZvDQ0_2),.din(w_dff_A_ENGhT1wc6_2),.clk(gclk));
	jdff dff_A_vm4mmnSs7_0(.dout(w_G137_1[0]),.din(w_dff_A_vm4mmnSs7_0),.clk(gclk));
	jdff dff_A_LW3Zr75J1_1(.dout(w_G137_1[1]),.din(w_dff_A_LW3Zr75J1_1),.clk(gclk));
	jdff dff_B_M7SHGnkw8_0(.din(n1342),.dout(w_dff_B_M7SHGnkw8_0),.clk(gclk));
	jdff dff_B_qtFJrn8I0_0(.din(w_dff_B_M7SHGnkw8_0),.dout(w_dff_B_qtFJrn8I0_0),.clk(gclk));
	jdff dff_B_8cBj3oOq5_0(.din(n1341),.dout(w_dff_B_8cBj3oOq5_0),.clk(gclk));
	jdff dff_B_5c0bILSV0_0(.din(w_dff_B_8cBj3oOq5_0),.dout(w_dff_B_5c0bILSV0_0),.clk(gclk));
	jdff dff_B_oTNeUFKQ7_0(.din(w_dff_B_5c0bILSV0_0),.dout(w_dff_B_oTNeUFKQ7_0),.clk(gclk));
	jdff dff_B_e8YAPToP2_0(.din(w_dff_B_oTNeUFKQ7_0),.dout(w_dff_B_e8YAPToP2_0),.clk(gclk));
	jdff dff_B_M4zknGzF3_0(.din(w_dff_B_e8YAPToP2_0),.dout(w_dff_B_M4zknGzF3_0),.clk(gclk));
	jdff dff_B_p9MjM4yu6_0(.din(w_dff_B_M4zknGzF3_0),.dout(w_dff_B_p9MjM4yu6_0),.clk(gclk));
	jdff dff_B_xf6O3MZo7_0(.din(w_dff_B_p9MjM4yu6_0),.dout(w_dff_B_xf6O3MZo7_0),.clk(gclk));
	jdff dff_B_YAPnp2Q61_0(.din(w_dff_B_xf6O3MZo7_0),.dout(w_dff_B_YAPnp2Q61_0),.clk(gclk));
	jdff dff_B_yy97jijI8_0(.din(w_dff_B_YAPnp2Q61_0),.dout(w_dff_B_yy97jijI8_0),.clk(gclk));
	jdff dff_B_VdR7OR9Q3_0(.din(n1340),.dout(w_dff_B_VdR7OR9Q3_0),.clk(gclk));
	jdff dff_B_2SbTkK094_2(.din(G161),.dout(w_dff_B_2SbTkK094_2),.clk(gclk));
	jdff dff_B_TiplbXo39_2(.din(G191),.dout(w_dff_B_TiplbXo39_2),.clk(gclk));
	jdff dff_B_cpaVajUF2_2(.din(w_dff_B_TiplbXo39_2),.dout(w_dff_B_cpaVajUF2_2),.clk(gclk));
	jdff dff_B_HfFaPkC65_0(.din(n1162),.dout(w_dff_B_HfFaPkC65_0),.clk(gclk));
	jdff dff_B_8XrlRDYx1_0(.din(w_dff_B_HfFaPkC65_0),.dout(w_dff_B_8XrlRDYx1_0),.clk(gclk));
	jdff dff_B_O1Otu4Kr7_0(.din(w_dff_B_8XrlRDYx1_0),.dout(w_dff_B_O1Otu4Kr7_0),.clk(gclk));
	jdff dff_B_ZkgHXbfY0_0(.din(w_dff_B_O1Otu4Kr7_0),.dout(w_dff_B_ZkgHXbfY0_0),.clk(gclk));
	jdff dff_B_BNivMpSa4_0(.din(w_dff_B_ZkgHXbfY0_0),.dout(w_dff_B_BNivMpSa4_0),.clk(gclk));
	jdff dff_B_tiF4XvPQ7_0(.din(w_dff_B_BNivMpSa4_0),.dout(w_dff_B_tiF4XvPQ7_0),.clk(gclk));
	jdff dff_B_qUG4y7cK7_0(.din(w_dff_B_tiF4XvPQ7_0),.dout(w_dff_B_qUG4y7cK7_0),.clk(gclk));
	jdff dff_B_OMwLOQoe0_1(.din(n1160),.dout(w_dff_B_OMwLOQoe0_1),.clk(gclk));
	jdff dff_A_1tQJNjSy6_1(.dout(w_n751_1[1]),.din(w_dff_A_1tQJNjSy6_1),.clk(gclk));
	jdff dff_A_Pny1KaRT0_0(.dout(w_G123_0[0]),.din(w_dff_A_Pny1KaRT0_0),.clk(gclk));
	jdff dff_B_PL0GQhlg7_2(.din(G123),.dout(w_dff_B_PL0GQhlg7_2),.clk(gclk));
	jdff dff_B_4bhq2NKq5_0(.din(n788),.dout(w_dff_B_4bhq2NKq5_0),.clk(gclk));
	jdff dff_A_8ttTp3Vi9_1(.dout(w_n633_1[1]),.din(w_dff_A_8ttTp3Vi9_1),.clk(gclk));
	jdff dff_A_gJmCSXsn7_0(.dout(w_G54_0[0]),.din(w_dff_A_gJmCSXsn7_0),.clk(gclk));
	jdff dff_A_StlX5KTO3_0(.dout(w_dff_A_gJmCSXsn7_0),.din(w_dff_A_StlX5KTO3_0),.clk(gclk));
	jdff dff_A_fw76MlPt4_0(.dout(w_dff_A_StlX5KTO3_0),.din(w_dff_A_fw76MlPt4_0),.clk(gclk));
	jdff dff_A_2pMiESGr0_0(.dout(w_dff_A_fw76MlPt4_0),.din(w_dff_A_2pMiESGr0_0),.clk(gclk));
	jdff dff_A_ro6qKbEt7_0(.dout(w_dff_A_2pMiESGr0_0),.din(w_dff_A_ro6qKbEt7_0),.clk(gclk));
	jdff dff_A_6Dvk6O510_0(.dout(w_dff_A_ro6qKbEt7_0),.din(w_dff_A_6Dvk6O510_0),.clk(gclk));
	jdff dff_A_J5FJNJKh7_0(.dout(w_n741_0[0]),.din(w_dff_A_J5FJNJKh7_0),.clk(gclk));
	jdff dff_B_jDCZofNF4_2(.din(n741),.dout(w_dff_B_jDCZofNF4_2),.clk(gclk));
	jdff dff_A_llMijzDi0_1(.dout(w_n747_2[1]),.din(w_dff_A_llMijzDi0_1),.clk(gclk));
	jdff dff_A_WSi3kZeY5_1(.dout(w_dff_A_llMijzDi0_1),.din(w_dff_A_WSi3kZeY5_1),.clk(gclk));
	jdff dff_B_kiRT4vhG2_0(.din(n1196),.dout(w_dff_B_kiRT4vhG2_0),.clk(gclk));
	jdff dff_B_g3wjCMSv3_0(.din(w_dff_B_kiRT4vhG2_0),.dout(w_dff_B_g3wjCMSv3_0),.clk(gclk));
	jdff dff_B_rsSuToCT0_0(.din(w_dff_B_g3wjCMSv3_0),.dout(w_dff_B_rsSuToCT0_0),.clk(gclk));
	jdff dff_B_3gfUOwFb5_0(.din(w_dff_B_rsSuToCT0_0),.dout(w_dff_B_3gfUOwFb5_0),.clk(gclk));
	jdff dff_B_OZTkSiqQ5_0(.din(w_dff_B_3gfUOwFb5_0),.dout(w_dff_B_OZTkSiqQ5_0),.clk(gclk));
	jdff dff_B_RiEGixy43_0(.din(w_dff_B_OZTkSiqQ5_0),.dout(w_dff_B_RiEGixy43_0),.clk(gclk));
	jdff dff_B_W7HNd5l65_0(.din(w_dff_B_RiEGixy43_0),.dout(w_dff_B_W7HNd5l65_0),.clk(gclk));
	jdff dff_B_J5kFLssw3_0(.din(w_dff_B_W7HNd5l65_0),.dout(w_dff_B_J5kFLssw3_0),.clk(gclk));
	jdff dff_B_RJFQge1i7_0(.din(n1195),.dout(w_dff_B_RJFQge1i7_0),.clk(gclk));
	jdff dff_B_e9P0BzYN6_0(.din(w_dff_B_RJFQge1i7_0),.dout(w_dff_B_e9P0BzYN6_0),.clk(gclk));
	jdff dff_B_0I6h65H62_1(.din(G115),.dout(w_dff_B_0I6h65H62_1),.clk(gclk));
	jdff dff_B_wxWIjnjD9_1(.din(w_dff_B_0I6h65H62_1),.dout(w_dff_B_wxWIjnjD9_1),.clk(gclk));
	jdff dff_A_ggzm7CIh2_2(.dout(w_n751_0[2]),.din(w_dff_A_ggzm7CIh2_2),.clk(gclk));
	jdff dff_A_SGJuPREI6_2(.dout(w_dff_A_ggzm7CIh2_2),.din(w_dff_A_SGJuPREI6_2),.clk(gclk));
	jdff dff_B_KTjZAv1M5_1(.din(n929),.dout(w_dff_B_KTjZAv1M5_1),.clk(gclk));
	jdff dff_B_vex8H1gp2_1(.din(w_dff_B_KTjZAv1M5_1),.dout(w_dff_B_vex8H1gp2_1),.clk(gclk));
	jdff dff_B_XZUn9BKN5_1(.din(w_dff_B_vex8H1gp2_1),.dout(w_dff_B_XZUn9BKN5_1),.clk(gclk));
	jdff dff_B_nrpAOopt1_1(.din(w_dff_B_XZUn9BKN5_1),.dout(w_dff_B_nrpAOopt1_1),.clk(gclk));
	jdff dff_B_9viapTLL6_1(.din(n931),.dout(w_dff_B_9viapTLL6_1),.clk(gclk));
	jdff dff_B_IjVSjQ8n3_1(.din(w_dff_B_9viapTLL6_1),.dout(w_dff_B_IjVSjQ8n3_1),.clk(gclk));
	jdff dff_B_6o6s6cOq5_1(.din(w_dff_B_IjVSjQ8n3_1),.dout(w_dff_B_6o6s6cOq5_1),.clk(gclk));
	jdff dff_B_zFkwWUqm1_1(.din(w_dff_B_6o6s6cOq5_1),.dout(w_dff_B_zFkwWUqm1_1),.clk(gclk));
	jdff dff_B_W6tnOw9y0_1(.din(w_dff_B_zFkwWUqm1_1),.dout(w_dff_B_W6tnOw9y0_1),.clk(gclk));
	jdff dff_B_fQWhak0j7_1(.din(w_dff_B_W6tnOw9y0_1),.dout(w_dff_B_fQWhak0j7_1),.clk(gclk));
	jdff dff_A_W5XI0bWh9_1(.dout(w_G4_0[1]),.din(w_dff_A_W5XI0bWh9_1),.clk(gclk));
	jdff dff_A_WCcbNtYi1_1(.dout(w_dff_A_W5XI0bWh9_1),.din(w_dff_A_WCcbNtYi1_1),.clk(gclk));
	jdff dff_A_9sdbsVg40_1(.dout(w_dff_A_WCcbNtYi1_1),.din(w_dff_A_9sdbsVg40_1),.clk(gclk));
	jdff dff_A_MNXxV7ES6_1(.dout(w_dff_A_9sdbsVg40_1),.din(w_dff_A_MNXxV7ES6_1),.clk(gclk));
	jdff dff_B_TibwFOW81_3(.din(G4),.dout(w_dff_B_TibwFOW81_3),.clk(gclk));
	jdff dff_B_pX7f7LqH6_3(.din(w_dff_B_TibwFOW81_3),.dout(w_dff_B_pX7f7LqH6_3),.clk(gclk));
	jdff dff_B_gTmA6XQD6_3(.din(w_dff_B_pX7f7LqH6_3),.dout(w_dff_B_gTmA6XQD6_3),.clk(gclk));
	jdff dff_B_QjCsz9SH9_2(.din(n932),.dout(w_dff_B_QjCsz9SH9_2),.clk(gclk));
	jdff dff_B_RcmgbfyC8_2(.din(w_dff_B_QjCsz9SH9_2),.dout(w_dff_B_RcmgbfyC8_2),.clk(gclk));
	jdff dff_B_9EKcqnJ09_2(.din(w_dff_B_RcmgbfyC8_2),.dout(w_dff_B_9EKcqnJ09_2),.clk(gclk));
	jdff dff_B_bzelxDXV2_2(.din(w_dff_B_9EKcqnJ09_2),.dout(w_dff_B_bzelxDXV2_2),.clk(gclk));
	jdff dff_B_VIoBQoCF0_2(.din(w_dff_B_bzelxDXV2_2),.dout(w_dff_B_VIoBQoCF0_2),.clk(gclk));
	jdff dff_B_N3N1Y1jD7_2(.din(w_dff_B_VIoBQoCF0_2),.dout(w_dff_B_N3N1Y1jD7_2),.clk(gclk));
	jdff dff_A_DxmC90yB9_1(.dout(w_n747_1[1]),.din(w_dff_A_DxmC90yB9_1),.clk(gclk));
	jdff dff_A_7X10HfUW9_2(.dout(w_n747_1[2]),.din(w_dff_A_7X10HfUW9_2),.clk(gclk));
	jdff dff_A_mgsbhz6J6_0(.dout(w_n747_0[0]),.din(w_dff_A_mgsbhz6J6_0),.clk(gclk));
	jdff dff_A_m7oKYewi8_0(.dout(w_dff_A_mgsbhz6J6_0),.din(w_dff_A_m7oKYewi8_0),.clk(gclk));
	jdff dff_A_JUZSiVxA0_0(.dout(w_dff_A_m7oKYewi8_0),.din(w_dff_A_JUZSiVxA0_0),.clk(gclk));
	jdff dff_A_7nP5QKik0_0(.dout(w_dff_A_JUZSiVxA0_0),.din(w_dff_A_7nP5QKik0_0),.clk(gclk));
	jdff dff_A_mgfZHYHO8_0(.dout(w_dff_A_7nP5QKik0_0),.din(w_dff_A_mgfZHYHO8_0),.clk(gclk));
	jdff dff_A_mxBuZMhX9_0(.dout(w_dff_A_mgfZHYHO8_0),.din(w_dff_A_mxBuZMhX9_0),.clk(gclk));
	jdff dff_A_6jB4SwTD5_0(.dout(w_dff_A_mxBuZMhX9_0),.din(w_dff_A_6jB4SwTD5_0),.clk(gclk));
	jdff dff_A_K7Di0Uvu6_0(.dout(w_dff_A_6jB4SwTD5_0),.din(w_dff_A_K7Di0Uvu6_0),.clk(gclk));
	jdff dff_A_cENZyIIS1_0(.dout(w_dff_A_K7Di0Uvu6_0),.din(w_dff_A_cENZyIIS1_0),.clk(gclk));
	jdff dff_A_HlGmURBk0_1(.dout(w_n747_0[1]),.din(w_dff_A_HlGmURBk0_1),.clk(gclk));
	jdff dff_A_HKYxXTwe9_1(.dout(w_dff_A_HlGmURBk0_1),.din(w_dff_A_HKYxXTwe9_1),.clk(gclk));
	jdff dff_A_fUcf2fqC9_1(.dout(w_dff_A_HKYxXTwe9_1),.din(w_dff_A_fUcf2fqC9_1),.clk(gclk));
	jdff dff_A_shtfT2Pp1_1(.dout(w_dff_A_fUcf2fqC9_1),.din(w_dff_A_shtfT2Pp1_1),.clk(gclk));
	jdff dff_A_93Tmmsg90_1(.dout(w_dff_A_shtfT2Pp1_1),.din(w_dff_A_93Tmmsg90_1),.clk(gclk));
	jdff dff_A_RIpPmYAd8_1(.dout(w_dff_A_93Tmmsg90_1),.din(w_dff_A_RIpPmYAd8_1),.clk(gclk));
	jdff dff_B_i3FsJUr95_1(.din(n1388),.dout(w_dff_B_i3FsJUr95_1),.clk(gclk));
	jdff dff_B_fFwXDLlc1_1(.din(w_dff_B_i3FsJUr95_1),.dout(w_dff_B_fFwXDLlc1_1),.clk(gclk));
	jdff dff_B_E3RDMGLX3_1(.din(w_dff_B_fFwXDLlc1_1),.dout(w_dff_B_E3RDMGLX3_1),.clk(gclk));
	jdff dff_B_uOuoRYtZ2_1(.din(w_dff_B_E3RDMGLX3_1),.dout(w_dff_B_uOuoRYtZ2_1),.clk(gclk));
	jdff dff_B_NUJRDPGh3_1(.din(w_dff_B_uOuoRYtZ2_1),.dout(w_dff_B_NUJRDPGh3_1),.clk(gclk));
	jdff dff_B_mtu0Bx9L3_1(.din(w_dff_B_NUJRDPGh3_1),.dout(w_dff_B_mtu0Bx9L3_1),.clk(gclk));
	jdff dff_B_UcVSyL2i5_1(.din(w_dff_B_mtu0Bx9L3_1),.dout(w_dff_B_UcVSyL2i5_1),.clk(gclk));
	jdff dff_B_e4YOXTGO5_1(.din(w_dff_B_UcVSyL2i5_1),.dout(w_dff_B_e4YOXTGO5_1),.clk(gclk));
	jdff dff_B_yxfhv4Fa6_1(.din(w_dff_B_e4YOXTGO5_1),.dout(w_dff_B_yxfhv4Fa6_1),.clk(gclk));
	jdff dff_B_5zC0WoXC2_1(.din(w_dff_B_yxfhv4Fa6_1),.dout(w_dff_B_5zC0WoXC2_1),.clk(gclk));
	jdff dff_B_LgoqLde44_1(.din(w_dff_B_5zC0WoXC2_1),.dout(w_dff_B_LgoqLde44_1),.clk(gclk));
	jdff dff_B_zAIAJcVN6_1(.din(w_dff_B_LgoqLde44_1),.dout(w_dff_B_zAIAJcVN6_1),.clk(gclk));
	jdff dff_B_B99ennDR0_0(.din(n1345),.dout(w_dff_B_B99ennDR0_0),.clk(gclk));
	jdff dff_B_bFOj7a0R4_1(.din(n1539),.dout(w_dff_B_bFOj7a0R4_1),.clk(gclk));
	jdff dff_B_6sM8oGHm0_1(.din(w_dff_B_bFOj7a0R4_1),.dout(w_dff_B_6sM8oGHm0_1),.clk(gclk));
	jdff dff_B_B1UYFk2o4_1(.din(w_dff_B_6sM8oGHm0_1),.dout(w_dff_B_B1UYFk2o4_1),.clk(gclk));
	jdff dff_B_Nq54T7Ky9_1(.din(w_dff_B_B1UYFk2o4_1),.dout(w_dff_B_Nq54T7Ky9_1),.clk(gclk));
	jdff dff_B_QPDnPbRd3_1(.din(w_dff_B_Nq54T7Ky9_1),.dout(w_dff_B_QPDnPbRd3_1),.clk(gclk));
	jdff dff_B_RauW5Vu18_1(.din(w_dff_B_QPDnPbRd3_1),.dout(w_dff_B_RauW5Vu18_1),.clk(gclk));
	jdff dff_B_MJdzDbaa6_1(.din(w_dff_B_RauW5Vu18_1),.dout(w_dff_B_MJdzDbaa6_1),.clk(gclk));
	jdff dff_B_EBoRtQx52_1(.din(w_dff_B_MJdzDbaa6_1),.dout(w_dff_B_EBoRtQx52_1),.clk(gclk));
	jdff dff_B_fuFAjgps1_1(.din(w_dff_B_EBoRtQx52_1),.dout(w_dff_B_fuFAjgps1_1),.clk(gclk));
	jdff dff_B_zgPyu6ru9_1(.din(w_dff_B_fuFAjgps1_1),.dout(w_dff_B_zgPyu6ru9_1),.clk(gclk));
	jdff dff_B_pbz0Cmqh4_1(.din(w_dff_B_zgPyu6ru9_1),.dout(w_dff_B_pbz0Cmqh4_1),.clk(gclk));
	jdff dff_B_FtthFBnC9_1(.din(w_dff_B_pbz0Cmqh4_1),.dout(w_dff_B_FtthFBnC9_1),.clk(gclk));
	jdff dff_B_fPpq6yDu9_1(.din(w_dff_B_FtthFBnC9_1),.dout(w_dff_B_fPpq6yDu9_1),.clk(gclk));
	jdff dff_B_wicwbTDi0_1(.din(w_dff_B_fPpq6yDu9_1),.dout(w_dff_B_wicwbTDi0_1),.clk(gclk));
	jdff dff_B_Pyyd8abY6_1(.din(w_dff_B_wicwbTDi0_1),.dout(w_dff_B_Pyyd8abY6_1),.clk(gclk));
	jdff dff_B_htnjqMlm6_0(.din(n1454),.dout(w_dff_B_htnjqMlm6_0),.clk(gclk));
	jdff dff_B_BGFZewS63_0(.din(n1615),.dout(w_dff_B_BGFZewS63_0),.clk(gclk));
	jdff dff_B_5ctXP9eo4_0(.din(w_dff_B_BGFZewS63_0),.dout(w_dff_B_5ctXP9eo4_0),.clk(gclk));
	jdff dff_B_VkhQF9W88_0(.din(w_dff_B_5ctXP9eo4_0),.dout(w_dff_B_VkhQF9W88_0),.clk(gclk));
	jdff dff_B_hdMl9aRK1_0(.din(w_dff_B_VkhQF9W88_0),.dout(w_dff_B_hdMl9aRK1_0),.clk(gclk));
	jdff dff_B_8sUGvrK17_0(.din(w_dff_B_hdMl9aRK1_0),.dout(w_dff_B_8sUGvrK17_0),.clk(gclk));
	jdff dff_B_nCk8U6TP4_0(.din(n1614),.dout(w_dff_B_nCk8U6TP4_0),.clk(gclk));
	jdff dff_B_PRMxhqAJ0_0(.din(w_dff_B_nCk8U6TP4_0),.dout(w_dff_B_PRMxhqAJ0_0),.clk(gclk));
	jdff dff_B_sjSsXpMB5_0(.din(w_dff_B_PRMxhqAJ0_0),.dout(w_dff_B_sjSsXpMB5_0),.clk(gclk));
	jdff dff_B_e6Z5c8AC5_0(.din(w_dff_B_sjSsXpMB5_0),.dout(w_dff_B_e6Z5c8AC5_0),.clk(gclk));
	jdff dff_B_JTD7njZr3_0(.din(w_dff_B_e6Z5c8AC5_0),.dout(w_dff_B_JTD7njZr3_0),.clk(gclk));
	jdff dff_B_FZlu4RZA7_0(.din(w_dff_B_JTD7njZr3_0),.dout(w_dff_B_FZlu4RZA7_0),.clk(gclk));
	jdff dff_B_1M3YZdXG6_0(.din(w_dff_B_FZlu4RZA7_0),.dout(w_dff_B_1M3YZdXG6_0),.clk(gclk));
	jdff dff_B_KHEGqgld8_0(.din(w_dff_B_1M3YZdXG6_0),.dout(w_dff_B_KHEGqgld8_0),.clk(gclk));
	jdff dff_B_qVVUs1qO2_0(.din(w_dff_B_KHEGqgld8_0),.dout(w_dff_B_qVVUs1qO2_0),.clk(gclk));
	jdff dff_B_7vOvb3sI0_0(.din(w_dff_B_qVVUs1qO2_0),.dout(w_dff_B_7vOvb3sI0_0),.clk(gclk));
	jdff dff_B_1A9Un1F09_0(.din(w_dff_B_7vOvb3sI0_0),.dout(w_dff_B_1A9Un1F09_0),.clk(gclk));
	jdff dff_B_VGR9opvU0_0(.din(n1613),.dout(w_dff_B_VGR9opvU0_0),.clk(gclk));
	jdff dff_A_Rhc3tDM80_1(.dout(w_n797_1[1]),.din(w_dff_A_Rhc3tDM80_1),.clk(gclk));
	jdff dff_A_H3oBqD3L7_1(.dout(w_dff_A_Rhc3tDM80_1),.din(w_dff_A_H3oBqD3L7_1),.clk(gclk));
	jdff dff_A_xerHdk6D7_1(.dout(w_dff_A_H3oBqD3L7_1),.din(w_dff_A_xerHdk6D7_1),.clk(gclk));
	jdff dff_A_ZgTFHJnh9_1(.dout(w_dff_A_xerHdk6D7_1),.din(w_dff_A_ZgTFHJnh9_1),.clk(gclk));
	jdff dff_A_f3qoZ7Cz7_1(.dout(w_dff_A_ZgTFHJnh9_1),.din(w_dff_A_f3qoZ7Cz7_1),.clk(gclk));
	jdff dff_A_MYL3Ibh64_1(.dout(w_dff_A_f3qoZ7Cz7_1),.din(w_dff_A_MYL3Ibh64_1),.clk(gclk));
	jdff dff_A_ZFvdDV6w3_1(.dout(w_dff_A_MYL3Ibh64_1),.din(w_dff_A_ZFvdDV6w3_1),.clk(gclk));
	jdff dff_A_RfCGG9Om0_2(.dout(w_n797_1[2]),.din(w_dff_A_RfCGG9Om0_2),.clk(gclk));
	jdff dff_A_wid5fOrc7_2(.dout(w_dff_A_RfCGG9Om0_2),.din(w_dff_A_wid5fOrc7_2),.clk(gclk));
	jdff dff_A_nVSbX7wO5_2(.dout(w_dff_A_wid5fOrc7_2),.din(w_dff_A_nVSbX7wO5_2),.clk(gclk));
	jdff dff_A_eTvjzC3E2_2(.dout(w_dff_A_nVSbX7wO5_2),.din(w_dff_A_eTvjzC3E2_2),.clk(gclk));
	jdff dff_A_llyazwr65_2(.dout(w_dff_A_eTvjzC3E2_2),.din(w_dff_A_llyazwr65_2),.clk(gclk));
	jdff dff_A_bAjPhM2N9_2(.dout(w_dff_A_llyazwr65_2),.din(w_dff_A_bAjPhM2N9_2),.clk(gclk));
	jdff dff_A_k3WV8kxG7_1(.dout(w_n797_0[1]),.din(w_dff_A_k3WV8kxG7_1),.clk(gclk));
	jdff dff_A_OYUtI3739_1(.dout(w_dff_A_k3WV8kxG7_1),.din(w_dff_A_OYUtI3739_1),.clk(gclk));
	jdff dff_A_rwkBpeNA8_1(.dout(w_dff_A_OYUtI3739_1),.din(w_dff_A_rwkBpeNA8_1),.clk(gclk));
	jdff dff_A_XqzPCH1w8_1(.dout(w_dff_A_rwkBpeNA8_1),.din(w_dff_A_XqzPCH1w8_1),.clk(gclk));
	jdff dff_A_QS2IeYwS3_1(.dout(w_dff_A_XqzPCH1w8_1),.din(w_dff_A_QS2IeYwS3_1),.clk(gclk));
	jdff dff_A_Zckhoghx0_2(.dout(w_n797_0[2]),.din(w_dff_A_Zckhoghx0_2),.clk(gclk));
	jdff dff_B_YSXjY3xx5_3(.din(n797),.dout(w_dff_B_YSXjY3xx5_3),.clk(gclk));
	jdff dff_B_HB2DzWmL0_3(.din(w_dff_B_YSXjY3xx5_3),.dout(w_dff_B_HB2DzWmL0_3),.clk(gclk));
	jdff dff_B_vpIeW4oQ2_3(.din(w_dff_B_HB2DzWmL0_3),.dout(w_dff_B_vpIeW4oQ2_3),.clk(gclk));
	jdff dff_B_7IGwgqcQ8_3(.din(w_dff_B_vpIeW4oQ2_3),.dout(w_dff_B_7IGwgqcQ8_3),.clk(gclk));
	jdff dff_A_iUZuXxWP7_1(.dout(w_n793_1[1]),.din(w_dff_A_iUZuXxWP7_1),.clk(gclk));
	jdff dff_A_VanVvJhj2_1(.dout(w_dff_A_iUZuXxWP7_1),.din(w_dff_A_VanVvJhj2_1),.clk(gclk));
	jdff dff_A_CxN3yo6u0_1(.dout(w_dff_A_VanVvJhj2_1),.din(w_dff_A_CxN3yo6u0_1),.clk(gclk));
	jdff dff_A_rFFwgffD7_1(.dout(w_dff_A_CxN3yo6u0_1),.din(w_dff_A_rFFwgffD7_1),.clk(gclk));
	jdff dff_A_I9MJSD190_1(.dout(w_dff_A_rFFwgffD7_1),.din(w_dff_A_I9MJSD190_1),.clk(gclk));
	jdff dff_A_QlZOPNq30_1(.dout(w_dff_A_I9MJSD190_1),.din(w_dff_A_QlZOPNq30_1),.clk(gclk));
	jdff dff_A_bHmzluzP8_1(.dout(w_dff_A_QlZOPNq30_1),.din(w_dff_A_bHmzluzP8_1),.clk(gclk));
	jdff dff_A_jpRvdR2a4_1(.dout(w_dff_A_bHmzluzP8_1),.din(w_dff_A_jpRvdR2a4_1),.clk(gclk));
	jdff dff_A_OqdiTg7f4_1(.dout(w_dff_A_jpRvdR2a4_1),.din(w_dff_A_OqdiTg7f4_1),.clk(gclk));
	jdff dff_A_2W8pSPwQ6_1(.dout(w_dff_A_OqdiTg7f4_1),.din(w_dff_A_2W8pSPwQ6_1),.clk(gclk));
	jdff dff_A_lnjU3B0F6_2(.dout(w_n793_1[2]),.din(w_dff_A_lnjU3B0F6_2),.clk(gclk));
	jdff dff_A_iq8ABI189_2(.dout(w_dff_A_lnjU3B0F6_2),.din(w_dff_A_iq8ABI189_2),.clk(gclk));
	jdff dff_A_E4OTRdCl7_2(.dout(w_dff_A_iq8ABI189_2),.din(w_dff_A_E4OTRdCl7_2),.clk(gclk));
	jdff dff_A_Uo3QZuGO4_2(.dout(w_dff_A_E4OTRdCl7_2),.din(w_dff_A_Uo3QZuGO4_2),.clk(gclk));
	jdff dff_A_jJ6AozAY6_2(.dout(w_dff_A_Uo3QZuGO4_2),.din(w_dff_A_jJ6AozAY6_2),.clk(gclk));
	jdff dff_A_8pvUP4jg8_2(.dout(w_dff_A_jJ6AozAY6_2),.din(w_dff_A_8pvUP4jg8_2),.clk(gclk));
	jdff dff_A_j7BaaYgz3_2(.dout(w_dff_A_8pvUP4jg8_2),.din(w_dff_A_j7BaaYgz3_2),.clk(gclk));
	jdff dff_A_1cCJGC275_1(.dout(w_n793_0[1]),.din(w_dff_A_1cCJGC275_1),.clk(gclk));
	jdff dff_A_tbNhpOKQ3_1(.dout(w_dff_A_1cCJGC275_1),.din(w_dff_A_tbNhpOKQ3_1),.clk(gclk));
	jdff dff_A_XbVu0WMF1_1(.dout(w_dff_A_tbNhpOKQ3_1),.din(w_dff_A_XbVu0WMF1_1),.clk(gclk));
	jdff dff_A_u2MqTlpg8_1(.dout(w_dff_A_XbVu0WMF1_1),.din(w_dff_A_u2MqTlpg8_1),.clk(gclk));
	jdff dff_A_CLCfiF5u8_1(.dout(w_dff_A_u2MqTlpg8_1),.din(w_dff_A_CLCfiF5u8_1),.clk(gclk));
	jdff dff_A_l6LMCiKm3_2(.dout(w_n793_0[2]),.din(w_dff_A_l6LMCiKm3_2),.clk(gclk));
	jdff dff_A_8Mno0JcQ7_2(.dout(w_dff_A_l6LMCiKm3_2),.din(w_dff_A_8Mno0JcQ7_2),.clk(gclk));
	jdff dff_A_PDsmLccJ7_2(.dout(w_dff_A_8Mno0JcQ7_2),.din(w_dff_A_PDsmLccJ7_2),.clk(gclk));
	jdff dff_A_1vCY42P70_2(.dout(w_dff_A_PDsmLccJ7_2),.din(w_dff_A_1vCY42P70_2),.clk(gclk));
	jdff dff_B_YmYQRpHf4_3(.din(n793),.dout(w_dff_B_YmYQRpHf4_3),.clk(gclk));
	jdff dff_B_B6H4VXy27_3(.din(w_dff_B_YmYQRpHf4_3),.dout(w_dff_B_B6H4VXy27_3),.clk(gclk));
	jdff dff_B_gqD19LCf9_3(.din(w_dff_B_B6H4VXy27_3),.dout(w_dff_B_gqD19LCf9_3),.clk(gclk));
	jdff dff_B_NpdFLm1V0_3(.din(w_dff_B_gqD19LCf9_3),.dout(w_dff_B_NpdFLm1V0_3),.clk(gclk));
	jdff dff_B_r4PTKkIp0_3(.din(w_dff_B_NpdFLm1V0_3),.dout(w_dff_B_r4PTKkIp0_3),.clk(gclk));
	jdff dff_B_W0wuerbt5_3(.din(w_dff_B_r4PTKkIp0_3),.dout(w_dff_B_W0wuerbt5_3),.clk(gclk));
	jdff dff_A_D88n27GW8_2(.dout(w_G4088_0[2]),.din(w_dff_A_D88n27GW8_2),.clk(gclk));
	jdff dff_A_PjTDWTfI7_1(.dout(w_G4087_0[1]),.din(w_dff_A_PjTDWTfI7_1),.clk(gclk));
	jdff dff_B_IyXlR4hY7_0(.din(n1622),.dout(w_dff_B_IyXlR4hY7_0),.clk(gclk));
	jdff dff_B_ZLtLf6e24_0(.din(w_dff_B_IyXlR4hY7_0),.dout(w_dff_B_ZLtLf6e24_0),.clk(gclk));
	jdff dff_B_qNgk59pk6_0(.din(w_dff_B_ZLtLf6e24_0),.dout(w_dff_B_qNgk59pk6_0),.clk(gclk));
	jdff dff_B_3WrV56Wd1_0(.din(w_dff_B_qNgk59pk6_0),.dout(w_dff_B_3WrV56Wd1_0),.clk(gclk));
	jdff dff_B_hOPT3Yyh1_0(.din(w_dff_B_3WrV56Wd1_0),.dout(w_dff_B_hOPT3Yyh1_0),.clk(gclk));
	jdff dff_B_wnElaByr2_0(.din(n1621),.dout(w_dff_B_wnElaByr2_0),.clk(gclk));
	jdff dff_B_JxVXYiaX8_0(.din(w_dff_B_wnElaByr2_0),.dout(w_dff_B_JxVXYiaX8_0),.clk(gclk));
	jdff dff_B_GV2db3OD6_0(.din(w_dff_B_JxVXYiaX8_0),.dout(w_dff_B_GV2db3OD6_0),.clk(gclk));
	jdff dff_B_V0ZsOrIP0_0(.din(w_dff_B_GV2db3OD6_0),.dout(w_dff_B_V0ZsOrIP0_0),.clk(gclk));
	jdff dff_B_pVj1v5wW0_0(.din(w_dff_B_V0ZsOrIP0_0),.dout(w_dff_B_pVj1v5wW0_0),.clk(gclk));
	jdff dff_B_YYdSncrK0_0(.din(w_dff_B_pVj1v5wW0_0),.dout(w_dff_B_YYdSncrK0_0),.clk(gclk));
	jdff dff_B_7ckjdnBU4_0(.din(w_dff_B_YYdSncrK0_0),.dout(w_dff_B_7ckjdnBU4_0),.clk(gclk));
	jdff dff_B_Gwk3KFCt9_0(.din(w_dff_B_7ckjdnBU4_0),.dout(w_dff_B_Gwk3KFCt9_0),.clk(gclk));
	jdff dff_B_p1sY2Bkz6_0(.din(w_dff_B_Gwk3KFCt9_0),.dout(w_dff_B_p1sY2Bkz6_0),.clk(gclk));
	jdff dff_B_AEdSkG510_0(.din(w_dff_B_p1sY2Bkz6_0),.dout(w_dff_B_AEdSkG510_0),.clk(gclk));
	jdff dff_B_2ozSsQQ30_0(.din(w_dff_B_AEdSkG510_0),.dout(w_dff_B_2ozSsQQ30_0),.clk(gclk));
	jdff dff_B_TbPXMdHi8_0(.din(n1620),.dout(w_dff_B_TbPXMdHi8_0),.clk(gclk));
	jdff dff_B_wYeNHq3I4_2(.din(G64),.dout(w_dff_B_wYeNHq3I4_2),.clk(gclk));
	jdff dff_B_goR4it6E5_2(.din(G14),.dout(w_dff_B_goR4it6E5_2),.clk(gclk));
	jdff dff_B_Vi4narfa5_2(.din(w_dff_B_goR4it6E5_2),.dout(w_dff_B_Vi4narfa5_2),.clk(gclk));
	jdff dff_A_4D4LeZGo5_1(.dout(w_n843_1[1]),.din(w_dff_A_4D4LeZGo5_1),.clk(gclk));
	jdff dff_A_zdEm43ho5_1(.dout(w_dff_A_4D4LeZGo5_1),.din(w_dff_A_zdEm43ho5_1),.clk(gclk));
	jdff dff_A_aOjiNL5O2_1(.dout(w_dff_A_zdEm43ho5_1),.din(w_dff_A_aOjiNL5O2_1),.clk(gclk));
	jdff dff_A_y6ed07EG4_1(.dout(w_dff_A_aOjiNL5O2_1),.din(w_dff_A_y6ed07EG4_1),.clk(gclk));
	jdff dff_A_gaCAXaqN9_1(.dout(w_dff_A_y6ed07EG4_1),.din(w_dff_A_gaCAXaqN9_1),.clk(gclk));
	jdff dff_A_fCefUJbV9_1(.dout(w_dff_A_gaCAXaqN9_1),.din(w_dff_A_fCefUJbV9_1),.clk(gclk));
	jdff dff_A_i6yV8PVe8_1(.dout(w_dff_A_fCefUJbV9_1),.din(w_dff_A_i6yV8PVe8_1),.clk(gclk));
	jdff dff_A_iYlu67LX7_2(.dout(w_n843_1[2]),.din(w_dff_A_iYlu67LX7_2),.clk(gclk));
	jdff dff_A_BalXCdcn6_2(.dout(w_dff_A_iYlu67LX7_2),.din(w_dff_A_BalXCdcn6_2),.clk(gclk));
	jdff dff_A_Gxfq656C7_2(.dout(w_dff_A_BalXCdcn6_2),.din(w_dff_A_Gxfq656C7_2),.clk(gclk));
	jdff dff_A_CoexmRvB7_2(.dout(w_dff_A_Gxfq656C7_2),.din(w_dff_A_CoexmRvB7_2),.clk(gclk));
	jdff dff_A_zJTbukgA4_2(.dout(w_dff_A_CoexmRvB7_2),.din(w_dff_A_zJTbukgA4_2),.clk(gclk));
	jdff dff_A_8m2i4gXb4_2(.dout(w_dff_A_zJTbukgA4_2),.din(w_dff_A_8m2i4gXb4_2),.clk(gclk));
	jdff dff_A_4joDZmYv9_1(.dout(w_n843_0[1]),.din(w_dff_A_4joDZmYv9_1),.clk(gclk));
	jdff dff_A_HnYLLHG05_1(.dout(w_dff_A_4joDZmYv9_1),.din(w_dff_A_HnYLLHG05_1),.clk(gclk));
	jdff dff_A_7Qp7UjoB4_1(.dout(w_dff_A_HnYLLHG05_1),.din(w_dff_A_7Qp7UjoB4_1),.clk(gclk));
	jdff dff_A_bramFFDL0_1(.dout(w_dff_A_7Qp7UjoB4_1),.din(w_dff_A_bramFFDL0_1),.clk(gclk));
	jdff dff_A_EWrfPdBv2_1(.dout(w_dff_A_bramFFDL0_1),.din(w_dff_A_EWrfPdBv2_1),.clk(gclk));
	jdff dff_A_pPhhY0IA6_2(.dout(w_n843_0[2]),.din(w_dff_A_pPhhY0IA6_2),.clk(gclk));
	jdff dff_B_IiAysqFu4_3(.din(n843),.dout(w_dff_B_IiAysqFu4_3),.clk(gclk));
	jdff dff_B_PYX2lF964_3(.din(w_dff_B_IiAysqFu4_3),.dout(w_dff_B_PYX2lF964_3),.clk(gclk));
	jdff dff_B_p5nMLCf24_3(.din(w_dff_B_PYX2lF964_3),.dout(w_dff_B_p5nMLCf24_3),.clk(gclk));
	jdff dff_B_otVDLEHT6_3(.din(w_dff_B_p5nMLCf24_3),.dout(w_dff_B_otVDLEHT6_3),.clk(gclk));
	jdff dff_A_7LYzfzSD1_1(.dout(w_n840_1[1]),.din(w_dff_A_7LYzfzSD1_1),.clk(gclk));
	jdff dff_A_3lQP8ya17_1(.dout(w_dff_A_7LYzfzSD1_1),.din(w_dff_A_3lQP8ya17_1),.clk(gclk));
	jdff dff_A_3kuZopJo7_1(.dout(w_dff_A_3lQP8ya17_1),.din(w_dff_A_3kuZopJo7_1),.clk(gclk));
	jdff dff_A_b5vc8FTZ1_1(.dout(w_dff_A_3kuZopJo7_1),.din(w_dff_A_b5vc8FTZ1_1),.clk(gclk));
	jdff dff_A_6fhnPVYK1_1(.dout(w_dff_A_b5vc8FTZ1_1),.din(w_dff_A_6fhnPVYK1_1),.clk(gclk));
	jdff dff_A_OdWhSluN0_1(.dout(w_dff_A_6fhnPVYK1_1),.din(w_dff_A_OdWhSluN0_1),.clk(gclk));
	jdff dff_A_HBrApsK97_1(.dout(w_dff_A_OdWhSluN0_1),.din(w_dff_A_HBrApsK97_1),.clk(gclk));
	jdff dff_A_m2wipF8h2_1(.dout(w_dff_A_HBrApsK97_1),.din(w_dff_A_m2wipF8h2_1),.clk(gclk));
	jdff dff_A_byVzplzN1_1(.dout(w_dff_A_m2wipF8h2_1),.din(w_dff_A_byVzplzN1_1),.clk(gclk));
	jdff dff_A_OAmdyT2Q3_1(.dout(w_dff_A_byVzplzN1_1),.din(w_dff_A_OAmdyT2Q3_1),.clk(gclk));
	jdff dff_A_V1sULonp0_2(.dout(w_n840_1[2]),.din(w_dff_A_V1sULonp0_2),.clk(gclk));
	jdff dff_A_LDDCOmTK7_2(.dout(w_dff_A_V1sULonp0_2),.din(w_dff_A_LDDCOmTK7_2),.clk(gclk));
	jdff dff_A_STwPZpN01_2(.dout(w_dff_A_LDDCOmTK7_2),.din(w_dff_A_STwPZpN01_2),.clk(gclk));
	jdff dff_A_w7rRNa1K2_2(.dout(w_dff_A_STwPZpN01_2),.din(w_dff_A_w7rRNa1K2_2),.clk(gclk));
	jdff dff_A_k8BHUIRL0_2(.dout(w_dff_A_w7rRNa1K2_2),.din(w_dff_A_k8BHUIRL0_2),.clk(gclk));
	jdff dff_A_6l0cAnec7_2(.dout(w_dff_A_k8BHUIRL0_2),.din(w_dff_A_6l0cAnec7_2),.clk(gclk));
	jdff dff_A_2csyo9hG7_2(.dout(w_dff_A_6l0cAnec7_2),.din(w_dff_A_2csyo9hG7_2),.clk(gclk));
	jdff dff_A_K2lEsZEX3_1(.dout(w_n840_0[1]),.din(w_dff_A_K2lEsZEX3_1),.clk(gclk));
	jdff dff_A_rOGRVMiY5_1(.dout(w_dff_A_K2lEsZEX3_1),.din(w_dff_A_rOGRVMiY5_1),.clk(gclk));
	jdff dff_A_YLqsyOWq0_1(.dout(w_dff_A_rOGRVMiY5_1),.din(w_dff_A_YLqsyOWq0_1),.clk(gclk));
	jdff dff_A_qr0LnxOY1_1(.dout(w_dff_A_YLqsyOWq0_1),.din(w_dff_A_qr0LnxOY1_1),.clk(gclk));
	jdff dff_A_uFGO2QA43_1(.dout(w_dff_A_qr0LnxOY1_1),.din(w_dff_A_uFGO2QA43_1),.clk(gclk));
	jdff dff_A_sCQiNn1o4_2(.dout(w_n840_0[2]),.din(w_dff_A_sCQiNn1o4_2),.clk(gclk));
	jdff dff_A_KFFPcOaf4_2(.dout(w_dff_A_sCQiNn1o4_2),.din(w_dff_A_KFFPcOaf4_2),.clk(gclk));
	jdff dff_A_xGvSj7hy3_2(.dout(w_dff_A_KFFPcOaf4_2),.din(w_dff_A_xGvSj7hy3_2),.clk(gclk));
	jdff dff_A_225P8l8c2_2(.dout(w_dff_A_xGvSj7hy3_2),.din(w_dff_A_225P8l8c2_2),.clk(gclk));
	jdff dff_B_tBgkUl0I6_3(.din(n840),.dout(w_dff_B_tBgkUl0I6_3),.clk(gclk));
	jdff dff_B_hr7FeO4t4_3(.din(w_dff_B_tBgkUl0I6_3),.dout(w_dff_B_hr7FeO4t4_3),.clk(gclk));
	jdff dff_B_VSUl2bQH4_3(.din(w_dff_B_hr7FeO4t4_3),.dout(w_dff_B_VSUl2bQH4_3),.clk(gclk));
	jdff dff_B_SwqRqUfg5_3(.din(w_dff_B_VSUl2bQH4_3),.dout(w_dff_B_SwqRqUfg5_3),.clk(gclk));
	jdff dff_B_eS2njwbW0_3(.din(w_dff_B_SwqRqUfg5_3),.dout(w_dff_B_eS2njwbW0_3),.clk(gclk));
	jdff dff_B_47vXz1si6_3(.din(w_dff_B_eS2njwbW0_3),.dout(w_dff_B_47vXz1si6_3),.clk(gclk));
	jdff dff_A_oD4ZL31J1_1(.dout(w_G4090_0[1]),.din(w_dff_A_oD4ZL31J1_1),.clk(gclk));
	jdff dff_A_CfNDWJtS0_2(.dout(w_G4089_0[2]),.din(w_dff_A_CfNDWJtS0_2),.clk(gclk));
	jdff dff_B_sNBr3ATY3_0(.din(n1638),.dout(w_dff_B_sNBr3ATY3_0),.clk(gclk));
	jdff dff_B_eBSRsZqY1_0(.din(w_dff_B_sNBr3ATY3_0),.dout(w_dff_B_eBSRsZqY1_0),.clk(gclk));
	jdff dff_B_okrWZa0i1_0(.din(n1637),.dout(w_dff_B_okrWZa0i1_0),.clk(gclk));
	jdff dff_B_OS5yAMzL9_0(.din(w_dff_B_okrWZa0i1_0),.dout(w_dff_B_OS5yAMzL9_0),.clk(gclk));
	jdff dff_B_uzvCX6Ce6_0(.din(w_dff_B_OS5yAMzL9_0),.dout(w_dff_B_uzvCX6Ce6_0),.clk(gclk));
	jdff dff_B_I8A9TEcj2_0(.din(w_dff_B_uzvCX6Ce6_0),.dout(w_dff_B_I8A9TEcj2_0),.clk(gclk));
	jdff dff_B_mcHwpzJl9_0(.din(w_dff_B_I8A9TEcj2_0),.dout(w_dff_B_mcHwpzJl9_0),.clk(gclk));
	jdff dff_B_mawCYAhC3_0(.din(w_dff_B_mcHwpzJl9_0),.dout(w_dff_B_mawCYAhC3_0),.clk(gclk));
	jdff dff_B_lzhpR4z89_0(.din(w_dff_B_mawCYAhC3_0),.dout(w_dff_B_lzhpR4z89_0),.clk(gclk));
	jdff dff_B_Y33MBaP45_0(.din(w_dff_B_lzhpR4z89_0),.dout(w_dff_B_Y33MBaP45_0),.clk(gclk));
	jdff dff_B_uGuT4d9i7_0(.din(w_dff_B_Y33MBaP45_0),.dout(w_dff_B_uGuT4d9i7_0),.clk(gclk));
	jdff dff_B_7OXd0QYL8_0(.din(w_dff_B_uGuT4d9i7_0),.dout(w_dff_B_7OXd0QYL8_0),.clk(gclk));
	jdff dff_B_iLAdrS1b7_1(.din(n1633),.dout(w_dff_B_iLAdrS1b7_1),.clk(gclk));
	jdff dff_B_BvUgjQVi0_1(.din(n1627),.dout(w_dff_B_BvUgjQVi0_1),.clk(gclk));
	jdff dff_B_hZ2QxyWZ5_1(.din(w_dff_B_BvUgjQVi0_1),.dout(w_dff_B_hZ2QxyWZ5_1),.clk(gclk));
	jdff dff_B_maOVicp01_1(.din(w_dff_B_hZ2QxyWZ5_1),.dout(w_dff_B_maOVicp01_1),.clk(gclk));
	jdff dff_B_ABCI4f7I3_1(.din(w_dff_B_maOVicp01_1),.dout(w_dff_B_ABCI4f7I3_1),.clk(gclk));
	jdff dff_B_HWHU7TwK8_1(.din(w_dff_B_ABCI4f7I3_1),.dout(w_dff_B_HWHU7TwK8_1),.clk(gclk));
	jdff dff_B_f0LutFs85_1(.din(w_dff_B_HWHU7TwK8_1),.dout(w_dff_B_f0LutFs85_1),.clk(gclk));
	jdff dff_B_o2ZrxLxI2_1(.din(w_dff_B_f0LutFs85_1),.dout(w_dff_B_o2ZrxLxI2_1),.clk(gclk));
	jdff dff_B_GfeBdrXb4_1(.din(w_dff_B_o2ZrxLxI2_1),.dout(w_dff_B_GfeBdrXb4_1),.clk(gclk));
	jdff dff_B_e89mvSKZ7_1(.din(w_dff_B_GfeBdrXb4_1),.dout(w_dff_B_e89mvSKZ7_1),.clk(gclk));
	jdff dff_B_fWsQXXrF4_1(.din(w_dff_B_e89mvSKZ7_1),.dout(w_dff_B_fWsQXXrF4_1),.clk(gclk));
	jdff dff_B_VaxEOFz65_1(.din(w_dff_B_fWsQXXrF4_1),.dout(w_dff_B_VaxEOFz65_1),.clk(gclk));
	jdff dff_A_2u9BSIhp7_0(.dout(w_n988_1[0]),.din(w_dff_A_2u9BSIhp7_0),.clk(gclk));
	jdff dff_A_DdmFGqHt5_0(.dout(w_dff_A_2u9BSIhp7_0),.din(w_dff_A_DdmFGqHt5_0),.clk(gclk));
	jdff dff_A_dJaYxjqo6_0(.dout(w_dff_A_DdmFGqHt5_0),.din(w_dff_A_dJaYxjqo6_0),.clk(gclk));
	jdff dff_A_pWkXD5lq7_0(.dout(w_dff_A_dJaYxjqo6_0),.din(w_dff_A_pWkXD5lq7_0),.clk(gclk));
	jdff dff_A_YGRwvE6t0_2(.dout(w_n988_1[2]),.din(w_dff_A_YGRwvE6t0_2),.clk(gclk));
	jdff dff_A_cw52e6LO7_2(.dout(w_dff_A_YGRwvE6t0_2),.din(w_dff_A_cw52e6LO7_2),.clk(gclk));
	jdff dff_A_pBaM6wMA7_2(.dout(w_dff_A_cw52e6LO7_2),.din(w_dff_A_pBaM6wMA7_2),.clk(gclk));
	jdff dff_A_z0Jg1tsc0_2(.dout(w_dff_A_pBaM6wMA7_2),.din(w_dff_A_z0Jg1tsc0_2),.clk(gclk));
	jdff dff_A_TjEuZVEy3_2(.dout(w_dff_A_z0Jg1tsc0_2),.din(w_dff_A_TjEuZVEy3_2),.clk(gclk));
	jdff dff_A_zWFcKXYn6_2(.dout(w_dff_A_TjEuZVEy3_2),.din(w_dff_A_zWFcKXYn6_2),.clk(gclk));
	jdff dff_A_82wkT1EN3_2(.dout(w_dff_A_zWFcKXYn6_2),.din(w_dff_A_82wkT1EN3_2),.clk(gclk));
	jdff dff_A_QsdVDy8B5_2(.dout(w_dff_A_82wkT1EN3_2),.din(w_dff_A_QsdVDy8B5_2),.clk(gclk));
	jdff dff_A_m3SICdOU5_2(.dout(w_dff_A_QsdVDy8B5_2),.din(w_dff_A_m3SICdOU5_2),.clk(gclk));
	jdff dff_A_7RiZXL4r0_1(.dout(w_n988_0[1]),.din(w_dff_A_7RiZXL4r0_1),.clk(gclk));
	jdff dff_A_ZItrffyO1_1(.dout(w_dff_A_7RiZXL4r0_1),.din(w_dff_A_ZItrffyO1_1),.clk(gclk));
	jdff dff_A_Cm1cGdOU7_1(.dout(w_dff_A_ZItrffyO1_1),.din(w_dff_A_Cm1cGdOU7_1),.clk(gclk));
	jdff dff_A_5o8TgSOR1_1(.dout(w_dff_A_Cm1cGdOU7_1),.din(w_dff_A_5o8TgSOR1_1),.clk(gclk));
	jdff dff_A_PknUmGKH2_1(.dout(w_dff_A_5o8TgSOR1_1),.din(w_dff_A_PknUmGKH2_1),.clk(gclk));
	jdff dff_A_Pl6plcCR9_1(.dout(w_dff_A_PknUmGKH2_1),.din(w_dff_A_Pl6plcCR9_1),.clk(gclk));
	jdff dff_A_Fo2TcyFP3_1(.dout(w_dff_A_Pl6plcCR9_1),.din(w_dff_A_Fo2TcyFP3_1),.clk(gclk));
	jdff dff_A_eKpMuOXE5_1(.dout(w_dff_A_Fo2TcyFP3_1),.din(w_dff_A_eKpMuOXE5_1),.clk(gclk));
	jdff dff_A_oWhN8KOx3_1(.dout(w_dff_A_eKpMuOXE5_1),.din(w_dff_A_oWhN8KOx3_1),.clk(gclk));
	jdff dff_A_052EMNkd0_2(.dout(w_n988_0[2]),.din(w_dff_A_052EMNkd0_2),.clk(gclk));
	jdff dff_A_fknCMaa94_2(.dout(w_dff_A_052EMNkd0_2),.din(w_dff_A_fknCMaa94_2),.clk(gclk));
	jdff dff_A_4rJKj9vY1_2(.dout(w_dff_A_fknCMaa94_2),.din(w_dff_A_4rJKj9vY1_2),.clk(gclk));
	jdff dff_A_1KKrVCTr9_2(.dout(w_dff_A_4rJKj9vY1_2),.din(w_dff_A_1KKrVCTr9_2),.clk(gclk));
	jdff dff_A_rMbDKlHt8_2(.dout(w_dff_A_1KKrVCTr9_2),.din(w_dff_A_rMbDKlHt8_2),.clk(gclk));
	jdff dff_B_0KlNMVYb2_1(.din(n1625),.dout(w_dff_B_0KlNMVYb2_1),.clk(gclk));
	jdff dff_B_aojd7tuv2_1(.din(w_dff_B_0KlNMVYb2_1),.dout(w_dff_B_aojd7tuv2_1),.clk(gclk));
	jdff dff_B_trfTZQBd9_1(.din(w_dff_B_aojd7tuv2_1),.dout(w_dff_B_trfTZQBd9_1),.clk(gclk));
	jdff dff_B_wxInqJFz6_1(.din(w_dff_B_trfTZQBd9_1),.dout(w_dff_B_wxInqJFz6_1),.clk(gclk));
	jdff dff_B_00lEdccQ8_1(.din(w_dff_B_wxInqJFz6_1),.dout(w_dff_B_00lEdccQ8_1),.clk(gclk));
	jdff dff_B_tlznQ9Nw9_1(.din(w_dff_B_00lEdccQ8_1),.dout(w_dff_B_tlznQ9Nw9_1),.clk(gclk));
	jdff dff_B_o4aJ5EZ73_1(.din(w_dff_B_tlznQ9Nw9_1),.dout(w_dff_B_o4aJ5EZ73_1),.clk(gclk));
	jdff dff_B_72JzGlTT8_1(.din(w_dff_B_o4aJ5EZ73_1),.dout(w_dff_B_72JzGlTT8_1),.clk(gclk));
	jdff dff_B_QeCboIuJ4_1(.din(w_dff_B_72JzGlTT8_1),.dout(w_dff_B_QeCboIuJ4_1),.clk(gclk));
	jdff dff_B_uKF5PvQs8_1(.din(w_dff_B_QeCboIuJ4_1),.dout(w_dff_B_uKF5PvQs8_1),.clk(gclk));
	jdff dff_B_Ft5VBjlW8_1(.din(w_dff_B_uKF5PvQs8_1),.dout(w_dff_B_Ft5VBjlW8_1),.clk(gclk));
	jdff dff_B_VBe4Pi9L6_1(.din(w_dff_B_Ft5VBjlW8_1),.dout(w_dff_B_VBe4Pi9L6_1),.clk(gclk));
	jdff dff_B_41iV7Vct0_1(.din(w_dff_B_VBe4Pi9L6_1),.dout(w_dff_B_41iV7Vct0_1),.clk(gclk));
	jdff dff_B_jecj7M9W1_1(.din(w_dff_B_41iV7Vct0_1),.dout(w_dff_B_jecj7M9W1_1),.clk(gclk));
	jdff dff_A_adHWuCeE4_0(.dout(w_n985_1[0]),.din(w_dff_A_adHWuCeE4_0),.clk(gclk));
	jdff dff_A_leLUn6aC2_0(.dout(w_dff_A_adHWuCeE4_0),.din(w_dff_A_leLUn6aC2_0),.clk(gclk));
	jdff dff_A_NMvM3QNc1_0(.dout(w_dff_A_leLUn6aC2_0),.din(w_dff_A_NMvM3QNc1_0),.clk(gclk));
	jdff dff_A_sHkldfAJ2_0(.dout(w_dff_A_NMvM3QNc1_0),.din(w_dff_A_sHkldfAJ2_0),.clk(gclk));
	jdff dff_A_kN3KSB2c5_0(.dout(w_dff_A_sHkldfAJ2_0),.din(w_dff_A_kN3KSB2c5_0),.clk(gclk));
	jdff dff_A_YSPdOOlB5_0(.dout(w_dff_A_kN3KSB2c5_0),.din(w_dff_A_YSPdOOlB5_0),.clk(gclk));
	jdff dff_A_oYXk3jmS2_2(.dout(w_n985_1[2]),.din(w_dff_A_oYXk3jmS2_2),.clk(gclk));
	jdff dff_A_OwsF0eaN9_2(.dout(w_dff_A_oYXk3jmS2_2),.din(w_dff_A_OwsF0eaN9_2),.clk(gclk));
	jdff dff_A_hNECWQIm3_2(.dout(w_dff_A_OwsF0eaN9_2),.din(w_dff_A_hNECWQIm3_2),.clk(gclk));
	jdff dff_A_GG3wOGg22_2(.dout(w_dff_A_hNECWQIm3_2),.din(w_dff_A_GG3wOGg22_2),.clk(gclk));
	jdff dff_A_dszaMtZc7_2(.dout(w_dff_A_GG3wOGg22_2),.din(w_dff_A_dszaMtZc7_2),.clk(gclk));
	jdff dff_A_NjS41Zuc0_2(.dout(w_dff_A_dszaMtZc7_2),.din(w_dff_A_NjS41Zuc0_2),.clk(gclk));
	jdff dff_A_BOsRK9m87_2(.dout(w_dff_A_NjS41Zuc0_2),.din(w_dff_A_BOsRK9m87_2),.clk(gclk));
	jdff dff_A_UclOCWtG6_2(.dout(w_dff_A_BOsRK9m87_2),.din(w_dff_A_UclOCWtG6_2),.clk(gclk));
	jdff dff_A_qiAxdV336_2(.dout(w_dff_A_UclOCWtG6_2),.din(w_dff_A_qiAxdV336_2),.clk(gclk));
	jdff dff_A_pVUEcUwf2_2(.dout(w_dff_A_qiAxdV336_2),.din(w_dff_A_pVUEcUwf2_2),.clk(gclk));
	jdff dff_A_YrOEY4DL7_2(.dout(w_dff_A_pVUEcUwf2_2),.din(w_dff_A_YrOEY4DL7_2),.clk(gclk));
	jdff dff_A_U60A0pOU2_1(.dout(w_n985_0[1]),.din(w_dff_A_U60A0pOU2_1),.clk(gclk));
	jdff dff_A_ePAM0KZN2_1(.dout(w_dff_A_U60A0pOU2_1),.din(w_dff_A_ePAM0KZN2_1),.clk(gclk));
	jdff dff_A_TbNVKSXl8_1(.dout(w_dff_A_ePAM0KZN2_1),.din(w_dff_A_TbNVKSXl8_1),.clk(gclk));
	jdff dff_A_czh8Ldbd9_1(.dout(w_dff_A_TbNVKSXl8_1),.din(w_dff_A_czh8Ldbd9_1),.clk(gclk));
	jdff dff_A_giM0K1t94_1(.dout(w_dff_A_czh8Ldbd9_1),.din(w_dff_A_giM0K1t94_1),.clk(gclk));
	jdff dff_A_RFGR9Min8_1(.dout(w_dff_A_giM0K1t94_1),.din(w_dff_A_RFGR9Min8_1),.clk(gclk));
	jdff dff_A_uQhfEnFK9_1(.dout(w_dff_A_RFGR9Min8_1),.din(w_dff_A_uQhfEnFK9_1),.clk(gclk));
	jdff dff_A_LPO3o2Em8_1(.dout(w_dff_A_uQhfEnFK9_1),.din(w_dff_A_LPO3o2Em8_1),.clk(gclk));
	jdff dff_A_4Kcgv1au1_1(.dout(w_dff_A_LPO3o2Em8_1),.din(w_dff_A_4Kcgv1au1_1),.clk(gclk));
	jdff dff_A_FcxtTaGY8_1(.dout(w_dff_A_4Kcgv1au1_1),.din(w_dff_A_FcxtTaGY8_1),.clk(gclk));
	jdff dff_A_PWutiuU86_1(.dout(w_dff_A_FcxtTaGY8_1),.din(w_dff_A_PWutiuU86_1),.clk(gclk));
	jdff dff_A_CHXxb75R2_2(.dout(w_n985_0[2]),.din(w_dff_A_CHXxb75R2_2),.clk(gclk));
	jdff dff_A_lhKde5el0_2(.dout(w_dff_A_CHXxb75R2_2),.din(w_dff_A_lhKde5el0_2),.clk(gclk));
	jdff dff_A_fqSfXrmM9_2(.dout(w_dff_A_lhKde5el0_2),.din(w_dff_A_fqSfXrmM9_2),.clk(gclk));
	jdff dff_A_edZWuZD80_2(.dout(w_dff_A_fqSfXrmM9_2),.din(w_dff_A_edZWuZD80_2),.clk(gclk));
	jdff dff_A_0fzo63Xs3_2(.dout(w_dff_A_edZWuZD80_2),.din(w_dff_A_0fzo63Xs3_2),.clk(gclk));
	jdff dff_A_eDqHULD71_2(.dout(w_dff_A_0fzo63Xs3_2),.din(w_dff_A_eDqHULD71_2),.clk(gclk));
	jdff dff_A_zlirVD4t1_2(.dout(w_dff_A_eDqHULD71_2),.din(w_dff_A_zlirVD4t1_2),.clk(gclk));
	jdff dff_A_hyaNnRaW1_2(.dout(w_dff_A_zlirVD4t1_2),.din(w_dff_A_hyaNnRaW1_2),.clk(gclk));
	jdff dff_A_FKlsEDyB0_2(.dout(w_dff_A_hyaNnRaW1_2),.din(w_dff_A_FKlsEDyB0_2),.clk(gclk));
	jdff dff_A_AL1UiXwR6_2(.dout(w_dff_A_FKlsEDyB0_2),.din(w_dff_A_AL1UiXwR6_2),.clk(gclk));
	jdff dff_A_qzXADXbr4_1(.dout(w_G1690_0[1]),.din(w_dff_A_qzXADXbr4_1),.clk(gclk));
	jdff dff_A_URGcx6v34_2(.dout(w_G1689_0[2]),.din(w_dff_A_URGcx6v34_2),.clk(gclk));
	jdff dff_B_fqWouHea6_0(.din(n1650),.dout(w_dff_B_fqWouHea6_0),.clk(gclk));
	jdff dff_B_vBojNKb56_0(.din(w_dff_B_fqWouHea6_0),.dout(w_dff_B_vBojNKb56_0),.clk(gclk));
	jdff dff_B_WM1tHPGa7_0(.din(n1649),.dout(w_dff_B_WM1tHPGa7_0),.clk(gclk));
	jdff dff_B_FaABieyl2_0(.din(w_dff_B_WM1tHPGa7_0),.dout(w_dff_B_FaABieyl2_0),.clk(gclk));
	jdff dff_B_u7LXajn30_0(.din(w_dff_B_FaABieyl2_0),.dout(w_dff_B_u7LXajn30_0),.clk(gclk));
	jdff dff_B_bbJzPE2w9_0(.din(w_dff_B_u7LXajn30_0),.dout(w_dff_B_bbJzPE2w9_0),.clk(gclk));
	jdff dff_B_UzxBI4C67_0(.din(w_dff_B_bbJzPE2w9_0),.dout(w_dff_B_UzxBI4C67_0),.clk(gclk));
	jdff dff_B_agNzetIO5_0(.din(w_dff_B_UzxBI4C67_0),.dout(w_dff_B_agNzetIO5_0),.clk(gclk));
	jdff dff_B_Tnf8RmDr2_0(.din(w_dff_B_agNzetIO5_0),.dout(w_dff_B_Tnf8RmDr2_0),.clk(gclk));
	jdff dff_B_f8Xw0BPk7_0(.din(w_dff_B_Tnf8RmDr2_0),.dout(w_dff_B_f8Xw0BPk7_0),.clk(gclk));
	jdff dff_B_7l4zDyOq7_0(.din(w_dff_B_f8Xw0BPk7_0),.dout(w_dff_B_7l4zDyOq7_0),.clk(gclk));
	jdff dff_B_c0kWm8PA4_0(.din(w_dff_B_7l4zDyOq7_0),.dout(w_dff_B_c0kWm8PA4_0),.clk(gclk));
	jdff dff_B_j1RoE3pl4_1(.din(n1646),.dout(w_dff_B_j1RoE3pl4_1),.clk(gclk));
	jdff dff_B_OYLwbySd3_2(.din(n1634),.dout(w_dff_B_OYLwbySd3_2),.clk(gclk));
	jdff dff_B_IijeVrdw9_2(.din(w_dff_B_OYLwbySd3_2),.dout(w_dff_B_IijeVrdw9_2),.clk(gclk));
	jdff dff_B_yuVHT2KF9_2(.din(n1631),.dout(w_dff_B_yuVHT2KF9_2),.clk(gclk));
	jdff dff_B_mfru56XC0_1(.din(n1643),.dout(w_dff_B_mfru56XC0_1),.clk(gclk));
	jdff dff_B_rtdV5vk31_1(.din(w_dff_B_mfru56XC0_1),.dout(w_dff_B_rtdV5vk31_1),.clk(gclk));
	jdff dff_B_5UTeVcWU8_1(.din(w_dff_B_rtdV5vk31_1),.dout(w_dff_B_5UTeVcWU8_1),.clk(gclk));
	jdff dff_B_jHTfRm792_1(.din(w_dff_B_5UTeVcWU8_1),.dout(w_dff_B_jHTfRm792_1),.clk(gclk));
	jdff dff_B_sVg7GnU89_1(.din(w_dff_B_jHTfRm792_1),.dout(w_dff_B_sVg7GnU89_1),.clk(gclk));
	jdff dff_B_fOBGt4Bz8_1(.din(w_dff_B_sVg7GnU89_1),.dout(w_dff_B_fOBGt4Bz8_1),.clk(gclk));
	jdff dff_B_ORhifE5o6_1(.din(w_dff_B_fOBGt4Bz8_1),.dout(w_dff_B_ORhifE5o6_1),.clk(gclk));
	jdff dff_B_0Aa7H1r13_1(.din(w_dff_B_ORhifE5o6_1),.dout(w_dff_B_0Aa7H1r13_1),.clk(gclk));
	jdff dff_B_Z5BzX2Ir7_1(.din(w_dff_B_0Aa7H1r13_1),.dout(w_dff_B_Z5BzX2Ir7_1),.clk(gclk));
	jdff dff_B_So66SSTL9_1(.din(w_dff_B_Z5BzX2Ir7_1),.dout(w_dff_B_So66SSTL9_1),.clk(gclk));
	jdff dff_B_fOlDPyLf2_1(.din(w_dff_B_So66SSTL9_1),.dout(w_dff_B_fOlDPyLf2_1),.clk(gclk));
	jdff dff_B_jFTjUPkQ1_0(.din(n1628),.dout(w_dff_B_jFTjUPkQ1_0),.clk(gclk));
	jdff dff_B_t7aTVRiG7_0(.din(w_dff_B_jFTjUPkQ1_0),.dout(w_dff_B_t7aTVRiG7_0),.clk(gclk));
	jdff dff_B_PUgWhadD3_0(.din(w_dff_B_t7aTVRiG7_0),.dout(w_dff_B_PUgWhadD3_0),.clk(gclk));
	jdff dff_B_Qu0lJpbU3_0(.din(w_dff_B_PUgWhadD3_0),.dout(w_dff_B_Qu0lJpbU3_0),.clk(gclk));
	jdff dff_B_xGlEeWWG5_0(.din(w_dff_B_Qu0lJpbU3_0),.dout(w_dff_B_xGlEeWWG5_0),.clk(gclk));
	jdff dff_B_ZnOInu1j7_0(.din(w_dff_B_xGlEeWWG5_0),.dout(w_dff_B_ZnOInu1j7_0),.clk(gclk));
	jdff dff_B_5lYKl7oa9_0(.din(w_dff_B_ZnOInu1j7_0),.dout(w_dff_B_5lYKl7oa9_0),.clk(gclk));
	jdff dff_B_hpEDnRyu5_0(.din(w_dff_B_5lYKl7oa9_0),.dout(w_dff_B_hpEDnRyu5_0),.clk(gclk));
	jdff dff_B_vcfHocrm7_0(.din(w_dff_B_hpEDnRyu5_0),.dout(w_dff_B_vcfHocrm7_0),.clk(gclk));
	jdff dff_B_PpfcEzsH6_0(.din(w_dff_B_vcfHocrm7_0),.dout(w_dff_B_PpfcEzsH6_0),.clk(gclk));
	jdff dff_B_YbeTSPWj2_0(.din(w_dff_B_PpfcEzsH6_0),.dout(w_dff_B_YbeTSPWj2_0),.clk(gclk));
	jdff dff_A_rCYBnmEg1_1(.dout(w_n1609_0[1]),.din(w_dff_A_rCYBnmEg1_1),.clk(gclk));
	jdff dff_A_lP26CVsM0_1(.dout(w_dff_A_rCYBnmEg1_1),.din(w_dff_A_lP26CVsM0_1),.clk(gclk));
	jdff dff_A_AhLdy75s1_1(.dout(w_dff_A_lP26CVsM0_1),.din(w_dff_A_AhLdy75s1_1),.clk(gclk));
	jdff dff_A_MTiQNhBQ7_1(.dout(w_dff_A_AhLdy75s1_1),.din(w_dff_A_MTiQNhBQ7_1),.clk(gclk));
	jdff dff_A_Pmj0bQon5_1(.dout(w_dff_A_MTiQNhBQ7_1),.din(w_dff_A_Pmj0bQon5_1),.clk(gclk));
	jdff dff_A_VDZLaOd94_1(.dout(w_dff_A_Pmj0bQon5_1),.din(w_dff_A_VDZLaOd94_1),.clk(gclk));
	jdff dff_A_2ABTlY0k5_1(.dout(w_dff_A_VDZLaOd94_1),.din(w_dff_A_2ABTlY0k5_1),.clk(gclk));
	jdff dff_A_SPpikRhb5_1(.dout(w_dff_A_2ABTlY0k5_1),.din(w_dff_A_SPpikRhb5_1),.clk(gclk));
	jdff dff_A_FHEEx5ER8_1(.dout(w_dff_A_SPpikRhb5_1),.din(w_dff_A_FHEEx5ER8_1),.clk(gclk));
	jdff dff_A_t8CA8yz12_1(.dout(w_dff_A_FHEEx5ER8_1),.din(w_dff_A_t8CA8yz12_1),.clk(gclk));
	jdff dff_A_6nFD0VXw5_1(.dout(w_dff_A_t8CA8yz12_1),.din(w_dff_A_6nFD0VXw5_1),.clk(gclk));
	jdff dff_A_DtNh0NaG6_1(.dout(w_dff_A_6nFD0VXw5_1),.din(w_dff_A_DtNh0NaG6_1),.clk(gclk));
	jdff dff_B_IaVweoaI3_1(.din(n1392),.dout(w_dff_B_IaVweoaI3_1),.clk(gclk));
	jdff dff_B_h1XvESGJ0_1(.din(w_dff_B_IaVweoaI3_1),.dout(w_dff_B_h1XvESGJ0_1),.clk(gclk));
	jdff dff_B_Zd4hGI9Q4_1(.din(w_dff_B_h1XvESGJ0_1),.dout(w_dff_B_Zd4hGI9Q4_1),.clk(gclk));
	jdff dff_A_D7xd73bS1_1(.dout(w_n1447_0[1]),.din(w_dff_A_D7xd73bS1_1),.clk(gclk));
	jdff dff_B_ydJ6yyv97_1(.din(n1412),.dout(w_dff_B_ydJ6yyv97_1),.clk(gclk));
	jdff dff_B_6MrwQT9Q8_1(.din(w_dff_B_ydJ6yyv97_1),.dout(w_dff_B_6MrwQT9Q8_1),.clk(gclk));
	jdff dff_B_QzR7Lzsn5_1(.din(w_dff_B_6MrwQT9Q8_1),.dout(w_dff_B_QzR7Lzsn5_1),.clk(gclk));
	jdff dff_B_3a1Rd7XP1_1(.din(w_dff_B_QzR7Lzsn5_1),.dout(w_dff_B_3a1Rd7XP1_1),.clk(gclk));
	jdff dff_B_ulOgNjix6_1(.din(w_dff_B_3a1Rd7XP1_1),.dout(w_dff_B_ulOgNjix6_1),.clk(gclk));
	jdff dff_B_F6BENzHa7_0(.din(n1442),.dout(w_dff_B_F6BENzHa7_0),.clk(gclk));
	jdff dff_A_pKuIPQC85_1(.dout(w_n1438_0[1]),.din(w_dff_A_pKuIPQC85_1),.clk(gclk));
	jdff dff_A_OosqPwxe4_1(.dout(w_dff_A_pKuIPQC85_1),.din(w_dff_A_OosqPwxe4_1),.clk(gclk));
	jdff dff_B_d48WTmlE2_1(.din(n1428),.dout(w_dff_B_d48WTmlE2_1),.clk(gclk));
	jdff dff_B_PoG6LbAh5_1(.din(w_dff_B_d48WTmlE2_1),.dout(w_dff_B_PoG6LbAh5_1),.clk(gclk));
	jdff dff_B_kcnU5YOQ8_1(.din(w_dff_B_PoG6LbAh5_1),.dout(w_dff_B_kcnU5YOQ8_1),.clk(gclk));
	jdff dff_B_tyFSTSqR1_1(.din(w_dff_B_kcnU5YOQ8_1),.dout(w_dff_B_tyFSTSqR1_1),.clk(gclk));
	jdff dff_B_n9yeWDR19_1(.din(w_dff_B_tyFSTSqR1_1),.dout(w_dff_B_n9yeWDR19_1),.clk(gclk));
	jdff dff_B_nnw0AT4Z5_1(.din(w_dff_B_n9yeWDR19_1),.dout(w_dff_B_nnw0AT4Z5_1),.clk(gclk));
	jdff dff_B_M8LVzLZV3_1(.din(w_dff_B_nnw0AT4Z5_1),.dout(w_dff_B_M8LVzLZV3_1),.clk(gclk));
	jdff dff_A_dKjpUH6t2_0(.dout(w_n1421_0[0]),.din(w_dff_A_dKjpUH6t2_0),.clk(gclk));
	jdff dff_B_kv5PswOs4_0(.din(n1418),.dout(w_dff_B_kv5PswOs4_0),.clk(gclk));
	jdff dff_A_NH7oi9Al9_1(.dout(w_n829_0[1]),.din(w_dff_A_NH7oi9Al9_1),.clk(gclk));
	jdff dff_A_BQYkyJkX0_0(.dout(w_n614_1[0]),.din(w_dff_A_BQYkyJkX0_0),.clk(gclk));
	jdff dff_A_M91kGm5M5_2(.dout(w_n614_1[2]),.din(w_dff_A_M91kGm5M5_2),.clk(gclk));
	jdff dff_A_Hr6ZOa831_1(.dout(w_n828_0[1]),.din(w_dff_A_Hr6ZOa831_1),.clk(gclk));
	jdff dff_A_9UO06Igl5_1(.dout(w_dff_A_Hr6ZOa831_1),.din(w_dff_A_9UO06Igl5_1),.clk(gclk));
	jdff dff_A_5tZlyRKT7_1(.dout(w_dff_A_9UO06Igl5_1),.din(w_dff_A_5tZlyRKT7_1),.clk(gclk));
	jdff dff_A_IUNeA1Eq8_2(.dout(w_n828_0[2]),.din(w_dff_A_IUNeA1Eq8_2),.clk(gclk));
	jdff dff_B_uzq9ZczS6_3(.din(n828),.dout(w_dff_B_uzq9ZczS6_3),.clk(gclk));
	jdff dff_A_EFYaffDo5_0(.dout(w_n787_0[0]),.din(w_dff_A_EFYaffDo5_0),.clk(gclk));
	jdff dff_B_Zp6fleZK1_2(.din(n787),.dout(w_dff_B_Zp6fleZK1_2),.clk(gclk));
	jdff dff_B_uDLjX3Wb0_2(.din(w_dff_B_Zp6fleZK1_2),.dout(w_dff_B_uDLjX3Wb0_2),.clk(gclk));
	jdff dff_A_OPaFR7er4_1(.dout(w_n779_0[1]),.din(w_dff_A_OPaFR7er4_1),.clk(gclk));
	jdff dff_A_hzaxWGKC6_1(.dout(w_dff_A_OPaFR7er4_1),.din(w_dff_A_hzaxWGKC6_1),.clk(gclk));
	jdff dff_A_IeQOYRoV6_1(.dout(w_dff_A_hzaxWGKC6_1),.din(w_dff_A_IeQOYRoV6_1),.clk(gclk));
	jdff dff_A_94AJ8mIn3_1(.dout(w_dff_A_IeQOYRoV6_1),.din(w_dff_A_94AJ8mIn3_1),.clk(gclk));
	jdff dff_A_5khHNIqZ3_1(.dout(w_dff_A_94AJ8mIn3_1),.din(w_dff_A_5khHNIqZ3_1),.clk(gclk));
	jdff dff_B_t1yzHTb16_2(.din(n779),.dout(w_dff_B_t1yzHTb16_2),.clk(gclk));
	jdff dff_A_zdmK2Fm59_1(.dout(w_n636_1[1]),.din(w_dff_A_zdmK2Fm59_1),.clk(gclk));
	jdff dff_A_9glmY7mj1_1(.dout(w_dff_A_zdmK2Fm59_1),.din(w_dff_A_9glmY7mj1_1),.clk(gclk));
	jdff dff_A_Hf5VxlTZ1_1(.dout(w_dff_A_9glmY7mj1_1),.din(w_dff_A_Hf5VxlTZ1_1),.clk(gclk));
	jdff dff_A_Kt22aKLs3_0(.dout(w_n1411_0[0]),.din(w_dff_A_Kt22aKLs3_0),.clk(gclk));
	jdff dff_A_9KwEno5i5_0(.dout(w_dff_A_Kt22aKLs3_0),.din(w_dff_A_9KwEno5i5_0),.clk(gclk));
	jdff dff_A_RCY82oFT2_0(.dout(w_dff_A_9KwEno5i5_0),.din(w_dff_A_RCY82oFT2_0),.clk(gclk));
	jdff dff_A_rgjTPVoo8_0(.dout(w_dff_A_RCY82oFT2_0),.din(w_dff_A_rgjTPVoo8_0),.clk(gclk));
	jdff dff_A_Km3aMFaw3_0(.dout(w_dff_A_rgjTPVoo8_0),.din(w_dff_A_Km3aMFaw3_0),.clk(gclk));
	jdff dff_A_1QglDTsf6_0(.dout(w_dff_A_Km3aMFaw3_0),.din(w_dff_A_1QglDTsf6_0),.clk(gclk));
	jdff dff_B_KpRwIewu3_2(.din(n1410),.dout(w_dff_B_KpRwIewu3_2),.clk(gclk));
	jdff dff_A_ixjBq7ey4_0(.dout(w_n1409_0[0]),.din(w_dff_A_ixjBq7ey4_0),.clk(gclk));
	jdff dff_A_0EqgIHIf3_0(.dout(w_dff_A_ixjBq7ey4_0),.din(w_dff_A_0EqgIHIf3_0),.clk(gclk));
	jdff dff_B_w1DKnOjX2_2(.din(n968),.dout(w_dff_B_w1DKnOjX2_2),.clk(gclk));
	jdff dff_B_Ocovon7m7_2(.din(w_dff_B_w1DKnOjX2_2),.dout(w_dff_B_Ocovon7m7_2),.clk(gclk));
	jdff dff_B_BeqW3IrJ0_2(.din(w_dff_B_Ocovon7m7_2),.dout(w_dff_B_BeqW3IrJ0_2),.clk(gclk));
	jdff dff_B_O8BSADvy1_2(.din(w_dff_B_BeqW3IrJ0_2),.dout(w_dff_B_O8BSADvy1_2),.clk(gclk));
	jdff dff_B_4snys8hk0_2(.din(w_dff_B_O8BSADvy1_2),.dout(w_dff_B_4snys8hk0_2),.clk(gclk));
	jdff dff_B_NI9LZYTr6_0(.din(n1403),.dout(w_dff_B_NI9LZYTr6_0),.clk(gclk));
	jdff dff_B_qJMIxHQY4_1(.din(n1401),.dout(w_dff_B_qJMIxHQY4_1),.clk(gclk));
	jdff dff_B_rufnpOUb5_1(.din(w_dff_B_qJMIxHQY4_1),.dout(w_dff_B_rufnpOUb5_1),.clk(gclk));
	jdff dff_A_bmnWK5Td5_1(.dout(w_n651_0[1]),.din(w_dff_A_bmnWK5Td5_1),.clk(gclk));
	jdff dff_A_u4jsXSRD5_2(.dout(w_n651_0[2]),.din(w_dff_A_u4jsXSRD5_2),.clk(gclk));
	jdff dff_B_i8UCO9ug3_3(.din(n651),.dout(w_dff_B_i8UCO9ug3_3),.clk(gclk));
	jdff dff_B_dnF49iJf3_3(.din(w_dff_B_i8UCO9ug3_3),.dout(w_dff_B_dnF49iJf3_3),.clk(gclk));
	jdff dff_A_CDRu5jLO8_0(.dout(w_n650_0[0]),.din(w_dff_A_CDRu5jLO8_0),.clk(gclk));
	jdff dff_A_9amyVOl78_0(.dout(w_dff_A_CDRu5jLO8_0),.din(w_dff_A_9amyVOl78_0),.clk(gclk));
	jdff dff_A_GUVM0xNJ5_0(.dout(w_dff_A_9amyVOl78_0),.din(w_dff_A_GUVM0xNJ5_0),.clk(gclk));
	jdff dff_A_0ufqH2QY2_0(.dout(w_dff_A_GUVM0xNJ5_0),.din(w_dff_A_0ufqH2QY2_0),.clk(gclk));
	jdff dff_B_PnB00RFh4_1(.din(n1395),.dout(w_dff_B_PnB00RFh4_1),.clk(gclk));
	jdff dff_B_cSHY93X78_2(.din(n740),.dout(w_dff_B_cSHY93X78_2),.clk(gclk));
	jdff dff_B_kFnoWgK29_2(.din(w_dff_B_cSHY93X78_2),.dout(w_dff_B_kFnoWgK29_2),.clk(gclk));
	jdff dff_A_K7OHIxSs5_0(.dout(w_n739_1[0]),.din(w_dff_A_K7OHIxSs5_0),.clk(gclk));
	jdff dff_A_UNWT6EtT7_0(.dout(w_dff_A_K7OHIxSs5_0),.din(w_dff_A_UNWT6EtT7_0),.clk(gclk));
	jdff dff_A_coU1vn0C6_0(.dout(w_dff_A_UNWT6EtT7_0),.din(w_dff_A_coU1vn0C6_0),.clk(gclk));
	jdff dff_A_etJHdBC44_0(.dout(w_dff_A_coU1vn0C6_0),.din(w_dff_A_etJHdBC44_0),.clk(gclk));
	jdff dff_A_v1RVEhNo4_2(.dout(w_n739_0[2]),.din(w_dff_A_v1RVEhNo4_2),.clk(gclk));
	jdff dff_A_BoGRGPrV2_2(.dout(w_dff_A_v1RVEhNo4_2),.din(w_dff_A_BoGRGPrV2_2),.clk(gclk));
	jdff dff_A_G3Y4nvfc4_2(.dout(w_dff_A_BoGRGPrV2_2),.din(w_dff_A_G3Y4nvfc4_2),.clk(gclk));
	jdff dff_A_EfhrMbP10_2(.dout(w_dff_A_G3Y4nvfc4_2),.din(w_dff_A_EfhrMbP10_2),.clk(gclk));
	jdff dff_A_EvXNODuB0_2(.dout(w_n649_0[2]),.din(w_dff_A_EvXNODuB0_2),.clk(gclk));
	jdff dff_B_QqwOgu0G4_0(.din(n648),.dout(w_dff_B_QqwOgu0G4_0),.clk(gclk));
	jdff dff_B_78eIDvzX2_1(.din(G323),.dout(w_dff_B_78eIDvzX2_1),.clk(gclk));
	jdff dff_A_mKm665x34_0(.dout(w_n640_1[0]),.din(w_dff_A_mKm665x34_0),.clk(gclk));
	jdff dff_A_Jr12Bcpi8_0(.dout(w_dff_A_mKm665x34_0),.din(w_dff_A_Jr12Bcpi8_0),.clk(gclk));
	jdff dff_A_LPSyP4Pt9_0(.dout(w_dff_A_Jr12Bcpi8_0),.din(w_dff_A_LPSyP4Pt9_0),.clk(gclk));
	jdff dff_A_AmHetrVC6_0(.dout(w_dff_A_LPSyP4Pt9_0),.din(w_dff_A_AmHetrVC6_0),.clk(gclk));
	jdff dff_A_XFlxTCG45_0(.dout(w_n646_0[0]),.din(w_dff_A_XFlxTCG45_0),.clk(gclk));
	jdff dff_A_4xVxefcF9_0(.dout(w_dff_A_XFlxTCG45_0),.din(w_dff_A_4xVxefcF9_0),.clk(gclk));
	jdff dff_B_2JsLxuzT3_0(.din(n644),.dout(w_dff_B_2JsLxuzT3_0),.clk(gclk));
	jdff dff_B_qtjpYBK03_1(.din(G315),.dout(w_dff_B_qtjpYBK03_1),.clk(gclk));
	jdff dff_A_wcmYu4qH4_2(.dout(w_n640_0[2]),.din(w_dff_A_wcmYu4qH4_2),.clk(gclk));
	jdff dff_A_QSWmYASL9_2(.dout(w_dff_A_wcmYu4qH4_2),.din(w_dff_A_QSWmYASL9_2),.clk(gclk));
	jdff dff_A_cXeHmrsK1_2(.dout(w_dff_A_QSWmYASL9_2),.din(w_dff_A_cXeHmrsK1_2),.clk(gclk));
	jdff dff_A_N2Dbv83U3_2(.dout(w_dff_A_cXeHmrsK1_2),.din(w_dff_A_N2Dbv83U3_2),.clk(gclk));
	jdff dff_B_PtTfgjsn3_1(.din(n637),.dout(w_dff_B_PtTfgjsn3_1),.clk(gclk));
	jdff dff_B_L47W1YaZ0_1(.din(w_dff_B_PtTfgjsn3_1),.dout(w_dff_B_L47W1YaZ0_1),.clk(gclk));
	jdff dff_B_AUXkLHfA1_1(.din(G307),.dout(w_dff_B_AUXkLHfA1_1),.clk(gclk));
	jdff dff_A_1ROaP6aB5_1(.dout(w_n1394_0[1]),.din(w_dff_A_1ROaP6aB5_1),.clk(gclk));
	jdff dff_A_Nx4u9VHS9_1(.dout(w_n633_0[1]),.din(w_dff_A_Nx4u9VHS9_1),.clk(gclk));
	jdff dff_B_N09eC2bC1_0(.din(n632),.dout(w_dff_B_N09eC2bC1_0),.clk(gclk));
	jdff dff_A_MyLlQ7YH5_0(.dout(w_n631_0[0]),.din(w_dff_A_MyLlQ7YH5_0),.clk(gclk));
	jdff dff_A_d1F1DZWd3_0(.dout(w_dff_A_MyLlQ7YH5_0),.din(w_dff_A_d1F1DZWd3_0),.clk(gclk));
	jdff dff_A_DUWzhjT65_1(.dout(w_n629_0[1]),.din(w_dff_A_DUWzhjT65_1),.clk(gclk));
	jdff dff_A_EW7Myzab6_1(.dout(w_dff_A_DUWzhjT65_1),.din(w_dff_A_EW7Myzab6_1),.clk(gclk));
	jdff dff_A_HsDMthT51_1(.dout(w_n628_0[1]),.din(w_dff_A_HsDMthT51_1),.clk(gclk));
	jdff dff_B_eHBdsIik4_0(.din(n627),.dout(w_dff_B_eHBdsIik4_0),.clk(gclk));
	jdff dff_A_JgTALPGG5_0(.dout(w_n623_0[0]),.din(w_dff_A_JgTALPGG5_0),.clk(gclk));
	jdff dff_B_IY0qRKJx2_0(.din(n616),.dout(w_dff_B_IY0qRKJx2_0),.clk(gclk));
	jdff dff_A_hwNTQuYx7_0(.dout(w_G2174_0[0]),.din(w_dff_A_hwNTQuYx7_0),.clk(gclk));
	jdff dff_A_63dm3p8a8_0(.dout(w_dff_A_hwNTQuYx7_0),.din(w_dff_A_63dm3p8a8_0),.clk(gclk));
	jdff dff_A_tfA75Vlz0_0(.dout(w_dff_A_63dm3p8a8_0),.din(w_dff_A_tfA75Vlz0_0),.clk(gclk));
	jdff dff_A_TXkRm9yv3_0(.dout(w_dff_A_tfA75Vlz0_0),.din(w_dff_A_TXkRm9yv3_0),.clk(gclk));
	jdff dff_A_MYJX4VXo0_0(.dout(w_dff_A_TXkRm9yv3_0),.din(w_dff_A_MYJX4VXo0_0),.clk(gclk));
	jdff dff_A_lwdxxGTz4_0(.dout(w_dff_A_MYJX4VXo0_0),.din(w_dff_A_lwdxxGTz4_0),.clk(gclk));
	jdff dff_A_STo9Voqn1_0(.dout(w_dff_A_lwdxxGTz4_0),.din(w_dff_A_STo9Voqn1_0),.clk(gclk));
	jdff dff_A_2jpO3pqG4_2(.dout(w_G2174_0[2]),.din(w_dff_A_2jpO3pqG4_2),.clk(gclk));
	jdff dff_A_45eAnUZd1_2(.dout(w_dff_A_2jpO3pqG4_2),.din(w_dff_A_45eAnUZd1_2),.clk(gclk));
	jdff dff_A_kUPfPcNI0_2(.dout(w_dff_A_45eAnUZd1_2),.din(w_dff_A_kUPfPcNI0_2),.clk(gclk));
	jdff dff_A_YbhPx2op1_2(.dout(w_dff_A_kUPfPcNI0_2),.din(w_dff_A_YbhPx2op1_2),.clk(gclk));
	jdff dff_A_WmAB5ocj6_2(.dout(w_dff_A_YbhPx2op1_2),.din(w_dff_A_WmAB5ocj6_2),.clk(gclk));
	jdff dff_A_AAsaCbbk5_2(.dout(w_dff_A_WmAB5ocj6_2),.din(w_dff_A_AAsaCbbk5_2),.clk(gclk));
	jdff dff_B_apOsHt3m3_1(.din(n711),.dout(w_dff_B_apOsHt3m3_1),.clk(gclk));
	jdff dff_B_uC2qMyA97_1(.din(w_dff_B_apOsHt3m3_1),.dout(w_dff_B_uC2qMyA97_1),.clk(gclk));
	jdff dff_B_ahL5F1aQ9_1(.din(n712),.dout(w_dff_B_ahL5F1aQ9_1),.clk(gclk));
	jdff dff_B_TEmQKGRc4_1(.din(w_dff_B_ahL5F1aQ9_1),.dout(w_dff_B_TEmQKGRc4_1),.clk(gclk));
	jdff dff_B_1ge2BBjr5_1(.din(n713),.dout(w_dff_B_1ge2BBjr5_1),.clk(gclk));
	jdff dff_A_cs8aPMXM3_0(.dout(w_n723_0[0]),.din(w_dff_A_cs8aPMXM3_0),.clk(gclk));
	jdff dff_A_HGohNdA72_0(.dout(w_n621_2[0]),.din(w_dff_A_HGohNdA72_0),.clk(gclk));
	jdff dff_A_ry2AKRK42_1(.dout(w_n721_0[1]),.din(w_dff_A_ry2AKRK42_1),.clk(gclk));
	jdff dff_A_DrPWSbRu9_1(.dout(w_dff_A_ry2AKRK42_1),.din(w_dff_A_DrPWSbRu9_1),.clk(gclk));
	jdff dff_A_y2ad8xAP5_1(.dout(w_dff_A_DrPWSbRu9_1),.din(w_dff_A_y2ad8xAP5_1),.clk(gclk));
	jdff dff_A_vPdbNkDr1_0(.dout(w_G358_0[0]),.din(w_dff_A_vPdbNkDr1_0),.clk(gclk));
	jdff dff_A_MLsveOjQ4_1(.dout(w_n717_0[1]),.din(w_dff_A_MLsveOjQ4_1),.clk(gclk));
	jdff dff_A_qauZ8gI89_1(.dout(w_dff_A_MLsveOjQ4_1),.din(w_dff_A_qauZ8gI89_1),.clk(gclk));
	jdff dff_A_2YaYhArt2_2(.dout(w_n717_0[2]),.din(w_dff_A_2YaYhArt2_2),.clk(gclk));
	jdff dff_A_mQjqQizc4_0(.dout(w_G348_0[0]),.din(w_dff_A_mQjqQizc4_0),.clk(gclk));
	jdff dff_A_C1ZAZGdu3_0(.dout(w_G332_2[0]),.din(w_dff_A_C1ZAZGdu3_0),.clk(gclk));
	jdff dff_A_Qh9JfHui7_0(.dout(w_G332_3[0]),.din(w_dff_A_Qh9JfHui7_0),.clk(gclk));
	jdff dff_A_SQnpHEaN0_2(.dout(w_G332_3[2]),.din(w_dff_A_SQnpHEaN0_2),.clk(gclk));
	jdff dff_A_GJhqp7rA4_0(.dout(w_n410_1[0]),.din(w_dff_A_GJhqp7rA4_0),.clk(gclk));
	jdff dff_A_BNmdF2OE6_0(.dout(w_n614_2[0]),.din(w_dff_A_BNmdF2OE6_0),.clk(gclk));
	jdff dff_B_qSdA76el8_1(.din(n610),.dout(w_dff_B_qSdA76el8_1),.clk(gclk));
	jdff dff_B_bBt0olEp2_1(.din(w_dff_B_qSdA76el8_1),.dout(w_dff_B_bBt0olEp2_1),.clk(gclk));
	jdff dff_A_XLxZLxTv8_0(.dout(w_G332_4[0]),.din(w_dff_A_XLxZLxTv8_0),.clk(gclk));
	jdff dff_A_GdXNJ0p72_2(.dout(w_G332_1[2]),.din(w_dff_A_GdXNJ0p72_2),.clk(gclk));
	jdff dff_A_ad3WK7eX1_1(.dout(w_G331_0[1]),.din(w_dff_A_ad3WK7eX1_1),.clk(gclk));
	jdff dff_A_xq5uLGyz1_0(.dout(w_n1391_0[0]),.din(w_dff_A_xq5uLGyz1_0),.clk(gclk));
	jdff dff_A_eQP8c7Jd2_0(.dout(w_dff_A_xq5uLGyz1_0),.din(w_dff_A_eQP8c7Jd2_0),.clk(gclk));
	jdff dff_A_o4GHBTC55_0(.dout(w_dff_A_eQP8c7Jd2_0),.din(w_dff_A_o4GHBTC55_0),.clk(gclk));
	jdff dff_B_ERBCSkDC7_1(.din(n1389),.dout(w_dff_B_ERBCSkDC7_1),.clk(gclk));
	jdff dff_A_XdoSacvi2_1(.dout(w_G4091_1[1]),.din(w_dff_A_XdoSacvi2_1),.clk(gclk));
	jdff dff_A_fCXREFVt6_1(.dout(w_dff_A_XdoSacvi2_1),.din(w_dff_A_fCXREFVt6_1),.clk(gclk));
	jdff dff_A_RZM6XJEj9_1(.dout(w_dff_A_fCXREFVt6_1),.din(w_dff_A_RZM6XJEj9_1),.clk(gclk));
	jdff dff_A_QxuUtuVM6_1(.dout(w_dff_A_RZM6XJEj9_1),.din(w_dff_A_QxuUtuVM6_1),.clk(gclk));
	jdff dff_A_DbdoA8zo3_1(.dout(w_dff_A_QxuUtuVM6_1),.din(w_dff_A_DbdoA8zo3_1),.clk(gclk));
	jdff dff_A_0fg3PRYx0_1(.dout(w_dff_A_DbdoA8zo3_1),.din(w_dff_A_0fg3PRYx0_1),.clk(gclk));
	jdff dff_A_vPlwieRL3_1(.dout(w_dff_A_0fg3PRYx0_1),.din(w_dff_A_vPlwieRL3_1),.clk(gclk));
	jdff dff_A_mFCRSRPz5_1(.dout(w_dff_A_vPlwieRL3_1),.din(w_dff_A_mFCRSRPz5_1),.clk(gclk));
	jdff dff_A_pwgMBxzc3_1(.dout(w_dff_A_mFCRSRPz5_1),.din(w_dff_A_pwgMBxzc3_1),.clk(gclk));
	jdff dff_A_rNNYK3CC2_1(.dout(w_dff_A_pwgMBxzc3_1),.din(w_dff_A_rNNYK3CC2_1),.clk(gclk));
	jdff dff_A_GsGWKxYK5_1(.dout(w_dff_A_rNNYK3CC2_1),.din(w_dff_A_GsGWKxYK5_1),.clk(gclk));
	jdff dff_A_B3StbEzu5_2(.dout(w_G4091_1[2]),.din(w_dff_A_B3StbEzu5_2),.clk(gclk));
	jdff dff_A_hAVoL98k3_2(.dout(w_dff_A_B3StbEzu5_2),.din(w_dff_A_hAVoL98k3_2),.clk(gclk));
	jdff dff_A_wLE58KEQ9_2(.dout(w_dff_A_hAVoL98k3_2),.din(w_dff_A_wLE58KEQ9_2),.clk(gclk));
	jdff dff_A_qB8LxgmY1_2(.dout(w_dff_A_wLE58KEQ9_2),.din(w_dff_A_qB8LxgmY1_2),.clk(gclk));
	jdff dff_A_AJ0pjxUi0_2(.dout(w_dff_A_qB8LxgmY1_2),.din(w_dff_A_AJ0pjxUi0_2),.clk(gclk));
	jdff dff_A_If7em4U27_2(.dout(w_dff_A_AJ0pjxUi0_2),.din(w_dff_A_If7em4U27_2),.clk(gclk));
	jdff dff_A_EMgxuTUe0_2(.dout(w_dff_A_If7em4U27_2),.din(w_dff_A_EMgxuTUe0_2),.clk(gclk));
	jdff dff_A_thHBqV6D1_2(.dout(w_dff_A_EMgxuTUe0_2),.din(w_dff_A_thHBqV6D1_2),.clk(gclk));
	jdff dff_A_qJ8L9seo0_0(.dout(w_n1383_0[0]),.din(w_dff_A_qJ8L9seo0_0),.clk(gclk));
	jdff dff_A_6wIWtBnV1_0(.dout(w_dff_A_qJ8L9seo0_0),.din(w_dff_A_6wIWtBnV1_0),.clk(gclk));
	jdff dff_B_Q4zcJ1XI4_1(.din(n1363),.dout(w_dff_B_Q4zcJ1XI4_1),.clk(gclk));
	jdff dff_B_5NGtMF6T2_0(.din(n1375),.dout(w_dff_B_5NGtMF6T2_0),.clk(gclk));
	jdff dff_A_CDFLFID79_1(.dout(w_n426_0[1]),.din(w_dff_A_CDFLFID79_1),.clk(gclk));
	jdff dff_A_kUrqyGKP4_0(.dout(w_G503_1[0]),.din(w_dff_A_kUrqyGKP4_0),.clk(gclk));
	jdff dff_A_Lwvf9oX12_0(.dout(w_dff_A_kUrqyGKP4_0),.din(w_dff_A_Lwvf9oX12_0),.clk(gclk));
	jdff dff_A_pBdrQaSq8_0(.dout(w_dff_A_Lwvf9oX12_0),.din(w_dff_A_pBdrQaSq8_0),.clk(gclk));
	jdff dff_A_FnOpcfzC2_0(.dout(w_dff_A_pBdrQaSq8_0),.din(w_dff_A_FnOpcfzC2_0),.clk(gclk));
	jdff dff_A_yCbNsVp33_1(.dout(w_G503_1[1]),.din(w_dff_A_yCbNsVp33_1),.clk(gclk));
	jdff dff_A_iPQ35uet1_1(.dout(w_G503_0[1]),.din(w_dff_A_iPQ35uet1_1),.clk(gclk));
	jdff dff_A_2TZ0HTV80_1(.dout(w_dff_A_iPQ35uet1_1),.din(w_dff_A_2TZ0HTV80_1),.clk(gclk));
	jdff dff_A_6NnNjB6v3_2(.dout(w_G503_0[2]),.din(w_dff_A_6NnNjB6v3_2),.clk(gclk));
	jdff dff_A_fbYWB9YI0_2(.dout(w_dff_A_6NnNjB6v3_2),.din(w_dff_A_fbYWB9YI0_2),.clk(gclk));
	jdff dff_A_RNhbJnaP4_2(.dout(w_dff_A_fbYWB9YI0_2),.din(w_dff_A_RNhbJnaP4_2),.clk(gclk));
	jdff dff_A_QtjbEeNI5_2(.dout(w_dff_A_RNhbJnaP4_2),.din(w_dff_A_QtjbEeNI5_2),.clk(gclk));
	jdff dff_A_na05WsST4_1(.dout(w_G324_1[1]),.din(w_dff_A_na05WsST4_1),.clk(gclk));
	jdff dff_A_0MXc5Cex0_1(.dout(w_G324_0[1]),.din(w_dff_A_0MXc5Cex0_1),.clk(gclk));
	jdff dff_B_MWMKD1DM0_1(.din(n1368),.dout(w_dff_B_MWMKD1DM0_1),.clk(gclk));
	jdff dff_B_mWIbgAuX5_1(.din(w_dff_B_MWMKD1DM0_1),.dout(w_dff_B_mWIbgAuX5_1),.clk(gclk));
	jdff dff_A_gxRtB9es3_0(.dout(w_n388_0[0]),.din(w_dff_A_gxRtB9es3_0),.clk(gclk));
	jdff dff_A_cLtBuRqT4_2(.dout(w_n388_0[2]),.din(w_dff_A_cLtBuRqT4_2),.clk(gclk));
	jdff dff_A_GcIbqoCF5_0(.dout(w_G534_1[0]),.din(w_dff_A_GcIbqoCF5_0),.clk(gclk));
	jdff dff_A_h3pchY909_0(.dout(w_dff_A_GcIbqoCF5_0),.din(w_dff_A_h3pchY909_0),.clk(gclk));
	jdff dff_A_sd7fZ1847_1(.dout(w_G534_1[1]),.din(w_dff_A_sd7fZ1847_1),.clk(gclk));
	jdff dff_B_aVuxNvvi6_1(.din(n1364),.dout(w_dff_B_aVuxNvvi6_1),.clk(gclk));
	jdff dff_A_5PM0iRLc9_1(.dout(w_G351_2[1]),.din(w_dff_A_5PM0iRLc9_1),.clk(gclk));
	jdff dff_A_gVDVdBJY9_1(.dout(w_G534_0[1]),.din(w_dff_A_gVDVdBJY9_1),.clk(gclk));
	jdff dff_A_2mwCsm4j6_2(.dout(w_G534_0[2]),.din(w_dff_A_2mwCsm4j6_2),.clk(gclk));
	jdff dff_A_NIGnlWba9_2(.dout(w_dff_A_2mwCsm4j6_2),.din(w_dff_A_NIGnlWba9_2),.clk(gclk));
	jdff dff_A_OGSlSAjg7_0(.dout(w_G351_1[0]),.din(w_dff_A_OGSlSAjg7_0),.clk(gclk));
	jdff dff_A_AnvJjx9h2_2(.dout(w_n410_0[2]),.din(w_dff_A_AnvJjx9h2_2),.clk(gclk));
	jdff dff_A_TQfhw9Mw6_1(.dout(w_G514_0[1]),.din(w_dff_A_TQfhw9Mw6_1),.clk(gclk));
	jdff dff_A_K6TAvHT69_2(.dout(w_G514_0[2]),.din(w_dff_A_K6TAvHT69_2),.clk(gclk));
	jdff dff_A_MLS9kANA5_2(.dout(w_dff_A_K6TAvHT69_2),.din(w_dff_A_MLS9kANA5_2),.clk(gclk));
	jdff dff_A_kj64doxa1_1(.dout(w_G361_0[1]),.din(w_dff_A_kj64doxa1_1),.clk(gclk));
	jdff dff_B_0n2IaQjd2_1(.din(n1354),.dout(w_dff_B_0n2IaQjd2_1),.clk(gclk));
	jdff dff_B_BboVEPTk3_1(.din(w_dff_B_0n2IaQjd2_1),.dout(w_dff_B_BboVEPTk3_1),.clk(gclk));
	jdff dff_B_MHBdHR0n1_0(.din(n377),.dout(w_dff_B_MHBdHR0n1_0),.clk(gclk));
	jdff dff_A_3hOdmrop4_0(.dout(w_G490_1[0]),.din(w_dff_A_3hOdmrop4_0),.clk(gclk));
	jdff dff_A_DyUcskyR5_0(.dout(w_dff_A_3hOdmrop4_0),.din(w_dff_A_DyUcskyR5_0),.clk(gclk));
	jdff dff_A_cO9Gr6OZ1_1(.dout(w_G490_1[1]),.din(w_dff_A_cO9Gr6OZ1_1),.clk(gclk));
	jdff dff_A_F0OTlOFe7_1(.dout(w_dff_A_cO9Gr6OZ1_1),.din(w_dff_A_F0OTlOFe7_1),.clk(gclk));
	jdff dff_A_Ac2yJfaK8_1(.dout(w_G490_0[1]),.din(w_dff_A_Ac2yJfaK8_1),.clk(gclk));
	jdff dff_A_MKWq9gVH1_1(.dout(w_dff_A_Ac2yJfaK8_1),.din(w_dff_A_MKWq9gVH1_1),.clk(gclk));
	jdff dff_A_P03s7JlX1_2(.dout(w_G490_0[2]),.din(w_dff_A_P03s7JlX1_2),.clk(gclk));
	jdff dff_A_atVKGEcb4_2(.dout(w_dff_A_P03s7JlX1_2),.din(w_dff_A_atVKGEcb4_2),.clk(gclk));
	jdff dff_A_0ZhmUMim8_0(.dout(w_G316_1[0]),.din(w_dff_A_0ZhmUMim8_0),.clk(gclk));
	jdff dff_B_e1go9qx96_0(.din(n364),.dout(w_dff_B_e1go9qx96_0),.clk(gclk));
	jdff dff_A_oXlSBaSx5_0(.dout(w_n362_0[0]),.din(w_dff_A_oXlSBaSx5_0),.clk(gclk));
	jdff dff_A_d5VI5gxX9_0(.dout(w_dff_A_oXlSBaSx5_0),.din(w_dff_A_d5VI5gxX9_0),.clk(gclk));
	jdff dff_A_6R23NZgw3_0(.dout(w_G479_1[0]),.din(w_dff_A_6R23NZgw3_0),.clk(gclk));
	jdff dff_A_gVYY9rGg0_0(.dout(w_dff_A_6R23NZgw3_0),.din(w_dff_A_gVYY9rGg0_0),.clk(gclk));
	jdff dff_A_eEayZ6AJ4_1(.dout(w_G479_0[1]),.din(w_dff_A_eEayZ6AJ4_1),.clk(gclk));
	jdff dff_A_fMXpPf7C0_1(.dout(w_dff_A_eEayZ6AJ4_1),.din(w_dff_A_fMXpPf7C0_1),.clk(gclk));
	jdff dff_A_FHY5TT1y0_2(.dout(w_G479_0[2]),.din(w_dff_A_FHY5TT1y0_2),.clk(gclk));
	jdff dff_A_0x3qhw4g3_2(.dout(w_dff_A_FHY5TT1y0_2),.din(w_dff_A_0x3qhw4g3_2),.clk(gclk));
	jdff dff_A_bZHPyQTY7_0(.dout(w_G308_1[0]),.din(w_dff_A_bZHPyQTY7_0),.clk(gclk));
	jdff dff_A_Jnph24Rg6_0(.dout(w_G302_0[0]),.din(w_dff_A_Jnph24Rg6_0),.clk(gclk));
	jdff dff_A_TNwFbmIf5_1(.dout(w_G302_0[1]),.din(w_dff_A_TNwFbmIf5_1),.clk(gclk));
	jdff dff_A_5kixj4V24_0(.dout(w_n401_0[0]),.din(w_dff_A_5kixj4V24_0),.clk(gclk));
	jdff dff_A_XsN8yS8u2_2(.dout(w_n401_0[2]),.din(w_dff_A_XsN8yS8u2_2),.clk(gclk));
	jdff dff_A_W8Mlyg2V4_1(.dout(w_G293_0[1]),.din(w_dff_A_W8Mlyg2V4_1),.clk(gclk));
	jdff dff_B_aHlrTtf12_0(.din(n1348),.dout(w_dff_B_aHlrTtf12_0),.clk(gclk));
	jdff dff_A_6dzRm1Bg9_0(.dout(w_n437_0[0]),.din(w_dff_A_6dzRm1Bg9_0),.clk(gclk));
	jdff dff_A_fDbBMFjd2_2(.dout(w_n437_0[2]),.din(w_dff_A_fDbBMFjd2_2),.clk(gclk));
	jdff dff_A_SM2qFWos7_0(.dout(w_G523_1[0]),.din(w_dff_A_SM2qFWos7_0),.clk(gclk));
	jdff dff_A_cu79otYr7_1(.dout(w_G523_0[1]),.din(w_dff_A_cu79otYr7_1),.clk(gclk));
	jdff dff_A_OzvjWbRM9_1(.dout(w_dff_A_cu79otYr7_1),.din(w_dff_A_OzvjWbRM9_1),.clk(gclk));
	jdff dff_A_KozyfIKl5_2(.dout(w_G523_0[2]),.din(w_dff_A_KozyfIKl5_2),.clk(gclk));
	jdff dff_A_jAj800uz2_2(.dout(w_dff_A_KozyfIKl5_2),.din(w_dff_A_jAj800uz2_2),.clk(gclk));
	jdff dff_A_S7x97lQ49_1(.dout(w_G341_2[1]),.din(w_dff_A_S7x97lQ49_1),.clk(gclk));
	jdff dff_A_Yk7dySkI4_2(.dout(w_G341_0[2]),.din(w_dff_A_Yk7dySkI4_2),.clk(gclk));
	jdff dff_A_TnGIPudw5_2(.dout(w_n746_0[2]),.din(w_dff_A_TnGIPudw5_2),.clk(gclk));
	jdff dff_A_6EVykQ313_2(.dout(w_dff_A_TnGIPudw5_2),.din(w_dff_A_6EVykQ313_2),.clk(gclk));
	jdff dff_A_1ajh71Lv4_2(.dout(w_dff_A_6EVykQ313_2),.din(w_dff_A_1ajh71Lv4_2),.clk(gclk));
	jdff dff_A_asEazgg44_2(.dout(w_dff_A_1ajh71Lv4_2),.din(w_dff_A_asEazgg44_2),.clk(gclk));
	jdff dff_A_9WMDtgRQ9_2(.dout(w_dff_A_asEazgg44_2),.din(w_dff_A_9WMDtgRQ9_2),.clk(gclk));
	jdff dff_A_YSMGR71D3_2(.dout(w_dff_A_9WMDtgRQ9_2),.din(w_dff_A_YSMGR71D3_2),.clk(gclk));
	jdff dff_A_MWIaVXE52_2(.dout(w_dff_A_YSMGR71D3_2),.din(w_dff_A_MWIaVXE52_2),.clk(gclk));
	jdff dff_A_7j0KxMEI6_0(.dout(w_n1002_1[0]),.din(w_dff_A_7j0KxMEI6_0),.clk(gclk));
	jdff dff_A_qzgnXvTw3_0(.dout(w_dff_A_7j0KxMEI6_0),.din(w_dff_A_qzgnXvTw3_0),.clk(gclk));
	jdff dff_A_SzPMDIlA3_0(.dout(w_dff_A_qzgnXvTw3_0),.din(w_dff_A_SzPMDIlA3_0),.clk(gclk));
	jdff dff_A_HgKl2ejf3_0(.dout(w_dff_A_SzPMDIlA3_0),.din(w_dff_A_HgKl2ejf3_0),.clk(gclk));
	jdff dff_A_hpWNJz8J2_2(.dout(w_n1002_1[2]),.din(w_dff_A_hpWNJz8J2_2),.clk(gclk));
	jdff dff_A_yUafKato1_2(.dout(w_dff_A_hpWNJz8J2_2),.din(w_dff_A_yUafKato1_2),.clk(gclk));
	jdff dff_A_OJM2wDhK4_2(.dout(w_dff_A_yUafKato1_2),.din(w_dff_A_OJM2wDhK4_2),.clk(gclk));
	jdff dff_A_8pQ9if736_2(.dout(w_dff_A_OJM2wDhK4_2),.din(w_dff_A_8pQ9if736_2),.clk(gclk));
	jdff dff_A_9EOsrfw04_2(.dout(w_dff_A_8pQ9if736_2),.din(w_dff_A_9EOsrfw04_2),.clk(gclk));
	jdff dff_A_ACt647wx5_2(.dout(w_dff_A_9EOsrfw04_2),.din(w_dff_A_ACt647wx5_2),.clk(gclk));
	jdff dff_A_pmETJqGf8_2(.dout(w_dff_A_ACt647wx5_2),.din(w_dff_A_pmETJqGf8_2),.clk(gclk));
	jdff dff_A_23xNqoGD4_2(.dout(w_dff_A_pmETJqGf8_2),.din(w_dff_A_23xNqoGD4_2),.clk(gclk));
	jdff dff_A_qqem33b11_2(.dout(w_dff_A_23xNqoGD4_2),.din(w_dff_A_qqem33b11_2),.clk(gclk));
	jdff dff_A_WcsxV8R50_1(.dout(w_n1002_0[1]),.din(w_dff_A_WcsxV8R50_1),.clk(gclk));
	jdff dff_A_MbGbA55Z6_1(.dout(w_dff_A_WcsxV8R50_1),.din(w_dff_A_MbGbA55Z6_1),.clk(gclk));
	jdff dff_A_IecQwGAt9_1(.dout(w_dff_A_MbGbA55Z6_1),.din(w_dff_A_IecQwGAt9_1),.clk(gclk));
	jdff dff_A_4w7RLAhu3_1(.dout(w_dff_A_IecQwGAt9_1),.din(w_dff_A_4w7RLAhu3_1),.clk(gclk));
	jdff dff_A_XMJJW0tL8_1(.dout(w_dff_A_4w7RLAhu3_1),.din(w_dff_A_XMJJW0tL8_1),.clk(gclk));
	jdff dff_A_nATH1QcU2_1(.dout(w_dff_A_XMJJW0tL8_1),.din(w_dff_A_nATH1QcU2_1),.clk(gclk));
	jdff dff_A_0abN5IuP0_1(.dout(w_dff_A_nATH1QcU2_1),.din(w_dff_A_0abN5IuP0_1),.clk(gclk));
	jdff dff_A_AlwHnu960_1(.dout(w_dff_A_0abN5IuP0_1),.din(w_dff_A_AlwHnu960_1),.clk(gclk));
	jdff dff_A_06tVJ6yW9_1(.dout(w_dff_A_AlwHnu960_1),.din(w_dff_A_06tVJ6yW9_1),.clk(gclk));
	jdff dff_A_M5ypYtmO1_2(.dout(w_n1002_0[2]),.din(w_dff_A_M5ypYtmO1_2),.clk(gclk));
	jdff dff_A_iXloacdp9_2(.dout(w_dff_A_M5ypYtmO1_2),.din(w_dff_A_iXloacdp9_2),.clk(gclk));
	jdff dff_A_LedMmay24_2(.dout(w_dff_A_iXloacdp9_2),.din(w_dff_A_LedMmay24_2),.clk(gclk));
	jdff dff_A_GeOtFvMz8_2(.dout(w_dff_A_LedMmay24_2),.din(w_dff_A_GeOtFvMz8_2),.clk(gclk));
	jdff dff_A_XrIU7Ouo9_2(.dout(w_dff_A_GeOtFvMz8_2),.din(w_dff_A_XrIU7Ouo9_2),.clk(gclk));
	jdff dff_B_a7NpkydQ0_1(.din(n1641),.dout(w_dff_B_a7NpkydQ0_1),.clk(gclk));
	jdff dff_B_TYsxJWRF4_1(.din(w_dff_B_a7NpkydQ0_1),.dout(w_dff_B_TYsxJWRF4_1),.clk(gclk));
	jdff dff_B_9wK0nXUx1_1(.din(w_dff_B_TYsxJWRF4_1),.dout(w_dff_B_9wK0nXUx1_1),.clk(gclk));
	jdff dff_B_hZbVmIT35_1(.din(w_dff_B_9wK0nXUx1_1),.dout(w_dff_B_hZbVmIT35_1),.clk(gclk));
	jdff dff_B_yrHkSmoJ3_1(.din(w_dff_B_hZbVmIT35_1),.dout(w_dff_B_yrHkSmoJ3_1),.clk(gclk));
	jdff dff_B_7Y4A6LGo2_1(.din(w_dff_B_yrHkSmoJ3_1),.dout(w_dff_B_7Y4A6LGo2_1),.clk(gclk));
	jdff dff_B_NghpbNt44_1(.din(w_dff_B_7Y4A6LGo2_1),.dout(w_dff_B_NghpbNt44_1),.clk(gclk));
	jdff dff_B_TPpiuW7q6_1(.din(w_dff_B_NghpbNt44_1),.dout(w_dff_B_TPpiuW7q6_1),.clk(gclk));
	jdff dff_B_Lmmcwpge6_1(.din(w_dff_B_TPpiuW7q6_1),.dout(w_dff_B_Lmmcwpge6_1),.clk(gclk));
	jdff dff_B_ce0KwDZg2_1(.din(w_dff_B_Lmmcwpge6_1),.dout(w_dff_B_ce0KwDZg2_1),.clk(gclk));
	jdff dff_B_60oi5j988_1(.din(w_dff_B_ce0KwDZg2_1),.dout(w_dff_B_60oi5j988_1),.clk(gclk));
	jdff dff_B_J4oyQ6Tf1_1(.din(w_dff_B_60oi5j988_1),.dout(w_dff_B_J4oyQ6Tf1_1),.clk(gclk));
	jdff dff_B_vd96JV3q7_1(.din(w_dff_B_J4oyQ6Tf1_1),.dout(w_dff_B_vd96JV3q7_1),.clk(gclk));
	jdff dff_B_r8TMHfw99_1(.din(w_dff_B_vd96JV3q7_1),.dout(w_dff_B_r8TMHfw99_1),.clk(gclk));
	jdff dff_B_puD2XYxx4_0(.din(n1600),.dout(w_dff_B_puD2XYxx4_0),.clk(gclk));
	jdff dff_B_EYBxdOib0_0(.din(w_dff_B_puD2XYxx4_0),.dout(w_dff_B_EYBxdOib0_0),.clk(gclk));
	jdff dff_B_rqj1dBHn1_0(.din(w_dff_B_EYBxdOib0_0),.dout(w_dff_B_rqj1dBHn1_0),.clk(gclk));
	jdff dff_B_Vk5lW8kJ2_0(.din(w_dff_B_rqj1dBHn1_0),.dout(w_dff_B_Vk5lW8kJ2_0),.clk(gclk));
	jdff dff_B_mEW6uHnO7_0(.din(w_dff_B_Vk5lW8kJ2_0),.dout(w_dff_B_mEW6uHnO7_0),.clk(gclk));
	jdff dff_B_W0Xf4Z5O5_0(.din(w_dff_B_mEW6uHnO7_0),.dout(w_dff_B_W0Xf4Z5O5_0),.clk(gclk));
	jdff dff_B_gPz1QXqV5_0(.din(w_dff_B_W0Xf4Z5O5_0),.dout(w_dff_B_gPz1QXqV5_0),.clk(gclk));
	jdff dff_B_3neDW6fj7_0(.din(w_dff_B_gPz1QXqV5_0),.dout(w_dff_B_3neDW6fj7_0),.clk(gclk));
	jdff dff_B_Nt2c5WbK8_0(.din(w_dff_B_3neDW6fj7_0),.dout(w_dff_B_Nt2c5WbK8_0),.clk(gclk));
	jdff dff_B_AenvPhnV0_0(.din(w_dff_B_Nt2c5WbK8_0),.dout(w_dff_B_AenvPhnV0_0),.clk(gclk));
	jdff dff_B_ZbWxVY6Z8_0(.din(w_dff_B_AenvPhnV0_0),.dout(w_dff_B_ZbWxVY6Z8_0),.clk(gclk));
	jdff dff_B_BYbj11AS2_0(.din(w_dff_B_ZbWxVY6Z8_0),.dout(w_dff_B_BYbj11AS2_0),.clk(gclk));
	jdff dff_B_uKJRfvDV7_0(.din(w_dff_B_BYbj11AS2_0),.dout(w_dff_B_uKJRfvDV7_0),.clk(gclk));
	jdff dff_B_Oddba9KG5_0(.din(w_dff_B_uKJRfvDV7_0),.dout(w_dff_B_Oddba9KG5_0),.clk(gclk));
	jdff dff_B_lyNzQbrW4_1(.din(n1540),.dout(w_dff_B_lyNzQbrW4_1),.clk(gclk));
	jdff dff_B_fVY8S10L6_1(.din(w_dff_B_lyNzQbrW4_1),.dout(w_dff_B_fVY8S10L6_1),.clk(gclk));
	jdff dff_B_fzbEwBZS2_1(.din(w_dff_B_fVY8S10L6_1),.dout(w_dff_B_fzbEwBZS2_1),.clk(gclk));
	jdff dff_B_Jl7gnC2Q1_1(.din(w_dff_B_fzbEwBZS2_1),.dout(w_dff_B_Jl7gnC2Q1_1),.clk(gclk));
	jdff dff_B_OFt7BEtg6_1(.din(w_dff_B_Jl7gnC2Q1_1),.dout(w_dff_B_OFt7BEtg6_1),.clk(gclk));
	jdff dff_B_KkBBRbQw1_1(.din(w_dff_B_OFt7BEtg6_1),.dout(w_dff_B_KkBBRbQw1_1),.clk(gclk));
	jdff dff_B_ruE9ChaX7_1(.din(w_dff_B_KkBBRbQw1_1),.dout(w_dff_B_ruE9ChaX7_1),.clk(gclk));
	jdff dff_B_AcB2ERIg3_0(.din(n1595),.dout(w_dff_B_AcB2ERIg3_0),.clk(gclk));
	jdff dff_B_Xe7C2mQ81_1(.din(n1566),.dout(w_dff_B_Xe7C2mQ81_1),.clk(gclk));
	jdff dff_B_9sqnuwhk9_1(.din(w_dff_B_Xe7C2mQ81_1),.dout(w_dff_B_9sqnuwhk9_1),.clk(gclk));
	jdff dff_B_28Ijl9f45_0(.din(n1589),.dout(w_dff_B_28Ijl9f45_0),.clk(gclk));
	jdff dff_B_AiB4gh4m8_0(.din(w_dff_B_28Ijl9f45_0),.dout(w_dff_B_AiB4gh4m8_0),.clk(gclk));
	jdff dff_B_MMoHMBXD7_0(.din(w_dff_B_AiB4gh4m8_0),.dout(w_dff_B_MMoHMBXD7_0),.clk(gclk));
	jdff dff_B_g3O8EnKR9_1(.din(n1579),.dout(w_dff_B_g3O8EnKR9_1),.clk(gclk));
	jdff dff_B_PwDiaseQ0_0(.din(n1584),.dout(w_dff_B_PwDiaseQ0_0),.clk(gclk));
	jdff dff_B_vmJBUhKe9_1(.din(n1567),.dout(w_dff_B_vmJBUhKe9_1),.clk(gclk));
	jdff dff_B_B1P9dUjr7_1(.din(w_dff_B_vmJBUhKe9_1),.dout(w_dff_B_B1P9dUjr7_1),.clk(gclk));
	jdff dff_B_dS49bua96_1(.din(w_dff_B_B1P9dUjr7_1),.dout(w_dff_B_dS49bua96_1),.clk(gclk));
	jdff dff_B_8sHUGYlX8_1(.din(w_dff_B_dS49bua96_1),.dout(w_dff_B_8sHUGYlX8_1),.clk(gclk));
	jdff dff_B_rbRekOsa1_1(.din(w_dff_B_8sHUGYlX8_1),.dout(w_dff_B_rbRekOsa1_1),.clk(gclk));
	jdff dff_B_cFzSoUsO2_1(.din(w_dff_B_rbRekOsa1_1),.dout(w_dff_B_cFzSoUsO2_1),.clk(gclk));
	jdff dff_B_vIv3LLS91_1(.din(w_dff_B_cFzSoUsO2_1),.dout(w_dff_B_vIv3LLS91_1),.clk(gclk));
	jdff dff_B_o40UGd8j8_1(.din(w_dff_B_vIv3LLS91_1),.dout(w_dff_B_o40UGd8j8_1),.clk(gclk));
	jdff dff_B_VkAZvjam5_1(.din(w_dff_B_o40UGd8j8_1),.dout(w_dff_B_VkAZvjam5_1),.clk(gclk));
	jdff dff_B_BMknLLvv6_1(.din(w_dff_B_VkAZvjam5_1),.dout(w_dff_B_BMknLLvv6_1),.clk(gclk));
	jdff dff_B_kgYAeSDA7_1(.din(n1570),.dout(w_dff_B_kgYAeSDA7_1),.clk(gclk));
	jdff dff_B_903H55d30_1(.din(w_dff_B_kgYAeSDA7_1),.dout(w_dff_B_903H55d30_1),.clk(gclk));
	jdff dff_B_Glpa9uIe1_1(.din(n1571),.dout(w_dff_B_Glpa9uIe1_1),.clk(gclk));
	jdff dff_B_hvNLbXMv0_1(.din(w_dff_B_Glpa9uIe1_1),.dout(w_dff_B_hvNLbXMv0_1),.clk(gclk));
	jdff dff_B_iCKgjrF94_1(.din(w_dff_B_hvNLbXMv0_1),.dout(w_dff_B_iCKgjrF94_1),.clk(gclk));
	jdff dff_B_4PpQDkje0_1(.din(w_dff_B_iCKgjrF94_1),.dout(w_dff_B_4PpQDkje0_1),.clk(gclk));
	jdff dff_B_ZkE0SPhO5_0(.din(n1574),.dout(w_dff_B_ZkE0SPhO5_0),.clk(gclk));
	jdff dff_A_pddUHG9k4_1(.dout(w_n853_0[1]),.din(w_dff_A_pddUHG9k4_1),.clk(gclk));
	jdff dff_B_h7Crkwla2_2(.din(n853),.dout(w_dff_B_h7Crkwla2_2),.clk(gclk));
	jdff dff_B_ID5YT5Fh9_2(.din(w_dff_B_h7Crkwla2_2),.dout(w_dff_B_ID5YT5Fh9_2),.clk(gclk));
	jdff dff_B_E3ZWldZh9_2(.din(w_dff_B_ID5YT5Fh9_2),.dout(w_dff_B_E3ZWldZh9_2),.clk(gclk));
	jdff dff_B_WzfnIOVU6_2(.din(w_dff_B_E3ZWldZh9_2),.dout(w_dff_B_WzfnIOVU6_2),.clk(gclk));
	jdff dff_A_mVU5x45s0_0(.dout(w_n681_1[0]),.din(w_dff_A_mVU5x45s0_0),.clk(gclk));
	jdff dff_A_2ebXTWkX1_0(.dout(w_dff_A_mVU5x45s0_0),.din(w_dff_A_2ebXTWkX1_0),.clk(gclk));
	jdff dff_A_50lyW5Wd4_1(.dout(w_n681_1[1]),.din(w_dff_A_50lyW5Wd4_1),.clk(gclk));
	jdff dff_A_DmbG28e35_1(.dout(w_n1568_0[1]),.din(w_dff_A_DmbG28e35_1),.clk(gclk));
	jdff dff_B_vMN4xilR7_2(.din(n1568),.dout(w_dff_B_vMN4xilR7_2),.clk(gclk));
	jdff dff_B_VBxjGP5o5_0(.din(n1563),.dout(w_dff_B_VBxjGP5o5_0),.clk(gclk));
	jdff dff_A_JfvCvCPd3_0(.dout(w_n1555_0[0]),.din(w_dff_A_JfvCvCPd3_0),.clk(gclk));
	jdff dff_B_OmSN4Hff7_2(.din(n1553),.dout(w_dff_B_OmSN4Hff7_2),.clk(gclk));
	jdff dff_B_IJ6EX7S53_2(.din(w_dff_B_OmSN4Hff7_2),.dout(w_dff_B_IJ6EX7S53_2),.clk(gclk));
	jdff dff_B_3dRmf2ut7_2(.din(w_dff_B_IJ6EX7S53_2),.dout(w_dff_B_3dRmf2ut7_2),.clk(gclk));
	jdff dff_B_3OqlOmy05_0(.din(n1551),.dout(w_dff_B_3OqlOmy05_0),.clk(gclk));
	jdff dff_B_8pmLg6vj4_0(.din(n1550),.dout(w_dff_B_8pmLg6vj4_0),.clk(gclk));
	jdff dff_B_O4SYiGmJ5_0(.din(w_dff_B_8pmLg6vj4_0),.dout(w_dff_B_O4SYiGmJ5_0),.clk(gclk));
	jdff dff_B_ULwlZ6nV6_0(.din(w_dff_B_O4SYiGmJ5_0),.dout(w_dff_B_ULwlZ6nV6_0),.clk(gclk));
	jdff dff_A_fMprN1J51_2(.dout(w_n605_1[2]),.din(w_dff_A_fMprN1J51_2),.clk(gclk));
	jdff dff_A_en7ad1Kn4_2(.dout(w_dff_A_fMprN1J51_2),.din(w_dff_A_en7ad1Kn4_2),.clk(gclk));
	jdff dff_A_WLOZ7s6Q0_2(.dout(w_dff_A_en7ad1Kn4_2),.din(w_dff_A_WLOZ7s6Q0_2),.clk(gclk));
	jdff dff_A_BuNbo8jw9_2(.dout(w_dff_A_WLOZ7s6Q0_2),.din(w_dff_A_BuNbo8jw9_2),.clk(gclk));
	jdff dff_A_56x25ONW9_2(.dout(w_dff_A_BuNbo8jw9_2),.din(w_dff_A_56x25ONW9_2),.clk(gclk));
	jdff dff_A_c6TOSdvJ3_2(.dout(w_dff_A_56x25ONW9_2),.din(w_dff_A_c6TOSdvJ3_2),.clk(gclk));
	jdff dff_A_56NzQtJd9_2(.dout(w_dff_A_c6TOSdvJ3_2),.din(w_dff_A_56NzQtJd9_2),.clk(gclk));
	jdff dff_A_GhjW42Og9_2(.dout(w_dff_A_56NzQtJd9_2),.din(w_dff_A_GhjW42Og9_2),.clk(gclk));
	jdff dff_A_GZztyjC65_0(.dout(w_n948_0[0]),.din(w_dff_A_GZztyjC65_0),.clk(gclk));
	jdff dff_A_o9kwGvjU0_1(.dout(w_n948_0[1]),.din(w_dff_A_o9kwGvjU0_1),.clk(gclk));
	jdff dff_A_RgqKSrrU3_1(.dout(w_n944_0[1]),.din(w_dff_A_RgqKSrrU3_1),.clk(gclk));
	jdff dff_A_mq9RuaIy5_1(.dout(w_dff_A_RgqKSrrU3_1),.din(w_dff_A_mq9RuaIy5_1),.clk(gclk));
	jdff dff_A_raj9x4Dl2_1(.dout(w_dff_A_mq9RuaIy5_1),.din(w_dff_A_raj9x4Dl2_1),.clk(gclk));
	jdff dff_A_9AA4jxtz7_1(.dout(w_dff_A_raj9x4Dl2_1),.din(w_dff_A_9AA4jxtz7_1),.clk(gclk));
	jdff dff_A_qTwRcuC64_1(.dout(w_dff_A_9AA4jxtz7_1),.din(w_dff_A_qTwRcuC64_1),.clk(gclk));
	jdff dff_A_t5vzpAcD6_2(.dout(w_n930_0[2]),.din(w_dff_A_t5vzpAcD6_2),.clk(gclk));
	jdff dff_A_XqPQdzNs6_2(.dout(w_dff_A_t5vzpAcD6_2),.din(w_dff_A_XqPQdzNs6_2),.clk(gclk));
	jdff dff_A_5hchiyYo2_2(.dout(w_dff_A_XqPQdzNs6_2),.din(w_dff_A_5hchiyYo2_2),.clk(gclk));
	jdff dff_A_DzwLaq156_2(.dout(w_dff_A_5hchiyYo2_2),.din(w_dff_A_DzwLaq156_2),.clk(gclk));
	jdff dff_A_iFfrMLOE4_2(.dout(w_dff_A_DzwLaq156_2),.din(w_dff_A_iFfrMLOE4_2),.clk(gclk));
	jdff dff_B_zYtFHTP31_3(.din(n930),.dout(w_dff_B_zYtFHTP31_3),.clk(gclk));
	jdff dff_B_E3phhCox2_3(.din(w_dff_B_zYtFHTP31_3),.dout(w_dff_B_E3phhCox2_3),.clk(gclk));
	jdff dff_A_zfuHo9Re4_1(.dout(w_n700_0[1]),.din(w_dff_A_zfuHo9Re4_1),.clk(gclk));
	jdff dff_A_K4XQ6b8l3_1(.dout(w_dff_A_zfuHo9Re4_1),.din(w_dff_A_K4XQ6b8l3_1),.clk(gclk));
	jdff dff_A_QuPSF2du9_0(.dout(w_n706_0[0]),.din(w_dff_A_QuPSF2du9_0),.clk(gclk));
	jdff dff_B_dsPbd1ZL5_1(.din(n701),.dout(w_dff_B_dsPbd1ZL5_1),.clk(gclk));
	jdff dff_B_G7uNY9om7_0(.din(n599),.dout(w_dff_B_G7uNY9om7_0),.clk(gclk));
	jdff dff_B_sWj5ZqZw4_1(.din(G233),.dout(w_dff_B_sWj5ZqZw4_1),.clk(gclk));
	jdff dff_B_c7Q5rMIL4_2(.din(n702),.dout(w_dff_B_c7Q5rMIL4_2),.clk(gclk));
	jdff dff_A_0QktJ4318_0(.dout(w_n604_0[0]),.din(w_dff_A_0QktJ4318_0),.clk(gclk));
	jdff dff_A_X9guJ0Ki5_0(.dout(w_dff_A_0QktJ4318_0),.din(w_dff_A_X9guJ0Ki5_0),.clk(gclk));
	jdff dff_B_IEvps7dX4_0(.din(n603),.dout(w_dff_B_IEvps7dX4_0),.clk(gclk));
	jdff dff_B_RwvYYWHM3_1(.din(G225),.dout(w_dff_B_RwvYYWHM3_1),.clk(gclk));
	jdff dff_A_JhNsed8J2_1(.dout(w_n928_0[1]),.din(w_dff_A_JhNsed8J2_1),.clk(gclk));
	jdff dff_A_9po5nfMh2_1(.dout(w_dff_A_JhNsed8J2_1),.din(w_dff_A_9po5nfMh2_1),.clk(gclk));
	jdff dff_A_fRsPcMSn4_1(.dout(w_dff_A_9po5nfMh2_1),.din(w_dff_A_fRsPcMSn4_1),.clk(gclk));
	jdff dff_A_kzBFYKwr1_1(.dout(w_dff_A_fRsPcMSn4_1),.din(w_dff_A_kzBFYKwr1_1),.clk(gclk));
	jdff dff_A_ElfGvmoY0_1(.dout(w_dff_A_kzBFYKwr1_1),.din(w_dff_A_ElfGvmoY0_1),.clk(gclk));
	jdff dff_A_Vrj1WP1J8_0(.dout(w_n596_0[0]),.din(w_dff_A_Vrj1WP1J8_0),.clk(gclk));
	jdff dff_B_w4lX7e4x9_1(.din(n592),.dout(w_dff_B_w4lX7e4x9_1),.clk(gclk));
	jdff dff_B_DFcrzi0Y8_1(.din(w_dff_B_w4lX7e4x9_1),.dout(w_dff_B_DFcrzi0Y8_1),.clk(gclk));
	jdff dff_B_MxggyYSc5_1(.din(G209),.dout(w_dff_B_MxggyYSc5_1),.clk(gclk));
	jdff dff_B_ZZh5tCdu9_0(.din(n584),.dout(w_dff_B_ZZh5tCdu9_0),.clk(gclk));
	jdff dff_B_OHyepcNP0_0(.din(w_dff_B_ZZh5tCdu9_0),.dout(w_dff_B_OHyepcNP0_0),.clk(gclk));
	jdff dff_B_U8qwk8bP1_0(.din(w_dff_B_OHyepcNP0_0),.dout(w_dff_B_U8qwk8bP1_0),.clk(gclk));
	jdff dff_A_MnCHQddv6_0(.dout(w_n583_1[0]),.din(w_dff_A_MnCHQddv6_0),.clk(gclk));
	jdff dff_A_kCz2zH7F5_0(.dout(w_dff_A_MnCHQddv6_0),.din(w_dff_A_kCz2zH7F5_0),.clk(gclk));
	jdff dff_A_f2LfcUUq5_0(.dout(w_dff_A_kCz2zH7F5_0),.din(w_dff_A_f2LfcUUq5_0),.clk(gclk));
	jdff dff_A_jG3uHNL70_0(.dout(w_n572_0[0]),.din(w_dff_A_jG3uHNL70_0),.clk(gclk));
	jdff dff_A_O923MLma9_1(.dout(w_n567_1[1]),.din(w_dff_A_O923MLma9_1),.clk(gclk));
	jdff dff_A_JgZzs1jo2_0(.dout(w_n562_0[0]),.din(w_dff_A_JgZzs1jo2_0),.clk(gclk));
	jdff dff_A_XWnsyk0Z9_0(.dout(w_dff_A_JgZzs1jo2_0),.din(w_dff_A_XWnsyk0Z9_0),.clk(gclk));
	jdff dff_A_zgU2YMnZ9_0(.dout(w_dff_A_XWnsyk0Z9_0),.din(w_dff_A_zgU2YMnZ9_0),.clk(gclk));
	jdff dff_A_Z9CoqXJ94_0(.dout(w_dff_A_zgU2YMnZ9_0),.din(w_dff_A_Z9CoqXJ94_0),.clk(gclk));
	jdff dff_A_nEV5xnJU2_1(.dout(w_n561_0[1]),.din(w_dff_A_nEV5xnJU2_1),.clk(gclk));
	jdff dff_A_khti5bYU3_1(.dout(w_dff_A_nEV5xnJU2_1),.din(w_dff_A_khti5bYU3_1),.clk(gclk));
	jdff dff_A_2P0wzb8F8_0(.dout(w_G1497_0[0]),.din(w_dff_A_2P0wzb8F8_0),.clk(gclk));
	jdff dff_A_LEr7TiXz9_0(.dout(w_dff_A_2P0wzb8F8_0),.din(w_dff_A_LEr7TiXz9_0),.clk(gclk));
	jdff dff_A_7oiQ3gwa3_0(.dout(w_dff_A_LEr7TiXz9_0),.din(w_dff_A_7oiQ3gwa3_0),.clk(gclk));
	jdff dff_A_qaAvJrj08_0(.dout(w_dff_A_7oiQ3gwa3_0),.din(w_dff_A_qaAvJrj08_0),.clk(gclk));
	jdff dff_A_vgJ2DXI13_0(.dout(w_dff_A_qaAvJrj08_0),.din(w_dff_A_vgJ2DXI13_0),.clk(gclk));
	jdff dff_A_Zf7vTtPH2_0(.dout(w_dff_A_vgJ2DXI13_0),.din(w_dff_A_Zf7vTtPH2_0),.clk(gclk));
	jdff dff_A_9ov1B3Sl8_0(.dout(w_dff_A_Zf7vTtPH2_0),.din(w_dff_A_9ov1B3Sl8_0),.clk(gclk));
	jdff dff_A_kdJh28BH4_0(.dout(w_dff_A_9ov1B3Sl8_0),.din(w_dff_A_kdJh28BH4_0),.clk(gclk));
	jdff dff_A_8BUd6CkQ8_2(.dout(w_G1497_0[2]),.din(w_dff_A_8BUd6CkQ8_2),.clk(gclk));
	jdff dff_A_jlzzTimf3_2(.dout(w_dff_A_8BUd6CkQ8_2),.din(w_dff_A_jlzzTimf3_2),.clk(gclk));
	jdff dff_A_eH6lPn1M8_2(.dout(w_dff_A_jlzzTimf3_2),.din(w_dff_A_eH6lPn1M8_2),.clk(gclk));
	jdff dff_A_VnWqJ54o4_2(.dout(w_dff_A_eH6lPn1M8_2),.din(w_dff_A_VnWqJ54o4_2),.clk(gclk));
	jdff dff_A_02evRjqD3_2(.dout(w_dff_A_VnWqJ54o4_2),.din(w_dff_A_02evRjqD3_2),.clk(gclk));
	jdff dff_A_h8mlJ5ry7_2(.dout(w_dff_A_02evRjqD3_2),.din(w_dff_A_h8mlJ5ry7_2),.clk(gclk));
	jdff dff_A_G5zBqwwm1_2(.dout(w_dff_A_h8mlJ5ry7_2),.din(w_dff_A_G5zBqwwm1_2),.clk(gclk));
	jdff dff_B_1EgBCTye7_0(.din(n695),.dout(w_dff_B_1EgBCTye7_0),.clk(gclk));
	jdff dff_B_cLKal65A0_1(.din(n676),.dout(w_dff_B_cLKal65A0_1),.clk(gclk));
	jdff dff_A_dhh6kTWW6_1(.dout(w_n693_0[1]),.din(w_dff_A_dhh6kTWW6_1),.clk(gclk));
	jdff dff_A_xtYlC6vM0_1(.dout(w_n691_0[1]),.din(w_dff_A_xtYlC6vM0_1),.clk(gclk));
	jdff dff_A_yUFvQGBe4_1(.dout(w_dff_A_xtYlC6vM0_1),.din(w_dff_A_yUFvQGBe4_1),.clk(gclk));
	jdff dff_A_kiTgCdMK9_0(.dout(w_n687_0[0]),.din(w_dff_A_kiTgCdMK9_0),.clk(gclk));
	jdff dff_A_ns7p0HW69_1(.dout(w_n687_0[1]),.din(w_dff_A_ns7p0HW69_1),.clk(gclk));
	jdff dff_A_tub42awF6_1(.dout(w_dff_A_ns7p0HW69_1),.din(w_dff_A_tub42awF6_1),.clk(gclk));
	jdff dff_A_yPXAgVCv6_1(.dout(w_dff_A_tub42awF6_1),.din(w_dff_A_yPXAgVCv6_1),.clk(gclk));
	jdff dff_A_qh2rtEy50_1(.dout(w_dff_A_yPXAgVCv6_1),.din(w_dff_A_qh2rtEy50_1),.clk(gclk));
	jdff dff_B_Q9etFRNv5_0(.din(n685),.dout(w_dff_B_Q9etFRNv5_0),.clk(gclk));
	jdff dff_A_KhdVihu96_2(.dout(w_n571_0[2]),.din(w_dff_A_KhdVihu96_2),.clk(gclk));
	jdff dff_A_jVOsbSPk5_2(.dout(w_dff_A_KhdVihu96_2),.din(w_dff_A_jVOsbSPk5_2),.clk(gclk));
	jdff dff_A_TzhCfWqV9_2(.dout(w_dff_A_jVOsbSPk5_2),.din(w_dff_A_TzhCfWqV9_2),.clk(gclk));
	jdff dff_A_p5UUECnV1_1(.dout(w_n569_0[1]),.din(w_dff_A_p5UUECnV1_1),.clk(gclk));
	jdff dff_A_ukhumN2q9_1(.dout(w_G280_0[1]),.din(w_dff_A_ukhumN2q9_1),.clk(gclk));
	jdff dff_A_1sgg50Vh5_0(.dout(w_n681_2[0]),.din(w_dff_A_1sgg50Vh5_0),.clk(gclk));
	jdff dff_A_FjXNNgSc6_0(.dout(w_dff_A_1sgg50Vh5_0),.din(w_dff_A_FjXNNgSc6_0),.clk(gclk));
	jdff dff_A_u58kNjAx0_0(.dout(w_n681_0[0]),.din(w_dff_A_u58kNjAx0_0),.clk(gclk));
	jdff dff_A_ejRfFmEt0_1(.dout(w_n681_0[1]),.din(w_dff_A_ejRfFmEt0_1),.clk(gclk));
	jdff dff_A_dN1kmbjE3_1(.dout(w_n680_0[1]),.din(w_dff_A_dN1kmbjE3_1),.clk(gclk));
	jdff dff_A_aMAMcnaI2_1(.dout(w_n679_0[1]),.din(w_dff_A_aMAMcnaI2_1),.clk(gclk));
	jdff dff_A_OWasprSn8_1(.dout(w_n678_0[1]),.din(w_dff_A_OWasprSn8_1),.clk(gclk));
	jdff dff_B_e8L57UDN4_1(.din(n557),.dout(w_dff_B_e8L57UDN4_1),.clk(gclk));
	jdff dff_B_aLPQmUoB9_1(.din(w_dff_B_e8L57UDN4_1),.dout(w_dff_B_aLPQmUoB9_1),.clk(gclk));
	jdff dff_B_KBLk7vCb4_1(.din(G241),.dout(w_dff_B_KBLk7vCb4_1),.clk(gclk));
	jdff dff_B_JVOrBYxW0_2(.din(n1543),.dout(w_dff_B_JVOrBYxW0_2),.clk(gclk));
	jdff dff_B_fNYVBgIL5_2(.din(w_dff_B_JVOrBYxW0_2),.dout(w_dff_B_fNYVBgIL5_2),.clk(gclk));
	jdff dff_B_Y6TYRwuO0_2(.din(w_dff_B_fNYVBgIL5_2),.dout(w_dff_B_Y6TYRwuO0_2),.clk(gclk));
	jdff dff_B_JiSN9Gy68_2(.din(w_dff_B_Y6TYRwuO0_2),.dout(w_dff_B_JiSN9Gy68_2),.clk(gclk));
	jdff dff_B_xUG6aHmB6_2(.din(w_dff_B_JiSN9Gy68_2),.dout(w_dff_B_xUG6aHmB6_2),.clk(gclk));
	jdff dff_B_vtY4jYEU8_2(.din(w_dff_B_xUG6aHmB6_2),.dout(w_dff_B_vtY4jYEU8_2),.clk(gclk));
	jdff dff_B_hPZshaVc0_2(.din(w_dff_B_vtY4jYEU8_2),.dout(w_dff_B_hPZshaVc0_2),.clk(gclk));
	jdff dff_A_f79kWhbe5_2(.dout(w_n583_0[2]),.din(w_dff_A_f79kWhbe5_2),.clk(gclk));
	jdff dff_A_pWeJZXtu1_2(.dout(w_dff_A_f79kWhbe5_2),.din(w_dff_A_pWeJZXtu1_2),.clk(gclk));
	jdff dff_A_bRfgWAj95_2(.dout(w_dff_A_pWeJZXtu1_2),.din(w_dff_A_bRfgWAj95_2),.clk(gclk));
	jdff dff_A_Yf2qE8Lp4_2(.dout(w_dff_A_bRfgWAj95_2),.din(w_dff_A_Yf2qE8Lp4_2),.clk(gclk));
	jdff dff_A_tIC1BynL9_1(.dout(w_n578_0[1]),.din(w_dff_A_tIC1BynL9_1),.clk(gclk));
	jdff dff_A_i76LOC2U0_1(.dout(w_dff_A_tIC1BynL9_1),.din(w_dff_A_i76LOC2U0_1),.clk(gclk));
	jdff dff_A_1Ub2jJXa3_1(.dout(w_dff_A_i76LOC2U0_1),.din(w_dff_A_1Ub2jJXa3_1),.clk(gclk));
	jdff dff_A_QykfMVeT2_1(.dout(w_dff_A_1Ub2jJXa3_1),.din(w_dff_A_QykfMVeT2_1),.clk(gclk));
	jdff dff_A_3ADiFjjj6_1(.dout(w_dff_A_QykfMVeT2_1),.din(w_dff_A_3ADiFjjj6_1),.clk(gclk));
	jdff dff_A_Vqq2KzBu3_1(.dout(w_dff_A_3ADiFjjj6_1),.din(w_dff_A_Vqq2KzBu3_1),.clk(gclk));
	jdff dff_B_pJf8iC144_0(.din(n576),.dout(w_dff_B_pJf8iC144_0),.clk(gclk));
	jdff dff_A_Osos0htW4_0(.dout(w_G335_3[0]),.din(w_dff_A_Osos0htW4_0),.clk(gclk));
	jdff dff_B_tcW54GU74_1(.din(G264),.dout(w_dff_B_tcW54GU74_1),.clk(gclk));
	jdff dff_A_p4y39Lw87_0(.dout(w_n473_1[0]),.din(w_dff_A_p4y39Lw87_0),.clk(gclk));
	jdff dff_A_vLeUpb2s1_1(.dout(w_n943_0[1]),.din(w_dff_A_vLeUpb2s1_1),.clk(gclk));
	jdff dff_A_9qwxkvpO9_1(.dout(w_dff_A_vLeUpb2s1_1),.din(w_dff_A_9qwxkvpO9_1),.clk(gclk));
	jdff dff_A_WSYdpcS13_1(.dout(w_dff_A_9qwxkvpO9_1),.din(w_dff_A_WSYdpcS13_1),.clk(gclk));
	jdff dff_A_clTPiQcX1_1(.dout(w_dff_A_WSYdpcS13_1),.din(w_dff_A_clTPiQcX1_1),.clk(gclk));
	jdff dff_A_6tWZHaJc8_1(.dout(w_dff_A_clTPiQcX1_1),.din(w_dff_A_6tWZHaJc8_1),.clk(gclk));
	jdff dff_A_KEeEvvGT0_1(.dout(w_dff_A_6tWZHaJc8_1),.din(w_dff_A_KEeEvvGT0_1),.clk(gclk));
	jdff dff_A_sk2iuow46_1(.dout(w_dff_A_KEeEvvGT0_1),.din(w_dff_A_sk2iuow46_1),.clk(gclk));
	jdff dff_A_c8k55u2I4_1(.dout(w_n591_0[1]),.din(w_dff_A_c8k55u2I4_1),.clk(gclk));
	jdff dff_A_ivFqTZDA0_1(.dout(w_dff_A_c8k55u2I4_1),.din(w_dff_A_ivFqTZDA0_1),.clk(gclk));
	jdff dff_A_vCI94uB73_1(.dout(w_n590_0[1]),.din(w_dff_A_vCI94uB73_1),.clk(gclk));
	jdff dff_A_zWJzag0i3_1(.dout(w_dff_A_vCI94uB73_1),.din(w_dff_A_zWJzag0i3_1),.clk(gclk));
	jdff dff_B_FFemuDfY4_0(.din(n589),.dout(w_dff_B_FFemuDfY4_0),.clk(gclk));
	jdff dff_B_BES1QqrZ5_1(.din(G217),.dout(w_dff_B_BES1QqrZ5_1),.clk(gclk));
	jdff dff_A_yd3URyCi7_0(.dout(w_G335_4[0]),.din(w_dff_A_yd3URyCi7_0),.clk(gclk));
	jdff dff_A_bjbwUG7M0_2(.dout(w_G335_1[2]),.din(w_dff_A_bjbwUG7M0_2),.clk(gclk));
	jdff dff_B_fZBBz8PT9_0(.din(n1537),.dout(w_dff_B_fZBBz8PT9_0),.clk(gclk));
	jdff dff_A_wUBAaK9o5_1(.dout(w_n750_0[1]),.din(w_dff_A_wUBAaK9o5_1),.clk(gclk));
	jdff dff_A_IRGXz4DO5_1(.dout(w_dff_A_wUBAaK9o5_1),.din(w_dff_A_IRGXz4DO5_1),.clk(gclk));
	jdff dff_A_99mLvw3T2_1(.dout(w_dff_A_IRGXz4DO5_1),.din(w_dff_A_99mLvw3T2_1),.clk(gclk));
	jdff dff_A_yfizk2VW9_1(.dout(w_dff_A_99mLvw3T2_1),.din(w_dff_A_yfizk2VW9_1),.clk(gclk));
	jdff dff_A_0tA7cmZF9_1(.dout(w_dff_A_yfizk2VW9_1),.din(w_dff_A_0tA7cmZF9_1),.clk(gclk));
	jdff dff_A_rUUA4veq5_1(.dout(w_dff_A_0tA7cmZF9_1),.din(w_dff_A_rUUA4veq5_1),.clk(gclk));
	jdff dff_A_3iL3Rmpg0_1(.dout(w_dff_A_rUUA4veq5_1),.din(w_dff_A_3iL3Rmpg0_1),.clk(gclk));
	jdff dff_A_sl7mnM717_1(.dout(w_dff_A_3iL3Rmpg0_1),.din(w_dff_A_sl7mnM717_1),.clk(gclk));
	jdff dff_A_klDAUInG2_1(.dout(w_dff_A_sl7mnM717_1),.din(w_dff_A_klDAUInG2_1),.clk(gclk));
	jdff dff_A_9CJp5tTw1_1(.dout(w_dff_A_klDAUInG2_1),.din(w_dff_A_9CJp5tTw1_1),.clk(gclk));
	jdff dff_A_ABuFr46p9_1(.dout(w_dff_A_9CJp5tTw1_1),.din(w_dff_A_ABuFr46p9_1),.clk(gclk));
	jdff dff_A_9MIa6QAY4_2(.dout(w_n750_0[2]),.din(w_dff_A_9MIa6QAY4_2),.clk(gclk));
	jdff dff_A_xYW9Q1cW3_2(.dout(w_dff_A_9MIa6QAY4_2),.din(w_dff_A_xYW9Q1cW3_2),.clk(gclk));
	jdff dff_A_w7fSKZSl7_2(.dout(w_dff_A_xYW9Q1cW3_2),.din(w_dff_A_w7fSKZSl7_2),.clk(gclk));
	jdff dff_A_wp8DNQnT5_2(.dout(w_dff_A_w7fSKZSl7_2),.din(w_dff_A_wp8DNQnT5_2),.clk(gclk));
	jdff dff_A_Lsd8e2ir4_2(.dout(w_dff_A_wp8DNQnT5_2),.din(w_dff_A_Lsd8e2ir4_2),.clk(gclk));
	jdff dff_A_vKBiK2D37_2(.dout(w_G4091_2[2]),.din(w_dff_A_vKBiK2D37_2),.clk(gclk));
	jdff dff_A_YIaTwVTq4_2(.dout(w_G4091_0[2]),.din(w_dff_A_YIaTwVTq4_2),.clk(gclk));
	jdff dff_A_H6bIqRMJ3_2(.dout(w_dff_A_YIaTwVTq4_2),.din(w_dff_A_H6bIqRMJ3_2),.clk(gclk));
	jdff dff_A_OXVi1ln21_2(.dout(w_dff_A_H6bIqRMJ3_2),.din(w_dff_A_OXVi1ln21_2),.clk(gclk));
	jdff dff_A_1YgcUGKM0_2(.dout(w_dff_A_OXVi1ln21_2),.din(w_dff_A_1YgcUGKM0_2),.clk(gclk));
	jdff dff_A_LEkVKVBX8_2(.dout(w_dff_A_1YgcUGKM0_2),.din(w_dff_A_LEkVKVBX8_2),.clk(gclk));
	jdff dff_A_aLyJPXB60_2(.dout(w_dff_A_LEkVKVBX8_2),.din(w_dff_A_aLyJPXB60_2),.clk(gclk));
	jdff dff_A_1WXVIlvZ0_2(.dout(w_dff_A_aLyJPXB60_2),.din(w_dff_A_1WXVIlvZ0_2),.clk(gclk));
	jdff dff_A_5aFFldOM1_2(.dout(w_dff_A_1WXVIlvZ0_2),.din(w_dff_A_5aFFldOM1_2),.clk(gclk));
	jdff dff_A_lYniwzhv0_2(.dout(w_dff_A_5aFFldOM1_2),.din(w_dff_A_lYniwzhv0_2),.clk(gclk));
	jdff dff_A_0WzQkEuT8_2(.dout(w_dff_A_lYniwzhv0_2),.din(w_dff_A_0WzQkEuT8_2),.clk(gclk));
	jdff dff_A_6AbCe3U21_2(.dout(w_dff_A_0WzQkEuT8_2),.din(w_dff_A_6AbCe3U21_2),.clk(gclk));
	jdff dff_A_yBX3zBhB4_2(.dout(w_dff_A_6AbCe3U21_2),.din(w_dff_A_yBX3zBhB4_2),.clk(gclk));
	jdff dff_A_LQkLYlbU9_2(.dout(w_dff_A_yBX3zBhB4_2),.din(w_dff_A_LQkLYlbU9_2),.clk(gclk));
	jdff dff_B_MCAgvn5H2_2(.din(n1533),.dout(w_dff_B_MCAgvn5H2_2),.clk(gclk));
	jdff dff_B_nuDczt3V7_0(.din(n1525),.dout(w_dff_B_nuDczt3V7_0),.clk(gclk));
	jdff dff_A_LAvEutKN7_0(.dout(w_n486_0[0]),.din(w_dff_A_LAvEutKN7_0),.clk(gclk));
	jdff dff_A_t4Wy8jsh4_2(.dout(w_n486_0[2]),.din(w_dff_A_t4Wy8jsh4_2),.clk(gclk));
	jdff dff_A_lofmVhhj3_0(.dout(w_G411_0[0]),.din(w_dff_A_lofmVhhj3_0),.clk(gclk));
	jdff dff_A_7sr0iuu30_0(.dout(w_dff_A_lofmVhhj3_0),.din(w_dff_A_7sr0iuu30_0),.clk(gclk));
	jdff dff_A_1Hs6LHY27_1(.dout(w_G411_0[1]),.din(w_dff_A_1Hs6LHY27_1),.clk(gclk));
	jdff dff_A_Fsw5FWWf3_1(.dout(w_G273_2[1]),.din(w_dff_A_Fsw5FWWf3_1),.clk(gclk));
	jdff dff_A_oG5mlAkU3_2(.dout(w_G273_0[2]),.din(w_dff_A_oG5mlAkU3_2),.clk(gclk));
	jdff dff_B_QpVmftZ76_1(.din(n1518),.dout(w_dff_B_QpVmftZ76_1),.clk(gclk));
	jdff dff_B_gegiqUQb2_1(.din(w_dff_B_QpVmftZ76_1),.dout(w_dff_B_gegiqUQb2_1),.clk(gclk));
	jdff dff_A_hd0J9uOv7_0(.dout(w_n473_0[0]),.din(w_dff_A_hd0J9uOv7_0),.clk(gclk));
	jdff dff_A_mYCOLQWJ5_2(.dout(w_n473_0[2]),.din(w_dff_A_mYCOLQWJ5_2),.clk(gclk));
	jdff dff_A_Cds4j2RZ3_2(.dout(w_dff_A_mYCOLQWJ5_2),.din(w_dff_A_Cds4j2RZ3_2),.clk(gclk));
	jdff dff_B_qAzlFbbr0_1(.din(n1514),.dout(w_dff_B_qAzlFbbr0_1),.clk(gclk));
	jdff dff_A_itVy6ivB7_1(.dout(w_G257_2[1]),.din(w_dff_A_itVy6ivB7_1),.clk(gclk));
	jdff dff_A_dVCXe1m09_0(.dout(w_G389_0[0]),.din(w_dff_A_dVCXe1m09_0),.clk(gclk));
	jdff dff_A_bMCTS3lh5_1(.dout(w_G389_0[1]),.din(w_dff_A_bMCTS3lh5_1),.clk(gclk));
	jdff dff_A_uLwLcYkQ5_0(.dout(w_G257_1[0]),.din(w_dff_A_uLwLcYkQ5_0),.clk(gclk));
	jdff dff_B_c7KuWy6q2_0(.din(n1506),.dout(w_dff_B_c7KuWy6q2_0),.clk(gclk));
	jdff dff_A_aX7Q3r0A3_0(.dout(w_n451_0[0]),.din(w_dff_A_aX7Q3r0A3_0),.clk(gclk));
	jdff dff_A_SIaOqvhL3_2(.dout(w_n451_0[2]),.din(w_dff_A_SIaOqvhL3_2),.clk(gclk));
	jdff dff_A_TIbKSzWp7_0(.dout(w_G400_1[0]),.din(w_dff_A_TIbKSzWp7_0),.clk(gclk));
	jdff dff_A_BDi6pTbm8_1(.dout(w_G400_0[1]),.din(w_dff_A_BDi6pTbm8_1),.clk(gclk));
	jdff dff_A_6BxukAJX7_1(.dout(w_dff_A_BDi6pTbm8_1),.din(w_dff_A_6BxukAJX7_1),.clk(gclk));
	jdff dff_A_Dkuju8IF0_2(.dout(w_G400_0[2]),.din(w_dff_A_Dkuju8IF0_2),.clk(gclk));
	jdff dff_A_2ZmmhUZk7_2(.dout(w_dff_A_Dkuju8IF0_2),.din(w_dff_A_2ZmmhUZk7_2),.clk(gclk));
	jdff dff_A_nh5h3Tpz4_0(.dout(w_G265_2[0]),.din(w_dff_A_nh5h3Tpz4_0),.clk(gclk));
	jdff dff_A_HsHNtB4R8_2(.dout(w_G265_0[2]),.din(w_dff_A_HsHNtB4R8_2),.clk(gclk));
	jdff dff_B_bIs2Ifyb2_0(.din(n1497),.dout(w_dff_B_bIs2Ifyb2_0),.clk(gclk));
	jdff dff_A_Gyr6Xdi39_0(.dout(w_n497_0[0]),.din(w_dff_A_Gyr6Xdi39_0),.clk(gclk));
	jdff dff_A_rUqn3KEZ1_2(.dout(w_n497_0[2]),.din(w_dff_A_rUqn3KEZ1_2),.clk(gclk));
	jdff dff_A_ywFPaaCB1_0(.dout(w_G374_0[0]),.din(w_dff_A_ywFPaaCB1_0),.clk(gclk));
	jdff dff_A_DU9og2s62_0(.dout(w_dff_A_ywFPaaCB1_0),.din(w_dff_A_DU9og2s62_0),.clk(gclk));
	jdff dff_A_IFGuyCP12_1(.dout(w_G374_0[1]),.din(w_dff_A_IFGuyCP12_1),.clk(gclk));
	jdff dff_A_x9Mga5Vo5_0(.dout(w_G281_2[0]),.din(w_dff_A_x9Mga5Vo5_0),.clk(gclk));
	jdff dff_A_92zf0YJc9_2(.dout(w_G281_0[2]),.din(w_dff_A_92zf0YJc9_2),.clk(gclk));
	jdff dff_B_qxKn9S912_1(.din(n1463),.dout(w_dff_B_qxKn9S912_1),.clk(gclk));
	jdff dff_B_1gVAaMPB9_1(.din(w_dff_B_qxKn9S912_1),.dout(w_dff_B_1gVAaMPB9_1),.clk(gclk));
	jdff dff_B_4jxE2WRh1_0(.din(n1485),.dout(w_dff_B_4jxE2WRh1_0),.clk(gclk));
	jdff dff_A_LRGG1Bdy9_1(.dout(w_G210_1[1]),.din(w_dff_A_LRGG1Bdy9_1),.clk(gclk));
	jdff dff_A_rQBGozHr8_1(.dout(w_n543_0[1]),.din(w_dff_A_rQBGozHr8_1),.clk(gclk));
	jdff dff_A_UjyjVKCa7_0(.dout(w_G457_2[0]),.din(w_dff_A_UjyjVKCa7_0),.clk(gclk));
	jdff dff_A_t7kWPFrr4_0(.dout(w_G457_0[0]),.din(w_dff_A_t7kWPFrr4_0),.clk(gclk));
	jdff dff_A_FTBFJaf07_0(.dout(w_dff_A_t7kWPFrr4_0),.din(w_dff_A_FTBFJaf07_0),.clk(gclk));
	jdff dff_A_am9HuM5N3_2(.dout(w_G457_0[2]),.din(w_dff_A_am9HuM5N3_2),.clk(gclk));
	jdff dff_A_XdkzTyra1_2(.dout(w_dff_A_am9HuM5N3_2),.din(w_dff_A_XdkzTyra1_2),.clk(gclk));
	jdff dff_A_oO8qcMEs4_1(.dout(w_G210_2[1]),.din(w_dff_A_oO8qcMEs4_1),.clk(gclk));
	jdff dff_A_dBgxT8vC6_2(.dout(w_G210_0[2]),.din(w_dff_A_dBgxT8vC6_2),.clk(gclk));
	jdff dff_B_UWRsh97v6_1(.din(n1478),.dout(w_dff_B_UWRsh97v6_1),.clk(gclk));
	jdff dff_B_ufvP6d3X3_1(.din(w_dff_B_UWRsh97v6_1),.dout(w_dff_B_ufvP6d3X3_1),.clk(gclk));
	jdff dff_A_kGhS7hCR3_1(.dout(w_n509_0[1]),.din(w_dff_A_kGhS7hCR3_1),.clk(gclk));
	jdff dff_A_OYzD7mj43_0(.dout(w_G468_1[0]),.din(w_dff_A_OYzD7mj43_0),.clk(gclk));
	jdff dff_A_vXbNci8I3_0(.dout(w_dff_A_OYzD7mj43_0),.din(w_dff_A_vXbNci8I3_0),.clk(gclk));
	jdff dff_A_Rwtbp0hX3_1(.dout(w_G468_1[1]),.din(w_dff_A_Rwtbp0hX3_1),.clk(gclk));
	jdff dff_B_rPkfXDut9_1(.din(n1474),.dout(w_dff_B_rPkfXDut9_1),.clk(gclk));
	jdff dff_A_7GTAHaeJ5_1(.dout(w_G218_2[1]),.din(w_dff_A_7GTAHaeJ5_1),.clk(gclk));
	jdff dff_A_jHQrua3D1_1(.dout(w_G468_0[1]),.din(w_dff_A_jHQrua3D1_1),.clk(gclk));
	jdff dff_A_pyWdyymZ4_2(.dout(w_G468_0[2]),.din(w_dff_A_pyWdyymZ4_2),.clk(gclk));
	jdff dff_A_Arb3f7to5_2(.dout(w_dff_A_pyWdyymZ4_2),.din(w_dff_A_Arb3f7to5_2),.clk(gclk));
	jdff dff_A_aMxlNGir1_0(.dout(w_G218_1[0]),.din(w_dff_A_aMxlNGir1_0),.clk(gclk));
	jdff dff_B_Wl0mEALJ0_1(.din(n1468),.dout(w_dff_B_Wl0mEALJ0_1),.clk(gclk));
	jdff dff_B_weVoAiYu5_1(.din(w_dff_B_Wl0mEALJ0_1),.dout(w_dff_B_weVoAiYu5_1),.clk(gclk));
	jdff dff_A_5h5lW8da8_1(.dout(w_n532_0[1]),.din(w_dff_A_5h5lW8da8_1),.clk(gclk));
	jdff dff_A_VqUJsa6V0_0(.dout(w_G422_2[0]),.din(w_dff_A_VqUJsa6V0_0),.clk(gclk));
	jdff dff_B_P4UFu9w18_1(.din(n1464),.dout(w_dff_B_P4UFu9w18_1),.clk(gclk));
	jdff dff_A_an3LtqQN4_1(.dout(w_G226_2[1]),.din(w_dff_A_an3LtqQN4_1),.clk(gclk));
	jdff dff_A_QTvnrDK57_0(.dout(w_G422_0[0]),.din(w_dff_A_QTvnrDK57_0),.clk(gclk));
	jdff dff_A_G3VvcAxt0_0(.dout(w_dff_A_QTvnrDK57_0),.din(w_dff_A_G3VvcAxt0_0),.clk(gclk));
	jdff dff_A_IKwuN2PV3_2(.dout(w_G422_0[2]),.din(w_dff_A_IKwuN2PV3_2),.clk(gclk));
	jdff dff_A_wyHVClMG1_1(.dout(w_G251_4[1]),.din(w_dff_A_wyHVClMG1_1),.clk(gclk));
	jdff dff_A_mssGpBpw2_2(.dout(w_G251_4[2]),.din(w_dff_A_mssGpBpw2_2),.clk(gclk));
	jdff dff_A_A6waiVFy5_1(.dout(w_G251_1[1]),.din(w_dff_A_A6waiVFy5_1),.clk(gclk));
	jdff dff_A_KqWzSVqx9_2(.dout(w_G251_1[2]),.din(w_dff_A_KqWzSVqx9_2),.clk(gclk));
	jdff dff_A_DvF0fMCl5_0(.dout(w_G226_1[0]),.din(w_dff_A_DvF0fMCl5_0),.clk(gclk));
	jdff dff_B_BcV4qtdl5_0(.din(n522),.dout(w_dff_B_BcV4qtdl5_0),.clk(gclk));
	jdff dff_A_Hu0gcDYA1_0(.dout(w_G446_1[0]),.din(w_dff_A_Hu0gcDYA1_0),.clk(gclk));
	jdff dff_A_jgz4A8ZC0_0(.dout(w_dff_A_Hu0gcDYA1_0),.din(w_dff_A_jgz4A8ZC0_0),.clk(gclk));
	jdff dff_A_GOsOZ2FX8_0(.dout(w_dff_A_jgz4A8ZC0_0),.din(w_dff_A_GOsOZ2FX8_0),.clk(gclk));
	jdff dff_A_8flNOkE21_0(.dout(w_dff_A_GOsOZ2FX8_0),.din(w_dff_A_8flNOkE21_0),.clk(gclk));
	jdff dff_A_JRghSMkZ4_1(.dout(w_G446_1[1]),.din(w_dff_A_JRghSMkZ4_1),.clk(gclk));
	jdff dff_A_iKiEC3sc5_1(.dout(w_dff_A_JRghSMkZ4_1),.din(w_dff_A_iKiEC3sc5_1),.clk(gclk));
	jdff dff_A_iaeHegeY5_1(.dout(w_G446_0[1]),.din(w_dff_A_iaeHegeY5_1),.clk(gclk));
	jdff dff_A_bmLrmGfX2_1(.dout(w_dff_A_iaeHegeY5_1),.din(w_dff_A_bmLrmGfX2_1),.clk(gclk));
	jdff dff_A_Tp4monOj8_1(.dout(w_dff_A_bmLrmGfX2_1),.din(w_dff_A_Tp4monOj8_1),.clk(gclk));
	jdff dff_A_oi8BN86S2_1(.dout(w_dff_A_Tp4monOj8_1),.din(w_dff_A_oi8BN86S2_1),.clk(gclk));
	jdff dff_A_UaTz9xX71_2(.dout(w_G446_0[2]),.din(w_dff_A_UaTz9xX71_2),.clk(gclk));
	jdff dff_A_akMWDiC57_2(.dout(w_dff_A_UaTz9xX71_2),.din(w_dff_A_akMWDiC57_2),.clk(gclk));
	jdff dff_A_DG9GqePC8_2(.dout(w_dff_A_akMWDiC57_2),.din(w_dff_A_DG9GqePC8_2),.clk(gclk));
	jdff dff_A_kfmutEPO3_2(.dout(w_dff_A_DG9GqePC8_2),.din(w_dff_A_kfmutEPO3_2),.clk(gclk));
	jdff dff_A_27FkoB2q8_0(.dout(w_G206_0[0]),.din(w_dff_A_27FkoB2q8_0),.clk(gclk));
	jdff dff_A_qoxOJcP88_0(.dout(w_G242_1[0]),.din(w_dff_A_qoxOJcP88_0),.clk(gclk));
	jdff dff_A_hmdwoiRC5_1(.dout(w_G242_1[1]),.din(w_dff_A_hmdwoiRC5_1),.clk(gclk));
	jdff dff_A_eq9gA4NK7_1(.dout(w_G242_0[1]),.din(w_dff_A_eq9gA4NK7_1),.clk(gclk));
	jdff dff_A_uf7O1jrH4_2(.dout(w_G242_0[2]),.din(w_dff_A_uf7O1jrH4_2),.clk(gclk));
	jdff dff_B_EYGPxgol6_0(.din(n1457),.dout(w_dff_B_EYGPxgol6_0),.clk(gclk));
	jdff dff_A_yj6NuqGK2_2(.dout(w_G248_3[2]),.din(w_dff_A_yj6NuqGK2_2),.clk(gclk));
	jdff dff_A_ZQjdUpdm1_1(.dout(w_n462_0[1]),.din(w_dff_A_ZQjdUpdm1_1),.clk(gclk));
	jdff dff_A_2qaOPaK74_1(.dout(w_dff_A_ZQjdUpdm1_1),.din(w_dff_A_2qaOPaK74_1),.clk(gclk));
	jdff dff_A_r5cUzes00_1(.dout(w_dff_A_2qaOPaK74_1),.din(w_dff_A_r5cUzes00_1),.clk(gclk));
	jdff dff_A_cXlOgeUS3_1(.dout(w_dff_A_r5cUzes00_1),.din(w_dff_A_cXlOgeUS3_1),.clk(gclk));
	jdff dff_A_tzs6aVif1_2(.dout(w_n462_0[2]),.din(w_dff_A_tzs6aVif1_2),.clk(gclk));
	jdff dff_A_ynQu8YKB0_0(.dout(w_G435_1[0]),.din(w_dff_A_ynQu8YKB0_0),.clk(gclk));
	jdff dff_A_VdwvlNOa8_0(.dout(w_dff_A_ynQu8YKB0_0),.din(w_dff_A_VdwvlNOa8_0),.clk(gclk));
	jdff dff_A_fSkY3zGm9_0(.dout(w_dff_A_VdwvlNOa8_0),.din(w_dff_A_fSkY3zGm9_0),.clk(gclk));
	jdff dff_A_olwED41o7_0(.dout(w_dff_A_fSkY3zGm9_0),.din(w_dff_A_olwED41o7_0),.clk(gclk));
	jdff dff_A_42D1ZSQZ3_1(.dout(w_G435_1[1]),.din(w_dff_A_42D1ZSQZ3_1),.clk(gclk));
	jdff dff_A_68LXjsIP1_1(.dout(w_G435_0[1]),.din(w_dff_A_68LXjsIP1_1),.clk(gclk));
	jdff dff_A_35cJy9Fu7_1(.dout(w_dff_A_68LXjsIP1_1),.din(w_dff_A_35cJy9Fu7_1),.clk(gclk));
	jdff dff_A_ZF4JHgGb1_2(.dout(w_G435_0[2]),.din(w_dff_A_ZF4JHgGb1_2),.clk(gclk));
	jdff dff_A_hXTgRgpi5_2(.dout(w_dff_A_ZF4JHgGb1_2),.din(w_dff_A_hXTgRgpi5_2),.clk(gclk));
	jdff dff_A_QQpdEMIz9_2(.dout(w_dff_A_hXTgRgpi5_2),.din(w_dff_A_QQpdEMIz9_2),.clk(gclk));
	jdff dff_A_bVfatrKy2_2(.dout(w_dff_A_QQpdEMIz9_2),.din(w_dff_A_bVfatrKy2_2),.clk(gclk));
	jdff dff_A_mImFSVqW2_1(.dout(w_G251_0[1]),.din(w_dff_A_mImFSVqW2_1),.clk(gclk));
	jdff dff_A_GOTqrNDj2_2(.dout(w_G251_0[2]),.din(w_dff_A_GOTqrNDj2_2),.clk(gclk));
	jdff dff_A_Qzss2TnV3_0(.dout(w_G234_2[0]),.din(w_dff_A_Qzss2TnV3_0),.clk(gclk));
	jdff dff_A_B2BOyBS42_2(.dout(w_G234_0[2]),.din(w_dff_A_B2BOyBS42_2),.clk(gclk));
	jdff dff_A_h6Bje0u85_0(.dout(w_G4092_1[0]),.din(w_dff_A_h6Bje0u85_0),.clk(gclk));
	jdff dff_A_8dtHPSLt3_0(.dout(w_dff_A_h6Bje0u85_0),.din(w_dff_A_8dtHPSLt3_0),.clk(gclk));
	jdff dff_A_0IBeB7vB8_0(.dout(w_dff_A_8dtHPSLt3_0),.din(w_dff_A_0IBeB7vB8_0),.clk(gclk));
	jdff dff_A_menPV4hY9_0(.dout(w_dff_A_0IBeB7vB8_0),.din(w_dff_A_menPV4hY9_0),.clk(gclk));
	jdff dff_A_qoCehplD0_0(.dout(w_dff_A_menPV4hY9_0),.din(w_dff_A_qoCehplD0_0),.clk(gclk));
	jdff dff_A_yJIV1UTL6_0(.dout(w_dff_A_qoCehplD0_0),.din(w_dff_A_yJIV1UTL6_0),.clk(gclk));
	jdff dff_A_DCktl07W6_0(.dout(w_dff_A_yJIV1UTL6_0),.din(w_dff_A_DCktl07W6_0),.clk(gclk));
	jdff dff_A_PqJjzx568_0(.dout(w_dff_A_DCktl07W6_0),.din(w_dff_A_PqJjzx568_0),.clk(gclk));
	jdff dff_A_Tka5TvuH0_0(.dout(w_dff_A_PqJjzx568_0),.din(w_dff_A_Tka5TvuH0_0),.clk(gclk));
	jdff dff_A_rRft9HIC6_1(.dout(w_G4092_1[1]),.din(w_dff_A_rRft9HIC6_1),.clk(gclk));
	jdff dff_A_jrDNxaWR0_0(.dout(w_n999_1[0]),.din(w_dff_A_jrDNxaWR0_0),.clk(gclk));
	jdff dff_A_pWVrn1Ru0_0(.dout(w_dff_A_jrDNxaWR0_0),.din(w_dff_A_pWVrn1Ru0_0),.clk(gclk));
	jdff dff_A_SqyQK0Um1_0(.dout(w_dff_A_pWVrn1Ru0_0),.din(w_dff_A_SqyQK0Um1_0),.clk(gclk));
	jdff dff_A_YaQijCGJ1_0(.dout(w_dff_A_SqyQK0Um1_0),.din(w_dff_A_YaQijCGJ1_0),.clk(gclk));
	jdff dff_A_xhZzeUGE6_0(.dout(w_dff_A_YaQijCGJ1_0),.din(w_dff_A_xhZzeUGE6_0),.clk(gclk));
	jdff dff_A_C7kY2QMG8_0(.dout(w_dff_A_xhZzeUGE6_0),.din(w_dff_A_C7kY2QMG8_0),.clk(gclk));
	jdff dff_A_GTWccmwW1_2(.dout(w_n999_1[2]),.din(w_dff_A_GTWccmwW1_2),.clk(gclk));
	jdff dff_A_SRr5tQVE7_2(.dout(w_dff_A_GTWccmwW1_2),.din(w_dff_A_SRr5tQVE7_2),.clk(gclk));
	jdff dff_A_KzBGOplm6_2(.dout(w_dff_A_SRr5tQVE7_2),.din(w_dff_A_KzBGOplm6_2),.clk(gclk));
	jdff dff_A_XEBab9VM6_2(.dout(w_dff_A_KzBGOplm6_2),.din(w_dff_A_XEBab9VM6_2),.clk(gclk));
	jdff dff_A_ZPP8Z6Ok2_2(.dout(w_dff_A_XEBab9VM6_2),.din(w_dff_A_ZPP8Z6Ok2_2),.clk(gclk));
	jdff dff_A_wOz1qlpK5_2(.dout(w_dff_A_ZPP8Z6Ok2_2),.din(w_dff_A_wOz1qlpK5_2),.clk(gclk));
	jdff dff_A_68Ycn3WV1_2(.dout(w_dff_A_wOz1qlpK5_2),.din(w_dff_A_68Ycn3WV1_2),.clk(gclk));
	jdff dff_A_oekBM2LI9_2(.dout(w_dff_A_68Ycn3WV1_2),.din(w_dff_A_oekBM2LI9_2),.clk(gclk));
	jdff dff_A_NMinA4VU9_2(.dout(w_dff_A_oekBM2LI9_2),.din(w_dff_A_NMinA4VU9_2),.clk(gclk));
	jdff dff_A_hzACrLF68_2(.dout(w_dff_A_NMinA4VU9_2),.din(w_dff_A_hzACrLF68_2),.clk(gclk));
	jdff dff_A_BW1HhNof2_2(.dout(w_dff_A_hzACrLF68_2),.din(w_dff_A_BW1HhNof2_2),.clk(gclk));
	jdff dff_A_2vzhdSBC8_1(.dout(w_n999_0[1]),.din(w_dff_A_2vzhdSBC8_1),.clk(gclk));
	jdff dff_A_yOFZhdsY9_1(.dout(w_dff_A_2vzhdSBC8_1),.din(w_dff_A_yOFZhdsY9_1),.clk(gclk));
	jdff dff_A_EOOm8Zae7_1(.dout(w_dff_A_yOFZhdsY9_1),.din(w_dff_A_EOOm8Zae7_1),.clk(gclk));
	jdff dff_A_W6SOQCUV2_1(.dout(w_dff_A_EOOm8Zae7_1),.din(w_dff_A_W6SOQCUV2_1),.clk(gclk));
	jdff dff_A_8zyiSCVZ6_1(.dout(w_dff_A_W6SOQCUV2_1),.din(w_dff_A_8zyiSCVZ6_1),.clk(gclk));
	jdff dff_A_73FL0xGj1_1(.dout(w_dff_A_8zyiSCVZ6_1),.din(w_dff_A_73FL0xGj1_1),.clk(gclk));
	jdff dff_A_i51OnKUc9_1(.dout(w_dff_A_73FL0xGj1_1),.din(w_dff_A_i51OnKUc9_1),.clk(gclk));
	jdff dff_A_roWUZvzK1_1(.dout(w_dff_A_i51OnKUc9_1),.din(w_dff_A_roWUZvzK1_1),.clk(gclk));
	jdff dff_A_nEMLz3Xv9_1(.dout(w_dff_A_roWUZvzK1_1),.din(w_dff_A_nEMLz3Xv9_1),.clk(gclk));
	jdff dff_A_3QYF7sbO8_1(.dout(w_dff_A_nEMLz3Xv9_1),.din(w_dff_A_3QYF7sbO8_1),.clk(gclk));
	jdff dff_A_fE3PXaSr1_1(.dout(w_dff_A_3QYF7sbO8_1),.din(w_dff_A_fE3PXaSr1_1),.clk(gclk));
	jdff dff_A_lVagmxix5_2(.dout(w_n999_0[2]),.din(w_dff_A_lVagmxix5_2),.clk(gclk));
	jdff dff_A_mseKgEfw7_2(.dout(w_dff_A_lVagmxix5_2),.din(w_dff_A_mseKgEfw7_2),.clk(gclk));
	jdff dff_A_hyrXHCH65_2(.dout(w_dff_A_mseKgEfw7_2),.din(w_dff_A_hyrXHCH65_2),.clk(gclk));
	jdff dff_A_4RrNPMzp2_2(.dout(w_dff_A_hyrXHCH65_2),.din(w_dff_A_4RrNPMzp2_2),.clk(gclk));
	jdff dff_A_Y3eirACm9_2(.dout(w_dff_A_4RrNPMzp2_2),.din(w_dff_A_Y3eirACm9_2),.clk(gclk));
	jdff dff_A_rfJtINS35_2(.dout(w_dff_A_Y3eirACm9_2),.din(w_dff_A_rfJtINS35_2),.clk(gclk));
	jdff dff_A_aNJli9L43_2(.dout(w_dff_A_rfJtINS35_2),.din(w_dff_A_aNJli9L43_2),.clk(gclk));
	jdff dff_A_15yWLHBU3_2(.dout(w_dff_A_aNJli9L43_2),.din(w_dff_A_15yWLHBU3_2),.clk(gclk));
	jdff dff_A_CzxrGben0_2(.dout(w_dff_A_15yWLHBU3_2),.din(w_dff_A_CzxrGben0_2),.clk(gclk));
	jdff dff_A_4Xqc6g2q8_2(.dout(w_dff_A_CzxrGben0_2),.din(w_dff_A_4Xqc6g2q8_2),.clk(gclk));
	jdff dff_A_RoRRi9D51_1(.dout(w_G1694_0[1]),.din(w_dff_A_RoRRi9D51_1),.clk(gclk));
	jdff dff_A_YqYBMRA82_2(.dout(w_G1691_0[2]),.din(w_dff_A_YqYBMRA82_2),.clk(gclk));
	jdff dff_B_hAsW1QNe5_2(.din(n1624),.dout(w_dff_B_hAsW1QNe5_2),.clk(gclk));
	jdff dff_B_e8lsLn8v4_2(.din(w_dff_B_hAsW1QNe5_2),.dout(w_dff_B_e8lsLn8v4_2),.clk(gclk));
	jdff dff_B_GhCQXu828_2(.din(w_dff_B_e8lsLn8v4_2),.dout(w_dff_B_GhCQXu828_2),.clk(gclk));
	jdff dff_B_DdSWIOmF9_2(.din(w_dff_B_GhCQXu828_2),.dout(w_dff_B_DdSWIOmF9_2),.clk(gclk));
	jdff dff_B_LE69BYv77_2(.din(w_dff_B_DdSWIOmF9_2),.dout(w_dff_B_LE69BYv77_2),.clk(gclk));
	jdff dff_B_ex6DH80C1_2(.din(w_dff_B_LE69BYv77_2),.dout(w_dff_B_ex6DH80C1_2),.clk(gclk));
	jdff dff_B_yFtCufYV9_2(.din(w_dff_B_ex6DH80C1_2),.dout(w_dff_B_yFtCufYV9_2),.clk(gclk));
	jdff dff_B_IOQQV4z05_2(.din(w_dff_B_yFtCufYV9_2),.dout(w_dff_B_IOQQV4z05_2),.clk(gclk));
	jdff dff_B_HYMfqDBi5_2(.din(w_dff_B_IOQQV4z05_2),.dout(w_dff_B_HYMfqDBi5_2),.clk(gclk));
	jdff dff_B_MfX2NhZT2_2(.din(w_dff_B_HYMfqDBi5_2),.dout(w_dff_B_MfX2NhZT2_2),.clk(gclk));
	jdff dff_B_E7iF19gs1_2(.din(w_dff_B_MfX2NhZT2_2),.dout(w_dff_B_E7iF19gs1_2),.clk(gclk));
	jdff dff_B_Vdc2STjF8_2(.din(w_dff_B_E7iF19gs1_2),.dout(w_dff_B_Vdc2STjF8_2),.clk(gclk));
	jdff dff_B_XJnI6Mjh4_2(.din(w_dff_B_Vdc2STjF8_2),.dout(w_dff_B_XJnI6Mjh4_2),.clk(gclk));
	jdff dff_B_TIr9kou64_2(.din(w_dff_B_XJnI6Mjh4_2),.dout(w_dff_B_TIr9kou64_2),.clk(gclk));
	jdff dff_B_O1MltaaW7_2(.din(w_dff_B_TIr9kou64_2),.dout(w_dff_B_O1MltaaW7_2),.clk(gclk));
	jdff dff_B_2TonRPCs2_2(.din(w_dff_B_O1MltaaW7_2),.dout(w_dff_B_2TonRPCs2_2),.clk(gclk));
	jdff dff_B_Zp36ZbYQ3_2(.din(w_dff_B_2TonRPCs2_2),.dout(w_dff_B_Zp36ZbYQ3_2),.clk(gclk));
	jdff dff_A_pSl7gS7l5_2(.dout(w_G137_3[2]),.din(w_dff_A_pSl7gS7l5_2),.clk(gclk));
	jdff dff_A_7tP8I1sh3_2(.dout(w_dff_A_pSl7gS7l5_2),.din(w_dff_A_7tP8I1sh3_2),.clk(gclk));
	jdff dff_A_aRuwM3Bt5_2(.dout(w_dff_A_7tP8I1sh3_2),.din(w_dff_A_aRuwM3Bt5_2),.clk(gclk));
	jdff dff_A_umpHbgv29_2(.dout(w_dff_A_aRuwM3Bt5_2),.din(w_dff_A_umpHbgv29_2),.clk(gclk));
	jdff dff_A_SCuXrD4p4_2(.dout(w_dff_A_umpHbgv29_2),.din(w_dff_A_SCuXrD4p4_2),.clk(gclk));
	jdff dff_A_al0XeZAo5_2(.dout(w_dff_A_SCuXrD4p4_2),.din(w_dff_A_al0XeZAo5_2),.clk(gclk));
	jdff dff_A_ULJw2YN13_2(.dout(w_dff_A_al0XeZAo5_2),.din(w_dff_A_ULJw2YN13_2),.clk(gclk));
	jdff dff_A_vJgwuPfK8_2(.dout(w_dff_A_ULJw2YN13_2),.din(w_dff_A_vJgwuPfK8_2),.clk(gclk));
	jdff dff_A_nOoVUVcn4_2(.dout(w_dff_A_vJgwuPfK8_2),.din(w_dff_A_nOoVUVcn4_2),.clk(gclk));
	jdff dff_A_oLSzWvxp9_2(.dout(w_dff_A_nOoVUVcn4_2),.din(w_dff_A_oLSzWvxp9_2),.clk(gclk));
	jdff dff_A_9Sn4SKqe4_2(.dout(w_dff_A_oLSzWvxp9_2),.din(w_dff_A_9Sn4SKqe4_2),.clk(gclk));
	jdff dff_A_IrsfRMPU8_2(.dout(w_dff_A_9Sn4SKqe4_2),.din(w_dff_A_IrsfRMPU8_2),.clk(gclk));
	jdff dff_A_uOeiWLTT8_2(.dout(w_dff_A_IrsfRMPU8_2),.din(w_dff_A_uOeiWLTT8_2),.clk(gclk));
	jdff dff_A_F3DBGDKX0_2(.dout(w_dff_A_uOeiWLTT8_2),.din(w_dff_A_F3DBGDKX0_2),.clk(gclk));
	jdff dff_A_OuvWcien5_0(.dout(w_G137_0[0]),.din(w_dff_A_OuvWcien5_0),.clk(gclk));
	jdff dff_A_AzByg08a7_0(.dout(w_dff_A_OuvWcien5_0),.din(w_dff_A_AzByg08a7_0),.clk(gclk));
	jdff dff_A_nu0SSnYp0_0(.dout(w_dff_A_AzByg08a7_0),.din(w_dff_A_nu0SSnYp0_0),.clk(gclk));
	jdff dff_A_hnC9rVHO7_0(.dout(w_dff_A_nu0SSnYp0_0),.din(w_dff_A_hnC9rVHO7_0),.clk(gclk));
	jdff dff_A_4jFUwV7r7_0(.dout(w_dff_A_hnC9rVHO7_0),.din(w_dff_A_4jFUwV7r7_0),.clk(gclk));
	jdff dff_A_TLgGqsiv1_0(.dout(w_dff_A_4jFUwV7r7_0),.din(w_dff_A_TLgGqsiv1_0),.clk(gclk));
	jdff dff_A_798Txwvh4_0(.dout(w_dff_A_TLgGqsiv1_0),.din(w_dff_A_798Txwvh4_0),.clk(gclk));
	jdff dff_A_nc50f9tC2_0(.dout(w_dff_A_798Txwvh4_0),.din(w_dff_A_nc50f9tC2_0),.clk(gclk));
	jdff dff_A_mHr5OAWm1_0(.dout(w_dff_A_nc50f9tC2_0),.din(w_dff_A_mHr5OAWm1_0),.clk(gclk));
	jdff dff_A_EP1eZVSK3_0(.dout(w_dff_A_mHr5OAWm1_0),.din(w_dff_A_EP1eZVSK3_0),.clk(gclk));
	jdff dff_A_jrhmiOFV1_0(.dout(w_dff_A_EP1eZVSK3_0),.din(w_dff_A_jrhmiOFV1_0),.clk(gclk));
	jdff dff_A_fhfniE1w6_0(.dout(w_dff_A_jrhmiOFV1_0),.din(w_dff_A_fhfniE1w6_0),.clk(gclk));
	jdff dff_A_a8ZdlOSK8_0(.dout(w_dff_A_fhfniE1w6_0),.din(w_dff_A_a8ZdlOSK8_0),.clk(gclk));
	jdff dff_A_tQ26enkn1_1(.dout(w_G137_0[1]),.din(w_dff_A_tQ26enkn1_1),.clk(gclk));
	jdff dff_A_9mTtV3JI1_1(.dout(w_dff_A_tQ26enkn1_1),.din(w_dff_A_9mTtV3JI1_1),.clk(gclk));
	jdff dff_A_hSn8K9yg3_1(.dout(w_dff_A_9mTtV3JI1_1),.din(w_dff_A_hSn8K9yg3_1),.clk(gclk));
	jdff dff_A_vf2EN9pX1_1(.dout(w_dff_A_hSn8K9yg3_1),.din(w_dff_A_vf2EN9pX1_1),.clk(gclk));
	jdff dff_A_S5OQd7Ct9_1(.dout(w_dff_A_vf2EN9pX1_1),.din(w_dff_A_S5OQd7Ct9_1),.clk(gclk));
	jdff dff_A_USVXLc106_1(.dout(w_dff_A_S5OQd7Ct9_1),.din(w_dff_A_USVXLc106_1),.clk(gclk));
	jdff dff_A_ipof18BS6_1(.dout(w_dff_A_USVXLc106_1),.din(w_dff_A_ipof18BS6_1),.clk(gclk));
	jdff dff_A_f3QZiukM0_1(.dout(w_dff_A_ipof18BS6_1),.din(w_dff_A_f3QZiukM0_1),.clk(gclk));
	jdff dff_A_WjS2D61k4_1(.dout(w_dff_A_f3QZiukM0_1),.din(w_dff_A_WjS2D61k4_1),.clk(gclk));
endmodule

